// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N619,N608,N605,N596,N614,N617,N616,N613,N618,N621;

or OR4 (N22, N5, N20, N14, N10);
or OR2 (N23, N21, N22);
not NOT1 (N24, N14);
xor XOR2 (N25, N15, N4);
nor NOR3 (N26, N13, N17, N7);
nand NAND2 (N27, N18, N7);
nor NOR4 (N28, N12, N19, N16, N7);
or OR4 (N29, N20, N9, N9, N16);
xor XOR2 (N30, N13, N13);
not NOT1 (N31, N30);
xor XOR2 (N32, N13, N17);
buf BUF1 (N33, N6);
and AND2 (N34, N33, N4);
nor NOR2 (N35, N32, N20);
nand NAND3 (N36, N31, N34, N4);
xor XOR2 (N37, N26, N32);
and AND4 (N38, N2, N19, N17, N30);
and AND3 (N39, N37, N31, N4);
not NOT1 (N40, N27);
nand NAND3 (N41, N29, N4, N15);
buf BUF1 (N42, N35);
buf BUF1 (N43, N38);
buf BUF1 (N44, N24);
nand NAND3 (N45, N42, N38, N22);
xor XOR2 (N46, N28, N27);
buf BUF1 (N47, N43);
xor XOR2 (N48, N47, N7);
nand NAND4 (N49, N23, N41, N26, N1);
or OR2 (N50, N32, N1);
xor XOR2 (N51, N48, N49);
and AND4 (N52, N31, N7, N4, N37);
or OR3 (N53, N25, N32, N20);
and AND3 (N54, N52, N10, N41);
or OR3 (N55, N44, N10, N23);
not NOT1 (N56, N55);
buf BUF1 (N57, N51);
buf BUF1 (N58, N45);
and AND2 (N59, N57, N4);
nand NAND3 (N60, N39, N25, N36);
buf BUF1 (N61, N26);
buf BUF1 (N62, N54);
not NOT1 (N63, N61);
buf BUF1 (N64, N40);
nand NAND3 (N65, N60, N64, N56);
or OR2 (N66, N14, N40);
xor XOR2 (N67, N1, N24);
xor XOR2 (N68, N46, N52);
xor XOR2 (N69, N65, N51);
buf BUF1 (N70, N62);
buf BUF1 (N71, N70);
and AND2 (N72, N71, N37);
not NOT1 (N73, N53);
xor XOR2 (N74, N63, N49);
not NOT1 (N75, N58);
buf BUF1 (N76, N50);
buf BUF1 (N77, N75);
not NOT1 (N78, N59);
buf BUF1 (N79, N77);
buf BUF1 (N80, N72);
and AND3 (N81, N69, N31, N55);
buf BUF1 (N82, N73);
nor NOR3 (N83, N68, N67, N20);
or OR2 (N84, N16, N46);
not NOT1 (N85, N82);
nand NAND2 (N86, N66, N46);
buf BUF1 (N87, N81);
and AND4 (N88, N83, N37, N84, N38);
or OR3 (N89, N87, N17, N43);
not NOT1 (N90, N61);
and AND3 (N91, N89, N77, N2);
nor NOR2 (N92, N80, N90);
or OR4 (N93, N8, N34, N89, N27);
and AND3 (N94, N91, N10, N90);
xor XOR2 (N95, N74, N35);
or OR4 (N96, N86, N63, N45, N40);
xor XOR2 (N97, N96, N30);
nor NOR4 (N98, N88, N9, N8, N25);
and AND3 (N99, N95, N90, N65);
xor XOR2 (N100, N93, N54);
xor XOR2 (N101, N76, N80);
nor NOR3 (N102, N100, N58, N97);
and AND4 (N103, N6, N11, N10, N92);
and AND3 (N104, N91, N17, N30);
and AND3 (N105, N103, N54, N88);
nand NAND2 (N106, N104, N72);
xor XOR2 (N107, N102, N34);
xor XOR2 (N108, N85, N54);
buf BUF1 (N109, N78);
nand NAND2 (N110, N98, N46);
not NOT1 (N111, N99);
not NOT1 (N112, N106);
not NOT1 (N113, N111);
or OR3 (N114, N110, N4, N19);
and AND3 (N115, N101, N76, N113);
buf BUF1 (N116, N75);
buf BUF1 (N117, N108);
or OR4 (N118, N107, N91, N40, N60);
nor NOR2 (N119, N109, N33);
xor XOR2 (N120, N94, N10);
xor XOR2 (N121, N120, N98);
nor NOR4 (N122, N118, N35, N88, N115);
nand NAND4 (N123, N51, N26, N14, N83);
and AND3 (N124, N116, N87, N16);
or OR3 (N125, N121, N9, N83);
buf BUF1 (N126, N114);
nor NOR3 (N127, N119, N64, N43);
buf BUF1 (N128, N112);
xor XOR2 (N129, N127, N75);
nor NOR3 (N130, N129, N1, N40);
buf BUF1 (N131, N123);
or OR3 (N132, N125, N124, N7);
nand NAND3 (N133, N22, N126, N125);
xor XOR2 (N134, N100, N131);
not NOT1 (N135, N60);
not NOT1 (N136, N132);
nand NAND2 (N137, N134, N96);
xor XOR2 (N138, N137, N66);
not NOT1 (N139, N133);
buf BUF1 (N140, N138);
nand NAND3 (N141, N105, N124, N106);
buf BUF1 (N142, N79);
and AND4 (N143, N141, N58, N44, N132);
and AND3 (N144, N128, N58, N59);
nor NOR2 (N145, N135, N83);
or OR2 (N146, N145, N104);
xor XOR2 (N147, N143, N131);
or OR2 (N148, N142, N129);
nand NAND4 (N149, N148, N145, N29, N134);
nor NOR4 (N150, N144, N123, N73, N26);
not NOT1 (N151, N122);
buf BUF1 (N152, N130);
xor XOR2 (N153, N136, N49);
not NOT1 (N154, N152);
buf BUF1 (N155, N154);
nand NAND4 (N156, N117, N127, N53, N29);
nor NOR3 (N157, N139, N24, N89);
and AND3 (N158, N157, N113, N16);
nor NOR4 (N159, N147, N41, N125, N10);
buf BUF1 (N160, N155);
xor XOR2 (N161, N156, N46);
not NOT1 (N162, N140);
nand NAND2 (N163, N151, N41);
and AND4 (N164, N159, N58, N27, N68);
not NOT1 (N165, N149);
buf BUF1 (N166, N163);
not NOT1 (N167, N146);
nand NAND3 (N168, N164, N122, N45);
not NOT1 (N169, N160);
buf BUF1 (N170, N162);
xor XOR2 (N171, N170, N142);
nand NAND2 (N172, N165, N33);
not NOT1 (N173, N171);
nor NOR3 (N174, N169, N119, N52);
nor NOR3 (N175, N168, N7, N40);
xor XOR2 (N176, N153, N118);
not NOT1 (N177, N158);
nor NOR3 (N178, N167, N59, N66);
and AND2 (N179, N166, N45);
xor XOR2 (N180, N174, N4);
nand NAND2 (N181, N178, N22);
nand NAND4 (N182, N176, N124, N172, N77);
buf BUF1 (N183, N162);
and AND3 (N184, N173, N65, N38);
nor NOR3 (N185, N150, N40, N151);
nand NAND2 (N186, N181, N28);
and AND3 (N187, N177, N153, N155);
nor NOR3 (N188, N180, N187, N30);
and AND4 (N189, N153, N173, N70, N107);
nand NAND2 (N190, N179, N146);
and AND4 (N191, N182, N118, N188, N88);
nand NAND4 (N192, N154, N19, N98, N131);
or OR3 (N193, N191, N103, N42);
nor NOR2 (N194, N175, N67);
nand NAND3 (N195, N192, N39, N47);
not NOT1 (N196, N184);
buf BUF1 (N197, N185);
buf BUF1 (N198, N193);
nor NOR2 (N199, N197, N132);
not NOT1 (N200, N189);
nand NAND2 (N201, N190, N184);
not NOT1 (N202, N196);
or OR4 (N203, N195, N151, N153, N74);
and AND3 (N204, N161, N169, N118);
nand NAND3 (N205, N204, N107, N95);
not NOT1 (N206, N194);
or OR3 (N207, N200, N72, N133);
not NOT1 (N208, N205);
xor XOR2 (N209, N199, N24);
nor NOR3 (N210, N198, N164, N98);
nor NOR4 (N211, N210, N42, N7, N55);
and AND4 (N212, N183, N211, N175, N172);
xor XOR2 (N213, N156, N82);
nor NOR4 (N214, N212, N56, N179, N106);
nor NOR3 (N215, N208, N152, N152);
nor NOR2 (N216, N202, N92);
not NOT1 (N217, N214);
buf BUF1 (N218, N216);
and AND3 (N219, N217, N79, N134);
xor XOR2 (N220, N186, N139);
not NOT1 (N221, N207);
buf BUF1 (N222, N215);
or OR2 (N223, N222, N144);
not NOT1 (N224, N213);
nand NAND4 (N225, N206, N158, N132, N12);
xor XOR2 (N226, N218, N47);
nand NAND2 (N227, N219, N190);
or OR4 (N228, N203, N170, N56, N34);
or OR3 (N229, N225, N173, N103);
and AND4 (N230, N224, N132, N163, N116);
not NOT1 (N231, N226);
nand NAND2 (N232, N231, N88);
buf BUF1 (N233, N201);
or OR3 (N234, N228, N111, N149);
or OR3 (N235, N232, N115, N115);
or OR2 (N236, N234, N12);
not NOT1 (N237, N220);
not NOT1 (N238, N229);
nand NAND3 (N239, N235, N150, N158);
nor NOR2 (N240, N221, N43);
not NOT1 (N241, N239);
xor XOR2 (N242, N238, N169);
nand NAND4 (N243, N209, N10, N129, N137);
buf BUF1 (N244, N237);
xor XOR2 (N245, N240, N201);
nand NAND4 (N246, N243, N231, N190, N26);
and AND2 (N247, N227, N45);
not NOT1 (N248, N246);
xor XOR2 (N249, N233, N130);
nor NOR4 (N250, N247, N22, N31, N112);
or OR4 (N251, N223, N119, N72, N36);
xor XOR2 (N252, N244, N145);
xor XOR2 (N253, N245, N149);
nand NAND3 (N254, N250, N144, N2);
not NOT1 (N255, N241);
and AND3 (N256, N255, N98, N6);
xor XOR2 (N257, N252, N249);
or OR2 (N258, N201, N59);
buf BUF1 (N259, N251);
buf BUF1 (N260, N248);
buf BUF1 (N261, N260);
nor NOR2 (N262, N254, N136);
buf BUF1 (N263, N253);
nor NOR2 (N264, N236, N146);
buf BUF1 (N265, N257);
not NOT1 (N266, N264);
nand NAND4 (N267, N259, N205, N161, N183);
not NOT1 (N268, N267);
nand NAND4 (N269, N261, N259, N174, N101);
nor NOR4 (N270, N266, N225, N57, N246);
not NOT1 (N271, N263);
nand NAND4 (N272, N230, N210, N178, N31);
nor NOR2 (N273, N271, N198);
xor XOR2 (N274, N268, N250);
not NOT1 (N275, N258);
xor XOR2 (N276, N275, N149);
or OR2 (N277, N265, N24);
nand NAND2 (N278, N256, N252);
and AND2 (N279, N278, N144);
nand NAND4 (N280, N274, N148, N121, N180);
and AND2 (N281, N279, N203);
nand NAND2 (N282, N276, N49);
xor XOR2 (N283, N280, N271);
buf BUF1 (N284, N277);
xor XOR2 (N285, N284, N107);
or OR4 (N286, N283, N141, N100, N121);
nor NOR2 (N287, N262, N225);
buf BUF1 (N288, N286);
nand NAND3 (N289, N285, N281, N71);
nand NAND3 (N290, N94, N96, N241);
and AND3 (N291, N289, N77, N134);
xor XOR2 (N292, N270, N224);
xor XOR2 (N293, N288, N113);
or OR4 (N294, N242, N165, N254, N248);
nand NAND2 (N295, N272, N42);
xor XOR2 (N296, N287, N119);
and AND3 (N297, N282, N121, N1);
xor XOR2 (N298, N269, N33);
nor NOR4 (N299, N273, N289, N41, N43);
not NOT1 (N300, N298);
nand NAND2 (N301, N292, N295);
nor NOR3 (N302, N152, N47, N240);
xor XOR2 (N303, N297, N225);
and AND4 (N304, N302, N157, N295, N40);
and AND2 (N305, N294, N66);
nand NAND3 (N306, N299, N298, N206);
or OR2 (N307, N296, N88);
and AND2 (N308, N301, N264);
buf BUF1 (N309, N304);
and AND2 (N310, N306, N14);
nor NOR2 (N311, N300, N288);
xor XOR2 (N312, N307, N307);
nor NOR2 (N313, N309, N199);
xor XOR2 (N314, N313, N274);
xor XOR2 (N315, N293, N151);
xor XOR2 (N316, N315, N130);
or OR2 (N317, N312, N37);
nor NOR2 (N318, N291, N183);
or OR4 (N319, N290, N314, N187, N246);
nor NOR4 (N320, N125, N141, N106, N123);
buf BUF1 (N321, N308);
buf BUF1 (N322, N318);
nand NAND3 (N323, N305, N141, N288);
or OR2 (N324, N319, N54);
nand NAND3 (N325, N321, N305, N10);
or OR3 (N326, N317, N240, N313);
not NOT1 (N327, N325);
or OR2 (N328, N310, N92);
nand NAND4 (N329, N323, N44, N171, N153);
xor XOR2 (N330, N311, N93);
xor XOR2 (N331, N328, N281);
or OR2 (N332, N330, N266);
nor NOR2 (N333, N316, N195);
xor XOR2 (N334, N320, N184);
or OR2 (N335, N303, N253);
nor NOR4 (N336, N329, N288, N20, N49);
xor XOR2 (N337, N327, N316);
nand NAND3 (N338, N334, N251, N204);
not NOT1 (N339, N331);
nand NAND2 (N340, N338, N242);
xor XOR2 (N341, N332, N56);
buf BUF1 (N342, N326);
nand NAND3 (N343, N337, N174, N84);
buf BUF1 (N344, N340);
not NOT1 (N345, N336);
xor XOR2 (N346, N344, N321);
buf BUF1 (N347, N346);
or OR4 (N348, N342, N25, N309, N29);
not NOT1 (N349, N341);
nand NAND3 (N350, N322, N2, N182);
nor NOR3 (N351, N335, N280, N58);
nor NOR4 (N352, N351, N26, N157, N59);
xor XOR2 (N353, N339, N62);
not NOT1 (N354, N345);
nor NOR2 (N355, N349, N168);
nand NAND2 (N356, N354, N253);
or OR3 (N357, N356, N187, N189);
and AND4 (N358, N353, N286, N293, N285);
and AND3 (N359, N355, N150, N303);
buf BUF1 (N360, N358);
nor NOR3 (N361, N343, N275, N247);
or OR4 (N362, N333, N168, N349, N206);
or OR2 (N363, N348, N336);
buf BUF1 (N364, N352);
not NOT1 (N365, N350);
or OR4 (N366, N357, N169, N299, N308);
and AND3 (N367, N361, N200, N140);
and AND4 (N368, N324, N40, N195, N359);
not NOT1 (N369, N147);
not NOT1 (N370, N367);
or OR4 (N371, N362, N364, N180, N175);
nand NAND2 (N372, N320, N185);
xor XOR2 (N373, N372, N371);
nand NAND2 (N374, N10, N347);
not NOT1 (N375, N195);
and AND4 (N376, N370, N31, N294, N114);
nand NAND2 (N377, N373, N237);
nand NAND3 (N378, N369, N245, N329);
or OR2 (N379, N368, N365);
xor XOR2 (N380, N63, N186);
nor NOR4 (N381, N376, N33, N155, N187);
xor XOR2 (N382, N375, N175);
nor NOR3 (N383, N379, N18, N302);
xor XOR2 (N384, N377, N152);
xor XOR2 (N385, N366, N175);
nand NAND3 (N386, N360, N220, N376);
buf BUF1 (N387, N382);
not NOT1 (N388, N378);
buf BUF1 (N389, N374);
and AND2 (N390, N386, N48);
nand NAND3 (N391, N383, N195, N200);
nor NOR2 (N392, N387, N349);
or OR2 (N393, N385, N168);
nand NAND3 (N394, N393, N365, N67);
nand NAND4 (N395, N390, N170, N336, N99);
and AND2 (N396, N394, N97);
nand NAND3 (N397, N384, N113, N228);
xor XOR2 (N398, N392, N44);
not NOT1 (N399, N389);
not NOT1 (N400, N380);
nor NOR3 (N401, N400, N5, N165);
not NOT1 (N402, N397);
or OR3 (N403, N388, N251, N373);
or OR3 (N404, N363, N211, N188);
nor NOR2 (N405, N391, N42);
nand NAND2 (N406, N398, N148);
not NOT1 (N407, N396);
and AND2 (N408, N399, N315);
and AND3 (N409, N381, N198, N166);
nor NOR4 (N410, N402, N99, N331, N260);
nand NAND2 (N411, N405, N146);
and AND3 (N412, N404, N16, N104);
xor XOR2 (N413, N407, N64);
xor XOR2 (N414, N406, N318);
or OR3 (N415, N414, N301, N143);
buf BUF1 (N416, N408);
xor XOR2 (N417, N412, N399);
or OR2 (N418, N403, N55);
buf BUF1 (N419, N413);
buf BUF1 (N420, N395);
xor XOR2 (N421, N415, N214);
nand NAND4 (N422, N410, N266, N380, N308);
not NOT1 (N423, N401);
nand NAND2 (N424, N418, N201);
or OR4 (N425, N424, N55, N324, N412);
or OR3 (N426, N411, N102, N413);
nor NOR2 (N427, N416, N331);
nor NOR3 (N428, N419, N246, N346);
or OR4 (N429, N409, N250, N332, N118);
not NOT1 (N430, N417);
and AND4 (N431, N429, N253, N212, N263);
or OR4 (N432, N422, N304, N19, N48);
or OR4 (N433, N426, N185, N242, N345);
xor XOR2 (N434, N425, N40);
xor XOR2 (N435, N427, N331);
buf BUF1 (N436, N432);
and AND3 (N437, N430, N361, N248);
buf BUF1 (N438, N428);
or OR2 (N439, N437, N83);
not NOT1 (N440, N423);
xor XOR2 (N441, N420, N70);
not NOT1 (N442, N440);
not NOT1 (N443, N442);
nor NOR3 (N444, N439, N212, N246);
not NOT1 (N445, N444);
xor XOR2 (N446, N421, N232);
xor XOR2 (N447, N446, N173);
not NOT1 (N448, N438);
or OR3 (N449, N441, N222, N101);
not NOT1 (N450, N447);
xor XOR2 (N451, N434, N373);
not NOT1 (N452, N443);
nor NOR3 (N453, N433, N110, N64);
and AND4 (N454, N445, N115, N179, N81);
not NOT1 (N455, N448);
or OR2 (N456, N451, N454);
xor XOR2 (N457, N257, N246);
buf BUF1 (N458, N456);
not NOT1 (N459, N453);
nand NAND2 (N460, N435, N401);
buf BUF1 (N461, N460);
not NOT1 (N462, N449);
nor NOR2 (N463, N452, N275);
nand NAND3 (N464, N436, N325, N345);
nor NOR2 (N465, N455, N336);
nor NOR4 (N466, N450, N405, N206, N6);
buf BUF1 (N467, N461);
or OR3 (N468, N466, N382, N14);
or OR2 (N469, N465, N359);
buf BUF1 (N470, N467);
xor XOR2 (N471, N468, N266);
not NOT1 (N472, N471);
xor XOR2 (N473, N458, N240);
not NOT1 (N474, N463);
xor XOR2 (N475, N473, N236);
and AND2 (N476, N462, N307);
xor XOR2 (N477, N476, N442);
buf BUF1 (N478, N431);
nor NOR2 (N479, N472, N337);
nor NOR4 (N480, N459, N20, N469, N406);
xor XOR2 (N481, N64, N3);
xor XOR2 (N482, N479, N61);
buf BUF1 (N483, N474);
xor XOR2 (N484, N464, N66);
nor NOR2 (N485, N484, N326);
not NOT1 (N486, N481);
or OR4 (N487, N485, N414, N404, N355);
not NOT1 (N488, N483);
buf BUF1 (N489, N486);
not NOT1 (N490, N477);
not NOT1 (N491, N482);
or OR4 (N492, N487, N22, N273, N278);
buf BUF1 (N493, N492);
not NOT1 (N494, N470);
xor XOR2 (N495, N490, N374);
or OR4 (N496, N488, N18, N283, N32);
buf BUF1 (N497, N494);
nand NAND2 (N498, N478, N26);
buf BUF1 (N499, N498);
not NOT1 (N500, N493);
xor XOR2 (N501, N491, N124);
nor NOR2 (N502, N497, N175);
not NOT1 (N503, N502);
and AND4 (N504, N500, N309, N478, N280);
buf BUF1 (N505, N457);
buf BUF1 (N506, N496);
xor XOR2 (N507, N503, N263);
not NOT1 (N508, N499);
nand NAND3 (N509, N505, N132, N78);
nand NAND4 (N510, N501, N342, N458, N218);
nor NOR2 (N511, N510, N85);
xor XOR2 (N512, N508, N231);
nor NOR3 (N513, N495, N197, N150);
nor NOR4 (N514, N504, N290, N464, N202);
xor XOR2 (N515, N511, N383);
nor NOR2 (N516, N513, N487);
and AND2 (N517, N506, N136);
and AND4 (N518, N475, N106, N203, N337);
and AND4 (N519, N489, N77, N435, N79);
nor NOR3 (N520, N517, N98, N15);
xor XOR2 (N521, N507, N495);
nand NAND2 (N522, N514, N500);
not NOT1 (N523, N516);
nand NAND3 (N524, N522, N121, N445);
or OR4 (N525, N524, N323, N239, N328);
and AND3 (N526, N525, N337, N136);
nor NOR2 (N527, N521, N283);
nor NOR2 (N528, N519, N3);
xor XOR2 (N529, N527, N259);
not NOT1 (N530, N528);
nor NOR4 (N531, N480, N123, N314, N343);
or OR2 (N532, N530, N198);
xor XOR2 (N533, N532, N117);
nor NOR4 (N534, N518, N147, N527, N245);
nand NAND3 (N535, N534, N478, N18);
or OR2 (N536, N535, N374);
not NOT1 (N537, N509);
or OR3 (N538, N533, N485, N436);
not NOT1 (N539, N512);
or OR4 (N540, N537, N317, N145, N120);
not NOT1 (N541, N539);
buf BUF1 (N542, N538);
and AND3 (N543, N526, N235, N539);
or OR3 (N544, N531, N509, N479);
nand NAND2 (N545, N544, N400);
buf BUF1 (N546, N543);
and AND2 (N547, N545, N97);
xor XOR2 (N548, N520, N23);
xor XOR2 (N549, N523, N59);
nor NOR2 (N550, N540, N190);
buf BUF1 (N551, N542);
xor XOR2 (N552, N536, N48);
nand NAND2 (N553, N529, N278);
not NOT1 (N554, N549);
not NOT1 (N555, N552);
and AND3 (N556, N541, N518, N126);
nor NOR4 (N557, N546, N5, N260, N225);
and AND2 (N558, N553, N515);
buf BUF1 (N559, N76);
and AND2 (N560, N555, N398);
and AND3 (N561, N558, N471, N29);
nand NAND2 (N562, N547, N154);
xor XOR2 (N563, N548, N484);
not NOT1 (N564, N550);
buf BUF1 (N565, N561);
and AND4 (N566, N556, N426, N195, N81);
xor XOR2 (N567, N563, N256);
buf BUF1 (N568, N562);
nor NOR3 (N569, N551, N90, N537);
or OR2 (N570, N567, N407);
and AND2 (N571, N566, N222);
and AND3 (N572, N560, N198, N209);
or OR4 (N573, N572, N64, N424, N295);
buf BUF1 (N574, N571);
and AND3 (N575, N559, N496, N298);
not NOT1 (N576, N575);
or OR2 (N577, N564, N386);
nand NAND2 (N578, N577, N511);
nor NOR2 (N579, N557, N484);
nand NAND3 (N580, N569, N214, N270);
xor XOR2 (N581, N576, N148);
and AND4 (N582, N580, N247, N430, N33);
or OR4 (N583, N554, N375, N322, N122);
buf BUF1 (N584, N579);
nand NAND4 (N585, N583, N434, N175, N292);
buf BUF1 (N586, N568);
nand NAND2 (N587, N581, N408);
and AND2 (N588, N582, N48);
and AND3 (N589, N570, N535, N579);
or OR4 (N590, N585, N275, N532, N11);
or OR3 (N591, N589, N193, N37);
nor NOR2 (N592, N591, N253);
xor XOR2 (N593, N573, N159);
buf BUF1 (N594, N584);
nand NAND3 (N595, N565, N75, N582);
nor NOR3 (N596, N595, N555, N558);
not NOT1 (N597, N594);
xor XOR2 (N598, N593, N520);
nand NAND2 (N599, N578, N175);
and AND4 (N600, N587, N36, N23, N302);
and AND2 (N601, N598, N347);
or OR3 (N602, N592, N97, N24);
buf BUF1 (N603, N599);
nor NOR4 (N604, N600, N36, N359, N495);
and AND2 (N605, N590, N315);
nand NAND2 (N606, N601, N170);
nand NAND4 (N607, N606, N127, N52, N154);
not NOT1 (N608, N574);
or OR2 (N609, N597, N300);
nor NOR4 (N610, N586, N501, N42, N434);
buf BUF1 (N611, N607);
not NOT1 (N612, N609);
and AND3 (N613, N604, N529, N507);
not NOT1 (N614, N603);
not NOT1 (N615, N612);
nand NAND2 (N616, N602, N469);
or OR2 (N617, N588, N12);
xor XOR2 (N618, N615, N113);
nor NOR2 (N619, N611, N174);
or OR2 (N620, N610, N299);
or OR2 (N621, N620, N12);
endmodule