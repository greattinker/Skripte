// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N2009,N2010,N2007,N2003,N2006,N2001,N2013,N2012,N2011,N2014;

or OR2 (N15, N8, N12);
xor XOR2 (N16, N11, N5);
or OR3 (N17, N16, N4, N11);
not NOT1 (N18, N1);
nor NOR2 (N19, N17, N7);
not NOT1 (N20, N14);
nor NOR4 (N21, N9, N12, N2, N20);
not NOT1 (N22, N5);
nand NAND3 (N23, N13, N20, N8);
buf BUF1 (N24, N22);
not NOT1 (N25, N5);
nand NAND3 (N26, N1, N25, N14);
nand NAND4 (N27, N26, N6, N2, N3);
xor XOR2 (N28, N10, N15);
nand NAND3 (N29, N16, N13, N24);
or OR3 (N30, N13, N27, N7);
nand NAND4 (N31, N3, N5, N6, N19);
and AND4 (N32, N17, N5, N22, N21);
xor XOR2 (N33, N23, N16);
xor XOR2 (N34, N23, N9);
buf BUF1 (N35, N22);
nor NOR2 (N36, N6, N29);
or OR4 (N37, N13, N15, N10, N6);
not NOT1 (N38, N18);
and AND2 (N39, N33, N20);
and AND3 (N40, N37, N6, N15);
or OR2 (N41, N30, N15);
nand NAND2 (N42, N38, N37);
nor NOR4 (N43, N28, N3, N23, N38);
or OR3 (N44, N39, N41, N35);
nor NOR2 (N45, N16, N22);
xor XOR2 (N46, N18, N32);
or OR3 (N47, N14, N43, N13);
xor XOR2 (N48, N29, N40);
or OR4 (N49, N4, N44, N16, N11);
and AND2 (N50, N10, N23);
xor XOR2 (N51, N49, N1);
nor NOR3 (N52, N46, N16, N18);
and AND4 (N53, N47, N10, N8, N14);
and AND2 (N54, N52, N14);
buf BUF1 (N55, N54);
buf BUF1 (N56, N48);
nand NAND3 (N57, N56, N32, N38);
nand NAND2 (N58, N31, N32);
not NOT1 (N59, N53);
nand NAND3 (N60, N57, N7, N4);
buf BUF1 (N61, N60);
buf BUF1 (N62, N59);
nand NAND4 (N63, N42, N59, N19, N13);
not NOT1 (N64, N50);
nor NOR3 (N65, N58, N43, N34);
and AND2 (N66, N7, N26);
and AND3 (N67, N55, N34, N61);
not NOT1 (N68, N28);
or OR2 (N69, N45, N50);
nor NOR4 (N70, N51, N38, N23, N36);
or OR4 (N71, N43, N62, N62, N55);
nor NOR2 (N72, N19, N66);
or OR4 (N73, N13, N35, N38, N51);
or OR3 (N74, N72, N58, N24);
buf BUF1 (N75, N64);
or OR4 (N76, N67, N71, N6, N2);
buf BUF1 (N77, N41);
and AND2 (N78, N69, N49);
and AND2 (N79, N74, N21);
not NOT1 (N80, N68);
or OR4 (N81, N73, N9, N41, N35);
nand NAND2 (N82, N80, N42);
nand NAND4 (N83, N79, N81, N78, N47);
buf BUF1 (N84, N21);
not NOT1 (N85, N18);
nand NAND3 (N86, N85, N28, N59);
and AND2 (N87, N63, N77);
or OR3 (N88, N29, N37, N33);
or OR2 (N89, N84, N12);
or OR4 (N90, N89, N75, N45, N50);
or OR2 (N91, N23, N41);
nor NOR4 (N92, N91, N14, N22, N57);
or OR4 (N93, N90, N55, N46, N78);
and AND2 (N94, N76, N23);
xor XOR2 (N95, N94, N37);
and AND2 (N96, N93, N42);
nor NOR3 (N97, N95, N58, N14);
not NOT1 (N98, N82);
buf BUF1 (N99, N65);
nor NOR3 (N100, N87, N43, N58);
or OR4 (N101, N96, N98, N1, N5);
buf BUF1 (N102, N98);
xor XOR2 (N103, N99, N61);
not NOT1 (N104, N70);
not NOT1 (N105, N103);
buf BUF1 (N106, N102);
nor NOR3 (N107, N105, N10, N24);
or OR4 (N108, N83, N10, N98, N82);
buf BUF1 (N109, N101);
not NOT1 (N110, N86);
buf BUF1 (N111, N104);
not NOT1 (N112, N107);
nor NOR4 (N113, N97, N112, N9, N3);
xor XOR2 (N114, N15, N92);
nor NOR4 (N115, N88, N40, N10, N71);
or OR4 (N116, N3, N37, N44, N16);
nand NAND4 (N117, N108, N80, N8, N88);
buf BUF1 (N118, N117);
nand NAND2 (N119, N111, N40);
and AND3 (N120, N118, N39, N51);
not NOT1 (N121, N106);
nand NAND2 (N122, N115, N110);
or OR2 (N123, N6, N13);
buf BUF1 (N124, N109);
nor NOR4 (N125, N121, N67, N80, N120);
not NOT1 (N126, N18);
and AND3 (N127, N100, N55, N57);
and AND2 (N128, N114, N98);
nor NOR3 (N129, N113, N109, N122);
xor XOR2 (N130, N64, N10);
or OR4 (N131, N123, N86, N65, N25);
not NOT1 (N132, N125);
buf BUF1 (N133, N132);
nand NAND2 (N134, N119, N54);
and AND3 (N135, N124, N55, N66);
or OR4 (N136, N116, N108, N62, N102);
and AND4 (N137, N135, N2, N43, N77);
not NOT1 (N138, N134);
nor NOR4 (N139, N126, N107, N55, N112);
and AND3 (N140, N136, N124, N83);
or OR4 (N141, N133, N23, N137, N117);
and AND2 (N142, N116, N1);
xor XOR2 (N143, N130, N30);
not NOT1 (N144, N142);
not NOT1 (N145, N141);
or OR3 (N146, N139, N65, N85);
nor NOR3 (N147, N129, N98, N124);
xor XOR2 (N148, N127, N44);
not NOT1 (N149, N128);
not NOT1 (N150, N144);
or OR4 (N151, N148, N105, N93, N111);
or OR3 (N152, N150, N83, N137);
not NOT1 (N153, N138);
xor XOR2 (N154, N147, N74);
buf BUF1 (N155, N146);
xor XOR2 (N156, N131, N154);
buf BUF1 (N157, N94);
nor NOR3 (N158, N156, N24, N132);
nand NAND2 (N159, N143, N106);
and AND3 (N160, N140, N150, N53);
and AND4 (N161, N145, N121, N144, N142);
not NOT1 (N162, N157);
and AND2 (N163, N151, N30);
nand NAND2 (N164, N163, N82);
nor NOR3 (N165, N153, N40, N138);
xor XOR2 (N166, N155, N160);
and AND2 (N167, N129, N20);
nand NAND2 (N168, N161, N139);
buf BUF1 (N169, N158);
buf BUF1 (N170, N162);
buf BUF1 (N171, N166);
and AND2 (N172, N171, N149);
and AND4 (N173, N145, N109, N135, N105);
nand NAND2 (N174, N159, N105);
and AND3 (N175, N165, N99, N26);
buf BUF1 (N176, N170);
or OR4 (N177, N167, N119, N30, N100);
buf BUF1 (N178, N175);
nand NAND2 (N179, N174, N82);
nand NAND4 (N180, N168, N101, N151, N173);
or OR3 (N181, N40, N59, N39);
nand NAND2 (N182, N169, N81);
and AND3 (N183, N164, N168, N94);
or OR2 (N184, N178, N12);
not NOT1 (N185, N181);
and AND2 (N186, N182, N90);
buf BUF1 (N187, N177);
buf BUF1 (N188, N152);
buf BUF1 (N189, N180);
or OR3 (N190, N184, N124, N182);
or OR3 (N191, N185, N26, N167);
not NOT1 (N192, N186);
and AND4 (N193, N187, N44, N18, N76);
not NOT1 (N194, N191);
and AND3 (N195, N179, N80, N110);
nand NAND3 (N196, N176, N136, N126);
or OR4 (N197, N172, N36, N175, N35);
not NOT1 (N198, N195);
buf BUF1 (N199, N183);
not NOT1 (N200, N190);
and AND2 (N201, N194, N143);
not NOT1 (N202, N192);
buf BUF1 (N203, N196);
or OR2 (N204, N197, N76);
nand NAND4 (N205, N199, N64, N92, N93);
and AND4 (N206, N188, N60, N177, N190);
buf BUF1 (N207, N202);
buf BUF1 (N208, N203);
nor NOR2 (N209, N206, N131);
nor NOR4 (N210, N201, N13, N55, N46);
nand NAND2 (N211, N200, N94);
nand NAND4 (N212, N207, N5, N117, N56);
or OR4 (N213, N211, N181, N174, N63);
xor XOR2 (N214, N193, N129);
not NOT1 (N215, N198);
buf BUF1 (N216, N210);
not NOT1 (N217, N205);
nand NAND4 (N218, N189, N37, N57, N44);
not NOT1 (N219, N216);
not NOT1 (N220, N219);
buf BUF1 (N221, N212);
nor NOR2 (N222, N218, N168);
not NOT1 (N223, N221);
and AND2 (N224, N220, N73);
nor NOR2 (N225, N214, N51);
nand NAND2 (N226, N204, N178);
nor NOR4 (N227, N213, N208, N202, N210);
not NOT1 (N228, N174);
buf BUF1 (N229, N226);
and AND4 (N230, N229, N175, N48, N122);
nor NOR2 (N231, N224, N48);
or OR3 (N232, N228, N102, N169);
buf BUF1 (N233, N209);
xor XOR2 (N234, N223, N115);
nor NOR4 (N235, N217, N149, N213, N85);
or OR3 (N236, N233, N93, N62);
xor XOR2 (N237, N232, N140);
and AND2 (N238, N215, N29);
or OR2 (N239, N235, N218);
or OR3 (N240, N239, N131, N131);
nand NAND4 (N241, N238, N189, N87, N178);
nand NAND4 (N242, N240, N120, N33, N37);
buf BUF1 (N243, N236);
or OR2 (N244, N243, N173);
and AND2 (N245, N230, N184);
xor XOR2 (N246, N241, N233);
not NOT1 (N247, N227);
buf BUF1 (N248, N247);
xor XOR2 (N249, N242, N193);
xor XOR2 (N250, N234, N16);
xor XOR2 (N251, N245, N69);
nor NOR2 (N252, N244, N185);
nand NAND3 (N253, N222, N193, N196);
or OR4 (N254, N237, N175, N248, N36);
nor NOR4 (N255, N28, N72, N60, N138);
and AND2 (N256, N254, N252);
nor NOR4 (N257, N251, N256, N114, N140);
nor NOR4 (N258, N231, N220, N42, N207);
nand NAND4 (N259, N70, N122, N154, N145);
nor NOR3 (N260, N182, N236, N1);
buf BUF1 (N261, N249);
nand NAND2 (N262, N257, N98);
nor NOR4 (N263, N262, N48, N160, N77);
nand NAND3 (N264, N263, N103, N15);
nor NOR2 (N265, N253, N134);
xor XOR2 (N266, N259, N230);
xor XOR2 (N267, N260, N2);
xor XOR2 (N268, N265, N157);
or OR4 (N269, N246, N45, N144, N161);
nor NOR4 (N270, N267, N240, N239, N57);
buf BUF1 (N271, N258);
and AND2 (N272, N270, N192);
nand NAND4 (N273, N264, N32, N74, N38);
nor NOR3 (N274, N266, N181, N52);
buf BUF1 (N275, N274);
xor XOR2 (N276, N272, N44);
nand NAND3 (N277, N273, N247, N11);
buf BUF1 (N278, N250);
xor XOR2 (N279, N255, N22);
nand NAND3 (N280, N225, N86, N141);
xor XOR2 (N281, N275, N53);
not NOT1 (N282, N268);
xor XOR2 (N283, N281, N239);
nand NAND3 (N284, N282, N142, N61);
and AND4 (N285, N261, N179, N132, N75);
and AND2 (N286, N271, N264);
or OR3 (N287, N279, N94, N279);
buf BUF1 (N288, N269);
and AND3 (N289, N288, N125, N118);
nand NAND4 (N290, N284, N119, N178, N15);
nand NAND2 (N291, N287, N1);
buf BUF1 (N292, N276);
buf BUF1 (N293, N285);
nor NOR3 (N294, N290, N167, N144);
nor NOR2 (N295, N277, N240);
not NOT1 (N296, N280);
not NOT1 (N297, N283);
buf BUF1 (N298, N286);
nand NAND2 (N299, N292, N147);
and AND3 (N300, N295, N140, N69);
nor NOR4 (N301, N296, N74, N217, N224);
or OR2 (N302, N297, N255);
and AND3 (N303, N293, N179, N106);
buf BUF1 (N304, N289);
nor NOR2 (N305, N299, N208);
nand NAND2 (N306, N300, N33);
not NOT1 (N307, N291);
and AND3 (N308, N306, N68, N286);
or OR3 (N309, N303, N245, N108);
buf BUF1 (N310, N309);
nand NAND4 (N311, N302, N89, N17, N112);
buf BUF1 (N312, N310);
and AND3 (N313, N304, N71, N86);
nor NOR3 (N314, N278, N130, N228);
or OR3 (N315, N311, N59, N159);
or OR4 (N316, N308, N93, N157, N295);
and AND3 (N317, N298, N102, N82);
buf BUF1 (N318, N294);
and AND3 (N319, N314, N82, N50);
not NOT1 (N320, N312);
and AND3 (N321, N320, N144, N41);
nand NAND3 (N322, N301, N176, N37);
buf BUF1 (N323, N315);
or OR3 (N324, N323, N1, N88);
nand NAND3 (N325, N317, N91, N245);
and AND2 (N326, N318, N185);
and AND3 (N327, N319, N182, N145);
buf BUF1 (N328, N326);
and AND2 (N329, N328, N94);
and AND3 (N330, N307, N7, N65);
nor NOR2 (N331, N305, N3);
or OR4 (N332, N316, N38, N154, N181);
buf BUF1 (N333, N327);
buf BUF1 (N334, N330);
and AND4 (N335, N324, N140, N304, N84);
and AND4 (N336, N331, N122, N308, N183);
xor XOR2 (N337, N313, N11);
nor NOR2 (N338, N332, N170);
nor NOR2 (N339, N338, N159);
nand NAND4 (N340, N329, N178, N195, N300);
xor XOR2 (N341, N337, N330);
nand NAND4 (N342, N340, N113, N57, N36);
buf BUF1 (N343, N321);
not NOT1 (N344, N339);
xor XOR2 (N345, N344, N172);
nand NAND3 (N346, N341, N210, N202);
not NOT1 (N347, N335);
buf BUF1 (N348, N345);
buf BUF1 (N349, N334);
and AND3 (N350, N325, N162, N99);
nand NAND4 (N351, N333, N22, N28, N21);
not NOT1 (N352, N350);
not NOT1 (N353, N351);
not NOT1 (N354, N349);
and AND2 (N355, N342, N110);
nand NAND4 (N356, N352, N153, N254, N92);
nand NAND4 (N357, N353, N315, N203, N203);
buf BUF1 (N358, N343);
xor XOR2 (N359, N322, N32);
or OR2 (N360, N359, N326);
not NOT1 (N361, N355);
nor NOR2 (N362, N336, N28);
nand NAND4 (N363, N362, N308, N276, N17);
not NOT1 (N364, N357);
nand NAND3 (N365, N356, N15, N139);
buf BUF1 (N366, N364);
or OR4 (N367, N363, N22, N308, N127);
not NOT1 (N368, N358);
nor NOR4 (N369, N367, N320, N134, N331);
nand NAND2 (N370, N366, N73);
nand NAND4 (N371, N348, N55, N293, N129);
nor NOR4 (N372, N361, N15, N80, N275);
nor NOR4 (N373, N347, N42, N279, N147);
nor NOR4 (N374, N346, N43, N56, N69);
buf BUF1 (N375, N354);
buf BUF1 (N376, N374);
buf BUF1 (N377, N376);
nand NAND2 (N378, N369, N18);
not NOT1 (N379, N377);
buf BUF1 (N380, N378);
and AND4 (N381, N380, N231, N363, N181);
nor NOR2 (N382, N365, N54);
or OR2 (N383, N372, N116);
or OR3 (N384, N375, N277, N319);
xor XOR2 (N385, N383, N368);
not NOT1 (N386, N140);
or OR2 (N387, N384, N349);
xor XOR2 (N388, N379, N360);
xor XOR2 (N389, N87, N310);
nand NAND3 (N390, N382, N268, N301);
xor XOR2 (N391, N381, N13);
nand NAND4 (N392, N387, N283, N46, N152);
or OR4 (N393, N391, N301, N340, N38);
buf BUF1 (N394, N370);
and AND4 (N395, N373, N178, N250, N348);
buf BUF1 (N396, N395);
and AND3 (N397, N393, N145, N324);
nor NOR2 (N398, N389, N29);
or OR4 (N399, N390, N76, N204, N85);
xor XOR2 (N400, N397, N188);
xor XOR2 (N401, N386, N93);
nand NAND2 (N402, N399, N342);
and AND2 (N403, N402, N363);
or OR2 (N404, N401, N254);
and AND4 (N405, N396, N82, N343, N219);
buf BUF1 (N406, N404);
nor NOR4 (N407, N406, N43, N120, N325);
nand NAND4 (N408, N407, N195, N370, N290);
or OR2 (N409, N398, N198);
xor XOR2 (N410, N408, N103);
or OR4 (N411, N371, N7, N27, N214);
xor XOR2 (N412, N409, N163);
xor XOR2 (N413, N405, N135);
nand NAND3 (N414, N388, N105, N104);
nand NAND2 (N415, N392, N380);
nand NAND3 (N416, N415, N257, N172);
not NOT1 (N417, N414);
not NOT1 (N418, N416);
not NOT1 (N419, N418);
and AND2 (N420, N413, N297);
not NOT1 (N421, N411);
or OR3 (N422, N410, N401, N5);
nor NOR2 (N423, N417, N114);
or OR3 (N424, N421, N55, N177);
xor XOR2 (N425, N422, N344);
buf BUF1 (N426, N400);
xor XOR2 (N427, N403, N332);
and AND2 (N428, N394, N300);
and AND4 (N429, N427, N423, N331, N59);
not NOT1 (N430, N335);
nor NOR2 (N431, N385, N232);
xor XOR2 (N432, N420, N403);
buf BUF1 (N433, N428);
not NOT1 (N434, N431);
nand NAND3 (N435, N425, N354, N166);
nand NAND3 (N436, N432, N176, N3);
nand NAND3 (N437, N419, N204, N348);
buf BUF1 (N438, N436);
or OR4 (N439, N435, N323, N260, N144);
buf BUF1 (N440, N424);
xor XOR2 (N441, N430, N239);
xor XOR2 (N442, N439, N103);
nor NOR2 (N443, N412, N265);
or OR3 (N444, N441, N49, N126);
and AND2 (N445, N437, N144);
xor XOR2 (N446, N429, N435);
or OR3 (N447, N443, N306, N135);
xor XOR2 (N448, N440, N431);
xor XOR2 (N449, N438, N287);
and AND3 (N450, N444, N405, N347);
or OR4 (N451, N426, N26, N415, N201);
xor XOR2 (N452, N446, N63);
or OR2 (N453, N452, N46);
and AND4 (N454, N433, N52, N446, N221);
buf BUF1 (N455, N453);
xor XOR2 (N456, N448, N306);
buf BUF1 (N457, N450);
xor XOR2 (N458, N457, N410);
nor NOR3 (N459, N451, N66, N441);
not NOT1 (N460, N458);
not NOT1 (N461, N456);
xor XOR2 (N462, N445, N416);
not NOT1 (N463, N442);
nor NOR3 (N464, N447, N164, N6);
and AND2 (N465, N461, N41);
nor NOR2 (N466, N459, N63);
nor NOR2 (N467, N465, N244);
not NOT1 (N468, N449);
and AND3 (N469, N468, N222, N343);
or OR3 (N470, N462, N257, N396);
or OR2 (N471, N454, N133);
nor NOR2 (N472, N463, N254);
xor XOR2 (N473, N434, N75);
buf BUF1 (N474, N467);
buf BUF1 (N475, N474);
and AND2 (N476, N471, N322);
xor XOR2 (N477, N460, N93);
nor NOR3 (N478, N477, N39, N266);
and AND3 (N479, N466, N49, N400);
or OR3 (N480, N475, N452, N321);
nand NAND4 (N481, N464, N225, N101, N196);
buf BUF1 (N482, N455);
buf BUF1 (N483, N470);
buf BUF1 (N484, N483);
and AND4 (N485, N478, N445, N39, N10);
nand NAND2 (N486, N479, N444);
or OR2 (N487, N485, N347);
xor XOR2 (N488, N469, N323);
nand NAND2 (N489, N484, N161);
xor XOR2 (N490, N487, N101);
buf BUF1 (N491, N486);
xor XOR2 (N492, N473, N280);
xor XOR2 (N493, N476, N489);
buf BUF1 (N494, N226);
not NOT1 (N495, N494);
nand NAND4 (N496, N482, N285, N305, N421);
xor XOR2 (N497, N495, N158);
xor XOR2 (N498, N496, N431);
and AND2 (N499, N492, N356);
buf BUF1 (N500, N472);
and AND3 (N501, N497, N483, N389);
nor NOR3 (N502, N480, N225, N473);
nor NOR3 (N503, N481, N65, N314);
nand NAND2 (N504, N501, N315);
xor XOR2 (N505, N498, N255);
nor NOR4 (N506, N503, N333, N234, N35);
not NOT1 (N507, N499);
xor XOR2 (N508, N488, N323);
nand NAND3 (N509, N500, N495, N130);
or OR4 (N510, N493, N351, N321, N320);
nand NAND2 (N511, N510, N464);
or OR3 (N512, N508, N421, N228);
not NOT1 (N513, N505);
nand NAND2 (N514, N509, N361);
and AND3 (N515, N490, N248, N313);
nand NAND2 (N516, N512, N108);
xor XOR2 (N517, N516, N420);
nand NAND2 (N518, N514, N305);
not NOT1 (N519, N506);
nor NOR2 (N520, N507, N133);
xor XOR2 (N521, N519, N409);
or OR4 (N522, N513, N63, N119, N324);
buf BUF1 (N523, N522);
and AND4 (N524, N491, N33, N60, N223);
and AND4 (N525, N511, N515, N284, N509);
nand NAND4 (N526, N19, N78, N173, N377);
nand NAND3 (N527, N517, N175, N212);
or OR3 (N528, N524, N150, N251);
buf BUF1 (N529, N504);
or OR2 (N530, N526, N99);
nand NAND4 (N531, N523, N434, N284, N351);
or OR3 (N532, N530, N4, N427);
xor XOR2 (N533, N520, N408);
xor XOR2 (N534, N527, N135);
and AND3 (N535, N531, N377, N302);
nand NAND4 (N536, N521, N476, N292, N192);
buf BUF1 (N537, N529);
and AND2 (N538, N534, N222);
nor NOR3 (N539, N532, N115, N423);
nor NOR3 (N540, N528, N142, N226);
xor XOR2 (N541, N536, N38);
buf BUF1 (N542, N541);
xor XOR2 (N543, N542, N415);
or OR3 (N544, N502, N66, N181);
nand NAND3 (N545, N544, N459, N58);
nor NOR3 (N546, N533, N67, N399);
not NOT1 (N547, N540);
and AND4 (N548, N518, N172, N126, N410);
nor NOR2 (N549, N546, N330);
and AND3 (N550, N537, N540, N466);
buf BUF1 (N551, N545);
or OR4 (N552, N548, N9, N409, N127);
or OR3 (N553, N552, N95, N99);
not NOT1 (N554, N549);
buf BUF1 (N555, N550);
not NOT1 (N556, N553);
nor NOR3 (N557, N543, N371, N3);
not NOT1 (N558, N535);
and AND4 (N559, N547, N85, N386, N344);
xor XOR2 (N560, N539, N299);
and AND2 (N561, N554, N15);
nor NOR3 (N562, N558, N127, N214);
not NOT1 (N563, N559);
not NOT1 (N564, N555);
buf BUF1 (N565, N561);
xor XOR2 (N566, N563, N325);
or OR4 (N567, N557, N453, N138, N7);
not NOT1 (N568, N564);
nand NAND3 (N569, N538, N203, N429);
xor XOR2 (N570, N525, N282);
and AND4 (N571, N566, N57, N304, N180);
buf BUF1 (N572, N567);
nand NAND4 (N573, N568, N319, N17, N212);
and AND2 (N574, N565, N185);
nand NAND2 (N575, N569, N247);
or OR2 (N576, N571, N251);
or OR3 (N577, N551, N478, N434);
not NOT1 (N578, N562);
not NOT1 (N579, N577);
not NOT1 (N580, N573);
or OR3 (N581, N572, N284, N195);
xor XOR2 (N582, N556, N575);
buf BUF1 (N583, N574);
and AND4 (N584, N251, N418, N174, N130);
or OR3 (N585, N560, N536, N18);
not NOT1 (N586, N585);
xor XOR2 (N587, N584, N415);
or OR3 (N588, N570, N158, N203);
buf BUF1 (N589, N587);
nand NAND2 (N590, N578, N505);
not NOT1 (N591, N588);
xor XOR2 (N592, N591, N400);
nor NOR3 (N593, N583, N547, N436);
xor XOR2 (N594, N593, N305);
buf BUF1 (N595, N594);
nand NAND4 (N596, N581, N457, N260, N120);
or OR3 (N597, N592, N456, N140);
xor XOR2 (N598, N597, N249);
or OR2 (N599, N598, N153);
or OR2 (N600, N576, N138);
not NOT1 (N601, N595);
and AND3 (N602, N579, N298, N449);
and AND2 (N603, N596, N195);
not NOT1 (N604, N586);
buf BUF1 (N605, N603);
xor XOR2 (N606, N582, N428);
and AND3 (N607, N606, N457, N605);
and AND4 (N608, N393, N565, N135, N359);
not NOT1 (N609, N599);
not NOT1 (N610, N589);
and AND3 (N611, N601, N23, N488);
nand NAND4 (N612, N590, N452, N13, N4);
nor NOR2 (N613, N610, N251);
xor XOR2 (N614, N608, N74);
and AND3 (N615, N614, N442, N199);
or OR2 (N616, N600, N472);
and AND2 (N617, N611, N22);
nor NOR4 (N618, N615, N164, N315, N483);
nor NOR2 (N619, N604, N15);
or OR4 (N620, N616, N517, N116, N117);
and AND4 (N621, N620, N591, N245, N606);
buf BUF1 (N622, N613);
nand NAND2 (N623, N607, N118);
and AND2 (N624, N619, N295);
buf BUF1 (N625, N609);
or OR4 (N626, N624, N46, N295, N314);
not NOT1 (N627, N626);
and AND2 (N628, N625, N602);
and AND4 (N629, N39, N31, N469, N168);
nand NAND4 (N630, N629, N212, N525, N403);
nor NOR4 (N631, N623, N166, N461, N108);
xor XOR2 (N632, N617, N161);
and AND4 (N633, N618, N425, N632, N2);
nand NAND3 (N634, N470, N592, N633);
not NOT1 (N635, N415);
not NOT1 (N636, N621);
and AND4 (N637, N631, N444, N33, N347);
and AND3 (N638, N580, N306, N602);
and AND3 (N639, N612, N161, N151);
and AND3 (N640, N622, N628, N259);
nand NAND2 (N641, N617, N193);
or OR2 (N642, N639, N497);
xor XOR2 (N643, N627, N216);
or OR4 (N644, N642, N533, N127, N87);
not NOT1 (N645, N636);
and AND2 (N646, N635, N443);
or OR2 (N647, N638, N224);
nor NOR4 (N648, N630, N540, N34, N385);
buf BUF1 (N649, N646);
xor XOR2 (N650, N643, N247);
nor NOR3 (N651, N640, N483, N334);
nand NAND4 (N652, N648, N197, N318, N557);
nand NAND2 (N653, N647, N509);
xor XOR2 (N654, N637, N322);
nand NAND2 (N655, N652, N284);
or OR4 (N656, N644, N633, N633, N268);
xor XOR2 (N657, N654, N309);
buf BUF1 (N658, N655);
nand NAND2 (N659, N649, N368);
not NOT1 (N660, N653);
and AND2 (N661, N660, N194);
buf BUF1 (N662, N634);
nor NOR2 (N663, N641, N236);
and AND3 (N664, N662, N167, N610);
nand NAND4 (N665, N658, N628, N433, N315);
buf BUF1 (N666, N659);
buf BUF1 (N667, N661);
or OR4 (N668, N664, N49, N379, N623);
buf BUF1 (N669, N657);
and AND2 (N670, N668, N331);
and AND4 (N671, N669, N617, N224, N6);
xor XOR2 (N672, N651, N668);
nand NAND3 (N673, N667, N544, N517);
nand NAND4 (N674, N656, N56, N149, N314);
and AND4 (N675, N673, N242, N128, N471);
xor XOR2 (N676, N665, N469);
not NOT1 (N677, N674);
not NOT1 (N678, N672);
and AND4 (N679, N663, N74, N87, N210);
nor NOR2 (N680, N650, N302);
nor NOR3 (N681, N680, N112, N161);
and AND3 (N682, N671, N286, N206);
nor NOR2 (N683, N676, N196);
xor XOR2 (N684, N645, N393);
or OR4 (N685, N666, N135, N456, N313);
or OR2 (N686, N683, N382);
or OR3 (N687, N685, N510, N521);
nand NAND4 (N688, N681, N233, N273, N578);
not NOT1 (N689, N687);
and AND2 (N690, N682, N208);
nand NAND2 (N691, N688, N90);
buf BUF1 (N692, N675);
or OR4 (N693, N689, N276, N536, N366);
xor XOR2 (N694, N670, N28);
nand NAND4 (N695, N691, N671, N95, N317);
and AND3 (N696, N690, N318, N588);
and AND3 (N697, N686, N343, N112);
or OR3 (N698, N684, N503, N267);
nor NOR3 (N699, N693, N383, N211);
buf BUF1 (N700, N696);
not NOT1 (N701, N700);
xor XOR2 (N702, N699, N123);
xor XOR2 (N703, N698, N597);
or OR2 (N704, N677, N69);
not NOT1 (N705, N695);
nand NAND2 (N706, N704, N673);
xor XOR2 (N707, N678, N99);
or OR4 (N708, N694, N66, N261, N422);
xor XOR2 (N709, N679, N689);
not NOT1 (N710, N701);
nand NAND3 (N711, N709, N285, N248);
and AND3 (N712, N710, N532, N501);
nor NOR2 (N713, N692, N262);
or OR2 (N714, N706, N3);
or OR2 (N715, N713, N474);
and AND2 (N716, N707, N334);
nand NAND3 (N717, N703, N11, N679);
not NOT1 (N718, N715);
or OR3 (N719, N702, N255, N514);
xor XOR2 (N720, N718, N568);
not NOT1 (N721, N711);
nor NOR2 (N722, N717, N346);
nor NOR2 (N723, N720, N464);
not NOT1 (N724, N705);
xor XOR2 (N725, N712, N240);
nand NAND3 (N726, N722, N242, N287);
xor XOR2 (N727, N716, N245);
xor XOR2 (N728, N708, N393);
nand NAND4 (N729, N719, N655, N333, N483);
or OR4 (N730, N725, N218, N192, N121);
not NOT1 (N731, N727);
and AND2 (N732, N730, N329);
nand NAND3 (N733, N724, N710, N655);
nor NOR3 (N734, N726, N345, N449);
nor NOR3 (N735, N733, N37, N386);
or OR2 (N736, N697, N186);
not NOT1 (N737, N714);
nor NOR4 (N738, N723, N67, N640, N78);
buf BUF1 (N739, N729);
xor XOR2 (N740, N732, N642);
and AND2 (N741, N728, N565);
buf BUF1 (N742, N721);
buf BUF1 (N743, N735);
nor NOR3 (N744, N739, N247, N477);
xor XOR2 (N745, N744, N294);
buf BUF1 (N746, N737);
or OR2 (N747, N731, N686);
nor NOR3 (N748, N745, N331, N407);
nand NAND3 (N749, N748, N217, N29);
nand NAND4 (N750, N741, N502, N385, N68);
nand NAND4 (N751, N734, N179, N516, N356);
and AND3 (N752, N746, N65, N162);
nor NOR4 (N753, N738, N78, N549, N207);
buf BUF1 (N754, N742);
and AND2 (N755, N753, N237);
or OR2 (N756, N743, N48);
nand NAND3 (N757, N752, N270, N29);
xor XOR2 (N758, N747, N546);
nand NAND4 (N759, N758, N98, N569, N713);
or OR3 (N760, N757, N93, N291);
nor NOR4 (N761, N754, N97, N659, N12);
xor XOR2 (N762, N751, N633);
nand NAND3 (N763, N761, N60, N589);
and AND3 (N764, N756, N588, N572);
and AND3 (N765, N749, N445, N700);
and AND4 (N766, N750, N603, N2, N435);
or OR3 (N767, N755, N327, N604);
nor NOR2 (N768, N760, N30);
xor XOR2 (N769, N736, N386);
and AND2 (N770, N762, N559);
or OR4 (N771, N767, N725, N483, N451);
not NOT1 (N772, N740);
nand NAND4 (N773, N768, N147, N332, N307);
not NOT1 (N774, N770);
or OR3 (N775, N769, N733, N258);
nand NAND2 (N776, N763, N64);
xor XOR2 (N777, N766, N156);
buf BUF1 (N778, N776);
and AND4 (N779, N765, N475, N172, N291);
or OR4 (N780, N779, N127, N643, N224);
and AND2 (N781, N759, N701);
and AND2 (N782, N778, N80);
or OR2 (N783, N781, N522);
xor XOR2 (N784, N780, N124);
and AND3 (N785, N777, N115, N260);
nor NOR3 (N786, N773, N247, N719);
or OR4 (N787, N782, N218, N295, N235);
nor NOR3 (N788, N771, N340, N595);
and AND3 (N789, N783, N592, N253);
or OR2 (N790, N789, N315);
buf BUF1 (N791, N787);
xor XOR2 (N792, N788, N545);
and AND4 (N793, N791, N243, N525, N705);
xor XOR2 (N794, N792, N759);
nand NAND4 (N795, N764, N170, N482, N11);
nand NAND4 (N796, N793, N594, N668, N579);
xor XOR2 (N797, N785, N417);
and AND2 (N798, N786, N782);
nor NOR3 (N799, N796, N254, N126);
and AND4 (N800, N772, N364, N765, N589);
xor XOR2 (N801, N794, N89);
buf BUF1 (N802, N795);
buf BUF1 (N803, N799);
and AND4 (N804, N800, N321, N733, N360);
buf BUF1 (N805, N797);
xor XOR2 (N806, N804, N124);
buf BUF1 (N807, N775);
xor XOR2 (N808, N802, N654);
or OR3 (N809, N790, N725, N321);
or OR4 (N810, N806, N588, N606, N474);
xor XOR2 (N811, N803, N473);
nor NOR3 (N812, N784, N727, N704);
buf BUF1 (N813, N809);
and AND4 (N814, N810, N469, N622, N710);
xor XOR2 (N815, N805, N535);
not NOT1 (N816, N807);
and AND2 (N817, N815, N43);
xor XOR2 (N818, N817, N174);
and AND4 (N819, N801, N451, N83, N185);
xor XOR2 (N820, N811, N784);
nor NOR4 (N821, N813, N566, N277, N231);
or OR2 (N822, N774, N619);
nor NOR2 (N823, N820, N16);
nor NOR4 (N824, N816, N240, N195, N161);
xor XOR2 (N825, N808, N758);
nor NOR2 (N826, N812, N195);
buf BUF1 (N827, N798);
buf BUF1 (N828, N827);
and AND3 (N829, N822, N266, N294);
nand NAND3 (N830, N823, N15, N748);
not NOT1 (N831, N830);
not NOT1 (N832, N821);
nor NOR4 (N833, N826, N728, N204, N35);
nor NOR2 (N834, N833, N605);
nor NOR2 (N835, N829, N129);
xor XOR2 (N836, N824, N777);
or OR2 (N837, N828, N512);
or OR3 (N838, N814, N231, N38);
nor NOR3 (N839, N836, N90, N423);
xor XOR2 (N840, N819, N227);
not NOT1 (N841, N838);
nand NAND3 (N842, N818, N261, N396);
buf BUF1 (N843, N831);
xor XOR2 (N844, N837, N592);
and AND3 (N845, N832, N236, N722);
or OR3 (N846, N834, N360, N597);
xor XOR2 (N847, N841, N801);
not NOT1 (N848, N840);
not NOT1 (N849, N835);
buf BUF1 (N850, N848);
nand NAND4 (N851, N843, N533, N80, N619);
or OR3 (N852, N839, N562, N829);
nand NAND3 (N853, N852, N626, N455);
xor XOR2 (N854, N849, N339);
buf BUF1 (N855, N853);
and AND4 (N856, N845, N13, N627, N758);
or OR2 (N857, N856, N677);
or OR3 (N858, N855, N818, N671);
buf BUF1 (N859, N851);
and AND2 (N860, N859, N5);
nor NOR4 (N861, N844, N324, N369, N441);
and AND2 (N862, N854, N607);
and AND4 (N863, N850, N226, N314, N741);
xor XOR2 (N864, N858, N852);
nand NAND4 (N865, N842, N44, N509, N585);
xor XOR2 (N866, N864, N538);
and AND2 (N867, N847, N502);
not NOT1 (N868, N865);
and AND4 (N869, N868, N406, N362, N695);
buf BUF1 (N870, N867);
xor XOR2 (N871, N825, N49);
or OR2 (N872, N862, N617);
xor XOR2 (N873, N860, N713);
or OR2 (N874, N870, N662);
or OR3 (N875, N866, N237, N386);
buf BUF1 (N876, N857);
not NOT1 (N877, N871);
buf BUF1 (N878, N876);
or OR2 (N879, N861, N463);
not NOT1 (N880, N869);
not NOT1 (N881, N874);
not NOT1 (N882, N878);
not NOT1 (N883, N872);
nor NOR2 (N884, N880, N429);
not NOT1 (N885, N877);
nor NOR4 (N886, N885, N73, N112, N689);
buf BUF1 (N887, N846);
not NOT1 (N888, N887);
nand NAND2 (N889, N873, N315);
nor NOR2 (N890, N879, N556);
or OR3 (N891, N875, N713, N652);
not NOT1 (N892, N890);
or OR4 (N893, N892, N133, N763, N481);
or OR2 (N894, N881, N391);
and AND3 (N895, N884, N274, N515);
buf BUF1 (N896, N894);
buf BUF1 (N897, N889);
and AND2 (N898, N882, N863);
buf BUF1 (N899, N894);
nand NAND4 (N900, N895, N133, N373, N297);
xor XOR2 (N901, N899, N639);
nand NAND4 (N902, N898, N198, N735, N665);
buf BUF1 (N903, N883);
nor NOR3 (N904, N900, N619, N372);
nor NOR4 (N905, N903, N225, N793, N94);
or OR3 (N906, N897, N274, N215);
nand NAND4 (N907, N896, N513, N354, N835);
not NOT1 (N908, N905);
or OR4 (N909, N907, N517, N12, N636);
or OR4 (N910, N901, N344, N216, N130);
and AND2 (N911, N909, N553);
nand NAND3 (N912, N911, N727, N537);
or OR4 (N913, N886, N339, N535, N210);
nand NAND2 (N914, N906, N223);
nor NOR2 (N915, N893, N159);
buf BUF1 (N916, N902);
and AND4 (N917, N891, N153, N63, N899);
and AND3 (N918, N910, N417, N743);
and AND4 (N919, N888, N167, N125, N791);
and AND4 (N920, N914, N415, N365, N26);
buf BUF1 (N921, N916);
buf BUF1 (N922, N913);
and AND2 (N923, N915, N869);
and AND3 (N924, N908, N868, N245);
and AND3 (N925, N918, N281, N444);
not NOT1 (N926, N919);
buf BUF1 (N927, N924);
nand NAND3 (N928, N926, N558, N510);
nor NOR4 (N929, N922, N417, N50, N130);
nand NAND2 (N930, N925, N836);
not NOT1 (N931, N927);
xor XOR2 (N932, N928, N354);
xor XOR2 (N933, N904, N369);
nor NOR3 (N934, N929, N563, N679);
or OR3 (N935, N934, N335, N576);
nor NOR4 (N936, N930, N726, N92, N115);
buf BUF1 (N937, N921);
nand NAND2 (N938, N932, N195);
nor NOR4 (N939, N933, N771, N875, N45);
or OR3 (N940, N937, N484, N461);
xor XOR2 (N941, N938, N874);
and AND4 (N942, N923, N889, N231, N365);
nor NOR4 (N943, N942, N287, N864, N839);
nor NOR4 (N944, N917, N20, N85, N643);
buf BUF1 (N945, N920);
nand NAND3 (N946, N940, N821, N799);
or OR2 (N947, N936, N401);
buf BUF1 (N948, N943);
not NOT1 (N949, N935);
or OR2 (N950, N946, N280);
buf BUF1 (N951, N939);
or OR2 (N952, N945, N751);
and AND2 (N953, N952, N539);
nor NOR4 (N954, N947, N914, N641, N439);
and AND4 (N955, N941, N680, N107, N433);
buf BUF1 (N956, N931);
nand NAND4 (N957, N954, N590, N344, N651);
not NOT1 (N958, N948);
nor NOR2 (N959, N953, N561);
and AND3 (N960, N958, N909, N559);
xor XOR2 (N961, N959, N551);
and AND4 (N962, N950, N333, N803, N134);
nand NAND2 (N963, N949, N653);
not NOT1 (N964, N912);
nand NAND4 (N965, N957, N710, N342, N819);
buf BUF1 (N966, N962);
buf BUF1 (N967, N964);
or OR3 (N968, N966, N622, N661);
xor XOR2 (N969, N951, N922);
nand NAND2 (N970, N963, N320);
xor XOR2 (N971, N960, N277);
xor XOR2 (N972, N961, N350);
xor XOR2 (N973, N944, N317);
nand NAND2 (N974, N969, N188);
not NOT1 (N975, N967);
buf BUF1 (N976, N956);
or OR3 (N977, N968, N498, N861);
nor NOR4 (N978, N970, N101, N462, N308);
buf BUF1 (N979, N976);
nand NAND2 (N980, N974, N263);
nand NAND2 (N981, N971, N505);
and AND2 (N982, N980, N973);
xor XOR2 (N983, N488, N423);
not NOT1 (N984, N975);
xor XOR2 (N985, N965, N753);
buf BUF1 (N986, N983);
nand NAND3 (N987, N985, N909, N391);
and AND2 (N988, N984, N831);
buf BUF1 (N989, N972);
or OR2 (N990, N978, N365);
not NOT1 (N991, N982);
and AND4 (N992, N979, N133, N715, N35);
xor XOR2 (N993, N955, N9);
xor XOR2 (N994, N993, N681);
or OR2 (N995, N987, N879);
not NOT1 (N996, N977);
xor XOR2 (N997, N989, N269);
nor NOR3 (N998, N995, N366, N851);
nor NOR2 (N999, N992, N468);
xor XOR2 (N1000, N990, N57);
or OR4 (N1001, N999, N649, N531, N844);
buf BUF1 (N1002, N1001);
and AND2 (N1003, N1000, N196);
buf BUF1 (N1004, N986);
buf BUF1 (N1005, N988);
not NOT1 (N1006, N981);
xor XOR2 (N1007, N1004, N408);
or OR4 (N1008, N1003, N572, N63, N3);
not NOT1 (N1009, N1002);
nand NAND2 (N1010, N1009, N492);
not NOT1 (N1011, N998);
xor XOR2 (N1012, N996, N78);
not NOT1 (N1013, N1010);
nor NOR4 (N1014, N1012, N841, N21, N959);
or OR2 (N1015, N1005, N558);
buf BUF1 (N1016, N1011);
and AND3 (N1017, N994, N885, N401);
nor NOR4 (N1018, N1017, N414, N619, N287);
nor NOR3 (N1019, N1014, N446, N370);
and AND3 (N1020, N1016, N39, N589);
or OR3 (N1021, N1020, N725, N637);
nor NOR3 (N1022, N997, N621, N81);
nand NAND2 (N1023, N1007, N243);
xor XOR2 (N1024, N1023, N64);
not NOT1 (N1025, N1013);
not NOT1 (N1026, N1024);
buf BUF1 (N1027, N1018);
nand NAND4 (N1028, N1006, N383, N219, N189);
nand NAND2 (N1029, N991, N462);
not NOT1 (N1030, N1027);
xor XOR2 (N1031, N1021, N673);
or OR3 (N1032, N1031, N630, N551);
not NOT1 (N1033, N1028);
nor NOR4 (N1034, N1032, N284, N49, N828);
nor NOR2 (N1035, N1033, N776);
nor NOR3 (N1036, N1015, N796, N524);
buf BUF1 (N1037, N1022);
nor NOR3 (N1038, N1036, N822, N94);
not NOT1 (N1039, N1038);
buf BUF1 (N1040, N1026);
buf BUF1 (N1041, N1019);
nor NOR4 (N1042, N1037, N66, N524, N460);
and AND2 (N1043, N1042, N775);
nor NOR2 (N1044, N1030, N343);
nand NAND3 (N1045, N1040, N776, N587);
nor NOR3 (N1046, N1025, N663, N497);
nand NAND3 (N1047, N1039, N1039, N142);
buf BUF1 (N1048, N1043);
or OR4 (N1049, N1046, N781, N549, N766);
buf BUF1 (N1050, N1049);
buf BUF1 (N1051, N1048);
or OR2 (N1052, N1050, N480);
not NOT1 (N1053, N1041);
and AND3 (N1054, N1045, N327, N193);
or OR2 (N1055, N1047, N327);
buf BUF1 (N1056, N1044);
and AND2 (N1057, N1029, N197);
nand NAND4 (N1058, N1008, N918, N721, N530);
nor NOR4 (N1059, N1055, N982, N657, N28);
and AND4 (N1060, N1059, N398, N718, N986);
nand NAND3 (N1061, N1035, N824, N436);
nand NAND2 (N1062, N1034, N491);
buf BUF1 (N1063, N1057);
nor NOR4 (N1064, N1051, N615, N1036, N295);
buf BUF1 (N1065, N1052);
xor XOR2 (N1066, N1062, N414);
xor XOR2 (N1067, N1058, N870);
nor NOR3 (N1068, N1053, N113, N1017);
nand NAND3 (N1069, N1054, N450, N194);
or OR3 (N1070, N1056, N98, N385);
or OR2 (N1071, N1067, N714);
xor XOR2 (N1072, N1064, N117);
nor NOR3 (N1073, N1061, N1020, N356);
xor XOR2 (N1074, N1068, N967);
nor NOR3 (N1075, N1070, N10, N262);
nand NAND3 (N1076, N1075, N482, N968);
and AND2 (N1077, N1063, N999);
xor XOR2 (N1078, N1071, N23);
or OR3 (N1079, N1066, N868, N687);
and AND2 (N1080, N1076, N572);
xor XOR2 (N1081, N1072, N566);
buf BUF1 (N1082, N1060);
nor NOR4 (N1083, N1078, N572, N141, N335);
buf BUF1 (N1084, N1080);
and AND3 (N1085, N1065, N857, N946);
buf BUF1 (N1086, N1081);
not NOT1 (N1087, N1073);
nor NOR2 (N1088, N1087, N189);
not NOT1 (N1089, N1082);
nand NAND3 (N1090, N1084, N507, N989);
not NOT1 (N1091, N1077);
and AND3 (N1092, N1090, N278, N1014);
not NOT1 (N1093, N1091);
buf BUF1 (N1094, N1069);
xor XOR2 (N1095, N1088, N360);
xor XOR2 (N1096, N1074, N474);
not NOT1 (N1097, N1086);
xor XOR2 (N1098, N1079, N997);
nor NOR2 (N1099, N1096, N789);
or OR2 (N1100, N1089, N571);
nand NAND2 (N1101, N1092, N757);
xor XOR2 (N1102, N1098, N1021);
and AND4 (N1103, N1085, N473, N657, N208);
buf BUF1 (N1104, N1103);
nor NOR4 (N1105, N1099, N1024, N118, N497);
or OR3 (N1106, N1102, N446, N361);
xor XOR2 (N1107, N1097, N954);
or OR2 (N1108, N1083, N699);
not NOT1 (N1109, N1105);
xor XOR2 (N1110, N1104, N997);
nor NOR4 (N1111, N1107, N305, N765, N876);
and AND4 (N1112, N1109, N937, N702, N622);
not NOT1 (N1113, N1094);
or OR4 (N1114, N1111, N626, N537, N805);
nand NAND4 (N1115, N1095, N123, N302, N176);
xor XOR2 (N1116, N1115, N925);
not NOT1 (N1117, N1112);
and AND3 (N1118, N1110, N594, N922);
buf BUF1 (N1119, N1093);
xor XOR2 (N1120, N1116, N910);
not NOT1 (N1121, N1119);
or OR4 (N1122, N1108, N383, N1109, N443);
buf BUF1 (N1123, N1101);
buf BUF1 (N1124, N1122);
or OR2 (N1125, N1120, N471);
not NOT1 (N1126, N1118);
nand NAND3 (N1127, N1123, N229, N248);
and AND3 (N1128, N1100, N930, N854);
and AND4 (N1129, N1106, N728, N831, N370);
and AND3 (N1130, N1126, N339, N153);
nor NOR3 (N1131, N1117, N765, N701);
buf BUF1 (N1132, N1125);
and AND2 (N1133, N1121, N791);
and AND3 (N1134, N1129, N240, N1123);
not NOT1 (N1135, N1133);
or OR2 (N1136, N1134, N463);
nand NAND2 (N1137, N1130, N68);
buf BUF1 (N1138, N1124);
and AND2 (N1139, N1136, N1010);
not NOT1 (N1140, N1113);
buf BUF1 (N1141, N1140);
nand NAND2 (N1142, N1141, N108);
xor XOR2 (N1143, N1127, N46);
nor NOR4 (N1144, N1132, N551, N256, N648);
xor XOR2 (N1145, N1131, N988);
and AND4 (N1146, N1139, N736, N796, N938);
not NOT1 (N1147, N1144);
nor NOR2 (N1148, N1128, N359);
not NOT1 (N1149, N1142);
not NOT1 (N1150, N1147);
xor XOR2 (N1151, N1114, N336);
buf BUF1 (N1152, N1138);
or OR2 (N1153, N1145, N2);
not NOT1 (N1154, N1151);
not NOT1 (N1155, N1146);
xor XOR2 (N1156, N1154, N377);
not NOT1 (N1157, N1148);
or OR4 (N1158, N1152, N205, N538, N738);
and AND2 (N1159, N1156, N895);
buf BUF1 (N1160, N1157);
nor NOR2 (N1161, N1135, N828);
nand NAND3 (N1162, N1153, N295, N935);
or OR4 (N1163, N1159, N729, N979, N961);
nand NAND2 (N1164, N1158, N894);
xor XOR2 (N1165, N1149, N188);
or OR3 (N1166, N1165, N995, N1066);
xor XOR2 (N1167, N1137, N65);
not NOT1 (N1168, N1163);
nor NOR2 (N1169, N1161, N509);
nor NOR2 (N1170, N1167, N826);
buf BUF1 (N1171, N1162);
or OR4 (N1172, N1143, N564, N744, N144);
not NOT1 (N1173, N1170);
not NOT1 (N1174, N1173);
not NOT1 (N1175, N1174);
nor NOR2 (N1176, N1169, N654);
or OR3 (N1177, N1172, N992, N607);
or OR4 (N1178, N1164, N777, N453, N1027);
buf BUF1 (N1179, N1155);
nand NAND3 (N1180, N1160, N630, N305);
and AND2 (N1181, N1179, N171);
nor NOR2 (N1182, N1171, N252);
nor NOR3 (N1183, N1175, N83, N120);
or OR2 (N1184, N1182, N683);
xor XOR2 (N1185, N1166, N42);
nor NOR4 (N1186, N1180, N905, N330, N629);
xor XOR2 (N1187, N1185, N859);
nor NOR4 (N1188, N1168, N817, N820, N988);
xor XOR2 (N1189, N1188, N172);
buf BUF1 (N1190, N1183);
xor XOR2 (N1191, N1177, N921);
not NOT1 (N1192, N1178);
nand NAND4 (N1193, N1191, N729, N238, N951);
not NOT1 (N1194, N1150);
nor NOR3 (N1195, N1186, N251, N129);
xor XOR2 (N1196, N1190, N1042);
or OR2 (N1197, N1196, N2);
buf BUF1 (N1198, N1193);
nor NOR3 (N1199, N1189, N754, N840);
buf BUF1 (N1200, N1195);
nor NOR3 (N1201, N1176, N836, N1035);
xor XOR2 (N1202, N1199, N1117);
nand NAND2 (N1203, N1192, N702);
xor XOR2 (N1204, N1198, N470);
not NOT1 (N1205, N1203);
xor XOR2 (N1206, N1197, N1045);
and AND3 (N1207, N1184, N187, N714);
or OR4 (N1208, N1181, N643, N532, N635);
nor NOR4 (N1209, N1202, N870, N1065, N898);
xor XOR2 (N1210, N1207, N898);
nor NOR4 (N1211, N1206, N76, N976, N127);
not NOT1 (N1212, N1201);
buf BUF1 (N1213, N1205);
buf BUF1 (N1214, N1211);
or OR2 (N1215, N1209, N958);
nand NAND3 (N1216, N1213, N1090, N981);
nand NAND3 (N1217, N1216, N792, N918);
nor NOR4 (N1218, N1212, N366, N1157, N756);
xor XOR2 (N1219, N1215, N815);
nor NOR3 (N1220, N1218, N15, N1043);
nor NOR4 (N1221, N1220, N68, N486, N1121);
nand NAND3 (N1222, N1219, N596, N765);
not NOT1 (N1223, N1222);
nor NOR3 (N1224, N1214, N459, N706);
nand NAND2 (N1225, N1210, N21);
and AND4 (N1226, N1208, N920, N528, N986);
nor NOR4 (N1227, N1221, N215, N276, N860);
nand NAND4 (N1228, N1224, N272, N1048, N570);
buf BUF1 (N1229, N1204);
or OR3 (N1230, N1225, N1031, N260);
not NOT1 (N1231, N1227);
nor NOR3 (N1232, N1217, N153, N123);
nand NAND3 (N1233, N1230, N306, N1213);
or OR2 (N1234, N1233, N862);
xor XOR2 (N1235, N1200, N1037);
nand NAND3 (N1236, N1223, N698, N173);
xor XOR2 (N1237, N1234, N9);
buf BUF1 (N1238, N1235);
nor NOR2 (N1239, N1238, N612);
and AND4 (N1240, N1187, N830, N723, N120);
nand NAND3 (N1241, N1232, N220, N829);
xor XOR2 (N1242, N1241, N940);
and AND2 (N1243, N1228, N1177);
nand NAND3 (N1244, N1237, N1242, N1181);
xor XOR2 (N1245, N165, N794);
xor XOR2 (N1246, N1226, N802);
nand NAND3 (N1247, N1243, N1050, N253);
not NOT1 (N1248, N1246);
buf BUF1 (N1249, N1231);
xor XOR2 (N1250, N1229, N223);
nand NAND3 (N1251, N1249, N1095, N147);
nor NOR2 (N1252, N1236, N4);
xor XOR2 (N1253, N1252, N623);
nand NAND3 (N1254, N1253, N868, N774);
and AND2 (N1255, N1254, N409);
buf BUF1 (N1256, N1239);
xor XOR2 (N1257, N1250, N969);
nor NOR4 (N1258, N1244, N1232, N405, N509);
xor XOR2 (N1259, N1248, N1167);
or OR4 (N1260, N1255, N512, N1188, N285);
nor NOR4 (N1261, N1245, N1155, N990, N206);
xor XOR2 (N1262, N1258, N833);
not NOT1 (N1263, N1247);
or OR2 (N1264, N1261, N720);
not NOT1 (N1265, N1240);
buf BUF1 (N1266, N1264);
buf BUF1 (N1267, N1262);
buf BUF1 (N1268, N1251);
buf BUF1 (N1269, N1256);
nand NAND2 (N1270, N1268, N798);
buf BUF1 (N1271, N1269);
nor NOR2 (N1272, N1259, N1018);
or OR3 (N1273, N1267, N530, N869);
nand NAND4 (N1274, N1260, N415, N535, N76);
xor XOR2 (N1275, N1274, N769);
xor XOR2 (N1276, N1270, N1152);
not NOT1 (N1277, N1194);
and AND3 (N1278, N1263, N334, N586);
not NOT1 (N1279, N1272);
not NOT1 (N1280, N1278);
nor NOR4 (N1281, N1266, N140, N153, N1257);
or OR3 (N1282, N724, N301, N286);
nor NOR2 (N1283, N1281, N590);
or OR2 (N1284, N1282, N91);
nand NAND4 (N1285, N1275, N561, N646, N92);
and AND3 (N1286, N1284, N402, N697);
xor XOR2 (N1287, N1276, N1059);
not NOT1 (N1288, N1279);
buf BUF1 (N1289, N1280);
or OR3 (N1290, N1283, N874, N1000);
or OR4 (N1291, N1277, N639, N1112, N168);
buf BUF1 (N1292, N1285);
nor NOR4 (N1293, N1291, N7, N700, N280);
or OR2 (N1294, N1290, N395);
and AND4 (N1295, N1287, N752, N1033, N68);
buf BUF1 (N1296, N1292);
and AND2 (N1297, N1271, N185);
nor NOR3 (N1298, N1294, N262, N1215);
nor NOR4 (N1299, N1298, N549, N68, N248);
nand NAND4 (N1300, N1286, N689, N134, N515);
buf BUF1 (N1301, N1289);
nor NOR4 (N1302, N1299, N379, N1090, N882);
or OR3 (N1303, N1301, N22, N188);
xor XOR2 (N1304, N1273, N56);
and AND4 (N1305, N1297, N900, N556, N880);
or OR4 (N1306, N1288, N381, N15, N951);
nor NOR4 (N1307, N1302, N527, N139, N375);
buf BUF1 (N1308, N1307);
or OR4 (N1309, N1265, N128, N300, N803);
buf BUF1 (N1310, N1306);
nor NOR2 (N1311, N1295, N948);
and AND4 (N1312, N1309, N720, N842, N1177);
xor XOR2 (N1313, N1296, N797);
buf BUF1 (N1314, N1310);
xor XOR2 (N1315, N1314, N264);
nand NAND2 (N1316, N1303, N430);
xor XOR2 (N1317, N1304, N1227);
or OR3 (N1318, N1312, N439, N359);
nand NAND4 (N1319, N1313, N925, N1210, N775);
and AND2 (N1320, N1311, N110);
and AND4 (N1321, N1316, N838, N1181, N1256);
not NOT1 (N1322, N1315);
not NOT1 (N1323, N1293);
and AND2 (N1324, N1305, N252);
and AND2 (N1325, N1322, N539);
and AND3 (N1326, N1318, N1186, N530);
xor XOR2 (N1327, N1319, N806);
or OR3 (N1328, N1324, N424, N701);
nor NOR4 (N1329, N1320, N936, N1287, N1313);
xor XOR2 (N1330, N1321, N1180);
and AND2 (N1331, N1330, N220);
not NOT1 (N1332, N1329);
and AND3 (N1333, N1308, N362, N164);
not NOT1 (N1334, N1327);
buf BUF1 (N1335, N1333);
not NOT1 (N1336, N1323);
or OR4 (N1337, N1328, N331, N411, N770);
nor NOR2 (N1338, N1336, N581);
buf BUF1 (N1339, N1325);
xor XOR2 (N1340, N1326, N939);
or OR3 (N1341, N1339, N766, N646);
or OR4 (N1342, N1337, N39, N735, N263);
nor NOR4 (N1343, N1300, N1275, N426, N1133);
or OR4 (N1344, N1331, N1166, N1016, N844);
or OR3 (N1345, N1335, N489, N965);
buf BUF1 (N1346, N1345);
nand NAND2 (N1347, N1340, N92);
xor XOR2 (N1348, N1342, N712);
nand NAND3 (N1349, N1338, N1060, N285);
buf BUF1 (N1350, N1348);
or OR4 (N1351, N1332, N281, N1298, N616);
buf BUF1 (N1352, N1344);
nand NAND3 (N1353, N1352, N305, N639);
not NOT1 (N1354, N1349);
buf BUF1 (N1355, N1350);
and AND4 (N1356, N1341, N71, N1141, N812);
and AND2 (N1357, N1343, N200);
nor NOR2 (N1358, N1357, N650);
nand NAND2 (N1359, N1358, N417);
nand NAND2 (N1360, N1334, N353);
nor NOR2 (N1361, N1360, N1134);
not NOT1 (N1362, N1354);
nand NAND2 (N1363, N1351, N871);
xor XOR2 (N1364, N1347, N964);
nor NOR3 (N1365, N1356, N735, N416);
buf BUF1 (N1366, N1364);
xor XOR2 (N1367, N1355, N172);
not NOT1 (N1368, N1367);
not NOT1 (N1369, N1368);
buf BUF1 (N1370, N1359);
nor NOR2 (N1371, N1346, N185);
nand NAND2 (N1372, N1361, N1365);
buf BUF1 (N1373, N543);
and AND3 (N1374, N1373, N911, N488);
buf BUF1 (N1375, N1371);
xor XOR2 (N1376, N1366, N174);
nor NOR4 (N1377, N1353, N783, N780, N1075);
buf BUF1 (N1378, N1369);
not NOT1 (N1379, N1370);
xor XOR2 (N1380, N1363, N1039);
and AND3 (N1381, N1377, N1092, N1335);
and AND4 (N1382, N1317, N1075, N653, N683);
and AND4 (N1383, N1375, N716, N704, N449);
not NOT1 (N1384, N1382);
nor NOR3 (N1385, N1378, N423, N297);
nand NAND4 (N1386, N1385, N122, N345, N226);
nand NAND4 (N1387, N1362, N136, N753, N1043);
not NOT1 (N1388, N1376);
not NOT1 (N1389, N1388);
not NOT1 (N1390, N1389);
buf BUF1 (N1391, N1390);
xor XOR2 (N1392, N1379, N859);
or OR3 (N1393, N1381, N92, N252);
xor XOR2 (N1394, N1380, N1199);
and AND3 (N1395, N1387, N593, N1339);
nand NAND4 (N1396, N1374, N833, N890, N865);
and AND4 (N1397, N1395, N81, N567, N490);
buf BUF1 (N1398, N1372);
nand NAND2 (N1399, N1383, N801);
and AND3 (N1400, N1392, N1358, N800);
or OR3 (N1401, N1393, N1223, N996);
buf BUF1 (N1402, N1397);
nand NAND2 (N1403, N1402, N284);
nor NOR2 (N1404, N1394, N1211);
not NOT1 (N1405, N1403);
nor NOR2 (N1406, N1401, N1041);
buf BUF1 (N1407, N1405);
or OR4 (N1408, N1399, N1125, N826, N106);
and AND2 (N1409, N1408, N878);
buf BUF1 (N1410, N1396);
nor NOR2 (N1411, N1391, N20);
buf BUF1 (N1412, N1400);
nor NOR2 (N1413, N1386, N462);
and AND2 (N1414, N1398, N694);
nand NAND3 (N1415, N1406, N1065, N1040);
and AND2 (N1416, N1414, N329);
buf BUF1 (N1417, N1416);
nor NOR3 (N1418, N1417, N1250, N1367);
nand NAND2 (N1419, N1412, N416);
buf BUF1 (N1420, N1415);
xor XOR2 (N1421, N1411, N222);
xor XOR2 (N1422, N1410, N674);
or OR3 (N1423, N1421, N1124, N279);
or OR4 (N1424, N1407, N1209, N425, N782);
nor NOR3 (N1425, N1413, N539, N8);
nor NOR2 (N1426, N1422, N189);
and AND2 (N1427, N1424, N239);
buf BUF1 (N1428, N1404);
xor XOR2 (N1429, N1423, N1329);
xor XOR2 (N1430, N1419, N933);
and AND3 (N1431, N1428, N1120, N823);
buf BUF1 (N1432, N1427);
nand NAND4 (N1433, N1418, N403, N1307, N465);
and AND3 (N1434, N1429, N284, N1280);
and AND2 (N1435, N1431, N1285);
nor NOR2 (N1436, N1384, N1199);
not NOT1 (N1437, N1436);
nor NOR2 (N1438, N1420, N328);
buf BUF1 (N1439, N1409);
xor XOR2 (N1440, N1426, N498);
buf BUF1 (N1441, N1425);
buf BUF1 (N1442, N1440);
not NOT1 (N1443, N1434);
and AND2 (N1444, N1430, N543);
or OR2 (N1445, N1442, N493);
or OR3 (N1446, N1443, N527, N1378);
buf BUF1 (N1447, N1435);
not NOT1 (N1448, N1441);
not NOT1 (N1449, N1432);
buf BUF1 (N1450, N1433);
nor NOR4 (N1451, N1447, N1138, N1359, N210);
nor NOR2 (N1452, N1444, N321);
nand NAND4 (N1453, N1452, N345, N1016, N842);
nand NAND2 (N1454, N1448, N995);
xor XOR2 (N1455, N1451, N1330);
and AND3 (N1456, N1446, N460, N978);
buf BUF1 (N1457, N1456);
and AND4 (N1458, N1453, N231, N602, N900);
xor XOR2 (N1459, N1449, N574);
nor NOR4 (N1460, N1439, N1075, N1311, N430);
xor XOR2 (N1461, N1457, N1145);
nand NAND4 (N1462, N1458, N1301, N966, N458);
xor XOR2 (N1463, N1460, N262);
xor XOR2 (N1464, N1445, N1418);
nand NAND3 (N1465, N1438, N399, N1204);
nor NOR3 (N1466, N1454, N4, N1117);
xor XOR2 (N1467, N1464, N360);
xor XOR2 (N1468, N1466, N863);
and AND3 (N1469, N1465, N334, N870);
or OR2 (N1470, N1461, N783);
nor NOR4 (N1471, N1459, N1387, N1385, N619);
not NOT1 (N1472, N1470);
nand NAND4 (N1473, N1467, N627, N268, N178);
nand NAND4 (N1474, N1450, N689, N1416, N197);
buf BUF1 (N1475, N1455);
or OR4 (N1476, N1472, N675, N59, N756);
nand NAND2 (N1477, N1476, N1234);
xor XOR2 (N1478, N1475, N328);
nand NAND3 (N1479, N1469, N671, N300);
buf BUF1 (N1480, N1474);
and AND3 (N1481, N1480, N1451, N1419);
not NOT1 (N1482, N1462);
not NOT1 (N1483, N1482);
nand NAND4 (N1484, N1471, N1422, N860, N98);
nor NOR2 (N1485, N1478, N388);
nand NAND3 (N1486, N1479, N259, N1188);
and AND4 (N1487, N1477, N1265, N646, N141);
xor XOR2 (N1488, N1484, N1158);
nor NOR4 (N1489, N1481, N95, N1312, N186);
xor XOR2 (N1490, N1437, N1470);
and AND4 (N1491, N1468, N818, N671, N494);
nor NOR4 (N1492, N1488, N258, N993, N548);
nand NAND4 (N1493, N1487, N927, N327, N614);
xor XOR2 (N1494, N1490, N210);
and AND4 (N1495, N1463, N638, N802, N1169);
xor XOR2 (N1496, N1494, N162);
xor XOR2 (N1497, N1495, N892);
nor NOR4 (N1498, N1493, N805, N322, N1042);
xor XOR2 (N1499, N1497, N110);
buf BUF1 (N1500, N1473);
not NOT1 (N1501, N1492);
buf BUF1 (N1502, N1496);
xor XOR2 (N1503, N1499, N15);
nor NOR4 (N1504, N1491, N200, N1425, N929);
nand NAND2 (N1505, N1503, N160);
nor NOR2 (N1506, N1489, N1446);
buf BUF1 (N1507, N1502);
nand NAND2 (N1508, N1505, N918);
or OR4 (N1509, N1483, N390, N1254, N452);
buf BUF1 (N1510, N1498);
or OR2 (N1511, N1500, N980);
and AND2 (N1512, N1511, N584);
xor XOR2 (N1513, N1506, N1161);
nand NAND4 (N1514, N1507, N305, N538, N847);
nand NAND2 (N1515, N1512, N939);
nor NOR4 (N1516, N1486, N681, N234, N969);
and AND4 (N1517, N1509, N130, N44, N761);
buf BUF1 (N1518, N1514);
xor XOR2 (N1519, N1513, N63);
or OR2 (N1520, N1517, N1095);
xor XOR2 (N1521, N1516, N265);
buf BUF1 (N1522, N1515);
nand NAND3 (N1523, N1504, N888, N1283);
xor XOR2 (N1524, N1518, N1367);
and AND4 (N1525, N1519, N499, N1169, N562);
nand NAND2 (N1526, N1521, N181);
and AND4 (N1527, N1524, N1516, N1020, N698);
nand NAND3 (N1528, N1520, N978, N879);
not NOT1 (N1529, N1522);
nor NOR4 (N1530, N1529, N89, N1263, N1037);
or OR3 (N1531, N1527, N70, N1111);
buf BUF1 (N1532, N1530);
and AND3 (N1533, N1531, N713, N582);
nor NOR4 (N1534, N1525, N1131, N280, N663);
xor XOR2 (N1535, N1534, N624);
buf BUF1 (N1536, N1528);
not NOT1 (N1537, N1532);
nor NOR2 (N1538, N1526, N15);
nand NAND2 (N1539, N1485, N979);
buf BUF1 (N1540, N1510);
and AND2 (N1541, N1508, N707);
not NOT1 (N1542, N1538);
buf BUF1 (N1543, N1533);
not NOT1 (N1544, N1535);
xor XOR2 (N1545, N1541, N352);
buf BUF1 (N1546, N1539);
nor NOR2 (N1547, N1542, N521);
or OR4 (N1548, N1547, N391, N101, N1012);
or OR4 (N1549, N1536, N1102, N273, N868);
nand NAND3 (N1550, N1540, N325, N177);
and AND3 (N1551, N1546, N533, N774);
or OR3 (N1552, N1550, N1390, N644);
nor NOR2 (N1553, N1543, N296);
or OR3 (N1554, N1551, N1390, N478);
nor NOR2 (N1555, N1548, N1203);
nor NOR3 (N1556, N1537, N1524, N1521);
or OR3 (N1557, N1544, N181, N294);
not NOT1 (N1558, N1553);
nor NOR4 (N1559, N1552, N109, N344, N1171);
not NOT1 (N1560, N1549);
or OR4 (N1561, N1559, N1466, N1456, N490);
xor XOR2 (N1562, N1557, N1250);
nor NOR2 (N1563, N1554, N193);
nor NOR3 (N1564, N1563, N1544, N649);
or OR4 (N1565, N1501, N90, N51, N1019);
xor XOR2 (N1566, N1556, N1160);
nor NOR3 (N1567, N1545, N290, N1230);
not NOT1 (N1568, N1567);
buf BUF1 (N1569, N1523);
buf BUF1 (N1570, N1565);
nor NOR4 (N1571, N1568, N1363, N858, N114);
nand NAND3 (N1572, N1564, N934, N518);
not NOT1 (N1573, N1560);
nor NOR3 (N1574, N1562, N984, N801);
buf BUF1 (N1575, N1571);
nor NOR3 (N1576, N1566, N1287, N422);
and AND3 (N1577, N1558, N1418, N991);
nor NOR2 (N1578, N1576, N595);
nor NOR2 (N1579, N1555, N621);
not NOT1 (N1580, N1561);
nand NAND3 (N1581, N1580, N875, N75);
not NOT1 (N1582, N1574);
and AND3 (N1583, N1572, N934, N525);
nand NAND2 (N1584, N1577, N701);
and AND2 (N1585, N1581, N1149);
xor XOR2 (N1586, N1575, N708);
not NOT1 (N1587, N1569);
nor NOR2 (N1588, N1587, N1106);
buf BUF1 (N1589, N1584);
not NOT1 (N1590, N1585);
buf BUF1 (N1591, N1583);
xor XOR2 (N1592, N1586, N1101);
not NOT1 (N1593, N1570);
nor NOR2 (N1594, N1592, N1463);
buf BUF1 (N1595, N1589);
not NOT1 (N1596, N1590);
nand NAND3 (N1597, N1593, N750, N32);
nand NAND3 (N1598, N1597, N330, N822);
nor NOR2 (N1599, N1582, N89);
or OR4 (N1600, N1595, N696, N1553, N1533);
nand NAND3 (N1601, N1598, N1419, N1354);
nor NOR3 (N1602, N1599, N249, N1320);
nor NOR3 (N1603, N1596, N136, N674);
nand NAND3 (N1604, N1591, N302, N972);
buf BUF1 (N1605, N1588);
nand NAND4 (N1606, N1600, N536, N1587, N812);
xor XOR2 (N1607, N1601, N1220);
xor XOR2 (N1608, N1604, N829);
xor XOR2 (N1609, N1603, N1310);
not NOT1 (N1610, N1594);
and AND4 (N1611, N1610, N849, N1596, N932);
and AND4 (N1612, N1611, N231, N1458, N133);
or OR3 (N1613, N1608, N1022, N681);
nand NAND2 (N1614, N1612, N1588);
not NOT1 (N1615, N1605);
not NOT1 (N1616, N1573);
or OR2 (N1617, N1578, N726);
or OR4 (N1618, N1613, N925, N1418, N363);
and AND4 (N1619, N1616, N431, N1245, N1222);
or OR2 (N1620, N1579, N710);
nand NAND2 (N1621, N1620, N1525);
buf BUF1 (N1622, N1615);
or OR4 (N1623, N1614, N310, N197, N10);
xor XOR2 (N1624, N1618, N1157);
not NOT1 (N1625, N1607);
xor XOR2 (N1626, N1625, N1409);
nor NOR4 (N1627, N1606, N1305, N874, N814);
nand NAND2 (N1628, N1621, N217);
nand NAND2 (N1629, N1627, N772);
nand NAND2 (N1630, N1609, N1434);
and AND3 (N1631, N1626, N93, N604);
or OR3 (N1632, N1602, N1150, N1106);
not NOT1 (N1633, N1619);
xor XOR2 (N1634, N1617, N842);
not NOT1 (N1635, N1623);
nand NAND3 (N1636, N1622, N1171, N1278);
not NOT1 (N1637, N1629);
or OR4 (N1638, N1631, N1231, N1544, N1556);
and AND4 (N1639, N1636, N1134, N637, N823);
nand NAND4 (N1640, N1639, N766, N1262, N361);
xor XOR2 (N1641, N1635, N1570);
buf BUF1 (N1642, N1633);
xor XOR2 (N1643, N1641, N59);
buf BUF1 (N1644, N1634);
or OR3 (N1645, N1644, N830, N1140);
or OR3 (N1646, N1645, N1101, N464);
not NOT1 (N1647, N1643);
not NOT1 (N1648, N1638);
buf BUF1 (N1649, N1630);
not NOT1 (N1650, N1640);
not NOT1 (N1651, N1642);
nor NOR4 (N1652, N1648, N90, N1334, N152);
xor XOR2 (N1653, N1624, N1390);
or OR3 (N1654, N1646, N544, N1097);
or OR3 (N1655, N1649, N1302, N560);
nand NAND4 (N1656, N1655, N952, N734, N642);
not NOT1 (N1657, N1653);
nor NOR4 (N1658, N1654, N133, N883, N1052);
nor NOR2 (N1659, N1628, N588);
not NOT1 (N1660, N1658);
xor XOR2 (N1661, N1632, N431);
not NOT1 (N1662, N1647);
nand NAND4 (N1663, N1650, N538, N1062, N756);
xor XOR2 (N1664, N1660, N938);
xor XOR2 (N1665, N1662, N797);
xor XOR2 (N1666, N1637, N757);
buf BUF1 (N1667, N1665);
xor XOR2 (N1668, N1659, N402);
xor XOR2 (N1669, N1663, N632);
nor NOR3 (N1670, N1667, N1217, N219);
and AND3 (N1671, N1657, N1277, N942);
buf BUF1 (N1672, N1668);
xor XOR2 (N1673, N1672, N1546);
nor NOR2 (N1674, N1664, N799);
buf BUF1 (N1675, N1661);
and AND3 (N1676, N1669, N204, N442);
xor XOR2 (N1677, N1671, N839);
buf BUF1 (N1678, N1651);
or OR3 (N1679, N1678, N1592, N187);
and AND2 (N1680, N1675, N439);
xor XOR2 (N1681, N1679, N1216);
nor NOR2 (N1682, N1652, N1376);
nand NAND4 (N1683, N1670, N914, N1324, N1064);
buf BUF1 (N1684, N1680);
buf BUF1 (N1685, N1681);
nor NOR3 (N1686, N1673, N514, N557);
and AND4 (N1687, N1682, N1507, N1243, N1107);
buf BUF1 (N1688, N1676);
and AND4 (N1689, N1688, N1432, N127, N105);
and AND2 (N1690, N1689, N782);
nor NOR3 (N1691, N1683, N879, N1494);
not NOT1 (N1692, N1677);
not NOT1 (N1693, N1685);
not NOT1 (N1694, N1687);
nand NAND4 (N1695, N1693, N1666, N1366, N463);
nor NOR4 (N1696, N634, N48, N232, N1182);
and AND4 (N1697, N1695, N1684, N278, N1487);
not NOT1 (N1698, N1074);
xor XOR2 (N1699, N1686, N1291);
or OR4 (N1700, N1691, N203, N1186, N566);
or OR4 (N1701, N1698, N1545, N1107, N238);
nand NAND4 (N1702, N1700, N198, N1217, N459);
buf BUF1 (N1703, N1696);
and AND3 (N1704, N1692, N102, N1294);
buf BUF1 (N1705, N1697);
nand NAND2 (N1706, N1656, N881);
xor XOR2 (N1707, N1690, N995);
and AND2 (N1708, N1703, N1051);
xor XOR2 (N1709, N1701, N1680);
nand NAND3 (N1710, N1706, N854, N34);
nand NAND3 (N1711, N1694, N798, N931);
nand NAND3 (N1712, N1702, N19, N1627);
or OR4 (N1713, N1711, N625, N509, N1680);
nand NAND2 (N1714, N1705, N1620);
not NOT1 (N1715, N1707);
xor XOR2 (N1716, N1714, N768);
or OR2 (N1717, N1708, N164);
nor NOR4 (N1718, N1704, N1171, N114, N1545);
nor NOR2 (N1719, N1712, N1428);
or OR4 (N1720, N1718, N992, N1241, N1542);
xor XOR2 (N1721, N1715, N685);
xor XOR2 (N1722, N1720, N1012);
or OR4 (N1723, N1722, N880, N1075, N902);
not NOT1 (N1724, N1709);
nand NAND4 (N1725, N1719, N867, N420, N684);
nand NAND2 (N1726, N1674, N1342);
or OR3 (N1727, N1713, N134, N1322);
and AND3 (N1728, N1699, N1242, N319);
not NOT1 (N1729, N1710);
and AND2 (N1730, N1724, N1612);
buf BUF1 (N1731, N1726);
not NOT1 (N1732, N1730);
nor NOR3 (N1733, N1732, N923, N392);
or OR2 (N1734, N1731, N588);
or OR2 (N1735, N1723, N1455);
buf BUF1 (N1736, N1728);
and AND2 (N1737, N1735, N588);
and AND4 (N1738, N1734, N542, N900, N617);
xor XOR2 (N1739, N1738, N809);
xor XOR2 (N1740, N1717, N1463);
nand NAND4 (N1741, N1736, N1149, N178, N593);
nand NAND2 (N1742, N1727, N1047);
buf BUF1 (N1743, N1721);
not NOT1 (N1744, N1729);
buf BUF1 (N1745, N1741);
and AND3 (N1746, N1744, N157, N654);
xor XOR2 (N1747, N1716, N35);
or OR2 (N1748, N1737, N168);
and AND2 (N1749, N1746, N717);
and AND3 (N1750, N1742, N664, N1703);
buf BUF1 (N1751, N1749);
xor XOR2 (N1752, N1745, N417);
nand NAND2 (N1753, N1733, N142);
nor NOR3 (N1754, N1752, N285, N912);
not NOT1 (N1755, N1739);
buf BUF1 (N1756, N1755);
buf BUF1 (N1757, N1754);
nor NOR2 (N1758, N1725, N188);
nor NOR3 (N1759, N1750, N1003, N1733);
or OR2 (N1760, N1743, N1106);
nand NAND3 (N1761, N1753, N876, N721);
xor XOR2 (N1762, N1751, N1702);
nand NAND4 (N1763, N1756, N823, N738, N938);
xor XOR2 (N1764, N1763, N571);
or OR2 (N1765, N1758, N165);
nand NAND2 (N1766, N1764, N601);
xor XOR2 (N1767, N1766, N1203);
xor XOR2 (N1768, N1759, N1532);
nand NAND3 (N1769, N1761, N1377, N1746);
xor XOR2 (N1770, N1760, N703);
xor XOR2 (N1771, N1762, N1149);
and AND2 (N1772, N1747, N1294);
not NOT1 (N1773, N1771);
buf BUF1 (N1774, N1769);
buf BUF1 (N1775, N1740);
xor XOR2 (N1776, N1768, N1426);
nand NAND2 (N1777, N1757, N191);
not NOT1 (N1778, N1777);
not NOT1 (N1779, N1774);
xor XOR2 (N1780, N1778, N1580);
not NOT1 (N1781, N1779);
or OR3 (N1782, N1780, N871, N768);
xor XOR2 (N1783, N1765, N1134);
nand NAND4 (N1784, N1781, N828, N635, N258);
nor NOR3 (N1785, N1775, N201, N889);
or OR4 (N1786, N1776, N500, N1255, N911);
or OR2 (N1787, N1770, N835);
not NOT1 (N1788, N1785);
xor XOR2 (N1789, N1772, N700);
and AND4 (N1790, N1789, N1177, N1359, N1322);
not NOT1 (N1791, N1782);
buf BUF1 (N1792, N1790);
nor NOR4 (N1793, N1748, N1568, N1005, N985);
nand NAND3 (N1794, N1788, N887, N835);
nand NAND3 (N1795, N1787, N1515, N1595);
nor NOR3 (N1796, N1767, N519, N2);
buf BUF1 (N1797, N1784);
and AND2 (N1798, N1783, N111);
xor XOR2 (N1799, N1796, N1266);
not NOT1 (N1800, N1792);
xor XOR2 (N1801, N1773, N1657);
buf BUF1 (N1802, N1799);
buf BUF1 (N1803, N1797);
nand NAND4 (N1804, N1793, N304, N762, N1063);
or OR3 (N1805, N1794, N1576, N302);
not NOT1 (N1806, N1798);
xor XOR2 (N1807, N1804, N927);
not NOT1 (N1808, N1801);
nor NOR3 (N1809, N1786, N1729, N979);
nand NAND3 (N1810, N1803, N401, N231);
and AND3 (N1811, N1791, N344, N1633);
nor NOR2 (N1812, N1807, N1331);
and AND4 (N1813, N1806, N608, N729, N941);
nor NOR4 (N1814, N1813, N567, N1115, N229);
not NOT1 (N1815, N1800);
or OR2 (N1816, N1795, N796);
or OR4 (N1817, N1810, N650, N971, N471);
nand NAND4 (N1818, N1812, N885, N382, N58);
not NOT1 (N1819, N1809);
not NOT1 (N1820, N1808);
nor NOR3 (N1821, N1805, N102, N1352);
buf BUF1 (N1822, N1814);
nor NOR3 (N1823, N1821, N324, N841);
not NOT1 (N1824, N1802);
nor NOR2 (N1825, N1815, N1603);
and AND2 (N1826, N1820, N1532);
nand NAND2 (N1827, N1822, N446);
nor NOR3 (N1828, N1811, N410, N1183);
nor NOR4 (N1829, N1824, N1264, N1006, N566);
and AND2 (N1830, N1829, N1674);
or OR3 (N1831, N1818, N1151, N1585);
buf BUF1 (N1832, N1816);
nor NOR2 (N1833, N1817, N645);
or OR2 (N1834, N1828, N449);
not NOT1 (N1835, N1826);
buf BUF1 (N1836, N1834);
nor NOR2 (N1837, N1823, N162);
or OR2 (N1838, N1827, N462);
or OR3 (N1839, N1825, N1005, N696);
or OR3 (N1840, N1838, N582, N176);
and AND4 (N1841, N1837, N526, N228, N630);
and AND4 (N1842, N1833, N1302, N55, N1436);
xor XOR2 (N1843, N1835, N815);
or OR3 (N1844, N1830, N1069, N1516);
nor NOR4 (N1845, N1831, N151, N1644, N1608);
nor NOR2 (N1846, N1842, N162);
or OR2 (N1847, N1840, N711);
or OR4 (N1848, N1844, N1376, N728, N277);
nor NOR4 (N1849, N1832, N1365, N26, N1716);
not NOT1 (N1850, N1845);
not NOT1 (N1851, N1819);
buf BUF1 (N1852, N1847);
and AND3 (N1853, N1846, N22, N1296);
nor NOR4 (N1854, N1852, N1785, N1584, N1582);
xor XOR2 (N1855, N1836, N450);
xor XOR2 (N1856, N1855, N553);
nor NOR4 (N1857, N1850, N274, N1317, N1207);
or OR2 (N1858, N1856, N1848);
xor XOR2 (N1859, N1039, N947);
buf BUF1 (N1860, N1859);
not NOT1 (N1861, N1849);
or OR2 (N1862, N1858, N1205);
nor NOR4 (N1863, N1854, N275, N1823, N1622);
not NOT1 (N1864, N1839);
nand NAND2 (N1865, N1841, N1408);
not NOT1 (N1866, N1865);
buf BUF1 (N1867, N1843);
buf BUF1 (N1868, N1867);
and AND4 (N1869, N1851, N1170, N231, N816);
and AND2 (N1870, N1864, N798);
nand NAND3 (N1871, N1862, N2, N1527);
nor NOR3 (N1872, N1869, N626, N1353);
nand NAND4 (N1873, N1853, N415, N982, N1312);
buf BUF1 (N1874, N1860);
nand NAND2 (N1875, N1857, N627);
and AND3 (N1876, N1863, N107, N11);
xor XOR2 (N1877, N1866, N1370);
not NOT1 (N1878, N1875);
and AND4 (N1879, N1861, N505, N608, N1733);
and AND3 (N1880, N1873, N711, N1716);
xor XOR2 (N1881, N1880, N1397);
or OR2 (N1882, N1868, N1356);
nand NAND2 (N1883, N1872, N834);
buf BUF1 (N1884, N1877);
xor XOR2 (N1885, N1870, N385);
or OR3 (N1886, N1879, N60, N372);
nand NAND4 (N1887, N1882, N391, N116, N562);
xor XOR2 (N1888, N1884, N1478);
nor NOR2 (N1889, N1881, N1572);
xor XOR2 (N1890, N1871, N842);
nor NOR4 (N1891, N1885, N1108, N1750, N621);
and AND3 (N1892, N1874, N1231, N742);
and AND2 (N1893, N1876, N107);
nand NAND2 (N1894, N1886, N971);
xor XOR2 (N1895, N1883, N527);
xor XOR2 (N1896, N1890, N717);
and AND2 (N1897, N1887, N684);
or OR2 (N1898, N1895, N428);
and AND3 (N1899, N1892, N812, N818);
xor XOR2 (N1900, N1888, N886);
not NOT1 (N1901, N1891);
or OR3 (N1902, N1900, N242, N1681);
or OR4 (N1903, N1898, N424, N129, N1398);
nand NAND2 (N1904, N1878, N1353);
buf BUF1 (N1905, N1901);
buf BUF1 (N1906, N1893);
buf BUF1 (N1907, N1903);
not NOT1 (N1908, N1894);
and AND4 (N1909, N1897, N807, N486, N947);
not NOT1 (N1910, N1905);
buf BUF1 (N1911, N1904);
not NOT1 (N1912, N1910);
and AND2 (N1913, N1909, N642);
nand NAND2 (N1914, N1906, N1491);
nand NAND2 (N1915, N1914, N1045);
xor XOR2 (N1916, N1912, N769);
buf BUF1 (N1917, N1907);
and AND2 (N1918, N1915, N1093);
and AND4 (N1919, N1913, N464, N1056, N777);
or OR3 (N1920, N1918, N1248, N1023);
and AND3 (N1921, N1916, N1600, N568);
not NOT1 (N1922, N1899);
buf BUF1 (N1923, N1917);
buf BUF1 (N1924, N1908);
not NOT1 (N1925, N1920);
nor NOR4 (N1926, N1902, N606, N1553, N1088);
or OR4 (N1927, N1911, N1535, N1265, N1122);
nor NOR3 (N1928, N1921, N1687, N1612);
nand NAND2 (N1929, N1927, N1090);
or OR4 (N1930, N1925, N681, N529, N976);
nor NOR4 (N1931, N1923, N717, N1063, N567);
xor XOR2 (N1932, N1919, N880);
and AND4 (N1933, N1922, N1828, N801, N149);
xor XOR2 (N1934, N1929, N1358);
nand NAND3 (N1935, N1932, N1699, N1911);
nor NOR2 (N1936, N1934, N388);
not NOT1 (N1937, N1889);
xor XOR2 (N1938, N1935, N1911);
nand NAND3 (N1939, N1924, N1390, N1554);
xor XOR2 (N1940, N1936, N1584);
buf BUF1 (N1941, N1930);
nor NOR2 (N1942, N1931, N533);
or OR4 (N1943, N1939, N1855, N1343, N534);
xor XOR2 (N1944, N1942, N731);
or OR2 (N1945, N1896, N4);
nor NOR4 (N1946, N1940, N477, N1296, N1421);
xor XOR2 (N1947, N1926, N58);
and AND4 (N1948, N1938, N711, N1342, N1141);
or OR2 (N1949, N1946, N1554);
xor XOR2 (N1950, N1933, N1898);
xor XOR2 (N1951, N1945, N844);
or OR2 (N1952, N1928, N1651);
nor NOR3 (N1953, N1950, N65, N1719);
buf BUF1 (N1954, N1949);
buf BUF1 (N1955, N1954);
xor XOR2 (N1956, N1947, N1868);
and AND4 (N1957, N1943, N1060, N153, N26);
nor NOR2 (N1958, N1944, N1368);
xor XOR2 (N1959, N1958, N728);
xor XOR2 (N1960, N1948, N372);
not NOT1 (N1961, N1951);
not NOT1 (N1962, N1953);
and AND3 (N1963, N1941, N583, N535);
and AND3 (N1964, N1957, N1256, N1108);
nor NOR3 (N1965, N1960, N1844, N38);
buf BUF1 (N1966, N1963);
nor NOR3 (N1967, N1965, N1497, N1077);
nand NAND4 (N1968, N1966, N806, N1348, N933);
nand NAND3 (N1969, N1956, N1059, N511);
buf BUF1 (N1970, N1952);
buf BUF1 (N1971, N1962);
nand NAND4 (N1972, N1964, N1680, N905, N671);
and AND2 (N1973, N1967, N593);
not NOT1 (N1974, N1971);
xor XOR2 (N1975, N1959, N83);
nand NAND2 (N1976, N1973, N1033);
xor XOR2 (N1977, N1961, N423);
and AND3 (N1978, N1974, N93, N630);
buf BUF1 (N1979, N1969);
nor NOR3 (N1980, N1977, N347, N1417);
buf BUF1 (N1981, N1980);
or OR4 (N1982, N1968, N1, N473, N1879);
and AND4 (N1983, N1981, N1760, N441, N258);
xor XOR2 (N1984, N1970, N583);
nor NOR2 (N1985, N1984, N1492);
and AND4 (N1986, N1985, N768, N1950, N241);
nor NOR4 (N1987, N1955, N1948, N815, N878);
and AND2 (N1988, N1978, N1443);
not NOT1 (N1989, N1979);
buf BUF1 (N1990, N1972);
nor NOR2 (N1991, N1976, N856);
buf BUF1 (N1992, N1991);
xor XOR2 (N1993, N1987, N630);
and AND2 (N1994, N1990, N1449);
buf BUF1 (N1995, N1988);
nor NOR2 (N1996, N1937, N806);
and AND2 (N1997, N1983, N1176);
xor XOR2 (N1998, N1996, N225);
not NOT1 (N1999, N1986);
not NOT1 (N2000, N1994);
or OR2 (N2001, N1993, N524);
buf BUF1 (N2002, N1989);
xor XOR2 (N2003, N2002, N1207);
nor NOR4 (N2004, N1995, N1283, N810, N66);
and AND4 (N2005, N1975, N1539, N980, N1939);
not NOT1 (N2006, N2005);
not NOT1 (N2007, N1998);
nand NAND4 (N2008, N1992, N883, N432, N1437);
xor XOR2 (N2009, N2000, N144);
not NOT1 (N2010, N1982);
or OR4 (N2011, N2004, N19, N1343, N165);
not NOT1 (N2012, N1997);
and AND3 (N2013, N1999, N779, N1978);
not NOT1 (N2014, N2008);
endmodule