// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N7994,N8004,N7999,N7988,N8001,N8000,N8005,N8008,N8010,N8011;

buf BUF1 (N12, N6);
or OR3 (N13, N4, N11, N10);
and AND3 (N14, N5, N10, N3);
buf BUF1 (N15, N12);
nand NAND2 (N16, N7, N12);
buf BUF1 (N17, N13);
nand NAND3 (N18, N1, N6, N3);
or OR2 (N19, N1, N14);
xor XOR2 (N20, N11, N13);
and AND4 (N21, N15, N3, N6, N12);
or OR4 (N22, N2, N20, N17, N18);
nor NOR4 (N23, N15, N21, N19, N10);
xor XOR2 (N24, N6, N16);
nor NOR3 (N25, N1, N20, N11);
or OR4 (N26, N9, N3, N3, N23);
or OR4 (N27, N24, N10, N7, N8);
buf BUF1 (N28, N8);
and AND2 (N29, N15, N20);
buf BUF1 (N30, N11);
and AND2 (N31, N20, N17);
and AND3 (N32, N23, N18, N24);
not NOT1 (N33, N14);
not NOT1 (N34, N26);
not NOT1 (N35, N27);
xor XOR2 (N36, N28, N26);
not NOT1 (N37, N22);
and AND4 (N38, N25, N6, N7, N21);
or OR4 (N39, N31, N36, N7, N17);
or OR4 (N40, N29, N6, N29, N11);
or OR2 (N41, N36, N1);
or OR3 (N42, N33, N34, N34);
and AND2 (N43, N42, N24);
buf BUF1 (N44, N10);
and AND3 (N45, N40, N18, N23);
buf BUF1 (N46, N39);
nand NAND3 (N47, N41, N44, N31);
not NOT1 (N48, N15);
nand NAND2 (N49, N32, N2);
nand NAND2 (N50, N43, N45);
or OR3 (N51, N45, N12, N17);
and AND4 (N52, N30, N21, N8, N15);
and AND2 (N53, N47, N42);
xor XOR2 (N54, N53, N46);
and AND3 (N55, N17, N26, N11);
buf BUF1 (N56, N49);
nand NAND2 (N57, N54, N45);
not NOT1 (N58, N38);
not NOT1 (N59, N50);
not NOT1 (N60, N35);
nor NOR2 (N61, N58, N12);
nand NAND4 (N62, N56, N40, N51, N36);
nand NAND2 (N63, N61, N31);
nor NOR4 (N64, N11, N21, N17, N22);
and AND3 (N65, N59, N9, N44);
nand NAND3 (N66, N62, N63, N44);
not NOT1 (N67, N54);
nand NAND2 (N68, N37, N44);
xor XOR2 (N69, N60, N54);
or OR3 (N70, N67, N37, N48);
buf BUF1 (N71, N63);
xor XOR2 (N72, N71, N48);
or OR3 (N73, N57, N25, N72);
and AND4 (N74, N66, N13, N60, N72);
nand NAND2 (N75, N58, N17);
xor XOR2 (N76, N64, N23);
and AND3 (N77, N74, N70, N63);
xor XOR2 (N78, N51, N54);
not NOT1 (N79, N73);
nor NOR2 (N80, N52, N22);
and AND3 (N81, N78, N68, N52);
not NOT1 (N82, N14);
xor XOR2 (N83, N80, N56);
xor XOR2 (N84, N82, N38);
or OR4 (N85, N65, N67, N48, N18);
xor XOR2 (N86, N69, N1);
buf BUF1 (N87, N76);
nor NOR2 (N88, N83, N14);
not NOT1 (N89, N55);
not NOT1 (N90, N89);
buf BUF1 (N91, N75);
nor NOR2 (N92, N79, N50);
nor NOR2 (N93, N87, N27);
not NOT1 (N94, N81);
and AND2 (N95, N86, N33);
nor NOR3 (N96, N88, N47, N77);
and AND4 (N97, N37, N52, N10, N54);
buf BUF1 (N98, N95);
or OR3 (N99, N98, N58, N40);
not NOT1 (N100, N91);
not NOT1 (N101, N92);
and AND4 (N102, N93, N51, N30, N71);
not NOT1 (N103, N101);
nand NAND3 (N104, N100, N61, N89);
not NOT1 (N105, N90);
not NOT1 (N106, N103);
and AND3 (N107, N105, N76, N30);
and AND2 (N108, N102, N58);
xor XOR2 (N109, N97, N42);
nor NOR3 (N110, N109, N9, N3);
nor NOR4 (N111, N106, N91, N9, N29);
and AND3 (N112, N84, N18, N38);
nand NAND3 (N113, N111, N81, N71);
buf BUF1 (N114, N112);
not NOT1 (N115, N104);
nand NAND4 (N116, N94, N31, N5, N114);
or OR2 (N117, N46, N50);
not NOT1 (N118, N99);
not NOT1 (N119, N110);
xor XOR2 (N120, N96, N96);
or OR3 (N121, N117, N53, N21);
not NOT1 (N122, N113);
or OR3 (N123, N122, N61, N9);
nand NAND4 (N124, N107, N67, N100, N94);
nor NOR3 (N125, N118, N93, N60);
not NOT1 (N126, N124);
and AND2 (N127, N115, N67);
buf BUF1 (N128, N116);
nand NAND2 (N129, N119, N114);
buf BUF1 (N130, N108);
or OR3 (N131, N128, N21, N88);
xor XOR2 (N132, N127, N43);
and AND4 (N133, N123, N118, N90, N122);
not NOT1 (N134, N121);
xor XOR2 (N135, N120, N98);
nand NAND4 (N136, N134, N94, N38, N57);
or OR4 (N137, N132, N68, N45, N76);
xor XOR2 (N138, N130, N90);
or OR4 (N139, N126, N89, N32, N129);
or OR2 (N140, N90, N40);
nor NOR2 (N141, N135, N131);
not NOT1 (N142, N85);
and AND2 (N143, N12, N56);
buf BUF1 (N144, N141);
xor XOR2 (N145, N140, N2);
buf BUF1 (N146, N139);
nor NOR2 (N147, N144, N2);
or OR2 (N148, N136, N86);
buf BUF1 (N149, N148);
not NOT1 (N150, N147);
nand NAND2 (N151, N125, N124);
nor NOR2 (N152, N138, N88);
buf BUF1 (N153, N137);
and AND2 (N154, N143, N64);
and AND2 (N155, N152, N140);
or OR4 (N156, N145, N132, N9, N16);
xor XOR2 (N157, N156, N34);
or OR3 (N158, N155, N7, N130);
and AND2 (N159, N154, N29);
nand NAND4 (N160, N150, N136, N131, N148);
or OR4 (N161, N146, N15, N83, N13);
xor XOR2 (N162, N158, N56);
xor XOR2 (N163, N160, N31);
and AND4 (N164, N163, N26, N133, N72);
not NOT1 (N165, N23);
nand NAND4 (N166, N149, N101, N46, N114);
not NOT1 (N167, N164);
or OR2 (N168, N161, N113);
xor XOR2 (N169, N142, N93);
nand NAND3 (N170, N169, N124, N154);
and AND2 (N171, N162, N135);
nor NOR4 (N172, N153, N156, N149, N43);
buf BUF1 (N173, N159);
and AND3 (N174, N167, N17, N116);
nand NAND3 (N175, N165, N6, N147);
and AND4 (N176, N174, N105, N172, N136);
nor NOR2 (N177, N125, N142);
not NOT1 (N178, N157);
nor NOR3 (N179, N170, N151, N149);
buf BUF1 (N180, N26);
xor XOR2 (N181, N168, N146);
and AND3 (N182, N179, N172, N140);
or OR3 (N183, N166, N160, N11);
not NOT1 (N184, N171);
xor XOR2 (N185, N181, N32);
xor XOR2 (N186, N177, N164);
nor NOR4 (N187, N186, N94, N93, N138);
not NOT1 (N188, N176);
xor XOR2 (N189, N182, N29);
xor XOR2 (N190, N189, N132);
nor NOR3 (N191, N188, N183, N65);
nor NOR4 (N192, N76, N55, N15, N82);
buf BUF1 (N193, N175);
xor XOR2 (N194, N191, N55);
nor NOR4 (N195, N190, N82, N123, N38);
xor XOR2 (N196, N193, N135);
nand NAND4 (N197, N192, N169, N60, N12);
nor NOR3 (N198, N195, N75, N58);
and AND2 (N199, N178, N31);
nand NAND3 (N200, N173, N44, N46);
nor NOR3 (N201, N199, N95, N81);
and AND2 (N202, N197, N17);
xor XOR2 (N203, N202, N83);
and AND3 (N204, N185, N34, N30);
or OR3 (N205, N198, N93, N112);
nor NOR4 (N206, N194, N51, N9, N114);
xor XOR2 (N207, N201, N107);
not NOT1 (N208, N200);
or OR4 (N209, N203, N133, N40, N57);
not NOT1 (N210, N207);
xor XOR2 (N211, N204, N102);
xor XOR2 (N212, N180, N101);
and AND2 (N213, N205, N180);
or OR2 (N214, N209, N150);
nor NOR2 (N215, N211, N150);
buf BUF1 (N216, N184);
nor NOR4 (N217, N216, N210, N37, N21);
buf BUF1 (N218, N179);
xor XOR2 (N219, N215, N209);
not NOT1 (N220, N208);
buf BUF1 (N221, N187);
buf BUF1 (N222, N219);
nand NAND2 (N223, N221, N14);
nor NOR3 (N224, N218, N21, N160);
not NOT1 (N225, N196);
nand NAND4 (N226, N225, N130, N92, N113);
and AND3 (N227, N226, N206, N126);
nor NOR4 (N228, N202, N168, N8, N177);
buf BUF1 (N229, N223);
xor XOR2 (N230, N217, N224);
xor XOR2 (N231, N165, N118);
not NOT1 (N232, N212);
nand NAND4 (N233, N220, N30, N136, N31);
nor NOR2 (N234, N231, N203);
xor XOR2 (N235, N222, N183);
nor NOR3 (N236, N230, N23, N201);
not NOT1 (N237, N236);
or OR2 (N238, N228, N52);
nor NOR2 (N239, N232, N11);
nor NOR2 (N240, N229, N238);
xor XOR2 (N241, N61, N13);
xor XOR2 (N242, N233, N185);
nor NOR3 (N243, N214, N137, N112);
nor NOR3 (N244, N234, N56, N125);
buf BUF1 (N245, N237);
nand NAND2 (N246, N242, N78);
or OR2 (N247, N241, N56);
or OR2 (N248, N243, N226);
xor XOR2 (N249, N235, N214);
buf BUF1 (N250, N246);
and AND3 (N251, N227, N74, N158);
xor XOR2 (N252, N244, N195);
not NOT1 (N253, N247);
buf BUF1 (N254, N251);
nand NAND2 (N255, N245, N168);
nor NOR4 (N256, N252, N201, N16, N52);
or OR4 (N257, N250, N194, N71, N226);
xor XOR2 (N258, N255, N138);
or OR4 (N259, N258, N186, N216, N204);
xor XOR2 (N260, N254, N61);
xor XOR2 (N261, N239, N13);
not NOT1 (N262, N240);
xor XOR2 (N263, N248, N35);
or OR4 (N264, N256, N235, N132, N215);
xor XOR2 (N265, N213, N161);
nand NAND4 (N266, N253, N6, N13, N97);
buf BUF1 (N267, N261);
xor XOR2 (N268, N263, N190);
not NOT1 (N269, N264);
nand NAND2 (N270, N257, N172);
not NOT1 (N271, N267);
or OR2 (N272, N266, N171);
buf BUF1 (N273, N272);
nand NAND4 (N274, N249, N96, N66, N48);
nor NOR3 (N275, N262, N200, N61);
buf BUF1 (N276, N268);
or OR2 (N277, N273, N204);
nor NOR2 (N278, N271, N250);
not NOT1 (N279, N260);
nand NAND2 (N280, N277, N123);
or OR4 (N281, N274, N33, N233, N163);
nand NAND2 (N282, N280, N79);
nor NOR3 (N283, N278, N105, N208);
and AND4 (N284, N279, N223, N201, N121);
nand NAND3 (N285, N281, N229, N90);
or OR4 (N286, N282, N50, N199, N164);
buf BUF1 (N287, N269);
or OR2 (N288, N283, N197);
nand NAND4 (N289, N286, N285, N213, N25);
nor NOR3 (N290, N79, N199, N76);
or OR3 (N291, N275, N3, N141);
buf BUF1 (N292, N290);
and AND3 (N293, N259, N288, N201);
or OR3 (N294, N12, N24, N174);
nand NAND2 (N295, N270, N143);
nand NAND4 (N296, N294, N60, N156, N75);
or OR4 (N297, N284, N16, N208, N118);
not NOT1 (N298, N293);
and AND2 (N299, N276, N89);
and AND3 (N300, N295, N24, N129);
nand NAND2 (N301, N265, N119);
and AND2 (N302, N298, N61);
buf BUF1 (N303, N302);
buf BUF1 (N304, N300);
nor NOR4 (N305, N289, N260, N59, N260);
not NOT1 (N306, N299);
nor NOR2 (N307, N287, N86);
not NOT1 (N308, N305);
and AND4 (N309, N301, N227, N259, N14);
not NOT1 (N310, N304);
nor NOR4 (N311, N292, N172, N90, N234);
nor NOR3 (N312, N303, N5, N138);
xor XOR2 (N313, N309, N152);
or OR4 (N314, N312, N79, N96, N305);
nand NAND3 (N315, N314, N101, N244);
and AND2 (N316, N310, N227);
not NOT1 (N317, N307);
nor NOR4 (N318, N306, N284, N215, N92);
buf BUF1 (N319, N291);
buf BUF1 (N320, N319);
buf BUF1 (N321, N316);
not NOT1 (N322, N317);
xor XOR2 (N323, N313, N252);
and AND4 (N324, N321, N275, N173, N136);
buf BUF1 (N325, N311);
xor XOR2 (N326, N324, N207);
not NOT1 (N327, N326);
xor XOR2 (N328, N315, N316);
nand NAND4 (N329, N296, N7, N215, N127);
nor NOR4 (N330, N328, N329, N319, N30);
nor NOR3 (N331, N257, N57, N251);
xor XOR2 (N332, N320, N42);
and AND3 (N333, N331, N68, N187);
buf BUF1 (N334, N330);
nand NAND2 (N335, N327, N306);
not NOT1 (N336, N308);
not NOT1 (N337, N325);
not NOT1 (N338, N297);
xor XOR2 (N339, N334, N202);
buf BUF1 (N340, N335);
or OR3 (N341, N340, N214, N74);
and AND2 (N342, N341, N81);
not NOT1 (N343, N332);
not NOT1 (N344, N337);
or OR3 (N345, N344, N266, N163);
and AND3 (N346, N342, N202, N42);
nor NOR4 (N347, N322, N159, N318, N5);
not NOT1 (N348, N139);
not NOT1 (N349, N338);
nor NOR3 (N350, N343, N165, N139);
nand NAND2 (N351, N345, N95);
and AND4 (N352, N349, N248, N7, N329);
nand NAND3 (N353, N348, N161, N35);
or OR4 (N354, N353, N289, N21, N26);
not NOT1 (N355, N323);
and AND3 (N356, N333, N89, N26);
xor XOR2 (N357, N352, N254);
xor XOR2 (N358, N356, N302);
nor NOR2 (N359, N336, N154);
nor NOR4 (N360, N351, N249, N233, N303);
and AND4 (N361, N354, N306, N156, N45);
buf BUF1 (N362, N350);
buf BUF1 (N363, N346);
and AND3 (N364, N359, N200, N113);
nor NOR3 (N365, N357, N23, N84);
not NOT1 (N366, N361);
not NOT1 (N367, N360);
and AND2 (N368, N367, N284);
not NOT1 (N369, N339);
or OR4 (N370, N369, N321, N136, N131);
buf BUF1 (N371, N355);
nor NOR2 (N372, N363, N126);
xor XOR2 (N373, N368, N241);
xor XOR2 (N374, N373, N358);
and AND3 (N375, N293, N366, N356);
not NOT1 (N376, N36);
or OR3 (N377, N347, N120, N344);
buf BUF1 (N378, N376);
and AND4 (N379, N374, N373, N247, N345);
and AND3 (N380, N370, N105, N93);
not NOT1 (N381, N362);
not NOT1 (N382, N377);
nand NAND3 (N383, N380, N68, N79);
nor NOR3 (N384, N365, N208, N265);
nand NAND3 (N385, N378, N247, N239);
xor XOR2 (N386, N382, N318);
or OR2 (N387, N385, N374);
buf BUF1 (N388, N372);
nor NOR4 (N389, N381, N99, N157, N188);
or OR2 (N390, N389, N355);
buf BUF1 (N391, N383);
or OR3 (N392, N388, N27, N111);
not NOT1 (N393, N371);
xor XOR2 (N394, N379, N3);
not NOT1 (N395, N394);
buf BUF1 (N396, N390);
not NOT1 (N397, N393);
or OR3 (N398, N397, N393, N163);
or OR4 (N399, N391, N98, N109, N115);
or OR4 (N400, N395, N190, N51, N87);
and AND3 (N401, N392, N364, N143);
not NOT1 (N402, N11);
not NOT1 (N403, N387);
nor NOR2 (N404, N400, N322);
buf BUF1 (N405, N404);
not NOT1 (N406, N396);
and AND3 (N407, N402, N205, N134);
nand NAND4 (N408, N406, N111, N98, N158);
and AND3 (N409, N398, N180, N198);
nand NAND4 (N410, N407, N94, N115, N152);
not NOT1 (N411, N403);
nand NAND3 (N412, N410, N5, N283);
or OR3 (N413, N412, N410, N264);
nor NOR4 (N414, N413, N196, N322, N397);
buf BUF1 (N415, N409);
buf BUF1 (N416, N408);
xor XOR2 (N417, N375, N382);
and AND3 (N418, N405, N42, N341);
or OR4 (N419, N401, N131, N34, N282);
or OR3 (N420, N417, N311, N1);
not NOT1 (N421, N399);
and AND3 (N422, N411, N18, N232);
and AND3 (N423, N414, N373, N95);
nor NOR2 (N424, N420, N36);
not NOT1 (N425, N384);
buf BUF1 (N426, N422);
nor NOR3 (N427, N419, N348, N264);
nand NAND2 (N428, N425, N252);
buf BUF1 (N429, N424);
and AND2 (N430, N427, N328);
not NOT1 (N431, N415);
buf BUF1 (N432, N429);
nand NAND3 (N433, N426, N161, N7);
and AND2 (N434, N428, N103);
not NOT1 (N435, N423);
xor XOR2 (N436, N432, N278);
or OR3 (N437, N431, N384, N41);
nor NOR2 (N438, N421, N347);
or OR3 (N439, N438, N395, N314);
xor XOR2 (N440, N433, N132);
not NOT1 (N441, N435);
and AND4 (N442, N434, N387, N185, N397);
and AND4 (N443, N442, N85, N66, N332);
buf BUF1 (N444, N443);
and AND2 (N445, N440, N45);
nand NAND4 (N446, N416, N117, N262, N287);
nor NOR4 (N447, N436, N84, N74, N419);
nand NAND3 (N448, N418, N380, N119);
nor NOR3 (N449, N441, N11, N25);
or OR2 (N450, N430, N39);
nand NAND2 (N451, N444, N345);
nand NAND4 (N452, N450, N327, N215, N367);
nand NAND4 (N453, N448, N285, N402, N163);
buf BUF1 (N454, N445);
not NOT1 (N455, N449);
xor XOR2 (N456, N446, N448);
nor NOR4 (N457, N386, N138, N336, N350);
buf BUF1 (N458, N451);
and AND2 (N459, N439, N379);
nor NOR2 (N460, N452, N49);
nand NAND2 (N461, N447, N362);
xor XOR2 (N462, N461, N62);
not NOT1 (N463, N453);
nor NOR3 (N464, N459, N64, N8);
and AND2 (N465, N458, N224);
and AND3 (N466, N463, N218, N146);
xor XOR2 (N467, N455, N431);
nor NOR4 (N468, N456, N76, N80, N115);
buf BUF1 (N469, N454);
not NOT1 (N470, N437);
xor XOR2 (N471, N467, N45);
xor XOR2 (N472, N465, N37);
buf BUF1 (N473, N470);
nand NAND2 (N474, N472, N190);
and AND3 (N475, N473, N66, N185);
not NOT1 (N476, N475);
and AND4 (N477, N462, N174, N138, N259);
buf BUF1 (N478, N477);
and AND3 (N479, N469, N248, N44);
and AND3 (N480, N466, N42, N9);
nand NAND3 (N481, N478, N31, N340);
nand NAND3 (N482, N480, N442, N473);
and AND2 (N483, N468, N188);
buf BUF1 (N484, N474);
nand NAND2 (N485, N457, N77);
or OR4 (N486, N464, N143, N239, N227);
nor NOR2 (N487, N485, N382);
or OR3 (N488, N481, N99, N173);
not NOT1 (N489, N483);
not NOT1 (N490, N460);
and AND3 (N491, N487, N394, N203);
or OR4 (N492, N482, N313, N361, N342);
and AND2 (N493, N489, N173);
not NOT1 (N494, N492);
nor NOR4 (N495, N486, N87, N260, N124);
not NOT1 (N496, N490);
and AND3 (N497, N476, N167, N435);
buf BUF1 (N498, N496);
not NOT1 (N499, N479);
nor NOR3 (N500, N488, N91, N429);
buf BUF1 (N501, N500);
or OR3 (N502, N484, N322, N336);
not NOT1 (N503, N494);
nand NAND2 (N504, N491, N54);
or OR4 (N505, N493, N98, N88, N44);
not NOT1 (N506, N498);
buf BUF1 (N507, N501);
buf BUF1 (N508, N502);
and AND2 (N509, N499, N68);
nor NOR2 (N510, N471, N323);
not NOT1 (N511, N504);
or OR2 (N512, N505, N394);
or OR3 (N513, N509, N244, N213);
not NOT1 (N514, N511);
nand NAND2 (N515, N503, N38);
nor NOR4 (N516, N514, N151, N273, N406);
nand NAND3 (N517, N516, N237, N472);
buf BUF1 (N518, N497);
buf BUF1 (N519, N508);
and AND4 (N520, N513, N438, N199, N388);
xor XOR2 (N521, N520, N349);
not NOT1 (N522, N507);
and AND2 (N523, N519, N136);
xor XOR2 (N524, N510, N345);
or OR4 (N525, N521, N497, N282, N211);
nand NAND2 (N526, N517, N151);
xor XOR2 (N527, N515, N226);
not NOT1 (N528, N522);
nor NOR2 (N529, N506, N442);
and AND2 (N530, N527, N128);
xor XOR2 (N531, N525, N53);
and AND2 (N532, N530, N374);
or OR4 (N533, N531, N157, N3, N16);
buf BUF1 (N534, N495);
or OR4 (N535, N523, N357, N272, N84);
nand NAND2 (N536, N524, N63);
buf BUF1 (N537, N533);
buf BUF1 (N538, N535);
xor XOR2 (N539, N538, N518);
and AND3 (N540, N49, N73, N4);
and AND2 (N541, N539, N119);
buf BUF1 (N542, N540);
or OR3 (N543, N534, N451, N521);
or OR4 (N544, N529, N346, N346, N165);
xor XOR2 (N545, N528, N410);
or OR4 (N546, N536, N267, N195, N253);
and AND3 (N547, N544, N128, N241);
not NOT1 (N548, N543);
or OR3 (N549, N541, N536, N482);
or OR3 (N550, N547, N179, N389);
xor XOR2 (N551, N545, N415);
nand NAND3 (N552, N537, N52, N66);
or OR3 (N553, N532, N88, N506);
buf BUF1 (N554, N550);
nor NOR3 (N555, N554, N278, N227);
buf BUF1 (N556, N555);
nand NAND3 (N557, N552, N412, N147);
and AND4 (N558, N542, N256, N319, N325);
xor XOR2 (N559, N557, N259);
buf BUF1 (N560, N526);
nand NAND3 (N561, N559, N474, N519);
nand NAND4 (N562, N551, N530, N204, N363);
and AND3 (N563, N562, N468, N198);
buf BUF1 (N564, N561);
nand NAND2 (N565, N512, N271);
nand NAND2 (N566, N553, N123);
not NOT1 (N567, N556);
nor NOR4 (N568, N560, N316, N91, N258);
or OR3 (N569, N567, N368, N350);
not NOT1 (N570, N568);
not NOT1 (N571, N563);
or OR4 (N572, N558, N23, N34, N35);
xor XOR2 (N573, N564, N306);
nor NOR3 (N574, N548, N467, N8);
buf BUF1 (N575, N571);
nand NAND4 (N576, N549, N144, N291, N389);
xor XOR2 (N577, N576, N223);
and AND2 (N578, N572, N155);
and AND2 (N579, N575, N345);
xor XOR2 (N580, N569, N504);
xor XOR2 (N581, N580, N552);
nor NOR2 (N582, N574, N298);
buf BUF1 (N583, N577);
or OR2 (N584, N582, N497);
nor NOR4 (N585, N565, N308, N42, N254);
nor NOR3 (N586, N581, N17, N354);
or OR3 (N587, N570, N298, N491);
buf BUF1 (N588, N585);
or OR2 (N589, N583, N581);
not NOT1 (N590, N587);
buf BUF1 (N591, N546);
xor XOR2 (N592, N584, N20);
not NOT1 (N593, N592);
xor XOR2 (N594, N578, N96);
xor XOR2 (N595, N588, N302);
nor NOR4 (N596, N586, N389, N46, N122);
nand NAND2 (N597, N590, N115);
and AND2 (N598, N589, N469);
xor XOR2 (N599, N594, N351);
not NOT1 (N600, N599);
xor XOR2 (N601, N600, N541);
xor XOR2 (N602, N591, N591);
nor NOR2 (N603, N596, N54);
nand NAND2 (N604, N573, N438);
nand NAND4 (N605, N602, N5, N200, N352);
not NOT1 (N606, N579);
nor NOR4 (N607, N605, N23, N519, N313);
or OR4 (N608, N597, N130, N497, N33);
and AND2 (N609, N604, N532);
xor XOR2 (N610, N607, N188);
or OR2 (N611, N603, N125);
nor NOR2 (N612, N610, N386);
and AND2 (N613, N601, N435);
xor XOR2 (N614, N593, N542);
nand NAND4 (N615, N611, N37, N142, N265);
xor XOR2 (N616, N608, N142);
or OR4 (N617, N614, N351, N221, N262);
nor NOR4 (N618, N613, N465, N50, N565);
not NOT1 (N619, N566);
buf BUF1 (N620, N615);
xor XOR2 (N621, N619, N379);
xor XOR2 (N622, N609, N178);
buf BUF1 (N623, N618);
nor NOR3 (N624, N595, N141, N12);
xor XOR2 (N625, N617, N571);
nand NAND3 (N626, N622, N95, N338);
or OR4 (N627, N598, N584, N226, N131);
and AND3 (N628, N625, N75, N376);
and AND4 (N629, N626, N117, N370, N619);
xor XOR2 (N630, N621, N139);
buf BUF1 (N631, N620);
or OR4 (N632, N606, N59, N10, N394);
not NOT1 (N633, N629);
nor NOR4 (N634, N623, N300, N1, N498);
or OR3 (N635, N634, N362, N396);
nand NAND3 (N636, N632, N393, N547);
nor NOR4 (N637, N635, N591, N50, N307);
not NOT1 (N638, N631);
and AND2 (N639, N638, N130);
not NOT1 (N640, N630);
nor NOR3 (N641, N624, N311, N517);
nor NOR3 (N642, N627, N263, N336);
xor XOR2 (N643, N637, N410);
buf BUF1 (N644, N640);
xor XOR2 (N645, N639, N30);
nand NAND4 (N646, N641, N74, N340, N251);
buf BUF1 (N647, N612);
nand NAND2 (N648, N644, N51);
nand NAND4 (N649, N616, N260, N445, N460);
not NOT1 (N650, N633);
nor NOR3 (N651, N628, N413, N164);
and AND4 (N652, N636, N322, N567, N426);
nor NOR2 (N653, N651, N318);
or OR2 (N654, N645, N356);
buf BUF1 (N655, N647);
xor XOR2 (N656, N654, N15);
buf BUF1 (N657, N656);
nand NAND2 (N658, N657, N558);
nand NAND3 (N659, N650, N171, N100);
buf BUF1 (N660, N649);
buf BUF1 (N661, N643);
nor NOR3 (N662, N648, N526, N295);
nand NAND2 (N663, N661, N352);
nor NOR2 (N664, N658, N60);
nor NOR4 (N665, N664, N554, N289, N181);
nand NAND3 (N666, N660, N108, N571);
nand NAND2 (N667, N659, N609);
not NOT1 (N668, N666);
xor XOR2 (N669, N665, N615);
nand NAND2 (N670, N668, N14);
or OR4 (N671, N652, N371, N68, N659);
xor XOR2 (N672, N653, N361);
or OR3 (N673, N662, N464, N519);
nor NOR4 (N674, N671, N518, N402, N414);
buf BUF1 (N675, N670);
and AND4 (N676, N672, N209, N331, N286);
buf BUF1 (N677, N673);
xor XOR2 (N678, N663, N604);
and AND4 (N679, N678, N227, N121, N569);
and AND4 (N680, N667, N104, N114, N635);
nor NOR2 (N681, N674, N318);
or OR2 (N682, N675, N95);
not NOT1 (N683, N676);
or OR2 (N684, N682, N235);
nand NAND3 (N685, N642, N22, N292);
nor NOR3 (N686, N684, N35, N353);
nand NAND4 (N687, N680, N473, N79, N295);
nor NOR3 (N688, N685, N174, N68);
and AND3 (N689, N683, N70, N221);
and AND3 (N690, N646, N447, N220);
not NOT1 (N691, N689);
not NOT1 (N692, N655);
xor XOR2 (N693, N687, N88);
not NOT1 (N694, N679);
not NOT1 (N695, N690);
nand NAND2 (N696, N688, N42);
buf BUF1 (N697, N694);
nor NOR3 (N698, N691, N89, N244);
buf BUF1 (N699, N686);
nor NOR3 (N700, N697, N315, N60);
xor XOR2 (N701, N692, N185);
buf BUF1 (N702, N696);
nand NAND2 (N703, N698, N139);
nor NOR2 (N704, N695, N314);
not NOT1 (N705, N693);
nand NAND3 (N706, N701, N517, N442);
not NOT1 (N707, N677);
and AND3 (N708, N699, N381, N427);
and AND3 (N709, N669, N413, N343);
or OR4 (N710, N681, N652, N502, N407);
not NOT1 (N711, N708);
and AND4 (N712, N709, N40, N570, N305);
nor NOR4 (N713, N711, N200, N366, N183);
nand NAND4 (N714, N712, N91, N646, N202);
or OR2 (N715, N713, N267);
not NOT1 (N716, N704);
and AND3 (N717, N714, N245, N614);
not NOT1 (N718, N705);
nand NAND2 (N719, N710, N703);
not NOT1 (N720, N319);
buf BUF1 (N721, N700);
or OR3 (N722, N702, N147, N560);
and AND4 (N723, N715, N266, N393, N542);
buf BUF1 (N724, N721);
and AND3 (N725, N717, N70, N662);
and AND4 (N726, N725, N273, N615, N85);
nand NAND3 (N727, N726, N93, N120);
or OR2 (N728, N723, N598);
nor NOR4 (N729, N724, N88, N132, N229);
not NOT1 (N730, N706);
not NOT1 (N731, N720);
or OR4 (N732, N716, N423, N288, N100);
not NOT1 (N733, N731);
buf BUF1 (N734, N722);
nand NAND4 (N735, N728, N133, N411, N188);
buf BUF1 (N736, N733);
and AND2 (N737, N727, N202);
or OR2 (N738, N737, N356);
not NOT1 (N739, N707);
and AND2 (N740, N719, N55);
buf BUF1 (N741, N732);
buf BUF1 (N742, N718);
nand NAND2 (N743, N739, N375);
and AND3 (N744, N741, N533, N325);
not NOT1 (N745, N736);
or OR4 (N746, N743, N687, N308, N185);
not NOT1 (N747, N744);
buf BUF1 (N748, N735);
nor NOR3 (N749, N745, N515, N509);
not NOT1 (N750, N748);
buf BUF1 (N751, N747);
not NOT1 (N752, N729);
not NOT1 (N753, N742);
not NOT1 (N754, N746);
nor NOR2 (N755, N752, N479);
not NOT1 (N756, N750);
nor NOR2 (N757, N734, N696);
xor XOR2 (N758, N756, N209);
nand NAND2 (N759, N758, N240);
and AND2 (N760, N757, N183);
nor NOR2 (N761, N760, N492);
and AND2 (N762, N754, N418);
and AND4 (N763, N755, N178, N624, N417);
not NOT1 (N764, N730);
not NOT1 (N765, N759);
and AND4 (N766, N763, N430, N176, N348);
xor XOR2 (N767, N766, N763);
nor NOR3 (N768, N749, N438, N655);
and AND3 (N769, N764, N665, N234);
or OR3 (N770, N765, N559, N173);
xor XOR2 (N771, N769, N624);
not NOT1 (N772, N738);
buf BUF1 (N773, N772);
xor XOR2 (N774, N753, N747);
buf BUF1 (N775, N774);
buf BUF1 (N776, N740);
nor NOR4 (N777, N762, N423, N744, N26);
buf BUF1 (N778, N761);
nor NOR2 (N779, N773, N775);
nor NOR3 (N780, N27, N45, N460);
and AND3 (N781, N778, N204, N136);
nand NAND3 (N782, N777, N189, N753);
not NOT1 (N783, N779);
buf BUF1 (N784, N780);
or OR3 (N785, N770, N276, N653);
nor NOR4 (N786, N784, N468, N356, N192);
xor XOR2 (N787, N781, N91);
or OR4 (N788, N776, N771, N154, N592);
xor XOR2 (N789, N26, N172);
buf BUF1 (N790, N788);
buf BUF1 (N791, N782);
not NOT1 (N792, N767);
not NOT1 (N793, N792);
or OR3 (N794, N751, N89, N295);
or OR2 (N795, N793, N778);
not NOT1 (N796, N785);
xor XOR2 (N797, N768, N199);
or OR3 (N798, N786, N242, N257);
nor NOR3 (N799, N796, N646, N771);
nor NOR2 (N800, N799, N110);
nand NAND4 (N801, N795, N630, N96, N636);
buf BUF1 (N802, N798);
buf BUF1 (N803, N797);
or OR3 (N804, N789, N444, N44);
or OR4 (N805, N801, N616, N677, N678);
or OR2 (N806, N804, N717);
nand NAND3 (N807, N803, N163, N759);
xor XOR2 (N808, N802, N655);
nand NAND4 (N809, N787, N497, N581, N329);
and AND2 (N810, N807, N700);
buf BUF1 (N811, N808);
not NOT1 (N812, N783);
xor XOR2 (N813, N805, N531);
or OR4 (N814, N813, N371, N666, N168);
buf BUF1 (N815, N809);
nand NAND2 (N816, N806, N413);
and AND2 (N817, N816, N117);
buf BUF1 (N818, N817);
not NOT1 (N819, N794);
buf BUF1 (N820, N819);
or OR2 (N821, N820, N487);
and AND3 (N822, N791, N246, N251);
nand NAND4 (N823, N814, N287, N797, N232);
buf BUF1 (N824, N823);
nand NAND2 (N825, N810, N130);
or OR3 (N826, N790, N673, N447);
buf BUF1 (N827, N821);
nor NOR3 (N828, N822, N437, N47);
and AND3 (N829, N818, N271, N51);
nor NOR4 (N830, N828, N515, N671, N224);
or OR2 (N831, N800, N546);
nor NOR2 (N832, N829, N526);
not NOT1 (N833, N825);
and AND2 (N834, N815, N578);
nor NOR4 (N835, N824, N562, N820, N526);
nand NAND3 (N836, N835, N770, N345);
nand NAND2 (N837, N836, N773);
nor NOR3 (N838, N830, N604, N212);
nor NOR4 (N839, N837, N472, N424, N141);
nand NAND3 (N840, N811, N416, N283);
or OR2 (N841, N839, N115);
or OR4 (N842, N838, N806, N766, N516);
nor NOR2 (N843, N831, N185);
nor NOR2 (N844, N826, N499);
nand NAND3 (N845, N812, N17, N606);
xor XOR2 (N846, N834, N305);
buf BUF1 (N847, N845);
nor NOR2 (N848, N846, N181);
and AND4 (N849, N844, N772, N551, N18);
xor XOR2 (N850, N842, N50);
and AND4 (N851, N850, N54, N518, N230);
and AND3 (N852, N827, N821, N31);
nand NAND3 (N853, N851, N477, N525);
nor NOR4 (N854, N848, N736, N277, N1);
not NOT1 (N855, N832);
nor NOR3 (N856, N852, N844, N761);
not NOT1 (N857, N849);
and AND2 (N858, N833, N443);
and AND4 (N859, N843, N831, N339, N411);
buf BUF1 (N860, N853);
nand NAND2 (N861, N854, N38);
buf BUF1 (N862, N840);
nand NAND2 (N863, N847, N596);
nand NAND3 (N864, N857, N49, N287);
or OR2 (N865, N858, N722);
or OR3 (N866, N860, N763, N114);
nand NAND4 (N867, N863, N197, N825, N190);
not NOT1 (N868, N855);
or OR3 (N869, N867, N573, N20);
not NOT1 (N870, N864);
and AND4 (N871, N868, N184, N216, N460);
buf BUF1 (N872, N870);
or OR2 (N873, N869, N302);
xor XOR2 (N874, N866, N762);
and AND2 (N875, N874, N708);
buf BUF1 (N876, N856);
buf BUF1 (N877, N859);
nand NAND2 (N878, N876, N417);
not NOT1 (N879, N841);
nand NAND3 (N880, N879, N616, N453);
nand NAND2 (N881, N871, N660);
nand NAND2 (N882, N880, N428);
and AND3 (N883, N877, N783, N293);
buf BUF1 (N884, N861);
nor NOR4 (N885, N882, N802, N390, N313);
or OR2 (N886, N865, N867);
xor XOR2 (N887, N862, N879);
nand NAND2 (N888, N878, N173);
nor NOR3 (N889, N884, N603, N44);
not NOT1 (N890, N875);
not NOT1 (N891, N885);
nor NOR3 (N892, N888, N344, N351);
or OR2 (N893, N872, N805);
and AND4 (N894, N883, N461, N685, N254);
buf BUF1 (N895, N887);
or OR4 (N896, N881, N884, N52, N492);
not NOT1 (N897, N892);
xor XOR2 (N898, N889, N560);
nand NAND4 (N899, N873, N721, N127, N842);
or OR4 (N900, N890, N600, N48, N194);
nor NOR3 (N901, N894, N307, N30);
nand NAND3 (N902, N897, N834, N586);
buf BUF1 (N903, N900);
buf BUF1 (N904, N896);
and AND4 (N905, N886, N555, N703, N724);
xor XOR2 (N906, N901, N472);
buf BUF1 (N907, N893);
and AND4 (N908, N899, N743, N61, N653);
or OR2 (N909, N905, N747);
nand NAND4 (N910, N895, N164, N504, N384);
xor XOR2 (N911, N906, N19);
nor NOR3 (N912, N907, N374, N112);
or OR3 (N913, N911, N162, N35);
not NOT1 (N914, N903);
and AND4 (N915, N898, N67, N412, N736);
not NOT1 (N916, N910);
and AND4 (N917, N908, N96, N164, N284);
buf BUF1 (N918, N916);
nor NOR3 (N919, N914, N791, N541);
and AND4 (N920, N918, N418, N405, N77);
nand NAND4 (N921, N913, N244, N394, N692);
buf BUF1 (N922, N917);
nand NAND3 (N923, N912, N677, N354);
or OR3 (N924, N904, N447, N356);
nand NAND4 (N925, N923, N783, N507, N572);
and AND4 (N926, N915, N529, N666, N704);
nand NAND4 (N927, N920, N68, N181, N89);
xor XOR2 (N928, N926, N267);
not NOT1 (N929, N925);
buf BUF1 (N930, N928);
and AND2 (N931, N921, N594);
buf BUF1 (N932, N922);
or OR2 (N933, N931, N724);
or OR2 (N934, N909, N405);
xor XOR2 (N935, N932, N266);
xor XOR2 (N936, N934, N912);
xor XOR2 (N937, N933, N839);
not NOT1 (N938, N936);
buf BUF1 (N939, N919);
buf BUF1 (N940, N924);
or OR3 (N941, N937, N183, N759);
or OR2 (N942, N940, N26);
nand NAND3 (N943, N935, N457, N741);
buf BUF1 (N944, N891);
nand NAND4 (N945, N902, N363, N5, N461);
nand NAND3 (N946, N927, N245, N216);
xor XOR2 (N947, N945, N899);
and AND4 (N948, N946, N895, N432, N350);
or OR3 (N949, N938, N615, N817);
nand NAND4 (N950, N947, N92, N218, N826);
and AND2 (N951, N942, N660);
not NOT1 (N952, N929);
or OR4 (N953, N949, N265, N194, N905);
buf BUF1 (N954, N950);
buf BUF1 (N955, N952);
and AND4 (N956, N939, N406, N644, N157);
nand NAND4 (N957, N953, N396, N477, N132);
and AND3 (N958, N955, N675, N86);
xor XOR2 (N959, N944, N80);
or OR2 (N960, N951, N837);
nor NOR3 (N961, N948, N852, N129);
buf BUF1 (N962, N943);
buf BUF1 (N963, N954);
nand NAND3 (N964, N956, N468, N321);
not NOT1 (N965, N963);
nor NOR3 (N966, N964, N622, N734);
and AND4 (N967, N966, N934, N349, N341);
and AND4 (N968, N967, N18, N477, N280);
and AND4 (N969, N961, N422, N585, N893);
buf BUF1 (N970, N959);
or OR3 (N971, N969, N200, N44);
buf BUF1 (N972, N960);
and AND3 (N973, N962, N418, N847);
nand NAND2 (N974, N965, N727);
and AND3 (N975, N974, N780, N905);
nor NOR4 (N976, N970, N705, N632, N277);
not NOT1 (N977, N968);
and AND2 (N978, N975, N613);
not NOT1 (N979, N971);
or OR2 (N980, N930, N715);
nand NAND2 (N981, N957, N429);
buf BUF1 (N982, N980);
and AND2 (N983, N977, N688);
or OR4 (N984, N958, N845, N135, N739);
buf BUF1 (N985, N982);
and AND3 (N986, N984, N186, N260);
buf BUF1 (N987, N985);
and AND3 (N988, N972, N117, N784);
and AND3 (N989, N986, N206, N207);
or OR4 (N990, N987, N777, N312, N385);
nand NAND4 (N991, N941, N219, N682, N696);
nor NOR3 (N992, N991, N305, N456);
buf BUF1 (N993, N990);
or OR4 (N994, N983, N273, N95, N286);
or OR3 (N995, N994, N317, N298);
not NOT1 (N996, N992);
xor XOR2 (N997, N973, N79);
and AND2 (N998, N981, N713);
xor XOR2 (N999, N997, N108);
nor NOR2 (N1000, N996, N605);
or OR3 (N1001, N995, N219, N417);
not NOT1 (N1002, N989);
and AND2 (N1003, N979, N979);
and AND4 (N1004, N978, N702, N728, N214);
nor NOR3 (N1005, N1004, N643, N239);
nand NAND4 (N1006, N999, N849, N394, N918);
xor XOR2 (N1007, N988, N337);
xor XOR2 (N1008, N1003, N474);
not NOT1 (N1009, N976);
nand NAND4 (N1010, N993, N338, N756, N232);
and AND4 (N1011, N1009, N234, N733, N51);
nor NOR4 (N1012, N1002, N174, N421, N718);
xor XOR2 (N1013, N1001, N540);
nor NOR2 (N1014, N1013, N826);
buf BUF1 (N1015, N1006);
xor XOR2 (N1016, N1010, N130);
not NOT1 (N1017, N1014);
nor NOR3 (N1018, N1017, N434, N1004);
or OR3 (N1019, N1000, N526, N900);
nand NAND2 (N1020, N1015, N894);
or OR4 (N1021, N1005, N138, N925, N964);
and AND2 (N1022, N1020, N255);
nand NAND4 (N1023, N1019, N949, N360, N551);
buf BUF1 (N1024, N1012);
buf BUF1 (N1025, N1018);
buf BUF1 (N1026, N1016);
buf BUF1 (N1027, N1011);
xor XOR2 (N1028, N1024, N228);
or OR2 (N1029, N1008, N682);
or OR3 (N1030, N1027, N376, N469);
and AND4 (N1031, N1022, N576, N22, N1017);
buf BUF1 (N1032, N1030);
nor NOR4 (N1033, N1032, N564, N1003, N320);
nand NAND2 (N1034, N1026, N535);
not NOT1 (N1035, N1023);
nor NOR2 (N1036, N1029, N52);
xor XOR2 (N1037, N998, N366);
or OR2 (N1038, N1034, N267);
xor XOR2 (N1039, N1036, N208);
not NOT1 (N1040, N1037);
or OR2 (N1041, N1021, N122);
not NOT1 (N1042, N1031);
and AND2 (N1043, N1038, N923);
or OR3 (N1044, N1033, N275, N420);
or OR4 (N1045, N1039, N859, N302, N84);
not NOT1 (N1046, N1044);
buf BUF1 (N1047, N1041);
nor NOR4 (N1048, N1028, N1028, N175, N836);
xor XOR2 (N1049, N1007, N472);
and AND3 (N1050, N1048, N832, N581);
xor XOR2 (N1051, N1049, N999);
buf BUF1 (N1052, N1050);
xor XOR2 (N1053, N1043, N395);
xor XOR2 (N1054, N1035, N956);
not NOT1 (N1055, N1047);
nor NOR4 (N1056, N1054, N471, N474, N525);
or OR3 (N1057, N1042, N887, N95);
nor NOR3 (N1058, N1052, N208, N345);
nand NAND2 (N1059, N1056, N45);
nor NOR2 (N1060, N1025, N897);
buf BUF1 (N1061, N1053);
xor XOR2 (N1062, N1060, N209);
and AND3 (N1063, N1061, N85, N912);
and AND2 (N1064, N1057, N134);
buf BUF1 (N1065, N1064);
nand NAND4 (N1066, N1051, N356, N360, N137);
and AND4 (N1067, N1055, N95, N543, N297);
nand NAND2 (N1068, N1058, N84);
not NOT1 (N1069, N1062);
buf BUF1 (N1070, N1059);
nor NOR4 (N1071, N1066, N123, N156, N609);
xor XOR2 (N1072, N1071, N244);
nor NOR3 (N1073, N1063, N973, N774);
nor NOR2 (N1074, N1045, N30);
not NOT1 (N1075, N1070);
or OR3 (N1076, N1075, N141, N768);
xor XOR2 (N1077, N1072, N581);
nor NOR2 (N1078, N1040, N19);
buf BUF1 (N1079, N1078);
nand NAND4 (N1080, N1074, N1060, N262, N1062);
or OR3 (N1081, N1046, N502, N899);
nand NAND4 (N1082, N1068, N656, N737, N600);
xor XOR2 (N1083, N1076, N831);
nand NAND3 (N1084, N1083, N536, N969);
not NOT1 (N1085, N1084);
nand NAND4 (N1086, N1079, N652, N566, N999);
or OR3 (N1087, N1073, N982, N924);
buf BUF1 (N1088, N1081);
nor NOR3 (N1089, N1085, N335, N399);
not NOT1 (N1090, N1082);
nor NOR4 (N1091, N1069, N914, N811, N174);
or OR2 (N1092, N1088, N806);
nor NOR4 (N1093, N1089, N599, N633, N261);
or OR4 (N1094, N1065, N499, N530, N48);
and AND3 (N1095, N1093, N452, N9);
xor XOR2 (N1096, N1095, N314);
xor XOR2 (N1097, N1092, N906);
nor NOR3 (N1098, N1096, N552, N200);
xor XOR2 (N1099, N1080, N943);
or OR2 (N1100, N1086, N189);
and AND4 (N1101, N1094, N1018, N271, N368);
not NOT1 (N1102, N1097);
nand NAND3 (N1103, N1098, N592, N510);
nand NAND3 (N1104, N1087, N124, N362);
xor XOR2 (N1105, N1104, N914);
buf BUF1 (N1106, N1077);
and AND3 (N1107, N1106, N720, N1007);
nand NAND2 (N1108, N1099, N25);
or OR2 (N1109, N1102, N812);
nor NOR4 (N1110, N1103, N1012, N186, N147);
nand NAND4 (N1111, N1108, N1082, N276, N103);
nor NOR4 (N1112, N1110, N665, N456, N421);
xor XOR2 (N1113, N1109, N834);
nand NAND4 (N1114, N1100, N132, N1087, N666);
or OR2 (N1115, N1091, N582);
nand NAND3 (N1116, N1101, N657, N1080);
buf BUF1 (N1117, N1111);
nor NOR2 (N1118, N1114, N636);
or OR2 (N1119, N1112, N847);
not NOT1 (N1120, N1067);
nor NOR3 (N1121, N1118, N1101, N511);
xor XOR2 (N1122, N1120, N825);
nor NOR3 (N1123, N1115, N1113, N561);
and AND4 (N1124, N1000, N752, N556, N746);
and AND4 (N1125, N1107, N416, N697, N959);
or OR3 (N1126, N1105, N173, N1094);
nand NAND4 (N1127, N1117, N844, N9, N841);
and AND3 (N1128, N1124, N948, N225);
nor NOR4 (N1129, N1121, N476, N527, N95);
nor NOR2 (N1130, N1119, N1018);
or OR3 (N1131, N1125, N524, N531);
nand NAND4 (N1132, N1126, N569, N729, N205);
buf BUF1 (N1133, N1132);
and AND3 (N1134, N1130, N1097, N22);
or OR3 (N1135, N1128, N273, N408);
and AND4 (N1136, N1090, N109, N687, N989);
xor XOR2 (N1137, N1134, N826);
nor NOR3 (N1138, N1135, N306, N182);
not NOT1 (N1139, N1133);
nand NAND2 (N1140, N1139, N513);
buf BUF1 (N1141, N1131);
xor XOR2 (N1142, N1136, N530);
not NOT1 (N1143, N1142);
buf BUF1 (N1144, N1127);
buf BUF1 (N1145, N1138);
nor NOR3 (N1146, N1116, N91, N268);
nand NAND4 (N1147, N1123, N517, N642, N191);
buf BUF1 (N1148, N1141);
or OR2 (N1149, N1143, N381);
nor NOR2 (N1150, N1129, N787);
nor NOR2 (N1151, N1145, N862);
nor NOR3 (N1152, N1151, N249, N640);
nand NAND2 (N1153, N1149, N236);
buf BUF1 (N1154, N1122);
xor XOR2 (N1155, N1153, N829);
xor XOR2 (N1156, N1146, N631);
and AND4 (N1157, N1154, N578, N610, N1146);
buf BUF1 (N1158, N1144);
buf BUF1 (N1159, N1157);
or OR2 (N1160, N1158, N832);
nor NOR3 (N1161, N1140, N697, N368);
nor NOR3 (N1162, N1161, N372, N1139);
not NOT1 (N1163, N1159);
nor NOR4 (N1164, N1150, N131, N484, N123);
or OR4 (N1165, N1163, N863, N735, N333);
and AND2 (N1166, N1165, N565);
and AND4 (N1167, N1156, N1109, N504, N399);
xor XOR2 (N1168, N1167, N540);
and AND3 (N1169, N1166, N1035, N1132);
or OR2 (N1170, N1137, N963);
and AND4 (N1171, N1164, N150, N1049, N27);
or OR3 (N1172, N1162, N37, N737);
nand NAND2 (N1173, N1169, N763);
buf BUF1 (N1174, N1148);
nand NAND2 (N1175, N1171, N399);
xor XOR2 (N1176, N1172, N207);
xor XOR2 (N1177, N1176, N778);
and AND2 (N1178, N1170, N491);
or OR2 (N1179, N1174, N1170);
xor XOR2 (N1180, N1152, N592);
and AND4 (N1181, N1155, N983, N433, N1093);
nor NOR4 (N1182, N1180, N745, N255, N1031);
buf BUF1 (N1183, N1175);
nor NOR4 (N1184, N1179, N303, N703, N1099);
nor NOR2 (N1185, N1178, N634);
or OR3 (N1186, N1173, N1059, N754);
not NOT1 (N1187, N1168);
xor XOR2 (N1188, N1182, N619);
not NOT1 (N1189, N1160);
buf BUF1 (N1190, N1187);
nor NOR2 (N1191, N1186, N951);
nand NAND2 (N1192, N1190, N563);
or OR3 (N1193, N1185, N644, N212);
buf BUF1 (N1194, N1192);
nor NOR3 (N1195, N1193, N509, N975);
or OR3 (N1196, N1177, N650, N246);
or OR3 (N1197, N1183, N385, N1015);
nand NAND3 (N1198, N1195, N343, N153);
nand NAND4 (N1199, N1189, N515, N380, N538);
or OR2 (N1200, N1198, N974);
xor XOR2 (N1201, N1191, N991);
nor NOR4 (N1202, N1184, N809, N138, N147);
or OR4 (N1203, N1181, N225, N169, N515);
nand NAND4 (N1204, N1196, N1014, N594, N995);
buf BUF1 (N1205, N1202);
and AND2 (N1206, N1204, N440);
not NOT1 (N1207, N1203);
and AND2 (N1208, N1201, N1112);
nor NOR4 (N1209, N1194, N1141, N639, N30);
xor XOR2 (N1210, N1200, N837);
and AND3 (N1211, N1205, N320, N576);
xor XOR2 (N1212, N1207, N578);
nor NOR3 (N1213, N1210, N167, N1203);
and AND3 (N1214, N1206, N953, N446);
buf BUF1 (N1215, N1197);
xor XOR2 (N1216, N1208, N726);
nor NOR4 (N1217, N1188, N1168, N803, N697);
nand NAND3 (N1218, N1214, N469, N112);
buf BUF1 (N1219, N1147);
not NOT1 (N1220, N1213);
buf BUF1 (N1221, N1212);
xor XOR2 (N1222, N1215, N632);
not NOT1 (N1223, N1211);
nand NAND4 (N1224, N1221, N939, N188, N1002);
not NOT1 (N1225, N1209);
nor NOR3 (N1226, N1223, N765, N1201);
nor NOR4 (N1227, N1224, N848, N795, N1146);
buf BUF1 (N1228, N1219);
xor XOR2 (N1229, N1228, N647);
not NOT1 (N1230, N1216);
not NOT1 (N1231, N1220);
nor NOR3 (N1232, N1227, N557, N708);
or OR4 (N1233, N1199, N1029, N778, N1200);
nor NOR3 (N1234, N1231, N941, N523);
nor NOR4 (N1235, N1225, N84, N908, N111);
buf BUF1 (N1236, N1235);
nor NOR3 (N1237, N1233, N371, N746);
and AND4 (N1238, N1229, N574, N784, N884);
nor NOR4 (N1239, N1238, N1119, N295, N1020);
or OR3 (N1240, N1217, N931, N313);
or OR2 (N1241, N1222, N204);
xor XOR2 (N1242, N1237, N398);
buf BUF1 (N1243, N1242);
and AND2 (N1244, N1226, N294);
nand NAND2 (N1245, N1244, N286);
and AND4 (N1246, N1232, N164, N83, N697);
nand NAND4 (N1247, N1243, N405, N1018, N125);
nand NAND4 (N1248, N1239, N1114, N547, N1226);
nor NOR2 (N1249, N1234, N947);
and AND4 (N1250, N1218, N319, N931, N699);
nor NOR3 (N1251, N1250, N450, N892);
or OR4 (N1252, N1246, N383, N47, N1151);
nor NOR4 (N1253, N1249, N1043, N1118, N10);
and AND2 (N1254, N1248, N246);
and AND2 (N1255, N1240, N1214);
or OR3 (N1256, N1247, N1134, N997);
not NOT1 (N1257, N1254);
nor NOR4 (N1258, N1257, N668, N463, N1028);
buf BUF1 (N1259, N1255);
buf BUF1 (N1260, N1256);
nand NAND2 (N1261, N1258, N402);
nor NOR2 (N1262, N1259, N873);
xor XOR2 (N1263, N1261, N838);
or OR2 (N1264, N1262, N1169);
buf BUF1 (N1265, N1241);
buf BUF1 (N1266, N1253);
nand NAND3 (N1267, N1245, N971, N906);
and AND3 (N1268, N1263, N1122, N403);
nor NOR2 (N1269, N1252, N1099);
buf BUF1 (N1270, N1264);
and AND4 (N1271, N1270, N135, N406, N533);
buf BUF1 (N1272, N1267);
xor XOR2 (N1273, N1230, N338);
and AND3 (N1274, N1271, N1159, N948);
not NOT1 (N1275, N1272);
xor XOR2 (N1276, N1273, N1214);
buf BUF1 (N1277, N1260);
xor XOR2 (N1278, N1265, N553);
xor XOR2 (N1279, N1269, N963);
nor NOR3 (N1280, N1274, N236, N764);
nor NOR4 (N1281, N1266, N1034, N894, N728);
xor XOR2 (N1282, N1268, N1011);
buf BUF1 (N1283, N1251);
nand NAND4 (N1284, N1275, N1177, N671, N881);
xor XOR2 (N1285, N1280, N157);
not NOT1 (N1286, N1283);
and AND4 (N1287, N1282, N109, N506, N385);
buf BUF1 (N1288, N1278);
or OR3 (N1289, N1277, N316, N943);
nand NAND3 (N1290, N1289, N1056, N799);
buf BUF1 (N1291, N1279);
nand NAND4 (N1292, N1286, N727, N243, N58);
nor NOR3 (N1293, N1284, N855, N885);
nor NOR3 (N1294, N1281, N556, N513);
xor XOR2 (N1295, N1236, N253);
nand NAND4 (N1296, N1287, N185, N21, N1141);
nand NAND4 (N1297, N1291, N21, N456, N748);
not NOT1 (N1298, N1296);
nor NOR2 (N1299, N1294, N1290);
xor XOR2 (N1300, N1277, N674);
nand NAND4 (N1301, N1298, N1094, N1248, N183);
buf BUF1 (N1302, N1292);
or OR3 (N1303, N1276, N807, N1047);
and AND3 (N1304, N1303, N1020, N1288);
buf BUF1 (N1305, N62);
buf BUF1 (N1306, N1304);
nor NOR3 (N1307, N1297, N1225, N593);
xor XOR2 (N1308, N1307, N223);
nand NAND3 (N1309, N1301, N513, N1297);
not NOT1 (N1310, N1308);
not NOT1 (N1311, N1285);
xor XOR2 (N1312, N1299, N920);
xor XOR2 (N1313, N1312, N798);
and AND3 (N1314, N1311, N694, N129);
nand NAND4 (N1315, N1314, N332, N121, N555);
buf BUF1 (N1316, N1315);
or OR3 (N1317, N1305, N776, N182);
or OR2 (N1318, N1295, N1122);
or OR2 (N1319, N1300, N768);
nand NAND4 (N1320, N1318, N342, N1047, N1178);
nand NAND2 (N1321, N1320, N285);
not NOT1 (N1322, N1302);
nand NAND3 (N1323, N1322, N948, N356);
not NOT1 (N1324, N1317);
buf BUF1 (N1325, N1321);
not NOT1 (N1326, N1324);
buf BUF1 (N1327, N1325);
not NOT1 (N1328, N1323);
not NOT1 (N1329, N1327);
nand NAND3 (N1330, N1306, N495, N589);
nand NAND4 (N1331, N1329, N881, N1013, N206);
buf BUF1 (N1332, N1310);
and AND4 (N1333, N1313, N53, N758, N894);
not NOT1 (N1334, N1328);
buf BUF1 (N1335, N1331);
xor XOR2 (N1336, N1335, N15);
and AND3 (N1337, N1330, N708, N1059);
and AND2 (N1338, N1326, N1178);
xor XOR2 (N1339, N1337, N983);
or OR3 (N1340, N1319, N917, N430);
not NOT1 (N1341, N1332);
nand NAND2 (N1342, N1316, N490);
buf BUF1 (N1343, N1293);
nor NOR2 (N1344, N1333, N339);
buf BUF1 (N1345, N1342);
and AND3 (N1346, N1344, N577, N1072);
xor XOR2 (N1347, N1339, N172);
and AND2 (N1348, N1343, N1046);
nor NOR3 (N1349, N1341, N781, N907);
not NOT1 (N1350, N1309);
or OR4 (N1351, N1349, N228, N440, N239);
xor XOR2 (N1352, N1338, N1290);
or OR2 (N1353, N1351, N731);
nor NOR3 (N1354, N1353, N135, N1275);
and AND3 (N1355, N1354, N1198, N503);
nor NOR4 (N1356, N1336, N1195, N209, N224);
xor XOR2 (N1357, N1356, N609);
nor NOR2 (N1358, N1357, N1317);
xor XOR2 (N1359, N1355, N1286);
nor NOR3 (N1360, N1358, N663, N594);
not NOT1 (N1361, N1340);
and AND3 (N1362, N1352, N634, N360);
nand NAND2 (N1363, N1334, N465);
buf BUF1 (N1364, N1345);
buf BUF1 (N1365, N1350);
not NOT1 (N1366, N1359);
or OR4 (N1367, N1348, N1299, N184, N1242);
buf BUF1 (N1368, N1363);
or OR2 (N1369, N1367, N804);
nor NOR2 (N1370, N1369, N1029);
or OR2 (N1371, N1368, N327);
or OR2 (N1372, N1366, N850);
nor NOR2 (N1373, N1364, N710);
nor NOR3 (N1374, N1371, N541, N57);
nor NOR2 (N1375, N1361, N1301);
nand NAND4 (N1376, N1370, N671, N433, N731);
and AND2 (N1377, N1362, N856);
and AND4 (N1378, N1375, N791, N930, N454);
and AND4 (N1379, N1376, N469, N1031, N544);
or OR2 (N1380, N1373, N44);
and AND3 (N1381, N1372, N687, N1123);
nor NOR4 (N1382, N1346, N984, N882, N1311);
xor XOR2 (N1383, N1377, N367);
nand NAND2 (N1384, N1383, N810);
or OR3 (N1385, N1365, N1220, N574);
nand NAND3 (N1386, N1380, N1165, N1384);
or OR3 (N1387, N1061, N1096, N519);
not NOT1 (N1388, N1385);
nand NAND4 (N1389, N1379, N561, N392, N3);
and AND2 (N1390, N1360, N165);
xor XOR2 (N1391, N1390, N108);
buf BUF1 (N1392, N1391);
nand NAND3 (N1393, N1388, N1174, N1091);
buf BUF1 (N1394, N1378);
nor NOR4 (N1395, N1394, N1371, N117, N1290);
xor XOR2 (N1396, N1389, N808);
xor XOR2 (N1397, N1393, N761);
nor NOR3 (N1398, N1396, N152, N551);
nand NAND4 (N1399, N1347, N1089, N588, N380);
and AND4 (N1400, N1395, N927, N897, N234);
nor NOR3 (N1401, N1387, N1165, N99);
xor XOR2 (N1402, N1382, N1135);
xor XOR2 (N1403, N1399, N1006);
not NOT1 (N1404, N1401);
buf BUF1 (N1405, N1392);
and AND4 (N1406, N1402, N851, N645, N879);
xor XOR2 (N1407, N1397, N351);
or OR2 (N1408, N1374, N411);
and AND4 (N1409, N1406, N726, N918, N1275);
nand NAND3 (N1410, N1408, N129, N1198);
nand NAND4 (N1411, N1407, N129, N371, N688);
nor NOR4 (N1412, N1386, N163, N1398, N554);
nand NAND2 (N1413, N461, N153);
nor NOR2 (N1414, N1411, N420);
and AND2 (N1415, N1413, N927);
or OR2 (N1416, N1403, N210);
not NOT1 (N1417, N1415);
nor NOR2 (N1418, N1416, N180);
buf BUF1 (N1419, N1417);
and AND2 (N1420, N1400, N273);
xor XOR2 (N1421, N1404, N18);
not NOT1 (N1422, N1419);
nor NOR4 (N1423, N1410, N929, N176, N452);
or OR3 (N1424, N1405, N1423, N161);
or OR4 (N1425, N306, N902, N262, N886);
or OR3 (N1426, N1409, N377, N1102);
not NOT1 (N1427, N1414);
or OR4 (N1428, N1426, N145, N636, N76);
or OR2 (N1429, N1421, N810);
buf BUF1 (N1430, N1418);
buf BUF1 (N1431, N1412);
not NOT1 (N1432, N1424);
nor NOR2 (N1433, N1429, N188);
nand NAND3 (N1434, N1427, N914, N1267);
xor XOR2 (N1435, N1428, N1064);
not NOT1 (N1436, N1420);
nand NAND4 (N1437, N1434, N788, N205, N459);
and AND2 (N1438, N1430, N1099);
not NOT1 (N1439, N1435);
nand NAND3 (N1440, N1422, N1032, N829);
not NOT1 (N1441, N1432);
not NOT1 (N1442, N1437);
nor NOR2 (N1443, N1439, N348);
nand NAND3 (N1444, N1425, N60, N464);
buf BUF1 (N1445, N1381);
not NOT1 (N1446, N1440);
nand NAND3 (N1447, N1446, N1100, N683);
xor XOR2 (N1448, N1442, N354);
or OR2 (N1449, N1441, N439);
not NOT1 (N1450, N1449);
or OR2 (N1451, N1444, N808);
and AND2 (N1452, N1431, N811);
and AND2 (N1453, N1438, N1024);
nor NOR2 (N1454, N1443, N1374);
not NOT1 (N1455, N1445);
nor NOR2 (N1456, N1450, N289);
and AND4 (N1457, N1451, N1063, N419, N358);
and AND2 (N1458, N1447, N1136);
buf BUF1 (N1459, N1452);
nor NOR4 (N1460, N1459, N451, N1001, N239);
buf BUF1 (N1461, N1453);
buf BUF1 (N1462, N1457);
nor NOR2 (N1463, N1460, N58);
nand NAND2 (N1464, N1456, N266);
or OR2 (N1465, N1454, N1415);
xor XOR2 (N1466, N1455, N236);
xor XOR2 (N1467, N1464, N145);
xor XOR2 (N1468, N1463, N1396);
xor XOR2 (N1469, N1468, N821);
buf BUF1 (N1470, N1461);
nand NAND3 (N1471, N1469, N582, N891);
and AND4 (N1472, N1467, N394, N785, N1288);
xor XOR2 (N1473, N1470, N876);
xor XOR2 (N1474, N1466, N635);
buf BUF1 (N1475, N1448);
not NOT1 (N1476, N1472);
and AND4 (N1477, N1465, N358, N684, N55);
not NOT1 (N1478, N1436);
xor XOR2 (N1479, N1433, N53);
buf BUF1 (N1480, N1477);
and AND3 (N1481, N1471, N179, N580);
nor NOR3 (N1482, N1474, N1121, N811);
and AND2 (N1483, N1475, N637);
buf BUF1 (N1484, N1458);
xor XOR2 (N1485, N1482, N863);
not NOT1 (N1486, N1480);
nor NOR4 (N1487, N1481, N727, N782, N29);
not NOT1 (N1488, N1479);
not NOT1 (N1489, N1487);
and AND4 (N1490, N1473, N122, N961, N547);
buf BUF1 (N1491, N1483);
and AND3 (N1492, N1485, N1076, N1042);
xor XOR2 (N1493, N1491, N438);
nand NAND2 (N1494, N1486, N766);
not NOT1 (N1495, N1492);
nor NOR3 (N1496, N1495, N1220, N725);
xor XOR2 (N1497, N1493, N174);
not NOT1 (N1498, N1462);
buf BUF1 (N1499, N1488);
and AND3 (N1500, N1484, N952, N1416);
or OR4 (N1501, N1498, N651, N825, N336);
or OR3 (N1502, N1496, N811, N1401);
buf BUF1 (N1503, N1501);
and AND2 (N1504, N1489, N374);
nor NOR4 (N1505, N1478, N1177, N420, N488);
xor XOR2 (N1506, N1505, N390);
nor NOR3 (N1507, N1494, N449, N1182);
buf BUF1 (N1508, N1476);
xor XOR2 (N1509, N1508, N569);
nor NOR2 (N1510, N1502, N547);
buf BUF1 (N1511, N1510);
buf BUF1 (N1512, N1503);
nor NOR2 (N1513, N1497, N401);
nand NAND3 (N1514, N1512, N1281, N290);
or OR4 (N1515, N1514, N321, N557, N1463);
and AND2 (N1516, N1515, N1128);
buf BUF1 (N1517, N1490);
buf BUF1 (N1518, N1507);
nor NOR4 (N1519, N1511, N238, N1267, N75);
xor XOR2 (N1520, N1504, N1188);
and AND3 (N1521, N1519, N1214, N397);
xor XOR2 (N1522, N1500, N932);
buf BUF1 (N1523, N1516);
not NOT1 (N1524, N1522);
xor XOR2 (N1525, N1524, N1302);
xor XOR2 (N1526, N1499, N1186);
buf BUF1 (N1527, N1513);
buf BUF1 (N1528, N1525);
nor NOR4 (N1529, N1520, N807, N90, N546);
buf BUF1 (N1530, N1529);
and AND4 (N1531, N1527, N314, N1315, N1158);
or OR2 (N1532, N1506, N535);
nor NOR3 (N1533, N1532, N971, N1423);
or OR4 (N1534, N1531, N80, N920, N1054);
not NOT1 (N1535, N1533);
and AND3 (N1536, N1530, N913, N299);
nor NOR2 (N1537, N1526, N1487);
buf BUF1 (N1538, N1535);
nor NOR4 (N1539, N1509, N1382, N1043, N907);
not NOT1 (N1540, N1536);
xor XOR2 (N1541, N1528, N740);
xor XOR2 (N1542, N1541, N1514);
buf BUF1 (N1543, N1542);
nand NAND4 (N1544, N1538, N1391, N586, N281);
nand NAND4 (N1545, N1517, N926, N1436, N624);
nand NAND2 (N1546, N1539, N753);
xor XOR2 (N1547, N1518, N13);
nand NAND4 (N1548, N1540, N1188, N1448, N775);
nor NOR3 (N1549, N1545, N121, N1300);
buf BUF1 (N1550, N1534);
nand NAND3 (N1551, N1521, N719, N1491);
xor XOR2 (N1552, N1551, N1181);
nand NAND4 (N1553, N1537, N1089, N1369, N776);
buf BUF1 (N1554, N1549);
buf BUF1 (N1555, N1554);
nand NAND3 (N1556, N1552, N712, N1278);
xor XOR2 (N1557, N1548, N984);
xor XOR2 (N1558, N1546, N254);
nand NAND2 (N1559, N1550, N272);
buf BUF1 (N1560, N1559);
xor XOR2 (N1561, N1555, N810);
buf BUF1 (N1562, N1544);
and AND4 (N1563, N1543, N334, N165, N1240);
and AND3 (N1564, N1558, N1159, N431);
buf BUF1 (N1565, N1563);
buf BUF1 (N1566, N1553);
nor NOR4 (N1567, N1557, N658, N439, N871);
or OR4 (N1568, N1566, N601, N1436, N808);
nor NOR3 (N1569, N1567, N900, N1488);
xor XOR2 (N1570, N1562, N596);
buf BUF1 (N1571, N1564);
buf BUF1 (N1572, N1565);
and AND2 (N1573, N1569, N1557);
xor XOR2 (N1574, N1556, N777);
buf BUF1 (N1575, N1523);
nor NOR3 (N1576, N1572, N57, N600);
nand NAND4 (N1577, N1576, N1048, N968, N443);
buf BUF1 (N1578, N1560);
or OR4 (N1579, N1575, N597, N1251, N252);
xor XOR2 (N1580, N1561, N236);
nor NOR2 (N1581, N1577, N1130);
nor NOR2 (N1582, N1581, N1131);
xor XOR2 (N1583, N1573, N1247);
and AND4 (N1584, N1568, N963, N1443, N1564);
xor XOR2 (N1585, N1582, N358);
buf BUF1 (N1586, N1578);
xor XOR2 (N1587, N1585, N72);
nand NAND3 (N1588, N1547, N794, N771);
or OR3 (N1589, N1588, N412, N1432);
and AND4 (N1590, N1583, N543, N629, N1335);
xor XOR2 (N1591, N1570, N521);
xor XOR2 (N1592, N1579, N707);
nor NOR3 (N1593, N1571, N1003, N34);
nor NOR2 (N1594, N1590, N891);
and AND3 (N1595, N1589, N405, N764);
and AND2 (N1596, N1580, N8);
xor XOR2 (N1597, N1592, N522);
or OR4 (N1598, N1595, N875, N1305, N1110);
xor XOR2 (N1599, N1587, N991);
xor XOR2 (N1600, N1574, N369);
nand NAND3 (N1601, N1597, N774, N262);
nand NAND4 (N1602, N1594, N1005, N584, N1515);
or OR3 (N1603, N1599, N1209, N1328);
not NOT1 (N1604, N1593);
not NOT1 (N1605, N1600);
nand NAND2 (N1606, N1603, N1346);
nor NOR3 (N1607, N1604, N75, N1003);
xor XOR2 (N1608, N1598, N1586);
xor XOR2 (N1609, N840, N1090);
buf BUF1 (N1610, N1608);
buf BUF1 (N1611, N1596);
and AND4 (N1612, N1602, N738, N915, N747);
and AND3 (N1613, N1609, N1569, N688);
nand NAND2 (N1614, N1612, N943);
or OR4 (N1615, N1601, N580, N1273, N1544);
buf BUF1 (N1616, N1591);
nand NAND4 (N1617, N1616, N1427, N1234, N806);
or OR3 (N1618, N1605, N1143, N79);
and AND2 (N1619, N1617, N377);
and AND2 (N1620, N1606, N1515);
and AND3 (N1621, N1611, N892, N1597);
xor XOR2 (N1622, N1621, N1058);
xor XOR2 (N1623, N1620, N1483);
not NOT1 (N1624, N1613);
nor NOR3 (N1625, N1619, N1349, N260);
buf BUF1 (N1626, N1614);
and AND3 (N1627, N1615, N1376, N902);
and AND4 (N1628, N1622, N1209, N352, N589);
and AND3 (N1629, N1584, N1068, N615);
buf BUF1 (N1630, N1627);
or OR2 (N1631, N1610, N623);
not NOT1 (N1632, N1623);
xor XOR2 (N1633, N1628, N976);
nor NOR4 (N1634, N1629, N1322, N112, N1355);
nor NOR3 (N1635, N1633, N610, N635);
and AND4 (N1636, N1607, N93, N575, N330);
or OR3 (N1637, N1631, N1305, N202);
buf BUF1 (N1638, N1636);
not NOT1 (N1639, N1625);
nand NAND2 (N1640, N1638, N798);
nand NAND4 (N1641, N1639, N1328, N1537, N1025);
nor NOR4 (N1642, N1626, N102, N573, N661);
nor NOR4 (N1643, N1634, N1207, N903, N1301);
and AND2 (N1644, N1635, N1211);
nor NOR4 (N1645, N1642, N452, N372, N801);
buf BUF1 (N1646, N1645);
or OR2 (N1647, N1644, N1088);
buf BUF1 (N1648, N1624);
and AND4 (N1649, N1640, N170, N1578, N1364);
or OR4 (N1650, N1649, N879, N1498, N972);
not NOT1 (N1651, N1632);
not NOT1 (N1652, N1646);
or OR3 (N1653, N1650, N1110, N1061);
nor NOR3 (N1654, N1652, N538, N619);
or OR2 (N1655, N1647, N1595);
nand NAND4 (N1656, N1653, N1132, N1012, N1087);
or OR4 (N1657, N1618, N20, N119, N236);
buf BUF1 (N1658, N1643);
xor XOR2 (N1659, N1655, N466);
or OR4 (N1660, N1641, N595, N496, N11);
nor NOR3 (N1661, N1654, N443, N189);
buf BUF1 (N1662, N1656);
and AND4 (N1663, N1651, N1386, N701, N818);
xor XOR2 (N1664, N1658, N349);
buf BUF1 (N1665, N1660);
nor NOR4 (N1666, N1664, N750, N846, N199);
not NOT1 (N1667, N1665);
xor XOR2 (N1668, N1630, N398);
buf BUF1 (N1669, N1648);
xor XOR2 (N1670, N1669, N1336);
buf BUF1 (N1671, N1659);
nand NAND4 (N1672, N1670, N1601, N526, N180);
buf BUF1 (N1673, N1668);
nor NOR4 (N1674, N1672, N1419, N7, N289);
xor XOR2 (N1675, N1657, N559);
buf BUF1 (N1676, N1674);
xor XOR2 (N1677, N1666, N1346);
nor NOR4 (N1678, N1667, N1422, N631, N980);
nand NAND4 (N1679, N1675, N394, N494, N642);
buf BUF1 (N1680, N1662);
nor NOR3 (N1681, N1671, N1461, N1558);
not NOT1 (N1682, N1673);
or OR3 (N1683, N1680, N586, N1544);
nand NAND4 (N1684, N1677, N900, N142, N639);
not NOT1 (N1685, N1663);
nor NOR2 (N1686, N1685, N280);
nor NOR4 (N1687, N1678, N1289, N836, N341);
nor NOR2 (N1688, N1676, N1124);
not NOT1 (N1689, N1637);
xor XOR2 (N1690, N1689, N1194);
xor XOR2 (N1691, N1679, N1151);
and AND2 (N1692, N1687, N530);
and AND2 (N1693, N1661, N1146);
nand NAND3 (N1694, N1684, N218, N519);
not NOT1 (N1695, N1692);
xor XOR2 (N1696, N1694, N349);
nor NOR2 (N1697, N1683, N1545);
not NOT1 (N1698, N1693);
xor XOR2 (N1699, N1695, N1306);
or OR3 (N1700, N1691, N996, N1549);
nand NAND3 (N1701, N1681, N328, N620);
buf BUF1 (N1702, N1700);
nor NOR4 (N1703, N1696, N1226, N94, N501);
and AND4 (N1704, N1702, N320, N637, N1240);
and AND4 (N1705, N1686, N168, N516, N1602);
nor NOR4 (N1706, N1697, N814, N404, N1457);
nand NAND3 (N1707, N1682, N554, N606);
xor XOR2 (N1708, N1701, N485);
and AND3 (N1709, N1698, N344, N326);
or OR4 (N1710, N1688, N153, N499, N1662);
or OR3 (N1711, N1710, N1601, N1294);
not NOT1 (N1712, N1703);
or OR4 (N1713, N1707, N1545, N272, N1144);
and AND2 (N1714, N1704, N360);
buf BUF1 (N1715, N1709);
buf BUF1 (N1716, N1712);
xor XOR2 (N1717, N1716, N352);
not NOT1 (N1718, N1714);
and AND3 (N1719, N1713, N1350, N591);
nor NOR3 (N1720, N1711, N863, N1657);
and AND2 (N1721, N1717, N1163);
buf BUF1 (N1722, N1720);
buf BUF1 (N1723, N1690);
and AND3 (N1724, N1721, N1401, N908);
and AND4 (N1725, N1718, N873, N587, N329);
nand NAND4 (N1726, N1719, N405, N897, N340);
or OR3 (N1727, N1699, N610, N684);
nand NAND4 (N1728, N1706, N1170, N1443, N1035);
buf BUF1 (N1729, N1728);
buf BUF1 (N1730, N1725);
not NOT1 (N1731, N1727);
nand NAND3 (N1732, N1708, N284, N7);
nor NOR4 (N1733, N1731, N166, N1457, N46);
xor XOR2 (N1734, N1715, N1404);
nor NOR3 (N1735, N1729, N1055, N1109);
and AND4 (N1736, N1735, N560, N1438, N725);
buf BUF1 (N1737, N1733);
not NOT1 (N1738, N1705);
buf BUF1 (N1739, N1736);
or OR2 (N1740, N1737, N1118);
buf BUF1 (N1741, N1734);
and AND3 (N1742, N1723, N1249, N1724);
xor XOR2 (N1743, N270, N484);
or OR4 (N1744, N1740, N918, N1208, N1272);
nand NAND4 (N1745, N1741, N1593, N141, N1221);
xor XOR2 (N1746, N1730, N674);
xor XOR2 (N1747, N1739, N1312);
buf BUF1 (N1748, N1743);
nor NOR3 (N1749, N1747, N859, N731);
nor NOR2 (N1750, N1726, N696);
nand NAND3 (N1751, N1746, N1303, N1609);
or OR3 (N1752, N1751, N293, N1470);
and AND2 (N1753, N1748, N1136);
not NOT1 (N1754, N1742);
or OR4 (N1755, N1738, N844, N1024, N1221);
buf BUF1 (N1756, N1754);
xor XOR2 (N1757, N1732, N860);
buf BUF1 (N1758, N1755);
or OR4 (N1759, N1745, N849, N803, N543);
not NOT1 (N1760, N1752);
and AND3 (N1761, N1756, N1214, N482);
nor NOR2 (N1762, N1749, N476);
buf BUF1 (N1763, N1753);
buf BUF1 (N1764, N1762);
nand NAND2 (N1765, N1758, N1653);
or OR4 (N1766, N1744, N598, N1623, N1345);
or OR3 (N1767, N1759, N1743, N1431);
not NOT1 (N1768, N1757);
nand NAND3 (N1769, N1764, N1194, N587);
nand NAND2 (N1770, N1767, N749);
nor NOR4 (N1771, N1765, N1310, N1730, N42);
nand NAND2 (N1772, N1768, N1722);
and AND4 (N1773, N1121, N461, N802, N1286);
buf BUF1 (N1774, N1773);
xor XOR2 (N1775, N1761, N446);
and AND2 (N1776, N1771, N1458);
and AND3 (N1777, N1775, N222, N1743);
nor NOR2 (N1778, N1774, N1497);
buf BUF1 (N1779, N1763);
not NOT1 (N1780, N1750);
nor NOR2 (N1781, N1778, N451);
and AND4 (N1782, N1770, N389, N1681, N1635);
xor XOR2 (N1783, N1769, N1);
nor NOR3 (N1784, N1766, N103, N48);
buf BUF1 (N1785, N1772);
buf BUF1 (N1786, N1785);
nand NAND3 (N1787, N1781, N1451, N294);
and AND4 (N1788, N1787, N588, N1259, N387);
buf BUF1 (N1789, N1786);
buf BUF1 (N1790, N1788);
nor NOR4 (N1791, N1784, N103, N648, N1649);
and AND4 (N1792, N1790, N628, N1617, N1363);
nand NAND3 (N1793, N1777, N1368, N889);
nor NOR2 (N1794, N1782, N805);
or OR2 (N1795, N1776, N1262);
xor XOR2 (N1796, N1795, N1606);
buf BUF1 (N1797, N1760);
nor NOR2 (N1798, N1779, N650);
nand NAND3 (N1799, N1793, N1097, N1423);
nand NAND3 (N1800, N1780, N1674, N613);
and AND2 (N1801, N1789, N347);
or OR2 (N1802, N1796, N373);
nand NAND4 (N1803, N1802, N1445, N717, N1641);
and AND3 (N1804, N1803, N492, N582);
not NOT1 (N1805, N1783);
nand NAND3 (N1806, N1797, N420, N1016);
buf BUF1 (N1807, N1792);
and AND2 (N1808, N1799, N1626);
or OR3 (N1809, N1807, N1492, N1678);
buf BUF1 (N1810, N1809);
or OR2 (N1811, N1794, N1366);
nand NAND3 (N1812, N1810, N1441, N1258);
and AND3 (N1813, N1808, N991, N493);
not NOT1 (N1814, N1801);
buf BUF1 (N1815, N1798);
not NOT1 (N1816, N1805);
not NOT1 (N1817, N1804);
nor NOR4 (N1818, N1811, N221, N1345, N276);
not NOT1 (N1819, N1816);
not NOT1 (N1820, N1813);
and AND3 (N1821, N1820, N194, N554);
buf BUF1 (N1822, N1819);
and AND4 (N1823, N1821, N767, N140, N974);
not NOT1 (N1824, N1817);
or OR2 (N1825, N1823, N1601);
buf BUF1 (N1826, N1800);
nor NOR2 (N1827, N1824, N695);
not NOT1 (N1828, N1822);
nand NAND3 (N1829, N1826, N1823, N627);
and AND3 (N1830, N1791, N1175, N691);
and AND3 (N1831, N1812, N1806, N589);
or OR3 (N1832, N647, N1736, N649);
not NOT1 (N1833, N1831);
buf BUF1 (N1834, N1832);
nand NAND4 (N1835, N1818, N1004, N322, N788);
buf BUF1 (N1836, N1833);
not NOT1 (N1837, N1828);
and AND2 (N1838, N1815, N1747);
buf BUF1 (N1839, N1814);
not NOT1 (N1840, N1838);
buf BUF1 (N1841, N1835);
buf BUF1 (N1842, N1841);
nor NOR2 (N1843, N1830, N398);
not NOT1 (N1844, N1840);
buf BUF1 (N1845, N1839);
buf BUF1 (N1846, N1843);
xor XOR2 (N1847, N1846, N585);
nor NOR4 (N1848, N1844, N1333, N878, N91);
not NOT1 (N1849, N1834);
xor XOR2 (N1850, N1836, N945);
nor NOR3 (N1851, N1849, N1567, N1252);
and AND3 (N1852, N1847, N1047, N59);
not NOT1 (N1853, N1837);
or OR3 (N1854, N1852, N1551, N684);
nor NOR3 (N1855, N1850, N562, N777);
or OR4 (N1856, N1854, N682, N1434, N805);
not NOT1 (N1857, N1825);
nand NAND4 (N1858, N1857, N456, N1755, N252);
and AND2 (N1859, N1848, N953);
nand NAND3 (N1860, N1845, N553, N1178);
xor XOR2 (N1861, N1855, N834);
nand NAND2 (N1862, N1829, N398);
not NOT1 (N1863, N1851);
and AND4 (N1864, N1861, N993, N1704, N601);
and AND4 (N1865, N1853, N1706, N830, N1200);
nor NOR4 (N1866, N1862, N691, N673, N1741);
not NOT1 (N1867, N1842);
or OR2 (N1868, N1863, N1588);
not NOT1 (N1869, N1856);
xor XOR2 (N1870, N1858, N448);
nor NOR2 (N1871, N1859, N225);
xor XOR2 (N1872, N1866, N651);
nor NOR2 (N1873, N1869, N178);
and AND4 (N1874, N1827, N1255, N24, N716);
not NOT1 (N1875, N1867);
nor NOR2 (N1876, N1860, N172);
or OR2 (N1877, N1865, N241);
and AND2 (N1878, N1872, N1227);
buf BUF1 (N1879, N1878);
not NOT1 (N1880, N1873);
xor XOR2 (N1881, N1864, N46);
and AND2 (N1882, N1870, N568);
nand NAND4 (N1883, N1871, N153, N1497, N1584);
or OR2 (N1884, N1882, N922);
nor NOR2 (N1885, N1874, N269);
nand NAND4 (N1886, N1885, N1050, N841, N1665);
and AND3 (N1887, N1886, N27, N721);
or OR4 (N1888, N1876, N1679, N896, N431);
not NOT1 (N1889, N1887);
or OR2 (N1890, N1880, N1819);
xor XOR2 (N1891, N1879, N1576);
or OR4 (N1892, N1877, N1886, N1084, N373);
and AND2 (N1893, N1889, N287);
buf BUF1 (N1894, N1890);
not NOT1 (N1895, N1883);
or OR3 (N1896, N1895, N1415, N36);
buf BUF1 (N1897, N1894);
nand NAND4 (N1898, N1896, N1631, N1012, N1858);
nor NOR4 (N1899, N1898, N597, N821, N29);
and AND4 (N1900, N1892, N542, N783, N287);
nand NAND4 (N1901, N1891, N617, N1027, N522);
nor NOR3 (N1902, N1900, N888, N322);
nand NAND3 (N1903, N1884, N1685, N156);
nand NAND2 (N1904, N1897, N1012);
nand NAND3 (N1905, N1868, N1410, N455);
buf BUF1 (N1906, N1905);
xor XOR2 (N1907, N1881, N1799);
buf BUF1 (N1908, N1899);
or OR2 (N1909, N1888, N663);
xor XOR2 (N1910, N1906, N1305);
nor NOR4 (N1911, N1901, N1282, N1668, N1505);
and AND4 (N1912, N1907, N1739, N29, N208);
and AND2 (N1913, N1909, N664);
xor XOR2 (N1914, N1902, N1868);
nor NOR3 (N1915, N1912, N588, N1309);
buf BUF1 (N1916, N1914);
xor XOR2 (N1917, N1904, N1436);
nand NAND4 (N1918, N1875, N507, N1258, N1603);
and AND3 (N1919, N1908, N903, N1222);
not NOT1 (N1920, N1903);
nand NAND3 (N1921, N1913, N578, N290);
not NOT1 (N1922, N1919);
not NOT1 (N1923, N1917);
nand NAND2 (N1924, N1893, N1191);
nand NAND2 (N1925, N1921, N615);
not NOT1 (N1926, N1922);
nor NOR4 (N1927, N1918, N567, N274, N1730);
buf BUF1 (N1928, N1915);
nand NAND2 (N1929, N1924, N1284);
nand NAND2 (N1930, N1928, N873);
not NOT1 (N1931, N1929);
and AND2 (N1932, N1931, N1124);
not NOT1 (N1933, N1925);
buf BUF1 (N1934, N1910);
buf BUF1 (N1935, N1923);
and AND3 (N1936, N1932, N1540, N618);
or OR4 (N1937, N1927, N689, N941, N1158);
nor NOR2 (N1938, N1935, N755);
xor XOR2 (N1939, N1938, N529);
or OR4 (N1940, N1933, N1227, N1012, N1263);
nor NOR2 (N1941, N1930, N1169);
buf BUF1 (N1942, N1940);
buf BUF1 (N1943, N1916);
xor XOR2 (N1944, N1939, N1332);
buf BUF1 (N1945, N1944);
and AND2 (N1946, N1943, N935);
nor NOR2 (N1947, N1937, N1162);
xor XOR2 (N1948, N1946, N1263);
nor NOR2 (N1949, N1942, N823);
or OR4 (N1950, N1941, N1946, N202, N1658);
not NOT1 (N1951, N1934);
and AND3 (N1952, N1950, N1297, N107);
or OR4 (N1953, N1949, N206, N1385, N286);
not NOT1 (N1954, N1926);
xor XOR2 (N1955, N1952, N1272);
xor XOR2 (N1956, N1947, N957);
and AND2 (N1957, N1951, N1236);
nor NOR2 (N1958, N1936, N1951);
not NOT1 (N1959, N1920);
not NOT1 (N1960, N1948);
and AND4 (N1961, N1956, N1733, N1763, N1209);
not NOT1 (N1962, N1953);
xor XOR2 (N1963, N1961, N1370);
not NOT1 (N1964, N1960);
nand NAND4 (N1965, N1959, N1597, N450, N1621);
nand NAND4 (N1966, N1955, N136, N556, N1862);
buf BUF1 (N1967, N1911);
nand NAND4 (N1968, N1962, N920, N510, N292);
xor XOR2 (N1969, N1945, N1806);
nand NAND3 (N1970, N1957, N987, N819);
nand NAND4 (N1971, N1963, N363, N920, N1258);
or OR4 (N1972, N1965, N1733, N839, N1478);
nor NOR4 (N1973, N1968, N1831, N1867, N324);
or OR3 (N1974, N1954, N523, N88);
buf BUF1 (N1975, N1972);
nand NAND2 (N1976, N1970, N1487);
not NOT1 (N1977, N1964);
buf BUF1 (N1978, N1958);
or OR3 (N1979, N1978, N453, N55);
nor NOR2 (N1980, N1974, N1751);
and AND4 (N1981, N1969, N1786, N64, N336);
buf BUF1 (N1982, N1980);
nor NOR4 (N1983, N1966, N1331, N1662, N1484);
or OR4 (N1984, N1981, N1556, N329, N1594);
nor NOR2 (N1985, N1976, N1629);
and AND2 (N1986, N1973, N108);
and AND4 (N1987, N1975, N127, N1605, N1111);
nand NAND2 (N1988, N1984, N692);
nand NAND2 (N1989, N1967, N1536);
nor NOR2 (N1990, N1983, N143);
nand NAND3 (N1991, N1985, N123, N164);
buf BUF1 (N1992, N1989);
xor XOR2 (N1993, N1971, N1345);
nor NOR2 (N1994, N1986, N350);
or OR3 (N1995, N1994, N1071, N468);
and AND4 (N1996, N1992, N1046, N1940, N822);
and AND4 (N1997, N1982, N1425, N609, N103);
not NOT1 (N1998, N1997);
nor NOR4 (N1999, N1995, N72, N199, N415);
nand NAND4 (N2000, N1990, N263, N1436, N1937);
not NOT1 (N2001, N2000);
nand NAND4 (N2002, N1993, N294, N66, N1871);
buf BUF1 (N2003, N2002);
not NOT1 (N2004, N1998);
and AND4 (N2005, N2003, N1682, N248, N1738);
not NOT1 (N2006, N2004);
not NOT1 (N2007, N1987);
not NOT1 (N2008, N1988);
nand NAND3 (N2009, N2008, N1959, N1531);
nor NOR2 (N2010, N2001, N1788);
xor XOR2 (N2011, N1996, N1238);
and AND4 (N2012, N1999, N1417, N1269, N681);
xor XOR2 (N2013, N2010, N1890);
nand NAND2 (N2014, N2013, N1552);
nand NAND3 (N2015, N2005, N639, N490);
not NOT1 (N2016, N1977);
nor NOR3 (N2017, N1991, N1576, N585);
nand NAND4 (N2018, N2007, N986, N898, N348);
nand NAND2 (N2019, N2015, N1753);
xor XOR2 (N2020, N2009, N87);
xor XOR2 (N2021, N2011, N98);
buf BUF1 (N2022, N2012);
or OR4 (N2023, N2014, N1814, N635, N657);
not NOT1 (N2024, N2020);
nor NOR2 (N2025, N2017, N580);
nor NOR3 (N2026, N2025, N1977, N792);
xor XOR2 (N2027, N2018, N246);
nor NOR2 (N2028, N2021, N1288);
not NOT1 (N2029, N2022);
and AND3 (N2030, N2023, N445, N1877);
nand NAND4 (N2031, N2024, N1964, N1499, N974);
nand NAND2 (N2032, N2019, N1249);
nand NAND3 (N2033, N2030, N376, N1679);
xor XOR2 (N2034, N2031, N1880);
xor XOR2 (N2035, N2034, N1637);
not NOT1 (N2036, N2026);
nand NAND3 (N2037, N2029, N7, N40);
not NOT1 (N2038, N2027);
and AND2 (N2039, N1979, N254);
nand NAND3 (N2040, N2016, N1355, N1449);
not NOT1 (N2041, N2036);
buf BUF1 (N2042, N2041);
and AND2 (N2043, N2039, N826);
and AND3 (N2044, N2033, N1676, N541);
and AND4 (N2045, N2043, N1174, N339, N1817);
or OR2 (N2046, N2037, N488);
or OR2 (N2047, N2032, N743);
not NOT1 (N2048, N2040);
nor NOR3 (N2049, N2042, N650, N1037);
buf BUF1 (N2050, N2038);
xor XOR2 (N2051, N2006, N444);
not NOT1 (N2052, N2048);
buf BUF1 (N2053, N2051);
xor XOR2 (N2054, N2028, N891);
buf BUF1 (N2055, N2044);
buf BUF1 (N2056, N2053);
or OR4 (N2057, N2050, N1562, N486, N70);
buf BUF1 (N2058, N2046);
nor NOR4 (N2059, N2054, N1521, N1954, N27);
or OR2 (N2060, N2057, N1623);
not NOT1 (N2061, N2059);
nand NAND3 (N2062, N2058, N1439, N1590);
nand NAND3 (N2063, N2047, N1851, N2017);
nor NOR2 (N2064, N2049, N956);
xor XOR2 (N2065, N2035, N1564);
and AND3 (N2066, N2063, N1548, N1000);
buf BUF1 (N2067, N2045);
buf BUF1 (N2068, N2065);
xor XOR2 (N2069, N2066, N227);
not NOT1 (N2070, N2067);
or OR4 (N2071, N2062, N1225, N909, N120);
and AND3 (N2072, N2056, N407, N1481);
nor NOR2 (N2073, N2052, N568);
and AND3 (N2074, N2061, N1148, N1259);
and AND4 (N2075, N2072, N623, N1834, N828);
buf BUF1 (N2076, N2064);
and AND2 (N2077, N2076, N1627);
and AND3 (N2078, N2071, N461, N1675);
nand NAND2 (N2079, N2074, N1840);
nand NAND4 (N2080, N2073, N1976, N1515, N610);
buf BUF1 (N2081, N2075);
or OR3 (N2082, N2078, N1204, N1833);
and AND2 (N2083, N2077, N1005);
and AND3 (N2084, N2068, N890, N2063);
nand NAND2 (N2085, N2082, N415);
and AND4 (N2086, N2060, N673, N101, N1587);
or OR2 (N2087, N2084, N1793);
xor XOR2 (N2088, N2070, N817);
or OR2 (N2089, N2085, N603);
nor NOR3 (N2090, N2080, N22, N1994);
nand NAND2 (N2091, N2087, N177);
xor XOR2 (N2092, N2069, N1481);
and AND2 (N2093, N2055, N1657);
nor NOR4 (N2094, N2081, N801, N1944, N74);
xor XOR2 (N2095, N2083, N677);
or OR2 (N2096, N2088, N465);
or OR3 (N2097, N2096, N1773, N1429);
nand NAND3 (N2098, N2097, N750, N854);
not NOT1 (N2099, N2090);
not NOT1 (N2100, N2094);
xor XOR2 (N2101, N2093, N1706);
or OR2 (N2102, N2101, N1819);
buf BUF1 (N2103, N2089);
not NOT1 (N2104, N2098);
xor XOR2 (N2105, N2103, N1955);
xor XOR2 (N2106, N2099, N1370);
and AND4 (N2107, N2105, N1134, N293, N1565);
not NOT1 (N2108, N2091);
or OR3 (N2109, N2092, N1913, N878);
not NOT1 (N2110, N2109);
buf BUF1 (N2111, N2102);
not NOT1 (N2112, N2104);
nor NOR3 (N2113, N2086, N1136, N1032);
nand NAND4 (N2114, N2095, N725, N1434, N1326);
xor XOR2 (N2115, N2100, N1512);
or OR4 (N2116, N2111, N1106, N1411, N1612);
not NOT1 (N2117, N2115);
and AND4 (N2118, N2117, N1895, N13, N998);
not NOT1 (N2119, N2108);
or OR4 (N2120, N2106, N1042, N1811, N595);
nor NOR2 (N2121, N2116, N1062);
xor XOR2 (N2122, N2120, N664);
nand NAND4 (N2123, N2118, N1811, N240, N1272);
nor NOR4 (N2124, N2107, N1038, N716, N965);
buf BUF1 (N2125, N2112);
nand NAND4 (N2126, N2113, N1465, N2033, N1686);
and AND2 (N2127, N2114, N996);
and AND2 (N2128, N2079, N1988);
not NOT1 (N2129, N2124);
xor XOR2 (N2130, N2121, N2005);
nor NOR2 (N2131, N2129, N951);
and AND4 (N2132, N2110, N913, N8, N617);
nor NOR2 (N2133, N2125, N1594);
and AND2 (N2134, N2119, N706);
buf BUF1 (N2135, N2127);
xor XOR2 (N2136, N2122, N353);
or OR4 (N2137, N2136, N1056, N393, N1406);
and AND4 (N2138, N2130, N1117, N236, N638);
and AND2 (N2139, N2133, N2001);
xor XOR2 (N2140, N2135, N773);
nand NAND2 (N2141, N2123, N888);
not NOT1 (N2142, N2140);
and AND3 (N2143, N2126, N1392, N1166);
not NOT1 (N2144, N2137);
nor NOR4 (N2145, N2144, N1625, N1011, N1999);
xor XOR2 (N2146, N2134, N164);
nor NOR2 (N2147, N2128, N1795);
not NOT1 (N2148, N2143);
xor XOR2 (N2149, N2139, N749);
nand NAND2 (N2150, N2131, N1335);
buf BUF1 (N2151, N2132);
and AND3 (N2152, N2141, N637, N449);
xor XOR2 (N2153, N2150, N689);
nand NAND3 (N2154, N2148, N806, N1459);
nor NOR3 (N2155, N2151, N2084, N73);
buf BUF1 (N2156, N2147);
and AND4 (N2157, N2145, N395, N1900, N519);
or OR3 (N2158, N2153, N1644, N1836);
nand NAND4 (N2159, N2138, N807, N1250, N1207);
not NOT1 (N2160, N2142);
and AND3 (N2161, N2159, N1560, N1969);
nand NAND4 (N2162, N2157, N263, N473, N351);
nor NOR4 (N2163, N2149, N2068, N1013, N830);
xor XOR2 (N2164, N2162, N1616);
buf BUF1 (N2165, N2160);
xor XOR2 (N2166, N2146, N1628);
nor NOR2 (N2167, N2152, N697);
xor XOR2 (N2168, N2163, N1595);
nor NOR2 (N2169, N2155, N1851);
not NOT1 (N2170, N2156);
nand NAND4 (N2171, N2161, N2047, N1600, N1747);
buf BUF1 (N2172, N2168);
nand NAND2 (N2173, N2169, N825);
nand NAND2 (N2174, N2170, N1956);
and AND2 (N2175, N2158, N359);
and AND2 (N2176, N2164, N21);
xor XOR2 (N2177, N2173, N169);
nor NOR2 (N2178, N2172, N174);
xor XOR2 (N2179, N2165, N455);
or OR2 (N2180, N2176, N420);
nand NAND2 (N2181, N2166, N401);
not NOT1 (N2182, N2180);
nand NAND3 (N2183, N2177, N817, N47);
and AND4 (N2184, N2171, N525, N441, N2056);
buf BUF1 (N2185, N2184);
not NOT1 (N2186, N2178);
and AND3 (N2187, N2181, N29, N1992);
or OR3 (N2188, N2183, N370, N341);
nor NOR2 (N2189, N2167, N2083);
or OR3 (N2190, N2187, N1378, N1442);
buf BUF1 (N2191, N2185);
nor NOR2 (N2192, N2154, N404);
nor NOR3 (N2193, N2174, N1677, N1152);
nor NOR3 (N2194, N2175, N332, N248);
not NOT1 (N2195, N2179);
nand NAND2 (N2196, N2191, N1911);
not NOT1 (N2197, N2189);
or OR3 (N2198, N2195, N1045, N436);
xor XOR2 (N2199, N2190, N1007);
and AND2 (N2200, N2194, N2135);
nor NOR4 (N2201, N2198, N1932, N738, N161);
not NOT1 (N2202, N2192);
buf BUF1 (N2203, N2200);
nand NAND2 (N2204, N2202, N1063);
and AND4 (N2205, N2182, N455, N1952, N1264);
and AND3 (N2206, N2199, N2115, N728);
and AND2 (N2207, N2197, N1220);
buf BUF1 (N2208, N2201);
or OR4 (N2209, N2208, N65, N2118, N1380);
and AND2 (N2210, N2205, N1651);
or OR4 (N2211, N2209, N1595, N1729, N365);
xor XOR2 (N2212, N2204, N262);
nor NOR4 (N2213, N2212, N2006, N2057, N139);
nand NAND4 (N2214, N2186, N2111, N967, N1868);
nor NOR4 (N2215, N2210, N581, N390, N1501);
not NOT1 (N2216, N2213);
buf BUF1 (N2217, N2216);
nand NAND2 (N2218, N2206, N442);
xor XOR2 (N2219, N2203, N2185);
buf BUF1 (N2220, N2207);
nor NOR3 (N2221, N2211, N1168, N211);
and AND4 (N2222, N2214, N537, N364, N1101);
or OR4 (N2223, N2188, N1107, N1833, N963);
nand NAND2 (N2224, N2219, N1432);
nand NAND4 (N2225, N2215, N2193, N161, N985);
nand NAND2 (N2226, N1647, N880);
and AND2 (N2227, N2223, N674);
nand NAND2 (N2228, N2225, N383);
xor XOR2 (N2229, N2220, N932);
or OR3 (N2230, N2218, N1524, N1954);
buf BUF1 (N2231, N2222);
and AND4 (N2232, N2221, N552, N1272, N1970);
or OR4 (N2233, N2230, N508, N1301, N845);
and AND2 (N2234, N2217, N467);
not NOT1 (N2235, N2232);
xor XOR2 (N2236, N2226, N673);
or OR3 (N2237, N2234, N910, N389);
buf BUF1 (N2238, N2227);
nand NAND4 (N2239, N2196, N1071, N1653, N302);
xor XOR2 (N2240, N2236, N6);
nand NAND3 (N2241, N2229, N1508, N776);
or OR4 (N2242, N2224, N699, N546, N560);
buf BUF1 (N2243, N2237);
xor XOR2 (N2244, N2239, N1959);
buf BUF1 (N2245, N2235);
and AND4 (N2246, N2245, N643, N1197, N1077);
nor NOR2 (N2247, N2240, N2022);
or OR3 (N2248, N2241, N2019, N265);
and AND4 (N2249, N2243, N2048, N1907, N1185);
buf BUF1 (N2250, N2233);
and AND4 (N2251, N2246, N1718, N1838, N1289);
and AND4 (N2252, N2251, N1721, N249, N2023);
or OR2 (N2253, N2242, N301);
not NOT1 (N2254, N2244);
or OR3 (N2255, N2252, N576, N1749);
not NOT1 (N2256, N2247);
and AND3 (N2257, N2248, N1636, N1481);
xor XOR2 (N2258, N2254, N312);
nor NOR4 (N2259, N2228, N1546, N494, N562);
xor XOR2 (N2260, N2231, N590);
buf BUF1 (N2261, N2258);
buf BUF1 (N2262, N2257);
or OR2 (N2263, N2256, N611);
and AND4 (N2264, N2259, N1518, N1571, N319);
or OR2 (N2265, N2249, N1941);
nand NAND3 (N2266, N2238, N1131, N1415);
nor NOR3 (N2267, N2253, N116, N1093);
nand NAND2 (N2268, N2250, N104);
nor NOR3 (N2269, N2255, N974, N1499);
buf BUF1 (N2270, N2265);
nand NAND4 (N2271, N2263, N595, N147, N2064);
or OR2 (N2272, N2261, N1827);
or OR2 (N2273, N2272, N1918);
nor NOR4 (N2274, N2266, N1658, N1124, N1955);
not NOT1 (N2275, N2271);
or OR2 (N2276, N2270, N822);
and AND2 (N2277, N2276, N238);
xor XOR2 (N2278, N2274, N973);
not NOT1 (N2279, N2277);
nand NAND3 (N2280, N2264, N395, N1025);
not NOT1 (N2281, N2268);
not NOT1 (N2282, N2280);
and AND3 (N2283, N2275, N2232, N1327);
nand NAND4 (N2284, N2267, N2205, N615, N1443);
xor XOR2 (N2285, N2282, N166);
nor NOR3 (N2286, N2284, N1222, N1781);
and AND4 (N2287, N2281, N502, N894, N391);
and AND3 (N2288, N2260, N127, N1401);
xor XOR2 (N2289, N2287, N503);
buf BUF1 (N2290, N2262);
buf BUF1 (N2291, N2279);
xor XOR2 (N2292, N2269, N2267);
nor NOR2 (N2293, N2273, N613);
not NOT1 (N2294, N2291);
and AND2 (N2295, N2286, N1891);
and AND3 (N2296, N2289, N888, N1060);
nor NOR3 (N2297, N2292, N1072, N1013);
and AND2 (N2298, N2294, N1359);
not NOT1 (N2299, N2296);
and AND3 (N2300, N2283, N1737, N882);
and AND4 (N2301, N2293, N823, N1769, N1820);
nor NOR3 (N2302, N2278, N1927, N2278);
or OR2 (N2303, N2301, N2082);
or OR3 (N2304, N2297, N748, N1577);
nand NAND2 (N2305, N2300, N1533);
buf BUF1 (N2306, N2298);
not NOT1 (N2307, N2303);
and AND2 (N2308, N2288, N1388);
or OR2 (N2309, N2306, N620);
nand NAND3 (N2310, N2309, N1441, N290);
and AND2 (N2311, N2295, N712);
and AND4 (N2312, N2304, N508, N1608, N1069);
not NOT1 (N2313, N2305);
and AND2 (N2314, N2285, N59);
nand NAND2 (N2315, N2307, N1135);
and AND2 (N2316, N2310, N713);
xor XOR2 (N2317, N2308, N331);
nor NOR4 (N2318, N2316, N1971, N1520, N1091);
nor NOR3 (N2319, N2315, N1559, N2199);
nand NAND3 (N2320, N2290, N835, N577);
nand NAND3 (N2321, N2317, N173, N1071);
buf BUF1 (N2322, N2313);
nand NAND2 (N2323, N2299, N933);
and AND4 (N2324, N2302, N409, N1534, N2150);
not NOT1 (N2325, N2318);
or OR4 (N2326, N2320, N825, N1842, N1117);
nand NAND4 (N2327, N2322, N685, N154, N193);
nor NOR3 (N2328, N2324, N96, N2228);
or OR3 (N2329, N2314, N445, N1841);
nand NAND2 (N2330, N2321, N1111);
nand NAND3 (N2331, N2319, N798, N2274);
nand NAND4 (N2332, N2331, N2202, N1226, N770);
and AND2 (N2333, N2325, N1614);
or OR4 (N2334, N2311, N1983, N640, N70);
xor XOR2 (N2335, N2323, N716);
and AND3 (N2336, N2312, N2040, N858);
nor NOR2 (N2337, N2332, N1199);
nand NAND4 (N2338, N2335, N1027, N1989, N865);
buf BUF1 (N2339, N2337);
or OR4 (N2340, N2328, N52, N1029, N393);
xor XOR2 (N2341, N2330, N1604);
not NOT1 (N2342, N2340);
nor NOR3 (N2343, N2333, N336, N838);
nor NOR3 (N2344, N2334, N2287, N2034);
nand NAND4 (N2345, N2343, N817, N1687, N1446);
nand NAND4 (N2346, N2344, N1289, N1048, N1547);
and AND3 (N2347, N2345, N934, N173);
xor XOR2 (N2348, N2326, N1161);
or OR4 (N2349, N2339, N1538, N1269, N1977);
or OR3 (N2350, N2346, N646, N375);
or OR4 (N2351, N2338, N1824, N418, N1515);
nor NOR2 (N2352, N2342, N816);
nor NOR2 (N2353, N2352, N1279);
buf BUF1 (N2354, N2348);
nand NAND3 (N2355, N2349, N1885, N1823);
nor NOR3 (N2356, N2336, N1868, N155);
nor NOR3 (N2357, N2354, N583, N101);
nand NAND4 (N2358, N2351, N619, N251, N748);
and AND3 (N2359, N2329, N1494, N103);
buf BUF1 (N2360, N2350);
nand NAND3 (N2361, N2327, N1707, N1987);
and AND4 (N2362, N2347, N597, N1575, N1991);
buf BUF1 (N2363, N2360);
and AND2 (N2364, N2355, N1747);
nand NAND3 (N2365, N2359, N839, N1279);
nand NAND4 (N2366, N2357, N2026, N146, N276);
or OR4 (N2367, N2356, N233, N1742, N1225);
or OR2 (N2368, N2367, N1028);
and AND2 (N2369, N2363, N421);
nand NAND3 (N2370, N2353, N478, N1315);
nor NOR2 (N2371, N2366, N826);
xor XOR2 (N2372, N2341, N1129);
or OR4 (N2373, N2362, N196, N1443, N2067);
buf BUF1 (N2374, N2370);
not NOT1 (N2375, N2371);
or OR3 (N2376, N2372, N1068, N310);
nor NOR4 (N2377, N2368, N1417, N141, N2013);
xor XOR2 (N2378, N2376, N565);
not NOT1 (N2379, N2373);
nor NOR2 (N2380, N2379, N368);
or OR2 (N2381, N2375, N2337);
xor XOR2 (N2382, N2377, N1151);
nand NAND4 (N2383, N2361, N1532, N160, N1702);
and AND3 (N2384, N2358, N1190, N550);
or OR4 (N2385, N2365, N823, N1115, N2064);
and AND2 (N2386, N2374, N915);
nand NAND3 (N2387, N2381, N2190, N2042);
and AND4 (N2388, N2378, N1828, N1748, N898);
nor NOR4 (N2389, N2364, N1925, N1130, N2103);
or OR2 (N2390, N2382, N1965);
nor NOR4 (N2391, N2383, N2306, N57, N848);
not NOT1 (N2392, N2387);
not NOT1 (N2393, N2385);
xor XOR2 (N2394, N2380, N452);
xor XOR2 (N2395, N2388, N634);
not NOT1 (N2396, N2393);
buf BUF1 (N2397, N2396);
or OR2 (N2398, N2394, N358);
nand NAND2 (N2399, N2395, N2299);
nor NOR2 (N2400, N2392, N1575);
xor XOR2 (N2401, N2390, N238);
not NOT1 (N2402, N2369);
or OR3 (N2403, N2400, N1892, N891);
and AND2 (N2404, N2401, N868);
and AND3 (N2405, N2397, N1071, N2323);
nand NAND2 (N2406, N2398, N1107);
buf BUF1 (N2407, N2386);
not NOT1 (N2408, N2384);
buf BUF1 (N2409, N2399);
nor NOR4 (N2410, N2406, N1807, N1315, N1196);
xor XOR2 (N2411, N2404, N1631);
nand NAND4 (N2412, N2405, N1499, N1655, N11);
xor XOR2 (N2413, N2412, N758);
not NOT1 (N2414, N2389);
not NOT1 (N2415, N2402);
nor NOR3 (N2416, N2414, N1062, N642);
nor NOR4 (N2417, N2415, N1967, N1908, N70);
xor XOR2 (N2418, N2407, N1897);
and AND2 (N2419, N2413, N1749);
nand NAND2 (N2420, N2416, N2283);
nor NOR4 (N2421, N2409, N467, N578, N1218);
xor XOR2 (N2422, N2410, N1175);
buf BUF1 (N2423, N2418);
xor XOR2 (N2424, N2391, N2068);
and AND3 (N2425, N2419, N2280, N1005);
nand NAND4 (N2426, N2411, N1385, N284, N2390);
and AND4 (N2427, N2403, N666, N2406, N1824);
or OR2 (N2428, N2424, N1273);
and AND4 (N2429, N2425, N2048, N1937, N1906);
xor XOR2 (N2430, N2427, N1147);
and AND3 (N2431, N2421, N426, N2142);
buf BUF1 (N2432, N2431);
nand NAND4 (N2433, N2432, N1502, N1178, N114);
xor XOR2 (N2434, N2429, N808);
or OR4 (N2435, N2422, N1050, N941, N2185);
nand NAND2 (N2436, N2428, N1546);
nor NOR2 (N2437, N2434, N1368);
nand NAND2 (N2438, N2408, N1252);
nand NAND4 (N2439, N2436, N1700, N2165, N1434);
nor NOR3 (N2440, N2423, N993, N2021);
nand NAND4 (N2441, N2435, N575, N1317, N1899);
nand NAND4 (N2442, N2433, N1370, N1924, N1294);
nor NOR2 (N2443, N2440, N1095);
buf BUF1 (N2444, N2426);
and AND4 (N2445, N2417, N2022, N1868, N863);
or OR3 (N2446, N2420, N15, N1227);
or OR2 (N2447, N2438, N1856);
buf BUF1 (N2448, N2446);
xor XOR2 (N2449, N2444, N164);
nand NAND3 (N2450, N2442, N155, N1251);
nand NAND2 (N2451, N2450, N1484);
or OR4 (N2452, N2447, N81, N876, N238);
nand NAND4 (N2453, N2451, N173, N1083, N2049);
and AND2 (N2454, N2453, N1034);
or OR4 (N2455, N2452, N1272, N1600, N755);
buf BUF1 (N2456, N2448);
nand NAND2 (N2457, N2441, N1968);
or OR4 (N2458, N2455, N1405, N938, N2096);
or OR3 (N2459, N2456, N2254, N2413);
and AND4 (N2460, N2458, N1925, N2165, N1911);
or OR4 (N2461, N2449, N756, N387, N1735);
nand NAND2 (N2462, N2460, N2334);
buf BUF1 (N2463, N2439);
nand NAND4 (N2464, N2463, N1545, N151, N570);
nand NAND2 (N2465, N2464, N1200);
nor NOR2 (N2466, N2461, N357);
nand NAND4 (N2467, N2445, N2461, N329, N484);
nor NOR3 (N2468, N2457, N460, N2378);
not NOT1 (N2469, N2459);
nor NOR3 (N2470, N2462, N1764, N558);
xor XOR2 (N2471, N2454, N1770);
xor XOR2 (N2472, N2465, N513);
and AND2 (N2473, N2470, N2183);
and AND3 (N2474, N2430, N1660, N2127);
nor NOR2 (N2475, N2443, N2189);
nor NOR3 (N2476, N2471, N2273, N462);
nand NAND4 (N2477, N2467, N1788, N1791, N494);
and AND2 (N2478, N2473, N2266);
nor NOR2 (N2479, N2468, N927);
buf BUF1 (N2480, N2479);
or OR4 (N2481, N2477, N202, N1778, N1550);
or OR3 (N2482, N2476, N1188, N544);
nor NOR2 (N2483, N2474, N471);
and AND3 (N2484, N2469, N1568, N50);
xor XOR2 (N2485, N2472, N1457);
or OR2 (N2486, N2478, N175);
or OR3 (N2487, N2480, N1814, N95);
xor XOR2 (N2488, N2486, N173);
buf BUF1 (N2489, N2466);
xor XOR2 (N2490, N2483, N1237);
nor NOR3 (N2491, N2481, N215, N1641);
and AND4 (N2492, N2485, N97, N384, N1832);
not NOT1 (N2493, N2482);
nor NOR4 (N2494, N2437, N1328, N2261, N1660);
buf BUF1 (N2495, N2490);
buf BUF1 (N2496, N2491);
nor NOR3 (N2497, N2489, N862, N866);
nand NAND2 (N2498, N2484, N2184);
not NOT1 (N2499, N2475);
xor XOR2 (N2500, N2495, N1742);
nor NOR2 (N2501, N2498, N518);
buf BUF1 (N2502, N2500);
buf BUF1 (N2503, N2497);
buf BUF1 (N2504, N2499);
nor NOR3 (N2505, N2501, N60, N2272);
nor NOR2 (N2506, N2502, N1896);
xor XOR2 (N2507, N2492, N2249);
or OR4 (N2508, N2493, N2401, N1634, N462);
and AND2 (N2509, N2504, N1727);
not NOT1 (N2510, N2506);
buf BUF1 (N2511, N2488);
buf BUF1 (N2512, N2507);
and AND3 (N2513, N2510, N1487, N1304);
or OR3 (N2514, N2513, N1448, N1148);
or OR4 (N2515, N2503, N1085, N2243, N1988);
nand NAND4 (N2516, N2487, N501, N1993, N2222);
not NOT1 (N2517, N2509);
nand NAND3 (N2518, N2511, N6, N1821);
xor XOR2 (N2519, N2496, N1833);
and AND4 (N2520, N2508, N361, N812, N1830);
nor NOR3 (N2521, N2518, N25, N228);
or OR4 (N2522, N2512, N1055, N1678, N169);
or OR3 (N2523, N2521, N286, N1044);
and AND3 (N2524, N2519, N176, N1439);
xor XOR2 (N2525, N2515, N658);
and AND3 (N2526, N2514, N213, N2027);
nor NOR3 (N2527, N2516, N229, N1107);
or OR4 (N2528, N2525, N366, N1999, N1041);
or OR4 (N2529, N2517, N268, N1874, N1108);
xor XOR2 (N2530, N2523, N1510);
buf BUF1 (N2531, N2522);
or OR3 (N2532, N2524, N2244, N769);
and AND2 (N2533, N2505, N1585);
not NOT1 (N2534, N2526);
nand NAND2 (N2535, N2531, N404);
nand NAND3 (N2536, N2533, N1755, N2355);
nand NAND4 (N2537, N2529, N1765, N628, N332);
and AND3 (N2538, N2535, N1734, N350);
not NOT1 (N2539, N2520);
or OR2 (N2540, N2538, N2062);
xor XOR2 (N2541, N2528, N1892);
nand NAND2 (N2542, N2541, N1288);
nand NAND3 (N2543, N2494, N1453, N969);
or OR3 (N2544, N2543, N2126, N1946);
and AND3 (N2545, N2540, N1722, N2094);
nor NOR4 (N2546, N2527, N1995, N165, N2192);
or OR2 (N2547, N2534, N716);
buf BUF1 (N2548, N2545);
and AND3 (N2549, N2547, N601, N1706);
or OR2 (N2550, N2537, N953);
not NOT1 (N2551, N2539);
xor XOR2 (N2552, N2532, N2352);
not NOT1 (N2553, N2549);
xor XOR2 (N2554, N2548, N1654);
xor XOR2 (N2555, N2530, N2178);
nor NOR4 (N2556, N2553, N1113, N661, N1469);
not NOT1 (N2557, N2552);
nor NOR2 (N2558, N2555, N608);
or OR2 (N2559, N2557, N1442);
not NOT1 (N2560, N2558);
buf BUF1 (N2561, N2554);
nand NAND3 (N2562, N2556, N1373, N1764);
buf BUF1 (N2563, N2536);
nand NAND2 (N2564, N2544, N2194);
nor NOR4 (N2565, N2546, N2437, N780, N1321);
nand NAND4 (N2566, N2551, N1529, N407, N1106);
and AND3 (N2567, N2564, N2197, N1060);
and AND2 (N2568, N2562, N238);
or OR2 (N2569, N2550, N2352);
xor XOR2 (N2570, N2565, N335);
not NOT1 (N2571, N2559);
or OR3 (N2572, N2571, N1818, N1273);
xor XOR2 (N2573, N2569, N922);
buf BUF1 (N2574, N2568);
buf BUF1 (N2575, N2566);
xor XOR2 (N2576, N2572, N2080);
buf BUF1 (N2577, N2567);
or OR3 (N2578, N2575, N2427, N869);
nor NOR3 (N2579, N2561, N1496, N1350);
nor NOR3 (N2580, N2542, N2373, N671);
or OR2 (N2581, N2580, N1453);
or OR4 (N2582, N2577, N2183, N2006, N1493);
buf BUF1 (N2583, N2573);
and AND2 (N2584, N2576, N2168);
xor XOR2 (N2585, N2560, N198);
buf BUF1 (N2586, N2578);
not NOT1 (N2587, N2570);
xor XOR2 (N2588, N2574, N176);
or OR2 (N2589, N2586, N2451);
not NOT1 (N2590, N2583);
or OR2 (N2591, N2590, N1603);
or OR4 (N2592, N2589, N1493, N2396, N930);
not NOT1 (N2593, N2587);
and AND3 (N2594, N2588, N1442, N2001);
and AND3 (N2595, N2579, N1524, N1069);
or OR2 (N2596, N2591, N829);
buf BUF1 (N2597, N2593);
xor XOR2 (N2598, N2594, N1025);
and AND2 (N2599, N2598, N1271);
xor XOR2 (N2600, N2596, N2288);
xor XOR2 (N2601, N2600, N696);
nor NOR4 (N2602, N2582, N1258, N919, N1972);
nor NOR2 (N2603, N2592, N1050);
xor XOR2 (N2604, N2599, N2193);
or OR4 (N2605, N2563, N1374, N2268, N378);
nor NOR4 (N2606, N2604, N1073, N2064, N1864);
and AND2 (N2607, N2603, N1465);
not NOT1 (N2608, N2601);
nor NOR2 (N2609, N2607, N1736);
or OR4 (N2610, N2606, N2065, N706, N477);
nor NOR2 (N2611, N2609, N1693);
buf BUF1 (N2612, N2595);
xor XOR2 (N2613, N2611, N1540);
or OR2 (N2614, N2610, N1810);
not NOT1 (N2615, N2581);
nand NAND2 (N2616, N2615, N149);
or OR2 (N2617, N2602, N1304);
and AND4 (N2618, N2613, N929, N1488, N950);
or OR3 (N2619, N2597, N1813, N150);
not NOT1 (N2620, N2612);
buf BUF1 (N2621, N2618);
nor NOR3 (N2622, N2585, N2195, N2209);
not NOT1 (N2623, N2616);
nand NAND2 (N2624, N2621, N1317);
buf BUF1 (N2625, N2605);
nor NOR3 (N2626, N2617, N2170, N1472);
nand NAND4 (N2627, N2620, N554, N1763, N209);
nor NOR3 (N2628, N2614, N211, N30);
not NOT1 (N2629, N2619);
nor NOR2 (N2630, N2624, N2459);
buf BUF1 (N2631, N2584);
and AND2 (N2632, N2628, N2532);
nor NOR2 (N2633, N2632, N975);
and AND3 (N2634, N2629, N1034, N662);
nand NAND4 (N2635, N2634, N974, N2476, N2316);
nand NAND3 (N2636, N2627, N17, N359);
not NOT1 (N2637, N2622);
not NOT1 (N2638, N2631);
buf BUF1 (N2639, N2636);
nand NAND3 (N2640, N2630, N856, N629);
or OR2 (N2641, N2638, N239);
or OR2 (N2642, N2635, N1678);
and AND3 (N2643, N2626, N469, N85);
xor XOR2 (N2644, N2608, N68);
nor NOR2 (N2645, N2643, N608);
and AND4 (N2646, N2637, N257, N918, N788);
nor NOR2 (N2647, N2646, N1795);
buf BUF1 (N2648, N2647);
not NOT1 (N2649, N2633);
and AND3 (N2650, N2623, N1427, N2229);
or OR4 (N2651, N2640, N292, N1269, N297);
xor XOR2 (N2652, N2641, N1286);
and AND2 (N2653, N2642, N1807);
not NOT1 (N2654, N2651);
or OR3 (N2655, N2653, N1853, N466);
not NOT1 (N2656, N2655);
not NOT1 (N2657, N2645);
buf BUF1 (N2658, N2644);
or OR4 (N2659, N2654, N1378, N676, N2395);
or OR4 (N2660, N2650, N1287, N1243, N2185);
or OR4 (N2661, N2656, N448, N1757, N439);
nor NOR2 (N2662, N2661, N1280);
nand NAND4 (N2663, N2639, N860, N44, N1433);
and AND4 (N2664, N2652, N306, N2479, N779);
xor XOR2 (N2665, N2658, N1713);
nand NAND3 (N2666, N2649, N1827, N909);
xor XOR2 (N2667, N2659, N679);
buf BUF1 (N2668, N2667);
nor NOR2 (N2669, N2648, N1909);
nand NAND3 (N2670, N2657, N45, N1137);
or OR2 (N2671, N2669, N412);
and AND4 (N2672, N2625, N1221, N701, N1219);
not NOT1 (N2673, N2664);
nor NOR3 (N2674, N2660, N2158, N559);
not NOT1 (N2675, N2672);
buf BUF1 (N2676, N2670);
nand NAND4 (N2677, N2674, N1624, N1250, N1487);
not NOT1 (N2678, N2665);
nand NAND3 (N2679, N2675, N2268, N1998);
nor NOR3 (N2680, N2677, N488, N1589);
or OR2 (N2681, N2662, N517);
xor XOR2 (N2682, N2681, N1115);
or OR3 (N2683, N2676, N324, N33);
buf BUF1 (N2684, N2673);
nor NOR3 (N2685, N2678, N49, N567);
and AND4 (N2686, N2671, N2508, N1622, N532);
or OR2 (N2687, N2685, N2680);
buf BUF1 (N2688, N489);
nand NAND3 (N2689, N2686, N1562, N2630);
and AND2 (N2690, N2682, N720);
and AND2 (N2691, N2690, N1556);
xor XOR2 (N2692, N2663, N287);
xor XOR2 (N2693, N2683, N2149);
nand NAND2 (N2694, N2688, N2058);
xor XOR2 (N2695, N2693, N528);
nand NAND3 (N2696, N2692, N2388, N897);
or OR3 (N2697, N2687, N2597, N2205);
not NOT1 (N2698, N2666);
nand NAND3 (N2699, N2698, N954, N1426);
nor NOR3 (N2700, N2684, N940, N1086);
and AND3 (N2701, N2694, N1118, N26);
nor NOR3 (N2702, N2699, N1765, N1241);
buf BUF1 (N2703, N2691);
and AND2 (N2704, N2701, N946);
nor NOR2 (N2705, N2668, N2333);
buf BUF1 (N2706, N2704);
or OR3 (N2707, N2689, N1305, N2401);
and AND4 (N2708, N2707, N571, N1288, N699);
or OR4 (N2709, N2705, N2355, N2163, N320);
buf BUF1 (N2710, N2696);
not NOT1 (N2711, N2708);
or OR3 (N2712, N2697, N2575, N2305);
buf BUF1 (N2713, N2710);
nor NOR4 (N2714, N2679, N765, N293, N1231);
and AND3 (N2715, N2700, N198, N2348);
and AND4 (N2716, N2706, N1275, N1018, N2684);
or OR2 (N2717, N2711, N2319);
and AND4 (N2718, N2713, N2253, N2220, N1451);
nand NAND4 (N2719, N2716, N1427, N1363, N34);
xor XOR2 (N2720, N2718, N1335);
nand NAND3 (N2721, N2695, N2480, N1747);
xor XOR2 (N2722, N2703, N362);
or OR3 (N2723, N2721, N2012, N1410);
nor NOR2 (N2724, N2719, N1588);
and AND4 (N2725, N2702, N955, N2454, N1703);
nand NAND3 (N2726, N2709, N152, N617);
or OR2 (N2727, N2726, N1305);
or OR2 (N2728, N2724, N542);
not NOT1 (N2729, N2722);
or OR3 (N2730, N2723, N1173, N850);
and AND4 (N2731, N2720, N732, N621, N488);
not NOT1 (N2732, N2727);
xor XOR2 (N2733, N2725, N2523);
and AND4 (N2734, N2728, N2391, N2407, N1000);
or OR2 (N2735, N2730, N2043);
and AND3 (N2736, N2714, N2635, N1673);
or OR4 (N2737, N2732, N535, N1041, N1670);
nand NAND4 (N2738, N2735, N42, N1712, N271);
not NOT1 (N2739, N2729);
or OR3 (N2740, N2736, N852, N2331);
nand NAND3 (N2741, N2734, N675, N939);
not NOT1 (N2742, N2733);
nand NAND3 (N2743, N2742, N287, N2254);
and AND2 (N2744, N2741, N1631);
and AND4 (N2745, N2712, N2150, N1826, N558);
or OR4 (N2746, N2743, N2574, N1217, N362);
or OR4 (N2747, N2717, N1093, N1549, N989);
nor NOR3 (N2748, N2746, N1707, N1380);
or OR2 (N2749, N2739, N1845);
nand NAND4 (N2750, N2749, N1980, N1924, N926);
not NOT1 (N2751, N2737);
not NOT1 (N2752, N2738);
xor XOR2 (N2753, N2747, N1850);
and AND3 (N2754, N2744, N2094, N2244);
nor NOR4 (N2755, N2753, N21, N2168, N399);
and AND4 (N2756, N2731, N2740, N50, N2048);
nand NAND2 (N2757, N334, N2450);
nor NOR3 (N2758, N2752, N31, N1930);
nor NOR4 (N2759, N2745, N1721, N2702, N1094);
nor NOR3 (N2760, N2759, N1832, N1424);
xor XOR2 (N2761, N2760, N1801);
buf BUF1 (N2762, N2757);
not NOT1 (N2763, N2750);
nor NOR3 (N2764, N2762, N1721, N2432);
not NOT1 (N2765, N2763);
nor NOR2 (N2766, N2758, N1227);
buf BUF1 (N2767, N2765);
and AND4 (N2768, N2756, N290, N1978, N1776);
nor NOR3 (N2769, N2754, N2265, N1407);
nor NOR3 (N2770, N2751, N1558, N744);
and AND2 (N2771, N2748, N1253);
or OR2 (N2772, N2771, N411);
not NOT1 (N2773, N2772);
not NOT1 (N2774, N2773);
nand NAND2 (N2775, N2769, N2424);
or OR3 (N2776, N2768, N718, N1467);
buf BUF1 (N2777, N2766);
xor XOR2 (N2778, N2764, N969);
not NOT1 (N2779, N2770);
xor XOR2 (N2780, N2715, N588);
nand NAND3 (N2781, N2767, N427, N842);
xor XOR2 (N2782, N2778, N26);
xor XOR2 (N2783, N2781, N963);
or OR4 (N2784, N2782, N623, N2353, N1075);
not NOT1 (N2785, N2783);
or OR3 (N2786, N2784, N1410, N1173);
and AND3 (N2787, N2785, N2536, N909);
buf BUF1 (N2788, N2777);
xor XOR2 (N2789, N2779, N80);
buf BUF1 (N2790, N2786);
xor XOR2 (N2791, N2775, N1041);
xor XOR2 (N2792, N2776, N1324);
nor NOR3 (N2793, N2755, N2503, N130);
buf BUF1 (N2794, N2793);
nand NAND2 (N2795, N2794, N167);
nand NAND3 (N2796, N2780, N469, N1624);
buf BUF1 (N2797, N2790);
and AND3 (N2798, N2761, N2642, N1366);
or OR3 (N2799, N2797, N959, N2133);
not NOT1 (N2800, N2789);
or OR3 (N2801, N2792, N2087, N2137);
nand NAND4 (N2802, N2801, N636, N1517, N1520);
not NOT1 (N2803, N2788);
not NOT1 (N2804, N2802);
buf BUF1 (N2805, N2800);
nor NOR3 (N2806, N2795, N1414, N813);
xor XOR2 (N2807, N2774, N711);
buf BUF1 (N2808, N2804);
buf BUF1 (N2809, N2796);
or OR2 (N2810, N2809, N2404);
or OR4 (N2811, N2799, N2622, N177, N583);
not NOT1 (N2812, N2805);
xor XOR2 (N2813, N2791, N300);
xor XOR2 (N2814, N2807, N974);
xor XOR2 (N2815, N2806, N977);
not NOT1 (N2816, N2803);
or OR2 (N2817, N2816, N826);
nand NAND4 (N2818, N2813, N28, N2256, N1201);
nand NAND3 (N2819, N2812, N1072, N1245);
nor NOR2 (N2820, N2815, N1436);
xor XOR2 (N2821, N2814, N1045);
or OR3 (N2822, N2819, N590, N2102);
buf BUF1 (N2823, N2787);
nand NAND2 (N2824, N2808, N2237);
buf BUF1 (N2825, N2821);
not NOT1 (N2826, N2820);
buf BUF1 (N2827, N2824);
not NOT1 (N2828, N2823);
nor NOR4 (N2829, N2817, N1899, N1727, N1238);
buf BUF1 (N2830, N2818);
nor NOR3 (N2831, N2810, N1639, N1245);
not NOT1 (N2832, N2822);
xor XOR2 (N2833, N2827, N1187);
nor NOR2 (N2834, N2825, N2551);
nand NAND3 (N2835, N2830, N1160, N1939);
nor NOR3 (N2836, N2811, N1357, N1093);
and AND4 (N2837, N2834, N672, N1244, N2712);
nand NAND3 (N2838, N2836, N2549, N1183);
or OR4 (N2839, N2837, N2318, N1191, N160);
xor XOR2 (N2840, N2829, N504);
not NOT1 (N2841, N2833);
and AND3 (N2842, N2841, N32, N2197);
nand NAND4 (N2843, N2840, N336, N481, N2252);
xor XOR2 (N2844, N2842, N2210);
and AND4 (N2845, N2839, N2831, N1333, N184);
or OR4 (N2846, N1338, N2441, N2490, N2);
and AND4 (N2847, N2835, N2214, N34, N2187);
or OR2 (N2848, N2846, N320);
and AND2 (N2849, N2845, N690);
xor XOR2 (N2850, N2844, N634);
or OR2 (N2851, N2832, N2500);
not NOT1 (N2852, N2826);
buf BUF1 (N2853, N2843);
nor NOR2 (N2854, N2853, N1448);
xor XOR2 (N2855, N2847, N625);
not NOT1 (N2856, N2848);
nand NAND3 (N2857, N2855, N253, N1536);
or OR4 (N2858, N2857, N2074, N2129, N2450);
and AND4 (N2859, N2828, N2416, N402, N1147);
nor NOR4 (N2860, N2851, N187, N600, N1591);
and AND2 (N2861, N2852, N2635);
buf BUF1 (N2862, N2854);
and AND4 (N2863, N2861, N1225, N770, N2623);
and AND4 (N2864, N2859, N725, N2486, N75);
buf BUF1 (N2865, N2798);
not NOT1 (N2866, N2849);
and AND2 (N2867, N2858, N638);
buf BUF1 (N2868, N2866);
buf BUF1 (N2869, N2860);
or OR4 (N2870, N2838, N951, N573, N2008);
buf BUF1 (N2871, N2864);
nor NOR3 (N2872, N2869, N1781, N340);
or OR2 (N2873, N2863, N1719);
nand NAND3 (N2874, N2873, N316, N2765);
or OR4 (N2875, N2865, N897, N860, N302);
and AND4 (N2876, N2856, N1749, N267, N1712);
buf BUF1 (N2877, N2850);
not NOT1 (N2878, N2867);
and AND4 (N2879, N2868, N1991, N1131, N1070);
buf BUF1 (N2880, N2870);
nor NOR4 (N2881, N2876, N1332, N6, N843);
xor XOR2 (N2882, N2880, N589);
nand NAND3 (N2883, N2871, N2775, N2607);
buf BUF1 (N2884, N2862);
not NOT1 (N2885, N2878);
nor NOR2 (N2886, N2881, N1572);
or OR4 (N2887, N2879, N1797, N519, N2034);
not NOT1 (N2888, N2886);
xor XOR2 (N2889, N2885, N755);
and AND2 (N2890, N2884, N989);
and AND4 (N2891, N2875, N2807, N2744, N297);
not NOT1 (N2892, N2888);
nand NAND3 (N2893, N2883, N1385, N270);
not NOT1 (N2894, N2893);
nand NAND4 (N2895, N2894, N759, N2604, N1799);
or OR3 (N2896, N2892, N43, N645);
and AND2 (N2897, N2882, N2534);
not NOT1 (N2898, N2872);
nor NOR2 (N2899, N2874, N309);
not NOT1 (N2900, N2877);
xor XOR2 (N2901, N2899, N740);
buf BUF1 (N2902, N2887);
or OR4 (N2903, N2896, N665, N2111, N1939);
or OR4 (N2904, N2903, N233, N1988, N1311);
and AND3 (N2905, N2901, N166, N502);
nand NAND3 (N2906, N2895, N2363, N2740);
xor XOR2 (N2907, N2906, N2869);
and AND2 (N2908, N2904, N1679);
xor XOR2 (N2909, N2891, N1950);
buf BUF1 (N2910, N2897);
not NOT1 (N2911, N2909);
or OR2 (N2912, N2908, N2158);
not NOT1 (N2913, N2911);
not NOT1 (N2914, N2905);
and AND4 (N2915, N2898, N726, N2335, N446);
and AND2 (N2916, N2912, N1841);
or OR4 (N2917, N2913, N2736, N929, N2839);
and AND2 (N2918, N2916, N1950);
xor XOR2 (N2919, N2917, N2272);
xor XOR2 (N2920, N2889, N1126);
or OR4 (N2921, N2890, N1406, N1, N635);
not NOT1 (N2922, N2900);
and AND3 (N2923, N2914, N1063, N585);
nand NAND3 (N2924, N2923, N2540, N2208);
xor XOR2 (N2925, N2918, N1897);
and AND4 (N2926, N2925, N1193, N733, N2112);
nor NOR2 (N2927, N2920, N272);
xor XOR2 (N2928, N2915, N445);
and AND4 (N2929, N2919, N384, N1918, N2315);
nor NOR2 (N2930, N2902, N2898);
nor NOR3 (N2931, N2930, N2905, N2221);
nand NAND3 (N2932, N2929, N2840, N62);
not NOT1 (N2933, N2921);
nand NAND3 (N2934, N2932, N1455, N1337);
not NOT1 (N2935, N2924);
buf BUF1 (N2936, N2910);
and AND3 (N2937, N2926, N217, N475);
not NOT1 (N2938, N2907);
nor NOR4 (N2939, N2934, N1967, N927, N950);
buf BUF1 (N2940, N2939);
nand NAND3 (N2941, N2928, N1802, N1472);
not NOT1 (N2942, N2935);
xor XOR2 (N2943, N2931, N2901);
and AND2 (N2944, N2922, N1695);
xor XOR2 (N2945, N2936, N2576);
not NOT1 (N2946, N2933);
and AND4 (N2947, N2937, N7, N460, N1230);
and AND2 (N2948, N2943, N2404);
buf BUF1 (N2949, N2944);
or OR2 (N2950, N2940, N2511);
nand NAND4 (N2951, N2947, N98, N2048, N263);
buf BUF1 (N2952, N2942);
xor XOR2 (N2953, N2941, N2148);
and AND3 (N2954, N2927, N1346, N402);
not NOT1 (N2955, N2950);
nor NOR3 (N2956, N2945, N1112, N1440);
xor XOR2 (N2957, N2951, N2775);
nor NOR4 (N2958, N2946, N2102, N2545, N2052);
nand NAND3 (N2959, N2957, N1076, N1293);
buf BUF1 (N2960, N2953);
nor NOR4 (N2961, N2949, N2618, N6, N1702);
xor XOR2 (N2962, N2961, N1015);
and AND4 (N2963, N2955, N663, N538, N866);
buf BUF1 (N2964, N2956);
buf BUF1 (N2965, N2958);
xor XOR2 (N2966, N2938, N2849);
and AND2 (N2967, N2966, N507);
not NOT1 (N2968, N2963);
xor XOR2 (N2969, N2965, N1497);
and AND3 (N2970, N2948, N246, N2423);
xor XOR2 (N2971, N2954, N1463);
xor XOR2 (N2972, N2971, N1413);
not NOT1 (N2973, N2970);
not NOT1 (N2974, N2967);
buf BUF1 (N2975, N2962);
not NOT1 (N2976, N2974);
buf BUF1 (N2977, N2976);
and AND3 (N2978, N2973, N1300, N310);
and AND2 (N2979, N2978, N662);
nor NOR4 (N2980, N2969, N1310, N1646, N752);
and AND4 (N2981, N2959, N1429, N1202, N1003);
and AND4 (N2982, N2980, N1795, N1207, N1622);
not NOT1 (N2983, N2968);
nor NOR4 (N2984, N2982, N303, N2864, N2223);
and AND4 (N2985, N2972, N2924, N1171, N2101);
nor NOR2 (N2986, N2979, N2979);
or OR3 (N2987, N2960, N2664, N650);
or OR4 (N2988, N2975, N1922, N486, N2825);
not NOT1 (N2989, N2985);
xor XOR2 (N2990, N2988, N1400);
nor NOR2 (N2991, N2952, N2910);
nor NOR3 (N2992, N2984, N1501, N955);
and AND2 (N2993, N2977, N2321);
xor XOR2 (N2994, N2990, N10);
nor NOR4 (N2995, N2983, N2759, N1121, N495);
not NOT1 (N2996, N2994);
buf BUF1 (N2997, N2987);
or OR2 (N2998, N2986, N561);
not NOT1 (N2999, N2996);
and AND2 (N3000, N2993, N539);
not NOT1 (N3001, N2964);
buf BUF1 (N3002, N2992);
buf BUF1 (N3003, N2998);
nand NAND4 (N3004, N3003, N694, N1505, N2983);
buf BUF1 (N3005, N2981);
or OR4 (N3006, N2991, N2406, N1738, N359);
buf BUF1 (N3007, N3004);
buf BUF1 (N3008, N3005);
or OR3 (N3009, N2997, N382, N2318);
buf BUF1 (N3010, N3008);
or OR2 (N3011, N2995, N1228);
nor NOR2 (N3012, N3002, N686);
nand NAND3 (N3013, N3011, N2126, N1626);
buf BUF1 (N3014, N3007);
xor XOR2 (N3015, N3014, N2561);
buf BUF1 (N3016, N3009);
buf BUF1 (N3017, N3015);
xor XOR2 (N3018, N3000, N1399);
buf BUF1 (N3019, N3013);
buf BUF1 (N3020, N2999);
nand NAND3 (N3021, N3012, N1963, N1798);
xor XOR2 (N3022, N3017, N1873);
or OR3 (N3023, N3018, N309, N632);
xor XOR2 (N3024, N3021, N2140);
and AND2 (N3025, N3024, N38);
nand NAND3 (N3026, N3022, N2480, N747);
xor XOR2 (N3027, N3006, N2889);
nand NAND2 (N3028, N3023, N2608);
xor XOR2 (N3029, N3016, N1198);
nand NAND4 (N3030, N3019, N219, N2590, N2264);
buf BUF1 (N3031, N3026);
not NOT1 (N3032, N3025);
not NOT1 (N3033, N3027);
or OR3 (N3034, N3029, N195, N2823);
nor NOR3 (N3035, N3020, N1817, N365);
not NOT1 (N3036, N3001);
xor XOR2 (N3037, N3030, N1540);
not NOT1 (N3038, N3035);
not NOT1 (N3039, N3033);
nor NOR3 (N3040, N3010, N149, N81);
not NOT1 (N3041, N3032);
and AND2 (N3042, N3041, N1864);
or OR2 (N3043, N3031, N839);
or OR3 (N3044, N3039, N1353, N1170);
and AND3 (N3045, N3038, N10, N2192);
not NOT1 (N3046, N3040);
nor NOR2 (N3047, N3042, N1686);
and AND3 (N3048, N3036, N736, N1706);
or OR2 (N3049, N3034, N1479);
not NOT1 (N3050, N2989);
nand NAND2 (N3051, N3046, N824);
nor NOR3 (N3052, N3028, N2644, N2244);
nand NAND4 (N3053, N3052, N884, N1650, N394);
not NOT1 (N3054, N3049);
buf BUF1 (N3055, N3048);
xor XOR2 (N3056, N3055, N2099);
not NOT1 (N3057, N3051);
xor XOR2 (N3058, N3057, N1903);
not NOT1 (N3059, N3056);
xor XOR2 (N3060, N3044, N2574);
nor NOR4 (N3061, N3050, N1439, N865, N988);
or OR2 (N3062, N3060, N994);
or OR3 (N3063, N3061, N551, N290);
xor XOR2 (N3064, N3047, N1368);
nand NAND3 (N3065, N3058, N24, N1016);
xor XOR2 (N3066, N3062, N373);
not NOT1 (N3067, N3053);
or OR2 (N3068, N3037, N802);
nor NOR4 (N3069, N3067, N2272, N622, N2786);
or OR3 (N3070, N3069, N1422, N349);
buf BUF1 (N3071, N3059);
and AND4 (N3072, N3065, N1215, N2415, N1435);
or OR4 (N3073, N3071, N1758, N2064, N1226);
not NOT1 (N3074, N3045);
and AND4 (N3075, N3068, N1820, N2024, N2321);
and AND3 (N3076, N3066, N1808, N330);
and AND3 (N3077, N3074, N139, N2563);
nor NOR2 (N3078, N3077, N2819);
buf BUF1 (N3079, N3075);
and AND2 (N3080, N3078, N2292);
nand NAND4 (N3081, N3064, N3073, N2112, N167);
nand NAND3 (N3082, N666, N763, N1394);
nand NAND4 (N3083, N3079, N1093, N1098, N2520);
nand NAND4 (N3084, N3043, N546, N2436, N1515);
not NOT1 (N3085, N3083);
nand NAND2 (N3086, N3084, N875);
not NOT1 (N3087, N3076);
buf BUF1 (N3088, N3086);
not NOT1 (N3089, N3054);
or OR2 (N3090, N3063, N1407);
not NOT1 (N3091, N3082);
xor XOR2 (N3092, N3090, N171);
not NOT1 (N3093, N3085);
nand NAND4 (N3094, N3070, N907, N466, N70);
nand NAND4 (N3095, N3092, N1061, N812, N30);
xor XOR2 (N3096, N3080, N1215);
nand NAND3 (N3097, N3095, N1088, N2992);
nor NOR2 (N3098, N3087, N696);
nor NOR2 (N3099, N3094, N1648);
buf BUF1 (N3100, N3089);
buf BUF1 (N3101, N3098);
and AND2 (N3102, N3072, N3025);
nor NOR4 (N3103, N3093, N2228, N1306, N2533);
and AND2 (N3104, N3100, N79);
xor XOR2 (N3105, N3081, N1202);
not NOT1 (N3106, N3103);
xor XOR2 (N3107, N3104, N42);
buf BUF1 (N3108, N3097);
not NOT1 (N3109, N3101);
nor NOR2 (N3110, N3109, N2991);
not NOT1 (N3111, N3099);
or OR3 (N3112, N3091, N2771, N2309);
xor XOR2 (N3113, N3108, N1443);
nand NAND4 (N3114, N3113, N2079, N2187, N424);
nor NOR4 (N3115, N3105, N1716, N2412, N604);
nor NOR3 (N3116, N3088, N1859, N2286);
and AND3 (N3117, N3114, N2237, N2964);
buf BUF1 (N3118, N3110);
nor NOR4 (N3119, N3118, N1533, N1214, N1301);
and AND4 (N3120, N3106, N1568, N1232, N335);
xor XOR2 (N3121, N3117, N2593);
buf BUF1 (N3122, N3119);
nor NOR4 (N3123, N3120, N2073, N1634, N2490);
nor NOR2 (N3124, N3112, N875);
not NOT1 (N3125, N3111);
nand NAND2 (N3126, N3121, N421);
xor XOR2 (N3127, N3125, N2588);
nor NOR3 (N3128, N3123, N539, N1353);
and AND3 (N3129, N3128, N2111, N1908);
nand NAND3 (N3130, N3126, N2474, N312);
nor NOR2 (N3131, N3115, N872);
not NOT1 (N3132, N3096);
xor XOR2 (N3133, N3107, N529);
not NOT1 (N3134, N3127);
nand NAND4 (N3135, N3102, N1500, N219, N1403);
nand NAND2 (N3136, N3129, N1084);
xor XOR2 (N3137, N3135, N622);
xor XOR2 (N3138, N3136, N72);
and AND2 (N3139, N3116, N2307);
nand NAND4 (N3140, N3134, N2963, N1630, N2670);
nand NAND2 (N3141, N3138, N2982);
buf BUF1 (N3142, N3132);
nor NOR3 (N3143, N3139, N225, N753);
nor NOR2 (N3144, N3124, N3054);
buf BUF1 (N3145, N3131);
xor XOR2 (N3146, N3133, N2812);
nand NAND2 (N3147, N3143, N2346);
xor XOR2 (N3148, N3122, N2561);
nand NAND3 (N3149, N3137, N1827, N486);
nand NAND2 (N3150, N3147, N522);
nor NOR3 (N3151, N3140, N2188, N2837);
buf BUF1 (N3152, N3144);
buf BUF1 (N3153, N3146);
and AND4 (N3154, N3142, N2072, N1041, N991);
or OR2 (N3155, N3148, N747);
or OR2 (N3156, N3153, N1221);
nor NOR3 (N3157, N3149, N2788, N2215);
nand NAND3 (N3158, N3145, N968, N2235);
or OR2 (N3159, N3141, N2550);
and AND2 (N3160, N3156, N1536);
xor XOR2 (N3161, N3155, N2774);
nor NOR2 (N3162, N3160, N36);
buf BUF1 (N3163, N3161);
buf BUF1 (N3164, N3159);
nand NAND2 (N3165, N3150, N2462);
nor NOR2 (N3166, N3154, N1514);
or OR4 (N3167, N3164, N1791, N2703, N1763);
nor NOR2 (N3168, N3163, N799);
nand NAND4 (N3169, N3158, N921, N1099, N1860);
or OR4 (N3170, N3166, N799, N276, N180);
nand NAND3 (N3171, N3167, N2670, N1557);
nand NAND3 (N3172, N3152, N2412, N2121);
nor NOR4 (N3173, N3157, N109, N2333, N75);
not NOT1 (N3174, N3130);
not NOT1 (N3175, N3171);
xor XOR2 (N3176, N3170, N825);
and AND2 (N3177, N3169, N35);
and AND4 (N3178, N3177, N1301, N2526, N1855);
buf BUF1 (N3179, N3172);
nand NAND3 (N3180, N3165, N1697, N2326);
not NOT1 (N3181, N3179);
xor XOR2 (N3182, N3174, N1649);
nor NOR4 (N3183, N3168, N898, N817, N1663);
nor NOR3 (N3184, N3176, N895, N853);
xor XOR2 (N3185, N3182, N2238);
or OR4 (N3186, N3183, N2675, N2701, N2319);
buf BUF1 (N3187, N3173);
xor XOR2 (N3188, N3181, N1270);
not NOT1 (N3189, N3162);
xor XOR2 (N3190, N3184, N1347);
not NOT1 (N3191, N3189);
xor XOR2 (N3192, N3178, N936);
nor NOR4 (N3193, N3188, N864, N1845, N1749);
and AND4 (N3194, N3187, N950, N2762, N2854);
or OR2 (N3195, N3191, N2505);
buf BUF1 (N3196, N3192);
buf BUF1 (N3197, N3180);
and AND4 (N3198, N3193, N414, N2397, N1645);
and AND2 (N3199, N3196, N451);
nor NOR3 (N3200, N3185, N457, N2255);
xor XOR2 (N3201, N3194, N144);
not NOT1 (N3202, N3190);
nor NOR2 (N3203, N3198, N2416);
buf BUF1 (N3204, N3186);
xor XOR2 (N3205, N3201, N2971);
nor NOR2 (N3206, N3151, N760);
nand NAND4 (N3207, N3202, N1492, N833, N1375);
and AND4 (N3208, N3204, N676, N277, N2288);
xor XOR2 (N3209, N3203, N179);
or OR4 (N3210, N3200, N1429, N2611, N2652);
and AND2 (N3211, N3207, N2256);
or OR2 (N3212, N3205, N380);
nand NAND2 (N3213, N3197, N3035);
buf BUF1 (N3214, N3208);
not NOT1 (N3215, N3214);
nand NAND2 (N3216, N3211, N1431);
buf BUF1 (N3217, N3216);
nand NAND2 (N3218, N3175, N2435);
not NOT1 (N3219, N3217);
xor XOR2 (N3220, N3199, N439);
buf BUF1 (N3221, N3218);
nand NAND4 (N3222, N3195, N1999, N935, N2822);
buf BUF1 (N3223, N3206);
and AND2 (N3224, N3222, N1084);
xor XOR2 (N3225, N3223, N2545);
nand NAND4 (N3226, N3225, N1899, N2920, N785);
nor NOR2 (N3227, N3221, N898);
buf BUF1 (N3228, N3210);
nand NAND2 (N3229, N3213, N226);
xor XOR2 (N3230, N3212, N2595);
and AND2 (N3231, N3230, N678);
not NOT1 (N3232, N3215);
nor NOR4 (N3233, N3231, N616, N1448, N1118);
and AND4 (N3234, N3229, N1209, N2053, N2063);
nor NOR2 (N3235, N3232, N1004);
xor XOR2 (N3236, N3235, N768);
xor XOR2 (N3237, N3227, N1378);
nor NOR4 (N3238, N3228, N2190, N2465, N1077);
nor NOR4 (N3239, N3234, N456, N2437, N2099);
not NOT1 (N3240, N3239);
xor XOR2 (N3241, N3240, N2824);
nand NAND4 (N3242, N3224, N1580, N311, N1760);
nor NOR4 (N3243, N3220, N2210, N970, N914);
xor XOR2 (N3244, N3241, N1434);
not NOT1 (N3245, N3209);
nor NOR4 (N3246, N3233, N2739, N2530, N1498);
buf BUF1 (N3247, N3236);
nand NAND3 (N3248, N3226, N114, N2955);
not NOT1 (N3249, N3248);
nor NOR4 (N3250, N3249, N15, N1203, N3104);
nor NOR2 (N3251, N3245, N2658);
nor NOR3 (N3252, N3246, N2556, N2327);
or OR4 (N3253, N3247, N400, N1256, N2250);
xor XOR2 (N3254, N3244, N2716);
buf BUF1 (N3255, N3238);
buf BUF1 (N3256, N3254);
buf BUF1 (N3257, N3237);
nand NAND2 (N3258, N3257, N2623);
xor XOR2 (N3259, N3250, N2832);
or OR4 (N3260, N3258, N2082, N2208, N1402);
buf BUF1 (N3261, N3256);
not NOT1 (N3262, N3242);
nand NAND3 (N3263, N3262, N263, N2512);
nor NOR4 (N3264, N3252, N1467, N2720, N3037);
buf BUF1 (N3265, N3259);
or OR4 (N3266, N3261, N2806, N1888, N918);
and AND3 (N3267, N3264, N1121, N945);
not NOT1 (N3268, N3260);
or OR4 (N3269, N3251, N1081, N2515, N3009);
not NOT1 (N3270, N3253);
nand NAND4 (N3271, N3268, N1013, N2906, N177);
nand NAND2 (N3272, N3269, N240);
or OR2 (N3273, N3255, N2873);
and AND4 (N3274, N3266, N562, N3226, N2737);
not NOT1 (N3275, N3243);
nor NOR4 (N3276, N3219, N3168, N1999, N996);
buf BUF1 (N3277, N3265);
nand NAND2 (N3278, N3276, N3146);
xor XOR2 (N3279, N3275, N2666);
or OR4 (N3280, N3273, N2296, N3201, N3188);
nor NOR3 (N3281, N3278, N1123, N2679);
not NOT1 (N3282, N3277);
xor XOR2 (N3283, N3274, N1900);
nor NOR3 (N3284, N3283, N453, N166);
not NOT1 (N3285, N3263);
nor NOR3 (N3286, N3267, N744, N1816);
xor XOR2 (N3287, N3270, N744);
not NOT1 (N3288, N3284);
or OR3 (N3289, N3288, N1146, N2157);
nor NOR3 (N3290, N3279, N941, N1407);
or OR4 (N3291, N3289, N2621, N1027, N2815);
nand NAND4 (N3292, N3291, N2776, N278, N1842);
or OR2 (N3293, N3292, N1585);
nand NAND3 (N3294, N3285, N305, N118);
xor XOR2 (N3295, N3286, N1881);
nand NAND3 (N3296, N3280, N1782, N2237);
nand NAND3 (N3297, N3294, N1891, N2051);
buf BUF1 (N3298, N3295);
nand NAND4 (N3299, N3290, N3173, N3204, N1704);
not NOT1 (N3300, N3297);
or OR3 (N3301, N3272, N3164, N876);
or OR3 (N3302, N3301, N2520, N166);
not NOT1 (N3303, N3302);
xor XOR2 (N3304, N3293, N1625);
nand NAND3 (N3305, N3298, N1710, N2604);
xor XOR2 (N3306, N3282, N1386);
not NOT1 (N3307, N3299);
or OR4 (N3308, N3307, N1318, N546, N2);
xor XOR2 (N3309, N3287, N303);
xor XOR2 (N3310, N3281, N768);
and AND4 (N3311, N3304, N1864, N3073, N2803);
and AND3 (N3312, N3296, N3250, N1228);
nand NAND4 (N3313, N3308, N1523, N1243, N3003);
nor NOR3 (N3314, N3303, N861, N2166);
not NOT1 (N3315, N3314);
and AND2 (N3316, N3309, N2661);
buf BUF1 (N3317, N3306);
xor XOR2 (N3318, N3271, N1899);
nand NAND3 (N3319, N3318, N546, N126);
and AND2 (N3320, N3315, N1105);
not NOT1 (N3321, N3300);
not NOT1 (N3322, N3321);
xor XOR2 (N3323, N3305, N1411);
xor XOR2 (N3324, N3310, N1331);
nor NOR3 (N3325, N3319, N2205, N1616);
nor NOR3 (N3326, N3317, N175, N1483);
nor NOR3 (N3327, N3320, N2129, N3042);
buf BUF1 (N3328, N3324);
xor XOR2 (N3329, N3328, N1080);
xor XOR2 (N3330, N3327, N19);
and AND3 (N3331, N3325, N1307, N3131);
nand NAND2 (N3332, N3311, N1889);
xor XOR2 (N3333, N3316, N2246);
nand NAND3 (N3334, N3312, N1130, N482);
nor NOR3 (N3335, N3330, N1539, N586);
and AND4 (N3336, N3332, N379, N2691, N271);
or OR4 (N3337, N3326, N2729, N3248, N1578);
nand NAND2 (N3338, N3336, N131);
nand NAND3 (N3339, N3338, N609, N1403);
and AND2 (N3340, N3323, N311);
nor NOR2 (N3341, N3334, N42);
not NOT1 (N3342, N3333);
buf BUF1 (N3343, N3322);
nor NOR2 (N3344, N3329, N2915);
nand NAND2 (N3345, N3313, N972);
not NOT1 (N3346, N3344);
not NOT1 (N3347, N3340);
nor NOR3 (N3348, N3342, N2425, N1101);
and AND2 (N3349, N3348, N1134);
or OR2 (N3350, N3339, N1577);
nor NOR3 (N3351, N3331, N2360, N1080);
or OR3 (N3352, N3337, N2186, N2502);
nor NOR3 (N3353, N3350, N1848, N1663);
xor XOR2 (N3354, N3353, N880);
nand NAND4 (N3355, N3352, N3121, N37, N52);
nand NAND4 (N3356, N3351, N508, N674, N841);
and AND4 (N3357, N3341, N2401, N2652, N2259);
nor NOR4 (N3358, N3355, N1618, N450, N1592);
or OR2 (N3359, N3346, N3133);
nor NOR2 (N3360, N3349, N813);
nand NAND4 (N3361, N3335, N1067, N1371, N251);
and AND3 (N3362, N3345, N1187, N3101);
nor NOR2 (N3363, N3347, N2077);
buf BUF1 (N3364, N3361);
nor NOR2 (N3365, N3354, N566);
or OR4 (N3366, N3360, N2318, N472, N1894);
xor XOR2 (N3367, N3363, N884);
nor NOR4 (N3368, N3367, N2907, N2676, N1228);
or OR4 (N3369, N3357, N319, N2375, N1009);
buf BUF1 (N3370, N3368);
not NOT1 (N3371, N3362);
xor XOR2 (N3372, N3358, N259);
or OR2 (N3373, N3369, N1900);
buf BUF1 (N3374, N3359);
not NOT1 (N3375, N3370);
xor XOR2 (N3376, N3375, N1028);
or OR4 (N3377, N3364, N1954, N2800, N466);
nor NOR3 (N3378, N3343, N1929, N1836);
and AND4 (N3379, N3374, N3220, N1944, N2949);
not NOT1 (N3380, N3376);
nor NOR2 (N3381, N3379, N1211);
not NOT1 (N3382, N3365);
nor NOR2 (N3383, N3356, N2582);
xor XOR2 (N3384, N3381, N1516);
nor NOR4 (N3385, N3377, N2772, N2987, N52);
not NOT1 (N3386, N3385);
or OR3 (N3387, N3366, N2926, N3012);
nor NOR2 (N3388, N3387, N3236);
or OR4 (N3389, N3378, N2829, N1966, N1537);
or OR4 (N3390, N3382, N1631, N2821, N877);
not NOT1 (N3391, N3372);
not NOT1 (N3392, N3371);
nand NAND2 (N3393, N3391, N2524);
not NOT1 (N3394, N3392);
not NOT1 (N3395, N3389);
or OR4 (N3396, N3390, N645, N3261, N2336);
buf BUF1 (N3397, N3388);
xor XOR2 (N3398, N3384, N343);
nor NOR2 (N3399, N3383, N2764);
xor XOR2 (N3400, N3397, N695);
nand NAND4 (N3401, N3380, N1514, N2079, N1899);
nor NOR3 (N3402, N3386, N1826, N554);
not NOT1 (N3403, N3399);
buf BUF1 (N3404, N3396);
nand NAND3 (N3405, N3404, N1530, N2482);
not NOT1 (N3406, N3403);
not NOT1 (N3407, N3394);
xor XOR2 (N3408, N3402, N2868);
buf BUF1 (N3409, N3406);
nand NAND3 (N3410, N3401, N3111, N1165);
or OR2 (N3411, N3410, N2292);
xor XOR2 (N3412, N3400, N2815);
buf BUF1 (N3413, N3412);
nor NOR4 (N3414, N3408, N1936, N552, N3012);
buf BUF1 (N3415, N3393);
not NOT1 (N3416, N3414);
xor XOR2 (N3417, N3407, N2544);
nand NAND4 (N3418, N3373, N3332, N3240, N2408);
and AND4 (N3419, N3417, N2256, N2128, N1222);
and AND2 (N3420, N3416, N1672);
xor XOR2 (N3421, N3419, N1628);
buf BUF1 (N3422, N3405);
buf BUF1 (N3423, N3398);
nor NOR2 (N3424, N3395, N1289);
nand NAND2 (N3425, N3423, N33);
or OR2 (N3426, N3420, N1584);
nand NAND4 (N3427, N3426, N1458, N2989, N1530);
buf BUF1 (N3428, N3418);
buf BUF1 (N3429, N3422);
nor NOR3 (N3430, N3415, N109, N65);
nor NOR4 (N3431, N3425, N470, N1000, N1174);
nor NOR3 (N3432, N3429, N132, N2835);
xor XOR2 (N3433, N3424, N1042);
xor XOR2 (N3434, N3409, N2614);
nand NAND3 (N3435, N3430, N2339, N1235);
xor XOR2 (N3436, N3413, N3178);
nand NAND4 (N3437, N3434, N1622, N2063, N2731);
and AND2 (N3438, N3431, N151);
or OR4 (N3439, N3437, N2288, N2585, N1630);
and AND3 (N3440, N3435, N2563, N2259);
buf BUF1 (N3441, N3428);
and AND3 (N3442, N3436, N1315, N816);
nor NOR4 (N3443, N3439, N3351, N168, N2191);
not NOT1 (N3444, N3441);
nand NAND2 (N3445, N3442, N2943);
and AND4 (N3446, N3438, N2546, N2840, N2800);
nor NOR4 (N3447, N3446, N1392, N1357, N1691);
and AND3 (N3448, N3443, N2743, N3447);
not NOT1 (N3449, N1056);
buf BUF1 (N3450, N3411);
buf BUF1 (N3451, N3449);
or OR3 (N3452, N3448, N1648, N1151);
xor XOR2 (N3453, N3440, N818);
nor NOR2 (N3454, N3453, N118);
nand NAND3 (N3455, N3427, N904, N3063);
nor NOR4 (N3456, N3444, N1251, N2866, N2989);
buf BUF1 (N3457, N3456);
buf BUF1 (N3458, N3454);
and AND4 (N3459, N3421, N1366, N2613, N1226);
not NOT1 (N3460, N3450);
buf BUF1 (N3461, N3460);
or OR2 (N3462, N3451, N955);
not NOT1 (N3463, N3433);
or OR3 (N3464, N3458, N1530, N2319);
and AND4 (N3465, N3463, N3393, N464, N884);
and AND3 (N3466, N3432, N602, N2161);
nand NAND3 (N3467, N3464, N2415, N2501);
and AND2 (N3468, N3455, N1902);
or OR3 (N3469, N3468, N206, N470);
nand NAND2 (N3470, N3461, N2671);
nor NOR4 (N3471, N3469, N3253, N2932, N2047);
nor NOR2 (N3472, N3465, N803);
not NOT1 (N3473, N3471);
not NOT1 (N3474, N3470);
and AND2 (N3475, N3459, N2810);
nand NAND3 (N3476, N3445, N925, N2604);
and AND2 (N3477, N3466, N379);
nor NOR4 (N3478, N3474, N3406, N1310, N2066);
xor XOR2 (N3479, N3472, N3466);
buf BUF1 (N3480, N3452);
not NOT1 (N3481, N3467);
or OR3 (N3482, N3475, N352, N1416);
xor XOR2 (N3483, N3476, N2508);
xor XOR2 (N3484, N3483, N2181);
nor NOR3 (N3485, N3481, N3349, N2460);
nand NAND2 (N3486, N3484, N1570);
xor XOR2 (N3487, N3457, N1993);
and AND3 (N3488, N3477, N255, N2839);
xor XOR2 (N3489, N3487, N2348);
nor NOR3 (N3490, N3478, N2700, N533);
nor NOR3 (N3491, N3490, N3093, N1473);
or OR4 (N3492, N3486, N902, N2667, N573);
or OR4 (N3493, N3485, N231, N1997, N3320);
not NOT1 (N3494, N3479);
buf BUF1 (N3495, N3492);
nand NAND3 (N3496, N3494, N135, N835);
buf BUF1 (N3497, N3488);
buf BUF1 (N3498, N3493);
xor XOR2 (N3499, N3462, N649);
and AND2 (N3500, N3482, N2121);
or OR3 (N3501, N3500, N204, N929);
nor NOR2 (N3502, N3489, N1303);
and AND4 (N3503, N3495, N434, N3414, N263);
and AND3 (N3504, N3491, N577, N609);
buf BUF1 (N3505, N3480);
not NOT1 (N3506, N3501);
buf BUF1 (N3507, N3503);
xor XOR2 (N3508, N3506, N1987);
and AND4 (N3509, N3504, N2481, N2915, N3377);
nor NOR4 (N3510, N3473, N885, N1966, N1150);
xor XOR2 (N3511, N3509, N1443);
nand NAND2 (N3512, N3510, N1750);
buf BUF1 (N3513, N3511);
not NOT1 (N3514, N3499);
buf BUF1 (N3515, N3497);
not NOT1 (N3516, N3507);
buf BUF1 (N3517, N3508);
xor XOR2 (N3518, N3502, N2226);
or OR3 (N3519, N3514, N545, N342);
nand NAND2 (N3520, N3505, N2053);
buf BUF1 (N3521, N3516);
or OR4 (N3522, N3498, N1761, N2986, N2881);
nand NAND4 (N3523, N3520, N1483, N3077, N2210);
buf BUF1 (N3524, N3518);
or OR2 (N3525, N3513, N945);
nand NAND2 (N3526, N3522, N93);
nand NAND4 (N3527, N3526, N687, N340, N3176);
or OR2 (N3528, N3519, N98);
xor XOR2 (N3529, N3517, N3235);
xor XOR2 (N3530, N3512, N778);
xor XOR2 (N3531, N3527, N524);
and AND2 (N3532, N3525, N2958);
xor XOR2 (N3533, N3524, N1687);
buf BUF1 (N3534, N3496);
xor XOR2 (N3535, N3515, N3169);
xor XOR2 (N3536, N3533, N3193);
not NOT1 (N3537, N3528);
or OR4 (N3538, N3537, N198, N470, N2798);
and AND4 (N3539, N3529, N3505, N3033, N2412);
xor XOR2 (N3540, N3523, N925);
nor NOR4 (N3541, N3532, N2950, N2660, N2821);
not NOT1 (N3542, N3538);
buf BUF1 (N3543, N3542);
nand NAND2 (N3544, N3540, N1097);
not NOT1 (N3545, N3535);
xor XOR2 (N3546, N3531, N1019);
not NOT1 (N3547, N3530);
buf BUF1 (N3548, N3539);
not NOT1 (N3549, N3545);
nor NOR3 (N3550, N3543, N812, N1888);
and AND3 (N3551, N3546, N1529, N2977);
buf BUF1 (N3552, N3551);
nor NOR2 (N3553, N3550, N2020);
nand NAND3 (N3554, N3544, N1823, N3305);
nand NAND4 (N3555, N3553, N1011, N1294, N272);
nand NAND2 (N3556, N3521, N1328);
and AND3 (N3557, N3547, N299, N1437);
buf BUF1 (N3558, N3552);
nor NOR3 (N3559, N3556, N392, N1584);
nor NOR2 (N3560, N3554, N2415);
or OR2 (N3561, N3555, N96);
nand NAND3 (N3562, N3541, N1685, N631);
not NOT1 (N3563, N3549);
or OR4 (N3564, N3559, N448, N2028, N2921);
or OR2 (N3565, N3548, N1351);
nand NAND2 (N3566, N3562, N3105);
nor NOR3 (N3567, N3560, N264, N621);
nor NOR2 (N3568, N3564, N1723);
and AND3 (N3569, N3565, N1727, N2773);
buf BUF1 (N3570, N3563);
nor NOR4 (N3571, N3558, N479, N3332, N3535);
nand NAND3 (N3572, N3567, N1051, N572);
nand NAND2 (N3573, N3566, N323);
nor NOR4 (N3574, N3572, N3372, N3288, N329);
or OR2 (N3575, N3574, N1964);
nand NAND2 (N3576, N3573, N1859);
not NOT1 (N3577, N3536);
not NOT1 (N3578, N3561);
nor NOR3 (N3579, N3570, N48, N2380);
nor NOR4 (N3580, N3568, N3306, N3067, N305);
nand NAND4 (N3581, N3580, N3331, N3267, N1633);
nor NOR3 (N3582, N3569, N3390, N87);
xor XOR2 (N3583, N3579, N1646);
and AND4 (N3584, N3581, N1671, N1710, N308);
not NOT1 (N3585, N3575);
xor XOR2 (N3586, N3584, N2570);
buf BUF1 (N3587, N3571);
nand NAND3 (N3588, N3576, N3322, N2432);
and AND2 (N3589, N3583, N1713);
or OR4 (N3590, N3588, N1275, N1573, N831);
or OR3 (N3591, N3587, N3558, N1403);
and AND2 (N3592, N3589, N1308);
not NOT1 (N3593, N3577);
not NOT1 (N3594, N3534);
nand NAND3 (N3595, N3578, N3370, N227);
and AND4 (N3596, N3592, N645, N110, N3044);
xor XOR2 (N3597, N3593, N470);
buf BUF1 (N3598, N3595);
or OR2 (N3599, N3582, N1619);
or OR2 (N3600, N3557, N2159);
or OR3 (N3601, N3586, N130, N1680);
nor NOR2 (N3602, N3591, N1411);
nand NAND2 (N3603, N3585, N1319);
xor XOR2 (N3604, N3601, N584);
not NOT1 (N3605, N3597);
xor XOR2 (N3606, N3599, N841);
nor NOR4 (N3607, N3600, N1239, N398, N515);
or OR2 (N3608, N3602, N1946);
nor NOR2 (N3609, N3608, N977);
nor NOR4 (N3610, N3609, N2076, N2548, N317);
nand NAND3 (N3611, N3590, N3285, N1250);
nand NAND2 (N3612, N3605, N1955);
buf BUF1 (N3613, N3603);
not NOT1 (N3614, N3610);
nand NAND3 (N3615, N3612, N693, N3079);
or OR4 (N3616, N3606, N2422, N3586, N1666);
nand NAND4 (N3617, N3594, N1078, N984, N3089);
and AND2 (N3618, N3598, N362);
and AND4 (N3619, N3611, N814, N719, N2046);
nor NOR3 (N3620, N3616, N2040, N727);
and AND2 (N3621, N3614, N1689);
nand NAND3 (N3622, N3607, N21, N3518);
and AND2 (N3623, N3619, N2257);
xor XOR2 (N3624, N3613, N3506);
buf BUF1 (N3625, N3624);
nor NOR3 (N3626, N3617, N3271, N3598);
nor NOR4 (N3627, N3622, N1732, N1403, N1519);
or OR2 (N3628, N3621, N1861);
not NOT1 (N3629, N3615);
buf BUF1 (N3630, N3620);
and AND3 (N3631, N3630, N1845, N3587);
xor XOR2 (N3632, N3627, N2382);
not NOT1 (N3633, N3604);
and AND4 (N3634, N3596, N2199, N2160, N3158);
and AND2 (N3635, N3631, N2894);
buf BUF1 (N3636, N3635);
or OR2 (N3637, N3618, N46);
nand NAND3 (N3638, N3628, N535, N2830);
xor XOR2 (N3639, N3625, N2205);
nor NOR2 (N3640, N3634, N2457);
xor XOR2 (N3641, N3633, N1176);
nand NAND3 (N3642, N3626, N252, N2561);
and AND2 (N3643, N3640, N410);
not NOT1 (N3644, N3642);
or OR4 (N3645, N3623, N1091, N1623, N3394);
or OR2 (N3646, N3637, N2359);
and AND2 (N3647, N3636, N2302);
buf BUF1 (N3648, N3647);
nand NAND4 (N3649, N3643, N646, N2986, N1214);
or OR4 (N3650, N3648, N2175, N3638, N533);
and AND2 (N3651, N460, N2257);
and AND4 (N3652, N3649, N2676, N1521, N2116);
or OR3 (N3653, N3641, N592, N1139);
or OR3 (N3654, N3632, N3545, N1588);
nand NAND4 (N3655, N3650, N31, N3237, N2319);
buf BUF1 (N3656, N3639);
xor XOR2 (N3657, N3652, N2192);
buf BUF1 (N3658, N3654);
and AND4 (N3659, N3651, N1999, N1697, N1448);
nand NAND4 (N3660, N3655, N2508, N2287, N1828);
and AND2 (N3661, N3659, N3042);
and AND4 (N3662, N3656, N3131, N3532, N3600);
nor NOR2 (N3663, N3661, N1500);
nand NAND3 (N3664, N3646, N1875, N223);
nand NAND2 (N3665, N3657, N2602);
not NOT1 (N3666, N3629);
buf BUF1 (N3667, N3653);
xor XOR2 (N3668, N3662, N2182);
xor XOR2 (N3669, N3644, N2335);
nor NOR4 (N3670, N3664, N2530, N970, N2172);
xor XOR2 (N3671, N3663, N3214);
nor NOR4 (N3672, N3670, N3022, N1292, N3398);
nand NAND2 (N3673, N3667, N243);
nor NOR2 (N3674, N3668, N1097);
or OR2 (N3675, N3660, N1842);
buf BUF1 (N3676, N3673);
buf BUF1 (N3677, N3674);
xor XOR2 (N3678, N3677, N3503);
and AND2 (N3679, N3669, N426);
nor NOR4 (N3680, N3645, N2417, N3073, N2064);
nor NOR2 (N3681, N3666, N2456);
nor NOR4 (N3682, N3681, N3005, N3264, N272);
not NOT1 (N3683, N3672);
nand NAND3 (N3684, N3671, N1152, N2771);
buf BUF1 (N3685, N3683);
not NOT1 (N3686, N3685);
not NOT1 (N3687, N3679);
buf BUF1 (N3688, N3665);
xor XOR2 (N3689, N3687, N345);
nand NAND2 (N3690, N3689, N1069);
and AND2 (N3691, N3690, N2929);
buf BUF1 (N3692, N3688);
xor XOR2 (N3693, N3686, N930);
nand NAND2 (N3694, N3691, N2216);
nand NAND4 (N3695, N3658, N352, N3019, N1223);
nor NOR4 (N3696, N3695, N1651, N2066, N2985);
nand NAND4 (N3697, N3696, N58, N1151, N1891);
and AND2 (N3698, N3697, N2107);
or OR3 (N3699, N3692, N674, N1976);
nor NOR2 (N3700, N3699, N803);
xor XOR2 (N3701, N3682, N615);
nor NOR4 (N3702, N3680, N444, N2881, N309);
not NOT1 (N3703, N3700);
and AND4 (N3704, N3678, N183, N3006, N432);
nand NAND3 (N3705, N3693, N1805, N3666);
nor NOR4 (N3706, N3694, N1678, N3031, N2675);
buf BUF1 (N3707, N3684);
and AND2 (N3708, N3705, N1336);
or OR4 (N3709, N3707, N956, N524, N140);
xor XOR2 (N3710, N3675, N2035);
nor NOR4 (N3711, N3702, N1270, N1147, N870);
and AND4 (N3712, N3706, N2706, N1757, N915);
not NOT1 (N3713, N3676);
nor NOR2 (N3714, N3710, N3110);
nand NAND3 (N3715, N3714, N3181, N3303);
nor NOR3 (N3716, N3715, N3428, N760);
and AND2 (N3717, N3712, N1110);
nand NAND2 (N3718, N3711, N3019);
nor NOR3 (N3719, N3716, N462, N1209);
not NOT1 (N3720, N3701);
xor XOR2 (N3721, N3709, N3120);
xor XOR2 (N3722, N3704, N667);
or OR2 (N3723, N3717, N2074);
not NOT1 (N3724, N3713);
xor XOR2 (N3725, N3720, N3019);
xor XOR2 (N3726, N3722, N401);
and AND2 (N3727, N3721, N3385);
not NOT1 (N3728, N3718);
nand NAND4 (N3729, N3719, N1072, N1889, N2548);
nand NAND2 (N3730, N3726, N2301);
or OR3 (N3731, N3728, N2097, N668);
or OR2 (N3732, N3708, N283);
buf BUF1 (N3733, N3724);
xor XOR2 (N3734, N3723, N2298);
nor NOR3 (N3735, N3727, N1018, N3624);
nor NOR3 (N3736, N3734, N537, N2833);
buf BUF1 (N3737, N3735);
nor NOR3 (N3738, N3736, N2418, N3652);
buf BUF1 (N3739, N3703);
and AND4 (N3740, N3725, N66, N2541, N132);
xor XOR2 (N3741, N3739, N827);
not NOT1 (N3742, N3731);
or OR4 (N3743, N3730, N379, N3019, N2724);
nand NAND2 (N3744, N3741, N190);
nor NOR2 (N3745, N3742, N3542);
or OR4 (N3746, N3732, N2808, N3745, N1812);
buf BUF1 (N3747, N944);
not NOT1 (N3748, N3737);
not NOT1 (N3749, N3738);
nand NAND3 (N3750, N3743, N1050, N3128);
buf BUF1 (N3751, N3746);
or OR3 (N3752, N3748, N1770, N1942);
nor NOR2 (N3753, N3752, N627);
or OR3 (N3754, N3751, N1432, N1866);
nor NOR2 (N3755, N3744, N3355);
nor NOR3 (N3756, N3733, N2575, N2808);
nor NOR4 (N3757, N3755, N1558, N1970, N1374);
and AND2 (N3758, N3698, N3357);
nor NOR3 (N3759, N3754, N2161, N2730);
nand NAND2 (N3760, N3749, N1309);
or OR3 (N3761, N3758, N2968, N1801);
buf BUF1 (N3762, N3757);
or OR2 (N3763, N3753, N1183);
buf BUF1 (N3764, N3740);
not NOT1 (N3765, N3763);
xor XOR2 (N3766, N3759, N3458);
nand NAND4 (N3767, N3766, N1376, N18, N2667);
buf BUF1 (N3768, N3764);
and AND2 (N3769, N3761, N2503);
buf BUF1 (N3770, N3729);
or OR3 (N3771, N3747, N1868, N1505);
or OR4 (N3772, N3769, N1474, N48, N2520);
and AND3 (N3773, N3772, N3446, N581);
not NOT1 (N3774, N3768);
nand NAND4 (N3775, N3760, N1106, N3084, N3195);
buf BUF1 (N3776, N3756);
xor XOR2 (N3777, N3767, N1411);
xor XOR2 (N3778, N3774, N581);
nand NAND4 (N3779, N3762, N729, N3460, N3368);
or OR2 (N3780, N3750, N287);
xor XOR2 (N3781, N3771, N2006);
xor XOR2 (N3782, N3765, N2598);
nand NAND2 (N3783, N3777, N263);
or OR2 (N3784, N3773, N1995);
not NOT1 (N3785, N3775);
not NOT1 (N3786, N3785);
nand NAND3 (N3787, N3783, N2182, N2798);
and AND4 (N3788, N3784, N1055, N2625, N49);
and AND4 (N3789, N3786, N267, N3701, N1400);
xor XOR2 (N3790, N3779, N561);
nor NOR2 (N3791, N3781, N640);
or OR3 (N3792, N3791, N910, N3038);
nand NAND2 (N3793, N3778, N1232);
or OR3 (N3794, N3770, N2252, N1051);
xor XOR2 (N3795, N3782, N726);
not NOT1 (N3796, N3794);
nor NOR4 (N3797, N3789, N2907, N1751, N1457);
nand NAND3 (N3798, N3787, N2479, N67);
nand NAND4 (N3799, N3793, N3096, N3403, N1772);
not NOT1 (N3800, N3776);
buf BUF1 (N3801, N3799);
nand NAND4 (N3802, N3795, N1783, N1617, N1520);
or OR2 (N3803, N3790, N1596);
or OR2 (N3804, N3798, N1661);
buf BUF1 (N3805, N3788);
xor XOR2 (N3806, N3805, N3520);
nor NOR4 (N3807, N3802, N296, N3197, N2402);
nand NAND2 (N3808, N3804, N1021);
or OR3 (N3809, N3806, N2617, N15);
nor NOR3 (N3810, N3807, N1926, N1267);
nor NOR3 (N3811, N3780, N1922, N1645);
nor NOR3 (N3812, N3800, N602, N3102);
nand NAND2 (N3813, N3796, N942);
buf BUF1 (N3814, N3811);
nand NAND3 (N3815, N3808, N2726, N3160);
and AND4 (N3816, N3797, N2903, N3761, N2744);
xor XOR2 (N3817, N3801, N1117);
and AND2 (N3818, N3813, N2763);
buf BUF1 (N3819, N3815);
buf BUF1 (N3820, N3817);
not NOT1 (N3821, N3809);
buf BUF1 (N3822, N3816);
nor NOR2 (N3823, N3819, N466);
or OR2 (N3824, N3803, N2269);
and AND4 (N3825, N3812, N1449, N3352, N3585);
xor XOR2 (N3826, N3810, N1733);
nand NAND3 (N3827, N3823, N1252, N265);
or OR4 (N3828, N3822, N2936, N1951, N122);
not NOT1 (N3829, N3792);
xor XOR2 (N3830, N3814, N2189);
or OR4 (N3831, N3828, N1084, N3052, N2041);
or OR3 (N3832, N3820, N1459, N2387);
nor NOR2 (N3833, N3831, N3669);
not NOT1 (N3834, N3826);
xor XOR2 (N3835, N3833, N3043);
buf BUF1 (N3836, N3832);
nor NOR3 (N3837, N3835, N2764, N3607);
nor NOR2 (N3838, N3827, N2341);
and AND3 (N3839, N3824, N1448, N3211);
xor XOR2 (N3840, N3836, N1446);
nor NOR3 (N3841, N3840, N846, N762);
xor XOR2 (N3842, N3841, N3129);
nor NOR4 (N3843, N3839, N529, N1574, N2890);
nor NOR2 (N3844, N3838, N3566);
buf BUF1 (N3845, N3842);
nor NOR3 (N3846, N3834, N598, N3117);
not NOT1 (N3847, N3837);
not NOT1 (N3848, N3845);
or OR3 (N3849, N3830, N2028, N1217);
or OR4 (N3850, N3848, N2331, N3684, N964);
or OR2 (N3851, N3821, N1855);
nand NAND4 (N3852, N3847, N653, N2563, N1689);
nand NAND4 (N3853, N3852, N76, N1993, N2140);
nor NOR2 (N3854, N3849, N19);
xor XOR2 (N3855, N3853, N3159);
and AND2 (N3856, N3851, N16);
not NOT1 (N3857, N3855);
or OR3 (N3858, N3850, N872, N1630);
buf BUF1 (N3859, N3858);
buf BUF1 (N3860, N3856);
not NOT1 (N3861, N3860);
nand NAND3 (N3862, N3844, N3329, N2739);
or OR4 (N3863, N3862, N973, N552, N2423);
or OR2 (N3864, N3863, N2239);
or OR4 (N3865, N3843, N759, N879, N409);
or OR3 (N3866, N3825, N904, N2004);
nor NOR4 (N3867, N3866, N3387, N112, N279);
not NOT1 (N3868, N3864);
and AND3 (N3869, N3865, N2325, N597);
xor XOR2 (N3870, N3829, N703);
or OR4 (N3871, N3818, N337, N3376, N3556);
not NOT1 (N3872, N3859);
buf BUF1 (N3873, N3868);
and AND3 (N3874, N3869, N1840, N3366);
or OR3 (N3875, N3871, N2202, N3625);
buf BUF1 (N3876, N3872);
buf BUF1 (N3877, N3857);
nor NOR2 (N3878, N3876, N2132);
buf BUF1 (N3879, N3867);
xor XOR2 (N3880, N3878, N1915);
not NOT1 (N3881, N3870);
nand NAND2 (N3882, N3879, N1707);
or OR2 (N3883, N3873, N2645);
buf BUF1 (N3884, N3875);
buf BUF1 (N3885, N3854);
buf BUF1 (N3886, N3846);
nand NAND3 (N3887, N3874, N2810, N1987);
not NOT1 (N3888, N3885);
not NOT1 (N3889, N3886);
not NOT1 (N3890, N3881);
xor XOR2 (N3891, N3882, N1051);
and AND3 (N3892, N3861, N703, N2841);
or OR4 (N3893, N3889, N3855, N3877, N2897);
or OR2 (N3894, N2106, N980);
and AND2 (N3895, N3893, N2695);
buf BUF1 (N3896, N3888);
nand NAND3 (N3897, N3891, N3451, N2299);
nor NOR2 (N3898, N3897, N2790);
and AND3 (N3899, N3896, N2694, N1630);
xor XOR2 (N3900, N3890, N1396);
nand NAND2 (N3901, N3899, N393);
or OR4 (N3902, N3880, N2080, N1940, N1920);
nand NAND3 (N3903, N3887, N3051, N2520);
nand NAND2 (N3904, N3883, N3515);
buf BUF1 (N3905, N3898);
nand NAND4 (N3906, N3900, N2897, N465, N1684);
xor XOR2 (N3907, N3906, N3149);
not NOT1 (N3908, N3892);
or OR2 (N3909, N3904, N1065);
and AND2 (N3910, N3895, N3609);
xor XOR2 (N3911, N3894, N2732);
not NOT1 (N3912, N3905);
and AND2 (N3913, N3908, N1120);
nor NOR2 (N3914, N3907, N748);
xor XOR2 (N3915, N3902, N432);
buf BUF1 (N3916, N3909);
or OR4 (N3917, N3915, N3527, N2717, N438);
buf BUF1 (N3918, N3912);
or OR3 (N3919, N3901, N2262, N1987);
buf BUF1 (N3920, N3917);
nor NOR2 (N3921, N3916, N1431);
nand NAND2 (N3922, N3919, N2951);
buf BUF1 (N3923, N3914);
nor NOR2 (N3924, N3884, N3901);
or OR2 (N3925, N3921, N3209);
not NOT1 (N3926, N3911);
nand NAND4 (N3927, N3922, N2663, N671, N1569);
buf BUF1 (N3928, N3910);
or OR2 (N3929, N3918, N215);
nand NAND4 (N3930, N3913, N3316, N426, N1297);
or OR3 (N3931, N3924, N3292, N1080);
buf BUF1 (N3932, N3925);
not NOT1 (N3933, N3929);
nand NAND2 (N3934, N3931, N1309);
or OR4 (N3935, N3926, N168, N391, N1932);
nand NAND2 (N3936, N3930, N1308);
xor XOR2 (N3937, N3928, N253);
and AND4 (N3938, N3932, N2709, N2361, N1667);
nor NOR2 (N3939, N3903, N397);
xor XOR2 (N3940, N3939, N3633);
and AND4 (N3941, N3938, N218, N1902, N2702);
and AND4 (N3942, N3937, N3350, N1366, N511);
not NOT1 (N3943, N3934);
buf BUF1 (N3944, N3923);
buf BUF1 (N3945, N3941);
or OR4 (N3946, N3933, N2024, N1364, N2124);
nand NAND4 (N3947, N3946, N1829, N1721, N1172);
xor XOR2 (N3948, N3945, N2837);
buf BUF1 (N3949, N3943);
nand NAND3 (N3950, N3920, N1547, N3713);
nor NOR3 (N3951, N3927, N878, N1828);
nor NOR3 (N3952, N3950, N1165, N721);
xor XOR2 (N3953, N3947, N2253);
nand NAND4 (N3954, N3944, N2254, N3118, N2440);
buf BUF1 (N3955, N3954);
xor XOR2 (N3956, N3935, N3127);
nor NOR2 (N3957, N3955, N3490);
buf BUF1 (N3958, N3952);
not NOT1 (N3959, N3949);
nand NAND4 (N3960, N3953, N1999, N1293, N3709);
nand NAND3 (N3961, N3960, N3326, N610);
buf BUF1 (N3962, N3961);
xor XOR2 (N3963, N3948, N1005);
or OR2 (N3964, N3956, N95);
not NOT1 (N3965, N3936);
nor NOR3 (N3966, N3942, N1527, N1572);
and AND3 (N3967, N3958, N1292, N514);
xor XOR2 (N3968, N3957, N300);
nor NOR3 (N3969, N3968, N1718, N904);
or OR3 (N3970, N3964, N3305, N558);
and AND3 (N3971, N3963, N2348, N2117);
or OR3 (N3972, N3965, N2520, N2657);
nand NAND3 (N3973, N3951, N2393, N3965);
not NOT1 (N3974, N3970);
nand NAND3 (N3975, N3971, N534, N408);
buf BUF1 (N3976, N3973);
nor NOR4 (N3977, N3975, N3915, N3550, N2211);
not NOT1 (N3978, N3966);
nor NOR4 (N3979, N3969, N2160, N2135, N1022);
buf BUF1 (N3980, N3978);
buf BUF1 (N3981, N3976);
or OR4 (N3982, N3981, N3527, N297, N1532);
nand NAND2 (N3983, N3940, N1527);
and AND2 (N3984, N3962, N1807);
nor NOR2 (N3985, N3959, N1431);
not NOT1 (N3986, N3983);
or OR2 (N3987, N3982, N1975);
nand NAND3 (N3988, N3986, N3048, N3020);
not NOT1 (N3989, N3977);
not NOT1 (N3990, N3972);
nand NAND4 (N3991, N3984, N1136, N15, N1209);
buf BUF1 (N3992, N3990);
xor XOR2 (N3993, N3992, N122);
buf BUF1 (N3994, N3987);
nand NAND4 (N3995, N3974, N3714, N3825, N1582);
nand NAND4 (N3996, N3985, N1620, N132, N3243);
nand NAND4 (N3997, N3979, N2106, N68, N1846);
nand NAND2 (N3998, N3991, N2332);
or OR4 (N3999, N3989, N2602, N714, N519);
nor NOR3 (N4000, N3999, N2944, N1309);
and AND2 (N4001, N3993, N3866);
or OR4 (N4002, N4001, N2439, N3689, N1);
and AND2 (N4003, N3980, N606);
nor NOR2 (N4004, N3988, N2344);
nand NAND4 (N4005, N3998, N779, N2607, N2030);
nand NAND2 (N4006, N4003, N3272);
not NOT1 (N4007, N3967);
not NOT1 (N4008, N4002);
xor XOR2 (N4009, N4006, N3192);
or OR4 (N4010, N3994, N1827, N3681, N3754);
buf BUF1 (N4011, N4004);
not NOT1 (N4012, N4008);
not NOT1 (N4013, N3996);
or OR2 (N4014, N3995, N3664);
buf BUF1 (N4015, N4009);
nand NAND4 (N4016, N4011, N3292, N766, N2229);
nor NOR2 (N4017, N4007, N3068);
or OR3 (N4018, N4013, N605, N2459);
and AND2 (N4019, N4000, N2378);
and AND2 (N4020, N4015, N3212);
xor XOR2 (N4021, N4012, N2371);
buf BUF1 (N4022, N4016);
xor XOR2 (N4023, N3997, N1399);
nor NOR2 (N4024, N4014, N2943);
xor XOR2 (N4025, N4010, N1155);
nor NOR3 (N4026, N4021, N2675, N704);
not NOT1 (N4027, N4023);
nand NAND3 (N4028, N4024, N3677, N1428);
or OR4 (N4029, N4028, N3221, N437, N65);
buf BUF1 (N4030, N4019);
or OR4 (N4031, N4017, N1058, N1952, N2108);
nand NAND2 (N4032, N4029, N3542);
xor XOR2 (N4033, N4005, N3056);
nor NOR3 (N4034, N4018, N482, N1051);
and AND2 (N4035, N4031, N325);
not NOT1 (N4036, N4032);
not NOT1 (N4037, N4030);
and AND2 (N4038, N4020, N1650);
and AND3 (N4039, N4033, N3771, N639);
nand NAND3 (N4040, N4036, N3544, N2395);
not NOT1 (N4041, N4039);
and AND4 (N4042, N4025, N3218, N150, N2783);
buf BUF1 (N4043, N4035);
nand NAND2 (N4044, N4034, N1867);
nor NOR4 (N4045, N4038, N1097, N642, N2339);
buf BUF1 (N4046, N4041);
buf BUF1 (N4047, N4043);
nand NAND3 (N4048, N4026, N2684, N3827);
nor NOR2 (N4049, N4048, N3435);
and AND3 (N4050, N4045, N2883, N1780);
or OR4 (N4051, N4037, N1810, N1781, N953);
xor XOR2 (N4052, N4047, N2554);
buf BUF1 (N4053, N4049);
nor NOR3 (N4054, N4044, N2672, N1648);
and AND4 (N4055, N4040, N654, N982, N2617);
nor NOR4 (N4056, N4022, N687, N13, N308);
and AND3 (N4057, N4050, N1172, N2062);
nor NOR3 (N4058, N4051, N802, N1803);
nand NAND3 (N4059, N4027, N1310, N3235);
buf BUF1 (N4060, N4057);
not NOT1 (N4061, N4052);
xor XOR2 (N4062, N4053, N1553);
and AND4 (N4063, N4056, N104, N2566, N767);
buf BUF1 (N4064, N4061);
nand NAND2 (N4065, N4042, N3261);
nand NAND4 (N4066, N4064, N900, N1382, N1568);
xor XOR2 (N4067, N4066, N2738);
buf BUF1 (N4068, N4046);
nor NOR2 (N4069, N4062, N655);
and AND3 (N4070, N4054, N330, N392);
and AND2 (N4071, N4058, N2488);
nor NOR3 (N4072, N4067, N627, N998);
not NOT1 (N4073, N4069);
nand NAND4 (N4074, N4071, N1441, N2597, N4046);
nand NAND4 (N4075, N4059, N3809, N3288, N3459);
or OR3 (N4076, N4073, N2537, N2750);
buf BUF1 (N4077, N4076);
xor XOR2 (N4078, N4055, N2347);
xor XOR2 (N4079, N4070, N2091);
buf BUF1 (N4080, N4065);
not NOT1 (N4081, N4077);
not NOT1 (N4082, N4072);
nor NOR3 (N4083, N4068, N675, N1814);
and AND3 (N4084, N4060, N673, N1073);
xor XOR2 (N4085, N4079, N2816);
and AND3 (N4086, N4085, N1666, N1662);
or OR2 (N4087, N4078, N1668);
not NOT1 (N4088, N4081);
or OR3 (N4089, N4083, N1087, N2523);
xor XOR2 (N4090, N4075, N3618);
buf BUF1 (N4091, N4090);
not NOT1 (N4092, N4082);
or OR2 (N4093, N4088, N3772);
buf BUF1 (N4094, N4092);
nor NOR2 (N4095, N4063, N3889);
buf BUF1 (N4096, N4087);
nand NAND4 (N4097, N4086, N680, N895, N332);
buf BUF1 (N4098, N4091);
nand NAND3 (N4099, N4096, N66, N3543);
nor NOR2 (N4100, N4074, N1341);
xor XOR2 (N4101, N4095, N1390);
and AND3 (N4102, N4097, N1832, N829);
or OR3 (N4103, N4102, N2735, N1835);
nor NOR2 (N4104, N4100, N3448);
buf BUF1 (N4105, N4093);
and AND3 (N4106, N4105, N18, N3122);
buf BUF1 (N4107, N4104);
buf BUF1 (N4108, N4099);
and AND2 (N4109, N4094, N4015);
not NOT1 (N4110, N4103);
xor XOR2 (N4111, N4106, N4059);
or OR3 (N4112, N4108, N3052, N2968);
xor XOR2 (N4113, N4110, N1231);
nor NOR3 (N4114, N4080, N891, N2592);
nand NAND3 (N4115, N4109, N1033, N3990);
and AND2 (N4116, N4111, N2986);
and AND2 (N4117, N4114, N3378);
buf BUF1 (N4118, N4107);
xor XOR2 (N4119, N4115, N682);
and AND4 (N4120, N4084, N1984, N562, N2235);
xor XOR2 (N4121, N4119, N165);
nand NAND4 (N4122, N4113, N3638, N92, N1064);
not NOT1 (N4123, N4116);
buf BUF1 (N4124, N4112);
not NOT1 (N4125, N4117);
not NOT1 (N4126, N4121);
not NOT1 (N4127, N4118);
nor NOR4 (N4128, N4126, N1599, N1586, N303);
nor NOR3 (N4129, N4125, N2786, N2653);
not NOT1 (N4130, N4127);
not NOT1 (N4131, N4129);
or OR3 (N4132, N4124, N2444, N115);
xor XOR2 (N4133, N4101, N944);
nand NAND4 (N4134, N4128, N357, N3163, N3112);
and AND4 (N4135, N4123, N3471, N557, N400);
or OR2 (N4136, N4089, N3254);
or OR2 (N4137, N4120, N1435);
xor XOR2 (N4138, N4130, N3175);
xor XOR2 (N4139, N4135, N2656);
nor NOR2 (N4140, N4131, N2216);
and AND4 (N4141, N4133, N1971, N3086, N3359);
xor XOR2 (N4142, N4140, N1255);
nand NAND3 (N4143, N4122, N3849, N3958);
or OR2 (N4144, N4142, N409);
and AND2 (N4145, N4136, N2123);
xor XOR2 (N4146, N4132, N4010);
or OR3 (N4147, N4143, N175, N2614);
not NOT1 (N4148, N4145);
or OR2 (N4149, N4148, N1342);
nand NAND4 (N4150, N4138, N2971, N4099, N610);
and AND4 (N4151, N4139, N3674, N3125, N804);
and AND2 (N4152, N4134, N3581);
and AND3 (N4153, N4151, N2575, N590);
and AND2 (N4154, N4141, N2751);
or OR2 (N4155, N4098, N2441);
not NOT1 (N4156, N4150);
nor NOR3 (N4157, N4153, N2633, N3183);
buf BUF1 (N4158, N4152);
buf BUF1 (N4159, N4155);
or OR4 (N4160, N4154, N3811, N3323, N1492);
buf BUF1 (N4161, N4144);
nor NOR4 (N4162, N4146, N4128, N1231, N326);
and AND4 (N4163, N4159, N3011, N1172, N3370);
not NOT1 (N4164, N4160);
xor XOR2 (N4165, N4164, N3121);
xor XOR2 (N4166, N4161, N2144);
or OR2 (N4167, N4147, N2139);
or OR2 (N4168, N4167, N2341);
or OR3 (N4169, N4137, N1235, N515);
or OR3 (N4170, N4165, N2568, N794);
xor XOR2 (N4171, N4169, N2663);
xor XOR2 (N4172, N4149, N514);
and AND3 (N4173, N4171, N3053, N1774);
nor NOR3 (N4174, N4168, N611, N2379);
xor XOR2 (N4175, N4170, N635);
xor XOR2 (N4176, N4173, N2779);
nand NAND2 (N4177, N4172, N3331);
buf BUF1 (N4178, N4174);
buf BUF1 (N4179, N4163);
or OR2 (N4180, N4179, N3199);
not NOT1 (N4181, N4162);
xor XOR2 (N4182, N4157, N1411);
buf BUF1 (N4183, N4176);
or OR3 (N4184, N4180, N3386, N184);
buf BUF1 (N4185, N4181);
not NOT1 (N4186, N4166);
nand NAND2 (N4187, N4177, N1777);
xor XOR2 (N4188, N4158, N135);
xor XOR2 (N4189, N4156, N1221);
not NOT1 (N4190, N4178);
xor XOR2 (N4191, N4189, N2710);
or OR3 (N4192, N4184, N2723, N3507);
nand NAND2 (N4193, N4183, N1445);
nand NAND3 (N4194, N4191, N3098, N1042);
not NOT1 (N4195, N4175);
nand NAND4 (N4196, N4195, N3928, N448, N4174);
buf BUF1 (N4197, N4190);
nand NAND3 (N4198, N4187, N4189, N3409);
or OR3 (N4199, N4193, N1401, N2256);
xor XOR2 (N4200, N4186, N88);
not NOT1 (N4201, N4194);
not NOT1 (N4202, N4200);
nor NOR3 (N4203, N4202, N3165, N3540);
nand NAND2 (N4204, N4192, N3626);
not NOT1 (N4205, N4204);
buf BUF1 (N4206, N4198);
nor NOR4 (N4207, N4182, N874, N3523, N3661);
nor NOR3 (N4208, N4197, N2156, N260);
buf BUF1 (N4209, N4203);
not NOT1 (N4210, N4185);
not NOT1 (N4211, N4209);
buf BUF1 (N4212, N4205);
nand NAND3 (N4213, N4210, N3636, N652);
not NOT1 (N4214, N4188);
xor XOR2 (N4215, N4214, N604);
and AND3 (N4216, N4208, N1756, N1778);
nor NOR2 (N4217, N4199, N989);
and AND2 (N4218, N4212, N2612);
not NOT1 (N4219, N4218);
or OR4 (N4220, N4219, N2421, N3895, N2149);
not NOT1 (N4221, N4217);
nand NAND4 (N4222, N4196, N3682, N3151, N1804);
and AND3 (N4223, N4221, N3983, N877);
buf BUF1 (N4224, N4220);
not NOT1 (N4225, N4207);
nor NOR3 (N4226, N4222, N2272, N2454);
and AND2 (N4227, N4216, N557);
and AND4 (N4228, N4206, N160, N274, N3535);
xor XOR2 (N4229, N4201, N825);
and AND2 (N4230, N4213, N2761);
nand NAND3 (N4231, N4230, N875, N2827);
or OR3 (N4232, N4224, N888, N2261);
nor NOR4 (N4233, N4227, N256, N1969, N2050);
or OR4 (N4234, N4215, N3474, N1432, N1063);
not NOT1 (N4235, N4228);
nor NOR2 (N4236, N4226, N1577);
and AND3 (N4237, N4211, N3634, N2731);
and AND4 (N4238, N4235, N1808, N142, N2959);
and AND4 (N4239, N4233, N465, N2069, N2709);
nor NOR2 (N4240, N4239, N1896);
xor XOR2 (N4241, N4223, N2521);
and AND2 (N4242, N4225, N516);
buf BUF1 (N4243, N4236);
and AND4 (N4244, N4240, N2269, N2890, N3169);
buf BUF1 (N4245, N4243);
buf BUF1 (N4246, N4232);
nand NAND2 (N4247, N4231, N2527);
nor NOR4 (N4248, N4244, N1586, N1657, N584);
xor XOR2 (N4249, N4245, N2268);
or OR4 (N4250, N4249, N3230, N3418, N718);
nor NOR3 (N4251, N4238, N310, N1079);
buf BUF1 (N4252, N4247);
buf BUF1 (N4253, N4248);
buf BUF1 (N4254, N4251);
buf BUF1 (N4255, N4253);
nand NAND2 (N4256, N4229, N2865);
nor NOR4 (N4257, N4252, N4234, N3913, N3631);
nor NOR3 (N4258, N2143, N282, N3357);
xor XOR2 (N4259, N4256, N2799);
nand NAND3 (N4260, N4250, N3739, N3149);
nand NAND4 (N4261, N4254, N3013, N2223, N2257);
and AND4 (N4262, N4257, N1080, N1938, N579);
and AND4 (N4263, N4242, N3043, N191, N1442);
nand NAND4 (N4264, N4255, N175, N609, N1357);
buf BUF1 (N4265, N4261);
not NOT1 (N4266, N4258);
xor XOR2 (N4267, N4266, N1132);
nor NOR3 (N4268, N4237, N115, N3700);
not NOT1 (N4269, N4267);
buf BUF1 (N4270, N4241);
not NOT1 (N4271, N4264);
not NOT1 (N4272, N4260);
nand NAND2 (N4273, N4246, N2868);
not NOT1 (N4274, N4265);
not NOT1 (N4275, N4273);
buf BUF1 (N4276, N4271);
nor NOR3 (N4277, N4268, N2407, N3950);
nand NAND3 (N4278, N4263, N1905, N14);
buf BUF1 (N4279, N4270);
buf BUF1 (N4280, N4259);
nor NOR2 (N4281, N4278, N2416);
nor NOR2 (N4282, N4277, N3080);
buf BUF1 (N4283, N4280);
xor XOR2 (N4284, N4276, N682);
xor XOR2 (N4285, N4279, N4275);
or OR2 (N4286, N2375, N1012);
xor XOR2 (N4287, N4269, N2967);
nand NAND3 (N4288, N4287, N799, N4133);
buf BUF1 (N4289, N4288);
buf BUF1 (N4290, N4282);
xor XOR2 (N4291, N4283, N1022);
nor NOR4 (N4292, N4284, N2940, N1428, N4229);
nor NOR4 (N4293, N4286, N298, N2051, N2545);
nand NAND2 (N4294, N4262, N2283);
xor XOR2 (N4295, N4293, N91);
nand NAND4 (N4296, N4274, N3187, N4222, N164);
or OR2 (N4297, N4295, N2685);
xor XOR2 (N4298, N4281, N2718);
xor XOR2 (N4299, N4290, N1077);
and AND3 (N4300, N4299, N32, N2539);
xor XOR2 (N4301, N4298, N2335);
buf BUF1 (N4302, N4294);
not NOT1 (N4303, N4296);
and AND2 (N4304, N4291, N2200);
not NOT1 (N4305, N4303);
nand NAND4 (N4306, N4304, N2237, N917, N2944);
nor NOR4 (N4307, N4272, N3376, N1362, N2791);
xor XOR2 (N4308, N4285, N1479);
buf BUF1 (N4309, N4301);
nand NAND2 (N4310, N4300, N2405);
and AND3 (N4311, N4306, N556, N2354);
and AND4 (N4312, N4302, N4193, N1825, N3803);
nor NOR3 (N4313, N4308, N3645, N815);
not NOT1 (N4314, N4311);
and AND2 (N4315, N4297, N3820);
nand NAND3 (N4316, N4310, N2511, N2485);
not NOT1 (N4317, N4289);
nor NOR2 (N4318, N4307, N2354);
nand NAND3 (N4319, N4317, N3360, N1736);
xor XOR2 (N4320, N4316, N1980);
or OR4 (N4321, N4318, N3424, N263, N1411);
nand NAND4 (N4322, N4314, N3003, N3610, N578);
not NOT1 (N4323, N4322);
and AND2 (N4324, N4319, N784);
not NOT1 (N4325, N4315);
nand NAND4 (N4326, N4312, N3395, N2988, N3357);
or OR3 (N4327, N4320, N2741, N1482);
nand NAND2 (N4328, N4326, N1238);
and AND4 (N4329, N4323, N2864, N7, N1960);
nor NOR3 (N4330, N4292, N4059, N3192);
nand NAND2 (N4331, N4305, N2773);
buf BUF1 (N4332, N4328);
or OR2 (N4333, N4331, N1396);
and AND4 (N4334, N4309, N2985, N845, N1752);
and AND2 (N4335, N4327, N2345);
buf BUF1 (N4336, N4329);
nand NAND4 (N4337, N4313, N3821, N106, N3925);
xor XOR2 (N4338, N4334, N1415);
or OR3 (N4339, N4338, N111, N276);
buf BUF1 (N4340, N4335);
or OR4 (N4341, N4321, N2884, N3647, N2330);
not NOT1 (N4342, N4324);
buf BUF1 (N4343, N4339);
or OR4 (N4344, N4336, N1304, N2125, N3615);
and AND4 (N4345, N4344, N3091, N3692, N1131);
not NOT1 (N4346, N4343);
and AND4 (N4347, N4340, N470, N3094, N4268);
xor XOR2 (N4348, N4330, N2779);
not NOT1 (N4349, N4333);
nor NOR2 (N4350, N4337, N4280);
nor NOR2 (N4351, N4348, N938);
xor XOR2 (N4352, N4332, N2668);
buf BUF1 (N4353, N4342);
not NOT1 (N4354, N4346);
xor XOR2 (N4355, N4325, N3579);
nand NAND4 (N4356, N4347, N215, N3845, N261);
and AND3 (N4357, N4353, N1873, N3945);
xor XOR2 (N4358, N4345, N3669);
nand NAND3 (N4359, N4341, N746, N482);
or OR4 (N4360, N4351, N3086, N931, N2104);
not NOT1 (N4361, N4355);
xor XOR2 (N4362, N4358, N1061);
buf BUF1 (N4363, N4361);
nor NOR4 (N4364, N4349, N232, N2613, N3775);
nor NOR4 (N4365, N4363, N750, N3403, N2647);
and AND4 (N4366, N4350, N2951, N801, N3550);
and AND4 (N4367, N4357, N3239, N1670, N400);
not NOT1 (N4368, N4367);
and AND4 (N4369, N4364, N1208, N1302, N2122);
nand NAND4 (N4370, N4352, N3272, N1650, N2618);
nor NOR2 (N4371, N4354, N2624);
nor NOR2 (N4372, N4370, N1124);
nor NOR3 (N4373, N4371, N4266, N3160);
buf BUF1 (N4374, N4356);
not NOT1 (N4375, N4374);
nor NOR4 (N4376, N4366, N3640, N1942, N4135);
xor XOR2 (N4377, N4362, N196);
xor XOR2 (N4378, N4375, N2142);
or OR2 (N4379, N4360, N369);
buf BUF1 (N4380, N4376);
nand NAND4 (N4381, N4380, N3090, N3385, N4353);
nor NOR3 (N4382, N4372, N2350, N838);
not NOT1 (N4383, N4368);
or OR2 (N4384, N4377, N1742);
not NOT1 (N4385, N4382);
and AND2 (N4386, N4373, N3041);
xor XOR2 (N4387, N4383, N90);
or OR2 (N4388, N4365, N4212);
buf BUF1 (N4389, N4386);
xor XOR2 (N4390, N4388, N2575);
and AND3 (N4391, N4387, N2200, N3325);
nand NAND3 (N4392, N4379, N3556, N209);
not NOT1 (N4393, N4378);
or OR4 (N4394, N4369, N3143, N3336, N4138);
not NOT1 (N4395, N4390);
not NOT1 (N4396, N4395);
and AND3 (N4397, N4391, N3844, N1096);
buf BUF1 (N4398, N4393);
or OR3 (N4399, N4385, N2776, N2151);
or OR4 (N4400, N4381, N1588, N4303, N27);
or OR3 (N4401, N4399, N11, N950);
nor NOR4 (N4402, N4392, N3244, N2700, N3759);
nand NAND2 (N4403, N4389, N2246);
or OR4 (N4404, N4359, N2543, N2792, N4381);
buf BUF1 (N4405, N4394);
or OR3 (N4406, N4404, N3690, N3944);
buf BUF1 (N4407, N4405);
nor NOR3 (N4408, N4402, N3768, N3180);
and AND4 (N4409, N4398, N2659, N1303, N1847);
xor XOR2 (N4410, N4396, N3666);
buf BUF1 (N4411, N4407);
not NOT1 (N4412, N4403);
nand NAND2 (N4413, N4409, N1166);
nand NAND4 (N4414, N4401, N3495, N1452, N2205);
xor XOR2 (N4415, N4412, N2070);
buf BUF1 (N4416, N4410);
xor XOR2 (N4417, N4406, N537);
nand NAND4 (N4418, N4408, N2966, N1726, N3819);
and AND4 (N4419, N4400, N818, N1984, N2568);
or OR4 (N4420, N4418, N2487, N1627, N1803);
not NOT1 (N4421, N4415);
not NOT1 (N4422, N4420);
nor NOR4 (N4423, N4416, N2641, N505, N3962);
nor NOR2 (N4424, N4397, N4205);
nor NOR2 (N4425, N4422, N2575);
or OR4 (N4426, N4384, N1042, N1618, N1438);
and AND2 (N4427, N4419, N668);
nand NAND2 (N4428, N4411, N1466);
nor NOR4 (N4429, N4423, N2605, N2881, N997);
nand NAND3 (N4430, N4424, N1765, N3428);
nand NAND4 (N4431, N4425, N4079, N1341, N3173);
nand NAND3 (N4432, N4430, N2144, N2738);
nand NAND3 (N4433, N4417, N2463, N916);
nand NAND3 (N4434, N4432, N3684, N2995);
nor NOR4 (N4435, N4414, N3485, N3546, N2425);
not NOT1 (N4436, N4431);
and AND4 (N4437, N4435, N275, N2817, N4347);
xor XOR2 (N4438, N4429, N1257);
or OR3 (N4439, N4437, N1269, N1354);
buf BUF1 (N4440, N4426);
buf BUF1 (N4441, N4436);
nor NOR3 (N4442, N4439, N1841, N4276);
buf BUF1 (N4443, N4427);
not NOT1 (N4444, N4433);
xor XOR2 (N4445, N4444, N458);
not NOT1 (N4446, N4428);
nor NOR2 (N4447, N4443, N2328);
not NOT1 (N4448, N4434);
xor XOR2 (N4449, N4448, N1077);
nor NOR2 (N4450, N4438, N3420);
nand NAND4 (N4451, N4446, N4030, N5, N1921);
and AND4 (N4452, N4451, N515, N2057, N949);
or OR3 (N4453, N4421, N63, N2266);
nor NOR4 (N4454, N4452, N623, N3908, N838);
buf BUF1 (N4455, N4440);
buf BUF1 (N4456, N4442);
or OR4 (N4457, N4449, N2098, N3641, N2980);
and AND2 (N4458, N4447, N4220);
and AND3 (N4459, N4454, N1708, N2101);
and AND2 (N4460, N4457, N4093);
and AND2 (N4461, N4460, N1621);
not NOT1 (N4462, N4413);
buf BUF1 (N4463, N4450);
nand NAND2 (N4464, N4463, N212);
xor XOR2 (N4465, N4445, N3929);
buf BUF1 (N4466, N4464);
not NOT1 (N4467, N4466);
xor XOR2 (N4468, N4467, N1059);
buf BUF1 (N4469, N4459);
not NOT1 (N4470, N4461);
buf BUF1 (N4471, N4468);
or OR4 (N4472, N4455, N2318, N1034, N1568);
not NOT1 (N4473, N4471);
nand NAND2 (N4474, N4465, N466);
or OR2 (N4475, N4456, N2426);
xor XOR2 (N4476, N4469, N3912);
buf BUF1 (N4477, N4441);
buf BUF1 (N4478, N4458);
nor NOR4 (N4479, N4476, N1107, N2789, N1506);
nor NOR2 (N4480, N4477, N4325);
nand NAND2 (N4481, N4475, N3995);
buf BUF1 (N4482, N4481);
buf BUF1 (N4483, N4479);
not NOT1 (N4484, N4474);
or OR2 (N4485, N4472, N2235);
or OR4 (N4486, N4484, N593, N974, N4081);
or OR2 (N4487, N4485, N949);
not NOT1 (N4488, N4480);
nor NOR4 (N4489, N4482, N1365, N4223, N4307);
not NOT1 (N4490, N4473);
or OR3 (N4491, N4483, N641, N3395);
not NOT1 (N4492, N4487);
and AND3 (N4493, N4478, N3955, N2658);
nor NOR2 (N4494, N4492, N3715);
buf BUF1 (N4495, N4490);
and AND3 (N4496, N4489, N2462, N3421);
and AND3 (N4497, N4495, N4363, N342);
nand NAND2 (N4498, N4486, N193);
xor XOR2 (N4499, N4462, N1314);
not NOT1 (N4500, N4494);
not NOT1 (N4501, N4470);
buf BUF1 (N4502, N4453);
and AND3 (N4503, N4498, N469, N4121);
nand NAND4 (N4504, N4502, N2266, N1757, N4369);
not NOT1 (N4505, N4504);
and AND2 (N4506, N4488, N3260);
buf BUF1 (N4507, N4496);
nor NOR4 (N4508, N4493, N1390, N60, N3703);
and AND2 (N4509, N4505, N393);
or OR2 (N4510, N4497, N194);
and AND4 (N4511, N4503, N4201, N1187, N3784);
xor XOR2 (N4512, N4511, N386);
nor NOR2 (N4513, N4500, N1980);
or OR2 (N4514, N4499, N1126);
and AND4 (N4515, N4491, N2377, N2229, N3311);
buf BUF1 (N4516, N4515);
not NOT1 (N4517, N4501);
or OR2 (N4518, N4512, N4515);
not NOT1 (N4519, N4518);
not NOT1 (N4520, N4507);
not NOT1 (N4521, N4509);
xor XOR2 (N4522, N4519, N2156);
nor NOR2 (N4523, N4521, N3613);
not NOT1 (N4524, N4522);
not NOT1 (N4525, N4510);
buf BUF1 (N4526, N4514);
nand NAND3 (N4527, N4516, N4017, N1060);
not NOT1 (N4528, N4524);
nor NOR2 (N4529, N4517, N2990);
xor XOR2 (N4530, N4508, N4307);
nand NAND2 (N4531, N4526, N2475);
or OR2 (N4532, N4525, N3269);
or OR4 (N4533, N4527, N1011, N1530, N1802);
buf BUF1 (N4534, N4532);
not NOT1 (N4535, N4530);
xor XOR2 (N4536, N4533, N2272);
buf BUF1 (N4537, N4520);
buf BUF1 (N4538, N4528);
not NOT1 (N4539, N4537);
xor XOR2 (N4540, N4513, N1851);
nand NAND3 (N4541, N4531, N2313, N1742);
nor NOR3 (N4542, N4538, N1148, N2891);
and AND3 (N4543, N4529, N2110, N1677);
or OR2 (N4544, N4539, N2064);
and AND2 (N4545, N4541, N3440);
nand NAND4 (N4546, N4544, N1713, N4081, N3662);
nor NOR2 (N4547, N4536, N1575);
buf BUF1 (N4548, N4546);
xor XOR2 (N4549, N4523, N4437);
xor XOR2 (N4550, N4543, N2645);
xor XOR2 (N4551, N4506, N2215);
not NOT1 (N4552, N4545);
buf BUF1 (N4553, N4542);
nor NOR4 (N4554, N4549, N1155, N1854, N683);
and AND2 (N4555, N4552, N1101);
buf BUF1 (N4556, N4553);
xor XOR2 (N4557, N4534, N605);
buf BUF1 (N4558, N4556);
buf BUF1 (N4559, N4555);
nand NAND4 (N4560, N4547, N2316, N652, N4330);
buf BUF1 (N4561, N4554);
buf BUF1 (N4562, N4535);
or OR2 (N4563, N4557, N248);
not NOT1 (N4564, N4563);
buf BUF1 (N4565, N4562);
nor NOR4 (N4566, N4565, N1349, N4163, N2157);
and AND4 (N4567, N4540, N544, N2538, N2434);
or OR3 (N4568, N4559, N1137, N197);
and AND2 (N4569, N4561, N337);
nor NOR4 (N4570, N4550, N2207, N2602, N3228);
and AND3 (N4571, N4558, N4201, N1183);
and AND2 (N4572, N4570, N3555);
buf BUF1 (N4573, N4560);
or OR3 (N4574, N4548, N1154, N359);
nor NOR2 (N4575, N4573, N1674);
and AND3 (N4576, N4564, N2420, N3902);
nor NOR3 (N4577, N4566, N3481, N580);
not NOT1 (N4578, N4576);
and AND3 (N4579, N4577, N3365, N4428);
nand NAND3 (N4580, N4568, N2370, N1425);
and AND3 (N4581, N4578, N2952, N4394);
and AND3 (N4582, N4569, N4325, N492);
and AND4 (N4583, N4575, N1423, N2334, N1407);
or OR2 (N4584, N4572, N837);
not NOT1 (N4585, N4583);
not NOT1 (N4586, N4567);
and AND3 (N4587, N4551, N2206, N1718);
buf BUF1 (N4588, N4586);
not NOT1 (N4589, N4585);
buf BUF1 (N4590, N4584);
not NOT1 (N4591, N4582);
xor XOR2 (N4592, N4587, N3495);
nor NOR2 (N4593, N4592, N1958);
nand NAND3 (N4594, N4574, N2033, N3354);
nor NOR3 (N4595, N4590, N2766, N1003);
or OR2 (N4596, N4580, N3424);
nand NAND2 (N4597, N4581, N2416);
xor XOR2 (N4598, N4597, N4401);
buf BUF1 (N4599, N4594);
nor NOR4 (N4600, N4589, N3814, N3654, N1728);
not NOT1 (N4601, N4598);
not NOT1 (N4602, N4595);
nor NOR3 (N4603, N4601, N1610, N4023);
nor NOR4 (N4604, N4602, N3237, N976, N3102);
not NOT1 (N4605, N4604);
buf BUF1 (N4606, N4603);
or OR3 (N4607, N4600, N608, N3294);
or OR3 (N4608, N4596, N1146, N2209);
and AND2 (N4609, N4599, N96);
xor XOR2 (N4610, N4579, N4345);
not NOT1 (N4611, N4593);
buf BUF1 (N4612, N4588);
buf BUF1 (N4613, N4591);
xor XOR2 (N4614, N4571, N3707);
xor XOR2 (N4615, N4610, N2857);
and AND2 (N4616, N4609, N3686);
xor XOR2 (N4617, N4608, N4186);
or OR2 (N4618, N4615, N4451);
nor NOR4 (N4619, N4606, N3144, N1333, N1321);
or OR2 (N4620, N4619, N160);
and AND4 (N4621, N4613, N3104, N2217, N2047);
buf BUF1 (N4622, N4621);
not NOT1 (N4623, N4612);
nor NOR2 (N4624, N4607, N2991);
or OR3 (N4625, N4616, N4079, N2611);
nor NOR3 (N4626, N4618, N637, N1595);
and AND3 (N4627, N4605, N4392, N581);
buf BUF1 (N4628, N4626);
and AND3 (N4629, N4622, N3112, N215);
or OR2 (N4630, N4617, N3213);
and AND3 (N4631, N4614, N795, N4132);
nor NOR4 (N4632, N4620, N3447, N523, N1058);
not NOT1 (N4633, N4623);
nor NOR2 (N4634, N4624, N2949);
and AND3 (N4635, N4611, N3670, N672);
or OR4 (N4636, N4631, N2893, N4612, N4423);
nand NAND2 (N4637, N4632, N2674);
buf BUF1 (N4638, N4629);
buf BUF1 (N4639, N4625);
and AND2 (N4640, N4627, N2865);
and AND4 (N4641, N4640, N1916, N2037, N1946);
xor XOR2 (N4642, N4636, N2980);
not NOT1 (N4643, N4638);
nor NOR3 (N4644, N4628, N3744, N4546);
nand NAND2 (N4645, N4630, N2306);
xor XOR2 (N4646, N4642, N1428);
nor NOR3 (N4647, N4643, N1718, N2552);
not NOT1 (N4648, N4634);
nor NOR4 (N4649, N4633, N4258, N2420, N4345);
nor NOR4 (N4650, N4639, N4631, N4479, N2609);
and AND4 (N4651, N4648, N2220, N1608, N1692);
not NOT1 (N4652, N4650);
buf BUF1 (N4653, N4651);
or OR3 (N4654, N4641, N3563, N3246);
nand NAND4 (N4655, N4637, N3983, N1892, N3075);
not NOT1 (N4656, N4647);
xor XOR2 (N4657, N4646, N3841);
xor XOR2 (N4658, N4635, N3508);
nand NAND3 (N4659, N4655, N1249, N1195);
nand NAND4 (N4660, N4659, N4222, N2148, N2368);
buf BUF1 (N4661, N4654);
buf BUF1 (N4662, N4645);
xor XOR2 (N4663, N4652, N3736);
or OR4 (N4664, N4649, N4205, N19, N3524);
buf BUF1 (N4665, N4664);
xor XOR2 (N4666, N4658, N1353);
and AND4 (N4667, N4661, N2729, N41, N2553);
xor XOR2 (N4668, N4657, N4575);
nand NAND3 (N4669, N4662, N1010, N3063);
xor XOR2 (N4670, N4656, N1996);
or OR4 (N4671, N4666, N2368, N3035, N625);
or OR3 (N4672, N4669, N1779, N1553);
not NOT1 (N4673, N4663);
and AND3 (N4674, N4673, N3066, N4524);
or OR2 (N4675, N4644, N3463);
xor XOR2 (N4676, N4675, N4393);
buf BUF1 (N4677, N4674);
nor NOR3 (N4678, N4660, N3371, N1861);
nor NOR4 (N4679, N4677, N463, N1557, N3889);
not NOT1 (N4680, N4653);
not NOT1 (N4681, N4680);
and AND4 (N4682, N4676, N4206, N3937, N2232);
not NOT1 (N4683, N4681);
not NOT1 (N4684, N4671);
buf BUF1 (N4685, N4667);
nor NOR4 (N4686, N4670, N2168, N1302, N1191);
nor NOR2 (N4687, N4682, N1441);
nor NOR2 (N4688, N4686, N4373);
or OR4 (N4689, N4672, N1834, N1550, N3164);
and AND3 (N4690, N4665, N3610, N2827);
nor NOR3 (N4691, N4668, N2291, N1459);
or OR4 (N4692, N4691, N31, N2158, N4197);
nor NOR3 (N4693, N4688, N2396, N2550);
nor NOR2 (N4694, N4679, N1983);
nand NAND2 (N4695, N4692, N432);
and AND4 (N4696, N4693, N4602, N3740, N1140);
buf BUF1 (N4697, N4687);
xor XOR2 (N4698, N4694, N2510);
and AND4 (N4699, N4697, N2983, N618, N4525);
buf BUF1 (N4700, N4683);
xor XOR2 (N4701, N4698, N1277);
or OR4 (N4702, N4701, N851, N4528, N2181);
or OR3 (N4703, N4702, N4211, N998);
nand NAND3 (N4704, N4690, N4691, N92);
not NOT1 (N4705, N4704);
and AND4 (N4706, N4696, N4318, N3881, N4128);
and AND3 (N4707, N4703, N2355, N2629);
xor XOR2 (N4708, N4695, N3656);
buf BUF1 (N4709, N4678);
xor XOR2 (N4710, N4705, N1641);
nor NOR4 (N4711, N4684, N4645, N4389, N4371);
xor XOR2 (N4712, N4685, N1084);
buf BUF1 (N4713, N4689);
buf BUF1 (N4714, N4709);
nor NOR4 (N4715, N4712, N1364, N2925, N3369);
not NOT1 (N4716, N4708);
nor NOR3 (N4717, N4699, N700, N964);
or OR4 (N4718, N4716, N340, N902, N1808);
xor XOR2 (N4719, N4706, N2213);
or OR2 (N4720, N4718, N3417);
nor NOR3 (N4721, N4713, N2091, N3643);
nor NOR3 (N4722, N4715, N4159, N2990);
not NOT1 (N4723, N4720);
nand NAND4 (N4724, N4710, N2694, N832, N2186);
not NOT1 (N4725, N4714);
xor XOR2 (N4726, N4717, N2881);
nand NAND3 (N4727, N4721, N2358, N3342);
or OR2 (N4728, N4719, N1881);
xor XOR2 (N4729, N4728, N322);
nand NAND2 (N4730, N4707, N2069);
nand NAND4 (N4731, N4729, N4109, N560, N900);
nand NAND2 (N4732, N4711, N4205);
or OR2 (N4733, N4722, N3324);
or OR3 (N4734, N4732, N2196, N1443);
nand NAND2 (N4735, N4731, N3586);
nor NOR3 (N4736, N4733, N314, N1978);
or OR2 (N4737, N4736, N2339);
and AND3 (N4738, N4727, N1977, N4442);
xor XOR2 (N4739, N4734, N4207);
nor NOR3 (N4740, N4739, N4387, N3006);
buf BUF1 (N4741, N4737);
buf BUF1 (N4742, N4741);
not NOT1 (N4743, N4735);
buf BUF1 (N4744, N4730);
buf BUF1 (N4745, N4700);
and AND3 (N4746, N4742, N1988, N3674);
nor NOR4 (N4747, N4746, N1028, N2484, N3158);
nand NAND2 (N4748, N4744, N575);
nand NAND4 (N4749, N4740, N1748, N2602, N2671);
nor NOR3 (N4750, N4749, N576, N2306);
not NOT1 (N4751, N4725);
or OR4 (N4752, N4748, N4683, N1121, N596);
nor NOR3 (N4753, N4724, N2443, N12);
buf BUF1 (N4754, N4726);
nor NOR3 (N4755, N4745, N3560, N1941);
not NOT1 (N4756, N4752);
xor XOR2 (N4757, N4723, N1652);
buf BUF1 (N4758, N4743);
not NOT1 (N4759, N4750);
or OR2 (N4760, N4756, N2525);
and AND3 (N4761, N4758, N405, N951);
nor NOR3 (N4762, N4759, N2330, N3307);
nor NOR3 (N4763, N4754, N3791, N4327);
xor XOR2 (N4764, N4757, N1751);
nand NAND4 (N4765, N4764, N516, N2084, N337);
buf BUF1 (N4766, N4751);
or OR2 (N4767, N4765, N3198);
buf BUF1 (N4768, N4766);
and AND4 (N4769, N4768, N2441, N1798, N1387);
xor XOR2 (N4770, N4747, N3027);
xor XOR2 (N4771, N4753, N507);
nand NAND4 (N4772, N4771, N1401, N233, N4130);
nor NOR4 (N4773, N4761, N3753, N4062, N4269);
nor NOR3 (N4774, N4762, N3695, N3659);
xor XOR2 (N4775, N4774, N4166);
xor XOR2 (N4776, N4760, N2048);
nor NOR3 (N4777, N4770, N4016, N2894);
nand NAND4 (N4778, N4773, N3471, N3326, N4554);
buf BUF1 (N4779, N4776);
and AND4 (N4780, N4777, N2392, N89, N3165);
and AND2 (N4781, N4755, N177);
and AND4 (N4782, N4772, N2923, N4148, N277);
xor XOR2 (N4783, N4778, N2457);
xor XOR2 (N4784, N4767, N636);
buf BUF1 (N4785, N4763);
xor XOR2 (N4786, N4779, N2148);
nand NAND4 (N4787, N4780, N814, N3131, N481);
not NOT1 (N4788, N4786);
nand NAND3 (N4789, N4783, N3009, N1407);
nor NOR4 (N4790, N4782, N2545, N4464, N2908);
nand NAND4 (N4791, N4785, N3383, N1244, N1360);
xor XOR2 (N4792, N4775, N2090);
buf BUF1 (N4793, N4787);
and AND2 (N4794, N4781, N3565);
buf BUF1 (N4795, N4791);
or OR2 (N4796, N4792, N1176);
not NOT1 (N4797, N4790);
or OR2 (N4798, N4784, N3956);
xor XOR2 (N4799, N4797, N4405);
and AND3 (N4800, N4789, N436, N3174);
nor NOR2 (N4801, N4795, N1320);
and AND3 (N4802, N4788, N1502, N2714);
or OR3 (N4803, N4802, N922, N3400);
nor NOR4 (N4804, N4796, N1543, N2065, N2253);
xor XOR2 (N4805, N4801, N1367);
or OR3 (N4806, N4805, N2755, N1012);
buf BUF1 (N4807, N4738);
nor NOR4 (N4808, N4806, N4024, N2873, N2765);
xor XOR2 (N4809, N4807, N2315);
or OR2 (N4810, N4809, N1905);
nor NOR3 (N4811, N4800, N3803, N2790);
not NOT1 (N4812, N4794);
nor NOR2 (N4813, N4810, N4170);
or OR2 (N4814, N4803, N2477);
nor NOR2 (N4815, N4793, N750);
and AND4 (N4816, N4811, N531, N3403, N4545);
and AND3 (N4817, N4815, N1111, N4698);
xor XOR2 (N4818, N4814, N1277);
or OR2 (N4819, N4769, N2964);
or OR2 (N4820, N4798, N1803);
and AND3 (N4821, N4816, N1242, N1679);
xor XOR2 (N4822, N4820, N4774);
nand NAND3 (N4823, N4813, N4017, N3619);
or OR2 (N4824, N4812, N1449);
or OR4 (N4825, N4808, N4678, N624, N4033);
buf BUF1 (N4826, N4825);
or OR2 (N4827, N4819, N3025);
nor NOR3 (N4828, N4818, N1931, N1694);
xor XOR2 (N4829, N4824, N4567);
nor NOR3 (N4830, N4823, N950, N618);
nand NAND4 (N4831, N4826, N2609, N771, N3124);
nor NOR4 (N4832, N4827, N2258, N2228, N4797);
buf BUF1 (N4833, N4821);
nand NAND2 (N4834, N4829, N2911);
or OR2 (N4835, N4799, N803);
or OR3 (N4836, N4831, N4495, N1672);
and AND4 (N4837, N4828, N3457, N675, N1862);
and AND4 (N4838, N4837, N1747, N1544, N2586);
and AND2 (N4839, N4832, N4300);
xor XOR2 (N4840, N4833, N621);
and AND2 (N4841, N4822, N3896);
not NOT1 (N4842, N4840);
or OR3 (N4843, N4835, N1802, N3734);
or OR3 (N4844, N4841, N4057, N3030);
nand NAND4 (N4845, N4842, N513, N1770, N3278);
not NOT1 (N4846, N4817);
buf BUF1 (N4847, N4834);
not NOT1 (N4848, N4843);
nor NOR3 (N4849, N4804, N660, N558);
buf BUF1 (N4850, N4846);
buf BUF1 (N4851, N4850);
nor NOR2 (N4852, N4847, N3505);
not NOT1 (N4853, N4851);
nand NAND2 (N4854, N4852, N81);
buf BUF1 (N4855, N4853);
not NOT1 (N4856, N4844);
not NOT1 (N4857, N4855);
nand NAND4 (N4858, N4854, N1269, N2019, N3068);
and AND2 (N4859, N4858, N1752);
and AND3 (N4860, N4830, N4382, N1095);
not NOT1 (N4861, N4848);
and AND3 (N4862, N4849, N1471, N2252);
nor NOR3 (N4863, N4845, N4746, N4526);
xor XOR2 (N4864, N4857, N3012);
nand NAND3 (N4865, N4861, N344, N1153);
and AND4 (N4866, N4863, N1255, N495, N2264);
buf BUF1 (N4867, N4865);
or OR3 (N4868, N4867, N3963, N1555);
nand NAND3 (N4869, N4836, N2220, N3613);
xor XOR2 (N4870, N4868, N4812);
or OR3 (N4871, N4869, N2025, N487);
not NOT1 (N4872, N4870);
or OR2 (N4873, N4860, N1255);
and AND4 (N4874, N4873, N1111, N3166, N2315);
buf BUF1 (N4875, N4838);
xor XOR2 (N4876, N4871, N280);
and AND3 (N4877, N4864, N2322, N4639);
nor NOR3 (N4878, N4872, N4545, N2396);
not NOT1 (N4879, N4874);
and AND3 (N4880, N4877, N4149, N872);
nand NAND4 (N4881, N4839, N4495, N661, N3849);
xor XOR2 (N4882, N4859, N3077);
nor NOR2 (N4883, N4880, N174);
buf BUF1 (N4884, N4875);
or OR4 (N4885, N4884, N728, N611, N3332);
xor XOR2 (N4886, N4878, N939);
xor XOR2 (N4887, N4876, N2725);
and AND3 (N4888, N4856, N4784, N1729);
nor NOR3 (N4889, N4862, N1073, N2669);
xor XOR2 (N4890, N4889, N45);
nand NAND4 (N4891, N4888, N1547, N4295, N2303);
or OR2 (N4892, N4890, N1075);
and AND3 (N4893, N4882, N2833, N1650);
xor XOR2 (N4894, N4886, N4234);
or OR2 (N4895, N4879, N2239);
xor XOR2 (N4896, N4887, N2783);
nand NAND4 (N4897, N4891, N339, N4694, N4095);
and AND3 (N4898, N4892, N347, N2925);
nand NAND3 (N4899, N4896, N2865, N176);
nor NOR2 (N4900, N4899, N4370);
buf BUF1 (N4901, N4900);
buf BUF1 (N4902, N4898);
and AND3 (N4903, N4883, N3196, N3841);
not NOT1 (N4904, N4901);
or OR2 (N4905, N4894, N3919);
nand NAND2 (N4906, N4905, N2817);
nand NAND2 (N4907, N4897, N3612);
or OR4 (N4908, N4866, N1724, N1801, N4227);
or OR4 (N4909, N4904, N718, N2658, N3391);
or OR3 (N4910, N4881, N3919, N4381);
not NOT1 (N4911, N4893);
and AND2 (N4912, N4909, N1358);
not NOT1 (N4913, N4910);
not NOT1 (N4914, N4908);
buf BUF1 (N4915, N4895);
buf BUF1 (N4916, N4911);
nand NAND2 (N4917, N4913, N306);
or OR2 (N4918, N4916, N368);
and AND3 (N4919, N4917, N2804, N3103);
buf BUF1 (N4920, N4918);
xor XOR2 (N4921, N4906, N4886);
xor XOR2 (N4922, N4903, N1579);
and AND3 (N4923, N4912, N4303, N4096);
xor XOR2 (N4924, N4885, N156);
xor XOR2 (N4925, N4902, N3620);
not NOT1 (N4926, N4914);
xor XOR2 (N4927, N4926, N48);
nor NOR2 (N4928, N4921, N1609);
and AND3 (N4929, N4920, N495, N3484);
nand NAND2 (N4930, N4907, N776);
nand NAND3 (N4931, N4928, N3958, N2150);
and AND4 (N4932, N4930, N3826, N4078, N3915);
nor NOR4 (N4933, N4923, N4238, N3422, N1814);
buf BUF1 (N4934, N4932);
buf BUF1 (N4935, N4933);
not NOT1 (N4936, N4935);
or OR4 (N4937, N4922, N1581, N1875, N2037);
nor NOR4 (N4938, N4919, N1965, N4265, N4100);
nand NAND2 (N4939, N4929, N2179);
not NOT1 (N4940, N4927);
buf BUF1 (N4941, N4925);
and AND2 (N4942, N4941, N4177);
buf BUF1 (N4943, N4937);
or OR3 (N4944, N4940, N134, N1892);
nor NOR2 (N4945, N4936, N1467);
nand NAND2 (N4946, N4939, N4448);
and AND2 (N4947, N4931, N3960);
not NOT1 (N4948, N4924);
not NOT1 (N4949, N4942);
not NOT1 (N4950, N4948);
nand NAND2 (N4951, N4944, N1439);
xor XOR2 (N4952, N4947, N2565);
not NOT1 (N4953, N4934);
buf BUF1 (N4954, N4943);
not NOT1 (N4955, N4951);
xor XOR2 (N4956, N4949, N2703);
xor XOR2 (N4957, N4954, N4405);
or OR3 (N4958, N4957, N1434, N913);
and AND4 (N4959, N4915, N24, N4830, N546);
not NOT1 (N4960, N4956);
not NOT1 (N4961, N4953);
and AND4 (N4962, N4945, N4013, N3819, N2930);
xor XOR2 (N4963, N4961, N1391);
xor XOR2 (N4964, N4952, N3290);
nand NAND2 (N4965, N4950, N3051);
or OR4 (N4966, N4964, N3627, N2668, N4267);
nor NOR4 (N4967, N4960, N744, N3680, N477);
or OR3 (N4968, N4962, N3452, N2150);
nor NOR4 (N4969, N4963, N3776, N452, N4465);
not NOT1 (N4970, N4946);
nor NOR4 (N4971, N4959, N30, N3527, N1181);
and AND2 (N4972, N4968, N1301);
and AND2 (N4973, N4971, N178);
buf BUF1 (N4974, N4965);
nand NAND2 (N4975, N4974, N1023);
nor NOR2 (N4976, N4966, N2717);
or OR3 (N4977, N4967, N2210, N755);
or OR4 (N4978, N4977, N2537, N2178, N799);
and AND3 (N4979, N4938, N1410, N3358);
buf BUF1 (N4980, N4972);
nand NAND4 (N4981, N4978, N3626, N2272, N3872);
nand NAND3 (N4982, N4981, N2689, N1047);
not NOT1 (N4983, N4976);
and AND4 (N4984, N4973, N972, N1449, N4882);
or OR2 (N4985, N4980, N2564);
nor NOR4 (N4986, N4979, N3333, N2336, N2214);
not NOT1 (N4987, N4955);
nor NOR3 (N4988, N4986, N3326, N4596);
and AND3 (N4989, N4975, N1440, N81);
buf BUF1 (N4990, N4969);
nor NOR4 (N4991, N4970, N914, N1751, N849);
and AND2 (N4992, N4983, N4429);
or OR4 (N4993, N4985, N393, N3871, N1233);
nor NOR4 (N4994, N4992, N2520, N3212, N866);
and AND3 (N4995, N4990, N1825, N3648);
or OR3 (N4996, N4993, N4423, N3263);
not NOT1 (N4997, N4982);
not NOT1 (N4998, N4987);
xor XOR2 (N4999, N4997, N3493);
nor NOR3 (N5000, N4958, N4351, N2978);
nand NAND2 (N5001, N4984, N902);
buf BUF1 (N5002, N4994);
nor NOR4 (N5003, N4989, N860, N1587, N186);
xor XOR2 (N5004, N5001, N2973);
nand NAND3 (N5005, N5004, N4101, N1650);
xor XOR2 (N5006, N5002, N778);
nand NAND2 (N5007, N4996, N383);
buf BUF1 (N5008, N4998);
xor XOR2 (N5009, N4999, N2888);
not NOT1 (N5010, N4991);
nor NOR4 (N5011, N5009, N3946, N652, N3342);
or OR2 (N5012, N5005, N2520);
and AND4 (N5013, N4988, N4176, N2550, N5012);
or OR3 (N5014, N5002, N4610, N1739);
and AND3 (N5015, N5010, N4857, N2424);
not NOT1 (N5016, N5003);
xor XOR2 (N5017, N5013, N3982);
nor NOR4 (N5018, N5016, N1456, N5012, N3874);
buf BUF1 (N5019, N5007);
buf BUF1 (N5020, N5018);
or OR3 (N5021, N5020, N3724, N3658);
nand NAND4 (N5022, N4995, N1180, N3128, N4033);
nand NAND4 (N5023, N5011, N3236, N4729, N10);
or OR2 (N5024, N5008, N2343);
nor NOR4 (N5025, N5006, N4810, N1169, N1740);
nand NAND2 (N5026, N5023, N2262);
not NOT1 (N5027, N5015);
xor XOR2 (N5028, N5017, N597);
buf BUF1 (N5029, N5026);
nand NAND4 (N5030, N5019, N2706, N1087, N3024);
nor NOR2 (N5031, N5022, N3591);
buf BUF1 (N5032, N5030);
not NOT1 (N5033, N5014);
nand NAND2 (N5034, N5033, N369);
or OR4 (N5035, N5029, N625, N3791, N1906);
not NOT1 (N5036, N5028);
and AND2 (N5037, N5024, N4613);
nor NOR4 (N5038, N5037, N4573, N2008, N1669);
not NOT1 (N5039, N5000);
not NOT1 (N5040, N5039);
or OR3 (N5041, N5036, N3090, N3941);
nor NOR2 (N5042, N5040, N4436);
not NOT1 (N5043, N5032);
xor XOR2 (N5044, N5043, N4028);
buf BUF1 (N5045, N5041);
or OR2 (N5046, N5042, N1545);
not NOT1 (N5047, N5046);
xor XOR2 (N5048, N5045, N4569);
buf BUF1 (N5049, N5027);
buf BUF1 (N5050, N5038);
nor NOR4 (N5051, N5025, N4097, N1645, N4917);
not NOT1 (N5052, N5044);
xor XOR2 (N5053, N5047, N618);
xor XOR2 (N5054, N5035, N4600);
or OR2 (N5055, N5034, N1956);
buf BUF1 (N5056, N5050);
nand NAND3 (N5057, N5048, N3622, N190);
nor NOR4 (N5058, N5057, N1128, N2234, N1304);
or OR4 (N5059, N5021, N2304, N3966, N1590);
not NOT1 (N5060, N5058);
not NOT1 (N5061, N5060);
xor XOR2 (N5062, N5053, N2272);
xor XOR2 (N5063, N5052, N1280);
not NOT1 (N5064, N5056);
nand NAND4 (N5065, N5064, N3125, N3234, N4251);
not NOT1 (N5066, N5065);
buf BUF1 (N5067, N5061);
or OR3 (N5068, N5063, N2210, N3861);
nor NOR4 (N5069, N5062, N1470, N354, N4056);
buf BUF1 (N5070, N5049);
not NOT1 (N5071, N5051);
and AND2 (N5072, N5071, N2543);
nor NOR3 (N5073, N5054, N28, N1455);
xor XOR2 (N5074, N5069, N2137);
nor NOR4 (N5075, N5055, N2934, N3485, N209);
nor NOR2 (N5076, N5068, N1288);
nand NAND4 (N5077, N5067, N1007, N401, N2467);
nand NAND2 (N5078, N5076, N2880);
nand NAND3 (N5079, N5077, N4618, N1811);
and AND2 (N5080, N5031, N2416);
nand NAND3 (N5081, N5066, N210, N547);
not NOT1 (N5082, N5075);
and AND3 (N5083, N5082, N4195, N2870);
not NOT1 (N5084, N5079);
nor NOR4 (N5085, N5074, N4833, N3012, N1275);
buf BUF1 (N5086, N5084);
nor NOR2 (N5087, N5072, N1047);
xor XOR2 (N5088, N5073, N4064);
not NOT1 (N5089, N5080);
and AND4 (N5090, N5059, N814, N2758, N1553);
buf BUF1 (N5091, N5085);
buf BUF1 (N5092, N5070);
nor NOR4 (N5093, N5088, N2240, N3454, N395);
or OR2 (N5094, N5083, N2401);
xor XOR2 (N5095, N5081, N2908);
nand NAND2 (N5096, N5090, N1211);
nand NAND4 (N5097, N5086, N2757, N4165, N2396);
not NOT1 (N5098, N5087);
and AND3 (N5099, N5092, N4085, N1881);
buf BUF1 (N5100, N5098);
and AND4 (N5101, N5078, N4362, N4075, N4738);
nand NAND2 (N5102, N5099, N2432);
nand NAND2 (N5103, N5101, N1221);
buf BUF1 (N5104, N5097);
nor NOR3 (N5105, N5091, N5049, N4979);
xor XOR2 (N5106, N5104, N2391);
and AND2 (N5107, N5106, N4123);
or OR2 (N5108, N5105, N2881);
xor XOR2 (N5109, N5102, N3877);
buf BUF1 (N5110, N5089);
or OR4 (N5111, N5107, N138, N3371, N2679);
and AND3 (N5112, N5096, N1239, N408);
xor XOR2 (N5113, N5093, N4478);
nor NOR3 (N5114, N5113, N1032, N3904);
xor XOR2 (N5115, N5100, N3590);
xor XOR2 (N5116, N5110, N4687);
nor NOR3 (N5117, N5108, N3065, N2536);
nand NAND2 (N5118, N5103, N1360);
buf BUF1 (N5119, N5109);
xor XOR2 (N5120, N5115, N19);
xor XOR2 (N5121, N5119, N3782);
or OR4 (N5122, N5116, N3723, N4159, N3648);
or OR2 (N5123, N5121, N4744);
nor NOR2 (N5124, N5117, N3755);
not NOT1 (N5125, N5118);
xor XOR2 (N5126, N5111, N2671);
or OR4 (N5127, N5112, N3021, N4054, N4829);
xor XOR2 (N5128, N5126, N2139);
nand NAND2 (N5129, N5094, N485);
not NOT1 (N5130, N5129);
xor XOR2 (N5131, N5114, N2268);
nor NOR2 (N5132, N5124, N1280);
buf BUF1 (N5133, N5123);
xor XOR2 (N5134, N5133, N3530);
nor NOR3 (N5135, N5120, N4768, N4668);
xor XOR2 (N5136, N5125, N500);
or OR3 (N5137, N5136, N909, N2541);
nand NAND3 (N5138, N5137, N4586, N1172);
not NOT1 (N5139, N5128);
not NOT1 (N5140, N5138);
not NOT1 (N5141, N5135);
nand NAND2 (N5142, N5132, N4592);
buf BUF1 (N5143, N5134);
xor XOR2 (N5144, N5142, N2516);
xor XOR2 (N5145, N5140, N2360);
buf BUF1 (N5146, N5143);
or OR3 (N5147, N5095, N3798, N3951);
xor XOR2 (N5148, N5127, N2775);
nor NOR4 (N5149, N5147, N3659, N2781, N4746);
or OR3 (N5150, N5148, N1218, N4202);
not NOT1 (N5151, N5150);
or OR4 (N5152, N5149, N224, N2921, N3971);
not NOT1 (N5153, N5139);
buf BUF1 (N5154, N5144);
nand NAND4 (N5155, N5151, N3614, N4454, N476);
or OR2 (N5156, N5155, N335);
nor NOR2 (N5157, N5130, N4027);
nand NAND4 (N5158, N5156, N1392, N3458, N3223);
and AND4 (N5159, N5153, N830, N3985, N332);
xor XOR2 (N5160, N5154, N720);
nor NOR2 (N5161, N5122, N252);
nor NOR2 (N5162, N5145, N172);
nand NAND4 (N5163, N5159, N3765, N3244, N3300);
nand NAND3 (N5164, N5146, N2286, N2373);
and AND2 (N5165, N5163, N1378);
nand NAND3 (N5166, N5158, N3320, N3364);
xor XOR2 (N5167, N5152, N3180);
and AND3 (N5168, N5164, N3146, N2984);
nand NAND2 (N5169, N5141, N5118);
or OR4 (N5170, N5169, N3612, N1803, N1222);
and AND2 (N5171, N5160, N1185);
and AND2 (N5172, N5131, N2743);
nor NOR4 (N5173, N5157, N3385, N4706, N1942);
and AND3 (N5174, N5165, N2957, N4662);
and AND4 (N5175, N5166, N3758, N4338, N2566);
not NOT1 (N5176, N5172);
nor NOR2 (N5177, N5161, N3250);
and AND4 (N5178, N5171, N39, N741, N4956);
nor NOR2 (N5179, N5168, N4010);
and AND4 (N5180, N5178, N4232, N3415, N3442);
or OR4 (N5181, N5175, N3251, N1828, N3649);
nor NOR3 (N5182, N5177, N2002, N525);
and AND2 (N5183, N5162, N20);
buf BUF1 (N5184, N5180);
not NOT1 (N5185, N5167);
not NOT1 (N5186, N5185);
xor XOR2 (N5187, N5170, N3332);
xor XOR2 (N5188, N5176, N4097);
xor XOR2 (N5189, N5184, N260);
nand NAND3 (N5190, N5173, N4758, N3488);
and AND3 (N5191, N5183, N4645, N3757);
and AND3 (N5192, N5190, N1656, N2962);
and AND3 (N5193, N5192, N524, N43);
nor NOR4 (N5194, N5179, N1035, N317, N1238);
and AND4 (N5195, N5191, N3432, N1261, N2816);
buf BUF1 (N5196, N5188);
and AND4 (N5197, N5193, N3427, N2677, N5005);
nor NOR3 (N5198, N5187, N3213, N2549);
and AND2 (N5199, N5181, N5074);
and AND2 (N5200, N5196, N2338);
xor XOR2 (N5201, N5182, N2063);
nor NOR4 (N5202, N5197, N1392, N2431, N2781);
or OR2 (N5203, N5200, N439);
nand NAND4 (N5204, N5194, N4477, N923, N5154);
or OR3 (N5205, N5186, N2106, N1210);
not NOT1 (N5206, N5198);
and AND3 (N5207, N5205, N4248, N4560);
and AND2 (N5208, N5204, N3242);
not NOT1 (N5209, N5207);
or OR2 (N5210, N5189, N4681);
xor XOR2 (N5211, N5209, N4249);
nand NAND2 (N5212, N5211, N940);
nor NOR3 (N5213, N5195, N198, N4321);
or OR2 (N5214, N5202, N3087);
nor NOR4 (N5215, N5174, N2377, N2262, N1529);
xor XOR2 (N5216, N5208, N2009);
and AND2 (N5217, N5203, N4476);
buf BUF1 (N5218, N5212);
and AND2 (N5219, N5217, N4930);
or OR2 (N5220, N5218, N296);
and AND4 (N5221, N5213, N3039, N1888, N1432);
buf BUF1 (N5222, N5214);
and AND2 (N5223, N5220, N910);
xor XOR2 (N5224, N5199, N2671);
xor XOR2 (N5225, N5216, N2885);
nor NOR3 (N5226, N5224, N4405, N732);
nand NAND3 (N5227, N5210, N1191, N2163);
buf BUF1 (N5228, N5227);
nand NAND4 (N5229, N5228, N3161, N3030, N4292);
nor NOR4 (N5230, N5206, N1068, N5148, N1578);
not NOT1 (N5231, N5223);
or OR4 (N5232, N5201, N437, N2295, N4243);
or OR4 (N5233, N5221, N2643, N2957, N4373);
and AND2 (N5234, N5230, N699);
or OR2 (N5235, N5225, N89);
xor XOR2 (N5236, N5215, N3683);
or OR3 (N5237, N5231, N2217, N3605);
not NOT1 (N5238, N5235);
buf BUF1 (N5239, N5237);
not NOT1 (N5240, N5222);
not NOT1 (N5241, N5229);
nor NOR3 (N5242, N5241, N3285, N780);
buf BUF1 (N5243, N5226);
and AND4 (N5244, N5238, N1652, N672, N4244);
nand NAND3 (N5245, N5243, N833, N1339);
nor NOR2 (N5246, N5219, N2236);
xor XOR2 (N5247, N5246, N2838);
or OR4 (N5248, N5240, N4635, N2594, N4770);
nor NOR4 (N5249, N5248, N5114, N3099, N1089);
buf BUF1 (N5250, N5249);
nor NOR2 (N5251, N5244, N2151);
xor XOR2 (N5252, N5236, N912);
buf BUF1 (N5253, N5252);
nand NAND2 (N5254, N5232, N4992);
buf BUF1 (N5255, N5239);
buf BUF1 (N5256, N5251);
not NOT1 (N5257, N5242);
and AND2 (N5258, N5250, N4284);
and AND2 (N5259, N5255, N1257);
buf BUF1 (N5260, N5257);
or OR3 (N5261, N5245, N4249, N4694);
buf BUF1 (N5262, N5234);
or OR4 (N5263, N5260, N3103, N943, N911);
xor XOR2 (N5264, N5256, N3270);
and AND4 (N5265, N5254, N5221, N1179, N1582);
xor XOR2 (N5266, N5253, N974);
buf BUF1 (N5267, N5263);
and AND4 (N5268, N5266, N3576, N4253, N1074);
or OR3 (N5269, N5259, N964, N1408);
and AND2 (N5270, N5261, N3534);
not NOT1 (N5271, N5270);
buf BUF1 (N5272, N5268);
nand NAND3 (N5273, N5272, N530, N3401);
or OR4 (N5274, N5233, N1711, N4125, N4635);
nor NOR4 (N5275, N5269, N1796, N468, N1069);
buf BUF1 (N5276, N5258);
or OR2 (N5277, N5262, N4623);
or OR3 (N5278, N5277, N2359, N4862);
buf BUF1 (N5279, N5274);
nand NAND2 (N5280, N5275, N2212);
xor XOR2 (N5281, N5271, N821);
buf BUF1 (N5282, N5280);
nor NOR4 (N5283, N5282, N3898, N3409, N2763);
or OR3 (N5284, N5279, N3508, N1093);
xor XOR2 (N5285, N5283, N4088);
and AND2 (N5286, N5267, N1203);
nand NAND4 (N5287, N5284, N3569, N722, N4261);
buf BUF1 (N5288, N5285);
nor NOR3 (N5289, N5276, N3196, N2502);
buf BUF1 (N5290, N5287);
nand NAND4 (N5291, N5286, N4840, N3935, N1373);
or OR3 (N5292, N5291, N220, N2192);
or OR3 (N5293, N5281, N1278, N3790);
not NOT1 (N5294, N5289);
and AND2 (N5295, N5278, N1021);
not NOT1 (N5296, N5292);
and AND4 (N5297, N5294, N3878, N3993, N3044);
or OR3 (N5298, N5295, N281, N5224);
nand NAND2 (N5299, N5288, N2094);
and AND2 (N5300, N5265, N3174);
not NOT1 (N5301, N5264);
xor XOR2 (N5302, N5247, N4507);
not NOT1 (N5303, N5290);
buf BUF1 (N5304, N5296);
not NOT1 (N5305, N5303);
nor NOR2 (N5306, N5298, N744);
buf BUF1 (N5307, N5293);
nor NOR2 (N5308, N5307, N3996);
buf BUF1 (N5309, N5301);
buf BUF1 (N5310, N5305);
xor XOR2 (N5311, N5273, N1457);
and AND2 (N5312, N5306, N1799);
or OR3 (N5313, N5311, N814, N1548);
or OR4 (N5314, N5310, N4774, N1030, N2640);
not NOT1 (N5315, N5313);
not NOT1 (N5316, N5308);
and AND3 (N5317, N5309, N1957, N1519);
not NOT1 (N5318, N5312);
xor XOR2 (N5319, N5300, N1665);
nand NAND3 (N5320, N5297, N1374, N532);
and AND4 (N5321, N5315, N2132, N2080, N1311);
or OR4 (N5322, N5302, N3626, N1209, N1535);
nor NOR4 (N5323, N5321, N4112, N1573, N20);
xor XOR2 (N5324, N5299, N4384);
xor XOR2 (N5325, N5323, N3405);
or OR4 (N5326, N5319, N1632, N5104, N4843);
not NOT1 (N5327, N5304);
not NOT1 (N5328, N5314);
nor NOR2 (N5329, N5318, N5126);
xor XOR2 (N5330, N5328, N728);
nor NOR4 (N5331, N5317, N5104, N2350, N5313);
buf BUF1 (N5332, N5329);
or OR2 (N5333, N5327, N3011);
nor NOR4 (N5334, N5332, N928, N2548, N894);
and AND4 (N5335, N5333, N2464, N2506, N4306);
and AND4 (N5336, N5320, N1830, N967, N5073);
not NOT1 (N5337, N5326);
xor XOR2 (N5338, N5335, N3807);
and AND4 (N5339, N5322, N2107, N4135, N4551);
nor NOR2 (N5340, N5325, N2597);
xor XOR2 (N5341, N5338, N3463);
nand NAND2 (N5342, N5334, N3745);
or OR4 (N5343, N5342, N2081, N4156, N303);
or OR4 (N5344, N5341, N175, N4783, N2081);
or OR2 (N5345, N5336, N447);
buf BUF1 (N5346, N5331);
nor NOR2 (N5347, N5330, N3083);
nor NOR3 (N5348, N5346, N5256, N1490);
nand NAND3 (N5349, N5340, N4730, N2380);
or OR4 (N5350, N5349, N3417, N3619, N3451);
and AND4 (N5351, N5350, N1635, N3168, N3404);
xor XOR2 (N5352, N5339, N2560);
buf BUF1 (N5353, N5316);
nor NOR4 (N5354, N5337, N60, N4080, N983);
or OR4 (N5355, N5352, N693, N4049, N4019);
nand NAND2 (N5356, N5353, N1053);
and AND2 (N5357, N5344, N2834);
not NOT1 (N5358, N5357);
nor NOR4 (N5359, N5348, N17, N3510, N1374);
nor NOR4 (N5360, N5345, N2880, N195, N2377);
and AND3 (N5361, N5356, N729, N2264);
nand NAND2 (N5362, N5361, N3548);
xor XOR2 (N5363, N5362, N148);
nand NAND3 (N5364, N5360, N1801, N564);
not NOT1 (N5365, N5355);
xor XOR2 (N5366, N5363, N4249);
buf BUF1 (N5367, N5358);
nor NOR4 (N5368, N5343, N1497, N3664, N1882);
not NOT1 (N5369, N5351);
not NOT1 (N5370, N5359);
buf BUF1 (N5371, N5347);
or OR3 (N5372, N5371, N703, N277);
nor NOR3 (N5373, N5365, N4858, N1367);
buf BUF1 (N5374, N5370);
nand NAND2 (N5375, N5324, N1752);
and AND2 (N5376, N5364, N1834);
xor XOR2 (N5377, N5367, N1740);
xor XOR2 (N5378, N5375, N3133);
xor XOR2 (N5379, N5372, N2582);
not NOT1 (N5380, N5374);
nand NAND3 (N5381, N5380, N4234, N3475);
nand NAND2 (N5382, N5373, N4921);
buf BUF1 (N5383, N5368);
nand NAND3 (N5384, N5379, N5003, N1592);
buf BUF1 (N5385, N5366);
xor XOR2 (N5386, N5376, N3525);
not NOT1 (N5387, N5386);
nor NOR3 (N5388, N5383, N3006, N1503);
nand NAND2 (N5389, N5369, N3255);
not NOT1 (N5390, N5378);
nor NOR3 (N5391, N5387, N2526, N4064);
and AND4 (N5392, N5391, N1387, N2852, N3494);
nor NOR2 (N5393, N5392, N4061);
xor XOR2 (N5394, N5388, N4311);
xor XOR2 (N5395, N5377, N4048);
nor NOR4 (N5396, N5389, N3959, N3004, N2357);
nor NOR4 (N5397, N5354, N144, N3124, N575);
nor NOR4 (N5398, N5395, N2775, N4973, N4710);
and AND2 (N5399, N5396, N2770);
xor XOR2 (N5400, N5390, N2012);
buf BUF1 (N5401, N5382);
nand NAND3 (N5402, N5385, N18, N642);
or OR2 (N5403, N5393, N5138);
and AND2 (N5404, N5403, N4677);
not NOT1 (N5405, N5404);
nor NOR2 (N5406, N5398, N904);
nor NOR4 (N5407, N5394, N2840, N4730, N1442);
or OR4 (N5408, N5384, N2648, N2232, N1965);
buf BUF1 (N5409, N5405);
nand NAND2 (N5410, N5381, N1763);
buf BUF1 (N5411, N5399);
nand NAND4 (N5412, N5402, N5110, N1887, N1193);
or OR3 (N5413, N5407, N2230, N1751);
or OR2 (N5414, N5412, N641);
nor NOR2 (N5415, N5401, N5067);
or OR2 (N5416, N5410, N3796);
and AND2 (N5417, N5406, N4248);
nor NOR3 (N5418, N5408, N3564, N1203);
buf BUF1 (N5419, N5414);
nand NAND4 (N5420, N5418, N4312, N3386, N2044);
or OR3 (N5421, N5397, N4641, N1520);
nand NAND2 (N5422, N5409, N3823);
not NOT1 (N5423, N5420);
xor XOR2 (N5424, N5411, N180);
or OR4 (N5425, N5423, N5396, N2915, N3557);
buf BUF1 (N5426, N5421);
buf BUF1 (N5427, N5419);
not NOT1 (N5428, N5426);
and AND4 (N5429, N5422, N713, N1014, N4654);
or OR3 (N5430, N5416, N2525, N752);
nand NAND4 (N5431, N5417, N1451, N2753, N3378);
buf BUF1 (N5432, N5429);
or OR3 (N5433, N5431, N148, N1305);
nand NAND2 (N5434, N5400, N2320);
and AND2 (N5435, N5413, N3316);
xor XOR2 (N5436, N5427, N3947);
buf BUF1 (N5437, N5433);
xor XOR2 (N5438, N5425, N595);
and AND3 (N5439, N5430, N1183, N3934);
or OR3 (N5440, N5437, N132, N3261);
or OR3 (N5441, N5432, N5082, N815);
and AND4 (N5442, N5439, N198, N2295, N854);
not NOT1 (N5443, N5440);
not NOT1 (N5444, N5442);
and AND4 (N5445, N5444, N40, N2142, N3821);
xor XOR2 (N5446, N5436, N925);
nand NAND2 (N5447, N5434, N5151);
not NOT1 (N5448, N5445);
and AND2 (N5449, N5415, N4082);
buf BUF1 (N5450, N5424);
buf BUF1 (N5451, N5443);
not NOT1 (N5452, N5441);
nand NAND3 (N5453, N5446, N3694, N2532);
xor XOR2 (N5454, N5438, N3450);
buf BUF1 (N5455, N5435);
nor NOR3 (N5456, N5428, N1855, N3453);
or OR4 (N5457, N5452, N5002, N1411, N4070);
buf BUF1 (N5458, N5453);
buf BUF1 (N5459, N5455);
nand NAND2 (N5460, N5456, N5079);
not NOT1 (N5461, N5454);
xor XOR2 (N5462, N5459, N4582);
and AND2 (N5463, N5448, N470);
not NOT1 (N5464, N5449);
not NOT1 (N5465, N5462);
and AND4 (N5466, N5447, N2226, N3614, N1628);
xor XOR2 (N5467, N5451, N921);
buf BUF1 (N5468, N5450);
buf BUF1 (N5469, N5460);
nand NAND3 (N5470, N5463, N3370, N1141);
nand NAND3 (N5471, N5467, N953, N1718);
nand NAND3 (N5472, N5468, N2568, N467);
nor NOR3 (N5473, N5471, N3580, N4145);
not NOT1 (N5474, N5473);
or OR3 (N5475, N5458, N4278, N310);
nand NAND3 (N5476, N5472, N1246, N316);
xor XOR2 (N5477, N5457, N1373);
nand NAND4 (N5478, N5470, N606, N1969, N1214);
buf BUF1 (N5479, N5461);
xor XOR2 (N5480, N5478, N2309);
and AND2 (N5481, N5475, N4351);
xor XOR2 (N5482, N5474, N2339);
nor NOR3 (N5483, N5465, N5408, N4755);
nor NOR3 (N5484, N5476, N4858, N4293);
nand NAND4 (N5485, N5481, N1942, N1183, N2066);
and AND4 (N5486, N5485, N3413, N2528, N2664);
nand NAND4 (N5487, N5477, N340, N38, N4550);
nand NAND3 (N5488, N5484, N5308, N846);
xor XOR2 (N5489, N5469, N4282);
buf BUF1 (N5490, N5479);
and AND4 (N5491, N5489, N173, N5020, N957);
not NOT1 (N5492, N5491);
or OR3 (N5493, N5480, N2222, N1545);
buf BUF1 (N5494, N5483);
nand NAND4 (N5495, N5487, N822, N730, N1271);
buf BUF1 (N5496, N5493);
xor XOR2 (N5497, N5464, N2262);
not NOT1 (N5498, N5492);
or OR4 (N5499, N5496, N4318, N3329, N5073);
and AND3 (N5500, N5488, N1117, N140);
not NOT1 (N5501, N5486);
buf BUF1 (N5502, N5490);
nor NOR2 (N5503, N5500, N4142);
and AND2 (N5504, N5503, N1830);
or OR3 (N5505, N5504, N103, N3980);
not NOT1 (N5506, N5495);
and AND4 (N5507, N5466, N4339, N4154, N951);
not NOT1 (N5508, N5494);
not NOT1 (N5509, N5501);
and AND2 (N5510, N5507, N5481);
buf BUF1 (N5511, N5482);
xor XOR2 (N5512, N5509, N1569);
not NOT1 (N5513, N5499);
xor XOR2 (N5514, N5510, N2327);
xor XOR2 (N5515, N5497, N4334);
nor NOR4 (N5516, N5513, N2084, N4956, N4112);
xor XOR2 (N5517, N5516, N3731);
and AND2 (N5518, N5505, N5127);
and AND2 (N5519, N5515, N1695);
or OR3 (N5520, N5508, N5442, N3820);
xor XOR2 (N5521, N5520, N51);
nor NOR3 (N5522, N5502, N1532, N926);
xor XOR2 (N5523, N5512, N4175);
nor NOR4 (N5524, N5522, N4670, N2486, N4876);
and AND3 (N5525, N5524, N1234, N4477);
not NOT1 (N5526, N5498);
not NOT1 (N5527, N5517);
xor XOR2 (N5528, N5525, N1843);
not NOT1 (N5529, N5523);
xor XOR2 (N5530, N5528, N3729);
nor NOR3 (N5531, N5519, N1029, N3441);
buf BUF1 (N5532, N5521);
or OR2 (N5533, N5532, N3804);
or OR3 (N5534, N5529, N219, N540);
buf BUF1 (N5535, N5534);
nand NAND2 (N5536, N5527, N986);
nor NOR2 (N5537, N5531, N999);
and AND2 (N5538, N5533, N231);
nor NOR2 (N5539, N5536, N3782);
or OR2 (N5540, N5514, N4611);
nor NOR2 (N5541, N5506, N4127);
xor XOR2 (N5542, N5511, N2671);
buf BUF1 (N5543, N5538);
and AND3 (N5544, N5540, N2223, N4744);
and AND4 (N5545, N5543, N2296, N4821, N3759);
buf BUF1 (N5546, N5545);
or OR3 (N5547, N5539, N608, N1772);
or OR3 (N5548, N5530, N5066, N2699);
not NOT1 (N5549, N5537);
and AND4 (N5550, N5526, N1376, N2270, N435);
buf BUF1 (N5551, N5546);
nor NOR4 (N5552, N5547, N5192, N258, N5536);
buf BUF1 (N5553, N5550);
or OR4 (N5554, N5542, N3400, N3471, N5493);
xor XOR2 (N5555, N5552, N2784);
buf BUF1 (N5556, N5535);
nor NOR4 (N5557, N5556, N532, N822, N5092);
xor XOR2 (N5558, N5554, N3238);
nor NOR2 (N5559, N5548, N4503);
or OR4 (N5560, N5518, N3169, N2004, N5238);
or OR4 (N5561, N5541, N3306, N5367, N4003);
buf BUF1 (N5562, N5559);
not NOT1 (N5563, N5549);
buf BUF1 (N5564, N5560);
xor XOR2 (N5565, N5561, N4235);
xor XOR2 (N5566, N5555, N456);
not NOT1 (N5567, N5558);
xor XOR2 (N5568, N5553, N3017);
and AND4 (N5569, N5565, N2539, N3859, N2421);
not NOT1 (N5570, N5551);
buf BUF1 (N5571, N5563);
buf BUF1 (N5572, N5557);
buf BUF1 (N5573, N5571);
or OR4 (N5574, N5569, N1121, N97, N2128);
or OR2 (N5575, N5572, N4907);
not NOT1 (N5576, N5574);
xor XOR2 (N5577, N5566, N4796);
and AND4 (N5578, N5544, N3009, N4445, N1768);
and AND3 (N5579, N5562, N2003, N4133);
nor NOR3 (N5580, N5570, N108, N3763);
and AND4 (N5581, N5568, N2722, N5108, N1324);
nor NOR4 (N5582, N5573, N4336, N4495, N2411);
and AND4 (N5583, N5564, N674, N4675, N114);
not NOT1 (N5584, N5581);
not NOT1 (N5585, N5576);
buf BUF1 (N5586, N5575);
buf BUF1 (N5587, N5580);
not NOT1 (N5588, N5579);
buf BUF1 (N5589, N5584);
or OR2 (N5590, N5583, N2521);
and AND3 (N5591, N5589, N1589, N4640);
nand NAND4 (N5592, N5567, N177, N276, N3049);
nor NOR4 (N5593, N5587, N4927, N922, N3556);
not NOT1 (N5594, N5592);
xor XOR2 (N5595, N5594, N4286);
or OR3 (N5596, N5591, N4209, N2447);
nand NAND4 (N5597, N5585, N2141, N5338, N651);
buf BUF1 (N5598, N5578);
nand NAND3 (N5599, N5598, N1087, N5485);
nand NAND2 (N5600, N5588, N2034);
and AND4 (N5601, N5596, N4659, N3585, N2001);
nor NOR2 (N5602, N5599, N87);
and AND4 (N5603, N5590, N1816, N844, N3949);
not NOT1 (N5604, N5603);
and AND4 (N5605, N5593, N792, N2945, N5364);
and AND2 (N5606, N5577, N5267);
nand NAND2 (N5607, N5601, N2523);
not NOT1 (N5608, N5600);
nand NAND3 (N5609, N5605, N3325, N779);
or OR3 (N5610, N5595, N1695, N1079);
xor XOR2 (N5611, N5604, N483);
or OR2 (N5612, N5582, N2150);
xor XOR2 (N5613, N5612, N4814);
or OR4 (N5614, N5586, N2937, N3112, N5349);
nand NAND3 (N5615, N5611, N61, N3410);
nor NOR2 (N5616, N5610, N902);
or OR2 (N5617, N5607, N385);
or OR4 (N5618, N5606, N4758, N2660, N3743);
nand NAND2 (N5619, N5597, N3264);
buf BUF1 (N5620, N5614);
xor XOR2 (N5621, N5608, N2677);
nor NOR4 (N5622, N5609, N3741, N3078, N788);
nor NOR3 (N5623, N5616, N2664, N3509);
not NOT1 (N5624, N5615);
or OR4 (N5625, N5618, N215, N4905, N3786);
and AND3 (N5626, N5625, N3991, N362);
and AND4 (N5627, N5621, N3149, N4195, N232);
nor NOR4 (N5628, N5617, N1654, N3142, N1523);
xor XOR2 (N5629, N5624, N2068);
buf BUF1 (N5630, N5628);
xor XOR2 (N5631, N5623, N4762);
nor NOR3 (N5632, N5629, N1324, N232);
or OR4 (N5633, N5602, N2414, N222, N1527);
nor NOR2 (N5634, N5633, N3667);
not NOT1 (N5635, N5613);
and AND4 (N5636, N5635, N4533, N3290, N2242);
and AND3 (N5637, N5620, N876, N102);
nor NOR3 (N5638, N5631, N863, N1305);
nand NAND4 (N5639, N5637, N1032, N86, N780);
xor XOR2 (N5640, N5632, N4378);
nor NOR3 (N5641, N5626, N1605, N736);
or OR2 (N5642, N5627, N5429);
or OR2 (N5643, N5641, N537);
xor XOR2 (N5644, N5638, N3902);
nand NAND4 (N5645, N5644, N1741, N662, N716);
buf BUF1 (N5646, N5634);
nand NAND2 (N5647, N5622, N3073);
nor NOR4 (N5648, N5640, N4416, N3172, N3864);
buf BUF1 (N5649, N5630);
nand NAND3 (N5650, N5649, N3743, N2053);
not NOT1 (N5651, N5619);
or OR4 (N5652, N5642, N178, N827, N2852);
not NOT1 (N5653, N5647);
and AND4 (N5654, N5650, N3402, N5524, N5131);
nand NAND2 (N5655, N5639, N3244);
buf BUF1 (N5656, N5654);
buf BUF1 (N5657, N5656);
xor XOR2 (N5658, N5646, N4132);
nand NAND3 (N5659, N5655, N3054, N839);
or OR4 (N5660, N5645, N4734, N5348, N2368);
nand NAND3 (N5661, N5657, N1035, N4126);
nor NOR3 (N5662, N5651, N4394, N1370);
not NOT1 (N5663, N5652);
buf BUF1 (N5664, N5658);
or OR3 (N5665, N5648, N1204, N1696);
xor XOR2 (N5666, N5662, N2426);
nand NAND4 (N5667, N5643, N2273, N4446, N3095);
nand NAND2 (N5668, N5660, N3088);
nand NAND3 (N5669, N5666, N4216, N1360);
not NOT1 (N5670, N5668);
buf BUF1 (N5671, N5661);
nand NAND2 (N5672, N5653, N4498);
buf BUF1 (N5673, N5670);
and AND3 (N5674, N5659, N1688, N3494);
nand NAND3 (N5675, N5667, N1428, N2318);
or OR3 (N5676, N5671, N4046, N3288);
nand NAND2 (N5677, N5675, N3332);
nand NAND3 (N5678, N5664, N3545, N3358);
nor NOR4 (N5679, N5676, N2141, N4420, N976);
not NOT1 (N5680, N5636);
and AND2 (N5681, N5665, N5151);
buf BUF1 (N5682, N5680);
not NOT1 (N5683, N5673);
not NOT1 (N5684, N5677);
nor NOR3 (N5685, N5672, N3030, N4805);
xor XOR2 (N5686, N5674, N5527);
or OR3 (N5687, N5678, N2662, N708);
xor XOR2 (N5688, N5686, N2811);
not NOT1 (N5689, N5681);
xor XOR2 (N5690, N5684, N1026);
buf BUF1 (N5691, N5685);
nor NOR4 (N5692, N5682, N262, N389, N3440);
xor XOR2 (N5693, N5688, N1152);
and AND2 (N5694, N5691, N5396);
nand NAND2 (N5695, N5692, N1880);
nor NOR3 (N5696, N5663, N1230, N1028);
buf BUF1 (N5697, N5669);
and AND2 (N5698, N5689, N4347);
xor XOR2 (N5699, N5687, N3749);
nand NAND3 (N5700, N5679, N4050, N3057);
or OR2 (N5701, N5695, N5619);
or OR3 (N5702, N5700, N1632, N246);
nand NAND3 (N5703, N5690, N5695, N3033);
or OR4 (N5704, N5699, N424, N2479, N1093);
and AND3 (N5705, N5696, N1401, N4835);
xor XOR2 (N5706, N5703, N5698);
or OR3 (N5707, N5356, N1150, N4824);
xor XOR2 (N5708, N5706, N2622);
nand NAND4 (N5709, N5701, N2765, N4222, N3149);
nand NAND4 (N5710, N5702, N441, N4668, N5407);
not NOT1 (N5711, N5708);
nand NAND4 (N5712, N5694, N3218, N3328, N2260);
and AND4 (N5713, N5710, N4061, N5683, N2640);
xor XOR2 (N5714, N3281, N3133);
xor XOR2 (N5715, N5711, N201);
nor NOR2 (N5716, N5712, N4669);
nor NOR2 (N5717, N5715, N2517);
nor NOR2 (N5718, N5705, N1144);
and AND2 (N5719, N5717, N419);
not NOT1 (N5720, N5718);
buf BUF1 (N5721, N5697);
nand NAND3 (N5722, N5709, N4571, N4628);
buf BUF1 (N5723, N5719);
nand NAND4 (N5724, N5704, N3975, N4891, N5446);
or OR2 (N5725, N5724, N3795);
xor XOR2 (N5726, N5713, N2312);
or OR4 (N5727, N5716, N3379, N71, N2286);
nor NOR4 (N5728, N5727, N5512, N1975, N2264);
or OR2 (N5729, N5728, N5488);
and AND2 (N5730, N5721, N1491);
xor XOR2 (N5731, N5722, N5334);
or OR3 (N5732, N5730, N5326, N2476);
or OR3 (N5733, N5731, N3323, N23);
not NOT1 (N5734, N5725);
not NOT1 (N5735, N5734);
or OR2 (N5736, N5733, N1250);
or OR2 (N5737, N5729, N5069);
nand NAND2 (N5738, N5737, N3070);
not NOT1 (N5739, N5707);
buf BUF1 (N5740, N5714);
buf BUF1 (N5741, N5738);
xor XOR2 (N5742, N5720, N2539);
and AND3 (N5743, N5739, N5452, N2372);
not NOT1 (N5744, N5742);
and AND2 (N5745, N5723, N613);
xor XOR2 (N5746, N5693, N632);
nand NAND4 (N5747, N5744, N4921, N904, N5416);
nor NOR3 (N5748, N5736, N2276, N2090);
nor NOR3 (N5749, N5732, N3888, N2879);
and AND3 (N5750, N5735, N1478, N955);
and AND2 (N5751, N5746, N2361);
not NOT1 (N5752, N5748);
not NOT1 (N5753, N5751);
xor XOR2 (N5754, N5745, N3675);
nor NOR2 (N5755, N5754, N1864);
nor NOR2 (N5756, N5740, N1733);
and AND4 (N5757, N5741, N2625, N3044, N5355);
nand NAND2 (N5758, N5752, N127);
not NOT1 (N5759, N5755);
nor NOR3 (N5760, N5747, N5053, N3596);
or OR4 (N5761, N5756, N5326, N3737, N5668);
not NOT1 (N5762, N5743);
not NOT1 (N5763, N5757);
nor NOR2 (N5764, N5749, N4937);
xor XOR2 (N5765, N5750, N4571);
or OR4 (N5766, N5760, N5550, N4744, N5575);
xor XOR2 (N5767, N5764, N2090);
and AND2 (N5768, N5726, N32);
not NOT1 (N5769, N5759);
nand NAND4 (N5770, N5753, N1208, N3662, N3895);
and AND4 (N5771, N5762, N1064, N1288, N1777);
nand NAND2 (N5772, N5763, N5716);
xor XOR2 (N5773, N5772, N2517);
xor XOR2 (N5774, N5773, N5323);
not NOT1 (N5775, N5767);
or OR2 (N5776, N5769, N3589);
nand NAND4 (N5777, N5776, N5643, N1953, N2584);
nand NAND2 (N5778, N5765, N1494);
not NOT1 (N5779, N5771);
not NOT1 (N5780, N5768);
and AND4 (N5781, N5758, N1776, N2069, N337);
or OR3 (N5782, N5781, N2129, N431);
nor NOR4 (N5783, N5766, N2762, N108, N2922);
buf BUF1 (N5784, N5780);
or OR4 (N5785, N5777, N5588, N2685, N4306);
not NOT1 (N5786, N5761);
nor NOR4 (N5787, N5784, N5438, N1368, N2176);
not NOT1 (N5788, N5786);
xor XOR2 (N5789, N5774, N3585);
nand NAND4 (N5790, N5787, N5142, N4428, N4669);
not NOT1 (N5791, N5788);
and AND4 (N5792, N5783, N4390, N4823, N3366);
not NOT1 (N5793, N5782);
nor NOR3 (N5794, N5791, N2881, N2287);
and AND2 (N5795, N5778, N2393);
nand NAND3 (N5796, N5775, N2845, N790);
nand NAND2 (N5797, N5794, N1322);
nor NOR3 (N5798, N5770, N1168, N5716);
xor XOR2 (N5799, N5795, N2407);
not NOT1 (N5800, N5792);
nand NAND2 (N5801, N5796, N1093);
nor NOR2 (N5802, N5801, N5117);
xor XOR2 (N5803, N5789, N3101);
not NOT1 (N5804, N5798);
xor XOR2 (N5805, N5803, N496);
buf BUF1 (N5806, N5785);
not NOT1 (N5807, N5793);
buf BUF1 (N5808, N5799);
and AND3 (N5809, N5779, N429, N5043);
nor NOR4 (N5810, N5809, N4296, N1653, N4231);
xor XOR2 (N5811, N5805, N4417);
nor NOR4 (N5812, N5797, N4943, N539, N670);
buf BUF1 (N5813, N5811);
or OR3 (N5814, N5804, N82, N1325);
nor NOR2 (N5815, N5813, N3899);
buf BUF1 (N5816, N5807);
nor NOR4 (N5817, N5816, N4890, N2478, N4152);
nor NOR4 (N5818, N5806, N1874, N1877, N5714);
not NOT1 (N5819, N5817);
not NOT1 (N5820, N5815);
xor XOR2 (N5821, N5808, N1041);
and AND3 (N5822, N5790, N696, N3698);
xor XOR2 (N5823, N5810, N3743);
or OR3 (N5824, N5819, N410, N424);
buf BUF1 (N5825, N5802);
buf BUF1 (N5826, N5825);
and AND4 (N5827, N5812, N4716, N2752, N2254);
buf BUF1 (N5828, N5827);
buf BUF1 (N5829, N5821);
and AND4 (N5830, N5826, N1735, N3895, N2345);
or OR3 (N5831, N5800, N312, N2104);
nor NOR3 (N5832, N5831, N2415, N764);
and AND3 (N5833, N5820, N2578, N1531);
or OR2 (N5834, N5814, N2573);
not NOT1 (N5835, N5818);
xor XOR2 (N5836, N5833, N4102);
not NOT1 (N5837, N5836);
buf BUF1 (N5838, N5824);
buf BUF1 (N5839, N5838);
nor NOR3 (N5840, N5835, N5478, N3996);
and AND2 (N5841, N5837, N716);
not NOT1 (N5842, N5830);
buf BUF1 (N5843, N5839);
nand NAND2 (N5844, N5841, N444);
buf BUF1 (N5845, N5842);
xor XOR2 (N5846, N5844, N4154);
or OR2 (N5847, N5840, N147);
and AND2 (N5848, N5828, N885);
xor XOR2 (N5849, N5823, N4400);
and AND2 (N5850, N5846, N1681);
and AND2 (N5851, N5845, N5770);
buf BUF1 (N5852, N5822);
buf BUF1 (N5853, N5851);
buf BUF1 (N5854, N5832);
or OR3 (N5855, N5849, N455, N1919);
not NOT1 (N5856, N5847);
buf BUF1 (N5857, N5855);
and AND2 (N5858, N5834, N3798);
buf BUF1 (N5859, N5854);
xor XOR2 (N5860, N5858, N3046);
not NOT1 (N5861, N5856);
nor NOR2 (N5862, N5848, N1463);
or OR4 (N5863, N5860, N1792, N2098, N3066);
nand NAND2 (N5864, N5857, N396);
nor NOR2 (N5865, N5863, N4483);
nand NAND4 (N5866, N5852, N3374, N2871, N1522);
nand NAND3 (N5867, N5850, N3631, N4563);
and AND4 (N5868, N5843, N4795, N2856, N3475);
nor NOR2 (N5869, N5867, N36);
or OR4 (N5870, N5861, N5436, N5577, N3162);
buf BUF1 (N5871, N5829);
nor NOR2 (N5872, N5866, N376);
buf BUF1 (N5873, N5864);
or OR4 (N5874, N5865, N5374, N5722, N231);
nand NAND3 (N5875, N5869, N1279, N485);
or OR4 (N5876, N5853, N2814, N549, N2440);
and AND3 (N5877, N5870, N3616, N4511);
nor NOR2 (N5878, N5876, N1797);
and AND2 (N5879, N5874, N5346);
xor XOR2 (N5880, N5871, N5023);
buf BUF1 (N5881, N5859);
or OR3 (N5882, N5868, N4929, N4856);
and AND4 (N5883, N5875, N4253, N677, N986);
or OR4 (N5884, N5880, N4373, N3853, N4172);
buf BUF1 (N5885, N5872);
buf BUF1 (N5886, N5862);
xor XOR2 (N5887, N5873, N55);
or OR3 (N5888, N5879, N4264, N5830);
not NOT1 (N5889, N5885);
not NOT1 (N5890, N5883);
not NOT1 (N5891, N5889);
xor XOR2 (N5892, N5881, N5085);
or OR3 (N5893, N5888, N5278, N5796);
xor XOR2 (N5894, N5884, N4608);
and AND4 (N5895, N5891, N5886, N4408, N1061);
buf BUF1 (N5896, N1589);
and AND3 (N5897, N5893, N3023, N3539);
and AND3 (N5898, N5896, N4336, N3293);
not NOT1 (N5899, N5892);
nand NAND2 (N5900, N5890, N1563);
nand NAND3 (N5901, N5895, N4408, N522);
xor XOR2 (N5902, N5898, N4533);
nand NAND4 (N5903, N5894, N5654, N4273, N3624);
nor NOR4 (N5904, N5899, N4930, N5107, N2201);
and AND4 (N5905, N5897, N5708, N4721, N3424);
nor NOR2 (N5906, N5900, N4330);
or OR3 (N5907, N5903, N3900, N649);
buf BUF1 (N5908, N5878);
or OR3 (N5909, N5905, N5797, N834);
xor XOR2 (N5910, N5909, N2385);
buf BUF1 (N5911, N5904);
nand NAND3 (N5912, N5908, N2667, N4321);
not NOT1 (N5913, N5907);
nor NOR2 (N5914, N5887, N410);
buf BUF1 (N5915, N5901);
nor NOR2 (N5916, N5913, N939);
buf BUF1 (N5917, N5906);
nand NAND3 (N5918, N5917, N5619, N3945);
buf BUF1 (N5919, N5914);
nor NOR4 (N5920, N5877, N553, N4484, N5566);
or OR4 (N5921, N5911, N4258, N5148, N354);
and AND4 (N5922, N5882, N2051, N5850, N2543);
nor NOR2 (N5923, N5922, N967);
not NOT1 (N5924, N5920);
xor XOR2 (N5925, N5902, N5202);
buf BUF1 (N5926, N5924);
nand NAND4 (N5927, N5923, N5309, N5534, N3284);
xor XOR2 (N5928, N5925, N919);
nand NAND4 (N5929, N5915, N4925, N3498, N4421);
xor XOR2 (N5930, N5919, N5687);
and AND2 (N5931, N5916, N3999);
or OR3 (N5932, N5921, N3411, N1024);
and AND3 (N5933, N5926, N4392, N5301);
or OR4 (N5934, N5912, N1774, N1712, N2329);
xor XOR2 (N5935, N5927, N4618);
and AND3 (N5936, N5935, N3265, N2355);
nor NOR4 (N5937, N5932, N4475, N3685, N1805);
xor XOR2 (N5938, N5933, N2626);
not NOT1 (N5939, N5938);
and AND3 (N5940, N5910, N3656, N571);
not NOT1 (N5941, N5934);
xor XOR2 (N5942, N5941, N154);
buf BUF1 (N5943, N5942);
and AND3 (N5944, N5931, N828, N2434);
and AND4 (N5945, N5936, N3482, N1255, N769);
not NOT1 (N5946, N5945);
nand NAND4 (N5947, N5944, N5109, N3690, N173);
buf BUF1 (N5948, N5940);
not NOT1 (N5949, N5943);
nand NAND3 (N5950, N5948, N2245, N617);
not NOT1 (N5951, N5949);
nor NOR4 (N5952, N5937, N3244, N2455, N3711);
xor XOR2 (N5953, N5918, N848);
nand NAND2 (N5954, N5930, N1636);
not NOT1 (N5955, N5947);
buf BUF1 (N5956, N5952);
buf BUF1 (N5957, N5928);
xor XOR2 (N5958, N5957, N3188);
nor NOR3 (N5959, N5950, N5586, N5932);
buf BUF1 (N5960, N5929);
and AND2 (N5961, N5959, N4845);
buf BUF1 (N5962, N5951);
buf BUF1 (N5963, N5946);
nor NOR3 (N5964, N5958, N738, N1059);
nand NAND4 (N5965, N5955, N1436, N1816, N3419);
not NOT1 (N5966, N5964);
nand NAND2 (N5967, N5966, N3570);
xor XOR2 (N5968, N5953, N3732);
xor XOR2 (N5969, N5967, N3876);
nand NAND3 (N5970, N5962, N1823, N4372);
and AND2 (N5971, N5965, N4051);
buf BUF1 (N5972, N5956);
and AND2 (N5973, N5961, N674);
or OR4 (N5974, N5954, N8, N4865, N4566);
nand NAND2 (N5975, N5974, N462);
or OR4 (N5976, N5968, N1245, N33, N4321);
or OR2 (N5977, N5969, N3661);
xor XOR2 (N5978, N5963, N1251);
nand NAND3 (N5979, N5960, N22, N3676);
and AND2 (N5980, N5975, N1100);
nand NAND4 (N5981, N5973, N3058, N2310, N766);
nor NOR2 (N5982, N5970, N2467);
nand NAND3 (N5983, N5980, N4922, N2141);
buf BUF1 (N5984, N5977);
or OR4 (N5985, N5972, N3975, N5908, N5511);
and AND3 (N5986, N5984, N2504, N4011);
and AND3 (N5987, N5976, N222, N482);
and AND4 (N5988, N5971, N3498, N3456, N3479);
xor XOR2 (N5989, N5979, N2273);
not NOT1 (N5990, N5987);
or OR4 (N5991, N5989, N1373, N2346, N5677);
buf BUF1 (N5992, N5978);
xor XOR2 (N5993, N5992, N4980);
nor NOR4 (N5994, N5985, N972, N2580, N3622);
not NOT1 (N5995, N5986);
nor NOR2 (N5996, N5983, N4908);
xor XOR2 (N5997, N5995, N1567);
not NOT1 (N5998, N5991);
and AND3 (N5999, N5990, N1984, N2820);
nand NAND3 (N6000, N5994, N1697, N4971);
not NOT1 (N6001, N5996);
or OR4 (N6002, N6000, N1460, N5186, N4912);
or OR2 (N6003, N6001, N1331);
nor NOR2 (N6004, N5993, N5818);
buf BUF1 (N6005, N5997);
xor XOR2 (N6006, N5982, N1984);
buf BUF1 (N6007, N6002);
nor NOR4 (N6008, N6005, N5341, N703, N2280);
nand NAND2 (N6009, N5999, N3630);
nor NOR2 (N6010, N5988, N763);
nor NOR3 (N6011, N6010, N919, N5725);
nor NOR2 (N6012, N6006, N608);
xor XOR2 (N6013, N5939, N4789);
and AND4 (N6014, N5998, N2315, N870, N1750);
or OR4 (N6015, N6012, N4164, N1202, N303);
and AND4 (N6016, N6008, N4462, N1285, N4587);
nand NAND4 (N6017, N6009, N4325, N3634, N2413);
or OR3 (N6018, N6007, N3297, N1795);
buf BUF1 (N6019, N6011);
nand NAND4 (N6020, N6019, N4021, N5559, N3121);
or OR2 (N6021, N6015, N4886);
or OR4 (N6022, N6020, N1151, N2597, N707);
nand NAND3 (N6023, N6013, N3146, N1422);
xor XOR2 (N6024, N6003, N211);
nor NOR2 (N6025, N6004, N1894);
buf BUF1 (N6026, N6024);
and AND2 (N6027, N6016, N3015);
xor XOR2 (N6028, N6021, N945);
or OR3 (N6029, N6018, N4640, N5048);
nand NAND4 (N6030, N6029, N5693, N3281, N1797);
nor NOR4 (N6031, N6028, N4950, N2258, N4113);
buf BUF1 (N6032, N6023);
xor XOR2 (N6033, N6032, N1909);
xor XOR2 (N6034, N6025, N1197);
buf BUF1 (N6035, N6014);
nor NOR4 (N6036, N6026, N392, N3623, N3136);
xor XOR2 (N6037, N6031, N2451);
buf BUF1 (N6038, N6027);
and AND3 (N6039, N6030, N547, N4362);
nor NOR2 (N6040, N6037, N2221);
and AND4 (N6041, N6033, N2182, N1782, N5398);
nand NAND3 (N6042, N6041, N1078, N3727);
and AND4 (N6043, N6035, N4085, N557, N918);
nand NAND2 (N6044, N6042, N4003);
and AND2 (N6045, N6043, N3150);
buf BUF1 (N6046, N6017);
xor XOR2 (N6047, N6036, N426);
nor NOR2 (N6048, N6040, N739);
or OR3 (N6049, N6048, N4512, N3807);
buf BUF1 (N6050, N5981);
nand NAND2 (N6051, N6049, N1225);
not NOT1 (N6052, N6050);
and AND4 (N6053, N6022, N4121, N2276, N3034);
and AND2 (N6054, N6044, N1790);
nor NOR3 (N6055, N6053, N2386, N4799);
xor XOR2 (N6056, N6047, N4905);
buf BUF1 (N6057, N6051);
or OR2 (N6058, N6052, N5763);
xor XOR2 (N6059, N6034, N3508);
buf BUF1 (N6060, N6039);
or OR4 (N6061, N6056, N3756, N285, N4350);
and AND2 (N6062, N6057, N3689);
nor NOR4 (N6063, N6038, N2586, N1645, N4539);
and AND4 (N6064, N6060, N2734, N3963, N4629);
not NOT1 (N6065, N6055);
or OR4 (N6066, N6061, N2821, N3144, N2496);
or OR3 (N6067, N6066, N211, N4085);
nand NAND3 (N6068, N6045, N3025, N717);
and AND4 (N6069, N6058, N382, N475, N558);
not NOT1 (N6070, N6067);
xor XOR2 (N6071, N6065, N4592);
xor XOR2 (N6072, N6063, N2030);
and AND4 (N6073, N6069, N5030, N950, N3740);
and AND2 (N6074, N6072, N3204);
or OR4 (N6075, N6074, N1373, N2617, N4611);
or OR4 (N6076, N6075, N1761, N198, N4875);
or OR4 (N6077, N6068, N2862, N682, N484);
xor XOR2 (N6078, N6046, N3743);
and AND4 (N6079, N6059, N5319, N477, N5069);
and AND4 (N6080, N6070, N2616, N3103, N2095);
or OR3 (N6081, N6062, N1227, N404);
or OR3 (N6082, N6076, N2502, N1013);
buf BUF1 (N6083, N6078);
not NOT1 (N6084, N6082);
not NOT1 (N6085, N6081);
and AND4 (N6086, N6054, N5637, N5007, N1033);
and AND3 (N6087, N6084, N2081, N2711);
not NOT1 (N6088, N6080);
buf BUF1 (N6089, N6079);
nor NOR3 (N6090, N6071, N797, N2235);
nor NOR3 (N6091, N6088, N4161, N1901);
or OR3 (N6092, N6090, N2849, N1236);
xor XOR2 (N6093, N6064, N90);
not NOT1 (N6094, N6087);
nand NAND4 (N6095, N6092, N4113, N3792, N5754);
not NOT1 (N6096, N6073);
and AND2 (N6097, N6083, N3792);
or OR2 (N6098, N6077, N3352);
or OR2 (N6099, N6097, N1183);
nor NOR2 (N6100, N6086, N3900);
not NOT1 (N6101, N6089);
xor XOR2 (N6102, N6099, N1275);
buf BUF1 (N6103, N6091);
buf BUF1 (N6104, N6095);
not NOT1 (N6105, N6096);
nor NOR4 (N6106, N6101, N5875, N368, N6067);
or OR3 (N6107, N6102, N1577, N2993);
nor NOR2 (N6108, N6100, N678);
buf BUF1 (N6109, N6098);
buf BUF1 (N6110, N6104);
and AND2 (N6111, N6085, N3341);
and AND3 (N6112, N6109, N20, N858);
not NOT1 (N6113, N6103);
and AND2 (N6114, N6113, N4884);
nand NAND2 (N6115, N6108, N4887);
not NOT1 (N6116, N6093);
and AND4 (N6117, N6112, N1029, N5519, N3755);
not NOT1 (N6118, N6105);
nand NAND4 (N6119, N6117, N1051, N118, N4871);
not NOT1 (N6120, N6118);
nand NAND2 (N6121, N6116, N317);
buf BUF1 (N6122, N6094);
nand NAND3 (N6123, N6114, N717, N3400);
and AND3 (N6124, N6110, N5265, N1745);
buf BUF1 (N6125, N6106);
and AND2 (N6126, N6115, N4316);
and AND2 (N6127, N6107, N5406);
nor NOR4 (N6128, N6126, N639, N3875, N3113);
xor XOR2 (N6129, N6128, N920);
buf BUF1 (N6130, N6127);
nor NOR4 (N6131, N6124, N1658, N3227, N954);
nand NAND4 (N6132, N6121, N601, N3166, N1564);
nand NAND4 (N6133, N6123, N439, N5169, N5396);
and AND3 (N6134, N6132, N334, N2885);
xor XOR2 (N6135, N6111, N1144);
not NOT1 (N6136, N6133);
not NOT1 (N6137, N6130);
xor XOR2 (N6138, N6135, N3512);
xor XOR2 (N6139, N6125, N5477);
buf BUF1 (N6140, N6131);
nand NAND4 (N6141, N6129, N3971, N2068, N6015);
nand NAND3 (N6142, N6119, N1225, N4338);
nor NOR4 (N6143, N6138, N2079, N705, N5744);
not NOT1 (N6144, N6134);
or OR2 (N6145, N6141, N2643);
nand NAND3 (N6146, N6120, N3108, N4447);
nor NOR4 (N6147, N6122, N4257, N1281, N3723);
nor NOR4 (N6148, N6136, N4932, N1259, N1780);
and AND2 (N6149, N6147, N320);
buf BUF1 (N6150, N6143);
buf BUF1 (N6151, N6149);
nand NAND3 (N6152, N6137, N5455, N1242);
nand NAND2 (N6153, N6148, N5396);
nor NOR2 (N6154, N6151, N1329);
nand NAND4 (N6155, N6153, N1448, N5701, N1480);
nand NAND3 (N6156, N6142, N3600, N1228);
nand NAND3 (N6157, N6140, N5343, N4626);
nand NAND2 (N6158, N6156, N6058);
and AND2 (N6159, N6146, N5330);
or OR4 (N6160, N6158, N4005, N2867, N4207);
and AND3 (N6161, N6145, N5516, N828);
or OR2 (N6162, N6150, N1604);
nor NOR3 (N6163, N6157, N4171, N5991);
not NOT1 (N6164, N6163);
not NOT1 (N6165, N6152);
or OR2 (N6166, N6144, N3446);
or OR4 (N6167, N6154, N5315, N4201, N2640);
or OR2 (N6168, N6162, N4838);
nand NAND4 (N6169, N6159, N4391, N1601, N2231);
xor XOR2 (N6170, N6161, N3833);
xor XOR2 (N6171, N6168, N2093);
buf BUF1 (N6172, N6167);
nand NAND2 (N6173, N6165, N2056);
not NOT1 (N6174, N6173);
nand NAND3 (N6175, N6160, N5939, N1451);
nor NOR2 (N6176, N6166, N41);
nor NOR3 (N6177, N6139, N236, N904);
buf BUF1 (N6178, N6174);
buf BUF1 (N6179, N6172);
not NOT1 (N6180, N6176);
and AND2 (N6181, N6179, N5066);
nor NOR3 (N6182, N6169, N3022, N256);
nand NAND3 (N6183, N6171, N3674, N2343);
buf BUF1 (N6184, N6180);
or OR4 (N6185, N6170, N2396, N5680, N3519);
nand NAND2 (N6186, N6175, N3655);
not NOT1 (N6187, N6181);
buf BUF1 (N6188, N6183);
nand NAND4 (N6189, N6186, N115, N4036, N4087);
not NOT1 (N6190, N6155);
xor XOR2 (N6191, N6190, N2776);
xor XOR2 (N6192, N6188, N3450);
nand NAND4 (N6193, N6192, N2312, N5741, N259);
nand NAND3 (N6194, N6182, N230, N1286);
xor XOR2 (N6195, N6185, N3706);
nor NOR3 (N6196, N6178, N534, N3815);
not NOT1 (N6197, N6195);
buf BUF1 (N6198, N6164);
or OR4 (N6199, N6191, N1451, N4989, N1359);
and AND3 (N6200, N6199, N235, N3707);
and AND2 (N6201, N6198, N1770);
xor XOR2 (N6202, N6184, N5780);
xor XOR2 (N6203, N6189, N5113);
or OR4 (N6204, N6203, N4833, N240, N4816);
not NOT1 (N6205, N6187);
buf BUF1 (N6206, N6202);
not NOT1 (N6207, N6196);
buf BUF1 (N6208, N6201);
not NOT1 (N6209, N6204);
or OR2 (N6210, N6200, N5145);
xor XOR2 (N6211, N6209, N1847);
buf BUF1 (N6212, N6177);
or OR2 (N6213, N6197, N1709);
nand NAND2 (N6214, N6210, N4877);
buf BUF1 (N6215, N6207);
and AND2 (N6216, N6213, N988);
xor XOR2 (N6217, N6208, N2636);
not NOT1 (N6218, N6205);
and AND4 (N6219, N6217, N3904, N1670, N2317);
not NOT1 (N6220, N6215);
xor XOR2 (N6221, N6212, N6092);
and AND2 (N6222, N6219, N3231);
or OR2 (N6223, N6193, N4502);
xor XOR2 (N6224, N6206, N1690);
and AND4 (N6225, N6223, N1759, N4064, N1848);
buf BUF1 (N6226, N6225);
xor XOR2 (N6227, N6218, N2138);
or OR2 (N6228, N6194, N3848);
or OR2 (N6229, N6216, N5341);
not NOT1 (N6230, N6227);
or OR3 (N6231, N6226, N1069, N1643);
nand NAND3 (N6232, N6229, N1382, N4202);
nand NAND2 (N6233, N6228, N1759);
nor NOR4 (N6234, N6214, N5863, N4063, N4177);
not NOT1 (N6235, N6211);
nand NAND4 (N6236, N6222, N764, N2661, N3672);
or OR3 (N6237, N6233, N4970, N988);
nor NOR4 (N6238, N6236, N4864, N4383, N255);
not NOT1 (N6239, N6232);
nor NOR2 (N6240, N6221, N1719);
xor XOR2 (N6241, N6240, N3174);
nand NAND4 (N6242, N6241, N1036, N261, N2026);
or OR3 (N6243, N6242, N2901, N5886);
nand NAND2 (N6244, N6234, N5379);
or OR3 (N6245, N6235, N658, N1279);
xor XOR2 (N6246, N6243, N5758);
not NOT1 (N6247, N6246);
and AND2 (N6248, N6245, N2200);
nor NOR2 (N6249, N6237, N2713);
buf BUF1 (N6250, N6247);
not NOT1 (N6251, N6224);
buf BUF1 (N6252, N6248);
not NOT1 (N6253, N6231);
buf BUF1 (N6254, N6244);
or OR3 (N6255, N6252, N3628, N4227);
and AND4 (N6256, N6220, N4915, N4788, N2643);
nand NAND3 (N6257, N6250, N2548, N1939);
nand NAND2 (N6258, N6255, N605);
nand NAND3 (N6259, N6258, N3137, N3222);
nand NAND4 (N6260, N6239, N5236, N3018, N3872);
or OR2 (N6261, N6260, N2017);
nand NAND4 (N6262, N6238, N1356, N934, N2286);
not NOT1 (N6263, N6230);
nor NOR3 (N6264, N6249, N5222, N1746);
and AND4 (N6265, N6259, N2178, N2835, N4004);
buf BUF1 (N6266, N6251);
and AND2 (N6267, N6261, N632);
buf BUF1 (N6268, N6264);
and AND2 (N6269, N6268, N4085);
not NOT1 (N6270, N6254);
nor NOR2 (N6271, N6266, N1733);
nor NOR3 (N6272, N6269, N2659, N5770);
buf BUF1 (N6273, N6253);
nor NOR2 (N6274, N6272, N1386);
and AND2 (N6275, N6274, N5871);
or OR3 (N6276, N6273, N1161, N4729);
not NOT1 (N6277, N6257);
buf BUF1 (N6278, N6262);
nor NOR2 (N6279, N6265, N5691);
buf BUF1 (N6280, N6278);
xor XOR2 (N6281, N6270, N4912);
nand NAND2 (N6282, N6275, N1501);
nor NOR3 (N6283, N6279, N2892, N5992);
buf BUF1 (N6284, N6283);
and AND3 (N6285, N6256, N2760, N2819);
and AND2 (N6286, N6285, N2868);
not NOT1 (N6287, N6280);
nor NOR4 (N6288, N6276, N4708, N5794, N2180);
and AND4 (N6289, N6263, N2643, N4308, N1799);
nor NOR4 (N6290, N6282, N6165, N389, N1644);
not NOT1 (N6291, N6267);
or OR2 (N6292, N6287, N5220);
not NOT1 (N6293, N6288);
or OR2 (N6294, N6291, N4731);
and AND2 (N6295, N6294, N2970);
not NOT1 (N6296, N6293);
not NOT1 (N6297, N6271);
nand NAND3 (N6298, N6286, N1516, N405);
and AND2 (N6299, N6281, N737);
buf BUF1 (N6300, N6277);
and AND3 (N6301, N6292, N2579, N3243);
xor XOR2 (N6302, N6297, N2283);
not NOT1 (N6303, N6290);
nand NAND4 (N6304, N6295, N958, N6017, N5163);
nand NAND3 (N6305, N6298, N1396, N1097);
nand NAND3 (N6306, N6289, N3843, N3447);
buf BUF1 (N6307, N6301);
nand NAND3 (N6308, N6304, N1871, N2136);
buf BUF1 (N6309, N6300);
buf BUF1 (N6310, N6308);
buf BUF1 (N6311, N6302);
xor XOR2 (N6312, N6310, N3142);
nor NOR3 (N6313, N6296, N6251, N2052);
or OR4 (N6314, N6309, N2542, N802, N1474);
nor NOR3 (N6315, N6299, N2974, N267);
not NOT1 (N6316, N6314);
buf BUF1 (N6317, N6313);
and AND4 (N6318, N6312, N1736, N2883, N4341);
not NOT1 (N6319, N6315);
buf BUF1 (N6320, N6305);
nand NAND4 (N6321, N6316, N3287, N2139, N2790);
or OR4 (N6322, N6317, N2064, N6252, N448);
buf BUF1 (N6323, N6311);
or OR3 (N6324, N6306, N3906, N4135);
not NOT1 (N6325, N6323);
not NOT1 (N6326, N6303);
not NOT1 (N6327, N6321);
nor NOR4 (N6328, N6284, N5451, N4001, N4945);
nor NOR2 (N6329, N6324, N501);
xor XOR2 (N6330, N6307, N4327);
not NOT1 (N6331, N6319);
xor XOR2 (N6332, N6328, N3639);
xor XOR2 (N6333, N6327, N2072);
not NOT1 (N6334, N6331);
xor XOR2 (N6335, N6334, N1122);
not NOT1 (N6336, N6329);
buf BUF1 (N6337, N6332);
nor NOR2 (N6338, N6326, N4327);
and AND4 (N6339, N6322, N4311, N891, N3239);
and AND4 (N6340, N6336, N310, N4831, N2378);
buf BUF1 (N6341, N6330);
nor NOR4 (N6342, N6335, N1637, N5120, N5200);
and AND4 (N6343, N6340, N4336, N2580, N3648);
not NOT1 (N6344, N6338);
nand NAND2 (N6345, N6342, N2084);
not NOT1 (N6346, N6337);
nor NOR2 (N6347, N6320, N4624);
or OR4 (N6348, N6346, N609, N3848, N4744);
not NOT1 (N6349, N6348);
xor XOR2 (N6350, N6345, N6065);
buf BUF1 (N6351, N6349);
or OR2 (N6352, N6343, N5784);
not NOT1 (N6353, N6341);
and AND2 (N6354, N6333, N462);
and AND3 (N6355, N6318, N4581, N5304);
buf BUF1 (N6356, N6325);
nand NAND2 (N6357, N6351, N519);
nor NOR2 (N6358, N6357, N3067);
or OR3 (N6359, N6352, N4195, N1916);
not NOT1 (N6360, N6354);
buf BUF1 (N6361, N6350);
nor NOR2 (N6362, N6339, N3590);
nor NOR2 (N6363, N6347, N5987);
not NOT1 (N6364, N6344);
not NOT1 (N6365, N6364);
buf BUF1 (N6366, N6353);
nor NOR4 (N6367, N6366, N766, N6213, N5052);
or OR3 (N6368, N6356, N698, N364);
not NOT1 (N6369, N6361);
not NOT1 (N6370, N6363);
or OR4 (N6371, N6367, N262, N4421, N1647);
not NOT1 (N6372, N6371);
nor NOR2 (N6373, N6360, N4184);
or OR2 (N6374, N6362, N6178);
or OR2 (N6375, N6368, N5281);
not NOT1 (N6376, N6372);
nand NAND2 (N6377, N6365, N1944);
nor NOR4 (N6378, N6358, N4986, N3035, N5310);
and AND4 (N6379, N6359, N169, N3163, N5292);
and AND3 (N6380, N6376, N3326, N4153);
or OR4 (N6381, N6369, N4563, N5918, N755);
nor NOR4 (N6382, N6381, N2662, N6053, N6325);
not NOT1 (N6383, N6379);
or OR4 (N6384, N6383, N4517, N4917, N1828);
and AND2 (N6385, N6382, N4031);
buf BUF1 (N6386, N6355);
xor XOR2 (N6387, N6380, N5706);
or OR4 (N6388, N6370, N6115, N2191, N1631);
buf BUF1 (N6389, N6386);
nand NAND2 (N6390, N6378, N5379);
not NOT1 (N6391, N6375);
nand NAND2 (N6392, N6377, N6106);
or OR2 (N6393, N6390, N266);
not NOT1 (N6394, N6391);
xor XOR2 (N6395, N6385, N591);
buf BUF1 (N6396, N6374);
or OR3 (N6397, N6396, N3457, N4364);
or OR3 (N6398, N6388, N3982, N1443);
not NOT1 (N6399, N6387);
or OR3 (N6400, N6392, N6023, N4721);
nand NAND4 (N6401, N6398, N6138, N4629, N5125);
nor NOR4 (N6402, N6400, N2185, N4160, N4747);
and AND4 (N6403, N6373, N1741, N3864, N2184);
not NOT1 (N6404, N6401);
or OR4 (N6405, N6389, N2300, N3922, N5721);
and AND2 (N6406, N6404, N4504);
nor NOR3 (N6407, N6406, N3452, N5441);
xor XOR2 (N6408, N6395, N5442);
not NOT1 (N6409, N6393);
xor XOR2 (N6410, N6403, N5441);
not NOT1 (N6411, N6394);
or OR4 (N6412, N6410, N1837, N4715, N5249);
nand NAND4 (N6413, N6399, N4909, N5296, N19);
nor NOR3 (N6414, N6412, N1287, N1272);
xor XOR2 (N6415, N6405, N6298);
xor XOR2 (N6416, N6407, N5877);
buf BUF1 (N6417, N6402);
and AND2 (N6418, N6384, N5315);
nor NOR4 (N6419, N6408, N5221, N5963, N6416);
nor NOR2 (N6420, N528, N3316);
xor XOR2 (N6421, N6409, N4352);
and AND2 (N6422, N6397, N4464);
or OR3 (N6423, N6415, N2318, N2098);
not NOT1 (N6424, N6423);
nand NAND2 (N6425, N6414, N6418);
nand NAND2 (N6426, N1141, N6244);
not NOT1 (N6427, N6424);
nor NOR3 (N6428, N6422, N2222, N2658);
not NOT1 (N6429, N6413);
xor XOR2 (N6430, N6425, N1662);
and AND2 (N6431, N6417, N2616);
or OR2 (N6432, N6419, N5624);
not NOT1 (N6433, N6432);
xor XOR2 (N6434, N6428, N2645);
and AND3 (N6435, N6427, N1247, N4514);
nand NAND4 (N6436, N6434, N3256, N4629, N3534);
buf BUF1 (N6437, N6436);
buf BUF1 (N6438, N6435);
nor NOR4 (N6439, N6433, N4555, N2471, N4446);
xor XOR2 (N6440, N6411, N4166);
or OR2 (N6441, N6438, N334);
or OR3 (N6442, N6439, N1280, N1907);
nand NAND2 (N6443, N6437, N3174);
xor XOR2 (N6444, N6442, N5146);
nand NAND3 (N6445, N6429, N904, N771);
nor NOR2 (N6446, N6443, N670);
nor NOR3 (N6447, N6445, N358, N4858);
not NOT1 (N6448, N6446);
xor XOR2 (N6449, N6421, N148);
and AND2 (N6450, N6444, N3851);
nor NOR2 (N6451, N6441, N6272);
and AND4 (N6452, N6451, N888, N6187, N985);
buf BUF1 (N6453, N6450);
nand NAND4 (N6454, N6453, N2283, N4914, N5300);
nand NAND2 (N6455, N6420, N4722);
nand NAND3 (N6456, N6449, N1078, N103);
and AND4 (N6457, N6426, N4202, N3823, N1076);
nand NAND4 (N6458, N6448, N2559, N5106, N1745);
and AND4 (N6459, N6457, N3942, N5523, N5692);
and AND3 (N6460, N6459, N4445, N5974);
not NOT1 (N6461, N6456);
or OR2 (N6462, N6458, N5729);
or OR2 (N6463, N6454, N723);
nor NOR2 (N6464, N6447, N2681);
nor NOR4 (N6465, N6462, N5980, N12, N736);
not NOT1 (N6466, N6464);
nand NAND3 (N6467, N6455, N4007, N4747);
nand NAND2 (N6468, N6467, N2601);
or OR4 (N6469, N6466, N3289, N623, N6115);
and AND3 (N6470, N6431, N36, N2825);
not NOT1 (N6471, N6469);
nor NOR3 (N6472, N6452, N5485, N3800);
and AND4 (N6473, N6430, N4289, N1564, N143);
nand NAND3 (N6474, N6471, N3736, N6374);
nor NOR4 (N6475, N6463, N3160, N3497, N2690);
buf BUF1 (N6476, N6473);
or OR2 (N6477, N6472, N3176);
nand NAND2 (N6478, N6460, N4220);
nand NAND2 (N6479, N6465, N5405);
or OR4 (N6480, N6476, N3377, N1803, N4113);
not NOT1 (N6481, N6478);
xor XOR2 (N6482, N6477, N6077);
and AND3 (N6483, N6481, N1524, N1682);
nand NAND3 (N6484, N6440, N5048, N3058);
buf BUF1 (N6485, N6482);
xor XOR2 (N6486, N6480, N795);
not NOT1 (N6487, N6468);
xor XOR2 (N6488, N6486, N5994);
nor NOR4 (N6489, N6479, N1643, N2986, N1391);
xor XOR2 (N6490, N6461, N2249);
buf BUF1 (N6491, N6485);
nor NOR3 (N6492, N6470, N5747, N1600);
and AND3 (N6493, N6488, N3839, N794);
not NOT1 (N6494, N6493);
nor NOR3 (N6495, N6475, N3897, N1825);
nor NOR3 (N6496, N6474, N5807, N6395);
buf BUF1 (N6497, N6496);
nor NOR3 (N6498, N6487, N931, N1612);
and AND3 (N6499, N6495, N4154, N4585);
nor NOR2 (N6500, N6494, N6276);
nor NOR4 (N6501, N6490, N3221, N808, N409);
xor XOR2 (N6502, N6492, N1788);
nor NOR3 (N6503, N6501, N2420, N4203);
buf BUF1 (N6504, N6497);
not NOT1 (N6505, N6483);
and AND3 (N6506, N6500, N3609, N5093);
nand NAND4 (N6507, N6499, N3800, N4127, N856);
buf BUF1 (N6508, N6507);
or OR4 (N6509, N6508, N3388, N6067, N130);
and AND4 (N6510, N6489, N3000, N5428, N3029);
nand NAND2 (N6511, N6509, N4755);
or OR2 (N6512, N6484, N1841);
not NOT1 (N6513, N6491);
nand NAND2 (N6514, N6510, N3360);
or OR3 (N6515, N6512, N2137, N6159);
not NOT1 (N6516, N6511);
nand NAND4 (N6517, N6503, N5246, N1484, N4550);
buf BUF1 (N6518, N6517);
not NOT1 (N6519, N6514);
buf BUF1 (N6520, N6518);
buf BUF1 (N6521, N6506);
not NOT1 (N6522, N6515);
not NOT1 (N6523, N6502);
nor NOR4 (N6524, N6520, N5188, N365, N4205);
or OR3 (N6525, N6505, N1456, N5736);
nand NAND4 (N6526, N6525, N3825, N4165, N2431);
or OR3 (N6527, N6523, N4509, N3362);
or OR3 (N6528, N6498, N4026, N6188);
and AND3 (N6529, N6504, N4447, N4348);
nor NOR3 (N6530, N6526, N6112, N2294);
nor NOR2 (N6531, N6529, N6495);
and AND3 (N6532, N6519, N5650, N6002);
nor NOR4 (N6533, N6528, N4805, N2778, N3583);
and AND3 (N6534, N6513, N1147, N2490);
buf BUF1 (N6535, N6533);
not NOT1 (N6536, N6521);
nand NAND2 (N6537, N6527, N6300);
and AND2 (N6538, N6536, N2444);
nand NAND3 (N6539, N6530, N5593, N1780);
buf BUF1 (N6540, N6537);
not NOT1 (N6541, N6538);
or OR2 (N6542, N6516, N1261);
nor NOR2 (N6543, N6532, N3275);
and AND2 (N6544, N6535, N824);
xor XOR2 (N6545, N6543, N4957);
nor NOR2 (N6546, N6531, N3945);
or OR3 (N6547, N6534, N3003, N6083);
and AND2 (N6548, N6524, N4239);
buf BUF1 (N6549, N6544);
or OR4 (N6550, N6541, N1762, N3058, N3141);
or OR3 (N6551, N6546, N368, N1516);
buf BUF1 (N6552, N6522);
nand NAND2 (N6553, N6542, N4542);
nor NOR3 (N6554, N6548, N5630, N2499);
nand NAND3 (N6555, N6553, N1830, N4849);
and AND4 (N6556, N6551, N4575, N1616, N3366);
xor XOR2 (N6557, N6539, N328);
or OR4 (N6558, N6550, N4650, N2132, N3262);
xor XOR2 (N6559, N6558, N5003);
not NOT1 (N6560, N6556);
buf BUF1 (N6561, N6547);
nand NAND4 (N6562, N6540, N4681, N3011, N6362);
nor NOR2 (N6563, N6545, N3034);
xor XOR2 (N6564, N6560, N5315);
or OR2 (N6565, N6549, N2664);
nor NOR2 (N6566, N6565, N6207);
nand NAND2 (N6567, N6555, N5630);
not NOT1 (N6568, N6559);
not NOT1 (N6569, N6566);
xor XOR2 (N6570, N6554, N6403);
not NOT1 (N6571, N6561);
not NOT1 (N6572, N6564);
and AND4 (N6573, N6567, N1636, N1433, N2968);
or OR2 (N6574, N6562, N4046);
nor NOR3 (N6575, N6570, N1743, N4349);
buf BUF1 (N6576, N6572);
nand NAND2 (N6577, N6552, N6477);
not NOT1 (N6578, N6571);
buf BUF1 (N6579, N6576);
nor NOR2 (N6580, N6575, N6038);
and AND3 (N6581, N6573, N1093, N3792);
not NOT1 (N6582, N6577);
and AND2 (N6583, N6578, N5882);
or OR2 (N6584, N6569, N5063);
buf BUF1 (N6585, N6582);
and AND2 (N6586, N6574, N3191);
buf BUF1 (N6587, N6584);
nor NOR2 (N6588, N6586, N4836);
or OR4 (N6589, N6557, N2695, N4478, N6303);
nand NAND4 (N6590, N6589, N4521, N88, N619);
or OR3 (N6591, N6579, N3018, N6499);
nand NAND4 (N6592, N6563, N3106, N5642, N656);
or OR3 (N6593, N6583, N3370, N613);
nor NOR3 (N6594, N6590, N2507, N3888);
nor NOR3 (N6595, N6594, N2696, N1614);
not NOT1 (N6596, N6593);
xor XOR2 (N6597, N6591, N4096);
not NOT1 (N6598, N6587);
buf BUF1 (N6599, N6585);
xor XOR2 (N6600, N6597, N5091);
nand NAND2 (N6601, N6581, N6060);
nand NAND4 (N6602, N6580, N1661, N978, N4282);
and AND4 (N6603, N6588, N4393, N3349, N6080);
and AND4 (N6604, N6603, N5015, N4053, N5859);
buf BUF1 (N6605, N6604);
nand NAND2 (N6606, N6596, N2219);
or OR2 (N6607, N6599, N1931);
and AND3 (N6608, N6598, N6539, N2402);
nor NOR4 (N6609, N6605, N1681, N5425, N5582);
and AND2 (N6610, N6609, N2625);
xor XOR2 (N6611, N6608, N6218);
nor NOR4 (N6612, N6602, N2636, N3741, N419);
buf BUF1 (N6613, N6607);
and AND4 (N6614, N6613, N5635, N2575, N5403);
buf BUF1 (N6615, N6606);
not NOT1 (N6616, N6601);
nor NOR3 (N6617, N6611, N1935, N4662);
and AND2 (N6618, N6592, N4702);
nand NAND3 (N6619, N6615, N2933, N3966);
and AND2 (N6620, N6600, N3770);
and AND4 (N6621, N6618, N3481, N1962, N6151);
buf BUF1 (N6622, N6614);
xor XOR2 (N6623, N6619, N4171);
nor NOR4 (N6624, N6622, N2852, N6292, N3824);
or OR3 (N6625, N6621, N5063, N3515);
and AND2 (N6626, N6616, N1915);
or OR4 (N6627, N6612, N1075, N3958, N3948);
buf BUF1 (N6628, N6626);
and AND4 (N6629, N6628, N2032, N3005, N3442);
nor NOR2 (N6630, N6625, N1908);
xor XOR2 (N6631, N6610, N1002);
nand NAND4 (N6632, N6620, N3622, N1894, N5079);
and AND3 (N6633, N6595, N4216, N122);
nor NOR4 (N6634, N6568, N857, N4358, N5230);
xor XOR2 (N6635, N6630, N5748);
xor XOR2 (N6636, N6634, N1334);
nand NAND3 (N6637, N6627, N6048, N2933);
xor XOR2 (N6638, N6636, N391);
buf BUF1 (N6639, N6637);
nor NOR4 (N6640, N6624, N4608, N5189, N3264);
buf BUF1 (N6641, N6629);
buf BUF1 (N6642, N6632);
nor NOR4 (N6643, N6638, N3143, N5561, N3328);
and AND2 (N6644, N6617, N3946);
or OR4 (N6645, N6631, N5397, N3348, N4867);
xor XOR2 (N6646, N6644, N1353);
buf BUF1 (N6647, N6623);
and AND3 (N6648, N6635, N4656, N890);
buf BUF1 (N6649, N6643);
and AND4 (N6650, N6641, N6322, N6510, N1973);
xor XOR2 (N6651, N6650, N3140);
nor NOR4 (N6652, N6646, N2746, N4944, N3570);
nor NOR3 (N6653, N6652, N983, N5440);
and AND4 (N6654, N6645, N1181, N6062, N4435);
not NOT1 (N6655, N6648);
or OR3 (N6656, N6649, N2005, N4685);
nor NOR2 (N6657, N6642, N1817);
nand NAND2 (N6658, N6653, N360);
nand NAND2 (N6659, N6640, N5097);
not NOT1 (N6660, N6647);
or OR4 (N6661, N6656, N4062, N1185, N1732);
or OR4 (N6662, N6639, N2106, N2394, N1076);
nor NOR4 (N6663, N6651, N2219, N4434, N4455);
buf BUF1 (N6664, N6659);
xor XOR2 (N6665, N6661, N3187);
xor XOR2 (N6666, N6657, N5603);
nor NOR4 (N6667, N6665, N2958, N282, N6016);
and AND3 (N6668, N6666, N1116, N5099);
and AND3 (N6669, N6664, N61, N4020);
and AND4 (N6670, N6662, N6595, N893, N5639);
xor XOR2 (N6671, N6667, N220);
or OR4 (N6672, N6658, N1690, N3166, N1550);
nor NOR4 (N6673, N6672, N2634, N1144, N3374);
xor XOR2 (N6674, N6668, N4328);
nand NAND4 (N6675, N6655, N2046, N5792, N6620);
or OR2 (N6676, N6660, N335);
buf BUF1 (N6677, N6673);
buf BUF1 (N6678, N6633);
nor NOR3 (N6679, N6669, N2201, N2138);
xor XOR2 (N6680, N6679, N964);
nand NAND3 (N6681, N6654, N3930, N1348);
xor XOR2 (N6682, N6678, N1130);
or OR2 (N6683, N6670, N5933);
xor XOR2 (N6684, N6683, N2423);
or OR4 (N6685, N6663, N2154, N1962, N4761);
xor XOR2 (N6686, N6676, N30);
and AND2 (N6687, N6682, N4781);
and AND4 (N6688, N6675, N2983, N2666, N4957);
nand NAND2 (N6689, N6674, N421);
buf BUF1 (N6690, N6677);
and AND4 (N6691, N6680, N3292, N822, N5143);
nand NAND4 (N6692, N6691, N4470, N3958, N5717);
and AND4 (N6693, N6684, N667, N1715, N2116);
or OR4 (N6694, N6685, N773, N2518, N2431);
xor XOR2 (N6695, N6688, N5380);
or OR4 (N6696, N6671, N1441, N5271, N3812);
buf BUF1 (N6697, N6687);
not NOT1 (N6698, N6692);
buf BUF1 (N6699, N6681);
buf BUF1 (N6700, N6694);
xor XOR2 (N6701, N6699, N5244);
or OR4 (N6702, N6700, N1862, N2862, N6486);
nand NAND4 (N6703, N6695, N3176, N1119, N3427);
or OR4 (N6704, N6703, N2091, N2121, N2540);
or OR2 (N6705, N6701, N1371);
and AND3 (N6706, N6702, N6403, N5237);
buf BUF1 (N6707, N6697);
or OR4 (N6708, N6706, N6358, N5874, N3676);
or OR2 (N6709, N6708, N883);
buf BUF1 (N6710, N6709);
nor NOR3 (N6711, N6704, N4137, N5272);
xor XOR2 (N6712, N6705, N5172);
or OR3 (N6713, N6696, N2303, N5911);
or OR4 (N6714, N6707, N208, N445, N1135);
nand NAND2 (N6715, N6689, N2985);
nand NAND2 (N6716, N6712, N4047);
buf BUF1 (N6717, N6715);
buf BUF1 (N6718, N6710);
or OR4 (N6719, N6690, N1297, N5023, N5832);
or OR2 (N6720, N6686, N1125);
nand NAND2 (N6721, N6713, N1369);
xor XOR2 (N6722, N6698, N2951);
not NOT1 (N6723, N6722);
not NOT1 (N6724, N6717);
nor NOR3 (N6725, N6693, N3062, N2986);
xor XOR2 (N6726, N6720, N2738);
nor NOR2 (N6727, N6711, N2892);
nor NOR3 (N6728, N6716, N4369, N668);
or OR2 (N6729, N6719, N5168);
xor XOR2 (N6730, N6714, N2165);
and AND3 (N6731, N6729, N4702, N2194);
nor NOR3 (N6732, N6731, N3646, N5131);
nor NOR4 (N6733, N6723, N2645, N4037, N6677);
xor XOR2 (N6734, N6733, N296);
buf BUF1 (N6735, N6732);
not NOT1 (N6736, N6730);
and AND4 (N6737, N6718, N696, N5460, N3214);
nand NAND3 (N6738, N6728, N6255, N5110);
nand NAND4 (N6739, N6736, N4117, N3130, N4584);
buf BUF1 (N6740, N6738);
nor NOR2 (N6741, N6739, N5547);
xor XOR2 (N6742, N6726, N4731);
xor XOR2 (N6743, N6741, N5115);
and AND3 (N6744, N6737, N3923, N1029);
nor NOR2 (N6745, N6727, N5632);
and AND2 (N6746, N6742, N1275);
nand NAND3 (N6747, N6721, N5347, N5208);
nor NOR2 (N6748, N6724, N2557);
xor XOR2 (N6749, N6747, N2088);
nand NAND3 (N6750, N6745, N3549, N6347);
not NOT1 (N6751, N6748);
or OR3 (N6752, N6735, N5921, N453);
and AND4 (N6753, N6749, N6140, N3959, N5397);
or OR2 (N6754, N6743, N5350);
nor NOR3 (N6755, N6746, N5589, N6697);
nor NOR3 (N6756, N6734, N86, N4022);
not NOT1 (N6757, N6725);
and AND2 (N6758, N6757, N3095);
and AND3 (N6759, N6744, N2170, N5944);
nand NAND4 (N6760, N6740, N1729, N131, N4637);
nor NOR2 (N6761, N6758, N3014);
nor NOR3 (N6762, N6754, N460, N417);
nand NAND2 (N6763, N6761, N4479);
nor NOR4 (N6764, N6755, N4628, N2890, N4985);
nand NAND2 (N6765, N6759, N5891);
or OR2 (N6766, N6751, N6585);
nand NAND3 (N6767, N6752, N6280, N2486);
or OR4 (N6768, N6750, N2086, N2460, N5019);
xor XOR2 (N6769, N6767, N1877);
nand NAND4 (N6770, N6756, N1748, N4669, N1045);
nor NOR4 (N6771, N6765, N6555, N4351, N4497);
or OR4 (N6772, N6763, N5635, N1612, N3994);
xor XOR2 (N6773, N6753, N6188);
nor NOR3 (N6774, N6769, N1761, N3018);
and AND4 (N6775, N6762, N1558, N1165, N603);
nor NOR4 (N6776, N6773, N459, N1628, N6761);
or OR4 (N6777, N6760, N131, N5172, N1322);
or OR2 (N6778, N6775, N4360);
nor NOR2 (N6779, N6776, N5633);
xor XOR2 (N6780, N6770, N3597);
nand NAND3 (N6781, N6768, N1874, N2804);
and AND4 (N6782, N6766, N2367, N4191, N3784);
or OR3 (N6783, N6778, N3607, N4803);
xor XOR2 (N6784, N6781, N1175);
xor XOR2 (N6785, N6777, N1516);
not NOT1 (N6786, N6779);
buf BUF1 (N6787, N6783);
and AND3 (N6788, N6784, N1366, N3507);
and AND3 (N6789, N6774, N1719, N2691);
xor XOR2 (N6790, N6785, N5020);
buf BUF1 (N6791, N6771);
and AND4 (N6792, N6782, N1040, N3935, N324);
xor XOR2 (N6793, N6792, N3647);
or OR4 (N6794, N6789, N6344, N252, N5054);
and AND3 (N6795, N6791, N4225, N4848);
buf BUF1 (N6796, N6794);
and AND3 (N6797, N6795, N5404, N1444);
not NOT1 (N6798, N6796);
or OR4 (N6799, N6793, N3895, N6557, N5869);
or OR4 (N6800, N6764, N1825, N3778, N362);
nand NAND4 (N6801, N6800, N1868, N1633, N5154);
not NOT1 (N6802, N6790);
buf BUF1 (N6803, N6802);
nor NOR2 (N6804, N6799, N5230);
not NOT1 (N6805, N6801);
not NOT1 (N6806, N6805);
nand NAND2 (N6807, N6786, N3477);
not NOT1 (N6808, N6798);
xor XOR2 (N6809, N6804, N271);
nand NAND4 (N6810, N6787, N4143, N246, N5168);
or OR4 (N6811, N6788, N1300, N2731, N5252);
nor NOR3 (N6812, N6797, N2542, N1888);
not NOT1 (N6813, N6807);
or OR3 (N6814, N6780, N1030, N4984);
nor NOR4 (N6815, N6806, N1184, N3356, N1984);
nor NOR3 (N6816, N6811, N4700, N732);
or OR4 (N6817, N6810, N4415, N1694, N5414);
not NOT1 (N6818, N6817);
nor NOR2 (N6819, N6816, N4554);
nor NOR3 (N6820, N6772, N887, N343);
xor XOR2 (N6821, N6803, N108);
not NOT1 (N6822, N6808);
and AND4 (N6823, N6820, N5853, N5238, N3854);
not NOT1 (N6824, N6823);
or OR2 (N6825, N6812, N3021);
nor NOR4 (N6826, N6825, N4603, N2864, N1489);
and AND4 (N6827, N6815, N322, N3458, N5068);
buf BUF1 (N6828, N6821);
xor XOR2 (N6829, N6809, N1061);
not NOT1 (N6830, N6824);
nor NOR3 (N6831, N6813, N6084, N2053);
xor XOR2 (N6832, N6826, N6092);
xor XOR2 (N6833, N6829, N955);
or OR3 (N6834, N6828, N5455, N140);
nand NAND2 (N6835, N6818, N4616);
and AND2 (N6836, N6831, N804);
nand NAND3 (N6837, N6835, N4646, N6357);
xor XOR2 (N6838, N6830, N3345);
or OR4 (N6839, N6837, N6241, N2594, N75);
and AND3 (N6840, N6827, N4246, N3025);
buf BUF1 (N6841, N6822);
buf BUF1 (N6842, N6840);
buf BUF1 (N6843, N6834);
and AND3 (N6844, N6838, N6707, N5912);
buf BUF1 (N6845, N6819);
or OR4 (N6846, N6845, N5185, N621, N755);
or OR3 (N6847, N6839, N650, N5998);
or OR3 (N6848, N6844, N5023, N1010);
buf BUF1 (N6849, N6841);
or OR3 (N6850, N6814, N413, N3795);
nand NAND4 (N6851, N6833, N1353, N807, N3579);
nand NAND4 (N6852, N6850, N2979, N899, N4978);
nand NAND4 (N6853, N6847, N1471, N3601, N4583);
or OR4 (N6854, N6853, N2331, N1512, N4604);
buf BUF1 (N6855, N6852);
not NOT1 (N6856, N6832);
xor XOR2 (N6857, N6836, N1971);
or OR4 (N6858, N6854, N4380, N5773, N4530);
or OR2 (N6859, N6849, N6107);
and AND4 (N6860, N6859, N3554, N78, N6088);
xor XOR2 (N6861, N6860, N3798);
and AND2 (N6862, N6848, N1772);
and AND2 (N6863, N6842, N814);
buf BUF1 (N6864, N6858);
or OR2 (N6865, N6843, N4139);
buf BUF1 (N6866, N6857);
nor NOR2 (N6867, N6866, N1689);
and AND4 (N6868, N6861, N4799, N4307, N1574);
not NOT1 (N6869, N6862);
not NOT1 (N6870, N6868);
nor NOR4 (N6871, N6851, N5517, N3695, N5603);
xor XOR2 (N6872, N6856, N1);
nor NOR3 (N6873, N6864, N2955, N172);
nand NAND4 (N6874, N6871, N5010, N3351, N2149);
xor XOR2 (N6875, N6872, N1622);
nand NAND3 (N6876, N6867, N4184, N2488);
xor XOR2 (N6877, N6846, N5884);
nand NAND3 (N6878, N6870, N4319, N5766);
not NOT1 (N6879, N6878);
buf BUF1 (N6880, N6865);
nor NOR3 (N6881, N6869, N6558, N4293);
not NOT1 (N6882, N6863);
buf BUF1 (N6883, N6881);
nand NAND3 (N6884, N6879, N2713, N2772);
and AND2 (N6885, N6875, N3139);
not NOT1 (N6886, N6880);
or OR3 (N6887, N6874, N610, N3811);
xor XOR2 (N6888, N6885, N6819);
or OR2 (N6889, N6877, N5240);
nor NOR3 (N6890, N6876, N1298, N2522);
and AND4 (N6891, N6873, N2833, N2384, N4359);
not NOT1 (N6892, N6855);
xor XOR2 (N6893, N6890, N666);
xor XOR2 (N6894, N6884, N2913);
xor XOR2 (N6895, N6882, N3925);
xor XOR2 (N6896, N6892, N6436);
nand NAND4 (N6897, N6888, N4857, N1937, N657);
or OR2 (N6898, N6894, N4419);
not NOT1 (N6899, N6887);
or OR2 (N6900, N6895, N5865);
nor NOR2 (N6901, N6889, N4100);
and AND4 (N6902, N6883, N3846, N3484, N3128);
nor NOR2 (N6903, N6891, N1520);
and AND2 (N6904, N6897, N4290);
not NOT1 (N6905, N6886);
buf BUF1 (N6906, N6898);
nor NOR3 (N6907, N6899, N4586, N2595);
nor NOR4 (N6908, N6904, N5820, N4373, N5003);
nand NAND2 (N6909, N6903, N3253);
nand NAND4 (N6910, N6907, N3685, N793, N4471);
buf BUF1 (N6911, N6902);
and AND4 (N6912, N6908, N5738, N6413, N1700);
buf BUF1 (N6913, N6911);
and AND3 (N6914, N6896, N5843, N1640);
xor XOR2 (N6915, N6910, N3508);
not NOT1 (N6916, N6915);
xor XOR2 (N6917, N6916, N1445);
nor NOR4 (N6918, N6912, N5998, N6730, N2680);
buf BUF1 (N6919, N6901);
or OR4 (N6920, N6913, N3893, N6752, N6736);
buf BUF1 (N6921, N6900);
and AND2 (N6922, N6917, N4250);
buf BUF1 (N6923, N6919);
not NOT1 (N6924, N6923);
nor NOR2 (N6925, N6922, N4546);
and AND2 (N6926, N6918, N3953);
buf BUF1 (N6927, N6905);
or OR3 (N6928, N6924, N5444, N6044);
not NOT1 (N6929, N6893);
or OR3 (N6930, N6925, N2301, N195);
xor XOR2 (N6931, N6921, N358);
nor NOR2 (N6932, N6920, N6264);
xor XOR2 (N6933, N6928, N127);
and AND4 (N6934, N6927, N230, N6371, N574);
nor NOR4 (N6935, N6926, N539, N6178, N3112);
buf BUF1 (N6936, N6914);
or OR4 (N6937, N6932, N2897, N613, N1627);
nor NOR2 (N6938, N6909, N4145);
nor NOR4 (N6939, N6937, N4461, N1234, N170);
xor XOR2 (N6940, N6934, N2086);
xor XOR2 (N6941, N6931, N6142);
buf BUF1 (N6942, N6935);
buf BUF1 (N6943, N6906);
buf BUF1 (N6944, N6941);
not NOT1 (N6945, N6943);
or OR4 (N6946, N6929, N6753, N3762, N6738);
nand NAND4 (N6947, N6930, N134, N1303, N6097);
not NOT1 (N6948, N6944);
or OR2 (N6949, N6945, N3847);
and AND4 (N6950, N6940, N258, N2093, N6945);
nand NAND3 (N6951, N6950, N2225, N4016);
and AND2 (N6952, N6947, N236);
or OR3 (N6953, N6951, N1649, N5044);
not NOT1 (N6954, N6933);
and AND2 (N6955, N6946, N1640);
or OR2 (N6956, N6953, N4848);
xor XOR2 (N6957, N6942, N3615);
and AND3 (N6958, N6954, N1630, N6690);
xor XOR2 (N6959, N6949, N6285);
xor XOR2 (N6960, N6958, N891);
xor XOR2 (N6961, N6956, N1202);
nor NOR4 (N6962, N6939, N2876, N753, N4770);
not NOT1 (N6963, N6936);
nor NOR2 (N6964, N6955, N5621);
not NOT1 (N6965, N6963);
nor NOR4 (N6966, N6960, N5495, N3082, N4964);
buf BUF1 (N6967, N6964);
not NOT1 (N6968, N6962);
xor XOR2 (N6969, N6959, N2243);
or OR4 (N6970, N6938, N3311, N6450, N5648);
xor XOR2 (N6971, N6961, N208);
not NOT1 (N6972, N6968);
or OR3 (N6973, N6965, N1426, N5097);
nor NOR2 (N6974, N6966, N6968);
nor NOR4 (N6975, N6957, N2104, N3002, N2091);
nand NAND2 (N6976, N6975, N6038);
xor XOR2 (N6977, N6948, N2181);
and AND4 (N6978, N6970, N1211, N4479, N190);
buf BUF1 (N6979, N6974);
not NOT1 (N6980, N6973);
buf BUF1 (N6981, N6971);
or OR3 (N6982, N6969, N4976, N3982);
nor NOR4 (N6983, N6972, N480, N4375, N359);
nor NOR3 (N6984, N6978, N6056, N1769);
nor NOR2 (N6985, N6981, N2589);
xor XOR2 (N6986, N6967, N4063);
buf BUF1 (N6987, N6980);
nand NAND4 (N6988, N6986, N1196, N61, N5926);
nand NAND4 (N6989, N6982, N236, N6276, N2015);
not NOT1 (N6990, N6984);
buf BUF1 (N6991, N6989);
nor NOR3 (N6992, N6976, N5661, N4180);
xor XOR2 (N6993, N6979, N2706);
nand NAND3 (N6994, N6990, N1164, N6445);
buf BUF1 (N6995, N6994);
nand NAND3 (N6996, N6992, N120, N4807);
not NOT1 (N6997, N6993);
xor XOR2 (N6998, N6996, N4372);
buf BUF1 (N6999, N6952);
not NOT1 (N7000, N6995);
nor NOR4 (N7001, N7000, N1877, N604, N3405);
xor XOR2 (N7002, N6985, N2759);
xor XOR2 (N7003, N6988, N4879);
buf BUF1 (N7004, N6977);
nor NOR3 (N7005, N6983, N3210, N1244);
xor XOR2 (N7006, N6998, N2665);
nor NOR2 (N7007, N6997, N2570);
nor NOR4 (N7008, N6991, N3288, N5194, N5542);
nor NOR2 (N7009, N7003, N5117);
and AND2 (N7010, N7009, N3632);
or OR4 (N7011, N6987, N2173, N6323, N744);
and AND2 (N7012, N7011, N440);
xor XOR2 (N7013, N7004, N5413);
nand NAND2 (N7014, N7001, N6763);
nand NAND3 (N7015, N7013, N455, N2020);
nand NAND2 (N7016, N7015, N1594);
nor NOR2 (N7017, N6999, N5686);
nand NAND2 (N7018, N7016, N4699);
or OR2 (N7019, N7014, N4581);
not NOT1 (N7020, N7012);
buf BUF1 (N7021, N7008);
or OR2 (N7022, N7005, N567);
nand NAND4 (N7023, N7006, N806, N1885, N2817);
buf BUF1 (N7024, N7017);
not NOT1 (N7025, N7023);
not NOT1 (N7026, N7010);
xor XOR2 (N7027, N7026, N4550);
and AND3 (N7028, N7018, N4807, N875);
nor NOR4 (N7029, N7022, N1898, N765, N5536);
not NOT1 (N7030, N7019);
nand NAND2 (N7031, N7029, N2829);
nor NOR4 (N7032, N7024, N2141, N6252, N5493);
or OR2 (N7033, N7007, N2718);
not NOT1 (N7034, N7032);
xor XOR2 (N7035, N7030, N88);
and AND3 (N7036, N7002, N6225, N3220);
nor NOR2 (N7037, N7033, N2876);
xor XOR2 (N7038, N7028, N2370);
or OR4 (N7039, N7034, N4361, N1354, N3527);
xor XOR2 (N7040, N7025, N5979);
nand NAND2 (N7041, N7031, N17);
xor XOR2 (N7042, N7027, N2805);
nor NOR3 (N7043, N7037, N1943, N485);
nand NAND2 (N7044, N7040, N5761);
nor NOR4 (N7045, N7044, N5249, N6627, N6382);
nor NOR3 (N7046, N7045, N6936, N2684);
or OR4 (N7047, N7036, N5217, N6241, N6831);
nor NOR4 (N7048, N7035, N1302, N3239, N3274);
nor NOR2 (N7049, N7048, N4192);
nor NOR3 (N7050, N7020, N2249, N4217);
or OR2 (N7051, N7021, N2629);
not NOT1 (N7052, N7038);
or OR3 (N7053, N7046, N4518, N1141);
not NOT1 (N7054, N7051);
not NOT1 (N7055, N7039);
and AND3 (N7056, N7052, N6393, N92);
and AND3 (N7057, N7053, N3655, N2261);
or OR3 (N7058, N7049, N4003, N145);
nor NOR4 (N7059, N7050, N2549, N3572, N1127);
xor XOR2 (N7060, N7059, N6706);
xor XOR2 (N7061, N7043, N5194);
not NOT1 (N7062, N7057);
buf BUF1 (N7063, N7047);
or OR4 (N7064, N7063, N4891, N1130, N600);
nand NAND2 (N7065, N7042, N4354);
or OR4 (N7066, N7055, N6464, N1721, N521);
and AND4 (N7067, N7064, N171, N6093, N2822);
buf BUF1 (N7068, N7061);
and AND3 (N7069, N7065, N6810, N1767);
buf BUF1 (N7070, N7068);
nor NOR4 (N7071, N7070, N5274, N4990, N6145);
buf BUF1 (N7072, N7062);
nand NAND2 (N7073, N7066, N6019);
nor NOR3 (N7074, N7060, N4801, N5979);
not NOT1 (N7075, N7069);
or OR3 (N7076, N7075, N2070, N6329);
nor NOR4 (N7077, N7071, N2224, N4550, N84);
nand NAND2 (N7078, N7067, N1517);
buf BUF1 (N7079, N7078);
not NOT1 (N7080, N7058);
not NOT1 (N7081, N7041);
not NOT1 (N7082, N7080);
nor NOR2 (N7083, N7072, N6684);
nand NAND4 (N7084, N7079, N6494, N1158, N6449);
nor NOR4 (N7085, N7083, N677, N1784, N4089);
nor NOR3 (N7086, N7073, N2374, N3313);
buf BUF1 (N7087, N7082);
nor NOR4 (N7088, N7084, N6008, N6799, N3969);
buf BUF1 (N7089, N7056);
or OR4 (N7090, N7088, N2136, N5265, N6752);
nand NAND3 (N7091, N7054, N1714, N2068);
xor XOR2 (N7092, N7076, N6702);
xor XOR2 (N7093, N7090, N1296);
xor XOR2 (N7094, N7093, N5992);
nand NAND3 (N7095, N7074, N117, N5480);
not NOT1 (N7096, N7091);
nor NOR3 (N7097, N7094, N3318, N2596);
and AND3 (N7098, N7077, N6916, N555);
nand NAND4 (N7099, N7097, N825, N1689, N4838);
nand NAND4 (N7100, N7089, N6581, N3482, N1344);
or OR4 (N7101, N7086, N781, N2099, N2836);
buf BUF1 (N7102, N7092);
and AND4 (N7103, N7085, N3744, N3977, N5772);
nand NAND3 (N7104, N7096, N5723, N4635);
not NOT1 (N7105, N7103);
xor XOR2 (N7106, N7100, N6074);
and AND3 (N7107, N7101, N6876, N1286);
not NOT1 (N7108, N7107);
and AND4 (N7109, N7105, N6098, N5317, N1431);
and AND2 (N7110, N7104, N6864);
nor NOR3 (N7111, N7081, N2445, N1886);
xor XOR2 (N7112, N7102, N188);
and AND4 (N7113, N7098, N4612, N5988, N6771);
or OR3 (N7114, N7095, N221, N3067);
or OR3 (N7115, N7110, N6062, N530);
or OR4 (N7116, N7111, N1745, N6624, N1867);
buf BUF1 (N7117, N7108);
nand NAND4 (N7118, N7113, N237, N2346, N3173);
buf BUF1 (N7119, N7117);
buf BUF1 (N7120, N7099);
not NOT1 (N7121, N7109);
or OR2 (N7122, N7114, N1026);
buf BUF1 (N7123, N7087);
xor XOR2 (N7124, N7115, N6209);
buf BUF1 (N7125, N7106);
not NOT1 (N7126, N7121);
buf BUF1 (N7127, N7112);
xor XOR2 (N7128, N7119, N3579);
nand NAND2 (N7129, N7127, N6489);
not NOT1 (N7130, N7124);
xor XOR2 (N7131, N7128, N4060);
nand NAND4 (N7132, N7130, N377, N4069, N4600);
xor XOR2 (N7133, N7131, N2442);
or OR3 (N7134, N7126, N1817, N3701);
buf BUF1 (N7135, N7116);
and AND4 (N7136, N7132, N5503, N5389, N6756);
and AND3 (N7137, N7118, N1197, N2034);
buf BUF1 (N7138, N7137);
or OR2 (N7139, N7138, N644);
nand NAND4 (N7140, N7120, N1870, N2127, N711);
nand NAND2 (N7141, N7123, N870);
buf BUF1 (N7142, N7122);
xor XOR2 (N7143, N7139, N6769);
nand NAND3 (N7144, N7133, N2794, N5101);
buf BUF1 (N7145, N7142);
or OR2 (N7146, N7125, N2165);
and AND3 (N7147, N7135, N2540, N3171);
not NOT1 (N7148, N7145);
not NOT1 (N7149, N7148);
and AND2 (N7150, N7136, N5232);
nor NOR3 (N7151, N7141, N2107, N4571);
or OR4 (N7152, N7144, N5889, N6575, N6483);
or OR4 (N7153, N7150, N5273, N90, N5457);
or OR3 (N7154, N7134, N6758, N5510);
not NOT1 (N7155, N7147);
not NOT1 (N7156, N7151);
xor XOR2 (N7157, N7154, N1021);
xor XOR2 (N7158, N7156, N4931);
not NOT1 (N7159, N7146);
nor NOR4 (N7160, N7159, N4207, N5880, N4636);
or OR3 (N7161, N7158, N377, N5752);
not NOT1 (N7162, N7149);
not NOT1 (N7163, N7162);
xor XOR2 (N7164, N7161, N2217);
buf BUF1 (N7165, N7157);
or OR4 (N7166, N7160, N406, N5200, N3605);
not NOT1 (N7167, N7166);
buf BUF1 (N7168, N7153);
or OR2 (N7169, N7143, N4615);
not NOT1 (N7170, N7155);
xor XOR2 (N7171, N7167, N2489);
or OR4 (N7172, N7171, N1511, N2674, N5086);
nor NOR3 (N7173, N7152, N5241, N1617);
or OR3 (N7174, N7140, N499, N230);
nand NAND2 (N7175, N7168, N5731);
nor NOR3 (N7176, N7163, N1721, N776);
buf BUF1 (N7177, N7174);
xor XOR2 (N7178, N7173, N4876);
or OR4 (N7179, N7164, N1479, N7011, N4593);
not NOT1 (N7180, N7172);
nor NOR3 (N7181, N7170, N3526, N1717);
or OR2 (N7182, N7177, N204);
and AND2 (N7183, N7169, N3521);
nor NOR3 (N7184, N7178, N661, N3243);
buf BUF1 (N7185, N7175);
or OR2 (N7186, N7129, N7170);
nor NOR3 (N7187, N7179, N749, N1025);
nand NAND3 (N7188, N7185, N3188, N6592);
buf BUF1 (N7189, N7181);
xor XOR2 (N7190, N7176, N72);
or OR4 (N7191, N7184, N4469, N4483, N5945);
and AND3 (N7192, N7191, N1057, N2753);
xor XOR2 (N7193, N7182, N4115);
nor NOR4 (N7194, N7183, N4632, N4243, N2985);
nand NAND4 (N7195, N7190, N4060, N2263, N718);
and AND3 (N7196, N7186, N6970, N4745);
nor NOR4 (N7197, N7194, N2023, N5773, N128);
nor NOR3 (N7198, N7187, N928, N599);
and AND4 (N7199, N7188, N318, N7058, N6858);
nor NOR4 (N7200, N7195, N1011, N1135, N2335);
not NOT1 (N7201, N7189);
nor NOR2 (N7202, N7192, N5467);
xor XOR2 (N7203, N7201, N5400);
and AND3 (N7204, N7165, N4159, N412);
xor XOR2 (N7205, N7198, N1419);
nand NAND4 (N7206, N7204, N1764, N6054, N3693);
or OR4 (N7207, N7193, N268, N6231, N4312);
or OR4 (N7208, N7203, N169, N1425, N2100);
nand NAND4 (N7209, N7196, N3857, N2413, N6603);
nand NAND2 (N7210, N7207, N6094);
buf BUF1 (N7211, N7197);
or OR2 (N7212, N7209, N3995);
and AND2 (N7213, N7208, N2632);
nor NOR4 (N7214, N7206, N3762, N3956, N4995);
buf BUF1 (N7215, N7214);
and AND2 (N7216, N7215, N4595);
nor NOR4 (N7217, N7199, N5354, N1474, N1290);
xor XOR2 (N7218, N7211, N4830);
and AND2 (N7219, N7216, N2311);
nand NAND4 (N7220, N7202, N2983, N4993, N1401);
nor NOR2 (N7221, N7220, N5926);
xor XOR2 (N7222, N7205, N2355);
and AND3 (N7223, N7217, N3008, N7044);
and AND3 (N7224, N7200, N5792, N5991);
and AND2 (N7225, N7219, N3174);
or OR4 (N7226, N7213, N3443, N2230, N6418);
nor NOR3 (N7227, N7221, N909, N4391);
nor NOR2 (N7228, N7210, N1915);
and AND3 (N7229, N7223, N2535, N670);
and AND2 (N7230, N7228, N2719);
nand NAND3 (N7231, N7230, N4106, N2708);
nand NAND2 (N7232, N7225, N2759);
nor NOR3 (N7233, N7231, N4815, N264);
nor NOR2 (N7234, N7232, N285);
not NOT1 (N7235, N7224);
buf BUF1 (N7236, N7235);
not NOT1 (N7237, N7212);
and AND2 (N7238, N7227, N1605);
nor NOR2 (N7239, N7234, N5740);
xor XOR2 (N7240, N7218, N3536);
or OR3 (N7241, N7240, N1263, N6057);
nand NAND4 (N7242, N7226, N1725, N5115, N5882);
and AND2 (N7243, N7233, N1247);
or OR2 (N7244, N7238, N1525);
nor NOR4 (N7245, N7242, N3679, N3039, N7094);
buf BUF1 (N7246, N7236);
and AND2 (N7247, N7229, N4029);
nand NAND2 (N7248, N7239, N4338);
or OR3 (N7249, N7241, N6277, N4393);
and AND4 (N7250, N7246, N892, N2880, N5964);
and AND2 (N7251, N7249, N1746);
buf BUF1 (N7252, N7245);
or OR3 (N7253, N7248, N6353, N6720);
not NOT1 (N7254, N7251);
not NOT1 (N7255, N7254);
buf BUF1 (N7256, N7253);
xor XOR2 (N7257, N7250, N2013);
buf BUF1 (N7258, N7243);
nand NAND3 (N7259, N7244, N5271, N7173);
not NOT1 (N7260, N7259);
buf BUF1 (N7261, N7255);
nand NAND2 (N7262, N7261, N2301);
not NOT1 (N7263, N7247);
not NOT1 (N7264, N7222);
nor NOR2 (N7265, N7263, N1657);
nor NOR4 (N7266, N7257, N4114, N1780, N3952);
buf BUF1 (N7267, N7265);
not NOT1 (N7268, N7237);
not NOT1 (N7269, N7266);
xor XOR2 (N7270, N7258, N3505);
xor XOR2 (N7271, N7268, N3850);
buf BUF1 (N7272, N7271);
nor NOR3 (N7273, N7180, N1530, N6859);
not NOT1 (N7274, N7269);
xor XOR2 (N7275, N7274, N2515);
not NOT1 (N7276, N7252);
nor NOR4 (N7277, N7273, N2998, N256, N28);
nor NOR2 (N7278, N7262, N6743);
xor XOR2 (N7279, N7275, N20);
buf BUF1 (N7280, N7276);
nor NOR4 (N7281, N7279, N598, N5203, N6283);
nor NOR4 (N7282, N7272, N6472, N6010, N2543);
and AND4 (N7283, N7278, N5333, N1224, N2274);
or OR3 (N7284, N7281, N6266, N5850);
or OR2 (N7285, N7282, N5235);
nand NAND3 (N7286, N7267, N2262, N308);
or OR4 (N7287, N7285, N3927, N1076, N1499);
nor NOR3 (N7288, N7280, N272, N856);
not NOT1 (N7289, N7256);
or OR4 (N7290, N7260, N3751, N284, N3457);
nand NAND2 (N7291, N7264, N1546);
not NOT1 (N7292, N7277);
not NOT1 (N7293, N7270);
buf BUF1 (N7294, N7283);
xor XOR2 (N7295, N7288, N5258);
nor NOR4 (N7296, N7287, N4179, N2793, N3972);
nor NOR2 (N7297, N7286, N3537);
or OR4 (N7298, N7291, N5527, N3585, N6826);
xor XOR2 (N7299, N7284, N6582);
xor XOR2 (N7300, N7293, N2032);
not NOT1 (N7301, N7298);
buf BUF1 (N7302, N7301);
buf BUF1 (N7303, N7300);
or OR4 (N7304, N7294, N4232, N3319, N2468);
or OR2 (N7305, N7290, N234);
nand NAND4 (N7306, N7304, N3519, N730, N2404);
buf BUF1 (N7307, N7296);
nand NAND2 (N7308, N7297, N4702);
and AND2 (N7309, N7302, N3828);
not NOT1 (N7310, N7307);
nand NAND3 (N7311, N7299, N1008, N5645);
nor NOR3 (N7312, N7310, N4061, N6225);
and AND3 (N7313, N7312, N6121, N102);
or OR3 (N7314, N7309, N2099, N1421);
and AND2 (N7315, N7308, N2154);
and AND4 (N7316, N7303, N2978, N6824, N3743);
buf BUF1 (N7317, N7306);
and AND3 (N7318, N7315, N4363, N4806);
nor NOR3 (N7319, N7292, N5018, N7309);
nand NAND2 (N7320, N7314, N1051);
nor NOR2 (N7321, N7318, N5135);
nand NAND3 (N7322, N7321, N1832, N7234);
nand NAND4 (N7323, N7295, N4836, N1598, N3419);
or OR4 (N7324, N7317, N1893, N1361, N6621);
or OR4 (N7325, N7322, N488, N6345, N3013);
or OR2 (N7326, N7313, N6452);
or OR4 (N7327, N7311, N6910, N3810, N2441);
or OR2 (N7328, N7325, N3632);
buf BUF1 (N7329, N7320);
and AND3 (N7330, N7329, N6683, N681);
buf BUF1 (N7331, N7326);
nand NAND3 (N7332, N7316, N4100, N5926);
buf BUF1 (N7333, N7331);
or OR4 (N7334, N7323, N6453, N6953, N3219);
or OR2 (N7335, N7319, N6838);
or OR3 (N7336, N7289, N2703, N3677);
or OR2 (N7337, N7334, N1890);
xor XOR2 (N7338, N7335, N6380);
buf BUF1 (N7339, N7336);
nor NOR3 (N7340, N7327, N7153, N6829);
xor XOR2 (N7341, N7330, N802);
buf BUF1 (N7342, N7339);
not NOT1 (N7343, N7305);
or OR4 (N7344, N7340, N3354, N4664, N2549);
and AND4 (N7345, N7342, N5993, N1072, N2173);
and AND3 (N7346, N7344, N7119, N3132);
not NOT1 (N7347, N7346);
buf BUF1 (N7348, N7343);
buf BUF1 (N7349, N7333);
buf BUF1 (N7350, N7338);
nand NAND2 (N7351, N7347, N365);
not NOT1 (N7352, N7341);
nor NOR2 (N7353, N7337, N1807);
xor XOR2 (N7354, N7353, N6643);
nand NAND2 (N7355, N7352, N1710);
nor NOR3 (N7356, N7354, N4728, N6662);
xor XOR2 (N7357, N7355, N1670);
not NOT1 (N7358, N7351);
nor NOR2 (N7359, N7324, N3816);
buf BUF1 (N7360, N7348);
nand NAND4 (N7361, N7357, N2002, N3119, N755);
nand NAND2 (N7362, N7356, N5424);
nor NOR3 (N7363, N7349, N2397, N2484);
and AND4 (N7364, N7332, N6622, N2935, N599);
nand NAND4 (N7365, N7328, N4090, N5896, N5052);
buf BUF1 (N7366, N7363);
not NOT1 (N7367, N7361);
or OR2 (N7368, N7366, N5014);
nor NOR3 (N7369, N7359, N4294, N1921);
buf BUF1 (N7370, N7345);
nand NAND2 (N7371, N7365, N4606);
or OR2 (N7372, N7371, N7032);
nor NOR4 (N7373, N7367, N3453, N3048, N668);
and AND2 (N7374, N7362, N6128);
nor NOR2 (N7375, N7372, N588);
xor XOR2 (N7376, N7360, N1727);
xor XOR2 (N7377, N7350, N5668);
and AND4 (N7378, N7368, N5330, N3253, N2611);
nor NOR3 (N7379, N7378, N6249, N6260);
or OR4 (N7380, N7379, N1560, N4281, N4769);
buf BUF1 (N7381, N7377);
or OR3 (N7382, N7376, N4397, N3134);
nand NAND2 (N7383, N7370, N2160);
nor NOR2 (N7384, N7358, N3884);
xor XOR2 (N7385, N7381, N264);
or OR3 (N7386, N7364, N7384, N5411);
and AND4 (N7387, N4209, N6134, N4505, N4238);
not NOT1 (N7388, N7380);
xor XOR2 (N7389, N7388, N981);
xor XOR2 (N7390, N7389, N4727);
nor NOR4 (N7391, N7382, N2795, N7171, N1741);
xor XOR2 (N7392, N7387, N6395);
and AND4 (N7393, N7392, N1438, N4557, N863);
nand NAND4 (N7394, N7383, N590, N1824, N4366);
and AND3 (N7395, N7375, N1565, N6534);
not NOT1 (N7396, N7395);
not NOT1 (N7397, N7396);
nor NOR3 (N7398, N7369, N4803, N3808);
or OR3 (N7399, N7398, N4558, N6048);
and AND4 (N7400, N7394, N3329, N6186, N4172);
xor XOR2 (N7401, N7374, N4688);
xor XOR2 (N7402, N7373, N2611);
nand NAND4 (N7403, N7386, N6785, N5124, N2008);
xor XOR2 (N7404, N7385, N2473);
and AND3 (N7405, N7397, N2730, N7061);
nand NAND4 (N7406, N7393, N3854, N6159, N1);
and AND3 (N7407, N7406, N783, N6979);
or OR2 (N7408, N7400, N1923);
or OR4 (N7409, N7402, N442, N990, N6537);
xor XOR2 (N7410, N7409, N6891);
not NOT1 (N7411, N7399);
not NOT1 (N7412, N7405);
nor NOR2 (N7413, N7403, N5769);
not NOT1 (N7414, N7410);
xor XOR2 (N7415, N7404, N4487);
or OR4 (N7416, N7411, N6056, N6389, N1316);
not NOT1 (N7417, N7413);
buf BUF1 (N7418, N7412);
and AND3 (N7419, N7416, N4663, N416);
not NOT1 (N7420, N7401);
or OR2 (N7421, N7414, N2175);
and AND3 (N7422, N7418, N7023, N6792);
or OR2 (N7423, N7407, N4067);
not NOT1 (N7424, N7421);
and AND2 (N7425, N7417, N739);
buf BUF1 (N7426, N7408);
nor NOR4 (N7427, N7390, N2883, N5576, N6308);
nand NAND4 (N7428, N7419, N5176, N4617, N579);
xor XOR2 (N7429, N7425, N6179);
or OR3 (N7430, N7424, N7350, N2385);
nor NOR3 (N7431, N7428, N5721, N6326);
buf BUF1 (N7432, N7431);
or OR4 (N7433, N7423, N2784, N6825, N1665);
buf BUF1 (N7434, N7422);
and AND2 (N7435, N7420, N286);
xor XOR2 (N7436, N7429, N931);
buf BUF1 (N7437, N7436);
not NOT1 (N7438, N7434);
nor NOR3 (N7439, N7437, N507, N7312);
nand NAND4 (N7440, N7432, N5983, N5414, N3773);
nand NAND4 (N7441, N7433, N5226, N6435, N6088);
nor NOR3 (N7442, N7435, N2588, N2518);
and AND2 (N7443, N7415, N3471);
not NOT1 (N7444, N7441);
nand NAND3 (N7445, N7439, N5385, N4179);
and AND4 (N7446, N7444, N1558, N5693, N6501);
xor XOR2 (N7447, N7442, N1469);
not NOT1 (N7448, N7427);
buf BUF1 (N7449, N7445);
buf BUF1 (N7450, N7448);
or OR3 (N7451, N7450, N6892, N137);
nor NOR3 (N7452, N7447, N7341, N61);
xor XOR2 (N7453, N7438, N6672);
or OR3 (N7454, N7430, N5326, N5949);
and AND2 (N7455, N7452, N733);
or OR4 (N7456, N7455, N7099, N1548, N1329);
nor NOR3 (N7457, N7453, N1068, N4512);
nand NAND4 (N7458, N7440, N706, N1256, N1505);
nand NAND4 (N7459, N7426, N5326, N296, N4181);
or OR2 (N7460, N7459, N4911);
buf BUF1 (N7461, N7443);
nor NOR2 (N7462, N7454, N2748);
nand NAND2 (N7463, N7391, N4617);
xor XOR2 (N7464, N7456, N5959);
nand NAND4 (N7465, N7451, N6788, N1978, N6326);
and AND4 (N7466, N7446, N3268, N2051, N7405);
nor NOR2 (N7467, N7462, N119);
and AND3 (N7468, N7466, N2636, N5839);
nand NAND2 (N7469, N7467, N6480);
not NOT1 (N7470, N7458);
not NOT1 (N7471, N7460);
buf BUF1 (N7472, N7461);
buf BUF1 (N7473, N7470);
not NOT1 (N7474, N7457);
nand NAND2 (N7475, N7468, N7052);
xor XOR2 (N7476, N7463, N409);
xor XOR2 (N7477, N7469, N923);
not NOT1 (N7478, N7472);
or OR2 (N7479, N7464, N4756);
xor XOR2 (N7480, N7449, N4087);
and AND3 (N7481, N7475, N6843, N3479);
buf BUF1 (N7482, N7471);
nor NOR3 (N7483, N7465, N5247, N3230);
xor XOR2 (N7484, N7477, N3859);
xor XOR2 (N7485, N7482, N6164);
nand NAND3 (N7486, N7478, N4581, N2629);
nand NAND4 (N7487, N7485, N2033, N215, N4772);
not NOT1 (N7488, N7476);
nor NOR2 (N7489, N7480, N3346);
or OR4 (N7490, N7486, N5410, N2575, N916);
buf BUF1 (N7491, N7481);
xor XOR2 (N7492, N7490, N2534);
buf BUF1 (N7493, N7483);
nand NAND2 (N7494, N7479, N3598);
and AND4 (N7495, N7473, N3867, N7117, N4099);
nand NAND4 (N7496, N7487, N232, N1584, N5497);
and AND4 (N7497, N7488, N1030, N5768, N3047);
nand NAND3 (N7498, N7493, N5073, N2580);
nor NOR2 (N7499, N7494, N6516);
and AND4 (N7500, N7491, N3991, N958, N4096);
nor NOR4 (N7501, N7474, N7230, N1005, N3135);
nor NOR3 (N7502, N7498, N3879, N5431);
nand NAND2 (N7503, N7499, N3389);
and AND3 (N7504, N7503, N1464, N7338);
buf BUF1 (N7505, N7484);
or OR3 (N7506, N7501, N2954, N128);
nand NAND2 (N7507, N7495, N7414);
or OR4 (N7508, N7506, N4017, N177, N1517);
and AND3 (N7509, N7502, N2852, N2465);
or OR3 (N7510, N7505, N6958, N2190);
xor XOR2 (N7511, N7510, N326);
not NOT1 (N7512, N7504);
and AND3 (N7513, N7512, N6758, N2641);
xor XOR2 (N7514, N7489, N4195);
or OR2 (N7515, N7509, N6459);
or OR4 (N7516, N7497, N7215, N1619, N533);
buf BUF1 (N7517, N7508);
nor NOR2 (N7518, N7513, N5719);
not NOT1 (N7519, N7514);
nand NAND2 (N7520, N7516, N6157);
buf BUF1 (N7521, N7507);
and AND4 (N7522, N7517, N6685, N3346, N3617);
buf BUF1 (N7523, N7496);
xor XOR2 (N7524, N7511, N6921);
not NOT1 (N7525, N7524);
and AND3 (N7526, N7523, N6214, N4243);
or OR3 (N7527, N7519, N5584, N6624);
or OR3 (N7528, N7525, N981, N5274);
xor XOR2 (N7529, N7527, N109);
xor XOR2 (N7530, N7492, N312);
nor NOR3 (N7531, N7515, N5292, N2731);
and AND2 (N7532, N7528, N4063);
or OR2 (N7533, N7529, N3717);
and AND2 (N7534, N7520, N6028);
buf BUF1 (N7535, N7531);
not NOT1 (N7536, N7535);
nand NAND3 (N7537, N7500, N2706, N2483);
nor NOR4 (N7538, N7522, N2203, N2673, N1913);
and AND3 (N7539, N7530, N600, N6782);
nor NOR3 (N7540, N7521, N707, N4451);
and AND2 (N7541, N7518, N3813);
nand NAND2 (N7542, N7539, N1039);
buf BUF1 (N7543, N7540);
not NOT1 (N7544, N7533);
nor NOR3 (N7545, N7534, N4712, N3853);
not NOT1 (N7546, N7543);
and AND4 (N7547, N7546, N4267, N1542, N1588);
not NOT1 (N7548, N7545);
and AND4 (N7549, N7541, N2962, N3394, N4703);
and AND2 (N7550, N7548, N871);
xor XOR2 (N7551, N7532, N3696);
nor NOR2 (N7552, N7526, N1008);
buf BUF1 (N7553, N7537);
and AND2 (N7554, N7547, N1060);
not NOT1 (N7555, N7551);
buf BUF1 (N7556, N7542);
xor XOR2 (N7557, N7552, N6609);
not NOT1 (N7558, N7555);
nor NOR4 (N7559, N7556, N3036, N2475, N728);
nor NOR3 (N7560, N7549, N1156, N392);
or OR2 (N7561, N7536, N868);
not NOT1 (N7562, N7560);
nor NOR4 (N7563, N7558, N7559, N938, N2634);
or OR4 (N7564, N4861, N7444, N2938, N6462);
buf BUF1 (N7565, N7564);
nor NOR3 (N7566, N7562, N5622, N2578);
not NOT1 (N7567, N7553);
and AND2 (N7568, N7544, N3919);
not NOT1 (N7569, N7568);
nand NAND2 (N7570, N7566, N6447);
buf BUF1 (N7571, N7561);
not NOT1 (N7572, N7565);
and AND2 (N7573, N7569, N1231);
nor NOR3 (N7574, N7554, N3580, N4029);
xor XOR2 (N7575, N7572, N3394);
nand NAND3 (N7576, N7570, N6486, N3026);
nand NAND3 (N7577, N7563, N7352, N956);
nor NOR2 (N7578, N7573, N1361);
or OR3 (N7579, N7550, N6675, N6431);
nor NOR3 (N7580, N7571, N3979, N4729);
nand NAND2 (N7581, N7577, N5254);
not NOT1 (N7582, N7574);
not NOT1 (N7583, N7538);
not NOT1 (N7584, N7582);
not NOT1 (N7585, N7584);
buf BUF1 (N7586, N7567);
and AND3 (N7587, N7579, N2686, N2094);
buf BUF1 (N7588, N7585);
and AND2 (N7589, N7580, N2638);
nor NOR3 (N7590, N7575, N6953, N2170);
nor NOR3 (N7591, N7583, N1542, N6328);
not NOT1 (N7592, N7557);
buf BUF1 (N7593, N7589);
nand NAND4 (N7594, N7581, N3052, N5235, N2179);
and AND2 (N7595, N7578, N121);
and AND4 (N7596, N7594, N1168, N1154, N5860);
not NOT1 (N7597, N7590);
not NOT1 (N7598, N7587);
xor XOR2 (N7599, N7586, N6141);
nor NOR3 (N7600, N7597, N5033, N372);
nor NOR3 (N7601, N7596, N4404, N2864);
nor NOR2 (N7602, N7595, N3411);
or OR3 (N7603, N7591, N829, N5634);
not NOT1 (N7604, N7601);
nor NOR3 (N7605, N7593, N7177, N5450);
xor XOR2 (N7606, N7598, N5423);
or OR3 (N7607, N7600, N4884, N151);
not NOT1 (N7608, N7604);
nor NOR3 (N7609, N7608, N668, N7445);
nor NOR4 (N7610, N7607, N726, N7464, N1412);
nor NOR4 (N7611, N7603, N6366, N1785, N2715);
not NOT1 (N7612, N7602);
nand NAND4 (N7613, N7610, N7125, N1046, N1973);
buf BUF1 (N7614, N7611);
nand NAND2 (N7615, N7599, N2748);
buf BUF1 (N7616, N7612);
or OR3 (N7617, N7592, N4142, N3019);
and AND3 (N7618, N7616, N1963, N1078);
xor XOR2 (N7619, N7618, N571);
xor XOR2 (N7620, N7619, N5536);
or OR3 (N7621, N7620, N732, N6459);
and AND2 (N7622, N7614, N3575);
and AND3 (N7623, N7588, N1469, N425);
xor XOR2 (N7624, N7615, N5610);
or OR2 (N7625, N7622, N7454);
nor NOR4 (N7626, N7613, N4547, N1806, N1914);
buf BUF1 (N7627, N7623);
nand NAND3 (N7628, N7617, N1267, N2410);
buf BUF1 (N7629, N7625);
xor XOR2 (N7630, N7629, N1461);
not NOT1 (N7631, N7606);
and AND4 (N7632, N7626, N1094, N5130, N3456);
nor NOR3 (N7633, N7605, N1391, N5030);
and AND2 (N7634, N7576, N3576);
xor XOR2 (N7635, N7627, N70);
xor XOR2 (N7636, N7635, N248);
xor XOR2 (N7637, N7631, N4966);
not NOT1 (N7638, N7637);
and AND3 (N7639, N7630, N5280, N5559);
nand NAND2 (N7640, N7621, N5549);
or OR4 (N7641, N7628, N3567, N5032, N1353);
xor XOR2 (N7642, N7624, N2054);
nor NOR2 (N7643, N7641, N6111);
xor XOR2 (N7644, N7634, N2223);
not NOT1 (N7645, N7640);
not NOT1 (N7646, N7632);
and AND2 (N7647, N7645, N5965);
or OR2 (N7648, N7636, N6363);
xor XOR2 (N7649, N7643, N5054);
and AND2 (N7650, N7648, N2736);
nor NOR4 (N7651, N7633, N1326, N6526, N4071);
not NOT1 (N7652, N7646);
or OR4 (N7653, N7651, N5616, N2274, N7328);
or OR4 (N7654, N7638, N2048, N1847, N2264);
buf BUF1 (N7655, N7649);
xor XOR2 (N7656, N7653, N3755);
xor XOR2 (N7657, N7654, N1978);
not NOT1 (N7658, N7650);
nand NAND4 (N7659, N7644, N1285, N1802, N5998);
xor XOR2 (N7660, N7639, N6214);
nor NOR2 (N7661, N7652, N5783);
not NOT1 (N7662, N7657);
buf BUF1 (N7663, N7661);
xor XOR2 (N7664, N7662, N4944);
not NOT1 (N7665, N7658);
not NOT1 (N7666, N7647);
xor XOR2 (N7667, N7642, N796);
not NOT1 (N7668, N7656);
nand NAND2 (N7669, N7659, N6671);
and AND2 (N7670, N7655, N3764);
or OR3 (N7671, N7665, N1581, N2916);
xor XOR2 (N7672, N7660, N5063);
nand NAND4 (N7673, N7667, N4438, N5881, N6203);
nor NOR4 (N7674, N7669, N3768, N130, N1077);
xor XOR2 (N7675, N7664, N2576);
or OR3 (N7676, N7671, N6257, N253);
xor XOR2 (N7677, N7673, N7010);
buf BUF1 (N7678, N7674);
and AND4 (N7679, N7609, N5851, N529, N5350);
nor NOR3 (N7680, N7679, N1556, N6362);
nor NOR2 (N7681, N7678, N1406);
buf BUF1 (N7682, N7677);
or OR2 (N7683, N7668, N426);
and AND2 (N7684, N7666, N2761);
nor NOR2 (N7685, N7672, N2147);
nand NAND4 (N7686, N7675, N5676, N1502, N5520);
and AND2 (N7687, N7680, N7575);
nand NAND4 (N7688, N7686, N4602, N4731, N1977);
xor XOR2 (N7689, N7687, N418);
or OR3 (N7690, N7684, N5212, N1597);
and AND4 (N7691, N7681, N1041, N5757, N562);
or OR2 (N7692, N7688, N5160);
nor NOR2 (N7693, N7682, N6415);
xor XOR2 (N7694, N7685, N3254);
xor XOR2 (N7695, N7670, N1198);
and AND4 (N7696, N7683, N932, N7361, N7564);
or OR4 (N7697, N7676, N2805, N7682, N7341);
nand NAND4 (N7698, N7689, N2241, N3265, N1354);
xor XOR2 (N7699, N7695, N482);
xor XOR2 (N7700, N7692, N5478);
not NOT1 (N7701, N7694);
nand NAND2 (N7702, N7701, N2685);
nand NAND2 (N7703, N7699, N7525);
buf BUF1 (N7704, N7703);
nor NOR3 (N7705, N7702, N5213, N2593);
not NOT1 (N7706, N7663);
and AND3 (N7707, N7693, N5739, N6001);
nand NAND4 (N7708, N7690, N3423, N7580, N1384);
and AND4 (N7709, N7706, N3148, N6282, N7020);
and AND3 (N7710, N7696, N3377, N2770);
nand NAND3 (N7711, N7704, N400, N7119);
and AND3 (N7712, N7709, N7458, N2834);
nand NAND4 (N7713, N7705, N5303, N4431, N1082);
not NOT1 (N7714, N7712);
nand NAND4 (N7715, N7707, N1515, N4935, N3462);
nand NAND3 (N7716, N7708, N1207, N3632);
nand NAND3 (N7717, N7697, N1950, N928);
nor NOR3 (N7718, N7716, N260, N2964);
xor XOR2 (N7719, N7713, N3856);
nand NAND2 (N7720, N7710, N6007);
buf BUF1 (N7721, N7711);
buf BUF1 (N7722, N7718);
not NOT1 (N7723, N7717);
xor XOR2 (N7724, N7700, N4197);
buf BUF1 (N7725, N7691);
nand NAND3 (N7726, N7724, N1427, N64);
or OR4 (N7727, N7698, N1350, N5491, N1480);
buf BUF1 (N7728, N7722);
nand NAND4 (N7729, N7719, N4417, N2764, N2937);
buf BUF1 (N7730, N7726);
nor NOR2 (N7731, N7728, N3197);
not NOT1 (N7732, N7714);
xor XOR2 (N7733, N7732, N3407);
nor NOR2 (N7734, N7721, N5750);
xor XOR2 (N7735, N7725, N6170);
xor XOR2 (N7736, N7715, N4282);
and AND4 (N7737, N7730, N6525, N3109, N7563);
buf BUF1 (N7738, N7727);
nor NOR2 (N7739, N7729, N2028);
nand NAND4 (N7740, N7733, N2815, N3734, N4485);
nand NAND4 (N7741, N7737, N2931, N5732, N3265);
nor NOR4 (N7742, N7720, N5160, N6531, N5462);
or OR3 (N7743, N7734, N5213, N696);
buf BUF1 (N7744, N7738);
or OR3 (N7745, N7742, N3721, N5520);
or OR2 (N7746, N7723, N7642);
nor NOR3 (N7747, N7735, N1276, N2203);
nand NAND2 (N7748, N7741, N1568);
and AND4 (N7749, N7747, N1924, N966, N2124);
nor NOR3 (N7750, N7740, N7467, N7111);
and AND2 (N7751, N7750, N4824);
xor XOR2 (N7752, N7746, N6867);
xor XOR2 (N7753, N7752, N662);
xor XOR2 (N7754, N7739, N1345);
not NOT1 (N7755, N7731);
or OR2 (N7756, N7736, N1955);
and AND2 (N7757, N7753, N1477);
not NOT1 (N7758, N7754);
buf BUF1 (N7759, N7757);
or OR2 (N7760, N7759, N670);
not NOT1 (N7761, N7751);
buf BUF1 (N7762, N7745);
xor XOR2 (N7763, N7761, N2774);
nor NOR4 (N7764, N7749, N7235, N5011, N5441);
nor NOR3 (N7765, N7748, N1697, N2413);
xor XOR2 (N7766, N7765, N2243);
or OR4 (N7767, N7764, N2849, N3835, N7542);
not NOT1 (N7768, N7758);
and AND2 (N7769, N7756, N738);
buf BUF1 (N7770, N7763);
or OR3 (N7771, N7768, N2066, N77);
nand NAND4 (N7772, N7771, N2002, N6220, N3438);
and AND2 (N7773, N7767, N6406);
and AND2 (N7774, N7755, N3367);
nor NOR4 (N7775, N7762, N7017, N5853, N6931);
xor XOR2 (N7776, N7772, N1588);
not NOT1 (N7777, N7766);
buf BUF1 (N7778, N7770);
xor XOR2 (N7779, N7760, N6563);
xor XOR2 (N7780, N7743, N5981);
or OR4 (N7781, N7780, N4571, N6792, N6392);
nor NOR4 (N7782, N7773, N6580, N6573, N6324);
and AND2 (N7783, N7781, N3573);
nor NOR2 (N7784, N7769, N7202);
nand NAND2 (N7785, N7777, N4785);
or OR3 (N7786, N7744, N3807, N2280);
nor NOR3 (N7787, N7776, N4145, N4331);
and AND2 (N7788, N7785, N7546);
buf BUF1 (N7789, N7774);
nand NAND3 (N7790, N7789, N1430, N4790);
or OR4 (N7791, N7778, N7236, N772, N4554);
nor NOR2 (N7792, N7791, N6627);
nand NAND3 (N7793, N7792, N6372, N4407);
and AND4 (N7794, N7790, N5358, N1785, N7627);
not NOT1 (N7795, N7784);
xor XOR2 (N7796, N7783, N1978);
or OR4 (N7797, N7786, N2775, N6737, N3297);
nand NAND3 (N7798, N7793, N7748, N3788);
nand NAND3 (N7799, N7798, N341, N3005);
buf BUF1 (N7800, N7796);
xor XOR2 (N7801, N7787, N639);
nor NOR4 (N7802, N7788, N921, N5699, N1808);
buf BUF1 (N7803, N7775);
not NOT1 (N7804, N7802);
or OR2 (N7805, N7795, N2650);
buf BUF1 (N7806, N7779);
xor XOR2 (N7807, N7801, N1926);
not NOT1 (N7808, N7804);
buf BUF1 (N7809, N7805);
nor NOR4 (N7810, N7807, N6655, N182, N699);
and AND3 (N7811, N7809, N4106, N6251);
or OR3 (N7812, N7794, N7422, N6790);
and AND2 (N7813, N7812, N1683);
nor NOR3 (N7814, N7811, N2480, N6918);
xor XOR2 (N7815, N7814, N7112);
xor XOR2 (N7816, N7813, N813);
xor XOR2 (N7817, N7806, N899);
not NOT1 (N7818, N7808);
nand NAND2 (N7819, N7782, N1553);
xor XOR2 (N7820, N7797, N5178);
buf BUF1 (N7821, N7819);
nor NOR4 (N7822, N7810, N4239, N3120, N5179);
or OR4 (N7823, N7816, N5174, N3061, N467);
buf BUF1 (N7824, N7818);
buf BUF1 (N7825, N7822);
and AND2 (N7826, N7803, N6192);
and AND4 (N7827, N7815, N3246, N1091, N6853);
not NOT1 (N7828, N7823);
not NOT1 (N7829, N7820);
xor XOR2 (N7830, N7817, N2519);
and AND4 (N7831, N7799, N6093, N2025, N2929);
buf BUF1 (N7832, N7821);
not NOT1 (N7833, N7829);
nor NOR2 (N7834, N7833, N7089);
not NOT1 (N7835, N7828);
nor NOR3 (N7836, N7800, N6591, N1258);
or OR4 (N7837, N7836, N2298, N4215, N2756);
and AND4 (N7838, N7826, N2272, N1870, N2539);
nor NOR3 (N7839, N7831, N5631, N7274);
nor NOR3 (N7840, N7830, N6148, N3237);
and AND2 (N7841, N7824, N592);
and AND2 (N7842, N7839, N2357);
and AND4 (N7843, N7832, N1622, N3626, N2661);
and AND2 (N7844, N7835, N1733);
nor NOR2 (N7845, N7837, N3524);
or OR4 (N7846, N7841, N1385, N7322, N3618);
nor NOR2 (N7847, N7840, N7124);
nor NOR3 (N7848, N7845, N5835, N6455);
nor NOR4 (N7849, N7844, N6994, N7005, N6283);
and AND4 (N7850, N7848, N662, N5585, N6113);
and AND2 (N7851, N7843, N7751);
not NOT1 (N7852, N7846);
and AND4 (N7853, N7827, N7238, N5833, N7653);
and AND2 (N7854, N7852, N7405);
nor NOR4 (N7855, N7854, N6776, N7402, N596);
buf BUF1 (N7856, N7850);
nor NOR3 (N7857, N7825, N1334, N3715);
not NOT1 (N7858, N7855);
xor XOR2 (N7859, N7857, N3414);
nor NOR3 (N7860, N7851, N6938, N6941);
nor NOR3 (N7861, N7842, N6304, N4341);
and AND3 (N7862, N7853, N1838, N3361);
or OR2 (N7863, N7858, N5476);
buf BUF1 (N7864, N7861);
or OR4 (N7865, N7847, N4649, N1109, N2962);
or OR4 (N7866, N7849, N5859, N5250, N124);
not NOT1 (N7867, N7864);
xor XOR2 (N7868, N7838, N7601);
and AND4 (N7869, N7865, N2794, N3784, N2460);
not NOT1 (N7870, N7834);
buf BUF1 (N7871, N7856);
nor NOR3 (N7872, N7871, N1213, N3823);
or OR2 (N7873, N7860, N4908);
nand NAND2 (N7874, N7863, N6826);
or OR4 (N7875, N7873, N3983, N1398, N4201);
or OR2 (N7876, N7874, N5508);
buf BUF1 (N7877, N7875);
and AND4 (N7878, N7876, N5542, N4532, N5637);
or OR4 (N7879, N7867, N6620, N3679, N6238);
nand NAND4 (N7880, N7879, N2124, N6086, N6019);
nand NAND4 (N7881, N7866, N684, N7045, N1331);
not NOT1 (N7882, N7868);
nand NAND2 (N7883, N7862, N7403);
xor XOR2 (N7884, N7859, N732);
nand NAND2 (N7885, N7877, N6098);
buf BUF1 (N7886, N7869);
buf BUF1 (N7887, N7870);
nor NOR3 (N7888, N7882, N7755, N3354);
nor NOR3 (N7889, N7881, N3745, N881);
xor XOR2 (N7890, N7878, N6074);
xor XOR2 (N7891, N7883, N1902);
and AND4 (N7892, N7890, N335, N3056, N6459);
or OR4 (N7893, N7888, N3728, N7661, N2262);
nor NOR2 (N7894, N7889, N7825);
and AND4 (N7895, N7892, N3330, N4891, N1290);
nand NAND4 (N7896, N7893, N11, N3034, N7333);
buf BUF1 (N7897, N7896);
not NOT1 (N7898, N7886);
or OR2 (N7899, N7880, N2843);
nor NOR4 (N7900, N7885, N838, N1734, N4970);
or OR4 (N7901, N7872, N6962, N5730, N4618);
buf BUF1 (N7902, N7898);
buf BUF1 (N7903, N7884);
xor XOR2 (N7904, N7901, N2869);
and AND2 (N7905, N7900, N4128);
buf BUF1 (N7906, N7897);
xor XOR2 (N7907, N7906, N1953);
nand NAND3 (N7908, N7904, N3582, N917);
and AND4 (N7909, N7895, N3243, N7703, N6723);
buf BUF1 (N7910, N7905);
nand NAND2 (N7911, N7909, N4794);
not NOT1 (N7912, N7903);
and AND2 (N7913, N7887, N7007);
nor NOR2 (N7914, N7913, N4736);
buf BUF1 (N7915, N7911);
and AND3 (N7916, N7910, N6489, N6138);
buf BUF1 (N7917, N7908);
nand NAND4 (N7918, N7916, N7444, N3098, N1301);
xor XOR2 (N7919, N7917, N945);
buf BUF1 (N7920, N7902);
or OR2 (N7921, N7891, N1245);
not NOT1 (N7922, N7899);
buf BUF1 (N7923, N7894);
buf BUF1 (N7924, N7919);
buf BUF1 (N7925, N7920);
not NOT1 (N7926, N7907);
xor XOR2 (N7927, N7925, N830);
xor XOR2 (N7928, N7921, N6827);
and AND4 (N7929, N7923, N3039, N455, N1851);
nand NAND4 (N7930, N7927, N5882, N2326, N5103);
buf BUF1 (N7931, N7912);
not NOT1 (N7932, N7928);
xor XOR2 (N7933, N7914, N5318);
nand NAND3 (N7934, N7931, N870, N7316);
or OR3 (N7935, N7934, N4563, N3860);
or OR4 (N7936, N7926, N2649, N6202, N7667);
nand NAND4 (N7937, N7935, N6893, N3020, N5873);
or OR4 (N7938, N7915, N7619, N4857, N582);
and AND3 (N7939, N7930, N7137, N6813);
and AND3 (N7940, N7924, N2634, N4662);
nor NOR4 (N7941, N7918, N3714, N5742, N1252);
buf BUF1 (N7942, N7940);
and AND4 (N7943, N7942, N7552, N4772, N6686);
nor NOR3 (N7944, N7929, N2897, N2686);
xor XOR2 (N7945, N7936, N401);
nor NOR3 (N7946, N7933, N614, N845);
buf BUF1 (N7947, N7922);
and AND2 (N7948, N7932, N2476);
not NOT1 (N7949, N7947);
buf BUF1 (N7950, N7944);
nand NAND3 (N7951, N7939, N5170, N3914);
xor XOR2 (N7952, N7943, N5259);
or OR3 (N7953, N7937, N1316, N3896);
not NOT1 (N7954, N7950);
nor NOR2 (N7955, N7954, N6104);
buf BUF1 (N7956, N7949);
xor XOR2 (N7957, N7952, N6610);
nor NOR3 (N7958, N7946, N4952, N1854);
nor NOR2 (N7959, N7958, N7329);
xor XOR2 (N7960, N7955, N2238);
xor XOR2 (N7961, N7948, N2337);
nor NOR3 (N7962, N7938, N2252, N6028);
and AND2 (N7963, N7941, N1024);
nand NAND4 (N7964, N7963, N3737, N2414, N2742);
or OR4 (N7965, N7945, N34, N3409, N4042);
buf BUF1 (N7966, N7964);
and AND2 (N7967, N7957, N7276);
nor NOR3 (N7968, N7966, N1221, N1539);
xor XOR2 (N7969, N7961, N3844);
and AND4 (N7970, N7951, N1593, N7588, N6356);
nand NAND2 (N7971, N7965, N6576);
nand NAND2 (N7972, N7970, N3712);
buf BUF1 (N7973, N7962);
nand NAND2 (N7974, N7960, N4052);
buf BUF1 (N7975, N7972);
buf BUF1 (N7976, N7968);
or OR3 (N7977, N7971, N1543, N7947);
and AND3 (N7978, N7967, N2578, N4154);
nor NOR4 (N7979, N7973, N5187, N2527, N4627);
buf BUF1 (N7980, N7979);
or OR4 (N7981, N7975, N1096, N52, N2214);
nand NAND4 (N7982, N7956, N7714, N7858, N7227);
not NOT1 (N7983, N7978);
or OR4 (N7984, N7953, N6514, N4839, N1168);
and AND4 (N7985, N7959, N5304, N4033, N1506);
not NOT1 (N7986, N7977);
nand NAND3 (N7987, N7985, N4937, N2903);
xor XOR2 (N7988, N7980, N778);
buf BUF1 (N7989, N7986);
or OR4 (N7990, N7974, N1528, N3100, N5632);
nor NOR3 (N7991, N7983, N3214, N1343);
or OR4 (N7992, N7984, N1699, N661, N5021);
nand NAND4 (N7993, N7981, N292, N7059, N1743);
buf BUF1 (N7994, N7993);
xor XOR2 (N7995, N7992, N2614);
nand NAND2 (N7996, N7991, N773);
nor NOR4 (N7997, N7982, N7317, N4454, N7981);
or OR4 (N7998, N7976, N3152, N1174, N7193);
and AND2 (N7999, N7990, N6090);
xor XOR2 (N8000, N7995, N5742);
and AND4 (N8001, N7987, N6730, N71, N5167);
or OR2 (N8002, N7989, N1182);
xor XOR2 (N8003, N7969, N729);
and AND3 (N8004, N8003, N6640, N4993);
nand NAND3 (N8005, N7998, N2116, N20);
nand NAND3 (N8006, N8002, N6823, N2425);
nand NAND2 (N8007, N8006, N5432);
not NOT1 (N8008, N7997);
buf BUF1 (N8009, N8007);
or OR3 (N8010, N7996, N2541, N5535);
xor XOR2 (N8011, N8009, N777);
endmodule