// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N903,N917,N915,N911,N916,N910,N900,N918,N914,N919;

nand NAND4 (N20, N14, N6, N11, N8);
nor NOR3 (N21, N13, N10, N7);
or OR3 (N22, N5, N19, N12);
or OR2 (N23, N12, N22);
nand NAND3 (N24, N8, N20, N19);
or OR2 (N25, N20, N5);
xor XOR2 (N26, N14, N7);
not NOT1 (N27, N1);
and AND4 (N28, N21, N15, N10, N7);
not NOT1 (N29, N23);
or OR4 (N30, N28, N11, N17, N24);
or OR2 (N31, N28, N1);
and AND2 (N32, N26, N11);
not NOT1 (N33, N6);
nand NAND4 (N34, N30, N4, N10, N26);
nor NOR4 (N35, N12, N32, N13, N6);
nand NAND3 (N36, N4, N3, N20);
xor XOR2 (N37, N33, N13);
not NOT1 (N38, N19);
nand NAND3 (N39, N24, N10, N38);
buf BUF1 (N40, N2);
nor NOR4 (N41, N34, N33, N10, N15);
xor XOR2 (N42, N25, N21);
nor NOR3 (N43, N41, N41, N7);
nor NOR2 (N44, N40, N10);
buf BUF1 (N45, N43);
nand NAND4 (N46, N42, N37, N35, N12);
not NOT1 (N47, N23);
not NOT1 (N48, N21);
xor XOR2 (N49, N48, N12);
or OR2 (N50, N29, N30);
not NOT1 (N51, N36);
not NOT1 (N52, N49);
xor XOR2 (N53, N31, N15);
or OR2 (N54, N27, N14);
nand NAND3 (N55, N39, N37, N50);
xor XOR2 (N56, N32, N46);
buf BUF1 (N57, N52);
buf BUF1 (N58, N53);
and AND4 (N59, N34, N53, N40, N35);
nor NOR2 (N60, N57, N1);
nor NOR4 (N61, N58, N51, N58, N33);
buf BUF1 (N62, N13);
nor NOR3 (N63, N59, N5, N27);
nor NOR4 (N64, N56, N43, N31, N12);
and AND4 (N65, N44, N46, N64, N59);
nand NAND4 (N66, N31, N48, N16, N64);
and AND4 (N67, N61, N60, N1, N9);
or OR2 (N68, N8, N3);
and AND3 (N69, N55, N44, N16);
or OR3 (N70, N66, N57, N27);
and AND2 (N71, N69, N32);
nand NAND2 (N72, N62, N71);
nor NOR2 (N73, N43, N27);
and AND3 (N74, N65, N65, N2);
buf BUF1 (N75, N72);
and AND4 (N76, N45, N28, N70, N48);
nand NAND4 (N77, N56, N68, N42, N53);
not NOT1 (N78, N8);
not NOT1 (N79, N67);
xor XOR2 (N80, N47, N66);
nand NAND4 (N81, N77, N57, N23, N34);
and AND4 (N82, N75, N10, N64, N72);
xor XOR2 (N83, N63, N65);
not NOT1 (N84, N54);
xor XOR2 (N85, N80, N1);
nor NOR4 (N86, N74, N27, N48, N11);
or OR2 (N87, N76, N3);
nand NAND2 (N88, N78, N54);
or OR3 (N89, N73, N28, N83);
nand NAND2 (N90, N83, N38);
xor XOR2 (N91, N88, N69);
buf BUF1 (N92, N84);
not NOT1 (N93, N91);
buf BUF1 (N94, N92);
and AND4 (N95, N82, N72, N7, N11);
buf BUF1 (N96, N79);
or OR3 (N97, N89, N76, N19);
xor XOR2 (N98, N86, N82);
nor NOR3 (N99, N94, N8, N65);
nor NOR4 (N100, N93, N1, N17, N66);
xor XOR2 (N101, N100, N94);
and AND4 (N102, N87, N7, N16, N79);
nor NOR2 (N103, N97, N63);
xor XOR2 (N104, N103, N7);
or OR2 (N105, N101, N89);
nand NAND3 (N106, N99, N17, N53);
nand NAND4 (N107, N106, N50, N52, N67);
and AND2 (N108, N95, N37);
not NOT1 (N109, N104);
and AND2 (N110, N105, N106);
and AND4 (N111, N107, N100, N107, N21);
nand NAND3 (N112, N85, N38, N14);
nor NOR4 (N113, N90, N96, N33, N109);
xor XOR2 (N114, N78, N15);
and AND4 (N115, N17, N61, N45, N16);
buf BUF1 (N116, N81);
buf BUF1 (N117, N114);
nand NAND2 (N118, N111, N35);
not NOT1 (N119, N102);
buf BUF1 (N120, N119);
buf BUF1 (N121, N110);
not NOT1 (N122, N115);
not NOT1 (N123, N112);
nand NAND4 (N124, N120, N88, N110, N45);
and AND4 (N125, N123, N61, N26, N82);
nand NAND3 (N126, N108, N54, N124);
and AND3 (N127, N22, N1, N91);
nand NAND4 (N128, N113, N65, N55, N125);
and AND2 (N129, N122, N111);
or OR4 (N130, N69, N19, N17, N36);
xor XOR2 (N131, N117, N4);
buf BUF1 (N132, N127);
nand NAND3 (N133, N98, N49, N119);
or OR4 (N134, N133, N38, N56, N45);
or OR4 (N135, N118, N4, N68, N26);
nand NAND2 (N136, N128, N87);
xor XOR2 (N137, N126, N46);
nand NAND2 (N138, N121, N26);
and AND4 (N139, N132, N64, N26, N126);
nor NOR3 (N140, N139, N113, N55);
nor NOR2 (N141, N131, N50);
and AND3 (N142, N135, N22, N94);
buf BUF1 (N143, N116);
nor NOR4 (N144, N140, N15, N42, N100);
not NOT1 (N145, N136);
not NOT1 (N146, N129);
buf BUF1 (N147, N134);
or OR2 (N148, N145, N68);
xor XOR2 (N149, N143, N29);
and AND2 (N150, N147, N64);
nor NOR2 (N151, N149, N43);
nand NAND3 (N152, N151, N83, N47);
not NOT1 (N153, N130);
and AND2 (N154, N141, N118);
nand NAND3 (N155, N152, N79, N81);
nor NOR2 (N156, N148, N125);
buf BUF1 (N157, N137);
nor NOR3 (N158, N154, N128, N44);
nand NAND2 (N159, N157, N149);
or OR2 (N160, N144, N22);
not NOT1 (N161, N156);
xor XOR2 (N162, N159, N61);
not NOT1 (N163, N162);
xor XOR2 (N164, N161, N97);
xor XOR2 (N165, N150, N41);
or OR3 (N166, N165, N47, N117);
not NOT1 (N167, N155);
buf BUF1 (N168, N160);
nand NAND2 (N169, N164, N103);
not NOT1 (N170, N158);
and AND4 (N171, N146, N145, N95, N33);
nand NAND2 (N172, N142, N34);
not NOT1 (N173, N153);
not NOT1 (N174, N163);
nor NOR3 (N175, N173, N78, N108);
nor NOR2 (N176, N168, N145);
nand NAND3 (N177, N175, N159, N82);
or OR4 (N178, N177, N171, N93, N132);
xor XOR2 (N179, N124, N23);
or OR2 (N180, N166, N94);
and AND4 (N181, N138, N83, N15, N158);
not NOT1 (N182, N170);
not NOT1 (N183, N174);
nand NAND2 (N184, N178, N30);
or OR4 (N185, N180, N64, N51, N103);
nand NAND2 (N186, N183, N34);
and AND3 (N187, N172, N136, N90);
xor XOR2 (N188, N167, N111);
buf BUF1 (N189, N184);
and AND4 (N190, N186, N36, N9, N66);
not NOT1 (N191, N185);
not NOT1 (N192, N182);
not NOT1 (N193, N188);
or OR4 (N194, N191, N100, N184, N75);
xor XOR2 (N195, N169, N182);
nand NAND2 (N196, N194, N3);
buf BUF1 (N197, N192);
nor NOR4 (N198, N179, N193, N193, N47);
buf BUF1 (N199, N75);
buf BUF1 (N200, N199);
not NOT1 (N201, N196);
buf BUF1 (N202, N200);
nand NAND3 (N203, N190, N58, N20);
xor XOR2 (N204, N195, N179);
xor XOR2 (N205, N203, N101);
nor NOR3 (N206, N201, N205, N85);
xor XOR2 (N207, N91, N83);
xor XOR2 (N208, N197, N197);
not NOT1 (N209, N208);
or OR3 (N210, N204, N41, N181);
nand NAND3 (N211, N131, N69, N60);
and AND4 (N212, N187, N1, N10, N178);
not NOT1 (N213, N212);
or OR2 (N214, N189, N193);
nand NAND2 (N215, N207, N43);
and AND4 (N216, N215, N98, N109, N45);
or OR3 (N217, N209, N124, N136);
and AND3 (N218, N216, N80, N99);
not NOT1 (N219, N211);
xor XOR2 (N220, N214, N114);
or OR2 (N221, N220, N82);
nand NAND4 (N222, N213, N117, N108, N78);
nor NOR4 (N223, N176, N103, N145, N2);
nor NOR4 (N224, N198, N35, N173, N170);
xor XOR2 (N225, N219, N5);
and AND4 (N226, N222, N110, N17, N60);
nor NOR3 (N227, N206, N166, N13);
nand NAND3 (N228, N218, N98, N210);
or OR2 (N229, N209, N146);
and AND4 (N230, N224, N157, N138, N44);
nor NOR2 (N231, N223, N111);
nand NAND2 (N232, N230, N55);
and AND2 (N233, N202, N27);
xor XOR2 (N234, N233, N1);
not NOT1 (N235, N226);
or OR3 (N236, N227, N91, N232);
or OR2 (N237, N157, N155);
nand NAND2 (N238, N236, N3);
or OR2 (N239, N221, N54);
not NOT1 (N240, N237);
nor NOR3 (N241, N239, N184, N109);
not NOT1 (N242, N231);
or OR3 (N243, N225, N32, N42);
nor NOR2 (N244, N228, N116);
xor XOR2 (N245, N234, N188);
nor NOR2 (N246, N245, N105);
nor NOR4 (N247, N238, N243, N35, N42);
not NOT1 (N248, N17);
buf BUF1 (N249, N217);
and AND2 (N250, N242, N66);
or OR4 (N251, N244, N216, N132, N126);
xor XOR2 (N252, N241, N27);
buf BUF1 (N253, N252);
not NOT1 (N254, N248);
or OR4 (N255, N247, N46, N28, N40);
or OR3 (N256, N253, N130, N163);
and AND4 (N257, N229, N97, N186, N170);
nand NAND3 (N258, N235, N223, N129);
and AND3 (N259, N258, N144, N26);
or OR3 (N260, N256, N4, N127);
and AND4 (N261, N255, N137, N36, N90);
buf BUF1 (N262, N250);
buf BUF1 (N263, N260);
not NOT1 (N264, N240);
xor XOR2 (N265, N263, N35);
and AND3 (N266, N259, N254, N118);
nor NOR4 (N267, N98, N156, N135, N185);
buf BUF1 (N268, N262);
xor XOR2 (N269, N268, N206);
xor XOR2 (N270, N249, N89);
nand NAND2 (N271, N261, N35);
not NOT1 (N272, N257);
and AND4 (N273, N264, N245, N258, N171);
or OR4 (N274, N251, N236, N235, N101);
xor XOR2 (N275, N271, N141);
and AND2 (N276, N265, N160);
or OR3 (N277, N246, N199, N107);
not NOT1 (N278, N274);
xor XOR2 (N279, N276, N120);
and AND4 (N280, N279, N51, N73, N138);
not NOT1 (N281, N277);
nand NAND3 (N282, N272, N31, N93);
buf BUF1 (N283, N278);
and AND4 (N284, N273, N64, N25, N273);
not NOT1 (N285, N275);
buf BUF1 (N286, N270);
buf BUF1 (N287, N284);
buf BUF1 (N288, N267);
xor XOR2 (N289, N281, N268);
and AND4 (N290, N288, N199, N8, N151);
nand NAND4 (N291, N287, N35, N148, N133);
xor XOR2 (N292, N280, N109);
not NOT1 (N293, N291);
or OR3 (N294, N269, N180, N255);
nand NAND4 (N295, N293, N185, N27, N25);
buf BUF1 (N296, N286);
nand NAND4 (N297, N296, N274, N266, N149);
nor NOR2 (N298, N222, N134);
buf BUF1 (N299, N290);
nor NOR3 (N300, N285, N232, N298);
nand NAND4 (N301, N224, N96, N81, N71);
not NOT1 (N302, N295);
nand NAND4 (N303, N300, N249, N218, N17);
xor XOR2 (N304, N294, N286);
nand NAND4 (N305, N283, N118, N225, N290);
not NOT1 (N306, N289);
nand NAND4 (N307, N297, N103, N113, N149);
buf BUF1 (N308, N307);
buf BUF1 (N309, N303);
nor NOR3 (N310, N282, N197, N204);
and AND3 (N311, N309, N70, N133);
and AND3 (N312, N304, N277, N202);
and AND2 (N313, N299, N186);
or OR2 (N314, N311, N274);
buf BUF1 (N315, N305);
nor NOR4 (N316, N314, N176, N71, N254);
nor NOR3 (N317, N292, N189, N74);
and AND3 (N318, N301, N139, N205);
buf BUF1 (N319, N306);
nand NAND4 (N320, N313, N108, N286, N287);
and AND4 (N321, N320, N82, N150, N119);
and AND4 (N322, N321, N194, N29, N219);
not NOT1 (N323, N318);
and AND2 (N324, N323, N175);
or OR2 (N325, N310, N237);
and AND3 (N326, N325, N206, N213);
and AND3 (N327, N315, N110, N171);
not NOT1 (N328, N322);
nand NAND4 (N329, N312, N120, N112, N211);
or OR4 (N330, N327, N142, N275, N198);
nand NAND4 (N331, N319, N204, N156, N197);
not NOT1 (N332, N302);
not NOT1 (N333, N331);
nand NAND4 (N334, N333, N247, N211, N137);
nor NOR4 (N335, N329, N221, N147, N59);
nand NAND3 (N336, N308, N165, N215);
or OR4 (N337, N317, N46, N107, N220);
nor NOR3 (N338, N330, N68, N285);
buf BUF1 (N339, N326);
not NOT1 (N340, N334);
or OR3 (N341, N339, N24, N331);
xor XOR2 (N342, N335, N93);
nand NAND2 (N343, N340, N62);
not NOT1 (N344, N332);
nand NAND2 (N345, N344, N335);
buf BUF1 (N346, N345);
nand NAND2 (N347, N342, N254);
nor NOR4 (N348, N343, N322, N178, N187);
not NOT1 (N349, N316);
not NOT1 (N350, N346);
not NOT1 (N351, N341);
nor NOR3 (N352, N324, N43, N206);
buf BUF1 (N353, N351);
xor XOR2 (N354, N352, N19);
buf BUF1 (N355, N336);
xor XOR2 (N356, N354, N246);
not NOT1 (N357, N356);
nand NAND3 (N358, N350, N127, N126);
nand NAND2 (N359, N337, N231);
not NOT1 (N360, N328);
not NOT1 (N361, N358);
not NOT1 (N362, N338);
buf BUF1 (N363, N362);
not NOT1 (N364, N359);
or OR4 (N365, N357, N289, N252, N16);
nand NAND3 (N366, N365, N253, N273);
not NOT1 (N367, N355);
or OR3 (N368, N348, N87, N186);
nand NAND4 (N369, N353, N238, N148, N289);
not NOT1 (N370, N349);
not NOT1 (N371, N364);
and AND4 (N372, N360, N161, N100, N144);
buf BUF1 (N373, N372);
nor NOR2 (N374, N361, N350);
and AND2 (N375, N374, N132);
and AND4 (N376, N366, N120, N189, N347);
xor XOR2 (N377, N122, N253);
and AND3 (N378, N375, N253, N290);
xor XOR2 (N379, N369, N280);
nor NOR2 (N380, N367, N181);
or OR4 (N381, N363, N272, N351, N257);
not NOT1 (N382, N378);
xor XOR2 (N383, N382, N336);
or OR4 (N384, N379, N319, N237, N364);
nand NAND4 (N385, N384, N376, N327, N205);
not NOT1 (N386, N3);
not NOT1 (N387, N385);
nand NAND4 (N388, N381, N203, N236, N104);
not NOT1 (N389, N373);
and AND4 (N390, N371, N240, N309, N119);
nor NOR2 (N391, N380, N196);
not NOT1 (N392, N368);
xor XOR2 (N393, N388, N336);
xor XOR2 (N394, N386, N229);
not NOT1 (N395, N393);
xor XOR2 (N396, N387, N238);
xor XOR2 (N397, N394, N162);
or OR4 (N398, N389, N377, N114, N300);
nor NOR2 (N399, N256, N126);
buf BUF1 (N400, N383);
nor NOR3 (N401, N398, N289, N192);
buf BUF1 (N402, N397);
not NOT1 (N403, N390);
xor XOR2 (N404, N396, N80);
and AND4 (N405, N403, N219, N143, N56);
not NOT1 (N406, N392);
nand NAND2 (N407, N404, N353);
not NOT1 (N408, N402);
not NOT1 (N409, N407);
not NOT1 (N410, N391);
or OR4 (N411, N401, N123, N282, N363);
or OR2 (N412, N406, N403);
xor XOR2 (N413, N395, N365);
nor NOR4 (N414, N412, N72, N121, N401);
buf BUF1 (N415, N410);
and AND3 (N416, N409, N380, N346);
not NOT1 (N417, N400);
buf BUF1 (N418, N411);
nand NAND4 (N419, N417, N258, N247, N162);
nand NAND3 (N420, N370, N208, N78);
nand NAND2 (N421, N416, N310);
xor XOR2 (N422, N405, N376);
nand NAND2 (N423, N413, N70);
buf BUF1 (N424, N415);
not NOT1 (N425, N419);
nand NAND4 (N426, N420, N208, N114, N35);
nand NAND3 (N427, N424, N43, N37);
and AND3 (N428, N399, N348, N35);
and AND2 (N429, N423, N319);
not NOT1 (N430, N429);
or OR3 (N431, N414, N84, N291);
xor XOR2 (N432, N422, N38);
or OR4 (N433, N427, N347, N288, N355);
nand NAND3 (N434, N425, N163, N150);
buf BUF1 (N435, N432);
and AND3 (N436, N433, N430, N203);
nor NOR2 (N437, N63, N144);
nand NAND3 (N438, N435, N74, N34);
nor NOR4 (N439, N421, N388, N345, N259);
xor XOR2 (N440, N437, N420);
not NOT1 (N441, N418);
not NOT1 (N442, N431);
nand NAND2 (N443, N408, N21);
not NOT1 (N444, N440);
or OR3 (N445, N439, N259, N134);
xor XOR2 (N446, N443, N121);
buf BUF1 (N447, N441);
xor XOR2 (N448, N434, N409);
nand NAND4 (N449, N426, N109, N140, N123);
or OR4 (N450, N447, N176, N285, N315);
xor XOR2 (N451, N436, N87);
and AND3 (N452, N445, N71, N410);
buf BUF1 (N453, N442);
buf BUF1 (N454, N452);
buf BUF1 (N455, N454);
nand NAND2 (N456, N450, N14);
or OR4 (N457, N446, N223, N256, N160);
buf BUF1 (N458, N428);
nand NAND4 (N459, N451, N77, N367, N406);
and AND4 (N460, N455, N104, N263, N293);
nor NOR2 (N461, N453, N365);
buf BUF1 (N462, N444);
and AND2 (N463, N459, N216);
nand NAND2 (N464, N438, N268);
buf BUF1 (N465, N461);
buf BUF1 (N466, N456);
nor NOR3 (N467, N457, N94, N406);
not NOT1 (N468, N464);
buf BUF1 (N469, N467);
not NOT1 (N470, N449);
nor NOR3 (N471, N463, N435, N301);
xor XOR2 (N472, N465, N85);
not NOT1 (N473, N469);
nand NAND3 (N474, N471, N251, N211);
or OR4 (N475, N462, N274, N335, N210);
not NOT1 (N476, N472);
nor NOR4 (N477, N466, N280, N327, N108);
or OR4 (N478, N460, N245, N275, N254);
nand NAND4 (N479, N475, N174, N121, N257);
or OR2 (N480, N470, N155);
or OR3 (N481, N468, N44, N123);
xor XOR2 (N482, N448, N394);
and AND3 (N483, N481, N389, N361);
not NOT1 (N484, N476);
xor XOR2 (N485, N478, N170);
buf BUF1 (N486, N483);
xor XOR2 (N487, N480, N242);
nand NAND3 (N488, N487, N447, N59);
buf BUF1 (N489, N479);
nand NAND2 (N490, N485, N259);
buf BUF1 (N491, N474);
nor NOR4 (N492, N489, N185, N402, N339);
or OR4 (N493, N488, N430, N51, N301);
nand NAND3 (N494, N458, N404, N465);
and AND3 (N495, N492, N355, N277);
nand NAND3 (N496, N473, N371, N30);
nor NOR4 (N497, N496, N337, N69, N311);
nand NAND4 (N498, N491, N346, N27, N262);
nor NOR2 (N499, N497, N252);
buf BUF1 (N500, N486);
not NOT1 (N501, N494);
nand NAND3 (N502, N499, N420, N400);
or OR2 (N503, N498, N353);
and AND4 (N504, N482, N6, N446, N301);
or OR4 (N505, N504, N238, N485, N22);
or OR3 (N506, N490, N153, N246);
not NOT1 (N507, N495);
xor XOR2 (N508, N505, N460);
not NOT1 (N509, N500);
and AND3 (N510, N503, N302, N456);
nor NOR4 (N511, N502, N222, N455, N400);
or OR2 (N512, N506, N91);
not NOT1 (N513, N507);
nand NAND3 (N514, N510, N472, N235);
and AND3 (N515, N514, N435, N110);
not NOT1 (N516, N515);
nor NOR2 (N517, N513, N255);
or OR4 (N518, N509, N342, N423, N517);
xor XOR2 (N519, N484, N365);
and AND2 (N520, N271, N328);
xor XOR2 (N521, N516, N452);
buf BUF1 (N522, N518);
nor NOR4 (N523, N493, N477, N60, N225);
nor NOR2 (N524, N228, N303);
or OR2 (N525, N523, N360);
xor XOR2 (N526, N524, N458);
and AND3 (N527, N512, N218, N139);
not NOT1 (N528, N525);
or OR2 (N529, N521, N302);
xor XOR2 (N530, N520, N322);
not NOT1 (N531, N519);
xor XOR2 (N532, N508, N123);
xor XOR2 (N533, N532, N40);
not NOT1 (N534, N531);
not NOT1 (N535, N511);
or OR2 (N536, N530, N381);
buf BUF1 (N537, N501);
buf BUF1 (N538, N529);
nor NOR2 (N539, N528, N489);
nor NOR4 (N540, N522, N505, N304, N411);
buf BUF1 (N541, N533);
or OR4 (N542, N534, N221, N212, N196);
nand NAND3 (N543, N540, N262, N372);
xor XOR2 (N544, N542, N251);
nor NOR4 (N545, N543, N264, N493, N541);
not NOT1 (N546, N252);
nand NAND4 (N547, N535, N426, N56, N419);
or OR2 (N548, N546, N276);
xor XOR2 (N549, N527, N58);
nor NOR3 (N550, N539, N446, N146);
and AND2 (N551, N547, N83);
xor XOR2 (N552, N536, N14);
nor NOR2 (N553, N545, N144);
not NOT1 (N554, N538);
and AND2 (N555, N526, N127);
and AND4 (N556, N549, N538, N437, N297);
and AND3 (N557, N548, N98, N291);
xor XOR2 (N558, N557, N269);
or OR4 (N559, N551, N397, N474, N77);
and AND3 (N560, N556, N49, N296);
or OR4 (N561, N555, N348, N161, N486);
not NOT1 (N562, N553);
and AND4 (N563, N562, N293, N208, N279);
xor XOR2 (N564, N561, N143);
and AND3 (N565, N560, N384, N63);
or OR2 (N566, N544, N91);
nor NOR4 (N567, N537, N113, N54, N482);
xor XOR2 (N568, N565, N298);
xor XOR2 (N569, N566, N167);
and AND2 (N570, N558, N116);
xor XOR2 (N571, N559, N460);
or OR3 (N572, N564, N150, N510);
and AND4 (N573, N570, N478, N83, N323);
and AND2 (N574, N571, N89);
or OR4 (N575, N568, N387, N566, N462);
nand NAND3 (N576, N575, N161, N551);
nand NAND4 (N577, N567, N153, N412, N55);
buf BUF1 (N578, N574);
and AND3 (N579, N572, N412, N504);
nor NOR3 (N580, N579, N120, N337);
not NOT1 (N581, N577);
nor NOR3 (N582, N554, N161, N326);
xor XOR2 (N583, N569, N582);
and AND2 (N584, N550, N208);
or OR2 (N585, N154, N13);
and AND4 (N586, N581, N61, N428, N548);
buf BUF1 (N587, N552);
nand NAND4 (N588, N563, N287, N117, N538);
xor XOR2 (N589, N578, N142);
nor NOR3 (N590, N573, N503, N104);
buf BUF1 (N591, N590);
or OR4 (N592, N587, N28, N178, N438);
or OR3 (N593, N576, N213, N335);
xor XOR2 (N594, N589, N94);
and AND2 (N595, N585, N89);
and AND3 (N596, N583, N155, N355);
buf BUF1 (N597, N586);
and AND3 (N598, N584, N509, N257);
buf BUF1 (N599, N596);
or OR2 (N600, N598, N178);
xor XOR2 (N601, N592, N596);
or OR2 (N602, N599, N166);
or OR2 (N603, N597, N25);
nand NAND2 (N604, N601, N100);
or OR4 (N605, N604, N70, N427, N152);
and AND3 (N606, N594, N142, N59);
and AND4 (N607, N600, N606, N528, N275);
nor NOR4 (N608, N331, N552, N186, N400);
or OR4 (N609, N607, N573, N342, N525);
and AND4 (N610, N595, N519, N487, N557);
nor NOR2 (N611, N602, N147);
or OR2 (N612, N603, N105);
and AND2 (N613, N580, N583);
xor XOR2 (N614, N612, N520);
not NOT1 (N615, N588);
buf BUF1 (N616, N611);
nor NOR3 (N617, N605, N59, N395);
buf BUF1 (N618, N610);
buf BUF1 (N619, N614);
buf BUF1 (N620, N608);
or OR4 (N621, N617, N416, N259, N97);
buf BUF1 (N622, N618);
buf BUF1 (N623, N619);
buf BUF1 (N624, N622);
not NOT1 (N625, N593);
not NOT1 (N626, N621);
buf BUF1 (N627, N616);
xor XOR2 (N628, N627, N144);
xor XOR2 (N629, N620, N247);
nor NOR4 (N630, N628, N473, N559, N582);
buf BUF1 (N631, N623);
xor XOR2 (N632, N629, N241);
nand NAND2 (N633, N609, N2);
nand NAND4 (N634, N632, N419, N191, N515);
and AND4 (N635, N615, N257, N294, N268);
nand NAND3 (N636, N613, N574, N339);
or OR2 (N637, N631, N562);
not NOT1 (N638, N591);
or OR3 (N639, N637, N20, N441);
or OR2 (N640, N626, N419);
not NOT1 (N641, N633);
and AND2 (N642, N641, N198);
nor NOR3 (N643, N636, N513, N415);
nand NAND2 (N644, N639, N508);
nand NAND2 (N645, N624, N389);
nand NAND4 (N646, N640, N28, N172, N237);
nand NAND3 (N647, N642, N304, N312);
and AND4 (N648, N638, N379, N111, N242);
or OR2 (N649, N647, N186);
nor NOR2 (N650, N625, N189);
not NOT1 (N651, N630);
and AND4 (N652, N650, N600, N153, N184);
buf BUF1 (N653, N649);
nor NOR3 (N654, N652, N561, N619);
nor NOR2 (N655, N643, N196);
not NOT1 (N656, N646);
buf BUF1 (N657, N655);
buf BUF1 (N658, N653);
buf BUF1 (N659, N656);
nor NOR4 (N660, N644, N513, N578, N72);
buf BUF1 (N661, N659);
xor XOR2 (N662, N657, N465);
not NOT1 (N663, N635);
xor XOR2 (N664, N645, N134);
and AND3 (N665, N664, N264, N212);
or OR3 (N666, N658, N126, N504);
not NOT1 (N667, N648);
xor XOR2 (N668, N661, N498);
nor NOR4 (N669, N651, N163, N517, N262);
buf BUF1 (N670, N663);
or OR4 (N671, N662, N40, N296, N606);
nor NOR3 (N672, N660, N668, N183);
xor XOR2 (N673, N371, N354);
xor XOR2 (N674, N654, N302);
nor NOR4 (N675, N667, N468, N539, N208);
and AND3 (N676, N669, N165, N58);
xor XOR2 (N677, N665, N395);
nor NOR4 (N678, N674, N128, N265, N226);
nand NAND3 (N679, N676, N435, N312);
or OR4 (N680, N671, N185, N569, N90);
buf BUF1 (N681, N677);
buf BUF1 (N682, N672);
or OR3 (N683, N679, N453, N314);
buf BUF1 (N684, N683);
xor XOR2 (N685, N673, N578);
or OR4 (N686, N670, N158, N311, N381);
or OR3 (N687, N634, N261, N326);
or OR2 (N688, N666, N132);
nand NAND4 (N689, N687, N38, N564, N444);
not NOT1 (N690, N684);
buf BUF1 (N691, N680);
or OR2 (N692, N686, N683);
nand NAND2 (N693, N685, N103);
xor XOR2 (N694, N675, N632);
not NOT1 (N695, N688);
nand NAND2 (N696, N682, N384);
buf BUF1 (N697, N692);
not NOT1 (N698, N695);
nand NAND2 (N699, N694, N664);
buf BUF1 (N700, N678);
buf BUF1 (N701, N698);
xor XOR2 (N702, N697, N698);
nand NAND3 (N703, N700, N505, N352);
and AND3 (N704, N690, N292, N538);
buf BUF1 (N705, N691);
nor NOR3 (N706, N689, N504, N285);
or OR4 (N707, N704, N700, N105, N93);
xor XOR2 (N708, N693, N402);
buf BUF1 (N709, N707);
xor XOR2 (N710, N699, N221);
nand NAND3 (N711, N701, N194, N41);
nand NAND2 (N712, N710, N45);
or OR2 (N713, N703, N252);
and AND4 (N714, N713, N22, N218, N170);
nand NAND2 (N715, N708, N466);
and AND4 (N716, N711, N312, N707, N340);
nand NAND3 (N717, N714, N61, N704);
or OR4 (N718, N709, N654, N314, N362);
not NOT1 (N719, N696);
xor XOR2 (N720, N718, N151);
and AND4 (N721, N719, N193, N304, N72);
and AND4 (N722, N721, N518, N74, N590);
not NOT1 (N723, N720);
not NOT1 (N724, N681);
nor NOR2 (N725, N723, N699);
or OR4 (N726, N717, N476, N248, N448);
buf BUF1 (N727, N706);
nand NAND2 (N728, N727, N153);
buf BUF1 (N729, N716);
not NOT1 (N730, N725);
and AND2 (N731, N730, N510);
buf BUF1 (N732, N731);
nor NOR4 (N733, N726, N194, N246, N2);
xor XOR2 (N734, N732, N569);
buf BUF1 (N735, N705);
or OR3 (N736, N724, N243, N235);
or OR4 (N737, N733, N323, N262, N415);
nor NOR3 (N738, N728, N598, N564);
nor NOR2 (N739, N737, N451);
and AND3 (N740, N729, N570, N513);
nor NOR2 (N741, N738, N538);
not NOT1 (N742, N739);
nand NAND4 (N743, N702, N227, N181, N633);
or OR2 (N744, N736, N125);
and AND4 (N745, N742, N605, N98, N725);
and AND4 (N746, N715, N400, N160, N556);
buf BUF1 (N747, N743);
or OR3 (N748, N735, N16, N667);
buf BUF1 (N749, N748);
and AND2 (N750, N746, N112);
nand NAND3 (N751, N741, N302, N658);
buf BUF1 (N752, N740);
and AND2 (N753, N749, N84);
and AND2 (N754, N752, N667);
or OR4 (N755, N745, N432, N288, N181);
nand NAND4 (N756, N755, N61, N316, N227);
xor XOR2 (N757, N747, N7);
and AND4 (N758, N722, N34, N736, N316);
nand NAND3 (N759, N751, N597, N671);
nand NAND4 (N760, N759, N329, N270, N437);
nor NOR3 (N761, N734, N336, N133);
nor NOR2 (N762, N756, N246);
and AND4 (N763, N754, N567, N304, N197);
xor XOR2 (N764, N753, N625);
nand NAND2 (N765, N744, N585);
buf BUF1 (N766, N762);
xor XOR2 (N767, N765, N470);
not NOT1 (N768, N712);
and AND2 (N769, N757, N39);
not NOT1 (N770, N761);
and AND3 (N771, N760, N757, N271);
xor XOR2 (N772, N766, N113);
nor NOR2 (N773, N750, N756);
xor XOR2 (N774, N772, N195);
xor XOR2 (N775, N764, N345);
or OR3 (N776, N775, N230, N121);
or OR3 (N777, N769, N447, N33);
buf BUF1 (N778, N771);
and AND4 (N779, N774, N328, N289, N777);
nor NOR2 (N780, N582, N456);
nor NOR4 (N781, N770, N265, N187, N280);
buf BUF1 (N782, N767);
buf BUF1 (N783, N780);
and AND2 (N784, N782, N617);
buf BUF1 (N785, N763);
xor XOR2 (N786, N784, N136);
and AND2 (N787, N781, N597);
not NOT1 (N788, N758);
xor XOR2 (N789, N786, N693);
nand NAND3 (N790, N785, N508, N717);
nand NAND2 (N791, N788, N425);
not NOT1 (N792, N776);
or OR4 (N793, N768, N217, N225, N455);
nor NOR2 (N794, N793, N630);
nor NOR4 (N795, N783, N313, N734, N11);
xor XOR2 (N796, N773, N780);
and AND3 (N797, N778, N384, N763);
nand NAND3 (N798, N790, N603, N664);
nand NAND4 (N799, N797, N578, N793, N404);
nor NOR3 (N800, N795, N623, N710);
and AND3 (N801, N791, N424, N81);
nand NAND2 (N802, N796, N628);
nand NAND4 (N803, N787, N106, N286, N289);
nor NOR2 (N804, N801, N347);
or OR3 (N805, N779, N589, N224);
nand NAND4 (N806, N800, N273, N687, N139);
xor XOR2 (N807, N802, N334);
not NOT1 (N808, N789);
nor NOR4 (N809, N808, N353, N544, N235);
buf BUF1 (N810, N792);
or OR4 (N811, N804, N254, N646, N78);
not NOT1 (N812, N810);
xor XOR2 (N813, N799, N99);
nor NOR2 (N814, N809, N470);
nor NOR4 (N815, N812, N286, N386, N714);
xor XOR2 (N816, N794, N542);
xor XOR2 (N817, N813, N774);
or OR2 (N818, N814, N304);
xor XOR2 (N819, N805, N528);
xor XOR2 (N820, N816, N431);
and AND4 (N821, N806, N35, N486, N25);
or OR4 (N822, N807, N294, N5, N157);
and AND4 (N823, N821, N275, N176, N143);
nand NAND2 (N824, N818, N376);
xor XOR2 (N825, N798, N376);
buf BUF1 (N826, N822);
or OR2 (N827, N820, N582);
xor XOR2 (N828, N819, N706);
or OR4 (N829, N811, N796, N229, N783);
nor NOR3 (N830, N827, N104, N251);
nor NOR2 (N831, N826, N249);
xor XOR2 (N832, N815, N128);
nand NAND4 (N833, N823, N228, N106, N207);
nor NOR2 (N834, N831, N810);
xor XOR2 (N835, N824, N265);
and AND4 (N836, N817, N531, N226, N631);
and AND4 (N837, N834, N171, N148, N356);
not NOT1 (N838, N829);
nor NOR2 (N839, N833, N794);
nor NOR4 (N840, N830, N372, N520, N133);
nand NAND3 (N841, N828, N346, N39);
or OR4 (N842, N835, N466, N319, N601);
nor NOR2 (N843, N842, N695);
buf BUF1 (N844, N832);
and AND2 (N845, N837, N396);
and AND2 (N846, N844, N381);
nor NOR2 (N847, N839, N605);
buf BUF1 (N848, N825);
nand NAND2 (N849, N846, N15);
nand NAND2 (N850, N840, N709);
and AND2 (N851, N849, N564);
buf BUF1 (N852, N850);
buf BUF1 (N853, N845);
nand NAND4 (N854, N852, N715, N159, N588);
buf BUF1 (N855, N843);
xor XOR2 (N856, N853, N628);
nor NOR3 (N857, N803, N622, N106);
not NOT1 (N858, N847);
xor XOR2 (N859, N838, N372);
or OR4 (N860, N848, N224, N586, N545);
buf BUF1 (N861, N855);
xor XOR2 (N862, N841, N489);
buf BUF1 (N863, N857);
not NOT1 (N864, N854);
buf BUF1 (N865, N836);
and AND3 (N866, N862, N278, N577);
nor NOR2 (N867, N861, N100);
or OR2 (N868, N858, N590);
or OR4 (N869, N856, N699, N18, N503);
buf BUF1 (N870, N869);
and AND3 (N871, N870, N361, N468);
nor NOR4 (N872, N851, N818, N392, N616);
nor NOR2 (N873, N859, N672);
xor XOR2 (N874, N863, N247);
buf BUF1 (N875, N874);
buf BUF1 (N876, N871);
and AND4 (N877, N864, N840, N725, N481);
nand NAND3 (N878, N876, N805, N135);
or OR4 (N879, N877, N248, N243, N503);
and AND3 (N880, N878, N410, N607);
and AND3 (N881, N875, N87, N197);
buf BUF1 (N882, N860);
nand NAND3 (N883, N880, N791, N303);
and AND2 (N884, N865, N4);
or OR4 (N885, N868, N276, N489, N654);
nand NAND3 (N886, N881, N300, N452);
nor NOR4 (N887, N872, N7, N532, N231);
buf BUF1 (N888, N882);
buf BUF1 (N889, N867);
nor NOR2 (N890, N884, N627);
or OR2 (N891, N866, N176);
or OR2 (N892, N886, N530);
buf BUF1 (N893, N889);
and AND4 (N894, N888, N870, N213, N480);
or OR2 (N895, N891, N413);
buf BUF1 (N896, N885);
buf BUF1 (N897, N890);
buf BUF1 (N898, N883);
nor NOR4 (N899, N887, N80, N321, N373);
and AND2 (N900, N899, N10);
xor XOR2 (N901, N879, N248);
buf BUF1 (N902, N898);
and AND4 (N903, N873, N109, N403, N48);
buf BUF1 (N904, N902);
nand NAND3 (N905, N892, N714, N647);
or OR3 (N906, N901, N86, N480);
xor XOR2 (N907, N906, N243);
xor XOR2 (N908, N895, N551);
xor XOR2 (N909, N907, N254);
or OR2 (N910, N897, N149);
nand NAND3 (N911, N904, N536, N574);
nor NOR2 (N912, N894, N697);
nand NAND4 (N913, N893, N454, N311, N618);
nor NOR2 (N914, N905, N530);
and AND2 (N915, N913, N641);
buf BUF1 (N916, N909);
nor NOR2 (N917, N912, N799);
nand NAND3 (N918, N908, N222, N327);
not NOT1 (N919, N896);
endmodule