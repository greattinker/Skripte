// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N401,N359,N409,N405,N408,N402,N400,N396,N397,N411;

nor NOR3 (N12, N8, N4, N6);
nor NOR3 (N13, N7, N10, N7);
nor NOR3 (N14, N5, N11, N5);
buf BUF1 (N15, N2);
and AND3 (N16, N10, N11, N7);
and AND2 (N17, N15, N7);
xor XOR2 (N18, N12, N12);
not NOT1 (N19, N1);
and AND3 (N20, N8, N8, N8);
buf BUF1 (N21, N14);
nand NAND4 (N22, N10, N12, N8, N17);
nand NAND4 (N23, N20, N15, N9, N19);
nand NAND3 (N24, N10, N15, N12);
nand NAND2 (N25, N24, N14);
or OR4 (N26, N11, N11, N21, N1);
and AND3 (N27, N16, N18, N18);
or OR4 (N28, N25, N19, N3, N26);
not NOT1 (N29, N22);
not NOT1 (N30, N13);
nand NAND2 (N31, N12, N13);
xor XOR2 (N32, N16, N16);
nand NAND4 (N33, N17, N25, N29, N4);
buf BUF1 (N34, N19);
or OR4 (N35, N7, N20, N33, N30);
xor XOR2 (N36, N35, N32);
and AND2 (N37, N4, N36);
nor NOR4 (N38, N11, N24, N16, N21);
xor XOR2 (N39, N37, N15);
xor XOR2 (N40, N1, N14);
and AND4 (N41, N25, N15, N6, N36);
nor NOR4 (N42, N35, N19, N28, N26);
buf BUF1 (N43, N35);
buf BUF1 (N44, N39);
or OR3 (N45, N44, N13, N30);
and AND4 (N46, N31, N12, N4, N42);
nor NOR3 (N47, N21, N41, N40);
and AND4 (N48, N1, N46, N10, N27);
not NOT1 (N49, N42);
not NOT1 (N50, N40);
xor XOR2 (N51, N8, N50);
nor NOR4 (N52, N4, N9, N40, N41);
and AND4 (N53, N23, N34, N26, N19);
xor XOR2 (N54, N31, N26);
xor XOR2 (N55, N38, N24);
xor XOR2 (N56, N48, N52);
or OR3 (N57, N55, N52, N37);
not NOT1 (N58, N18);
nor NOR3 (N59, N47, N29, N3);
xor XOR2 (N60, N49, N7);
xor XOR2 (N61, N45, N50);
and AND2 (N62, N43, N34);
nand NAND3 (N63, N60, N8, N25);
nor NOR2 (N64, N56, N17);
xor XOR2 (N65, N63, N30);
and AND4 (N66, N64, N25, N52, N33);
or OR2 (N67, N65, N66);
buf BUF1 (N68, N41);
or OR3 (N69, N51, N37, N55);
buf BUF1 (N70, N68);
not NOT1 (N71, N58);
buf BUF1 (N72, N69);
buf BUF1 (N73, N57);
or OR3 (N74, N54, N5, N42);
not NOT1 (N75, N53);
buf BUF1 (N76, N62);
or OR4 (N77, N72, N51, N20, N70);
buf BUF1 (N78, N57);
not NOT1 (N79, N73);
or OR4 (N80, N74, N63, N54, N17);
not NOT1 (N81, N59);
nor NOR3 (N82, N78, N68, N40);
or OR4 (N83, N75, N28, N55, N17);
and AND3 (N84, N79, N26, N41);
nor NOR2 (N85, N71, N70);
buf BUF1 (N86, N84);
not NOT1 (N87, N83);
and AND2 (N88, N86, N35);
or OR3 (N89, N61, N20, N42);
nor NOR4 (N90, N77, N27, N27, N64);
buf BUF1 (N91, N89);
nor NOR3 (N92, N87, N88, N87);
nand NAND2 (N93, N84, N22);
buf BUF1 (N94, N81);
or OR3 (N95, N92, N64, N33);
nor NOR2 (N96, N80, N26);
buf BUF1 (N97, N76);
xor XOR2 (N98, N85, N24);
and AND2 (N99, N91, N13);
nor NOR4 (N100, N98, N6, N55, N91);
nor NOR3 (N101, N95, N2, N41);
or OR3 (N102, N96, N32, N79);
buf BUF1 (N103, N99);
not NOT1 (N104, N67);
xor XOR2 (N105, N102, N56);
and AND2 (N106, N90, N70);
and AND4 (N107, N82, N5, N32, N29);
xor XOR2 (N108, N107, N5);
buf BUF1 (N109, N97);
nor NOR4 (N110, N100, N22, N3, N69);
and AND4 (N111, N101, N37, N106, N101);
not NOT1 (N112, N92);
not NOT1 (N113, N103);
and AND4 (N114, N105, N28, N101, N103);
not NOT1 (N115, N114);
nand NAND4 (N116, N93, N104, N89, N72);
buf BUF1 (N117, N100);
xor XOR2 (N118, N117, N15);
and AND4 (N119, N113, N86, N113, N18);
nor NOR2 (N120, N94, N77);
or OR4 (N121, N120, N85, N12, N46);
or OR4 (N122, N121, N5, N117, N53);
nor NOR4 (N123, N118, N37, N12, N80);
not NOT1 (N124, N122);
nand NAND4 (N125, N110, N7, N7, N82);
and AND3 (N126, N125, N115, N73);
nand NAND3 (N127, N64, N113, N105);
nand NAND4 (N128, N124, N61, N46, N9);
nand NAND4 (N129, N109, N75, N68, N48);
or OR4 (N130, N123, N20, N122, N89);
buf BUF1 (N131, N111);
xor XOR2 (N132, N112, N55);
nor NOR2 (N133, N129, N1);
and AND2 (N134, N127, N95);
nand NAND3 (N135, N116, N31, N131);
nor NOR4 (N136, N112, N42, N40, N56);
nor NOR3 (N137, N128, N63, N28);
not NOT1 (N138, N130);
or OR2 (N139, N134, N114);
or OR4 (N140, N132, N28, N19, N120);
xor XOR2 (N141, N139, N73);
nor NOR2 (N142, N133, N82);
not NOT1 (N143, N142);
buf BUF1 (N144, N126);
buf BUF1 (N145, N141);
nor NOR2 (N146, N143, N114);
nor NOR4 (N147, N145, N125, N61, N121);
and AND4 (N148, N146, N100, N124, N134);
buf BUF1 (N149, N138);
nor NOR3 (N150, N147, N49, N52);
nor NOR4 (N151, N108, N92, N7, N67);
nor NOR4 (N152, N148, N41, N47, N109);
buf BUF1 (N153, N152);
buf BUF1 (N154, N151);
not NOT1 (N155, N137);
buf BUF1 (N156, N149);
and AND2 (N157, N135, N100);
buf BUF1 (N158, N157);
xor XOR2 (N159, N156, N35);
not NOT1 (N160, N153);
nand NAND2 (N161, N154, N77);
and AND4 (N162, N119, N146, N160, N134);
nand NAND2 (N163, N158, N64);
and AND2 (N164, N71, N67);
not NOT1 (N165, N155);
nand NAND2 (N166, N165, N132);
nor NOR3 (N167, N144, N142, N65);
and AND2 (N168, N162, N69);
nand NAND4 (N169, N167, N59, N43, N54);
not NOT1 (N170, N159);
not NOT1 (N171, N168);
nor NOR3 (N172, N169, N54, N77);
nand NAND3 (N173, N150, N134, N106);
or OR3 (N174, N140, N138, N126);
buf BUF1 (N175, N174);
nor NOR3 (N176, N166, N111, N76);
buf BUF1 (N177, N171);
or OR3 (N178, N164, N55, N144);
buf BUF1 (N179, N136);
buf BUF1 (N180, N177);
buf BUF1 (N181, N180);
or OR2 (N182, N173, N179);
not NOT1 (N183, N100);
and AND4 (N184, N183, N104, N136, N157);
nand NAND4 (N185, N178, N164, N72, N149);
nor NOR2 (N186, N161, N9);
or OR2 (N187, N186, N72);
nor NOR3 (N188, N175, N99, N139);
nor NOR4 (N189, N163, N40, N50, N61);
xor XOR2 (N190, N181, N66);
and AND3 (N191, N184, N151, N169);
and AND3 (N192, N189, N179, N117);
or OR4 (N193, N188, N68, N165, N191);
not NOT1 (N194, N193);
nand NAND3 (N195, N98, N162, N176);
nand NAND4 (N196, N161, N183, N172, N15);
buf BUF1 (N197, N172);
xor XOR2 (N198, N182, N132);
xor XOR2 (N199, N190, N29);
buf BUF1 (N200, N195);
xor XOR2 (N201, N196, N78);
or OR3 (N202, N200, N23, N129);
or OR2 (N203, N202, N64);
buf BUF1 (N204, N199);
nand NAND3 (N205, N170, N116, N74);
xor XOR2 (N206, N205, N182);
or OR4 (N207, N203, N117, N172, N103);
or OR4 (N208, N187, N192, N51, N81);
not NOT1 (N209, N13);
or OR4 (N210, N194, N153, N29, N124);
nand NAND2 (N211, N198, N40);
nand NAND2 (N212, N210, N77);
and AND2 (N213, N201, N105);
nor NOR3 (N214, N207, N15, N76);
buf BUF1 (N215, N206);
and AND4 (N216, N185, N111, N198, N158);
or OR3 (N217, N209, N52, N174);
not NOT1 (N218, N197);
or OR2 (N219, N214, N80);
xor XOR2 (N220, N219, N73);
not NOT1 (N221, N216);
buf BUF1 (N222, N218);
nor NOR4 (N223, N212, N187, N96, N157);
xor XOR2 (N224, N221, N37);
xor XOR2 (N225, N222, N66);
xor XOR2 (N226, N204, N187);
not NOT1 (N227, N225);
nor NOR2 (N228, N208, N41);
buf BUF1 (N229, N215);
not NOT1 (N230, N226);
not NOT1 (N231, N220);
nor NOR4 (N232, N228, N113, N128, N3);
and AND3 (N233, N223, N28, N103);
nand NAND4 (N234, N213, N83, N182, N89);
buf BUF1 (N235, N217);
not NOT1 (N236, N230);
and AND2 (N237, N231, N198);
or OR2 (N238, N224, N221);
not NOT1 (N239, N235);
or OR3 (N240, N229, N234, N228);
buf BUF1 (N241, N205);
and AND4 (N242, N241, N212, N69, N133);
not NOT1 (N243, N233);
or OR3 (N244, N242, N50, N43);
and AND3 (N245, N237, N37, N23);
and AND2 (N246, N211, N124);
and AND4 (N247, N244, N204, N49, N88);
nor NOR3 (N248, N227, N38, N124);
buf BUF1 (N249, N246);
xor XOR2 (N250, N247, N54);
nand NAND3 (N251, N236, N243, N122);
or OR2 (N252, N46, N225);
nor NOR3 (N253, N250, N221, N100);
not NOT1 (N254, N232);
not NOT1 (N255, N252);
nor NOR3 (N256, N238, N73, N103);
xor XOR2 (N257, N240, N155);
or OR3 (N258, N249, N148, N74);
not NOT1 (N259, N253);
xor XOR2 (N260, N248, N25);
and AND3 (N261, N255, N236, N225);
nor NOR4 (N262, N245, N10, N217, N51);
or OR4 (N263, N257, N146, N68, N131);
or OR3 (N264, N263, N190, N22);
or OR4 (N265, N258, N109, N237, N121);
xor XOR2 (N266, N256, N79);
or OR3 (N267, N260, N124, N136);
or OR2 (N268, N259, N258);
xor XOR2 (N269, N239, N139);
and AND2 (N270, N262, N77);
nor NOR3 (N271, N264, N3, N89);
nor NOR3 (N272, N268, N172, N178);
buf BUF1 (N273, N251);
not NOT1 (N274, N265);
xor XOR2 (N275, N273, N150);
not NOT1 (N276, N254);
or OR3 (N277, N269, N174, N237);
and AND4 (N278, N276, N150, N26, N34);
or OR4 (N279, N272, N92, N91, N171);
or OR4 (N280, N261, N100, N233, N26);
and AND4 (N281, N279, N31, N17, N66);
or OR3 (N282, N277, N181, N111);
or OR3 (N283, N266, N47, N275);
or OR3 (N284, N148, N126, N124);
or OR4 (N285, N283, N119, N254, N72);
buf BUF1 (N286, N271);
not NOT1 (N287, N270);
buf BUF1 (N288, N282);
or OR4 (N289, N281, N210, N276, N120);
nor NOR4 (N290, N274, N281, N251, N142);
buf BUF1 (N291, N286);
not NOT1 (N292, N287);
or OR4 (N293, N288, N88, N257, N152);
buf BUF1 (N294, N267);
xor XOR2 (N295, N291, N162);
not NOT1 (N296, N284);
not NOT1 (N297, N290);
xor XOR2 (N298, N293, N198);
buf BUF1 (N299, N297);
nand NAND3 (N300, N289, N215, N258);
nor NOR4 (N301, N299, N222, N42, N33);
or OR2 (N302, N301, N150);
buf BUF1 (N303, N298);
xor XOR2 (N304, N296, N27);
nand NAND3 (N305, N303, N85, N280);
nand NAND4 (N306, N245, N118, N108, N165);
and AND3 (N307, N300, N25, N38);
and AND4 (N308, N285, N127, N132, N66);
and AND4 (N309, N292, N254, N299, N15);
or OR4 (N310, N302, N240, N298, N112);
nor NOR2 (N311, N278, N210);
not NOT1 (N312, N311);
xor XOR2 (N313, N304, N80);
nand NAND3 (N314, N295, N136, N215);
not NOT1 (N315, N305);
nor NOR2 (N316, N312, N51);
buf BUF1 (N317, N313);
nand NAND4 (N318, N316, N129, N313, N13);
nand NAND3 (N319, N314, N277, N287);
and AND2 (N320, N319, N10);
xor XOR2 (N321, N294, N195);
nor NOR3 (N322, N321, N195, N108);
xor XOR2 (N323, N308, N282);
and AND4 (N324, N310, N318, N298, N227);
buf BUF1 (N325, N301);
and AND2 (N326, N307, N257);
xor XOR2 (N327, N325, N30);
not NOT1 (N328, N317);
not NOT1 (N329, N324);
nand NAND3 (N330, N323, N75, N154);
buf BUF1 (N331, N326);
buf BUF1 (N332, N329);
not NOT1 (N333, N330);
not NOT1 (N334, N327);
not NOT1 (N335, N331);
or OR3 (N336, N333, N102, N250);
and AND3 (N337, N322, N79, N22);
or OR2 (N338, N332, N102);
nor NOR4 (N339, N334, N185, N309, N240);
not NOT1 (N340, N33);
not NOT1 (N341, N337);
or OR4 (N342, N320, N38, N237, N296);
or OR3 (N343, N341, N113, N99);
nand NAND3 (N344, N315, N341, N88);
or OR4 (N345, N340, N31, N294, N61);
not NOT1 (N346, N328);
nor NOR2 (N347, N342, N262);
and AND2 (N348, N336, N168);
or OR2 (N349, N348, N184);
nor NOR2 (N350, N349, N100);
nor NOR2 (N351, N339, N303);
nor NOR3 (N352, N351, N182, N273);
xor XOR2 (N353, N352, N234);
not NOT1 (N354, N347);
or OR4 (N355, N344, N59, N23, N224);
buf BUF1 (N356, N353);
not NOT1 (N357, N356);
and AND3 (N358, N343, N294, N109);
nand NAND4 (N359, N338, N161, N323, N260);
not NOT1 (N360, N358);
and AND3 (N361, N360, N122, N270);
or OR3 (N362, N346, N329, N146);
not NOT1 (N363, N306);
nand NAND4 (N364, N350, N150, N208, N128);
not NOT1 (N365, N345);
not NOT1 (N366, N354);
nor NOR4 (N367, N335, N126, N276, N94);
and AND2 (N368, N362, N76);
xor XOR2 (N369, N364, N79);
and AND2 (N370, N355, N3);
or OR3 (N371, N369, N25, N367);
or OR2 (N372, N135, N294);
xor XOR2 (N373, N371, N308);
not NOT1 (N374, N368);
buf BUF1 (N375, N373);
or OR4 (N376, N365, N39, N316, N283);
nor NOR2 (N377, N357, N198);
or OR4 (N378, N375, N252, N183, N75);
not NOT1 (N379, N374);
xor XOR2 (N380, N363, N68);
nand NAND2 (N381, N376, N40);
nor NOR4 (N382, N377, N292, N330, N56);
nor NOR4 (N383, N361, N7, N103, N301);
nor NOR3 (N384, N382, N288, N6);
buf BUF1 (N385, N383);
xor XOR2 (N386, N380, N154);
not NOT1 (N387, N385);
and AND2 (N388, N384, N6);
or OR2 (N389, N388, N256);
and AND4 (N390, N366, N63, N183, N309);
xor XOR2 (N391, N389, N272);
nor NOR4 (N392, N391, N287, N33, N77);
and AND3 (N393, N386, N120, N87);
buf BUF1 (N394, N392);
not NOT1 (N395, N372);
xor XOR2 (N396, N378, N191);
not NOT1 (N397, N379);
or OR2 (N398, N390, N304);
nand NAND2 (N399, N387, N380);
buf BUF1 (N400, N381);
nor NOR4 (N401, N395, N250, N399, N160);
not NOT1 (N402, N26);
not NOT1 (N403, N370);
nand NAND3 (N404, N393, N237, N52);
xor XOR2 (N405, N394, N19);
nand NAND4 (N406, N403, N60, N48, N395);
nand NAND2 (N407, N406, N101);
or OR3 (N408, N404, N140, N247);
buf BUF1 (N409, N407);
nand NAND2 (N410, N398, N170);
or OR4 (N411, N410, N305, N317, N131);
endmodule