// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N608,N588,N601,N612,N607,N609,N613,N615,N605,N616;

not NOT1 (N17, N5);
not NOT1 (N18, N10);
not NOT1 (N19, N16);
nor NOR3 (N20, N12, N4, N11);
nor NOR2 (N21, N10, N9);
nand NAND2 (N22, N19, N7);
not NOT1 (N23, N1);
xor XOR2 (N24, N23, N10);
nor NOR2 (N25, N16, N23);
buf BUF1 (N26, N6);
buf BUF1 (N27, N18);
buf BUF1 (N28, N20);
nor NOR3 (N29, N1, N2, N17);
nor NOR4 (N30, N9, N20, N1, N17);
or OR3 (N31, N22, N14, N2);
buf BUF1 (N32, N5);
nand NAND3 (N33, N26, N21, N3);
nor NOR3 (N34, N4, N25, N33);
nor NOR2 (N35, N9, N20);
or OR4 (N36, N5, N14, N14, N33);
not NOT1 (N37, N28);
not NOT1 (N38, N27);
xor XOR2 (N39, N29, N9);
xor XOR2 (N40, N24, N13);
buf BUF1 (N41, N37);
xor XOR2 (N42, N34, N7);
buf BUF1 (N43, N35);
not NOT1 (N44, N31);
buf BUF1 (N45, N30);
nor NOR4 (N46, N39, N40, N35, N11);
xor XOR2 (N47, N38, N1);
xor XOR2 (N48, N42, N21);
not NOT1 (N49, N16);
nand NAND3 (N50, N46, N37, N15);
nand NAND3 (N51, N43, N44, N41);
nor NOR2 (N52, N1, N20);
not NOT1 (N53, N43);
not NOT1 (N54, N48);
nor NOR4 (N55, N50, N10, N28, N18);
not NOT1 (N56, N45);
nand NAND4 (N57, N51, N56, N6, N2);
and AND2 (N58, N12, N38);
or OR3 (N59, N36, N29, N44);
xor XOR2 (N60, N55, N37);
and AND4 (N61, N58, N23, N28, N5);
and AND2 (N62, N53, N27);
buf BUF1 (N63, N54);
xor XOR2 (N64, N49, N54);
buf BUF1 (N65, N59);
or OR2 (N66, N60, N17);
buf BUF1 (N67, N62);
not NOT1 (N68, N65);
and AND4 (N69, N63, N15, N7, N35);
not NOT1 (N70, N66);
not NOT1 (N71, N57);
buf BUF1 (N72, N32);
not NOT1 (N73, N61);
buf BUF1 (N74, N52);
and AND2 (N75, N47, N56);
buf BUF1 (N76, N67);
or OR3 (N77, N72, N67, N56);
nor NOR2 (N78, N64, N70);
or OR4 (N79, N48, N16, N4, N40);
nand NAND4 (N80, N69, N27, N4, N39);
and AND3 (N81, N78, N16, N71);
or OR2 (N82, N53, N36);
nor NOR2 (N83, N68, N21);
not NOT1 (N84, N82);
xor XOR2 (N85, N73, N66);
nand NAND2 (N86, N74, N4);
not NOT1 (N87, N86);
or OR4 (N88, N84, N56, N28, N42);
or OR2 (N89, N77, N84);
not NOT1 (N90, N80);
nor NOR4 (N91, N75, N58, N23, N82);
buf BUF1 (N92, N76);
or OR2 (N93, N81, N51);
not NOT1 (N94, N91);
nor NOR4 (N95, N79, N64, N73, N81);
not NOT1 (N96, N93);
or OR3 (N97, N95, N23, N8);
nor NOR4 (N98, N90, N45, N1, N67);
nor NOR2 (N99, N98, N98);
xor XOR2 (N100, N94, N1);
nand NAND3 (N101, N88, N19, N90);
buf BUF1 (N102, N96);
or OR3 (N103, N83, N6, N77);
nand NAND2 (N104, N99, N5);
or OR3 (N105, N101, N18, N98);
xor XOR2 (N106, N105, N81);
xor XOR2 (N107, N89, N63);
buf BUF1 (N108, N92);
nand NAND3 (N109, N108, N59, N20);
xor XOR2 (N110, N97, N75);
nor NOR3 (N111, N102, N103, N100);
nand NAND2 (N112, N64, N6);
nand NAND4 (N113, N44, N57, N100, N83);
and AND3 (N114, N107, N84, N51);
nor NOR3 (N115, N106, N68, N48);
or OR3 (N116, N109, N44, N27);
and AND4 (N117, N116, N109, N93, N8);
buf BUF1 (N118, N117);
or OR4 (N119, N104, N92, N39, N7);
xor XOR2 (N120, N111, N96);
nor NOR2 (N121, N115, N41);
not NOT1 (N122, N110);
buf BUF1 (N123, N87);
and AND2 (N124, N119, N22);
nand NAND3 (N125, N124, N43, N60);
nor NOR2 (N126, N85, N23);
buf BUF1 (N127, N126);
buf BUF1 (N128, N113);
nand NAND4 (N129, N112, N17, N22, N108);
not NOT1 (N130, N120);
nand NAND4 (N131, N114, N9, N3, N49);
or OR3 (N132, N131, N99, N115);
or OR4 (N133, N122, N64, N11, N91);
not NOT1 (N134, N118);
xor XOR2 (N135, N123, N133);
or OR4 (N136, N72, N79, N97, N35);
nor NOR4 (N137, N121, N110, N42, N119);
xor XOR2 (N138, N137, N133);
buf BUF1 (N139, N136);
nand NAND4 (N140, N135, N76, N103, N48);
nand NAND4 (N141, N130, N71, N60, N17);
not NOT1 (N142, N138);
or OR4 (N143, N134, N21, N93, N31);
or OR4 (N144, N132, N52, N62, N105);
nand NAND3 (N145, N141, N52, N6);
xor XOR2 (N146, N127, N35);
not NOT1 (N147, N145);
xor XOR2 (N148, N144, N30);
buf BUF1 (N149, N129);
xor XOR2 (N150, N125, N42);
nand NAND2 (N151, N143, N122);
nor NOR2 (N152, N148, N63);
buf BUF1 (N153, N150);
not NOT1 (N154, N146);
nor NOR4 (N155, N147, N136, N147, N30);
not NOT1 (N156, N155);
nand NAND3 (N157, N149, N143, N32);
or OR3 (N158, N139, N145, N30);
xor XOR2 (N159, N158, N83);
not NOT1 (N160, N153);
nand NAND4 (N161, N157, N37, N57, N68);
and AND4 (N162, N152, N49, N155, N69);
buf BUF1 (N163, N140);
or OR4 (N164, N163, N59, N118, N42);
and AND4 (N165, N156, N79, N81, N162);
xor XOR2 (N166, N38, N45);
or OR3 (N167, N164, N76, N118);
buf BUF1 (N168, N165);
nor NOR3 (N169, N159, N14, N104);
buf BUF1 (N170, N168);
nand NAND4 (N171, N160, N161, N24, N27);
and AND2 (N172, N102, N53);
xor XOR2 (N173, N170, N139);
and AND4 (N174, N172, N127, N22, N71);
and AND4 (N175, N174, N151, N130, N23);
xor XOR2 (N176, N170, N157);
nor NOR2 (N177, N176, N101);
not NOT1 (N178, N175);
and AND3 (N179, N128, N128, N120);
not NOT1 (N180, N179);
xor XOR2 (N181, N167, N61);
or OR2 (N182, N178, N93);
buf BUF1 (N183, N181);
nor NOR4 (N184, N169, N64, N95, N25);
buf BUF1 (N185, N173);
buf BUF1 (N186, N184);
nor NOR4 (N187, N183, N71, N35, N8);
nand NAND2 (N188, N187, N122);
nand NAND3 (N189, N186, N20, N72);
not NOT1 (N190, N177);
and AND2 (N191, N171, N186);
buf BUF1 (N192, N189);
and AND2 (N193, N192, N191);
buf BUF1 (N194, N164);
and AND4 (N195, N166, N158, N131, N159);
or OR4 (N196, N190, N178, N185, N142);
nor NOR4 (N197, N89, N122, N87, N178);
nor NOR3 (N198, N101, N118, N114);
nor NOR3 (N199, N195, N158, N47);
nand NAND3 (N200, N198, N31, N47);
xor XOR2 (N201, N197, N12);
not NOT1 (N202, N154);
nand NAND2 (N203, N199, N183);
xor XOR2 (N204, N188, N117);
and AND3 (N205, N180, N181, N77);
and AND2 (N206, N193, N119);
or OR2 (N207, N201, N36);
nand NAND2 (N208, N204, N155);
nor NOR4 (N209, N208, N182, N195, N28);
not NOT1 (N210, N165);
buf BUF1 (N211, N209);
nor NOR2 (N212, N207, N199);
nor NOR4 (N213, N210, N136, N205, N97);
not NOT1 (N214, N36);
buf BUF1 (N215, N213);
or OR2 (N216, N206, N96);
or OR2 (N217, N211, N92);
and AND4 (N218, N194, N119, N183, N16);
not NOT1 (N219, N214);
not NOT1 (N220, N196);
xor XOR2 (N221, N220, N144);
not NOT1 (N222, N203);
or OR2 (N223, N202, N187);
xor XOR2 (N224, N212, N76);
and AND2 (N225, N218, N94);
nor NOR3 (N226, N219, N140, N4);
xor XOR2 (N227, N216, N174);
buf BUF1 (N228, N222);
nor NOR2 (N229, N224, N3);
xor XOR2 (N230, N229, N9);
or OR3 (N231, N223, N89, N210);
and AND4 (N232, N228, N145, N209, N98);
buf BUF1 (N233, N217);
not NOT1 (N234, N227);
buf BUF1 (N235, N200);
not NOT1 (N236, N221);
nand NAND4 (N237, N236, N217, N107, N58);
nor NOR3 (N238, N215, N159, N122);
buf BUF1 (N239, N237);
or OR2 (N240, N231, N48);
xor XOR2 (N241, N234, N155);
and AND4 (N242, N232, N199, N192, N34);
or OR2 (N243, N230, N167);
xor XOR2 (N244, N235, N102);
xor XOR2 (N245, N226, N206);
nand NAND4 (N246, N238, N224, N132, N40);
nor NOR2 (N247, N246, N132);
not NOT1 (N248, N242);
and AND2 (N249, N248, N85);
nand NAND2 (N250, N240, N32);
nor NOR4 (N251, N249, N72, N138, N102);
and AND2 (N252, N239, N205);
not NOT1 (N253, N247);
xor XOR2 (N254, N245, N107);
buf BUF1 (N255, N252);
not NOT1 (N256, N233);
or OR2 (N257, N225, N234);
xor XOR2 (N258, N251, N78);
and AND2 (N259, N257, N223);
xor XOR2 (N260, N253, N258);
not NOT1 (N261, N6);
buf BUF1 (N262, N255);
xor XOR2 (N263, N262, N108);
and AND2 (N264, N241, N163);
buf BUF1 (N265, N244);
xor XOR2 (N266, N263, N82);
not NOT1 (N267, N250);
nor NOR2 (N268, N256, N154);
nand NAND2 (N269, N267, N160);
nand NAND3 (N270, N266, N262, N37);
buf BUF1 (N271, N269);
or OR4 (N272, N265, N19, N12, N94);
nand NAND3 (N273, N271, N184, N123);
or OR2 (N274, N268, N238);
nor NOR3 (N275, N274, N260, N138);
and AND2 (N276, N148, N193);
or OR3 (N277, N273, N53, N103);
not NOT1 (N278, N277);
nor NOR2 (N279, N259, N71);
not NOT1 (N280, N272);
nor NOR4 (N281, N270, N168, N120, N10);
nor NOR4 (N282, N280, N213, N209, N50);
nor NOR2 (N283, N279, N67);
nor NOR4 (N284, N283, N84, N137, N38);
not NOT1 (N285, N278);
nand NAND3 (N286, N285, N105, N22);
and AND3 (N287, N276, N155, N130);
and AND3 (N288, N284, N18, N78);
nor NOR4 (N289, N264, N3, N282, N33);
or OR4 (N290, N216, N232, N236, N17);
nor NOR3 (N291, N275, N109, N201);
buf BUF1 (N292, N281);
not NOT1 (N293, N287);
or OR3 (N294, N293, N132, N122);
nor NOR2 (N295, N261, N186);
nand NAND4 (N296, N286, N96, N140, N65);
not NOT1 (N297, N292);
and AND3 (N298, N288, N13, N59);
nor NOR4 (N299, N290, N261, N249, N288);
buf BUF1 (N300, N243);
not NOT1 (N301, N298);
or OR2 (N302, N254, N280);
xor XOR2 (N303, N302, N151);
nor NOR2 (N304, N295, N41);
buf BUF1 (N305, N297);
nor NOR4 (N306, N299, N218, N281, N100);
xor XOR2 (N307, N306, N198);
not NOT1 (N308, N300);
xor XOR2 (N309, N304, N198);
nand NAND3 (N310, N307, N17, N111);
and AND4 (N311, N303, N300, N273, N231);
nor NOR2 (N312, N308, N252);
xor XOR2 (N313, N294, N120);
or OR4 (N314, N296, N113, N287, N93);
nand NAND3 (N315, N309, N291, N103);
nand NAND3 (N316, N161, N128, N134);
nand NAND4 (N317, N311, N33, N305, N170);
and AND2 (N318, N75, N14);
xor XOR2 (N319, N318, N173);
not NOT1 (N320, N314);
xor XOR2 (N321, N312, N62);
buf BUF1 (N322, N310);
not NOT1 (N323, N301);
nand NAND2 (N324, N322, N260);
not NOT1 (N325, N323);
or OR4 (N326, N313, N244, N282, N124);
nand NAND2 (N327, N315, N281);
and AND2 (N328, N327, N96);
nand NAND2 (N329, N324, N307);
nor NOR2 (N330, N317, N95);
or OR2 (N331, N289, N130);
and AND2 (N332, N320, N132);
and AND2 (N333, N316, N183);
nor NOR4 (N334, N333, N212, N263, N270);
buf BUF1 (N335, N319);
buf BUF1 (N336, N332);
nor NOR2 (N337, N331, N128);
xor XOR2 (N338, N326, N229);
or OR4 (N339, N328, N90, N288, N4);
nor NOR3 (N340, N335, N163, N173);
nor NOR3 (N341, N338, N203, N212);
not NOT1 (N342, N334);
and AND3 (N343, N342, N143, N288);
buf BUF1 (N344, N325);
nor NOR4 (N345, N329, N14, N34, N10);
and AND3 (N346, N341, N230, N180);
xor XOR2 (N347, N340, N104);
xor XOR2 (N348, N337, N86);
nand NAND4 (N349, N343, N234, N27, N138);
and AND4 (N350, N336, N27, N162, N327);
nor NOR2 (N351, N344, N119);
or OR4 (N352, N351, N220, N61, N175);
or OR4 (N353, N352, N258, N350, N87);
not NOT1 (N354, N293);
and AND2 (N355, N345, N221);
nand NAND2 (N356, N346, N110);
and AND3 (N357, N349, N150, N104);
not NOT1 (N358, N330);
not NOT1 (N359, N347);
xor XOR2 (N360, N359, N16);
nand NAND3 (N361, N356, N249, N249);
not NOT1 (N362, N357);
nor NOR4 (N363, N321, N171, N10, N24);
nor NOR4 (N364, N348, N352, N145, N101);
not NOT1 (N365, N362);
nor NOR2 (N366, N354, N229);
nand NAND4 (N367, N358, N349, N173, N169);
xor XOR2 (N368, N365, N232);
buf BUF1 (N369, N360);
nand NAND4 (N370, N361, N81, N167, N204);
or OR3 (N371, N367, N309, N174);
nand NAND2 (N372, N364, N361);
not NOT1 (N373, N370);
or OR2 (N374, N353, N200);
buf BUF1 (N375, N371);
and AND4 (N376, N366, N239, N36, N13);
buf BUF1 (N377, N373);
nor NOR4 (N378, N363, N85, N299, N24);
not NOT1 (N379, N377);
xor XOR2 (N380, N379, N23);
nor NOR3 (N381, N376, N354, N290);
and AND4 (N382, N381, N208, N9, N110);
and AND2 (N383, N368, N124);
and AND3 (N384, N375, N108, N57);
or OR4 (N385, N378, N155, N35, N264);
nand NAND4 (N386, N383, N154, N221, N178);
and AND2 (N387, N339, N15);
buf BUF1 (N388, N369);
and AND2 (N389, N386, N78);
and AND3 (N390, N380, N104, N116);
xor XOR2 (N391, N390, N316);
nand NAND4 (N392, N355, N120, N11, N26);
or OR3 (N393, N389, N283, N351);
buf BUF1 (N394, N374);
nor NOR4 (N395, N391, N112, N336, N85);
buf BUF1 (N396, N382);
not NOT1 (N397, N394);
nor NOR2 (N398, N396, N173);
nand NAND2 (N399, N392, N155);
not NOT1 (N400, N372);
buf BUF1 (N401, N387);
not NOT1 (N402, N399);
xor XOR2 (N403, N397, N327);
nand NAND3 (N404, N403, N280, N269);
not NOT1 (N405, N395);
xor XOR2 (N406, N402, N191);
and AND2 (N407, N384, N371);
xor XOR2 (N408, N385, N154);
xor XOR2 (N409, N407, N198);
buf BUF1 (N410, N405);
or OR4 (N411, N400, N332, N127, N378);
buf BUF1 (N412, N401);
or OR3 (N413, N409, N191, N342);
not NOT1 (N414, N404);
not NOT1 (N415, N414);
nand NAND4 (N416, N410, N83, N360, N381);
nor NOR2 (N417, N412, N199);
and AND4 (N418, N406, N350, N297, N298);
xor XOR2 (N419, N415, N64);
or OR4 (N420, N418, N152, N314, N233);
or OR2 (N421, N416, N153);
buf BUF1 (N422, N417);
buf BUF1 (N423, N421);
or OR2 (N424, N393, N132);
nor NOR4 (N425, N420, N85, N235, N89);
and AND2 (N426, N413, N169);
xor XOR2 (N427, N422, N383);
or OR2 (N428, N424, N258);
or OR2 (N429, N426, N345);
and AND2 (N430, N388, N54);
or OR2 (N431, N398, N247);
nand NAND3 (N432, N419, N10, N245);
or OR4 (N433, N432, N423, N399, N332);
xor XOR2 (N434, N249, N426);
buf BUF1 (N435, N425);
or OR2 (N436, N429, N414);
nor NOR3 (N437, N427, N194, N59);
or OR2 (N438, N437, N191);
and AND2 (N439, N428, N112);
nand NAND4 (N440, N411, N160, N8, N28);
nand NAND2 (N441, N436, N180);
not NOT1 (N442, N430);
nand NAND3 (N443, N435, N101, N232);
or OR2 (N444, N441, N104);
not NOT1 (N445, N443);
nand NAND2 (N446, N433, N122);
not NOT1 (N447, N434);
not NOT1 (N448, N445);
buf BUF1 (N449, N446);
and AND4 (N450, N442, N200, N104, N116);
buf BUF1 (N451, N448);
and AND4 (N452, N450, N303, N369, N283);
buf BUF1 (N453, N438);
and AND2 (N454, N440, N403);
nor NOR3 (N455, N451, N220, N266);
buf BUF1 (N456, N452);
or OR2 (N457, N431, N354);
xor XOR2 (N458, N439, N275);
buf BUF1 (N459, N447);
buf BUF1 (N460, N457);
and AND4 (N461, N444, N213, N218, N313);
nor NOR2 (N462, N460, N143);
xor XOR2 (N463, N449, N458);
and AND4 (N464, N8, N442, N379, N440);
and AND4 (N465, N454, N294, N441, N215);
or OR3 (N466, N463, N138, N265);
nor NOR4 (N467, N453, N354, N460, N342);
or OR3 (N468, N462, N271, N330);
buf BUF1 (N469, N455);
or OR4 (N470, N466, N8, N57, N61);
buf BUF1 (N471, N470);
not NOT1 (N472, N468);
not NOT1 (N473, N456);
and AND2 (N474, N467, N212);
xor XOR2 (N475, N408, N9);
nor NOR3 (N476, N474, N240, N235);
nor NOR4 (N477, N461, N221, N223, N280);
not NOT1 (N478, N475);
not NOT1 (N479, N473);
buf BUF1 (N480, N471);
and AND2 (N481, N476, N299);
nor NOR2 (N482, N478, N116);
or OR4 (N483, N459, N185, N53, N479);
xor XOR2 (N484, N464, N84);
and AND2 (N485, N457, N379);
nand NAND4 (N486, N469, N480, N248, N345);
nor NOR4 (N487, N156, N282, N385, N285);
nand NAND4 (N488, N481, N352, N36, N201);
buf BUF1 (N489, N477);
or OR4 (N490, N482, N309, N258, N437);
nor NOR2 (N491, N487, N248);
nand NAND3 (N492, N465, N378, N74);
nor NOR4 (N493, N483, N188, N56, N308);
and AND4 (N494, N485, N275, N273, N325);
and AND4 (N495, N493, N55, N394, N449);
nor NOR4 (N496, N484, N446, N361, N213);
or OR4 (N497, N472, N309, N428, N166);
buf BUF1 (N498, N489);
xor XOR2 (N499, N491, N182);
buf BUF1 (N500, N488);
buf BUF1 (N501, N499);
not NOT1 (N502, N501);
nand NAND2 (N503, N490, N395);
or OR3 (N504, N500, N221, N83);
nand NAND2 (N505, N496, N285);
or OR3 (N506, N503, N226, N100);
nor NOR3 (N507, N502, N88, N476);
buf BUF1 (N508, N495);
buf BUF1 (N509, N506);
or OR2 (N510, N486, N317);
xor XOR2 (N511, N510, N185);
nor NOR2 (N512, N508, N164);
not NOT1 (N513, N494);
not NOT1 (N514, N507);
xor XOR2 (N515, N498, N430);
not NOT1 (N516, N511);
nand NAND4 (N517, N516, N429, N234, N488);
or OR4 (N518, N512, N252, N429, N133);
and AND3 (N519, N509, N111, N264);
and AND4 (N520, N504, N464, N389, N518);
buf BUF1 (N521, N74);
buf BUF1 (N522, N515);
and AND4 (N523, N505, N489, N292, N214);
and AND4 (N524, N519, N492, N283, N361);
and AND3 (N525, N434, N301, N517);
nor NOR3 (N526, N328, N343, N388);
nor NOR3 (N527, N523, N204, N130);
xor XOR2 (N528, N520, N290);
or OR2 (N529, N527, N285);
buf BUF1 (N530, N529);
and AND3 (N531, N522, N17, N503);
not NOT1 (N532, N514);
nor NOR3 (N533, N521, N426, N363);
and AND4 (N534, N497, N292, N66, N462);
xor XOR2 (N535, N531, N145);
buf BUF1 (N536, N526);
nand NAND4 (N537, N535, N197, N272, N143);
and AND4 (N538, N536, N353, N379, N412);
or OR3 (N539, N524, N110, N310);
buf BUF1 (N540, N537);
xor XOR2 (N541, N538, N28);
and AND4 (N542, N513, N271, N419, N352);
nor NOR3 (N543, N542, N537, N306);
and AND2 (N544, N541, N210);
xor XOR2 (N545, N544, N525);
or OR2 (N546, N36, N233);
or OR4 (N547, N539, N92, N54, N251);
not NOT1 (N548, N530);
buf BUF1 (N549, N547);
nand NAND2 (N550, N540, N419);
and AND2 (N551, N533, N452);
buf BUF1 (N552, N545);
or OR2 (N553, N546, N211);
nand NAND4 (N554, N553, N455, N138, N112);
not NOT1 (N555, N548);
nand NAND2 (N556, N551, N303);
xor XOR2 (N557, N555, N90);
nor NOR4 (N558, N557, N479, N510, N421);
nor NOR3 (N559, N554, N42, N46);
not NOT1 (N560, N532);
not NOT1 (N561, N549);
xor XOR2 (N562, N543, N499);
nor NOR3 (N563, N559, N363, N488);
or OR3 (N564, N561, N288, N492);
not NOT1 (N565, N552);
and AND3 (N566, N556, N521, N298);
nor NOR3 (N567, N558, N435, N117);
nand NAND3 (N568, N562, N99, N389);
not NOT1 (N569, N528);
nor NOR4 (N570, N563, N458, N59, N361);
not NOT1 (N571, N564);
not NOT1 (N572, N550);
not NOT1 (N573, N565);
nor NOR2 (N574, N570, N380);
xor XOR2 (N575, N574, N377);
not NOT1 (N576, N566);
nor NOR4 (N577, N560, N211, N477, N374);
nor NOR2 (N578, N572, N403);
and AND3 (N579, N577, N496, N441);
xor XOR2 (N580, N567, N311);
nor NOR2 (N581, N580, N399);
xor XOR2 (N582, N568, N323);
or OR3 (N583, N578, N550, N67);
nand NAND3 (N584, N534, N94, N210);
nand NAND3 (N585, N576, N574, N283);
nor NOR4 (N586, N571, N527, N332, N294);
and AND3 (N587, N586, N299, N87);
nand NAND3 (N588, N581, N202, N378);
and AND2 (N589, N575, N138);
buf BUF1 (N590, N584);
nor NOR4 (N591, N590, N134, N110, N424);
or OR2 (N592, N579, N238);
buf BUF1 (N593, N589);
not NOT1 (N594, N583);
or OR4 (N595, N587, N227, N368, N157);
nand NAND4 (N596, N573, N305, N362, N489);
nor NOR2 (N597, N594, N191);
nor NOR3 (N598, N569, N225, N459);
or OR4 (N599, N597, N506, N151, N191);
nand NAND3 (N600, N591, N310, N137);
nor NOR3 (N601, N595, N526, N385);
xor XOR2 (N602, N585, N84);
nor NOR2 (N603, N602, N9);
nand NAND4 (N604, N592, N251, N171, N586);
buf BUF1 (N605, N582);
xor XOR2 (N606, N598, N14);
nor NOR2 (N607, N596, N394);
and AND2 (N608, N600, N570);
buf BUF1 (N609, N604);
not NOT1 (N610, N599);
nor NOR2 (N611, N606, N570);
xor XOR2 (N612, N611, N174);
nand NAND3 (N613, N610, N535, N168);
and AND2 (N614, N593, N150);
buf BUF1 (N615, N614);
buf BUF1 (N616, N603);
endmodule