// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N2510,N2504,N2521,N2493,N2520,N2517,N2509,N2516,N2514,N2522;

nor NOR3 (N23, N21, N12, N14);
xor XOR2 (N24, N17, N18);
nor NOR3 (N25, N13, N23, N14);
xor XOR2 (N26, N25, N19);
nor NOR2 (N27, N2, N22);
or OR3 (N28, N18, N24, N10);
or OR3 (N29, N25, N9, N2);
nor NOR4 (N30, N21, N12, N7, N21);
not NOT1 (N31, N10);
nand NAND2 (N32, N16, N25);
nand NAND2 (N33, N26, N32);
nor NOR2 (N34, N4, N19);
buf BUF1 (N35, N17);
not NOT1 (N36, N10);
and AND2 (N37, N29, N21);
not NOT1 (N38, N30);
not NOT1 (N39, N37);
xor XOR2 (N40, N38, N10);
xor XOR2 (N41, N25, N34);
nor NOR3 (N42, N1, N13, N27);
xor XOR2 (N43, N40, N14);
not NOT1 (N44, N10);
buf BUF1 (N45, N31);
buf BUF1 (N46, N41);
xor XOR2 (N47, N46, N9);
buf BUF1 (N48, N33);
buf BUF1 (N49, N39);
or OR4 (N50, N49, N17, N41, N21);
or OR3 (N51, N42, N50, N35);
and AND2 (N52, N44, N22);
or OR2 (N53, N45, N40);
or OR2 (N54, N30, N19);
nand NAND2 (N55, N12, N48);
not NOT1 (N56, N9);
not NOT1 (N57, N47);
or OR2 (N58, N54, N1);
buf BUF1 (N59, N58);
xor XOR2 (N60, N53, N25);
xor XOR2 (N61, N57, N37);
and AND3 (N62, N52, N48, N11);
buf BUF1 (N63, N28);
xor XOR2 (N64, N61, N34);
not NOT1 (N65, N43);
or OR2 (N66, N60, N60);
nor NOR3 (N67, N64, N42, N13);
nor NOR3 (N68, N67, N5, N2);
or OR3 (N69, N65, N39, N14);
not NOT1 (N70, N66);
or OR2 (N71, N68, N37);
buf BUF1 (N72, N63);
and AND3 (N73, N59, N55, N57);
nor NOR4 (N74, N21, N38, N57, N65);
buf BUF1 (N75, N56);
not NOT1 (N76, N75);
or OR3 (N77, N70, N66, N45);
or OR2 (N78, N71, N23);
nor NOR3 (N79, N73, N58, N56);
nand NAND4 (N80, N69, N3, N49, N61);
nor NOR2 (N81, N77, N8);
xor XOR2 (N82, N79, N21);
not NOT1 (N83, N51);
not NOT1 (N84, N83);
nor NOR4 (N85, N84, N2, N63, N10);
or OR4 (N86, N85, N44, N80, N31);
nor NOR4 (N87, N25, N70, N74, N58);
buf BUF1 (N88, N26);
not NOT1 (N89, N76);
and AND2 (N90, N72, N48);
and AND4 (N91, N81, N12, N50, N35);
nand NAND2 (N92, N86, N36);
nor NOR4 (N93, N41, N32, N92, N89);
not NOT1 (N94, N66);
not NOT1 (N95, N8);
xor XOR2 (N96, N78, N46);
xor XOR2 (N97, N91, N50);
buf BUF1 (N98, N87);
nand NAND3 (N99, N96, N20, N80);
buf BUF1 (N100, N88);
buf BUF1 (N101, N90);
buf BUF1 (N102, N99);
nor NOR2 (N103, N102, N47);
nand NAND3 (N104, N94, N65, N8);
buf BUF1 (N105, N95);
not NOT1 (N106, N103);
not NOT1 (N107, N82);
xor XOR2 (N108, N98, N95);
nand NAND2 (N109, N97, N81);
buf BUF1 (N110, N105);
xor XOR2 (N111, N62, N91);
xor XOR2 (N112, N110, N104);
and AND4 (N113, N91, N83, N53, N38);
buf BUF1 (N114, N108);
nand NAND3 (N115, N107, N71, N104);
or OR2 (N116, N101, N83);
nand NAND3 (N117, N116, N85, N40);
not NOT1 (N118, N93);
not NOT1 (N119, N115);
not NOT1 (N120, N113);
and AND3 (N121, N106, N42, N74);
nor NOR3 (N122, N111, N69, N27);
not NOT1 (N123, N117);
buf BUF1 (N124, N121);
nor NOR4 (N125, N123, N41, N26, N36);
buf BUF1 (N126, N114);
nand NAND4 (N127, N122, N3, N85, N6);
xor XOR2 (N128, N112, N102);
buf BUF1 (N129, N124);
not NOT1 (N130, N127);
or OR4 (N131, N126, N22, N120, N13);
and AND3 (N132, N92, N104, N79);
xor XOR2 (N133, N118, N10);
nor NOR3 (N134, N132, N27, N121);
xor XOR2 (N135, N119, N110);
and AND2 (N136, N100, N53);
nand NAND4 (N137, N130, N49, N36, N30);
and AND4 (N138, N133, N80, N70, N10);
nor NOR2 (N139, N125, N32);
or OR2 (N140, N128, N5);
not NOT1 (N141, N140);
nand NAND2 (N142, N129, N59);
not NOT1 (N143, N109);
xor XOR2 (N144, N131, N66);
or OR3 (N145, N139, N80, N78);
nand NAND3 (N146, N138, N47, N52);
xor XOR2 (N147, N142, N84);
not NOT1 (N148, N145);
buf BUF1 (N149, N134);
nor NOR3 (N150, N149, N129, N99);
xor XOR2 (N151, N136, N130);
nor NOR2 (N152, N141, N4);
nor NOR4 (N153, N147, N94, N100, N92);
xor XOR2 (N154, N153, N114);
and AND3 (N155, N154, N78, N70);
not NOT1 (N156, N151);
or OR2 (N157, N146, N140);
not NOT1 (N158, N135);
not NOT1 (N159, N152);
and AND3 (N160, N159, N133, N49);
or OR4 (N161, N148, N53, N101, N104);
xor XOR2 (N162, N161, N72);
and AND2 (N163, N156, N64);
xor XOR2 (N164, N163, N50);
xor XOR2 (N165, N158, N19);
nand NAND3 (N166, N157, N126, N18);
or OR4 (N167, N164, N77, N134, N139);
xor XOR2 (N168, N155, N40);
nand NAND2 (N169, N165, N158);
xor XOR2 (N170, N162, N59);
nand NAND2 (N171, N137, N12);
or OR3 (N172, N143, N35, N121);
not NOT1 (N173, N144);
buf BUF1 (N174, N167);
nor NOR3 (N175, N172, N44, N162);
and AND2 (N176, N160, N140);
nor NOR2 (N177, N168, N146);
xor XOR2 (N178, N176, N15);
not NOT1 (N179, N171);
buf BUF1 (N180, N150);
xor XOR2 (N181, N175, N2);
not NOT1 (N182, N174);
xor XOR2 (N183, N170, N14);
buf BUF1 (N184, N173);
nand NAND4 (N185, N184, N155, N92, N21);
buf BUF1 (N186, N177);
not NOT1 (N187, N178);
xor XOR2 (N188, N180, N134);
and AND4 (N189, N182, N36, N60, N40);
not NOT1 (N190, N179);
nor NOR4 (N191, N181, N51, N176, N154);
and AND2 (N192, N169, N12);
not NOT1 (N193, N183);
xor XOR2 (N194, N193, N77);
or OR4 (N195, N188, N108, N184, N186);
not NOT1 (N196, N72);
xor XOR2 (N197, N191, N93);
nor NOR4 (N198, N197, N158, N37, N178);
and AND4 (N199, N195, N4, N19, N26);
not NOT1 (N200, N196);
not NOT1 (N201, N192);
buf BUF1 (N202, N190);
or OR4 (N203, N185, N193, N64, N147);
nand NAND3 (N204, N202, N170, N36);
nand NAND2 (N205, N204, N3);
nor NOR3 (N206, N166, N23, N188);
buf BUF1 (N207, N194);
xor XOR2 (N208, N201, N109);
buf BUF1 (N209, N208);
not NOT1 (N210, N198);
and AND3 (N211, N205, N61, N115);
nand NAND3 (N212, N203, N176, N158);
nand NAND3 (N213, N206, N165, N64);
xor XOR2 (N214, N207, N207);
not NOT1 (N215, N213);
and AND4 (N216, N200, N161, N158, N137);
nand NAND3 (N217, N211, N89, N5);
nor NOR2 (N218, N210, N216);
and AND3 (N219, N192, N7, N119);
xor XOR2 (N220, N212, N102);
xor XOR2 (N221, N209, N191);
buf BUF1 (N222, N187);
buf BUF1 (N223, N215);
nor NOR2 (N224, N221, N176);
and AND3 (N225, N199, N205, N166);
nand NAND4 (N226, N223, N220, N124, N179);
or OR3 (N227, N137, N66, N158);
nor NOR3 (N228, N189, N10, N18);
nand NAND4 (N229, N228, N213, N220, N119);
xor XOR2 (N230, N229, N104);
not NOT1 (N231, N222);
and AND4 (N232, N219, N169, N1, N50);
xor XOR2 (N233, N224, N189);
and AND3 (N234, N226, N17, N40);
xor XOR2 (N235, N217, N29);
nor NOR4 (N236, N230, N41, N76, N158);
nand NAND2 (N237, N233, N131);
nor NOR2 (N238, N214, N32);
xor XOR2 (N239, N227, N74);
not NOT1 (N240, N238);
not NOT1 (N241, N232);
xor XOR2 (N242, N237, N195);
and AND3 (N243, N240, N81, N35);
xor XOR2 (N244, N243, N204);
xor XOR2 (N245, N234, N213);
xor XOR2 (N246, N235, N210);
buf BUF1 (N247, N236);
xor XOR2 (N248, N246, N218);
nand NAND3 (N249, N186, N186, N34);
nand NAND2 (N250, N231, N194);
or OR2 (N251, N248, N64);
buf BUF1 (N252, N241);
or OR3 (N253, N249, N44, N139);
nand NAND3 (N254, N252, N8, N13);
and AND4 (N255, N247, N89, N117, N124);
nand NAND4 (N256, N253, N137, N111, N64);
xor XOR2 (N257, N239, N157);
xor XOR2 (N258, N254, N224);
and AND3 (N259, N242, N171, N51);
nand NAND2 (N260, N255, N186);
or OR3 (N261, N259, N198, N55);
and AND2 (N262, N225, N99);
xor XOR2 (N263, N251, N21);
nand NAND4 (N264, N245, N256, N215, N190);
not NOT1 (N265, N248);
nand NAND2 (N266, N263, N173);
xor XOR2 (N267, N250, N133);
buf BUF1 (N268, N265);
nand NAND2 (N269, N260, N69);
not NOT1 (N270, N264);
not NOT1 (N271, N261);
not NOT1 (N272, N244);
or OR3 (N273, N266, N69, N121);
nor NOR2 (N274, N273, N192);
not NOT1 (N275, N269);
not NOT1 (N276, N270);
or OR3 (N277, N275, N160, N159);
buf BUF1 (N278, N268);
nand NAND2 (N279, N271, N97);
or OR2 (N280, N279, N271);
not NOT1 (N281, N262);
xor XOR2 (N282, N280, N189);
not NOT1 (N283, N278);
buf BUF1 (N284, N277);
buf BUF1 (N285, N258);
nand NAND2 (N286, N281, N107);
buf BUF1 (N287, N276);
nor NOR3 (N288, N283, N159, N46);
nand NAND3 (N289, N288, N9, N181);
xor XOR2 (N290, N274, N188);
buf BUF1 (N291, N287);
buf BUF1 (N292, N272);
nand NAND3 (N293, N284, N79, N222);
xor XOR2 (N294, N282, N287);
nand NAND3 (N295, N291, N17, N111);
nor NOR3 (N296, N293, N57, N167);
nand NAND3 (N297, N285, N225, N15);
nand NAND3 (N298, N292, N224, N286);
buf BUF1 (N299, N150);
xor XOR2 (N300, N294, N243);
or OR4 (N301, N257, N204, N139, N270);
or OR4 (N302, N298, N127, N10, N93);
or OR4 (N303, N267, N112, N204, N215);
nor NOR4 (N304, N303, N294, N146, N9);
and AND3 (N305, N304, N277, N192);
nand NAND4 (N306, N300, N1, N295, N28);
and AND2 (N307, N209, N272);
nand NAND4 (N308, N306, N277, N119, N267);
buf BUF1 (N309, N297);
and AND3 (N310, N305, N37, N15);
xor XOR2 (N311, N299, N259);
nor NOR4 (N312, N310, N109, N97, N86);
nor NOR3 (N313, N309, N249, N30);
or OR4 (N314, N308, N197, N89, N229);
xor XOR2 (N315, N313, N72);
or OR2 (N316, N307, N258);
buf BUF1 (N317, N312);
xor XOR2 (N318, N302, N8);
nor NOR3 (N319, N317, N22, N83);
not NOT1 (N320, N315);
nand NAND4 (N321, N289, N199, N94, N265);
nand NAND3 (N322, N301, N137, N89);
buf BUF1 (N323, N318);
not NOT1 (N324, N319);
nand NAND4 (N325, N314, N267, N60, N70);
buf BUF1 (N326, N324);
and AND2 (N327, N290, N31);
buf BUF1 (N328, N320);
and AND3 (N329, N328, N295, N73);
nand NAND4 (N330, N327, N216, N215, N264);
nor NOR4 (N331, N330, N219, N53, N202);
not NOT1 (N332, N325);
not NOT1 (N333, N321);
or OR2 (N334, N326, N328);
or OR2 (N335, N334, N27);
xor XOR2 (N336, N332, N12);
not NOT1 (N337, N296);
xor XOR2 (N338, N322, N36);
and AND4 (N339, N329, N186, N211, N261);
xor XOR2 (N340, N311, N65);
xor XOR2 (N341, N339, N226);
and AND4 (N342, N335, N168, N161, N157);
nor NOR3 (N343, N323, N25, N306);
and AND2 (N344, N338, N5);
buf BUF1 (N345, N333);
buf BUF1 (N346, N331);
nor NOR3 (N347, N316, N233, N108);
nor NOR3 (N348, N344, N54, N174);
or OR4 (N349, N341, N334, N177, N238);
not NOT1 (N350, N347);
or OR4 (N351, N346, N146, N140, N71);
buf BUF1 (N352, N336);
not NOT1 (N353, N337);
buf BUF1 (N354, N348);
nor NOR2 (N355, N345, N244);
buf BUF1 (N356, N342);
nor NOR3 (N357, N356, N52, N336);
and AND3 (N358, N352, N159, N178);
or OR3 (N359, N350, N342, N11);
nor NOR2 (N360, N359, N46);
buf BUF1 (N361, N357);
not NOT1 (N362, N349);
nand NAND3 (N363, N351, N49, N180);
nand NAND4 (N364, N355, N158, N251, N58);
or OR3 (N365, N358, N254, N115);
buf BUF1 (N366, N362);
not NOT1 (N367, N366);
xor XOR2 (N368, N363, N189);
not NOT1 (N369, N353);
nand NAND2 (N370, N369, N241);
nor NOR2 (N371, N340, N254);
not NOT1 (N372, N361);
not NOT1 (N373, N371);
nand NAND2 (N374, N373, N204);
or OR3 (N375, N365, N348, N374);
nor NOR2 (N376, N285, N275);
xor XOR2 (N377, N372, N326);
nand NAND2 (N378, N370, N91);
and AND3 (N379, N376, N106, N15);
and AND4 (N380, N367, N345, N167, N365);
nand NAND4 (N381, N360, N113, N369, N7);
nor NOR4 (N382, N379, N194, N106, N304);
or OR2 (N383, N380, N63);
nor NOR3 (N384, N364, N179, N267);
buf BUF1 (N385, N377);
nor NOR2 (N386, N385, N238);
and AND2 (N387, N386, N140);
buf BUF1 (N388, N381);
buf BUF1 (N389, N343);
and AND4 (N390, N383, N187, N317, N386);
buf BUF1 (N391, N390);
xor XOR2 (N392, N389, N321);
or OR2 (N393, N382, N344);
not NOT1 (N394, N392);
xor XOR2 (N395, N378, N289);
nand NAND3 (N396, N354, N49, N156);
not NOT1 (N397, N388);
nand NAND3 (N398, N395, N319, N86);
and AND4 (N399, N384, N244, N249, N288);
and AND4 (N400, N391, N100, N327, N314);
nor NOR4 (N401, N368, N354, N92, N164);
and AND2 (N402, N397, N269);
buf BUF1 (N403, N400);
buf BUF1 (N404, N401);
buf BUF1 (N405, N387);
xor XOR2 (N406, N402, N247);
not NOT1 (N407, N406);
buf BUF1 (N408, N405);
xor XOR2 (N409, N407, N334);
nor NOR3 (N410, N396, N143, N261);
xor XOR2 (N411, N393, N355);
or OR3 (N412, N411, N4, N336);
nand NAND3 (N413, N412, N370, N304);
or OR4 (N414, N394, N203, N210, N303);
nor NOR4 (N415, N410, N301, N311, N53);
and AND4 (N416, N414, N179, N109, N157);
buf BUF1 (N417, N415);
not NOT1 (N418, N408);
buf BUF1 (N419, N409);
and AND4 (N420, N419, N297, N187, N328);
nor NOR2 (N421, N404, N404);
not NOT1 (N422, N399);
nor NOR4 (N423, N420, N76, N211, N132);
not NOT1 (N424, N417);
not NOT1 (N425, N416);
and AND4 (N426, N418, N356, N152, N150);
xor XOR2 (N427, N426, N9);
not NOT1 (N428, N413);
buf BUF1 (N429, N424);
not NOT1 (N430, N427);
and AND3 (N431, N421, N394, N363);
and AND4 (N432, N422, N155, N388, N136);
buf BUF1 (N433, N428);
xor XOR2 (N434, N433, N321);
buf BUF1 (N435, N398);
buf BUF1 (N436, N434);
nor NOR2 (N437, N432, N255);
or OR4 (N438, N430, N223, N280, N377);
not NOT1 (N439, N429);
nand NAND4 (N440, N425, N106, N281, N88);
nand NAND3 (N441, N423, N337, N192);
buf BUF1 (N442, N438);
nor NOR2 (N443, N437, N434);
nand NAND2 (N444, N375, N171);
nor NOR4 (N445, N436, N310, N406, N147);
or OR3 (N446, N445, N298, N54);
xor XOR2 (N447, N439, N173);
nor NOR3 (N448, N442, N259, N415);
and AND4 (N449, N440, N20, N103, N260);
or OR3 (N450, N449, N223, N114);
not NOT1 (N451, N403);
not NOT1 (N452, N451);
not NOT1 (N453, N447);
buf BUF1 (N454, N452);
not NOT1 (N455, N443);
nor NOR2 (N456, N453, N160);
xor XOR2 (N457, N448, N264);
xor XOR2 (N458, N444, N50);
nand NAND2 (N459, N441, N343);
xor XOR2 (N460, N458, N140);
xor XOR2 (N461, N456, N70);
nor NOR4 (N462, N435, N75, N333, N445);
and AND3 (N463, N462, N138, N145);
not NOT1 (N464, N461);
nor NOR2 (N465, N463, N461);
nor NOR3 (N466, N457, N362, N267);
nor NOR4 (N467, N455, N285, N252, N159);
nor NOR3 (N468, N459, N213, N49);
nor NOR2 (N469, N465, N190);
buf BUF1 (N470, N460);
xor XOR2 (N471, N431, N289);
or OR2 (N472, N470, N444);
buf BUF1 (N473, N472);
nand NAND2 (N474, N468, N220);
xor XOR2 (N475, N469, N233);
nand NAND2 (N476, N454, N419);
nor NOR3 (N477, N466, N382, N84);
and AND2 (N478, N471, N128);
or OR4 (N479, N467, N169, N72, N137);
nand NAND4 (N480, N474, N383, N371, N252);
nand NAND3 (N481, N473, N389, N135);
nor NOR3 (N482, N476, N210, N432);
or OR2 (N483, N450, N457);
buf BUF1 (N484, N478);
buf BUF1 (N485, N484);
xor XOR2 (N486, N479, N481);
nor NOR4 (N487, N421, N138, N64, N105);
and AND3 (N488, N480, N223, N387);
nand NAND3 (N489, N488, N457, N473);
or OR2 (N490, N482, N87);
nand NAND3 (N491, N483, N178, N47);
and AND2 (N492, N486, N364);
and AND2 (N493, N475, N474);
and AND3 (N494, N487, N45, N305);
nand NAND2 (N495, N489, N53);
not NOT1 (N496, N477);
not NOT1 (N497, N494);
nor NOR2 (N498, N485, N106);
and AND4 (N499, N496, N237, N434, N482);
buf BUF1 (N500, N498);
or OR4 (N501, N492, N464, N159, N138);
nand NAND2 (N502, N496, N66);
or OR2 (N503, N490, N407);
xor XOR2 (N504, N497, N401);
xor XOR2 (N505, N503, N330);
buf BUF1 (N506, N501);
nand NAND3 (N507, N495, N14, N424);
xor XOR2 (N508, N499, N480);
xor XOR2 (N509, N500, N176);
nor NOR2 (N510, N508, N492);
nor NOR3 (N511, N446, N342, N409);
nor NOR2 (N512, N510, N117);
and AND2 (N513, N493, N265);
and AND2 (N514, N502, N136);
nand NAND2 (N515, N491, N255);
nor NOR2 (N516, N507, N103);
or OR2 (N517, N512, N20);
not NOT1 (N518, N515);
nor NOR2 (N519, N506, N133);
not NOT1 (N520, N505);
and AND2 (N521, N519, N138);
buf BUF1 (N522, N514);
or OR2 (N523, N513, N207);
buf BUF1 (N524, N523);
not NOT1 (N525, N509);
not NOT1 (N526, N518);
or OR3 (N527, N525, N25, N45);
nand NAND4 (N528, N516, N402, N135, N244);
not NOT1 (N529, N528);
not NOT1 (N530, N526);
and AND4 (N531, N524, N101, N81, N454);
xor XOR2 (N532, N517, N122);
or OR2 (N533, N532, N145);
and AND3 (N534, N504, N118, N435);
xor XOR2 (N535, N527, N351);
and AND3 (N536, N530, N216, N204);
xor XOR2 (N537, N536, N399);
xor XOR2 (N538, N521, N21);
not NOT1 (N539, N538);
nor NOR4 (N540, N537, N30, N460, N140);
buf BUF1 (N541, N511);
xor XOR2 (N542, N541, N441);
nor NOR2 (N543, N522, N223);
and AND3 (N544, N529, N334, N179);
nand NAND4 (N545, N534, N535, N373, N104);
and AND3 (N546, N124, N452, N281);
nor NOR4 (N547, N543, N479, N424, N512);
not NOT1 (N548, N540);
not NOT1 (N549, N545);
buf BUF1 (N550, N549);
not NOT1 (N551, N546);
nand NAND2 (N552, N539, N306);
not NOT1 (N553, N520);
nand NAND2 (N554, N552, N242);
not NOT1 (N555, N531);
buf BUF1 (N556, N554);
or OR3 (N557, N544, N329, N468);
not NOT1 (N558, N553);
nand NAND4 (N559, N551, N180, N203, N75);
nand NAND4 (N560, N555, N109, N275, N180);
and AND2 (N561, N548, N480);
xor XOR2 (N562, N542, N376);
nand NAND3 (N563, N558, N262, N117);
not NOT1 (N564, N563);
nand NAND2 (N565, N560, N309);
xor XOR2 (N566, N564, N388);
and AND2 (N567, N556, N73);
and AND2 (N568, N565, N116);
buf BUF1 (N569, N550);
nor NOR4 (N570, N547, N557, N207, N25);
not NOT1 (N571, N393);
buf BUF1 (N572, N562);
or OR4 (N573, N569, N449, N291, N262);
not NOT1 (N574, N573);
and AND4 (N575, N559, N524, N538, N46);
xor XOR2 (N576, N566, N465);
buf BUF1 (N577, N572);
xor XOR2 (N578, N533, N293);
nand NAND2 (N579, N574, N556);
nand NAND4 (N580, N561, N345, N9, N448);
xor XOR2 (N581, N579, N87);
or OR2 (N582, N575, N109);
or OR3 (N583, N576, N321, N236);
buf BUF1 (N584, N577);
nor NOR3 (N585, N571, N88, N392);
or OR4 (N586, N582, N344, N402, N282);
or OR2 (N587, N578, N348);
or OR4 (N588, N570, N171, N218, N337);
buf BUF1 (N589, N567);
xor XOR2 (N590, N585, N210);
or OR2 (N591, N583, N526);
nand NAND2 (N592, N589, N120);
or OR4 (N593, N592, N136, N557, N281);
buf BUF1 (N594, N588);
nand NAND3 (N595, N590, N44, N338);
buf BUF1 (N596, N568);
and AND2 (N597, N593, N486);
and AND3 (N598, N591, N133, N563);
nand NAND4 (N599, N584, N122, N226, N410);
or OR4 (N600, N581, N542, N232, N128);
or OR4 (N601, N597, N469, N100, N98);
nor NOR2 (N602, N599, N492);
not NOT1 (N603, N594);
xor XOR2 (N604, N595, N513);
xor XOR2 (N605, N600, N140);
nor NOR3 (N606, N602, N207, N1);
and AND2 (N607, N598, N178);
and AND2 (N608, N586, N340);
nor NOR3 (N609, N601, N464, N588);
nand NAND3 (N610, N609, N92, N45);
buf BUF1 (N611, N587);
or OR3 (N612, N596, N431, N271);
nor NOR2 (N613, N605, N435);
not NOT1 (N614, N606);
xor XOR2 (N615, N612, N334);
not NOT1 (N616, N580);
nand NAND2 (N617, N610, N149);
buf BUF1 (N618, N614);
and AND3 (N619, N608, N276, N398);
nor NOR3 (N620, N604, N455, N68);
buf BUF1 (N621, N615);
or OR2 (N622, N611, N50);
or OR4 (N623, N607, N432, N576, N139);
and AND3 (N624, N617, N198, N450);
xor XOR2 (N625, N619, N402);
nand NAND3 (N626, N618, N26, N494);
nor NOR2 (N627, N621, N227);
and AND3 (N628, N622, N623, N399);
nand NAND3 (N629, N622, N594, N510);
not NOT1 (N630, N626);
and AND4 (N631, N603, N41, N13, N289);
or OR4 (N632, N620, N591, N156, N370);
not NOT1 (N633, N625);
not NOT1 (N634, N630);
and AND4 (N635, N613, N451, N587, N44);
nand NAND4 (N636, N616, N16, N291, N57);
nand NAND2 (N637, N629, N65);
not NOT1 (N638, N624);
not NOT1 (N639, N631);
nand NAND2 (N640, N627, N159);
not NOT1 (N641, N636);
and AND2 (N642, N637, N288);
buf BUF1 (N643, N639);
buf BUF1 (N644, N635);
xor XOR2 (N645, N643, N34);
and AND2 (N646, N638, N302);
nand NAND2 (N647, N645, N404);
or OR2 (N648, N633, N433);
buf BUF1 (N649, N634);
nand NAND3 (N650, N632, N608, N534);
nand NAND4 (N651, N648, N96, N312, N179);
nand NAND4 (N652, N640, N349, N648, N583);
or OR3 (N653, N651, N150, N482);
nor NOR4 (N654, N646, N424, N143, N500);
not NOT1 (N655, N654);
or OR2 (N656, N642, N593);
not NOT1 (N657, N647);
or OR3 (N658, N649, N338, N634);
xor XOR2 (N659, N650, N330);
or OR3 (N660, N657, N645, N465);
not NOT1 (N661, N658);
or OR3 (N662, N644, N27, N653);
and AND2 (N663, N348, N219);
nand NAND4 (N664, N641, N118, N149, N407);
nor NOR3 (N665, N661, N92, N503);
nand NAND4 (N666, N662, N363, N57, N125);
and AND4 (N667, N660, N395, N67, N48);
not NOT1 (N668, N667);
not NOT1 (N669, N656);
nor NOR4 (N670, N664, N573, N579, N559);
buf BUF1 (N671, N655);
not NOT1 (N672, N666);
not NOT1 (N673, N663);
or OR3 (N674, N672, N51, N504);
not NOT1 (N675, N665);
not NOT1 (N676, N675);
and AND3 (N677, N659, N484, N565);
or OR3 (N678, N676, N165, N573);
nor NOR2 (N679, N669, N107);
not NOT1 (N680, N677);
xor XOR2 (N681, N652, N654);
not NOT1 (N682, N628);
buf BUF1 (N683, N682);
buf BUF1 (N684, N678);
nor NOR3 (N685, N684, N341, N579);
or OR2 (N686, N680, N92);
nand NAND3 (N687, N673, N527, N32);
xor XOR2 (N688, N687, N468);
and AND3 (N689, N679, N100, N442);
and AND2 (N690, N683, N149);
and AND2 (N691, N668, N405);
buf BUF1 (N692, N688);
nor NOR3 (N693, N689, N183, N662);
or OR2 (N694, N691, N454);
and AND2 (N695, N686, N80);
and AND3 (N696, N692, N179, N250);
nor NOR3 (N697, N690, N627, N493);
and AND3 (N698, N670, N591, N373);
nor NOR4 (N699, N696, N178, N178, N202);
or OR4 (N700, N685, N458, N139, N480);
and AND3 (N701, N697, N394, N503);
xor XOR2 (N702, N698, N41);
and AND2 (N703, N700, N449);
buf BUF1 (N704, N681);
buf BUF1 (N705, N671);
buf BUF1 (N706, N694);
nand NAND2 (N707, N704, N467);
nor NOR2 (N708, N695, N521);
nor NOR2 (N709, N707, N425);
not NOT1 (N710, N709);
nor NOR2 (N711, N701, N37);
not NOT1 (N712, N693);
nand NAND2 (N713, N699, N188);
xor XOR2 (N714, N703, N187);
nor NOR2 (N715, N706, N410);
xor XOR2 (N716, N705, N277);
not NOT1 (N717, N713);
or OR3 (N718, N716, N228, N137);
nand NAND4 (N719, N717, N519, N169, N1);
nand NAND2 (N720, N718, N46);
or OR3 (N721, N674, N203, N340);
buf BUF1 (N722, N712);
buf BUF1 (N723, N708);
nand NAND3 (N724, N722, N254, N527);
nand NAND4 (N725, N702, N253, N295, N660);
buf BUF1 (N726, N715);
xor XOR2 (N727, N719, N280);
nor NOR2 (N728, N721, N367);
nand NAND4 (N729, N726, N38, N147, N210);
nor NOR2 (N730, N729, N708);
buf BUF1 (N731, N724);
or OR3 (N732, N711, N413, N375);
and AND4 (N733, N731, N599, N281, N84);
nand NAND2 (N734, N727, N189);
buf BUF1 (N735, N710);
or OR3 (N736, N732, N271, N647);
not NOT1 (N737, N728);
or OR2 (N738, N725, N714);
or OR4 (N739, N99, N610, N524, N170);
not NOT1 (N740, N738);
nand NAND4 (N741, N730, N540, N645, N412);
and AND2 (N742, N734, N148);
and AND4 (N743, N720, N437, N486, N154);
nand NAND2 (N744, N737, N584);
and AND2 (N745, N723, N71);
buf BUF1 (N746, N745);
buf BUF1 (N747, N740);
xor XOR2 (N748, N746, N124);
not NOT1 (N749, N743);
nand NAND2 (N750, N736, N615);
nand NAND3 (N751, N742, N553, N98);
buf BUF1 (N752, N744);
buf BUF1 (N753, N747);
nor NOR2 (N754, N749, N96);
and AND3 (N755, N733, N699, N555);
xor XOR2 (N756, N752, N677);
buf BUF1 (N757, N750);
and AND3 (N758, N756, N75, N746);
buf BUF1 (N759, N735);
nand NAND3 (N760, N758, N444, N275);
xor XOR2 (N761, N739, N660);
buf BUF1 (N762, N751);
nor NOR2 (N763, N753, N677);
xor XOR2 (N764, N760, N645);
and AND2 (N765, N764, N402);
xor XOR2 (N766, N762, N432);
nand NAND2 (N767, N766, N209);
nor NOR3 (N768, N759, N700, N39);
buf BUF1 (N769, N757);
nand NAND3 (N770, N754, N591, N157);
xor XOR2 (N771, N748, N71);
buf BUF1 (N772, N768);
buf BUF1 (N773, N741);
nand NAND2 (N774, N767, N771);
xor XOR2 (N775, N632, N652);
xor XOR2 (N776, N772, N53);
nor NOR3 (N777, N775, N272, N634);
xor XOR2 (N778, N769, N195);
xor XOR2 (N779, N755, N661);
buf BUF1 (N780, N770);
buf BUF1 (N781, N776);
not NOT1 (N782, N780);
and AND3 (N783, N765, N93, N430);
nor NOR4 (N784, N779, N754, N639, N295);
not NOT1 (N785, N763);
or OR4 (N786, N783, N299, N466, N458);
buf BUF1 (N787, N781);
buf BUF1 (N788, N777);
nand NAND2 (N789, N785, N4);
and AND2 (N790, N774, N163);
not NOT1 (N791, N786);
not NOT1 (N792, N761);
xor XOR2 (N793, N792, N709);
nor NOR2 (N794, N791, N423);
nand NAND2 (N795, N778, N221);
not NOT1 (N796, N787);
not NOT1 (N797, N784);
nor NOR3 (N798, N794, N549, N402);
nor NOR2 (N799, N789, N164);
nor NOR3 (N800, N790, N248, N410);
nand NAND3 (N801, N788, N769, N272);
buf BUF1 (N802, N795);
buf BUF1 (N803, N799);
and AND3 (N804, N798, N723, N604);
and AND2 (N805, N773, N180);
not NOT1 (N806, N796);
or OR3 (N807, N806, N679, N50);
not NOT1 (N808, N800);
nor NOR3 (N809, N801, N786, N709);
and AND4 (N810, N803, N589, N681, N407);
and AND4 (N811, N804, N2, N641, N627);
nor NOR3 (N812, N793, N485, N528);
not NOT1 (N813, N782);
not NOT1 (N814, N805);
nor NOR4 (N815, N810, N134, N117, N489);
xor XOR2 (N816, N797, N296);
nand NAND4 (N817, N807, N449, N690, N765);
nor NOR3 (N818, N802, N724, N761);
or OR2 (N819, N816, N807);
xor XOR2 (N820, N814, N79);
xor XOR2 (N821, N817, N89);
not NOT1 (N822, N818);
or OR3 (N823, N811, N505, N690);
and AND3 (N824, N808, N168, N19);
buf BUF1 (N825, N824);
xor XOR2 (N826, N813, N440);
xor XOR2 (N827, N819, N793);
and AND4 (N828, N826, N631, N95, N503);
nor NOR4 (N829, N828, N396, N463, N704);
and AND2 (N830, N823, N197);
and AND3 (N831, N815, N553, N461);
not NOT1 (N832, N827);
nor NOR3 (N833, N825, N631, N651);
nor NOR3 (N834, N812, N203, N229);
or OR2 (N835, N820, N235);
and AND3 (N836, N832, N824, N616);
xor XOR2 (N837, N821, N549);
and AND3 (N838, N835, N616, N166);
xor XOR2 (N839, N834, N293);
and AND3 (N840, N809, N89, N698);
buf BUF1 (N841, N839);
nand NAND4 (N842, N836, N568, N84, N583);
nand NAND3 (N843, N831, N368, N161);
buf BUF1 (N844, N842);
and AND3 (N845, N844, N216, N630);
buf BUF1 (N846, N845);
nor NOR4 (N847, N830, N817, N545, N740);
not NOT1 (N848, N833);
or OR3 (N849, N848, N660, N269);
not NOT1 (N850, N838);
buf BUF1 (N851, N846);
and AND3 (N852, N840, N662, N497);
nor NOR2 (N853, N837, N468);
nor NOR3 (N854, N851, N541, N561);
nand NAND4 (N855, N854, N126, N668, N451);
xor XOR2 (N856, N850, N708);
xor XOR2 (N857, N852, N720);
buf BUF1 (N858, N822);
nand NAND2 (N859, N849, N766);
nand NAND4 (N860, N857, N65, N292, N516);
xor XOR2 (N861, N841, N370);
and AND2 (N862, N860, N640);
not NOT1 (N863, N847);
buf BUF1 (N864, N853);
xor XOR2 (N865, N862, N379);
nor NOR2 (N866, N864, N258);
not NOT1 (N867, N865);
buf BUF1 (N868, N859);
or OR2 (N869, N866, N478);
buf BUF1 (N870, N868);
nand NAND2 (N871, N858, N814);
or OR2 (N872, N855, N309);
and AND2 (N873, N863, N327);
nor NOR3 (N874, N873, N25, N648);
xor XOR2 (N875, N861, N681);
nand NAND4 (N876, N843, N210, N57, N128);
and AND2 (N877, N872, N679);
buf BUF1 (N878, N875);
xor XOR2 (N879, N871, N64);
and AND4 (N880, N829, N852, N389, N195);
nand NAND3 (N881, N869, N772, N343);
xor XOR2 (N882, N878, N805);
buf BUF1 (N883, N879);
not NOT1 (N884, N870);
or OR3 (N885, N882, N505, N434);
and AND4 (N886, N874, N135, N499, N690);
or OR3 (N887, N886, N663, N250);
nand NAND4 (N888, N881, N663, N336, N323);
and AND4 (N889, N884, N268, N709, N452);
nor NOR4 (N890, N887, N24, N236, N834);
and AND2 (N891, N877, N513);
and AND3 (N892, N891, N44, N58);
xor XOR2 (N893, N883, N177);
buf BUF1 (N894, N867);
not NOT1 (N895, N894);
buf BUF1 (N896, N895);
or OR3 (N897, N880, N218, N540);
nor NOR4 (N898, N856, N465, N152, N597);
buf BUF1 (N899, N896);
or OR2 (N900, N876, N866);
and AND4 (N901, N899, N30, N493, N877);
nor NOR4 (N902, N885, N169, N171, N519);
xor XOR2 (N903, N900, N385);
and AND4 (N904, N902, N29, N555, N735);
xor XOR2 (N905, N889, N866);
xor XOR2 (N906, N897, N375);
or OR2 (N907, N904, N129);
or OR4 (N908, N907, N261, N537, N586);
or OR4 (N909, N892, N859, N565, N115);
and AND2 (N910, N888, N354);
and AND2 (N911, N901, N889);
xor XOR2 (N912, N911, N16);
not NOT1 (N913, N908);
nor NOR2 (N914, N890, N581);
nor NOR3 (N915, N913, N711, N905);
and AND3 (N916, N368, N779, N751);
buf BUF1 (N917, N903);
not NOT1 (N918, N915);
and AND3 (N919, N918, N468, N142);
and AND3 (N920, N909, N520, N284);
buf BUF1 (N921, N917);
nand NAND3 (N922, N912, N763, N369);
not NOT1 (N923, N916);
xor XOR2 (N924, N920, N789);
or OR2 (N925, N923, N247);
buf BUF1 (N926, N921);
buf BUF1 (N927, N922);
nor NOR4 (N928, N927, N588, N590, N732);
xor XOR2 (N929, N928, N646);
or OR3 (N930, N926, N99, N733);
not NOT1 (N931, N930);
and AND3 (N932, N931, N728, N397);
or OR3 (N933, N932, N190, N574);
nand NAND4 (N934, N924, N46, N784, N768);
xor XOR2 (N935, N914, N476);
buf BUF1 (N936, N919);
or OR4 (N937, N936, N230, N921, N663);
buf BUF1 (N938, N935);
nand NAND3 (N939, N925, N13, N285);
and AND3 (N940, N898, N888, N612);
not NOT1 (N941, N939);
buf BUF1 (N942, N910);
and AND2 (N943, N934, N850);
buf BUF1 (N944, N933);
not NOT1 (N945, N893);
or OR3 (N946, N906, N16, N330);
or OR3 (N947, N938, N595, N221);
nor NOR3 (N948, N946, N122, N753);
or OR3 (N949, N944, N133, N537);
not NOT1 (N950, N941);
xor XOR2 (N951, N943, N493);
not NOT1 (N952, N929);
xor XOR2 (N953, N950, N93);
not NOT1 (N954, N953);
nor NOR3 (N955, N947, N582, N929);
and AND4 (N956, N942, N605, N560, N793);
nor NOR2 (N957, N955, N624);
or OR2 (N958, N949, N537);
xor XOR2 (N959, N958, N570);
or OR2 (N960, N951, N185);
or OR2 (N961, N956, N698);
or OR2 (N962, N937, N650);
nand NAND2 (N963, N940, N307);
xor XOR2 (N964, N952, N36);
buf BUF1 (N965, N948);
or OR2 (N966, N959, N3);
not NOT1 (N967, N965);
nor NOR4 (N968, N961, N607, N754, N79);
and AND3 (N969, N966, N173, N847);
nand NAND4 (N970, N954, N66, N442, N744);
and AND2 (N971, N970, N811);
nor NOR2 (N972, N969, N815);
nor NOR2 (N973, N945, N18);
or OR4 (N974, N960, N82, N150, N784);
and AND4 (N975, N968, N201, N613, N75);
nand NAND4 (N976, N975, N75, N147, N334);
or OR4 (N977, N971, N708, N877, N744);
or OR2 (N978, N963, N883);
buf BUF1 (N979, N973);
xor XOR2 (N980, N977, N45);
xor XOR2 (N981, N979, N325);
or OR3 (N982, N967, N664, N195);
not NOT1 (N983, N957);
xor XOR2 (N984, N981, N386);
buf BUF1 (N985, N972);
xor XOR2 (N986, N962, N108);
nor NOR2 (N987, N974, N913);
or OR3 (N988, N976, N572, N211);
or OR3 (N989, N985, N401, N963);
not NOT1 (N990, N988);
nor NOR4 (N991, N987, N22, N150, N645);
nor NOR2 (N992, N986, N549);
and AND3 (N993, N984, N595, N870);
and AND4 (N994, N989, N332, N391, N745);
not NOT1 (N995, N991);
nor NOR3 (N996, N982, N539, N518);
buf BUF1 (N997, N992);
or OR2 (N998, N996, N791);
not NOT1 (N999, N997);
and AND3 (N1000, N978, N800, N295);
and AND3 (N1001, N964, N437, N790);
buf BUF1 (N1002, N1001);
not NOT1 (N1003, N983);
buf BUF1 (N1004, N995);
xor XOR2 (N1005, N999, N533);
not NOT1 (N1006, N1002);
xor XOR2 (N1007, N990, N373);
xor XOR2 (N1008, N1000, N263);
buf BUF1 (N1009, N994);
and AND2 (N1010, N1007, N781);
or OR3 (N1011, N1003, N26, N145);
nand NAND3 (N1012, N993, N998, N370);
nand NAND2 (N1013, N930, N482);
xor XOR2 (N1014, N1012, N57);
buf BUF1 (N1015, N1009);
and AND4 (N1016, N1005, N172, N431, N841);
nor NOR2 (N1017, N1014, N742);
or OR2 (N1018, N980, N140);
not NOT1 (N1019, N1017);
nor NOR3 (N1020, N1015, N112, N815);
nor NOR3 (N1021, N1018, N16, N665);
nand NAND2 (N1022, N1006, N315);
buf BUF1 (N1023, N1013);
nand NAND4 (N1024, N1004, N146, N821, N109);
nand NAND3 (N1025, N1019, N920, N605);
nor NOR4 (N1026, N1011, N4, N492, N970);
xor XOR2 (N1027, N1024, N31);
buf BUF1 (N1028, N1016);
xor XOR2 (N1029, N1020, N96);
buf BUF1 (N1030, N1028);
nand NAND3 (N1031, N1029, N845, N766);
buf BUF1 (N1032, N1022);
or OR2 (N1033, N1031, N629);
or OR2 (N1034, N1021, N692);
nor NOR2 (N1035, N1030, N790);
not NOT1 (N1036, N1033);
nand NAND3 (N1037, N1023, N225, N103);
nor NOR2 (N1038, N1032, N530);
or OR4 (N1039, N1008, N234, N281, N80);
nor NOR4 (N1040, N1034, N791, N260, N465);
xor XOR2 (N1041, N1036, N113);
buf BUF1 (N1042, N1039);
xor XOR2 (N1043, N1035, N321);
or OR3 (N1044, N1041, N507, N1021);
not NOT1 (N1045, N1038);
nor NOR4 (N1046, N1042, N140, N1043, N164);
or OR3 (N1047, N508, N677, N758);
xor XOR2 (N1048, N1044, N96);
and AND4 (N1049, N1048, N240, N183, N169);
or OR4 (N1050, N1010, N643, N1025, N419);
nand NAND3 (N1051, N203, N710, N278);
nand NAND4 (N1052, N1040, N991, N39, N213);
and AND2 (N1053, N1049, N301);
buf BUF1 (N1054, N1053);
xor XOR2 (N1055, N1052, N476);
or OR3 (N1056, N1046, N485, N818);
not NOT1 (N1057, N1055);
and AND3 (N1058, N1057, N572, N693);
xor XOR2 (N1059, N1027, N423);
not NOT1 (N1060, N1045);
and AND3 (N1061, N1060, N816, N737);
buf BUF1 (N1062, N1050);
not NOT1 (N1063, N1058);
and AND3 (N1064, N1026, N1001, N496);
not NOT1 (N1065, N1062);
nor NOR3 (N1066, N1037, N353, N556);
buf BUF1 (N1067, N1051);
nand NAND3 (N1068, N1054, N964, N995);
and AND4 (N1069, N1068, N88, N301, N684);
not NOT1 (N1070, N1061);
nor NOR4 (N1071, N1059, N417, N740, N742);
not NOT1 (N1072, N1063);
nor NOR3 (N1073, N1071, N753, N458);
nand NAND4 (N1074, N1067, N284, N919, N376);
not NOT1 (N1075, N1073);
nand NAND2 (N1076, N1056, N204);
xor XOR2 (N1077, N1070, N483);
or OR2 (N1078, N1065, N1072);
buf BUF1 (N1079, N638);
nor NOR2 (N1080, N1074, N128);
or OR4 (N1081, N1075, N97, N570, N22);
xor XOR2 (N1082, N1076, N690);
or OR3 (N1083, N1080, N14, N1012);
buf BUF1 (N1084, N1077);
or OR3 (N1085, N1078, N1067, N860);
nor NOR3 (N1086, N1047, N1006, N447);
xor XOR2 (N1087, N1082, N802);
and AND3 (N1088, N1087, N322, N1081);
buf BUF1 (N1089, N158);
nand NAND4 (N1090, N1066, N23, N281, N456);
nand NAND4 (N1091, N1090, N172, N839, N126);
and AND4 (N1092, N1088, N382, N602, N662);
not NOT1 (N1093, N1069);
nand NAND4 (N1094, N1092, N1039, N1019, N957);
or OR4 (N1095, N1086, N912, N685, N101);
and AND4 (N1096, N1089, N518, N974, N130);
buf BUF1 (N1097, N1085);
xor XOR2 (N1098, N1091, N681);
xor XOR2 (N1099, N1083, N894);
nand NAND3 (N1100, N1093, N414, N814);
not NOT1 (N1101, N1084);
nor NOR2 (N1102, N1097, N525);
xor XOR2 (N1103, N1094, N46);
nor NOR2 (N1104, N1095, N559);
not NOT1 (N1105, N1101);
buf BUF1 (N1106, N1099);
and AND3 (N1107, N1104, N116, N821);
xor XOR2 (N1108, N1079, N643);
nor NOR4 (N1109, N1100, N935, N137, N498);
nor NOR2 (N1110, N1106, N870);
buf BUF1 (N1111, N1107);
buf BUF1 (N1112, N1105);
and AND4 (N1113, N1109, N217, N131, N230);
buf BUF1 (N1114, N1102);
not NOT1 (N1115, N1110);
nor NOR2 (N1116, N1064, N1073);
not NOT1 (N1117, N1111);
nand NAND3 (N1118, N1112, N623, N417);
xor XOR2 (N1119, N1115, N430);
buf BUF1 (N1120, N1113);
or OR4 (N1121, N1098, N323, N153, N503);
or OR2 (N1122, N1114, N703);
and AND3 (N1123, N1103, N836, N745);
and AND3 (N1124, N1116, N232, N896);
and AND3 (N1125, N1124, N281, N782);
nand NAND4 (N1126, N1119, N48, N823, N357);
xor XOR2 (N1127, N1108, N1053);
buf BUF1 (N1128, N1126);
not NOT1 (N1129, N1121);
not NOT1 (N1130, N1096);
buf BUF1 (N1131, N1125);
nand NAND4 (N1132, N1127, N134, N979, N347);
buf BUF1 (N1133, N1130);
xor XOR2 (N1134, N1123, N48);
nor NOR2 (N1135, N1118, N608);
xor XOR2 (N1136, N1122, N243);
nor NOR2 (N1137, N1136, N825);
and AND3 (N1138, N1134, N979, N433);
xor XOR2 (N1139, N1117, N250);
nor NOR4 (N1140, N1120, N402, N793, N629);
and AND2 (N1141, N1128, N634);
and AND2 (N1142, N1129, N684);
nand NAND4 (N1143, N1139, N559, N384, N705);
and AND3 (N1144, N1141, N453, N726);
and AND3 (N1145, N1144, N1, N805);
and AND2 (N1146, N1132, N608);
and AND2 (N1147, N1145, N32);
xor XOR2 (N1148, N1142, N556);
nor NOR2 (N1149, N1140, N296);
and AND3 (N1150, N1131, N1066, N1002);
not NOT1 (N1151, N1148);
nor NOR3 (N1152, N1147, N403, N449);
xor XOR2 (N1153, N1151, N135);
nand NAND2 (N1154, N1143, N834);
not NOT1 (N1155, N1149);
or OR2 (N1156, N1133, N461);
xor XOR2 (N1157, N1154, N457);
nor NOR4 (N1158, N1152, N309, N25, N804);
and AND2 (N1159, N1153, N891);
or OR3 (N1160, N1135, N826, N35);
and AND2 (N1161, N1137, N940);
or OR4 (N1162, N1146, N248, N256, N263);
nor NOR2 (N1163, N1156, N722);
xor XOR2 (N1164, N1159, N259);
not NOT1 (N1165, N1160);
nor NOR4 (N1166, N1161, N219, N348, N1073);
and AND2 (N1167, N1162, N868);
not NOT1 (N1168, N1166);
buf BUF1 (N1169, N1164);
xor XOR2 (N1170, N1155, N152);
xor XOR2 (N1171, N1163, N666);
nand NAND3 (N1172, N1167, N661, N659);
buf BUF1 (N1173, N1169);
not NOT1 (N1174, N1171);
and AND3 (N1175, N1170, N243, N404);
or OR3 (N1176, N1174, N413, N851);
nor NOR3 (N1177, N1150, N412, N322);
and AND3 (N1178, N1157, N563, N785);
nor NOR4 (N1179, N1178, N943, N122, N985);
and AND3 (N1180, N1158, N620, N471);
buf BUF1 (N1181, N1173);
nor NOR2 (N1182, N1180, N1061);
not NOT1 (N1183, N1179);
nor NOR3 (N1184, N1176, N700, N1141);
and AND4 (N1185, N1183, N1017, N547, N951);
nand NAND2 (N1186, N1181, N821);
not NOT1 (N1187, N1172);
nand NAND4 (N1188, N1168, N1047, N429, N345);
xor XOR2 (N1189, N1182, N790);
buf BUF1 (N1190, N1185);
nand NAND4 (N1191, N1188, N808, N570, N471);
and AND4 (N1192, N1191, N768, N272, N741);
nor NOR2 (N1193, N1184, N173);
buf BUF1 (N1194, N1177);
buf BUF1 (N1195, N1190);
xor XOR2 (N1196, N1195, N578);
buf BUF1 (N1197, N1186);
and AND4 (N1198, N1192, N752, N289, N735);
buf BUF1 (N1199, N1138);
nor NOR3 (N1200, N1196, N655, N111);
not NOT1 (N1201, N1200);
nand NAND2 (N1202, N1165, N301);
nor NOR2 (N1203, N1189, N794);
or OR4 (N1204, N1187, N467, N51, N788);
nor NOR3 (N1205, N1199, N1011, N763);
and AND4 (N1206, N1204, N1065, N44, N1031);
not NOT1 (N1207, N1202);
buf BUF1 (N1208, N1207);
and AND2 (N1209, N1194, N908);
and AND2 (N1210, N1193, N1135);
nand NAND3 (N1211, N1203, N625, N639);
nand NAND3 (N1212, N1175, N865, N696);
or OR3 (N1213, N1201, N67, N491);
buf BUF1 (N1214, N1209);
xor XOR2 (N1215, N1205, N677);
and AND4 (N1216, N1215, N548, N635, N629);
not NOT1 (N1217, N1212);
or OR4 (N1218, N1197, N619, N1065, N110);
not NOT1 (N1219, N1214);
nor NOR3 (N1220, N1218, N1175, N258);
xor XOR2 (N1221, N1213, N503);
not NOT1 (N1222, N1210);
or OR3 (N1223, N1221, N377, N842);
nand NAND2 (N1224, N1222, N463);
xor XOR2 (N1225, N1223, N1063);
buf BUF1 (N1226, N1220);
nand NAND3 (N1227, N1198, N616, N453);
or OR3 (N1228, N1206, N772, N231);
not NOT1 (N1229, N1219);
nor NOR3 (N1230, N1211, N1205, N517);
nand NAND4 (N1231, N1229, N567, N1076, N664);
and AND4 (N1232, N1231, N65, N1050, N529);
nor NOR4 (N1233, N1225, N110, N377, N324);
nand NAND2 (N1234, N1217, N1191);
not NOT1 (N1235, N1227);
nand NAND4 (N1236, N1232, N635, N799, N118);
or OR4 (N1237, N1216, N1030, N159, N685);
buf BUF1 (N1238, N1235);
nand NAND3 (N1239, N1236, N842, N569);
buf BUF1 (N1240, N1228);
xor XOR2 (N1241, N1226, N853);
and AND3 (N1242, N1234, N564, N343);
nor NOR2 (N1243, N1233, N257);
or OR4 (N1244, N1240, N159, N134, N379);
not NOT1 (N1245, N1208);
and AND4 (N1246, N1243, N239, N229, N650);
nand NAND3 (N1247, N1242, N1205, N99);
buf BUF1 (N1248, N1238);
buf BUF1 (N1249, N1241);
buf BUF1 (N1250, N1246);
or OR3 (N1251, N1249, N290, N448);
not NOT1 (N1252, N1247);
nand NAND2 (N1253, N1230, N1222);
not NOT1 (N1254, N1224);
and AND4 (N1255, N1254, N1005, N129, N173);
xor XOR2 (N1256, N1255, N193);
and AND3 (N1257, N1248, N302, N1112);
and AND4 (N1258, N1250, N620, N1102, N1136);
and AND2 (N1259, N1239, N436);
buf BUF1 (N1260, N1245);
nor NOR3 (N1261, N1253, N1128, N631);
xor XOR2 (N1262, N1257, N689);
and AND4 (N1263, N1261, N501, N457, N959);
xor XOR2 (N1264, N1252, N499);
and AND3 (N1265, N1263, N929, N94);
nor NOR2 (N1266, N1260, N957);
buf BUF1 (N1267, N1264);
and AND4 (N1268, N1259, N674, N1009, N19);
nand NAND3 (N1269, N1268, N29, N910);
buf BUF1 (N1270, N1237);
and AND4 (N1271, N1267, N548, N723, N898);
xor XOR2 (N1272, N1266, N24);
nand NAND2 (N1273, N1251, N219);
buf BUF1 (N1274, N1265);
nand NAND3 (N1275, N1258, N474, N680);
nor NOR4 (N1276, N1270, N401, N122, N1233);
not NOT1 (N1277, N1244);
or OR3 (N1278, N1275, N710, N464);
nor NOR3 (N1279, N1271, N687, N1210);
xor XOR2 (N1280, N1269, N537);
and AND3 (N1281, N1276, N372, N281);
nand NAND4 (N1282, N1262, N491, N1087, N476);
and AND4 (N1283, N1256, N308, N492, N963);
not NOT1 (N1284, N1272);
xor XOR2 (N1285, N1283, N1250);
or OR4 (N1286, N1284, N1040, N874, N83);
not NOT1 (N1287, N1273);
xor XOR2 (N1288, N1286, N874);
xor XOR2 (N1289, N1274, N285);
and AND2 (N1290, N1287, N208);
nand NAND4 (N1291, N1290, N466, N39, N1279);
not NOT1 (N1292, N1085);
not NOT1 (N1293, N1280);
xor XOR2 (N1294, N1291, N887);
not NOT1 (N1295, N1293);
nor NOR2 (N1296, N1278, N39);
or OR2 (N1297, N1285, N364);
buf BUF1 (N1298, N1292);
and AND4 (N1299, N1295, N1288, N910, N49);
buf BUF1 (N1300, N435);
and AND3 (N1301, N1297, N919, N385);
nand NAND3 (N1302, N1282, N208, N195);
buf BUF1 (N1303, N1301);
nand NAND4 (N1304, N1289, N612, N515, N959);
not NOT1 (N1305, N1302);
and AND4 (N1306, N1300, N71, N470, N1240);
buf BUF1 (N1307, N1303);
xor XOR2 (N1308, N1281, N612);
nor NOR3 (N1309, N1277, N1147, N47);
nand NAND4 (N1310, N1296, N81, N222, N1267);
and AND2 (N1311, N1298, N1152);
nand NAND3 (N1312, N1311, N873, N303);
nor NOR4 (N1313, N1306, N418, N466, N835);
xor XOR2 (N1314, N1299, N225);
buf BUF1 (N1315, N1305);
and AND4 (N1316, N1310, N1011, N836, N629);
nor NOR3 (N1317, N1316, N741, N1131);
not NOT1 (N1318, N1304);
nand NAND2 (N1319, N1315, N189);
nor NOR4 (N1320, N1318, N688, N150, N791);
buf BUF1 (N1321, N1309);
or OR4 (N1322, N1314, N1311, N821, N469);
buf BUF1 (N1323, N1320);
or OR3 (N1324, N1319, N32, N404);
nor NOR4 (N1325, N1294, N1115, N189, N598);
and AND3 (N1326, N1308, N228, N867);
nand NAND2 (N1327, N1313, N559);
or OR2 (N1328, N1327, N957);
buf BUF1 (N1329, N1322);
nor NOR4 (N1330, N1326, N595, N171, N718);
nand NAND3 (N1331, N1330, N62, N1037);
nor NOR3 (N1332, N1325, N989, N48);
nand NAND4 (N1333, N1329, N1208, N585, N1069);
nand NAND4 (N1334, N1317, N657, N568, N1140);
and AND4 (N1335, N1307, N923, N621, N324);
or OR4 (N1336, N1333, N186, N19, N939);
or OR4 (N1337, N1321, N335, N1289, N1275);
and AND2 (N1338, N1323, N1154);
nand NAND3 (N1339, N1312, N573, N987);
and AND2 (N1340, N1336, N703);
nand NAND2 (N1341, N1324, N1265);
and AND3 (N1342, N1335, N357, N1091);
xor XOR2 (N1343, N1339, N341);
and AND2 (N1344, N1337, N387);
or OR4 (N1345, N1344, N196, N298, N909);
nor NOR4 (N1346, N1342, N16, N783, N572);
and AND3 (N1347, N1338, N373, N27);
xor XOR2 (N1348, N1328, N778);
nor NOR3 (N1349, N1345, N1118, N61);
nand NAND2 (N1350, N1343, N852);
not NOT1 (N1351, N1340);
and AND3 (N1352, N1348, N560, N1101);
not NOT1 (N1353, N1334);
nand NAND3 (N1354, N1331, N493, N549);
nand NAND3 (N1355, N1352, N67, N11);
nor NOR3 (N1356, N1332, N381, N591);
not NOT1 (N1357, N1353);
not NOT1 (N1358, N1354);
xor XOR2 (N1359, N1351, N925);
not NOT1 (N1360, N1358);
buf BUF1 (N1361, N1349);
nand NAND3 (N1362, N1347, N965, N1161);
and AND3 (N1363, N1341, N1078, N885);
or OR4 (N1364, N1360, N140, N837, N429);
or OR2 (N1365, N1361, N639);
xor XOR2 (N1366, N1362, N1053);
or OR3 (N1367, N1346, N1366, N364);
or OR2 (N1368, N79, N236);
nand NAND4 (N1369, N1350, N925, N1336, N11);
not NOT1 (N1370, N1357);
nor NOR2 (N1371, N1364, N1221);
and AND4 (N1372, N1355, N414, N193, N1254);
nand NAND2 (N1373, N1370, N963);
and AND2 (N1374, N1363, N685);
nor NOR4 (N1375, N1365, N567, N79, N1311);
xor XOR2 (N1376, N1372, N142);
nor NOR2 (N1377, N1371, N64);
nor NOR4 (N1378, N1369, N1145, N883, N1228);
nand NAND3 (N1379, N1378, N9, N1221);
buf BUF1 (N1380, N1377);
or OR2 (N1381, N1375, N208);
xor XOR2 (N1382, N1379, N898);
and AND4 (N1383, N1359, N1129, N872, N1310);
xor XOR2 (N1384, N1383, N269);
nor NOR2 (N1385, N1356, N839);
not NOT1 (N1386, N1382);
xor XOR2 (N1387, N1385, N527);
or OR2 (N1388, N1386, N1248);
nor NOR2 (N1389, N1381, N608);
or OR3 (N1390, N1387, N553, N173);
and AND4 (N1391, N1388, N576, N1173, N718);
and AND4 (N1392, N1374, N175, N798, N499);
or OR4 (N1393, N1368, N93, N605, N1374);
or OR3 (N1394, N1380, N1047, N1142);
not NOT1 (N1395, N1393);
nor NOR2 (N1396, N1367, N1327);
not NOT1 (N1397, N1392);
buf BUF1 (N1398, N1390);
nand NAND3 (N1399, N1384, N330, N46);
not NOT1 (N1400, N1395);
and AND3 (N1401, N1391, N1231, N1228);
or OR4 (N1402, N1376, N468, N70, N124);
buf BUF1 (N1403, N1402);
not NOT1 (N1404, N1403);
nor NOR4 (N1405, N1394, N1363, N1075, N643);
xor XOR2 (N1406, N1389, N842);
buf BUF1 (N1407, N1396);
not NOT1 (N1408, N1401);
nand NAND3 (N1409, N1397, N887, N921);
buf BUF1 (N1410, N1400);
and AND2 (N1411, N1373, N965);
or OR4 (N1412, N1398, N843, N1207, N253);
not NOT1 (N1413, N1404);
nand NAND3 (N1414, N1406, N40, N92);
buf BUF1 (N1415, N1408);
nor NOR2 (N1416, N1409, N652);
or OR4 (N1417, N1415, N830, N975, N922);
xor XOR2 (N1418, N1405, N635);
or OR4 (N1419, N1418, N391, N1009, N1330);
or OR3 (N1420, N1417, N643, N951);
or OR4 (N1421, N1411, N81, N562, N1161);
and AND2 (N1422, N1420, N420);
or OR2 (N1423, N1407, N217);
or OR3 (N1424, N1399, N70, N1060);
buf BUF1 (N1425, N1419);
nor NOR4 (N1426, N1422, N1171, N1166, N224);
xor XOR2 (N1427, N1413, N600);
nand NAND4 (N1428, N1424, N1232, N976, N547);
and AND2 (N1429, N1428, N684);
nor NOR4 (N1430, N1423, N411, N1119, N47);
and AND3 (N1431, N1410, N7, N797);
nand NAND4 (N1432, N1431, N901, N592, N819);
nand NAND4 (N1433, N1427, N723, N920, N799);
nor NOR2 (N1434, N1433, N1392);
and AND3 (N1435, N1434, N1069, N497);
nand NAND4 (N1436, N1429, N276, N698, N1064);
not NOT1 (N1437, N1421);
or OR3 (N1438, N1416, N4, N583);
xor XOR2 (N1439, N1430, N549);
nand NAND2 (N1440, N1435, N779);
and AND3 (N1441, N1432, N687, N332);
or OR3 (N1442, N1441, N216, N187);
not NOT1 (N1443, N1442);
or OR3 (N1444, N1412, N61, N327);
xor XOR2 (N1445, N1425, N917);
buf BUF1 (N1446, N1445);
buf BUF1 (N1447, N1446);
nand NAND3 (N1448, N1437, N1240, N197);
nor NOR2 (N1449, N1440, N715);
or OR2 (N1450, N1448, N794);
not NOT1 (N1451, N1436);
buf BUF1 (N1452, N1450);
and AND3 (N1453, N1426, N499, N750);
nor NOR2 (N1454, N1444, N712);
nor NOR3 (N1455, N1449, N152, N1312);
and AND2 (N1456, N1443, N8);
nor NOR4 (N1457, N1451, N212, N122, N907);
nor NOR3 (N1458, N1457, N1007, N839);
nor NOR3 (N1459, N1447, N1306, N1404);
not NOT1 (N1460, N1455);
nand NAND2 (N1461, N1454, N214);
nor NOR3 (N1462, N1458, N722, N1015);
xor XOR2 (N1463, N1453, N1078);
and AND3 (N1464, N1463, N174, N1116);
nor NOR4 (N1465, N1462, N757, N655, N1106);
nor NOR4 (N1466, N1439, N1045, N1332, N815);
xor XOR2 (N1467, N1456, N844);
nand NAND3 (N1468, N1460, N535, N723);
not NOT1 (N1469, N1464);
nor NOR4 (N1470, N1465, N474, N1344, N784);
buf BUF1 (N1471, N1466);
buf BUF1 (N1472, N1459);
nand NAND4 (N1473, N1472, N774, N1029, N1464);
and AND3 (N1474, N1414, N11, N1464);
buf BUF1 (N1475, N1469);
not NOT1 (N1476, N1467);
not NOT1 (N1477, N1474);
and AND4 (N1478, N1468, N411, N525, N997);
nand NAND2 (N1479, N1461, N966);
nor NOR2 (N1480, N1452, N444);
not NOT1 (N1481, N1438);
buf BUF1 (N1482, N1470);
buf BUF1 (N1483, N1480);
nand NAND3 (N1484, N1476, N1107, N570);
nor NOR2 (N1485, N1475, N226);
xor XOR2 (N1486, N1471, N528);
xor XOR2 (N1487, N1484, N796);
nor NOR2 (N1488, N1485, N195);
not NOT1 (N1489, N1477);
not NOT1 (N1490, N1487);
xor XOR2 (N1491, N1483, N1127);
nor NOR4 (N1492, N1488, N280, N483, N969);
buf BUF1 (N1493, N1482);
buf BUF1 (N1494, N1493);
nor NOR3 (N1495, N1486, N378, N958);
xor XOR2 (N1496, N1491, N137);
buf BUF1 (N1497, N1492);
or OR4 (N1498, N1494, N1107, N1432, N848);
or OR2 (N1499, N1495, N29);
or OR2 (N1500, N1473, N663);
not NOT1 (N1501, N1490);
and AND3 (N1502, N1498, N716, N1433);
nor NOR2 (N1503, N1499, N209);
nand NAND3 (N1504, N1502, N1384, N235);
or OR3 (N1505, N1496, N945, N678);
and AND4 (N1506, N1501, N1344, N646, N391);
xor XOR2 (N1507, N1478, N1040);
nor NOR3 (N1508, N1506, N1115, N1381);
not NOT1 (N1509, N1505);
and AND2 (N1510, N1508, N979);
buf BUF1 (N1511, N1479);
nor NOR2 (N1512, N1497, N1203);
xor XOR2 (N1513, N1489, N217);
nand NAND3 (N1514, N1504, N549, N200);
nor NOR2 (N1515, N1513, N1439);
not NOT1 (N1516, N1500);
not NOT1 (N1517, N1515);
or OR3 (N1518, N1511, N905, N1131);
buf BUF1 (N1519, N1514);
xor XOR2 (N1520, N1510, N1450);
or OR4 (N1521, N1517, N556, N1435, N732);
and AND3 (N1522, N1512, N905, N1197);
nand NAND2 (N1523, N1481, N131);
and AND3 (N1524, N1521, N214, N854);
and AND3 (N1525, N1524, N249, N1186);
nor NOR3 (N1526, N1507, N693, N1318);
not NOT1 (N1527, N1518);
nor NOR3 (N1528, N1519, N362, N1364);
xor XOR2 (N1529, N1516, N84);
nor NOR2 (N1530, N1526, N961);
or OR2 (N1531, N1527, N652);
and AND2 (N1532, N1503, N1027);
xor XOR2 (N1533, N1528, N150);
not NOT1 (N1534, N1525);
and AND4 (N1535, N1520, N1328, N530, N477);
nor NOR2 (N1536, N1532, N20);
and AND3 (N1537, N1522, N212, N224);
nand NAND4 (N1538, N1531, N429, N650, N488);
buf BUF1 (N1539, N1533);
buf BUF1 (N1540, N1535);
not NOT1 (N1541, N1537);
or OR3 (N1542, N1536, N764, N559);
not NOT1 (N1543, N1529);
nand NAND3 (N1544, N1530, N797, N1171);
and AND4 (N1545, N1541, N1006, N255, N611);
nor NOR3 (N1546, N1534, N633, N1064);
nand NAND3 (N1547, N1543, N1526, N1452);
buf BUF1 (N1548, N1547);
and AND4 (N1549, N1542, N862, N1275, N572);
and AND4 (N1550, N1509, N570, N728, N1406);
or OR2 (N1551, N1549, N665);
xor XOR2 (N1552, N1545, N673);
buf BUF1 (N1553, N1548);
nor NOR4 (N1554, N1550, N1477, N1486, N305);
buf BUF1 (N1555, N1540);
not NOT1 (N1556, N1539);
buf BUF1 (N1557, N1551);
not NOT1 (N1558, N1546);
nand NAND3 (N1559, N1553, N1476, N1124);
and AND4 (N1560, N1556, N407, N1542, N238);
not NOT1 (N1561, N1559);
and AND3 (N1562, N1552, N893, N454);
xor XOR2 (N1563, N1544, N583);
buf BUF1 (N1564, N1560);
xor XOR2 (N1565, N1561, N1110);
or OR4 (N1566, N1563, N629, N852, N1329);
nor NOR4 (N1567, N1562, N975, N1015, N1376);
buf BUF1 (N1568, N1554);
nor NOR4 (N1569, N1557, N959, N909, N634);
nand NAND4 (N1570, N1569, N414, N352, N1181);
buf BUF1 (N1571, N1565);
not NOT1 (N1572, N1564);
not NOT1 (N1573, N1567);
buf BUF1 (N1574, N1573);
buf BUF1 (N1575, N1523);
nor NOR3 (N1576, N1538, N57, N599);
or OR4 (N1577, N1570, N364, N1484, N1493);
and AND4 (N1578, N1566, N755, N447, N424);
or OR3 (N1579, N1578, N1073, N1075);
and AND4 (N1580, N1576, N1019, N1337, N196);
not NOT1 (N1581, N1579);
nor NOR2 (N1582, N1555, N682);
nor NOR4 (N1583, N1571, N124, N1446, N636);
and AND3 (N1584, N1575, N1504, N258);
and AND2 (N1585, N1577, N1378);
buf BUF1 (N1586, N1582);
and AND3 (N1587, N1558, N748, N407);
or OR3 (N1588, N1587, N1313, N703);
xor XOR2 (N1589, N1572, N436);
or OR2 (N1590, N1586, N1041);
or OR2 (N1591, N1580, N1271);
nor NOR3 (N1592, N1591, N727, N1522);
or OR3 (N1593, N1592, N1274, N1013);
nor NOR2 (N1594, N1583, N568);
or OR3 (N1595, N1593, N455, N658);
nand NAND3 (N1596, N1588, N588, N762);
not NOT1 (N1597, N1585);
buf BUF1 (N1598, N1574);
nor NOR3 (N1599, N1581, N1191, N669);
or OR2 (N1600, N1568, N849);
buf BUF1 (N1601, N1598);
nand NAND3 (N1602, N1584, N428, N211);
and AND4 (N1603, N1597, N539, N53, N950);
and AND2 (N1604, N1599, N842);
nor NOR4 (N1605, N1602, N1344, N519, N799);
and AND2 (N1606, N1601, N366);
nor NOR4 (N1607, N1600, N57, N1095, N812);
buf BUF1 (N1608, N1589);
or OR4 (N1609, N1603, N1075, N779, N1544);
xor XOR2 (N1610, N1594, N642);
or OR4 (N1611, N1605, N485, N1218, N600);
nand NAND2 (N1612, N1610, N1123);
nor NOR2 (N1613, N1595, N1571);
buf BUF1 (N1614, N1590);
or OR3 (N1615, N1613, N1213, N60);
and AND4 (N1616, N1596, N617, N425, N516);
nand NAND4 (N1617, N1615, N1412, N1355, N513);
nand NAND2 (N1618, N1616, N327);
nor NOR2 (N1619, N1612, N440);
and AND3 (N1620, N1614, N707, N1228);
not NOT1 (N1621, N1620);
buf BUF1 (N1622, N1606);
nand NAND2 (N1623, N1618, N1294);
nand NAND3 (N1624, N1621, N1616, N1278);
buf BUF1 (N1625, N1622);
nand NAND4 (N1626, N1624, N111, N1462, N174);
nand NAND3 (N1627, N1609, N1339, N75);
xor XOR2 (N1628, N1607, N1282);
buf BUF1 (N1629, N1604);
and AND4 (N1630, N1629, N1407, N43, N896);
nand NAND3 (N1631, N1608, N1269, N1128);
and AND2 (N1632, N1623, N218);
nor NOR4 (N1633, N1625, N1255, N522, N1495);
nor NOR4 (N1634, N1627, N1200, N1188, N1358);
nand NAND4 (N1635, N1630, N1254, N1325, N845);
nand NAND4 (N1636, N1611, N1322, N796, N1075);
buf BUF1 (N1637, N1617);
nor NOR3 (N1638, N1637, N256, N483);
and AND4 (N1639, N1631, N915, N492, N1049);
buf BUF1 (N1640, N1636);
nand NAND4 (N1641, N1626, N1547, N1272, N1382);
nor NOR4 (N1642, N1638, N1580, N809, N1235);
nand NAND4 (N1643, N1639, N1249, N417, N1383);
xor XOR2 (N1644, N1640, N527);
or OR2 (N1645, N1642, N288);
buf BUF1 (N1646, N1644);
or OR3 (N1647, N1645, N1556, N1154);
not NOT1 (N1648, N1643);
nor NOR4 (N1649, N1647, N1392, N625, N613);
xor XOR2 (N1650, N1648, N1463);
nor NOR3 (N1651, N1632, N1574, N1437);
not NOT1 (N1652, N1650);
xor XOR2 (N1653, N1646, N919);
xor XOR2 (N1654, N1635, N1628);
and AND4 (N1655, N1255, N1, N613, N606);
buf BUF1 (N1656, N1634);
nor NOR3 (N1657, N1655, N142, N1304);
xor XOR2 (N1658, N1657, N1300);
nor NOR2 (N1659, N1649, N642);
nand NAND2 (N1660, N1619, N1324);
buf BUF1 (N1661, N1659);
nand NAND3 (N1662, N1641, N891, N1089);
and AND2 (N1663, N1653, N1385);
and AND4 (N1664, N1663, N253, N645, N47);
and AND3 (N1665, N1656, N534, N687);
or OR4 (N1666, N1662, N737, N604, N595);
xor XOR2 (N1667, N1665, N156);
nor NOR4 (N1668, N1667, N1423, N344, N938);
not NOT1 (N1669, N1633);
and AND4 (N1670, N1652, N422, N1298, N299);
buf BUF1 (N1671, N1669);
xor XOR2 (N1672, N1670, N1259);
buf BUF1 (N1673, N1654);
buf BUF1 (N1674, N1660);
not NOT1 (N1675, N1672);
nand NAND4 (N1676, N1674, N1480, N417, N1453);
xor XOR2 (N1677, N1671, N1647);
nor NOR2 (N1678, N1661, N1550);
xor XOR2 (N1679, N1666, N1416);
nor NOR3 (N1680, N1664, N326, N178);
nor NOR3 (N1681, N1678, N586, N241);
nand NAND2 (N1682, N1679, N301);
not NOT1 (N1683, N1651);
buf BUF1 (N1684, N1682);
nor NOR4 (N1685, N1676, N1507, N615, N785);
nor NOR4 (N1686, N1673, N1224, N470, N107);
and AND2 (N1687, N1685, N1682);
or OR4 (N1688, N1687, N350, N845, N949);
nand NAND2 (N1689, N1658, N826);
xor XOR2 (N1690, N1689, N1515);
nor NOR2 (N1691, N1690, N581);
not NOT1 (N1692, N1686);
or OR3 (N1693, N1675, N466, N624);
and AND3 (N1694, N1692, N914, N1338);
xor XOR2 (N1695, N1668, N990);
not NOT1 (N1696, N1694);
or OR4 (N1697, N1681, N1233, N1488, N596);
not NOT1 (N1698, N1697);
or OR3 (N1699, N1677, N592, N1456);
buf BUF1 (N1700, N1699);
or OR2 (N1701, N1691, N783);
nand NAND2 (N1702, N1688, N705);
and AND3 (N1703, N1695, N728, N161);
or OR4 (N1704, N1684, N368, N1619, N536);
buf BUF1 (N1705, N1700);
xor XOR2 (N1706, N1705, N1408);
nor NOR4 (N1707, N1704, N894, N1333, N915);
or OR4 (N1708, N1701, N448, N954, N496);
not NOT1 (N1709, N1708);
or OR4 (N1710, N1706, N578, N1628, N234);
nor NOR2 (N1711, N1707, N365);
xor XOR2 (N1712, N1680, N299);
and AND2 (N1713, N1683, N995);
or OR3 (N1714, N1710, N1614, N522);
buf BUF1 (N1715, N1712);
buf BUF1 (N1716, N1703);
xor XOR2 (N1717, N1709, N728);
and AND2 (N1718, N1713, N948);
or OR4 (N1719, N1718, N1268, N693, N1286);
not NOT1 (N1720, N1698);
nor NOR2 (N1721, N1714, N1318);
xor XOR2 (N1722, N1693, N538);
not NOT1 (N1723, N1720);
nand NAND3 (N1724, N1719, N1427, N1713);
nor NOR4 (N1725, N1716, N421, N1217, N51);
nand NAND2 (N1726, N1711, N93);
nor NOR3 (N1727, N1721, N360, N1434);
nand NAND4 (N1728, N1724, N365, N100, N1408);
and AND3 (N1729, N1702, N1153, N332);
not NOT1 (N1730, N1722);
and AND4 (N1731, N1725, N1249, N833, N1608);
and AND2 (N1732, N1730, N135);
not NOT1 (N1733, N1717);
xor XOR2 (N1734, N1696, N554);
nand NAND4 (N1735, N1727, N699, N497, N341);
and AND4 (N1736, N1732, N915, N596, N121);
xor XOR2 (N1737, N1728, N1069);
nand NAND4 (N1738, N1733, N886, N332, N1027);
not NOT1 (N1739, N1723);
not NOT1 (N1740, N1734);
buf BUF1 (N1741, N1715);
buf BUF1 (N1742, N1738);
xor XOR2 (N1743, N1736, N1013);
or OR3 (N1744, N1737, N377, N1587);
nand NAND4 (N1745, N1740, N937, N1114, N1467);
and AND3 (N1746, N1729, N216, N818);
buf BUF1 (N1747, N1726);
or OR2 (N1748, N1747, N1451);
not NOT1 (N1749, N1744);
buf BUF1 (N1750, N1731);
nor NOR4 (N1751, N1735, N1482, N117, N1609);
buf BUF1 (N1752, N1743);
nor NOR3 (N1753, N1750, N592, N86);
xor XOR2 (N1754, N1745, N1739);
nor NOR4 (N1755, N609, N182, N1047, N581);
and AND3 (N1756, N1751, N437, N416);
or OR3 (N1757, N1754, N1485, N643);
or OR3 (N1758, N1741, N1733, N61);
buf BUF1 (N1759, N1758);
xor XOR2 (N1760, N1757, N816);
nand NAND3 (N1761, N1749, N469, N817);
buf BUF1 (N1762, N1760);
nor NOR2 (N1763, N1752, N946);
nor NOR2 (N1764, N1755, N1758);
or OR3 (N1765, N1759, N343, N996);
nand NAND2 (N1766, N1748, N681);
or OR3 (N1767, N1762, N31, N1636);
nor NOR3 (N1768, N1756, N1128, N1656);
nor NOR4 (N1769, N1761, N45, N554, N1597);
and AND4 (N1770, N1753, N905, N89, N125);
or OR2 (N1771, N1769, N1219);
buf BUF1 (N1772, N1764);
or OR2 (N1773, N1768, N1578);
nor NOR4 (N1774, N1771, N358, N1339, N1024);
or OR2 (N1775, N1774, N651);
nor NOR2 (N1776, N1746, N271);
nor NOR3 (N1777, N1742, N604, N1015);
and AND4 (N1778, N1772, N965, N446, N990);
not NOT1 (N1779, N1767);
xor XOR2 (N1780, N1776, N781);
not NOT1 (N1781, N1775);
nor NOR2 (N1782, N1780, N70);
buf BUF1 (N1783, N1765);
nand NAND4 (N1784, N1770, N1181, N1348, N116);
not NOT1 (N1785, N1782);
or OR4 (N1786, N1785, N1093, N325, N1410);
xor XOR2 (N1787, N1777, N1524);
nor NOR3 (N1788, N1787, N1729, N451);
or OR4 (N1789, N1778, N1470, N1672, N468);
nor NOR3 (N1790, N1789, N137, N734);
nand NAND3 (N1791, N1784, N1699, N414);
buf BUF1 (N1792, N1790);
and AND2 (N1793, N1763, N1069);
nand NAND4 (N1794, N1786, N118, N1293, N1455);
xor XOR2 (N1795, N1773, N565);
and AND2 (N1796, N1783, N1503);
nand NAND4 (N1797, N1788, N666, N1597, N899);
or OR4 (N1798, N1779, N1235, N702, N607);
and AND4 (N1799, N1795, N1578, N1013, N1227);
and AND2 (N1800, N1796, N1413);
xor XOR2 (N1801, N1791, N1756);
or OR4 (N1802, N1799, N831, N641, N523);
or OR4 (N1803, N1793, N320, N655, N626);
and AND4 (N1804, N1798, N52, N810, N1175);
nand NAND2 (N1805, N1794, N1615);
not NOT1 (N1806, N1797);
nor NOR4 (N1807, N1802, N1403, N1477, N775);
not NOT1 (N1808, N1801);
nand NAND3 (N1809, N1800, N1231, N1021);
xor XOR2 (N1810, N1803, N1680);
xor XOR2 (N1811, N1808, N1103);
xor XOR2 (N1812, N1781, N253);
buf BUF1 (N1813, N1766);
nand NAND2 (N1814, N1810, N291);
nand NAND3 (N1815, N1806, N541, N743);
buf BUF1 (N1816, N1814);
buf BUF1 (N1817, N1812);
and AND2 (N1818, N1792, N1159);
nor NOR2 (N1819, N1813, N828);
not NOT1 (N1820, N1804);
nor NOR4 (N1821, N1818, N1633, N1563, N610);
nor NOR4 (N1822, N1816, N969, N178, N113);
xor XOR2 (N1823, N1811, N1807);
nor NOR2 (N1824, N347, N1350);
buf BUF1 (N1825, N1815);
nand NAND2 (N1826, N1809, N1143);
nor NOR3 (N1827, N1821, N663, N1772);
and AND2 (N1828, N1820, N1306);
nor NOR3 (N1829, N1824, N1512, N1294);
and AND2 (N1830, N1819, N786);
buf BUF1 (N1831, N1823);
not NOT1 (N1832, N1825);
buf BUF1 (N1833, N1828);
not NOT1 (N1834, N1831);
and AND3 (N1835, N1827, N72, N1609);
xor XOR2 (N1836, N1822, N891);
not NOT1 (N1837, N1817);
or OR2 (N1838, N1835, N1544);
not NOT1 (N1839, N1830);
or OR3 (N1840, N1832, N240, N252);
buf BUF1 (N1841, N1838);
and AND4 (N1842, N1805, N1504, N619, N233);
not NOT1 (N1843, N1840);
nand NAND2 (N1844, N1826, N76);
not NOT1 (N1845, N1836);
buf BUF1 (N1846, N1834);
nor NOR3 (N1847, N1833, N1069, N354);
nand NAND2 (N1848, N1843, N619);
or OR2 (N1849, N1847, N435);
nand NAND4 (N1850, N1846, N41, N1363, N947);
xor XOR2 (N1851, N1839, N1721);
or OR4 (N1852, N1844, N1670, N1258, N1428);
xor XOR2 (N1853, N1848, N1765);
and AND2 (N1854, N1849, N1256);
nor NOR2 (N1855, N1854, N239);
buf BUF1 (N1856, N1852);
nor NOR4 (N1857, N1829, N1243, N1773, N567);
not NOT1 (N1858, N1851);
xor XOR2 (N1859, N1837, N833);
not NOT1 (N1860, N1856);
nand NAND3 (N1861, N1855, N803, N1227);
and AND4 (N1862, N1861, N970, N420, N352);
nor NOR2 (N1863, N1850, N1646);
nand NAND4 (N1864, N1841, N601, N288, N325);
not NOT1 (N1865, N1853);
nor NOR4 (N1866, N1863, N1009, N850, N1600);
not NOT1 (N1867, N1862);
not NOT1 (N1868, N1860);
buf BUF1 (N1869, N1864);
xor XOR2 (N1870, N1845, N815);
or OR3 (N1871, N1859, N970, N527);
and AND4 (N1872, N1869, N855, N220, N1560);
or OR3 (N1873, N1872, N307, N382);
or OR2 (N1874, N1870, N1024);
xor XOR2 (N1875, N1858, N1589);
nand NAND3 (N1876, N1871, N382, N1582);
xor XOR2 (N1877, N1865, N1786);
not NOT1 (N1878, N1868);
nand NAND2 (N1879, N1876, N394);
or OR4 (N1880, N1877, N550, N67, N1752);
not NOT1 (N1881, N1867);
not NOT1 (N1882, N1842);
not NOT1 (N1883, N1866);
not NOT1 (N1884, N1875);
buf BUF1 (N1885, N1873);
not NOT1 (N1886, N1885);
and AND4 (N1887, N1881, N192, N1565, N1784);
buf BUF1 (N1888, N1887);
buf BUF1 (N1889, N1883);
and AND4 (N1890, N1857, N551, N2, N617);
and AND4 (N1891, N1886, N1723, N558, N376);
and AND4 (N1892, N1878, N1670, N888, N548);
nor NOR4 (N1893, N1889, N771, N1619, N1328);
nand NAND2 (N1894, N1888, N1056);
nor NOR2 (N1895, N1880, N24);
xor XOR2 (N1896, N1891, N990);
buf BUF1 (N1897, N1896);
nand NAND2 (N1898, N1892, N1076);
nor NOR3 (N1899, N1894, N629, N18);
not NOT1 (N1900, N1898);
nand NAND3 (N1901, N1874, N1272, N1003);
buf BUF1 (N1902, N1879);
not NOT1 (N1903, N1882);
or OR3 (N1904, N1884, N1016, N1811);
nor NOR4 (N1905, N1904, N380, N568, N1787);
or OR3 (N1906, N1903, N291, N130);
or OR2 (N1907, N1901, N1678);
nor NOR3 (N1908, N1899, N1729, N474);
and AND4 (N1909, N1906, N1080, N911, N952);
xor XOR2 (N1910, N1908, N1388);
nand NAND4 (N1911, N1902, N804, N1110, N616);
and AND3 (N1912, N1895, N1696, N808);
nand NAND4 (N1913, N1909, N1557, N971, N285);
or OR3 (N1914, N1913, N1212, N1606);
xor XOR2 (N1915, N1912, N1657);
xor XOR2 (N1916, N1893, N978);
xor XOR2 (N1917, N1907, N359);
nand NAND3 (N1918, N1890, N616, N175);
or OR2 (N1919, N1917, N1679);
nand NAND3 (N1920, N1918, N1683, N86);
xor XOR2 (N1921, N1905, N578);
and AND3 (N1922, N1911, N1467, N1141);
and AND4 (N1923, N1914, N745, N766, N1059);
or OR4 (N1924, N1900, N326, N107, N975);
and AND2 (N1925, N1922, N462);
or OR4 (N1926, N1925, N230, N614, N1641);
and AND2 (N1927, N1919, N733);
or OR4 (N1928, N1916, N732, N817, N784);
and AND2 (N1929, N1921, N531);
nand NAND2 (N1930, N1923, N232);
buf BUF1 (N1931, N1910);
buf BUF1 (N1932, N1924);
buf BUF1 (N1933, N1931);
or OR2 (N1934, N1897, N1883);
or OR2 (N1935, N1929, N672);
or OR4 (N1936, N1934, N1163, N626, N293);
xor XOR2 (N1937, N1915, N18);
or OR3 (N1938, N1926, N1731, N1571);
buf BUF1 (N1939, N1920);
not NOT1 (N1940, N1927);
buf BUF1 (N1941, N1935);
xor XOR2 (N1942, N1940, N1116);
nor NOR2 (N1943, N1938, N1264);
nand NAND3 (N1944, N1943, N1360, N674);
or OR4 (N1945, N1942, N1686, N19, N1838);
buf BUF1 (N1946, N1944);
or OR3 (N1947, N1939, N1437, N1811);
xor XOR2 (N1948, N1933, N1769);
buf BUF1 (N1949, N1946);
and AND3 (N1950, N1945, N438, N1666);
nor NOR4 (N1951, N1937, N1769, N385, N201);
nor NOR3 (N1952, N1947, N962, N1842);
xor XOR2 (N1953, N1951, N49);
buf BUF1 (N1954, N1930);
nand NAND4 (N1955, N1932, N1790, N1075, N595);
nand NAND2 (N1956, N1952, N1324);
nand NAND3 (N1957, N1948, N1243, N623);
nand NAND3 (N1958, N1936, N1342, N461);
and AND4 (N1959, N1954, N1693, N1537, N598);
xor XOR2 (N1960, N1953, N433);
nor NOR3 (N1961, N1941, N1003, N909);
nand NAND3 (N1962, N1928, N1078, N1460);
and AND4 (N1963, N1956, N708, N1, N1166);
not NOT1 (N1964, N1959);
not NOT1 (N1965, N1957);
buf BUF1 (N1966, N1950);
not NOT1 (N1967, N1966);
xor XOR2 (N1968, N1961, N327);
buf BUF1 (N1969, N1962);
not NOT1 (N1970, N1960);
or OR2 (N1971, N1970, N179);
and AND3 (N1972, N1969, N188, N75);
nand NAND3 (N1973, N1965, N1587, N1260);
and AND4 (N1974, N1971, N1664, N1122, N272);
or OR3 (N1975, N1967, N785, N1056);
nor NOR3 (N1976, N1972, N1444, N840);
or OR2 (N1977, N1973, N1840);
nand NAND3 (N1978, N1974, N1769, N1971);
nand NAND3 (N1979, N1963, N754, N316);
and AND2 (N1980, N1979, N1939);
nand NAND4 (N1981, N1949, N1110, N637, N1177);
or OR4 (N1982, N1977, N1959, N807, N350);
buf BUF1 (N1983, N1968);
not NOT1 (N1984, N1976);
and AND3 (N1985, N1958, N1396, N1923);
buf BUF1 (N1986, N1983);
buf BUF1 (N1987, N1955);
not NOT1 (N1988, N1984);
and AND2 (N1989, N1986, N1182);
or OR3 (N1990, N1978, N983, N186);
or OR2 (N1991, N1990, N1469);
buf BUF1 (N1992, N1987);
nor NOR2 (N1993, N1985, N740);
not NOT1 (N1994, N1975);
xor XOR2 (N1995, N1982, N212);
buf BUF1 (N1996, N1993);
nor NOR4 (N1997, N1995, N1744, N1719, N1231);
nand NAND3 (N1998, N1980, N1833, N818);
buf BUF1 (N1999, N1964);
not NOT1 (N2000, N1997);
xor XOR2 (N2001, N1996, N492);
nand NAND2 (N2002, N1991, N777);
xor XOR2 (N2003, N1988, N1232);
or OR3 (N2004, N2003, N1414, N676);
xor XOR2 (N2005, N2002, N1313);
not NOT1 (N2006, N2004);
not NOT1 (N2007, N1989);
xor XOR2 (N2008, N2000, N1140);
nand NAND2 (N2009, N2005, N550);
xor XOR2 (N2010, N2006, N1609);
nand NAND3 (N2011, N2008, N1247, N1426);
buf BUF1 (N2012, N2009);
buf BUF1 (N2013, N2007);
nand NAND2 (N2014, N1994, N1754);
nor NOR2 (N2015, N1998, N1603);
and AND2 (N2016, N2013, N1905);
xor XOR2 (N2017, N2012, N381);
not NOT1 (N2018, N1999);
nand NAND2 (N2019, N2010, N1195);
nand NAND2 (N2020, N2001, N336);
nand NAND3 (N2021, N2019, N1889, N954);
buf BUF1 (N2022, N2021);
nor NOR3 (N2023, N1992, N1134, N274);
and AND4 (N2024, N1981, N660, N282, N856);
buf BUF1 (N2025, N2015);
xor XOR2 (N2026, N2024, N1689);
or OR3 (N2027, N2016, N1192, N747);
or OR4 (N2028, N2026, N1561, N72, N58);
nor NOR4 (N2029, N2028, N912, N1012, N170);
or OR3 (N2030, N2020, N145, N1767);
xor XOR2 (N2031, N2018, N1654);
buf BUF1 (N2032, N2011);
xor XOR2 (N2033, N2025, N627);
xor XOR2 (N2034, N2023, N650);
nor NOR3 (N2035, N2031, N994, N1744);
or OR4 (N2036, N2017, N1106, N1542, N839);
nand NAND3 (N2037, N2036, N1249, N1888);
or OR3 (N2038, N2030, N1520, N1016);
not NOT1 (N2039, N2035);
nand NAND4 (N2040, N2022, N718, N1606, N517);
or OR4 (N2041, N2040, N1293, N1069, N940);
not NOT1 (N2042, N2014);
not NOT1 (N2043, N2042);
nor NOR2 (N2044, N2037, N121);
and AND3 (N2045, N2038, N1184, N757);
or OR2 (N2046, N2029, N1128);
not NOT1 (N2047, N2027);
or OR3 (N2048, N2039, N845, N1571);
not NOT1 (N2049, N2046);
and AND3 (N2050, N2033, N826, N1088);
or OR3 (N2051, N2047, N1588, N1442);
and AND4 (N2052, N2051, N1343, N1260, N1140);
nor NOR3 (N2053, N2043, N79, N1736);
nor NOR3 (N2054, N2050, N611, N881);
nand NAND2 (N2055, N2044, N1659);
not NOT1 (N2056, N2048);
and AND3 (N2057, N2041, N616, N1126);
nor NOR3 (N2058, N2032, N1131, N584);
xor XOR2 (N2059, N2045, N1587);
nand NAND2 (N2060, N2049, N543);
and AND4 (N2061, N2057, N1243, N728, N1635);
or OR3 (N2062, N2055, N1795, N1855);
nor NOR2 (N2063, N2052, N1717);
not NOT1 (N2064, N2059);
nand NAND3 (N2065, N2058, N1139, N1956);
xor XOR2 (N2066, N2065, N264);
or OR3 (N2067, N2064, N268, N90);
and AND4 (N2068, N2060, N1759, N477, N1088);
xor XOR2 (N2069, N2062, N1883);
not NOT1 (N2070, N2061);
nand NAND3 (N2071, N2067, N1097, N1716);
xor XOR2 (N2072, N2034, N1123);
or OR2 (N2073, N2053, N1986);
not NOT1 (N2074, N2063);
nor NOR4 (N2075, N2069, N400, N1377, N1981);
buf BUF1 (N2076, N2072);
and AND2 (N2077, N2066, N312);
buf BUF1 (N2078, N2077);
or OR4 (N2079, N2068, N882, N107, N607);
xor XOR2 (N2080, N2074, N1254);
nor NOR4 (N2081, N2054, N1972, N1642, N1677);
and AND2 (N2082, N2071, N872);
not NOT1 (N2083, N2075);
and AND4 (N2084, N2073, N1948, N1354, N958);
or OR4 (N2085, N2081, N1303, N947, N296);
or OR3 (N2086, N2079, N1869, N1727);
not NOT1 (N2087, N2084);
xor XOR2 (N2088, N2078, N1338);
not NOT1 (N2089, N2085);
nand NAND2 (N2090, N2088, N946);
nand NAND2 (N2091, N2089, N996);
buf BUF1 (N2092, N2083);
nand NAND4 (N2093, N2076, N958, N1913, N809);
xor XOR2 (N2094, N2093, N71);
nor NOR4 (N2095, N2080, N38, N1527, N1618);
and AND2 (N2096, N2091, N1838);
and AND4 (N2097, N2087, N1004, N562, N1749);
not NOT1 (N2098, N2092);
nand NAND4 (N2099, N2094, N1088, N1968, N1351);
or OR4 (N2100, N2095, N1888, N200, N1498);
nor NOR4 (N2101, N2082, N754, N1104, N1125);
or OR2 (N2102, N2090, N1808);
buf BUF1 (N2103, N2099);
nand NAND3 (N2104, N2070, N1714, N1835);
nor NOR2 (N2105, N2102, N798);
buf BUF1 (N2106, N2104);
xor XOR2 (N2107, N2103, N440);
and AND4 (N2108, N2096, N498, N1786, N851);
or OR3 (N2109, N2056, N762, N201);
or OR3 (N2110, N2109, N250, N1942);
not NOT1 (N2111, N2097);
or OR4 (N2112, N2098, N582, N1671, N1186);
buf BUF1 (N2113, N2101);
xor XOR2 (N2114, N2112, N1748);
xor XOR2 (N2115, N2110, N1527);
nand NAND3 (N2116, N2107, N534, N1972);
not NOT1 (N2117, N2116);
xor XOR2 (N2118, N2108, N1145);
and AND3 (N2119, N2118, N937, N92);
not NOT1 (N2120, N2105);
nand NAND3 (N2121, N2114, N670, N1598);
buf BUF1 (N2122, N2111);
buf BUF1 (N2123, N2113);
and AND3 (N2124, N2119, N618, N109);
or OR2 (N2125, N2100, N357);
and AND2 (N2126, N2120, N504);
or OR3 (N2127, N2124, N1709, N340);
or OR2 (N2128, N2127, N1138);
nand NAND4 (N2129, N2123, N1193, N451, N1490);
nand NAND4 (N2130, N2128, N806, N256, N1678);
nand NAND3 (N2131, N2126, N1922, N2032);
nand NAND3 (N2132, N2130, N758, N1764);
and AND4 (N2133, N2086, N2109, N1230, N429);
or OR2 (N2134, N2133, N1671);
nand NAND4 (N2135, N2106, N330, N1829, N1353);
xor XOR2 (N2136, N2125, N480);
and AND4 (N2137, N2134, N687, N1084, N1451);
xor XOR2 (N2138, N2121, N1410);
nand NAND4 (N2139, N2138, N118, N2014, N1848);
not NOT1 (N2140, N2131);
buf BUF1 (N2141, N2140);
buf BUF1 (N2142, N2136);
buf BUF1 (N2143, N2137);
xor XOR2 (N2144, N2139, N1176);
nor NOR4 (N2145, N2142, N2043, N724, N1324);
buf BUF1 (N2146, N2144);
nor NOR4 (N2147, N2135, N1525, N451, N1994);
or OR3 (N2148, N2122, N1896, N653);
buf BUF1 (N2149, N2129);
and AND2 (N2150, N2145, N1376);
nand NAND2 (N2151, N2146, N125);
and AND3 (N2152, N2143, N717, N1510);
and AND2 (N2153, N2115, N953);
or OR3 (N2154, N2141, N1581, N1470);
nor NOR3 (N2155, N2148, N1312, N167);
not NOT1 (N2156, N2150);
nand NAND2 (N2157, N2147, N78);
nand NAND4 (N2158, N2154, N738, N818, N462);
not NOT1 (N2159, N2152);
not NOT1 (N2160, N2117);
or OR3 (N2161, N2155, N738, N1984);
not NOT1 (N2162, N2160);
or OR2 (N2163, N2149, N184);
xor XOR2 (N2164, N2163, N168);
not NOT1 (N2165, N2162);
not NOT1 (N2166, N2159);
not NOT1 (N2167, N2151);
xor XOR2 (N2168, N2153, N1167);
nor NOR3 (N2169, N2132, N144, N2115);
nand NAND2 (N2170, N2161, N952);
and AND4 (N2171, N2167, N1656, N15, N312);
or OR2 (N2172, N2170, N1318);
or OR2 (N2173, N2172, N825);
buf BUF1 (N2174, N2158);
nand NAND4 (N2175, N2166, N1584, N4, N816);
and AND4 (N2176, N2156, N755, N732, N141);
nor NOR4 (N2177, N2174, N333, N1536, N1514);
and AND3 (N2178, N2168, N1434, N1483);
buf BUF1 (N2179, N2165);
nand NAND2 (N2180, N2178, N1192);
nand NAND3 (N2181, N2171, N1495, N1276);
or OR2 (N2182, N2177, N298);
nor NOR4 (N2183, N2173, N1543, N1842, N417);
xor XOR2 (N2184, N2179, N360);
nand NAND4 (N2185, N2184, N2152, N1303, N728);
or OR4 (N2186, N2176, N1924, N1429, N1593);
nor NOR2 (N2187, N2175, N1049);
not NOT1 (N2188, N2185);
or OR3 (N2189, N2187, N891, N1084);
and AND3 (N2190, N2180, N1365, N690);
not NOT1 (N2191, N2181);
xor XOR2 (N2192, N2157, N167);
not NOT1 (N2193, N2164);
buf BUF1 (N2194, N2193);
and AND2 (N2195, N2192, N1750);
and AND3 (N2196, N2189, N2055, N1991);
or OR2 (N2197, N2188, N718);
and AND4 (N2198, N2196, N1432, N1766, N620);
or OR3 (N2199, N2186, N1539, N1981);
nor NOR3 (N2200, N2190, N1550, N578);
xor XOR2 (N2201, N2197, N1437);
not NOT1 (N2202, N2201);
or OR2 (N2203, N2195, N1560);
or OR2 (N2204, N2200, N220);
xor XOR2 (N2205, N2199, N1439);
or OR3 (N2206, N2205, N2012, N970);
buf BUF1 (N2207, N2182);
or OR4 (N2208, N2198, N1769, N278, N2038);
buf BUF1 (N2209, N2202);
not NOT1 (N2210, N2207);
and AND2 (N2211, N2204, N726);
nor NOR3 (N2212, N2194, N1359, N152);
nand NAND4 (N2213, N2203, N1675, N1700, N419);
nand NAND3 (N2214, N2210, N1766, N1331);
and AND3 (N2215, N2191, N1174, N1957);
or OR3 (N2216, N2209, N1366, N433);
nor NOR4 (N2217, N2211, N1812, N1032, N967);
xor XOR2 (N2218, N2214, N1610);
and AND4 (N2219, N2213, N14, N886, N749);
and AND3 (N2220, N2183, N595, N1630);
buf BUF1 (N2221, N2219);
nand NAND2 (N2222, N2216, N1459);
xor XOR2 (N2223, N2218, N873);
nor NOR4 (N2224, N2212, N466, N1196, N1448);
or OR4 (N2225, N2208, N1300, N272, N524);
nand NAND4 (N2226, N2221, N1588, N1693, N1809);
buf BUF1 (N2227, N2206);
buf BUF1 (N2228, N2217);
or OR2 (N2229, N2224, N1042);
xor XOR2 (N2230, N2222, N829);
nand NAND2 (N2231, N2227, N96);
nor NOR2 (N2232, N2229, N723);
and AND2 (N2233, N2220, N1539);
buf BUF1 (N2234, N2226);
nand NAND4 (N2235, N2228, N474, N1258, N2081);
nor NOR2 (N2236, N2233, N1641);
nor NOR3 (N2237, N2234, N221, N1704);
nand NAND3 (N2238, N2169, N1982, N1357);
nor NOR4 (N2239, N2236, N1525, N1338, N404);
nor NOR4 (N2240, N2230, N760, N147, N2149);
buf BUF1 (N2241, N2231);
buf BUF1 (N2242, N2238);
and AND2 (N2243, N2241, N1127);
nor NOR4 (N2244, N2232, N136, N827, N154);
xor XOR2 (N2245, N2225, N1346);
and AND3 (N2246, N2242, N872, N217);
not NOT1 (N2247, N2246);
buf BUF1 (N2248, N2237);
nand NAND3 (N2249, N2223, N926, N1062);
and AND4 (N2250, N2245, N753, N1508, N1368);
nor NOR2 (N2251, N2215, N179);
nor NOR2 (N2252, N2248, N1827);
not NOT1 (N2253, N2250);
and AND4 (N2254, N2239, N81, N56, N1294);
buf BUF1 (N2255, N2249);
not NOT1 (N2256, N2255);
and AND2 (N2257, N2256, N1781);
nand NAND4 (N2258, N2244, N202, N1159, N479);
not NOT1 (N2259, N2247);
xor XOR2 (N2260, N2258, N150);
xor XOR2 (N2261, N2235, N763);
nand NAND2 (N2262, N2257, N1319);
xor XOR2 (N2263, N2259, N483);
xor XOR2 (N2264, N2263, N1831);
or OR3 (N2265, N2251, N264, N854);
buf BUF1 (N2266, N2240);
and AND4 (N2267, N2253, N731, N412, N1369);
and AND4 (N2268, N2254, N1625, N1752, N63);
nor NOR2 (N2269, N2267, N404);
and AND4 (N2270, N2252, N1329, N1980, N1141);
not NOT1 (N2271, N2261);
xor XOR2 (N2272, N2264, N426);
or OR2 (N2273, N2269, N2186);
or OR2 (N2274, N2272, N1744);
nor NOR4 (N2275, N2262, N1575, N778, N821);
and AND2 (N2276, N2268, N1816);
buf BUF1 (N2277, N2271);
buf BUF1 (N2278, N2266);
xor XOR2 (N2279, N2243, N661);
and AND4 (N2280, N2274, N968, N1087, N593);
or OR3 (N2281, N2279, N2072, N1755);
or OR4 (N2282, N2275, N2146, N1395, N2178);
nor NOR3 (N2283, N2280, N368, N2179);
nand NAND3 (N2284, N2278, N283, N76);
or OR2 (N2285, N2260, N1301);
or OR2 (N2286, N2285, N1000);
nand NAND4 (N2287, N2277, N1210, N2274, N580);
or OR3 (N2288, N2265, N143, N1617);
not NOT1 (N2289, N2276);
xor XOR2 (N2290, N2270, N2166);
nor NOR2 (N2291, N2290, N2089);
or OR3 (N2292, N2284, N371, N217);
or OR4 (N2293, N2292, N1359, N1666, N712);
xor XOR2 (N2294, N2273, N850);
and AND2 (N2295, N2289, N1443);
and AND3 (N2296, N2294, N468, N806);
buf BUF1 (N2297, N2293);
or OR4 (N2298, N2295, N1466, N870, N235);
xor XOR2 (N2299, N2288, N2072);
not NOT1 (N2300, N2296);
xor XOR2 (N2301, N2283, N986);
nand NAND2 (N2302, N2286, N2037);
and AND2 (N2303, N2298, N1275);
or OR3 (N2304, N2301, N1740, N707);
nand NAND2 (N2305, N2299, N1589);
buf BUF1 (N2306, N2300);
xor XOR2 (N2307, N2302, N719);
and AND2 (N2308, N2297, N85);
xor XOR2 (N2309, N2282, N1418);
nand NAND3 (N2310, N2307, N726, N178);
and AND3 (N2311, N2305, N875, N945);
buf BUF1 (N2312, N2287);
buf BUF1 (N2313, N2310);
nand NAND2 (N2314, N2306, N1149);
and AND4 (N2315, N2309, N1651, N1140, N840);
nand NAND3 (N2316, N2315, N1494, N752);
and AND4 (N2317, N2311, N1906, N1070, N1652);
not NOT1 (N2318, N2317);
xor XOR2 (N2319, N2303, N1359);
not NOT1 (N2320, N2281);
not NOT1 (N2321, N2314);
buf BUF1 (N2322, N2308);
or OR3 (N2323, N2291, N492, N592);
buf BUF1 (N2324, N2320);
nand NAND2 (N2325, N2316, N186);
or OR4 (N2326, N2323, N784, N2304, N1556);
nor NOR4 (N2327, N922, N2034, N701, N2269);
buf BUF1 (N2328, N2327);
buf BUF1 (N2329, N2312);
buf BUF1 (N2330, N2321);
xor XOR2 (N2331, N2326, N738);
xor XOR2 (N2332, N2325, N256);
or OR2 (N2333, N2328, N1871);
buf BUF1 (N2334, N2319);
xor XOR2 (N2335, N2332, N1075);
nor NOR4 (N2336, N2313, N2225, N1526, N226);
not NOT1 (N2337, N2334);
nor NOR2 (N2338, N2322, N1535);
not NOT1 (N2339, N2333);
and AND3 (N2340, N2330, N938, N751);
nor NOR4 (N2341, N2336, N2193, N1789, N1612);
not NOT1 (N2342, N2331);
nor NOR4 (N2343, N2338, N391, N1773, N4);
buf BUF1 (N2344, N2342);
nand NAND3 (N2345, N2318, N303, N227);
nand NAND2 (N2346, N2337, N1021);
not NOT1 (N2347, N2343);
xor XOR2 (N2348, N2341, N312);
xor XOR2 (N2349, N2348, N925);
buf BUF1 (N2350, N2324);
and AND2 (N2351, N2346, N1456);
or OR3 (N2352, N2335, N1032, N27);
xor XOR2 (N2353, N2349, N1928);
not NOT1 (N2354, N2350);
and AND3 (N2355, N2329, N664, N1871);
nor NOR3 (N2356, N2355, N1055, N1717);
and AND4 (N2357, N2340, N1220, N1516, N1529);
not NOT1 (N2358, N2352);
and AND2 (N2359, N2344, N1776);
not NOT1 (N2360, N2359);
or OR2 (N2361, N2356, N759);
not NOT1 (N2362, N2345);
not NOT1 (N2363, N2339);
and AND4 (N2364, N2353, N730, N2062, N88);
nand NAND2 (N2365, N2360, N1538);
buf BUF1 (N2366, N2354);
and AND2 (N2367, N2366, N2146);
nor NOR3 (N2368, N2358, N19, N2);
or OR4 (N2369, N2365, N764, N610, N675);
nor NOR3 (N2370, N2361, N1043, N1225);
not NOT1 (N2371, N2368);
and AND3 (N2372, N2363, N1691, N679);
buf BUF1 (N2373, N2364);
or OR4 (N2374, N2369, N2003, N34, N855);
and AND3 (N2375, N2372, N15, N657);
and AND3 (N2376, N2362, N1111, N234);
xor XOR2 (N2377, N2375, N1223);
buf BUF1 (N2378, N2367);
not NOT1 (N2379, N2370);
xor XOR2 (N2380, N2357, N1961);
not NOT1 (N2381, N2373);
nand NAND4 (N2382, N2378, N999, N1049, N1357);
not NOT1 (N2383, N2374);
nand NAND4 (N2384, N2383, N1828, N1962, N878);
not NOT1 (N2385, N2381);
nor NOR4 (N2386, N2380, N925, N158, N242);
nand NAND4 (N2387, N2379, N1737, N1448, N1246);
xor XOR2 (N2388, N2347, N2109);
and AND2 (N2389, N2384, N2179);
nand NAND4 (N2390, N2382, N518, N750, N701);
or OR4 (N2391, N2371, N2009, N707, N162);
nand NAND2 (N2392, N2385, N1747);
not NOT1 (N2393, N2386);
xor XOR2 (N2394, N2388, N2384);
nand NAND3 (N2395, N2377, N1906, N2282);
nor NOR3 (N2396, N2393, N1856, N258);
buf BUF1 (N2397, N2389);
xor XOR2 (N2398, N2397, N1900);
and AND3 (N2399, N2390, N666, N1168);
buf BUF1 (N2400, N2394);
xor XOR2 (N2401, N2392, N2133);
or OR4 (N2402, N2401, N1566, N1063, N1729);
buf BUF1 (N2403, N2351);
or OR2 (N2404, N2376, N837);
xor XOR2 (N2405, N2403, N1515);
nor NOR2 (N2406, N2391, N2216);
nand NAND4 (N2407, N2395, N637, N2381, N1484);
or OR2 (N2408, N2402, N1440);
and AND3 (N2409, N2398, N1319, N1617);
or OR4 (N2410, N2387, N1251, N1558, N750);
not NOT1 (N2411, N2404);
or OR4 (N2412, N2407, N2001, N1224, N1684);
nand NAND4 (N2413, N2406, N2353, N1502, N2016);
nand NAND2 (N2414, N2411, N1897);
xor XOR2 (N2415, N2399, N2211);
nand NAND4 (N2416, N2408, N551, N226, N29);
not NOT1 (N2417, N2414);
nand NAND3 (N2418, N2409, N465, N2378);
nor NOR4 (N2419, N2410, N1978, N1029, N1004);
not NOT1 (N2420, N2412);
buf BUF1 (N2421, N2405);
xor XOR2 (N2422, N2413, N1442);
buf BUF1 (N2423, N2418);
xor XOR2 (N2424, N2416, N2151);
xor XOR2 (N2425, N2421, N2043);
not NOT1 (N2426, N2415);
nand NAND4 (N2427, N2396, N1056, N2162, N796);
xor XOR2 (N2428, N2419, N980);
or OR3 (N2429, N2417, N866, N1386);
and AND3 (N2430, N2400, N833, N1388);
or OR3 (N2431, N2427, N883, N644);
nor NOR4 (N2432, N2428, N878, N2125, N271);
not NOT1 (N2433, N2426);
not NOT1 (N2434, N2425);
or OR4 (N2435, N2422, N709, N1238, N610);
nand NAND2 (N2436, N2433, N1336);
nand NAND2 (N2437, N2420, N484);
buf BUF1 (N2438, N2435);
nand NAND4 (N2439, N2431, N2147, N1947, N1522);
not NOT1 (N2440, N2438);
nor NOR4 (N2441, N2432, N1738, N1635, N150);
not NOT1 (N2442, N2434);
not NOT1 (N2443, N2437);
xor XOR2 (N2444, N2423, N1930);
xor XOR2 (N2445, N2430, N1916);
and AND2 (N2446, N2436, N1829);
nand NAND2 (N2447, N2443, N200);
buf BUF1 (N2448, N2445);
xor XOR2 (N2449, N2424, N1664);
not NOT1 (N2450, N2444);
not NOT1 (N2451, N2440);
buf BUF1 (N2452, N2447);
nand NAND3 (N2453, N2439, N2032, N2223);
nor NOR4 (N2454, N2450, N2004, N2034, N393);
buf BUF1 (N2455, N2453);
xor XOR2 (N2456, N2442, N1303);
nand NAND3 (N2457, N2449, N890, N2077);
nor NOR2 (N2458, N2452, N1358);
buf BUF1 (N2459, N2441);
and AND4 (N2460, N2429, N2081, N227, N52);
nand NAND4 (N2461, N2451, N2157, N1821, N2313);
buf BUF1 (N2462, N2458);
nor NOR2 (N2463, N2457, N569);
buf BUF1 (N2464, N2461);
or OR2 (N2465, N2455, N1712);
or OR2 (N2466, N2454, N1922);
xor XOR2 (N2467, N2462, N1023);
nand NAND2 (N2468, N2463, N152);
or OR2 (N2469, N2468, N1775);
buf BUF1 (N2470, N2469);
not NOT1 (N2471, N2466);
or OR2 (N2472, N2465, N1466);
nor NOR4 (N2473, N2464, N1573, N747, N2463);
or OR2 (N2474, N2446, N1158);
buf BUF1 (N2475, N2460);
nand NAND2 (N2476, N2472, N1437);
not NOT1 (N2477, N2475);
xor XOR2 (N2478, N2467, N1844);
nor NOR3 (N2479, N2459, N2232, N2332);
and AND3 (N2480, N2479, N2056, N1961);
buf BUF1 (N2481, N2471);
or OR3 (N2482, N2448, N87, N2143);
not NOT1 (N2483, N2470);
or OR4 (N2484, N2478, N2154, N921, N2184);
or OR3 (N2485, N2477, N2472, N217);
nor NOR4 (N2486, N2482, N1183, N1947, N1159);
nor NOR3 (N2487, N2476, N1430, N649);
not NOT1 (N2488, N2485);
nor NOR3 (N2489, N2487, N905, N2218);
nor NOR2 (N2490, N2456, N395);
nor NOR4 (N2491, N2474, N946, N261, N2488);
nor NOR4 (N2492, N5, N1536, N920, N317);
and AND4 (N2493, N2481, N1130, N298, N219);
not NOT1 (N2494, N2480);
and AND3 (N2495, N2491, N1621, N45);
buf BUF1 (N2496, N2486);
or OR2 (N2497, N2492, N570);
buf BUF1 (N2498, N2483);
not NOT1 (N2499, N2484);
buf BUF1 (N2500, N2497);
or OR4 (N2501, N2490, N1738, N1725, N338);
and AND2 (N2502, N2494, N533);
nor NOR3 (N2503, N2499, N1299, N2409);
or OR3 (N2504, N2502, N283, N590);
or OR4 (N2505, N2489, N520, N2483, N463);
xor XOR2 (N2506, N2495, N738);
nor NOR3 (N2507, N2500, N2121, N358);
nand NAND3 (N2508, N2503, N1400, N1332);
or OR2 (N2509, N2505, N249);
buf BUF1 (N2510, N2506);
not NOT1 (N2511, N2498);
buf BUF1 (N2512, N2511);
and AND4 (N2513, N2473, N478, N1432, N306);
not NOT1 (N2514, N2496);
or OR2 (N2515, N2512, N2422);
buf BUF1 (N2516, N2508);
xor XOR2 (N2517, N2507, N2512);
or OR2 (N2518, N2515, N806);
xor XOR2 (N2519, N2513, N1949);
or OR2 (N2520, N2519, N2214);
xor XOR2 (N2521, N2518, N2124);
xor XOR2 (N2522, N2501, N1380);
endmodule