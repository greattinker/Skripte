// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N1001,N1009,N1010,N1005,N1002,N994,N978,N1008,N999,N1011;

nor NOR3 (N12, N3, N11, N4);
not NOT1 (N13, N10);
buf BUF1 (N14, N9);
or OR2 (N15, N5, N10);
and AND4 (N16, N9, N5, N2, N6);
or OR3 (N17, N2, N8, N7);
or OR3 (N18, N1, N11, N11);
nor NOR3 (N19, N7, N9, N4);
buf BUF1 (N20, N18);
nor NOR2 (N21, N4, N16);
buf BUF1 (N22, N9);
not NOT1 (N23, N2);
buf BUF1 (N24, N12);
and AND4 (N25, N22, N9, N19, N22);
or OR2 (N26, N3, N19);
nor NOR4 (N27, N14, N1, N25, N23);
buf BUF1 (N28, N14);
buf BUF1 (N29, N6);
or OR2 (N30, N26, N4);
and AND4 (N31, N20, N25, N24, N14);
and AND3 (N32, N7, N29, N4);
and AND3 (N33, N13, N30, N15);
nor NOR4 (N34, N9, N16, N22, N3);
or OR4 (N35, N3, N4, N6, N6);
xor XOR2 (N36, N2, N31);
xor XOR2 (N37, N9, N2);
nor NOR4 (N38, N21, N11, N37, N12);
or OR2 (N39, N29, N18);
xor XOR2 (N40, N36, N8);
nand NAND4 (N41, N32, N15, N38, N19);
or OR3 (N42, N20, N4, N35);
nand NAND4 (N43, N37, N32, N2, N29);
and AND2 (N44, N39, N6);
not NOT1 (N45, N33);
xor XOR2 (N46, N28, N12);
xor XOR2 (N47, N44, N7);
buf BUF1 (N48, N41);
not NOT1 (N49, N34);
or OR3 (N50, N42, N19, N11);
xor XOR2 (N51, N17, N6);
or OR4 (N52, N47, N23, N44, N51);
and AND2 (N53, N52, N34);
nor NOR4 (N54, N31, N43, N19, N17);
nand NAND3 (N55, N4, N9, N6);
and AND2 (N56, N53, N27);
nor NOR4 (N57, N5, N18, N23, N19);
xor XOR2 (N58, N56, N31);
xor XOR2 (N59, N46, N54);
or OR3 (N60, N3, N6, N15);
not NOT1 (N61, N59);
buf BUF1 (N62, N45);
not NOT1 (N63, N57);
and AND4 (N64, N55, N45, N4, N8);
and AND3 (N65, N63, N34, N22);
nor NOR4 (N66, N48, N29, N16, N40);
or OR3 (N67, N53, N49, N50);
xor XOR2 (N68, N63, N56);
not NOT1 (N69, N39);
not NOT1 (N70, N66);
and AND4 (N71, N67, N1, N50, N60);
nand NAND4 (N72, N29, N25, N16, N35);
xor XOR2 (N73, N61, N44);
xor XOR2 (N74, N64, N45);
nand NAND2 (N75, N73, N58);
nand NAND2 (N76, N64, N18);
nor NOR2 (N77, N69, N33);
and AND2 (N78, N62, N41);
or OR2 (N79, N72, N17);
or OR4 (N80, N77, N42, N8, N30);
not NOT1 (N81, N80);
xor XOR2 (N82, N68, N72);
xor XOR2 (N83, N81, N11);
nand NAND3 (N84, N76, N14, N48);
or OR3 (N85, N79, N45, N73);
xor XOR2 (N86, N84, N29);
and AND4 (N87, N82, N36, N23, N8);
not NOT1 (N88, N75);
nand NAND3 (N89, N87, N75, N58);
buf BUF1 (N90, N85);
buf BUF1 (N91, N65);
or OR4 (N92, N83, N70, N53, N13);
and AND4 (N93, N14, N8, N86, N90);
nand NAND4 (N94, N90, N28, N12, N7);
and AND3 (N95, N74, N24, N48);
nor NOR2 (N96, N36, N83);
and AND4 (N97, N93, N70, N94, N87);
and AND4 (N98, N71, N58, N48, N32);
xor XOR2 (N99, N13, N8);
xor XOR2 (N100, N88, N86);
nand NAND2 (N101, N96, N34);
buf BUF1 (N102, N98);
and AND3 (N103, N78, N87, N87);
not NOT1 (N104, N101);
not NOT1 (N105, N104);
buf BUF1 (N106, N89);
not NOT1 (N107, N97);
nor NOR3 (N108, N103, N29, N6);
and AND3 (N109, N105, N95, N96);
xor XOR2 (N110, N69, N50);
not NOT1 (N111, N100);
xor XOR2 (N112, N110, N13);
nand NAND4 (N113, N99, N51, N104, N28);
nand NAND3 (N114, N91, N65, N66);
not NOT1 (N115, N113);
not NOT1 (N116, N92);
or OR2 (N117, N106, N11);
buf BUF1 (N118, N102);
buf BUF1 (N119, N117);
or OR3 (N120, N115, N79, N45);
xor XOR2 (N121, N119, N38);
nor NOR2 (N122, N118, N42);
nor NOR3 (N123, N111, N52, N20);
nor NOR2 (N124, N107, N100);
not NOT1 (N125, N108);
xor XOR2 (N126, N123, N28);
or OR3 (N127, N121, N61, N43);
xor XOR2 (N128, N120, N67);
buf BUF1 (N129, N122);
buf BUF1 (N130, N116);
nor NOR2 (N131, N112, N10);
or OR2 (N132, N130, N101);
xor XOR2 (N133, N109, N52);
buf BUF1 (N134, N132);
nor NOR2 (N135, N129, N131);
and AND2 (N136, N30, N38);
xor XOR2 (N137, N124, N57);
nand NAND2 (N138, N127, N98);
xor XOR2 (N139, N136, N100);
not NOT1 (N140, N114);
nor NOR4 (N141, N137, N88, N44, N48);
xor XOR2 (N142, N139, N10);
buf BUF1 (N143, N134);
and AND3 (N144, N141, N126, N107);
nand NAND3 (N145, N6, N93, N96);
nand NAND3 (N146, N140, N132, N64);
not NOT1 (N147, N145);
nand NAND4 (N148, N125, N72, N96, N45);
nor NOR3 (N149, N148, N148, N125);
not NOT1 (N150, N138);
not NOT1 (N151, N146);
nor NOR3 (N152, N133, N106, N78);
buf BUF1 (N153, N151);
and AND4 (N154, N128, N85, N97, N133);
buf BUF1 (N155, N144);
buf BUF1 (N156, N135);
xor XOR2 (N157, N150, N53);
not NOT1 (N158, N149);
xor XOR2 (N159, N154, N79);
nor NOR4 (N160, N159, N131, N40, N87);
buf BUF1 (N161, N147);
or OR4 (N162, N153, N108, N38, N77);
xor XOR2 (N163, N155, N92);
not NOT1 (N164, N142);
nor NOR3 (N165, N160, N128, N134);
xor XOR2 (N166, N143, N56);
buf BUF1 (N167, N157);
nand NAND3 (N168, N161, N129, N2);
not NOT1 (N169, N164);
xor XOR2 (N170, N169, N113);
and AND3 (N171, N158, N100, N2);
nor NOR3 (N172, N166, N63, N61);
buf BUF1 (N173, N156);
and AND4 (N174, N162, N53, N126, N86);
buf BUF1 (N175, N172);
buf BUF1 (N176, N163);
or OR2 (N177, N168, N34);
not NOT1 (N178, N174);
buf BUF1 (N179, N178);
nor NOR2 (N180, N152, N150);
xor XOR2 (N181, N170, N134);
not NOT1 (N182, N175);
buf BUF1 (N183, N167);
xor XOR2 (N184, N179, N54);
not NOT1 (N185, N177);
not NOT1 (N186, N185);
not NOT1 (N187, N165);
or OR2 (N188, N176, N24);
xor XOR2 (N189, N183, N68);
not NOT1 (N190, N184);
not NOT1 (N191, N173);
not NOT1 (N192, N189);
nor NOR3 (N193, N191, N165, N190);
nor NOR4 (N194, N117, N187, N105, N14);
not NOT1 (N195, N21);
not NOT1 (N196, N186);
buf BUF1 (N197, N192);
nor NOR2 (N198, N180, N4);
nor NOR2 (N199, N197, N71);
xor XOR2 (N200, N198, N191);
nand NAND4 (N201, N196, N97, N142, N44);
not NOT1 (N202, N171);
or OR3 (N203, N182, N100, N33);
xor XOR2 (N204, N200, N61);
nor NOR3 (N205, N203, N145, N56);
and AND3 (N206, N199, N19, N88);
and AND2 (N207, N204, N31);
nor NOR4 (N208, N206, N40, N36, N57);
and AND3 (N209, N194, N169, N162);
xor XOR2 (N210, N209, N10);
nor NOR3 (N211, N202, N118, N149);
nor NOR3 (N212, N208, N5, N140);
nand NAND4 (N213, N193, N190, N189, N86);
buf BUF1 (N214, N213);
nor NOR3 (N215, N181, N92, N6);
nor NOR3 (N216, N211, N215, N168);
nand NAND4 (N217, N40, N129, N162, N31);
buf BUF1 (N218, N207);
and AND4 (N219, N201, N43, N91, N126);
nor NOR4 (N220, N217, N146, N31, N65);
buf BUF1 (N221, N218);
xor XOR2 (N222, N212, N194);
not NOT1 (N223, N214);
or OR3 (N224, N220, N146, N132);
xor XOR2 (N225, N216, N134);
nand NAND4 (N226, N219, N132, N119, N86);
and AND4 (N227, N226, N133, N72, N154);
xor XOR2 (N228, N195, N212);
nor NOR4 (N229, N221, N2, N153, N87);
buf BUF1 (N230, N227);
xor XOR2 (N231, N223, N192);
buf BUF1 (N232, N225);
buf BUF1 (N233, N232);
xor XOR2 (N234, N233, N27);
not NOT1 (N235, N229);
nor NOR4 (N236, N224, N128, N227, N43);
buf BUF1 (N237, N231);
not NOT1 (N238, N205);
not NOT1 (N239, N228);
not NOT1 (N240, N236);
xor XOR2 (N241, N239, N39);
buf BUF1 (N242, N237);
xor XOR2 (N243, N188, N161);
nand NAND4 (N244, N210, N44, N23, N120);
not NOT1 (N245, N235);
and AND2 (N246, N234, N116);
buf BUF1 (N247, N245);
buf BUF1 (N248, N243);
or OR2 (N249, N244, N21);
nor NOR3 (N250, N238, N236, N86);
nor NOR4 (N251, N250, N133, N165, N167);
nor NOR4 (N252, N249, N167, N27, N234);
nand NAND3 (N253, N230, N69, N190);
or OR3 (N254, N246, N109, N250);
not NOT1 (N255, N254);
nor NOR3 (N256, N252, N22, N133);
nor NOR4 (N257, N248, N36, N238, N97);
nand NAND3 (N258, N241, N161, N225);
and AND2 (N259, N258, N103);
nand NAND4 (N260, N256, N230, N225, N259);
buf BUF1 (N261, N156);
and AND4 (N262, N251, N191, N84, N174);
buf BUF1 (N263, N260);
buf BUF1 (N264, N263);
and AND3 (N265, N240, N98, N27);
buf BUF1 (N266, N253);
buf BUF1 (N267, N242);
xor XOR2 (N268, N266, N169);
or OR4 (N269, N262, N241, N84, N247);
or OR2 (N270, N115, N103);
buf BUF1 (N271, N264);
xor XOR2 (N272, N261, N63);
and AND3 (N273, N268, N234, N53);
not NOT1 (N274, N272);
not NOT1 (N275, N267);
or OR4 (N276, N265, N102, N174, N258);
nand NAND3 (N277, N273, N15, N8);
xor XOR2 (N278, N255, N110);
and AND2 (N279, N276, N8);
and AND2 (N280, N274, N125);
not NOT1 (N281, N257);
not NOT1 (N282, N269);
xor XOR2 (N283, N280, N278);
or OR4 (N284, N162, N255, N145, N18);
or OR2 (N285, N270, N87);
buf BUF1 (N286, N277);
not NOT1 (N287, N222);
nor NOR3 (N288, N282, N77, N70);
buf BUF1 (N289, N283);
xor XOR2 (N290, N287, N208);
not NOT1 (N291, N275);
buf BUF1 (N292, N285);
buf BUF1 (N293, N288);
or OR3 (N294, N293, N37, N259);
not NOT1 (N295, N292);
xor XOR2 (N296, N281, N250);
or OR3 (N297, N294, N280, N22);
and AND4 (N298, N296, N189, N208, N261);
not NOT1 (N299, N279);
buf BUF1 (N300, N286);
nor NOR2 (N301, N298, N14);
not NOT1 (N302, N291);
nor NOR4 (N303, N299, N124, N71, N281);
nor NOR4 (N304, N271, N110, N129, N176);
nor NOR3 (N305, N290, N169, N74);
or OR3 (N306, N289, N296, N24);
or OR2 (N307, N297, N213);
xor XOR2 (N308, N301, N182);
nand NAND4 (N309, N305, N76, N282, N168);
or OR3 (N310, N295, N260, N129);
nand NAND2 (N311, N309, N310);
buf BUF1 (N312, N253);
and AND3 (N313, N306, N234, N18);
buf BUF1 (N314, N303);
and AND2 (N315, N312, N50);
or OR4 (N316, N313, N52, N81, N251);
nand NAND2 (N317, N315, N175);
and AND2 (N318, N317, N228);
xor XOR2 (N319, N284, N153);
not NOT1 (N320, N302);
nor NOR2 (N321, N318, N299);
buf BUF1 (N322, N308);
and AND2 (N323, N322, N137);
buf BUF1 (N324, N311);
not NOT1 (N325, N319);
not NOT1 (N326, N325);
and AND2 (N327, N326, N314);
or OR4 (N328, N91, N319, N102, N57);
or OR3 (N329, N323, N206, N223);
nor NOR2 (N330, N320, N280);
and AND3 (N331, N321, N222, N15);
nand NAND4 (N332, N316, N290, N265, N163);
and AND4 (N333, N329, N41, N217, N137);
xor XOR2 (N334, N328, N112);
nor NOR2 (N335, N304, N139);
and AND4 (N336, N324, N223, N123, N162);
and AND2 (N337, N336, N161);
and AND4 (N338, N333, N118, N6, N141);
and AND3 (N339, N331, N152, N327);
not NOT1 (N340, N77);
nor NOR2 (N341, N334, N42);
nor NOR3 (N342, N340, N17, N86);
nor NOR2 (N343, N330, N239);
xor XOR2 (N344, N337, N261);
nand NAND2 (N345, N307, N185);
nand NAND2 (N346, N300, N189);
and AND3 (N347, N343, N243, N195);
nand NAND3 (N348, N338, N336, N28);
and AND2 (N349, N346, N78);
not NOT1 (N350, N339);
nand NAND2 (N351, N349, N233);
nand NAND4 (N352, N345, N146, N187, N314);
not NOT1 (N353, N344);
or OR4 (N354, N351, N113, N212, N205);
buf BUF1 (N355, N342);
nand NAND2 (N356, N350, N109);
nor NOR3 (N357, N347, N338, N356);
nand NAND3 (N358, N25, N262, N347);
nor NOR2 (N359, N352, N21);
not NOT1 (N360, N359);
not NOT1 (N361, N353);
or OR3 (N362, N332, N39, N313);
xor XOR2 (N363, N335, N70);
xor XOR2 (N364, N362, N32);
and AND2 (N365, N358, N175);
and AND2 (N366, N341, N267);
nand NAND4 (N367, N355, N248, N208, N343);
xor XOR2 (N368, N354, N54);
not NOT1 (N369, N357);
or OR3 (N370, N369, N152, N87);
or OR3 (N371, N368, N65, N176);
not NOT1 (N372, N370);
or OR4 (N373, N363, N219, N318, N108);
or OR3 (N374, N365, N141, N34);
not NOT1 (N375, N373);
nor NOR3 (N376, N348, N20, N78);
xor XOR2 (N377, N375, N294);
or OR2 (N378, N374, N92);
and AND4 (N379, N378, N202, N189, N210);
nor NOR2 (N380, N379, N189);
and AND2 (N381, N371, N196);
or OR4 (N382, N361, N92, N330, N32);
nor NOR2 (N383, N381, N10);
nor NOR2 (N384, N377, N120);
or OR2 (N385, N367, N262);
and AND3 (N386, N372, N164, N241);
not NOT1 (N387, N360);
and AND2 (N388, N383, N328);
or OR2 (N389, N366, N252);
xor XOR2 (N390, N376, N254);
nand NAND3 (N391, N388, N278, N221);
not NOT1 (N392, N389);
or OR4 (N393, N384, N164, N370, N29);
xor XOR2 (N394, N391, N18);
or OR4 (N395, N364, N24, N362, N138);
and AND2 (N396, N395, N236);
or OR2 (N397, N393, N241);
not NOT1 (N398, N392);
nand NAND4 (N399, N397, N2, N29, N192);
xor XOR2 (N400, N386, N302);
nand NAND3 (N401, N390, N294, N194);
or OR3 (N402, N400, N181, N64);
and AND4 (N403, N401, N83, N129, N74);
not NOT1 (N404, N385);
xor XOR2 (N405, N396, N335);
and AND4 (N406, N405, N198, N211, N238);
not NOT1 (N407, N387);
xor XOR2 (N408, N403, N342);
and AND2 (N409, N382, N157);
nor NOR4 (N410, N409, N398, N59, N266);
nand NAND4 (N411, N98, N302, N126, N39);
nor NOR3 (N412, N407, N156, N228);
buf BUF1 (N413, N408);
nand NAND2 (N414, N413, N375);
or OR2 (N415, N402, N303);
nand NAND3 (N416, N406, N380, N122);
and AND3 (N417, N199, N290, N8);
nor NOR2 (N418, N412, N269);
not NOT1 (N419, N399);
nor NOR4 (N420, N418, N134, N340, N35);
and AND2 (N421, N417, N327);
nor NOR4 (N422, N420, N59, N114, N171);
or OR3 (N423, N416, N365, N304);
xor XOR2 (N424, N415, N318);
nand NAND3 (N425, N394, N304, N107);
or OR3 (N426, N414, N67, N4);
and AND3 (N427, N410, N124, N371);
buf BUF1 (N428, N424);
or OR4 (N429, N423, N96, N393, N221);
nand NAND2 (N430, N425, N28);
nand NAND2 (N431, N428, N162);
or OR3 (N432, N431, N341, N260);
nand NAND4 (N433, N429, N418, N221, N264);
not NOT1 (N434, N433);
nand NAND3 (N435, N421, N11, N115);
and AND3 (N436, N422, N369, N7);
nor NOR3 (N437, N404, N227, N394);
not NOT1 (N438, N436);
or OR2 (N439, N419, N300);
buf BUF1 (N440, N426);
and AND2 (N441, N435, N103);
and AND2 (N442, N439, N157);
or OR4 (N443, N411, N374, N108, N286);
nand NAND4 (N444, N432, N196, N423, N267);
nand NAND4 (N445, N440, N224, N297, N271);
nor NOR2 (N446, N443, N325);
nor NOR4 (N447, N430, N335, N175, N405);
xor XOR2 (N448, N437, N97);
nor NOR2 (N449, N442, N48);
xor XOR2 (N450, N444, N68);
or OR3 (N451, N447, N303, N309);
not NOT1 (N452, N451);
nor NOR4 (N453, N448, N36, N114, N380);
not NOT1 (N454, N449);
xor XOR2 (N455, N454, N386);
and AND2 (N456, N455, N307);
or OR2 (N457, N456, N313);
not NOT1 (N458, N452);
or OR3 (N459, N453, N179, N365);
xor XOR2 (N460, N445, N129);
nor NOR4 (N461, N438, N241, N204, N286);
xor XOR2 (N462, N458, N151);
nand NAND2 (N463, N457, N193);
nand NAND2 (N464, N446, N381);
nand NAND2 (N465, N434, N234);
nor NOR3 (N466, N463, N179, N181);
xor XOR2 (N467, N460, N395);
not NOT1 (N468, N461);
nand NAND4 (N469, N468, N385, N190, N122);
and AND3 (N470, N441, N241, N63);
nand NAND3 (N471, N469, N9, N166);
and AND4 (N472, N466, N360, N433, N108);
nor NOR3 (N473, N470, N442, N165);
nor NOR4 (N474, N473, N242, N370, N35);
buf BUF1 (N475, N450);
and AND4 (N476, N475, N35, N276, N402);
or OR4 (N477, N464, N380, N144, N272);
buf BUF1 (N478, N474);
nor NOR3 (N479, N477, N52, N70);
xor XOR2 (N480, N478, N18);
or OR3 (N481, N462, N52, N11);
nand NAND4 (N482, N481, N414, N266, N418);
nor NOR4 (N483, N459, N120, N156, N372);
not NOT1 (N484, N467);
nor NOR2 (N485, N482, N449);
buf BUF1 (N486, N476);
nor NOR2 (N487, N486, N363);
buf BUF1 (N488, N480);
xor XOR2 (N489, N471, N377);
xor XOR2 (N490, N484, N211);
or OR2 (N491, N485, N21);
buf BUF1 (N492, N491);
buf BUF1 (N493, N472);
or OR2 (N494, N483, N128);
xor XOR2 (N495, N465, N394);
not NOT1 (N496, N427);
or OR2 (N497, N495, N138);
not NOT1 (N498, N487);
or OR3 (N499, N492, N1, N431);
not NOT1 (N500, N498);
and AND3 (N501, N499, N309, N495);
or OR2 (N502, N496, N280);
buf BUF1 (N503, N494);
nand NAND2 (N504, N479, N259);
xor XOR2 (N505, N500, N484);
and AND4 (N506, N504, N349, N186, N463);
xor XOR2 (N507, N506, N429);
buf BUF1 (N508, N503);
nor NOR3 (N509, N507, N464, N438);
nor NOR3 (N510, N490, N310, N72);
xor XOR2 (N511, N501, N277);
xor XOR2 (N512, N488, N117);
nor NOR4 (N513, N509, N215, N176, N27);
xor XOR2 (N514, N497, N369);
xor XOR2 (N515, N514, N173);
and AND4 (N516, N512, N510, N22, N210);
or OR3 (N517, N98, N296, N156);
or OR4 (N518, N515, N31, N310, N321);
nor NOR3 (N519, N505, N122, N482);
buf BUF1 (N520, N513);
nand NAND3 (N521, N508, N202, N256);
nor NOR4 (N522, N502, N444, N492, N107);
and AND4 (N523, N516, N370, N173, N278);
and AND2 (N524, N493, N290);
buf BUF1 (N525, N524);
nand NAND2 (N526, N522, N110);
not NOT1 (N527, N511);
nor NOR2 (N528, N523, N166);
and AND3 (N529, N519, N365, N336);
buf BUF1 (N530, N526);
or OR3 (N531, N521, N137, N474);
or OR2 (N532, N489, N235);
and AND2 (N533, N530, N45);
and AND4 (N534, N525, N165, N300, N222);
nand NAND4 (N535, N528, N84, N13, N381);
nand NAND3 (N536, N533, N12, N212);
buf BUF1 (N537, N535);
nor NOR3 (N538, N534, N366, N282);
or OR2 (N539, N538, N147);
not NOT1 (N540, N537);
or OR3 (N541, N518, N115, N146);
not NOT1 (N542, N536);
xor XOR2 (N543, N529, N299);
nor NOR2 (N544, N520, N354);
nor NOR2 (N545, N531, N288);
or OR3 (N546, N544, N539, N129);
or OR3 (N547, N367, N441, N460);
nor NOR4 (N548, N541, N93, N49, N200);
or OR2 (N549, N540, N221);
xor XOR2 (N550, N543, N290);
nor NOR4 (N551, N548, N502, N497, N288);
nand NAND2 (N552, N532, N4);
or OR2 (N553, N549, N244);
nor NOR2 (N554, N527, N519);
and AND4 (N555, N517, N97, N85, N321);
or OR2 (N556, N546, N537);
and AND3 (N557, N554, N451, N228);
and AND3 (N558, N542, N509, N238);
not NOT1 (N559, N551);
buf BUF1 (N560, N550);
nor NOR3 (N561, N555, N280, N521);
and AND3 (N562, N553, N310, N49);
xor XOR2 (N563, N552, N169);
not NOT1 (N564, N560);
nand NAND2 (N565, N562, N5);
xor XOR2 (N566, N557, N391);
or OR3 (N567, N563, N556, N245);
or OR4 (N568, N160, N437, N139, N423);
nor NOR3 (N569, N559, N349, N354);
or OR2 (N570, N561, N192);
buf BUF1 (N571, N565);
and AND3 (N572, N567, N368, N200);
and AND4 (N573, N566, N389, N548, N563);
xor XOR2 (N574, N564, N458);
or OR3 (N575, N571, N491, N529);
nand NAND2 (N576, N572, N429);
nor NOR3 (N577, N569, N412, N15);
xor XOR2 (N578, N574, N292);
nand NAND2 (N579, N573, N368);
nand NAND4 (N580, N576, N570, N115, N124);
nand NAND3 (N581, N192, N105, N461);
or OR3 (N582, N579, N180, N313);
nor NOR3 (N583, N582, N464, N345);
not NOT1 (N584, N583);
buf BUF1 (N585, N584);
or OR3 (N586, N558, N414, N69);
buf BUF1 (N587, N585);
buf BUF1 (N588, N587);
or OR2 (N589, N547, N164);
or OR2 (N590, N577, N433);
nand NAND2 (N591, N589, N92);
buf BUF1 (N592, N590);
nand NAND4 (N593, N575, N77, N100, N6);
not NOT1 (N594, N586);
or OR3 (N595, N588, N271, N38);
buf BUF1 (N596, N593);
not NOT1 (N597, N581);
not NOT1 (N598, N597);
xor XOR2 (N599, N596, N357);
buf BUF1 (N600, N594);
nor NOR2 (N601, N545, N5);
nor NOR2 (N602, N580, N90);
nand NAND3 (N603, N592, N596, N96);
nor NOR3 (N604, N599, N577, N343);
xor XOR2 (N605, N604, N580);
nand NAND3 (N606, N601, N600, N293);
nor NOR4 (N607, N532, N267, N603, N227);
buf BUF1 (N608, N488);
or OR4 (N609, N578, N228, N359, N401);
not NOT1 (N610, N608);
nand NAND4 (N611, N602, N207, N533, N508);
or OR2 (N612, N598, N563);
buf BUF1 (N613, N607);
buf BUF1 (N614, N611);
nor NOR4 (N615, N606, N240, N378, N444);
nand NAND3 (N616, N612, N530, N571);
or OR4 (N617, N609, N190, N613, N237);
or OR3 (N618, N393, N571, N24);
not NOT1 (N619, N615);
not NOT1 (N620, N619);
and AND4 (N621, N618, N26, N255, N497);
nand NAND3 (N622, N620, N249, N81);
and AND3 (N623, N622, N574, N35);
and AND2 (N624, N610, N541);
nor NOR3 (N625, N605, N219, N156);
not NOT1 (N626, N616);
buf BUF1 (N627, N568);
xor XOR2 (N628, N626, N212);
nand NAND3 (N629, N591, N156, N430);
nor NOR3 (N630, N595, N48, N532);
nor NOR3 (N631, N621, N627, N137);
not NOT1 (N632, N550);
nor NOR2 (N633, N624, N311);
and AND4 (N634, N630, N259, N451, N620);
nor NOR3 (N635, N628, N575, N29);
or OR3 (N636, N633, N582, N462);
buf BUF1 (N637, N629);
xor XOR2 (N638, N637, N279);
not NOT1 (N639, N631);
nor NOR4 (N640, N639, N559, N200, N136);
and AND3 (N641, N635, N115, N332);
buf BUF1 (N642, N623);
and AND2 (N643, N642, N510);
or OR2 (N644, N617, N165);
or OR2 (N645, N636, N326);
buf BUF1 (N646, N625);
buf BUF1 (N647, N634);
nand NAND2 (N648, N644, N153);
nand NAND4 (N649, N648, N317, N626, N204);
and AND2 (N650, N649, N619);
buf BUF1 (N651, N647);
nor NOR2 (N652, N643, N586);
xor XOR2 (N653, N638, N502);
not NOT1 (N654, N641);
nand NAND2 (N655, N653, N405);
xor XOR2 (N656, N646, N187);
xor XOR2 (N657, N651, N19);
xor XOR2 (N658, N640, N316);
xor XOR2 (N659, N655, N231);
buf BUF1 (N660, N650);
nor NOR2 (N661, N632, N593);
nand NAND2 (N662, N656, N113);
not NOT1 (N663, N652);
xor XOR2 (N664, N661, N443);
xor XOR2 (N665, N658, N662);
xor XOR2 (N666, N70, N219);
buf BUF1 (N667, N659);
and AND4 (N668, N645, N288, N579, N556);
buf BUF1 (N669, N654);
xor XOR2 (N670, N660, N481);
or OR2 (N671, N664, N218);
xor XOR2 (N672, N668, N415);
xor XOR2 (N673, N671, N651);
and AND2 (N674, N667, N641);
buf BUF1 (N675, N669);
and AND4 (N676, N672, N99, N20, N572);
nor NOR4 (N677, N675, N184, N106, N181);
xor XOR2 (N678, N666, N565);
not NOT1 (N679, N663);
and AND3 (N680, N665, N78, N543);
and AND2 (N681, N678, N613);
and AND3 (N682, N677, N590, N607);
and AND4 (N683, N676, N553, N321, N175);
and AND4 (N684, N679, N227, N503, N492);
buf BUF1 (N685, N681);
xor XOR2 (N686, N614, N211);
or OR2 (N687, N686, N184);
nand NAND4 (N688, N674, N299, N176, N6);
or OR2 (N689, N685, N406);
and AND4 (N690, N673, N591, N455, N450);
xor XOR2 (N691, N687, N404);
and AND2 (N692, N683, N369);
not NOT1 (N693, N657);
nor NOR3 (N694, N682, N455, N90);
buf BUF1 (N695, N692);
xor XOR2 (N696, N694, N302);
buf BUF1 (N697, N695);
xor XOR2 (N698, N684, N406);
nor NOR2 (N699, N680, N427);
not NOT1 (N700, N691);
nand NAND3 (N701, N700, N58, N647);
nor NOR2 (N702, N693, N269);
not NOT1 (N703, N688);
and AND3 (N704, N689, N185, N603);
xor XOR2 (N705, N701, N323);
nor NOR3 (N706, N704, N600, N103);
buf BUF1 (N707, N670);
xor XOR2 (N708, N703, N478);
or OR4 (N709, N699, N457, N544, N49);
nand NAND3 (N710, N709, N638, N217);
not NOT1 (N711, N705);
or OR4 (N712, N698, N402, N687, N271);
and AND3 (N713, N711, N589, N152);
and AND4 (N714, N710, N230, N664, N172);
and AND4 (N715, N696, N199, N208, N303);
and AND4 (N716, N714, N443, N117, N151);
buf BUF1 (N717, N713);
not NOT1 (N718, N716);
or OR4 (N719, N697, N86, N482, N331);
or OR2 (N720, N717, N83);
nor NOR3 (N721, N708, N587, N385);
not NOT1 (N722, N718);
or OR2 (N723, N702, N708);
nand NAND4 (N724, N707, N406, N117, N328);
and AND3 (N725, N720, N228, N456);
or OR2 (N726, N722, N564);
nor NOR3 (N727, N690, N299, N345);
and AND2 (N728, N719, N283);
xor XOR2 (N729, N706, N243);
xor XOR2 (N730, N726, N230);
xor XOR2 (N731, N712, N267);
and AND3 (N732, N724, N338, N272);
not NOT1 (N733, N728);
buf BUF1 (N734, N727);
nand NAND3 (N735, N731, N694, N566);
buf BUF1 (N736, N732);
nor NOR2 (N737, N723, N5);
not NOT1 (N738, N730);
xor XOR2 (N739, N738, N628);
nor NOR4 (N740, N729, N237, N620, N306);
buf BUF1 (N741, N721);
not NOT1 (N742, N739);
nor NOR4 (N743, N734, N627, N141, N712);
and AND4 (N744, N741, N624, N202, N385);
not NOT1 (N745, N740);
xor XOR2 (N746, N745, N430);
not NOT1 (N747, N746);
or OR3 (N748, N737, N687, N159);
buf BUF1 (N749, N735);
or OR2 (N750, N725, N622);
xor XOR2 (N751, N744, N73);
buf BUF1 (N752, N715);
nor NOR2 (N753, N742, N342);
not NOT1 (N754, N733);
and AND3 (N755, N750, N581, N722);
not NOT1 (N756, N747);
nand NAND4 (N757, N753, N81, N537, N199);
nor NOR3 (N758, N752, N175, N623);
or OR2 (N759, N749, N618);
nand NAND3 (N760, N736, N543, N224);
and AND3 (N761, N756, N386, N634);
not NOT1 (N762, N760);
and AND3 (N763, N757, N174, N332);
not NOT1 (N764, N761);
not NOT1 (N765, N759);
nand NAND4 (N766, N765, N49, N17, N303);
nor NOR2 (N767, N758, N101);
nand NAND3 (N768, N754, N540, N262);
xor XOR2 (N769, N767, N57);
xor XOR2 (N770, N766, N132);
xor XOR2 (N771, N748, N97);
buf BUF1 (N772, N771);
and AND3 (N773, N762, N522, N94);
xor XOR2 (N774, N751, N763);
nor NOR4 (N775, N623, N667, N252, N158);
nand NAND2 (N776, N768, N84);
and AND3 (N777, N773, N550, N160);
and AND2 (N778, N743, N60);
and AND3 (N779, N776, N700, N99);
nand NAND2 (N780, N778, N401);
not NOT1 (N781, N777);
nand NAND3 (N782, N764, N448, N698);
buf BUF1 (N783, N779);
xor XOR2 (N784, N775, N106);
nor NOR4 (N785, N755, N592, N740, N583);
nand NAND4 (N786, N770, N673, N22, N132);
nor NOR4 (N787, N786, N650, N78, N428);
xor XOR2 (N788, N781, N272);
buf BUF1 (N789, N772);
nand NAND3 (N790, N774, N378, N123);
nor NOR2 (N791, N769, N658);
not NOT1 (N792, N784);
and AND3 (N793, N790, N731, N760);
xor XOR2 (N794, N793, N699);
and AND2 (N795, N783, N124);
nand NAND2 (N796, N785, N386);
and AND3 (N797, N792, N227, N177);
and AND3 (N798, N796, N14, N528);
not NOT1 (N799, N782);
xor XOR2 (N800, N780, N756);
not NOT1 (N801, N794);
buf BUF1 (N802, N789);
nor NOR2 (N803, N800, N245);
and AND2 (N804, N795, N531);
or OR4 (N805, N802, N591, N727, N432);
nand NAND2 (N806, N797, N171);
xor XOR2 (N807, N787, N729);
or OR2 (N808, N798, N521);
buf BUF1 (N809, N804);
and AND3 (N810, N803, N426, N259);
or OR3 (N811, N791, N498, N692);
and AND2 (N812, N801, N41);
xor XOR2 (N813, N807, N180);
buf BUF1 (N814, N811);
xor XOR2 (N815, N813, N522);
nand NAND2 (N816, N808, N172);
or OR3 (N817, N809, N4, N469);
buf BUF1 (N818, N812);
not NOT1 (N819, N817);
nor NOR3 (N820, N805, N568, N27);
nand NAND2 (N821, N819, N583);
and AND2 (N822, N810, N636);
buf BUF1 (N823, N814);
nor NOR3 (N824, N823, N76, N802);
xor XOR2 (N825, N820, N691);
not NOT1 (N826, N816);
xor XOR2 (N827, N806, N76);
or OR2 (N828, N815, N212);
and AND3 (N829, N799, N305, N189);
buf BUF1 (N830, N821);
nand NAND4 (N831, N827, N692, N375, N643);
buf BUF1 (N832, N831);
and AND4 (N833, N788, N519, N718, N815);
and AND3 (N834, N824, N280, N324);
nor NOR4 (N835, N828, N88, N70, N750);
or OR3 (N836, N818, N550, N321);
nor NOR4 (N837, N835, N5, N124, N17);
xor XOR2 (N838, N832, N372);
not NOT1 (N839, N829);
not NOT1 (N840, N822);
nor NOR4 (N841, N826, N539, N434, N256);
xor XOR2 (N842, N839, N134);
xor XOR2 (N843, N840, N639);
buf BUF1 (N844, N833);
buf BUF1 (N845, N837);
or OR4 (N846, N844, N138, N356, N381);
or OR3 (N847, N830, N42, N808);
buf BUF1 (N848, N845);
or OR2 (N849, N841, N679);
nand NAND4 (N850, N848, N438, N653, N743);
nor NOR4 (N851, N836, N520, N733, N420);
and AND2 (N852, N846, N751);
nand NAND4 (N853, N834, N492, N150, N104);
and AND2 (N854, N847, N553);
nor NOR2 (N855, N843, N649);
or OR2 (N856, N842, N509);
not NOT1 (N857, N854);
nand NAND2 (N858, N850, N409);
nand NAND4 (N859, N853, N378, N588, N222);
nand NAND3 (N860, N858, N350, N244);
not NOT1 (N861, N851);
or OR4 (N862, N860, N675, N723, N22);
buf BUF1 (N863, N852);
nand NAND4 (N864, N862, N134, N149, N293);
not NOT1 (N865, N838);
or OR4 (N866, N857, N504, N527, N84);
or OR4 (N867, N864, N617, N564, N832);
or OR2 (N868, N859, N658);
or OR2 (N869, N861, N178);
and AND3 (N870, N866, N402, N127);
not NOT1 (N871, N825);
nand NAND2 (N872, N865, N755);
buf BUF1 (N873, N870);
or OR4 (N874, N849, N807, N663, N551);
xor XOR2 (N875, N874, N283);
buf BUF1 (N876, N868);
xor XOR2 (N877, N873, N436);
buf BUF1 (N878, N872);
and AND4 (N879, N878, N303, N165, N258);
buf BUF1 (N880, N879);
or OR3 (N881, N856, N47, N818);
not NOT1 (N882, N881);
buf BUF1 (N883, N875);
or OR4 (N884, N863, N219, N222, N222);
nand NAND4 (N885, N883, N367, N559, N325);
and AND2 (N886, N880, N686);
nand NAND2 (N887, N867, N54);
or OR3 (N888, N884, N553, N81);
nand NAND2 (N889, N877, N528);
or OR4 (N890, N886, N827, N669, N633);
not NOT1 (N891, N871);
nand NAND2 (N892, N888, N32);
and AND3 (N893, N876, N767, N66);
nor NOR4 (N894, N892, N264, N492, N765);
xor XOR2 (N895, N890, N573);
xor XOR2 (N896, N869, N520);
not NOT1 (N897, N896);
nand NAND2 (N898, N895, N709);
nand NAND3 (N899, N894, N21, N252);
nand NAND4 (N900, N898, N146, N144, N556);
not NOT1 (N901, N855);
nand NAND2 (N902, N891, N798);
nand NAND2 (N903, N902, N137);
buf BUF1 (N904, N893);
not NOT1 (N905, N887);
not NOT1 (N906, N903);
buf BUF1 (N907, N889);
nor NOR4 (N908, N885, N1, N103, N367);
or OR4 (N909, N899, N780, N828, N843);
or OR3 (N910, N882, N725, N241);
nand NAND3 (N911, N897, N215, N389);
buf BUF1 (N912, N901);
buf BUF1 (N913, N912);
nand NAND2 (N914, N906, N582);
xor XOR2 (N915, N905, N71);
xor XOR2 (N916, N913, N13);
nor NOR4 (N917, N914, N584, N589, N731);
xor XOR2 (N918, N916, N84);
buf BUF1 (N919, N908);
nand NAND2 (N920, N910, N6);
nor NOR4 (N921, N919, N509, N795, N396);
buf BUF1 (N922, N920);
nor NOR3 (N923, N911, N348, N916);
xor XOR2 (N924, N915, N408);
nor NOR4 (N925, N923, N746, N794, N422);
buf BUF1 (N926, N924);
nand NAND4 (N927, N918, N407, N718, N746);
not NOT1 (N928, N927);
not NOT1 (N929, N909);
xor XOR2 (N930, N926, N483);
nor NOR2 (N931, N928, N150);
nand NAND3 (N932, N917, N326, N113);
not NOT1 (N933, N929);
or OR4 (N934, N907, N521, N930, N201);
nand NAND3 (N935, N584, N160, N659);
or OR3 (N936, N931, N762, N188);
nand NAND3 (N937, N936, N654, N93);
nand NAND2 (N938, N937, N178);
or OR4 (N939, N935, N494, N281, N425);
or OR4 (N940, N922, N646, N680, N731);
or OR2 (N941, N904, N505);
not NOT1 (N942, N941);
nand NAND2 (N943, N921, N739);
xor XOR2 (N944, N939, N429);
xor XOR2 (N945, N944, N282);
or OR2 (N946, N938, N712);
and AND2 (N947, N946, N707);
not NOT1 (N948, N900);
and AND2 (N949, N948, N297);
and AND2 (N950, N942, N551);
nor NOR4 (N951, N932, N324, N354, N26);
not NOT1 (N952, N940);
buf BUF1 (N953, N945);
buf BUF1 (N954, N925);
nand NAND3 (N955, N933, N655, N197);
not NOT1 (N956, N955);
or OR2 (N957, N954, N127);
nor NOR4 (N958, N943, N35, N828, N757);
or OR4 (N959, N934, N543, N571, N7);
and AND3 (N960, N953, N287, N136);
buf BUF1 (N961, N952);
nor NOR4 (N962, N947, N577, N229, N726);
or OR4 (N963, N961, N151, N68, N657);
and AND2 (N964, N958, N445);
xor XOR2 (N965, N949, N44);
nor NOR2 (N966, N957, N42);
or OR3 (N967, N963, N393, N872);
nand NAND3 (N968, N960, N190, N622);
buf BUF1 (N969, N951);
nand NAND3 (N970, N966, N738, N668);
or OR3 (N971, N959, N721, N946);
buf BUF1 (N972, N969);
nor NOR4 (N973, N956, N694, N216, N163);
buf BUF1 (N974, N973);
or OR2 (N975, N950, N952);
or OR4 (N976, N968, N267, N278, N554);
buf BUF1 (N977, N976);
xor XOR2 (N978, N967, N619);
not NOT1 (N979, N970);
xor XOR2 (N980, N965, N611);
nand NAND2 (N981, N977, N67);
and AND3 (N982, N971, N11, N57);
xor XOR2 (N983, N974, N88);
and AND4 (N984, N975, N609, N77, N179);
or OR3 (N985, N979, N650, N379);
nand NAND3 (N986, N980, N99, N473);
nor NOR3 (N987, N981, N539, N809);
nor NOR3 (N988, N972, N229, N651);
and AND2 (N989, N983, N741);
nor NOR2 (N990, N986, N974);
nor NOR2 (N991, N982, N143);
and AND3 (N992, N991, N346, N938);
xor XOR2 (N993, N990, N811);
xor XOR2 (N994, N993, N478);
not NOT1 (N995, N964);
or OR2 (N996, N995, N788);
buf BUF1 (N997, N992);
not NOT1 (N998, N984);
xor XOR2 (N999, N987, N420);
buf BUF1 (N1000, N996);
nand NAND4 (N1001, N989, N64, N562, N859);
not NOT1 (N1002, N985);
and AND2 (N1003, N962, N143);
nand NAND2 (N1004, N1003, N311);
not NOT1 (N1005, N1004);
xor XOR2 (N1006, N997, N320);
and AND3 (N1007, N998, N672, N826);
nor NOR3 (N1008, N1007, N925, N558);
buf BUF1 (N1009, N1006);
not NOT1 (N1010, N1000);
nand NAND3 (N1011, N988, N280, N860);
endmodule