// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N211,N212,N188,N209,N210,N195,N205,N206,N200,N213;

or OR2 (N14, N4, N11);
nor NOR4 (N15, N10, N11, N13, N2);
nor NOR3 (N16, N11, N4, N8);
not NOT1 (N17, N8);
buf BUF1 (N18, N11);
not NOT1 (N19, N6);
xor XOR2 (N20, N4, N7);
xor XOR2 (N21, N6, N14);
not NOT1 (N22, N7);
not NOT1 (N23, N19);
and AND4 (N24, N9, N4, N23, N6);
not NOT1 (N25, N21);
and AND3 (N26, N18, N2, N10);
not NOT1 (N27, N21);
nand NAND3 (N28, N19, N3, N9);
or OR3 (N29, N15, N6, N20);
nand NAND2 (N30, N4, N14);
or OR2 (N31, N16, N1);
buf BUF1 (N32, N29);
not NOT1 (N33, N28);
nor NOR2 (N34, N24, N31);
not NOT1 (N35, N30);
buf BUF1 (N36, N35);
nor NOR4 (N37, N4, N6, N31, N16);
xor XOR2 (N38, N33, N12);
or OR3 (N39, N17, N11, N20);
xor XOR2 (N40, N38, N11);
buf BUF1 (N41, N26);
nand NAND3 (N42, N41, N6, N38);
and AND4 (N43, N37, N23, N28, N40);
xor XOR2 (N44, N19, N18);
not NOT1 (N45, N34);
nor NOR4 (N46, N36, N11, N37, N22);
xor XOR2 (N47, N1, N28);
or OR3 (N48, N27, N5, N33);
or OR2 (N49, N46, N29);
xor XOR2 (N50, N47, N14);
nor NOR3 (N51, N42, N50, N10);
nor NOR2 (N52, N3, N28);
buf BUF1 (N53, N45);
or OR2 (N54, N51, N23);
and AND3 (N55, N39, N30, N18);
or OR4 (N56, N55, N34, N46, N50);
not NOT1 (N57, N53);
xor XOR2 (N58, N56, N10);
nand NAND4 (N59, N43, N9, N1, N44);
buf BUF1 (N60, N3);
or OR4 (N61, N52, N33, N41, N54);
nand NAND2 (N62, N12, N2);
nor NOR4 (N63, N59, N59, N51, N30);
and AND2 (N64, N48, N60);
nand NAND3 (N65, N61, N59, N51);
not NOT1 (N66, N47);
and AND4 (N67, N64, N43, N28, N4);
nor NOR4 (N68, N66, N27, N54, N3);
nand NAND2 (N69, N67, N66);
nor NOR4 (N70, N62, N40, N65, N4);
or OR3 (N71, N66, N38, N31);
or OR3 (N72, N58, N12, N36);
or OR3 (N73, N25, N70, N16);
xor XOR2 (N74, N68, N37);
xor XOR2 (N75, N61, N59);
buf BUF1 (N76, N49);
nor NOR4 (N77, N75, N71, N50, N33);
nand NAND4 (N78, N75, N27, N25, N1);
not NOT1 (N79, N32);
buf BUF1 (N80, N63);
nor NOR2 (N81, N74, N24);
nor NOR4 (N82, N78, N29, N78, N42);
or OR4 (N83, N73, N71, N13, N32);
or OR3 (N84, N81, N52, N11);
nor NOR2 (N85, N84, N56);
and AND4 (N86, N79, N73, N62, N65);
and AND2 (N87, N77, N72);
nand NAND3 (N88, N55, N84, N11);
xor XOR2 (N89, N57, N53);
xor XOR2 (N90, N87, N36);
not NOT1 (N91, N90);
nor NOR2 (N92, N91, N51);
and AND3 (N93, N83, N39, N44);
nand NAND2 (N94, N89, N40);
not NOT1 (N95, N85);
or OR2 (N96, N82, N73);
not NOT1 (N97, N92);
buf BUF1 (N98, N86);
not NOT1 (N99, N76);
and AND3 (N100, N80, N67, N40);
nor NOR2 (N101, N98, N91);
xor XOR2 (N102, N88, N74);
not NOT1 (N103, N96);
xor XOR2 (N104, N103, N42);
nor NOR4 (N105, N95, N92, N54, N19);
and AND3 (N106, N104, N83, N68);
and AND4 (N107, N106, N46, N74, N77);
or OR2 (N108, N107, N78);
nand NAND4 (N109, N69, N107, N60, N85);
nand NAND2 (N110, N108, N8);
nor NOR3 (N111, N94, N85, N81);
xor XOR2 (N112, N111, N56);
or OR3 (N113, N102, N15, N15);
xor XOR2 (N114, N97, N80);
xor XOR2 (N115, N112, N112);
and AND3 (N116, N99, N106, N84);
xor XOR2 (N117, N110, N73);
nor NOR3 (N118, N117, N48, N93);
nand NAND2 (N119, N28, N80);
nor NOR2 (N120, N114, N64);
nor NOR2 (N121, N113, N24);
or OR4 (N122, N119, N116, N103, N49);
or OR4 (N123, N7, N40, N35, N39);
nor NOR2 (N124, N115, N117);
not NOT1 (N125, N118);
xor XOR2 (N126, N122, N24);
xor XOR2 (N127, N109, N17);
nor NOR2 (N128, N125, N11);
nand NAND3 (N129, N128, N34, N124);
buf BUF1 (N130, N97);
nor NOR3 (N131, N126, N43, N77);
or OR3 (N132, N131, N34, N70);
buf BUF1 (N133, N129);
xor XOR2 (N134, N100, N50);
and AND2 (N135, N130, N90);
and AND3 (N136, N121, N57, N123);
and AND3 (N137, N70, N18, N49);
buf BUF1 (N138, N105);
buf BUF1 (N139, N127);
nor NOR2 (N140, N136, N58);
buf BUF1 (N141, N132);
and AND2 (N142, N135, N96);
and AND2 (N143, N138, N103);
xor XOR2 (N144, N137, N104);
xor XOR2 (N145, N133, N132);
nor NOR2 (N146, N141, N92);
or OR3 (N147, N134, N140, N77);
xor XOR2 (N148, N14, N48);
or OR3 (N149, N146, N36, N66);
xor XOR2 (N150, N139, N95);
buf BUF1 (N151, N149);
nor NOR4 (N152, N150, N6, N109, N20);
nand NAND3 (N153, N120, N123, N15);
not NOT1 (N154, N152);
not NOT1 (N155, N154);
or OR2 (N156, N101, N121);
not NOT1 (N157, N144);
xor XOR2 (N158, N147, N126);
buf BUF1 (N159, N155);
or OR3 (N160, N145, N20, N92);
and AND3 (N161, N148, N26, N78);
nand NAND4 (N162, N142, N31, N129, N34);
buf BUF1 (N163, N158);
and AND2 (N164, N151, N13);
nor NOR4 (N165, N153, N101, N54, N22);
or OR3 (N166, N162, N112, N32);
buf BUF1 (N167, N143);
buf BUF1 (N168, N164);
buf BUF1 (N169, N159);
and AND4 (N170, N165, N69, N64, N38);
xor XOR2 (N171, N160, N140);
nor NOR3 (N172, N170, N9, N157);
and AND4 (N173, N60, N151, N23, N68);
or OR3 (N174, N168, N137, N58);
and AND2 (N175, N156, N107);
not NOT1 (N176, N161);
and AND2 (N177, N163, N158);
nand NAND4 (N178, N175, N83, N8, N33);
and AND3 (N179, N174, N57, N5);
not NOT1 (N180, N166);
not NOT1 (N181, N169);
or OR4 (N182, N177, N40, N168, N130);
xor XOR2 (N183, N173, N115);
xor XOR2 (N184, N183, N87);
and AND3 (N185, N167, N86, N8);
xor XOR2 (N186, N178, N148);
buf BUF1 (N187, N179);
nand NAND2 (N188, N186, N35);
and AND3 (N189, N182, N103, N73);
not NOT1 (N190, N180);
or OR2 (N191, N176, N118);
buf BUF1 (N192, N181);
or OR3 (N193, N187, N64, N185);
or OR4 (N194, N122, N68, N48, N85);
nor NOR3 (N195, N184, N152, N140);
xor XOR2 (N196, N194, N118);
and AND4 (N197, N189, N19, N26, N141);
and AND2 (N198, N197, N116);
nor NOR3 (N199, N190, N140, N172);
nor NOR4 (N200, N27, N194, N10, N133);
buf BUF1 (N201, N198);
and AND3 (N202, N199, N11, N177);
buf BUF1 (N203, N192);
buf BUF1 (N204, N191);
xor XOR2 (N205, N201, N5);
xor XOR2 (N206, N196, N179);
nor NOR2 (N207, N203, N141);
xor XOR2 (N208, N204, N17);
nand NAND4 (N209, N193, N187, N60, N108);
nor NOR4 (N210, N207, N26, N12, N51);
buf BUF1 (N211, N208);
nor NOR4 (N212, N202, N42, N126, N23);
and AND2 (N213, N171, N116);
endmodule