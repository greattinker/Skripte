// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N601,N609,N610,N581,N599,N598,N586,N608,N612;

buf BUF1 (N13, N11);
xor XOR2 (N14, N7, N11);
not NOT1 (N15, N13);
buf BUF1 (N16, N7);
not NOT1 (N17, N4);
nand NAND3 (N18, N6, N6, N14);
not NOT1 (N19, N1);
nor NOR3 (N20, N19, N1, N19);
buf BUF1 (N21, N20);
nand NAND2 (N22, N10, N13);
not NOT1 (N23, N14);
and AND2 (N24, N1, N19);
buf BUF1 (N25, N19);
nor NOR3 (N26, N20, N16, N16);
not NOT1 (N27, N1);
and AND3 (N28, N26, N22, N8);
buf BUF1 (N29, N10);
buf BUF1 (N30, N21);
not NOT1 (N31, N24);
nor NOR3 (N32, N28, N8, N15);
and AND2 (N33, N13, N21);
nor NOR2 (N34, N25, N19);
xor XOR2 (N35, N29, N28);
nand NAND2 (N36, N35, N11);
or OR2 (N37, N31, N3);
buf BUF1 (N38, N37);
nor NOR2 (N39, N34, N31);
or OR2 (N40, N38, N37);
and AND3 (N41, N36, N36, N16);
or OR3 (N42, N27, N17, N10);
nor NOR3 (N43, N38, N7, N17);
xor XOR2 (N44, N43, N12);
xor XOR2 (N45, N18, N31);
not NOT1 (N46, N41);
and AND4 (N47, N33, N30, N19, N6);
nand NAND2 (N48, N12, N39);
or OR2 (N49, N16, N5);
xor XOR2 (N50, N48, N7);
xor XOR2 (N51, N46, N35);
or OR2 (N52, N47, N5);
nor NOR4 (N53, N45, N29, N30, N34);
or OR2 (N54, N52, N5);
not NOT1 (N55, N49);
xor XOR2 (N56, N44, N46);
and AND2 (N57, N51, N48);
not NOT1 (N58, N55);
or OR2 (N59, N42, N57);
not NOT1 (N60, N51);
xor XOR2 (N61, N23, N9);
buf BUF1 (N62, N53);
buf BUF1 (N63, N32);
and AND4 (N64, N58, N45, N3, N38);
xor XOR2 (N65, N62, N22);
nor NOR3 (N66, N59, N1, N51);
xor XOR2 (N67, N56, N53);
buf BUF1 (N68, N61);
and AND3 (N69, N63, N33, N45);
not NOT1 (N70, N66);
nand NAND2 (N71, N65, N69);
and AND3 (N72, N68, N1, N30);
not NOT1 (N73, N45);
or OR4 (N74, N71, N45, N12, N59);
buf BUF1 (N75, N54);
or OR2 (N76, N75, N47);
or OR4 (N77, N74, N36, N23, N49);
nand NAND3 (N78, N60, N13, N43);
buf BUF1 (N79, N50);
nor NOR3 (N80, N40, N57, N32);
buf BUF1 (N81, N76);
or OR2 (N82, N78, N54);
not NOT1 (N83, N73);
or OR4 (N84, N72, N51, N69, N23);
buf BUF1 (N85, N77);
or OR3 (N86, N81, N66, N83);
not NOT1 (N87, N15);
nor NOR4 (N88, N84, N22, N65, N19);
nand NAND2 (N89, N82, N12);
or OR3 (N90, N79, N52, N24);
buf BUF1 (N91, N67);
buf BUF1 (N92, N89);
or OR3 (N93, N80, N30, N77);
nand NAND3 (N94, N88, N87, N46);
and AND4 (N95, N42, N93, N27, N70);
xor XOR2 (N96, N27, N6);
buf BUF1 (N97, N91);
and AND4 (N98, N5, N27, N80, N78);
and AND4 (N99, N92, N51, N96, N67);
buf BUF1 (N100, N5);
or OR4 (N101, N95, N5, N36, N64);
xor XOR2 (N102, N96, N97);
xor XOR2 (N103, N90, N54);
and AND2 (N104, N38, N53);
buf BUF1 (N105, N102);
buf BUF1 (N106, N105);
xor XOR2 (N107, N85, N45);
or OR2 (N108, N99, N51);
not NOT1 (N109, N104);
buf BUF1 (N110, N106);
or OR2 (N111, N108, N22);
nor NOR4 (N112, N98, N82, N92, N89);
and AND4 (N113, N110, N60, N23, N80);
and AND2 (N114, N107, N36);
buf BUF1 (N115, N112);
and AND2 (N116, N94, N18);
or OR3 (N117, N109, N77, N101);
not NOT1 (N118, N3);
nand NAND4 (N119, N113, N81, N62, N52);
nand NAND2 (N120, N115, N35);
or OR2 (N121, N114, N72);
or OR3 (N122, N86, N43, N94);
nor NOR2 (N123, N117, N65);
and AND2 (N124, N121, N37);
or OR4 (N125, N118, N114, N98, N66);
not NOT1 (N126, N111);
nor NOR3 (N127, N120, N34, N4);
not NOT1 (N128, N126);
xor XOR2 (N129, N125, N60);
or OR4 (N130, N127, N127, N7, N54);
nor NOR2 (N131, N116, N127);
nand NAND3 (N132, N131, N7, N120);
nor NOR3 (N133, N130, N109, N113);
xor XOR2 (N134, N123, N62);
nand NAND4 (N135, N124, N40, N54, N32);
not NOT1 (N136, N128);
and AND2 (N137, N129, N105);
and AND2 (N138, N132, N6);
or OR2 (N139, N134, N38);
or OR4 (N140, N119, N42, N54, N65);
or OR2 (N141, N122, N65);
nor NOR3 (N142, N103, N13, N61);
nand NAND4 (N143, N133, N101, N48, N126);
and AND2 (N144, N140, N121);
nand NAND4 (N145, N135, N35, N94, N25);
xor XOR2 (N146, N100, N12);
and AND4 (N147, N136, N79, N81, N12);
buf BUF1 (N148, N143);
buf BUF1 (N149, N145);
xor XOR2 (N150, N141, N124);
and AND2 (N151, N148, N28);
or OR2 (N152, N151, N54);
buf BUF1 (N153, N150);
nand NAND3 (N154, N138, N120, N61);
not NOT1 (N155, N142);
nor NOR4 (N156, N146, N23, N119, N23);
buf BUF1 (N157, N155);
not NOT1 (N158, N153);
and AND3 (N159, N147, N109, N156);
and AND3 (N160, N105, N44, N70);
nor NOR2 (N161, N159, N31);
xor XOR2 (N162, N161, N97);
xor XOR2 (N163, N149, N122);
or OR3 (N164, N158, N81, N101);
or OR4 (N165, N162, N19, N65, N42);
nor NOR4 (N166, N163, N24, N84, N1);
not NOT1 (N167, N139);
nor NOR4 (N168, N164, N140, N102, N53);
buf BUF1 (N169, N168);
nand NAND2 (N170, N160, N166);
or OR3 (N171, N44, N29, N51);
nand NAND2 (N172, N157, N32);
not NOT1 (N173, N169);
buf BUF1 (N174, N154);
buf BUF1 (N175, N170);
xor XOR2 (N176, N167, N5);
and AND3 (N177, N137, N94, N25);
and AND3 (N178, N165, N118, N146);
and AND2 (N179, N144, N121);
not NOT1 (N180, N175);
nor NOR4 (N181, N180, N135, N55, N71);
or OR2 (N182, N152, N8);
and AND3 (N183, N182, N59, N123);
or OR4 (N184, N176, N38, N10, N116);
nand NAND4 (N185, N174, N140, N143, N151);
not NOT1 (N186, N177);
not NOT1 (N187, N178);
not NOT1 (N188, N184);
xor XOR2 (N189, N186, N62);
nor NOR2 (N190, N185, N41);
or OR3 (N191, N183, N64, N106);
nor NOR2 (N192, N191, N58);
buf BUF1 (N193, N189);
or OR2 (N194, N179, N110);
or OR3 (N195, N190, N184, N41);
nand NAND4 (N196, N171, N14, N188, N10);
buf BUF1 (N197, N54);
buf BUF1 (N198, N181);
nand NAND4 (N199, N197, N140, N54, N185);
nor NOR4 (N200, N199, N115, N108, N44);
nand NAND2 (N201, N196, N14);
or OR2 (N202, N172, N2);
buf BUF1 (N203, N200);
nand NAND3 (N204, N203, N80, N65);
nor NOR3 (N205, N187, N178, N57);
or OR3 (N206, N195, N34, N79);
or OR3 (N207, N205, N195, N111);
not NOT1 (N208, N198);
not NOT1 (N209, N194);
xor XOR2 (N210, N208, N42);
xor XOR2 (N211, N206, N184);
and AND2 (N212, N202, N157);
not NOT1 (N213, N201);
and AND4 (N214, N210, N92, N106, N195);
not NOT1 (N215, N211);
xor XOR2 (N216, N209, N151);
nand NAND2 (N217, N214, N65);
or OR4 (N218, N173, N78, N3, N35);
and AND4 (N219, N204, N89, N75, N112);
xor XOR2 (N220, N215, N16);
xor XOR2 (N221, N219, N91);
nor NOR2 (N222, N212, N23);
nor NOR4 (N223, N217, N190, N133, N205);
buf BUF1 (N224, N221);
not NOT1 (N225, N207);
buf BUF1 (N226, N192);
xor XOR2 (N227, N225, N95);
nand NAND2 (N228, N223, N27);
xor XOR2 (N229, N226, N152);
nor NOR2 (N230, N224, N212);
xor XOR2 (N231, N216, N56);
nand NAND4 (N232, N228, N144, N134, N31);
xor XOR2 (N233, N231, N47);
buf BUF1 (N234, N227);
buf BUF1 (N235, N218);
not NOT1 (N236, N229);
or OR2 (N237, N233, N151);
not NOT1 (N238, N232);
and AND2 (N239, N235, N49);
not NOT1 (N240, N237);
xor XOR2 (N241, N213, N199);
not NOT1 (N242, N239);
nand NAND3 (N243, N193, N137, N177);
not NOT1 (N244, N234);
buf BUF1 (N245, N241);
not NOT1 (N246, N240);
nand NAND4 (N247, N230, N155, N112, N63);
nor NOR4 (N248, N242, N201, N82, N123);
xor XOR2 (N249, N243, N122);
not NOT1 (N250, N244);
and AND4 (N251, N245, N233, N162, N218);
or OR4 (N252, N220, N201, N77, N156);
and AND2 (N253, N246, N154);
xor XOR2 (N254, N238, N204);
nor NOR3 (N255, N247, N242, N107);
and AND2 (N256, N248, N38);
nand NAND2 (N257, N222, N234);
not NOT1 (N258, N253);
nand NAND2 (N259, N255, N159);
not NOT1 (N260, N256);
or OR2 (N261, N249, N13);
xor XOR2 (N262, N250, N205);
buf BUF1 (N263, N254);
buf BUF1 (N264, N257);
and AND3 (N265, N260, N141, N26);
nand NAND4 (N266, N264, N3, N59, N42);
or OR3 (N267, N265, N113, N60);
xor XOR2 (N268, N262, N213);
and AND4 (N269, N267, N249, N3, N211);
and AND3 (N270, N266, N2, N236);
nand NAND4 (N271, N98, N45, N68, N238);
xor XOR2 (N272, N268, N166);
or OR4 (N273, N271, N37, N6, N118);
not NOT1 (N274, N259);
and AND3 (N275, N272, N250, N162);
and AND3 (N276, N270, N157, N19);
buf BUF1 (N277, N251);
and AND2 (N278, N269, N56);
nand NAND3 (N279, N261, N48, N156);
and AND3 (N280, N263, N147, N55);
and AND4 (N281, N274, N232, N216, N272);
or OR4 (N282, N276, N276, N275, N35);
nand NAND4 (N283, N45, N129, N23, N100);
nand NAND3 (N284, N252, N62, N178);
nand NAND3 (N285, N284, N58, N38);
or OR4 (N286, N277, N61, N36, N68);
and AND4 (N287, N280, N231, N223, N13);
nand NAND3 (N288, N258, N168, N233);
not NOT1 (N289, N288);
or OR3 (N290, N285, N53, N213);
and AND2 (N291, N281, N173);
not NOT1 (N292, N279);
nand NAND3 (N293, N283, N136, N34);
nand NAND3 (N294, N282, N275, N37);
buf BUF1 (N295, N293);
and AND2 (N296, N286, N136);
not NOT1 (N297, N291);
xor XOR2 (N298, N290, N43);
and AND4 (N299, N289, N192, N165, N126);
and AND3 (N300, N296, N201, N236);
and AND3 (N301, N287, N204, N151);
nand NAND4 (N302, N294, N147, N45, N137);
xor XOR2 (N303, N295, N72);
and AND2 (N304, N278, N151);
nor NOR2 (N305, N292, N142);
not NOT1 (N306, N305);
or OR4 (N307, N306, N144, N32, N272);
and AND4 (N308, N297, N26, N8, N94);
xor XOR2 (N309, N303, N117);
or OR4 (N310, N309, N239, N52, N48);
and AND4 (N311, N307, N162, N194, N302);
nor NOR3 (N312, N227, N29, N99);
xor XOR2 (N313, N301, N91);
buf BUF1 (N314, N308);
or OR2 (N315, N314, N227);
nor NOR4 (N316, N311, N200, N168, N308);
buf BUF1 (N317, N310);
not NOT1 (N318, N317);
or OR2 (N319, N318, N7);
nand NAND2 (N320, N316, N304);
not NOT1 (N321, N111);
not NOT1 (N322, N319);
nand NAND4 (N323, N312, N211, N118, N93);
not NOT1 (N324, N300);
not NOT1 (N325, N323);
nand NAND3 (N326, N313, N52, N239);
or OR2 (N327, N299, N140);
nand NAND4 (N328, N273, N150, N325, N320);
and AND2 (N329, N214, N118);
nand NAND4 (N330, N90, N236, N146, N301);
or OR3 (N331, N322, N5, N186);
not NOT1 (N332, N326);
nor NOR3 (N333, N331, N77, N267);
or OR3 (N334, N333, N93, N224);
and AND2 (N335, N324, N170);
not NOT1 (N336, N330);
or OR3 (N337, N298, N13, N268);
nand NAND4 (N338, N321, N240, N32, N176);
and AND3 (N339, N336, N66, N146);
not NOT1 (N340, N339);
xor XOR2 (N341, N338, N319);
not NOT1 (N342, N315);
buf BUF1 (N343, N332);
nand NAND4 (N344, N327, N206, N106, N117);
or OR3 (N345, N337, N232, N270);
xor XOR2 (N346, N342, N41);
or OR3 (N347, N346, N164, N73);
not NOT1 (N348, N334);
nand NAND3 (N349, N348, N301, N198);
buf BUF1 (N350, N341);
or OR3 (N351, N335, N178, N227);
or OR2 (N352, N350, N80);
nor NOR3 (N353, N349, N16, N299);
nor NOR2 (N354, N344, N334);
or OR4 (N355, N354, N138, N342, N198);
and AND3 (N356, N353, N108, N76);
buf BUF1 (N357, N355);
not NOT1 (N358, N329);
buf BUF1 (N359, N356);
not NOT1 (N360, N347);
or OR3 (N361, N357, N282, N197);
xor XOR2 (N362, N351, N291);
or OR3 (N363, N343, N280, N144);
or OR3 (N364, N340, N350, N217);
or OR3 (N365, N359, N73, N194);
or OR2 (N366, N352, N38);
or OR2 (N367, N365, N359);
not NOT1 (N368, N364);
and AND2 (N369, N358, N251);
nand NAND3 (N370, N367, N36, N90);
xor XOR2 (N371, N369, N355);
xor XOR2 (N372, N370, N364);
nand NAND3 (N373, N361, N330, N3);
or OR2 (N374, N360, N287);
xor XOR2 (N375, N374, N195);
or OR3 (N376, N368, N6, N354);
buf BUF1 (N377, N371);
or OR3 (N378, N363, N222, N132);
or OR3 (N379, N372, N321, N288);
nand NAND3 (N380, N376, N306, N11);
or OR3 (N381, N380, N6, N163);
nand NAND4 (N382, N373, N264, N40, N117);
nor NOR4 (N383, N378, N279, N298, N357);
and AND2 (N384, N382, N299);
and AND4 (N385, N383, N364, N372, N275);
or OR3 (N386, N384, N10, N41);
nand NAND3 (N387, N366, N65, N270);
xor XOR2 (N388, N328, N142);
or OR2 (N389, N362, N326);
nor NOR2 (N390, N381, N62);
and AND2 (N391, N389, N94);
buf BUF1 (N392, N391);
nor NOR3 (N393, N385, N194, N363);
and AND2 (N394, N375, N224);
not NOT1 (N395, N388);
not NOT1 (N396, N379);
or OR4 (N397, N390, N365, N72, N93);
not NOT1 (N398, N397);
nor NOR3 (N399, N394, N30, N336);
not NOT1 (N400, N345);
buf BUF1 (N401, N377);
xor XOR2 (N402, N395, N27);
or OR4 (N403, N396, N313, N223, N257);
and AND2 (N404, N387, N202);
or OR3 (N405, N399, N81, N388);
or OR2 (N406, N400, N243);
nor NOR3 (N407, N386, N144, N99);
xor XOR2 (N408, N401, N5);
and AND3 (N409, N405, N212, N406);
buf BUF1 (N410, N91);
and AND3 (N411, N408, N208, N290);
buf BUF1 (N412, N398);
and AND2 (N413, N410, N378);
not NOT1 (N414, N392);
xor XOR2 (N415, N403, N329);
nand NAND3 (N416, N414, N89, N78);
xor XOR2 (N417, N407, N302);
buf BUF1 (N418, N409);
nand NAND3 (N419, N402, N112, N45);
and AND3 (N420, N415, N349, N90);
not NOT1 (N421, N411);
buf BUF1 (N422, N419);
and AND4 (N423, N422, N262, N276, N225);
not NOT1 (N424, N421);
xor XOR2 (N425, N423, N319);
nor NOR4 (N426, N413, N151, N62, N337);
nor NOR2 (N427, N416, N351);
or OR4 (N428, N393, N231, N154, N93);
or OR2 (N429, N427, N133);
buf BUF1 (N430, N425);
xor XOR2 (N431, N420, N7);
nor NOR4 (N432, N428, N240, N263, N201);
not NOT1 (N433, N431);
or OR2 (N434, N424, N159);
xor XOR2 (N435, N434, N386);
nand NAND2 (N436, N435, N240);
xor XOR2 (N437, N418, N408);
xor XOR2 (N438, N429, N302);
not NOT1 (N439, N426);
xor XOR2 (N440, N438, N376);
not NOT1 (N441, N404);
buf BUF1 (N442, N441);
buf BUF1 (N443, N433);
or OR4 (N444, N432, N427, N217, N180);
nand NAND3 (N445, N440, N367, N19);
nor NOR2 (N446, N443, N123);
xor XOR2 (N447, N437, N327);
buf BUF1 (N448, N445);
not NOT1 (N449, N436);
not NOT1 (N450, N442);
buf BUF1 (N451, N448);
or OR3 (N452, N450, N15, N65);
not NOT1 (N453, N417);
and AND3 (N454, N451, N193, N264);
nand NAND3 (N455, N444, N381, N327);
nand NAND4 (N456, N452, N236, N245, N90);
nand NAND4 (N457, N456, N19, N47, N38);
nand NAND3 (N458, N446, N245, N298);
not NOT1 (N459, N453);
and AND4 (N460, N457, N43, N262, N424);
nand NAND2 (N461, N455, N173);
not NOT1 (N462, N412);
buf BUF1 (N463, N454);
or OR4 (N464, N463, N18, N172, N415);
xor XOR2 (N465, N460, N151);
nor NOR4 (N466, N464, N231, N436, N32);
and AND2 (N467, N458, N300);
or OR3 (N468, N459, N308, N440);
nor NOR2 (N469, N439, N206);
buf BUF1 (N470, N468);
buf BUF1 (N471, N449);
xor XOR2 (N472, N469, N357);
xor XOR2 (N473, N466, N53);
not NOT1 (N474, N462);
nor NOR3 (N475, N430, N121, N34);
buf BUF1 (N476, N473);
buf BUF1 (N477, N447);
xor XOR2 (N478, N472, N390);
buf BUF1 (N479, N470);
not NOT1 (N480, N471);
not NOT1 (N481, N477);
nor NOR4 (N482, N475, N49, N445, N456);
and AND2 (N483, N482, N164);
or OR4 (N484, N461, N317, N77, N427);
buf BUF1 (N485, N478);
not NOT1 (N486, N467);
nor NOR2 (N487, N485, N238);
nor NOR2 (N488, N481, N208);
not NOT1 (N489, N483);
nor NOR2 (N490, N474, N347);
nor NOR2 (N491, N479, N476);
nand NAND3 (N492, N11, N121, N430);
or OR4 (N493, N491, N398, N335, N249);
xor XOR2 (N494, N484, N95);
or OR3 (N495, N487, N16, N182);
buf BUF1 (N496, N489);
and AND3 (N497, N490, N169, N134);
buf BUF1 (N498, N480);
nor NOR3 (N499, N486, N130, N454);
or OR4 (N500, N465, N103, N84, N83);
buf BUF1 (N501, N500);
buf BUF1 (N502, N499);
or OR3 (N503, N494, N94, N257);
or OR2 (N504, N492, N450);
xor XOR2 (N505, N497, N271);
buf BUF1 (N506, N493);
not NOT1 (N507, N506);
not NOT1 (N508, N505);
not NOT1 (N509, N503);
buf BUF1 (N510, N496);
not NOT1 (N511, N488);
buf BUF1 (N512, N498);
buf BUF1 (N513, N510);
nand NAND2 (N514, N504, N149);
nor NOR2 (N515, N495, N193);
or OR3 (N516, N515, N52, N495);
buf BUF1 (N517, N511);
xor XOR2 (N518, N509, N70);
not NOT1 (N519, N512);
buf BUF1 (N520, N514);
not NOT1 (N521, N501);
buf BUF1 (N522, N521);
not NOT1 (N523, N508);
buf BUF1 (N524, N518);
not NOT1 (N525, N516);
buf BUF1 (N526, N502);
and AND2 (N527, N523, N154);
buf BUF1 (N528, N513);
buf BUF1 (N529, N522);
buf BUF1 (N530, N529);
nand NAND4 (N531, N520, N465, N96, N320);
buf BUF1 (N532, N526);
buf BUF1 (N533, N519);
nor NOR3 (N534, N525, N454, N323);
not NOT1 (N535, N528);
nor NOR3 (N536, N531, N353, N119);
and AND2 (N537, N535, N80);
nor NOR4 (N538, N517, N179, N214, N13);
and AND3 (N539, N533, N164, N226);
xor XOR2 (N540, N507, N220);
xor XOR2 (N541, N534, N133);
xor XOR2 (N542, N530, N457);
nand NAND2 (N543, N541, N64);
and AND3 (N544, N542, N274, N387);
nand NAND4 (N545, N524, N328, N357, N469);
buf BUF1 (N546, N527);
not NOT1 (N547, N539);
nor NOR4 (N548, N546, N179, N284, N404);
nor NOR2 (N549, N543, N297);
not NOT1 (N550, N548);
nand NAND2 (N551, N550, N545);
xor XOR2 (N552, N396, N427);
or OR2 (N553, N540, N514);
nor NOR2 (N554, N551, N15);
not NOT1 (N555, N537);
xor XOR2 (N556, N538, N380);
nor NOR4 (N557, N532, N503, N321, N371);
nand NAND4 (N558, N552, N118, N16, N178);
nand NAND4 (N559, N556, N53, N211, N356);
xor XOR2 (N560, N549, N317);
nand NAND4 (N561, N553, N224, N523, N481);
xor XOR2 (N562, N547, N228);
not NOT1 (N563, N544);
not NOT1 (N564, N560);
nor NOR2 (N565, N555, N272);
xor XOR2 (N566, N558, N546);
nor NOR3 (N567, N559, N232, N381);
and AND3 (N568, N562, N552, N177);
nor NOR4 (N569, N565, N548, N563, N231);
buf BUF1 (N570, N552);
and AND3 (N571, N536, N204, N73);
nand NAND4 (N572, N571, N512, N139, N124);
or OR3 (N573, N568, N387, N403);
and AND3 (N574, N554, N197, N15);
not NOT1 (N575, N561);
or OR4 (N576, N567, N501, N190, N496);
nor NOR4 (N577, N575, N95, N442, N104);
or OR2 (N578, N557, N549);
not NOT1 (N579, N573);
and AND3 (N580, N574, N343, N558);
not NOT1 (N581, N578);
buf BUF1 (N582, N577);
or OR3 (N583, N572, N570, N143);
or OR4 (N584, N215, N221, N244, N221);
not NOT1 (N585, N569);
xor XOR2 (N586, N585, N241);
nor NOR4 (N587, N584, N110, N269, N577);
or OR3 (N588, N582, N18, N146);
and AND2 (N589, N583, N222);
not NOT1 (N590, N579);
and AND4 (N591, N564, N109, N455, N188);
nor NOR2 (N592, N587, N483);
buf BUF1 (N593, N588);
not NOT1 (N594, N591);
nand NAND3 (N595, N594, N75, N492);
not NOT1 (N596, N593);
buf BUF1 (N597, N589);
nand NAND3 (N598, N590, N468, N558);
xor XOR2 (N599, N592, N496);
xor XOR2 (N600, N576, N194);
not NOT1 (N601, N596);
not NOT1 (N602, N595);
xor XOR2 (N603, N597, N57);
nand NAND2 (N604, N580, N8);
or OR2 (N605, N603, N94);
xor XOR2 (N606, N605, N533);
nor NOR3 (N607, N602, N537, N34);
nand NAND4 (N608, N566, N205, N337, N188);
buf BUF1 (N609, N600);
buf BUF1 (N610, N607);
and AND2 (N611, N604, N486);
or OR4 (N612, N611, N499, N486, N606);
endmodule