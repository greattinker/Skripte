// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N314,N303,N316,N256,N270,N279,N304,N309,N315,N317;

not NOT1 (N18, N4);
and AND3 (N19, N4, N17, N6);
nand NAND3 (N20, N14, N10, N11);
nor NOR4 (N21, N8, N6, N6, N4);
not NOT1 (N22, N6);
and AND3 (N23, N9, N5, N20);
nor NOR4 (N24, N22, N19, N13, N20);
and AND3 (N25, N18, N11, N13);
buf BUF1 (N26, N19);
nor NOR2 (N27, N26, N25);
buf BUF1 (N28, N9);
or OR2 (N29, N4, N15);
xor XOR2 (N30, N28, N25);
nor NOR3 (N31, N11, N25, N15);
nor NOR4 (N32, N3, N10, N1, N13);
not NOT1 (N33, N13);
nand NAND4 (N34, N21, N33, N30, N14);
or OR3 (N35, N29, N26, N8);
xor XOR2 (N36, N7, N31);
buf BUF1 (N37, N9);
buf BUF1 (N38, N31);
buf BUF1 (N39, N16);
xor XOR2 (N40, N27, N4);
xor XOR2 (N41, N40, N12);
xor XOR2 (N42, N38, N3);
or OR4 (N43, N39, N13, N40, N14);
nor NOR3 (N44, N36, N41, N16);
nand NAND2 (N45, N39, N26);
or OR4 (N46, N32, N22, N1, N18);
nand NAND3 (N47, N46, N13, N24);
not NOT1 (N48, N12);
not NOT1 (N49, N34);
buf BUF1 (N50, N47);
not NOT1 (N51, N44);
and AND3 (N52, N35, N22, N20);
buf BUF1 (N53, N43);
or OR2 (N54, N49, N16);
and AND3 (N55, N54, N50, N27);
buf BUF1 (N56, N10);
nor NOR4 (N57, N51, N36, N28, N3);
not NOT1 (N58, N56);
nand NAND2 (N59, N48, N31);
nand NAND3 (N60, N52, N32, N29);
nand NAND3 (N61, N55, N39, N15);
and AND3 (N62, N42, N3, N30);
and AND3 (N63, N61, N55, N9);
or OR2 (N64, N23, N57);
buf BUF1 (N65, N15);
nor NOR4 (N66, N37, N50, N20, N47);
buf BUF1 (N67, N53);
not NOT1 (N68, N62);
not NOT1 (N69, N65);
not NOT1 (N70, N68);
and AND4 (N71, N69, N63, N13, N60);
nor NOR2 (N72, N28, N19);
not NOT1 (N73, N50);
nor NOR3 (N74, N70, N23, N72);
not NOT1 (N75, N66);
or OR2 (N76, N15, N58);
and AND4 (N77, N40, N13, N8, N35);
nand NAND2 (N78, N67, N26);
xor XOR2 (N79, N75, N6);
or OR4 (N80, N64, N63, N26, N78);
or OR4 (N81, N57, N20, N38, N49);
and AND4 (N82, N74, N2, N77, N23);
not NOT1 (N83, N58);
or OR2 (N84, N83, N77);
nor NOR4 (N85, N76, N62, N65, N28);
xor XOR2 (N86, N79, N83);
or OR4 (N87, N82, N67, N69, N66);
nor NOR4 (N88, N73, N69, N82, N33);
not NOT1 (N89, N59);
xor XOR2 (N90, N84, N4);
buf BUF1 (N91, N80);
not NOT1 (N92, N45);
not NOT1 (N93, N90);
nand NAND4 (N94, N86, N54, N11, N65);
buf BUF1 (N95, N81);
nand NAND3 (N96, N88, N79, N24);
or OR4 (N97, N92, N57, N86, N37);
buf BUF1 (N98, N85);
xor XOR2 (N99, N96, N45);
or OR2 (N100, N94, N56);
not NOT1 (N101, N95);
nor NOR4 (N102, N93, N95, N4, N25);
or OR4 (N103, N102, N73, N81, N21);
and AND3 (N104, N99, N45, N47);
and AND2 (N105, N103, N76);
not NOT1 (N106, N71);
xor XOR2 (N107, N105, N9);
buf BUF1 (N108, N97);
xor XOR2 (N109, N100, N102);
nand NAND4 (N110, N89, N66, N70, N35);
nor NOR2 (N111, N109, N46);
xor XOR2 (N112, N110, N70);
nor NOR2 (N113, N87, N14);
or OR4 (N114, N91, N101, N99, N19);
buf BUF1 (N115, N71);
and AND2 (N116, N114, N113);
buf BUF1 (N117, N98);
nand NAND2 (N118, N52, N47);
nand NAND3 (N119, N106, N60, N20);
xor XOR2 (N120, N119, N50);
nand NAND4 (N121, N117, N107, N27, N10);
buf BUF1 (N122, N35);
buf BUF1 (N123, N122);
xor XOR2 (N124, N123, N25);
not NOT1 (N125, N108);
or OR4 (N126, N104, N125, N29, N1);
xor XOR2 (N127, N92, N38);
xor XOR2 (N128, N115, N102);
xor XOR2 (N129, N128, N67);
buf BUF1 (N130, N111);
nor NOR4 (N131, N118, N103, N12, N6);
nand NAND2 (N132, N129, N83);
xor XOR2 (N133, N132, N84);
nand NAND4 (N134, N116, N20, N101, N76);
xor XOR2 (N135, N126, N56);
not NOT1 (N136, N130);
not NOT1 (N137, N124);
and AND3 (N138, N137, N94, N128);
not NOT1 (N139, N133);
nand NAND2 (N140, N131, N93);
nand NAND4 (N141, N138, N96, N86, N29);
and AND4 (N142, N140, N54, N48, N11);
or OR4 (N143, N121, N29, N120, N10);
nand NAND4 (N144, N113, N101, N81, N25);
and AND2 (N145, N144, N71);
nor NOR4 (N146, N139, N108, N78, N28);
buf BUF1 (N147, N136);
nor NOR4 (N148, N146, N137, N56, N118);
buf BUF1 (N149, N141);
buf BUF1 (N150, N148);
buf BUF1 (N151, N142);
nor NOR3 (N152, N149, N76, N22);
xor XOR2 (N153, N150, N3);
nor NOR2 (N154, N152, N97);
nand NAND4 (N155, N145, N148, N95, N83);
and AND4 (N156, N134, N54, N18, N106);
not NOT1 (N157, N156);
nand NAND3 (N158, N143, N56, N69);
not NOT1 (N159, N155);
not NOT1 (N160, N147);
not NOT1 (N161, N127);
not NOT1 (N162, N160);
and AND3 (N163, N153, N63, N139);
xor XOR2 (N164, N112, N153);
nor NOR3 (N165, N163, N11, N28);
nand NAND3 (N166, N135, N105, N164);
not NOT1 (N167, N125);
buf BUF1 (N168, N167);
nand NAND3 (N169, N158, N168, N62);
and AND4 (N170, N15, N120, N118, N169);
nand NAND3 (N171, N165, N64, N141);
or OR4 (N172, N122, N67, N17, N93);
not NOT1 (N173, N171);
and AND4 (N174, N173, N22, N145, N69);
or OR3 (N175, N166, N123, N100);
and AND2 (N176, N175, N113);
buf BUF1 (N177, N176);
buf BUF1 (N178, N172);
and AND2 (N179, N161, N142);
not NOT1 (N180, N174);
buf BUF1 (N181, N177);
nor NOR4 (N182, N181, N166, N17, N146);
and AND3 (N183, N162, N17, N88);
xor XOR2 (N184, N179, N41);
nor NOR4 (N185, N151, N11, N98, N39);
or OR4 (N186, N180, N99, N168, N80);
nor NOR4 (N187, N183, N138, N103, N122);
or OR2 (N188, N178, N185);
nand NAND4 (N189, N14, N159, N175, N150);
buf BUF1 (N190, N85);
and AND2 (N191, N190, N185);
nand NAND2 (N192, N157, N73);
and AND3 (N193, N187, N7, N86);
nor NOR3 (N194, N189, N55, N108);
nand NAND3 (N195, N186, N63, N121);
buf BUF1 (N196, N192);
xor XOR2 (N197, N193, N164);
nor NOR4 (N198, N170, N127, N70, N129);
nand NAND3 (N199, N198, N155, N23);
nor NOR4 (N200, N188, N50, N118, N93);
nand NAND2 (N201, N195, N148);
not NOT1 (N202, N197);
and AND2 (N203, N196, N133);
nand NAND4 (N204, N184, N24, N73, N24);
not NOT1 (N205, N154);
and AND4 (N206, N191, N168, N47, N174);
and AND2 (N207, N204, N60);
nor NOR2 (N208, N202, N48);
nand NAND3 (N209, N207, N204, N79);
buf BUF1 (N210, N209);
buf BUF1 (N211, N203);
not NOT1 (N212, N199);
buf BUF1 (N213, N200);
buf BUF1 (N214, N201);
buf BUF1 (N215, N205);
nor NOR2 (N216, N215, N60);
nand NAND3 (N217, N216, N164, N183);
xor XOR2 (N218, N194, N210);
nor NOR3 (N219, N207, N74, N121);
or OR3 (N220, N211, N213, N82);
xor XOR2 (N221, N205, N127);
nand NAND2 (N222, N221, N205);
nor NOR3 (N223, N220, N153, N185);
xor XOR2 (N224, N214, N127);
or OR3 (N225, N219, N87, N21);
and AND4 (N226, N225, N112, N224, N105);
buf BUF1 (N227, N221);
and AND2 (N228, N227, N186);
and AND4 (N229, N206, N209, N113, N24);
nor NOR3 (N230, N228, N68, N220);
xor XOR2 (N231, N182, N89);
nor NOR3 (N232, N226, N217, N164);
nor NOR4 (N233, N97, N103, N73, N46);
not NOT1 (N234, N229);
xor XOR2 (N235, N222, N106);
nor NOR2 (N236, N208, N77);
nor NOR2 (N237, N218, N118);
not NOT1 (N238, N223);
buf BUF1 (N239, N236);
or OR2 (N240, N232, N21);
nor NOR3 (N241, N237, N207, N34);
nand NAND4 (N242, N238, N113, N230, N13);
not NOT1 (N243, N38);
and AND2 (N244, N239, N162);
and AND3 (N245, N240, N112, N167);
buf BUF1 (N246, N212);
nand NAND3 (N247, N242, N134, N129);
buf BUF1 (N248, N246);
and AND3 (N249, N233, N200, N167);
and AND2 (N250, N231, N75);
buf BUF1 (N251, N248);
not NOT1 (N252, N244);
not NOT1 (N253, N241);
nor NOR4 (N254, N243, N244, N138, N96);
xor XOR2 (N255, N253, N90);
nor NOR2 (N256, N249, N49);
buf BUF1 (N257, N235);
and AND4 (N258, N250, N218, N193, N229);
xor XOR2 (N259, N245, N13);
xor XOR2 (N260, N234, N124);
buf BUF1 (N261, N260);
and AND2 (N262, N255, N105);
nand NAND4 (N263, N261, N146, N147, N180);
not NOT1 (N264, N247);
xor XOR2 (N265, N264, N208);
not NOT1 (N266, N252);
nand NAND4 (N267, N251, N242, N33, N117);
xor XOR2 (N268, N265, N56);
or OR2 (N269, N267, N197);
or OR3 (N270, N268, N149, N6);
buf BUF1 (N271, N269);
and AND2 (N272, N271, N101);
nor NOR2 (N273, N254, N176);
not NOT1 (N274, N257);
xor XOR2 (N275, N259, N74);
xor XOR2 (N276, N272, N91);
xor XOR2 (N277, N276, N271);
xor XOR2 (N278, N262, N95);
buf BUF1 (N279, N258);
not NOT1 (N280, N275);
buf BUF1 (N281, N263);
xor XOR2 (N282, N278, N184);
xor XOR2 (N283, N280, N98);
nand NAND2 (N284, N282, N195);
xor XOR2 (N285, N273, N239);
buf BUF1 (N286, N281);
nand NAND4 (N287, N283, N191, N131, N29);
nand NAND2 (N288, N266, N274);
or OR2 (N289, N285, N220);
or OR4 (N290, N189, N134, N230, N73);
buf BUF1 (N291, N286);
nor NOR4 (N292, N284, N53, N281, N228);
and AND3 (N293, N289, N238, N91);
nand NAND4 (N294, N293, N32, N278, N264);
and AND3 (N295, N287, N147, N190);
or OR3 (N296, N288, N294, N53);
not NOT1 (N297, N294);
or OR2 (N298, N291, N242);
nand NAND3 (N299, N290, N77, N217);
not NOT1 (N300, N292);
xor XOR2 (N301, N297, N239);
xor XOR2 (N302, N299, N50);
xor XOR2 (N303, N298, N68);
not NOT1 (N304, N301);
nand NAND2 (N305, N302, N295);
buf BUF1 (N306, N227);
nor NOR3 (N307, N277, N76, N283);
xor XOR2 (N308, N300, N122);
buf BUF1 (N309, N305);
buf BUF1 (N310, N307);
not NOT1 (N311, N310);
not NOT1 (N312, N311);
nor NOR3 (N313, N296, N147, N152);
buf BUF1 (N314, N306);
or OR2 (N315, N312, N111);
nor NOR2 (N316, N308, N299);
or OR2 (N317, N313, N135);
endmodule