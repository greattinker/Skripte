// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N8023,N8009,N8013,N8020,N8012,N8022,N8021,N8014,N8017,N8024;

buf BUF1 (N25, N6);
and AND2 (N26, N2, N2);
nand NAND4 (N27, N7, N10, N3, N18);
or OR3 (N28, N4, N9, N5);
nand NAND3 (N29, N3, N13, N26);
buf BUF1 (N30, N8);
not NOT1 (N31, N21);
or OR4 (N32, N31, N11, N15, N20);
xor XOR2 (N33, N3, N6);
xor XOR2 (N34, N1, N1);
nand NAND2 (N35, N3, N9);
and AND3 (N36, N22, N11, N30);
or OR3 (N37, N14, N22, N23);
or OR4 (N38, N37, N17, N9, N24);
nor NOR3 (N39, N33, N33, N9);
and AND4 (N40, N25, N3, N1, N7);
or OR3 (N41, N39, N22, N40);
nand NAND4 (N42, N6, N22, N11, N39);
nand NAND3 (N43, N29, N28, N39);
or OR3 (N44, N4, N43, N31);
or OR4 (N45, N23, N1, N8, N30);
or OR2 (N46, N41, N17);
or OR2 (N47, N36, N5);
or OR4 (N48, N45, N46, N39, N28);
buf BUF1 (N49, N9);
nand NAND3 (N50, N49, N23, N15);
nand NAND2 (N51, N32, N42);
nand NAND4 (N52, N44, N5, N1, N39);
or OR2 (N53, N32, N32);
nor NOR4 (N54, N48, N5, N11, N39);
and AND3 (N55, N51, N7, N12);
not NOT1 (N56, N27);
nand NAND4 (N57, N53, N42, N11, N18);
nand NAND4 (N58, N57, N51, N28, N40);
nand NAND4 (N59, N52, N41, N35, N40);
nor NOR2 (N60, N59, N49);
not NOT1 (N61, N22);
not NOT1 (N62, N38);
not NOT1 (N63, N61);
nand NAND3 (N64, N60, N60, N47);
buf BUF1 (N65, N22);
nor NOR3 (N66, N55, N33, N58);
nand NAND4 (N67, N51, N47, N52, N51);
and AND2 (N68, N67, N67);
nor NOR4 (N69, N68, N14, N68, N27);
nor NOR2 (N70, N63, N59);
nand NAND3 (N71, N64, N43, N34);
xor XOR2 (N72, N54, N28);
and AND3 (N73, N26, N48, N68);
or OR2 (N74, N56, N25);
not NOT1 (N75, N71);
xor XOR2 (N76, N74, N54);
nand NAND2 (N77, N73, N15);
buf BUF1 (N78, N65);
nor NOR4 (N79, N76, N75, N67, N39);
or OR3 (N80, N17, N9, N48);
and AND4 (N81, N50, N31, N59, N53);
and AND2 (N82, N72, N69);
xor XOR2 (N83, N33, N59);
and AND3 (N84, N80, N57, N64);
nand NAND3 (N85, N78, N42, N11);
nand NAND4 (N86, N81, N37, N39, N1);
or OR3 (N87, N70, N28, N41);
nor NOR2 (N88, N62, N36);
xor XOR2 (N89, N66, N64);
buf BUF1 (N90, N87);
and AND4 (N91, N88, N9, N48, N46);
buf BUF1 (N92, N91);
nor NOR4 (N93, N77, N65, N47, N72);
xor XOR2 (N94, N92, N13);
or OR3 (N95, N84, N23, N59);
nand NAND3 (N96, N89, N63, N45);
nor NOR4 (N97, N86, N38, N53, N58);
and AND4 (N98, N85, N94, N96, N21);
nor NOR2 (N99, N12, N73);
or OR3 (N100, N5, N70, N33);
nor NOR3 (N101, N98, N34, N54);
buf BUF1 (N102, N83);
buf BUF1 (N103, N90);
xor XOR2 (N104, N82, N36);
nand NAND4 (N105, N97, N104, N36, N79);
nor NOR3 (N106, N105, N51, N76);
nor NOR4 (N107, N83, N32, N18, N40);
nand NAND4 (N108, N101, N81, N90, N76);
buf BUF1 (N109, N49);
and AND2 (N110, N103, N19);
nor NOR3 (N111, N93, N34, N77);
nor NOR3 (N112, N99, N34, N20);
or OR3 (N113, N95, N111, N81);
nor NOR3 (N114, N3, N46, N23);
not NOT1 (N115, N112);
buf BUF1 (N116, N113);
buf BUF1 (N117, N116);
buf BUF1 (N118, N117);
not NOT1 (N119, N114);
or OR2 (N120, N102, N59);
nand NAND3 (N121, N107, N63, N119);
or OR3 (N122, N3, N86, N4);
xor XOR2 (N123, N121, N52);
or OR4 (N124, N108, N67, N106, N43);
nand NAND2 (N125, N3, N90);
or OR2 (N126, N122, N21);
not NOT1 (N127, N118);
buf BUF1 (N128, N109);
not NOT1 (N129, N126);
nand NAND3 (N130, N110, N56, N126);
not NOT1 (N131, N124);
buf BUF1 (N132, N130);
buf BUF1 (N133, N100);
buf BUF1 (N134, N127);
not NOT1 (N135, N120);
buf BUF1 (N136, N129);
and AND4 (N137, N131, N105, N93, N71);
xor XOR2 (N138, N134, N65);
nand NAND3 (N139, N138, N98, N41);
buf BUF1 (N140, N139);
nor NOR4 (N141, N137, N110, N124, N91);
and AND4 (N142, N132, N113, N86, N42);
and AND4 (N143, N140, N82, N15, N131);
or OR4 (N144, N136, N104, N98, N125);
or OR3 (N145, N31, N37, N17);
xor XOR2 (N146, N145, N129);
or OR4 (N147, N123, N73, N15, N120);
not NOT1 (N148, N115);
nor NOR2 (N149, N143, N133);
or OR3 (N150, N45, N91, N93);
buf BUF1 (N151, N148);
xor XOR2 (N152, N135, N65);
xor XOR2 (N153, N144, N53);
not NOT1 (N154, N141);
xor XOR2 (N155, N149, N33);
buf BUF1 (N156, N128);
or OR2 (N157, N155, N16);
or OR2 (N158, N146, N2);
nand NAND4 (N159, N147, N54, N139, N13);
nor NOR3 (N160, N157, N66, N154);
not NOT1 (N161, N26);
nand NAND2 (N162, N159, N24);
nand NAND3 (N163, N158, N87, N112);
buf BUF1 (N164, N160);
buf BUF1 (N165, N161);
nor NOR4 (N166, N165, N51, N84, N24);
not NOT1 (N167, N163);
or OR3 (N168, N153, N148, N96);
nor NOR2 (N169, N168, N27);
xor XOR2 (N170, N151, N42);
not NOT1 (N171, N164);
and AND2 (N172, N162, N63);
xor XOR2 (N173, N150, N36);
nand NAND4 (N174, N172, N134, N167, N152);
xor XOR2 (N175, N52, N136);
xor XOR2 (N176, N30, N21);
nor NOR4 (N177, N176, N99, N67, N94);
not NOT1 (N178, N166);
and AND3 (N179, N142, N155, N64);
or OR3 (N180, N175, N114, N45);
not NOT1 (N181, N177);
xor XOR2 (N182, N169, N90);
not NOT1 (N183, N182);
nand NAND3 (N184, N174, N106, N65);
nor NOR3 (N185, N173, N119, N103);
nand NAND3 (N186, N181, N135, N161);
nand NAND4 (N187, N186, N1, N74, N11);
or OR2 (N188, N185, N130);
buf BUF1 (N189, N179);
xor XOR2 (N190, N189, N85);
buf BUF1 (N191, N170);
xor XOR2 (N192, N171, N180);
buf BUF1 (N193, N13);
and AND2 (N194, N187, N116);
and AND3 (N195, N178, N6, N17);
nand NAND2 (N196, N193, N157);
not NOT1 (N197, N194);
nor NOR2 (N198, N188, N11);
not NOT1 (N199, N183);
not NOT1 (N200, N192);
nor NOR4 (N201, N184, N139, N38, N185);
and AND4 (N202, N198, N143, N7, N91);
buf BUF1 (N203, N156);
or OR2 (N204, N200, N192);
xor XOR2 (N205, N199, N143);
nand NAND3 (N206, N196, N29, N97);
buf BUF1 (N207, N206);
or OR4 (N208, N204, N25, N87, N66);
or OR3 (N209, N207, N94, N3);
or OR2 (N210, N203, N162);
or OR4 (N211, N197, N159, N129, N138);
and AND3 (N212, N201, N55, N197);
not NOT1 (N213, N191);
nand NAND2 (N214, N208, N172);
nor NOR3 (N215, N214, N68, N66);
nor NOR3 (N216, N213, N52, N113);
nand NAND4 (N217, N210, N108, N208, N9);
xor XOR2 (N218, N211, N204);
and AND3 (N219, N209, N115, N176);
or OR4 (N220, N195, N174, N14, N92);
and AND2 (N221, N218, N71);
nand NAND2 (N222, N220, N105);
or OR3 (N223, N190, N198, N188);
and AND2 (N224, N217, N61);
and AND4 (N225, N219, N102, N216, N208);
nand NAND2 (N226, N152, N52);
nor NOR4 (N227, N212, N66, N3, N57);
nor NOR2 (N228, N225, N108);
or OR4 (N229, N202, N140, N212, N200);
xor XOR2 (N230, N221, N108);
not NOT1 (N231, N222);
nor NOR3 (N232, N231, N123, N224);
xor XOR2 (N233, N182, N140);
xor XOR2 (N234, N227, N80);
and AND2 (N235, N232, N158);
nand NAND4 (N236, N223, N77, N18, N164);
nand NAND3 (N237, N233, N233, N174);
or OR4 (N238, N230, N195, N197, N52);
not NOT1 (N239, N234);
xor XOR2 (N240, N215, N144);
nand NAND2 (N241, N238, N129);
buf BUF1 (N242, N226);
not NOT1 (N243, N236);
xor XOR2 (N244, N228, N60);
nand NAND4 (N245, N240, N51, N21, N165);
xor XOR2 (N246, N237, N183);
xor XOR2 (N247, N243, N78);
not NOT1 (N248, N245);
buf BUF1 (N249, N235);
and AND2 (N250, N242, N245);
buf BUF1 (N251, N239);
buf BUF1 (N252, N249);
nor NOR3 (N253, N250, N74, N33);
xor XOR2 (N254, N244, N70);
or OR2 (N255, N251, N192);
nor NOR2 (N256, N253, N93);
not NOT1 (N257, N229);
nand NAND2 (N258, N255, N146);
xor XOR2 (N259, N241, N180);
or OR2 (N260, N254, N96);
buf BUF1 (N261, N256);
buf BUF1 (N262, N205);
nand NAND2 (N263, N259, N223);
nor NOR3 (N264, N246, N58, N40);
xor XOR2 (N265, N261, N91);
nand NAND2 (N266, N258, N100);
buf BUF1 (N267, N248);
xor XOR2 (N268, N260, N138);
not NOT1 (N269, N264);
nand NAND3 (N270, N266, N258, N214);
not NOT1 (N271, N262);
nor NOR4 (N272, N269, N151, N241, N9);
xor XOR2 (N273, N263, N185);
not NOT1 (N274, N247);
and AND4 (N275, N265, N257, N81, N69);
nor NOR3 (N276, N60, N29, N264);
xor XOR2 (N277, N268, N72);
not NOT1 (N278, N271);
and AND4 (N279, N267, N162, N259, N79);
buf BUF1 (N280, N274);
or OR3 (N281, N278, N185, N231);
or OR2 (N282, N270, N235);
and AND4 (N283, N280, N273, N139, N69);
nor NOR2 (N284, N86, N162);
not NOT1 (N285, N281);
buf BUF1 (N286, N272);
and AND2 (N287, N286, N159);
nand NAND4 (N288, N285, N101, N181, N40);
or OR3 (N289, N276, N263, N203);
buf BUF1 (N290, N283);
buf BUF1 (N291, N284);
not NOT1 (N292, N290);
nor NOR4 (N293, N275, N247, N232, N46);
or OR2 (N294, N292, N259);
not NOT1 (N295, N291);
nor NOR3 (N296, N252, N292, N139);
or OR3 (N297, N295, N262, N293);
not NOT1 (N298, N269);
or OR3 (N299, N288, N212, N153);
not NOT1 (N300, N294);
buf BUF1 (N301, N300);
nand NAND2 (N302, N296, N143);
or OR2 (N303, N287, N208);
nor NOR2 (N304, N297, N26);
or OR4 (N305, N298, N124, N253, N67);
buf BUF1 (N306, N289);
not NOT1 (N307, N277);
and AND3 (N308, N303, N54, N153);
xor XOR2 (N309, N308, N78);
xor XOR2 (N310, N302, N274);
buf BUF1 (N311, N299);
and AND3 (N312, N305, N252, N24);
xor XOR2 (N313, N307, N5);
or OR2 (N314, N310, N19);
buf BUF1 (N315, N306);
xor XOR2 (N316, N282, N111);
not NOT1 (N317, N315);
buf BUF1 (N318, N314);
and AND4 (N319, N301, N264, N296, N18);
xor XOR2 (N320, N311, N165);
not NOT1 (N321, N317);
xor XOR2 (N322, N318, N9);
nor NOR4 (N323, N279, N300, N102, N253);
buf BUF1 (N324, N323);
or OR3 (N325, N312, N23, N121);
nor NOR4 (N326, N309, N17, N212, N101);
or OR2 (N327, N304, N26);
xor XOR2 (N328, N321, N91);
nand NAND4 (N329, N327, N110, N295, N129);
and AND4 (N330, N320, N43, N239, N197);
or OR4 (N331, N319, N239, N238, N130);
and AND3 (N332, N322, N1, N286);
xor XOR2 (N333, N330, N312);
buf BUF1 (N334, N333);
and AND3 (N335, N334, N206, N217);
and AND2 (N336, N325, N166);
or OR4 (N337, N324, N103, N103, N271);
nand NAND4 (N338, N336, N19, N283, N24);
or OR4 (N339, N329, N121, N334, N309);
nor NOR2 (N340, N316, N126);
or OR3 (N341, N338, N8, N158);
buf BUF1 (N342, N313);
xor XOR2 (N343, N328, N81);
nor NOR4 (N344, N335, N126, N21, N53);
or OR3 (N345, N342, N307, N184);
nand NAND2 (N346, N343, N50);
not NOT1 (N347, N345);
nor NOR4 (N348, N337, N151, N35, N198);
nand NAND2 (N349, N326, N185);
nand NAND2 (N350, N348, N326);
and AND4 (N351, N349, N138, N12, N347);
not NOT1 (N352, N314);
xor XOR2 (N353, N340, N230);
or OR4 (N354, N332, N85, N247, N93);
nand NAND2 (N355, N353, N85);
buf BUF1 (N356, N352);
and AND4 (N357, N341, N141, N177, N199);
not NOT1 (N358, N354);
not NOT1 (N359, N350);
and AND4 (N360, N346, N214, N53, N321);
and AND4 (N361, N360, N219, N17, N248);
or OR4 (N362, N355, N123, N118, N289);
not NOT1 (N363, N356);
nand NAND3 (N364, N339, N294, N314);
buf BUF1 (N365, N362);
not NOT1 (N366, N351);
not NOT1 (N367, N344);
xor XOR2 (N368, N361, N100);
and AND3 (N369, N358, N231, N135);
nand NAND2 (N370, N367, N173);
not NOT1 (N371, N366);
and AND4 (N372, N359, N278, N31, N200);
not NOT1 (N373, N369);
nor NOR2 (N374, N373, N193);
nand NAND3 (N375, N371, N297, N64);
xor XOR2 (N376, N372, N76);
not NOT1 (N377, N370);
xor XOR2 (N378, N364, N119);
nor NOR4 (N379, N357, N372, N63, N127);
or OR3 (N380, N375, N92, N17);
nand NAND3 (N381, N331, N278, N36);
nor NOR4 (N382, N365, N6, N240, N109);
xor XOR2 (N383, N374, N161);
nor NOR2 (N384, N380, N341);
nand NAND3 (N385, N376, N343, N362);
not NOT1 (N386, N379);
and AND3 (N387, N381, N30, N31);
buf BUF1 (N388, N368);
nor NOR2 (N389, N378, N132);
xor XOR2 (N390, N384, N188);
or OR4 (N391, N387, N351, N48, N86);
nand NAND3 (N392, N389, N271, N252);
xor XOR2 (N393, N363, N269);
and AND4 (N394, N385, N187, N127, N321);
buf BUF1 (N395, N392);
buf BUF1 (N396, N394);
xor XOR2 (N397, N393, N84);
xor XOR2 (N398, N386, N167);
not NOT1 (N399, N398);
and AND2 (N400, N382, N171);
xor XOR2 (N401, N388, N4);
nand NAND4 (N402, N377, N4, N393, N198);
not NOT1 (N403, N390);
xor XOR2 (N404, N391, N32);
not NOT1 (N405, N400);
buf BUF1 (N406, N395);
not NOT1 (N407, N406);
xor XOR2 (N408, N402, N180);
not NOT1 (N409, N397);
nand NAND3 (N410, N407, N120, N340);
xor XOR2 (N411, N403, N157);
buf BUF1 (N412, N399);
or OR3 (N413, N409, N395, N370);
not NOT1 (N414, N405);
not NOT1 (N415, N404);
not NOT1 (N416, N410);
and AND3 (N417, N411, N228, N176);
buf BUF1 (N418, N413);
not NOT1 (N419, N416);
nor NOR3 (N420, N401, N361, N155);
not NOT1 (N421, N415);
buf BUF1 (N422, N419);
and AND2 (N423, N383, N158);
not NOT1 (N424, N422);
nor NOR4 (N425, N396, N281, N167, N341);
nand NAND3 (N426, N408, N403, N279);
buf BUF1 (N427, N414);
buf BUF1 (N428, N412);
nand NAND3 (N429, N426, N309, N253);
buf BUF1 (N430, N427);
buf BUF1 (N431, N421);
nor NOR4 (N432, N418, N385, N74, N402);
or OR2 (N433, N417, N424);
buf BUF1 (N434, N29);
nor NOR4 (N435, N425, N42, N70, N376);
nor NOR3 (N436, N420, N397, N163);
or OR2 (N437, N436, N259);
buf BUF1 (N438, N435);
and AND4 (N439, N432, N53, N378, N384);
nand NAND2 (N440, N431, N375);
xor XOR2 (N441, N438, N182);
nor NOR3 (N442, N440, N84, N187);
and AND2 (N443, N428, N167);
buf BUF1 (N444, N437);
nand NAND4 (N445, N429, N329, N110, N158);
or OR4 (N446, N433, N302, N328, N282);
xor XOR2 (N447, N441, N234);
xor XOR2 (N448, N443, N165);
nor NOR3 (N449, N445, N407, N59);
nor NOR2 (N450, N444, N60);
and AND2 (N451, N447, N62);
buf BUF1 (N452, N442);
xor XOR2 (N453, N450, N193);
or OR4 (N454, N449, N50, N204, N29);
or OR3 (N455, N434, N401, N19);
xor XOR2 (N456, N430, N374);
nand NAND4 (N457, N455, N119, N43, N144);
and AND3 (N458, N454, N294, N224);
xor XOR2 (N459, N446, N203);
or OR3 (N460, N451, N347, N141);
nor NOR2 (N461, N453, N177);
not NOT1 (N462, N461);
nand NAND2 (N463, N460, N31);
nand NAND2 (N464, N452, N193);
or OR3 (N465, N439, N410, N83);
nor NOR2 (N466, N465, N365);
buf BUF1 (N467, N462);
buf BUF1 (N468, N457);
nand NAND3 (N469, N463, N342, N466);
nor NOR3 (N470, N170, N326, N91);
buf BUF1 (N471, N423);
buf BUF1 (N472, N459);
nand NAND2 (N473, N468, N183);
not NOT1 (N474, N469);
nor NOR3 (N475, N456, N362, N220);
nor NOR2 (N476, N448, N259);
or OR3 (N477, N471, N142, N27);
and AND3 (N478, N470, N103, N469);
nor NOR3 (N479, N474, N7, N38);
not NOT1 (N480, N478);
nor NOR3 (N481, N476, N276, N302);
xor XOR2 (N482, N467, N396);
nand NAND4 (N483, N481, N172, N335, N304);
or OR4 (N484, N472, N210, N359, N220);
nand NAND3 (N485, N483, N424, N135);
nor NOR4 (N486, N484, N116, N408, N440);
xor XOR2 (N487, N479, N418);
xor XOR2 (N488, N482, N5);
xor XOR2 (N489, N475, N212);
not NOT1 (N490, N487);
buf BUF1 (N491, N458);
and AND2 (N492, N480, N312);
buf BUF1 (N493, N464);
nor NOR2 (N494, N490, N50);
xor XOR2 (N495, N473, N434);
nand NAND4 (N496, N492, N67, N53, N421);
not NOT1 (N497, N485);
nand NAND2 (N498, N497, N62);
xor XOR2 (N499, N493, N11);
xor XOR2 (N500, N488, N225);
nor NOR4 (N501, N496, N4, N71, N117);
not NOT1 (N502, N495);
and AND2 (N503, N486, N431);
buf BUF1 (N504, N498);
xor XOR2 (N505, N501, N116);
nand NAND3 (N506, N491, N231, N134);
and AND2 (N507, N502, N200);
nand NAND2 (N508, N494, N181);
not NOT1 (N509, N503);
buf BUF1 (N510, N499);
and AND4 (N511, N504, N145, N290, N291);
buf BUF1 (N512, N508);
or OR3 (N513, N509, N422, N183);
nand NAND2 (N514, N512, N292);
xor XOR2 (N515, N506, N187);
not NOT1 (N516, N500);
or OR2 (N517, N515, N446);
xor XOR2 (N518, N517, N405);
xor XOR2 (N519, N477, N497);
xor XOR2 (N520, N513, N165);
nand NAND2 (N521, N510, N22);
buf BUF1 (N522, N521);
nand NAND4 (N523, N505, N384, N16, N459);
nor NOR3 (N524, N520, N260, N452);
nand NAND3 (N525, N522, N493, N480);
and AND2 (N526, N514, N144);
nor NOR3 (N527, N525, N94, N267);
or OR2 (N528, N511, N87);
buf BUF1 (N529, N489);
nor NOR3 (N530, N524, N488, N458);
and AND2 (N531, N526, N458);
not NOT1 (N532, N527);
buf BUF1 (N533, N518);
and AND2 (N534, N533, N163);
xor XOR2 (N535, N507, N47);
xor XOR2 (N536, N516, N524);
buf BUF1 (N537, N535);
nor NOR3 (N538, N530, N198, N494);
nor NOR3 (N539, N534, N323, N317);
or OR4 (N540, N519, N378, N188, N124);
or OR2 (N541, N528, N363);
or OR4 (N542, N523, N30, N245, N342);
nand NAND4 (N543, N542, N461, N15, N328);
not NOT1 (N544, N532);
nand NAND4 (N545, N543, N489, N290, N446);
buf BUF1 (N546, N545);
nand NAND3 (N547, N537, N445, N434);
nor NOR4 (N548, N546, N221, N195, N230);
not NOT1 (N549, N531);
nor NOR2 (N550, N548, N127);
nand NAND2 (N551, N536, N515);
xor XOR2 (N552, N550, N10);
nand NAND2 (N553, N540, N286);
buf BUF1 (N554, N544);
xor XOR2 (N555, N541, N149);
not NOT1 (N556, N539);
or OR4 (N557, N529, N522, N307, N469);
and AND2 (N558, N547, N511);
not NOT1 (N559, N554);
buf BUF1 (N560, N555);
buf BUF1 (N561, N552);
xor XOR2 (N562, N560, N84);
not NOT1 (N563, N553);
nor NOR4 (N564, N559, N245, N129, N368);
and AND3 (N565, N556, N441, N90);
buf BUF1 (N566, N561);
nor NOR4 (N567, N558, N151, N423, N475);
or OR3 (N568, N567, N42, N356);
or OR3 (N569, N557, N355, N361);
not NOT1 (N570, N568);
or OR2 (N571, N538, N506);
nor NOR3 (N572, N570, N504, N359);
and AND4 (N573, N563, N378, N9, N185);
or OR3 (N574, N549, N261, N96);
and AND3 (N575, N562, N532, N567);
nand NAND4 (N576, N571, N162, N564, N462);
nor NOR4 (N577, N188, N147, N274, N414);
xor XOR2 (N578, N551, N417);
not NOT1 (N579, N566);
buf BUF1 (N580, N565);
not NOT1 (N581, N576);
nand NAND3 (N582, N578, N321, N580);
nand NAND2 (N583, N260, N391);
nor NOR4 (N584, N569, N273, N186, N235);
buf BUF1 (N585, N581);
buf BUF1 (N586, N572);
nand NAND2 (N587, N577, N473);
buf BUF1 (N588, N587);
or OR2 (N589, N585, N312);
or OR4 (N590, N584, N366, N375, N107);
nor NOR3 (N591, N582, N385, N417);
or OR4 (N592, N573, N188, N188, N361);
nand NAND4 (N593, N591, N195, N515, N306);
not NOT1 (N594, N588);
xor XOR2 (N595, N593, N410);
nand NAND2 (N596, N579, N27);
xor XOR2 (N597, N575, N83);
buf BUF1 (N598, N586);
or OR2 (N599, N574, N382);
xor XOR2 (N600, N594, N491);
buf BUF1 (N601, N592);
nor NOR4 (N602, N589, N326, N390, N530);
not NOT1 (N603, N600);
nand NAND4 (N604, N590, N449, N593, N225);
xor XOR2 (N605, N604, N60);
nor NOR3 (N606, N596, N278, N188);
not NOT1 (N607, N602);
or OR4 (N608, N606, N477, N476, N412);
not NOT1 (N609, N595);
buf BUF1 (N610, N609);
or OR2 (N611, N597, N455);
xor XOR2 (N612, N603, N222);
xor XOR2 (N613, N605, N510);
or OR3 (N614, N612, N257, N200);
buf BUF1 (N615, N608);
or OR4 (N616, N598, N311, N173, N575);
and AND4 (N617, N611, N536, N325, N591);
and AND4 (N618, N607, N280, N444, N74);
buf BUF1 (N619, N599);
nor NOR3 (N620, N619, N54, N9);
buf BUF1 (N621, N618);
buf BUF1 (N622, N620);
or OR3 (N623, N615, N243, N290);
and AND2 (N624, N621, N375);
and AND3 (N625, N614, N222, N90);
nor NOR4 (N626, N625, N237, N479, N471);
or OR2 (N627, N622, N546);
nand NAND2 (N628, N627, N453);
xor XOR2 (N629, N626, N381);
buf BUF1 (N630, N583);
xor XOR2 (N631, N610, N77);
buf BUF1 (N632, N628);
nand NAND3 (N633, N623, N480, N577);
or OR2 (N634, N629, N580);
not NOT1 (N635, N617);
nor NOR3 (N636, N631, N298, N474);
xor XOR2 (N637, N616, N130);
xor XOR2 (N638, N633, N238);
nor NOR2 (N639, N638, N101);
xor XOR2 (N640, N636, N66);
not NOT1 (N641, N632);
nand NAND2 (N642, N634, N332);
nand NAND4 (N643, N637, N271, N94, N320);
nand NAND2 (N644, N643, N75);
or OR3 (N645, N630, N266, N8);
xor XOR2 (N646, N635, N455);
buf BUF1 (N647, N645);
xor XOR2 (N648, N642, N216);
and AND2 (N649, N639, N35);
nor NOR2 (N650, N646, N355);
nor NOR4 (N651, N647, N12, N539, N167);
or OR3 (N652, N641, N485, N295);
xor XOR2 (N653, N648, N541);
not NOT1 (N654, N624);
or OR3 (N655, N613, N100, N520);
buf BUF1 (N656, N654);
or OR3 (N657, N644, N423, N635);
buf BUF1 (N658, N651);
or OR4 (N659, N650, N122, N82, N246);
nor NOR3 (N660, N649, N109, N570);
not NOT1 (N661, N658);
or OR4 (N662, N657, N99, N137, N499);
nand NAND4 (N663, N640, N30, N261, N442);
or OR4 (N664, N661, N518, N125, N408);
or OR2 (N665, N663, N10);
nand NAND3 (N666, N653, N232, N508);
xor XOR2 (N667, N664, N419);
nand NAND3 (N668, N652, N3, N571);
nand NAND2 (N669, N668, N390);
buf BUF1 (N670, N656);
or OR3 (N671, N667, N223, N630);
buf BUF1 (N672, N601);
and AND3 (N673, N672, N399, N130);
xor XOR2 (N674, N660, N568);
nand NAND4 (N675, N666, N461, N195, N184);
xor XOR2 (N676, N655, N417);
buf BUF1 (N677, N675);
not NOT1 (N678, N673);
nor NOR3 (N679, N662, N70, N13);
nand NAND2 (N680, N659, N288);
and AND2 (N681, N676, N391);
nand NAND4 (N682, N679, N132, N300, N241);
nand NAND2 (N683, N674, N355);
not NOT1 (N684, N681);
buf BUF1 (N685, N680);
nand NAND2 (N686, N670, N482);
nor NOR4 (N687, N682, N208, N307, N536);
nor NOR4 (N688, N685, N541, N424, N374);
nor NOR4 (N689, N678, N446, N392, N11);
and AND3 (N690, N684, N305, N32);
nand NAND2 (N691, N688, N424);
nor NOR3 (N692, N665, N348, N653);
not NOT1 (N693, N683);
nand NAND4 (N694, N669, N418, N669, N489);
not NOT1 (N695, N689);
xor XOR2 (N696, N686, N497);
buf BUF1 (N697, N687);
not NOT1 (N698, N690);
nand NAND4 (N699, N696, N535, N445, N449);
buf BUF1 (N700, N693);
nand NAND3 (N701, N699, N313, N618);
buf BUF1 (N702, N701);
buf BUF1 (N703, N698);
nand NAND4 (N704, N694, N504, N242, N657);
nor NOR4 (N705, N700, N131, N577, N699);
nor NOR3 (N706, N677, N668, N251);
and AND3 (N707, N671, N504, N656);
nor NOR2 (N708, N695, N7);
not NOT1 (N709, N707);
and AND2 (N710, N706, N36);
nor NOR4 (N711, N709, N110, N36, N70);
buf BUF1 (N712, N692);
not NOT1 (N713, N703);
buf BUF1 (N714, N697);
nor NOR4 (N715, N713, N392, N79, N677);
nand NAND2 (N716, N708, N575);
nor NOR3 (N717, N710, N246, N303);
nand NAND4 (N718, N691, N66, N61, N284);
or OR4 (N719, N711, N261, N271, N118);
or OR2 (N720, N705, N336);
or OR4 (N721, N702, N648, N583, N376);
xor XOR2 (N722, N716, N441);
xor XOR2 (N723, N721, N464);
not NOT1 (N724, N719);
or OR4 (N725, N720, N126, N390, N672);
xor XOR2 (N726, N724, N190);
not NOT1 (N727, N704);
or OR2 (N728, N714, N179);
buf BUF1 (N729, N728);
nor NOR3 (N730, N717, N282, N185);
xor XOR2 (N731, N725, N173);
or OR3 (N732, N726, N651, N497);
nor NOR4 (N733, N715, N659, N45, N502);
xor XOR2 (N734, N718, N140);
buf BUF1 (N735, N733);
xor XOR2 (N736, N729, N296);
xor XOR2 (N737, N723, N127);
and AND2 (N738, N735, N20);
xor XOR2 (N739, N730, N669);
nand NAND2 (N740, N731, N341);
and AND3 (N741, N727, N54, N361);
xor XOR2 (N742, N734, N435);
and AND2 (N743, N740, N686);
xor XOR2 (N744, N712, N718);
or OR4 (N745, N738, N64, N171, N378);
nor NOR2 (N746, N742, N467);
buf BUF1 (N747, N744);
and AND2 (N748, N732, N131);
and AND4 (N749, N722, N457, N49, N724);
and AND2 (N750, N739, N256);
buf BUF1 (N751, N747);
xor XOR2 (N752, N736, N263);
xor XOR2 (N753, N751, N387);
xor XOR2 (N754, N750, N535);
nor NOR3 (N755, N746, N305, N261);
xor XOR2 (N756, N741, N614);
and AND4 (N757, N749, N666, N370, N60);
nand NAND3 (N758, N756, N679, N94);
xor XOR2 (N759, N755, N401);
nand NAND3 (N760, N752, N487, N478);
not NOT1 (N761, N754);
not NOT1 (N762, N758);
and AND2 (N763, N761, N76);
or OR4 (N764, N763, N142, N486, N610);
buf BUF1 (N765, N764);
or OR4 (N766, N743, N658, N676, N117);
or OR3 (N767, N759, N601, N556);
nand NAND4 (N768, N745, N387, N701, N110);
nor NOR3 (N769, N748, N117, N662);
not NOT1 (N770, N753);
and AND2 (N771, N767, N725);
nor NOR4 (N772, N766, N8, N191, N505);
and AND3 (N773, N762, N558, N213);
not NOT1 (N774, N770);
and AND4 (N775, N769, N569, N312, N328);
xor XOR2 (N776, N771, N488);
not NOT1 (N777, N737);
buf BUF1 (N778, N757);
not NOT1 (N779, N760);
buf BUF1 (N780, N774);
buf BUF1 (N781, N778);
or OR2 (N782, N765, N255);
nand NAND2 (N783, N779, N468);
xor XOR2 (N784, N780, N409);
or OR4 (N785, N768, N540, N86, N244);
or OR2 (N786, N773, N137);
nand NAND2 (N787, N782, N346);
buf BUF1 (N788, N786);
nand NAND2 (N789, N788, N560);
not NOT1 (N790, N789);
buf BUF1 (N791, N772);
nor NOR2 (N792, N776, N396);
and AND2 (N793, N775, N369);
xor XOR2 (N794, N792, N330);
xor XOR2 (N795, N791, N782);
and AND4 (N796, N790, N640, N554, N761);
and AND3 (N797, N777, N216, N622);
or OR4 (N798, N783, N201, N368, N168);
xor XOR2 (N799, N796, N155);
not NOT1 (N800, N781);
or OR2 (N801, N793, N470);
xor XOR2 (N802, N795, N44);
buf BUF1 (N803, N802);
not NOT1 (N804, N798);
nand NAND3 (N805, N785, N554, N581);
or OR3 (N806, N799, N734, N5);
xor XOR2 (N807, N784, N343);
not NOT1 (N808, N797);
nand NAND2 (N809, N794, N539);
and AND4 (N810, N803, N608, N265, N100);
nor NOR3 (N811, N801, N530, N694);
buf BUF1 (N812, N787);
nand NAND4 (N813, N810, N55, N763, N550);
nand NAND2 (N814, N808, N588);
not NOT1 (N815, N805);
buf BUF1 (N816, N807);
nor NOR4 (N817, N800, N177, N738, N291);
not NOT1 (N818, N804);
or OR3 (N819, N811, N444, N227);
not NOT1 (N820, N817);
xor XOR2 (N821, N816, N364);
xor XOR2 (N822, N813, N583);
buf BUF1 (N823, N822);
and AND4 (N824, N809, N201, N768, N147);
or OR3 (N825, N824, N681, N243);
xor XOR2 (N826, N821, N793);
buf BUF1 (N827, N812);
not NOT1 (N828, N820);
and AND3 (N829, N827, N86, N98);
buf BUF1 (N830, N826);
nor NOR2 (N831, N823, N257);
nor NOR3 (N832, N829, N778, N149);
buf BUF1 (N833, N828);
nor NOR4 (N834, N818, N419, N190, N75);
xor XOR2 (N835, N819, N656);
not NOT1 (N836, N806);
or OR2 (N837, N830, N187);
or OR4 (N838, N836, N704, N12, N701);
xor XOR2 (N839, N835, N318);
nand NAND4 (N840, N825, N327, N554, N546);
or OR3 (N841, N814, N122, N689);
buf BUF1 (N842, N839);
buf BUF1 (N843, N842);
nand NAND4 (N844, N815, N596, N496, N679);
xor XOR2 (N845, N840, N178);
and AND4 (N846, N833, N446, N558, N795);
nand NAND2 (N847, N843, N602);
nor NOR4 (N848, N837, N41, N608, N168);
or OR2 (N849, N831, N696);
or OR2 (N850, N841, N96);
or OR3 (N851, N846, N537, N176);
not NOT1 (N852, N848);
not NOT1 (N853, N832);
nand NAND3 (N854, N851, N240, N785);
buf BUF1 (N855, N847);
buf BUF1 (N856, N854);
or OR3 (N857, N838, N258, N808);
buf BUF1 (N858, N853);
and AND4 (N859, N850, N743, N118, N587);
xor XOR2 (N860, N834, N514);
xor XOR2 (N861, N849, N746);
xor XOR2 (N862, N859, N281);
or OR4 (N863, N862, N375, N641, N670);
buf BUF1 (N864, N852);
nand NAND4 (N865, N858, N111, N183, N320);
buf BUF1 (N866, N857);
buf BUF1 (N867, N865);
not NOT1 (N868, N844);
nor NOR2 (N869, N855, N543);
or OR2 (N870, N845, N536);
nand NAND3 (N871, N869, N145, N365);
nor NOR3 (N872, N856, N6, N198);
buf BUF1 (N873, N867);
nand NAND2 (N874, N866, N641);
nand NAND3 (N875, N873, N122, N83);
nand NAND4 (N876, N871, N485, N752, N293);
not NOT1 (N877, N872);
not NOT1 (N878, N863);
buf BUF1 (N879, N874);
nand NAND2 (N880, N878, N791);
nor NOR4 (N881, N879, N248, N864, N609);
xor XOR2 (N882, N30, N269);
or OR3 (N883, N880, N633, N12);
nand NAND4 (N884, N876, N328, N315, N493);
xor XOR2 (N885, N861, N585);
buf BUF1 (N886, N881);
nand NAND2 (N887, N884, N800);
nand NAND2 (N888, N875, N700);
or OR3 (N889, N883, N879, N186);
xor XOR2 (N890, N887, N91);
not NOT1 (N891, N888);
nand NAND3 (N892, N885, N354, N874);
buf BUF1 (N893, N882);
xor XOR2 (N894, N890, N582);
and AND2 (N895, N886, N374);
and AND4 (N896, N889, N584, N449, N295);
not NOT1 (N897, N870);
buf BUF1 (N898, N868);
buf BUF1 (N899, N893);
or OR4 (N900, N897, N637, N571, N149);
and AND2 (N901, N860, N450);
nor NOR2 (N902, N895, N608);
nor NOR2 (N903, N900, N241);
and AND4 (N904, N902, N228, N805, N18);
nand NAND4 (N905, N898, N219, N501, N18);
nor NOR3 (N906, N905, N546, N100);
xor XOR2 (N907, N896, N762);
not NOT1 (N908, N907);
or OR4 (N909, N904, N17, N589, N579);
nor NOR2 (N910, N901, N755);
nand NAND2 (N911, N910, N753);
nor NOR2 (N912, N903, N131);
xor XOR2 (N913, N906, N518);
xor XOR2 (N914, N913, N569);
and AND3 (N915, N891, N841, N538);
nor NOR4 (N916, N894, N221, N680, N587);
buf BUF1 (N917, N909);
nand NAND3 (N918, N912, N884, N3);
xor XOR2 (N919, N916, N548);
not NOT1 (N920, N877);
nor NOR3 (N921, N917, N533, N671);
xor XOR2 (N922, N915, N557);
nand NAND3 (N923, N918, N502, N553);
xor XOR2 (N924, N920, N409);
nor NOR4 (N925, N919, N367, N760, N42);
nand NAND3 (N926, N914, N798, N498);
buf BUF1 (N927, N925);
not NOT1 (N928, N924);
nor NOR4 (N929, N911, N599, N540, N522);
nand NAND4 (N930, N921, N270, N103, N426);
nor NOR3 (N931, N928, N785, N662);
buf BUF1 (N932, N922);
xor XOR2 (N933, N892, N299);
and AND4 (N934, N908, N661, N832, N283);
or OR2 (N935, N933, N233);
xor XOR2 (N936, N935, N817);
buf BUF1 (N937, N899);
nor NOR3 (N938, N923, N605, N345);
and AND3 (N939, N927, N156, N88);
or OR4 (N940, N937, N131, N760, N125);
and AND2 (N941, N934, N626);
nor NOR2 (N942, N938, N614);
and AND3 (N943, N926, N277, N765);
not NOT1 (N944, N932);
not NOT1 (N945, N942);
not NOT1 (N946, N945);
nor NOR2 (N947, N941, N155);
buf BUF1 (N948, N940);
and AND4 (N949, N929, N451, N219, N684);
nand NAND4 (N950, N931, N516, N360, N329);
buf BUF1 (N951, N950);
xor XOR2 (N952, N930, N840);
xor XOR2 (N953, N951, N649);
nand NAND2 (N954, N949, N375);
not NOT1 (N955, N953);
or OR3 (N956, N936, N848, N125);
not NOT1 (N957, N948);
nand NAND3 (N958, N954, N254, N683);
nor NOR3 (N959, N939, N578, N500);
and AND3 (N960, N952, N453, N865);
not NOT1 (N961, N947);
and AND2 (N962, N960, N588);
nand NAND3 (N963, N959, N840, N631);
nor NOR3 (N964, N958, N620, N200);
nand NAND2 (N965, N957, N336);
nor NOR4 (N966, N963, N154, N90, N854);
and AND4 (N967, N965, N77, N122, N446);
or OR4 (N968, N964, N924, N572, N766);
not NOT1 (N969, N955);
nand NAND4 (N970, N967, N380, N502, N856);
or OR2 (N971, N969, N223);
or OR4 (N972, N944, N739, N322, N725);
xor XOR2 (N973, N943, N861);
xor XOR2 (N974, N956, N576);
or OR2 (N975, N961, N678);
or OR2 (N976, N962, N410);
nor NOR2 (N977, N946, N437);
nand NAND4 (N978, N976, N134, N879, N589);
not NOT1 (N979, N975);
or OR2 (N980, N979, N276);
buf BUF1 (N981, N973);
xor XOR2 (N982, N978, N689);
buf BUF1 (N983, N966);
xor XOR2 (N984, N981, N749);
nand NAND4 (N985, N971, N364, N297, N890);
xor XOR2 (N986, N972, N857);
nand NAND2 (N987, N974, N124);
nor NOR3 (N988, N970, N343, N488);
xor XOR2 (N989, N984, N314);
not NOT1 (N990, N977);
or OR4 (N991, N983, N196, N306, N877);
or OR3 (N992, N988, N96, N317);
or OR2 (N993, N990, N321);
not NOT1 (N994, N968);
buf BUF1 (N995, N994);
and AND2 (N996, N992, N439);
buf BUF1 (N997, N995);
buf BUF1 (N998, N987);
and AND3 (N999, N982, N413, N29);
not NOT1 (N1000, N989);
nor NOR3 (N1001, N986, N34, N399);
xor XOR2 (N1002, N997, N45);
not NOT1 (N1003, N991);
not NOT1 (N1004, N1002);
nor NOR2 (N1005, N985, N235);
nand NAND4 (N1006, N999, N278, N331, N362);
and AND3 (N1007, N980, N354, N789);
xor XOR2 (N1008, N993, N197);
xor XOR2 (N1009, N998, N178);
not NOT1 (N1010, N1004);
xor XOR2 (N1011, N1010, N655);
nor NOR4 (N1012, N1008, N147, N266, N679);
xor XOR2 (N1013, N996, N528);
or OR2 (N1014, N1007, N702);
not NOT1 (N1015, N1013);
xor XOR2 (N1016, N1012, N180);
not NOT1 (N1017, N1006);
and AND4 (N1018, N1005, N582, N101, N574);
xor XOR2 (N1019, N1009, N958);
and AND3 (N1020, N1003, N871, N137);
and AND3 (N1021, N1014, N779, N118);
and AND4 (N1022, N1011, N942, N48, N716);
nand NAND4 (N1023, N1001, N566, N755, N447);
and AND3 (N1024, N1016, N390, N159);
buf BUF1 (N1025, N1022);
not NOT1 (N1026, N1019);
xor XOR2 (N1027, N1024, N294);
nand NAND4 (N1028, N1017, N538, N940, N22);
or OR4 (N1029, N1020, N525, N5, N899);
nand NAND3 (N1030, N1023, N681, N292);
not NOT1 (N1031, N1025);
nand NAND2 (N1032, N1028, N24);
and AND4 (N1033, N1031, N173, N416, N458);
or OR4 (N1034, N1030, N565, N627, N204);
buf BUF1 (N1035, N1033);
buf BUF1 (N1036, N1015);
nand NAND2 (N1037, N1029, N126);
nor NOR3 (N1038, N1026, N986, N950);
nand NAND4 (N1039, N1027, N175, N119, N166);
and AND4 (N1040, N1038, N308, N363, N1032);
nand NAND3 (N1041, N593, N886, N736);
not NOT1 (N1042, N1040);
not NOT1 (N1043, N1035);
and AND4 (N1044, N1021, N219, N215, N564);
and AND3 (N1045, N1042, N640, N883);
buf BUF1 (N1046, N1045);
and AND4 (N1047, N1018, N336, N314, N761);
xor XOR2 (N1048, N1043, N1013);
and AND4 (N1049, N1037, N215, N1042, N13);
or OR4 (N1050, N1036, N232, N705, N829);
xor XOR2 (N1051, N1049, N868);
nor NOR2 (N1052, N1047, N757);
and AND4 (N1053, N1039, N612, N792, N692);
not NOT1 (N1054, N1052);
xor XOR2 (N1055, N1041, N885);
nor NOR4 (N1056, N1034, N567, N510, N987);
nand NAND3 (N1057, N1055, N980, N141);
not NOT1 (N1058, N1050);
nor NOR2 (N1059, N1051, N283);
not NOT1 (N1060, N1054);
buf BUF1 (N1061, N1000);
or OR4 (N1062, N1061, N278, N141, N895);
xor XOR2 (N1063, N1057, N384);
nand NAND4 (N1064, N1048, N267, N865, N548);
not NOT1 (N1065, N1046);
and AND3 (N1066, N1053, N394, N286);
xor XOR2 (N1067, N1063, N677);
and AND3 (N1068, N1059, N568, N194);
buf BUF1 (N1069, N1065);
buf BUF1 (N1070, N1066);
and AND3 (N1071, N1068, N656, N650);
nand NAND4 (N1072, N1064, N623, N1063, N106);
xor XOR2 (N1073, N1058, N309);
and AND3 (N1074, N1060, N73, N129);
or OR2 (N1075, N1073, N64);
buf BUF1 (N1076, N1062);
or OR4 (N1077, N1044, N1053, N269, N955);
xor XOR2 (N1078, N1075, N887);
not NOT1 (N1079, N1069);
nor NOR3 (N1080, N1076, N549, N851);
nand NAND4 (N1081, N1056, N168, N230, N829);
not NOT1 (N1082, N1072);
and AND3 (N1083, N1081, N990, N193);
nor NOR2 (N1084, N1070, N460);
or OR2 (N1085, N1067, N566);
or OR3 (N1086, N1085, N167, N732);
buf BUF1 (N1087, N1078);
not NOT1 (N1088, N1080);
and AND3 (N1089, N1074, N606, N792);
and AND4 (N1090, N1089, N620, N867, N654);
xor XOR2 (N1091, N1083, N931);
not NOT1 (N1092, N1079);
or OR3 (N1093, N1086, N847, N235);
xor XOR2 (N1094, N1077, N317);
xor XOR2 (N1095, N1087, N24);
and AND3 (N1096, N1091, N883, N665);
nor NOR4 (N1097, N1092, N548, N511, N187);
not NOT1 (N1098, N1096);
not NOT1 (N1099, N1082);
not NOT1 (N1100, N1071);
or OR4 (N1101, N1098, N1020, N560, N709);
nand NAND2 (N1102, N1100, N220);
or OR4 (N1103, N1094, N1049, N289, N688);
xor XOR2 (N1104, N1088, N440);
nand NAND4 (N1105, N1101, N313, N780, N609);
or OR2 (N1106, N1093, N965);
xor XOR2 (N1107, N1099, N141);
and AND3 (N1108, N1106, N101, N565);
buf BUF1 (N1109, N1084);
or OR3 (N1110, N1107, N280, N847);
nor NOR2 (N1111, N1095, N196);
nand NAND2 (N1112, N1090, N962);
buf BUF1 (N1113, N1105);
buf BUF1 (N1114, N1111);
nor NOR3 (N1115, N1114, N84, N599);
xor XOR2 (N1116, N1115, N124);
not NOT1 (N1117, N1103);
xor XOR2 (N1118, N1108, N506);
not NOT1 (N1119, N1104);
nor NOR2 (N1120, N1116, N1012);
and AND2 (N1121, N1097, N145);
or OR3 (N1122, N1113, N920, N1042);
nand NAND4 (N1123, N1121, N272, N493, N639);
not NOT1 (N1124, N1123);
nand NAND2 (N1125, N1119, N557);
nor NOR2 (N1126, N1112, N503);
not NOT1 (N1127, N1110);
not NOT1 (N1128, N1109);
and AND4 (N1129, N1128, N355, N644, N749);
nor NOR2 (N1130, N1120, N344);
buf BUF1 (N1131, N1102);
xor XOR2 (N1132, N1129, N683);
nor NOR2 (N1133, N1131, N563);
and AND4 (N1134, N1117, N594, N727, N508);
buf BUF1 (N1135, N1124);
nor NOR4 (N1136, N1132, N961, N1056, N1116);
and AND4 (N1137, N1133, N499, N1113, N893);
and AND2 (N1138, N1136, N736);
and AND4 (N1139, N1135, N449, N162, N1034);
not NOT1 (N1140, N1137);
or OR3 (N1141, N1140, N378, N230);
not NOT1 (N1142, N1122);
or OR2 (N1143, N1138, N560);
not NOT1 (N1144, N1143);
xor XOR2 (N1145, N1126, N545);
or OR3 (N1146, N1118, N737, N881);
nand NAND3 (N1147, N1125, N396, N378);
buf BUF1 (N1148, N1134);
nor NOR4 (N1149, N1141, N504, N46, N13);
nand NAND4 (N1150, N1148, N908, N1047, N202);
xor XOR2 (N1151, N1149, N585);
or OR4 (N1152, N1144, N867, N923, N1140);
nor NOR3 (N1153, N1152, N1023, N965);
xor XOR2 (N1154, N1139, N1002);
not NOT1 (N1155, N1130);
or OR3 (N1156, N1155, N78, N405);
or OR2 (N1157, N1150, N204);
buf BUF1 (N1158, N1142);
not NOT1 (N1159, N1154);
or OR3 (N1160, N1158, N926, N90);
not NOT1 (N1161, N1146);
or OR2 (N1162, N1153, N872);
not NOT1 (N1163, N1127);
nand NAND4 (N1164, N1163, N791, N309, N159);
and AND4 (N1165, N1145, N266, N1051, N93);
or OR3 (N1166, N1159, N947, N566);
nand NAND4 (N1167, N1165, N916, N998, N525);
or OR2 (N1168, N1147, N586);
not NOT1 (N1169, N1162);
and AND3 (N1170, N1151, N125, N502);
or OR4 (N1171, N1157, N843, N793, N666);
nor NOR2 (N1172, N1167, N869);
nor NOR4 (N1173, N1156, N1069, N411, N785);
or OR3 (N1174, N1164, N1030, N381);
buf BUF1 (N1175, N1170);
nor NOR2 (N1176, N1169, N11);
or OR3 (N1177, N1161, N658, N598);
nor NOR3 (N1178, N1160, N193, N541);
or OR2 (N1179, N1172, N629);
nand NAND3 (N1180, N1166, N716, N360);
buf BUF1 (N1181, N1175);
and AND2 (N1182, N1168, N1166);
and AND3 (N1183, N1181, N401, N1036);
not NOT1 (N1184, N1183);
nand NAND2 (N1185, N1173, N1141);
and AND2 (N1186, N1180, N609);
nand NAND2 (N1187, N1186, N227);
and AND4 (N1188, N1178, N977, N343, N883);
or OR4 (N1189, N1177, N961, N609, N81);
not NOT1 (N1190, N1187);
buf BUF1 (N1191, N1184);
not NOT1 (N1192, N1174);
not NOT1 (N1193, N1176);
not NOT1 (N1194, N1171);
and AND2 (N1195, N1191, N130);
buf BUF1 (N1196, N1190);
buf BUF1 (N1197, N1185);
buf BUF1 (N1198, N1179);
or OR2 (N1199, N1182, N767);
not NOT1 (N1200, N1194);
xor XOR2 (N1201, N1197, N921);
xor XOR2 (N1202, N1201, N490);
and AND3 (N1203, N1188, N293, N471);
not NOT1 (N1204, N1195);
buf BUF1 (N1205, N1202);
nand NAND2 (N1206, N1196, N1197);
not NOT1 (N1207, N1200);
nand NAND3 (N1208, N1192, N641, N200);
buf BUF1 (N1209, N1199);
nand NAND4 (N1210, N1203, N446, N95, N368);
nand NAND3 (N1211, N1189, N113, N686);
nand NAND3 (N1212, N1209, N547, N41);
or OR2 (N1213, N1205, N1211);
or OR4 (N1214, N882, N379, N457, N168);
buf BUF1 (N1215, N1204);
or OR2 (N1216, N1210, N263);
not NOT1 (N1217, N1213);
or OR2 (N1218, N1217, N121);
buf BUF1 (N1219, N1214);
buf BUF1 (N1220, N1208);
and AND2 (N1221, N1193, N291);
nand NAND2 (N1222, N1216, N1008);
or OR3 (N1223, N1220, N1161, N593);
nor NOR2 (N1224, N1222, N980);
and AND3 (N1225, N1215, N414, N97);
not NOT1 (N1226, N1219);
nand NAND4 (N1227, N1198, N854, N1016, N619);
and AND4 (N1228, N1207, N610, N195, N897);
nor NOR3 (N1229, N1221, N529, N988);
or OR4 (N1230, N1227, N1122, N749, N1172);
buf BUF1 (N1231, N1228);
not NOT1 (N1232, N1229);
nor NOR4 (N1233, N1212, N231, N353, N661);
buf BUF1 (N1234, N1223);
or OR3 (N1235, N1226, N416, N39);
buf BUF1 (N1236, N1218);
buf BUF1 (N1237, N1234);
nand NAND2 (N1238, N1231, N624);
or OR2 (N1239, N1225, N505);
buf BUF1 (N1240, N1238);
nand NAND4 (N1241, N1237, N637, N287, N707);
or OR3 (N1242, N1235, N512, N87);
not NOT1 (N1243, N1233);
nand NAND2 (N1244, N1243, N364);
buf BUF1 (N1245, N1206);
or OR2 (N1246, N1239, N856);
nor NOR4 (N1247, N1232, N864, N612, N110);
nor NOR2 (N1248, N1247, N771);
buf BUF1 (N1249, N1242);
buf BUF1 (N1250, N1246);
nor NOR2 (N1251, N1224, N373);
nor NOR3 (N1252, N1244, N484, N662);
or OR3 (N1253, N1251, N1246, N566);
or OR2 (N1254, N1241, N324);
nand NAND4 (N1255, N1254, N846, N379, N37);
buf BUF1 (N1256, N1230);
buf BUF1 (N1257, N1255);
not NOT1 (N1258, N1250);
buf BUF1 (N1259, N1258);
buf BUF1 (N1260, N1252);
buf BUF1 (N1261, N1260);
or OR4 (N1262, N1261, N880, N506, N705);
nand NAND4 (N1263, N1253, N837, N442, N738);
and AND2 (N1264, N1245, N1164);
buf BUF1 (N1265, N1262);
buf BUF1 (N1266, N1264);
and AND3 (N1267, N1263, N951, N1250);
buf BUF1 (N1268, N1249);
or OR4 (N1269, N1267, N1061, N511, N204);
not NOT1 (N1270, N1248);
nor NOR4 (N1271, N1240, N755, N884, N275);
nor NOR3 (N1272, N1270, N1116, N792);
nor NOR2 (N1273, N1266, N1008);
or OR4 (N1274, N1273, N1196, N243, N190);
nand NAND2 (N1275, N1257, N261);
xor XOR2 (N1276, N1271, N1051);
or OR4 (N1277, N1268, N1166, N19, N580);
not NOT1 (N1278, N1256);
buf BUF1 (N1279, N1236);
nor NOR4 (N1280, N1276, N161, N553, N467);
or OR4 (N1281, N1265, N507, N471, N729);
nand NAND3 (N1282, N1259, N521, N37);
and AND3 (N1283, N1281, N712, N493);
nor NOR2 (N1284, N1283, N514);
xor XOR2 (N1285, N1282, N690);
and AND4 (N1286, N1285, N722, N708, N732);
xor XOR2 (N1287, N1279, N943);
nand NAND3 (N1288, N1277, N619, N1255);
or OR2 (N1289, N1278, N139);
and AND4 (N1290, N1280, N1027, N775, N294);
nor NOR2 (N1291, N1286, N434);
nand NAND2 (N1292, N1287, N1082);
or OR2 (N1293, N1272, N1143);
xor XOR2 (N1294, N1288, N1262);
nor NOR2 (N1295, N1275, N1091);
and AND4 (N1296, N1284, N40, N658, N988);
and AND4 (N1297, N1290, N185, N495, N601);
nand NAND3 (N1298, N1293, N1179, N63);
nand NAND4 (N1299, N1292, N395, N1111, N270);
nor NOR4 (N1300, N1298, N945, N638, N1149);
nand NAND3 (N1301, N1295, N457, N173);
nor NOR2 (N1302, N1291, N104);
and AND3 (N1303, N1289, N887, N806);
buf BUF1 (N1304, N1301);
buf BUF1 (N1305, N1274);
nor NOR2 (N1306, N1303, N1290);
not NOT1 (N1307, N1269);
xor XOR2 (N1308, N1297, N1056);
nand NAND4 (N1309, N1299, N8, N54, N460);
xor XOR2 (N1310, N1304, N991);
and AND4 (N1311, N1294, N31, N1157, N934);
and AND3 (N1312, N1307, N89, N1127);
or OR2 (N1313, N1302, N144);
or OR2 (N1314, N1310, N1099);
not NOT1 (N1315, N1308);
and AND2 (N1316, N1311, N83);
or OR4 (N1317, N1316, N929, N670, N1118);
or OR2 (N1318, N1315, N778);
and AND3 (N1319, N1313, N207, N528);
not NOT1 (N1320, N1309);
buf BUF1 (N1321, N1312);
nand NAND4 (N1322, N1306, N237, N232, N497);
nor NOR4 (N1323, N1319, N135, N778, N871);
not NOT1 (N1324, N1314);
not NOT1 (N1325, N1305);
nand NAND4 (N1326, N1322, N194, N255, N1018);
not NOT1 (N1327, N1296);
nor NOR3 (N1328, N1318, N797, N859);
xor XOR2 (N1329, N1321, N375);
xor XOR2 (N1330, N1300, N1106);
nand NAND3 (N1331, N1326, N1147, N1100);
nor NOR4 (N1332, N1330, N495, N91, N1079);
or OR3 (N1333, N1331, N556, N725);
or OR2 (N1334, N1332, N250);
xor XOR2 (N1335, N1320, N1059);
nand NAND4 (N1336, N1327, N396, N1055, N1144);
nand NAND4 (N1337, N1333, N825, N351, N674);
buf BUF1 (N1338, N1323);
nand NAND4 (N1339, N1337, N522, N977, N1124);
xor XOR2 (N1340, N1325, N1089);
buf BUF1 (N1341, N1329);
nor NOR4 (N1342, N1341, N778, N942, N249);
nor NOR3 (N1343, N1317, N166, N130);
not NOT1 (N1344, N1342);
not NOT1 (N1345, N1336);
nor NOR2 (N1346, N1335, N906);
xor XOR2 (N1347, N1334, N549);
not NOT1 (N1348, N1339);
buf BUF1 (N1349, N1344);
and AND3 (N1350, N1349, N866, N1101);
nor NOR4 (N1351, N1328, N919, N802, N854);
or OR4 (N1352, N1324, N1011, N660, N901);
nor NOR2 (N1353, N1346, N1311);
nor NOR3 (N1354, N1351, N2, N1195);
or OR3 (N1355, N1343, N1350, N6);
xor XOR2 (N1356, N741, N171);
buf BUF1 (N1357, N1345);
or OR3 (N1358, N1352, N772, N357);
xor XOR2 (N1359, N1338, N292);
nor NOR2 (N1360, N1354, N143);
or OR4 (N1361, N1360, N1262, N863, N282);
nor NOR4 (N1362, N1358, N1119, N393, N428);
xor XOR2 (N1363, N1361, N9);
not NOT1 (N1364, N1340);
not NOT1 (N1365, N1363);
nor NOR3 (N1366, N1364, N422, N281);
xor XOR2 (N1367, N1357, N74);
buf BUF1 (N1368, N1362);
and AND4 (N1369, N1353, N1008, N734, N322);
not NOT1 (N1370, N1347);
not NOT1 (N1371, N1369);
not NOT1 (N1372, N1359);
nor NOR2 (N1373, N1371, N990);
nor NOR3 (N1374, N1365, N762, N39);
nor NOR2 (N1375, N1373, N1055);
buf BUF1 (N1376, N1355);
buf BUF1 (N1377, N1366);
nand NAND3 (N1378, N1370, N852, N1171);
buf BUF1 (N1379, N1378);
not NOT1 (N1380, N1375);
or OR3 (N1381, N1379, N86, N629);
nand NAND4 (N1382, N1381, N1067, N58, N1053);
xor XOR2 (N1383, N1377, N545);
nand NAND2 (N1384, N1382, N536);
nor NOR3 (N1385, N1372, N313, N1129);
xor XOR2 (N1386, N1384, N761);
buf BUF1 (N1387, N1376);
nor NOR4 (N1388, N1367, N336, N207, N13);
or OR3 (N1389, N1374, N525, N794);
or OR4 (N1390, N1388, N1113, N1099, N479);
nor NOR4 (N1391, N1386, N481, N578, N377);
nand NAND4 (N1392, N1391, N1124, N1237, N1382);
and AND4 (N1393, N1348, N247, N561, N1352);
nand NAND3 (N1394, N1380, N54, N117);
not NOT1 (N1395, N1393);
or OR3 (N1396, N1395, N244, N1313);
xor XOR2 (N1397, N1356, N285);
xor XOR2 (N1398, N1368, N254);
xor XOR2 (N1399, N1385, N408);
nor NOR4 (N1400, N1398, N904, N557, N588);
nand NAND2 (N1401, N1400, N894);
and AND4 (N1402, N1401, N462, N780, N568);
not NOT1 (N1403, N1399);
and AND4 (N1404, N1390, N1286, N794, N765);
nand NAND2 (N1405, N1396, N482);
xor XOR2 (N1406, N1394, N628);
and AND3 (N1407, N1387, N1179, N1340);
xor XOR2 (N1408, N1389, N553);
or OR3 (N1409, N1392, N1011, N163);
and AND3 (N1410, N1405, N909, N1322);
and AND2 (N1411, N1407, N524);
or OR3 (N1412, N1408, N270, N540);
or OR3 (N1413, N1404, N41, N40);
not NOT1 (N1414, N1411);
or OR2 (N1415, N1414, N684);
and AND4 (N1416, N1410, N1131, N290, N964);
nor NOR4 (N1417, N1403, N997, N580, N243);
and AND3 (N1418, N1397, N50, N597);
or OR4 (N1419, N1416, N688, N1188, N1013);
nand NAND2 (N1420, N1418, N323);
buf BUF1 (N1421, N1412);
not NOT1 (N1422, N1417);
or OR4 (N1423, N1415, N1264, N616, N859);
buf BUF1 (N1424, N1419);
buf BUF1 (N1425, N1423);
nor NOR3 (N1426, N1406, N940, N481);
and AND3 (N1427, N1424, N802, N236);
buf BUF1 (N1428, N1422);
not NOT1 (N1429, N1427);
xor XOR2 (N1430, N1429, N168);
and AND4 (N1431, N1428, N594, N439, N1253);
buf BUF1 (N1432, N1426);
and AND4 (N1433, N1420, N356, N989, N214);
xor XOR2 (N1434, N1433, N1228);
or OR3 (N1435, N1425, N1350, N1196);
xor XOR2 (N1436, N1431, N898);
or OR4 (N1437, N1430, N272, N205, N112);
not NOT1 (N1438, N1434);
nor NOR3 (N1439, N1437, N281, N1141);
nand NAND2 (N1440, N1432, N1059);
nor NOR3 (N1441, N1440, N918, N931);
and AND2 (N1442, N1383, N904);
and AND4 (N1443, N1435, N881, N352, N1080);
nor NOR3 (N1444, N1439, N236, N1405);
nand NAND4 (N1445, N1444, N907, N1201, N1164);
xor XOR2 (N1446, N1436, N908);
xor XOR2 (N1447, N1421, N571);
nor NOR3 (N1448, N1409, N1269, N973);
buf BUF1 (N1449, N1447);
and AND3 (N1450, N1442, N929, N1146);
or OR2 (N1451, N1413, N37);
or OR2 (N1452, N1451, N1023);
or OR3 (N1453, N1452, N42, N1202);
buf BUF1 (N1454, N1448);
not NOT1 (N1455, N1443);
buf BUF1 (N1456, N1402);
nand NAND4 (N1457, N1441, N439, N586, N402);
nor NOR2 (N1458, N1457, N1206);
or OR4 (N1459, N1455, N1107, N61, N821);
not NOT1 (N1460, N1445);
not NOT1 (N1461, N1460);
or OR4 (N1462, N1438, N962, N868, N597);
nor NOR2 (N1463, N1450, N594);
nor NOR4 (N1464, N1461, N1069, N275, N1300);
and AND3 (N1465, N1459, N33, N83);
xor XOR2 (N1466, N1464, N530);
and AND2 (N1467, N1453, N1357);
buf BUF1 (N1468, N1463);
and AND4 (N1469, N1456, N862, N920, N1334);
buf BUF1 (N1470, N1465);
nor NOR3 (N1471, N1470, N29, N60);
buf BUF1 (N1472, N1471);
nor NOR3 (N1473, N1472, N1168, N38);
or OR2 (N1474, N1462, N1384);
nand NAND4 (N1475, N1446, N727, N745, N434);
xor XOR2 (N1476, N1449, N1126);
or OR2 (N1477, N1468, N101);
buf BUF1 (N1478, N1458);
not NOT1 (N1479, N1474);
nor NOR3 (N1480, N1469, N615, N166);
not NOT1 (N1481, N1454);
and AND4 (N1482, N1467, N1170, N431, N1136);
xor XOR2 (N1483, N1476, N132);
not NOT1 (N1484, N1466);
buf BUF1 (N1485, N1481);
and AND4 (N1486, N1484, N721, N200, N883);
or OR2 (N1487, N1483, N543);
nor NOR4 (N1488, N1486, N974, N88, N547);
nand NAND3 (N1489, N1477, N119, N1276);
buf BUF1 (N1490, N1479);
and AND3 (N1491, N1478, N1064, N1171);
or OR2 (N1492, N1475, N1294);
nor NOR4 (N1493, N1492, N652, N1358, N318);
or OR3 (N1494, N1485, N777, N1117);
xor XOR2 (N1495, N1487, N354);
and AND3 (N1496, N1495, N915, N737);
buf BUF1 (N1497, N1480);
buf BUF1 (N1498, N1482);
nand NAND4 (N1499, N1493, N819, N872, N877);
and AND2 (N1500, N1498, N681);
nor NOR4 (N1501, N1473, N342, N772, N18);
or OR3 (N1502, N1490, N806, N605);
or OR3 (N1503, N1499, N153, N993);
buf BUF1 (N1504, N1503);
not NOT1 (N1505, N1489);
or OR4 (N1506, N1504, N646, N69, N840);
nand NAND4 (N1507, N1497, N297, N1288, N157);
buf BUF1 (N1508, N1488);
buf BUF1 (N1509, N1496);
nor NOR4 (N1510, N1507, N751, N1172, N867);
not NOT1 (N1511, N1494);
nand NAND4 (N1512, N1511, N384, N850, N1403);
and AND3 (N1513, N1510, N1398, N758);
nand NAND3 (N1514, N1501, N317, N1046);
nand NAND2 (N1515, N1513, N668);
or OR4 (N1516, N1512, N1154, N778, N135);
not NOT1 (N1517, N1514);
xor XOR2 (N1518, N1509, N1363);
nand NAND3 (N1519, N1508, N1412, N923);
not NOT1 (N1520, N1517);
or OR2 (N1521, N1500, N543);
nor NOR2 (N1522, N1516, N404);
nor NOR2 (N1523, N1502, N82);
or OR3 (N1524, N1521, N1131, N1049);
nor NOR3 (N1525, N1518, N570, N1097);
not NOT1 (N1526, N1524);
not NOT1 (N1527, N1505);
xor XOR2 (N1528, N1491, N1242);
nand NAND2 (N1529, N1528, N549);
nand NAND4 (N1530, N1526, N728, N122, N677);
buf BUF1 (N1531, N1523);
not NOT1 (N1532, N1530);
nor NOR2 (N1533, N1532, N1200);
nand NAND2 (N1534, N1529, N712);
xor XOR2 (N1535, N1531, N34);
and AND4 (N1536, N1535, N1505, N1209, N164);
nand NAND4 (N1537, N1515, N1422, N1034, N829);
nand NAND3 (N1538, N1527, N1322, N776);
nand NAND3 (N1539, N1533, N809, N95);
nor NOR2 (N1540, N1519, N653);
or OR4 (N1541, N1537, N1234, N969, N1266);
or OR2 (N1542, N1540, N283);
nor NOR2 (N1543, N1522, N522);
not NOT1 (N1544, N1536);
nand NAND3 (N1545, N1506, N592, N459);
nor NOR4 (N1546, N1534, N361, N429, N435);
xor XOR2 (N1547, N1544, N1115);
nor NOR2 (N1548, N1543, N270);
nor NOR2 (N1549, N1546, N301);
not NOT1 (N1550, N1542);
buf BUF1 (N1551, N1545);
nand NAND3 (N1552, N1525, N738, N99);
or OR3 (N1553, N1550, N133, N939);
or OR3 (N1554, N1549, N1326, N1346);
nor NOR4 (N1555, N1554, N437, N1380, N1018);
xor XOR2 (N1556, N1547, N948);
not NOT1 (N1557, N1548);
and AND4 (N1558, N1552, N1254, N714, N1236);
and AND3 (N1559, N1558, N1031, N602);
not NOT1 (N1560, N1556);
xor XOR2 (N1561, N1560, N17);
and AND4 (N1562, N1520, N238, N287, N1311);
not NOT1 (N1563, N1553);
not NOT1 (N1564, N1559);
nor NOR2 (N1565, N1539, N952);
xor XOR2 (N1566, N1538, N1380);
buf BUF1 (N1567, N1564);
xor XOR2 (N1568, N1557, N1107);
nand NAND3 (N1569, N1562, N181, N369);
nand NAND2 (N1570, N1551, N611);
and AND4 (N1571, N1563, N519, N1051, N513);
xor XOR2 (N1572, N1568, N456);
xor XOR2 (N1573, N1570, N1336);
xor XOR2 (N1574, N1572, N13);
xor XOR2 (N1575, N1567, N715);
or OR2 (N1576, N1573, N551);
or OR2 (N1577, N1555, N1395);
buf BUF1 (N1578, N1541);
not NOT1 (N1579, N1565);
not NOT1 (N1580, N1571);
nor NOR4 (N1581, N1561, N217, N235, N836);
not NOT1 (N1582, N1578);
and AND4 (N1583, N1580, N988, N1383, N129);
and AND2 (N1584, N1569, N776);
buf BUF1 (N1585, N1576);
nand NAND2 (N1586, N1585, N1496);
buf BUF1 (N1587, N1575);
or OR4 (N1588, N1586, N843, N1212, N469);
nor NOR2 (N1589, N1581, N39);
nand NAND2 (N1590, N1579, N563);
and AND2 (N1591, N1590, N886);
not NOT1 (N1592, N1566);
xor XOR2 (N1593, N1587, N1115);
buf BUF1 (N1594, N1574);
nand NAND2 (N1595, N1589, N156);
nor NOR4 (N1596, N1584, N926, N1464, N302);
buf BUF1 (N1597, N1596);
or OR2 (N1598, N1594, N915);
not NOT1 (N1599, N1577);
and AND2 (N1600, N1583, N1003);
and AND2 (N1601, N1591, N239);
and AND4 (N1602, N1599, N304, N801, N1213);
or OR3 (N1603, N1600, N1054, N1152);
and AND2 (N1604, N1598, N1337);
xor XOR2 (N1605, N1595, N815);
buf BUF1 (N1606, N1601);
buf BUF1 (N1607, N1604);
and AND4 (N1608, N1588, N1122, N330, N1096);
xor XOR2 (N1609, N1605, N401);
xor XOR2 (N1610, N1603, N1281);
nand NAND3 (N1611, N1597, N515, N1487);
or OR2 (N1612, N1592, N912);
buf BUF1 (N1613, N1608);
or OR4 (N1614, N1593, N301, N561, N1274);
not NOT1 (N1615, N1611);
nor NOR3 (N1616, N1613, N1328, N904);
nor NOR4 (N1617, N1582, N162, N193, N728);
nand NAND3 (N1618, N1614, N1489, N15);
not NOT1 (N1619, N1609);
nand NAND2 (N1620, N1607, N1490);
buf BUF1 (N1621, N1620);
xor XOR2 (N1622, N1615, N1177);
buf BUF1 (N1623, N1622);
and AND2 (N1624, N1616, N786);
xor XOR2 (N1625, N1618, N1096);
nand NAND3 (N1626, N1623, N363, N1111);
not NOT1 (N1627, N1625);
nor NOR2 (N1628, N1602, N911);
and AND3 (N1629, N1626, N817, N797);
nand NAND2 (N1630, N1627, N92);
buf BUF1 (N1631, N1628);
xor XOR2 (N1632, N1629, N784);
and AND4 (N1633, N1610, N1322, N583, N643);
nor NOR4 (N1634, N1617, N516, N744, N1170);
xor XOR2 (N1635, N1606, N376);
or OR4 (N1636, N1634, N1564, N1049, N513);
buf BUF1 (N1637, N1633);
or OR3 (N1638, N1621, N792, N540);
and AND2 (N1639, N1619, N282);
or OR3 (N1640, N1637, N165, N247);
xor XOR2 (N1641, N1624, N1411);
xor XOR2 (N1642, N1640, N1575);
xor XOR2 (N1643, N1641, N1280);
not NOT1 (N1644, N1631);
xor XOR2 (N1645, N1642, N502);
or OR3 (N1646, N1639, N170, N1147);
and AND2 (N1647, N1638, N878);
buf BUF1 (N1648, N1632);
or OR3 (N1649, N1644, N285, N1570);
xor XOR2 (N1650, N1630, N27);
and AND3 (N1651, N1635, N1403, N272);
not NOT1 (N1652, N1646);
nand NAND4 (N1653, N1647, N1452, N226, N1134);
buf BUF1 (N1654, N1645);
xor XOR2 (N1655, N1649, N1150);
and AND2 (N1656, N1654, N1500);
and AND3 (N1657, N1652, N1209, N1000);
buf BUF1 (N1658, N1612);
not NOT1 (N1659, N1636);
not NOT1 (N1660, N1656);
nor NOR4 (N1661, N1643, N1119, N1565, N178);
or OR2 (N1662, N1657, N307);
xor XOR2 (N1663, N1662, N448);
not NOT1 (N1664, N1663);
buf BUF1 (N1665, N1648);
nor NOR4 (N1666, N1658, N1016, N897, N1520);
and AND4 (N1667, N1664, N374, N420, N1169);
not NOT1 (N1668, N1655);
nand NAND3 (N1669, N1667, N242, N414);
xor XOR2 (N1670, N1650, N1623);
xor XOR2 (N1671, N1669, N33);
nor NOR2 (N1672, N1660, N146);
not NOT1 (N1673, N1653);
or OR4 (N1674, N1659, N1416, N1547, N159);
not NOT1 (N1675, N1668);
not NOT1 (N1676, N1665);
not NOT1 (N1677, N1666);
not NOT1 (N1678, N1670);
xor XOR2 (N1679, N1674, N716);
xor XOR2 (N1680, N1672, N1457);
and AND4 (N1681, N1651, N225, N615, N450);
not NOT1 (N1682, N1673);
xor XOR2 (N1683, N1675, N50);
or OR2 (N1684, N1680, N1154);
not NOT1 (N1685, N1681);
buf BUF1 (N1686, N1684);
nand NAND4 (N1687, N1685, N673, N663, N1578);
nand NAND3 (N1688, N1676, N1254, N956);
nand NAND4 (N1689, N1678, N1175, N1072, N941);
not NOT1 (N1690, N1689);
xor XOR2 (N1691, N1688, N1268);
not NOT1 (N1692, N1661);
or OR2 (N1693, N1686, N1527);
or OR3 (N1694, N1690, N666, N1033);
buf BUF1 (N1695, N1683);
nor NOR2 (N1696, N1679, N882);
buf BUF1 (N1697, N1677);
nand NAND2 (N1698, N1695, N590);
xor XOR2 (N1699, N1687, N1518);
not NOT1 (N1700, N1697);
nor NOR2 (N1701, N1700, N1233);
nor NOR4 (N1702, N1682, N1290, N1436, N983);
nand NAND4 (N1703, N1693, N1280, N1629, N37);
or OR2 (N1704, N1671, N1624);
and AND4 (N1705, N1702, N1326, N1606, N170);
nor NOR2 (N1706, N1691, N63);
nor NOR3 (N1707, N1698, N181, N1587);
xor XOR2 (N1708, N1704, N233);
and AND4 (N1709, N1708, N1424, N998, N1047);
and AND2 (N1710, N1699, N691);
nor NOR2 (N1711, N1692, N994);
xor XOR2 (N1712, N1711, N133);
and AND3 (N1713, N1705, N253, N456);
nand NAND4 (N1714, N1712, N1030, N1432, N1396);
and AND2 (N1715, N1713, N658);
and AND3 (N1716, N1707, N269, N1594);
not NOT1 (N1717, N1706);
xor XOR2 (N1718, N1710, N1188);
and AND2 (N1719, N1715, N330);
buf BUF1 (N1720, N1719);
buf BUF1 (N1721, N1696);
or OR2 (N1722, N1720, N319);
or OR2 (N1723, N1694, N1056);
nor NOR4 (N1724, N1701, N1305, N642, N890);
buf BUF1 (N1725, N1717);
not NOT1 (N1726, N1723);
buf BUF1 (N1727, N1709);
and AND2 (N1728, N1703, N750);
and AND2 (N1729, N1726, N1456);
or OR2 (N1730, N1718, N970);
nand NAND2 (N1731, N1722, N1308);
nor NOR4 (N1732, N1731, N717, N1124, N845);
nand NAND4 (N1733, N1729, N1553, N831, N513);
nand NAND2 (N1734, N1724, N263);
or OR2 (N1735, N1714, N814);
xor XOR2 (N1736, N1733, N456);
nor NOR2 (N1737, N1716, N600);
xor XOR2 (N1738, N1735, N281);
xor XOR2 (N1739, N1728, N1687);
xor XOR2 (N1740, N1732, N12);
not NOT1 (N1741, N1734);
not NOT1 (N1742, N1739);
nand NAND2 (N1743, N1740, N1230);
not NOT1 (N1744, N1730);
buf BUF1 (N1745, N1744);
not NOT1 (N1746, N1745);
and AND4 (N1747, N1743, N1576, N1742, N598);
or OR3 (N1748, N776, N319, N70);
not NOT1 (N1749, N1725);
nor NOR3 (N1750, N1727, N1586, N1395);
and AND2 (N1751, N1749, N396);
nor NOR3 (N1752, N1737, N1579, N837);
buf BUF1 (N1753, N1721);
buf BUF1 (N1754, N1738);
nor NOR3 (N1755, N1747, N937, N1624);
nand NAND4 (N1756, N1755, N1703, N1337, N168);
or OR2 (N1757, N1750, N745);
buf BUF1 (N1758, N1754);
and AND3 (N1759, N1756, N591, N722);
buf BUF1 (N1760, N1758);
not NOT1 (N1761, N1759);
or OR4 (N1762, N1736, N1544, N860, N508);
nand NAND2 (N1763, N1748, N1305);
and AND2 (N1764, N1761, N85);
xor XOR2 (N1765, N1760, N1141);
and AND3 (N1766, N1751, N1765, N1752);
nor NOR3 (N1767, N1663, N970, N952);
nor NOR2 (N1768, N884, N507);
nand NAND3 (N1769, N1762, N1074, N25);
not NOT1 (N1770, N1767);
and AND4 (N1771, N1757, N1693, N742, N1097);
or OR2 (N1772, N1771, N709);
not NOT1 (N1773, N1741);
nor NOR4 (N1774, N1764, N54, N16, N692);
and AND3 (N1775, N1763, N258, N362);
nand NAND4 (N1776, N1770, N313, N1767, N577);
and AND4 (N1777, N1746, N1539, N963, N1773);
xor XOR2 (N1778, N655, N873);
not NOT1 (N1779, N1769);
or OR2 (N1780, N1775, N716);
or OR3 (N1781, N1753, N703, N1708);
buf BUF1 (N1782, N1781);
or OR4 (N1783, N1768, N606, N1584, N1150);
not NOT1 (N1784, N1774);
not NOT1 (N1785, N1779);
nor NOR2 (N1786, N1777, N169);
buf BUF1 (N1787, N1782);
nand NAND4 (N1788, N1787, N1301, N792, N542);
nand NAND3 (N1789, N1780, N232, N1446);
nor NOR2 (N1790, N1786, N1635);
or OR2 (N1791, N1772, N405);
or OR4 (N1792, N1783, N84, N1657, N900);
buf BUF1 (N1793, N1785);
nand NAND4 (N1794, N1776, N293, N1380, N92);
or OR2 (N1795, N1793, N13);
or OR3 (N1796, N1789, N679, N825);
nand NAND3 (N1797, N1796, N1635, N1157);
buf BUF1 (N1798, N1791);
or OR4 (N1799, N1790, N1106, N1734, N45);
not NOT1 (N1800, N1799);
and AND2 (N1801, N1778, N458);
and AND4 (N1802, N1794, N412, N477, N1428);
buf BUF1 (N1803, N1792);
nand NAND3 (N1804, N1803, N1036, N51);
nand NAND4 (N1805, N1801, N1231, N1578, N364);
or OR3 (N1806, N1802, N803, N517);
and AND2 (N1807, N1795, N1028);
buf BUF1 (N1808, N1807);
buf BUF1 (N1809, N1798);
and AND3 (N1810, N1788, N156, N388);
nand NAND4 (N1811, N1797, N1461, N504, N1648);
buf BUF1 (N1812, N1811);
buf BUF1 (N1813, N1784);
buf BUF1 (N1814, N1813);
or OR4 (N1815, N1809, N1712, N1382, N1167);
or OR3 (N1816, N1805, N1781, N1671);
nor NOR4 (N1817, N1808, N1267, N407, N342);
nor NOR2 (N1818, N1800, N848);
buf BUF1 (N1819, N1816);
and AND4 (N1820, N1812, N1455, N838, N1279);
buf BUF1 (N1821, N1815);
xor XOR2 (N1822, N1766, N1406);
not NOT1 (N1823, N1810);
nor NOR3 (N1824, N1817, N738, N1064);
nand NAND4 (N1825, N1822, N798, N1759, N1469);
buf BUF1 (N1826, N1814);
xor XOR2 (N1827, N1821, N104);
nand NAND3 (N1828, N1818, N1095, N1512);
or OR2 (N1829, N1823, N460);
and AND2 (N1830, N1828, N642);
and AND3 (N1831, N1826, N1147, N1758);
nand NAND3 (N1832, N1824, N1723, N787);
nand NAND4 (N1833, N1827, N237, N1184, N920);
not NOT1 (N1834, N1819);
nand NAND2 (N1835, N1825, N783);
buf BUF1 (N1836, N1834);
and AND4 (N1837, N1829, N134, N823, N1068);
or OR2 (N1838, N1831, N1385);
xor XOR2 (N1839, N1804, N1273);
or OR4 (N1840, N1835, N1066, N843, N1687);
not NOT1 (N1841, N1830);
xor XOR2 (N1842, N1806, N1546);
nor NOR2 (N1843, N1839, N1739);
not NOT1 (N1844, N1820);
buf BUF1 (N1845, N1841);
and AND3 (N1846, N1836, N1768, N784);
xor XOR2 (N1847, N1842, N639);
nand NAND4 (N1848, N1837, N1463, N519, N516);
and AND4 (N1849, N1845, N972, N512, N1022);
not NOT1 (N1850, N1838);
nor NOR3 (N1851, N1843, N1161, N372);
nand NAND4 (N1852, N1847, N1276, N806, N884);
or OR4 (N1853, N1851, N390, N466, N977);
and AND2 (N1854, N1832, N885);
not NOT1 (N1855, N1844);
nand NAND3 (N1856, N1854, N1492, N1735);
not NOT1 (N1857, N1855);
nand NAND4 (N1858, N1846, N223, N768, N1010);
or OR4 (N1859, N1853, N879, N141, N1275);
xor XOR2 (N1860, N1840, N1311);
xor XOR2 (N1861, N1857, N354);
xor XOR2 (N1862, N1852, N1358);
nor NOR4 (N1863, N1862, N828, N682, N657);
or OR4 (N1864, N1849, N1326, N564, N1434);
nor NOR3 (N1865, N1861, N1196, N1611);
not NOT1 (N1866, N1859);
and AND4 (N1867, N1850, N81, N1070, N1743);
xor XOR2 (N1868, N1856, N1167);
xor XOR2 (N1869, N1867, N602);
nor NOR4 (N1870, N1865, N230, N1418, N56);
nor NOR3 (N1871, N1866, N979, N1144);
nand NAND3 (N1872, N1864, N1054, N795);
or OR4 (N1873, N1860, N421, N264, N903);
and AND2 (N1874, N1870, N517);
nor NOR3 (N1875, N1863, N456, N49);
nor NOR2 (N1876, N1868, N1174);
and AND2 (N1877, N1872, N1118);
and AND4 (N1878, N1871, N458, N1335, N1487);
nand NAND3 (N1879, N1876, N1205, N314);
buf BUF1 (N1880, N1874);
and AND2 (N1881, N1869, N1774);
buf BUF1 (N1882, N1879);
nand NAND3 (N1883, N1848, N1238, N1156);
buf BUF1 (N1884, N1878);
xor XOR2 (N1885, N1877, N1660);
nor NOR3 (N1886, N1882, N634, N508);
not NOT1 (N1887, N1875);
not NOT1 (N1888, N1887);
not NOT1 (N1889, N1883);
xor XOR2 (N1890, N1881, N1332);
and AND3 (N1891, N1886, N881, N962);
xor XOR2 (N1892, N1873, N1173);
or OR3 (N1893, N1858, N846, N1754);
buf BUF1 (N1894, N1889);
nor NOR4 (N1895, N1880, N467, N1350, N1675);
nand NAND4 (N1896, N1891, N31, N1154, N39);
or OR3 (N1897, N1833, N172, N939);
or OR4 (N1898, N1885, N1875, N301, N1626);
nor NOR4 (N1899, N1894, N12, N368, N1867);
nand NAND4 (N1900, N1896, N703, N972, N421);
not NOT1 (N1901, N1898);
not NOT1 (N1902, N1884);
xor XOR2 (N1903, N1900, N1253);
xor XOR2 (N1904, N1901, N157);
buf BUF1 (N1905, N1899);
xor XOR2 (N1906, N1895, N273);
nor NOR2 (N1907, N1905, N283);
xor XOR2 (N1908, N1892, N918);
xor XOR2 (N1909, N1906, N286);
nor NOR3 (N1910, N1890, N841, N769);
not NOT1 (N1911, N1910);
or OR4 (N1912, N1911, N12, N1253, N718);
or OR3 (N1913, N1902, N504, N846);
buf BUF1 (N1914, N1897);
nand NAND4 (N1915, N1893, N1557, N778, N320);
and AND4 (N1916, N1913, N576, N778, N869);
not NOT1 (N1917, N1907);
xor XOR2 (N1918, N1888, N993);
or OR4 (N1919, N1904, N1542, N1027, N409);
or OR3 (N1920, N1916, N55, N1172);
and AND4 (N1921, N1909, N1206, N895, N1410);
xor XOR2 (N1922, N1915, N395);
and AND4 (N1923, N1917, N1133, N1071, N97);
nor NOR2 (N1924, N1922, N747);
buf BUF1 (N1925, N1914);
nand NAND4 (N1926, N1918, N1099, N1797, N742);
and AND3 (N1927, N1924, N1178, N276);
or OR2 (N1928, N1912, N1903);
buf BUF1 (N1929, N1248);
not NOT1 (N1930, N1928);
and AND2 (N1931, N1926, N424);
and AND3 (N1932, N1930, N974, N799);
nand NAND3 (N1933, N1927, N1135, N1904);
nand NAND4 (N1934, N1929, N869, N1788, N1379);
nand NAND4 (N1935, N1921, N1223, N118, N1193);
xor XOR2 (N1936, N1932, N1448);
buf BUF1 (N1937, N1935);
not NOT1 (N1938, N1933);
buf BUF1 (N1939, N1908);
nor NOR3 (N1940, N1925, N50, N396);
buf BUF1 (N1941, N1934);
nor NOR3 (N1942, N1940, N379, N1728);
nor NOR2 (N1943, N1942, N1338);
nand NAND3 (N1944, N1936, N1271, N1114);
nor NOR4 (N1945, N1920, N1905, N290, N666);
or OR3 (N1946, N1923, N1890, N1864);
not NOT1 (N1947, N1938);
nor NOR2 (N1948, N1937, N1248);
buf BUF1 (N1949, N1939);
and AND4 (N1950, N1948, N35, N1137, N754);
xor XOR2 (N1951, N1931, N655);
xor XOR2 (N1952, N1946, N1491);
nand NAND2 (N1953, N1952, N1260);
xor XOR2 (N1954, N1953, N691);
or OR4 (N1955, N1949, N1474, N625, N1728);
buf BUF1 (N1956, N1955);
nor NOR3 (N1957, N1945, N1003, N67);
and AND2 (N1958, N1947, N830);
and AND4 (N1959, N1954, N459, N1448, N1534);
nand NAND2 (N1960, N1959, N692);
nand NAND4 (N1961, N1951, N3, N78, N1479);
nand NAND2 (N1962, N1950, N1701);
nor NOR4 (N1963, N1956, N1317, N861, N1904);
not NOT1 (N1964, N1960);
buf BUF1 (N1965, N1962);
buf BUF1 (N1966, N1965);
xor XOR2 (N1967, N1957, N1825);
nand NAND3 (N1968, N1966, N880, N1861);
xor XOR2 (N1969, N1964, N935);
nor NOR3 (N1970, N1961, N377, N1518);
nand NAND3 (N1971, N1967, N78, N1326);
not NOT1 (N1972, N1963);
buf BUF1 (N1973, N1970);
not NOT1 (N1974, N1969);
xor XOR2 (N1975, N1974, N640);
nor NOR3 (N1976, N1944, N740, N1152);
and AND3 (N1977, N1976, N3, N770);
and AND2 (N1978, N1919, N1630);
xor XOR2 (N1979, N1977, N1019);
nor NOR4 (N1980, N1943, N563, N434, N1501);
xor XOR2 (N1981, N1971, N1610);
and AND2 (N1982, N1968, N1829);
and AND2 (N1983, N1981, N58);
not NOT1 (N1984, N1983);
not NOT1 (N1985, N1984);
not NOT1 (N1986, N1972);
and AND2 (N1987, N1973, N867);
or OR2 (N1988, N1978, N1827);
or OR2 (N1989, N1988, N1382);
buf BUF1 (N1990, N1986);
nor NOR4 (N1991, N1980, N38, N343, N1223);
xor XOR2 (N1992, N1975, N119);
or OR2 (N1993, N1990, N699);
or OR2 (N1994, N1991, N1423);
buf BUF1 (N1995, N1982);
buf BUF1 (N1996, N1995);
or OR3 (N1997, N1979, N1773, N937);
xor XOR2 (N1998, N1987, N15);
buf BUF1 (N1999, N1989);
xor XOR2 (N2000, N1993, N1043);
and AND4 (N2001, N1992, N1971, N723, N454);
nor NOR3 (N2002, N1996, N1481, N187);
not NOT1 (N2003, N1999);
and AND3 (N2004, N1941, N1997, N540);
nor NOR3 (N2005, N120, N533, N1606);
buf BUF1 (N2006, N2004);
or OR4 (N2007, N2003, N1512, N1541, N483);
and AND2 (N2008, N2006, N1958);
nor NOR3 (N2009, N225, N76, N432);
nor NOR3 (N2010, N2000, N1100, N2007);
and AND4 (N2011, N163, N307, N1560, N346);
xor XOR2 (N2012, N2001, N939);
nand NAND4 (N2013, N2010, N403, N1471, N1495);
not NOT1 (N2014, N2012);
xor XOR2 (N2015, N1994, N145);
nand NAND3 (N2016, N2002, N114, N1669);
not NOT1 (N2017, N2009);
nor NOR2 (N2018, N2016, N436);
not NOT1 (N2019, N2008);
or OR4 (N2020, N1998, N124, N1386, N1968);
or OR4 (N2021, N1985, N1306, N226, N420);
xor XOR2 (N2022, N2014, N1825);
not NOT1 (N2023, N2022);
not NOT1 (N2024, N2005);
buf BUF1 (N2025, N2018);
and AND4 (N2026, N2013, N1444, N278, N1251);
and AND2 (N2027, N2017, N1496);
or OR3 (N2028, N2026, N522, N1960);
and AND2 (N2029, N2015, N390);
buf BUF1 (N2030, N2029);
buf BUF1 (N2031, N2028);
nor NOR3 (N2032, N2024, N946, N1793);
or OR3 (N2033, N2023, N394, N1369);
or OR2 (N2034, N2030, N587);
nand NAND2 (N2035, N2020, N442);
nand NAND3 (N2036, N2034, N1078, N650);
not NOT1 (N2037, N2032);
and AND4 (N2038, N2027, N666, N1680, N1681);
nor NOR2 (N2039, N2033, N657);
nand NAND2 (N2040, N2021, N1257);
buf BUF1 (N2041, N2039);
buf BUF1 (N2042, N2040);
xor XOR2 (N2043, N2041, N238);
xor XOR2 (N2044, N2025, N964);
buf BUF1 (N2045, N2019);
buf BUF1 (N2046, N2038);
and AND3 (N2047, N2031, N1301, N954);
nor NOR3 (N2048, N2036, N924, N1012);
and AND4 (N2049, N2044, N1643, N1716, N1501);
xor XOR2 (N2050, N2035, N228);
nand NAND4 (N2051, N2043, N602, N550, N1989);
nor NOR3 (N2052, N2045, N1686, N1338);
nand NAND2 (N2053, N2052, N284);
and AND3 (N2054, N2042, N1750, N346);
buf BUF1 (N2055, N2053);
not NOT1 (N2056, N2047);
or OR2 (N2057, N2049, N1901);
xor XOR2 (N2058, N2050, N35);
nand NAND4 (N2059, N2046, N1856, N1306, N576);
or OR4 (N2060, N2037, N347, N45, N1444);
nand NAND4 (N2061, N2011, N1156, N604, N1045);
nand NAND2 (N2062, N2061, N1256);
nand NAND3 (N2063, N2060, N587, N1678);
not NOT1 (N2064, N2048);
or OR3 (N2065, N2063, N1251, N299);
or OR3 (N2066, N2059, N1176, N1001);
nor NOR3 (N2067, N2065, N719, N186);
nand NAND3 (N2068, N2064, N460, N1603);
nor NOR3 (N2069, N2066, N1213, N1851);
xor XOR2 (N2070, N2069, N598);
and AND4 (N2071, N2057, N1048, N996, N1280);
not NOT1 (N2072, N2070);
buf BUF1 (N2073, N2068);
nor NOR4 (N2074, N2073, N140, N854, N715);
not NOT1 (N2075, N2067);
xor XOR2 (N2076, N2072, N171);
buf BUF1 (N2077, N2075);
not NOT1 (N2078, N2054);
not NOT1 (N2079, N2062);
buf BUF1 (N2080, N2077);
buf BUF1 (N2081, N2058);
nand NAND4 (N2082, N2071, N1809, N826, N1340);
or OR4 (N2083, N2082, N1325, N910, N748);
and AND4 (N2084, N2079, N977, N143, N681);
xor XOR2 (N2085, N2056, N1965);
nand NAND2 (N2086, N2074, N758);
and AND4 (N2087, N2051, N1257, N121, N1442);
nor NOR4 (N2088, N2078, N1400, N643, N2001);
nor NOR4 (N2089, N2055, N1608, N512, N1985);
buf BUF1 (N2090, N2080);
and AND2 (N2091, N2088, N1568);
buf BUF1 (N2092, N2085);
not NOT1 (N2093, N2076);
and AND2 (N2094, N2081, N1298);
buf BUF1 (N2095, N2093);
xor XOR2 (N2096, N2091, N914);
xor XOR2 (N2097, N2094, N1030);
or OR3 (N2098, N2097, N383, N1477);
nor NOR4 (N2099, N2083, N509, N1015, N556);
xor XOR2 (N2100, N2098, N873);
or OR2 (N2101, N2095, N1841);
not NOT1 (N2102, N2089);
and AND2 (N2103, N2086, N1197);
nand NAND4 (N2104, N2084, N748, N944, N968);
not NOT1 (N2105, N2101);
or OR3 (N2106, N2099, N2034, N1686);
buf BUF1 (N2107, N2104);
nor NOR4 (N2108, N2092, N147, N893, N1451);
buf BUF1 (N2109, N2106);
nor NOR3 (N2110, N2109, N489, N1217);
nor NOR2 (N2111, N2102, N1021);
not NOT1 (N2112, N2096);
xor XOR2 (N2113, N2090, N1204);
and AND2 (N2114, N2112, N1318);
and AND2 (N2115, N2107, N1078);
buf BUF1 (N2116, N2100);
and AND4 (N2117, N2110, N1439, N1853, N771);
not NOT1 (N2118, N2117);
nor NOR3 (N2119, N2087, N1826, N653);
or OR4 (N2120, N2108, N661, N896, N979);
not NOT1 (N2121, N2105);
and AND3 (N2122, N2119, N378, N943);
xor XOR2 (N2123, N2111, N263);
buf BUF1 (N2124, N2114);
xor XOR2 (N2125, N2120, N1099);
nand NAND2 (N2126, N2118, N514);
not NOT1 (N2127, N2103);
and AND3 (N2128, N2125, N2090, N1228);
buf BUF1 (N2129, N2122);
buf BUF1 (N2130, N2127);
not NOT1 (N2131, N2121);
or OR3 (N2132, N2130, N1374, N1360);
nor NOR4 (N2133, N2113, N416, N1406, N519);
nor NOR4 (N2134, N2133, N1084, N1779, N1621);
not NOT1 (N2135, N2132);
and AND3 (N2136, N2129, N928, N882);
and AND4 (N2137, N2136, N2039, N22, N1144);
not NOT1 (N2138, N2134);
buf BUF1 (N2139, N2128);
not NOT1 (N2140, N2126);
and AND3 (N2141, N2116, N1868, N2013);
not NOT1 (N2142, N2115);
nor NOR3 (N2143, N2131, N1071, N1380);
buf BUF1 (N2144, N2137);
xor XOR2 (N2145, N2143, N15);
nand NAND4 (N2146, N2138, N1465, N971, N1633);
buf BUF1 (N2147, N2140);
or OR3 (N2148, N2145, N835, N496);
nor NOR2 (N2149, N2135, N677);
xor XOR2 (N2150, N2142, N661);
or OR3 (N2151, N2147, N1279, N905);
buf BUF1 (N2152, N2124);
not NOT1 (N2153, N2123);
and AND4 (N2154, N2141, N487, N814, N1845);
or OR4 (N2155, N2149, N1561, N1513, N933);
and AND3 (N2156, N2150, N1484, N47);
buf BUF1 (N2157, N2151);
xor XOR2 (N2158, N2153, N1344);
nor NOR2 (N2159, N2157, N1068);
and AND2 (N2160, N2144, N583);
nor NOR4 (N2161, N2156, N1855, N498, N306);
nor NOR3 (N2162, N2161, N337, N1680);
nor NOR2 (N2163, N2160, N1095);
nand NAND2 (N2164, N2148, N735);
and AND2 (N2165, N2152, N2079);
and AND2 (N2166, N2158, N2110);
and AND2 (N2167, N2165, N844);
not NOT1 (N2168, N2163);
nor NOR3 (N2169, N2154, N1885, N959);
nor NOR3 (N2170, N2155, N1510, N1544);
nand NAND3 (N2171, N2168, N369, N1633);
or OR4 (N2172, N2139, N1015, N990, N1177);
nor NOR4 (N2173, N2167, N819, N1898, N1206);
or OR4 (N2174, N2170, N139, N726, N1521);
nand NAND4 (N2175, N2166, N1950, N614, N836);
or OR2 (N2176, N2159, N725);
xor XOR2 (N2177, N2175, N174);
xor XOR2 (N2178, N2176, N221);
nor NOR3 (N2179, N2178, N1207, N1766);
buf BUF1 (N2180, N2162);
nor NOR2 (N2181, N2171, N1189);
not NOT1 (N2182, N2164);
not NOT1 (N2183, N2182);
xor XOR2 (N2184, N2169, N603);
buf BUF1 (N2185, N2174);
nand NAND4 (N2186, N2172, N2089, N1787, N2097);
nor NOR3 (N2187, N2181, N1795, N648);
or OR3 (N2188, N2173, N1603, N868);
not NOT1 (N2189, N2184);
buf BUF1 (N2190, N2177);
or OR4 (N2191, N2180, N1000, N1965, N2141);
and AND4 (N2192, N2187, N2025, N1306, N1496);
or OR3 (N2193, N2190, N2146, N1288);
xor XOR2 (N2194, N1260, N1271);
and AND3 (N2195, N2183, N696, N107);
or OR4 (N2196, N2192, N961, N1623, N1084);
xor XOR2 (N2197, N2196, N1301);
xor XOR2 (N2198, N2197, N1105);
nor NOR2 (N2199, N2195, N73);
or OR2 (N2200, N2199, N1530);
or OR3 (N2201, N2198, N1119, N158);
nand NAND3 (N2202, N2185, N1003, N1633);
or OR2 (N2203, N2186, N1110);
nand NAND3 (N2204, N2191, N2034, N1895);
and AND2 (N2205, N2201, N1057);
xor XOR2 (N2206, N2189, N1619);
and AND3 (N2207, N2205, N655, N1394);
and AND3 (N2208, N2200, N717, N14);
not NOT1 (N2209, N2203);
nand NAND4 (N2210, N2204, N1411, N937, N1300);
and AND4 (N2211, N2208, N1257, N703, N963);
xor XOR2 (N2212, N2188, N1896);
not NOT1 (N2213, N2179);
not NOT1 (N2214, N2212);
and AND2 (N2215, N2213, N1018);
and AND2 (N2216, N2209, N1623);
and AND4 (N2217, N2216, N941, N1471, N472);
or OR2 (N2218, N2215, N1022);
buf BUF1 (N2219, N2207);
or OR3 (N2220, N2217, N1925, N1713);
nor NOR2 (N2221, N2218, N324);
buf BUF1 (N2222, N2193);
or OR2 (N2223, N2211, N1901);
nand NAND2 (N2224, N2206, N1257);
and AND2 (N2225, N2223, N1713);
buf BUF1 (N2226, N2222);
not NOT1 (N2227, N2219);
buf BUF1 (N2228, N2226);
xor XOR2 (N2229, N2194, N1273);
buf BUF1 (N2230, N2227);
xor XOR2 (N2231, N2214, N1270);
nand NAND2 (N2232, N2228, N1660);
or OR4 (N2233, N2202, N875, N1807, N2137);
nor NOR4 (N2234, N2220, N507, N1393, N833);
nor NOR4 (N2235, N2233, N1296, N301, N1290);
and AND3 (N2236, N2225, N1951, N9);
nor NOR4 (N2237, N2232, N1867, N1142, N1835);
not NOT1 (N2238, N2229);
nor NOR2 (N2239, N2224, N297);
nor NOR2 (N2240, N2230, N2106);
and AND2 (N2241, N2210, N1785);
nor NOR4 (N2242, N2234, N128, N470, N1511);
or OR2 (N2243, N2221, N1747);
or OR2 (N2244, N2239, N337);
and AND3 (N2245, N2238, N223, N1845);
nand NAND3 (N2246, N2243, N1438, N1793);
xor XOR2 (N2247, N2242, N1919);
nor NOR4 (N2248, N2235, N1211, N815, N2009);
and AND2 (N2249, N2246, N1758);
nor NOR2 (N2250, N2240, N15);
nor NOR2 (N2251, N2244, N1437);
and AND3 (N2252, N2247, N1689, N914);
nor NOR4 (N2253, N2248, N272, N140, N1005);
not NOT1 (N2254, N2231);
not NOT1 (N2255, N2251);
xor XOR2 (N2256, N2237, N108);
nand NAND3 (N2257, N2236, N363, N1020);
not NOT1 (N2258, N2254);
or OR4 (N2259, N2257, N1546, N824, N631);
or OR2 (N2260, N2250, N1301);
xor XOR2 (N2261, N2249, N1546);
xor XOR2 (N2262, N2261, N488);
buf BUF1 (N2263, N2259);
or OR3 (N2264, N2260, N661, N298);
nand NAND2 (N2265, N2264, N212);
buf BUF1 (N2266, N2255);
nand NAND2 (N2267, N2263, N2088);
or OR4 (N2268, N2245, N808, N313, N2025);
buf BUF1 (N2269, N2256);
not NOT1 (N2270, N2241);
xor XOR2 (N2271, N2266, N374);
or OR2 (N2272, N2268, N1974);
not NOT1 (N2273, N2270);
xor XOR2 (N2274, N2271, N2114);
buf BUF1 (N2275, N2267);
xor XOR2 (N2276, N2269, N1194);
xor XOR2 (N2277, N2272, N1913);
and AND2 (N2278, N2277, N1381);
buf BUF1 (N2279, N2258);
nor NOR2 (N2280, N2252, N1313);
or OR4 (N2281, N2273, N1315, N960, N1815);
and AND2 (N2282, N2275, N521);
xor XOR2 (N2283, N2278, N230);
and AND2 (N2284, N2280, N1098);
buf BUF1 (N2285, N2283);
buf BUF1 (N2286, N2262);
buf BUF1 (N2287, N2253);
buf BUF1 (N2288, N2282);
nor NOR2 (N2289, N2284, N1811);
nor NOR3 (N2290, N2279, N1782, N1148);
buf BUF1 (N2291, N2289);
or OR3 (N2292, N2276, N1041, N2100);
xor XOR2 (N2293, N2265, N832);
buf BUF1 (N2294, N2281);
buf BUF1 (N2295, N2274);
or OR2 (N2296, N2293, N2150);
or OR2 (N2297, N2286, N1281);
or OR3 (N2298, N2285, N123, N407);
nand NAND4 (N2299, N2295, N1865, N2074, N1626);
and AND2 (N2300, N2294, N535);
not NOT1 (N2301, N2287);
nand NAND4 (N2302, N2299, N2026, N2158, N330);
nor NOR2 (N2303, N2302, N1970);
and AND2 (N2304, N2288, N1634);
buf BUF1 (N2305, N2297);
nor NOR4 (N2306, N2298, N484, N493, N2068);
nor NOR4 (N2307, N2305, N603, N1706, N2101);
nor NOR3 (N2308, N2301, N844, N1168);
or OR4 (N2309, N2308, N2284, N216, N1727);
not NOT1 (N2310, N2291);
nand NAND2 (N2311, N2303, N1452);
and AND2 (N2312, N2292, N1159);
nand NAND3 (N2313, N2310, N2210, N16);
and AND3 (N2314, N2311, N1061, N569);
and AND4 (N2315, N2312, N130, N28, N1742);
or OR4 (N2316, N2315, N370, N990, N2122);
nand NAND2 (N2317, N2296, N1214);
and AND2 (N2318, N2316, N1032);
not NOT1 (N2319, N2317);
or OR4 (N2320, N2314, N2034, N1805, N1090);
nand NAND2 (N2321, N2320, N2280);
and AND2 (N2322, N2304, N128);
nand NAND3 (N2323, N2309, N1950, N1760);
not NOT1 (N2324, N2319);
nand NAND4 (N2325, N2321, N169, N1750, N975);
or OR4 (N2326, N2323, N1985, N811, N267);
or OR3 (N2327, N2322, N1996, N464);
xor XOR2 (N2328, N2324, N1667);
nand NAND4 (N2329, N2327, N2129, N1521, N2102);
and AND3 (N2330, N2290, N1139, N947);
buf BUF1 (N2331, N2307);
not NOT1 (N2332, N2328);
not NOT1 (N2333, N2300);
not NOT1 (N2334, N2330);
not NOT1 (N2335, N2318);
buf BUF1 (N2336, N2325);
nand NAND2 (N2337, N2336, N2232);
or OR3 (N2338, N2306, N2239, N1444);
not NOT1 (N2339, N2326);
or OR3 (N2340, N2338, N634, N247);
not NOT1 (N2341, N2340);
nor NOR2 (N2342, N2331, N1580);
xor XOR2 (N2343, N2337, N1620);
not NOT1 (N2344, N2334);
or OR2 (N2345, N2344, N187);
xor XOR2 (N2346, N2313, N2224);
or OR2 (N2347, N2339, N175);
buf BUF1 (N2348, N2345);
nand NAND4 (N2349, N2332, N781, N917, N176);
not NOT1 (N2350, N2343);
not NOT1 (N2351, N2329);
buf BUF1 (N2352, N2342);
nor NOR2 (N2353, N2347, N1934);
buf BUF1 (N2354, N2351);
and AND3 (N2355, N2348, N752, N1537);
nor NOR4 (N2356, N2354, N1395, N1030, N432);
nand NAND4 (N2357, N2341, N1408, N1308, N1232);
buf BUF1 (N2358, N2352);
not NOT1 (N2359, N2358);
and AND2 (N2360, N2346, N391);
xor XOR2 (N2361, N2333, N618);
nand NAND2 (N2362, N2335, N341);
nand NAND3 (N2363, N2357, N1383, N720);
nand NAND2 (N2364, N2363, N478);
xor XOR2 (N2365, N2360, N399);
or OR3 (N2366, N2356, N1455, N2151);
nor NOR4 (N2367, N2355, N1449, N2168, N84);
and AND3 (N2368, N2364, N1294, N986);
nand NAND4 (N2369, N2349, N1463, N584, N1524);
and AND3 (N2370, N2353, N1801, N1723);
nor NOR3 (N2371, N2366, N929, N1647);
buf BUF1 (N2372, N2361);
buf BUF1 (N2373, N2350);
not NOT1 (N2374, N2359);
and AND4 (N2375, N2369, N923, N1452, N369);
and AND3 (N2376, N2365, N667, N1701);
nor NOR3 (N2377, N2373, N1016, N763);
not NOT1 (N2378, N2367);
nor NOR3 (N2379, N2372, N2050, N1939);
nand NAND4 (N2380, N2376, N567, N1453, N385);
nor NOR2 (N2381, N2371, N2103);
not NOT1 (N2382, N2380);
buf BUF1 (N2383, N2379);
nor NOR2 (N2384, N2362, N675);
buf BUF1 (N2385, N2382);
nor NOR4 (N2386, N2378, N885, N1967, N2018);
nand NAND2 (N2387, N2375, N2341);
or OR4 (N2388, N2368, N351, N1254, N258);
and AND3 (N2389, N2387, N2003, N444);
nor NOR4 (N2390, N2374, N4, N1131, N90);
nand NAND3 (N2391, N2385, N1232, N1535);
nor NOR3 (N2392, N2386, N1813, N1960);
nand NAND3 (N2393, N2389, N1208, N2132);
nand NAND4 (N2394, N2370, N1989, N1597, N1115);
not NOT1 (N2395, N2392);
or OR4 (N2396, N2388, N1799, N262, N1706);
buf BUF1 (N2397, N2393);
not NOT1 (N2398, N2390);
nand NAND4 (N2399, N2395, N243, N744, N1627);
xor XOR2 (N2400, N2394, N184);
nand NAND3 (N2401, N2377, N658, N2045);
nor NOR4 (N2402, N2397, N115, N676, N1618);
nor NOR2 (N2403, N2381, N357);
not NOT1 (N2404, N2391);
buf BUF1 (N2405, N2400);
nor NOR2 (N2406, N2404, N1481);
buf BUF1 (N2407, N2401);
or OR3 (N2408, N2396, N1191, N986);
and AND3 (N2409, N2403, N1859, N1794);
nand NAND2 (N2410, N2383, N217);
buf BUF1 (N2411, N2407);
nand NAND4 (N2412, N2411, N107, N391, N2087);
not NOT1 (N2413, N2405);
and AND3 (N2414, N2399, N189, N1148);
nand NAND2 (N2415, N2398, N1894);
and AND4 (N2416, N2402, N253, N703, N2318);
xor XOR2 (N2417, N2416, N643);
and AND3 (N2418, N2417, N352, N1160);
nor NOR4 (N2419, N2384, N2222, N487, N611);
nand NAND4 (N2420, N2408, N1302, N2298, N2136);
nand NAND4 (N2421, N2409, N2391, N945, N2269);
xor XOR2 (N2422, N2406, N850);
or OR3 (N2423, N2421, N996, N618);
buf BUF1 (N2424, N2413);
or OR3 (N2425, N2422, N18, N890);
nor NOR4 (N2426, N2412, N1679, N557, N2088);
nor NOR2 (N2427, N2425, N333);
buf BUF1 (N2428, N2418);
xor XOR2 (N2429, N2419, N1729);
and AND2 (N2430, N2414, N2040);
nand NAND3 (N2431, N2428, N2390, N877);
nand NAND4 (N2432, N2415, N183, N315, N2206);
nand NAND2 (N2433, N2423, N7);
nor NOR3 (N2434, N2432, N275, N1165);
or OR2 (N2435, N2434, N2092);
buf BUF1 (N2436, N2427);
or OR4 (N2437, N2426, N746, N162, N2332);
buf BUF1 (N2438, N2410);
xor XOR2 (N2439, N2438, N1820);
not NOT1 (N2440, N2435);
xor XOR2 (N2441, N2436, N2434);
buf BUF1 (N2442, N2424);
not NOT1 (N2443, N2440);
buf BUF1 (N2444, N2443);
xor XOR2 (N2445, N2420, N148);
xor XOR2 (N2446, N2437, N2196);
nand NAND3 (N2447, N2444, N1601, N2075);
not NOT1 (N2448, N2433);
xor XOR2 (N2449, N2446, N753);
not NOT1 (N2450, N2442);
xor XOR2 (N2451, N2430, N1953);
and AND4 (N2452, N2441, N360, N1359, N1237);
xor XOR2 (N2453, N2450, N2389);
buf BUF1 (N2454, N2453);
and AND4 (N2455, N2445, N1130, N683, N825);
or OR3 (N2456, N2448, N2249, N2295);
or OR2 (N2457, N2455, N1539);
not NOT1 (N2458, N2457);
or OR4 (N2459, N2447, N594, N440, N1270);
xor XOR2 (N2460, N2429, N2031);
or OR4 (N2461, N2454, N581, N2301, N1641);
not NOT1 (N2462, N2452);
or OR4 (N2463, N2431, N51, N2377, N1782);
nand NAND3 (N2464, N2456, N500, N424);
and AND2 (N2465, N2460, N1316);
nand NAND3 (N2466, N2461, N2006, N2245);
nand NAND2 (N2467, N2462, N1276);
buf BUF1 (N2468, N2467);
not NOT1 (N2469, N2465);
and AND2 (N2470, N2449, N2387);
nor NOR2 (N2471, N2458, N1920);
not NOT1 (N2472, N2469);
and AND2 (N2473, N2471, N1816);
buf BUF1 (N2474, N2466);
xor XOR2 (N2475, N2464, N40);
or OR3 (N2476, N2463, N684, N274);
nand NAND4 (N2477, N2459, N2224, N1552, N1761);
or OR4 (N2478, N2468, N1376, N635, N1624);
or OR2 (N2479, N2478, N1802);
or OR4 (N2480, N2451, N1260, N1695, N1881);
nand NAND4 (N2481, N2477, N1223, N978, N1813);
xor XOR2 (N2482, N2439, N183);
and AND4 (N2483, N2474, N1209, N531, N1019);
buf BUF1 (N2484, N2472);
nor NOR4 (N2485, N2481, N2095, N2426, N1476);
xor XOR2 (N2486, N2476, N2135);
xor XOR2 (N2487, N2480, N974);
not NOT1 (N2488, N2483);
and AND3 (N2489, N2475, N1031, N48);
not NOT1 (N2490, N2484);
and AND3 (N2491, N2485, N1822, N1191);
and AND4 (N2492, N2473, N1137, N1157, N1001);
nand NAND2 (N2493, N2470, N1356);
buf BUF1 (N2494, N2486);
or OR2 (N2495, N2493, N1755);
xor XOR2 (N2496, N2495, N1991);
xor XOR2 (N2497, N2488, N1906);
and AND4 (N2498, N2494, N1338, N1986, N153);
or OR2 (N2499, N2496, N717);
or OR3 (N2500, N2498, N1137, N189);
not NOT1 (N2501, N2489);
xor XOR2 (N2502, N2492, N1724);
not NOT1 (N2503, N2479);
buf BUF1 (N2504, N2500);
nand NAND2 (N2505, N2490, N1586);
and AND2 (N2506, N2497, N20);
or OR4 (N2507, N2506, N896, N2095, N666);
and AND2 (N2508, N2482, N127);
and AND4 (N2509, N2487, N509, N2384, N825);
nor NOR3 (N2510, N2508, N1884, N935);
xor XOR2 (N2511, N2510, N1217);
and AND3 (N2512, N2491, N13, N651);
xor XOR2 (N2513, N2499, N1369);
or OR2 (N2514, N2509, N1813);
buf BUF1 (N2515, N2504);
buf BUF1 (N2516, N2515);
not NOT1 (N2517, N2511);
or OR2 (N2518, N2501, N1538);
nand NAND4 (N2519, N2502, N522, N438, N2476);
or OR3 (N2520, N2517, N2345, N1271);
buf BUF1 (N2521, N2512);
nand NAND4 (N2522, N2516, N1107, N1478, N1007);
nor NOR4 (N2523, N2505, N58, N213, N551);
buf BUF1 (N2524, N2514);
buf BUF1 (N2525, N2519);
buf BUF1 (N2526, N2523);
or OR4 (N2527, N2526, N195, N1341, N1705);
nand NAND4 (N2528, N2507, N1883, N540, N601);
buf BUF1 (N2529, N2503);
buf BUF1 (N2530, N2527);
buf BUF1 (N2531, N2521);
or OR4 (N2532, N2513, N323, N2143, N2516);
xor XOR2 (N2533, N2524, N385);
nand NAND4 (N2534, N2518, N408, N1807, N753);
nand NAND3 (N2535, N2525, N1682, N915);
buf BUF1 (N2536, N2534);
not NOT1 (N2537, N2533);
or OR2 (N2538, N2532, N2369);
and AND3 (N2539, N2530, N696, N2439);
xor XOR2 (N2540, N2535, N1551);
nand NAND3 (N2541, N2540, N237, N56);
nor NOR2 (N2542, N2528, N526);
not NOT1 (N2543, N2538);
nand NAND4 (N2544, N2536, N2310, N925, N889);
nand NAND4 (N2545, N2529, N584, N388, N1254);
xor XOR2 (N2546, N2531, N1653);
not NOT1 (N2547, N2545);
and AND3 (N2548, N2522, N75, N1532);
nand NAND3 (N2549, N2541, N1759, N747);
or OR4 (N2550, N2543, N1813, N2304, N1627);
nand NAND4 (N2551, N2546, N1788, N1273, N1351);
nor NOR2 (N2552, N2520, N897);
not NOT1 (N2553, N2544);
nand NAND3 (N2554, N2551, N2136, N2447);
and AND3 (N2555, N2547, N1241, N1303);
or OR4 (N2556, N2553, N1922, N1512, N20);
nand NAND4 (N2557, N2552, N2071, N1206, N406);
and AND4 (N2558, N2555, N2016, N242, N1937);
buf BUF1 (N2559, N2539);
nand NAND3 (N2560, N2548, N714, N2169);
xor XOR2 (N2561, N2557, N516);
nor NOR2 (N2562, N2554, N306);
or OR4 (N2563, N2542, N2177, N1644, N1244);
buf BUF1 (N2564, N2560);
xor XOR2 (N2565, N2537, N639);
not NOT1 (N2566, N2558);
not NOT1 (N2567, N2561);
and AND3 (N2568, N2556, N2358, N1235);
and AND2 (N2569, N2559, N2239);
or OR3 (N2570, N2569, N335, N458);
not NOT1 (N2571, N2570);
or OR3 (N2572, N2568, N1866, N2483);
nand NAND3 (N2573, N2565, N966, N2089);
not NOT1 (N2574, N2567);
not NOT1 (N2575, N2562);
xor XOR2 (N2576, N2571, N145);
xor XOR2 (N2577, N2563, N1748);
buf BUF1 (N2578, N2564);
xor XOR2 (N2579, N2573, N1005);
nor NOR2 (N2580, N2566, N861);
nand NAND3 (N2581, N2550, N1605, N1273);
xor XOR2 (N2582, N2574, N1541);
xor XOR2 (N2583, N2572, N2175);
nand NAND4 (N2584, N2576, N1211, N1749, N2344);
xor XOR2 (N2585, N2584, N874);
xor XOR2 (N2586, N2579, N2350);
nand NAND3 (N2587, N2577, N762, N235);
not NOT1 (N2588, N2582);
or OR3 (N2589, N2587, N1175, N1860);
xor XOR2 (N2590, N2581, N851);
and AND2 (N2591, N2575, N2176);
and AND2 (N2592, N2580, N1152);
and AND4 (N2593, N2590, N754, N897, N478);
and AND3 (N2594, N2592, N109, N2155);
buf BUF1 (N2595, N2588);
nor NOR3 (N2596, N2583, N1883, N2051);
and AND4 (N2597, N2593, N277, N2021, N1930);
nor NOR4 (N2598, N2549, N1378, N72, N70);
not NOT1 (N2599, N2585);
nor NOR3 (N2600, N2597, N681, N1638);
or OR4 (N2601, N2599, N2338, N2004, N527);
and AND4 (N2602, N2591, N622, N395, N1426);
xor XOR2 (N2603, N2601, N1502);
nor NOR3 (N2604, N2596, N1682, N1750);
nor NOR3 (N2605, N2594, N2479, N565);
nor NOR2 (N2606, N2600, N1955);
not NOT1 (N2607, N2606);
and AND4 (N2608, N2604, N190, N1244, N382);
not NOT1 (N2609, N2608);
nand NAND4 (N2610, N2603, N1770, N1656, N1331);
or OR3 (N2611, N2610, N1706, N1876);
or OR4 (N2612, N2595, N1845, N2098, N1090);
xor XOR2 (N2613, N2612, N2348);
xor XOR2 (N2614, N2607, N1832);
and AND3 (N2615, N2611, N1405, N2555);
nor NOR2 (N2616, N2602, N1479);
or OR3 (N2617, N2589, N2172, N304);
not NOT1 (N2618, N2616);
nor NOR3 (N2619, N2618, N2574, N1754);
not NOT1 (N2620, N2614);
buf BUF1 (N2621, N2613);
and AND3 (N2622, N2615, N856, N461);
buf BUF1 (N2623, N2620);
nand NAND3 (N2624, N2623, N2096, N1946);
nand NAND3 (N2625, N2619, N2264, N1931);
buf BUF1 (N2626, N2621);
or OR3 (N2627, N2586, N323, N2432);
nor NOR2 (N2628, N2605, N2258);
not NOT1 (N2629, N2624);
not NOT1 (N2630, N2578);
nor NOR3 (N2631, N2628, N2317, N1486);
not NOT1 (N2632, N2622);
and AND3 (N2633, N2632, N2590, N1824);
buf BUF1 (N2634, N2631);
not NOT1 (N2635, N2634);
xor XOR2 (N2636, N2617, N43);
nand NAND3 (N2637, N2630, N1900, N284);
xor XOR2 (N2638, N2609, N361);
buf BUF1 (N2639, N2633);
buf BUF1 (N2640, N2637);
xor XOR2 (N2641, N2635, N680);
nand NAND4 (N2642, N2626, N1133, N1456, N2631);
nand NAND2 (N2643, N2640, N1320);
nand NAND4 (N2644, N2598, N2216, N2331, N476);
nor NOR3 (N2645, N2644, N1951, N2110);
not NOT1 (N2646, N2629);
xor XOR2 (N2647, N2642, N1785);
buf BUF1 (N2648, N2647);
buf BUF1 (N2649, N2638);
buf BUF1 (N2650, N2648);
not NOT1 (N2651, N2627);
buf BUF1 (N2652, N2625);
not NOT1 (N2653, N2645);
and AND4 (N2654, N2652, N610, N661, N1787);
not NOT1 (N2655, N2636);
not NOT1 (N2656, N2650);
buf BUF1 (N2657, N2649);
or OR3 (N2658, N2643, N789, N691);
xor XOR2 (N2659, N2656, N145);
and AND4 (N2660, N2641, N2073, N1696, N2188);
nor NOR3 (N2661, N2653, N320, N508);
not NOT1 (N2662, N2660);
not NOT1 (N2663, N2646);
and AND2 (N2664, N2657, N1833);
not NOT1 (N2665, N2663);
or OR3 (N2666, N2639, N2402, N1858);
not NOT1 (N2667, N2651);
xor XOR2 (N2668, N2654, N1874);
buf BUF1 (N2669, N2655);
nor NOR4 (N2670, N2664, N1725, N2102, N10);
xor XOR2 (N2671, N2669, N361);
or OR3 (N2672, N2671, N340, N1237);
and AND3 (N2673, N2672, N487, N2270);
and AND2 (N2674, N2659, N2524);
xor XOR2 (N2675, N2661, N698);
not NOT1 (N2676, N2670);
nand NAND3 (N2677, N2676, N1435, N2111);
nor NOR3 (N2678, N2673, N1738, N1241);
nor NOR4 (N2679, N2674, N2350, N1979, N1615);
not NOT1 (N2680, N2677);
nor NOR4 (N2681, N2668, N1960, N475, N1457);
or OR2 (N2682, N2678, N1750);
nand NAND4 (N2683, N2665, N1413, N974, N2586);
nand NAND3 (N2684, N2666, N1819, N2264);
nor NOR3 (N2685, N2658, N961, N2450);
not NOT1 (N2686, N2679);
buf BUF1 (N2687, N2681);
not NOT1 (N2688, N2680);
xor XOR2 (N2689, N2667, N1469);
buf BUF1 (N2690, N2683);
and AND4 (N2691, N2689, N1250, N981, N704);
xor XOR2 (N2692, N2685, N1755);
or OR2 (N2693, N2675, N1866);
nand NAND3 (N2694, N2688, N650, N223);
nand NAND2 (N2695, N2687, N378);
nor NOR4 (N2696, N2662, N1140, N928, N20);
or OR3 (N2697, N2694, N2420, N1634);
xor XOR2 (N2698, N2690, N808);
nor NOR4 (N2699, N2695, N921, N1266, N2298);
not NOT1 (N2700, N2686);
buf BUF1 (N2701, N2692);
xor XOR2 (N2702, N2701, N2695);
or OR4 (N2703, N2682, N1401, N2172, N344);
buf BUF1 (N2704, N2693);
buf BUF1 (N2705, N2684);
xor XOR2 (N2706, N2700, N1931);
not NOT1 (N2707, N2691);
xor XOR2 (N2708, N2696, N223);
not NOT1 (N2709, N2703);
buf BUF1 (N2710, N2706);
xor XOR2 (N2711, N2699, N1209);
nor NOR3 (N2712, N2708, N2111, N2019);
buf BUF1 (N2713, N2712);
buf BUF1 (N2714, N2707);
or OR3 (N2715, N2709, N2490, N1775);
nand NAND4 (N2716, N2704, N419, N1280, N2235);
not NOT1 (N2717, N2711);
nor NOR4 (N2718, N2715, N2040, N1884, N2684);
and AND2 (N2719, N2716, N1872);
xor XOR2 (N2720, N2698, N2270);
buf BUF1 (N2721, N2720);
buf BUF1 (N2722, N2705);
xor XOR2 (N2723, N2710, N732);
nor NOR4 (N2724, N2714, N2271, N1956, N2695);
xor XOR2 (N2725, N2718, N2567);
not NOT1 (N2726, N2719);
nor NOR4 (N2727, N2713, N2300, N936, N551);
nand NAND2 (N2728, N2702, N1183);
nand NAND3 (N2729, N2724, N1490, N510);
not NOT1 (N2730, N2717);
or OR3 (N2731, N2730, N2021, N91);
nand NAND3 (N2732, N2697, N648, N237);
or OR4 (N2733, N2721, N1570, N1455, N481);
and AND4 (N2734, N2733, N1330, N1734, N460);
nor NOR2 (N2735, N2728, N668);
not NOT1 (N2736, N2726);
nand NAND2 (N2737, N2729, N1722);
nor NOR4 (N2738, N2725, N2396, N2011, N57);
nand NAND2 (N2739, N2735, N1275);
nor NOR4 (N2740, N2731, N262, N1084, N2026);
buf BUF1 (N2741, N2736);
xor XOR2 (N2742, N2727, N2405);
buf BUF1 (N2743, N2737);
nor NOR3 (N2744, N2722, N1550, N1058);
not NOT1 (N2745, N2738);
buf BUF1 (N2746, N2744);
nor NOR3 (N2747, N2743, N2738, N655);
or OR2 (N2748, N2747, N476);
xor XOR2 (N2749, N2732, N748);
nand NAND2 (N2750, N2749, N1340);
buf BUF1 (N2751, N2748);
xor XOR2 (N2752, N2745, N2119);
not NOT1 (N2753, N2750);
nand NAND4 (N2754, N2751, N2169, N2664, N2393);
or OR4 (N2755, N2742, N1767, N2497, N90);
nor NOR2 (N2756, N2734, N104);
xor XOR2 (N2757, N2755, N200);
nand NAND4 (N2758, N2757, N1658, N1937, N1296);
xor XOR2 (N2759, N2754, N415);
nor NOR4 (N2760, N2741, N2615, N2496, N371);
or OR3 (N2761, N2752, N384, N2205);
nor NOR4 (N2762, N2740, N930, N916, N2511);
not NOT1 (N2763, N2758);
xor XOR2 (N2764, N2756, N1494);
nor NOR4 (N2765, N2763, N361, N783, N1183);
buf BUF1 (N2766, N2753);
or OR3 (N2767, N2760, N2646, N2693);
or OR2 (N2768, N2764, N958);
nor NOR4 (N2769, N2739, N1196, N1782, N712);
not NOT1 (N2770, N2746);
xor XOR2 (N2771, N2765, N2732);
nand NAND3 (N2772, N2768, N758, N720);
and AND2 (N2773, N2762, N1174);
buf BUF1 (N2774, N2772);
not NOT1 (N2775, N2769);
xor XOR2 (N2776, N2774, N1355);
and AND2 (N2777, N2723, N1383);
or OR3 (N2778, N2761, N1508, N1696);
nor NOR3 (N2779, N2770, N1801, N2681);
not NOT1 (N2780, N2779);
buf BUF1 (N2781, N2767);
buf BUF1 (N2782, N2771);
not NOT1 (N2783, N2782);
or OR3 (N2784, N2780, N2570, N747);
or OR3 (N2785, N2773, N432, N1565);
not NOT1 (N2786, N2759);
and AND3 (N2787, N2783, N1582, N2686);
nor NOR4 (N2788, N2781, N1482, N488, N1097);
xor XOR2 (N2789, N2787, N2770);
or OR3 (N2790, N2786, N609, N1986);
nor NOR4 (N2791, N2778, N460, N70, N2088);
buf BUF1 (N2792, N2775);
nand NAND3 (N2793, N2784, N1523, N472);
and AND2 (N2794, N2793, N1512);
or OR4 (N2795, N2785, N28, N2554, N570);
and AND4 (N2796, N2792, N2463, N1318, N1122);
buf BUF1 (N2797, N2795);
nor NOR3 (N2798, N2777, N1594, N2425);
buf BUF1 (N2799, N2791);
not NOT1 (N2800, N2789);
xor XOR2 (N2801, N2776, N777);
xor XOR2 (N2802, N2801, N1217);
buf BUF1 (N2803, N2790);
and AND4 (N2804, N2800, N1974, N2283, N1063);
nand NAND3 (N2805, N2796, N1351, N891);
or OR2 (N2806, N2788, N2675);
nand NAND3 (N2807, N2803, N1575, N1701);
not NOT1 (N2808, N2797);
nor NOR2 (N2809, N2808, N1854);
xor XOR2 (N2810, N2809, N2755);
not NOT1 (N2811, N2766);
nand NAND3 (N2812, N2810, N794, N185);
or OR4 (N2813, N2799, N297, N1406, N1722);
not NOT1 (N2814, N2805);
not NOT1 (N2815, N2804);
or OR2 (N2816, N2815, N2364);
xor XOR2 (N2817, N2812, N1014);
nand NAND2 (N2818, N2814, N2435);
or OR3 (N2819, N2816, N1880, N2344);
xor XOR2 (N2820, N2794, N736);
nor NOR3 (N2821, N2818, N652, N1472);
or OR3 (N2822, N2819, N740, N883);
and AND3 (N2823, N2806, N497, N1381);
buf BUF1 (N2824, N2820);
or OR2 (N2825, N2807, N71);
nand NAND3 (N2826, N2825, N84, N1423);
xor XOR2 (N2827, N2802, N363);
nor NOR4 (N2828, N2826, N696, N2422, N969);
not NOT1 (N2829, N2813);
nand NAND4 (N2830, N2823, N2162, N858, N2398);
xor XOR2 (N2831, N2817, N986);
nand NAND2 (N2832, N2824, N2621);
buf BUF1 (N2833, N2798);
or OR2 (N2834, N2829, N2762);
and AND4 (N2835, N2834, N2400, N2019, N413);
not NOT1 (N2836, N2811);
not NOT1 (N2837, N2836);
buf BUF1 (N2838, N2837);
or OR4 (N2839, N2832, N461, N2668, N2498);
nand NAND4 (N2840, N2833, N1524, N707, N1721);
or OR3 (N2841, N2839, N614, N1889);
not NOT1 (N2842, N2827);
or OR4 (N2843, N2841, N1880, N181, N907);
nor NOR4 (N2844, N2838, N2769, N1087, N225);
not NOT1 (N2845, N2830);
xor XOR2 (N2846, N2831, N881);
or OR2 (N2847, N2843, N2735);
or OR3 (N2848, N2846, N254, N675);
buf BUF1 (N2849, N2835);
and AND2 (N2850, N2848, N1846);
or OR4 (N2851, N2821, N641, N1351, N1947);
and AND4 (N2852, N2849, N2195, N2294, N2027);
xor XOR2 (N2853, N2852, N440);
xor XOR2 (N2854, N2853, N1093);
buf BUF1 (N2855, N2851);
nor NOR2 (N2856, N2850, N462);
nor NOR2 (N2857, N2854, N2530);
and AND2 (N2858, N2855, N1940);
or OR4 (N2859, N2847, N423, N214, N1783);
nand NAND2 (N2860, N2858, N2769);
not NOT1 (N2861, N2860);
nand NAND3 (N2862, N2842, N2506, N1948);
buf BUF1 (N2863, N2861);
buf BUF1 (N2864, N2859);
nand NAND2 (N2865, N2844, N2790);
buf BUF1 (N2866, N2863);
nand NAND4 (N2867, N2840, N664, N2626, N1813);
nor NOR2 (N2868, N2866, N1265);
not NOT1 (N2869, N2822);
or OR3 (N2870, N2856, N280, N1350);
and AND3 (N2871, N2865, N1945, N1536);
buf BUF1 (N2872, N2864);
or OR3 (N2873, N2867, N1617, N1447);
and AND2 (N2874, N2872, N875);
nand NAND4 (N2875, N2845, N635, N777, N502);
not NOT1 (N2876, N2869);
and AND2 (N2877, N2871, N2462);
xor XOR2 (N2878, N2868, N2231);
buf BUF1 (N2879, N2828);
and AND2 (N2880, N2874, N1097);
buf BUF1 (N2881, N2873);
and AND4 (N2882, N2876, N90, N1808, N2144);
buf BUF1 (N2883, N2877);
nor NOR4 (N2884, N2875, N1878, N903, N400);
or OR4 (N2885, N2870, N2824, N1164, N2757);
xor XOR2 (N2886, N2882, N2245);
buf BUF1 (N2887, N2857);
not NOT1 (N2888, N2887);
nand NAND4 (N2889, N2881, N1015, N2536, N1160);
nor NOR2 (N2890, N2886, N2170);
nor NOR3 (N2891, N2884, N2413, N2103);
and AND4 (N2892, N2889, N1439, N930, N1947);
buf BUF1 (N2893, N2888);
not NOT1 (N2894, N2890);
not NOT1 (N2895, N2880);
nor NOR4 (N2896, N2862, N2892, N461, N2798);
nor NOR4 (N2897, N1769, N1314, N1172, N133);
or OR2 (N2898, N2891, N446);
nand NAND2 (N2899, N2898, N2267);
or OR4 (N2900, N2895, N318, N998, N902);
nand NAND2 (N2901, N2896, N2094);
xor XOR2 (N2902, N2900, N153);
xor XOR2 (N2903, N2893, N702);
nand NAND4 (N2904, N2878, N2702, N2214, N1037);
nor NOR4 (N2905, N2904, N104, N402, N2448);
buf BUF1 (N2906, N2885);
nand NAND3 (N2907, N2903, N840, N988);
nor NOR4 (N2908, N2905, N2151, N2905, N1424);
not NOT1 (N2909, N2897);
nor NOR3 (N2910, N2906, N103, N2607);
not NOT1 (N2911, N2907);
xor XOR2 (N2912, N2899, N242);
buf BUF1 (N2913, N2883);
not NOT1 (N2914, N2894);
nor NOR2 (N2915, N2901, N908);
and AND4 (N2916, N2914, N2529, N2464, N2558);
buf BUF1 (N2917, N2909);
or OR3 (N2918, N2912, N1445, N161);
and AND2 (N2919, N2916, N687);
nor NOR2 (N2920, N2919, N1691);
or OR2 (N2921, N2913, N1509);
nor NOR4 (N2922, N2921, N1743, N2267, N848);
buf BUF1 (N2923, N2915);
nor NOR2 (N2924, N2879, N178);
nand NAND4 (N2925, N2911, N1306, N462, N1338);
buf BUF1 (N2926, N2902);
or OR2 (N2927, N2922, N1022);
or OR2 (N2928, N2926, N2747);
nand NAND2 (N2929, N2918, N1084);
nor NOR4 (N2930, N2908, N2775, N2925, N1705);
nand NAND2 (N2931, N581, N1488);
and AND3 (N2932, N2931, N535, N2683);
nor NOR4 (N2933, N2910, N1896, N974, N2209);
and AND3 (N2934, N2933, N1733, N2410);
not NOT1 (N2935, N2920);
not NOT1 (N2936, N2932);
or OR4 (N2937, N2936, N2577, N1306, N1040);
xor XOR2 (N2938, N2934, N2523);
and AND4 (N2939, N2917, N2173, N46, N2120);
buf BUF1 (N2940, N2923);
xor XOR2 (N2941, N2938, N2720);
nand NAND3 (N2942, N2929, N2708, N1113);
buf BUF1 (N2943, N2937);
or OR2 (N2944, N2924, N746);
xor XOR2 (N2945, N2939, N474);
xor XOR2 (N2946, N2940, N2277);
and AND3 (N2947, N2928, N1298, N2366);
nand NAND4 (N2948, N2944, N464, N613, N2202);
and AND2 (N2949, N2935, N2347);
xor XOR2 (N2950, N2927, N737);
not NOT1 (N2951, N2942);
or OR4 (N2952, N2930, N2815, N887, N2302);
xor XOR2 (N2953, N2945, N482);
not NOT1 (N2954, N2946);
buf BUF1 (N2955, N2948);
xor XOR2 (N2956, N2954, N258);
buf BUF1 (N2957, N2953);
and AND4 (N2958, N2957, N151, N2390, N1204);
xor XOR2 (N2959, N2951, N1816);
nand NAND4 (N2960, N2956, N1064, N1253, N1869);
nor NOR3 (N2961, N2959, N2157, N399);
buf BUF1 (N2962, N2961);
not NOT1 (N2963, N2949);
and AND4 (N2964, N2955, N2136, N1770, N2713);
nand NAND3 (N2965, N2964, N389, N1033);
or OR4 (N2966, N2958, N2571, N1874, N2320);
not NOT1 (N2967, N2947);
xor XOR2 (N2968, N2963, N2703);
not NOT1 (N2969, N2962);
buf BUF1 (N2970, N2941);
not NOT1 (N2971, N2965);
not NOT1 (N2972, N2966);
not NOT1 (N2973, N2970);
or OR3 (N2974, N2969, N1128, N2039);
or OR2 (N2975, N2967, N2654);
or OR2 (N2976, N2960, N1720);
buf BUF1 (N2977, N2950);
buf BUF1 (N2978, N2975);
and AND4 (N2979, N2952, N1339, N556, N1815);
nand NAND3 (N2980, N2978, N2822, N2564);
nand NAND4 (N2981, N2971, N1841, N1438, N2598);
or OR2 (N2982, N2981, N1152);
xor XOR2 (N2983, N2974, N2287);
nor NOR2 (N2984, N2979, N1890);
buf BUF1 (N2985, N2980);
buf BUF1 (N2986, N2976);
or OR4 (N2987, N2972, N356, N720, N726);
nor NOR2 (N2988, N2986, N2378);
or OR2 (N2989, N2968, N386);
nand NAND3 (N2990, N2983, N996, N1638);
and AND3 (N2991, N2990, N2014, N936);
and AND2 (N2992, N2985, N2363);
not NOT1 (N2993, N2943);
or OR3 (N2994, N2982, N2886, N2477);
or OR2 (N2995, N2989, N1016);
nor NOR4 (N2996, N2973, N2096, N1766, N1328);
xor XOR2 (N2997, N2988, N967);
or OR3 (N2998, N2977, N306, N2109);
buf BUF1 (N2999, N2998);
not NOT1 (N3000, N2996);
nand NAND3 (N3001, N2992, N2120, N697);
or OR3 (N3002, N3000, N416, N2272);
nor NOR4 (N3003, N2991, N1165, N1947, N2034);
buf BUF1 (N3004, N2995);
or OR3 (N3005, N2984, N3003, N2202);
nand NAND3 (N3006, N2162, N1797, N2950);
or OR2 (N3007, N3001, N957);
or OR4 (N3008, N3006, N1599, N346, N825);
buf BUF1 (N3009, N3007);
not NOT1 (N3010, N2999);
nand NAND4 (N3011, N2987, N972, N2669, N2172);
or OR3 (N3012, N3008, N50, N281);
or OR3 (N3013, N2994, N582, N2912);
and AND2 (N3014, N3002, N600);
buf BUF1 (N3015, N3010);
not NOT1 (N3016, N2993);
nand NAND2 (N3017, N3014, N1161);
xor XOR2 (N3018, N3004, N299);
xor XOR2 (N3019, N3005, N233);
and AND3 (N3020, N3015, N595, N2556);
nor NOR3 (N3021, N3012, N2372, N1712);
buf BUF1 (N3022, N3021);
nand NAND2 (N3023, N3013, N622);
or OR4 (N3024, N2997, N2407, N1992, N2794);
xor XOR2 (N3025, N3016, N403);
nor NOR3 (N3026, N3009, N492, N2091);
nand NAND2 (N3027, N3019, N1921);
nor NOR2 (N3028, N3024, N2106);
not NOT1 (N3029, N3022);
buf BUF1 (N3030, N3018);
not NOT1 (N3031, N3026);
nand NAND4 (N3032, N3017, N2429, N1502, N827);
xor XOR2 (N3033, N3011, N227);
and AND4 (N3034, N3031, N1114, N436, N2679);
nand NAND2 (N3035, N3032, N3029);
xor XOR2 (N3036, N745, N1756);
not NOT1 (N3037, N3027);
nand NAND2 (N3038, N3035, N956);
nand NAND4 (N3039, N3037, N1096, N2696, N2369);
xor XOR2 (N3040, N3030, N1229);
buf BUF1 (N3041, N3040);
nand NAND4 (N3042, N3028, N135, N1046, N679);
not NOT1 (N3043, N3038);
not NOT1 (N3044, N3034);
xor XOR2 (N3045, N3042, N2361);
nand NAND4 (N3046, N3041, N2158, N1022, N2671);
xor XOR2 (N3047, N3046, N2424);
not NOT1 (N3048, N3023);
buf BUF1 (N3049, N3044);
nand NAND4 (N3050, N3047, N2472, N2119, N777);
not NOT1 (N3051, N3033);
buf BUF1 (N3052, N3036);
or OR4 (N3053, N3039, N699, N1807, N1685);
not NOT1 (N3054, N3053);
nor NOR4 (N3055, N3045, N1878, N1477, N3023);
xor XOR2 (N3056, N3054, N2727);
or OR2 (N3057, N3048, N203);
xor XOR2 (N3058, N3051, N1915);
buf BUF1 (N3059, N3020);
nor NOR3 (N3060, N3059, N1331, N117);
buf BUF1 (N3061, N3058);
nand NAND3 (N3062, N3050, N2078, N1958);
nor NOR3 (N3063, N3043, N2462, N740);
nand NAND3 (N3064, N3063, N2614, N2095);
nand NAND3 (N3065, N3056, N1182, N585);
not NOT1 (N3066, N3057);
and AND2 (N3067, N3025, N1607);
nand NAND3 (N3068, N3055, N93, N1098);
nor NOR4 (N3069, N3067, N793, N1524, N2528);
nand NAND4 (N3070, N3065, N718, N1570, N91);
nand NAND4 (N3071, N3061, N2279, N1910, N356);
nor NOR4 (N3072, N3070, N214, N49, N2560);
not NOT1 (N3073, N3072);
or OR2 (N3074, N3060, N1281);
not NOT1 (N3075, N3073);
buf BUF1 (N3076, N3066);
buf BUF1 (N3077, N3049);
nand NAND4 (N3078, N3068, N1698, N1892, N3076);
or OR4 (N3079, N1619, N2670, N2287, N1526);
and AND4 (N3080, N3062, N1383, N1549, N2724);
buf BUF1 (N3081, N3075);
nand NAND3 (N3082, N3079, N759, N1849);
or OR4 (N3083, N3080, N1088, N2146, N128);
and AND3 (N3084, N3082, N618, N1566);
nor NOR3 (N3085, N3064, N538, N1583);
not NOT1 (N3086, N3084);
and AND4 (N3087, N3086, N944, N1335, N2259);
and AND3 (N3088, N3083, N2124, N640);
buf BUF1 (N3089, N3085);
xor XOR2 (N3090, N3077, N1392);
nand NAND2 (N3091, N3069, N1667);
nand NAND2 (N3092, N3087, N349);
not NOT1 (N3093, N3081);
nand NAND4 (N3094, N3074, N1198, N2482, N655);
xor XOR2 (N3095, N3094, N422);
or OR2 (N3096, N3091, N2064);
and AND2 (N3097, N3089, N2685);
or OR2 (N3098, N3092, N2950);
buf BUF1 (N3099, N3052);
nor NOR4 (N3100, N3097, N2751, N853, N2857);
nand NAND2 (N3101, N3100, N1004);
nor NOR4 (N3102, N3071, N2787, N2245, N1534);
xor XOR2 (N3103, N3090, N1878);
and AND2 (N3104, N3096, N2637);
nor NOR2 (N3105, N3098, N1185);
not NOT1 (N3106, N3104);
not NOT1 (N3107, N3095);
buf BUF1 (N3108, N3103);
or OR3 (N3109, N3108, N198, N1484);
or OR3 (N3110, N3105, N1651, N3051);
nor NOR4 (N3111, N3093, N2218, N1230, N2246);
nand NAND4 (N3112, N3110, N1266, N1181, N437);
buf BUF1 (N3113, N3107);
xor XOR2 (N3114, N3112, N2885);
nor NOR2 (N3115, N3109, N2402);
buf BUF1 (N3116, N3078);
and AND3 (N3117, N3111, N1800, N1838);
not NOT1 (N3118, N3113);
or OR2 (N3119, N3106, N2334);
or OR3 (N3120, N3119, N2806, N2136);
nand NAND4 (N3121, N3117, N30, N445, N2172);
not NOT1 (N3122, N3101);
xor XOR2 (N3123, N3088, N2672);
nand NAND4 (N3124, N3115, N1577, N1854, N1853);
and AND2 (N3125, N3124, N2035);
or OR4 (N3126, N3102, N2039, N2303, N568);
or OR2 (N3127, N3125, N812);
and AND2 (N3128, N3099, N690);
nor NOR4 (N3129, N3116, N2700, N2444, N25);
or OR2 (N3130, N3128, N2969);
and AND4 (N3131, N3118, N3014, N2631, N2991);
nand NAND4 (N3132, N3130, N161, N2326, N2167);
nand NAND4 (N3133, N3132, N2254, N1957, N2734);
nor NOR2 (N3134, N3129, N1725);
not NOT1 (N3135, N3122);
nand NAND4 (N3136, N3127, N2708, N3063, N2218);
nor NOR2 (N3137, N3135, N2668);
nand NAND4 (N3138, N3134, N1217, N1571, N2830);
xor XOR2 (N3139, N3120, N2497);
nor NOR2 (N3140, N3126, N1772);
nor NOR3 (N3141, N3139, N2656, N2763);
xor XOR2 (N3142, N3133, N2096);
not NOT1 (N3143, N3123);
buf BUF1 (N3144, N3131);
not NOT1 (N3145, N3136);
buf BUF1 (N3146, N3141);
nor NOR2 (N3147, N3140, N833);
and AND4 (N3148, N3143, N719, N2576, N252);
nor NOR2 (N3149, N3145, N2479);
not NOT1 (N3150, N3121);
buf BUF1 (N3151, N3146);
not NOT1 (N3152, N3144);
nand NAND3 (N3153, N3151, N2430, N259);
or OR2 (N3154, N3147, N1056);
nor NOR3 (N3155, N3149, N196, N1994);
nand NAND3 (N3156, N3148, N2409, N144);
xor XOR2 (N3157, N3142, N1838);
nor NOR3 (N3158, N3152, N557, N673);
nand NAND2 (N3159, N3157, N846);
xor XOR2 (N3160, N3156, N172);
xor XOR2 (N3161, N3158, N2833);
buf BUF1 (N3162, N3155);
and AND2 (N3163, N3162, N120);
xor XOR2 (N3164, N3159, N2038);
nand NAND4 (N3165, N3154, N383, N1, N2553);
or OR3 (N3166, N3137, N1225, N221);
or OR3 (N3167, N3161, N2691, N660);
buf BUF1 (N3168, N3114);
nand NAND4 (N3169, N3167, N344, N2948, N124);
nand NAND4 (N3170, N3160, N647, N2581, N1054);
not NOT1 (N3171, N3164);
nand NAND3 (N3172, N3169, N1913, N2805);
nor NOR3 (N3173, N3163, N2716, N943);
and AND4 (N3174, N3153, N2703, N1849, N1626);
not NOT1 (N3175, N3165);
or OR2 (N3176, N3175, N191);
nor NOR4 (N3177, N3150, N237, N1878, N2684);
nand NAND3 (N3178, N3166, N2656, N1094);
and AND2 (N3179, N3138, N1485);
xor XOR2 (N3180, N3170, N3059);
nand NAND3 (N3181, N3179, N2029, N2771);
nor NOR3 (N3182, N3180, N1071, N1843);
nand NAND4 (N3183, N3172, N2167, N1150, N264);
nor NOR4 (N3184, N3173, N1002, N108, N2955);
and AND3 (N3185, N3176, N598, N3066);
xor XOR2 (N3186, N3181, N1342);
or OR2 (N3187, N3174, N2115);
nand NAND4 (N3188, N3171, N375, N3177, N2717);
not NOT1 (N3189, N208);
buf BUF1 (N3190, N3189);
and AND3 (N3191, N3182, N932, N1840);
nor NOR4 (N3192, N3183, N167, N1527, N1651);
not NOT1 (N3193, N3192);
buf BUF1 (N3194, N3188);
or OR3 (N3195, N3190, N908, N3000);
nor NOR2 (N3196, N3191, N2324);
or OR2 (N3197, N3186, N1192);
nor NOR4 (N3198, N3197, N1426, N1727, N584);
nor NOR2 (N3199, N3168, N816);
or OR4 (N3200, N3194, N612, N3189, N1170);
nor NOR2 (N3201, N3178, N199);
or OR2 (N3202, N3196, N242);
nor NOR3 (N3203, N3199, N1946, N3008);
and AND3 (N3204, N3200, N300, N1808);
buf BUF1 (N3205, N3195);
nand NAND4 (N3206, N3198, N1606, N1127, N2233);
not NOT1 (N3207, N3202);
xor XOR2 (N3208, N3193, N892);
nand NAND3 (N3209, N3207, N563, N817);
not NOT1 (N3210, N3208);
xor XOR2 (N3211, N3185, N838);
xor XOR2 (N3212, N3204, N2539);
not NOT1 (N3213, N3205);
xor XOR2 (N3214, N3210, N188);
xor XOR2 (N3215, N3206, N2486);
and AND3 (N3216, N3209, N3084, N113);
not NOT1 (N3217, N3214);
nand NAND3 (N3218, N3217, N390, N359);
buf BUF1 (N3219, N3203);
nand NAND3 (N3220, N3184, N868, N843);
and AND3 (N3221, N3201, N1175, N811);
not NOT1 (N3222, N3216);
and AND3 (N3223, N3221, N3058, N1297);
nand NAND2 (N3224, N3212, N1251);
buf BUF1 (N3225, N3222);
not NOT1 (N3226, N3225);
xor XOR2 (N3227, N3220, N2763);
nor NOR2 (N3228, N3227, N683);
nand NAND4 (N3229, N3211, N320, N2348, N163);
or OR3 (N3230, N3219, N3228, N3162);
and AND2 (N3231, N1646, N1084);
buf BUF1 (N3232, N3187);
nand NAND3 (N3233, N3215, N2832, N2713);
and AND2 (N3234, N3223, N3022);
nand NAND4 (N3235, N3213, N1614, N2682, N998);
or OR2 (N3236, N3235, N1997);
nor NOR4 (N3237, N3236, N983, N71, N2419);
nand NAND2 (N3238, N3226, N772);
nand NAND4 (N3239, N3233, N2199, N2555, N2380);
nor NOR2 (N3240, N3230, N1306);
not NOT1 (N3241, N3240);
buf BUF1 (N3242, N3224);
xor XOR2 (N3243, N3238, N1113);
nand NAND2 (N3244, N3218, N503);
buf BUF1 (N3245, N3241);
not NOT1 (N3246, N3232);
nand NAND4 (N3247, N3242, N1406, N845, N2587);
nor NOR4 (N3248, N3245, N267, N266, N2182);
buf BUF1 (N3249, N3239);
nor NOR4 (N3250, N3246, N3206, N858, N2868);
nor NOR4 (N3251, N3244, N2890, N2334, N2099);
not NOT1 (N3252, N3251);
xor XOR2 (N3253, N3229, N177);
buf BUF1 (N3254, N3253);
nand NAND4 (N3255, N3254, N2980, N3010, N2831);
buf BUF1 (N3256, N3255);
nand NAND2 (N3257, N3243, N393);
nand NAND3 (N3258, N3234, N706, N1207);
nor NOR2 (N3259, N3257, N269);
and AND4 (N3260, N3249, N552, N2451, N2090);
not NOT1 (N3261, N3260);
or OR4 (N3262, N3256, N3004, N813, N74);
not NOT1 (N3263, N3248);
and AND3 (N3264, N3262, N3060, N2852);
or OR2 (N3265, N3263, N2534);
and AND2 (N3266, N3250, N395);
buf BUF1 (N3267, N3266);
nand NAND4 (N3268, N3237, N3196, N1343, N1612);
xor XOR2 (N3269, N3268, N1980);
xor XOR2 (N3270, N3258, N1122);
and AND2 (N3271, N3231, N2752);
and AND2 (N3272, N3270, N2133);
or OR2 (N3273, N3271, N3173);
nor NOR3 (N3274, N3247, N321, N649);
and AND2 (N3275, N3272, N2030);
or OR3 (N3276, N3264, N2473, N768);
nand NAND2 (N3277, N3274, N1905);
buf BUF1 (N3278, N3259);
and AND2 (N3279, N3278, N721);
not NOT1 (N3280, N3252);
and AND2 (N3281, N3275, N1380);
xor XOR2 (N3282, N3280, N468);
nand NAND3 (N3283, N3281, N1781, N2727);
nor NOR4 (N3284, N3265, N2623, N1155, N401);
and AND2 (N3285, N3276, N82);
buf BUF1 (N3286, N3269);
nand NAND4 (N3287, N3285, N380, N611, N1256);
buf BUF1 (N3288, N3284);
nand NAND4 (N3289, N3267, N1214, N2608, N3242);
buf BUF1 (N3290, N3283);
not NOT1 (N3291, N3288);
or OR2 (N3292, N3282, N2199);
buf BUF1 (N3293, N3261);
nand NAND3 (N3294, N3287, N2568, N1453);
buf BUF1 (N3295, N3290);
xor XOR2 (N3296, N3289, N2999);
nand NAND4 (N3297, N3291, N83, N2448, N1265);
buf BUF1 (N3298, N3277);
or OR3 (N3299, N3279, N1313, N1905);
and AND3 (N3300, N3286, N652, N2516);
or OR4 (N3301, N3296, N1826, N1951, N2819);
nor NOR2 (N3302, N3301, N2633);
xor XOR2 (N3303, N3292, N525);
not NOT1 (N3304, N3297);
nor NOR3 (N3305, N3295, N1300, N725);
buf BUF1 (N3306, N3302);
xor XOR2 (N3307, N3305, N2220);
or OR2 (N3308, N3306, N1938);
nand NAND4 (N3309, N3298, N1286, N1910, N2507);
or OR4 (N3310, N3304, N41, N562, N2522);
nand NAND4 (N3311, N3310, N2183, N645, N1311);
nor NOR4 (N3312, N3303, N1691, N1141, N1430);
or OR2 (N3313, N3312, N2864);
xor XOR2 (N3314, N3293, N2728);
xor XOR2 (N3315, N3273, N2281);
not NOT1 (N3316, N3315);
nand NAND3 (N3317, N3307, N2565, N2949);
not NOT1 (N3318, N3314);
or OR4 (N3319, N3309, N2920, N120, N60);
buf BUF1 (N3320, N3318);
and AND2 (N3321, N3294, N1554);
buf BUF1 (N3322, N3319);
buf BUF1 (N3323, N3317);
nor NOR3 (N3324, N3300, N925, N2869);
nand NAND4 (N3325, N3299, N1921, N2824, N1470);
or OR2 (N3326, N3316, N2415);
buf BUF1 (N3327, N3322);
xor XOR2 (N3328, N3323, N1586);
and AND3 (N3329, N3313, N578, N1776);
nor NOR2 (N3330, N3325, N600);
and AND2 (N3331, N3324, N471);
or OR4 (N3332, N3331, N2410, N3328, N1426);
nand NAND4 (N3333, N2325, N763, N1529, N865);
not NOT1 (N3334, N3330);
not NOT1 (N3335, N3320);
and AND2 (N3336, N3335, N2059);
or OR3 (N3337, N3327, N1822, N1219);
and AND3 (N3338, N3337, N2958, N722);
buf BUF1 (N3339, N3333);
or OR4 (N3340, N3321, N2526, N1401, N2992);
or OR4 (N3341, N3308, N3219, N1504, N2149);
not NOT1 (N3342, N3336);
buf BUF1 (N3343, N3311);
not NOT1 (N3344, N3326);
xor XOR2 (N3345, N3342, N1080);
nand NAND3 (N3346, N3341, N599, N3209);
or OR3 (N3347, N3345, N2871, N439);
and AND3 (N3348, N3339, N228, N2203);
and AND2 (N3349, N3332, N2733);
nor NOR4 (N3350, N3329, N3116, N2561, N2192);
xor XOR2 (N3351, N3334, N1448);
or OR4 (N3352, N3338, N1213, N1829, N467);
xor XOR2 (N3353, N3340, N2522);
xor XOR2 (N3354, N3352, N1567);
or OR4 (N3355, N3350, N2120, N698, N1152);
xor XOR2 (N3356, N3348, N3314);
buf BUF1 (N3357, N3343);
or OR3 (N3358, N3354, N947, N2499);
and AND4 (N3359, N3353, N1847, N229, N3004);
nand NAND3 (N3360, N3347, N1552, N2380);
buf BUF1 (N3361, N3359);
xor XOR2 (N3362, N3360, N1533);
xor XOR2 (N3363, N3358, N2004);
nand NAND3 (N3364, N3349, N3235, N2863);
xor XOR2 (N3365, N3356, N726);
and AND2 (N3366, N3361, N376);
xor XOR2 (N3367, N3346, N1249);
nand NAND4 (N3368, N3357, N2308, N3300, N735);
and AND4 (N3369, N3367, N2625, N1323, N888);
nand NAND2 (N3370, N3368, N843);
and AND3 (N3371, N3370, N2464, N3248);
not NOT1 (N3372, N3364);
or OR2 (N3373, N3344, N2033);
and AND3 (N3374, N3366, N391, N2938);
xor XOR2 (N3375, N3351, N319);
buf BUF1 (N3376, N3369);
and AND2 (N3377, N3371, N581);
buf BUF1 (N3378, N3373);
buf BUF1 (N3379, N3363);
or OR2 (N3380, N3375, N194);
nor NOR3 (N3381, N3380, N3125, N1826);
nand NAND2 (N3382, N3372, N3122);
nor NOR4 (N3383, N3374, N603, N3016, N1359);
nor NOR4 (N3384, N3365, N126, N2640, N461);
not NOT1 (N3385, N3383);
not NOT1 (N3386, N3355);
or OR2 (N3387, N3377, N1661);
nand NAND2 (N3388, N3376, N1095);
buf BUF1 (N3389, N3386);
nand NAND2 (N3390, N3378, N753);
nor NOR2 (N3391, N3389, N3125);
and AND4 (N3392, N3388, N376, N1009, N903);
and AND4 (N3393, N3362, N1185, N135, N1408);
nor NOR4 (N3394, N3382, N2181, N1320, N823);
xor XOR2 (N3395, N3394, N1194);
not NOT1 (N3396, N3381);
or OR3 (N3397, N3395, N266, N1529);
not NOT1 (N3398, N3391);
nor NOR3 (N3399, N3385, N3127, N1149);
nor NOR3 (N3400, N3399, N2874, N1244);
or OR2 (N3401, N3384, N3355);
and AND2 (N3402, N3393, N429);
nand NAND3 (N3403, N3392, N796, N274);
buf BUF1 (N3404, N3397);
nand NAND3 (N3405, N3400, N1563, N1838);
not NOT1 (N3406, N3403);
buf BUF1 (N3407, N3390);
and AND4 (N3408, N3379, N441, N496, N2056);
not NOT1 (N3409, N3396);
and AND4 (N3410, N3401, N1061, N821, N784);
buf BUF1 (N3411, N3409);
nand NAND2 (N3412, N3404, N1368);
xor XOR2 (N3413, N3412, N2864);
or OR4 (N3414, N3405, N1241, N482, N801);
nand NAND2 (N3415, N3398, N1593);
not NOT1 (N3416, N3411);
or OR3 (N3417, N3407, N3132, N3228);
and AND4 (N3418, N3415, N999, N1144, N1648);
nor NOR2 (N3419, N3406, N2228);
or OR4 (N3420, N3408, N1121, N1352, N985);
nand NAND4 (N3421, N3416, N2262, N2795, N399);
xor XOR2 (N3422, N3387, N464);
and AND2 (N3423, N3419, N1850);
buf BUF1 (N3424, N3420);
xor XOR2 (N3425, N3423, N2934);
and AND3 (N3426, N3424, N1253, N1922);
nor NOR4 (N3427, N3422, N1492, N2882, N3389);
or OR3 (N3428, N3427, N462, N980);
nand NAND2 (N3429, N3414, N2574);
and AND2 (N3430, N3425, N99);
buf BUF1 (N3431, N3430);
nand NAND2 (N3432, N3413, N1102);
and AND2 (N3433, N3432, N959);
or OR3 (N3434, N3410, N2001, N3184);
nand NAND4 (N3435, N3431, N2344, N397, N1704);
not NOT1 (N3436, N3429);
xor XOR2 (N3437, N3436, N1897);
or OR4 (N3438, N3426, N615, N1686, N2627);
not NOT1 (N3439, N3418);
xor XOR2 (N3440, N3402, N1313);
not NOT1 (N3441, N3440);
or OR4 (N3442, N3428, N785, N574, N830);
xor XOR2 (N3443, N3439, N2882);
nand NAND4 (N3444, N3421, N1439, N2532, N3101);
or OR3 (N3445, N3443, N2488, N2430);
nand NAND3 (N3446, N3435, N3169, N276);
or OR3 (N3447, N3433, N410, N3112);
nand NAND4 (N3448, N3447, N2865, N538, N4);
or OR3 (N3449, N3417, N2706, N2870);
xor XOR2 (N3450, N3444, N2773);
nand NAND4 (N3451, N3448, N867, N15, N1669);
or OR2 (N3452, N3445, N2633);
xor XOR2 (N3453, N3451, N1085);
not NOT1 (N3454, N3437);
buf BUF1 (N3455, N3450);
nor NOR3 (N3456, N3449, N1249, N3377);
or OR4 (N3457, N3454, N739, N1285, N3097);
and AND2 (N3458, N3453, N2203);
nor NOR4 (N3459, N3438, N2327, N1489, N1527);
nand NAND4 (N3460, N3458, N1053, N2001, N1856);
or OR3 (N3461, N3446, N2851, N1018);
or OR3 (N3462, N3441, N448, N3106);
and AND2 (N3463, N3462, N2532);
nor NOR2 (N3464, N3459, N3114);
nor NOR2 (N3465, N3464, N2636);
or OR3 (N3466, N3442, N654, N2942);
nor NOR2 (N3467, N3465, N1492);
nand NAND3 (N3468, N3452, N1993, N3316);
and AND4 (N3469, N3466, N97, N1014, N1401);
xor XOR2 (N3470, N3469, N2221);
xor XOR2 (N3471, N3461, N1469);
xor XOR2 (N3472, N3460, N2738);
or OR4 (N3473, N3472, N1776, N1135, N54);
nor NOR4 (N3474, N3457, N1759, N574, N155);
buf BUF1 (N3475, N3467);
not NOT1 (N3476, N3473);
buf BUF1 (N3477, N3463);
buf BUF1 (N3478, N3434);
and AND2 (N3479, N3468, N2952);
or OR4 (N3480, N3474, N581, N557, N1119);
xor XOR2 (N3481, N3478, N1785);
or OR4 (N3482, N3455, N3110, N165, N1778);
xor XOR2 (N3483, N3476, N3178);
buf BUF1 (N3484, N3481);
xor XOR2 (N3485, N3483, N2352);
not NOT1 (N3486, N3480);
or OR4 (N3487, N3477, N210, N2808, N1371);
and AND4 (N3488, N3486, N2655, N2777, N102);
or OR2 (N3489, N3479, N2817);
and AND4 (N3490, N3488, N2110, N982, N2835);
nor NOR2 (N3491, N3484, N1672);
xor XOR2 (N3492, N3456, N683);
buf BUF1 (N3493, N3485);
buf BUF1 (N3494, N3471);
and AND2 (N3495, N3482, N2133);
not NOT1 (N3496, N3487);
nor NOR3 (N3497, N3495, N2821, N2249);
and AND3 (N3498, N3470, N2984, N1911);
nor NOR4 (N3499, N3489, N3306, N3187, N3162);
nand NAND3 (N3500, N3494, N39, N3270);
buf BUF1 (N3501, N3475);
and AND2 (N3502, N3491, N584);
xor XOR2 (N3503, N3497, N2694);
xor XOR2 (N3504, N3501, N2802);
not NOT1 (N3505, N3492);
xor XOR2 (N3506, N3499, N399);
nand NAND2 (N3507, N3490, N315);
or OR4 (N3508, N3500, N966, N3395, N3297);
nor NOR3 (N3509, N3502, N1205, N2379);
nor NOR2 (N3510, N3498, N3250);
xor XOR2 (N3511, N3506, N2371);
xor XOR2 (N3512, N3507, N791);
or OR4 (N3513, N3504, N1752, N15, N3406);
or OR3 (N3514, N3509, N1069, N982);
or OR3 (N3515, N3496, N1178, N3360);
buf BUF1 (N3516, N3511);
nor NOR4 (N3517, N3503, N3113, N2563, N465);
and AND3 (N3518, N3517, N2380, N1664);
xor XOR2 (N3519, N3493, N2576);
buf BUF1 (N3520, N3505);
nor NOR3 (N3521, N3518, N1810, N180);
nor NOR3 (N3522, N3519, N2142, N2719);
nand NAND2 (N3523, N3515, N2121);
not NOT1 (N3524, N3516);
buf BUF1 (N3525, N3512);
or OR4 (N3526, N3514, N179, N2135, N1578);
nand NAND3 (N3527, N3523, N390, N2242);
and AND2 (N3528, N3510, N2977);
and AND2 (N3529, N3521, N2373);
xor XOR2 (N3530, N3513, N701);
and AND4 (N3531, N3527, N725, N3361, N2345);
not NOT1 (N3532, N3530);
nor NOR2 (N3533, N3525, N2316);
and AND4 (N3534, N3522, N2731, N2068, N528);
nor NOR2 (N3535, N3534, N39);
buf BUF1 (N3536, N3533);
nand NAND4 (N3537, N3536, N870, N2568, N3372);
or OR3 (N3538, N3508, N1531, N1107);
buf BUF1 (N3539, N3528);
xor XOR2 (N3540, N3520, N2708);
or OR3 (N3541, N3524, N278, N257);
nor NOR4 (N3542, N3532, N642, N1298, N474);
and AND2 (N3543, N3541, N2597);
or OR3 (N3544, N3529, N3333, N2702);
xor XOR2 (N3545, N3543, N1179);
buf BUF1 (N3546, N3535);
and AND4 (N3547, N3538, N3543, N1980, N1097);
not NOT1 (N3548, N3539);
and AND3 (N3549, N3540, N445, N1339);
or OR3 (N3550, N3547, N536, N2249);
nand NAND3 (N3551, N3544, N1348, N2386);
buf BUF1 (N3552, N3546);
and AND4 (N3553, N3545, N3283, N2786, N2827);
nand NAND2 (N3554, N3550, N2850);
and AND3 (N3555, N3526, N2054, N2953);
xor XOR2 (N3556, N3551, N2031);
buf BUF1 (N3557, N3531);
buf BUF1 (N3558, N3557);
buf BUF1 (N3559, N3537);
buf BUF1 (N3560, N3555);
buf BUF1 (N3561, N3558);
not NOT1 (N3562, N3549);
nand NAND3 (N3563, N3552, N1055, N443);
not NOT1 (N3564, N3559);
not NOT1 (N3565, N3554);
nor NOR3 (N3566, N3561, N2090, N949);
or OR3 (N3567, N3566, N1758, N1373);
nor NOR2 (N3568, N3553, N931);
or OR4 (N3569, N3567, N241, N1697, N159);
nand NAND4 (N3570, N3565, N1106, N2561, N1173);
and AND3 (N3571, N3560, N2969, N937);
nor NOR4 (N3572, N3548, N3504, N3506, N1582);
buf BUF1 (N3573, N3571);
buf BUF1 (N3574, N3564);
and AND2 (N3575, N3570, N580);
or OR3 (N3576, N3568, N2172, N1144);
not NOT1 (N3577, N3574);
nand NAND2 (N3578, N3542, N1613);
not NOT1 (N3579, N3573);
or OR3 (N3580, N3562, N970, N628);
buf BUF1 (N3581, N3580);
nand NAND2 (N3582, N3579, N2943);
not NOT1 (N3583, N3563);
xor XOR2 (N3584, N3575, N3399);
or OR4 (N3585, N3576, N3317, N1768, N1443);
not NOT1 (N3586, N3582);
xor XOR2 (N3587, N3569, N893);
or OR2 (N3588, N3578, N734);
and AND3 (N3589, N3585, N2082, N327);
xor XOR2 (N3590, N3588, N344);
nor NOR3 (N3591, N3581, N3344, N3321);
or OR3 (N3592, N3586, N1860, N354);
nor NOR4 (N3593, N3589, N3565, N1968, N509);
not NOT1 (N3594, N3592);
xor XOR2 (N3595, N3556, N3229);
nor NOR2 (N3596, N3577, N1493);
or OR3 (N3597, N3595, N2188, N1986);
nand NAND3 (N3598, N3591, N1722, N366);
and AND3 (N3599, N3584, N1818, N2513);
and AND4 (N3600, N3590, N1212, N1671, N948);
buf BUF1 (N3601, N3583);
xor XOR2 (N3602, N3600, N2383);
not NOT1 (N3603, N3572);
and AND2 (N3604, N3599, N217);
nor NOR2 (N3605, N3604, N3588);
nand NAND4 (N3606, N3598, N1676, N2419, N1263);
xor XOR2 (N3607, N3587, N615);
or OR2 (N3608, N3607, N1900);
xor XOR2 (N3609, N3606, N1468);
or OR3 (N3610, N3594, N1250, N2416);
not NOT1 (N3611, N3608);
xor XOR2 (N3612, N3597, N3346);
and AND3 (N3613, N3610, N1638, N1582);
not NOT1 (N3614, N3612);
nand NAND4 (N3615, N3602, N2933, N2263, N2078);
buf BUF1 (N3616, N3609);
buf BUF1 (N3617, N3614);
or OR2 (N3618, N3596, N653);
nor NOR2 (N3619, N3611, N1278);
or OR2 (N3620, N3617, N3515);
not NOT1 (N3621, N3603);
and AND4 (N3622, N3616, N2742, N3062, N2291);
not NOT1 (N3623, N3622);
nand NAND2 (N3624, N3618, N3008);
nand NAND3 (N3625, N3620, N2017, N1622);
nand NAND3 (N3626, N3593, N201, N1307);
not NOT1 (N3627, N3615);
or OR3 (N3628, N3624, N1502, N2973);
or OR4 (N3629, N3625, N153, N1174, N3089);
or OR2 (N3630, N3623, N1205);
or OR3 (N3631, N3626, N3625, N2015);
or OR2 (N3632, N3629, N67);
and AND2 (N3633, N3628, N2068);
or OR2 (N3634, N3630, N1165);
xor XOR2 (N3635, N3633, N2336);
and AND4 (N3636, N3605, N1273, N2009, N1238);
nand NAND4 (N3637, N3613, N1289, N1524, N3117);
nor NOR4 (N3638, N3637, N2013, N1897, N1334);
nand NAND3 (N3639, N3638, N1472, N3134);
buf BUF1 (N3640, N3634);
or OR3 (N3641, N3601, N1815, N2700);
not NOT1 (N3642, N3619);
nand NAND4 (N3643, N3635, N3219, N1044, N3350);
not NOT1 (N3644, N3640);
and AND2 (N3645, N3644, N65);
nand NAND3 (N3646, N3645, N2071, N1978);
xor XOR2 (N3647, N3643, N413);
nand NAND3 (N3648, N3632, N1956, N1330);
buf BUF1 (N3649, N3642);
nor NOR3 (N3650, N3639, N3576, N2108);
and AND2 (N3651, N3650, N426);
nand NAND2 (N3652, N3621, N1125);
xor XOR2 (N3653, N3652, N650);
xor XOR2 (N3654, N3627, N2235);
buf BUF1 (N3655, N3649);
buf BUF1 (N3656, N3631);
xor XOR2 (N3657, N3656, N1332);
not NOT1 (N3658, N3646);
or OR3 (N3659, N3657, N728, N1694);
nor NOR4 (N3660, N3658, N1964, N119, N542);
nand NAND4 (N3661, N3655, N2873, N1847, N3198);
not NOT1 (N3662, N3659);
or OR4 (N3663, N3653, N1118, N2969, N225);
not NOT1 (N3664, N3647);
nand NAND2 (N3665, N3663, N2705);
not NOT1 (N3666, N3641);
xor XOR2 (N3667, N3664, N2393);
and AND4 (N3668, N3660, N998, N1263, N1921);
and AND4 (N3669, N3662, N948, N2500, N715);
not NOT1 (N3670, N3654);
buf BUF1 (N3671, N3665);
buf BUF1 (N3672, N3661);
nand NAND3 (N3673, N3636, N2969, N1254);
not NOT1 (N3674, N3671);
not NOT1 (N3675, N3673);
or OR4 (N3676, N3670, N2137, N438, N95);
not NOT1 (N3677, N3668);
or OR3 (N3678, N3666, N1359, N2875);
buf BUF1 (N3679, N3674);
buf BUF1 (N3680, N3679);
and AND3 (N3681, N3667, N2699, N479);
xor XOR2 (N3682, N3681, N3075);
xor XOR2 (N3683, N3682, N143);
nor NOR4 (N3684, N3680, N2942, N430, N2675);
nand NAND3 (N3685, N3683, N2083, N434);
buf BUF1 (N3686, N3684);
and AND2 (N3687, N3686, N920);
buf BUF1 (N3688, N3648);
and AND2 (N3689, N3669, N1440);
nand NAND4 (N3690, N3688, N1822, N3334, N507);
nand NAND4 (N3691, N3690, N2392, N1473, N522);
not NOT1 (N3692, N3677);
buf BUF1 (N3693, N3691);
or OR4 (N3694, N3692, N70, N1336, N2686);
nor NOR4 (N3695, N3689, N3491, N3674, N697);
not NOT1 (N3696, N3694);
nor NOR3 (N3697, N3696, N556, N2420);
or OR3 (N3698, N3695, N2591, N1346);
xor XOR2 (N3699, N3651, N938);
or OR2 (N3700, N3687, N1392);
buf BUF1 (N3701, N3675);
nand NAND3 (N3702, N3676, N1216, N422);
or OR3 (N3703, N3672, N2865, N3622);
buf BUF1 (N3704, N3700);
not NOT1 (N3705, N3697);
not NOT1 (N3706, N3701);
buf BUF1 (N3707, N3685);
and AND4 (N3708, N3707, N715, N3696, N1782);
nand NAND3 (N3709, N3705, N2506, N1241);
nand NAND3 (N3710, N3693, N2920, N2846);
not NOT1 (N3711, N3704);
xor XOR2 (N3712, N3698, N797);
xor XOR2 (N3713, N3678, N2794);
buf BUF1 (N3714, N3710);
nor NOR2 (N3715, N3711, N504);
xor XOR2 (N3716, N3713, N1232);
and AND3 (N3717, N3716, N2802, N3667);
nor NOR2 (N3718, N3708, N867);
xor XOR2 (N3719, N3718, N838);
or OR4 (N3720, N3714, N3120, N1240, N1464);
nor NOR2 (N3721, N3703, N23);
nand NAND4 (N3722, N3721, N2673, N3016, N684);
or OR3 (N3723, N3715, N1280, N2772);
nor NOR3 (N3724, N3717, N3247, N1893);
xor XOR2 (N3725, N3699, N304);
nor NOR2 (N3726, N3719, N1725);
nor NOR3 (N3727, N3726, N1262, N2445);
xor XOR2 (N3728, N3706, N2364);
xor XOR2 (N3729, N3723, N1163);
or OR4 (N3730, N3729, N536, N2354, N1342);
not NOT1 (N3731, N3702);
nor NOR3 (N3732, N3725, N3238, N458);
nor NOR4 (N3733, N3727, N30, N1448, N1764);
nand NAND2 (N3734, N3733, N1797);
nand NAND4 (N3735, N3712, N208, N3666, N1771);
buf BUF1 (N3736, N3734);
xor XOR2 (N3737, N3736, N2649);
not NOT1 (N3738, N3737);
buf BUF1 (N3739, N3735);
not NOT1 (N3740, N3732);
not NOT1 (N3741, N3739);
nor NOR4 (N3742, N3728, N916, N3442, N2259);
and AND2 (N3743, N3742, N3359);
nand NAND2 (N3744, N3720, N1056);
xor XOR2 (N3745, N3731, N3317);
nor NOR3 (N3746, N3722, N290, N640);
buf BUF1 (N3747, N3744);
not NOT1 (N3748, N3709);
xor XOR2 (N3749, N3738, N2511);
or OR3 (N3750, N3749, N1342, N220);
and AND2 (N3751, N3746, N1553);
and AND3 (N3752, N3751, N229, N2781);
xor XOR2 (N3753, N3724, N119);
nor NOR3 (N3754, N3743, N2139, N2417);
and AND3 (N3755, N3745, N1577, N2244);
or OR3 (N3756, N3748, N977, N551);
not NOT1 (N3757, N3756);
not NOT1 (N3758, N3753);
buf BUF1 (N3759, N3747);
not NOT1 (N3760, N3754);
nor NOR4 (N3761, N3741, N3642, N353, N1118);
buf BUF1 (N3762, N3755);
not NOT1 (N3763, N3761);
not NOT1 (N3764, N3757);
or OR2 (N3765, N3752, N810);
not NOT1 (N3766, N3740);
nor NOR3 (N3767, N3763, N1019, N3155);
buf BUF1 (N3768, N3760);
xor XOR2 (N3769, N3759, N2069);
or OR4 (N3770, N3750, N495, N1815, N1906);
and AND2 (N3771, N3764, N1274);
and AND4 (N3772, N3766, N3729, N2410, N1844);
xor XOR2 (N3773, N3772, N2852);
not NOT1 (N3774, N3730);
or OR2 (N3775, N3765, N2766);
not NOT1 (N3776, N3769);
xor XOR2 (N3777, N3771, N197);
nor NOR2 (N3778, N3758, N1879);
and AND2 (N3779, N3770, N1571);
nand NAND3 (N3780, N3779, N5, N1012);
buf BUF1 (N3781, N3780);
xor XOR2 (N3782, N3768, N160);
not NOT1 (N3783, N3776);
and AND3 (N3784, N3777, N2197, N1161);
not NOT1 (N3785, N3782);
and AND3 (N3786, N3774, N3487, N1416);
and AND3 (N3787, N3762, N1909, N2983);
and AND2 (N3788, N3775, N975);
or OR2 (N3789, N3788, N1239);
and AND2 (N3790, N3786, N2477);
and AND3 (N3791, N3778, N1555, N2153);
not NOT1 (N3792, N3781);
and AND4 (N3793, N3787, N1948, N1088, N1285);
xor XOR2 (N3794, N3773, N436);
not NOT1 (N3795, N3792);
xor XOR2 (N3796, N3785, N2282);
or OR3 (N3797, N3791, N2452, N2309);
or OR3 (N3798, N3783, N997, N2415);
nand NAND3 (N3799, N3789, N1713, N2737);
buf BUF1 (N3800, N3797);
nand NAND2 (N3801, N3796, N884);
or OR4 (N3802, N3794, N1056, N1998, N1698);
xor XOR2 (N3803, N3798, N3735);
not NOT1 (N3804, N3795);
and AND2 (N3805, N3803, N3149);
nand NAND4 (N3806, N3790, N113, N332, N3118);
nand NAND3 (N3807, N3804, N3344, N3182);
and AND2 (N3808, N3784, N2444);
not NOT1 (N3809, N3802);
xor XOR2 (N3810, N3809, N660);
not NOT1 (N3811, N3807);
and AND2 (N3812, N3793, N897);
buf BUF1 (N3813, N3812);
or OR4 (N3814, N3805, N1456, N1869, N2041);
xor XOR2 (N3815, N3801, N2429);
nor NOR4 (N3816, N3815, N111, N3558, N1041);
xor XOR2 (N3817, N3767, N2189);
nor NOR2 (N3818, N3813, N456);
and AND3 (N3819, N3814, N2735, N435);
buf BUF1 (N3820, N3819);
or OR4 (N3821, N3820, N175, N1512, N2178);
or OR4 (N3822, N3800, N2950, N1991, N2143);
nor NOR4 (N3823, N3818, N30, N914, N381);
not NOT1 (N3824, N3811);
xor XOR2 (N3825, N3808, N543);
buf BUF1 (N3826, N3824);
nand NAND3 (N3827, N3823, N802, N1145);
and AND2 (N3828, N3799, N2990);
xor XOR2 (N3829, N3817, N2362);
xor XOR2 (N3830, N3829, N2460);
buf BUF1 (N3831, N3816);
nand NAND4 (N3832, N3806, N2229, N3309, N3596);
or OR4 (N3833, N3830, N2863, N1629, N1728);
or OR4 (N3834, N3826, N2790, N322, N3377);
and AND3 (N3835, N3821, N1738, N3701);
and AND4 (N3836, N3822, N262, N3333, N681);
nor NOR2 (N3837, N3836, N1298);
nor NOR4 (N3838, N3834, N120, N363, N1987);
and AND3 (N3839, N3825, N2126, N2627);
buf BUF1 (N3840, N3810);
and AND3 (N3841, N3835, N2049, N3314);
and AND2 (N3842, N3828, N2871);
and AND4 (N3843, N3831, N417, N2449, N2662);
xor XOR2 (N3844, N3833, N2796);
or OR4 (N3845, N3844, N65, N276, N1122);
buf BUF1 (N3846, N3842);
not NOT1 (N3847, N3839);
nor NOR4 (N3848, N3847, N3589, N1978, N533);
not NOT1 (N3849, N3848);
or OR4 (N3850, N3843, N185, N1330, N1925);
or OR4 (N3851, N3832, N3122, N609, N2917);
and AND4 (N3852, N3851, N1028, N2756, N781);
or OR2 (N3853, N3840, N1087);
xor XOR2 (N3854, N3852, N3099);
buf BUF1 (N3855, N3845);
and AND3 (N3856, N3854, N722, N1825);
not NOT1 (N3857, N3846);
or OR4 (N3858, N3841, N3401, N987, N2622);
and AND4 (N3859, N3856, N1227, N2210, N3837);
nand NAND4 (N3860, N3045, N1462, N799, N419);
xor XOR2 (N3861, N3853, N2767);
or OR3 (N3862, N3860, N1562, N3377);
nor NOR4 (N3863, N3850, N3478, N1898, N1104);
not NOT1 (N3864, N3861);
not NOT1 (N3865, N3849);
buf BUF1 (N3866, N3838);
nand NAND4 (N3867, N3859, N143, N3315, N308);
not NOT1 (N3868, N3827);
and AND3 (N3869, N3855, N1282, N1020);
xor XOR2 (N3870, N3864, N2038);
or OR4 (N3871, N3865, N1234, N1201, N1332);
nand NAND2 (N3872, N3858, N3592);
xor XOR2 (N3873, N3872, N521);
nor NOR2 (N3874, N3857, N1249);
nor NOR3 (N3875, N3863, N3031, N2649);
nand NAND4 (N3876, N3871, N277, N3024, N1431);
buf BUF1 (N3877, N3862);
not NOT1 (N3878, N3870);
and AND3 (N3879, N3878, N997, N1511);
not NOT1 (N3880, N3866);
xor XOR2 (N3881, N3869, N2653);
or OR4 (N3882, N3876, N95, N2779, N2066);
nor NOR2 (N3883, N3880, N1383);
buf BUF1 (N3884, N3875);
or OR2 (N3885, N3867, N2864);
buf BUF1 (N3886, N3884);
not NOT1 (N3887, N3879);
nand NAND3 (N3888, N3886, N1057, N2958);
nor NOR4 (N3889, N3888, N578, N1976, N2054);
and AND4 (N3890, N3868, N696, N495, N2329);
xor XOR2 (N3891, N3890, N2514);
xor XOR2 (N3892, N3874, N421);
and AND3 (N3893, N3889, N1653, N778);
and AND4 (N3894, N3877, N2833, N1714, N2556);
nor NOR2 (N3895, N3894, N2500);
and AND3 (N3896, N3887, N2376, N983);
and AND3 (N3897, N3883, N2697, N603);
nor NOR4 (N3898, N3873, N384, N2853, N995);
buf BUF1 (N3899, N3897);
and AND4 (N3900, N3885, N1667, N1332, N2628);
not NOT1 (N3901, N3882);
and AND3 (N3902, N3898, N2779, N2246);
buf BUF1 (N3903, N3891);
not NOT1 (N3904, N3896);
buf BUF1 (N3905, N3900);
nor NOR3 (N3906, N3899, N2335, N1101);
not NOT1 (N3907, N3895);
nor NOR4 (N3908, N3901, N2458, N2668, N425);
xor XOR2 (N3909, N3881, N1951);
buf BUF1 (N3910, N3893);
not NOT1 (N3911, N3903);
or OR4 (N3912, N3906, N2682, N2719, N2990);
xor XOR2 (N3913, N3907, N2400);
nand NAND4 (N3914, N3913, N3232, N1249, N1737);
or OR3 (N3915, N3912, N2091, N3761);
nor NOR4 (N3916, N3909, N1535, N796, N2700);
nand NAND3 (N3917, N3892, N2184, N1250);
xor XOR2 (N3918, N3911, N1304);
not NOT1 (N3919, N3905);
buf BUF1 (N3920, N3914);
buf BUF1 (N3921, N3910);
nand NAND4 (N3922, N3919, N3079, N3767, N2157);
xor XOR2 (N3923, N3916, N719);
nand NAND3 (N3924, N3920, N1426, N3894);
nand NAND2 (N3925, N3918, N1834);
xor XOR2 (N3926, N3902, N1928);
nor NOR3 (N3927, N3924, N3589, N2580);
not NOT1 (N3928, N3926);
or OR3 (N3929, N3921, N776, N1503);
not NOT1 (N3930, N3927);
not NOT1 (N3931, N3928);
xor XOR2 (N3932, N3904, N2983);
and AND4 (N3933, N3931, N1570, N3547, N1436);
buf BUF1 (N3934, N3932);
and AND2 (N3935, N3925, N1875);
and AND4 (N3936, N3930, N2597, N3373, N3232);
and AND3 (N3937, N3933, N927, N2507);
xor XOR2 (N3938, N3935, N892);
buf BUF1 (N3939, N3936);
xor XOR2 (N3940, N3915, N1976);
or OR3 (N3941, N3934, N2307, N674);
xor XOR2 (N3942, N3922, N254);
nand NAND4 (N3943, N3938, N3871, N1161, N1060);
and AND3 (N3944, N3939, N2838, N3930);
or OR2 (N3945, N3943, N2312);
not NOT1 (N3946, N3929);
not NOT1 (N3947, N3923);
buf BUF1 (N3948, N3942);
nand NAND2 (N3949, N3948, N1250);
nor NOR3 (N3950, N3947, N3251, N3481);
buf BUF1 (N3951, N3917);
xor XOR2 (N3952, N3940, N3468);
buf BUF1 (N3953, N3950);
and AND4 (N3954, N3945, N1607, N1086, N2412);
nor NOR4 (N3955, N3944, N1692, N523, N3183);
xor XOR2 (N3956, N3908, N2917);
and AND4 (N3957, N3956, N1538, N2317, N1436);
nor NOR4 (N3958, N3952, N319, N3418, N2274);
or OR3 (N3959, N3951, N628, N2092);
nand NAND3 (N3960, N3955, N2160, N3351);
nor NOR3 (N3961, N3959, N3117, N2380);
not NOT1 (N3962, N3946);
xor XOR2 (N3963, N3960, N2904);
and AND3 (N3964, N3954, N762, N3279);
not NOT1 (N3965, N3962);
nand NAND2 (N3966, N3957, N2971);
not NOT1 (N3967, N3966);
and AND2 (N3968, N3953, N154);
not NOT1 (N3969, N3941);
buf BUF1 (N3970, N3965);
xor XOR2 (N3971, N3970, N1271);
or OR3 (N3972, N3968, N982, N1792);
nor NOR3 (N3973, N3967, N2489, N880);
or OR3 (N3974, N3971, N2650, N759);
nand NAND2 (N3975, N3974, N984);
not NOT1 (N3976, N3964);
or OR4 (N3977, N3937, N2702, N1816, N1700);
buf BUF1 (N3978, N3963);
nand NAND4 (N3979, N3975, N97, N3862, N3789);
xor XOR2 (N3980, N3978, N2587);
or OR2 (N3981, N3980, N3153);
not NOT1 (N3982, N3977);
buf BUF1 (N3983, N3972);
or OR3 (N3984, N3961, N1223, N2806);
and AND2 (N3985, N3949, N2821);
not NOT1 (N3986, N3984);
buf BUF1 (N3987, N3976);
buf BUF1 (N3988, N3986);
xor XOR2 (N3989, N3958, N2097);
or OR2 (N3990, N3983, N3520);
xor XOR2 (N3991, N3988, N1973);
and AND4 (N3992, N3973, N530, N1214, N2812);
not NOT1 (N3993, N3989);
buf BUF1 (N3994, N3991);
not NOT1 (N3995, N3990);
not NOT1 (N3996, N3992);
nor NOR2 (N3997, N3985, N2547);
nor NOR4 (N3998, N3979, N2408, N2215, N705);
nor NOR3 (N3999, N3996, N512, N277);
not NOT1 (N4000, N3995);
nand NAND2 (N4001, N3994, N1585);
xor XOR2 (N4002, N3998, N2962);
nand NAND3 (N4003, N3993, N227, N3981);
not NOT1 (N4004, N789);
not NOT1 (N4005, N3982);
buf BUF1 (N4006, N4004);
xor XOR2 (N4007, N3969, N1007);
or OR2 (N4008, N4001, N1000);
or OR4 (N4009, N4005, N1688, N3861, N2557);
buf BUF1 (N4010, N3987);
buf BUF1 (N4011, N4006);
or OR3 (N4012, N4008, N294, N915);
nor NOR2 (N4013, N4009, N2945);
and AND2 (N4014, N4010, N426);
not NOT1 (N4015, N4007);
nor NOR2 (N4016, N4015, N244);
not NOT1 (N4017, N4002);
or OR3 (N4018, N4017, N3153, N3788);
xor XOR2 (N4019, N4012, N533);
nor NOR3 (N4020, N4014, N1311, N1242);
nand NAND3 (N4021, N4003, N1271, N1362);
buf BUF1 (N4022, N4013);
not NOT1 (N4023, N4000);
and AND3 (N4024, N4018, N3249, N3952);
and AND4 (N4025, N3999, N2687, N1570, N2306);
nor NOR2 (N4026, N3997, N1470);
nor NOR4 (N4027, N4026, N2161, N3484, N1833);
nor NOR2 (N4028, N4020, N3011);
nand NAND4 (N4029, N4027, N1673, N2506, N13);
nand NAND4 (N4030, N4019, N2941, N357, N1293);
xor XOR2 (N4031, N4023, N1982);
nand NAND4 (N4032, N4011, N3787, N1338, N681);
nor NOR4 (N4033, N4022, N487, N806, N1635);
or OR4 (N4034, N4029, N3817, N1698, N1142);
not NOT1 (N4035, N4030);
buf BUF1 (N4036, N4021);
nor NOR3 (N4037, N4032, N2882, N3292);
or OR4 (N4038, N4016, N3754, N1808, N1271);
and AND4 (N4039, N4025, N2965, N1796, N2813);
not NOT1 (N4040, N4037);
nor NOR4 (N4041, N4034, N3863, N330, N4007);
nand NAND3 (N4042, N4028, N3425, N1508);
nor NOR2 (N4043, N4033, N3313);
nand NAND3 (N4044, N4041, N2039, N895);
not NOT1 (N4045, N4036);
xor XOR2 (N4046, N4031, N2122);
xor XOR2 (N4047, N4045, N3605);
nor NOR3 (N4048, N4038, N3004, N2654);
not NOT1 (N4049, N4048);
and AND3 (N4050, N4024, N730, N2441);
and AND2 (N4051, N4047, N970);
nor NOR3 (N4052, N4035, N821, N1356);
nor NOR3 (N4053, N4052, N689, N2940);
buf BUF1 (N4054, N4044);
or OR2 (N4055, N4051, N2323);
and AND3 (N4056, N4046, N1131, N1167);
not NOT1 (N4057, N4042);
nor NOR2 (N4058, N4054, N12);
buf BUF1 (N4059, N4055);
xor XOR2 (N4060, N4050, N3026);
nor NOR4 (N4061, N4059, N2910, N370, N264);
or OR4 (N4062, N4053, N2618, N2409, N1383);
and AND3 (N4063, N4062, N3315, N2230);
nand NAND2 (N4064, N4058, N847);
xor XOR2 (N4065, N4039, N3113);
buf BUF1 (N4066, N4060);
and AND3 (N4067, N4057, N2762, N4028);
buf BUF1 (N4068, N4061);
xor XOR2 (N4069, N4043, N1974);
buf BUF1 (N4070, N4066);
nand NAND2 (N4071, N4067, N1657);
not NOT1 (N4072, N4065);
buf BUF1 (N4073, N4071);
xor XOR2 (N4074, N4068, N247);
xor XOR2 (N4075, N4070, N1595);
xor XOR2 (N4076, N4069, N1357);
or OR3 (N4077, N4049, N4064, N2616);
and AND2 (N4078, N1402, N3712);
and AND4 (N4079, N4073, N3384, N2690, N4073);
and AND2 (N4080, N4077, N2080);
or OR2 (N4081, N4072, N2416);
and AND3 (N4082, N4063, N1157, N3980);
nor NOR2 (N4083, N4040, N3306);
nand NAND3 (N4084, N4081, N2243, N1082);
or OR4 (N4085, N4083, N1251, N250, N1776);
xor XOR2 (N4086, N4084, N670);
and AND2 (N4087, N4082, N3782);
and AND3 (N4088, N4076, N1674, N392);
xor XOR2 (N4089, N4085, N3701);
xor XOR2 (N4090, N4088, N600);
or OR3 (N4091, N4089, N1232, N3302);
or OR2 (N4092, N4079, N2288);
nor NOR2 (N4093, N4056, N3017);
xor XOR2 (N4094, N4074, N997);
or OR4 (N4095, N4093, N248, N213, N2755);
not NOT1 (N4096, N4086);
buf BUF1 (N4097, N4092);
xor XOR2 (N4098, N4087, N334);
buf BUF1 (N4099, N4097);
xor XOR2 (N4100, N4095, N559);
not NOT1 (N4101, N4098);
nand NAND4 (N4102, N4080, N1284, N1431, N2063);
nand NAND3 (N4103, N4099, N3502, N2155);
nand NAND2 (N4104, N4090, N464);
nand NAND3 (N4105, N4091, N3378, N1770);
and AND2 (N4106, N4096, N481);
or OR4 (N4107, N4078, N473, N2537, N908);
or OR3 (N4108, N4107, N3959, N1435);
buf BUF1 (N4109, N4105);
and AND3 (N4110, N4109, N3511, N3669);
xor XOR2 (N4111, N4075, N3064);
xor XOR2 (N4112, N4100, N1779);
nor NOR3 (N4113, N4101, N2770, N967);
and AND3 (N4114, N4110, N2553, N931);
xor XOR2 (N4115, N4103, N1387);
and AND2 (N4116, N4112, N470);
or OR2 (N4117, N4108, N2497);
nand NAND4 (N4118, N4116, N3247, N3447, N1845);
or OR2 (N4119, N4094, N4115);
buf BUF1 (N4120, N2886);
nor NOR2 (N4121, N4120, N1923);
nor NOR2 (N4122, N4113, N468);
and AND2 (N4123, N4118, N1302);
and AND4 (N4124, N4104, N3806, N569, N3323);
nand NAND4 (N4125, N4114, N726, N2266, N202);
xor XOR2 (N4126, N4106, N1804);
nand NAND2 (N4127, N4102, N340);
nor NOR3 (N4128, N4127, N879, N1284);
nand NAND4 (N4129, N4124, N531, N1890, N3307);
not NOT1 (N4130, N4125);
nor NOR3 (N4131, N4111, N1404, N1268);
buf BUF1 (N4132, N4122);
xor XOR2 (N4133, N4119, N2889);
xor XOR2 (N4134, N4128, N2154);
xor XOR2 (N4135, N4117, N3748);
and AND2 (N4136, N4135, N4103);
nand NAND4 (N4137, N4130, N3128, N148, N2801);
xor XOR2 (N4138, N4137, N3515);
buf BUF1 (N4139, N4121);
nand NAND3 (N4140, N4131, N3771, N1027);
xor XOR2 (N4141, N4123, N2894);
and AND4 (N4142, N4134, N3188, N2483, N2520);
not NOT1 (N4143, N4140);
buf BUF1 (N4144, N4126);
or OR2 (N4145, N4132, N3939);
buf BUF1 (N4146, N4141);
nand NAND2 (N4147, N4144, N2921);
not NOT1 (N4148, N4147);
or OR2 (N4149, N4145, N1891);
nor NOR3 (N4150, N4148, N23, N1586);
and AND3 (N4151, N4139, N1717, N2902);
nor NOR2 (N4152, N4150, N3424);
or OR3 (N4153, N4146, N1072, N3417);
not NOT1 (N4154, N4138);
not NOT1 (N4155, N4129);
not NOT1 (N4156, N4142);
xor XOR2 (N4157, N4154, N1325);
and AND3 (N4158, N4133, N3747, N2410);
nor NOR4 (N4159, N4152, N3366, N430, N2391);
xor XOR2 (N4160, N4151, N138);
xor XOR2 (N4161, N4160, N3276);
not NOT1 (N4162, N4157);
nor NOR2 (N4163, N4159, N1232);
buf BUF1 (N4164, N4143);
or OR3 (N4165, N4153, N707, N3810);
not NOT1 (N4166, N4158);
nand NAND4 (N4167, N4162, N475, N3834, N3344);
buf BUF1 (N4168, N4167);
buf BUF1 (N4169, N4164);
not NOT1 (N4170, N4169);
nand NAND2 (N4171, N4155, N1566);
nand NAND3 (N4172, N4149, N830, N3398);
nor NOR3 (N4173, N4168, N3276, N2063);
nand NAND4 (N4174, N4170, N2871, N3472, N3785);
buf BUF1 (N4175, N4161);
or OR3 (N4176, N4165, N458, N24);
nor NOR4 (N4177, N4172, N666, N3547, N1725);
nand NAND3 (N4178, N4166, N1958, N1547);
nand NAND2 (N4179, N4174, N72);
buf BUF1 (N4180, N4177);
buf BUF1 (N4181, N4179);
xor XOR2 (N4182, N4163, N235);
buf BUF1 (N4183, N4171);
nand NAND2 (N4184, N4175, N2816);
and AND2 (N4185, N4183, N3738);
and AND3 (N4186, N4178, N2646, N3017);
nor NOR4 (N4187, N4180, N404, N1517, N3442);
xor XOR2 (N4188, N4181, N2234);
nand NAND3 (N4189, N4173, N1582, N2914);
buf BUF1 (N4190, N4176);
or OR4 (N4191, N4136, N2143, N3377, N2052);
not NOT1 (N4192, N4185);
not NOT1 (N4193, N4189);
xor XOR2 (N4194, N4190, N3804);
nand NAND3 (N4195, N4188, N1101, N2789);
and AND4 (N4196, N4187, N476, N2662, N1068);
xor XOR2 (N4197, N4195, N1259);
buf BUF1 (N4198, N4196);
not NOT1 (N4199, N4197);
nand NAND4 (N4200, N4194, N726, N813, N1403);
buf BUF1 (N4201, N4186);
or OR3 (N4202, N4198, N3748, N896);
buf BUF1 (N4203, N4156);
xor XOR2 (N4204, N4202, N1905);
nor NOR3 (N4205, N4193, N787, N716);
and AND2 (N4206, N4192, N3537);
buf BUF1 (N4207, N4205);
xor XOR2 (N4208, N4203, N684);
nor NOR4 (N4209, N4191, N2565, N668, N989);
nand NAND2 (N4210, N4184, N635);
and AND4 (N4211, N4210, N4069, N3234, N3093);
xor XOR2 (N4212, N4211, N415);
or OR4 (N4213, N4206, N1980, N1955, N3180);
xor XOR2 (N4214, N4213, N3008);
nand NAND4 (N4215, N4200, N1471, N3995, N444);
xor XOR2 (N4216, N4207, N1207);
buf BUF1 (N4217, N4212);
not NOT1 (N4218, N4214);
nand NAND3 (N4219, N4217, N1361, N1518);
nor NOR3 (N4220, N4208, N2565, N2100);
nor NOR3 (N4221, N4201, N2077, N2531);
buf BUF1 (N4222, N4221);
buf BUF1 (N4223, N4219);
nand NAND3 (N4224, N4222, N1622, N3149);
nor NOR2 (N4225, N4215, N24);
buf BUF1 (N4226, N4182);
nand NAND2 (N4227, N4204, N4190);
nor NOR2 (N4228, N4216, N2984);
nand NAND3 (N4229, N4218, N4220, N3330);
nor NOR3 (N4230, N2334, N3800, N1079);
buf BUF1 (N4231, N4229);
xor XOR2 (N4232, N4227, N542);
nor NOR4 (N4233, N4225, N2065, N2186, N1160);
nor NOR3 (N4234, N4199, N4087, N4061);
xor XOR2 (N4235, N4226, N2386);
and AND3 (N4236, N4209, N3435, N205);
or OR3 (N4237, N4224, N2806, N1671);
nor NOR4 (N4238, N4231, N2542, N3297, N3674);
buf BUF1 (N4239, N4233);
or OR4 (N4240, N4239, N1601, N1638, N3771);
not NOT1 (N4241, N4234);
xor XOR2 (N4242, N4232, N4120);
buf BUF1 (N4243, N4241);
and AND4 (N4244, N4236, N3582, N1763, N3224);
or OR3 (N4245, N4242, N1231, N4208);
or OR2 (N4246, N4240, N2257);
nor NOR4 (N4247, N4230, N1570, N2763, N1783);
nor NOR3 (N4248, N4247, N1548, N1063);
nand NAND3 (N4249, N4223, N2569, N3821);
xor XOR2 (N4250, N4243, N748);
or OR2 (N4251, N4238, N2421);
nor NOR2 (N4252, N4249, N3338);
or OR2 (N4253, N4235, N1991);
xor XOR2 (N4254, N4246, N3192);
or OR4 (N4255, N4251, N2098, N1111, N158);
and AND4 (N4256, N4248, N2755, N2094, N1757);
buf BUF1 (N4257, N4252);
nand NAND4 (N4258, N4256, N1483, N3837, N710);
buf BUF1 (N4259, N4254);
xor XOR2 (N4260, N4255, N403);
nand NAND3 (N4261, N4258, N3844, N719);
nor NOR4 (N4262, N4245, N1639, N1362, N254);
nor NOR3 (N4263, N4250, N810, N1675);
xor XOR2 (N4264, N4244, N1647);
buf BUF1 (N4265, N4259);
buf BUF1 (N4266, N4265);
or OR2 (N4267, N4260, N2779);
not NOT1 (N4268, N4264);
and AND4 (N4269, N4268, N325, N2442, N607);
xor XOR2 (N4270, N4262, N366);
xor XOR2 (N4271, N4263, N1009);
or OR3 (N4272, N4228, N2929, N2248);
not NOT1 (N4273, N4237);
nor NOR4 (N4274, N4253, N2937, N3547, N1365);
xor XOR2 (N4275, N4274, N3967);
not NOT1 (N4276, N4273);
or OR2 (N4277, N4257, N1625);
xor XOR2 (N4278, N4270, N3072);
or OR2 (N4279, N4277, N1777);
xor XOR2 (N4280, N4278, N1051);
nand NAND4 (N4281, N4279, N1276, N2054, N223);
nor NOR2 (N4282, N4280, N3817);
nor NOR2 (N4283, N4282, N1362);
and AND3 (N4284, N4281, N789, N4257);
not NOT1 (N4285, N4271);
xor XOR2 (N4286, N4275, N3536);
nor NOR4 (N4287, N4276, N1423, N1149, N1517);
nand NAND2 (N4288, N4287, N3211);
or OR3 (N4289, N4283, N1824, N1320);
xor XOR2 (N4290, N4269, N2978);
nor NOR3 (N4291, N4288, N3843, N424);
nand NAND2 (N4292, N4286, N2926);
xor XOR2 (N4293, N4266, N1580);
nand NAND2 (N4294, N4261, N2917);
nand NAND3 (N4295, N4292, N2449, N4265);
nor NOR3 (N4296, N4289, N1519, N3397);
buf BUF1 (N4297, N4284);
nand NAND4 (N4298, N4296, N1905, N1238, N3663);
not NOT1 (N4299, N4298);
and AND3 (N4300, N4295, N1808, N2456);
xor XOR2 (N4301, N4293, N846);
not NOT1 (N4302, N4294);
xor XOR2 (N4303, N4299, N223);
and AND2 (N4304, N4290, N424);
not NOT1 (N4305, N4272);
buf BUF1 (N4306, N4304);
not NOT1 (N4307, N4305);
nor NOR4 (N4308, N4306, N3732, N1193, N1959);
buf BUF1 (N4309, N4308);
and AND4 (N4310, N4307, N4281, N1957, N1696);
xor XOR2 (N4311, N4267, N3401);
and AND2 (N4312, N4302, N736);
or OR4 (N4313, N4301, N224, N3335, N3373);
or OR2 (N4314, N4300, N2814);
nor NOR3 (N4315, N4297, N308, N4234);
xor XOR2 (N4316, N4309, N128);
nand NAND2 (N4317, N4311, N4080);
buf BUF1 (N4318, N4314);
xor XOR2 (N4319, N4317, N849);
xor XOR2 (N4320, N4312, N1583);
or OR2 (N4321, N4291, N1801);
or OR4 (N4322, N4310, N1410, N2176, N3757);
buf BUF1 (N4323, N4285);
xor XOR2 (N4324, N4316, N4114);
or OR4 (N4325, N4313, N2978, N1328, N1758);
nor NOR2 (N4326, N4325, N3481);
not NOT1 (N4327, N4320);
buf BUF1 (N4328, N4326);
nor NOR2 (N4329, N4319, N1576);
not NOT1 (N4330, N4315);
or OR4 (N4331, N4323, N2845, N2884, N919);
nand NAND2 (N4332, N4328, N332);
not NOT1 (N4333, N4329);
not NOT1 (N4334, N4333);
and AND2 (N4335, N4331, N2875);
not NOT1 (N4336, N4322);
not NOT1 (N4337, N4334);
and AND2 (N4338, N4327, N281);
buf BUF1 (N4339, N4336);
xor XOR2 (N4340, N4321, N1124);
nand NAND4 (N4341, N4337, N417, N614, N4176);
not NOT1 (N4342, N4341);
nor NOR2 (N4343, N4339, N2876);
nor NOR4 (N4344, N4318, N3475, N3839, N3783);
not NOT1 (N4345, N4330);
or OR4 (N4346, N4343, N4071, N4087, N2926);
or OR4 (N4347, N4345, N1543, N2860, N2720);
buf BUF1 (N4348, N4346);
nand NAND3 (N4349, N4347, N838, N116);
nand NAND2 (N4350, N4332, N4054);
and AND2 (N4351, N4335, N2153);
or OR2 (N4352, N4340, N1731);
nand NAND4 (N4353, N4350, N1031, N3390, N951);
not NOT1 (N4354, N4353);
or OR3 (N4355, N4324, N451, N4262);
nor NOR3 (N4356, N4348, N2019, N2499);
nand NAND4 (N4357, N4342, N2898, N3551, N1929);
not NOT1 (N4358, N4357);
nand NAND4 (N4359, N4356, N3085, N784, N1013);
not NOT1 (N4360, N4359);
xor XOR2 (N4361, N4358, N3724);
and AND4 (N4362, N4303, N1312, N2247, N4285);
not NOT1 (N4363, N4354);
nor NOR2 (N4364, N4362, N3055);
and AND3 (N4365, N4355, N1434, N157);
and AND4 (N4366, N4344, N832, N2375, N4314);
buf BUF1 (N4367, N4363);
not NOT1 (N4368, N4364);
not NOT1 (N4369, N4361);
buf BUF1 (N4370, N4367);
xor XOR2 (N4371, N4366, N1755);
buf BUF1 (N4372, N4365);
or OR2 (N4373, N4338, N4196);
xor XOR2 (N4374, N4349, N3149);
or OR4 (N4375, N4374, N4199, N393, N4080);
xor XOR2 (N4376, N4369, N2399);
or OR4 (N4377, N4351, N1979, N1233, N111);
nand NAND4 (N4378, N4377, N150, N2750, N465);
nor NOR4 (N4379, N4376, N1536, N1806, N285);
and AND3 (N4380, N4360, N1533, N2298);
and AND2 (N4381, N4380, N1496);
or OR3 (N4382, N4379, N3378, N3352);
or OR3 (N4383, N4352, N3638, N3355);
nor NOR3 (N4384, N4375, N1555, N2948);
nor NOR3 (N4385, N4373, N2056, N1770);
xor XOR2 (N4386, N4381, N3498);
buf BUF1 (N4387, N4378);
or OR2 (N4388, N4372, N1299);
and AND3 (N4389, N4386, N3093, N696);
xor XOR2 (N4390, N4382, N2907);
or OR2 (N4391, N4370, N667);
or OR3 (N4392, N4385, N683, N1697);
buf BUF1 (N4393, N4390);
and AND4 (N4394, N4389, N1985, N1249, N547);
xor XOR2 (N4395, N4392, N1598);
nand NAND4 (N4396, N4383, N2153, N4058, N4178);
nor NOR4 (N4397, N4368, N3899, N325, N3351);
nand NAND2 (N4398, N4395, N151);
xor XOR2 (N4399, N4398, N62);
and AND3 (N4400, N4387, N1216, N2758);
nand NAND2 (N4401, N4396, N486);
nand NAND4 (N4402, N4391, N1231, N1112, N3295);
nand NAND2 (N4403, N4388, N2331);
buf BUF1 (N4404, N4397);
not NOT1 (N4405, N4384);
buf BUF1 (N4406, N4371);
xor XOR2 (N4407, N4406, N3375);
nand NAND3 (N4408, N4401, N3646, N3289);
or OR3 (N4409, N4399, N1698, N4112);
nor NOR4 (N4410, N4408, N56, N437, N3048);
not NOT1 (N4411, N4409);
buf BUF1 (N4412, N4410);
or OR2 (N4413, N4393, N3774);
nor NOR4 (N4414, N4412, N2005, N317, N1749);
not NOT1 (N4415, N4400);
not NOT1 (N4416, N4405);
nand NAND3 (N4417, N4416, N2035, N2900);
nor NOR4 (N4418, N4415, N3563, N485, N2971);
nor NOR2 (N4419, N4407, N369);
or OR3 (N4420, N4417, N3577, N848);
xor XOR2 (N4421, N4413, N4330);
and AND3 (N4422, N4414, N2357, N4058);
and AND3 (N4423, N4402, N4132, N516);
and AND2 (N4424, N4394, N2284);
xor XOR2 (N4425, N4411, N1589);
and AND2 (N4426, N4403, N3327);
and AND4 (N4427, N4418, N579, N1372, N55);
nor NOR2 (N4428, N4425, N3347);
not NOT1 (N4429, N4427);
and AND3 (N4430, N4429, N1493, N2318);
not NOT1 (N4431, N4419);
not NOT1 (N4432, N4428);
nand NAND4 (N4433, N4420, N1346, N1234, N929);
buf BUF1 (N4434, N4404);
or OR3 (N4435, N4434, N670, N2685);
buf BUF1 (N4436, N4435);
buf BUF1 (N4437, N4426);
xor XOR2 (N4438, N4431, N4050);
or OR4 (N4439, N4422, N1920, N560, N1349);
and AND4 (N4440, N4430, N3521, N1670, N1594);
xor XOR2 (N4441, N4437, N2701);
nor NOR3 (N4442, N4432, N3753, N3113);
or OR4 (N4443, N4423, N2759, N103, N2572);
and AND2 (N4444, N4438, N1051);
buf BUF1 (N4445, N4444);
xor XOR2 (N4446, N4442, N3832);
not NOT1 (N4447, N4446);
nor NOR3 (N4448, N4424, N2181, N2972);
and AND4 (N4449, N4436, N1043, N525, N1974);
or OR4 (N4450, N4443, N1587, N737, N3425);
buf BUF1 (N4451, N4449);
and AND3 (N4452, N4445, N675, N3207);
xor XOR2 (N4453, N4439, N2347);
nand NAND3 (N4454, N4453, N1793, N2566);
xor XOR2 (N4455, N4440, N3977);
buf BUF1 (N4456, N4455);
not NOT1 (N4457, N4441);
nor NOR4 (N4458, N4450, N3549, N3766, N1128);
xor XOR2 (N4459, N4448, N4366);
xor XOR2 (N4460, N4421, N3467);
nand NAND4 (N4461, N4447, N2762, N1411, N1491);
or OR2 (N4462, N4451, N1529);
nor NOR3 (N4463, N4458, N4143, N193);
nor NOR3 (N4464, N4457, N1505, N3225);
or OR3 (N4465, N4433, N3610, N1470);
or OR4 (N4466, N4465, N944, N943, N1123);
and AND2 (N4467, N4462, N1468);
not NOT1 (N4468, N4459);
nor NOR4 (N4469, N4466, N3202, N4326, N3042);
xor XOR2 (N4470, N4469, N1122);
xor XOR2 (N4471, N4454, N3454);
and AND4 (N4472, N4471, N3336, N3721, N4383);
buf BUF1 (N4473, N4472);
nand NAND4 (N4474, N4460, N338, N60, N417);
nor NOR2 (N4475, N4464, N121);
xor XOR2 (N4476, N4474, N1666);
not NOT1 (N4477, N4475);
and AND4 (N4478, N4473, N3869, N1671, N2010);
nand NAND4 (N4479, N4456, N4247, N3152, N3547);
xor XOR2 (N4480, N4468, N129);
buf BUF1 (N4481, N4478);
and AND2 (N4482, N4452, N3452);
nor NOR2 (N4483, N4470, N4087);
xor XOR2 (N4484, N4463, N1364);
or OR3 (N4485, N4477, N3020, N3825);
not NOT1 (N4486, N4485);
not NOT1 (N4487, N4481);
xor XOR2 (N4488, N4484, N1328);
or OR2 (N4489, N4487, N2560);
buf BUF1 (N4490, N4461);
xor XOR2 (N4491, N4467, N1752);
not NOT1 (N4492, N4489);
nand NAND4 (N4493, N4476, N3888, N1865, N1358);
xor XOR2 (N4494, N4486, N1145);
nor NOR4 (N4495, N4491, N3469, N254, N1195);
nand NAND4 (N4496, N4482, N1283, N2, N3994);
buf BUF1 (N4497, N4492);
not NOT1 (N4498, N4497);
buf BUF1 (N4499, N4493);
and AND4 (N4500, N4494, N168, N27, N4023);
buf BUF1 (N4501, N4496);
and AND3 (N4502, N4500, N1731, N2990);
nand NAND3 (N4503, N4479, N1337, N2266);
or OR2 (N4504, N4483, N3698);
nand NAND2 (N4505, N4504, N2746);
nand NAND4 (N4506, N4501, N1259, N2831, N1651);
or OR4 (N4507, N4480, N1001, N3862, N1160);
buf BUF1 (N4508, N4506);
and AND2 (N4509, N4495, N3770);
nor NOR4 (N4510, N4499, N2559, N2716, N950);
or OR2 (N4511, N4508, N4015);
nor NOR3 (N4512, N4510, N3468, N3550);
buf BUF1 (N4513, N4490);
and AND4 (N4514, N4488, N127, N325, N991);
and AND3 (N4515, N4505, N1243, N2888);
nand NAND2 (N4516, N4513, N694);
not NOT1 (N4517, N4498);
nor NOR4 (N4518, N4509, N3334, N4151, N73);
and AND4 (N4519, N4517, N3833, N2211, N3035);
buf BUF1 (N4520, N4518);
nor NOR4 (N4521, N4515, N701, N1638, N577);
nor NOR4 (N4522, N4519, N2609, N3135, N1820);
buf BUF1 (N4523, N4516);
buf BUF1 (N4524, N4522);
not NOT1 (N4525, N4523);
nand NAND3 (N4526, N4502, N1929, N1699);
not NOT1 (N4527, N4524);
or OR3 (N4528, N4521, N398, N3535);
not NOT1 (N4529, N4514);
and AND2 (N4530, N4507, N2754);
and AND2 (N4531, N4526, N347);
nor NOR3 (N4532, N4531, N484, N1523);
not NOT1 (N4533, N4520);
nand NAND4 (N4534, N4528, N1770, N783, N1250);
nand NAND3 (N4535, N4529, N3384, N1088);
not NOT1 (N4536, N4512);
xor XOR2 (N4537, N4533, N824);
buf BUF1 (N4538, N4536);
nand NAND4 (N4539, N4511, N3936, N3377, N171);
and AND4 (N4540, N4503, N1363, N2179, N4041);
xor XOR2 (N4541, N4539, N1440);
buf BUF1 (N4542, N4535);
nand NAND3 (N4543, N4532, N3104, N2592);
xor XOR2 (N4544, N4530, N613);
buf BUF1 (N4545, N4543);
buf BUF1 (N4546, N4538);
or OR4 (N4547, N4534, N167, N104, N2977);
or OR4 (N4548, N4541, N1717, N2766, N1902);
xor XOR2 (N4549, N4545, N1842);
not NOT1 (N4550, N4544);
buf BUF1 (N4551, N4527);
and AND3 (N4552, N4525, N2836, N1025);
nor NOR3 (N4553, N4549, N4533, N1525);
nand NAND4 (N4554, N4550, N3353, N4352, N4384);
buf BUF1 (N4555, N4553);
xor XOR2 (N4556, N4551, N2235);
nand NAND4 (N4557, N4537, N1174, N2482, N891);
or OR3 (N4558, N4540, N861, N350);
xor XOR2 (N4559, N4542, N505);
nor NOR2 (N4560, N4554, N1701);
not NOT1 (N4561, N4556);
and AND4 (N4562, N4546, N662, N231, N1339);
buf BUF1 (N4563, N4555);
nor NOR2 (N4564, N4548, N3217);
not NOT1 (N4565, N4547);
xor XOR2 (N4566, N4565, N921);
buf BUF1 (N4567, N4562);
nor NOR4 (N4568, N4558, N1986, N950, N2037);
and AND2 (N4569, N4566, N2664);
not NOT1 (N4570, N4567);
or OR4 (N4571, N4564, N217, N4239, N3662);
not NOT1 (N4572, N4559);
not NOT1 (N4573, N4570);
nor NOR3 (N4574, N4569, N4063, N3566);
nor NOR3 (N4575, N4572, N3386, N2306);
xor XOR2 (N4576, N4560, N3596);
or OR2 (N4577, N4557, N2626);
or OR3 (N4578, N4571, N3173, N151);
and AND3 (N4579, N4575, N2171, N1365);
xor XOR2 (N4580, N4579, N1251);
and AND3 (N4581, N4574, N2637, N2916);
xor XOR2 (N4582, N4552, N501);
buf BUF1 (N4583, N4563);
buf BUF1 (N4584, N4568);
not NOT1 (N4585, N4584);
or OR2 (N4586, N4580, N4261);
not NOT1 (N4587, N4576);
and AND4 (N4588, N4578, N4433, N2864, N2159);
not NOT1 (N4589, N4573);
nor NOR3 (N4590, N4561, N2374, N126);
not NOT1 (N4591, N4581);
buf BUF1 (N4592, N4586);
or OR4 (N4593, N4590, N4425, N3943, N4112);
buf BUF1 (N4594, N4591);
or OR3 (N4595, N4585, N1280, N1048);
nor NOR4 (N4596, N4589, N1166, N4307, N2765);
and AND4 (N4597, N4583, N3220, N2895, N3326);
or OR2 (N4598, N4587, N507);
not NOT1 (N4599, N4597);
and AND3 (N4600, N4595, N3616, N1318);
buf BUF1 (N4601, N4594);
nand NAND3 (N4602, N4577, N4592, N4245);
and AND2 (N4603, N425, N1549);
xor XOR2 (N4604, N4596, N3218);
or OR4 (N4605, N4601, N3422, N3010, N182);
and AND4 (N4606, N4602, N2004, N1747, N1563);
xor XOR2 (N4607, N4606, N1171);
and AND2 (N4608, N4603, N2547);
buf BUF1 (N4609, N4588);
and AND2 (N4610, N4582, N857);
xor XOR2 (N4611, N4609, N2055);
and AND4 (N4612, N4599, N3378, N3763, N4538);
xor XOR2 (N4613, N4598, N3791);
not NOT1 (N4614, N4610);
and AND4 (N4615, N4613, N3332, N718, N2420);
nand NAND4 (N4616, N4614, N4613, N2388, N1151);
buf BUF1 (N4617, N4593);
not NOT1 (N4618, N4611);
not NOT1 (N4619, N4608);
nor NOR3 (N4620, N4615, N677, N1338);
xor XOR2 (N4621, N4607, N1953);
not NOT1 (N4622, N4618);
or OR3 (N4623, N4620, N2109, N3006);
or OR4 (N4624, N4619, N2357, N1272, N492);
nand NAND4 (N4625, N4623, N4537, N2310, N3539);
not NOT1 (N4626, N4625);
not NOT1 (N4627, N4600);
buf BUF1 (N4628, N4624);
not NOT1 (N4629, N4627);
nand NAND4 (N4630, N4612, N3556, N2073, N2315);
nor NOR4 (N4631, N4628, N4410, N399, N3982);
and AND4 (N4632, N4605, N3166, N828, N2998);
not NOT1 (N4633, N4617);
and AND3 (N4634, N4622, N4326, N1679);
xor XOR2 (N4635, N4630, N869);
nor NOR2 (N4636, N4631, N2303);
or OR3 (N4637, N4632, N3033, N2236);
nor NOR4 (N4638, N4637, N4183, N3728, N602);
not NOT1 (N4639, N4638);
nand NAND2 (N4640, N4604, N888);
or OR3 (N4641, N4634, N1049, N4318);
buf BUF1 (N4642, N4633);
xor XOR2 (N4643, N4616, N1256);
or OR3 (N4644, N4642, N3305, N1289);
nor NOR4 (N4645, N4635, N2689, N341, N3420);
not NOT1 (N4646, N4640);
nand NAND4 (N4647, N4644, N152, N358, N567);
nor NOR4 (N4648, N4639, N1276, N2054, N2154);
or OR3 (N4649, N4647, N1057, N4041);
not NOT1 (N4650, N4648);
buf BUF1 (N4651, N4650);
buf BUF1 (N4652, N4641);
buf BUF1 (N4653, N4646);
buf BUF1 (N4654, N4621);
nand NAND4 (N4655, N4626, N2743, N4040, N4013);
xor XOR2 (N4656, N4655, N874);
nor NOR3 (N4657, N4656, N54, N1745);
or OR2 (N4658, N4643, N3191);
xor XOR2 (N4659, N4636, N24);
nand NAND2 (N4660, N4653, N2400);
nor NOR3 (N4661, N4658, N2131, N550);
nand NAND2 (N4662, N4661, N3318);
or OR4 (N4663, N4651, N4364, N4186, N802);
and AND2 (N4664, N4657, N3796);
buf BUF1 (N4665, N4652);
or OR4 (N4666, N4659, N2762, N3631, N3781);
nand NAND4 (N4667, N4662, N3165, N2635, N3812);
and AND3 (N4668, N4667, N2946, N290);
or OR2 (N4669, N4664, N419);
or OR3 (N4670, N4660, N1892, N3873);
not NOT1 (N4671, N4629);
xor XOR2 (N4672, N4668, N1809);
buf BUF1 (N4673, N4666);
or OR2 (N4674, N4671, N657);
not NOT1 (N4675, N4672);
not NOT1 (N4676, N4649);
buf BUF1 (N4677, N4663);
not NOT1 (N4678, N4676);
buf BUF1 (N4679, N4669);
xor XOR2 (N4680, N4673, N2177);
not NOT1 (N4681, N4675);
not NOT1 (N4682, N4678);
nand NAND3 (N4683, N4654, N4615, N1426);
nand NAND4 (N4684, N4674, N2543, N2183, N797);
nor NOR3 (N4685, N4680, N1598, N3107);
xor XOR2 (N4686, N4677, N3772);
and AND2 (N4687, N4685, N547);
buf BUF1 (N4688, N4684);
not NOT1 (N4689, N4665);
buf BUF1 (N4690, N4686);
and AND2 (N4691, N4690, N181);
xor XOR2 (N4692, N4688, N2595);
nand NAND4 (N4693, N4687, N1384, N2787, N1446);
nor NOR4 (N4694, N4682, N4476, N668, N1740);
and AND3 (N4695, N4692, N4299, N1168);
not NOT1 (N4696, N4670);
buf BUF1 (N4697, N4695);
xor XOR2 (N4698, N4679, N3669);
or OR4 (N4699, N4693, N3269, N2830, N40);
xor XOR2 (N4700, N4681, N4069);
and AND2 (N4701, N4689, N4308);
xor XOR2 (N4702, N4694, N805);
or OR4 (N4703, N4699, N868, N4477, N4198);
buf BUF1 (N4704, N4697);
not NOT1 (N4705, N4683);
nand NAND3 (N4706, N4645, N954, N1754);
buf BUF1 (N4707, N4703);
nand NAND2 (N4708, N4701, N3302);
nand NAND2 (N4709, N4707, N4337);
not NOT1 (N4710, N4705);
or OR4 (N4711, N4710, N1120, N4319, N1783);
xor XOR2 (N4712, N4691, N3435);
nand NAND2 (N4713, N4702, N1294);
or OR3 (N4714, N4700, N4239, N1606);
xor XOR2 (N4715, N4711, N3668);
nor NOR3 (N4716, N4704, N3063, N4461);
buf BUF1 (N4717, N4716);
nor NOR4 (N4718, N4706, N3399, N1844, N2588);
or OR4 (N4719, N4715, N3856, N2244, N1926);
xor XOR2 (N4720, N4714, N2728);
buf BUF1 (N4721, N4712);
nor NOR2 (N4722, N4709, N4298);
or OR3 (N4723, N4720, N3963, N3551);
buf BUF1 (N4724, N4722);
nand NAND4 (N4725, N4708, N217, N3753, N1563);
or OR2 (N4726, N4696, N4167);
buf BUF1 (N4727, N4723);
or OR3 (N4728, N4698, N2356, N3932);
and AND4 (N4729, N4713, N4594, N2167, N115);
nor NOR4 (N4730, N4721, N4665, N666, N4679);
or OR4 (N4731, N4725, N1429, N2308, N737);
or OR3 (N4732, N4727, N859, N2354);
nor NOR4 (N4733, N4724, N958, N3649, N2828);
or OR3 (N4734, N4728, N4510, N374);
xor XOR2 (N4735, N4730, N2023);
xor XOR2 (N4736, N4729, N3231);
buf BUF1 (N4737, N4726);
or OR4 (N4738, N4736, N3041, N14, N4130);
nand NAND2 (N4739, N4737, N1433);
nor NOR2 (N4740, N4731, N4619);
or OR4 (N4741, N4739, N2130, N3855, N4350);
and AND4 (N4742, N4717, N1539, N231, N215);
nand NAND2 (N4743, N4742, N1393);
not NOT1 (N4744, N4738);
or OR2 (N4745, N4743, N2621);
buf BUF1 (N4746, N4733);
buf BUF1 (N4747, N4719);
or OR2 (N4748, N4745, N765);
buf BUF1 (N4749, N4732);
nor NOR3 (N4750, N4735, N2913, N443);
nand NAND2 (N4751, N4749, N3470);
xor XOR2 (N4752, N4740, N1464);
nand NAND2 (N4753, N4746, N3992);
not NOT1 (N4754, N4751);
and AND3 (N4755, N4748, N2544, N2473);
and AND4 (N4756, N4750, N996, N3173, N4171);
and AND3 (N4757, N4756, N1298, N1224);
not NOT1 (N4758, N4747);
buf BUF1 (N4759, N4752);
and AND2 (N4760, N4718, N4031);
not NOT1 (N4761, N4755);
and AND2 (N4762, N4759, N76);
not NOT1 (N4763, N4734);
nand NAND3 (N4764, N4762, N379, N576);
buf BUF1 (N4765, N4753);
nor NOR4 (N4766, N4765, N3095, N4454, N2450);
nor NOR4 (N4767, N4764, N3888, N1766, N1866);
or OR3 (N4768, N4757, N2093, N4074);
and AND4 (N4769, N4754, N857, N2274, N4332);
nor NOR4 (N4770, N4758, N4536, N3588, N639);
nor NOR2 (N4771, N4770, N3494);
nand NAND3 (N4772, N4771, N416, N2848);
buf BUF1 (N4773, N4767);
and AND4 (N4774, N4766, N974, N988, N2848);
and AND4 (N4775, N4768, N3834, N1991, N982);
not NOT1 (N4776, N4769);
nand NAND4 (N4777, N4741, N3962, N1072, N136);
nor NOR2 (N4778, N4760, N418);
or OR3 (N4779, N4773, N4532, N27);
nand NAND2 (N4780, N4774, N1339);
not NOT1 (N4781, N4780);
xor XOR2 (N4782, N4776, N1170);
nor NOR3 (N4783, N4781, N4150, N1224);
not NOT1 (N4784, N4761);
nand NAND3 (N4785, N4778, N1408, N472);
nand NAND3 (N4786, N4775, N4536, N1511);
buf BUF1 (N4787, N4779);
nor NOR3 (N4788, N4782, N1471, N2548);
or OR3 (N4789, N4744, N603, N4060);
or OR2 (N4790, N4777, N4163);
xor XOR2 (N4791, N4788, N1218);
buf BUF1 (N4792, N4790);
nor NOR3 (N4793, N4783, N4676, N396);
nand NAND2 (N4794, N4772, N3950);
buf BUF1 (N4795, N4789);
not NOT1 (N4796, N4795);
not NOT1 (N4797, N4792);
and AND3 (N4798, N4763, N3390, N1019);
xor XOR2 (N4799, N4784, N2496);
buf BUF1 (N4800, N4786);
not NOT1 (N4801, N4800);
nor NOR2 (N4802, N4801, N1863);
not NOT1 (N4803, N4791);
and AND2 (N4804, N4793, N2361);
and AND2 (N4805, N4796, N3027);
xor XOR2 (N4806, N4804, N2307);
and AND2 (N4807, N4798, N734);
and AND2 (N4808, N4807, N4709);
nor NOR4 (N4809, N4787, N3787, N4485, N2839);
nand NAND3 (N4810, N4809, N1142, N4182);
xor XOR2 (N4811, N4805, N1848);
buf BUF1 (N4812, N4797);
buf BUF1 (N4813, N4785);
xor XOR2 (N4814, N4802, N3818);
buf BUF1 (N4815, N4803);
buf BUF1 (N4816, N4810);
nand NAND2 (N4817, N4794, N408);
xor XOR2 (N4818, N4812, N4445);
or OR2 (N4819, N4815, N2459);
xor XOR2 (N4820, N4817, N4323);
buf BUF1 (N4821, N4811);
nand NAND3 (N4822, N4820, N4076, N2133);
not NOT1 (N4823, N4814);
and AND3 (N4824, N4818, N4752, N1694);
not NOT1 (N4825, N4806);
not NOT1 (N4826, N4813);
not NOT1 (N4827, N4808);
and AND3 (N4828, N4821, N1015, N1002);
nand NAND3 (N4829, N4819, N89, N2157);
buf BUF1 (N4830, N4822);
or OR3 (N4831, N4816, N3181, N2486);
nor NOR2 (N4832, N4830, N2651);
or OR4 (N4833, N4832, N296, N3680, N133);
xor XOR2 (N4834, N4828, N83);
or OR3 (N4835, N4824, N1054, N1010);
not NOT1 (N4836, N4835);
nand NAND3 (N4837, N4834, N894, N3875);
xor XOR2 (N4838, N4833, N323);
buf BUF1 (N4839, N4823);
or OR4 (N4840, N4826, N2099, N72, N2858);
nor NOR4 (N4841, N4831, N3133, N4633, N852);
nor NOR4 (N4842, N4837, N4138, N1346, N3084);
not NOT1 (N4843, N4825);
buf BUF1 (N4844, N4799);
buf BUF1 (N4845, N4827);
buf BUF1 (N4846, N4836);
not NOT1 (N4847, N4844);
and AND2 (N4848, N4842, N1873);
or OR3 (N4849, N4840, N97, N2783);
not NOT1 (N4850, N4841);
xor XOR2 (N4851, N4848, N4539);
xor XOR2 (N4852, N4849, N1995);
nand NAND2 (N4853, N4851, N3441);
nor NOR3 (N4854, N4850, N4406, N3532);
and AND4 (N4855, N4852, N4431, N4672, N4735);
nor NOR2 (N4856, N4846, N1071);
or OR2 (N4857, N4839, N1822);
or OR4 (N4858, N4847, N2436, N1317, N4510);
and AND2 (N4859, N4857, N1091);
xor XOR2 (N4860, N4845, N2358);
xor XOR2 (N4861, N4843, N4409);
and AND2 (N4862, N4854, N558);
xor XOR2 (N4863, N4829, N3854);
buf BUF1 (N4864, N4858);
buf BUF1 (N4865, N4864);
xor XOR2 (N4866, N4860, N3428);
nor NOR3 (N4867, N4863, N4650, N3459);
nor NOR4 (N4868, N4856, N2112, N3793, N696);
not NOT1 (N4869, N4861);
nor NOR4 (N4870, N4855, N4654, N1497, N3560);
nor NOR2 (N4871, N4862, N1868);
buf BUF1 (N4872, N4866);
buf BUF1 (N4873, N4871);
not NOT1 (N4874, N4853);
or OR4 (N4875, N4859, N1935, N832, N3620);
not NOT1 (N4876, N4872);
not NOT1 (N4877, N4876);
nor NOR4 (N4878, N4877, N3239, N1109, N2307);
not NOT1 (N4879, N4878);
buf BUF1 (N4880, N4838);
xor XOR2 (N4881, N4865, N2444);
nand NAND2 (N4882, N4875, N4851);
xor XOR2 (N4883, N4869, N3843);
buf BUF1 (N4884, N4881);
not NOT1 (N4885, N4868);
nor NOR3 (N4886, N4874, N989, N3153);
and AND2 (N4887, N4885, N77);
buf BUF1 (N4888, N4873);
and AND4 (N4889, N4870, N61, N4340, N2638);
nor NOR2 (N4890, N4887, N11);
and AND2 (N4891, N4883, N1317);
nand NAND2 (N4892, N4882, N1602);
nand NAND3 (N4893, N4884, N4825, N1797);
xor XOR2 (N4894, N4888, N3300);
and AND2 (N4895, N4890, N796);
buf BUF1 (N4896, N4889);
nor NOR3 (N4897, N4896, N471, N2319);
not NOT1 (N4898, N4867);
buf BUF1 (N4899, N4892);
xor XOR2 (N4900, N4879, N4308);
not NOT1 (N4901, N4880);
xor XOR2 (N4902, N4886, N4450);
nor NOR3 (N4903, N4899, N3420, N2832);
and AND3 (N4904, N4895, N1023, N4267);
or OR4 (N4905, N4893, N3606, N1930, N2820);
nor NOR2 (N4906, N4903, N2601);
nor NOR3 (N4907, N4898, N2188, N3200);
nand NAND4 (N4908, N4907, N1861, N3601, N3842);
nor NOR2 (N4909, N4908, N662);
nor NOR3 (N4910, N4909, N375, N806);
buf BUF1 (N4911, N4901);
or OR3 (N4912, N4897, N4367, N3864);
and AND3 (N4913, N4904, N4181, N4869);
nand NAND4 (N4914, N4911, N643, N1791, N2767);
xor XOR2 (N4915, N4891, N364);
buf BUF1 (N4916, N4914);
nand NAND3 (N4917, N4912, N4189, N3979);
not NOT1 (N4918, N4902);
nor NOR2 (N4919, N4915, N2401);
nand NAND4 (N4920, N4910, N2876, N1549, N1439);
or OR3 (N4921, N4913, N3092, N2393);
and AND4 (N4922, N4920, N744, N2935, N524);
buf BUF1 (N4923, N4916);
nor NOR3 (N4924, N4905, N2998, N1428);
nor NOR4 (N4925, N4900, N2658, N2313, N4629);
xor XOR2 (N4926, N4924, N2115);
nand NAND2 (N4927, N4919, N2375);
nand NAND4 (N4928, N4925, N1640, N1921, N4137);
nand NAND3 (N4929, N4928, N66, N4156);
nand NAND4 (N4930, N4923, N3684, N1739, N3867);
buf BUF1 (N4931, N4929);
nor NOR2 (N4932, N4917, N4696);
nor NOR2 (N4933, N4921, N1103);
nor NOR4 (N4934, N4931, N912, N2920, N3377);
buf BUF1 (N4935, N4918);
nand NAND3 (N4936, N4932, N2654, N3166);
xor XOR2 (N4937, N4935, N4520);
or OR4 (N4938, N4936, N4524, N2135, N1598);
nor NOR3 (N4939, N4933, N67, N2604);
and AND3 (N4940, N4939, N810, N2429);
nand NAND3 (N4941, N4937, N1501, N4097);
not NOT1 (N4942, N4927);
buf BUF1 (N4943, N4942);
xor XOR2 (N4944, N4934, N2725);
buf BUF1 (N4945, N4922);
nor NOR3 (N4946, N4938, N4164, N2034);
xor XOR2 (N4947, N4930, N411);
and AND2 (N4948, N4947, N2665);
xor XOR2 (N4949, N4940, N78);
nor NOR3 (N4950, N4926, N1314, N4052);
buf BUF1 (N4951, N4944);
and AND4 (N4952, N4941, N4211, N3756, N946);
buf BUF1 (N4953, N4948);
nand NAND4 (N4954, N4894, N148, N1173, N3111);
nand NAND4 (N4955, N4950, N3573, N4254, N3527);
nand NAND2 (N4956, N4943, N3862);
or OR3 (N4957, N4949, N603, N1376);
or OR3 (N4958, N4956, N3412, N857);
not NOT1 (N4959, N4946);
and AND4 (N4960, N4954, N408, N4519, N1943);
nor NOR4 (N4961, N4960, N4792, N103, N1288);
or OR3 (N4962, N4953, N2805, N378);
or OR3 (N4963, N4962, N1915, N1924);
xor XOR2 (N4964, N4961, N3285);
not NOT1 (N4965, N4963);
nand NAND3 (N4966, N4965, N1820, N4906);
or OR3 (N4967, N4267, N2444, N622);
xor XOR2 (N4968, N4952, N3214);
nor NOR3 (N4969, N4959, N1008, N1068);
not NOT1 (N4970, N4967);
xor XOR2 (N4971, N4958, N305);
nor NOR3 (N4972, N4951, N746, N2828);
and AND4 (N4973, N4971, N4123, N2411, N2725);
not NOT1 (N4974, N4973);
nand NAND2 (N4975, N4974, N2387);
nand NAND4 (N4976, N4945, N1637, N2735, N676);
nand NAND3 (N4977, N4966, N3248, N4587);
not NOT1 (N4978, N4957);
nor NOR4 (N4979, N4969, N3277, N4660, N4375);
or OR2 (N4980, N4979, N530);
not NOT1 (N4981, N4970);
nand NAND3 (N4982, N4978, N4565, N3570);
not NOT1 (N4983, N4976);
nand NAND3 (N4984, N4980, N4525, N626);
nor NOR3 (N4985, N4955, N989, N1453);
buf BUF1 (N4986, N4984);
and AND4 (N4987, N4986, N4338, N1186, N1823);
buf BUF1 (N4988, N4977);
nor NOR3 (N4989, N4968, N3679, N34);
nand NAND2 (N4990, N4964, N1695);
buf BUF1 (N4991, N4982);
nand NAND3 (N4992, N4989, N402, N1337);
nor NOR4 (N4993, N4987, N194, N2237, N3676);
and AND3 (N4994, N4988, N40, N2086);
buf BUF1 (N4995, N4975);
not NOT1 (N4996, N4983);
or OR3 (N4997, N4991, N3038, N4831);
or OR3 (N4998, N4997, N4616, N3606);
buf BUF1 (N4999, N4990);
not NOT1 (N5000, N4985);
nor NOR4 (N5001, N4993, N2133, N3349, N2905);
and AND4 (N5002, N4981, N76, N1145, N2666);
or OR2 (N5003, N4996, N2759);
or OR2 (N5004, N5002, N2539);
nor NOR2 (N5005, N5001, N1128);
or OR2 (N5006, N4992, N1112);
nor NOR2 (N5007, N5000, N3778);
or OR3 (N5008, N5003, N3038, N3498);
buf BUF1 (N5009, N5006);
and AND4 (N5010, N4998, N1023, N3621, N1981);
or OR3 (N5011, N5004, N4068, N3226);
buf BUF1 (N5012, N4999);
or OR4 (N5013, N5005, N2020, N3317, N3185);
buf BUF1 (N5014, N5009);
buf BUF1 (N5015, N4994);
xor XOR2 (N5016, N5010, N4183);
or OR3 (N5017, N5014, N4155, N456);
nand NAND3 (N5018, N5008, N4905, N4913);
or OR2 (N5019, N5011, N729);
nand NAND2 (N5020, N5012, N3084);
nor NOR4 (N5021, N5007, N3465, N4001, N2438);
and AND4 (N5022, N5019, N313, N2107, N180);
and AND3 (N5023, N5013, N723, N2485);
nor NOR2 (N5024, N5015, N3126);
not NOT1 (N5025, N4972);
nor NOR3 (N5026, N5021, N600, N3911);
not NOT1 (N5027, N5022);
nor NOR3 (N5028, N5026, N4520, N3102);
xor XOR2 (N5029, N4995, N354);
nor NOR2 (N5030, N5028, N4472);
or OR3 (N5031, N5029, N4129, N4807);
and AND3 (N5032, N5017, N1855, N1250);
xor XOR2 (N5033, N5030, N1806);
and AND3 (N5034, N5020, N4341, N269);
and AND3 (N5035, N5033, N429, N1004);
nor NOR3 (N5036, N5027, N4778, N147);
nor NOR3 (N5037, N5018, N1404, N3693);
or OR4 (N5038, N5032, N1265, N2568, N3893);
not NOT1 (N5039, N5016);
not NOT1 (N5040, N5038);
nor NOR2 (N5041, N5031, N1799);
and AND2 (N5042, N5036, N3288);
nand NAND4 (N5043, N5037, N2641, N798, N3415);
and AND2 (N5044, N5040, N629);
nand NAND2 (N5045, N5044, N4522);
and AND3 (N5046, N5035, N1855, N984);
and AND3 (N5047, N5041, N4987, N1157);
buf BUF1 (N5048, N5023);
or OR3 (N5049, N5048, N1083, N1899);
or OR3 (N5050, N5045, N448, N2626);
nand NAND4 (N5051, N5049, N2723, N3859, N988);
xor XOR2 (N5052, N5050, N2490);
xor XOR2 (N5053, N5025, N1324);
not NOT1 (N5054, N5039);
nand NAND2 (N5055, N5047, N2415);
or OR4 (N5056, N5055, N3493, N1173, N1577);
and AND2 (N5057, N5056, N9);
and AND2 (N5058, N5051, N299);
xor XOR2 (N5059, N5043, N1239);
xor XOR2 (N5060, N5058, N2182);
not NOT1 (N5061, N5042);
buf BUF1 (N5062, N5057);
not NOT1 (N5063, N5054);
nor NOR3 (N5064, N5059, N3766, N4680);
not NOT1 (N5065, N5052);
nor NOR4 (N5066, N5046, N2648, N4278, N1551);
not NOT1 (N5067, N5024);
and AND2 (N5068, N5060, N4930);
nand NAND2 (N5069, N5062, N1939);
nor NOR4 (N5070, N5066, N1705, N2924, N2088);
xor XOR2 (N5071, N5061, N665);
xor XOR2 (N5072, N5070, N1847);
not NOT1 (N5073, N5064);
and AND4 (N5074, N5068, N531, N3485, N2020);
and AND2 (N5075, N5053, N2077);
and AND4 (N5076, N5074, N667, N3999, N2031);
not NOT1 (N5077, N5067);
xor XOR2 (N5078, N5034, N3162);
and AND4 (N5079, N5075, N4098, N1090, N2102);
nor NOR3 (N5080, N5079, N996, N4603);
xor XOR2 (N5081, N5077, N3914);
xor XOR2 (N5082, N5069, N2630);
not NOT1 (N5083, N5078);
or OR3 (N5084, N5072, N4587, N2177);
and AND2 (N5085, N5084, N813);
buf BUF1 (N5086, N5063);
buf BUF1 (N5087, N5085);
nand NAND4 (N5088, N5087, N3937, N4960, N3753);
xor XOR2 (N5089, N5080, N4947);
and AND3 (N5090, N5089, N3873, N2953);
not NOT1 (N5091, N5088);
or OR3 (N5092, N5086, N1651, N1298);
xor XOR2 (N5093, N5065, N960);
or OR3 (N5094, N5090, N4257, N4022);
nand NAND3 (N5095, N5094, N4518, N998);
nor NOR3 (N5096, N5091, N3117, N3913);
and AND3 (N5097, N5082, N3558, N3017);
or OR4 (N5098, N5092, N3863, N286, N4953);
nor NOR4 (N5099, N5095, N4477, N796, N2230);
xor XOR2 (N5100, N5099, N3046);
not NOT1 (N5101, N5083);
not NOT1 (N5102, N5096);
buf BUF1 (N5103, N5097);
buf BUF1 (N5104, N5101);
and AND4 (N5105, N5103, N4174, N1897, N21);
xor XOR2 (N5106, N5100, N2987);
buf BUF1 (N5107, N5104);
buf BUF1 (N5108, N5105);
xor XOR2 (N5109, N5098, N4149);
buf BUF1 (N5110, N5093);
or OR3 (N5111, N5106, N751, N1476);
buf BUF1 (N5112, N5108);
nor NOR2 (N5113, N5102, N1086);
or OR4 (N5114, N5081, N460, N3513, N4572);
nand NAND2 (N5115, N5076, N3865);
buf BUF1 (N5116, N5113);
nand NAND2 (N5117, N5110, N2223);
xor XOR2 (N5118, N5114, N4391);
xor XOR2 (N5119, N5116, N359);
buf BUF1 (N5120, N5119);
and AND2 (N5121, N5118, N25);
buf BUF1 (N5122, N5111);
nor NOR2 (N5123, N5107, N1896);
and AND3 (N5124, N5071, N3416, N173);
nand NAND4 (N5125, N5109, N1557, N3127, N3361);
xor XOR2 (N5126, N5122, N3663);
nor NOR3 (N5127, N5115, N2853, N1535);
not NOT1 (N5128, N5123);
nor NOR3 (N5129, N5128, N3068, N2648);
nand NAND2 (N5130, N5117, N4938);
xor XOR2 (N5131, N5126, N1401);
buf BUF1 (N5132, N5121);
or OR4 (N5133, N5073, N3067, N2608, N3494);
and AND3 (N5134, N5130, N4695, N1306);
buf BUF1 (N5135, N5112);
buf BUF1 (N5136, N5132);
nand NAND4 (N5137, N5120, N842, N2276, N4459);
xor XOR2 (N5138, N5133, N2563);
not NOT1 (N5139, N5137);
and AND2 (N5140, N5139, N1465);
or OR4 (N5141, N5127, N1733, N491, N162);
xor XOR2 (N5142, N5141, N3267);
or OR2 (N5143, N5124, N1739);
nand NAND2 (N5144, N5142, N5077);
not NOT1 (N5145, N5136);
and AND2 (N5146, N5145, N896);
buf BUF1 (N5147, N5144);
not NOT1 (N5148, N5146);
or OR2 (N5149, N5143, N3142);
or OR4 (N5150, N5148, N4328, N3956, N4775);
or OR3 (N5151, N5131, N2154, N2308);
xor XOR2 (N5152, N5134, N1832);
not NOT1 (N5153, N5129);
xor XOR2 (N5154, N5150, N2938);
or OR3 (N5155, N5152, N4320, N2024);
not NOT1 (N5156, N5151);
or OR2 (N5157, N5153, N1700);
xor XOR2 (N5158, N5157, N143);
and AND3 (N5159, N5125, N3761, N409);
buf BUF1 (N5160, N5140);
nand NAND3 (N5161, N5155, N4586, N3051);
not NOT1 (N5162, N5159);
nor NOR3 (N5163, N5162, N2194, N2741);
buf BUF1 (N5164, N5160);
xor XOR2 (N5165, N5163, N2871);
nor NOR3 (N5166, N5147, N2859, N1222);
and AND4 (N5167, N5161, N124, N5060, N3868);
or OR4 (N5168, N5158, N1005, N1168, N2494);
buf BUF1 (N5169, N5154);
and AND4 (N5170, N5149, N2426, N1687, N2663);
or OR3 (N5171, N5156, N2844, N961);
nand NAND2 (N5172, N5169, N4703);
and AND3 (N5173, N5172, N3291, N4870);
and AND2 (N5174, N5170, N4479);
and AND4 (N5175, N5166, N619, N3379, N3792);
buf BUF1 (N5176, N5173);
and AND4 (N5177, N5135, N2631, N1779, N775);
or OR2 (N5178, N5174, N2970);
and AND2 (N5179, N5168, N3990);
nor NOR4 (N5180, N5178, N1511, N4063, N3342);
nand NAND4 (N5181, N5165, N4817, N4432, N4815);
not NOT1 (N5182, N5180);
buf BUF1 (N5183, N5138);
xor XOR2 (N5184, N5171, N594);
and AND3 (N5185, N5182, N4319, N3900);
nor NOR4 (N5186, N5181, N1341, N1140, N3750);
nand NAND3 (N5187, N5184, N2868, N2328);
nand NAND2 (N5188, N5183, N2191);
and AND3 (N5189, N5175, N1676, N502);
or OR4 (N5190, N5177, N2141, N781, N1353);
and AND4 (N5191, N5167, N3124, N2758, N630);
and AND3 (N5192, N5179, N4886, N1900);
nor NOR2 (N5193, N5176, N2502);
nor NOR4 (N5194, N5189, N3114, N4034, N4057);
or OR2 (N5195, N5191, N566);
and AND4 (N5196, N5188, N3978, N29, N509);
nand NAND4 (N5197, N5190, N1248, N4738, N1594);
nor NOR2 (N5198, N5197, N3311);
buf BUF1 (N5199, N5196);
nor NOR2 (N5200, N5195, N1621);
and AND3 (N5201, N5194, N3156, N1206);
buf BUF1 (N5202, N5187);
nand NAND2 (N5203, N5200, N1337);
xor XOR2 (N5204, N5193, N3513);
nand NAND4 (N5205, N5164, N82, N2750, N3847);
nand NAND3 (N5206, N5185, N1052, N1956);
xor XOR2 (N5207, N5204, N2677);
nor NOR3 (N5208, N5198, N1174, N2539);
not NOT1 (N5209, N5202);
or OR2 (N5210, N5203, N3769);
not NOT1 (N5211, N5208);
xor XOR2 (N5212, N5199, N4789);
nor NOR3 (N5213, N5211, N2809, N1577);
xor XOR2 (N5214, N5186, N610);
xor XOR2 (N5215, N5210, N2005);
nand NAND4 (N5216, N5206, N4196, N2561, N955);
and AND4 (N5217, N5213, N2227, N3256, N1327);
and AND2 (N5218, N5192, N4837);
or OR4 (N5219, N5205, N757, N4736, N4372);
or OR2 (N5220, N5218, N5110);
xor XOR2 (N5221, N5217, N608);
not NOT1 (N5222, N5215);
nand NAND4 (N5223, N5222, N2380, N5150, N4029);
xor XOR2 (N5224, N5219, N2695);
or OR2 (N5225, N5221, N3731);
buf BUF1 (N5226, N5207);
nand NAND4 (N5227, N5225, N2992, N916, N983);
nand NAND3 (N5228, N5201, N3243, N5021);
and AND3 (N5229, N5209, N4209, N2719);
nand NAND3 (N5230, N5216, N2721, N1758);
or OR2 (N5231, N5228, N5107);
or OR4 (N5232, N5214, N2273, N257, N1951);
xor XOR2 (N5233, N5223, N3730);
not NOT1 (N5234, N5229);
and AND3 (N5235, N5224, N3948, N546);
xor XOR2 (N5236, N5227, N2);
xor XOR2 (N5237, N5233, N1929);
or OR2 (N5238, N5220, N929);
buf BUF1 (N5239, N5237);
nor NOR4 (N5240, N5232, N1444, N3580, N4639);
and AND4 (N5241, N5236, N1638, N2649, N4090);
xor XOR2 (N5242, N5239, N2244);
not NOT1 (N5243, N5234);
or OR3 (N5244, N5235, N3893, N3409);
or OR3 (N5245, N5244, N4153, N2582);
and AND3 (N5246, N5243, N2736, N1040);
not NOT1 (N5247, N5240);
nor NOR2 (N5248, N5246, N347);
or OR2 (N5249, N5242, N457);
not NOT1 (N5250, N5241);
and AND2 (N5251, N5212, N3077);
nor NOR2 (N5252, N5249, N468);
buf BUF1 (N5253, N5226);
or OR3 (N5254, N5253, N4472, N3447);
nor NOR2 (N5255, N5230, N2015);
and AND4 (N5256, N5252, N5141, N5177, N5164);
or OR3 (N5257, N5255, N3721, N1590);
not NOT1 (N5258, N5238);
and AND4 (N5259, N5251, N2788, N2266, N1669);
and AND2 (N5260, N5259, N2083);
or OR2 (N5261, N5248, N2115);
nand NAND3 (N5262, N5247, N2310, N4593);
not NOT1 (N5263, N5256);
nand NAND4 (N5264, N5250, N3078, N4160, N88);
not NOT1 (N5265, N5245);
nor NOR2 (N5266, N5231, N3296);
not NOT1 (N5267, N5260);
not NOT1 (N5268, N5258);
buf BUF1 (N5269, N5263);
xor XOR2 (N5270, N5262, N3161);
not NOT1 (N5271, N5265);
buf BUF1 (N5272, N5268);
not NOT1 (N5273, N5270);
nor NOR2 (N5274, N5271, N3149);
xor XOR2 (N5275, N5257, N2212);
xor XOR2 (N5276, N5274, N3187);
and AND4 (N5277, N5267, N3351, N3133, N1986);
or OR2 (N5278, N5269, N2246);
not NOT1 (N5279, N5272);
nor NOR4 (N5280, N5279, N3764, N1506, N1732);
buf BUF1 (N5281, N5277);
nor NOR2 (N5282, N5276, N973);
nand NAND3 (N5283, N5281, N2253, N2920);
xor XOR2 (N5284, N5264, N2861);
nor NOR2 (N5285, N5278, N3229);
buf BUF1 (N5286, N5280);
nor NOR4 (N5287, N5284, N63, N3917, N5120);
or OR4 (N5288, N5285, N5145, N945, N4680);
or OR4 (N5289, N5283, N185, N236, N489);
and AND4 (N5290, N5282, N802, N1276, N3542);
and AND3 (N5291, N5254, N3663, N214);
or OR3 (N5292, N5290, N2642, N359);
nand NAND4 (N5293, N5289, N2661, N202, N2297);
and AND3 (N5294, N5292, N5174, N1179);
not NOT1 (N5295, N5261);
not NOT1 (N5296, N5266);
xor XOR2 (N5297, N5275, N4809);
and AND2 (N5298, N5287, N4998);
nand NAND3 (N5299, N5273, N339, N258);
or OR3 (N5300, N5298, N995, N2313);
buf BUF1 (N5301, N5300);
nand NAND4 (N5302, N5293, N3450, N5254, N3546);
xor XOR2 (N5303, N5299, N4912);
and AND2 (N5304, N5302, N231);
nand NAND3 (N5305, N5301, N2606, N3222);
nand NAND3 (N5306, N5303, N2183, N1698);
xor XOR2 (N5307, N5286, N972);
not NOT1 (N5308, N5305);
nor NOR2 (N5309, N5308, N3954);
nand NAND3 (N5310, N5304, N3040, N64);
or OR4 (N5311, N5295, N2629, N834, N3500);
and AND3 (N5312, N5294, N3988, N2164);
buf BUF1 (N5313, N5288);
xor XOR2 (N5314, N5311, N22);
xor XOR2 (N5315, N5307, N1346);
not NOT1 (N5316, N5297);
buf BUF1 (N5317, N5315);
or OR3 (N5318, N5316, N593, N4425);
nor NOR4 (N5319, N5296, N5111, N498, N1047);
nand NAND2 (N5320, N5312, N990);
nand NAND4 (N5321, N5320, N5130, N1625, N1336);
xor XOR2 (N5322, N5321, N1510);
not NOT1 (N5323, N5322);
not NOT1 (N5324, N5309);
nand NAND3 (N5325, N5323, N4270, N2566);
xor XOR2 (N5326, N5324, N2284);
or OR4 (N5327, N5310, N2818, N2486, N4886);
or OR3 (N5328, N5319, N622, N4852);
xor XOR2 (N5329, N5328, N2289);
not NOT1 (N5330, N5325);
or OR2 (N5331, N5329, N2390);
nand NAND2 (N5332, N5330, N2800);
not NOT1 (N5333, N5313);
and AND4 (N5334, N5314, N3149, N2024, N5289);
nor NOR3 (N5335, N5333, N3178, N4145);
nor NOR4 (N5336, N5331, N3136, N4493, N2981);
buf BUF1 (N5337, N5306);
buf BUF1 (N5338, N5336);
not NOT1 (N5339, N5337);
xor XOR2 (N5340, N5332, N1091);
and AND2 (N5341, N5326, N1486);
buf BUF1 (N5342, N5338);
not NOT1 (N5343, N5339);
nor NOR3 (N5344, N5327, N3162, N3943);
or OR2 (N5345, N5343, N2782);
or OR3 (N5346, N5344, N1353, N1266);
and AND2 (N5347, N5341, N3491);
not NOT1 (N5348, N5334);
and AND2 (N5349, N5318, N1735);
nand NAND3 (N5350, N5347, N561, N4533);
xor XOR2 (N5351, N5335, N4993);
nor NOR4 (N5352, N5342, N2177, N4219, N121);
xor XOR2 (N5353, N5352, N2830);
nand NAND4 (N5354, N5348, N4582, N4951, N1151);
xor XOR2 (N5355, N5291, N1170);
nor NOR2 (N5356, N5340, N3436);
not NOT1 (N5357, N5349);
nor NOR2 (N5358, N5346, N4598);
buf BUF1 (N5359, N5358);
buf BUF1 (N5360, N5350);
xor XOR2 (N5361, N5354, N2002);
and AND3 (N5362, N5356, N5319, N2375);
nand NAND4 (N5363, N5357, N2423, N3235, N1476);
or OR2 (N5364, N5360, N2237);
not NOT1 (N5365, N5359);
not NOT1 (N5366, N5317);
nor NOR4 (N5367, N5362, N2658, N2647, N2179);
and AND2 (N5368, N5355, N146);
xor XOR2 (N5369, N5361, N4761);
or OR3 (N5370, N5353, N1403, N2406);
nand NAND4 (N5371, N5364, N3546, N5312, N4708);
buf BUF1 (N5372, N5371);
and AND2 (N5373, N5351, N2789);
or OR2 (N5374, N5365, N5194);
xor XOR2 (N5375, N5370, N55);
and AND2 (N5376, N5372, N2451);
buf BUF1 (N5377, N5345);
nand NAND4 (N5378, N5363, N3865, N4812, N4244);
nand NAND3 (N5379, N5367, N3837, N4616);
buf BUF1 (N5380, N5378);
nor NOR4 (N5381, N5376, N4828, N2840, N258);
nand NAND3 (N5382, N5379, N2911, N4592);
or OR3 (N5383, N5382, N4295, N3383);
and AND3 (N5384, N5383, N4980, N3427);
xor XOR2 (N5385, N5381, N3790);
xor XOR2 (N5386, N5373, N4486);
nor NOR3 (N5387, N5368, N3443, N2776);
and AND4 (N5388, N5384, N2399, N2887, N1316);
or OR2 (N5389, N5369, N3117);
buf BUF1 (N5390, N5386);
nor NOR2 (N5391, N5374, N2613);
buf BUF1 (N5392, N5390);
nor NOR2 (N5393, N5392, N419);
or OR4 (N5394, N5375, N2823, N2340, N2185);
not NOT1 (N5395, N5366);
and AND2 (N5396, N5380, N1158);
buf BUF1 (N5397, N5387);
xor XOR2 (N5398, N5396, N815);
xor XOR2 (N5399, N5377, N4144);
xor XOR2 (N5400, N5388, N1387);
nand NAND2 (N5401, N5389, N1150);
xor XOR2 (N5402, N5400, N1950);
nor NOR3 (N5403, N5398, N106, N864);
not NOT1 (N5404, N5399);
nor NOR2 (N5405, N5393, N3698);
not NOT1 (N5406, N5397);
buf BUF1 (N5407, N5405);
xor XOR2 (N5408, N5406, N1650);
buf BUF1 (N5409, N5402);
and AND2 (N5410, N5385, N3324);
buf BUF1 (N5411, N5408);
buf BUF1 (N5412, N5391);
or OR3 (N5413, N5410, N1198, N880);
not NOT1 (N5414, N5394);
or OR4 (N5415, N5407, N2215, N1637, N1675);
and AND2 (N5416, N5403, N3757);
nor NOR3 (N5417, N5412, N332, N2028);
xor XOR2 (N5418, N5411, N1261);
nor NOR3 (N5419, N5413, N3384, N3142);
nor NOR4 (N5420, N5419, N633, N527, N269);
and AND4 (N5421, N5409, N290, N304, N3223);
buf BUF1 (N5422, N5395);
not NOT1 (N5423, N5420);
and AND3 (N5424, N5414, N1053, N1037);
nor NOR2 (N5425, N5417, N1993);
or OR4 (N5426, N5416, N3593, N1386, N5129);
not NOT1 (N5427, N5421);
nand NAND4 (N5428, N5401, N5094, N510, N4235);
not NOT1 (N5429, N5427);
xor XOR2 (N5430, N5426, N450);
nand NAND2 (N5431, N5429, N1889);
xor XOR2 (N5432, N5430, N5080);
nand NAND3 (N5433, N5404, N2930, N1832);
or OR3 (N5434, N5425, N621, N199);
nand NAND4 (N5435, N5418, N1537, N2498, N2550);
not NOT1 (N5436, N5435);
not NOT1 (N5437, N5424);
not NOT1 (N5438, N5423);
or OR3 (N5439, N5432, N2969, N2546);
xor XOR2 (N5440, N5438, N268);
and AND2 (N5441, N5439, N2584);
nor NOR3 (N5442, N5431, N2245, N1553);
nand NAND2 (N5443, N5434, N1271);
and AND2 (N5444, N5433, N1839);
not NOT1 (N5445, N5444);
and AND4 (N5446, N5422, N4387, N4433, N357);
nand NAND4 (N5447, N5440, N3169, N2549, N1281);
not NOT1 (N5448, N5428);
and AND4 (N5449, N5441, N4772, N2124, N4043);
nand NAND4 (N5450, N5436, N4509, N2477, N2087);
not NOT1 (N5451, N5447);
or OR3 (N5452, N5451, N4596, N2728);
buf BUF1 (N5453, N5446);
xor XOR2 (N5454, N5448, N1246);
xor XOR2 (N5455, N5415, N4171);
xor XOR2 (N5456, N5449, N2648);
xor XOR2 (N5457, N5454, N4909);
nor NOR3 (N5458, N5456, N5312, N5298);
and AND4 (N5459, N5453, N744, N5121, N3581);
buf BUF1 (N5460, N5450);
or OR3 (N5461, N5457, N511, N3342);
nor NOR4 (N5462, N5459, N4918, N3371, N3659);
or OR3 (N5463, N5445, N1397, N5173);
not NOT1 (N5464, N5460);
nor NOR4 (N5465, N5455, N799, N4797, N4617);
and AND4 (N5466, N5461, N681, N1153, N3356);
xor XOR2 (N5467, N5462, N2142);
buf BUF1 (N5468, N5443);
and AND3 (N5469, N5464, N97, N3576);
nand NAND2 (N5470, N5463, N5037);
xor XOR2 (N5471, N5458, N2194);
xor XOR2 (N5472, N5468, N4464);
and AND3 (N5473, N5465, N342, N2675);
and AND4 (N5474, N5442, N2087, N354, N1285);
and AND2 (N5475, N5437, N648);
nor NOR2 (N5476, N5470, N5022);
nor NOR3 (N5477, N5466, N3579, N515);
or OR4 (N5478, N5475, N1957, N1541, N2407);
or OR4 (N5479, N5467, N2957, N4077, N3223);
or OR4 (N5480, N5472, N3168, N693, N1965);
and AND3 (N5481, N5469, N3729, N4584);
not NOT1 (N5482, N5474);
xor XOR2 (N5483, N5480, N5107);
not NOT1 (N5484, N5476);
nand NAND4 (N5485, N5484, N4898, N80, N3125);
nor NOR4 (N5486, N5477, N2365, N73, N2782);
buf BUF1 (N5487, N5452);
and AND3 (N5488, N5486, N4882, N735);
and AND2 (N5489, N5485, N5461);
nor NOR4 (N5490, N5489, N4702, N1007, N1216);
or OR2 (N5491, N5481, N5222);
not NOT1 (N5492, N5471);
or OR4 (N5493, N5487, N1078, N4872, N4549);
nand NAND3 (N5494, N5490, N5387, N62);
nor NOR3 (N5495, N5492, N256, N422);
or OR4 (N5496, N5488, N3745, N3775, N3845);
not NOT1 (N5497, N5491);
xor XOR2 (N5498, N5497, N1782);
and AND3 (N5499, N5479, N2849, N3232);
not NOT1 (N5500, N5498);
or OR3 (N5501, N5496, N892, N5226);
xor XOR2 (N5502, N5495, N5282);
xor XOR2 (N5503, N5501, N2462);
buf BUF1 (N5504, N5483);
buf BUF1 (N5505, N5504);
xor XOR2 (N5506, N5482, N2268);
not NOT1 (N5507, N5499);
nand NAND3 (N5508, N5493, N377, N5332);
nand NAND2 (N5509, N5507, N2524);
or OR4 (N5510, N5478, N41, N5473, N4942);
nor NOR4 (N5511, N4308, N390, N3688, N5029);
buf BUF1 (N5512, N5494);
xor XOR2 (N5513, N5512, N5131);
not NOT1 (N5514, N5511);
xor XOR2 (N5515, N5513, N5442);
buf BUF1 (N5516, N5502);
and AND2 (N5517, N5510, N3949);
buf BUF1 (N5518, N5503);
xor XOR2 (N5519, N5506, N5409);
or OR3 (N5520, N5514, N2790, N2951);
and AND2 (N5521, N5518, N4152);
or OR4 (N5522, N5521, N2398, N314, N897);
and AND4 (N5523, N5517, N952, N25, N5498);
or OR4 (N5524, N5519, N5069, N46, N185);
and AND4 (N5525, N5523, N894, N2029, N54);
nand NAND3 (N5526, N5525, N2918, N3318);
xor XOR2 (N5527, N5509, N4181);
nand NAND3 (N5528, N5505, N1026, N809);
nor NOR4 (N5529, N5524, N104, N5467, N3957);
and AND2 (N5530, N5515, N130);
and AND3 (N5531, N5528, N1384, N392);
xor XOR2 (N5532, N5530, N2251);
nor NOR3 (N5533, N5500, N889, N836);
not NOT1 (N5534, N5531);
not NOT1 (N5535, N5508);
and AND2 (N5536, N5529, N865);
and AND4 (N5537, N5534, N523, N660, N1756);
and AND2 (N5538, N5535, N642);
nor NOR4 (N5539, N5533, N572, N1373, N386);
nand NAND2 (N5540, N5520, N4364);
and AND4 (N5541, N5527, N2158, N4582, N5234);
not NOT1 (N5542, N5536);
buf BUF1 (N5543, N5522);
buf BUF1 (N5544, N5539);
nor NOR2 (N5545, N5541, N4883);
nor NOR3 (N5546, N5538, N2251, N269);
not NOT1 (N5547, N5546);
nand NAND4 (N5548, N5547, N5249, N5295, N5489);
nor NOR4 (N5549, N5542, N3370, N4144, N4562);
buf BUF1 (N5550, N5549);
buf BUF1 (N5551, N5548);
nor NOR4 (N5552, N5545, N2828, N5422, N2239);
buf BUF1 (N5553, N5540);
or OR3 (N5554, N5552, N4016, N5453);
and AND2 (N5555, N5544, N1043);
nand NAND3 (N5556, N5551, N1003, N4108);
not NOT1 (N5557, N5516);
buf BUF1 (N5558, N5554);
buf BUF1 (N5559, N5553);
buf BUF1 (N5560, N5543);
buf BUF1 (N5561, N5532);
nand NAND4 (N5562, N5555, N754, N2475, N2713);
or OR2 (N5563, N5550, N2392);
not NOT1 (N5564, N5556);
and AND4 (N5565, N5559, N398, N959, N1070);
and AND4 (N5566, N5565, N2818, N369, N1004);
buf BUF1 (N5567, N5537);
not NOT1 (N5568, N5558);
xor XOR2 (N5569, N5560, N5057);
and AND2 (N5570, N5564, N973);
xor XOR2 (N5571, N5561, N1860);
or OR4 (N5572, N5568, N43, N2141, N3375);
nand NAND2 (N5573, N5572, N1722);
nor NOR3 (N5574, N5567, N4963, N2884);
xor XOR2 (N5575, N5573, N1380);
buf BUF1 (N5576, N5526);
not NOT1 (N5577, N5569);
xor XOR2 (N5578, N5562, N14);
and AND2 (N5579, N5576, N2973);
or OR4 (N5580, N5570, N2837, N380, N3602);
xor XOR2 (N5581, N5566, N2194);
buf BUF1 (N5582, N5563);
and AND4 (N5583, N5581, N1061, N4307, N1697);
nor NOR2 (N5584, N5583, N905);
and AND2 (N5585, N5579, N2919);
nand NAND2 (N5586, N5571, N3538);
nor NOR4 (N5587, N5574, N730, N4199, N979);
and AND2 (N5588, N5577, N5491);
or OR3 (N5589, N5585, N5223, N4480);
nor NOR2 (N5590, N5587, N1555);
xor XOR2 (N5591, N5589, N1570);
or OR2 (N5592, N5557, N4582);
nor NOR4 (N5593, N5586, N95, N2768, N4746);
and AND2 (N5594, N5592, N5455);
nand NAND4 (N5595, N5590, N4137, N1297, N1985);
or OR4 (N5596, N5584, N680, N4750, N4571);
nor NOR3 (N5597, N5578, N4219, N4343);
and AND2 (N5598, N5580, N4508);
nand NAND3 (N5599, N5596, N3534, N3653);
nand NAND3 (N5600, N5593, N3099, N2442);
buf BUF1 (N5601, N5599);
nor NOR3 (N5602, N5588, N3920, N193);
buf BUF1 (N5603, N5582);
and AND2 (N5604, N5602, N3267);
nor NOR3 (N5605, N5595, N4907, N1434);
nor NOR2 (N5606, N5604, N2889);
xor XOR2 (N5607, N5594, N1258);
nand NAND3 (N5608, N5601, N2548, N3543);
nor NOR4 (N5609, N5606, N2082, N2850, N3352);
nor NOR4 (N5610, N5600, N2687, N1238, N4580);
buf BUF1 (N5611, N5591);
or OR3 (N5612, N5598, N3470, N4264);
and AND2 (N5613, N5610, N939);
or OR2 (N5614, N5605, N4231);
or OR2 (N5615, N5607, N5163);
xor XOR2 (N5616, N5612, N873);
nor NOR4 (N5617, N5609, N3866, N1345, N82);
buf BUF1 (N5618, N5616);
nor NOR4 (N5619, N5613, N5334, N3018, N5285);
or OR2 (N5620, N5619, N3088);
and AND4 (N5621, N5614, N5467, N151, N1117);
not NOT1 (N5622, N5618);
nand NAND4 (N5623, N5615, N1897, N4063, N4715);
nor NOR2 (N5624, N5617, N2431);
nand NAND3 (N5625, N5623, N3988, N2285);
nor NOR2 (N5626, N5622, N2427);
buf BUF1 (N5627, N5608);
or OR4 (N5628, N5620, N5592, N2385, N1612);
nand NAND3 (N5629, N5575, N3051, N859);
nor NOR3 (N5630, N5624, N5025, N390);
nand NAND2 (N5631, N5625, N3991);
not NOT1 (N5632, N5597);
and AND3 (N5633, N5630, N3962, N3247);
and AND3 (N5634, N5611, N3225, N4465);
nand NAND2 (N5635, N5628, N1938);
and AND3 (N5636, N5629, N2833, N737);
or OR4 (N5637, N5633, N2134, N3992, N3461);
xor XOR2 (N5638, N5603, N1752);
nand NAND2 (N5639, N5635, N4084);
or OR3 (N5640, N5638, N4149, N5277);
and AND3 (N5641, N5621, N1331, N2410);
xor XOR2 (N5642, N5636, N5130);
or OR3 (N5643, N5642, N2420, N817);
nand NAND2 (N5644, N5627, N1584);
nor NOR3 (N5645, N5626, N2800, N1786);
buf BUF1 (N5646, N5643);
nand NAND4 (N5647, N5632, N199, N4726, N2078);
buf BUF1 (N5648, N5646);
and AND2 (N5649, N5637, N1493);
not NOT1 (N5650, N5648);
not NOT1 (N5651, N5639);
or OR3 (N5652, N5634, N278, N1941);
nor NOR3 (N5653, N5651, N3358, N1556);
and AND3 (N5654, N5645, N5458, N3076);
not NOT1 (N5655, N5641);
nor NOR3 (N5656, N5650, N3735, N5645);
xor XOR2 (N5657, N5653, N3174);
nor NOR3 (N5658, N5649, N4315, N909);
or OR4 (N5659, N5644, N518, N1601, N4218);
nand NAND2 (N5660, N5647, N3006);
nand NAND3 (N5661, N5656, N4339, N4487);
nor NOR4 (N5662, N5659, N510, N1634, N1662);
or OR2 (N5663, N5658, N4441);
xor XOR2 (N5664, N5640, N1481);
xor XOR2 (N5665, N5655, N5084);
nand NAND4 (N5666, N5662, N1170, N4888, N4082);
buf BUF1 (N5667, N5652);
not NOT1 (N5668, N5661);
not NOT1 (N5669, N5654);
not NOT1 (N5670, N5657);
xor XOR2 (N5671, N5660, N1282);
or OR2 (N5672, N5670, N1237);
nor NOR2 (N5673, N5664, N3071);
or OR4 (N5674, N5665, N4693, N4086, N3210);
or OR2 (N5675, N5672, N1398);
not NOT1 (N5676, N5667);
and AND2 (N5677, N5631, N4705);
xor XOR2 (N5678, N5676, N1100);
not NOT1 (N5679, N5666);
or OR3 (N5680, N5663, N2619, N800);
xor XOR2 (N5681, N5678, N1364);
xor XOR2 (N5682, N5669, N3583);
buf BUF1 (N5683, N5674);
or OR2 (N5684, N5679, N3657);
nor NOR3 (N5685, N5683, N4077, N1161);
xor XOR2 (N5686, N5685, N4539);
nor NOR4 (N5687, N5677, N247, N1486, N395);
xor XOR2 (N5688, N5687, N1718);
buf BUF1 (N5689, N5680);
nand NAND3 (N5690, N5688, N1271, N1556);
xor XOR2 (N5691, N5675, N1463);
nor NOR3 (N5692, N5690, N1187, N3634);
or OR4 (N5693, N5691, N1446, N4787, N2353);
xor XOR2 (N5694, N5681, N5363);
or OR3 (N5695, N5689, N97, N1783);
not NOT1 (N5696, N5692);
buf BUF1 (N5697, N5671);
or OR3 (N5698, N5696, N3888, N5382);
buf BUF1 (N5699, N5697);
xor XOR2 (N5700, N5694, N4512);
nor NOR3 (N5701, N5698, N3712, N5194);
or OR2 (N5702, N5686, N5507);
not NOT1 (N5703, N5693);
and AND2 (N5704, N5700, N46);
nor NOR4 (N5705, N5699, N2782, N2134, N2807);
xor XOR2 (N5706, N5695, N2445);
nand NAND3 (N5707, N5682, N3701, N5521);
or OR4 (N5708, N5673, N2511, N4426, N3254);
xor XOR2 (N5709, N5703, N547);
and AND4 (N5710, N5706, N4398, N2403, N1751);
xor XOR2 (N5711, N5708, N352);
xor XOR2 (N5712, N5707, N4360);
buf BUF1 (N5713, N5710);
buf BUF1 (N5714, N5709);
not NOT1 (N5715, N5701);
nand NAND2 (N5716, N5715, N58);
xor XOR2 (N5717, N5704, N3440);
not NOT1 (N5718, N5711);
not NOT1 (N5719, N5713);
and AND3 (N5720, N5714, N4290, N887);
nor NOR2 (N5721, N5702, N2395);
nor NOR3 (N5722, N5721, N23, N4220);
xor XOR2 (N5723, N5717, N5452);
xor XOR2 (N5724, N5718, N2872);
nand NAND3 (N5725, N5668, N3290, N2831);
nor NOR4 (N5726, N5720, N3566, N5599, N4265);
nand NAND4 (N5727, N5716, N3190, N325, N2504);
and AND2 (N5728, N5705, N218);
not NOT1 (N5729, N5728);
nand NAND4 (N5730, N5724, N3714, N2167, N1941);
nand NAND2 (N5731, N5727, N340);
buf BUF1 (N5732, N5712);
not NOT1 (N5733, N5725);
nand NAND4 (N5734, N5719, N5569, N1561, N2767);
nor NOR2 (N5735, N5726, N4128);
xor XOR2 (N5736, N5731, N5072);
xor XOR2 (N5737, N5684, N2220);
nand NAND4 (N5738, N5722, N332, N2234, N3817);
not NOT1 (N5739, N5730);
buf BUF1 (N5740, N5723);
nor NOR2 (N5741, N5736, N2176);
nor NOR3 (N5742, N5739, N24, N2219);
not NOT1 (N5743, N5732);
buf BUF1 (N5744, N5734);
nor NOR3 (N5745, N5729, N2754, N1159);
nand NAND3 (N5746, N5737, N2275, N319);
nand NAND4 (N5747, N5744, N1558, N2886, N3058);
and AND4 (N5748, N5745, N3145, N4434, N393);
or OR4 (N5749, N5735, N1083, N4422, N1900);
or OR2 (N5750, N5738, N275);
nand NAND4 (N5751, N5740, N862, N2245, N4220);
not NOT1 (N5752, N5749);
and AND2 (N5753, N5751, N3767);
or OR4 (N5754, N5753, N5665, N3958, N1273);
nand NAND2 (N5755, N5741, N4670);
nand NAND4 (N5756, N5733, N775, N5694, N1801);
nor NOR3 (N5757, N5755, N840, N3854);
nand NAND3 (N5758, N5757, N4248, N4977);
or OR4 (N5759, N5756, N5379, N279, N1241);
nor NOR4 (N5760, N5759, N2982, N3361, N3721);
xor XOR2 (N5761, N5750, N4635);
nand NAND4 (N5762, N5748, N432, N4730, N1450);
xor XOR2 (N5763, N5761, N1941);
and AND4 (N5764, N5760, N667, N3592, N5244);
buf BUF1 (N5765, N5758);
xor XOR2 (N5766, N5746, N1642);
buf BUF1 (N5767, N5764);
nor NOR4 (N5768, N5765, N1073, N2470, N1434);
not NOT1 (N5769, N5752);
not NOT1 (N5770, N5754);
nor NOR3 (N5771, N5770, N1334, N1233);
and AND4 (N5772, N5742, N5550, N155, N4928);
not NOT1 (N5773, N5769);
or OR2 (N5774, N5743, N1682);
or OR4 (N5775, N5774, N3367, N4399, N784);
buf BUF1 (N5776, N5747);
buf BUF1 (N5777, N5766);
buf BUF1 (N5778, N5768);
not NOT1 (N5779, N5772);
or OR3 (N5780, N5762, N5656, N2059);
nand NAND3 (N5781, N5767, N5486, N5476);
nor NOR4 (N5782, N5763, N405, N3845, N2532);
or OR2 (N5783, N5773, N5228);
nor NOR4 (N5784, N5776, N2279, N2044, N3628);
and AND4 (N5785, N5783, N2563, N4061, N2771);
buf BUF1 (N5786, N5781);
and AND4 (N5787, N5784, N2661, N3673, N3494);
and AND2 (N5788, N5778, N3615);
xor XOR2 (N5789, N5782, N4299);
nand NAND4 (N5790, N5786, N4336, N3261, N5524);
nor NOR4 (N5791, N5785, N1198, N2643, N5133);
nand NAND4 (N5792, N5771, N3513, N2031, N3073);
nand NAND3 (N5793, N5775, N5314, N40);
nor NOR3 (N5794, N5792, N1169, N339);
nor NOR2 (N5795, N5779, N2855);
xor XOR2 (N5796, N5780, N5563);
nor NOR3 (N5797, N5790, N1030, N4492);
nand NAND3 (N5798, N5795, N3815, N5548);
nor NOR2 (N5799, N5791, N3047);
not NOT1 (N5800, N5799);
not NOT1 (N5801, N5796);
nor NOR4 (N5802, N5793, N3002, N4556, N4385);
not NOT1 (N5803, N5802);
not NOT1 (N5804, N5800);
nor NOR3 (N5805, N5777, N2730, N3698);
nand NAND3 (N5806, N5787, N2745, N4670);
not NOT1 (N5807, N5805);
and AND3 (N5808, N5798, N2843, N5645);
or OR3 (N5809, N5807, N5362, N574);
and AND4 (N5810, N5789, N2815, N526, N4218);
buf BUF1 (N5811, N5810);
not NOT1 (N5812, N5788);
xor XOR2 (N5813, N5812, N1174);
and AND4 (N5814, N5809, N2834, N5364, N1621);
nand NAND4 (N5815, N5813, N3445, N1359, N4252);
and AND4 (N5816, N5808, N5434, N2512, N485);
nor NOR4 (N5817, N5803, N5369, N5248, N3524);
not NOT1 (N5818, N5801);
nand NAND2 (N5819, N5804, N5585);
not NOT1 (N5820, N5794);
nand NAND3 (N5821, N5797, N5045, N3351);
nand NAND3 (N5822, N5820, N1241, N1282);
xor XOR2 (N5823, N5821, N970);
not NOT1 (N5824, N5816);
not NOT1 (N5825, N5811);
nor NOR2 (N5826, N5815, N4788);
nand NAND2 (N5827, N5814, N1909);
and AND2 (N5828, N5818, N1196);
nand NAND2 (N5829, N5824, N5823);
nor NOR3 (N5830, N3443, N1213, N2925);
and AND2 (N5831, N5827, N4905);
or OR4 (N5832, N5826, N3346, N5441, N2512);
and AND3 (N5833, N5829, N1982, N5155);
xor XOR2 (N5834, N5806, N2899);
and AND2 (N5835, N5828, N4894);
not NOT1 (N5836, N5834);
buf BUF1 (N5837, N5825);
buf BUF1 (N5838, N5817);
nand NAND2 (N5839, N5832, N306);
and AND4 (N5840, N5835, N813, N5565, N4327);
xor XOR2 (N5841, N5838, N3497);
xor XOR2 (N5842, N5840, N3604);
xor XOR2 (N5843, N5839, N1355);
nor NOR2 (N5844, N5819, N1571);
nand NAND4 (N5845, N5822, N4613, N1994, N5538);
buf BUF1 (N5846, N5845);
nand NAND3 (N5847, N5842, N1717, N4409);
xor XOR2 (N5848, N5837, N3999);
nor NOR2 (N5849, N5847, N5345);
buf BUF1 (N5850, N5849);
nor NOR3 (N5851, N5831, N2770, N2587);
xor XOR2 (N5852, N5846, N1924);
nor NOR3 (N5853, N5830, N2215, N2367);
and AND4 (N5854, N5836, N4221, N2487, N4645);
and AND4 (N5855, N5850, N3367, N3263, N4481);
and AND3 (N5856, N5844, N717, N5671);
or OR3 (N5857, N5854, N5676, N4587);
nor NOR2 (N5858, N5853, N2045);
or OR4 (N5859, N5856, N3862, N426, N1120);
nand NAND2 (N5860, N5858, N2431);
or OR4 (N5861, N5841, N921, N4969, N4290);
not NOT1 (N5862, N5848);
not NOT1 (N5863, N5861);
buf BUF1 (N5864, N5863);
nand NAND3 (N5865, N5862, N5308, N947);
and AND3 (N5866, N5843, N4308, N5407);
or OR2 (N5867, N5855, N5865);
nand NAND4 (N5868, N4633, N829, N1833, N4326);
buf BUF1 (N5869, N5857);
nand NAND3 (N5870, N5868, N4506, N1562);
nand NAND2 (N5871, N5869, N1978);
buf BUF1 (N5872, N5866);
xor XOR2 (N5873, N5860, N5676);
and AND2 (N5874, N5864, N5296);
xor XOR2 (N5875, N5871, N4643);
nand NAND2 (N5876, N5873, N4882);
and AND4 (N5877, N5870, N4269, N4339, N3900);
and AND2 (N5878, N5874, N3241);
nand NAND4 (N5879, N5872, N1841, N3300, N79);
not NOT1 (N5880, N5877);
not NOT1 (N5881, N5852);
nand NAND2 (N5882, N5833, N1954);
nand NAND2 (N5883, N5867, N4207);
nor NOR2 (N5884, N5880, N5416);
not NOT1 (N5885, N5851);
buf BUF1 (N5886, N5882);
nor NOR2 (N5887, N5879, N2346);
or OR4 (N5888, N5878, N4542, N243, N4335);
or OR3 (N5889, N5888, N3344, N3059);
and AND3 (N5890, N5881, N1444, N3598);
not NOT1 (N5891, N5876);
xor XOR2 (N5892, N5886, N1292);
and AND2 (N5893, N5890, N5662);
or OR3 (N5894, N5885, N5254, N3843);
and AND4 (N5895, N5883, N4102, N876, N3343);
not NOT1 (N5896, N5859);
nand NAND3 (N5897, N5891, N2471, N3495);
nor NOR4 (N5898, N5896, N5399, N4146, N3844);
or OR4 (N5899, N5884, N336, N3084, N5332);
not NOT1 (N5900, N5875);
not NOT1 (N5901, N5893);
nand NAND3 (N5902, N5901, N181, N5424);
nand NAND3 (N5903, N5900, N3406, N3260);
or OR2 (N5904, N5895, N2027);
nand NAND3 (N5905, N5904, N229, N1398);
xor XOR2 (N5906, N5889, N2825);
buf BUF1 (N5907, N5902);
buf BUF1 (N5908, N5906);
not NOT1 (N5909, N5898);
buf BUF1 (N5910, N5892);
nand NAND4 (N5911, N5903, N868, N967, N1423);
and AND4 (N5912, N5910, N4270, N5688, N1074);
nand NAND4 (N5913, N5905, N4690, N4507, N397);
xor XOR2 (N5914, N5907, N4470);
buf BUF1 (N5915, N5909);
not NOT1 (N5916, N5887);
xor XOR2 (N5917, N5913, N4900);
and AND3 (N5918, N5917, N4143, N2092);
not NOT1 (N5919, N5915);
and AND2 (N5920, N5918, N100);
buf BUF1 (N5921, N5897);
not NOT1 (N5922, N5894);
and AND3 (N5923, N5911, N3910, N4301);
buf BUF1 (N5924, N5916);
buf BUF1 (N5925, N5920);
nor NOR4 (N5926, N5922, N1610, N5573, N4431);
or OR4 (N5927, N5912, N1266, N4571, N4076);
not NOT1 (N5928, N5921);
and AND4 (N5929, N5923, N4394, N3885, N2175);
and AND3 (N5930, N5914, N2398, N4256);
not NOT1 (N5931, N5929);
buf BUF1 (N5932, N5924);
not NOT1 (N5933, N5908);
nand NAND2 (N5934, N5919, N4626);
buf BUF1 (N5935, N5933);
not NOT1 (N5936, N5927);
xor XOR2 (N5937, N5936, N2840);
buf BUF1 (N5938, N5932);
or OR2 (N5939, N5938, N4240);
xor XOR2 (N5940, N5899, N3023);
not NOT1 (N5941, N5939);
nand NAND4 (N5942, N5930, N2944, N4228, N5273);
not NOT1 (N5943, N5942);
xor XOR2 (N5944, N5931, N982);
nand NAND2 (N5945, N5925, N1547);
not NOT1 (N5946, N5926);
nor NOR2 (N5947, N5928, N5278);
or OR3 (N5948, N5937, N3498, N3745);
nor NOR2 (N5949, N5943, N791);
or OR4 (N5950, N5940, N4296, N905, N5543);
and AND2 (N5951, N5934, N2748);
or OR3 (N5952, N5935, N2411, N707);
xor XOR2 (N5953, N5946, N3501);
not NOT1 (N5954, N5947);
nand NAND2 (N5955, N5948, N3341);
or OR2 (N5956, N5950, N1173);
nor NOR3 (N5957, N5953, N161, N4747);
nand NAND2 (N5958, N5956, N3216);
xor XOR2 (N5959, N5958, N2536);
or OR3 (N5960, N5945, N677, N394);
nand NAND4 (N5961, N5949, N5344, N3334, N5694);
buf BUF1 (N5962, N5960);
nand NAND4 (N5963, N5959, N703, N5245, N1402);
nand NAND3 (N5964, N5961, N5048, N177);
or OR4 (N5965, N5954, N1501, N2670, N4542);
and AND4 (N5966, N5963, N4234, N5307, N7);
not NOT1 (N5967, N5965);
xor XOR2 (N5968, N5944, N3029);
nand NAND2 (N5969, N5968, N1882);
nand NAND4 (N5970, N5957, N4680, N5039, N3950);
buf BUF1 (N5971, N5967);
or OR4 (N5972, N5955, N4391, N5246, N3124);
and AND2 (N5973, N5962, N3984);
not NOT1 (N5974, N5941);
not NOT1 (N5975, N5972);
xor XOR2 (N5976, N5971, N1201);
and AND3 (N5977, N5966, N1581, N2612);
xor XOR2 (N5978, N5977, N4637);
nor NOR4 (N5979, N5951, N2987, N2709, N754);
xor XOR2 (N5980, N5979, N5113);
xor XOR2 (N5981, N5978, N5704);
xor XOR2 (N5982, N5969, N1621);
not NOT1 (N5983, N5980);
nand NAND4 (N5984, N5981, N2073, N1983, N1071);
xor XOR2 (N5985, N5973, N1865);
nor NOR4 (N5986, N5970, N3194, N2954, N5128);
xor XOR2 (N5987, N5983, N5900);
or OR3 (N5988, N5985, N1985, N3211);
nand NAND2 (N5989, N5964, N5551);
and AND2 (N5990, N5982, N4136);
buf BUF1 (N5991, N5989);
buf BUF1 (N5992, N5988);
not NOT1 (N5993, N5991);
or OR2 (N5994, N5952, N526);
nand NAND3 (N5995, N5990, N2186, N2007);
or OR4 (N5996, N5976, N3290, N2275, N1615);
and AND4 (N5997, N5993, N2450, N2233, N3965);
not NOT1 (N5998, N5995);
xor XOR2 (N5999, N5994, N5501);
nand NAND3 (N6000, N5984, N153, N5731);
nand NAND2 (N6001, N5996, N5400);
nand NAND4 (N6002, N6000, N2592, N4955, N4117);
buf BUF1 (N6003, N5974);
not NOT1 (N6004, N5975);
or OR4 (N6005, N5997, N3477, N5779, N4475);
nor NOR3 (N6006, N6001, N583, N3755);
xor XOR2 (N6007, N6005, N1773);
nor NOR3 (N6008, N5999, N4079, N399);
buf BUF1 (N6009, N6008);
and AND2 (N6010, N5987, N3201);
or OR2 (N6011, N6007, N1040);
nor NOR2 (N6012, N5986, N326);
buf BUF1 (N6013, N6006);
buf BUF1 (N6014, N6003);
nor NOR2 (N6015, N6002, N3378);
buf BUF1 (N6016, N6012);
buf BUF1 (N6017, N6014);
buf BUF1 (N6018, N6013);
nand NAND3 (N6019, N5992, N5299, N5927);
and AND3 (N6020, N6018, N3939, N681);
nand NAND4 (N6021, N5998, N316, N3746, N3014);
nand NAND2 (N6022, N6019, N76);
not NOT1 (N6023, N6017);
not NOT1 (N6024, N6023);
buf BUF1 (N6025, N6015);
nor NOR2 (N6026, N6020, N1075);
and AND4 (N6027, N6010, N494, N5594, N699);
xor XOR2 (N6028, N6027, N1994);
buf BUF1 (N6029, N6025);
or OR3 (N6030, N6024, N3556, N5994);
not NOT1 (N6031, N6028);
nand NAND3 (N6032, N6031, N5783, N5432);
and AND2 (N6033, N6026, N3580);
xor XOR2 (N6034, N6029, N1805);
buf BUF1 (N6035, N6021);
or OR4 (N6036, N6033, N3604, N2859, N4427);
buf BUF1 (N6037, N6022);
xor XOR2 (N6038, N6016, N3243);
nor NOR2 (N6039, N6037, N962);
xor XOR2 (N6040, N6030, N5180);
and AND4 (N6041, N6038, N3526, N5318, N2564);
nor NOR3 (N6042, N6035, N357, N5961);
buf BUF1 (N6043, N6039);
not NOT1 (N6044, N6011);
buf BUF1 (N6045, N6009);
not NOT1 (N6046, N6034);
or OR4 (N6047, N6042, N1404, N1822, N109);
or OR2 (N6048, N6047, N2625);
buf BUF1 (N6049, N6043);
nor NOR4 (N6050, N6040, N831, N4240, N2790);
nand NAND4 (N6051, N6044, N3444, N2877, N961);
nor NOR3 (N6052, N6046, N4878, N2511);
buf BUF1 (N6053, N6036);
nand NAND3 (N6054, N6050, N2375, N435);
not NOT1 (N6055, N6054);
buf BUF1 (N6056, N6052);
nand NAND2 (N6057, N6056, N884);
or OR4 (N6058, N6057, N4050, N4216, N1050);
buf BUF1 (N6059, N6045);
and AND3 (N6060, N6032, N1408, N3564);
nand NAND4 (N6061, N6058, N354, N4529, N3202);
not NOT1 (N6062, N6061);
nand NAND3 (N6063, N6059, N524, N361);
not NOT1 (N6064, N6051);
nor NOR3 (N6065, N6004, N630, N640);
nand NAND3 (N6066, N6063, N4441, N2143);
not NOT1 (N6067, N6066);
nand NAND2 (N6068, N6049, N1556);
nor NOR3 (N6069, N6055, N1440, N1412);
buf BUF1 (N6070, N6069);
xor XOR2 (N6071, N6053, N1739);
nand NAND2 (N6072, N6060, N1561);
nand NAND2 (N6073, N6062, N2720);
not NOT1 (N6074, N6041);
nand NAND3 (N6075, N6071, N2933, N2966);
nor NOR3 (N6076, N6073, N3848, N2174);
nor NOR4 (N6077, N6075, N1958, N691, N2320);
or OR2 (N6078, N6064, N2140);
buf BUF1 (N6079, N6067);
and AND4 (N6080, N6072, N4410, N3729, N319);
xor XOR2 (N6081, N6070, N3057);
not NOT1 (N6082, N6074);
xor XOR2 (N6083, N6076, N3550);
or OR4 (N6084, N6068, N3430, N163, N4265);
nand NAND2 (N6085, N6079, N3789);
not NOT1 (N6086, N6080);
nand NAND4 (N6087, N6048, N1169, N3276, N4472);
not NOT1 (N6088, N6081);
buf BUF1 (N6089, N6082);
xor XOR2 (N6090, N6085, N26);
xor XOR2 (N6091, N6086, N4253);
nor NOR4 (N6092, N6077, N5477, N4756, N739);
nor NOR3 (N6093, N6087, N162, N4259);
and AND4 (N6094, N6092, N2781, N4339, N5125);
nor NOR3 (N6095, N6093, N2050, N550);
not NOT1 (N6096, N6088);
or OR3 (N6097, N6090, N846, N4662);
or OR4 (N6098, N6091, N978, N979, N1353);
or OR2 (N6099, N6065, N1326);
nor NOR3 (N6100, N6084, N276, N3235);
and AND3 (N6101, N6078, N3624, N1855);
buf BUF1 (N6102, N6098);
not NOT1 (N6103, N6102);
and AND3 (N6104, N6097, N2782, N749);
or OR3 (N6105, N6101, N299, N1486);
not NOT1 (N6106, N6096);
and AND2 (N6107, N6105, N1249);
and AND4 (N6108, N6083, N429, N3723, N315);
or OR2 (N6109, N6095, N5462);
not NOT1 (N6110, N6109);
xor XOR2 (N6111, N6103, N67);
xor XOR2 (N6112, N6094, N5870);
nor NOR2 (N6113, N6104, N6063);
nand NAND4 (N6114, N6112, N4140, N219, N1265);
or OR2 (N6115, N6106, N1859);
buf BUF1 (N6116, N6113);
not NOT1 (N6117, N6099);
and AND2 (N6118, N6100, N1810);
nor NOR4 (N6119, N6107, N62, N4139, N1096);
xor XOR2 (N6120, N6116, N3971);
nand NAND3 (N6121, N6118, N4097, N2879);
nand NAND3 (N6122, N6121, N867, N4561);
nand NAND3 (N6123, N6115, N543, N488);
nor NOR4 (N6124, N6122, N5950, N3243, N4581);
or OR4 (N6125, N6108, N1502, N2944, N4348);
or OR4 (N6126, N6123, N2284, N4681, N5038);
buf BUF1 (N6127, N6126);
not NOT1 (N6128, N6120);
xor XOR2 (N6129, N6127, N3534);
buf BUF1 (N6130, N6129);
or OR3 (N6131, N6125, N2321, N2355);
buf BUF1 (N6132, N6130);
not NOT1 (N6133, N6124);
and AND2 (N6134, N6133, N4270);
and AND3 (N6135, N6134, N2129, N2375);
buf BUF1 (N6136, N6110);
not NOT1 (N6137, N6111);
xor XOR2 (N6138, N6137, N792);
and AND2 (N6139, N6135, N5042);
and AND4 (N6140, N6114, N3619, N2455, N23);
or OR2 (N6141, N6136, N3995);
or OR3 (N6142, N6141, N2824, N2292);
and AND2 (N6143, N6117, N6075);
nand NAND2 (N6144, N6142, N5431);
xor XOR2 (N6145, N6089, N2017);
xor XOR2 (N6146, N6140, N4111);
nand NAND2 (N6147, N6146, N2004);
xor XOR2 (N6148, N6143, N3934);
buf BUF1 (N6149, N6119);
buf BUF1 (N6150, N6148);
buf BUF1 (N6151, N6149);
not NOT1 (N6152, N6151);
or OR3 (N6153, N6144, N1112, N2349);
nor NOR2 (N6154, N6147, N1067);
and AND2 (N6155, N6138, N817);
or OR3 (N6156, N6145, N4409, N5092);
nand NAND3 (N6157, N6132, N3065, N1329);
and AND4 (N6158, N6155, N2175, N3364, N5270);
nand NAND4 (N6159, N6131, N3307, N5638, N4140);
xor XOR2 (N6160, N6152, N5843);
and AND2 (N6161, N6154, N122);
or OR2 (N6162, N6128, N5611);
nor NOR4 (N6163, N6156, N960, N5377, N3948);
nor NOR2 (N6164, N6157, N343);
not NOT1 (N6165, N6160);
and AND4 (N6166, N6139, N3884, N2451, N3975);
or OR3 (N6167, N6163, N3948, N1249);
and AND2 (N6168, N6164, N4085);
nor NOR2 (N6169, N6161, N2720);
or OR2 (N6170, N6162, N2508);
nand NAND4 (N6171, N6168, N671, N6121, N330);
not NOT1 (N6172, N6171);
nand NAND2 (N6173, N6166, N624);
buf BUF1 (N6174, N6158);
nor NOR2 (N6175, N6150, N3119);
nand NAND3 (N6176, N6153, N5807, N3010);
buf BUF1 (N6177, N6174);
not NOT1 (N6178, N6173);
nor NOR2 (N6179, N6176, N4648);
xor XOR2 (N6180, N6175, N4598);
nor NOR3 (N6181, N6179, N319, N1872);
buf BUF1 (N6182, N6159);
not NOT1 (N6183, N6180);
xor XOR2 (N6184, N6183, N276);
xor XOR2 (N6185, N6170, N5712);
or OR4 (N6186, N6169, N482, N1847, N5019);
and AND3 (N6187, N6186, N6098, N726);
not NOT1 (N6188, N6187);
nand NAND2 (N6189, N6184, N4888);
and AND2 (N6190, N6189, N2946);
or OR4 (N6191, N6172, N765, N2809, N883);
xor XOR2 (N6192, N6165, N4962);
or OR2 (N6193, N6182, N609);
and AND4 (N6194, N6181, N2534, N89, N5150);
not NOT1 (N6195, N6192);
not NOT1 (N6196, N6178);
or OR3 (N6197, N6185, N3741, N2723);
nand NAND2 (N6198, N6196, N6109);
not NOT1 (N6199, N6167);
nor NOR2 (N6200, N6195, N3021);
xor XOR2 (N6201, N6191, N3160);
buf BUF1 (N6202, N6198);
nand NAND2 (N6203, N6188, N3798);
buf BUF1 (N6204, N6199);
xor XOR2 (N6205, N6194, N3021);
nor NOR3 (N6206, N6177, N631, N5009);
not NOT1 (N6207, N6206);
nor NOR3 (N6208, N6203, N1067, N4883);
or OR4 (N6209, N6193, N4527, N2801, N5193);
or OR4 (N6210, N6209, N1200, N5775, N4590);
and AND2 (N6211, N6207, N2919);
and AND3 (N6212, N6210, N1575, N1578);
xor XOR2 (N6213, N6205, N1926);
nor NOR3 (N6214, N6208, N2506, N3521);
not NOT1 (N6215, N6214);
xor XOR2 (N6216, N6204, N4178);
or OR2 (N6217, N6190, N5921);
or OR4 (N6218, N6197, N4357, N1154, N3985);
and AND3 (N6219, N6217, N2685, N1057);
not NOT1 (N6220, N6215);
or OR3 (N6221, N6216, N2512, N4364);
not NOT1 (N6222, N6220);
or OR2 (N6223, N6200, N3600);
xor XOR2 (N6224, N6201, N6110);
xor XOR2 (N6225, N6221, N1202);
buf BUF1 (N6226, N6222);
buf BUF1 (N6227, N6226);
not NOT1 (N6228, N6225);
buf BUF1 (N6229, N6224);
or OR2 (N6230, N6223, N1140);
buf BUF1 (N6231, N6229);
nand NAND4 (N6232, N6228, N984, N3196, N2860);
nor NOR4 (N6233, N6202, N3775, N4768, N2862);
not NOT1 (N6234, N6230);
or OR4 (N6235, N6211, N168, N4704, N2897);
not NOT1 (N6236, N6235);
not NOT1 (N6237, N6218);
not NOT1 (N6238, N6237);
buf BUF1 (N6239, N6236);
and AND3 (N6240, N6238, N925, N4438);
and AND2 (N6241, N6232, N342);
xor XOR2 (N6242, N6241, N2140);
and AND3 (N6243, N6234, N1964, N5859);
not NOT1 (N6244, N6227);
and AND3 (N6245, N6233, N1154, N2580);
nor NOR2 (N6246, N6212, N3032);
and AND2 (N6247, N6244, N5171);
and AND2 (N6248, N6246, N1752);
xor XOR2 (N6249, N6219, N5924);
xor XOR2 (N6250, N6249, N3497);
nor NOR2 (N6251, N6239, N5858);
xor XOR2 (N6252, N6240, N1954);
not NOT1 (N6253, N6213);
xor XOR2 (N6254, N6248, N1710);
or OR2 (N6255, N6247, N1062);
nand NAND2 (N6256, N6251, N3328);
not NOT1 (N6257, N6250);
buf BUF1 (N6258, N6254);
and AND2 (N6259, N6231, N2766);
not NOT1 (N6260, N6253);
xor XOR2 (N6261, N6256, N5090);
nor NOR2 (N6262, N6260, N582);
or OR3 (N6263, N6262, N5861, N4720);
nand NAND2 (N6264, N6263, N4766);
nand NAND4 (N6265, N6258, N2155, N5302, N5921);
xor XOR2 (N6266, N6242, N3451);
nand NAND4 (N6267, N6264, N6049, N4927, N1468);
buf BUF1 (N6268, N6257);
not NOT1 (N6269, N6252);
nor NOR4 (N6270, N6266, N18, N4930, N4057);
nor NOR2 (N6271, N6243, N3523);
nand NAND2 (N6272, N6267, N1113);
and AND4 (N6273, N6269, N1143, N1976, N10);
not NOT1 (N6274, N6265);
and AND2 (N6275, N6270, N2585);
xor XOR2 (N6276, N6245, N461);
buf BUF1 (N6277, N6268);
and AND4 (N6278, N6274, N1415, N4757, N6212);
or OR3 (N6279, N6278, N6266, N4298);
not NOT1 (N6280, N6279);
nand NAND4 (N6281, N6273, N4970, N1035, N5652);
or OR3 (N6282, N6259, N5188, N6213);
and AND3 (N6283, N6271, N2440, N811);
xor XOR2 (N6284, N6280, N5542);
xor XOR2 (N6285, N6281, N4209);
or OR2 (N6286, N6272, N4077);
nor NOR3 (N6287, N6283, N2346, N468);
nor NOR2 (N6288, N6276, N1501);
not NOT1 (N6289, N6282);
xor XOR2 (N6290, N6286, N3375);
nand NAND3 (N6291, N6290, N5553, N3588);
or OR2 (N6292, N6255, N3512);
not NOT1 (N6293, N6284);
or OR3 (N6294, N6275, N213, N617);
not NOT1 (N6295, N6288);
nand NAND4 (N6296, N6295, N4799, N5015, N734);
or OR4 (N6297, N6296, N4473, N5663, N5221);
and AND3 (N6298, N6261, N362, N2058);
and AND2 (N6299, N6289, N3991);
xor XOR2 (N6300, N6285, N4136);
and AND3 (N6301, N6292, N961, N3348);
nor NOR3 (N6302, N6301, N6131, N6094);
xor XOR2 (N6303, N6293, N672);
nand NAND4 (N6304, N6298, N1775, N1458, N369);
buf BUF1 (N6305, N6303);
and AND2 (N6306, N6305, N5496);
or OR4 (N6307, N6277, N2156, N4740, N5572);
and AND4 (N6308, N6299, N2295, N3851, N3835);
or OR2 (N6309, N6300, N307);
xor XOR2 (N6310, N6291, N4160);
buf BUF1 (N6311, N6310);
nor NOR3 (N6312, N6311, N5445, N4070);
xor XOR2 (N6313, N6302, N5021);
nor NOR2 (N6314, N6313, N3339);
buf BUF1 (N6315, N6304);
buf BUF1 (N6316, N6309);
xor XOR2 (N6317, N6294, N1562);
nand NAND3 (N6318, N6316, N910, N6246);
nand NAND2 (N6319, N6315, N4222);
xor XOR2 (N6320, N6318, N5980);
xor XOR2 (N6321, N6306, N3760);
buf BUF1 (N6322, N6321);
nand NAND3 (N6323, N6308, N5259, N4244);
or OR2 (N6324, N6287, N3351);
and AND3 (N6325, N6320, N1634, N848);
not NOT1 (N6326, N6314);
and AND3 (N6327, N6319, N4279, N2353);
xor XOR2 (N6328, N6317, N3134);
not NOT1 (N6329, N6327);
and AND3 (N6330, N6328, N4284, N3323);
not NOT1 (N6331, N6307);
nand NAND4 (N6332, N6325, N903, N325, N2879);
buf BUF1 (N6333, N6332);
and AND4 (N6334, N6312, N4356, N81, N5306);
nor NOR2 (N6335, N6323, N1274);
not NOT1 (N6336, N6331);
buf BUF1 (N6337, N6329);
nor NOR2 (N6338, N6326, N4887);
xor XOR2 (N6339, N6322, N1252);
nand NAND2 (N6340, N6333, N3569);
buf BUF1 (N6341, N6335);
nor NOR2 (N6342, N6297, N1253);
buf BUF1 (N6343, N6330);
not NOT1 (N6344, N6337);
nor NOR2 (N6345, N6338, N5817);
not NOT1 (N6346, N6334);
and AND2 (N6347, N6343, N3185);
buf BUF1 (N6348, N6336);
buf BUF1 (N6349, N6341);
nor NOR2 (N6350, N6340, N2516);
buf BUF1 (N6351, N6349);
and AND4 (N6352, N6350, N5163, N4044, N1086);
nand NAND2 (N6353, N6347, N4731);
nor NOR3 (N6354, N6344, N3581, N4194);
nor NOR3 (N6355, N6345, N2894, N1088);
buf BUF1 (N6356, N6339);
nor NOR4 (N6357, N6351, N818, N3597, N6291);
not NOT1 (N6358, N6356);
nor NOR2 (N6359, N6324, N6173);
or OR2 (N6360, N6357, N2219);
xor XOR2 (N6361, N6346, N761);
nor NOR4 (N6362, N6348, N2049, N3972, N1291);
buf BUF1 (N6363, N6361);
buf BUF1 (N6364, N6360);
nand NAND3 (N6365, N6362, N2255, N3395);
not NOT1 (N6366, N6352);
or OR4 (N6367, N6364, N2984, N1785, N1774);
buf BUF1 (N6368, N6365);
nand NAND3 (N6369, N6367, N2092, N3140);
not NOT1 (N6370, N6353);
not NOT1 (N6371, N6354);
or OR4 (N6372, N6370, N92, N1620, N3867);
and AND2 (N6373, N6363, N1048);
nand NAND2 (N6374, N6372, N665);
buf BUF1 (N6375, N6355);
or OR2 (N6376, N6342, N5173);
not NOT1 (N6377, N6375);
or OR4 (N6378, N6359, N566, N4167, N2289);
nand NAND2 (N6379, N6366, N2005);
nor NOR2 (N6380, N6368, N4210);
nor NOR2 (N6381, N6376, N6121);
or OR2 (N6382, N6373, N1246);
xor XOR2 (N6383, N6378, N1002);
xor XOR2 (N6384, N6369, N3633);
nand NAND4 (N6385, N6380, N156, N5559, N3255);
or OR3 (N6386, N6379, N3389, N3173);
nand NAND4 (N6387, N6381, N5880, N2654, N2632);
nand NAND3 (N6388, N6371, N3392, N5855);
nor NOR2 (N6389, N6385, N6084);
nor NOR4 (N6390, N6387, N5208, N1274, N1404);
nor NOR4 (N6391, N6386, N1571, N1343, N770);
not NOT1 (N6392, N6382);
or OR3 (N6393, N6389, N4620, N795);
nor NOR4 (N6394, N6392, N5620, N3242, N5117);
not NOT1 (N6395, N6388);
nor NOR4 (N6396, N6395, N6141, N3833, N3426);
or OR3 (N6397, N6393, N5144, N5726);
not NOT1 (N6398, N6384);
xor XOR2 (N6399, N6391, N5231);
xor XOR2 (N6400, N6390, N2840);
buf BUF1 (N6401, N6396);
nor NOR4 (N6402, N6377, N3557, N5864, N2882);
or OR3 (N6403, N6401, N3907, N5534);
buf BUF1 (N6404, N6358);
xor XOR2 (N6405, N6404, N4301);
nand NAND3 (N6406, N6397, N5733, N3792);
nand NAND3 (N6407, N6405, N1055, N542);
not NOT1 (N6408, N6402);
nand NAND2 (N6409, N6407, N4030);
nand NAND3 (N6410, N6403, N4355, N939);
not NOT1 (N6411, N6383);
buf BUF1 (N6412, N6406);
buf BUF1 (N6413, N6410);
not NOT1 (N6414, N6398);
buf BUF1 (N6415, N6399);
not NOT1 (N6416, N6413);
nand NAND2 (N6417, N6374, N5755);
buf BUF1 (N6418, N6417);
or OR3 (N6419, N6416, N3402, N2435);
and AND3 (N6420, N6411, N5614, N3086);
or OR3 (N6421, N6394, N36, N4787);
buf BUF1 (N6422, N6409);
and AND3 (N6423, N6412, N4929, N5415);
xor XOR2 (N6424, N6414, N3568);
and AND2 (N6425, N6400, N4757);
buf BUF1 (N6426, N6415);
xor XOR2 (N6427, N6424, N4952);
nor NOR4 (N6428, N6420, N1280, N1805, N274);
xor XOR2 (N6429, N6408, N1344);
buf BUF1 (N6430, N6428);
nor NOR4 (N6431, N6425, N2893, N2756, N1741);
or OR4 (N6432, N6418, N1691, N4560, N4982);
xor XOR2 (N6433, N6430, N5046);
and AND4 (N6434, N6429, N3615, N5581, N908);
nand NAND4 (N6435, N6432, N2477, N4968, N5240);
or OR4 (N6436, N6421, N2154, N3679, N1944);
buf BUF1 (N6437, N6426);
xor XOR2 (N6438, N6423, N3262);
and AND4 (N6439, N6419, N4074, N897, N228);
buf BUF1 (N6440, N6436);
buf BUF1 (N6441, N6438);
not NOT1 (N6442, N6441);
buf BUF1 (N6443, N6431);
buf BUF1 (N6444, N6437);
xor XOR2 (N6445, N6435, N718);
not NOT1 (N6446, N6439);
or OR2 (N6447, N6446, N1523);
xor XOR2 (N6448, N6427, N4158);
nand NAND2 (N6449, N6447, N211);
xor XOR2 (N6450, N6449, N4461);
xor XOR2 (N6451, N6442, N3123);
or OR3 (N6452, N6443, N4564, N5277);
nand NAND4 (N6453, N6433, N466, N5735, N5399);
or OR4 (N6454, N6450, N4136, N2146, N4966);
buf BUF1 (N6455, N6454);
or OR2 (N6456, N6445, N391);
buf BUF1 (N6457, N6448);
buf BUF1 (N6458, N6453);
nor NOR2 (N6459, N6434, N1815);
nor NOR3 (N6460, N6451, N903, N3387);
xor XOR2 (N6461, N6460, N3966);
or OR4 (N6462, N6444, N3999, N4063, N4718);
xor XOR2 (N6463, N6462, N2203);
nand NAND2 (N6464, N6458, N6122);
nand NAND4 (N6465, N6459, N3181, N665, N4295);
buf BUF1 (N6466, N6465);
xor XOR2 (N6467, N6440, N4172);
nor NOR3 (N6468, N6456, N1059, N2675);
not NOT1 (N6469, N6468);
or OR4 (N6470, N6452, N2624, N3057, N592);
xor XOR2 (N6471, N6470, N4510);
buf BUF1 (N6472, N6464);
nor NOR2 (N6473, N6469, N5286);
nor NOR2 (N6474, N6463, N5443);
nor NOR2 (N6475, N6422, N560);
nand NAND4 (N6476, N6461, N6385, N4762, N1656);
or OR2 (N6477, N6457, N6236);
nand NAND2 (N6478, N6473, N55);
nor NOR4 (N6479, N6467, N3702, N160, N2388);
nor NOR2 (N6480, N6475, N2292);
nor NOR2 (N6481, N6478, N6324);
nand NAND3 (N6482, N6455, N5042, N2132);
buf BUF1 (N6483, N6472);
or OR3 (N6484, N6480, N5228, N4875);
not NOT1 (N6485, N6477);
nand NAND3 (N6486, N6466, N530, N1416);
and AND4 (N6487, N6471, N4226, N4375, N5661);
or OR3 (N6488, N6482, N2930, N3268);
nand NAND4 (N6489, N6474, N6267, N1347, N315);
nand NAND2 (N6490, N6483, N4499);
not NOT1 (N6491, N6476);
nor NOR2 (N6492, N6481, N3754);
nand NAND4 (N6493, N6486, N5589, N2301, N4469);
xor XOR2 (N6494, N6491, N1791);
or OR4 (N6495, N6479, N599, N3201, N3086);
not NOT1 (N6496, N6493);
nand NAND3 (N6497, N6488, N5394, N5584);
nand NAND4 (N6498, N6489, N3122, N1183, N1196);
or OR3 (N6499, N6495, N1333, N1565);
nor NOR4 (N6500, N6498, N335, N3655, N3007);
nand NAND2 (N6501, N6484, N1059);
buf BUF1 (N6502, N6499);
and AND4 (N6503, N6485, N3798, N402, N4625);
not NOT1 (N6504, N6502);
not NOT1 (N6505, N6503);
nand NAND2 (N6506, N6497, N445);
and AND3 (N6507, N6506, N6439, N3345);
or OR3 (N6508, N6500, N4760, N5216);
buf BUF1 (N6509, N6494);
nand NAND4 (N6510, N6505, N2647, N5628, N4985);
xor XOR2 (N6511, N6496, N1157);
and AND2 (N6512, N6504, N1406);
nor NOR3 (N6513, N6508, N4189, N939);
buf BUF1 (N6514, N6510);
or OR4 (N6515, N6511, N4948, N2227, N4067);
nand NAND4 (N6516, N6514, N1701, N6309, N6226);
buf BUF1 (N6517, N6487);
and AND4 (N6518, N6515, N3520, N1044, N2779);
nor NOR2 (N6519, N6509, N2599);
nand NAND4 (N6520, N6490, N2163, N3628, N5733);
or OR2 (N6521, N6520, N3971);
not NOT1 (N6522, N6517);
nor NOR2 (N6523, N6512, N6359);
buf BUF1 (N6524, N6516);
and AND4 (N6525, N6524, N314, N5478, N4009);
or OR2 (N6526, N6519, N3181);
nor NOR2 (N6527, N6518, N4754);
and AND2 (N6528, N6527, N4207);
not NOT1 (N6529, N6501);
or OR3 (N6530, N6513, N4052, N2663);
and AND3 (N6531, N6521, N1034, N1466);
nand NAND4 (N6532, N6492, N5670, N91, N6202);
not NOT1 (N6533, N6531);
nor NOR4 (N6534, N6523, N2233, N5384, N4008);
or OR2 (N6535, N6532, N2566);
nor NOR2 (N6536, N6525, N103);
not NOT1 (N6537, N6533);
or OR4 (N6538, N6534, N6278, N1379, N2870);
xor XOR2 (N6539, N6536, N178);
nor NOR2 (N6540, N6522, N6174);
buf BUF1 (N6541, N6526);
or OR2 (N6542, N6538, N2326);
xor XOR2 (N6543, N6537, N706);
and AND4 (N6544, N6528, N975, N2849, N3469);
and AND4 (N6545, N6530, N4459, N4803, N2487);
buf BUF1 (N6546, N6545);
nand NAND2 (N6547, N6529, N1197);
or OR4 (N6548, N6543, N562, N4739, N1167);
nand NAND3 (N6549, N6547, N5847, N3371);
xor XOR2 (N6550, N6507, N1266);
nor NOR3 (N6551, N6539, N5691, N1867);
xor XOR2 (N6552, N6548, N5442);
nor NOR2 (N6553, N6551, N1853);
not NOT1 (N6554, N6549);
and AND4 (N6555, N6546, N4927, N5650, N4341);
not NOT1 (N6556, N6541);
and AND2 (N6557, N6535, N1328);
or OR2 (N6558, N6540, N883);
nand NAND3 (N6559, N6556, N4899, N5113);
buf BUF1 (N6560, N6552);
nor NOR2 (N6561, N6544, N375);
nor NOR4 (N6562, N6550, N1358, N396, N5275);
not NOT1 (N6563, N6562);
xor XOR2 (N6564, N6557, N65);
not NOT1 (N6565, N6553);
nor NOR3 (N6566, N6554, N1921, N2715);
xor XOR2 (N6567, N6566, N6062);
nand NAND4 (N6568, N6555, N4379, N2293, N5543);
xor XOR2 (N6569, N6561, N5523);
nor NOR2 (N6570, N6568, N467);
xor XOR2 (N6571, N6542, N4325);
buf BUF1 (N6572, N6559);
xor XOR2 (N6573, N6569, N1477);
nor NOR2 (N6574, N6560, N4296);
nor NOR3 (N6575, N6563, N6408, N3467);
buf BUF1 (N6576, N6570);
not NOT1 (N6577, N6571);
nor NOR3 (N6578, N6576, N1076, N6282);
and AND2 (N6579, N6558, N42);
and AND3 (N6580, N6575, N1423, N6371);
not NOT1 (N6581, N6572);
xor XOR2 (N6582, N6577, N3328);
buf BUF1 (N6583, N6582);
buf BUF1 (N6584, N6573);
nor NOR2 (N6585, N6578, N6272);
and AND2 (N6586, N6581, N442);
not NOT1 (N6587, N6584);
nor NOR3 (N6588, N6583, N2026, N414);
buf BUF1 (N6589, N6567);
nand NAND2 (N6590, N6574, N64);
buf BUF1 (N6591, N6587);
or OR3 (N6592, N6565, N4875, N4868);
nand NAND4 (N6593, N6591, N875, N4575, N5440);
and AND3 (N6594, N6593, N5889, N4801);
and AND4 (N6595, N6585, N4742, N3000, N3862);
nor NOR4 (N6596, N6589, N1492, N97, N6185);
and AND2 (N6597, N6596, N3788);
nor NOR4 (N6598, N6580, N5160, N4894, N3958);
and AND2 (N6599, N6590, N4080);
nand NAND3 (N6600, N6564, N5109, N5009);
xor XOR2 (N6601, N6600, N446);
xor XOR2 (N6602, N6594, N4436);
nand NAND2 (N6603, N6597, N1167);
or OR3 (N6604, N6599, N3504, N2429);
or OR3 (N6605, N6598, N1252, N4055);
xor XOR2 (N6606, N6586, N5352);
nand NAND3 (N6607, N6592, N2422, N6274);
buf BUF1 (N6608, N6601);
or OR2 (N6609, N6608, N267);
nand NAND4 (N6610, N6605, N204, N1505, N6414);
not NOT1 (N6611, N6579);
nor NOR3 (N6612, N6588, N1971, N1683);
not NOT1 (N6613, N6604);
not NOT1 (N6614, N6595);
nand NAND2 (N6615, N6609, N6363);
and AND3 (N6616, N6607, N1143, N6417);
xor XOR2 (N6617, N6614, N3295);
nand NAND3 (N6618, N6610, N5635, N1284);
nand NAND2 (N6619, N6617, N4368);
xor XOR2 (N6620, N6619, N1356);
nor NOR4 (N6621, N6602, N806, N1956, N3323);
nor NOR4 (N6622, N6612, N1188, N5587, N3654);
nand NAND4 (N6623, N6621, N3305, N3870, N5669);
xor XOR2 (N6624, N6615, N985);
nor NOR4 (N6625, N6623, N6221, N2294, N4047);
buf BUF1 (N6626, N6618);
not NOT1 (N6627, N6626);
not NOT1 (N6628, N6616);
nor NOR4 (N6629, N6620, N146, N1841, N4523);
nand NAND3 (N6630, N6611, N5775, N1962);
and AND4 (N6631, N6630, N959, N227, N4791);
nand NAND3 (N6632, N6613, N1748, N4753);
nor NOR3 (N6633, N6603, N1916, N4221);
or OR4 (N6634, N6632, N2477, N1482, N2915);
nor NOR4 (N6635, N6624, N4469, N4041, N4309);
or OR4 (N6636, N6606, N4706, N1202, N4876);
nor NOR4 (N6637, N6634, N3948, N6012, N5904);
nand NAND3 (N6638, N6625, N1226, N4685);
nor NOR3 (N6639, N6638, N2881, N66);
not NOT1 (N6640, N6635);
not NOT1 (N6641, N6628);
and AND3 (N6642, N6627, N2615, N1110);
nor NOR4 (N6643, N6633, N6221, N2402, N3488);
or OR4 (N6644, N6643, N665, N1681, N6092);
buf BUF1 (N6645, N6640);
not NOT1 (N6646, N6636);
nand NAND4 (N6647, N6645, N836, N1386, N1754);
and AND3 (N6648, N6637, N1652, N2901);
xor XOR2 (N6649, N6629, N2936);
nand NAND4 (N6650, N6631, N6196, N4899, N5709);
nor NOR2 (N6651, N6646, N1904);
buf BUF1 (N6652, N6641);
or OR2 (N6653, N6642, N742);
and AND4 (N6654, N6622, N4959, N6052, N2229);
not NOT1 (N6655, N6649);
buf BUF1 (N6656, N6639);
and AND2 (N6657, N6653, N3363);
not NOT1 (N6658, N6644);
xor XOR2 (N6659, N6657, N5997);
not NOT1 (N6660, N6656);
nor NOR3 (N6661, N6652, N4022, N3108);
and AND2 (N6662, N6647, N5746);
buf BUF1 (N6663, N6655);
nor NOR2 (N6664, N6658, N3189);
nand NAND4 (N6665, N6660, N5770, N3554, N5540);
buf BUF1 (N6666, N6650);
nor NOR3 (N6667, N6659, N2192, N5586);
nor NOR4 (N6668, N6665, N2263, N1472, N51);
or OR4 (N6669, N6664, N2673, N74, N3015);
and AND3 (N6670, N6661, N5395, N407);
nand NAND3 (N6671, N6663, N5458, N4925);
or OR4 (N6672, N6662, N3478, N2683, N2884);
nor NOR2 (N6673, N6648, N6188);
nor NOR3 (N6674, N6672, N36, N2238);
not NOT1 (N6675, N6673);
or OR3 (N6676, N6670, N1879, N1730);
not NOT1 (N6677, N6654);
buf BUF1 (N6678, N6668);
nor NOR3 (N6679, N6669, N1279, N4021);
buf BUF1 (N6680, N6666);
or OR3 (N6681, N6677, N1171, N3512);
buf BUF1 (N6682, N6671);
or OR2 (N6683, N6676, N5281);
xor XOR2 (N6684, N6675, N1947);
nor NOR3 (N6685, N6679, N2967, N316);
not NOT1 (N6686, N6674);
buf BUF1 (N6687, N6685);
nand NAND4 (N6688, N6667, N2573, N6277, N382);
nor NOR2 (N6689, N6680, N3948);
nor NOR4 (N6690, N6681, N786, N3789, N2305);
buf BUF1 (N6691, N6684);
or OR2 (N6692, N6683, N3434);
nor NOR2 (N6693, N6688, N2279);
and AND4 (N6694, N6689, N4925, N6650, N5621);
buf BUF1 (N6695, N6682);
xor XOR2 (N6696, N6651, N3111);
buf BUF1 (N6697, N6692);
xor XOR2 (N6698, N6678, N1052);
and AND3 (N6699, N6694, N3063, N2207);
xor XOR2 (N6700, N6695, N4896);
or OR4 (N6701, N6691, N3271, N4808, N5778);
nand NAND2 (N6702, N6690, N1514);
not NOT1 (N6703, N6693);
buf BUF1 (N6704, N6696);
buf BUF1 (N6705, N6698);
or OR2 (N6706, N6704, N2236);
or OR3 (N6707, N6702, N4117, N2635);
and AND3 (N6708, N6705, N1426, N3890);
and AND2 (N6709, N6701, N3307);
not NOT1 (N6710, N6706);
or OR4 (N6711, N6710, N337, N473, N734);
and AND2 (N6712, N6703, N4109);
buf BUF1 (N6713, N6687);
and AND2 (N6714, N6707, N637);
not NOT1 (N6715, N6711);
and AND4 (N6716, N6700, N3460, N3524, N1254);
buf BUF1 (N6717, N6714);
and AND3 (N6718, N6712, N3055, N5823);
xor XOR2 (N6719, N6708, N6173);
nand NAND4 (N6720, N6718, N6431, N2418, N6687);
not NOT1 (N6721, N6697);
or OR4 (N6722, N6699, N2611, N119, N5520);
xor XOR2 (N6723, N6719, N6703);
and AND3 (N6724, N6723, N6133, N2894);
nor NOR3 (N6725, N6709, N5834, N3313);
or OR4 (N6726, N6716, N2832, N1687, N73);
nand NAND2 (N6727, N6715, N5120);
or OR2 (N6728, N6720, N970);
or OR3 (N6729, N6717, N536, N3875);
or OR4 (N6730, N6729, N234, N6408, N6031);
xor XOR2 (N6731, N6726, N5478);
and AND3 (N6732, N6713, N1055, N933);
or OR3 (N6733, N6731, N6109, N3369);
not NOT1 (N6734, N6733);
xor XOR2 (N6735, N6686, N3144);
or OR2 (N6736, N6724, N6051);
nand NAND3 (N6737, N6728, N2383, N3537);
and AND4 (N6738, N6737, N2687, N4456, N2566);
and AND3 (N6739, N6722, N4733, N5397);
and AND4 (N6740, N6721, N6480, N4615, N6644);
xor XOR2 (N6741, N6736, N3893);
or OR2 (N6742, N6727, N5790);
not NOT1 (N6743, N6730);
nand NAND4 (N6744, N6738, N3054, N4010, N2279);
and AND3 (N6745, N6742, N5482, N1932);
xor XOR2 (N6746, N6735, N4464);
buf BUF1 (N6747, N6732);
or OR2 (N6748, N6734, N2573);
xor XOR2 (N6749, N6725, N6448);
xor XOR2 (N6750, N6743, N3811);
or OR2 (N6751, N6745, N6551);
nand NAND3 (N6752, N6746, N4038, N2738);
not NOT1 (N6753, N6752);
buf BUF1 (N6754, N6741);
xor XOR2 (N6755, N6748, N1610);
xor XOR2 (N6756, N6747, N5891);
not NOT1 (N6757, N6754);
or OR4 (N6758, N6749, N4040, N5825, N1420);
nor NOR2 (N6759, N6758, N1285);
not NOT1 (N6760, N6756);
nand NAND4 (N6761, N6759, N6048, N5067, N2689);
nor NOR4 (N6762, N6750, N5166, N760, N6252);
and AND4 (N6763, N6762, N5850, N5051, N1788);
or OR3 (N6764, N6763, N4679, N3488);
nor NOR2 (N6765, N6753, N5131);
buf BUF1 (N6766, N6740);
and AND3 (N6767, N6739, N4980, N2793);
xor XOR2 (N6768, N6760, N6153);
not NOT1 (N6769, N6744);
and AND2 (N6770, N6767, N2733);
nand NAND4 (N6771, N6761, N6160, N872, N3513);
xor XOR2 (N6772, N6771, N2292);
xor XOR2 (N6773, N6772, N1432);
and AND4 (N6774, N6765, N5565, N6511, N2666);
xor XOR2 (N6775, N6751, N4308);
buf BUF1 (N6776, N6757);
buf BUF1 (N6777, N6755);
or OR4 (N6778, N6775, N129, N357, N2645);
buf BUF1 (N6779, N6769);
and AND4 (N6780, N6776, N6078, N4292, N6724);
or OR3 (N6781, N6777, N3467, N5368);
nand NAND3 (N6782, N6781, N329, N127);
nor NOR3 (N6783, N6774, N3403, N1592);
or OR4 (N6784, N6764, N4153, N4113, N644);
xor XOR2 (N6785, N6770, N1852);
nand NAND2 (N6786, N6778, N6138);
xor XOR2 (N6787, N6784, N2317);
nand NAND3 (N6788, N6779, N1048, N4675);
nand NAND3 (N6789, N6768, N49, N773);
and AND3 (N6790, N6785, N1286, N5129);
nor NOR2 (N6791, N6789, N3281);
xor XOR2 (N6792, N6790, N4181);
or OR3 (N6793, N6782, N378, N2027);
and AND3 (N6794, N6788, N4103, N3604);
not NOT1 (N6795, N6773);
not NOT1 (N6796, N6766);
or OR4 (N6797, N6791, N1739, N5327, N1371);
not NOT1 (N6798, N6780);
or OR4 (N6799, N6792, N3852, N4985, N1536);
xor XOR2 (N6800, N6793, N6177);
and AND4 (N6801, N6787, N4415, N2791, N993);
buf BUF1 (N6802, N6796);
nor NOR2 (N6803, N6794, N2725);
nand NAND4 (N6804, N6786, N4527, N3738, N487);
xor XOR2 (N6805, N6803, N4844);
nand NAND3 (N6806, N6804, N6218, N4057);
xor XOR2 (N6807, N6800, N5382);
or OR2 (N6808, N6783, N1640);
nand NAND2 (N6809, N6797, N6005);
or OR4 (N6810, N6798, N6020, N6246, N4923);
nand NAND3 (N6811, N6795, N2763, N2735);
or OR2 (N6812, N6807, N4066);
xor XOR2 (N6813, N6810, N4874);
and AND3 (N6814, N6812, N2405, N3022);
and AND4 (N6815, N6813, N5400, N2683, N2006);
or OR3 (N6816, N6801, N6784, N3639);
and AND3 (N6817, N6802, N1683, N2364);
nor NOR4 (N6818, N6817, N5813, N1814, N1541);
nand NAND3 (N6819, N6806, N5819, N3592);
nand NAND2 (N6820, N6799, N5951);
buf BUF1 (N6821, N6820);
nor NOR4 (N6822, N6805, N1293, N5538, N4737);
nand NAND2 (N6823, N6821, N387);
xor XOR2 (N6824, N6809, N2175);
not NOT1 (N6825, N6823);
not NOT1 (N6826, N6814);
nand NAND2 (N6827, N6819, N6790);
nor NOR3 (N6828, N6824, N4105, N3795);
xor XOR2 (N6829, N6822, N5048);
not NOT1 (N6830, N6827);
not NOT1 (N6831, N6808);
nand NAND2 (N6832, N6831, N3018);
or OR3 (N6833, N6818, N69, N2161);
not NOT1 (N6834, N6832);
or OR4 (N6835, N6833, N5947, N896, N4532);
and AND2 (N6836, N6830, N2339);
nor NOR4 (N6837, N6825, N4658, N6528, N5349);
not NOT1 (N6838, N6829);
not NOT1 (N6839, N6811);
nand NAND3 (N6840, N6838, N6083, N1957);
nor NOR4 (N6841, N6840, N3895, N1863, N1597);
xor XOR2 (N6842, N6839, N2815);
and AND2 (N6843, N6837, N1110);
nor NOR4 (N6844, N6842, N4766, N6698, N5740);
xor XOR2 (N6845, N6835, N6579);
buf BUF1 (N6846, N6815);
not NOT1 (N6847, N6828);
and AND4 (N6848, N6836, N1139, N3219, N3613);
buf BUF1 (N6849, N6826);
nor NOR2 (N6850, N6845, N6111);
nand NAND3 (N6851, N6848, N4305, N951);
xor XOR2 (N6852, N6849, N98);
or OR2 (N6853, N6846, N2050);
nand NAND2 (N6854, N6841, N5512);
nand NAND4 (N6855, N6853, N6349, N3680, N3939);
not NOT1 (N6856, N6843);
or OR4 (N6857, N6847, N3370, N810, N5112);
nor NOR4 (N6858, N6856, N2821, N4402, N3102);
buf BUF1 (N6859, N6858);
or OR4 (N6860, N6851, N1745, N1515, N3585);
or OR3 (N6861, N6855, N2412, N6834);
buf BUF1 (N6862, N601);
nand NAND4 (N6863, N6852, N1898, N1704, N4327);
xor XOR2 (N6864, N6844, N6436);
or OR4 (N6865, N6859, N316, N3617, N6733);
nand NAND4 (N6866, N6816, N126, N5323, N1362);
nor NOR3 (N6867, N6866, N5896, N1982);
nor NOR4 (N6868, N6850, N4813, N2086, N2867);
buf BUF1 (N6869, N6865);
nand NAND2 (N6870, N6861, N6691);
nand NAND3 (N6871, N6862, N2165, N3657);
nand NAND2 (N6872, N6871, N5644);
nor NOR2 (N6873, N6854, N889);
and AND2 (N6874, N6860, N6132);
not NOT1 (N6875, N6874);
and AND3 (N6876, N6869, N5379, N1594);
nand NAND2 (N6877, N6875, N691);
and AND3 (N6878, N6863, N5628, N4524);
xor XOR2 (N6879, N6868, N6574);
nor NOR2 (N6880, N6857, N3749);
xor XOR2 (N6881, N6880, N4551);
not NOT1 (N6882, N6873);
nor NOR2 (N6883, N6867, N4233);
or OR3 (N6884, N6878, N318, N3894);
xor XOR2 (N6885, N6876, N5220);
nand NAND2 (N6886, N6881, N6499);
not NOT1 (N6887, N6872);
nand NAND2 (N6888, N6882, N496);
buf BUF1 (N6889, N6886);
buf BUF1 (N6890, N6870);
not NOT1 (N6891, N6877);
and AND3 (N6892, N6888, N3028, N3074);
or OR4 (N6893, N6889, N1388, N1434, N5890);
nand NAND2 (N6894, N6887, N261);
nor NOR3 (N6895, N6884, N6395, N2025);
and AND4 (N6896, N6894, N6623, N4772, N2210);
not NOT1 (N6897, N6885);
and AND3 (N6898, N6897, N4330, N3045);
xor XOR2 (N6899, N6892, N6538);
xor XOR2 (N6900, N6879, N5718);
and AND2 (N6901, N6890, N4985);
xor XOR2 (N6902, N6883, N3089);
nor NOR3 (N6903, N6895, N6267, N4376);
or OR3 (N6904, N6893, N80, N2542);
and AND2 (N6905, N6901, N1650);
nand NAND4 (N6906, N6902, N4201, N5657, N5372);
or OR3 (N6907, N6891, N6362, N138);
and AND3 (N6908, N6906, N300, N679);
xor XOR2 (N6909, N6898, N4877);
and AND3 (N6910, N6907, N3575, N6271);
xor XOR2 (N6911, N6904, N6844);
and AND4 (N6912, N6910, N403, N4676, N6304);
or OR2 (N6913, N6864, N6643);
buf BUF1 (N6914, N6912);
not NOT1 (N6915, N6903);
or OR4 (N6916, N6899, N1927, N6168, N556);
buf BUF1 (N6917, N6913);
nor NOR3 (N6918, N6909, N1503, N4404);
not NOT1 (N6919, N6905);
xor XOR2 (N6920, N6911, N3334);
not NOT1 (N6921, N6900);
nor NOR4 (N6922, N6914, N2651, N4651, N420);
nor NOR3 (N6923, N6916, N2437, N4739);
xor XOR2 (N6924, N6915, N1975);
or OR3 (N6925, N6917, N5962, N5305);
or OR3 (N6926, N6920, N1162, N3859);
nor NOR2 (N6927, N6926, N3004);
nand NAND2 (N6928, N6923, N5689);
nor NOR4 (N6929, N6928, N3738, N6828, N564);
nand NAND3 (N6930, N6919, N1452, N3927);
nor NOR2 (N6931, N6908, N2599);
not NOT1 (N6932, N6931);
nor NOR2 (N6933, N6896, N4231);
or OR3 (N6934, N6918, N2530, N2918);
not NOT1 (N6935, N6927);
not NOT1 (N6936, N6934);
nor NOR2 (N6937, N6929, N1688);
xor XOR2 (N6938, N6935, N1224);
not NOT1 (N6939, N6937);
and AND2 (N6940, N6932, N5784);
nor NOR2 (N6941, N6924, N3952);
xor XOR2 (N6942, N6941, N509);
nor NOR4 (N6943, N6939, N3832, N2347, N3971);
not NOT1 (N6944, N6930);
nor NOR2 (N6945, N6933, N3250);
or OR2 (N6946, N6936, N944);
buf BUF1 (N6947, N6946);
and AND2 (N6948, N6945, N4290);
xor XOR2 (N6949, N6942, N1684);
nor NOR4 (N6950, N6943, N6425, N1594, N6829);
not NOT1 (N6951, N6949);
nand NAND2 (N6952, N6951, N3198);
nor NOR4 (N6953, N6925, N1869, N4211, N5385);
buf BUF1 (N6954, N6952);
nand NAND2 (N6955, N6947, N5198);
buf BUF1 (N6956, N6953);
nand NAND4 (N6957, N6954, N5791, N5173, N5517);
nor NOR4 (N6958, N6944, N4288, N6379, N4891);
xor XOR2 (N6959, N6957, N4696);
xor XOR2 (N6960, N6955, N2400);
and AND2 (N6961, N6950, N3866);
not NOT1 (N6962, N6948);
or OR4 (N6963, N6962, N1512, N6949, N2351);
xor XOR2 (N6964, N6961, N3913);
nand NAND4 (N6965, N6959, N5938, N3718, N4635);
buf BUF1 (N6966, N6964);
xor XOR2 (N6967, N6966, N5595);
nand NAND2 (N6968, N6940, N2253);
xor XOR2 (N6969, N6921, N367);
buf BUF1 (N6970, N6958);
and AND2 (N6971, N6968, N343);
xor XOR2 (N6972, N6965, N1651);
xor XOR2 (N6973, N6967, N2719);
nor NOR3 (N6974, N6970, N2299, N5675);
buf BUF1 (N6975, N6922);
buf BUF1 (N6976, N6956);
buf BUF1 (N6977, N6974);
buf BUF1 (N6978, N6975);
not NOT1 (N6979, N6971);
nand NAND4 (N6980, N6976, N4813, N3179, N1980);
not NOT1 (N6981, N6960);
or OR3 (N6982, N6963, N6093, N5186);
xor XOR2 (N6983, N6969, N4790);
buf BUF1 (N6984, N6982);
or OR2 (N6985, N6981, N5895);
not NOT1 (N6986, N6984);
and AND3 (N6987, N6985, N3131, N4439);
buf BUF1 (N6988, N6987);
or OR4 (N6989, N6977, N2079, N54, N3977);
nor NOR4 (N6990, N6979, N2207, N6129, N6386);
nor NOR3 (N6991, N6972, N2509, N6301);
not NOT1 (N6992, N6938);
buf BUF1 (N6993, N6989);
not NOT1 (N6994, N6993);
buf BUF1 (N6995, N6978);
xor XOR2 (N6996, N6992, N2714);
and AND2 (N6997, N6990, N6816);
and AND4 (N6998, N6997, N5513, N2060, N5767);
xor XOR2 (N6999, N6998, N5157);
nand NAND4 (N7000, N6986, N5516, N3619, N4684);
buf BUF1 (N7001, N7000);
not NOT1 (N7002, N6996);
not NOT1 (N7003, N6973);
buf BUF1 (N7004, N7002);
buf BUF1 (N7005, N6995);
and AND3 (N7006, N7004, N1401, N3203);
nor NOR3 (N7007, N6999, N3900, N2399);
or OR3 (N7008, N6988, N3685, N4901);
nand NAND4 (N7009, N6980, N3993, N4955, N315);
xor XOR2 (N7010, N7008, N880);
and AND2 (N7011, N7005, N2279);
not NOT1 (N7012, N7007);
nor NOR4 (N7013, N7001, N3648, N6279, N4235);
xor XOR2 (N7014, N7011, N2354);
not NOT1 (N7015, N7003);
nor NOR3 (N7016, N7015, N4315, N4783);
nor NOR4 (N7017, N7014, N4404, N4738, N3060);
nand NAND2 (N7018, N7016, N3668);
or OR3 (N7019, N7010, N3919, N304);
nand NAND4 (N7020, N7018, N2851, N4618, N3062);
nand NAND2 (N7021, N6994, N6646);
or OR3 (N7022, N6991, N2615, N743);
and AND2 (N7023, N7009, N6472);
buf BUF1 (N7024, N7017);
buf BUF1 (N7025, N7023);
nor NOR3 (N7026, N7019, N860, N2236);
or OR3 (N7027, N7022, N1789, N2498);
and AND3 (N7028, N7027, N4523, N1471);
buf BUF1 (N7029, N7013);
and AND4 (N7030, N7012, N122, N2476, N3845);
not NOT1 (N7031, N7020);
and AND2 (N7032, N7026, N699);
buf BUF1 (N7033, N7029);
buf BUF1 (N7034, N6983);
and AND3 (N7035, N7030, N5562, N904);
nand NAND3 (N7036, N7033, N3878, N2512);
and AND3 (N7037, N7036, N6374, N4869);
buf BUF1 (N7038, N7025);
xor XOR2 (N7039, N7031, N3072);
nor NOR2 (N7040, N7028, N5635);
xor XOR2 (N7041, N7032, N5243);
and AND4 (N7042, N7035, N3763, N105, N5625);
nand NAND3 (N7043, N7034, N518, N1509);
or OR2 (N7044, N7006, N1531);
and AND2 (N7045, N7021, N3851);
xor XOR2 (N7046, N7024, N3152);
xor XOR2 (N7047, N7046, N1705);
nand NAND2 (N7048, N7042, N349);
not NOT1 (N7049, N7048);
nand NAND4 (N7050, N7049, N2867, N48, N6616);
buf BUF1 (N7051, N7044);
buf BUF1 (N7052, N7051);
and AND4 (N7053, N7043, N1242, N4583, N2010);
or OR3 (N7054, N7039, N1005, N6460);
nor NOR2 (N7055, N7045, N1875);
buf BUF1 (N7056, N7054);
nor NOR2 (N7057, N7041, N6754);
xor XOR2 (N7058, N7038, N793);
or OR4 (N7059, N7053, N2875, N3343, N207);
buf BUF1 (N7060, N7059);
xor XOR2 (N7061, N7047, N5612);
xor XOR2 (N7062, N7055, N1887);
nand NAND4 (N7063, N7061, N1867, N3863, N4114);
xor XOR2 (N7064, N7056, N4255);
or OR3 (N7065, N7052, N5449, N554);
nand NAND4 (N7066, N7064, N5830, N1577, N475);
xor XOR2 (N7067, N7065, N3298);
not NOT1 (N7068, N7063);
not NOT1 (N7069, N7037);
buf BUF1 (N7070, N7057);
nand NAND3 (N7071, N7069, N1615, N2118);
and AND3 (N7072, N7060, N5668, N5174);
not NOT1 (N7073, N7070);
nor NOR2 (N7074, N7072, N3402);
buf BUF1 (N7075, N7071);
not NOT1 (N7076, N7068);
buf BUF1 (N7077, N7058);
nand NAND3 (N7078, N7066, N2566, N1929);
buf BUF1 (N7079, N7074);
nor NOR3 (N7080, N7073, N4971, N1095);
nor NOR3 (N7081, N7050, N1629, N3983);
nand NAND4 (N7082, N7081, N1228, N3852, N5099);
nor NOR2 (N7083, N7082, N6051);
or OR3 (N7084, N7079, N3284, N5593);
and AND4 (N7085, N7084, N1359, N516, N4592);
buf BUF1 (N7086, N7083);
xor XOR2 (N7087, N7078, N1299);
nor NOR2 (N7088, N7067, N6191);
not NOT1 (N7089, N7088);
or OR2 (N7090, N7080, N2701);
or OR4 (N7091, N7086, N4394, N4018, N2102);
xor XOR2 (N7092, N7089, N6320);
buf BUF1 (N7093, N7092);
not NOT1 (N7094, N7090);
and AND4 (N7095, N7087, N1801, N3304, N6112);
or OR2 (N7096, N7040, N5624);
xor XOR2 (N7097, N7093, N4149);
not NOT1 (N7098, N7075);
xor XOR2 (N7099, N7094, N2835);
nand NAND3 (N7100, N7095, N4457, N565);
nor NOR3 (N7101, N7099, N4824, N666);
and AND3 (N7102, N7096, N2338, N2943);
xor XOR2 (N7103, N7101, N3138);
buf BUF1 (N7104, N7076);
nor NOR4 (N7105, N7085, N2160, N4664, N3514);
and AND3 (N7106, N7098, N5013, N3778);
not NOT1 (N7107, N7104);
nor NOR2 (N7108, N7103, N2318);
nor NOR4 (N7109, N7077, N2212, N2856, N6041);
and AND4 (N7110, N7100, N2330, N4491, N4133);
buf BUF1 (N7111, N7097);
xor XOR2 (N7112, N7105, N1617);
buf BUF1 (N7113, N7107);
nor NOR4 (N7114, N7112, N1356, N1219, N2990);
not NOT1 (N7115, N7106);
or OR2 (N7116, N7091, N2663);
buf BUF1 (N7117, N7108);
buf BUF1 (N7118, N7109);
or OR2 (N7119, N7118, N4789);
or OR4 (N7120, N7116, N1619, N3697, N5245);
and AND3 (N7121, N7062, N1868, N4825);
xor XOR2 (N7122, N7113, N6753);
xor XOR2 (N7123, N7119, N1144);
or OR3 (N7124, N7114, N4670, N2195);
and AND4 (N7125, N7124, N5947, N6375, N3553);
or OR4 (N7126, N7102, N5472, N5722, N3003);
buf BUF1 (N7127, N7122);
xor XOR2 (N7128, N7121, N5200);
buf BUF1 (N7129, N7128);
xor XOR2 (N7130, N7125, N977);
and AND2 (N7131, N7126, N6832);
and AND2 (N7132, N7110, N4531);
buf BUF1 (N7133, N7111);
nand NAND4 (N7134, N7117, N6047, N5000, N6136);
nand NAND3 (N7135, N7131, N442, N1473);
or OR3 (N7136, N7129, N7028, N4795);
xor XOR2 (N7137, N7127, N2736);
nand NAND2 (N7138, N7136, N2045);
nor NOR2 (N7139, N7137, N5370);
xor XOR2 (N7140, N7133, N3144);
xor XOR2 (N7141, N7135, N6216);
not NOT1 (N7142, N7130);
nor NOR3 (N7143, N7132, N1990, N4669);
not NOT1 (N7144, N7138);
nor NOR2 (N7145, N7142, N351);
nand NAND4 (N7146, N7139, N3995, N6294, N93);
xor XOR2 (N7147, N7123, N6221);
buf BUF1 (N7148, N7145);
nand NAND3 (N7149, N7146, N1742, N2430);
and AND2 (N7150, N7147, N5748);
or OR2 (N7151, N7150, N2384);
and AND2 (N7152, N7149, N6699);
or OR2 (N7153, N7120, N1567);
nand NAND4 (N7154, N7141, N1310, N4079, N4655);
or OR4 (N7155, N7154, N3033, N413, N280);
nor NOR4 (N7156, N7143, N1548, N1951, N3430);
nor NOR3 (N7157, N7115, N6668, N6846);
and AND4 (N7158, N7140, N5585, N966, N421);
or OR3 (N7159, N7157, N5613, N353);
not NOT1 (N7160, N7159);
buf BUF1 (N7161, N7134);
buf BUF1 (N7162, N7160);
or OR4 (N7163, N7151, N4715, N6616, N4616);
or OR2 (N7164, N7144, N5226);
nor NOR3 (N7165, N7158, N5457, N2270);
not NOT1 (N7166, N7155);
xor XOR2 (N7167, N7156, N3019);
buf BUF1 (N7168, N7148);
buf BUF1 (N7169, N7152);
nand NAND3 (N7170, N7168, N4992, N4550);
or OR2 (N7171, N7167, N3372);
nor NOR3 (N7172, N7162, N2345, N5442);
buf BUF1 (N7173, N7171);
buf BUF1 (N7174, N7170);
not NOT1 (N7175, N7173);
xor XOR2 (N7176, N7163, N3732);
nand NAND3 (N7177, N7153, N2485, N775);
buf BUF1 (N7178, N7177);
or OR3 (N7179, N7169, N9, N3697);
and AND4 (N7180, N7178, N954, N4130, N6404);
nor NOR2 (N7181, N7172, N3298);
nor NOR2 (N7182, N7175, N2868);
xor XOR2 (N7183, N7174, N5236);
and AND2 (N7184, N7165, N3291);
buf BUF1 (N7185, N7161);
xor XOR2 (N7186, N7181, N6905);
nand NAND2 (N7187, N7185, N2570);
xor XOR2 (N7188, N7184, N6134);
or OR2 (N7189, N7164, N1902);
nand NAND3 (N7190, N7179, N4607, N6960);
or OR4 (N7191, N7176, N235, N2366, N3340);
buf BUF1 (N7192, N7186);
xor XOR2 (N7193, N7183, N206);
nand NAND2 (N7194, N7187, N2313);
nor NOR2 (N7195, N7180, N846);
and AND2 (N7196, N7192, N2336);
not NOT1 (N7197, N7190);
buf BUF1 (N7198, N7195);
nand NAND2 (N7199, N7198, N5106);
xor XOR2 (N7200, N7166, N5998);
nand NAND3 (N7201, N7189, N4642, N1876);
or OR2 (N7202, N7193, N4470);
xor XOR2 (N7203, N7197, N2083);
and AND3 (N7204, N7194, N1337, N4005);
nand NAND4 (N7205, N7203, N4297, N4785, N2382);
and AND2 (N7206, N7199, N1351);
and AND4 (N7207, N7188, N3019, N4261, N4944);
buf BUF1 (N7208, N7200);
buf BUF1 (N7209, N7208);
buf BUF1 (N7210, N7206);
buf BUF1 (N7211, N7202);
nand NAND3 (N7212, N7182, N1335, N987);
and AND2 (N7213, N7191, N4171);
not NOT1 (N7214, N7209);
nor NOR3 (N7215, N7201, N1670, N273);
and AND3 (N7216, N7212, N5349, N5149);
and AND4 (N7217, N7210, N2061, N763, N6259);
nor NOR4 (N7218, N7196, N6652, N1779, N998);
or OR3 (N7219, N7218, N5950, N6060);
nand NAND4 (N7220, N7215, N2235, N2704, N748);
or OR3 (N7221, N7211, N1288, N2671);
nor NOR3 (N7222, N7219, N1600, N5336);
xor XOR2 (N7223, N7213, N5892);
nand NAND4 (N7224, N7222, N6815, N5929, N3784);
or OR3 (N7225, N7216, N6450, N2056);
or OR2 (N7226, N7214, N590);
and AND4 (N7227, N7224, N2633, N6862, N482);
xor XOR2 (N7228, N7205, N256);
nand NAND3 (N7229, N7220, N1351, N5278);
or OR2 (N7230, N7229, N4449);
xor XOR2 (N7231, N7225, N5546);
xor XOR2 (N7232, N7227, N4464);
nand NAND2 (N7233, N7231, N3624);
nand NAND3 (N7234, N7223, N5376, N68);
not NOT1 (N7235, N7204);
or OR4 (N7236, N7217, N2834, N6767, N3692);
xor XOR2 (N7237, N7230, N4493);
xor XOR2 (N7238, N7235, N3459);
xor XOR2 (N7239, N7237, N1974);
nand NAND4 (N7240, N7226, N4361, N5605, N978);
nor NOR3 (N7241, N7239, N394, N3193);
and AND4 (N7242, N7232, N952, N5569, N1997);
nand NAND3 (N7243, N7241, N5481, N4923);
nand NAND4 (N7244, N7228, N3124, N5026, N3374);
and AND2 (N7245, N7234, N554);
buf BUF1 (N7246, N7238);
nor NOR2 (N7247, N7236, N2552);
or OR2 (N7248, N7240, N2455);
nor NOR4 (N7249, N7221, N1478, N912, N1277);
or OR2 (N7250, N7242, N527);
buf BUF1 (N7251, N7248);
buf BUF1 (N7252, N7247);
nand NAND3 (N7253, N7244, N5428, N5801);
nand NAND2 (N7254, N7251, N1539);
nand NAND2 (N7255, N7243, N1559);
nand NAND4 (N7256, N7255, N3341, N2656, N136);
xor XOR2 (N7257, N7256, N6617);
or OR3 (N7258, N7246, N6739, N1271);
nand NAND3 (N7259, N7249, N4016, N2126);
and AND4 (N7260, N7253, N4694, N3879, N6210);
buf BUF1 (N7261, N7207);
xor XOR2 (N7262, N7261, N5738);
or OR4 (N7263, N7257, N4585, N7187, N3548);
not NOT1 (N7264, N7233);
xor XOR2 (N7265, N7262, N4879);
or OR2 (N7266, N7263, N3963);
or OR3 (N7267, N7265, N3881, N5405);
xor XOR2 (N7268, N7254, N1549);
buf BUF1 (N7269, N7267);
and AND2 (N7270, N7258, N413);
not NOT1 (N7271, N7259);
xor XOR2 (N7272, N7268, N3120);
not NOT1 (N7273, N7270);
nand NAND4 (N7274, N7272, N2580, N7094, N2497);
xor XOR2 (N7275, N7266, N3039);
not NOT1 (N7276, N7252);
and AND2 (N7277, N7245, N4516);
xor XOR2 (N7278, N7276, N2477);
xor XOR2 (N7279, N7278, N1199);
or OR3 (N7280, N7271, N4609, N4326);
buf BUF1 (N7281, N7275);
buf BUF1 (N7282, N7250);
or OR4 (N7283, N7269, N924, N1317, N6999);
or OR3 (N7284, N7260, N1398, N6213);
nor NOR2 (N7285, N7279, N1833);
or OR4 (N7286, N7283, N4305, N5029, N1280);
buf BUF1 (N7287, N7284);
nand NAND2 (N7288, N7286, N5033);
not NOT1 (N7289, N7264);
buf BUF1 (N7290, N7280);
nand NAND3 (N7291, N7289, N3941, N3031);
or OR4 (N7292, N7285, N1343, N7275, N3957);
and AND3 (N7293, N7288, N966, N4701);
buf BUF1 (N7294, N7290);
and AND4 (N7295, N7273, N2097, N6908, N1637);
nor NOR3 (N7296, N7287, N5438, N4163);
and AND3 (N7297, N7294, N7146, N4591);
or OR3 (N7298, N7296, N2146, N4501);
buf BUF1 (N7299, N7291);
not NOT1 (N7300, N7299);
xor XOR2 (N7301, N7293, N3237);
and AND3 (N7302, N7301, N518, N5976);
not NOT1 (N7303, N7274);
and AND2 (N7304, N7298, N4086);
not NOT1 (N7305, N7282);
xor XOR2 (N7306, N7277, N7026);
and AND4 (N7307, N7295, N481, N6268, N6854);
and AND3 (N7308, N7302, N362, N2609);
buf BUF1 (N7309, N7292);
buf BUF1 (N7310, N7300);
buf BUF1 (N7311, N7310);
buf BUF1 (N7312, N7308);
and AND3 (N7313, N7306, N4622, N3944);
nor NOR2 (N7314, N7297, N2072);
xor XOR2 (N7315, N7305, N3235);
or OR4 (N7316, N7312, N731, N1731, N4390);
or OR4 (N7317, N7313, N3165, N4726, N6459);
nor NOR3 (N7318, N7307, N37, N5629);
nor NOR4 (N7319, N7316, N5484, N3701, N6901);
nand NAND2 (N7320, N7311, N4051);
or OR3 (N7321, N7315, N1179, N3269);
xor XOR2 (N7322, N7314, N1689);
nand NAND4 (N7323, N7281, N6155, N2576, N2131);
not NOT1 (N7324, N7323);
and AND3 (N7325, N7303, N6794, N5337);
or OR3 (N7326, N7321, N5067, N5218);
buf BUF1 (N7327, N7309);
or OR2 (N7328, N7324, N2757);
buf BUF1 (N7329, N7322);
and AND3 (N7330, N7326, N6957, N4739);
buf BUF1 (N7331, N7325);
buf BUF1 (N7332, N7330);
buf BUF1 (N7333, N7304);
nand NAND3 (N7334, N7318, N4582, N2332);
nand NAND4 (N7335, N7331, N647, N1913, N3591);
nor NOR2 (N7336, N7329, N1751);
and AND2 (N7337, N7335, N6840);
xor XOR2 (N7338, N7333, N4562);
not NOT1 (N7339, N7332);
nand NAND4 (N7340, N7336, N3432, N770, N907);
xor XOR2 (N7341, N7334, N5254);
nor NOR2 (N7342, N7339, N4704);
or OR4 (N7343, N7328, N4109, N6587, N7064);
xor XOR2 (N7344, N7327, N2701);
and AND4 (N7345, N7338, N1186, N5710, N4577);
xor XOR2 (N7346, N7341, N5658);
buf BUF1 (N7347, N7337);
or OR3 (N7348, N7342, N4403, N5098);
xor XOR2 (N7349, N7343, N2897);
or OR2 (N7350, N7345, N1498);
buf BUF1 (N7351, N7317);
not NOT1 (N7352, N7344);
nand NAND2 (N7353, N7346, N4906);
buf BUF1 (N7354, N7320);
nand NAND4 (N7355, N7348, N496, N5671, N2919);
nand NAND2 (N7356, N7350, N1355);
or OR3 (N7357, N7349, N3213, N3011);
xor XOR2 (N7358, N7352, N6831);
nor NOR3 (N7359, N7347, N6617, N2281);
buf BUF1 (N7360, N7355);
buf BUF1 (N7361, N7354);
nand NAND2 (N7362, N7351, N3902);
or OR4 (N7363, N7359, N4933, N6627, N735);
nand NAND4 (N7364, N7361, N2617, N2688, N4001);
not NOT1 (N7365, N7360);
buf BUF1 (N7366, N7365);
buf BUF1 (N7367, N7366);
nand NAND2 (N7368, N7362, N5936);
buf BUF1 (N7369, N7319);
buf BUF1 (N7370, N7340);
nor NOR4 (N7371, N7370, N365, N4533, N4315);
or OR2 (N7372, N7357, N3312);
or OR2 (N7373, N7372, N4330);
xor XOR2 (N7374, N7353, N4944);
nor NOR4 (N7375, N7369, N5040, N5679, N4948);
and AND4 (N7376, N7368, N5804, N2996, N949);
buf BUF1 (N7377, N7356);
buf BUF1 (N7378, N7374);
buf BUF1 (N7379, N7364);
nand NAND2 (N7380, N7377, N2452);
nand NAND3 (N7381, N7367, N5559, N7201);
nor NOR4 (N7382, N7371, N4494, N255, N4440);
not NOT1 (N7383, N7378);
and AND3 (N7384, N7380, N6413, N3577);
nand NAND2 (N7385, N7381, N5683);
or OR4 (N7386, N7379, N1041, N6209, N5241);
buf BUF1 (N7387, N7385);
and AND3 (N7388, N7373, N1581, N4628);
and AND4 (N7389, N7386, N7304, N5716, N3404);
nand NAND2 (N7390, N7388, N4568);
buf BUF1 (N7391, N7384);
not NOT1 (N7392, N7358);
nor NOR3 (N7393, N7363, N792, N4948);
nand NAND4 (N7394, N7382, N5670, N960, N5383);
and AND4 (N7395, N7387, N426, N3257, N2989);
or OR4 (N7396, N7390, N2013, N2338, N5797);
and AND2 (N7397, N7383, N4882);
xor XOR2 (N7398, N7394, N779);
buf BUF1 (N7399, N7398);
and AND4 (N7400, N7395, N5247, N6504, N244);
and AND4 (N7401, N7400, N7273, N5831, N5242);
buf BUF1 (N7402, N7376);
nand NAND4 (N7403, N7389, N2716, N2696, N3356);
buf BUF1 (N7404, N7399);
nor NOR3 (N7405, N7404, N247, N6850);
not NOT1 (N7406, N7393);
and AND3 (N7407, N7397, N5742, N6377);
or OR4 (N7408, N7375, N1721, N1496, N4234);
nor NOR3 (N7409, N7407, N3302, N4825);
xor XOR2 (N7410, N7396, N6814);
and AND2 (N7411, N7392, N4777);
nand NAND2 (N7412, N7391, N7266);
buf BUF1 (N7413, N7412);
not NOT1 (N7414, N7410);
buf BUF1 (N7415, N7411);
or OR2 (N7416, N7415, N3216);
buf BUF1 (N7417, N7403);
nand NAND4 (N7418, N7402, N5605, N7391, N6908);
and AND4 (N7419, N7409, N5341, N1366, N33);
nand NAND3 (N7420, N7417, N1090, N1005);
nand NAND2 (N7421, N7406, N6499);
xor XOR2 (N7422, N7405, N2151);
not NOT1 (N7423, N7418);
buf BUF1 (N7424, N7420);
or OR2 (N7425, N7423, N3765);
xor XOR2 (N7426, N7422, N1316);
not NOT1 (N7427, N7426);
xor XOR2 (N7428, N7416, N344);
xor XOR2 (N7429, N7425, N6568);
buf BUF1 (N7430, N7419);
buf BUF1 (N7431, N7424);
and AND4 (N7432, N7429, N5252, N1793, N3370);
or OR4 (N7433, N7427, N1868, N2502, N5661);
not NOT1 (N7434, N7421);
and AND3 (N7435, N7432, N2694, N685);
nand NAND4 (N7436, N7433, N2089, N7355, N4995);
not NOT1 (N7437, N7431);
nand NAND2 (N7438, N7408, N681);
xor XOR2 (N7439, N7430, N1753);
or OR2 (N7440, N7401, N6520);
and AND4 (N7441, N7438, N4355, N6716, N827);
nand NAND4 (N7442, N7428, N483, N3031, N5420);
xor XOR2 (N7443, N7414, N4128);
nand NAND2 (N7444, N7436, N4377);
or OR4 (N7445, N7439, N96, N3167, N1402);
nand NAND3 (N7446, N7442, N1753, N7244);
nand NAND2 (N7447, N7435, N955);
nor NOR3 (N7448, N7413, N693, N806);
xor XOR2 (N7449, N7447, N5006);
xor XOR2 (N7450, N7443, N5436);
xor XOR2 (N7451, N7441, N4026);
and AND4 (N7452, N7446, N2006, N3418, N871);
or OR2 (N7453, N7448, N4536);
or OR3 (N7454, N7445, N5369, N3253);
nand NAND2 (N7455, N7434, N5250);
xor XOR2 (N7456, N7454, N5406);
or OR3 (N7457, N7455, N5820, N4033);
or OR3 (N7458, N7450, N3579, N5733);
nor NOR2 (N7459, N7456, N5609);
nor NOR3 (N7460, N7453, N6378, N5843);
or OR4 (N7461, N7440, N643, N375, N2494);
nor NOR4 (N7462, N7437, N1356, N587, N5962);
nand NAND4 (N7463, N7458, N464, N6201, N7172);
not NOT1 (N7464, N7452);
and AND4 (N7465, N7451, N4434, N6340, N4705);
not NOT1 (N7466, N7449);
xor XOR2 (N7467, N7465, N1341);
and AND4 (N7468, N7463, N5168, N6136, N5427);
or OR3 (N7469, N7468, N856, N884);
and AND2 (N7470, N7460, N3466);
xor XOR2 (N7471, N7464, N4120);
and AND3 (N7472, N7467, N5591, N5025);
buf BUF1 (N7473, N7469);
nor NOR4 (N7474, N7466, N1469, N2301, N1031);
or OR4 (N7475, N7461, N3516, N3325, N6144);
nor NOR4 (N7476, N7475, N711, N5527, N306);
buf BUF1 (N7477, N7471);
nor NOR3 (N7478, N7444, N1062, N4261);
nand NAND3 (N7479, N7474, N673, N6799);
xor XOR2 (N7480, N7476, N4752);
or OR3 (N7481, N7459, N5888, N6131);
nor NOR4 (N7482, N7479, N3580, N5177, N2189);
not NOT1 (N7483, N7473);
or OR2 (N7484, N7477, N2120);
and AND3 (N7485, N7462, N5320, N2140);
buf BUF1 (N7486, N7483);
buf BUF1 (N7487, N7486);
not NOT1 (N7488, N7481);
buf BUF1 (N7489, N7457);
or OR3 (N7490, N7478, N2555, N2646);
and AND4 (N7491, N7482, N3522, N2316, N2536);
not NOT1 (N7492, N7491);
nand NAND3 (N7493, N7480, N2707, N4010);
xor XOR2 (N7494, N7484, N1432);
nor NOR3 (N7495, N7492, N2898, N2842);
xor XOR2 (N7496, N7470, N6703);
xor XOR2 (N7497, N7490, N1986);
not NOT1 (N7498, N7495);
nand NAND3 (N7499, N7485, N885, N3522);
nand NAND4 (N7500, N7493, N4599, N836, N2942);
and AND3 (N7501, N7489, N619, N3483);
and AND3 (N7502, N7497, N91, N6007);
not NOT1 (N7503, N7501);
buf BUF1 (N7504, N7502);
buf BUF1 (N7505, N7503);
not NOT1 (N7506, N7487);
nand NAND4 (N7507, N7472, N3830, N5831, N7143);
xor XOR2 (N7508, N7505, N6487);
and AND2 (N7509, N7507, N2011);
or OR4 (N7510, N7504, N6070, N4016, N3551);
nor NOR2 (N7511, N7506, N4932);
nand NAND3 (N7512, N7508, N421, N237);
nand NAND4 (N7513, N7488, N4133, N3983, N104);
not NOT1 (N7514, N7511);
xor XOR2 (N7515, N7499, N1923);
buf BUF1 (N7516, N7494);
or OR4 (N7517, N7512, N6331, N2246, N603);
or OR4 (N7518, N7513, N4499, N5714, N726);
buf BUF1 (N7519, N7510);
and AND4 (N7520, N7516, N1596, N3026, N7292);
xor XOR2 (N7521, N7520, N691);
or OR3 (N7522, N7519, N3141, N694);
not NOT1 (N7523, N7509);
buf BUF1 (N7524, N7496);
buf BUF1 (N7525, N7524);
xor XOR2 (N7526, N7498, N341);
buf BUF1 (N7527, N7514);
xor XOR2 (N7528, N7518, N1913);
nand NAND3 (N7529, N7522, N1090, N689);
xor XOR2 (N7530, N7528, N6087);
nor NOR2 (N7531, N7500, N3684);
xor XOR2 (N7532, N7527, N4197);
nand NAND3 (N7533, N7525, N6076, N1073);
and AND4 (N7534, N7531, N1379, N2123, N5940);
or OR4 (N7535, N7517, N1787, N6360, N2702);
xor XOR2 (N7536, N7526, N5664);
buf BUF1 (N7537, N7523);
or OR4 (N7538, N7537, N966, N7074, N4664);
and AND2 (N7539, N7515, N2294);
buf BUF1 (N7540, N7535);
nor NOR3 (N7541, N7533, N44, N2260);
not NOT1 (N7542, N7538);
buf BUF1 (N7543, N7534);
not NOT1 (N7544, N7536);
or OR4 (N7545, N7532, N2274, N5918, N1596);
not NOT1 (N7546, N7530);
xor XOR2 (N7547, N7545, N5250);
buf BUF1 (N7548, N7543);
buf BUF1 (N7549, N7539);
and AND2 (N7550, N7549, N4044);
nand NAND2 (N7551, N7529, N5903);
or OR2 (N7552, N7547, N4649);
nor NOR4 (N7553, N7548, N3804, N3517, N778);
xor XOR2 (N7554, N7541, N7452);
or OR4 (N7555, N7552, N931, N6562, N736);
xor XOR2 (N7556, N7521, N2737);
buf BUF1 (N7557, N7553);
nor NOR3 (N7558, N7544, N233, N6332);
xor XOR2 (N7559, N7551, N2392);
buf BUF1 (N7560, N7556);
and AND3 (N7561, N7558, N974, N5383);
buf BUF1 (N7562, N7561);
buf BUF1 (N7563, N7542);
nand NAND3 (N7564, N7540, N275, N5009);
xor XOR2 (N7565, N7550, N1214);
xor XOR2 (N7566, N7562, N7073);
nor NOR2 (N7567, N7563, N7565);
not NOT1 (N7568, N7371);
buf BUF1 (N7569, N7555);
not NOT1 (N7570, N7566);
nand NAND4 (N7571, N7570, N1099, N526, N7407);
buf BUF1 (N7572, N7567);
or OR2 (N7573, N7571, N6781);
buf BUF1 (N7574, N7573);
and AND4 (N7575, N7564, N5706, N1017, N3806);
or OR4 (N7576, N7546, N5312, N7192, N6782);
not NOT1 (N7577, N7569);
and AND2 (N7578, N7577, N346);
xor XOR2 (N7579, N7572, N2521);
not NOT1 (N7580, N7560);
not NOT1 (N7581, N7575);
xor XOR2 (N7582, N7559, N552);
nand NAND4 (N7583, N7582, N3791, N5984, N1727);
buf BUF1 (N7584, N7557);
nand NAND3 (N7585, N7581, N4398, N6336);
buf BUF1 (N7586, N7574);
nand NAND2 (N7587, N7579, N6853);
xor XOR2 (N7588, N7578, N6209);
buf BUF1 (N7589, N7588);
and AND2 (N7590, N7554, N3859);
not NOT1 (N7591, N7584);
not NOT1 (N7592, N7589);
nand NAND4 (N7593, N7590, N787, N4563, N1971);
or OR3 (N7594, N7593, N3203, N4075);
nor NOR4 (N7595, N7580, N229, N3394, N5119);
xor XOR2 (N7596, N7591, N393);
and AND3 (N7597, N7583, N3570, N1885);
and AND2 (N7598, N7587, N3070);
buf BUF1 (N7599, N7595);
nor NOR2 (N7600, N7596, N4935);
nand NAND2 (N7601, N7586, N463);
buf BUF1 (N7602, N7598);
nor NOR3 (N7603, N7576, N3211, N4491);
not NOT1 (N7604, N7602);
buf BUF1 (N7605, N7603);
xor XOR2 (N7606, N7592, N7427);
or OR3 (N7607, N7599, N6256, N6397);
nor NOR2 (N7608, N7600, N7444);
nor NOR3 (N7609, N7601, N3843, N3117);
nor NOR4 (N7610, N7608, N3659, N7213, N5601);
or OR4 (N7611, N7610, N4585, N1147, N3230);
xor XOR2 (N7612, N7605, N5307);
xor XOR2 (N7613, N7568, N2105);
nand NAND4 (N7614, N7606, N3122, N4220, N6999);
xor XOR2 (N7615, N7614, N4805);
not NOT1 (N7616, N7594);
or OR2 (N7617, N7616, N4581);
not NOT1 (N7618, N7613);
not NOT1 (N7619, N7597);
xor XOR2 (N7620, N7611, N3689);
not NOT1 (N7621, N7618);
not NOT1 (N7622, N7612);
xor XOR2 (N7623, N7585, N869);
buf BUF1 (N7624, N7615);
xor XOR2 (N7625, N7624, N4429);
or OR2 (N7626, N7622, N6633);
nand NAND4 (N7627, N7604, N3072, N6460, N2434);
nand NAND4 (N7628, N7617, N4503, N2670, N5802);
buf BUF1 (N7629, N7625);
xor XOR2 (N7630, N7628, N4272);
xor XOR2 (N7631, N7621, N7509);
and AND3 (N7632, N7629, N4112, N1900);
not NOT1 (N7633, N7620);
xor XOR2 (N7634, N7607, N5133);
nand NAND2 (N7635, N7627, N7212);
buf BUF1 (N7636, N7635);
xor XOR2 (N7637, N7626, N6499);
xor XOR2 (N7638, N7609, N4458);
nand NAND4 (N7639, N7619, N6574, N1291, N2285);
and AND3 (N7640, N7632, N3532, N1066);
and AND4 (N7641, N7634, N6115, N2079, N128);
buf BUF1 (N7642, N7633);
xor XOR2 (N7643, N7637, N5922);
xor XOR2 (N7644, N7642, N5367);
buf BUF1 (N7645, N7640);
and AND2 (N7646, N7636, N1315);
nand NAND3 (N7647, N7630, N5607, N2426);
xor XOR2 (N7648, N7647, N3737);
and AND4 (N7649, N7623, N2552, N277, N7271);
and AND2 (N7650, N7638, N3733);
nor NOR2 (N7651, N7648, N4187);
nand NAND4 (N7652, N7641, N7280, N4178, N3511);
nor NOR2 (N7653, N7631, N3511);
buf BUF1 (N7654, N7644);
buf BUF1 (N7655, N7645);
not NOT1 (N7656, N7649);
xor XOR2 (N7657, N7654, N5094);
xor XOR2 (N7658, N7653, N648);
xor XOR2 (N7659, N7639, N4478);
nand NAND4 (N7660, N7656, N187, N4751, N2672);
nand NAND3 (N7661, N7655, N6217, N3557);
nand NAND2 (N7662, N7643, N2489);
nor NOR3 (N7663, N7646, N2036, N1652);
not NOT1 (N7664, N7661);
and AND4 (N7665, N7658, N5308, N2295, N2096);
buf BUF1 (N7666, N7660);
and AND2 (N7667, N7666, N2332);
nor NOR3 (N7668, N7650, N5974, N3558);
nand NAND3 (N7669, N7657, N4666, N915);
and AND2 (N7670, N7668, N4584);
buf BUF1 (N7671, N7664);
or OR3 (N7672, N7662, N7365, N3042);
and AND4 (N7673, N7672, N4244, N921, N5782);
nand NAND3 (N7674, N7663, N7670, N1915);
nor NOR3 (N7675, N3000, N530, N5438);
xor XOR2 (N7676, N7673, N4656);
nor NOR4 (N7677, N7667, N6740, N5021, N6537);
nor NOR3 (N7678, N7652, N7100, N5794);
xor XOR2 (N7679, N7665, N756);
nand NAND2 (N7680, N7659, N3434);
not NOT1 (N7681, N7675);
nor NOR4 (N7682, N7681, N5298, N2379, N1156);
or OR3 (N7683, N7680, N4294, N5470);
or OR3 (N7684, N7651, N300, N3791);
nand NAND2 (N7685, N7677, N2309);
buf BUF1 (N7686, N7678);
and AND4 (N7687, N7676, N7251, N2010, N3181);
and AND2 (N7688, N7669, N2634);
or OR2 (N7689, N7674, N5553);
nor NOR3 (N7690, N7682, N173, N6749);
nor NOR2 (N7691, N7684, N2591);
not NOT1 (N7692, N7686);
buf BUF1 (N7693, N7691);
not NOT1 (N7694, N7693);
not NOT1 (N7695, N7692);
xor XOR2 (N7696, N7695, N1840);
buf BUF1 (N7697, N7696);
xor XOR2 (N7698, N7689, N1242);
nand NAND3 (N7699, N7694, N1089, N3880);
or OR2 (N7700, N7690, N1245);
not NOT1 (N7701, N7699);
and AND4 (N7702, N7697, N3868, N5844, N5163);
or OR4 (N7703, N7685, N1944, N2143, N2661);
buf BUF1 (N7704, N7683);
buf BUF1 (N7705, N7679);
or OR4 (N7706, N7688, N2742, N6090, N5490);
nor NOR2 (N7707, N7671, N32);
or OR4 (N7708, N7698, N7276, N7262, N6926);
xor XOR2 (N7709, N7700, N975);
nand NAND2 (N7710, N7707, N7542);
buf BUF1 (N7711, N7701);
nor NOR3 (N7712, N7710, N5417, N2092);
buf BUF1 (N7713, N7706);
not NOT1 (N7714, N7704);
buf BUF1 (N7715, N7711);
nand NAND2 (N7716, N7705, N220);
nor NOR3 (N7717, N7709, N978, N6682);
or OR4 (N7718, N7687, N751, N4519, N2223);
or OR4 (N7719, N7702, N5602, N3112, N6606);
nor NOR2 (N7720, N7703, N691);
and AND2 (N7721, N7713, N3847);
nand NAND2 (N7722, N7714, N1955);
nand NAND2 (N7723, N7716, N7558);
or OR3 (N7724, N7720, N813, N309);
not NOT1 (N7725, N7721);
or OR2 (N7726, N7718, N4618);
nor NOR3 (N7727, N7717, N5701, N3684);
or OR2 (N7728, N7724, N8);
or OR3 (N7729, N7723, N6816, N5737);
buf BUF1 (N7730, N7708);
buf BUF1 (N7731, N7725);
or OR4 (N7732, N7728, N6949, N417, N3334);
not NOT1 (N7733, N7727);
buf BUF1 (N7734, N7729);
and AND2 (N7735, N7722, N1860);
xor XOR2 (N7736, N7730, N5444);
nand NAND4 (N7737, N7733, N2609, N528, N1044);
nand NAND4 (N7738, N7734, N6926, N2453, N4885);
nor NOR2 (N7739, N7715, N6807);
buf BUF1 (N7740, N7726);
and AND4 (N7741, N7719, N6464, N2919, N6370);
or OR2 (N7742, N7738, N351);
not NOT1 (N7743, N7741);
and AND2 (N7744, N7742, N1962);
not NOT1 (N7745, N7743);
nor NOR2 (N7746, N7712, N4719);
buf BUF1 (N7747, N7744);
buf BUF1 (N7748, N7739);
or OR3 (N7749, N7736, N4104, N1263);
nand NAND2 (N7750, N7749, N5384);
buf BUF1 (N7751, N7737);
xor XOR2 (N7752, N7750, N5551);
nor NOR2 (N7753, N7746, N5673);
nor NOR3 (N7754, N7732, N1301, N5088);
nand NAND3 (N7755, N7753, N2971, N4976);
nor NOR3 (N7756, N7735, N291, N6586);
or OR3 (N7757, N7751, N2485, N4885);
xor XOR2 (N7758, N7752, N1499);
and AND4 (N7759, N7745, N4274, N2587, N3540);
buf BUF1 (N7760, N7731);
xor XOR2 (N7761, N7760, N7223);
xor XOR2 (N7762, N7759, N686);
nor NOR3 (N7763, N7755, N24, N1495);
and AND4 (N7764, N7757, N1507, N4231, N1620);
xor XOR2 (N7765, N7762, N7687);
or OR3 (N7766, N7758, N6295, N4096);
nand NAND3 (N7767, N7765, N1750, N552);
not NOT1 (N7768, N7767);
nand NAND2 (N7769, N7761, N5726);
xor XOR2 (N7770, N7756, N1109);
not NOT1 (N7771, N7769);
nor NOR2 (N7772, N7766, N5979);
xor XOR2 (N7773, N7764, N1972);
not NOT1 (N7774, N7768);
xor XOR2 (N7775, N7747, N3851);
or OR2 (N7776, N7772, N1191);
or OR3 (N7777, N7775, N6070, N2323);
xor XOR2 (N7778, N7754, N7655);
xor XOR2 (N7779, N7777, N1622);
xor XOR2 (N7780, N7773, N3991);
xor XOR2 (N7781, N7763, N3047);
xor XOR2 (N7782, N7781, N1970);
and AND4 (N7783, N7748, N4515, N2643, N6422);
nor NOR3 (N7784, N7770, N5693, N7729);
not NOT1 (N7785, N7740);
xor XOR2 (N7786, N7779, N898);
and AND3 (N7787, N7783, N1617, N803);
or OR2 (N7788, N7778, N1497);
buf BUF1 (N7789, N7771);
or OR2 (N7790, N7774, N755);
buf BUF1 (N7791, N7782);
and AND4 (N7792, N7786, N682, N5202, N4963);
not NOT1 (N7793, N7780);
nor NOR3 (N7794, N7791, N1246, N3971);
nor NOR2 (N7795, N7794, N5095);
or OR4 (N7796, N7787, N7090, N4888, N4728);
buf BUF1 (N7797, N7789);
nor NOR3 (N7798, N7784, N3999, N3553);
and AND2 (N7799, N7788, N3046);
not NOT1 (N7800, N7798);
and AND4 (N7801, N7796, N1756, N12, N4572);
or OR2 (N7802, N7792, N5369);
and AND4 (N7803, N7785, N1953, N7308, N637);
not NOT1 (N7804, N7795);
buf BUF1 (N7805, N7797);
not NOT1 (N7806, N7802);
and AND3 (N7807, N7805, N5014, N7209);
not NOT1 (N7808, N7803);
not NOT1 (N7809, N7790);
not NOT1 (N7810, N7809);
or OR2 (N7811, N7804, N4115);
xor XOR2 (N7812, N7810, N139);
xor XOR2 (N7813, N7807, N4334);
buf BUF1 (N7814, N7799);
xor XOR2 (N7815, N7813, N3947);
and AND2 (N7816, N7800, N3164);
and AND3 (N7817, N7811, N5365, N1823);
buf BUF1 (N7818, N7806);
or OR3 (N7819, N7793, N6775, N6295);
nand NAND3 (N7820, N7817, N887, N827);
xor XOR2 (N7821, N7808, N4842);
buf BUF1 (N7822, N7818);
nand NAND2 (N7823, N7801, N3336);
nor NOR4 (N7824, N7822, N491, N1840, N1630);
nand NAND3 (N7825, N7823, N3385, N6701);
and AND4 (N7826, N7816, N7764, N4062, N1914);
or OR2 (N7827, N7814, N1986);
not NOT1 (N7828, N7821);
not NOT1 (N7829, N7819);
nor NOR3 (N7830, N7829, N2917, N5659);
and AND3 (N7831, N7812, N7435, N7529);
or OR4 (N7832, N7825, N400, N1294, N6136);
xor XOR2 (N7833, N7820, N754);
buf BUF1 (N7834, N7832);
not NOT1 (N7835, N7776);
nor NOR2 (N7836, N7834, N994);
xor XOR2 (N7837, N7827, N1880);
xor XOR2 (N7838, N7833, N2168);
nand NAND3 (N7839, N7831, N3131, N3976);
and AND4 (N7840, N7830, N3709, N1818, N612);
buf BUF1 (N7841, N7828);
not NOT1 (N7842, N7824);
nand NAND4 (N7843, N7836, N7621, N6017, N5746);
nor NOR3 (N7844, N7835, N3683, N7765);
xor XOR2 (N7845, N7837, N547);
or OR4 (N7846, N7841, N2677, N4532, N7804);
and AND3 (N7847, N7840, N1810, N6218);
or OR4 (N7848, N7844, N548, N3450, N3646);
not NOT1 (N7849, N7848);
nor NOR4 (N7850, N7826, N5010, N632, N3496);
buf BUF1 (N7851, N7847);
buf BUF1 (N7852, N7849);
nand NAND4 (N7853, N7851, N6085, N6305, N3427);
not NOT1 (N7854, N7839);
xor XOR2 (N7855, N7843, N6635);
buf BUF1 (N7856, N7853);
buf BUF1 (N7857, N7855);
and AND2 (N7858, N7815, N793);
or OR4 (N7859, N7838, N6900, N3725, N740);
nand NAND4 (N7860, N7859, N917, N134, N6455);
nand NAND4 (N7861, N7850, N1208, N5996, N5686);
nor NOR2 (N7862, N7852, N745);
nor NOR2 (N7863, N7854, N1034);
not NOT1 (N7864, N7856);
buf BUF1 (N7865, N7863);
nor NOR4 (N7866, N7858, N2626, N700, N6176);
or OR3 (N7867, N7861, N5963, N4788);
buf BUF1 (N7868, N7864);
not NOT1 (N7869, N7866);
and AND3 (N7870, N7862, N6880, N1000);
nor NOR2 (N7871, N7867, N967);
and AND3 (N7872, N7869, N4130, N1996);
not NOT1 (N7873, N7845);
not NOT1 (N7874, N7846);
nand NAND3 (N7875, N7860, N7757, N2177);
xor XOR2 (N7876, N7873, N4143);
buf BUF1 (N7877, N7870);
xor XOR2 (N7878, N7875, N994);
not NOT1 (N7879, N7857);
xor XOR2 (N7880, N7879, N4039);
and AND2 (N7881, N7876, N1578);
xor XOR2 (N7882, N7872, N2834);
nand NAND3 (N7883, N7842, N468, N321);
nor NOR3 (N7884, N7865, N6546, N251);
nand NAND2 (N7885, N7877, N4257);
nand NAND4 (N7886, N7885, N6385, N2086, N3763);
xor XOR2 (N7887, N7878, N4775);
nor NOR4 (N7888, N7871, N5792, N5006, N6565);
buf BUF1 (N7889, N7881);
and AND4 (N7890, N7868, N5693, N3593, N4542);
and AND4 (N7891, N7888, N7225, N3665, N1692);
not NOT1 (N7892, N7880);
or OR2 (N7893, N7891, N7353);
nand NAND4 (N7894, N7884, N3797, N3999, N107);
not NOT1 (N7895, N7882);
nand NAND3 (N7896, N7893, N3189, N43);
and AND2 (N7897, N7896, N2445);
xor XOR2 (N7898, N7874, N3352);
buf BUF1 (N7899, N7886);
buf BUF1 (N7900, N7889);
xor XOR2 (N7901, N7899, N4192);
nand NAND3 (N7902, N7900, N1271, N2597);
and AND2 (N7903, N7898, N3026);
buf BUF1 (N7904, N7895);
not NOT1 (N7905, N7883);
and AND4 (N7906, N7890, N5740, N3978, N7);
nor NOR4 (N7907, N7903, N6784, N4548, N2076);
nor NOR4 (N7908, N7902, N2924, N1455, N1807);
nand NAND4 (N7909, N7901, N5535, N6792, N1222);
and AND4 (N7910, N7909, N2843, N4866, N1257);
nand NAND2 (N7911, N7892, N2892);
not NOT1 (N7912, N7910);
xor XOR2 (N7913, N7904, N6311);
nor NOR4 (N7914, N7913, N2228, N6880, N2457);
nor NOR2 (N7915, N7905, N4841);
or OR4 (N7916, N7894, N7646, N1782, N302);
xor XOR2 (N7917, N7915, N1027);
or OR3 (N7918, N7897, N2925, N1024);
or OR3 (N7919, N7887, N1793, N3923);
nand NAND2 (N7920, N7914, N7551);
nor NOR2 (N7921, N7916, N1366);
and AND4 (N7922, N7917, N2396, N2109, N3979);
xor XOR2 (N7923, N7919, N1246);
or OR3 (N7924, N7918, N6582, N4609);
nor NOR4 (N7925, N7924, N6854, N6298, N1640);
not NOT1 (N7926, N7911);
xor XOR2 (N7927, N7912, N1190);
nor NOR2 (N7928, N7927, N596);
and AND2 (N7929, N7925, N4701);
nor NOR3 (N7930, N7928, N3407, N2192);
xor XOR2 (N7931, N7929, N1099);
nor NOR2 (N7932, N7926, N328);
not NOT1 (N7933, N7921);
xor XOR2 (N7934, N7933, N163);
nor NOR3 (N7935, N7931, N6926, N1562);
and AND3 (N7936, N7908, N6218, N528);
nor NOR4 (N7937, N7936, N3236, N7014, N3324);
xor XOR2 (N7938, N7922, N3785);
buf BUF1 (N7939, N7923);
not NOT1 (N7940, N7934);
or OR3 (N7941, N7930, N3548, N5017);
buf BUF1 (N7942, N7940);
nor NOR3 (N7943, N7935, N7826, N2538);
or OR4 (N7944, N7939, N6162, N2596, N2897);
buf BUF1 (N7945, N7942);
nand NAND4 (N7946, N7937, N5945, N6094, N2447);
nand NAND4 (N7947, N7932, N7448, N6246, N6944);
and AND4 (N7948, N7906, N5778, N6618, N2968);
and AND4 (N7949, N7907, N2293, N2472, N2771);
buf BUF1 (N7950, N7920);
xor XOR2 (N7951, N7949, N5793);
buf BUF1 (N7952, N7950);
nor NOR4 (N7953, N7951, N3275, N3763, N6958);
buf BUF1 (N7954, N7943);
xor XOR2 (N7955, N7945, N1109);
not NOT1 (N7956, N7952);
buf BUF1 (N7957, N7948);
and AND2 (N7958, N7944, N6919);
buf BUF1 (N7959, N7946);
nand NAND4 (N7960, N7955, N7010, N2705, N6866);
and AND2 (N7961, N7956, N7390);
or OR2 (N7962, N7947, N7357);
nand NAND4 (N7963, N7957, N5870, N5152, N3020);
not NOT1 (N7964, N7963);
nand NAND4 (N7965, N7958, N2584, N7224, N227);
nor NOR4 (N7966, N7961, N172, N2611, N6153);
nand NAND2 (N7967, N7960, N2261);
or OR3 (N7968, N7967, N5431, N3664);
xor XOR2 (N7969, N7962, N7680);
and AND3 (N7970, N7953, N2976, N7348);
nor NOR2 (N7971, N7954, N6060);
nand NAND2 (N7972, N7964, N4135);
and AND4 (N7973, N7968, N3248, N4944, N7822);
nor NOR2 (N7974, N7973, N5433);
nor NOR2 (N7975, N7974, N3333);
nand NAND4 (N7976, N7975, N5088, N1233, N7500);
nor NOR4 (N7977, N7969, N823, N5975, N1723);
nor NOR4 (N7978, N7938, N6082, N6507, N3798);
not NOT1 (N7979, N7971);
nor NOR4 (N7980, N7979, N7935, N6091, N3744);
not NOT1 (N7981, N7965);
or OR2 (N7982, N7977, N2075);
and AND4 (N7983, N7970, N5422, N1751, N3338);
not NOT1 (N7984, N7941);
xor XOR2 (N7985, N7966, N7832);
buf BUF1 (N7986, N7983);
or OR3 (N7987, N7982, N6509, N2659);
or OR3 (N7988, N7978, N2133, N6325);
or OR3 (N7989, N7985, N6474, N6872);
nand NAND2 (N7990, N7986, N1870);
buf BUF1 (N7991, N7972);
or OR3 (N7992, N7990, N7174, N3095);
and AND4 (N7993, N7981, N225, N579, N7970);
or OR4 (N7994, N7976, N2400, N2476, N1210);
nand NAND2 (N7995, N7991, N3311);
or OR2 (N7996, N7993, N4449);
xor XOR2 (N7997, N7988, N5021);
or OR2 (N7998, N7980, N2800);
xor XOR2 (N7999, N7995, N6785);
nor NOR3 (N8000, N7959, N7774, N7796);
nor NOR3 (N8001, N8000, N3171, N815);
and AND4 (N8002, N7992, N5154, N4902, N755);
nor NOR4 (N8003, N8001, N3987, N2084, N6385);
xor XOR2 (N8004, N7998, N3734);
xor XOR2 (N8005, N8003, N5700);
nor NOR3 (N8006, N7984, N5729, N4885);
not NOT1 (N8007, N8004);
and AND3 (N8008, N8007, N1881, N5397);
nor NOR4 (N8009, N7987, N3120, N6522, N2961);
or OR2 (N8010, N7997, N5693);
nor NOR3 (N8011, N8002, N3276, N5876);
or OR3 (N8012, N7996, N7863, N1948);
xor XOR2 (N8013, N8005, N4608);
not NOT1 (N8014, N8006);
xor XOR2 (N8015, N7989, N4010);
buf BUF1 (N8016, N8008);
nand NAND3 (N8017, N7994, N3594, N7548);
or OR4 (N8018, N8015, N5685, N5581, N7036);
buf BUF1 (N8019, N7999);
not NOT1 (N8020, N8018);
buf BUF1 (N8021, N8019);
not NOT1 (N8022, N8011);
xor XOR2 (N8023, N8010, N4195);
not NOT1 (N8024, N8016);
endmodule