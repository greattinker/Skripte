// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N809,N805,N797,N778,N803,N804,N806,N800,N807,N811;

xor XOR2 (N12, N11, N6);
not NOT1 (N13, N1);
nand NAND3 (N14, N7, N6, N10);
and AND2 (N15, N4, N1);
not NOT1 (N16, N1);
buf BUF1 (N17, N9);
or OR3 (N18, N15, N3, N3);
xor XOR2 (N19, N7, N11);
not NOT1 (N20, N7);
not NOT1 (N21, N15);
nor NOR2 (N22, N19, N21);
nor NOR2 (N23, N13, N17);
xor XOR2 (N24, N1, N22);
xor XOR2 (N25, N23, N24);
xor XOR2 (N26, N19, N11);
xor XOR2 (N27, N11, N24);
not NOT1 (N28, N3);
not NOT1 (N29, N9);
xor XOR2 (N30, N14, N16);
not NOT1 (N31, N11);
not NOT1 (N32, N29);
and AND2 (N33, N12, N27);
and AND3 (N34, N15, N13, N15);
nor NOR4 (N35, N18, N13, N32, N9);
buf BUF1 (N36, N11);
xor XOR2 (N37, N20, N33);
nor NOR3 (N38, N15, N25, N24);
and AND3 (N39, N31, N6, N18);
nor NOR2 (N40, N8, N26);
and AND2 (N41, N22, N15);
not NOT1 (N42, N35);
buf BUF1 (N43, N37);
nor NOR2 (N44, N30, N12);
or OR3 (N45, N42, N13, N24);
not NOT1 (N46, N40);
not NOT1 (N47, N34);
xor XOR2 (N48, N47, N12);
not NOT1 (N49, N28);
nand NAND4 (N50, N46, N43, N1, N21);
nor NOR3 (N51, N6, N10, N43);
buf BUF1 (N52, N36);
buf BUF1 (N53, N51);
xor XOR2 (N54, N50, N23);
and AND4 (N55, N49, N50, N39, N2);
buf BUF1 (N56, N17);
nand NAND3 (N57, N56, N25, N12);
nand NAND4 (N58, N38, N18, N19, N9);
buf BUF1 (N59, N45);
and AND4 (N60, N41, N4, N28, N49);
and AND3 (N61, N48, N38, N11);
xor XOR2 (N62, N59, N24);
nand NAND2 (N63, N60, N55);
and AND2 (N64, N42, N14);
buf BUF1 (N65, N63);
nand NAND4 (N66, N57, N2, N64, N30);
buf BUF1 (N67, N63);
or OR2 (N68, N66, N32);
buf BUF1 (N69, N68);
nor NOR3 (N70, N65, N19, N17);
buf BUF1 (N71, N58);
nor NOR4 (N72, N67, N30, N68, N61);
xor XOR2 (N73, N38, N71);
or OR4 (N74, N4, N33, N54, N13);
and AND2 (N75, N64, N11);
xor XOR2 (N76, N73, N33);
xor XOR2 (N77, N69, N51);
nor NOR3 (N78, N70, N7, N30);
buf BUF1 (N79, N74);
nand NAND3 (N80, N44, N74, N66);
not NOT1 (N81, N75);
and AND3 (N82, N62, N75, N6);
nand NAND3 (N83, N79, N4, N10);
or OR4 (N84, N81, N43, N50, N10);
and AND2 (N85, N77, N33);
xor XOR2 (N86, N85, N16);
or OR2 (N87, N86, N22);
buf BUF1 (N88, N84);
xor XOR2 (N89, N52, N75);
buf BUF1 (N90, N80);
nand NAND3 (N91, N90, N81, N77);
xor XOR2 (N92, N83, N4);
nand NAND2 (N93, N76, N50);
not NOT1 (N94, N53);
xor XOR2 (N95, N88, N77);
xor XOR2 (N96, N91, N49);
and AND2 (N97, N95, N63);
not NOT1 (N98, N72);
xor XOR2 (N99, N93, N17);
not NOT1 (N100, N98);
nand NAND3 (N101, N100, N25, N37);
and AND3 (N102, N94, N70, N7);
nand NAND4 (N103, N97, N64, N55, N21);
buf BUF1 (N104, N96);
buf BUF1 (N105, N101);
not NOT1 (N106, N92);
nor NOR3 (N107, N103, N36, N91);
buf BUF1 (N108, N107);
buf BUF1 (N109, N78);
buf BUF1 (N110, N104);
not NOT1 (N111, N105);
and AND2 (N112, N99, N77);
or OR2 (N113, N110, N59);
and AND4 (N114, N106, N34, N44, N40);
nor NOR3 (N115, N108, N72, N80);
xor XOR2 (N116, N89, N98);
not NOT1 (N117, N112);
and AND2 (N118, N111, N26);
xor XOR2 (N119, N117, N43);
and AND3 (N120, N102, N111, N94);
nor NOR3 (N121, N87, N116, N103);
buf BUF1 (N122, N52);
buf BUF1 (N123, N120);
xor XOR2 (N124, N118, N66);
nand NAND3 (N125, N123, N34, N98);
not NOT1 (N126, N109);
not NOT1 (N127, N115);
not NOT1 (N128, N121);
not NOT1 (N129, N128);
nand NAND3 (N130, N113, N35, N33);
nand NAND4 (N131, N119, N26, N13, N84);
xor XOR2 (N132, N126, N113);
xor XOR2 (N133, N125, N33);
nand NAND3 (N134, N122, N86, N108);
buf BUF1 (N135, N132);
xor XOR2 (N136, N124, N132);
buf BUF1 (N137, N127);
nand NAND3 (N138, N137, N73, N127);
xor XOR2 (N139, N135, N110);
and AND3 (N140, N82, N86, N58);
or OR4 (N141, N114, N100, N91, N94);
nor NOR4 (N142, N136, N93, N122, N103);
xor XOR2 (N143, N131, N89);
xor XOR2 (N144, N142, N112);
buf BUF1 (N145, N141);
nand NAND2 (N146, N130, N60);
xor XOR2 (N147, N129, N73);
xor XOR2 (N148, N139, N27);
or OR4 (N149, N145, N114, N16, N133);
nor NOR4 (N150, N102, N118, N61, N39);
xor XOR2 (N151, N143, N47);
and AND2 (N152, N146, N93);
buf BUF1 (N153, N151);
not NOT1 (N154, N149);
nand NAND2 (N155, N147, N126);
not NOT1 (N156, N155);
or OR4 (N157, N140, N14, N83, N25);
buf BUF1 (N158, N144);
nand NAND3 (N159, N152, N91, N91);
xor XOR2 (N160, N157, N88);
xor XOR2 (N161, N160, N136);
not NOT1 (N162, N138);
nand NAND3 (N163, N150, N42, N159);
or OR3 (N164, N105, N119, N73);
and AND3 (N165, N134, N24, N35);
and AND2 (N166, N158, N134);
nand NAND3 (N167, N156, N33, N139);
nor NOR2 (N168, N164, N128);
nand NAND2 (N169, N166, N99);
buf BUF1 (N170, N162);
and AND4 (N171, N148, N134, N135, N73);
buf BUF1 (N172, N153);
or OR4 (N173, N172, N159, N46, N49);
not NOT1 (N174, N171);
not NOT1 (N175, N173);
not NOT1 (N176, N163);
or OR4 (N177, N174, N160, N127, N172);
nor NOR2 (N178, N168, N40);
nand NAND4 (N179, N170, N105, N107, N72);
buf BUF1 (N180, N154);
buf BUF1 (N181, N176);
nor NOR3 (N182, N161, N38, N137);
nand NAND4 (N183, N167, N10, N89, N29);
nand NAND4 (N184, N181, N53, N13, N82);
not NOT1 (N185, N175);
not NOT1 (N186, N184);
nand NAND4 (N187, N182, N8, N30, N83);
nor NOR3 (N188, N183, N90, N115);
or OR4 (N189, N188, N84, N168, N50);
or OR4 (N190, N178, N129, N172, N130);
buf BUF1 (N191, N187);
and AND3 (N192, N165, N87, N33);
not NOT1 (N193, N169);
or OR2 (N194, N179, N147);
buf BUF1 (N195, N191);
nor NOR4 (N196, N190, N191, N30, N59);
or OR4 (N197, N194, N28, N176, N76);
and AND4 (N198, N195, N115, N90, N55);
or OR2 (N199, N186, N98);
buf BUF1 (N200, N177);
nor NOR2 (N201, N189, N8);
xor XOR2 (N202, N180, N127);
xor XOR2 (N203, N196, N103);
nor NOR2 (N204, N199, N12);
nand NAND4 (N205, N200, N95, N94, N115);
or OR3 (N206, N205, N99, N109);
or OR2 (N207, N193, N64);
buf BUF1 (N208, N185);
nand NAND2 (N209, N192, N197);
nand NAND3 (N210, N204, N26, N80);
buf BUF1 (N211, N11);
or OR3 (N212, N203, N66, N35);
or OR4 (N213, N211, N59, N13, N43);
and AND3 (N214, N209, N194, N198);
not NOT1 (N215, N182);
or OR3 (N216, N207, N20, N6);
nand NAND2 (N217, N212, N45);
xor XOR2 (N218, N217, N7);
or OR3 (N219, N218, N214, N10);
xor XOR2 (N220, N157, N102);
xor XOR2 (N221, N210, N91);
and AND4 (N222, N220, N9, N143, N49);
and AND2 (N223, N213, N143);
xor XOR2 (N224, N221, N69);
buf BUF1 (N225, N208);
and AND4 (N226, N223, N72, N89, N14);
and AND3 (N227, N202, N142, N204);
nor NOR2 (N228, N206, N92);
and AND3 (N229, N222, N220, N165);
not NOT1 (N230, N201);
not NOT1 (N231, N224);
and AND2 (N232, N227, N141);
nor NOR4 (N233, N215, N118, N84, N114);
xor XOR2 (N234, N219, N40);
nand NAND4 (N235, N233, N120, N106, N12);
not NOT1 (N236, N230);
nor NOR2 (N237, N235, N154);
or OR2 (N238, N234, N195);
buf BUF1 (N239, N238);
and AND2 (N240, N216, N141);
nor NOR4 (N241, N229, N14, N236, N19);
xor XOR2 (N242, N100, N235);
buf BUF1 (N243, N237);
or OR2 (N244, N231, N95);
buf BUF1 (N245, N240);
nor NOR4 (N246, N228, N230, N114, N17);
nand NAND3 (N247, N225, N141, N138);
xor XOR2 (N248, N242, N145);
and AND4 (N249, N232, N219, N6, N233);
not NOT1 (N250, N247);
nand NAND2 (N251, N246, N91);
or OR2 (N252, N249, N225);
nand NAND4 (N253, N248, N173, N150, N149);
and AND3 (N254, N226, N103, N222);
nor NOR2 (N255, N241, N215);
nand NAND3 (N256, N251, N181, N61);
not NOT1 (N257, N250);
xor XOR2 (N258, N243, N92);
nor NOR3 (N259, N253, N101, N204);
or OR4 (N260, N256, N243, N16, N231);
buf BUF1 (N261, N245);
nand NAND3 (N262, N244, N244, N195);
not NOT1 (N263, N255);
or OR2 (N264, N239, N45);
or OR4 (N265, N262, N39, N136, N20);
xor XOR2 (N266, N263, N20);
nand NAND3 (N267, N252, N129, N231);
and AND3 (N268, N265, N173, N97);
buf BUF1 (N269, N267);
or OR3 (N270, N264, N3, N180);
xor XOR2 (N271, N254, N10);
nand NAND4 (N272, N257, N27, N264, N102);
nand NAND2 (N273, N268, N173);
or OR4 (N274, N261, N244, N1, N70);
or OR2 (N275, N273, N99);
not NOT1 (N276, N275);
nor NOR3 (N277, N272, N227, N32);
and AND3 (N278, N277, N253, N57);
or OR2 (N279, N270, N232);
xor XOR2 (N280, N260, N56);
buf BUF1 (N281, N271);
and AND4 (N282, N259, N147, N114, N57);
buf BUF1 (N283, N278);
and AND2 (N284, N258, N90);
nor NOR3 (N285, N269, N188, N69);
or OR3 (N286, N282, N243, N264);
not NOT1 (N287, N266);
or OR4 (N288, N281, N98, N38, N206);
buf BUF1 (N289, N276);
and AND2 (N290, N286, N62);
nand NAND4 (N291, N289, N98, N106, N73);
not NOT1 (N292, N291);
nand NAND2 (N293, N279, N285);
and AND4 (N294, N115, N103, N74, N209);
not NOT1 (N295, N287);
nand NAND2 (N296, N284, N292);
nor NOR4 (N297, N108, N130, N100, N211);
not NOT1 (N298, N290);
nand NAND2 (N299, N295, N266);
or OR4 (N300, N297, N251, N120, N159);
xor XOR2 (N301, N300, N243);
nor NOR4 (N302, N298, N160, N29, N16);
or OR4 (N303, N293, N115, N112, N222);
nor NOR3 (N304, N283, N280, N150);
not NOT1 (N305, N260);
or OR3 (N306, N274, N261, N46);
nand NAND2 (N307, N301, N133);
xor XOR2 (N308, N288, N171);
and AND2 (N309, N296, N275);
not NOT1 (N310, N305);
nand NAND2 (N311, N304, N69);
or OR2 (N312, N302, N36);
nand NAND2 (N313, N303, N267);
xor XOR2 (N314, N310, N196);
nor NOR3 (N315, N308, N166, N140);
nor NOR4 (N316, N311, N15, N100, N286);
xor XOR2 (N317, N299, N215);
and AND4 (N318, N309, N96, N30, N266);
buf BUF1 (N319, N317);
nor NOR4 (N320, N314, N72, N111, N151);
nand NAND4 (N321, N306, N184, N176, N245);
or OR2 (N322, N320, N199);
xor XOR2 (N323, N315, N216);
not NOT1 (N324, N307);
xor XOR2 (N325, N321, N264);
not NOT1 (N326, N294);
or OR2 (N327, N316, N35);
nand NAND3 (N328, N325, N80, N41);
nand NAND2 (N329, N324, N16);
buf BUF1 (N330, N329);
xor XOR2 (N331, N330, N230);
or OR4 (N332, N323, N77, N231, N165);
or OR3 (N333, N318, N175, N46);
not NOT1 (N334, N331);
buf BUF1 (N335, N333);
or OR4 (N336, N334, N79, N238, N110);
or OR3 (N337, N336, N116, N188);
and AND2 (N338, N322, N2);
nor NOR3 (N339, N326, N42, N16);
nand NAND2 (N340, N327, N32);
nor NOR4 (N341, N313, N179, N92, N161);
buf BUF1 (N342, N339);
or OR4 (N343, N335, N156, N39, N35);
or OR4 (N344, N328, N120, N119, N262);
buf BUF1 (N345, N343);
and AND2 (N346, N312, N153);
nand NAND3 (N347, N340, N37, N227);
nand NAND2 (N348, N338, N253);
or OR2 (N349, N342, N282);
nor NOR4 (N350, N341, N245, N86, N221);
or OR2 (N351, N350, N187);
nand NAND3 (N352, N346, N131, N56);
nor NOR3 (N353, N348, N149, N137);
and AND2 (N354, N319, N128);
and AND4 (N355, N345, N274, N129, N39);
and AND3 (N356, N352, N178, N48);
and AND3 (N357, N332, N220, N298);
buf BUF1 (N358, N349);
buf BUF1 (N359, N351);
or OR4 (N360, N354, N87, N154, N98);
or OR4 (N361, N357, N201, N325, N240);
and AND2 (N362, N359, N154);
nand NAND4 (N363, N337, N13, N169, N196);
xor XOR2 (N364, N353, N15);
xor XOR2 (N365, N360, N342);
xor XOR2 (N366, N344, N113);
nand NAND4 (N367, N361, N123, N4, N293);
or OR3 (N368, N358, N152, N238);
buf BUF1 (N369, N368);
nand NAND2 (N370, N355, N277);
buf BUF1 (N371, N347);
xor XOR2 (N372, N363, N128);
nand NAND4 (N373, N369, N123, N206, N325);
xor XOR2 (N374, N367, N362);
not NOT1 (N375, N84);
buf BUF1 (N376, N370);
and AND2 (N377, N371, N204);
xor XOR2 (N378, N365, N146);
xor XOR2 (N379, N366, N163);
xor XOR2 (N380, N379, N267);
buf BUF1 (N381, N377);
xor XOR2 (N382, N376, N216);
not NOT1 (N383, N372);
nand NAND3 (N384, N381, N89, N99);
xor XOR2 (N385, N384, N202);
xor XOR2 (N386, N380, N65);
buf BUF1 (N387, N373);
nand NAND4 (N388, N386, N203, N16, N348);
nand NAND4 (N389, N388, N73, N231, N298);
nor NOR4 (N390, N383, N284, N316, N31);
buf BUF1 (N391, N387);
nand NAND2 (N392, N391, N381);
or OR2 (N393, N364, N215);
xor XOR2 (N394, N392, N340);
and AND4 (N395, N385, N138, N69, N278);
nand NAND4 (N396, N394, N90, N24, N189);
and AND4 (N397, N382, N278, N392, N356);
and AND2 (N398, N44, N331);
and AND4 (N399, N389, N83, N204, N92);
and AND4 (N400, N396, N332, N105, N62);
not NOT1 (N401, N393);
or OR4 (N402, N401, N300, N170, N310);
buf BUF1 (N403, N374);
and AND4 (N404, N378, N304, N217, N332);
buf BUF1 (N405, N402);
xor XOR2 (N406, N397, N358);
and AND3 (N407, N403, N85, N378);
or OR2 (N408, N405, N156);
buf BUF1 (N409, N406);
not NOT1 (N410, N409);
buf BUF1 (N411, N375);
buf BUF1 (N412, N400);
or OR3 (N413, N395, N85, N250);
nand NAND2 (N414, N407, N289);
nor NOR4 (N415, N414, N74, N47, N92);
nand NAND3 (N416, N411, N3, N264);
nand NAND4 (N417, N398, N249, N348, N218);
nand NAND2 (N418, N408, N179);
nor NOR3 (N419, N417, N17, N393);
nor NOR4 (N420, N415, N317, N295, N340);
or OR4 (N421, N399, N44, N180, N203);
nor NOR4 (N422, N413, N274, N309, N184);
or OR4 (N423, N422, N341, N373, N28);
xor XOR2 (N424, N421, N220);
not NOT1 (N425, N404);
and AND4 (N426, N416, N323, N235, N112);
and AND4 (N427, N420, N235, N50, N354);
nor NOR2 (N428, N424, N100);
and AND3 (N429, N423, N271, N339);
nor NOR4 (N430, N429, N269, N270, N163);
or OR3 (N431, N425, N297, N59);
and AND4 (N432, N410, N404, N250, N132);
or OR2 (N433, N412, N137);
nor NOR2 (N434, N433, N286);
nand NAND2 (N435, N430, N356);
not NOT1 (N436, N418);
nor NOR2 (N437, N436, N58);
nand NAND3 (N438, N431, N254, N242);
not NOT1 (N439, N428);
and AND3 (N440, N434, N106, N355);
buf BUF1 (N441, N439);
nand NAND2 (N442, N432, N70);
buf BUF1 (N443, N442);
nor NOR3 (N444, N440, N55, N179);
and AND2 (N445, N437, N107);
buf BUF1 (N446, N435);
or OR2 (N447, N443, N214);
buf BUF1 (N448, N427);
nand NAND2 (N449, N426, N377);
nand NAND4 (N450, N444, N438, N326, N306);
or OR2 (N451, N382, N233);
not NOT1 (N452, N448);
and AND4 (N453, N449, N171, N430, N180);
buf BUF1 (N454, N450);
nand NAND2 (N455, N445, N212);
nor NOR4 (N456, N454, N286, N356, N136);
nor NOR3 (N457, N455, N85, N311);
and AND4 (N458, N451, N421, N62, N89);
nand NAND2 (N459, N457, N329);
or OR4 (N460, N390, N295, N358, N295);
buf BUF1 (N461, N419);
nor NOR3 (N462, N452, N224, N194);
nor NOR3 (N463, N453, N395, N283);
nand NAND4 (N464, N456, N177, N298, N42);
and AND2 (N465, N464, N98);
buf BUF1 (N466, N461);
and AND4 (N467, N462, N344, N40, N18);
xor XOR2 (N468, N446, N22);
not NOT1 (N469, N463);
nand NAND4 (N470, N465, N22, N254, N252);
buf BUF1 (N471, N468);
buf BUF1 (N472, N458);
nand NAND4 (N473, N472, N50, N107, N2);
nor NOR3 (N474, N459, N364, N150);
xor XOR2 (N475, N447, N360);
buf BUF1 (N476, N467);
nand NAND4 (N477, N441, N250, N19, N68);
nand NAND4 (N478, N473, N22, N155, N368);
and AND2 (N479, N460, N377);
or OR4 (N480, N475, N129, N202, N347);
nand NAND3 (N481, N474, N385, N87);
or OR4 (N482, N480, N245, N340, N44);
and AND2 (N483, N479, N8);
or OR2 (N484, N477, N368);
or OR3 (N485, N469, N205, N224);
not NOT1 (N486, N470);
or OR2 (N487, N466, N236);
nand NAND4 (N488, N487, N477, N452, N427);
nand NAND3 (N489, N484, N37, N261);
not NOT1 (N490, N486);
or OR4 (N491, N481, N40, N226, N216);
xor XOR2 (N492, N490, N274);
nor NOR4 (N493, N476, N194, N196, N199);
buf BUF1 (N494, N482);
not NOT1 (N495, N478);
not NOT1 (N496, N485);
nand NAND3 (N497, N471, N104, N220);
and AND3 (N498, N496, N165, N227);
nand NAND3 (N499, N498, N258, N274);
not NOT1 (N500, N497);
and AND2 (N501, N488, N415);
nor NOR3 (N502, N492, N241, N72);
xor XOR2 (N503, N491, N238);
and AND2 (N504, N500, N111);
buf BUF1 (N505, N502);
and AND2 (N506, N503, N48);
and AND2 (N507, N499, N322);
nand NAND2 (N508, N493, N446);
nand NAND2 (N509, N483, N414);
not NOT1 (N510, N504);
nand NAND4 (N511, N510, N309, N47, N222);
and AND3 (N512, N506, N112, N426);
nand NAND2 (N513, N509, N162);
or OR4 (N514, N494, N294, N111, N196);
or OR3 (N515, N505, N324, N242);
or OR4 (N516, N507, N148, N174, N95);
nand NAND3 (N517, N501, N355, N349);
not NOT1 (N518, N511);
nor NOR3 (N519, N517, N138, N432);
nand NAND2 (N520, N514, N133);
or OR4 (N521, N519, N92, N163, N379);
and AND3 (N522, N516, N57, N298);
nand NAND4 (N523, N512, N369, N499, N153);
buf BUF1 (N524, N515);
not NOT1 (N525, N520);
xor XOR2 (N526, N521, N215);
and AND4 (N527, N495, N247, N518, N398);
xor XOR2 (N528, N69, N444);
xor XOR2 (N529, N526, N347);
xor XOR2 (N530, N522, N151);
or OR2 (N531, N508, N519);
and AND4 (N532, N531, N507, N66, N451);
xor XOR2 (N533, N532, N169);
not NOT1 (N534, N523);
nor NOR3 (N535, N534, N20, N156);
or OR2 (N536, N530, N335);
nand NAND3 (N537, N525, N196, N409);
nand NAND3 (N538, N524, N352, N432);
or OR2 (N539, N537, N370);
and AND3 (N540, N513, N462, N357);
nand NAND3 (N541, N529, N407, N335);
and AND4 (N542, N533, N260, N137, N269);
or OR2 (N543, N542, N395);
xor XOR2 (N544, N489, N445);
nand NAND3 (N545, N535, N284, N321);
buf BUF1 (N546, N536);
or OR3 (N547, N545, N199, N11);
not NOT1 (N548, N543);
and AND3 (N549, N541, N341, N390);
or OR2 (N550, N528, N133);
not NOT1 (N551, N546);
and AND3 (N552, N540, N166, N326);
xor XOR2 (N553, N527, N126);
nand NAND2 (N554, N544, N99);
buf BUF1 (N555, N551);
buf BUF1 (N556, N539);
and AND3 (N557, N549, N506, N174);
buf BUF1 (N558, N554);
xor XOR2 (N559, N550, N546);
nor NOR3 (N560, N558, N494, N210);
xor XOR2 (N561, N556, N288);
nor NOR2 (N562, N538, N450);
xor XOR2 (N563, N553, N33);
xor XOR2 (N564, N559, N46);
not NOT1 (N565, N547);
buf BUF1 (N566, N552);
or OR2 (N567, N563, N308);
or OR4 (N568, N567, N508, N51, N471);
xor XOR2 (N569, N561, N379);
not NOT1 (N570, N548);
nand NAND2 (N571, N564, N235);
and AND2 (N572, N566, N135);
and AND3 (N573, N570, N212, N332);
not NOT1 (N574, N571);
or OR4 (N575, N572, N528, N253, N170);
xor XOR2 (N576, N562, N487);
buf BUF1 (N577, N574);
and AND2 (N578, N575, N294);
and AND4 (N579, N569, N11, N410, N336);
or OR3 (N580, N577, N130, N261);
xor XOR2 (N581, N576, N185);
buf BUF1 (N582, N579);
nor NOR4 (N583, N555, N347, N530, N459);
not NOT1 (N584, N560);
and AND4 (N585, N580, N188, N396, N489);
nand NAND2 (N586, N583, N158);
not NOT1 (N587, N568);
buf BUF1 (N588, N585);
xor XOR2 (N589, N557, N41);
nand NAND2 (N590, N578, N525);
nor NOR3 (N591, N565, N59, N574);
xor XOR2 (N592, N590, N86);
buf BUF1 (N593, N573);
or OR2 (N594, N589, N586);
nor NOR3 (N595, N309, N218, N373);
not NOT1 (N596, N581);
xor XOR2 (N597, N592, N219);
nand NAND3 (N598, N597, N524, N215);
not NOT1 (N599, N596);
not NOT1 (N600, N593);
or OR3 (N601, N595, N496, N365);
nor NOR2 (N602, N600, N521);
and AND2 (N603, N582, N70);
nor NOR2 (N604, N587, N457);
and AND3 (N605, N588, N543, N11);
nand NAND2 (N606, N601, N344);
and AND2 (N607, N606, N319);
or OR3 (N608, N584, N109, N156);
and AND3 (N609, N599, N130, N540);
or OR4 (N610, N602, N359, N279, N558);
nand NAND3 (N611, N598, N402, N226);
buf BUF1 (N612, N608);
xor XOR2 (N613, N607, N609);
or OR4 (N614, N150, N379, N355, N325);
nand NAND2 (N615, N604, N226);
nor NOR2 (N616, N605, N421);
xor XOR2 (N617, N591, N231);
buf BUF1 (N618, N615);
and AND3 (N619, N614, N443, N565);
buf BUF1 (N620, N603);
nand NAND2 (N621, N617, N266);
nand NAND3 (N622, N611, N86, N542);
nand NAND4 (N623, N616, N328, N395, N213);
and AND3 (N624, N620, N211, N410);
buf BUF1 (N625, N610);
nor NOR3 (N626, N613, N86, N356);
nand NAND3 (N627, N626, N308, N39);
nor NOR4 (N628, N594, N436, N590, N194);
xor XOR2 (N629, N612, N79);
nor NOR2 (N630, N621, N591);
nor NOR2 (N631, N630, N333);
and AND2 (N632, N622, N558);
not NOT1 (N633, N627);
nand NAND2 (N634, N631, N366);
and AND4 (N635, N623, N147, N569, N93);
or OR4 (N636, N618, N527, N353, N557);
nand NAND4 (N637, N633, N226, N34, N110);
buf BUF1 (N638, N624);
xor XOR2 (N639, N634, N120);
and AND2 (N640, N619, N506);
and AND2 (N641, N629, N19);
xor XOR2 (N642, N638, N392);
buf BUF1 (N643, N635);
nand NAND4 (N644, N642, N597, N586, N438);
or OR3 (N645, N632, N286, N228);
nand NAND4 (N646, N641, N315, N217, N572);
xor XOR2 (N647, N628, N500);
or OR4 (N648, N636, N422, N540, N575);
nand NAND4 (N649, N637, N147, N120, N336);
nand NAND3 (N650, N643, N131, N499);
or OR3 (N651, N639, N441, N539);
and AND3 (N652, N650, N334, N209);
nor NOR2 (N653, N649, N646);
or OR2 (N654, N250, N607);
nor NOR4 (N655, N645, N433, N375, N595);
not NOT1 (N656, N652);
and AND3 (N657, N653, N486, N369);
or OR4 (N658, N625, N375, N619, N397);
nand NAND4 (N659, N656, N611, N591, N639);
or OR4 (N660, N655, N113, N582, N378);
not NOT1 (N661, N651);
xor XOR2 (N662, N658, N405);
xor XOR2 (N663, N648, N533);
xor XOR2 (N664, N640, N156);
nor NOR4 (N665, N657, N575, N370, N603);
xor XOR2 (N666, N647, N59);
and AND3 (N667, N660, N68, N624);
nand NAND3 (N668, N663, N260, N106);
xor XOR2 (N669, N654, N354);
nor NOR4 (N670, N664, N348, N226, N346);
not NOT1 (N671, N670);
and AND4 (N672, N666, N479, N563, N417);
and AND2 (N673, N672, N271);
nand NAND3 (N674, N644, N549, N303);
xor XOR2 (N675, N661, N509);
nand NAND2 (N676, N668, N327);
nand NAND2 (N677, N667, N204);
xor XOR2 (N678, N659, N630);
not NOT1 (N679, N673);
xor XOR2 (N680, N674, N81);
xor XOR2 (N681, N678, N60);
not NOT1 (N682, N680);
or OR2 (N683, N679, N16);
or OR2 (N684, N665, N673);
not NOT1 (N685, N671);
xor XOR2 (N686, N685, N156);
nand NAND4 (N687, N662, N438, N377, N175);
xor XOR2 (N688, N683, N368);
or OR3 (N689, N676, N128, N19);
nand NAND3 (N690, N669, N398, N521);
nor NOR2 (N691, N688, N359);
or OR3 (N692, N675, N539, N515);
not NOT1 (N693, N689);
nor NOR3 (N694, N690, N510, N380);
nand NAND2 (N695, N684, N118);
xor XOR2 (N696, N687, N665);
buf BUF1 (N697, N695);
xor XOR2 (N698, N693, N125);
xor XOR2 (N699, N696, N197);
or OR2 (N700, N682, N654);
or OR3 (N701, N686, N291, N468);
nor NOR3 (N702, N701, N364, N658);
not NOT1 (N703, N681);
or OR3 (N704, N691, N328, N117);
or OR4 (N705, N692, N539, N385, N437);
nor NOR4 (N706, N704, N676, N705, N3);
xor XOR2 (N707, N350, N598);
or OR4 (N708, N697, N165, N334, N172);
xor XOR2 (N709, N703, N351);
and AND2 (N710, N709, N668);
nor NOR2 (N711, N702, N370);
buf BUF1 (N712, N711);
or OR3 (N713, N677, N583, N90);
nand NAND2 (N714, N700, N316);
not NOT1 (N715, N707);
nor NOR2 (N716, N710, N387);
buf BUF1 (N717, N712);
xor XOR2 (N718, N717, N163);
nor NOR4 (N719, N714, N705, N583, N422);
not NOT1 (N720, N716);
buf BUF1 (N721, N718);
nand NAND3 (N722, N721, N120, N148);
buf BUF1 (N723, N719);
nor NOR2 (N724, N694, N169);
or OR4 (N725, N715, N533, N47, N686);
or OR2 (N726, N698, N116);
buf BUF1 (N727, N708);
and AND4 (N728, N713, N318, N143, N596);
nor NOR3 (N729, N724, N410, N173);
buf BUF1 (N730, N720);
buf BUF1 (N731, N728);
nor NOR2 (N732, N731, N260);
not NOT1 (N733, N730);
or OR4 (N734, N727, N266, N466, N314);
buf BUF1 (N735, N723);
nor NOR3 (N736, N706, N585, N508);
nand NAND4 (N737, N699, N329, N118, N634);
xor XOR2 (N738, N736, N93);
buf BUF1 (N739, N734);
nor NOR4 (N740, N739, N727, N248, N510);
nor NOR4 (N741, N740, N215, N456, N469);
nor NOR3 (N742, N733, N110, N663);
nor NOR3 (N743, N729, N344, N337);
not NOT1 (N744, N741);
or OR4 (N745, N735, N248, N142, N243);
and AND3 (N746, N725, N441, N144);
and AND4 (N747, N726, N4, N138, N745);
nand NAND4 (N748, N364, N642, N154, N535);
nand NAND4 (N749, N738, N67, N693, N631);
nand NAND2 (N750, N744, N13);
or OR2 (N751, N746, N466);
and AND4 (N752, N732, N137, N100, N87);
or OR3 (N753, N751, N233, N277);
xor XOR2 (N754, N750, N594);
nand NAND3 (N755, N748, N96, N63);
nand NAND4 (N756, N743, N298, N341, N714);
nor NOR4 (N757, N742, N643, N334, N61);
nor NOR3 (N758, N753, N101, N651);
nor NOR2 (N759, N747, N111);
nand NAND2 (N760, N756, N179);
xor XOR2 (N761, N722, N20);
nand NAND3 (N762, N758, N159, N33);
or OR4 (N763, N761, N280, N31, N382);
or OR2 (N764, N762, N126);
xor XOR2 (N765, N764, N736);
or OR4 (N766, N759, N381, N167, N636);
nand NAND3 (N767, N766, N765, N317);
or OR2 (N768, N599, N156);
buf BUF1 (N769, N755);
and AND3 (N770, N752, N26, N733);
or OR4 (N771, N767, N623, N354, N675);
nor NOR2 (N772, N757, N224);
or OR3 (N773, N737, N119, N449);
not NOT1 (N774, N769);
nor NOR3 (N775, N774, N163, N464);
buf BUF1 (N776, N773);
and AND2 (N777, N771, N711);
buf BUF1 (N778, N749);
nand NAND2 (N779, N772, N503);
buf BUF1 (N780, N763);
and AND3 (N781, N780, N724, N693);
not NOT1 (N782, N770);
nand NAND3 (N783, N777, N138, N346);
nand NAND2 (N784, N768, N708);
nand NAND2 (N785, N781, N402);
or OR2 (N786, N776, N654);
nor NOR3 (N787, N760, N80, N207);
or OR3 (N788, N775, N565, N353);
xor XOR2 (N789, N787, N589);
or OR4 (N790, N754, N361, N20, N690);
nor NOR3 (N791, N785, N447, N363);
buf BUF1 (N792, N783);
and AND4 (N793, N779, N729, N162, N14);
not NOT1 (N794, N789);
nand NAND2 (N795, N786, N534);
or OR3 (N796, N792, N300, N579);
and AND3 (N797, N796, N292, N136);
or OR3 (N798, N782, N131, N84);
xor XOR2 (N799, N790, N401);
nand NAND3 (N800, N795, N748, N347);
or OR2 (N801, N784, N246);
and AND4 (N802, N798, N361, N431, N490);
nor NOR3 (N803, N791, N732, N266);
xor XOR2 (N804, N788, N147);
nand NAND2 (N805, N799, N356);
buf BUF1 (N806, N794);
and AND3 (N807, N802, N621, N537);
and AND2 (N808, N793, N1);
and AND4 (N809, N808, N792, N128, N276);
xor XOR2 (N810, N801, N536);
or OR4 (N811, N810, N405, N184, N410);
endmodule