// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N881,N893,N899,N904,N908,N905,N907,N909,N897,N910;

not NOT1 (N11, N8);
xor XOR2 (N12, N1, N5);
nor NOR3 (N13, N9, N9, N1);
xor XOR2 (N14, N6, N7);
or OR2 (N15, N11, N12);
or OR3 (N16, N1, N6, N12);
not NOT1 (N17, N11);
nor NOR2 (N18, N14, N14);
xor XOR2 (N19, N9, N11);
or OR2 (N20, N8, N19);
buf BUF1 (N21, N2);
and AND4 (N22, N21, N14, N11, N9);
buf BUF1 (N23, N18);
xor XOR2 (N24, N1, N18);
nor NOR4 (N25, N13, N24, N14, N6);
and AND2 (N26, N14, N17);
or OR4 (N27, N20, N23, N20, N1);
and AND2 (N28, N25, N2);
nand NAND2 (N29, N19, N2);
nor NOR2 (N30, N16, N29);
xor XOR2 (N31, N4, N9);
nand NAND3 (N32, N9, N10, N10);
nand NAND2 (N33, N6, N31);
or OR2 (N34, N19, N25);
buf BUF1 (N35, N23);
or OR2 (N36, N34, N17);
or OR3 (N37, N15, N33, N13);
nor NOR3 (N38, N26, N26, N7);
xor XOR2 (N39, N23, N24);
buf BUF1 (N40, N39);
buf BUF1 (N41, N27);
or OR3 (N42, N35, N23, N27);
buf BUF1 (N43, N28);
and AND2 (N44, N32, N19);
or OR4 (N45, N40, N31, N41, N33);
or OR2 (N46, N28, N16);
buf BUF1 (N47, N44);
or OR3 (N48, N30, N3, N27);
xor XOR2 (N49, N48, N26);
nor NOR2 (N50, N43, N4);
nor NOR2 (N51, N38, N50);
and AND4 (N52, N32, N48, N38, N39);
or OR2 (N53, N37, N12);
nor NOR3 (N54, N22, N6, N28);
or OR3 (N55, N42, N8, N53);
xor XOR2 (N56, N52, N6);
and AND4 (N57, N20, N15, N29, N47);
nor NOR4 (N58, N57, N12, N54, N48);
or OR2 (N59, N19, N54);
or OR4 (N60, N14, N30, N48, N40);
or OR2 (N61, N60, N59);
nor NOR4 (N62, N1, N42, N18, N23);
buf BUF1 (N63, N36);
nor NOR2 (N64, N61, N58);
nand NAND2 (N65, N35, N61);
nor NOR3 (N66, N45, N44, N52);
nor NOR2 (N67, N56, N9);
nor NOR3 (N68, N51, N8, N16);
and AND4 (N69, N67, N54, N45, N67);
buf BUF1 (N70, N68);
nor NOR3 (N71, N70, N17, N28);
nor NOR4 (N72, N66, N14, N52, N27);
xor XOR2 (N73, N49, N18);
xor XOR2 (N74, N71, N51);
and AND2 (N75, N62, N35);
nor NOR3 (N76, N74, N70, N62);
and AND3 (N77, N69, N69, N7);
nand NAND2 (N78, N76, N36);
not NOT1 (N79, N65);
not NOT1 (N80, N46);
and AND4 (N81, N75, N51, N35, N41);
nor NOR4 (N82, N63, N14, N65, N56);
not NOT1 (N83, N80);
not NOT1 (N84, N77);
xor XOR2 (N85, N84, N40);
and AND2 (N86, N73, N34);
buf BUF1 (N87, N64);
nand NAND4 (N88, N55, N18, N64, N35);
or OR3 (N89, N81, N3, N66);
nand NAND2 (N90, N85, N33);
nand NAND2 (N91, N90, N53);
xor XOR2 (N92, N83, N60);
or OR4 (N93, N87, N4, N47, N17);
xor XOR2 (N94, N86, N50);
buf BUF1 (N95, N92);
or OR4 (N96, N89, N33, N56, N90);
and AND2 (N97, N91, N45);
xor XOR2 (N98, N95, N4);
not NOT1 (N99, N94);
and AND2 (N100, N78, N84);
and AND2 (N101, N82, N55);
nor NOR2 (N102, N93, N30);
nor NOR4 (N103, N97, N99, N83, N44);
nor NOR3 (N104, N67, N3, N37);
not NOT1 (N105, N98);
or OR4 (N106, N96, N16, N50, N48);
not NOT1 (N107, N100);
not NOT1 (N108, N107);
buf BUF1 (N109, N104);
nand NAND2 (N110, N105, N86);
and AND4 (N111, N103, N23, N97, N110);
buf BUF1 (N112, N34);
or OR2 (N113, N111, N59);
not NOT1 (N114, N109);
nor NOR2 (N115, N72, N96);
not NOT1 (N116, N102);
nor NOR4 (N117, N112, N32, N98, N11);
not NOT1 (N118, N115);
xor XOR2 (N119, N114, N45);
and AND4 (N120, N101, N8, N83, N112);
or OR3 (N121, N79, N107, N28);
xor XOR2 (N122, N121, N91);
nor NOR2 (N123, N113, N20);
xor XOR2 (N124, N119, N89);
or OR4 (N125, N124, N48, N94, N65);
nor NOR2 (N126, N117, N49);
xor XOR2 (N127, N116, N77);
not NOT1 (N128, N123);
buf BUF1 (N129, N126);
nand NAND4 (N130, N120, N67, N97, N73);
buf BUF1 (N131, N108);
and AND3 (N132, N122, N126, N93);
nand NAND3 (N133, N118, N124, N73);
nand NAND4 (N134, N132, N17, N14, N9);
or OR3 (N135, N133, N43, N22);
and AND3 (N136, N127, N99, N12);
xor XOR2 (N137, N128, N100);
not NOT1 (N138, N129);
and AND2 (N139, N131, N20);
or OR2 (N140, N139, N91);
or OR4 (N141, N140, N115, N17, N50);
xor XOR2 (N142, N134, N141);
and AND3 (N143, N124, N22, N61);
nand NAND2 (N144, N142, N92);
not NOT1 (N145, N88);
buf BUF1 (N146, N136);
nand NAND4 (N147, N138, N37, N70, N39);
or OR3 (N148, N143, N83, N116);
xor XOR2 (N149, N146, N53);
not NOT1 (N150, N145);
not NOT1 (N151, N147);
or OR2 (N152, N135, N90);
nor NOR2 (N153, N137, N71);
nor NOR2 (N154, N148, N82);
nand NAND2 (N155, N149, N87);
not NOT1 (N156, N106);
and AND4 (N157, N152, N146, N42, N100);
buf BUF1 (N158, N156);
nor NOR2 (N159, N154, N43);
or OR2 (N160, N157, N100);
not NOT1 (N161, N151);
or OR4 (N162, N158, N134, N33, N76);
not NOT1 (N163, N160);
and AND3 (N164, N155, N100, N150);
or OR2 (N165, N4, N141);
buf BUF1 (N166, N159);
not NOT1 (N167, N165);
xor XOR2 (N168, N164, N166);
or OR4 (N169, N141, N21, N35, N161);
nor NOR4 (N170, N127, N61, N75, N4);
xor XOR2 (N171, N167, N102);
and AND2 (N172, N130, N158);
buf BUF1 (N173, N169);
xor XOR2 (N174, N172, N23);
nor NOR4 (N175, N162, N136, N149, N92);
not NOT1 (N176, N125);
not NOT1 (N177, N173);
nand NAND2 (N178, N176, N91);
not NOT1 (N179, N171);
and AND2 (N180, N144, N46);
not NOT1 (N181, N153);
nand NAND2 (N182, N163, N160);
nor NOR2 (N183, N179, N93);
and AND3 (N184, N175, N114, N81);
and AND2 (N185, N177, N165);
buf BUF1 (N186, N178);
and AND3 (N187, N180, N46, N8);
or OR3 (N188, N170, N50, N22);
xor XOR2 (N189, N186, N27);
nand NAND4 (N190, N168, N70, N10, N9);
not NOT1 (N191, N174);
nand NAND3 (N192, N187, N58, N54);
and AND3 (N193, N182, N161, N3);
nand NAND2 (N194, N191, N168);
xor XOR2 (N195, N189, N186);
buf BUF1 (N196, N195);
nand NAND2 (N197, N196, N8);
or OR4 (N198, N183, N46, N55, N132);
and AND2 (N199, N190, N16);
buf BUF1 (N200, N194);
or OR2 (N201, N193, N167);
or OR4 (N202, N185, N173, N40, N137);
nand NAND2 (N203, N199, N40);
not NOT1 (N204, N181);
xor XOR2 (N205, N204, N185);
xor XOR2 (N206, N184, N122);
buf BUF1 (N207, N197);
xor XOR2 (N208, N205, N146);
or OR4 (N209, N200, N126, N180, N192);
not NOT1 (N210, N203);
nor NOR2 (N211, N50, N125);
xor XOR2 (N212, N188, N99);
or OR3 (N213, N211, N207, N61);
not NOT1 (N214, N154);
buf BUF1 (N215, N214);
buf BUF1 (N216, N213);
nand NAND2 (N217, N202, N39);
nand NAND3 (N218, N201, N32, N52);
xor XOR2 (N219, N208, N100);
nand NAND3 (N220, N209, N28, N75);
nand NAND3 (N221, N218, N204, N10);
nand NAND2 (N222, N216, N178);
not NOT1 (N223, N206);
or OR4 (N224, N215, N10, N184, N44);
xor XOR2 (N225, N212, N118);
buf BUF1 (N226, N198);
not NOT1 (N227, N226);
not NOT1 (N228, N220);
nand NAND2 (N229, N217, N20);
buf BUF1 (N230, N228);
xor XOR2 (N231, N229, N91);
xor XOR2 (N232, N221, N35);
buf BUF1 (N233, N222);
xor XOR2 (N234, N225, N38);
not NOT1 (N235, N230);
nand NAND4 (N236, N235, N185, N146, N118);
or OR4 (N237, N232, N63, N202, N47);
or OR2 (N238, N219, N44);
nor NOR4 (N239, N210, N41, N72, N43);
not NOT1 (N240, N233);
not NOT1 (N241, N236);
or OR4 (N242, N224, N33, N65, N43);
and AND2 (N243, N223, N63);
nor NOR2 (N244, N243, N80);
or OR4 (N245, N237, N185, N195, N128);
nand NAND2 (N246, N242, N176);
nor NOR2 (N247, N231, N123);
or OR2 (N248, N245, N14);
xor XOR2 (N249, N239, N233);
nand NAND2 (N250, N227, N53);
buf BUF1 (N251, N246);
nand NAND3 (N252, N249, N59, N208);
not NOT1 (N253, N238);
nor NOR2 (N254, N250, N253);
buf BUF1 (N255, N42);
not NOT1 (N256, N251);
and AND3 (N257, N248, N82, N164);
xor XOR2 (N258, N247, N240);
not NOT1 (N259, N190);
not NOT1 (N260, N259);
nor NOR3 (N261, N256, N84, N185);
and AND2 (N262, N258, N87);
buf BUF1 (N263, N262);
nand NAND3 (N264, N234, N169, N90);
nor NOR4 (N265, N261, N20, N85, N41);
xor XOR2 (N266, N241, N60);
or OR4 (N267, N263, N186, N171, N223);
xor XOR2 (N268, N265, N10);
not NOT1 (N269, N260);
xor XOR2 (N270, N268, N180);
and AND4 (N271, N252, N199, N125, N56);
and AND3 (N272, N270, N216, N8);
xor XOR2 (N273, N255, N96);
buf BUF1 (N274, N271);
buf BUF1 (N275, N269);
nor NOR3 (N276, N254, N67, N210);
not NOT1 (N277, N266);
or OR2 (N278, N267, N123);
nand NAND2 (N279, N264, N208);
and AND2 (N280, N279, N6);
not NOT1 (N281, N278);
and AND4 (N282, N244, N84, N64, N165);
buf BUF1 (N283, N257);
not NOT1 (N284, N281);
nand NAND2 (N285, N277, N4);
and AND4 (N286, N284, N271, N94, N20);
nor NOR2 (N287, N274, N73);
or OR2 (N288, N283, N266);
nand NAND3 (N289, N280, N31, N69);
buf BUF1 (N290, N288);
and AND3 (N291, N286, N177, N175);
and AND4 (N292, N287, N183, N266, N48);
not NOT1 (N293, N282);
nor NOR2 (N294, N272, N186);
not NOT1 (N295, N290);
nor NOR2 (N296, N293, N83);
or OR2 (N297, N296, N206);
nor NOR2 (N298, N292, N102);
xor XOR2 (N299, N285, N261);
or OR3 (N300, N294, N215, N180);
buf BUF1 (N301, N289);
or OR2 (N302, N273, N103);
buf BUF1 (N303, N302);
or OR3 (N304, N299, N215, N45);
not NOT1 (N305, N301);
buf BUF1 (N306, N305);
nor NOR4 (N307, N297, N211, N226, N231);
not NOT1 (N308, N298);
and AND4 (N309, N307, N155, N225, N190);
nand NAND4 (N310, N276, N57, N131, N186);
nand NAND4 (N311, N308, N143, N90, N37);
nor NOR3 (N312, N291, N129, N223);
nor NOR2 (N313, N300, N239);
xor XOR2 (N314, N275, N265);
not NOT1 (N315, N306);
buf BUF1 (N316, N310);
and AND4 (N317, N309, N123, N126, N56);
not NOT1 (N318, N311);
and AND3 (N319, N314, N128, N53);
nor NOR3 (N320, N317, N199, N220);
nor NOR4 (N321, N318, N302, N263, N130);
buf BUF1 (N322, N315);
and AND4 (N323, N303, N217, N80, N194);
not NOT1 (N324, N319);
buf BUF1 (N325, N321);
not NOT1 (N326, N316);
nand NAND2 (N327, N326, N78);
and AND3 (N328, N323, N220, N62);
and AND2 (N329, N324, N53);
not NOT1 (N330, N304);
or OR3 (N331, N329, N242, N161);
nand NAND4 (N332, N328, N30, N87, N305);
not NOT1 (N333, N312);
buf BUF1 (N334, N332);
nand NAND2 (N335, N325, N186);
not NOT1 (N336, N330);
nand NAND4 (N337, N327, N306, N14, N177);
nor NOR2 (N338, N333, N152);
not NOT1 (N339, N331);
and AND2 (N340, N336, N204);
or OR4 (N341, N338, N276, N307, N291);
xor XOR2 (N342, N341, N38);
xor XOR2 (N343, N320, N190);
or OR3 (N344, N295, N152, N291);
nor NOR2 (N345, N342, N203);
buf BUF1 (N346, N340);
xor XOR2 (N347, N334, N234);
or OR2 (N348, N313, N214);
nand NAND4 (N349, N339, N115, N98, N138);
not NOT1 (N350, N349);
and AND4 (N351, N345, N202, N1, N264);
xor XOR2 (N352, N347, N93);
nor NOR3 (N353, N350, N33, N3);
and AND4 (N354, N335, N110, N252, N26);
buf BUF1 (N355, N343);
nor NOR4 (N356, N344, N210, N147, N330);
xor XOR2 (N357, N346, N192);
or OR4 (N358, N322, N61, N71, N212);
nand NAND3 (N359, N354, N139, N105);
buf BUF1 (N360, N356);
buf BUF1 (N361, N353);
nor NOR4 (N362, N358, N259, N4, N358);
or OR3 (N363, N360, N178, N349);
nand NAND3 (N364, N351, N68, N293);
xor XOR2 (N365, N355, N159);
xor XOR2 (N366, N357, N46);
not NOT1 (N367, N365);
buf BUF1 (N368, N337);
not NOT1 (N369, N367);
buf BUF1 (N370, N364);
nor NOR3 (N371, N348, N198, N7);
buf BUF1 (N372, N371);
nor NOR4 (N373, N372, N336, N241, N315);
or OR2 (N374, N368, N267);
not NOT1 (N375, N370);
xor XOR2 (N376, N366, N84);
and AND4 (N377, N363, N97, N265, N141);
xor XOR2 (N378, N376, N225);
not NOT1 (N379, N377);
xor XOR2 (N380, N352, N341);
not NOT1 (N381, N378);
and AND2 (N382, N361, N306);
not NOT1 (N383, N369);
not NOT1 (N384, N362);
and AND2 (N385, N379, N332);
nor NOR3 (N386, N384, N363, N104);
buf BUF1 (N387, N386);
nand NAND3 (N388, N373, N227, N137);
or OR4 (N389, N359, N190, N294, N314);
and AND2 (N390, N375, N369);
nor NOR2 (N391, N390, N294);
nand NAND4 (N392, N374, N155, N205, N5);
and AND2 (N393, N391, N86);
nand NAND4 (N394, N388, N305, N1, N380);
nor NOR3 (N395, N118, N384, N137);
nand NAND3 (N396, N383, N80, N28);
buf BUF1 (N397, N385);
buf BUF1 (N398, N395);
or OR4 (N399, N396, N12, N70, N304);
and AND4 (N400, N387, N106, N60, N310);
xor XOR2 (N401, N392, N312);
nor NOR3 (N402, N382, N275, N364);
nand NAND2 (N403, N398, N140);
nor NOR2 (N404, N402, N55);
nor NOR3 (N405, N399, N324, N222);
nand NAND4 (N406, N403, N197, N155, N93);
nor NOR2 (N407, N394, N343);
xor XOR2 (N408, N393, N56);
nor NOR3 (N409, N406, N132, N106);
not NOT1 (N410, N405);
nand NAND4 (N411, N409, N347, N93, N50);
not NOT1 (N412, N397);
xor XOR2 (N413, N410, N6);
not NOT1 (N414, N411);
buf BUF1 (N415, N400);
and AND3 (N416, N407, N132, N223);
buf BUF1 (N417, N381);
or OR4 (N418, N401, N92, N103, N261);
or OR2 (N419, N417, N312);
not NOT1 (N420, N418);
xor XOR2 (N421, N416, N172);
nor NOR3 (N422, N414, N147, N25);
buf BUF1 (N423, N419);
nor NOR3 (N424, N404, N213, N121);
buf BUF1 (N425, N412);
not NOT1 (N426, N424);
buf BUF1 (N427, N425);
xor XOR2 (N428, N421, N138);
nor NOR3 (N429, N423, N13, N155);
xor XOR2 (N430, N420, N79);
and AND3 (N431, N408, N318, N238);
or OR3 (N432, N426, N325, N8);
buf BUF1 (N433, N389);
or OR3 (N434, N430, N229, N151);
nand NAND2 (N435, N422, N391);
xor XOR2 (N436, N413, N125);
xor XOR2 (N437, N431, N414);
and AND2 (N438, N432, N358);
and AND3 (N439, N434, N22, N134);
buf BUF1 (N440, N439);
xor XOR2 (N441, N436, N17);
or OR4 (N442, N427, N288, N401, N21);
buf BUF1 (N443, N428);
xor XOR2 (N444, N443, N106);
nor NOR4 (N445, N433, N153, N386, N277);
nand NAND3 (N446, N442, N133, N306);
nor NOR4 (N447, N446, N419, N371, N92);
nor NOR2 (N448, N429, N76);
and AND2 (N449, N448, N47);
nand NAND2 (N450, N440, N303);
nand NAND2 (N451, N444, N20);
xor XOR2 (N452, N437, N150);
nand NAND4 (N453, N445, N143, N341, N193);
and AND4 (N454, N453, N3, N140, N449);
and AND2 (N455, N387, N36);
nand NAND2 (N456, N415, N234);
buf BUF1 (N457, N455);
nand NAND4 (N458, N438, N106, N344, N445);
not NOT1 (N459, N435);
xor XOR2 (N460, N451, N242);
buf BUF1 (N461, N447);
not NOT1 (N462, N456);
buf BUF1 (N463, N452);
nand NAND3 (N464, N459, N121, N299);
xor XOR2 (N465, N462, N90);
and AND2 (N466, N465, N43);
not NOT1 (N467, N458);
buf BUF1 (N468, N460);
xor XOR2 (N469, N466, N456);
xor XOR2 (N470, N454, N449);
xor XOR2 (N471, N467, N83);
nor NOR4 (N472, N441, N147, N102, N379);
or OR4 (N473, N470, N204, N359, N142);
and AND4 (N474, N457, N119, N439, N178);
buf BUF1 (N475, N464);
and AND2 (N476, N469, N450);
not NOT1 (N477, N211);
nor NOR3 (N478, N468, N277, N360);
xor XOR2 (N479, N475, N102);
nor NOR4 (N480, N463, N185, N253, N206);
and AND2 (N481, N477, N188);
buf BUF1 (N482, N472);
nand NAND2 (N483, N480, N251);
not NOT1 (N484, N482);
not NOT1 (N485, N483);
or OR4 (N486, N481, N481, N318, N80);
and AND3 (N487, N473, N326, N229);
xor XOR2 (N488, N487, N487);
or OR3 (N489, N476, N244, N329);
xor XOR2 (N490, N478, N469);
nor NOR2 (N491, N485, N242);
buf BUF1 (N492, N490);
or OR4 (N493, N479, N263, N403, N241);
xor XOR2 (N494, N491, N226);
nor NOR4 (N495, N492, N234, N89, N332);
and AND4 (N496, N489, N209, N479, N164);
buf BUF1 (N497, N471);
nand NAND2 (N498, N474, N178);
xor XOR2 (N499, N484, N278);
nor NOR4 (N500, N461, N353, N26, N55);
buf BUF1 (N501, N497);
and AND4 (N502, N499, N306, N62, N330);
and AND4 (N503, N500, N315, N242, N289);
nor NOR2 (N504, N496, N310);
buf BUF1 (N505, N495);
or OR2 (N506, N503, N71);
and AND4 (N507, N502, N240, N119, N12);
buf BUF1 (N508, N493);
nor NOR3 (N509, N501, N280, N299);
buf BUF1 (N510, N506);
buf BUF1 (N511, N505);
or OR3 (N512, N509, N421, N171);
or OR4 (N513, N498, N76, N345, N76);
nor NOR4 (N514, N504, N139, N247, N160);
nand NAND2 (N515, N511, N441);
not NOT1 (N516, N514);
not NOT1 (N517, N507);
nor NOR4 (N518, N510, N202, N292, N509);
or OR2 (N519, N494, N39);
not NOT1 (N520, N486);
nand NAND2 (N521, N518, N251);
or OR3 (N522, N517, N93, N376);
xor XOR2 (N523, N488, N215);
or OR4 (N524, N508, N140, N72, N199);
nor NOR2 (N525, N513, N203);
nor NOR3 (N526, N522, N331, N520);
not NOT1 (N527, N318);
xor XOR2 (N528, N527, N350);
buf BUF1 (N529, N519);
buf BUF1 (N530, N529);
xor XOR2 (N531, N523, N422);
and AND2 (N532, N526, N115);
not NOT1 (N533, N532);
not NOT1 (N534, N524);
buf BUF1 (N535, N534);
not NOT1 (N536, N533);
nand NAND3 (N537, N536, N446, N263);
xor XOR2 (N538, N537, N10);
xor XOR2 (N539, N528, N17);
and AND4 (N540, N512, N202, N373, N131);
and AND2 (N541, N539, N126);
and AND4 (N542, N538, N171, N224, N212);
xor XOR2 (N543, N515, N427);
and AND2 (N544, N543, N161);
or OR4 (N545, N540, N202, N241, N311);
or OR3 (N546, N541, N422, N296);
nor NOR4 (N547, N535, N83, N196, N316);
buf BUF1 (N548, N521);
xor XOR2 (N549, N548, N13);
xor XOR2 (N550, N530, N179);
nor NOR4 (N551, N542, N332, N237, N550);
and AND4 (N552, N95, N112, N220, N210);
nor NOR2 (N553, N545, N122);
nand NAND4 (N554, N549, N419, N172, N501);
nand NAND2 (N555, N531, N502);
xor XOR2 (N556, N547, N269);
not NOT1 (N557, N555);
not NOT1 (N558, N516);
or OR3 (N559, N553, N284, N187);
and AND4 (N560, N554, N362, N54, N347);
nand NAND4 (N561, N552, N21, N65, N40);
buf BUF1 (N562, N556);
buf BUF1 (N563, N551);
or OR3 (N564, N557, N257, N75);
buf BUF1 (N565, N564);
xor XOR2 (N566, N563, N186);
or OR4 (N567, N566, N491, N7, N393);
nand NAND3 (N568, N546, N94, N257);
nor NOR4 (N569, N561, N156, N361, N266);
nor NOR3 (N570, N558, N304, N549);
or OR3 (N571, N560, N240, N276);
or OR4 (N572, N562, N141, N256, N481);
and AND2 (N573, N571, N507);
buf BUF1 (N574, N570);
nand NAND4 (N575, N559, N570, N503, N218);
and AND3 (N576, N573, N134, N274);
nor NOR2 (N577, N576, N451);
buf BUF1 (N578, N567);
and AND4 (N579, N578, N56, N329, N445);
not NOT1 (N580, N569);
xor XOR2 (N581, N575, N196);
nor NOR3 (N582, N580, N471, N52);
nor NOR3 (N583, N582, N56, N265);
and AND3 (N584, N577, N137, N355);
nor NOR2 (N585, N584, N220);
buf BUF1 (N586, N581);
nor NOR3 (N587, N586, N313, N543);
not NOT1 (N588, N574);
and AND3 (N589, N588, N231, N557);
and AND2 (N590, N565, N22);
nand NAND4 (N591, N585, N442, N350, N380);
nor NOR2 (N592, N583, N576);
not NOT1 (N593, N587);
buf BUF1 (N594, N525);
not NOT1 (N595, N594);
and AND3 (N596, N568, N311, N233);
xor XOR2 (N597, N592, N176);
nand NAND3 (N598, N589, N137, N266);
nor NOR3 (N599, N595, N36, N41);
nor NOR4 (N600, N598, N13, N173, N63);
not NOT1 (N601, N597);
xor XOR2 (N602, N600, N181);
or OR3 (N603, N602, N596, N567);
and AND2 (N604, N37, N171);
nand NAND3 (N605, N590, N52, N443);
xor XOR2 (N606, N544, N577);
xor XOR2 (N607, N606, N142);
buf BUF1 (N608, N603);
and AND4 (N609, N572, N260, N209, N591);
nand NAND2 (N610, N568, N93);
not NOT1 (N611, N609);
not NOT1 (N612, N608);
or OR3 (N613, N593, N469, N324);
not NOT1 (N614, N579);
nor NOR3 (N615, N605, N575, N301);
nand NAND2 (N616, N604, N137);
nand NAND4 (N617, N601, N52, N92, N121);
nand NAND4 (N618, N611, N197, N143, N247);
nor NOR4 (N619, N607, N197, N20, N507);
nor NOR2 (N620, N615, N380);
nor NOR4 (N621, N620, N328, N416, N224);
nand NAND4 (N622, N614, N357, N474, N528);
not NOT1 (N623, N617);
xor XOR2 (N624, N616, N183);
not NOT1 (N625, N624);
nand NAND4 (N626, N610, N10, N312, N519);
buf BUF1 (N627, N612);
not NOT1 (N628, N599);
nand NAND2 (N629, N622, N235);
nand NAND2 (N630, N625, N296);
or OR2 (N631, N613, N68);
nor NOR3 (N632, N626, N607, N328);
nor NOR4 (N633, N629, N119, N235, N406);
and AND4 (N634, N631, N520, N212, N111);
not NOT1 (N635, N633);
xor XOR2 (N636, N632, N490);
or OR4 (N637, N636, N129, N356, N265);
buf BUF1 (N638, N635);
or OR3 (N639, N637, N88, N359);
or OR3 (N640, N621, N453, N489);
xor XOR2 (N641, N627, N43);
xor XOR2 (N642, N638, N384);
nand NAND2 (N643, N623, N12);
xor XOR2 (N644, N619, N307);
xor XOR2 (N645, N618, N1);
xor XOR2 (N646, N643, N27);
not NOT1 (N647, N628);
nand NAND2 (N648, N644, N24);
nor NOR3 (N649, N642, N581, N247);
nor NOR4 (N650, N649, N154, N124, N366);
buf BUF1 (N651, N630);
nor NOR4 (N652, N651, N330, N197, N171);
nor NOR3 (N653, N652, N151, N242);
nand NAND3 (N654, N641, N309, N356);
xor XOR2 (N655, N634, N593);
and AND3 (N656, N653, N366, N327);
buf BUF1 (N657, N650);
not NOT1 (N658, N647);
and AND4 (N659, N655, N129, N504, N634);
buf BUF1 (N660, N654);
or OR4 (N661, N657, N603, N531, N160);
not NOT1 (N662, N656);
and AND2 (N663, N659, N373);
and AND3 (N664, N639, N585, N345);
nand NAND2 (N665, N640, N213);
nor NOR4 (N666, N648, N638, N408, N422);
nor NOR2 (N667, N666, N175);
nor NOR2 (N668, N661, N168);
nand NAND4 (N669, N668, N167, N171, N380);
nor NOR3 (N670, N665, N123, N304);
buf BUF1 (N671, N669);
buf BUF1 (N672, N664);
buf BUF1 (N673, N658);
xor XOR2 (N674, N670, N347);
not NOT1 (N675, N667);
and AND3 (N676, N674, N604, N466);
buf BUF1 (N677, N673);
nand NAND3 (N678, N672, N593, N325);
and AND2 (N679, N663, N656);
nor NOR4 (N680, N660, N158, N642, N258);
and AND2 (N681, N662, N186);
and AND4 (N682, N675, N18, N124, N511);
nor NOR3 (N683, N678, N54, N398);
or OR4 (N684, N645, N151, N483, N298);
nand NAND3 (N685, N646, N275, N65);
and AND2 (N686, N680, N312);
nand NAND2 (N687, N685, N584);
and AND2 (N688, N683, N534);
or OR4 (N689, N688, N451, N212, N399);
and AND3 (N690, N679, N413, N115);
nor NOR2 (N691, N690, N546);
nand NAND4 (N692, N684, N264, N54, N563);
xor XOR2 (N693, N692, N453);
and AND3 (N694, N691, N290, N201);
or OR2 (N695, N677, N621);
nor NOR2 (N696, N671, N615);
or OR3 (N697, N686, N419, N673);
nor NOR3 (N698, N681, N549, N690);
or OR3 (N699, N697, N507, N685);
buf BUF1 (N700, N693);
or OR2 (N701, N700, N338);
not NOT1 (N702, N676);
or OR4 (N703, N699, N3, N514, N183);
or OR3 (N704, N698, N77, N66);
not NOT1 (N705, N687);
and AND4 (N706, N703, N677, N418, N488);
nand NAND3 (N707, N696, N213, N216);
or OR3 (N708, N702, N308, N414);
not NOT1 (N709, N707);
or OR3 (N710, N701, N257, N145);
nor NOR3 (N711, N706, N333, N79);
nand NAND4 (N712, N709, N403, N133, N468);
nand NAND2 (N713, N695, N30);
and AND3 (N714, N712, N582, N153);
and AND3 (N715, N689, N119, N225);
or OR3 (N716, N713, N19, N600);
nand NAND4 (N717, N708, N348, N357, N206);
or OR3 (N718, N682, N562, N675);
nor NOR4 (N719, N705, N61, N195, N270);
or OR3 (N720, N718, N144, N166);
nand NAND4 (N721, N694, N657, N568, N398);
nand NAND3 (N722, N721, N330, N381);
buf BUF1 (N723, N720);
nand NAND2 (N724, N710, N219);
nand NAND3 (N725, N719, N172, N179);
and AND2 (N726, N716, N610);
nor NOR3 (N727, N714, N171, N220);
and AND3 (N728, N723, N349, N30);
and AND3 (N729, N725, N138, N343);
and AND2 (N730, N729, N710);
buf BUF1 (N731, N722);
nand NAND4 (N732, N724, N163, N407, N68);
not NOT1 (N733, N728);
not NOT1 (N734, N711);
or OR4 (N735, N731, N123, N143, N547);
buf BUF1 (N736, N727);
nand NAND3 (N737, N735, N569, N383);
buf BUF1 (N738, N733);
buf BUF1 (N739, N715);
nor NOR3 (N740, N737, N335, N68);
xor XOR2 (N741, N717, N609);
xor XOR2 (N742, N730, N445);
nand NAND3 (N743, N734, N596, N216);
buf BUF1 (N744, N742);
nand NAND4 (N745, N704, N523, N310, N630);
nand NAND3 (N746, N732, N251, N658);
or OR2 (N747, N746, N244);
buf BUF1 (N748, N745);
xor XOR2 (N749, N726, N159);
or OR3 (N750, N736, N79, N401);
buf BUF1 (N751, N741);
nand NAND4 (N752, N743, N154, N209, N579);
or OR4 (N753, N751, N377, N565, N622);
nand NAND2 (N754, N750, N213);
not NOT1 (N755, N748);
nor NOR4 (N756, N754, N174, N628, N167);
or OR2 (N757, N756, N177);
buf BUF1 (N758, N747);
or OR3 (N759, N738, N500, N113);
nand NAND3 (N760, N752, N407, N240);
or OR4 (N761, N753, N517, N736, N106);
buf BUF1 (N762, N757);
or OR2 (N763, N744, N440);
or OR2 (N764, N759, N129);
and AND3 (N765, N764, N621, N88);
nand NAND3 (N766, N755, N545, N161);
buf BUF1 (N767, N766);
buf BUF1 (N768, N765);
buf BUF1 (N769, N760);
and AND3 (N770, N763, N619, N661);
xor XOR2 (N771, N761, N304);
not NOT1 (N772, N770);
nand NAND2 (N773, N758, N21);
nand NAND4 (N774, N769, N298, N272, N42);
nor NOR4 (N775, N740, N604, N550, N428);
and AND2 (N776, N772, N736);
and AND4 (N777, N767, N87, N99, N125);
xor XOR2 (N778, N739, N536);
nor NOR2 (N779, N778, N452);
buf BUF1 (N780, N768);
not NOT1 (N781, N771);
not NOT1 (N782, N781);
nand NAND3 (N783, N775, N16, N170);
xor XOR2 (N784, N773, N637);
and AND2 (N785, N776, N134);
and AND3 (N786, N782, N359, N235);
buf BUF1 (N787, N762);
and AND4 (N788, N749, N754, N233, N447);
xor XOR2 (N789, N786, N189);
and AND4 (N790, N784, N29, N314, N355);
nand NAND2 (N791, N774, N426);
or OR3 (N792, N789, N372, N739);
and AND2 (N793, N787, N493);
nor NOR3 (N794, N791, N269, N711);
nor NOR3 (N795, N788, N748, N561);
and AND2 (N796, N794, N592);
nand NAND2 (N797, N796, N107);
or OR4 (N798, N777, N614, N72, N209);
xor XOR2 (N799, N785, N309);
xor XOR2 (N800, N799, N252);
nor NOR2 (N801, N797, N9);
not NOT1 (N802, N798);
nand NAND3 (N803, N783, N89, N139);
not NOT1 (N804, N795);
nand NAND2 (N805, N801, N160);
xor XOR2 (N806, N792, N309);
nor NOR4 (N807, N806, N558, N196, N426);
buf BUF1 (N808, N807);
or OR4 (N809, N803, N11, N58, N303);
xor XOR2 (N810, N805, N149);
nor NOR4 (N811, N780, N738, N596, N491);
or OR3 (N812, N790, N781, N641);
or OR4 (N813, N809, N32, N113, N544);
or OR2 (N814, N779, N271);
nor NOR2 (N815, N802, N653);
nor NOR3 (N816, N814, N272, N56);
buf BUF1 (N817, N812);
xor XOR2 (N818, N810, N305);
not NOT1 (N819, N800);
not NOT1 (N820, N815);
not NOT1 (N821, N817);
or OR4 (N822, N793, N663, N651, N313);
nand NAND4 (N823, N804, N118, N258, N490);
nor NOR3 (N824, N808, N232, N42);
buf BUF1 (N825, N816);
nor NOR4 (N826, N811, N489, N760, N238);
not NOT1 (N827, N822);
xor XOR2 (N828, N823, N588);
xor XOR2 (N829, N818, N33);
nor NOR4 (N830, N828, N515, N179, N244);
or OR3 (N831, N825, N132, N164);
nor NOR2 (N832, N829, N704);
or OR3 (N833, N819, N415, N802);
nor NOR2 (N834, N831, N380);
not NOT1 (N835, N830);
nor NOR4 (N836, N826, N30, N403, N534);
nor NOR2 (N837, N833, N179);
and AND2 (N838, N836, N426);
and AND3 (N839, N820, N619, N726);
or OR4 (N840, N824, N145, N68, N125);
not NOT1 (N841, N840);
or OR2 (N842, N835, N744);
nand NAND4 (N843, N838, N93, N352, N770);
or OR4 (N844, N839, N664, N25, N711);
or OR3 (N845, N832, N572, N142);
nor NOR4 (N846, N841, N781, N664, N19);
not NOT1 (N847, N843);
buf BUF1 (N848, N845);
and AND3 (N849, N847, N724, N244);
and AND3 (N850, N837, N331, N47);
and AND2 (N851, N844, N831);
buf BUF1 (N852, N813);
not NOT1 (N853, N821);
nor NOR3 (N854, N850, N654, N123);
xor XOR2 (N855, N846, N251);
not NOT1 (N856, N851);
xor XOR2 (N857, N834, N300);
buf BUF1 (N858, N853);
xor XOR2 (N859, N856, N806);
nor NOR2 (N860, N858, N341);
not NOT1 (N861, N849);
buf BUF1 (N862, N827);
nor NOR2 (N863, N862, N697);
xor XOR2 (N864, N842, N475);
nand NAND4 (N865, N863, N56, N533, N147);
nor NOR2 (N866, N857, N284);
xor XOR2 (N867, N865, N469);
xor XOR2 (N868, N867, N167);
nand NAND4 (N869, N855, N805, N201, N180);
or OR3 (N870, N864, N701, N331);
buf BUF1 (N871, N868);
nand NAND3 (N872, N848, N778, N627);
xor XOR2 (N873, N861, N76);
and AND2 (N874, N854, N769);
buf BUF1 (N875, N866);
or OR4 (N876, N852, N49, N226, N852);
nand NAND4 (N877, N876, N705, N337, N695);
or OR2 (N878, N870, N15);
nor NOR3 (N879, N859, N835, N372);
nor NOR3 (N880, N878, N692, N487);
xor XOR2 (N881, N874, N727);
not NOT1 (N882, N871);
buf BUF1 (N883, N860);
or OR3 (N884, N869, N575, N340);
or OR3 (N885, N882, N844, N374);
nor NOR4 (N886, N877, N189, N6, N647);
buf BUF1 (N887, N875);
and AND3 (N888, N879, N310, N495);
xor XOR2 (N889, N888, N64);
nor NOR3 (N890, N885, N349, N768);
not NOT1 (N891, N889);
nand NAND2 (N892, N873, N42);
buf BUF1 (N893, N880);
buf BUF1 (N894, N892);
buf BUF1 (N895, N872);
not NOT1 (N896, N883);
buf BUF1 (N897, N886);
nor NOR4 (N898, N895, N872, N658, N851);
and AND4 (N899, N894, N312, N488, N144);
buf BUF1 (N900, N887);
nand NAND3 (N901, N884, N27, N852);
or OR4 (N902, N891, N554, N172, N790);
xor XOR2 (N903, N896, N498);
or OR4 (N904, N900, N77, N708, N672);
buf BUF1 (N905, N902);
nand NAND3 (N906, N898, N14, N469);
nor NOR4 (N907, N890, N715, N663, N300);
xor XOR2 (N908, N906, N521);
nor NOR2 (N909, N903, N800);
not NOT1 (N910, N901);
endmodule