// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N16016,N16018,N16007,N15939,N16017,N16012,N16000,N16010,N16015,N16019;

nand NAND4 (N20, N19, N1, N16, N8);
and AND4 (N21, N2, N20, N10, N18);
buf BUF1 (N22, N21);
nand NAND2 (N23, N1, N8);
buf BUF1 (N24, N5);
nand NAND2 (N25, N7, N22);
buf BUF1 (N26, N19);
nor NOR3 (N27, N15, N20, N1);
nand NAND2 (N28, N17, N13);
nand NAND4 (N29, N11, N22, N6, N22);
and AND4 (N30, N15, N28, N17, N21);
nand NAND4 (N31, N22, N9, N26, N7);
xor XOR2 (N32, N1, N28);
xor XOR2 (N33, N6, N19);
xor XOR2 (N34, N21, N5);
nor NOR3 (N35, N27, N33, N30);
xor XOR2 (N36, N21, N17);
xor XOR2 (N37, N21, N15);
or OR3 (N38, N35, N11, N22);
xor XOR2 (N39, N37, N27);
xor XOR2 (N40, N31, N12);
nor NOR2 (N41, N34, N10);
buf BUF1 (N42, N24);
and AND4 (N43, N32, N8, N9, N35);
nand NAND4 (N44, N41, N19, N43, N11);
or OR2 (N45, N15, N30);
not NOT1 (N46, N25);
and AND3 (N47, N45, N45, N31);
and AND2 (N48, N40, N34);
xor XOR2 (N49, N36, N19);
nand NAND4 (N50, N23, N7, N48, N22);
not NOT1 (N51, N34);
buf BUF1 (N52, N44);
nand NAND3 (N53, N29, N17, N25);
not NOT1 (N54, N38);
and AND3 (N55, N42, N38, N50);
and AND4 (N56, N53, N52, N3, N43);
buf BUF1 (N57, N44);
buf BUF1 (N58, N27);
xor XOR2 (N59, N51, N17);
buf BUF1 (N60, N57);
xor XOR2 (N61, N58, N8);
or OR4 (N62, N39, N32, N61, N52);
buf BUF1 (N63, N57);
and AND3 (N64, N59, N47, N49);
and AND2 (N65, N47, N34);
or OR3 (N66, N61, N16, N25);
and AND2 (N67, N46, N5);
or OR3 (N68, N54, N12, N29);
and AND4 (N69, N56, N36, N37, N63);
nand NAND2 (N70, N8, N50);
buf BUF1 (N71, N70);
and AND4 (N72, N62, N37, N63, N34);
nand NAND4 (N73, N72, N49, N41, N60);
nand NAND4 (N74, N3, N2, N29, N49);
or OR3 (N75, N68, N68, N41);
and AND3 (N76, N69, N20, N6);
buf BUF1 (N77, N55);
and AND2 (N78, N64, N67);
and AND2 (N79, N58, N41);
nor NOR4 (N80, N71, N14, N37, N19);
and AND3 (N81, N78, N65, N40);
nand NAND2 (N82, N53, N27);
buf BUF1 (N83, N80);
and AND2 (N84, N74, N47);
nand NAND2 (N85, N82, N76);
nor NOR2 (N86, N64, N78);
not NOT1 (N87, N84);
nor NOR2 (N88, N86, N4);
and AND3 (N89, N66, N71, N52);
nor NOR4 (N90, N87, N8, N77, N76);
nor NOR3 (N91, N88, N21, N7);
nand NAND4 (N92, N14, N90, N85, N56);
or OR4 (N93, N73, N3, N92, N77);
or OR3 (N94, N44, N88, N14);
nor NOR3 (N95, N51, N83, N20);
nor NOR3 (N96, N21, N10, N37);
or OR4 (N97, N7, N42, N76, N20);
buf BUF1 (N98, N75);
xor XOR2 (N99, N94, N68);
nor NOR2 (N100, N96, N29);
nor NOR3 (N101, N91, N97, N81);
and AND2 (N102, N98, N15);
nor NOR3 (N103, N81, N21, N82);
not NOT1 (N104, N63);
nand NAND4 (N105, N95, N56, N49, N10);
buf BUF1 (N106, N89);
nor NOR3 (N107, N93, N2, N39);
nand NAND3 (N108, N99, N98, N98);
or OR4 (N109, N103, N101, N33, N23);
nor NOR4 (N110, N51, N31, N11, N58);
nand NAND2 (N111, N79, N62);
nor NOR3 (N112, N102, N106, N50);
buf BUF1 (N113, N65);
buf BUF1 (N114, N108);
or OR3 (N115, N114, N4, N59);
xor XOR2 (N116, N105, N86);
nand NAND4 (N117, N109, N40, N46, N98);
buf BUF1 (N118, N115);
or OR4 (N119, N118, N102, N74, N8);
nor NOR4 (N120, N107, N105, N15, N105);
nor NOR4 (N121, N112, N87, N71, N120);
and AND3 (N122, N39, N22, N113);
or OR3 (N123, N24, N95, N14);
nor NOR3 (N124, N104, N84, N16);
xor XOR2 (N125, N117, N79);
xor XOR2 (N126, N124, N100);
not NOT1 (N127, N22);
not NOT1 (N128, N119);
xor XOR2 (N129, N126, N49);
and AND4 (N130, N129, N71, N89, N50);
not NOT1 (N131, N123);
not NOT1 (N132, N111);
xor XOR2 (N133, N121, N57);
buf BUF1 (N134, N130);
nand NAND4 (N135, N116, N80, N67, N91);
and AND4 (N136, N110, N73, N79, N57);
not NOT1 (N137, N135);
xor XOR2 (N138, N128, N116);
and AND2 (N139, N138, N99);
and AND3 (N140, N136, N133, N69);
or OR3 (N141, N46, N81, N114);
xor XOR2 (N142, N140, N130);
and AND3 (N143, N141, N36, N23);
xor XOR2 (N144, N134, N90);
or OR3 (N145, N127, N30, N136);
xor XOR2 (N146, N143, N62);
nor NOR3 (N147, N137, N60, N43);
or OR2 (N148, N131, N111);
and AND3 (N149, N146, N38, N68);
nor NOR2 (N150, N148, N78);
xor XOR2 (N151, N125, N100);
nor NOR3 (N152, N150, N137, N70);
and AND2 (N153, N122, N12);
or OR3 (N154, N147, N16, N97);
nor NOR4 (N155, N151, N7, N87, N31);
or OR3 (N156, N153, N140, N140);
buf BUF1 (N157, N132);
buf BUF1 (N158, N155);
and AND4 (N159, N157, N90, N144, N55);
and AND2 (N160, N91, N158);
and AND3 (N161, N127, N150, N19);
buf BUF1 (N162, N161);
or OR2 (N163, N142, N120);
buf BUF1 (N164, N145);
buf BUF1 (N165, N163);
not NOT1 (N166, N139);
or OR4 (N167, N165, N105, N96, N79);
buf BUF1 (N168, N162);
and AND2 (N169, N149, N47);
not NOT1 (N170, N152);
not NOT1 (N171, N169);
or OR3 (N172, N168, N70, N85);
xor XOR2 (N173, N166, N76);
or OR3 (N174, N160, N127, N73);
xor XOR2 (N175, N156, N136);
nor NOR4 (N176, N164, N81, N32, N43);
xor XOR2 (N177, N174, N151);
xor XOR2 (N178, N159, N102);
or OR3 (N179, N177, N100, N128);
xor XOR2 (N180, N170, N138);
xor XOR2 (N181, N180, N124);
buf BUF1 (N182, N154);
xor XOR2 (N183, N182, N165);
nand NAND2 (N184, N179, N104);
and AND2 (N185, N181, N73);
xor XOR2 (N186, N175, N146);
buf BUF1 (N187, N186);
nor NOR4 (N188, N178, N115, N179, N184);
not NOT1 (N189, N133);
buf BUF1 (N190, N187);
or OR4 (N191, N185, N25, N102, N111);
nor NOR3 (N192, N191, N16, N185);
xor XOR2 (N193, N176, N65);
nand NAND2 (N194, N189, N36);
buf BUF1 (N195, N173);
nor NOR2 (N196, N192, N2);
and AND2 (N197, N171, N126);
nor NOR4 (N198, N167, N163, N154, N64);
or OR4 (N199, N194, N122, N176, N115);
and AND2 (N200, N197, N146);
xor XOR2 (N201, N188, N83);
and AND4 (N202, N200, N65, N35, N152);
and AND2 (N203, N190, N41);
or OR2 (N204, N199, N156);
not NOT1 (N205, N203);
nand NAND2 (N206, N204, N64);
not NOT1 (N207, N201);
not NOT1 (N208, N195);
and AND2 (N209, N183, N124);
nor NOR2 (N210, N207, N44);
or OR4 (N211, N172, N81, N76, N48);
and AND2 (N212, N206, N116);
nand NAND4 (N213, N209, N8, N64, N148);
and AND2 (N214, N205, N152);
nor NOR3 (N215, N212, N118, N208);
or OR3 (N216, N42, N128, N182);
buf BUF1 (N217, N216);
nand NAND2 (N218, N210, N11);
xor XOR2 (N219, N213, N12);
nand NAND3 (N220, N202, N167, N212);
nor NOR4 (N221, N211, N147, N209, N204);
nand NAND3 (N222, N220, N205, N133);
buf BUF1 (N223, N217);
buf BUF1 (N224, N215);
not NOT1 (N225, N193);
xor XOR2 (N226, N196, N147);
xor XOR2 (N227, N226, N70);
nor NOR3 (N228, N224, N40, N100);
not NOT1 (N229, N222);
or OR3 (N230, N227, N18, N175);
xor XOR2 (N231, N219, N173);
not NOT1 (N232, N221);
and AND4 (N233, N218, N177, N51, N43);
buf BUF1 (N234, N228);
xor XOR2 (N235, N231, N219);
and AND3 (N236, N230, N216, N73);
xor XOR2 (N237, N225, N110);
buf BUF1 (N238, N232);
or OR2 (N239, N233, N128);
and AND4 (N240, N223, N138, N226, N227);
xor XOR2 (N241, N234, N96);
not NOT1 (N242, N229);
nand NAND2 (N243, N241, N97);
or OR3 (N244, N239, N65, N149);
buf BUF1 (N245, N235);
nor NOR2 (N246, N198, N100);
nor NOR2 (N247, N245, N150);
and AND2 (N248, N246, N52);
buf BUF1 (N249, N237);
xor XOR2 (N250, N248, N182);
not NOT1 (N251, N249);
xor XOR2 (N252, N250, N56);
nand NAND3 (N253, N243, N220, N203);
not NOT1 (N254, N238);
nand NAND4 (N255, N214, N1, N178, N74);
not NOT1 (N256, N244);
xor XOR2 (N257, N253, N177);
nor NOR2 (N258, N252, N126);
not NOT1 (N259, N240);
or OR3 (N260, N257, N96, N19);
nor NOR4 (N261, N259, N126, N217, N211);
buf BUF1 (N262, N260);
nand NAND3 (N263, N256, N182, N153);
and AND4 (N264, N242, N227, N48, N153);
not NOT1 (N265, N254);
and AND3 (N266, N255, N240, N55);
buf BUF1 (N267, N247);
nor NOR4 (N268, N266, N215, N232, N262);
nor NOR4 (N269, N228, N160, N90, N33);
xor XOR2 (N270, N258, N166);
not NOT1 (N271, N265);
or OR2 (N272, N269, N145);
nand NAND3 (N273, N264, N98, N119);
not NOT1 (N274, N273);
nand NAND4 (N275, N261, N234, N250, N78);
nand NAND2 (N276, N271, N69);
nand NAND3 (N277, N276, N115, N12);
not NOT1 (N278, N251);
nand NAND2 (N279, N268, N195);
xor XOR2 (N280, N270, N75);
xor XOR2 (N281, N275, N62);
or OR4 (N282, N236, N204, N4, N190);
not NOT1 (N283, N280);
xor XOR2 (N284, N283, N263);
buf BUF1 (N285, N263);
not NOT1 (N286, N281);
buf BUF1 (N287, N286);
buf BUF1 (N288, N284);
buf BUF1 (N289, N274);
nand NAND2 (N290, N272, N83);
xor XOR2 (N291, N279, N173);
nor NOR4 (N292, N287, N150, N70, N163);
xor XOR2 (N293, N292, N59);
and AND3 (N294, N277, N11, N154);
or OR2 (N295, N290, N224);
buf BUF1 (N296, N289);
not NOT1 (N297, N291);
xor XOR2 (N298, N293, N201);
nand NAND3 (N299, N297, N25, N262);
buf BUF1 (N300, N295);
and AND3 (N301, N296, N79, N100);
nor NOR3 (N302, N299, N291, N203);
xor XOR2 (N303, N300, N273);
buf BUF1 (N304, N298);
and AND2 (N305, N288, N304);
buf BUF1 (N306, N154);
or OR2 (N307, N303, N284);
nand NAND3 (N308, N306, N193, N208);
buf BUF1 (N309, N267);
or OR3 (N310, N309, N165, N86);
nand NAND4 (N311, N278, N102, N86, N290);
nand NAND3 (N312, N305, N131, N269);
nor NOR2 (N313, N302, N110);
or OR3 (N314, N307, N141, N145);
buf BUF1 (N315, N310);
and AND3 (N316, N285, N119, N297);
nor NOR2 (N317, N312, N65);
nand NAND2 (N318, N313, N64);
buf BUF1 (N319, N301);
xor XOR2 (N320, N314, N237);
and AND3 (N321, N315, N277, N59);
xor XOR2 (N322, N311, N272);
or OR4 (N323, N316, N187, N180, N209);
nand NAND3 (N324, N323, N228, N153);
buf BUF1 (N325, N320);
or OR3 (N326, N294, N227, N124);
and AND4 (N327, N317, N234, N198, N47);
and AND4 (N328, N308, N221, N164, N71);
and AND2 (N329, N318, N145);
nor NOR4 (N330, N282, N298, N232, N194);
and AND2 (N331, N321, N176);
xor XOR2 (N332, N329, N62);
buf BUF1 (N333, N325);
nand NAND3 (N334, N327, N24, N313);
nor NOR4 (N335, N333, N107, N198, N227);
or OR4 (N336, N319, N215, N2, N291);
and AND2 (N337, N322, N336);
nor NOR4 (N338, N219, N289, N326, N142);
xor XOR2 (N339, N150, N155);
xor XOR2 (N340, N338, N248);
or OR4 (N341, N331, N305, N328, N3);
or OR4 (N342, N25, N31, N322, N203);
nor NOR3 (N343, N337, N327, N66);
buf BUF1 (N344, N342);
or OR4 (N345, N344, N143, N261, N160);
and AND4 (N346, N339, N97, N175, N81);
nand NAND2 (N347, N335, N114);
nand NAND3 (N348, N324, N128, N14);
xor XOR2 (N349, N348, N19);
not NOT1 (N350, N347);
nor NOR4 (N351, N343, N234, N35, N182);
or OR2 (N352, N349, N334);
nand NAND2 (N353, N206, N114);
buf BUF1 (N354, N345);
nand NAND3 (N355, N341, N133, N214);
and AND2 (N356, N340, N304);
and AND3 (N357, N355, N153, N157);
nor NOR4 (N358, N353, N251, N21, N91);
and AND3 (N359, N351, N210, N155);
and AND4 (N360, N346, N206, N11, N319);
not NOT1 (N361, N332);
nor NOR2 (N362, N354, N156);
or OR3 (N363, N361, N14, N183);
or OR3 (N364, N356, N269, N258);
and AND2 (N365, N364, N45);
and AND3 (N366, N358, N328, N221);
and AND3 (N367, N363, N347, N49);
not NOT1 (N368, N350);
xor XOR2 (N369, N366, N309);
and AND2 (N370, N360, N224);
nor NOR2 (N371, N359, N321);
or OR3 (N372, N369, N161, N296);
xor XOR2 (N373, N371, N18);
or OR4 (N374, N352, N222, N115, N235);
or OR2 (N375, N368, N3);
buf BUF1 (N376, N365);
buf BUF1 (N377, N367);
nor NOR4 (N378, N330, N134, N18, N170);
buf BUF1 (N379, N375);
xor XOR2 (N380, N362, N102);
nor NOR2 (N381, N376, N149);
nor NOR2 (N382, N381, N161);
or OR2 (N383, N382, N186);
buf BUF1 (N384, N374);
xor XOR2 (N385, N380, N304);
xor XOR2 (N386, N379, N339);
nand NAND3 (N387, N377, N152, N256);
nand NAND4 (N388, N372, N82, N387, N280);
xor XOR2 (N389, N15, N187);
buf BUF1 (N390, N373);
or OR4 (N391, N370, N306, N266, N364);
or OR4 (N392, N383, N250, N277, N223);
xor XOR2 (N393, N378, N305);
nand NAND4 (N394, N388, N389, N349, N209);
nand NAND3 (N395, N63, N290, N107);
or OR4 (N396, N391, N45, N136, N314);
or OR3 (N397, N393, N396, N54);
nand NAND4 (N398, N200, N228, N65, N88);
or OR4 (N399, N394, N154, N11, N285);
and AND4 (N400, N385, N22, N306, N311);
xor XOR2 (N401, N390, N100);
or OR2 (N402, N395, N297);
xor XOR2 (N403, N384, N5);
xor XOR2 (N404, N403, N100);
xor XOR2 (N405, N357, N309);
or OR2 (N406, N386, N78);
xor XOR2 (N407, N402, N306);
nand NAND3 (N408, N405, N52, N45);
xor XOR2 (N409, N399, N277);
nor NOR3 (N410, N401, N6, N173);
xor XOR2 (N411, N410, N174);
or OR3 (N412, N406, N65, N90);
buf BUF1 (N413, N404);
nor NOR4 (N414, N412, N73, N240, N160);
nand NAND3 (N415, N407, N14, N75);
buf BUF1 (N416, N397);
buf BUF1 (N417, N398);
nor NOR3 (N418, N415, N246, N182);
not NOT1 (N419, N413);
buf BUF1 (N420, N408);
nand NAND4 (N421, N409, N205, N109, N406);
nor NOR3 (N422, N416, N232, N227);
nor NOR4 (N423, N411, N165, N350, N108);
and AND2 (N424, N417, N59);
nor NOR4 (N425, N420, N71, N63, N341);
nand NAND2 (N426, N419, N26);
xor XOR2 (N427, N400, N179);
or OR3 (N428, N424, N249, N365);
and AND3 (N429, N422, N58, N271);
xor XOR2 (N430, N414, N131);
and AND3 (N431, N423, N282, N70);
not NOT1 (N432, N431);
nand NAND4 (N433, N392, N37, N191, N289);
or OR3 (N434, N418, N1, N260);
nand NAND3 (N435, N432, N239, N106);
or OR3 (N436, N435, N14, N424);
or OR4 (N437, N427, N328, N10, N222);
nor NOR4 (N438, N433, N53, N405, N282);
buf BUF1 (N439, N428);
or OR4 (N440, N434, N244, N318, N319);
or OR3 (N441, N436, N178, N118);
and AND3 (N442, N429, N124, N389);
or OR2 (N443, N426, N98);
or OR4 (N444, N442, N424, N13, N433);
not NOT1 (N445, N440);
not NOT1 (N446, N439);
xor XOR2 (N447, N430, N444);
nor NOR2 (N448, N19, N361);
xor XOR2 (N449, N448, N73);
or OR4 (N450, N445, N188, N327, N52);
or OR3 (N451, N425, N384, N129);
xor XOR2 (N452, N443, N314);
and AND2 (N453, N450, N235);
not NOT1 (N454, N441);
not NOT1 (N455, N437);
or OR2 (N456, N421, N139);
or OR4 (N457, N446, N70, N211, N132);
and AND4 (N458, N449, N152, N332, N186);
nand NAND2 (N459, N451, N324);
nand NAND4 (N460, N438, N444, N168, N161);
xor XOR2 (N461, N447, N125);
buf BUF1 (N462, N460);
or OR4 (N463, N455, N235, N281, N191);
not NOT1 (N464, N461);
not NOT1 (N465, N464);
nand NAND3 (N466, N462, N378, N166);
buf BUF1 (N467, N452);
or OR3 (N468, N453, N29, N188);
not NOT1 (N469, N466);
and AND3 (N470, N463, N375, N228);
buf BUF1 (N471, N469);
xor XOR2 (N472, N470, N62);
nand NAND4 (N473, N468, N417, N252, N400);
xor XOR2 (N474, N456, N315);
buf BUF1 (N475, N471);
xor XOR2 (N476, N475, N308);
or OR2 (N477, N467, N349);
nor NOR3 (N478, N472, N333, N211);
not NOT1 (N479, N476);
nand NAND2 (N480, N465, N161);
or OR2 (N481, N458, N208);
xor XOR2 (N482, N480, N434);
nand NAND2 (N483, N478, N241);
not NOT1 (N484, N479);
and AND3 (N485, N457, N149, N421);
not NOT1 (N486, N482);
not NOT1 (N487, N459);
nand NAND3 (N488, N481, N410, N112);
nor NOR4 (N489, N473, N8, N65, N61);
or OR2 (N490, N484, N246);
and AND3 (N491, N486, N472, N451);
xor XOR2 (N492, N489, N138);
and AND4 (N493, N474, N441, N114, N220);
xor XOR2 (N494, N483, N285);
and AND4 (N495, N487, N275, N70, N101);
or OR2 (N496, N454, N404);
not NOT1 (N497, N496);
or OR3 (N498, N492, N489, N86);
nor NOR4 (N499, N490, N494, N262, N403);
and AND4 (N500, N376, N246, N266, N471);
nand NAND2 (N501, N497, N118);
or OR2 (N502, N500, N24);
buf BUF1 (N503, N488);
nor NOR3 (N504, N503, N446, N393);
nor NOR3 (N505, N504, N442, N304);
nor NOR3 (N506, N485, N335, N418);
or OR2 (N507, N501, N429);
nor NOR3 (N508, N498, N271, N16);
xor XOR2 (N509, N491, N396);
xor XOR2 (N510, N502, N173);
buf BUF1 (N511, N493);
or OR4 (N512, N509, N174, N347, N498);
buf BUF1 (N513, N505);
nand NAND2 (N514, N495, N184);
xor XOR2 (N515, N477, N405);
or OR4 (N516, N513, N363, N492, N183);
nand NAND4 (N517, N510, N384, N109, N439);
xor XOR2 (N518, N516, N477);
or OR2 (N519, N514, N514);
not NOT1 (N520, N507);
xor XOR2 (N521, N499, N434);
nand NAND3 (N522, N506, N2, N161);
or OR4 (N523, N520, N337, N305, N317);
xor XOR2 (N524, N515, N459);
nor NOR3 (N525, N521, N374, N515);
not NOT1 (N526, N511);
nor NOR3 (N527, N517, N262, N107);
buf BUF1 (N528, N526);
and AND3 (N529, N518, N76, N364);
buf BUF1 (N530, N522);
nand NAND4 (N531, N519, N133, N330, N46);
nand NAND4 (N532, N524, N360, N5, N468);
not NOT1 (N533, N525);
not NOT1 (N534, N529);
nand NAND4 (N535, N532, N485, N188, N39);
and AND4 (N536, N527, N92, N273, N463);
nor NOR3 (N537, N535, N112, N158);
or OR4 (N538, N537, N201, N141, N475);
or OR2 (N539, N512, N531);
nand NAND4 (N540, N387, N205, N197, N277);
not NOT1 (N541, N536);
xor XOR2 (N542, N528, N74);
and AND2 (N543, N541, N75);
nand NAND4 (N544, N530, N230, N334, N55);
and AND4 (N545, N544, N319, N163, N17);
nor NOR2 (N546, N533, N475);
nor NOR2 (N547, N542, N508);
and AND3 (N548, N307, N1, N44);
nand NAND4 (N549, N538, N235, N363, N469);
and AND3 (N550, N539, N455, N75);
and AND4 (N551, N545, N37, N258, N275);
nor NOR2 (N552, N547, N352);
nand NAND2 (N553, N549, N471);
and AND4 (N554, N543, N280, N504, N133);
nor NOR2 (N555, N550, N319);
xor XOR2 (N556, N553, N126);
nor NOR3 (N557, N552, N99, N33);
nor NOR3 (N558, N555, N467, N97);
buf BUF1 (N559, N551);
xor XOR2 (N560, N546, N142);
xor XOR2 (N561, N560, N21);
nand NAND3 (N562, N561, N4, N196);
and AND4 (N563, N554, N229, N464, N15);
buf BUF1 (N564, N558);
or OR4 (N565, N562, N346, N149, N303);
and AND2 (N566, N557, N68);
buf BUF1 (N567, N565);
not NOT1 (N568, N559);
or OR3 (N569, N567, N294, N297);
not NOT1 (N570, N564);
or OR2 (N571, N534, N284);
or OR3 (N572, N556, N69, N152);
not NOT1 (N573, N523);
nand NAND2 (N574, N568, N207);
nor NOR4 (N575, N573, N557, N21, N325);
nand NAND3 (N576, N572, N114, N10);
nor NOR3 (N577, N575, N30, N533);
nor NOR4 (N578, N577, N296, N108, N335);
xor XOR2 (N579, N566, N44);
or OR3 (N580, N570, N548, N242);
nand NAND3 (N581, N248, N29, N270);
not NOT1 (N582, N540);
nand NAND2 (N583, N571, N223);
not NOT1 (N584, N582);
or OR3 (N585, N581, N376, N255);
not NOT1 (N586, N584);
nand NAND4 (N587, N576, N147, N321, N64);
nor NOR4 (N588, N586, N226, N187, N99);
buf BUF1 (N589, N588);
nand NAND3 (N590, N585, N102, N108);
and AND4 (N591, N574, N16, N171, N448);
xor XOR2 (N592, N590, N548);
xor XOR2 (N593, N569, N239);
buf BUF1 (N594, N589);
xor XOR2 (N595, N594, N81);
buf BUF1 (N596, N593);
nor NOR4 (N597, N578, N474, N168, N500);
not NOT1 (N598, N579);
nand NAND2 (N599, N592, N399);
and AND3 (N600, N597, N151, N421);
nand NAND4 (N601, N595, N435, N14, N485);
and AND2 (N602, N601, N273);
not NOT1 (N603, N599);
and AND3 (N604, N583, N580, N343);
or OR2 (N605, N183, N179);
nor NOR2 (N606, N603, N352);
xor XOR2 (N607, N602, N160);
buf BUF1 (N608, N587);
and AND2 (N609, N606, N411);
buf BUF1 (N610, N591);
and AND2 (N611, N604, N164);
nand NAND2 (N612, N563, N343);
and AND2 (N613, N611, N289);
not NOT1 (N614, N605);
nand NAND4 (N615, N610, N298, N468, N147);
not NOT1 (N616, N613);
buf BUF1 (N617, N598);
xor XOR2 (N618, N616, N233);
or OR3 (N619, N600, N483, N254);
nand NAND3 (N620, N608, N235, N556);
xor XOR2 (N621, N620, N92);
not NOT1 (N622, N596);
and AND3 (N623, N622, N307, N132);
buf BUF1 (N624, N607);
buf BUF1 (N625, N619);
nor NOR4 (N626, N618, N445, N155, N222);
nand NAND3 (N627, N609, N521, N173);
and AND2 (N628, N617, N591);
xor XOR2 (N629, N627, N497);
nor NOR3 (N630, N615, N507, N552);
or OR3 (N631, N630, N618, N512);
nand NAND2 (N632, N614, N221);
not NOT1 (N633, N621);
or OR4 (N634, N628, N317, N548, N586);
or OR2 (N635, N624, N134);
and AND3 (N636, N631, N164, N447);
nor NOR3 (N637, N623, N589, N218);
nand NAND4 (N638, N637, N35, N165, N11);
not NOT1 (N639, N636);
nand NAND2 (N640, N612, N187);
xor XOR2 (N641, N640, N210);
nor NOR4 (N642, N626, N110, N102, N427);
nand NAND3 (N643, N635, N64, N529);
not NOT1 (N644, N638);
nor NOR4 (N645, N634, N480, N58, N621);
nor NOR2 (N646, N632, N149);
not NOT1 (N647, N639);
buf BUF1 (N648, N644);
and AND3 (N649, N647, N483, N88);
not NOT1 (N650, N642);
or OR3 (N651, N649, N572, N500);
not NOT1 (N652, N646);
and AND2 (N653, N643, N275);
xor XOR2 (N654, N653, N397);
nand NAND2 (N655, N629, N497);
buf BUF1 (N656, N650);
buf BUF1 (N657, N625);
buf BUF1 (N658, N633);
nor NOR2 (N659, N654, N221);
xor XOR2 (N660, N657, N73);
or OR2 (N661, N651, N91);
nor NOR4 (N662, N656, N41, N24, N267);
not NOT1 (N663, N662);
or OR2 (N664, N652, N136);
buf BUF1 (N665, N660);
nand NAND3 (N666, N661, N45, N521);
and AND2 (N667, N666, N655);
and AND2 (N668, N258, N636);
and AND3 (N669, N658, N28, N531);
or OR3 (N670, N659, N469, N32);
nand NAND3 (N671, N641, N76, N661);
not NOT1 (N672, N671);
xor XOR2 (N673, N670, N545);
not NOT1 (N674, N672);
nand NAND2 (N675, N673, N96);
nand NAND3 (N676, N665, N80, N616);
nor NOR4 (N677, N669, N380, N454, N514);
buf BUF1 (N678, N648);
and AND3 (N679, N675, N515, N156);
or OR2 (N680, N674, N373);
nand NAND2 (N681, N677, N258);
nand NAND2 (N682, N681, N179);
buf BUF1 (N683, N682);
not NOT1 (N684, N679);
not NOT1 (N685, N676);
buf BUF1 (N686, N664);
and AND3 (N687, N686, N595, N86);
buf BUF1 (N688, N678);
nand NAND3 (N689, N668, N671, N403);
and AND2 (N690, N689, N49);
and AND3 (N691, N645, N257, N538);
nor NOR2 (N692, N690, N164);
not NOT1 (N693, N680);
nand NAND4 (N694, N691, N331, N285, N496);
xor XOR2 (N695, N667, N363);
or OR4 (N696, N687, N632, N376, N337);
nor NOR2 (N697, N683, N434);
or OR4 (N698, N688, N640, N285, N153);
not NOT1 (N699, N696);
xor XOR2 (N700, N685, N241);
or OR3 (N701, N684, N128, N287);
nand NAND4 (N702, N701, N636, N109, N108);
not NOT1 (N703, N697);
nand NAND4 (N704, N702, N574, N237, N451);
not NOT1 (N705, N692);
nand NAND2 (N706, N705, N346);
buf BUF1 (N707, N699);
nand NAND2 (N708, N707, N131);
nor NOR2 (N709, N703, N431);
nor NOR3 (N710, N708, N596, N646);
buf BUF1 (N711, N709);
not NOT1 (N712, N711);
or OR4 (N713, N663, N571, N690, N13);
or OR3 (N714, N710, N168, N656);
not NOT1 (N715, N712);
buf BUF1 (N716, N698);
not NOT1 (N717, N714);
buf BUF1 (N718, N693);
nand NAND3 (N719, N718, N565, N2);
and AND3 (N720, N713, N455, N183);
or OR4 (N721, N716, N588, N588, N263);
xor XOR2 (N722, N695, N650);
and AND4 (N723, N700, N337, N200, N262);
or OR2 (N724, N722, N59);
not NOT1 (N725, N694);
or OR3 (N726, N723, N133, N708);
nand NAND2 (N727, N704, N373);
not NOT1 (N728, N727);
and AND2 (N729, N717, N406);
xor XOR2 (N730, N729, N134);
or OR3 (N731, N726, N725, N336);
and AND3 (N732, N293, N402, N573);
and AND4 (N733, N730, N57, N124, N451);
or OR3 (N734, N720, N595, N295);
nand NAND2 (N735, N732, N674);
nor NOR2 (N736, N733, N365);
buf BUF1 (N737, N735);
xor XOR2 (N738, N706, N21);
nand NAND2 (N739, N721, N4);
or OR4 (N740, N736, N604, N495, N109);
nor NOR3 (N741, N737, N546, N204);
nand NAND4 (N742, N741, N101, N181, N145);
nand NAND4 (N743, N728, N350, N123, N618);
not NOT1 (N744, N715);
and AND4 (N745, N739, N143, N78, N42);
and AND3 (N746, N744, N456, N674);
buf BUF1 (N747, N740);
and AND3 (N748, N734, N208, N318);
nor NOR2 (N749, N719, N199);
xor XOR2 (N750, N742, N71);
or OR4 (N751, N750, N114, N563, N376);
buf BUF1 (N752, N749);
buf BUF1 (N753, N743);
xor XOR2 (N754, N751, N107);
xor XOR2 (N755, N738, N159);
xor XOR2 (N756, N747, N394);
buf BUF1 (N757, N731);
and AND2 (N758, N753, N327);
nor NOR3 (N759, N746, N166, N211);
buf BUF1 (N760, N745);
not NOT1 (N761, N755);
buf BUF1 (N762, N754);
buf BUF1 (N763, N724);
buf BUF1 (N764, N760);
not NOT1 (N765, N758);
and AND4 (N766, N748, N205, N227, N425);
nand NAND2 (N767, N761, N97);
buf BUF1 (N768, N752);
buf BUF1 (N769, N762);
xor XOR2 (N770, N765, N99);
nand NAND4 (N771, N757, N623, N51, N121);
xor XOR2 (N772, N767, N155);
nand NAND4 (N773, N756, N658, N369, N541);
and AND2 (N774, N771, N73);
buf BUF1 (N775, N770);
and AND2 (N776, N763, N570);
buf BUF1 (N777, N768);
nand NAND3 (N778, N776, N457, N516);
xor XOR2 (N779, N769, N125);
not NOT1 (N780, N777);
nand NAND2 (N781, N766, N541);
not NOT1 (N782, N773);
not NOT1 (N783, N781);
and AND2 (N784, N772, N426);
and AND4 (N785, N780, N66, N598, N106);
nand NAND4 (N786, N774, N618, N579, N436);
xor XOR2 (N787, N784, N145);
buf BUF1 (N788, N779);
or OR3 (N789, N775, N450, N456);
not NOT1 (N790, N789);
buf BUF1 (N791, N790);
xor XOR2 (N792, N764, N572);
buf BUF1 (N793, N783);
or OR2 (N794, N778, N191);
or OR3 (N795, N786, N757, N618);
xor XOR2 (N796, N785, N244);
or OR4 (N797, N787, N662, N592, N324);
buf BUF1 (N798, N788);
and AND2 (N799, N792, N587);
or OR2 (N800, N791, N448);
buf BUF1 (N801, N795);
buf BUF1 (N802, N800);
xor XOR2 (N803, N802, N51);
not NOT1 (N804, N803);
not NOT1 (N805, N759);
xor XOR2 (N806, N797, N748);
not NOT1 (N807, N796);
nand NAND2 (N808, N793, N163);
not NOT1 (N809, N799);
xor XOR2 (N810, N808, N9);
xor XOR2 (N811, N806, N610);
and AND3 (N812, N798, N752, N165);
xor XOR2 (N813, N782, N686);
not NOT1 (N814, N801);
buf BUF1 (N815, N812);
nand NAND2 (N816, N815, N617);
not NOT1 (N817, N811);
nand NAND2 (N818, N817, N79);
and AND4 (N819, N814, N316, N323, N361);
nand NAND2 (N820, N805, N523);
and AND4 (N821, N819, N274, N611, N752);
nor NOR4 (N822, N810, N358, N10, N356);
not NOT1 (N823, N809);
xor XOR2 (N824, N816, N725);
xor XOR2 (N825, N822, N130);
nor NOR3 (N826, N823, N545, N641);
xor XOR2 (N827, N804, N269);
nand NAND2 (N828, N820, N658);
nor NOR2 (N829, N825, N8);
nor NOR3 (N830, N824, N88, N644);
not NOT1 (N831, N807);
or OR2 (N832, N826, N421);
nand NAND3 (N833, N830, N694, N229);
buf BUF1 (N834, N813);
not NOT1 (N835, N794);
buf BUF1 (N836, N828);
buf BUF1 (N837, N832);
nand NAND3 (N838, N833, N52, N720);
and AND2 (N839, N821, N185);
not NOT1 (N840, N829);
nor NOR3 (N841, N840, N142, N339);
nand NAND4 (N842, N837, N634, N466, N328);
not NOT1 (N843, N818);
buf BUF1 (N844, N843);
buf BUF1 (N845, N831);
not NOT1 (N846, N838);
not NOT1 (N847, N836);
or OR4 (N848, N844, N29, N122, N321);
xor XOR2 (N849, N835, N32);
or OR3 (N850, N849, N171, N41);
xor XOR2 (N851, N842, N95);
not NOT1 (N852, N847);
not NOT1 (N853, N839);
xor XOR2 (N854, N846, N597);
nand NAND3 (N855, N841, N381, N18);
nand NAND4 (N856, N827, N45, N92, N736);
not NOT1 (N857, N850);
and AND2 (N858, N853, N649);
buf BUF1 (N859, N855);
buf BUF1 (N860, N834);
and AND2 (N861, N860, N100);
xor XOR2 (N862, N858, N768);
xor XOR2 (N863, N848, N322);
xor XOR2 (N864, N856, N711);
xor XOR2 (N865, N863, N463);
buf BUF1 (N866, N851);
buf BUF1 (N867, N866);
nor NOR3 (N868, N861, N674, N536);
buf BUF1 (N869, N862);
xor XOR2 (N870, N868, N274);
nand NAND4 (N871, N852, N115, N811, N634);
and AND2 (N872, N867, N647);
nand NAND2 (N873, N872, N649);
or OR4 (N874, N859, N167, N302, N353);
nor NOR2 (N875, N854, N308);
and AND3 (N876, N869, N378, N587);
nor NOR3 (N877, N870, N643, N627);
xor XOR2 (N878, N864, N539);
not NOT1 (N879, N871);
or OR3 (N880, N865, N112, N658);
not NOT1 (N881, N857);
not NOT1 (N882, N878);
nor NOR4 (N883, N875, N90, N624, N849);
xor XOR2 (N884, N883, N554);
buf BUF1 (N885, N884);
not NOT1 (N886, N874);
nor NOR3 (N887, N877, N611, N876);
and AND3 (N888, N604, N357, N495);
or OR3 (N889, N888, N8, N544);
nand NAND3 (N890, N873, N689, N216);
nor NOR4 (N891, N882, N702, N228, N348);
nand NAND2 (N892, N879, N500);
not NOT1 (N893, N845);
nand NAND2 (N894, N891, N819);
nor NOR3 (N895, N886, N484, N672);
buf BUF1 (N896, N889);
not NOT1 (N897, N894);
or OR3 (N898, N885, N512, N440);
buf BUF1 (N899, N881);
or OR4 (N900, N896, N449, N856, N422);
or OR3 (N901, N880, N900, N576);
and AND4 (N902, N852, N469, N774, N189);
and AND3 (N903, N901, N310, N565);
nand NAND4 (N904, N897, N898, N593, N200);
buf BUF1 (N905, N13);
and AND2 (N906, N905, N200);
and AND2 (N907, N904, N522);
buf BUF1 (N908, N899);
nor NOR4 (N909, N890, N834, N290, N546);
buf BUF1 (N910, N895);
xor XOR2 (N911, N893, N670);
buf BUF1 (N912, N903);
and AND2 (N913, N906, N770);
buf BUF1 (N914, N902);
or OR4 (N915, N908, N439, N829, N614);
xor XOR2 (N916, N887, N191);
nor NOR2 (N917, N915, N624);
or OR3 (N918, N910, N459, N860);
nor NOR3 (N919, N892, N599, N317);
nor NOR4 (N920, N919, N532, N816, N825);
buf BUF1 (N921, N911);
or OR3 (N922, N907, N863, N144);
xor XOR2 (N923, N918, N166);
or OR3 (N924, N916, N250, N274);
xor XOR2 (N925, N922, N105);
buf BUF1 (N926, N909);
and AND4 (N927, N926, N62, N880, N675);
and AND2 (N928, N913, N446);
nand NAND3 (N929, N914, N649, N560);
and AND2 (N930, N912, N205);
and AND4 (N931, N924, N639, N468, N11);
nand NAND4 (N932, N929, N102, N873, N411);
and AND3 (N933, N928, N377, N487);
or OR2 (N934, N927, N713);
xor XOR2 (N935, N923, N747);
nand NAND4 (N936, N934, N530, N335, N884);
or OR4 (N937, N925, N785, N629, N510);
nand NAND4 (N938, N921, N893, N531, N537);
nor NOR2 (N939, N917, N878);
not NOT1 (N940, N920);
xor XOR2 (N941, N938, N554);
nor NOR2 (N942, N940, N320);
not NOT1 (N943, N941);
xor XOR2 (N944, N936, N520);
not NOT1 (N945, N942);
nand NAND2 (N946, N935, N723);
nor NOR2 (N947, N945, N692);
buf BUF1 (N948, N937);
or OR4 (N949, N948, N473, N389, N924);
xor XOR2 (N950, N930, N935);
or OR2 (N951, N944, N75);
or OR2 (N952, N931, N470);
and AND4 (N953, N947, N833, N233, N942);
not NOT1 (N954, N939);
not NOT1 (N955, N954);
not NOT1 (N956, N946);
or OR4 (N957, N951, N855, N497, N711);
buf BUF1 (N958, N949);
or OR3 (N959, N957, N636, N613);
buf BUF1 (N960, N958);
xor XOR2 (N961, N932, N566);
or OR4 (N962, N933, N197, N462, N241);
not NOT1 (N963, N950);
and AND4 (N964, N959, N862, N670, N459);
not NOT1 (N965, N956);
xor XOR2 (N966, N960, N157);
and AND3 (N967, N961, N937, N546);
nor NOR2 (N968, N962, N22);
xor XOR2 (N969, N968, N19);
nor NOR3 (N970, N966, N616, N936);
not NOT1 (N971, N970);
buf BUF1 (N972, N963);
and AND2 (N973, N969, N493);
buf BUF1 (N974, N943);
not NOT1 (N975, N953);
or OR2 (N976, N952, N451);
buf BUF1 (N977, N975);
nand NAND2 (N978, N974, N420);
xor XOR2 (N979, N978, N789);
or OR4 (N980, N977, N636, N725, N292);
or OR4 (N981, N967, N61, N270, N589);
not NOT1 (N982, N972);
and AND2 (N983, N973, N438);
or OR2 (N984, N979, N738);
and AND2 (N985, N984, N855);
nand NAND3 (N986, N983, N395, N862);
not NOT1 (N987, N981);
not NOT1 (N988, N987);
buf BUF1 (N989, N971);
not NOT1 (N990, N986);
buf BUF1 (N991, N989);
not NOT1 (N992, N964);
xor XOR2 (N993, N980, N727);
nand NAND2 (N994, N990, N852);
and AND3 (N995, N985, N534, N774);
nor NOR2 (N996, N982, N511);
not NOT1 (N997, N991);
and AND3 (N998, N992, N460, N335);
and AND4 (N999, N997, N911, N608, N505);
or OR4 (N1000, N965, N444, N206, N303);
buf BUF1 (N1001, N996);
not NOT1 (N1002, N999);
nor NOR2 (N1003, N993, N179);
not NOT1 (N1004, N1000);
buf BUF1 (N1005, N988);
buf BUF1 (N1006, N994);
not NOT1 (N1007, N995);
nand NAND3 (N1008, N1001, N249, N652);
not NOT1 (N1009, N1008);
and AND2 (N1010, N955, N30);
or OR4 (N1011, N1005, N845, N228, N894);
xor XOR2 (N1012, N1003, N326);
nor NOR4 (N1013, N1009, N781, N29, N509);
nand NAND3 (N1014, N976, N240, N984);
and AND3 (N1015, N1014, N236, N53);
and AND2 (N1016, N1007, N784);
xor XOR2 (N1017, N1012, N309);
xor XOR2 (N1018, N1006, N281);
and AND2 (N1019, N1011, N70);
or OR2 (N1020, N1019, N243);
and AND3 (N1021, N1010, N564, N380);
and AND3 (N1022, N1013, N805, N703);
nand NAND3 (N1023, N1022, N744, N463);
xor XOR2 (N1024, N1020, N540);
or OR4 (N1025, N1004, N328, N613, N828);
and AND2 (N1026, N1025, N586);
not NOT1 (N1027, N1023);
and AND3 (N1028, N1026, N148, N652);
and AND2 (N1029, N998, N936);
nand NAND2 (N1030, N1021, N920);
nand NAND3 (N1031, N1017, N342, N291);
buf BUF1 (N1032, N1016);
buf BUF1 (N1033, N1024);
or OR2 (N1034, N1032, N267);
not NOT1 (N1035, N1027);
not NOT1 (N1036, N1002);
nor NOR3 (N1037, N1015, N271, N239);
not NOT1 (N1038, N1018);
or OR3 (N1039, N1031, N459, N624);
or OR4 (N1040, N1035, N805, N353, N694);
nor NOR2 (N1041, N1040, N59);
nand NAND4 (N1042, N1029, N671, N690, N350);
nor NOR4 (N1043, N1042, N518, N857, N589);
not NOT1 (N1044, N1043);
nand NAND3 (N1045, N1034, N133, N413);
nand NAND2 (N1046, N1045, N230);
nand NAND4 (N1047, N1037, N370, N303, N417);
nand NAND2 (N1048, N1047, N725);
nor NOR4 (N1049, N1036, N126, N54, N1005);
not NOT1 (N1050, N1038);
and AND2 (N1051, N1048, N902);
xor XOR2 (N1052, N1041, N867);
and AND2 (N1053, N1051, N994);
and AND2 (N1054, N1033, N651);
not NOT1 (N1055, N1053);
buf BUF1 (N1056, N1054);
nor NOR2 (N1057, N1049, N215);
or OR4 (N1058, N1052, N772, N178, N391);
or OR2 (N1059, N1046, N361);
not NOT1 (N1060, N1030);
and AND2 (N1061, N1055, N236);
xor XOR2 (N1062, N1058, N825);
xor XOR2 (N1063, N1059, N268);
and AND4 (N1064, N1044, N393, N419, N637);
nand NAND2 (N1065, N1061, N200);
and AND2 (N1066, N1050, N656);
and AND4 (N1067, N1065, N198, N846, N267);
buf BUF1 (N1068, N1066);
nor NOR2 (N1069, N1060, N405);
and AND4 (N1070, N1028, N303, N300, N774);
buf BUF1 (N1071, N1062);
xor XOR2 (N1072, N1057, N108);
xor XOR2 (N1073, N1068, N991);
nand NAND3 (N1074, N1073, N18, N309);
xor XOR2 (N1075, N1063, N351);
not NOT1 (N1076, N1070);
buf BUF1 (N1077, N1069);
or OR3 (N1078, N1072, N327, N860);
not NOT1 (N1079, N1078);
nor NOR3 (N1080, N1074, N40, N123);
buf BUF1 (N1081, N1071);
and AND3 (N1082, N1056, N325, N1016);
xor XOR2 (N1083, N1079, N1046);
buf BUF1 (N1084, N1076);
and AND2 (N1085, N1067, N15);
xor XOR2 (N1086, N1064, N188);
not NOT1 (N1087, N1077);
or OR3 (N1088, N1080, N60, N637);
not NOT1 (N1089, N1082);
or OR4 (N1090, N1075, N228, N791, N648);
buf BUF1 (N1091, N1085);
not NOT1 (N1092, N1090);
nor NOR4 (N1093, N1092, N805, N343, N943);
or OR3 (N1094, N1091, N654, N165);
not NOT1 (N1095, N1093);
xor XOR2 (N1096, N1083, N533);
xor XOR2 (N1097, N1088, N563);
xor XOR2 (N1098, N1039, N83);
or OR2 (N1099, N1096, N31);
nor NOR2 (N1100, N1099, N842);
nand NAND4 (N1101, N1086, N829, N109, N1079);
not NOT1 (N1102, N1101);
and AND4 (N1103, N1089, N864, N758, N518);
buf BUF1 (N1104, N1094);
xor XOR2 (N1105, N1098, N263);
or OR4 (N1106, N1081, N1002, N381, N30);
not NOT1 (N1107, N1106);
not NOT1 (N1108, N1107);
and AND3 (N1109, N1103, N185, N1065);
and AND4 (N1110, N1108, N226, N871, N843);
nand NAND2 (N1111, N1102, N274);
or OR2 (N1112, N1097, N463);
xor XOR2 (N1113, N1100, N448);
nor NOR4 (N1114, N1109, N324, N1029, N358);
or OR3 (N1115, N1104, N688, N265);
nor NOR3 (N1116, N1111, N1001, N888);
xor XOR2 (N1117, N1112, N672);
nor NOR2 (N1118, N1113, N1103);
nor NOR3 (N1119, N1087, N124, N5);
not NOT1 (N1120, N1105);
not NOT1 (N1121, N1119);
nand NAND4 (N1122, N1121, N1072, N635, N727);
nor NOR2 (N1123, N1084, N107);
buf BUF1 (N1124, N1122);
nand NAND3 (N1125, N1123, N719, N850);
buf BUF1 (N1126, N1125);
or OR2 (N1127, N1118, N385);
nor NOR2 (N1128, N1127, N399);
and AND4 (N1129, N1117, N333, N498, N936);
nor NOR2 (N1130, N1116, N629);
xor XOR2 (N1131, N1120, N775);
and AND2 (N1132, N1131, N1053);
nand NAND2 (N1133, N1126, N363);
buf BUF1 (N1134, N1128);
not NOT1 (N1135, N1132);
or OR4 (N1136, N1124, N79, N705, N952);
not NOT1 (N1137, N1129);
nor NOR4 (N1138, N1134, N581, N835, N947);
nor NOR2 (N1139, N1110, N750);
xor XOR2 (N1140, N1139, N610);
xor XOR2 (N1141, N1130, N351);
and AND4 (N1142, N1136, N831, N311, N886);
or OR3 (N1143, N1095, N296, N549);
xor XOR2 (N1144, N1138, N583);
nor NOR2 (N1145, N1141, N513);
or OR2 (N1146, N1133, N950);
or OR2 (N1147, N1114, N985);
and AND2 (N1148, N1145, N504);
xor XOR2 (N1149, N1135, N524);
not NOT1 (N1150, N1148);
not NOT1 (N1151, N1115);
nor NOR2 (N1152, N1137, N81);
nand NAND3 (N1153, N1146, N498, N649);
xor XOR2 (N1154, N1142, N664);
nor NOR4 (N1155, N1150, N1081, N1036, N752);
and AND4 (N1156, N1153, N570, N964, N187);
xor XOR2 (N1157, N1155, N218);
nand NAND3 (N1158, N1157, N290, N856);
and AND2 (N1159, N1143, N326);
and AND2 (N1160, N1149, N549);
not NOT1 (N1161, N1144);
nand NAND4 (N1162, N1152, N905, N854, N549);
nand NAND4 (N1163, N1147, N168, N1083, N1148);
or OR4 (N1164, N1159, N246, N910, N589);
nand NAND4 (N1165, N1163, N408, N728, N436);
not NOT1 (N1166, N1156);
xor XOR2 (N1167, N1162, N1149);
not NOT1 (N1168, N1160);
or OR2 (N1169, N1154, N117);
buf BUF1 (N1170, N1140);
buf BUF1 (N1171, N1161);
nor NOR3 (N1172, N1168, N638, N75);
or OR2 (N1173, N1158, N419);
nor NOR2 (N1174, N1169, N522);
nor NOR4 (N1175, N1172, N64, N291, N1149);
nand NAND3 (N1176, N1151, N816, N939);
or OR3 (N1177, N1164, N446, N1102);
xor XOR2 (N1178, N1167, N775);
not NOT1 (N1179, N1174);
or OR3 (N1180, N1165, N771, N313);
not NOT1 (N1181, N1170);
buf BUF1 (N1182, N1175);
nand NAND3 (N1183, N1166, N1089, N749);
nor NOR4 (N1184, N1176, N770, N1143, N298);
nor NOR3 (N1185, N1181, N266, N304);
buf BUF1 (N1186, N1177);
nor NOR2 (N1187, N1179, N245);
and AND2 (N1188, N1186, N1173);
or OR3 (N1189, N418, N49, N609);
not NOT1 (N1190, N1184);
not NOT1 (N1191, N1187);
not NOT1 (N1192, N1189);
buf BUF1 (N1193, N1188);
buf BUF1 (N1194, N1171);
and AND4 (N1195, N1194, N475, N1011, N493);
xor XOR2 (N1196, N1195, N548);
buf BUF1 (N1197, N1191);
nand NAND4 (N1198, N1192, N604, N156, N71);
xor XOR2 (N1199, N1198, N810);
buf BUF1 (N1200, N1190);
xor XOR2 (N1201, N1185, N8);
xor XOR2 (N1202, N1199, N444);
nor NOR4 (N1203, N1197, N240, N1145, N256);
and AND2 (N1204, N1202, N919);
nand NAND2 (N1205, N1204, N75);
nand NAND3 (N1206, N1193, N361, N921);
not NOT1 (N1207, N1182);
or OR4 (N1208, N1206, N608, N1046, N532);
and AND4 (N1209, N1180, N728, N1117, N172);
nand NAND2 (N1210, N1183, N237);
not NOT1 (N1211, N1203);
buf BUF1 (N1212, N1210);
or OR4 (N1213, N1209, N697, N279, N68);
xor XOR2 (N1214, N1208, N115);
xor XOR2 (N1215, N1201, N384);
and AND3 (N1216, N1212, N1190, N1082);
not NOT1 (N1217, N1216);
nand NAND2 (N1218, N1214, N799);
nor NOR3 (N1219, N1205, N1102, N779);
nor NOR4 (N1220, N1217, N267, N1, N1117);
buf BUF1 (N1221, N1196);
nand NAND3 (N1222, N1211, N148, N123);
not NOT1 (N1223, N1200);
or OR2 (N1224, N1219, N283);
nand NAND3 (N1225, N1222, N12, N838);
nor NOR2 (N1226, N1215, N618);
and AND4 (N1227, N1226, N64, N959, N396);
not NOT1 (N1228, N1221);
xor XOR2 (N1229, N1227, N1016);
or OR2 (N1230, N1178, N773);
nor NOR3 (N1231, N1218, N896, N1192);
nor NOR3 (N1232, N1231, N185, N989);
xor XOR2 (N1233, N1230, N707);
or OR4 (N1234, N1223, N692, N89, N79);
xor XOR2 (N1235, N1213, N65);
nand NAND4 (N1236, N1233, N1191, N883, N636);
xor XOR2 (N1237, N1207, N744);
and AND4 (N1238, N1220, N364, N919, N677);
xor XOR2 (N1239, N1234, N1218);
and AND3 (N1240, N1235, N994, N350);
nor NOR3 (N1241, N1238, N838, N46);
xor XOR2 (N1242, N1229, N812);
and AND3 (N1243, N1232, N346, N204);
nor NOR3 (N1244, N1243, N517, N869);
buf BUF1 (N1245, N1244);
nand NAND2 (N1246, N1225, N134);
nand NAND2 (N1247, N1242, N265);
nand NAND3 (N1248, N1239, N1, N459);
xor XOR2 (N1249, N1237, N628);
and AND2 (N1250, N1247, N998);
and AND4 (N1251, N1250, N807, N1079, N779);
xor XOR2 (N1252, N1241, N831);
not NOT1 (N1253, N1228);
or OR3 (N1254, N1252, N140, N548);
nor NOR2 (N1255, N1224, N823);
not NOT1 (N1256, N1248);
nand NAND2 (N1257, N1246, N550);
not NOT1 (N1258, N1255);
or OR3 (N1259, N1240, N195, N510);
xor XOR2 (N1260, N1251, N635);
and AND2 (N1261, N1245, N702);
xor XOR2 (N1262, N1257, N1123);
xor XOR2 (N1263, N1258, N34);
xor XOR2 (N1264, N1261, N841);
buf BUF1 (N1265, N1256);
or OR2 (N1266, N1262, N808);
nor NOR3 (N1267, N1263, N900, N923);
nor NOR2 (N1268, N1259, N817);
or OR2 (N1269, N1236, N202);
nor NOR4 (N1270, N1249, N648, N1106, N4);
nand NAND3 (N1271, N1265, N872, N985);
nand NAND3 (N1272, N1254, N646, N545);
and AND3 (N1273, N1270, N869, N1083);
nor NOR4 (N1274, N1260, N124, N1080, N422);
or OR2 (N1275, N1268, N921);
xor XOR2 (N1276, N1266, N994);
and AND4 (N1277, N1253, N329, N865, N518);
not NOT1 (N1278, N1273);
nand NAND4 (N1279, N1264, N126, N592, N452);
nand NAND2 (N1280, N1267, N1162);
buf BUF1 (N1281, N1277);
buf BUF1 (N1282, N1276);
nand NAND2 (N1283, N1279, N1119);
nand NAND3 (N1284, N1275, N1132, N954);
or OR4 (N1285, N1274, N391, N659, N749);
not NOT1 (N1286, N1269);
nor NOR2 (N1287, N1272, N342);
nand NAND2 (N1288, N1282, N602);
or OR2 (N1289, N1286, N918);
nor NOR4 (N1290, N1289, N708, N712, N1030);
buf BUF1 (N1291, N1288);
or OR2 (N1292, N1287, N1210);
nand NAND2 (N1293, N1278, N218);
and AND3 (N1294, N1285, N502, N982);
buf BUF1 (N1295, N1292);
not NOT1 (N1296, N1295);
xor XOR2 (N1297, N1293, N331);
nand NAND4 (N1298, N1271, N1245, N1099, N818);
nor NOR3 (N1299, N1280, N985, N762);
or OR2 (N1300, N1283, N8);
buf BUF1 (N1301, N1299);
xor XOR2 (N1302, N1291, N612);
or OR4 (N1303, N1300, N398, N526, N819);
nand NAND4 (N1304, N1294, N513, N1300, N943);
nand NAND2 (N1305, N1290, N118);
xor XOR2 (N1306, N1301, N519);
not NOT1 (N1307, N1305);
xor XOR2 (N1308, N1296, N774);
nor NOR4 (N1309, N1297, N995, N1010, N78);
nand NAND2 (N1310, N1284, N461);
or OR3 (N1311, N1304, N603, N1074);
and AND4 (N1312, N1310, N880, N1128, N712);
xor XOR2 (N1313, N1309, N523);
or OR4 (N1314, N1308, N540, N1165, N360);
and AND4 (N1315, N1311, N893, N539, N161);
xor XOR2 (N1316, N1302, N1220);
or OR2 (N1317, N1303, N1276);
or OR4 (N1318, N1281, N497, N275, N912);
buf BUF1 (N1319, N1312);
nor NOR4 (N1320, N1316, N978, N38, N605);
and AND3 (N1321, N1317, N696, N583);
or OR4 (N1322, N1318, N530, N202, N72);
or OR2 (N1323, N1321, N881);
nand NAND4 (N1324, N1313, N453, N815, N1176);
buf BUF1 (N1325, N1307);
buf BUF1 (N1326, N1323);
or OR2 (N1327, N1314, N977);
or OR2 (N1328, N1326, N790);
buf BUF1 (N1329, N1315);
nand NAND2 (N1330, N1319, N355);
buf BUF1 (N1331, N1328);
and AND2 (N1332, N1327, N695);
xor XOR2 (N1333, N1331, N828);
and AND4 (N1334, N1324, N1117, N1208, N295);
xor XOR2 (N1335, N1334, N623);
or OR3 (N1336, N1325, N678, N864);
buf BUF1 (N1337, N1322);
and AND2 (N1338, N1320, N548);
nor NOR2 (N1339, N1336, N536);
or OR4 (N1340, N1329, N625, N868, N690);
nand NAND2 (N1341, N1335, N267);
nor NOR2 (N1342, N1339, N1078);
xor XOR2 (N1343, N1332, N395);
and AND3 (N1344, N1338, N115, N1249);
buf BUF1 (N1345, N1341);
buf BUF1 (N1346, N1337);
and AND3 (N1347, N1340, N1030, N946);
and AND4 (N1348, N1345, N313, N218, N49);
not NOT1 (N1349, N1306);
or OR4 (N1350, N1330, N760, N97, N278);
not NOT1 (N1351, N1346);
nor NOR3 (N1352, N1350, N106, N773);
nand NAND3 (N1353, N1347, N1079, N817);
xor XOR2 (N1354, N1348, N879);
nor NOR3 (N1355, N1342, N328, N801);
nor NOR3 (N1356, N1353, N1220, N271);
nor NOR2 (N1357, N1344, N685);
nand NAND2 (N1358, N1298, N78);
nand NAND3 (N1359, N1355, N653, N207);
not NOT1 (N1360, N1358);
not NOT1 (N1361, N1352);
and AND2 (N1362, N1343, N525);
and AND4 (N1363, N1333, N464, N9, N1020);
or OR4 (N1364, N1360, N451, N362, N771);
not NOT1 (N1365, N1362);
nor NOR4 (N1366, N1364, N560, N38, N953);
and AND3 (N1367, N1357, N292, N1141);
not NOT1 (N1368, N1361);
nand NAND2 (N1369, N1363, N313);
and AND2 (N1370, N1356, N1316);
or OR3 (N1371, N1365, N302, N499);
not NOT1 (N1372, N1370);
not NOT1 (N1373, N1369);
nand NAND2 (N1374, N1349, N464);
nor NOR4 (N1375, N1374, N851, N75, N1259);
or OR3 (N1376, N1371, N1317, N166);
nand NAND3 (N1377, N1375, N194, N973);
nor NOR3 (N1378, N1359, N833, N811);
nand NAND4 (N1379, N1368, N3, N500, N468);
nor NOR4 (N1380, N1366, N731, N612, N510);
not NOT1 (N1381, N1367);
nand NAND2 (N1382, N1380, N677);
not NOT1 (N1383, N1379);
and AND4 (N1384, N1376, N209, N648, N351);
buf BUF1 (N1385, N1351);
nor NOR2 (N1386, N1381, N736);
nand NAND2 (N1387, N1354, N785);
buf BUF1 (N1388, N1373);
nor NOR2 (N1389, N1387, N1304);
not NOT1 (N1390, N1372);
nand NAND4 (N1391, N1385, N627, N1139, N1224);
or OR3 (N1392, N1390, N1039, N1225);
or OR4 (N1393, N1377, N1249, N173, N267);
or OR3 (N1394, N1389, N872, N222);
nor NOR2 (N1395, N1384, N1341);
or OR4 (N1396, N1393, N1138, N894, N464);
or OR3 (N1397, N1388, N818, N1256);
or OR2 (N1398, N1383, N720);
nand NAND2 (N1399, N1386, N1189);
nand NAND2 (N1400, N1392, N657);
not NOT1 (N1401, N1378);
or OR2 (N1402, N1400, N198);
nand NAND3 (N1403, N1399, N1378, N289);
nor NOR4 (N1404, N1403, N1191, N1334, N251);
buf BUF1 (N1405, N1401);
xor XOR2 (N1406, N1395, N955);
not NOT1 (N1407, N1391);
nor NOR4 (N1408, N1396, N192, N150, N1392);
not NOT1 (N1409, N1397);
and AND4 (N1410, N1404, N650, N132, N1257);
nand NAND2 (N1411, N1410, N1189);
nand NAND4 (N1412, N1406, N307, N468, N54);
nand NAND3 (N1413, N1411, N916, N1127);
buf BUF1 (N1414, N1409);
xor XOR2 (N1415, N1382, N151);
and AND2 (N1416, N1413, N639);
buf BUF1 (N1417, N1398);
nand NAND2 (N1418, N1407, N703);
nand NAND2 (N1419, N1415, N961);
and AND2 (N1420, N1408, N357);
or OR4 (N1421, N1414, N1296, N1302, N187);
nand NAND2 (N1422, N1419, N481);
nor NOR3 (N1423, N1416, N1229, N1259);
nor NOR3 (N1424, N1421, N30, N1178);
nor NOR4 (N1425, N1420, N626, N1261, N35);
nor NOR3 (N1426, N1412, N289, N1326);
or OR4 (N1427, N1417, N1355, N1125, N606);
buf BUF1 (N1428, N1394);
buf BUF1 (N1429, N1424);
not NOT1 (N1430, N1423);
nand NAND2 (N1431, N1430, N78);
nor NOR4 (N1432, N1428, N391, N896, N901);
nand NAND3 (N1433, N1402, N337, N741);
and AND4 (N1434, N1431, N521, N887, N696);
and AND4 (N1435, N1426, N682, N963, N933);
nor NOR4 (N1436, N1422, N1391, N150, N410);
buf BUF1 (N1437, N1432);
or OR4 (N1438, N1429, N110, N155, N69);
nand NAND3 (N1439, N1438, N15, N1230);
nand NAND4 (N1440, N1435, N1199, N596, N152);
xor XOR2 (N1441, N1433, N63);
nor NOR2 (N1442, N1441, N761);
xor XOR2 (N1443, N1425, N1072);
not NOT1 (N1444, N1440);
and AND2 (N1445, N1418, N1204);
and AND3 (N1446, N1439, N1302, N1062);
nor NOR4 (N1447, N1427, N261, N768, N1016);
not NOT1 (N1448, N1447);
nor NOR3 (N1449, N1442, N1429, N348);
or OR3 (N1450, N1448, N151, N588);
buf BUF1 (N1451, N1437);
xor XOR2 (N1452, N1451, N1141);
and AND2 (N1453, N1436, N1295);
or OR3 (N1454, N1450, N1181, N1337);
not NOT1 (N1455, N1449);
xor XOR2 (N1456, N1455, N11);
and AND2 (N1457, N1453, N180);
buf BUF1 (N1458, N1434);
nand NAND4 (N1459, N1456, N1188, N777, N1435);
not NOT1 (N1460, N1405);
and AND3 (N1461, N1459, N222, N283);
not NOT1 (N1462, N1458);
buf BUF1 (N1463, N1443);
not NOT1 (N1464, N1463);
xor XOR2 (N1465, N1464, N1193);
and AND4 (N1466, N1446, N1374, N45, N166);
or OR4 (N1467, N1462, N315, N715, N511);
or OR2 (N1468, N1466, N68);
and AND3 (N1469, N1465, N842, N1365);
nand NAND2 (N1470, N1444, N266);
nor NOR3 (N1471, N1452, N331, N726);
not NOT1 (N1472, N1470);
buf BUF1 (N1473, N1454);
nand NAND3 (N1474, N1471, N976, N1218);
not NOT1 (N1475, N1473);
buf BUF1 (N1476, N1475);
not NOT1 (N1477, N1468);
nor NOR2 (N1478, N1445, N993);
not NOT1 (N1479, N1476);
buf BUF1 (N1480, N1479);
nor NOR4 (N1481, N1457, N1334, N192, N538);
buf BUF1 (N1482, N1480);
and AND2 (N1483, N1477, N690);
and AND2 (N1484, N1483, N179);
nor NOR3 (N1485, N1481, N953, N650);
or OR2 (N1486, N1467, N1334);
not NOT1 (N1487, N1461);
and AND3 (N1488, N1460, N6, N1165);
buf BUF1 (N1489, N1472);
nor NOR2 (N1490, N1487, N737);
xor XOR2 (N1491, N1484, N219);
xor XOR2 (N1492, N1482, N143);
xor XOR2 (N1493, N1469, N690);
nand NAND2 (N1494, N1490, N1418);
xor XOR2 (N1495, N1474, N1464);
or OR2 (N1496, N1488, N1103);
or OR4 (N1497, N1493, N1097, N86, N1094);
xor XOR2 (N1498, N1491, N1432);
buf BUF1 (N1499, N1478);
nand NAND3 (N1500, N1486, N1336, N424);
nor NOR3 (N1501, N1498, N450, N1182);
xor XOR2 (N1502, N1492, N807);
buf BUF1 (N1503, N1496);
not NOT1 (N1504, N1494);
nor NOR3 (N1505, N1500, N1321, N186);
xor XOR2 (N1506, N1505, N964);
and AND2 (N1507, N1503, N16);
and AND2 (N1508, N1506, N495);
or OR4 (N1509, N1499, N55, N1469, N457);
not NOT1 (N1510, N1489);
not NOT1 (N1511, N1510);
or OR4 (N1512, N1509, N592, N107, N1164);
buf BUF1 (N1513, N1507);
not NOT1 (N1514, N1508);
buf BUF1 (N1515, N1514);
xor XOR2 (N1516, N1513, N564);
nor NOR4 (N1517, N1504, N857, N524, N1163);
or OR3 (N1518, N1516, N521, N675);
xor XOR2 (N1519, N1515, N402);
xor XOR2 (N1520, N1502, N1004);
or OR3 (N1521, N1495, N622, N1147);
nand NAND3 (N1522, N1519, N294, N373);
and AND2 (N1523, N1518, N784);
nor NOR3 (N1524, N1517, N1461, N871);
xor XOR2 (N1525, N1521, N1390);
and AND2 (N1526, N1524, N1360);
and AND4 (N1527, N1485, N428, N879, N147);
nor NOR4 (N1528, N1520, N1424, N276, N81);
and AND2 (N1529, N1511, N54);
or OR2 (N1530, N1523, N709);
xor XOR2 (N1531, N1522, N574);
not NOT1 (N1532, N1531);
nand NAND4 (N1533, N1526, N682, N516, N1326);
xor XOR2 (N1534, N1501, N935);
xor XOR2 (N1535, N1530, N919);
buf BUF1 (N1536, N1525);
or OR2 (N1537, N1532, N389);
or OR4 (N1538, N1528, N46, N116, N1372);
xor XOR2 (N1539, N1533, N1110);
nor NOR3 (N1540, N1497, N983, N336);
not NOT1 (N1541, N1537);
nor NOR2 (N1542, N1535, N1410);
not NOT1 (N1543, N1512);
nor NOR4 (N1544, N1538, N1433, N1316, N1046);
nor NOR4 (N1545, N1534, N959, N1313, N208);
buf BUF1 (N1546, N1543);
or OR4 (N1547, N1540, N745, N889, N367);
xor XOR2 (N1548, N1547, N283);
not NOT1 (N1549, N1536);
nor NOR3 (N1550, N1541, N1497, N1273);
and AND3 (N1551, N1548, N565, N794);
nand NAND3 (N1552, N1529, N41, N459);
and AND2 (N1553, N1542, N1101);
nor NOR3 (N1554, N1539, N1412, N1032);
nand NAND4 (N1555, N1554, N1434, N701, N1418);
or OR3 (N1556, N1551, N688, N541);
nand NAND3 (N1557, N1555, N419, N363);
and AND4 (N1558, N1556, N657, N1128, N595);
nor NOR2 (N1559, N1557, N214);
nand NAND3 (N1560, N1552, N1519, N906);
and AND4 (N1561, N1545, N770, N310, N1018);
nand NAND2 (N1562, N1559, N583);
nand NAND2 (N1563, N1553, N496);
or OR4 (N1564, N1562, N668, N366, N265);
buf BUF1 (N1565, N1558);
buf BUF1 (N1566, N1561);
or OR3 (N1567, N1560, N763, N1513);
not NOT1 (N1568, N1550);
xor XOR2 (N1569, N1568, N1397);
or OR3 (N1570, N1527, N912, N1215);
not NOT1 (N1571, N1544);
not NOT1 (N1572, N1563);
nor NOR3 (N1573, N1572, N704, N2);
nand NAND4 (N1574, N1571, N430, N829, N1016);
nand NAND2 (N1575, N1573, N570);
buf BUF1 (N1576, N1565);
and AND3 (N1577, N1570, N331, N674);
not NOT1 (N1578, N1549);
nand NAND3 (N1579, N1577, N1081, N172);
buf BUF1 (N1580, N1579);
buf BUF1 (N1581, N1566);
nand NAND4 (N1582, N1567, N818, N762, N897);
and AND2 (N1583, N1574, N891);
not NOT1 (N1584, N1564);
xor XOR2 (N1585, N1578, N928);
and AND4 (N1586, N1546, N902, N1002, N1528);
not NOT1 (N1587, N1576);
and AND3 (N1588, N1569, N191, N1269);
xor XOR2 (N1589, N1585, N921);
nor NOR4 (N1590, N1587, N1403, N1354, N530);
or OR4 (N1591, N1586, N207, N1053, N1505);
or OR2 (N1592, N1581, N180);
not NOT1 (N1593, N1591);
not NOT1 (N1594, N1580);
and AND3 (N1595, N1592, N842, N42);
buf BUF1 (N1596, N1594);
nand NAND3 (N1597, N1583, N1330, N1007);
buf BUF1 (N1598, N1595);
and AND2 (N1599, N1593, N870);
nand NAND3 (N1600, N1589, N1236, N602);
buf BUF1 (N1601, N1590);
nand NAND2 (N1602, N1588, N1057);
and AND2 (N1603, N1575, N888);
buf BUF1 (N1604, N1596);
nand NAND4 (N1605, N1599, N826, N1417, N339);
buf BUF1 (N1606, N1604);
buf BUF1 (N1607, N1584);
nor NOR2 (N1608, N1603, N991);
not NOT1 (N1609, N1608);
and AND2 (N1610, N1609, N987);
and AND2 (N1611, N1607, N202);
not NOT1 (N1612, N1601);
nand NAND2 (N1613, N1582, N1166);
buf BUF1 (N1614, N1613);
and AND2 (N1615, N1612, N1097);
nor NOR3 (N1616, N1611, N735, N642);
not NOT1 (N1617, N1606);
xor XOR2 (N1618, N1616, N1586);
xor XOR2 (N1619, N1597, N784);
nand NAND2 (N1620, N1598, N1238);
xor XOR2 (N1621, N1605, N1341);
nand NAND3 (N1622, N1600, N583, N385);
and AND3 (N1623, N1618, N80, N697);
or OR3 (N1624, N1614, N832, N1580);
not NOT1 (N1625, N1619);
xor XOR2 (N1626, N1617, N812);
not NOT1 (N1627, N1625);
buf BUF1 (N1628, N1623);
buf BUF1 (N1629, N1628);
nand NAND2 (N1630, N1610, N593);
not NOT1 (N1631, N1615);
xor XOR2 (N1632, N1622, N244);
buf BUF1 (N1633, N1629);
nand NAND4 (N1634, N1602, N219, N19, N280);
and AND2 (N1635, N1630, N1228);
and AND3 (N1636, N1635, N83, N1448);
buf BUF1 (N1637, N1624);
or OR2 (N1638, N1621, N196);
xor XOR2 (N1639, N1633, N1463);
xor XOR2 (N1640, N1634, N432);
nor NOR4 (N1641, N1631, N770, N987, N533);
or OR3 (N1642, N1636, N1398, N302);
or OR2 (N1643, N1642, N815);
nor NOR3 (N1644, N1640, N350, N208);
or OR2 (N1645, N1638, N556);
and AND3 (N1646, N1627, N786, N272);
or OR4 (N1647, N1637, N1041, N1332, N595);
not NOT1 (N1648, N1626);
or OR3 (N1649, N1646, N1079, N913);
nand NAND3 (N1650, N1641, N382, N1091);
or OR4 (N1651, N1643, N779, N555, N940);
buf BUF1 (N1652, N1644);
or OR4 (N1653, N1647, N520, N956, N870);
xor XOR2 (N1654, N1620, N178);
xor XOR2 (N1655, N1645, N650);
nand NAND4 (N1656, N1639, N29, N84, N1215);
or OR3 (N1657, N1656, N1154, N1454);
not NOT1 (N1658, N1653);
buf BUF1 (N1659, N1654);
buf BUF1 (N1660, N1659);
or OR4 (N1661, N1652, N923, N499, N961);
or OR3 (N1662, N1660, N575, N1555);
buf BUF1 (N1663, N1648);
xor XOR2 (N1664, N1657, N429);
nor NOR2 (N1665, N1632, N223);
nand NAND2 (N1666, N1658, N679);
nand NAND3 (N1667, N1661, N343, N1195);
buf BUF1 (N1668, N1662);
and AND2 (N1669, N1655, N174);
xor XOR2 (N1670, N1668, N443);
not NOT1 (N1671, N1651);
or OR4 (N1672, N1665, N1002, N193, N305);
nand NAND4 (N1673, N1672, N1652, N357, N964);
nor NOR3 (N1674, N1671, N31, N113);
nand NAND4 (N1675, N1650, N154, N20, N148);
not NOT1 (N1676, N1670);
and AND4 (N1677, N1666, N536, N727, N1551);
buf BUF1 (N1678, N1649);
buf BUF1 (N1679, N1673);
xor XOR2 (N1680, N1677, N1197);
buf BUF1 (N1681, N1678);
not NOT1 (N1682, N1675);
and AND3 (N1683, N1663, N49, N776);
buf BUF1 (N1684, N1683);
and AND2 (N1685, N1684, N688);
buf BUF1 (N1686, N1682);
xor XOR2 (N1687, N1676, N32);
nand NAND4 (N1688, N1680, N377, N1398, N1200);
and AND3 (N1689, N1679, N1246, N1110);
not NOT1 (N1690, N1688);
and AND3 (N1691, N1685, N1347, N314);
nand NAND3 (N1692, N1674, N1554, N1488);
and AND4 (N1693, N1687, N1400, N37, N1067);
buf BUF1 (N1694, N1667);
nand NAND3 (N1695, N1694, N629, N1527);
or OR4 (N1696, N1686, N1233, N857, N1371);
or OR4 (N1697, N1692, N627, N571, N1696);
and AND4 (N1698, N1432, N906, N254, N283);
nand NAND2 (N1699, N1691, N896);
nor NOR2 (N1700, N1690, N570);
or OR2 (N1701, N1700, N1692);
xor XOR2 (N1702, N1664, N1048);
buf BUF1 (N1703, N1681);
or OR2 (N1704, N1699, N1638);
nor NOR3 (N1705, N1702, N300, N654);
not NOT1 (N1706, N1705);
buf BUF1 (N1707, N1703);
nor NOR4 (N1708, N1697, N576, N865, N1095);
buf BUF1 (N1709, N1701);
and AND3 (N1710, N1698, N798, N121);
or OR2 (N1711, N1669, N1696);
nor NOR2 (N1712, N1689, N53);
and AND4 (N1713, N1710, N841, N1337, N317);
and AND2 (N1714, N1693, N637);
not NOT1 (N1715, N1714);
nand NAND4 (N1716, N1712, N1704, N615, N362);
nand NAND2 (N1717, N1395, N1671);
xor XOR2 (N1718, N1706, N1169);
not NOT1 (N1719, N1716);
not NOT1 (N1720, N1713);
buf BUF1 (N1721, N1718);
and AND2 (N1722, N1719, N379);
nand NAND4 (N1723, N1695, N1631, N1059, N371);
nand NAND4 (N1724, N1717, N1549, N1004, N393);
and AND4 (N1725, N1709, N988, N850, N1681);
nor NOR4 (N1726, N1711, N1327, N6, N108);
nand NAND3 (N1727, N1726, N1078, N1027);
not NOT1 (N1728, N1725);
not NOT1 (N1729, N1720);
or OR3 (N1730, N1728, N1219, N894);
nor NOR2 (N1731, N1722, N741);
and AND4 (N1732, N1715, N623, N241, N247);
buf BUF1 (N1733, N1724);
not NOT1 (N1734, N1732);
buf BUF1 (N1735, N1723);
not NOT1 (N1736, N1708);
nor NOR3 (N1737, N1735, N725, N308);
nand NAND4 (N1738, N1731, N1266, N183, N206);
buf BUF1 (N1739, N1730);
nor NOR3 (N1740, N1736, N853, N1700);
xor XOR2 (N1741, N1733, N494);
nand NAND3 (N1742, N1741, N1524, N1019);
or OR3 (N1743, N1738, N24, N993);
or OR3 (N1744, N1737, N416, N63);
nor NOR4 (N1745, N1729, N118, N1338, N593);
nand NAND2 (N1746, N1707, N1192);
buf BUF1 (N1747, N1727);
or OR4 (N1748, N1739, N836, N42, N466);
nand NAND3 (N1749, N1740, N769, N87);
or OR4 (N1750, N1742, N68, N1534, N1615);
or OR3 (N1751, N1746, N938, N138);
xor XOR2 (N1752, N1734, N18);
or OR4 (N1753, N1752, N234, N303, N603);
nand NAND3 (N1754, N1748, N1746, N1125);
nor NOR3 (N1755, N1745, N1015, N1712);
or OR3 (N1756, N1751, N122, N906);
not NOT1 (N1757, N1755);
and AND3 (N1758, N1756, N532, N403);
nor NOR2 (N1759, N1749, N4);
buf BUF1 (N1760, N1754);
and AND4 (N1761, N1721, N1298, N926, N1519);
nor NOR4 (N1762, N1753, N1627, N1715, N228);
or OR4 (N1763, N1747, N1293, N1615, N744);
and AND2 (N1764, N1750, N565);
not NOT1 (N1765, N1743);
buf BUF1 (N1766, N1757);
not NOT1 (N1767, N1764);
not NOT1 (N1768, N1765);
nand NAND2 (N1769, N1759, N963);
nor NOR3 (N1770, N1758, N1193, N999);
xor XOR2 (N1771, N1766, N1536);
and AND4 (N1772, N1760, N1160, N1652, N876);
buf BUF1 (N1773, N1769);
nor NOR2 (N1774, N1768, N812);
or OR4 (N1775, N1770, N1744, N561, N1128);
buf BUF1 (N1776, N1668);
nor NOR4 (N1777, N1774, N862, N838, N1064);
xor XOR2 (N1778, N1761, N1656);
and AND3 (N1779, N1776, N287, N987);
or OR2 (N1780, N1767, N419);
and AND2 (N1781, N1778, N1728);
not NOT1 (N1782, N1775);
nor NOR3 (N1783, N1780, N701, N997);
not NOT1 (N1784, N1771);
nand NAND2 (N1785, N1784, N181);
or OR3 (N1786, N1779, N1716, N1367);
buf BUF1 (N1787, N1777);
nor NOR2 (N1788, N1785, N184);
buf BUF1 (N1789, N1781);
nand NAND4 (N1790, N1762, N1580, N1237, N1392);
nor NOR4 (N1791, N1773, N995, N1005, N1657);
or OR2 (N1792, N1786, N288);
xor XOR2 (N1793, N1790, N528);
not NOT1 (N1794, N1782);
nand NAND2 (N1795, N1792, N1066);
not NOT1 (N1796, N1787);
nand NAND3 (N1797, N1772, N365, N972);
buf BUF1 (N1798, N1783);
or OR4 (N1799, N1791, N1169, N328, N1502);
and AND2 (N1800, N1763, N1113);
and AND3 (N1801, N1798, N49, N550);
not NOT1 (N1802, N1789);
buf BUF1 (N1803, N1794);
nand NAND2 (N1804, N1797, N164);
nor NOR2 (N1805, N1795, N1711);
buf BUF1 (N1806, N1800);
xor XOR2 (N1807, N1801, N1288);
xor XOR2 (N1808, N1799, N758);
not NOT1 (N1809, N1806);
and AND4 (N1810, N1796, N515, N1765, N1229);
not NOT1 (N1811, N1803);
and AND2 (N1812, N1807, N1545);
nor NOR2 (N1813, N1788, N404);
not NOT1 (N1814, N1811);
nor NOR3 (N1815, N1802, N1090, N1720);
and AND3 (N1816, N1808, N1726, N600);
xor XOR2 (N1817, N1812, N939);
buf BUF1 (N1818, N1815);
or OR4 (N1819, N1793, N424, N1560, N1361);
or OR3 (N1820, N1813, N82, N1064);
not NOT1 (N1821, N1814);
buf BUF1 (N1822, N1817);
not NOT1 (N1823, N1804);
nor NOR2 (N1824, N1809, N541);
buf BUF1 (N1825, N1818);
or OR2 (N1826, N1824, N942);
not NOT1 (N1827, N1819);
buf BUF1 (N1828, N1823);
buf BUF1 (N1829, N1810);
nand NAND2 (N1830, N1828, N1128);
buf BUF1 (N1831, N1829);
nor NOR4 (N1832, N1831, N1515, N1769, N1193);
or OR2 (N1833, N1822, N165);
nand NAND2 (N1834, N1805, N1004);
nor NOR2 (N1835, N1825, N1011);
not NOT1 (N1836, N1833);
xor XOR2 (N1837, N1827, N1123);
nor NOR3 (N1838, N1820, N1371, N746);
not NOT1 (N1839, N1838);
nand NAND2 (N1840, N1816, N1080);
xor XOR2 (N1841, N1839, N992);
nor NOR4 (N1842, N1834, N1077, N1029, N283);
buf BUF1 (N1843, N1842);
nor NOR4 (N1844, N1843, N1692, N442, N1331);
or OR4 (N1845, N1837, N274, N49, N1725);
or OR4 (N1846, N1845, N1617, N1341, N1440);
nor NOR3 (N1847, N1836, N1263, N1727);
or OR4 (N1848, N1830, N444, N1025, N826);
xor XOR2 (N1849, N1832, N1417);
and AND2 (N1850, N1847, N1421);
or OR2 (N1851, N1821, N17);
buf BUF1 (N1852, N1844);
not NOT1 (N1853, N1852);
xor XOR2 (N1854, N1849, N1694);
and AND4 (N1855, N1840, N1624, N198, N771);
nor NOR4 (N1856, N1826, N1663, N1449, N1790);
xor XOR2 (N1857, N1848, N620);
nand NAND4 (N1858, N1854, N1432, N1002, N1441);
nor NOR4 (N1859, N1856, N1540, N353, N37);
nand NAND2 (N1860, N1846, N1342);
not NOT1 (N1861, N1850);
nor NOR4 (N1862, N1859, N810, N45, N711);
or OR4 (N1863, N1862, N1797, N339, N1816);
not NOT1 (N1864, N1835);
nor NOR4 (N1865, N1857, N636, N1035, N838);
buf BUF1 (N1866, N1853);
or OR2 (N1867, N1866, N92);
xor XOR2 (N1868, N1861, N1572);
or OR4 (N1869, N1851, N131, N1727, N1673);
buf BUF1 (N1870, N1864);
not NOT1 (N1871, N1863);
nor NOR2 (N1872, N1855, N1336);
not NOT1 (N1873, N1841);
not NOT1 (N1874, N1871);
not NOT1 (N1875, N1867);
buf BUF1 (N1876, N1870);
nor NOR3 (N1877, N1873, N233, N1594);
and AND3 (N1878, N1869, N783, N1503);
buf BUF1 (N1879, N1877);
nand NAND4 (N1880, N1865, N324, N610, N1472);
buf BUF1 (N1881, N1868);
not NOT1 (N1882, N1860);
xor XOR2 (N1883, N1878, N1773);
xor XOR2 (N1884, N1876, N296);
nand NAND4 (N1885, N1875, N19, N15, N1177);
nand NAND2 (N1886, N1874, N1847);
nand NAND3 (N1887, N1858, N1102, N1381);
and AND3 (N1888, N1872, N232, N1420);
not NOT1 (N1889, N1885);
buf BUF1 (N1890, N1879);
not NOT1 (N1891, N1883);
nand NAND2 (N1892, N1884, N657);
buf BUF1 (N1893, N1880);
nand NAND2 (N1894, N1890, N393);
not NOT1 (N1895, N1881);
nor NOR3 (N1896, N1886, N804, N1658);
or OR3 (N1897, N1891, N1671, N1808);
and AND2 (N1898, N1889, N918);
buf BUF1 (N1899, N1887);
not NOT1 (N1900, N1892);
xor XOR2 (N1901, N1898, N1578);
buf BUF1 (N1902, N1896);
or OR2 (N1903, N1888, N475);
not NOT1 (N1904, N1902);
or OR4 (N1905, N1900, N342, N362, N737);
nor NOR4 (N1906, N1882, N400, N1464, N1408);
nor NOR4 (N1907, N1897, N1103, N1722, N271);
buf BUF1 (N1908, N1903);
nand NAND2 (N1909, N1894, N27);
or OR4 (N1910, N1908, N120, N1274, N852);
and AND3 (N1911, N1910, N737, N640);
and AND3 (N1912, N1901, N1444, N1047);
not NOT1 (N1913, N1893);
xor XOR2 (N1914, N1904, N1532);
or OR4 (N1915, N1914, N1906, N1526, N564);
or OR2 (N1916, N550, N1759);
or OR2 (N1917, N1912, N101);
nor NOR3 (N1918, N1899, N1548, N351);
nor NOR4 (N1919, N1916, N1463, N465, N1001);
xor XOR2 (N1920, N1895, N1750);
not NOT1 (N1921, N1911);
xor XOR2 (N1922, N1913, N1719);
nand NAND4 (N1923, N1921, N1526, N1639, N1291);
nand NAND2 (N1924, N1907, N660);
nand NAND2 (N1925, N1917, N1739);
nand NAND3 (N1926, N1925, N109, N1137);
not NOT1 (N1927, N1922);
xor XOR2 (N1928, N1924, N367);
not NOT1 (N1929, N1920);
or OR4 (N1930, N1928, N1460, N781, N1741);
nand NAND3 (N1931, N1918, N812, N1089);
nand NAND4 (N1932, N1929, N1170, N87, N1723);
xor XOR2 (N1933, N1919, N1384);
not NOT1 (N1934, N1905);
not NOT1 (N1935, N1931);
nor NOR3 (N1936, N1932, N1856, N313);
not NOT1 (N1937, N1923);
buf BUF1 (N1938, N1930);
nand NAND2 (N1939, N1915, N960);
buf BUF1 (N1940, N1909);
buf BUF1 (N1941, N1926);
nand NAND3 (N1942, N1938, N1660, N11);
or OR2 (N1943, N1936, N381);
buf BUF1 (N1944, N1940);
nand NAND2 (N1945, N1933, N1799);
xor XOR2 (N1946, N1927, N1091);
not NOT1 (N1947, N1935);
xor XOR2 (N1948, N1947, N369);
not NOT1 (N1949, N1941);
and AND3 (N1950, N1942, N1028, N686);
xor XOR2 (N1951, N1950, N585);
buf BUF1 (N1952, N1951);
nor NOR2 (N1953, N1943, N903);
and AND3 (N1954, N1934, N946, N1938);
xor XOR2 (N1955, N1948, N87);
xor XOR2 (N1956, N1946, N356);
not NOT1 (N1957, N1953);
nand NAND4 (N1958, N1949, N1410, N993, N1059);
buf BUF1 (N1959, N1957);
xor XOR2 (N1960, N1952, N23);
nor NOR2 (N1961, N1944, N1778);
nand NAND4 (N1962, N1959, N95, N51, N1638);
or OR3 (N1963, N1939, N428, N336);
xor XOR2 (N1964, N1954, N344);
nor NOR3 (N1965, N1961, N487, N1486);
xor XOR2 (N1966, N1963, N699);
buf BUF1 (N1967, N1945);
xor XOR2 (N1968, N1964, N704);
not NOT1 (N1969, N1955);
buf BUF1 (N1970, N1968);
xor XOR2 (N1971, N1965, N1926);
and AND4 (N1972, N1956, N427, N955, N1601);
nand NAND4 (N1973, N1937, N897, N307, N1404);
nand NAND4 (N1974, N1971, N533, N1314, N1932);
and AND3 (N1975, N1960, N601, N1323);
xor XOR2 (N1976, N1973, N496);
nor NOR3 (N1977, N1969, N1781, N1751);
buf BUF1 (N1978, N1958);
nor NOR2 (N1979, N1962, N1228);
or OR4 (N1980, N1972, N382, N581, N754);
and AND4 (N1981, N1976, N433, N398, N1927);
or OR3 (N1982, N1977, N1617, N1726);
nor NOR4 (N1983, N1974, N1294, N104, N617);
nor NOR4 (N1984, N1975, N523, N55, N1133);
buf BUF1 (N1985, N1984);
and AND2 (N1986, N1979, N317);
and AND2 (N1987, N1980, N1550);
or OR3 (N1988, N1981, N759, N867);
not NOT1 (N1989, N1983);
and AND3 (N1990, N1978, N538, N1076);
nor NOR3 (N1991, N1986, N1916, N1833);
xor XOR2 (N1992, N1990, N1083);
nor NOR3 (N1993, N1989, N696, N600);
nand NAND4 (N1994, N1982, N1489, N523, N51);
not NOT1 (N1995, N1988);
and AND4 (N1996, N1987, N176, N14, N962);
nor NOR2 (N1997, N1991, N1156);
not NOT1 (N1998, N1995);
nor NOR4 (N1999, N1994, N735, N1042, N1683);
xor XOR2 (N2000, N1967, N1154);
or OR2 (N2001, N1985, N117);
not NOT1 (N2002, N1966);
xor XOR2 (N2003, N1993, N1918);
nor NOR2 (N2004, N2002, N630);
buf BUF1 (N2005, N2000);
nor NOR4 (N2006, N2005, N458, N1279, N821);
nand NAND4 (N2007, N2004, N448, N431, N1420);
not NOT1 (N2008, N2007);
buf BUF1 (N2009, N2008);
not NOT1 (N2010, N2003);
nor NOR4 (N2011, N2006, N285, N501, N26);
and AND2 (N2012, N1970, N1379);
xor XOR2 (N2013, N2011, N887);
buf BUF1 (N2014, N2001);
or OR4 (N2015, N1998, N743, N1793, N1439);
nand NAND2 (N2016, N1996, N1273);
and AND2 (N2017, N2013, N1607);
nor NOR4 (N2018, N1997, N811, N387, N1906);
and AND4 (N2019, N2017, N1384, N1457, N24);
xor XOR2 (N2020, N2019, N1474);
buf BUF1 (N2021, N2015);
and AND2 (N2022, N1992, N757);
buf BUF1 (N2023, N2018);
and AND4 (N2024, N2023, N764, N80, N1016);
buf BUF1 (N2025, N2012);
nor NOR4 (N2026, N2020, N1766, N1970, N1375);
xor XOR2 (N2027, N2022, N935);
nor NOR2 (N2028, N2009, N1951);
or OR2 (N2029, N2024, N1532);
nor NOR2 (N2030, N2029, N1565);
or OR2 (N2031, N2016, N1619);
nor NOR4 (N2032, N2021, N1753, N199, N1474);
nand NAND4 (N2033, N2031, N276, N512, N1384);
or OR2 (N2034, N2030, N1957);
and AND2 (N2035, N2033, N740);
nor NOR4 (N2036, N2010, N1845, N662, N915);
buf BUF1 (N2037, N2027);
not NOT1 (N2038, N1999);
or OR2 (N2039, N2038, N448);
nand NAND4 (N2040, N2035, N1547, N1097, N1587);
or OR4 (N2041, N2039, N1661, N1635, N755);
not NOT1 (N2042, N2014);
and AND3 (N2043, N2041, N1090, N356);
buf BUF1 (N2044, N2026);
xor XOR2 (N2045, N2034, N127);
not NOT1 (N2046, N2028);
or OR3 (N2047, N2037, N1297, N1159);
xor XOR2 (N2048, N2025, N1584);
buf BUF1 (N2049, N2045);
nand NAND2 (N2050, N2040, N606);
nand NAND4 (N2051, N2044, N1447, N166, N711);
buf BUF1 (N2052, N2048);
and AND3 (N2053, N2032, N372, N1857);
nor NOR4 (N2054, N2053, N1725, N1382, N65);
nor NOR4 (N2055, N2046, N353, N1545, N1959);
and AND4 (N2056, N2036, N1013, N942, N1769);
not NOT1 (N2057, N2056);
or OR4 (N2058, N2051, N1651, N817, N1824);
or OR4 (N2059, N2042, N304, N1274, N338);
xor XOR2 (N2060, N2057, N895);
nor NOR3 (N2061, N2054, N579, N740);
nor NOR4 (N2062, N2052, N1608, N1710, N910);
buf BUF1 (N2063, N2043);
not NOT1 (N2064, N2059);
not NOT1 (N2065, N2063);
or OR2 (N2066, N2060, N1585);
and AND2 (N2067, N2065, N568);
nand NAND4 (N2068, N2067, N361, N1248, N241);
not NOT1 (N2069, N2068);
or OR2 (N2070, N2047, N1399);
and AND3 (N2071, N2055, N255, N226);
not NOT1 (N2072, N2070);
or OR4 (N2073, N2072, N1351, N1478, N1658);
buf BUF1 (N2074, N2062);
nor NOR3 (N2075, N2066, N1492, N424);
nor NOR2 (N2076, N2069, N1695);
nand NAND3 (N2077, N2049, N1045, N540);
buf BUF1 (N2078, N2061);
buf BUF1 (N2079, N2076);
nor NOR2 (N2080, N2078, N499);
and AND2 (N2081, N2073, N952);
or OR2 (N2082, N2075, N798);
xor XOR2 (N2083, N2081, N1865);
nand NAND2 (N2084, N2071, N1274);
nand NAND4 (N2085, N2079, N1122, N1826, N912);
not NOT1 (N2086, N2085);
buf BUF1 (N2087, N2058);
nor NOR4 (N2088, N2087, N670, N1304, N874);
nand NAND2 (N2089, N2080, N1245);
nor NOR4 (N2090, N2083, N190, N1423, N1774);
nor NOR2 (N2091, N2082, N1507);
buf BUF1 (N2092, N2077);
nor NOR2 (N2093, N2090, N1145);
nand NAND3 (N2094, N2093, N1814, N148);
not NOT1 (N2095, N2050);
buf BUF1 (N2096, N2091);
nor NOR3 (N2097, N2089, N64, N1572);
xor XOR2 (N2098, N2086, N645);
not NOT1 (N2099, N2098);
xor XOR2 (N2100, N2084, N2098);
buf BUF1 (N2101, N2095);
xor XOR2 (N2102, N2099, N54);
xor XOR2 (N2103, N2064, N1126);
not NOT1 (N2104, N2088);
nand NAND3 (N2105, N2101, N895, N933);
nand NAND2 (N2106, N2100, N915);
buf BUF1 (N2107, N2104);
xor XOR2 (N2108, N2096, N2005);
nand NAND3 (N2109, N2105, N1485, N1401);
buf BUF1 (N2110, N2074);
xor XOR2 (N2111, N2092, N1231);
nand NAND2 (N2112, N2106, N1082);
buf BUF1 (N2113, N2107);
not NOT1 (N2114, N2108);
not NOT1 (N2115, N2109);
nor NOR3 (N2116, N2112, N605, N1493);
or OR4 (N2117, N2097, N436, N1054, N178);
and AND4 (N2118, N2116, N224, N611, N1161);
xor XOR2 (N2119, N2113, N1383);
nand NAND3 (N2120, N2114, N585, N1558);
buf BUF1 (N2121, N2102);
and AND2 (N2122, N2103, N78);
xor XOR2 (N2123, N2115, N1022);
buf BUF1 (N2124, N2111);
or OR4 (N2125, N2110, N725, N334, N880);
buf BUF1 (N2126, N2124);
xor XOR2 (N2127, N2123, N59);
and AND4 (N2128, N2122, N1790, N1203, N411);
and AND3 (N2129, N2125, N1306, N997);
nand NAND3 (N2130, N2094, N769, N824);
not NOT1 (N2131, N2126);
buf BUF1 (N2132, N2131);
not NOT1 (N2133, N2129);
and AND4 (N2134, N2127, N1676, N643, N18);
xor XOR2 (N2135, N2117, N2118);
or OR2 (N2136, N871, N2111);
buf BUF1 (N2137, N2133);
buf BUF1 (N2138, N2134);
or OR2 (N2139, N2120, N357);
nand NAND2 (N2140, N2136, N1472);
nand NAND4 (N2141, N2128, N1441, N21, N2116);
nor NOR4 (N2142, N2130, N148, N2129, N937);
not NOT1 (N2143, N2121);
not NOT1 (N2144, N2142);
or OR3 (N2145, N2138, N1759, N1342);
nor NOR2 (N2146, N2141, N335);
or OR2 (N2147, N2132, N1911);
nor NOR4 (N2148, N2135, N759, N459, N1339);
and AND2 (N2149, N2147, N240);
buf BUF1 (N2150, N2143);
not NOT1 (N2151, N2140);
and AND2 (N2152, N2139, N1173);
not NOT1 (N2153, N2144);
nor NOR2 (N2154, N2148, N1854);
and AND4 (N2155, N2150, N1629, N1556, N148);
buf BUF1 (N2156, N2154);
and AND4 (N2157, N2146, N1369, N1642, N1799);
not NOT1 (N2158, N2156);
buf BUF1 (N2159, N2151);
not NOT1 (N2160, N2153);
not NOT1 (N2161, N2137);
and AND4 (N2162, N2152, N363, N2127, N605);
or OR4 (N2163, N2145, N170, N1190, N847);
or OR2 (N2164, N2159, N2058);
xor XOR2 (N2165, N2119, N1330);
and AND4 (N2166, N2155, N48, N1700, N1832);
nor NOR4 (N2167, N2162, N1098, N794, N1359);
buf BUF1 (N2168, N2157);
nand NAND4 (N2169, N2161, N841, N1342, N2135);
or OR4 (N2170, N2164, N723, N1824, N1901);
buf BUF1 (N2171, N2158);
buf BUF1 (N2172, N2149);
nand NAND4 (N2173, N2160, N828, N533, N933);
nand NAND3 (N2174, N2170, N2049, N1740);
nor NOR2 (N2175, N2166, N619);
or OR2 (N2176, N2171, N1218);
nand NAND3 (N2177, N2174, N1427, N2032);
or OR3 (N2178, N2167, N1614, N658);
buf BUF1 (N2179, N2169);
nor NOR3 (N2180, N2177, N820, N1972);
nor NOR3 (N2181, N2163, N338, N2027);
nand NAND3 (N2182, N2168, N746, N1964);
buf BUF1 (N2183, N2180);
xor XOR2 (N2184, N2178, N675);
nand NAND4 (N2185, N2183, N785, N640, N424);
or OR2 (N2186, N2176, N333);
and AND4 (N2187, N2173, N330, N1235, N1847);
and AND2 (N2188, N2186, N87);
nor NOR4 (N2189, N2172, N1366, N2079, N2101);
xor XOR2 (N2190, N2188, N1642);
nor NOR3 (N2191, N2182, N1592, N1909);
nand NAND3 (N2192, N2187, N1794, N712);
or OR3 (N2193, N2165, N1235, N152);
nor NOR4 (N2194, N2189, N1746, N84, N328);
and AND2 (N2195, N2179, N1715);
or OR3 (N2196, N2190, N747, N1475);
nand NAND4 (N2197, N2185, N66, N1821, N1736);
and AND3 (N2198, N2194, N499, N1273);
buf BUF1 (N2199, N2181);
not NOT1 (N2200, N2191);
or OR2 (N2201, N2195, N1498);
buf BUF1 (N2202, N2198);
or OR3 (N2203, N2175, N946, N1950);
and AND4 (N2204, N2197, N1047, N2193, N846);
xor XOR2 (N2205, N1250, N324);
nand NAND2 (N2206, N2199, N467);
or OR4 (N2207, N2204, N1429, N408, N1377);
nor NOR3 (N2208, N2202, N1411, N1683);
buf BUF1 (N2209, N2206);
and AND4 (N2210, N2200, N1704, N1910, N673);
nor NOR4 (N2211, N2201, N280, N2139, N1563);
and AND4 (N2212, N2211, N12, N1061, N1765);
xor XOR2 (N2213, N2184, N1306);
not NOT1 (N2214, N2207);
nand NAND3 (N2215, N2205, N1910, N91);
nand NAND3 (N2216, N2210, N973, N1855);
nand NAND4 (N2217, N2215, N269, N883, N70);
nor NOR3 (N2218, N2214, N422, N1554);
and AND3 (N2219, N2203, N872, N1846);
or OR2 (N2220, N2209, N547);
buf BUF1 (N2221, N2219);
xor XOR2 (N2222, N2208, N2035);
not NOT1 (N2223, N2213);
xor XOR2 (N2224, N2222, N1065);
xor XOR2 (N2225, N2196, N478);
or OR2 (N2226, N2212, N1859);
or OR2 (N2227, N2216, N96);
nor NOR3 (N2228, N2224, N1867, N1419);
nand NAND2 (N2229, N2225, N491);
xor XOR2 (N2230, N2192, N756);
buf BUF1 (N2231, N2226);
nand NAND3 (N2232, N2230, N582, N1157);
not NOT1 (N2233, N2218);
not NOT1 (N2234, N2233);
buf BUF1 (N2235, N2223);
buf BUF1 (N2236, N2229);
xor XOR2 (N2237, N2232, N1905);
and AND4 (N2238, N2227, N1001, N830, N1916);
nor NOR3 (N2239, N2234, N1662, N278);
or OR3 (N2240, N2228, N68, N2053);
xor XOR2 (N2241, N2239, N2089);
nand NAND2 (N2242, N2231, N746);
nor NOR2 (N2243, N2242, N1312);
nor NOR3 (N2244, N2243, N2196, N2127);
buf BUF1 (N2245, N2235);
nor NOR4 (N2246, N2238, N1130, N732, N1998);
nand NAND3 (N2247, N2246, N610, N1107);
buf BUF1 (N2248, N2221);
not NOT1 (N2249, N2248);
nand NAND4 (N2250, N2240, N1709, N828, N557);
nand NAND2 (N2251, N2236, N2229);
nand NAND3 (N2252, N2244, N1719, N133);
nor NOR4 (N2253, N2241, N1123, N840, N705);
buf BUF1 (N2254, N2220);
nand NAND4 (N2255, N2250, N1216, N2154, N594);
xor XOR2 (N2256, N2247, N1058);
nand NAND3 (N2257, N2252, N1014, N1123);
xor XOR2 (N2258, N2245, N1776);
nor NOR2 (N2259, N2217, N1682);
nor NOR4 (N2260, N2257, N1043, N1857, N828);
xor XOR2 (N2261, N2259, N2201);
or OR4 (N2262, N2254, N587, N1337, N2109);
nor NOR4 (N2263, N2255, N1873, N461, N1848);
nand NAND2 (N2264, N2263, N1053);
buf BUF1 (N2265, N2251);
and AND3 (N2266, N2262, N2063, N1134);
not NOT1 (N2267, N2264);
not NOT1 (N2268, N2260);
nor NOR4 (N2269, N2256, N395, N1556, N2134);
nand NAND3 (N2270, N2237, N1486, N1695);
xor XOR2 (N2271, N2267, N684);
buf BUF1 (N2272, N2261);
nand NAND2 (N2273, N2253, N1726);
and AND4 (N2274, N2271, N92, N1832, N1740);
nand NAND2 (N2275, N2266, N7);
buf BUF1 (N2276, N2273);
xor XOR2 (N2277, N2268, N1782);
or OR3 (N2278, N2270, N1056, N1724);
or OR4 (N2279, N2276, N931, N123, N869);
xor XOR2 (N2280, N2269, N921);
buf BUF1 (N2281, N2272);
not NOT1 (N2282, N2265);
or OR4 (N2283, N2282, N342, N1645, N869);
buf BUF1 (N2284, N2249);
buf BUF1 (N2285, N2279);
and AND2 (N2286, N2277, N555);
and AND2 (N2287, N2281, N2039);
and AND4 (N2288, N2283, N261, N408, N2073);
and AND4 (N2289, N2275, N2275, N2026, N754);
buf BUF1 (N2290, N2274);
xor XOR2 (N2291, N2288, N1926);
or OR2 (N2292, N2278, N1709);
nor NOR3 (N2293, N2291, N857, N835);
not NOT1 (N2294, N2290);
not NOT1 (N2295, N2258);
not NOT1 (N2296, N2285);
buf BUF1 (N2297, N2280);
and AND3 (N2298, N2292, N758, N1870);
nor NOR4 (N2299, N2297, N1412, N1001, N1201);
not NOT1 (N2300, N2293);
buf BUF1 (N2301, N2294);
nand NAND3 (N2302, N2296, N1147, N1411);
not NOT1 (N2303, N2289);
xor XOR2 (N2304, N2286, N175);
xor XOR2 (N2305, N2301, N1049);
and AND4 (N2306, N2298, N1100, N56, N1880);
and AND3 (N2307, N2299, N1653, N1324);
buf BUF1 (N2308, N2304);
nand NAND4 (N2309, N2308, N408, N1422, N1083);
xor XOR2 (N2310, N2302, N1205);
nand NAND2 (N2311, N2300, N2172);
xor XOR2 (N2312, N2303, N630);
nand NAND3 (N2313, N2295, N825, N776);
not NOT1 (N2314, N2310);
buf BUF1 (N2315, N2312);
nor NOR2 (N2316, N2306, N1661);
and AND4 (N2317, N2309, N2187, N1938, N1587);
nand NAND4 (N2318, N2313, N1375, N505, N861);
buf BUF1 (N2319, N2287);
nand NAND2 (N2320, N2318, N680);
nor NOR3 (N2321, N2319, N109, N1911);
nand NAND3 (N2322, N2316, N2137, N953);
or OR2 (N2323, N2311, N1036);
xor XOR2 (N2324, N2307, N121);
not NOT1 (N2325, N2305);
xor XOR2 (N2326, N2317, N321);
or OR4 (N2327, N2325, N1165, N1070, N581);
or OR4 (N2328, N2314, N942, N941, N578);
nor NOR3 (N2329, N2326, N1706, N1454);
nor NOR3 (N2330, N2321, N1810, N942);
or OR2 (N2331, N2330, N879);
xor XOR2 (N2332, N2284, N1288);
not NOT1 (N2333, N2323);
and AND2 (N2334, N2328, N997);
not NOT1 (N2335, N2327);
nand NAND3 (N2336, N2324, N1663, N838);
buf BUF1 (N2337, N2333);
not NOT1 (N2338, N2334);
nand NAND4 (N2339, N2331, N1787, N696, N1839);
or OR4 (N2340, N2339, N1181, N1476, N961);
buf BUF1 (N2341, N2315);
and AND4 (N2342, N2320, N763, N1757, N2050);
buf BUF1 (N2343, N2338);
buf BUF1 (N2344, N2341);
nor NOR3 (N2345, N2343, N1443, N633);
and AND2 (N2346, N2322, N2069);
buf BUF1 (N2347, N2345);
nor NOR4 (N2348, N2337, N662, N2271, N1049);
not NOT1 (N2349, N2342);
xor XOR2 (N2350, N2336, N307);
or OR4 (N2351, N2329, N1090, N2214, N1560);
or OR2 (N2352, N2349, N1283);
or OR4 (N2353, N2346, N113, N612, N1228);
not NOT1 (N2354, N2348);
or OR2 (N2355, N2347, N2159);
not NOT1 (N2356, N2350);
buf BUF1 (N2357, N2340);
or OR2 (N2358, N2351, N1689);
not NOT1 (N2359, N2354);
or OR3 (N2360, N2352, N1023, N1610);
and AND3 (N2361, N2359, N168, N1938);
nand NAND4 (N2362, N2344, N514, N765, N1442);
nand NAND4 (N2363, N2361, N1240, N21, N1579);
not NOT1 (N2364, N2332);
nor NOR2 (N2365, N2358, N2235);
not NOT1 (N2366, N2364);
not NOT1 (N2367, N2365);
nor NOR3 (N2368, N2335, N575, N141);
buf BUF1 (N2369, N2362);
nor NOR4 (N2370, N2353, N1711, N1191, N779);
xor XOR2 (N2371, N2357, N619);
not NOT1 (N2372, N2355);
and AND2 (N2373, N2369, N821);
buf BUF1 (N2374, N2372);
or OR2 (N2375, N2368, N2281);
xor XOR2 (N2376, N2370, N2331);
not NOT1 (N2377, N2366);
or OR4 (N2378, N2363, N71, N880, N730);
nand NAND2 (N2379, N2374, N195);
nand NAND3 (N2380, N2378, N1382, N1343);
nand NAND2 (N2381, N2376, N1551);
xor XOR2 (N2382, N2371, N282);
and AND4 (N2383, N2356, N244, N2090, N1213);
nand NAND2 (N2384, N2373, N683);
nand NAND2 (N2385, N2382, N1083);
xor XOR2 (N2386, N2380, N17);
or OR2 (N2387, N2385, N2030);
nand NAND4 (N2388, N2367, N1722, N355, N1956);
or OR4 (N2389, N2379, N1940, N2027, N1496);
xor XOR2 (N2390, N2386, N2298);
or OR4 (N2391, N2383, N1938, N1402, N2043);
nor NOR2 (N2392, N2375, N770);
nand NAND3 (N2393, N2388, N1323, N419);
or OR2 (N2394, N2387, N1539);
nor NOR3 (N2395, N2392, N1298, N2371);
and AND3 (N2396, N2390, N356, N284);
or OR4 (N2397, N2395, N43, N1859, N1365);
not NOT1 (N2398, N2396);
nor NOR2 (N2399, N2389, N536);
nand NAND2 (N2400, N2399, N1195);
not NOT1 (N2401, N2400);
buf BUF1 (N2402, N2398);
xor XOR2 (N2403, N2401, N1681);
or OR4 (N2404, N2377, N2086, N853, N1988);
and AND4 (N2405, N2394, N1482, N487, N264);
or OR3 (N2406, N2402, N866, N1037);
nand NAND4 (N2407, N2384, N735, N1160, N1288);
not NOT1 (N2408, N2403);
and AND2 (N2409, N2404, N6);
nand NAND2 (N2410, N2393, N789);
nand NAND2 (N2411, N2391, N1688);
xor XOR2 (N2412, N2381, N1563);
or OR4 (N2413, N2405, N1200, N1075, N1820);
and AND4 (N2414, N2411, N190, N1817, N387);
nand NAND4 (N2415, N2409, N1236, N1663, N329);
not NOT1 (N2416, N2397);
or OR3 (N2417, N2413, N2249, N1924);
buf BUF1 (N2418, N2414);
and AND3 (N2419, N2418, N1387, N1395);
and AND4 (N2420, N2415, N1410, N194, N2382);
nand NAND4 (N2421, N2408, N93, N1371, N508);
nand NAND3 (N2422, N2412, N636, N918);
xor XOR2 (N2423, N2421, N174);
nand NAND4 (N2424, N2422, N2038, N375, N2234);
not NOT1 (N2425, N2417);
nor NOR2 (N2426, N2423, N1690);
nand NAND3 (N2427, N2406, N622, N2000);
and AND2 (N2428, N2425, N1257);
buf BUF1 (N2429, N2426);
nand NAND2 (N2430, N2428, N330);
nor NOR3 (N2431, N2419, N1362, N1407);
or OR3 (N2432, N2407, N1149, N1299);
not NOT1 (N2433, N2431);
buf BUF1 (N2434, N2430);
nand NAND2 (N2435, N2433, N2258);
and AND2 (N2436, N2427, N1200);
and AND3 (N2437, N2424, N2055, N1591);
nand NAND2 (N2438, N2436, N2179);
or OR2 (N2439, N2429, N1469);
nor NOR4 (N2440, N2432, N42, N265, N347);
or OR3 (N2441, N2440, N766, N1998);
nor NOR2 (N2442, N2439, N1565);
and AND3 (N2443, N2441, N1883, N2052);
or OR3 (N2444, N2442, N184, N190);
xor XOR2 (N2445, N2444, N731);
or OR4 (N2446, N2445, N1557, N1244, N2183);
and AND4 (N2447, N2435, N1068, N546, N1066);
or OR3 (N2448, N2437, N507, N1907);
nand NAND4 (N2449, N2360, N1265, N1263, N1817);
not NOT1 (N2450, N2448);
not NOT1 (N2451, N2443);
nor NOR2 (N2452, N2434, N1755);
xor XOR2 (N2453, N2410, N917);
nor NOR3 (N2454, N2420, N2451, N1352);
or OR2 (N2455, N643, N1744);
and AND3 (N2456, N2455, N776, N1173);
not NOT1 (N2457, N2450);
xor XOR2 (N2458, N2456, N2219);
nor NOR2 (N2459, N2452, N276);
nor NOR2 (N2460, N2449, N402);
buf BUF1 (N2461, N2416);
not NOT1 (N2462, N2446);
buf BUF1 (N2463, N2462);
buf BUF1 (N2464, N2454);
not NOT1 (N2465, N2464);
not NOT1 (N2466, N2465);
nand NAND2 (N2467, N2460, N232);
xor XOR2 (N2468, N2447, N915);
nand NAND2 (N2469, N2467, N1503);
xor XOR2 (N2470, N2469, N1471);
not NOT1 (N2471, N2470);
not NOT1 (N2472, N2463);
nor NOR2 (N2473, N2457, N1185);
or OR4 (N2474, N2466, N521, N1622, N1234);
not NOT1 (N2475, N2468);
nand NAND3 (N2476, N2453, N1437, N1173);
or OR4 (N2477, N2461, N34, N257, N1160);
nor NOR4 (N2478, N2438, N1663, N205, N1924);
not NOT1 (N2479, N2458);
nor NOR4 (N2480, N2474, N850, N777, N2004);
and AND4 (N2481, N2473, N1673, N2388, N534);
xor XOR2 (N2482, N2479, N1742);
xor XOR2 (N2483, N2475, N658);
or OR2 (N2484, N2482, N121);
buf BUF1 (N2485, N2472);
or OR3 (N2486, N2480, N1122, N2049);
nor NOR2 (N2487, N2471, N2374);
nor NOR2 (N2488, N2477, N445);
not NOT1 (N2489, N2478);
nor NOR3 (N2490, N2485, N293, N1226);
xor XOR2 (N2491, N2476, N2395);
not NOT1 (N2492, N2483);
nor NOR4 (N2493, N2487, N1563, N658, N501);
nand NAND4 (N2494, N2484, N1832, N2041, N480);
not NOT1 (N2495, N2459);
or OR3 (N2496, N2489, N479, N1871);
nor NOR2 (N2497, N2490, N556);
not NOT1 (N2498, N2481);
and AND2 (N2499, N2493, N485);
nand NAND3 (N2500, N2494, N821, N1536);
nand NAND2 (N2501, N2488, N2350);
or OR4 (N2502, N2486, N777, N1778, N1499);
or OR2 (N2503, N2496, N1556);
nor NOR2 (N2504, N2501, N2307);
and AND3 (N2505, N2495, N1183, N1424);
nor NOR2 (N2506, N2502, N2491);
nand NAND4 (N2507, N1094, N1333, N1632, N1073);
or OR2 (N2508, N2499, N520);
xor XOR2 (N2509, N2492, N635);
xor XOR2 (N2510, N2497, N507);
and AND2 (N2511, N2509, N1879);
nor NOR2 (N2512, N2503, N970);
nand NAND3 (N2513, N2508, N1532, N1957);
nand NAND3 (N2514, N2507, N1914, N2194);
xor XOR2 (N2515, N2506, N637);
xor XOR2 (N2516, N2498, N788);
and AND3 (N2517, N2514, N1955, N1466);
xor XOR2 (N2518, N2504, N368);
and AND3 (N2519, N2510, N1653, N1024);
buf BUF1 (N2520, N2515);
not NOT1 (N2521, N2517);
buf BUF1 (N2522, N2500);
or OR2 (N2523, N2511, N94);
nor NOR4 (N2524, N2518, N2011, N1335, N2138);
or OR4 (N2525, N2523, N107, N2045, N900);
or OR2 (N2526, N2519, N2181);
nand NAND4 (N2527, N2516, N565, N179, N2251);
buf BUF1 (N2528, N2521);
or OR3 (N2529, N2520, N1086, N1030);
not NOT1 (N2530, N2529);
not NOT1 (N2531, N2525);
buf BUF1 (N2532, N2530);
nand NAND2 (N2533, N2524, N251);
nor NOR3 (N2534, N2513, N1859, N312);
not NOT1 (N2535, N2533);
nor NOR3 (N2536, N2512, N520, N1376);
not NOT1 (N2537, N2527);
or OR2 (N2538, N2505, N1970);
and AND4 (N2539, N2538, N147, N1962, N2097);
and AND3 (N2540, N2532, N1170, N1203);
or OR4 (N2541, N2528, N40, N1834, N2203);
and AND4 (N2542, N2535, N2222, N1311, N1883);
xor XOR2 (N2543, N2541, N266);
buf BUF1 (N2544, N2540);
buf BUF1 (N2545, N2534);
nand NAND3 (N2546, N2542, N1206, N759);
or OR2 (N2547, N2522, N2064);
buf BUF1 (N2548, N2536);
not NOT1 (N2549, N2547);
buf BUF1 (N2550, N2537);
or OR2 (N2551, N2546, N1608);
nand NAND2 (N2552, N2539, N1638);
xor XOR2 (N2553, N2544, N1843);
xor XOR2 (N2554, N2551, N225);
buf BUF1 (N2555, N2543);
buf BUF1 (N2556, N2552);
or OR4 (N2557, N2548, N1571, N1434, N312);
or OR4 (N2558, N2556, N2099, N1229, N526);
nand NAND3 (N2559, N2557, N1442, N1786);
and AND4 (N2560, N2554, N1001, N477, N545);
or OR2 (N2561, N2531, N353);
buf BUF1 (N2562, N2559);
nor NOR2 (N2563, N2558, N518);
not NOT1 (N2564, N2545);
and AND4 (N2565, N2526, N2085, N1226, N146);
or OR2 (N2566, N2565, N2091);
and AND2 (N2567, N2563, N1818);
not NOT1 (N2568, N2561);
nor NOR2 (N2569, N2568, N1971);
xor XOR2 (N2570, N2567, N603);
or OR4 (N2571, N2560, N1220, N127, N911);
or OR3 (N2572, N2564, N1871, N1403);
buf BUF1 (N2573, N2570);
xor XOR2 (N2574, N2569, N1955);
xor XOR2 (N2575, N2553, N422);
and AND2 (N2576, N2571, N536);
not NOT1 (N2577, N2562);
not NOT1 (N2578, N2575);
nand NAND2 (N2579, N2573, N328);
buf BUF1 (N2580, N2576);
nand NAND2 (N2581, N2549, N886);
and AND2 (N2582, N2566, N2492);
and AND4 (N2583, N2572, N1350, N1643, N867);
nor NOR2 (N2584, N2581, N37);
and AND4 (N2585, N2584, N675, N1286, N1804);
or OR3 (N2586, N2577, N1938, N2301);
and AND4 (N2587, N2555, N959, N1074, N470);
or OR2 (N2588, N2580, N1167);
not NOT1 (N2589, N2582);
and AND3 (N2590, N2585, N1535, N663);
nor NOR2 (N2591, N2579, N1752);
nor NOR2 (N2592, N2591, N1885);
not NOT1 (N2593, N2583);
buf BUF1 (N2594, N2587);
and AND3 (N2595, N2594, N458, N1508);
nand NAND2 (N2596, N2593, N381);
nor NOR2 (N2597, N2595, N168);
or OR4 (N2598, N2597, N1776, N2432, N795);
nand NAND2 (N2599, N2598, N2038);
nand NAND3 (N2600, N2589, N2536, N664);
xor XOR2 (N2601, N2588, N2120);
xor XOR2 (N2602, N2550, N472);
not NOT1 (N2603, N2586);
nand NAND4 (N2604, N2592, N1767, N1621, N2533);
and AND3 (N2605, N2600, N2304, N852);
nor NOR2 (N2606, N2578, N210);
nor NOR2 (N2607, N2590, N202);
buf BUF1 (N2608, N2574);
nor NOR3 (N2609, N2601, N1242, N1040);
and AND3 (N2610, N2604, N640, N1302);
or OR3 (N2611, N2603, N2546, N2422);
buf BUF1 (N2612, N2605);
xor XOR2 (N2613, N2599, N2051);
xor XOR2 (N2614, N2608, N1567);
nor NOR2 (N2615, N2614, N578);
or OR4 (N2616, N2611, N1105, N527, N1725);
not NOT1 (N2617, N2606);
and AND2 (N2618, N2615, N202);
nor NOR4 (N2619, N2616, N1893, N1175, N155);
nor NOR2 (N2620, N2609, N2214);
buf BUF1 (N2621, N2613);
not NOT1 (N2622, N2602);
nand NAND4 (N2623, N2621, N1716, N807, N2009);
and AND4 (N2624, N2596, N2509, N789, N1946);
or OR2 (N2625, N2619, N207);
nor NOR4 (N2626, N2607, N2011, N924, N1252);
buf BUF1 (N2627, N2625);
or OR4 (N2628, N2622, N2110, N1011, N1000);
not NOT1 (N2629, N2624);
and AND4 (N2630, N2617, N2253, N190, N1834);
not NOT1 (N2631, N2618);
or OR2 (N2632, N2623, N2187);
or OR2 (N2633, N2627, N352);
and AND3 (N2634, N2628, N415, N1793);
buf BUF1 (N2635, N2612);
and AND3 (N2636, N2634, N1408, N1123);
nand NAND4 (N2637, N2635, N1877, N1625, N2459);
and AND2 (N2638, N2620, N2164);
or OR2 (N2639, N2637, N2435);
nor NOR2 (N2640, N2629, N2478);
not NOT1 (N2641, N2632);
or OR3 (N2642, N2636, N1414, N1816);
nand NAND2 (N2643, N2640, N628);
nand NAND3 (N2644, N2642, N1262, N81);
nor NOR2 (N2645, N2626, N144);
or OR4 (N2646, N2630, N765, N307, N509);
xor XOR2 (N2647, N2610, N1948);
nor NOR4 (N2648, N2639, N19, N229, N80);
nor NOR4 (N2649, N2644, N952, N1901, N2274);
nand NAND4 (N2650, N2633, N1610, N1970, N32);
or OR3 (N2651, N2643, N129, N855);
or OR2 (N2652, N2651, N2145);
buf BUF1 (N2653, N2631);
and AND2 (N2654, N2641, N1478);
or OR2 (N2655, N2652, N358);
nor NOR3 (N2656, N2638, N814, N713);
or OR4 (N2657, N2649, N2042, N2469, N415);
or OR2 (N2658, N2655, N10);
and AND4 (N2659, N2645, N1617, N27, N993);
xor XOR2 (N2660, N2656, N14);
or OR4 (N2661, N2660, N830, N475, N687);
not NOT1 (N2662, N2653);
xor XOR2 (N2663, N2646, N927);
and AND3 (N2664, N2661, N368, N2363);
nor NOR4 (N2665, N2658, N497, N1153, N1750);
nand NAND2 (N2666, N2654, N2067);
and AND3 (N2667, N2659, N1421, N1528);
and AND4 (N2668, N2657, N703, N1834, N158);
and AND4 (N2669, N2668, N1106, N132, N921);
nor NOR4 (N2670, N2663, N1029, N2140, N782);
and AND3 (N2671, N2665, N2551, N61);
buf BUF1 (N2672, N2666);
and AND2 (N2673, N2671, N2060);
xor XOR2 (N2674, N2648, N2140);
buf BUF1 (N2675, N2647);
or OR3 (N2676, N2664, N1779, N1344);
not NOT1 (N2677, N2670);
and AND3 (N2678, N2673, N2248, N1338);
not NOT1 (N2679, N2675);
buf BUF1 (N2680, N2667);
not NOT1 (N2681, N2680);
nand NAND2 (N2682, N2677, N623);
or OR2 (N2683, N2669, N141);
and AND2 (N2684, N2678, N2572);
nor NOR2 (N2685, N2674, N1258);
not NOT1 (N2686, N2650);
buf BUF1 (N2687, N2672);
and AND3 (N2688, N2679, N1296, N2460);
xor XOR2 (N2689, N2662, N1806);
buf BUF1 (N2690, N2676);
nand NAND3 (N2691, N2689, N1435, N92);
or OR2 (N2692, N2685, N144);
and AND4 (N2693, N2692, N2528, N2377, N2691);
buf BUF1 (N2694, N1746);
nand NAND2 (N2695, N2693, N1571);
nand NAND3 (N2696, N2690, N485, N248);
and AND2 (N2697, N2688, N1825);
xor XOR2 (N2698, N2681, N2692);
nand NAND3 (N2699, N2698, N496, N1481);
xor XOR2 (N2700, N2683, N1653);
buf BUF1 (N2701, N2682);
buf BUF1 (N2702, N2684);
or OR2 (N2703, N2701, N482);
nor NOR2 (N2704, N2700, N952);
xor XOR2 (N2705, N2699, N1802);
xor XOR2 (N2706, N2704, N2506);
buf BUF1 (N2707, N2695);
buf BUF1 (N2708, N2687);
xor XOR2 (N2709, N2702, N212);
or OR2 (N2710, N2707, N1771);
and AND4 (N2711, N2694, N1645, N994, N62);
or OR2 (N2712, N2711, N1897);
or OR2 (N2713, N2709, N765);
xor XOR2 (N2714, N2712, N72);
nor NOR4 (N2715, N2703, N2603, N504, N1630);
or OR4 (N2716, N2715, N1282, N2083, N1150);
not NOT1 (N2717, N2708);
not NOT1 (N2718, N2713);
nand NAND3 (N2719, N2717, N2576, N883);
xor XOR2 (N2720, N2686, N1093);
not NOT1 (N2721, N2714);
and AND4 (N2722, N2716, N1003, N1201, N760);
and AND2 (N2723, N2710, N674);
nand NAND2 (N2724, N2718, N400);
and AND2 (N2725, N2720, N1594);
or OR3 (N2726, N2719, N445, N473);
buf BUF1 (N2727, N2697);
xor XOR2 (N2728, N2721, N2133);
and AND3 (N2729, N2724, N1047, N2044);
not NOT1 (N2730, N2728);
nand NAND2 (N2731, N2722, N2410);
buf BUF1 (N2732, N2726);
and AND3 (N2733, N2730, N428, N2566);
buf BUF1 (N2734, N2729);
nor NOR4 (N2735, N2731, N2651, N2396, N1943);
nand NAND2 (N2736, N2734, N2623);
xor XOR2 (N2737, N2696, N1938);
xor XOR2 (N2738, N2725, N2102);
nand NAND3 (N2739, N2705, N431, N1836);
buf BUF1 (N2740, N2706);
xor XOR2 (N2741, N2723, N493);
and AND3 (N2742, N2733, N1494, N1805);
or OR4 (N2743, N2738, N2063, N1100, N651);
buf BUF1 (N2744, N2739);
not NOT1 (N2745, N2737);
or OR2 (N2746, N2742, N1519);
nand NAND2 (N2747, N2736, N1455);
nor NOR4 (N2748, N2745, N2116, N1292, N1807);
xor XOR2 (N2749, N2748, N2106);
buf BUF1 (N2750, N2727);
nand NAND3 (N2751, N2744, N808, N660);
and AND3 (N2752, N2743, N963, N1425);
not NOT1 (N2753, N2749);
nor NOR2 (N2754, N2752, N230);
buf BUF1 (N2755, N2751);
or OR4 (N2756, N2750, N817, N2183, N1929);
xor XOR2 (N2757, N2732, N2491);
and AND2 (N2758, N2740, N2245);
nor NOR4 (N2759, N2746, N1595, N136, N1652);
buf BUF1 (N2760, N2757);
nor NOR3 (N2761, N2759, N2601, N2616);
nand NAND2 (N2762, N2761, N283);
not NOT1 (N2763, N2754);
nand NAND4 (N2764, N2760, N1577, N2651, N442);
nor NOR2 (N2765, N2756, N2608);
nor NOR3 (N2766, N2747, N2316, N2505);
nand NAND2 (N2767, N2741, N823);
nand NAND4 (N2768, N2766, N512, N1053, N2565);
not NOT1 (N2769, N2755);
nand NAND2 (N2770, N2767, N2133);
nor NOR3 (N2771, N2763, N1165, N127);
nand NAND4 (N2772, N2771, N1147, N1067, N2158);
nand NAND4 (N2773, N2758, N2391, N878, N1130);
xor XOR2 (N2774, N2770, N1);
buf BUF1 (N2775, N2774);
or OR3 (N2776, N2769, N2441, N704);
buf BUF1 (N2777, N2776);
or OR4 (N2778, N2765, N612, N2494, N1414);
xor XOR2 (N2779, N2772, N977);
xor XOR2 (N2780, N2753, N1161);
not NOT1 (N2781, N2775);
not NOT1 (N2782, N2778);
or OR3 (N2783, N2762, N792, N5);
buf BUF1 (N2784, N2735);
not NOT1 (N2785, N2764);
or OR2 (N2786, N2780, N259);
or OR3 (N2787, N2786, N2373, N2268);
and AND4 (N2788, N2784, N1433, N1139, N2313);
nand NAND3 (N2789, N2782, N2448, N2129);
nand NAND2 (N2790, N2785, N890);
or OR3 (N2791, N2783, N1224, N1688);
and AND3 (N2792, N2781, N1434, N1574);
or OR3 (N2793, N2788, N2499, N377);
and AND3 (N2794, N2790, N2340, N2330);
xor XOR2 (N2795, N2792, N1061);
xor XOR2 (N2796, N2795, N597);
nor NOR3 (N2797, N2791, N1294, N1351);
or OR2 (N2798, N2779, N1774);
buf BUF1 (N2799, N2787);
nand NAND4 (N2800, N2796, N1363, N998, N2387);
not NOT1 (N2801, N2789);
xor XOR2 (N2802, N2794, N725);
buf BUF1 (N2803, N2773);
or OR3 (N2804, N2801, N641, N2703);
or OR3 (N2805, N2798, N736, N335);
or OR4 (N2806, N2799, N370, N2192, N1894);
nor NOR2 (N2807, N2804, N1614);
nor NOR4 (N2808, N2797, N2528, N1910, N1617);
or OR3 (N2809, N2808, N1248, N148);
nor NOR4 (N2810, N2809, N2151, N102, N2414);
xor XOR2 (N2811, N2800, N1814);
not NOT1 (N2812, N2806);
nand NAND4 (N2813, N2807, N407, N395, N1444);
nand NAND2 (N2814, N2811, N2333);
nor NOR3 (N2815, N2777, N475, N1698);
buf BUF1 (N2816, N2814);
nand NAND2 (N2817, N2816, N2712);
not NOT1 (N2818, N2793);
nand NAND4 (N2819, N2812, N764, N2577, N547);
not NOT1 (N2820, N2815);
and AND2 (N2821, N2817, N1000);
xor XOR2 (N2822, N2813, N381);
or OR3 (N2823, N2818, N2576, N490);
buf BUF1 (N2824, N2821);
or OR4 (N2825, N2824, N2317, N105, N701);
nand NAND2 (N2826, N2819, N1936);
xor XOR2 (N2827, N2802, N76);
nand NAND2 (N2828, N2805, N624);
nor NOR2 (N2829, N2823, N1567);
and AND4 (N2830, N2810, N1493, N1187, N2296);
buf BUF1 (N2831, N2822);
nand NAND2 (N2832, N2826, N2553);
not NOT1 (N2833, N2831);
and AND4 (N2834, N2832, N1116, N1256, N1535);
or OR4 (N2835, N2833, N2809, N482, N144);
not NOT1 (N2836, N2830);
nand NAND2 (N2837, N2825, N1248);
xor XOR2 (N2838, N2828, N218);
or OR2 (N2839, N2836, N1835);
nand NAND3 (N2840, N2829, N1233, N518);
and AND4 (N2841, N2768, N1426, N1327, N1216);
buf BUF1 (N2842, N2837);
nor NOR2 (N2843, N2835, N342);
nor NOR3 (N2844, N2841, N1668, N2715);
not NOT1 (N2845, N2820);
not NOT1 (N2846, N2840);
buf BUF1 (N2847, N2839);
buf BUF1 (N2848, N2803);
and AND2 (N2849, N2838, N1776);
or OR4 (N2850, N2843, N915, N2352, N2756);
nor NOR3 (N2851, N2850, N1940, N2090);
buf BUF1 (N2852, N2842);
nor NOR3 (N2853, N2834, N807, N2817);
nor NOR2 (N2854, N2846, N1806);
not NOT1 (N2855, N2827);
and AND2 (N2856, N2855, N2434);
nor NOR4 (N2857, N2852, N138, N964, N1036);
xor XOR2 (N2858, N2853, N860);
xor XOR2 (N2859, N2845, N923);
or OR3 (N2860, N2857, N944, N2801);
not NOT1 (N2861, N2849);
nand NAND2 (N2862, N2859, N853);
and AND3 (N2863, N2851, N474, N1946);
nand NAND4 (N2864, N2854, N1621, N176, N2443);
and AND3 (N2865, N2860, N2818, N1658);
nor NOR3 (N2866, N2858, N1128, N696);
buf BUF1 (N2867, N2856);
xor XOR2 (N2868, N2864, N2100);
nand NAND3 (N2869, N2865, N413, N1719);
nor NOR2 (N2870, N2847, N1600);
buf BUF1 (N2871, N2861);
not NOT1 (N2872, N2871);
and AND2 (N2873, N2867, N825);
nand NAND3 (N2874, N2869, N895, N510);
nand NAND3 (N2875, N2872, N861, N848);
nand NAND2 (N2876, N2875, N2688);
nand NAND3 (N2877, N2848, N453, N1834);
not NOT1 (N2878, N2844);
xor XOR2 (N2879, N2868, N1462);
xor XOR2 (N2880, N2877, N860);
not NOT1 (N2881, N2876);
nor NOR4 (N2882, N2880, N1769, N2216, N2140);
or OR4 (N2883, N2879, N448, N2606, N1306);
not NOT1 (N2884, N2882);
not NOT1 (N2885, N2866);
not NOT1 (N2886, N2863);
or OR3 (N2887, N2881, N91, N2074);
nor NOR3 (N2888, N2874, N2580, N1197);
xor XOR2 (N2889, N2862, N843);
nor NOR2 (N2890, N2887, N153);
nor NOR3 (N2891, N2886, N976, N29);
xor XOR2 (N2892, N2891, N2563);
and AND3 (N2893, N2888, N2616, N69);
and AND4 (N2894, N2892, N140, N1549, N1987);
nor NOR3 (N2895, N2884, N2894, N2787);
and AND2 (N2896, N771, N2169);
nor NOR4 (N2897, N2873, N1180, N1363, N2700);
or OR3 (N2898, N2885, N2190, N316);
nand NAND3 (N2899, N2883, N1802, N1756);
or OR4 (N2900, N2889, N1296, N1895, N2122);
nor NOR4 (N2901, N2893, N470, N2039, N422);
buf BUF1 (N2902, N2890);
nand NAND3 (N2903, N2898, N317, N1981);
xor XOR2 (N2904, N2870, N2178);
or OR2 (N2905, N2901, N973);
or OR2 (N2906, N2904, N925);
or OR3 (N2907, N2897, N2523, N1305);
nor NOR3 (N2908, N2902, N2342, N81);
nor NOR4 (N2909, N2907, N1070, N2266, N1586);
nor NOR2 (N2910, N2905, N1605);
and AND4 (N2911, N2908, N2076, N1542, N2551);
xor XOR2 (N2912, N2911, N1802);
or OR4 (N2913, N2900, N831, N1630, N2151);
nand NAND2 (N2914, N2912, N1479);
xor XOR2 (N2915, N2878, N33);
not NOT1 (N2916, N2903);
not NOT1 (N2917, N2906);
or OR3 (N2918, N2910, N944, N1507);
nand NAND3 (N2919, N2918, N2243, N1013);
or OR2 (N2920, N2909, N2445);
buf BUF1 (N2921, N2920);
and AND4 (N2922, N2916, N813, N1554, N1200);
or OR4 (N2923, N2919, N2642, N1739, N2428);
xor XOR2 (N2924, N2914, N2796);
xor XOR2 (N2925, N2921, N1435);
xor XOR2 (N2926, N2913, N223);
nand NAND3 (N2927, N2895, N461, N829);
not NOT1 (N2928, N2923);
nor NOR2 (N2929, N2915, N2269);
not NOT1 (N2930, N2917);
nand NAND2 (N2931, N2927, N715);
or OR4 (N2932, N2925, N1135, N2268, N423);
nor NOR3 (N2933, N2928, N631, N101);
xor XOR2 (N2934, N2896, N1123);
not NOT1 (N2935, N2922);
and AND3 (N2936, N2934, N2761, N2802);
xor XOR2 (N2937, N2932, N633);
and AND3 (N2938, N2899, N1054, N633);
xor XOR2 (N2939, N2931, N2520);
not NOT1 (N2940, N2935);
not NOT1 (N2941, N2939);
and AND2 (N2942, N2926, N825);
xor XOR2 (N2943, N2933, N1958);
or OR2 (N2944, N2938, N2027);
nor NOR3 (N2945, N2943, N2510, N2221);
nor NOR2 (N2946, N2940, N2900);
buf BUF1 (N2947, N2945);
nand NAND3 (N2948, N2941, N1628, N1423);
nor NOR2 (N2949, N2937, N222);
nor NOR2 (N2950, N2949, N739);
and AND3 (N2951, N2924, N483, N2937);
and AND3 (N2952, N2936, N502, N140);
xor XOR2 (N2953, N2946, N1457);
buf BUF1 (N2954, N2952);
nand NAND3 (N2955, N2929, N2284, N702);
not NOT1 (N2956, N2951);
nand NAND3 (N2957, N2955, N618, N1452);
or OR4 (N2958, N2954, N1958, N285, N1752);
not NOT1 (N2959, N2950);
not NOT1 (N2960, N2948);
not NOT1 (N2961, N2959);
buf BUF1 (N2962, N2947);
nand NAND3 (N2963, N2953, N795, N2760);
buf BUF1 (N2964, N2962);
not NOT1 (N2965, N2960);
or OR4 (N2966, N2958, N874, N2039, N2889);
nor NOR3 (N2967, N2942, N2585, N2180);
nor NOR2 (N2968, N2957, N2451);
or OR2 (N2969, N2963, N2318);
nand NAND2 (N2970, N2967, N2799);
not NOT1 (N2971, N2970);
nor NOR4 (N2972, N2944, N1004, N1325, N2963);
or OR4 (N2973, N2969, N994, N1921, N2853);
nand NAND3 (N2974, N2956, N2615, N1181);
or OR4 (N2975, N2973, N767, N51, N2899);
nand NAND4 (N2976, N2974, N615, N512, N2437);
xor XOR2 (N2977, N2971, N2274);
not NOT1 (N2978, N2966);
xor XOR2 (N2979, N2976, N2467);
buf BUF1 (N2980, N2978);
not NOT1 (N2981, N2965);
or OR4 (N2982, N2979, N2502, N2470, N2528);
buf BUF1 (N2983, N2972);
xor XOR2 (N2984, N2977, N2641);
or OR3 (N2985, N2968, N496, N619);
not NOT1 (N2986, N2964);
and AND3 (N2987, N2975, N202, N372);
or OR2 (N2988, N2930, N784);
nand NAND2 (N2989, N2986, N2268);
not NOT1 (N2990, N2989);
nand NAND2 (N2991, N2982, N1864);
nand NAND3 (N2992, N2991, N5, N695);
nor NOR3 (N2993, N2988, N1594, N192);
and AND4 (N2994, N2983, N2606, N1222, N2392);
not NOT1 (N2995, N2984);
or OR4 (N2996, N2981, N1111, N246, N2604);
buf BUF1 (N2997, N2994);
nand NAND2 (N2998, N2997, N1836);
or OR3 (N2999, N2987, N1047, N491);
buf BUF1 (N3000, N2980);
xor XOR2 (N3001, N2996, N1393);
xor XOR2 (N3002, N3000, N726);
buf BUF1 (N3003, N2999);
buf BUF1 (N3004, N2992);
xor XOR2 (N3005, N2985, N1759);
xor XOR2 (N3006, N2995, N247);
or OR3 (N3007, N3006, N1472, N2118);
not NOT1 (N3008, N3007);
nand NAND2 (N3009, N3002, N136);
or OR2 (N3010, N2961, N1808);
buf BUF1 (N3011, N3001);
or OR3 (N3012, N3009, N1463, N2458);
nor NOR3 (N3013, N3005, N2795, N1840);
xor XOR2 (N3014, N3011, N1077);
nand NAND2 (N3015, N3008, N1343);
xor XOR2 (N3016, N2990, N942);
nand NAND2 (N3017, N3003, N1286);
xor XOR2 (N3018, N2993, N2306);
and AND2 (N3019, N3018, N2218);
and AND2 (N3020, N3013, N2342);
nand NAND2 (N3021, N3014, N242);
or OR4 (N3022, N3016, N207, N2958, N2312);
nand NAND2 (N3023, N3004, N1421);
and AND2 (N3024, N3012, N672);
buf BUF1 (N3025, N3019);
or OR2 (N3026, N3024, N51);
not NOT1 (N3027, N3010);
and AND4 (N3028, N3022, N1756, N2605, N2624);
nor NOR2 (N3029, N3017, N134);
and AND4 (N3030, N3029, N2260, N2506, N2190);
not NOT1 (N3031, N3015);
nand NAND2 (N3032, N2998, N510);
buf BUF1 (N3033, N3031);
buf BUF1 (N3034, N3026);
and AND4 (N3035, N3020, N516, N2990, N837);
and AND2 (N3036, N3035, N2359);
not NOT1 (N3037, N3023);
not NOT1 (N3038, N3036);
nor NOR3 (N3039, N3021, N323, N402);
xor XOR2 (N3040, N3037, N1412);
or OR2 (N3041, N3032, N3019);
xor XOR2 (N3042, N3027, N634);
xor XOR2 (N3043, N3042, N939);
nand NAND2 (N3044, N3043, N2932);
xor XOR2 (N3045, N3033, N1299);
nand NAND2 (N3046, N3028, N736);
or OR4 (N3047, N3025, N2942, N2416, N612);
and AND2 (N3048, N3041, N1395);
xor XOR2 (N3049, N3048, N878);
xor XOR2 (N3050, N3044, N2789);
nor NOR4 (N3051, N3045, N2418, N2565, N1985);
buf BUF1 (N3052, N3047);
nor NOR3 (N3053, N3051, N807, N2737);
xor XOR2 (N3054, N3053, N2401);
buf BUF1 (N3055, N3050);
and AND3 (N3056, N3046, N1624, N2429);
or OR3 (N3057, N3049, N2493, N2986);
xor XOR2 (N3058, N3056, N1268);
or OR4 (N3059, N3054, N1764, N408, N763);
nand NAND3 (N3060, N3038, N2218, N2940);
not NOT1 (N3061, N3055);
not NOT1 (N3062, N3058);
or OR2 (N3063, N3034, N2205);
buf BUF1 (N3064, N3060);
and AND4 (N3065, N3064, N238, N2158, N684);
not NOT1 (N3066, N3059);
nor NOR2 (N3067, N3040, N1408);
nand NAND3 (N3068, N3065, N1351, N490);
xor XOR2 (N3069, N3067, N636);
xor XOR2 (N3070, N3068, N2421);
xor XOR2 (N3071, N3057, N1538);
xor XOR2 (N3072, N3063, N81);
and AND4 (N3073, N3066, N804, N228, N2205);
and AND4 (N3074, N3061, N291, N334, N980);
or OR4 (N3075, N3062, N2072, N1203, N2421);
xor XOR2 (N3076, N3039, N1869);
not NOT1 (N3077, N3030);
or OR3 (N3078, N3071, N2753, N2545);
and AND4 (N3079, N3070, N513, N1079, N1234);
not NOT1 (N3080, N3077);
and AND2 (N3081, N3069, N2088);
and AND2 (N3082, N3080, N2912);
not NOT1 (N3083, N3082);
nand NAND3 (N3084, N3083, N1623, N485);
buf BUF1 (N3085, N3052);
nor NOR2 (N3086, N3076, N3015);
not NOT1 (N3087, N3079);
and AND3 (N3088, N3073, N2115, N418);
and AND3 (N3089, N3086, N1293, N3056);
nor NOR3 (N3090, N3078, N2765, N2894);
buf BUF1 (N3091, N3081);
buf BUF1 (N3092, N3087);
not NOT1 (N3093, N3092);
or OR3 (N3094, N3072, N640, N1449);
nand NAND4 (N3095, N3075, N1863, N1822, N2971);
or OR3 (N3096, N3084, N1149, N72);
buf BUF1 (N3097, N3088);
xor XOR2 (N3098, N3090, N2074);
nor NOR2 (N3099, N3094, N1773);
and AND4 (N3100, N3093, N3030, N2849, N1733);
not NOT1 (N3101, N3097);
not NOT1 (N3102, N3099);
buf BUF1 (N3103, N3100);
or OR3 (N3104, N3091, N2488, N46);
nor NOR2 (N3105, N3102, N722);
nor NOR2 (N3106, N3105, N588);
and AND2 (N3107, N3074, N3096);
buf BUF1 (N3108, N2462);
nand NAND2 (N3109, N3106, N2695);
nor NOR4 (N3110, N3101, N2883, N1999, N1377);
xor XOR2 (N3111, N3085, N905);
xor XOR2 (N3112, N3107, N184);
nor NOR3 (N3113, N3110, N2312, N2960);
xor XOR2 (N3114, N3113, N1497);
nand NAND2 (N3115, N3089, N1114);
xor XOR2 (N3116, N3103, N2510);
or OR2 (N3117, N3111, N165);
nand NAND3 (N3118, N3114, N1931, N993);
not NOT1 (N3119, N3112);
or OR2 (N3120, N3098, N650);
and AND2 (N3121, N3095, N680);
not NOT1 (N3122, N3118);
or OR3 (N3123, N3117, N3054, N249);
nand NAND3 (N3124, N3115, N1936, N255);
buf BUF1 (N3125, N3104);
nand NAND2 (N3126, N3121, N163);
nor NOR4 (N3127, N3125, N822, N890, N181);
xor XOR2 (N3128, N3124, N2654);
xor XOR2 (N3129, N3127, N411);
nor NOR4 (N3130, N3109, N774, N3118, N1317);
nor NOR3 (N3131, N3119, N880, N676);
buf BUF1 (N3132, N3130);
or OR2 (N3133, N3126, N1963);
buf BUF1 (N3134, N3123);
or OR4 (N3135, N3108, N1037, N1706, N1492);
and AND4 (N3136, N3134, N1567, N1076, N999);
or OR4 (N3137, N3131, N1272, N1721, N390);
nor NOR2 (N3138, N3135, N2239);
or OR3 (N3139, N3122, N638, N2078);
buf BUF1 (N3140, N3137);
xor XOR2 (N3141, N3116, N1911);
nand NAND3 (N3142, N3129, N1173, N940);
buf BUF1 (N3143, N3120);
not NOT1 (N3144, N3136);
nand NAND3 (N3145, N3140, N2991, N1529);
and AND3 (N3146, N3133, N338, N1451);
xor XOR2 (N3147, N3128, N1515);
buf BUF1 (N3148, N3147);
not NOT1 (N3149, N3146);
buf BUF1 (N3150, N3149);
or OR3 (N3151, N3148, N498, N2292);
or OR4 (N3152, N3142, N1060, N2679, N1118);
not NOT1 (N3153, N3144);
buf BUF1 (N3154, N3151);
or OR4 (N3155, N3138, N496, N730, N1279);
or OR2 (N3156, N3145, N2624);
xor XOR2 (N3157, N3153, N601);
and AND4 (N3158, N3157, N1290, N64, N3101);
or OR3 (N3159, N3141, N2429, N2325);
xor XOR2 (N3160, N3154, N3077);
nand NAND4 (N3161, N3156, N2248, N1248, N252);
xor XOR2 (N3162, N3158, N2153);
buf BUF1 (N3163, N3161);
buf BUF1 (N3164, N3139);
xor XOR2 (N3165, N3150, N501);
xor XOR2 (N3166, N3143, N1433);
or OR2 (N3167, N3132, N2342);
nand NAND4 (N3168, N3162, N1906, N1608, N802);
or OR4 (N3169, N3163, N1356, N2693, N2699);
nor NOR3 (N3170, N3155, N27, N2626);
or OR2 (N3171, N3152, N1673);
buf BUF1 (N3172, N3165);
nand NAND3 (N3173, N3160, N1842, N1340);
buf BUF1 (N3174, N3169);
nor NOR2 (N3175, N3167, N212);
not NOT1 (N3176, N3174);
not NOT1 (N3177, N3170);
xor XOR2 (N3178, N3164, N530);
nand NAND2 (N3179, N3176, N465);
buf BUF1 (N3180, N3159);
or OR3 (N3181, N3168, N1620, N2143);
xor XOR2 (N3182, N3177, N2589);
xor XOR2 (N3183, N3180, N2946);
nor NOR4 (N3184, N3178, N2985, N1501, N290);
or OR4 (N3185, N3181, N76, N2689, N87);
nor NOR4 (N3186, N3183, N647, N11, N248);
xor XOR2 (N3187, N3175, N3163);
nor NOR3 (N3188, N3185, N2752, N2538);
xor XOR2 (N3189, N3173, N2165);
buf BUF1 (N3190, N3172);
xor XOR2 (N3191, N3171, N323);
buf BUF1 (N3192, N3179);
nor NOR4 (N3193, N3191, N1524, N1406, N1404);
buf BUF1 (N3194, N3182);
and AND4 (N3195, N3188, N245, N950, N2810);
or OR2 (N3196, N3189, N1748);
buf BUF1 (N3197, N3193);
buf BUF1 (N3198, N3166);
buf BUF1 (N3199, N3195);
nor NOR2 (N3200, N3192, N1541);
xor XOR2 (N3201, N3199, N1482);
not NOT1 (N3202, N3184);
not NOT1 (N3203, N3200);
nand NAND3 (N3204, N3203, N182, N431);
xor XOR2 (N3205, N3187, N1462);
not NOT1 (N3206, N3205);
nand NAND3 (N3207, N3204, N988, N2176);
or OR4 (N3208, N3197, N379, N1997, N20);
nor NOR3 (N3209, N3190, N1465, N364);
buf BUF1 (N3210, N3194);
xor XOR2 (N3211, N3209, N391);
nand NAND4 (N3212, N3206, N299, N2725, N1372);
nand NAND3 (N3213, N3212, N2568, N2807);
nor NOR4 (N3214, N3196, N4, N3100, N1643);
not NOT1 (N3215, N3201);
not NOT1 (N3216, N3207);
not NOT1 (N3217, N3210);
nand NAND2 (N3218, N3213, N2346);
or OR2 (N3219, N3217, N2807);
xor XOR2 (N3220, N3215, N2748);
nand NAND3 (N3221, N3214, N207, N2814);
or OR4 (N3222, N3211, N2391, N1193, N2031);
buf BUF1 (N3223, N3198);
xor XOR2 (N3224, N3222, N2101);
and AND3 (N3225, N3220, N451, N792);
and AND3 (N3226, N3186, N758, N1267);
not NOT1 (N3227, N3225);
or OR4 (N3228, N3219, N1320, N1603, N1501);
and AND3 (N3229, N3216, N270, N1046);
nor NOR2 (N3230, N3221, N1612);
not NOT1 (N3231, N3229);
nor NOR4 (N3232, N3228, N2150, N435, N2802);
or OR4 (N3233, N3202, N744, N1006, N367);
not NOT1 (N3234, N3218);
nand NAND3 (N3235, N3227, N576, N2472);
nor NOR2 (N3236, N3230, N512);
xor XOR2 (N3237, N3233, N1936);
nor NOR4 (N3238, N3226, N644, N1310, N2482);
and AND4 (N3239, N3234, N2793, N1004, N1443);
not NOT1 (N3240, N3237);
or OR4 (N3241, N3239, N3145, N1287, N378);
buf BUF1 (N3242, N3241);
xor XOR2 (N3243, N3223, N1412);
xor XOR2 (N3244, N3238, N2691);
nand NAND3 (N3245, N3243, N387, N935);
and AND4 (N3246, N3232, N1516, N635, N2636);
nand NAND3 (N3247, N3244, N2361, N1720);
or OR3 (N3248, N3240, N2894, N272);
and AND2 (N3249, N3247, N2198);
buf BUF1 (N3250, N3208);
xor XOR2 (N3251, N3224, N2654);
nand NAND3 (N3252, N3242, N1773, N1058);
nand NAND2 (N3253, N3246, N253);
and AND4 (N3254, N3248, N1611, N2465, N184);
nor NOR3 (N3255, N3253, N1595, N2407);
nand NAND3 (N3256, N3250, N1177, N1082);
not NOT1 (N3257, N3254);
nor NOR2 (N3258, N3257, N2660);
or OR3 (N3259, N3249, N1451, N1719);
buf BUF1 (N3260, N3258);
nor NOR3 (N3261, N3235, N1978, N1304);
nand NAND3 (N3262, N3236, N3206, N2291);
buf BUF1 (N3263, N3255);
or OR3 (N3264, N3261, N1397, N2820);
nand NAND4 (N3265, N3260, N964, N2108, N1470);
xor XOR2 (N3266, N3251, N1606);
and AND3 (N3267, N3266, N832, N3208);
and AND4 (N3268, N3259, N241, N1703, N2058);
xor XOR2 (N3269, N3231, N1046);
nand NAND2 (N3270, N3265, N1251);
not NOT1 (N3271, N3264);
and AND4 (N3272, N3269, N1471, N2961, N3045);
nor NOR3 (N3273, N3270, N1488, N1216);
xor XOR2 (N3274, N3271, N1673);
and AND3 (N3275, N3252, N1065, N1463);
nor NOR4 (N3276, N3272, N1499, N1765, N2860);
and AND2 (N3277, N3268, N1224);
nand NAND4 (N3278, N3256, N1161, N1059, N533);
xor XOR2 (N3279, N3245, N288);
not NOT1 (N3280, N3273);
nor NOR4 (N3281, N3274, N798, N974, N318);
and AND4 (N3282, N3263, N212, N1760, N2979);
nor NOR2 (N3283, N3262, N2027);
and AND3 (N3284, N3275, N1972, N1736);
and AND4 (N3285, N3276, N1211, N2229, N2453);
or OR3 (N3286, N3267, N1729, N1352);
not NOT1 (N3287, N3286);
buf BUF1 (N3288, N3280);
and AND4 (N3289, N3288, N1973, N423, N253);
and AND2 (N3290, N3277, N1301);
nor NOR2 (N3291, N3282, N1683);
not NOT1 (N3292, N3279);
xor XOR2 (N3293, N3284, N2263);
not NOT1 (N3294, N3287);
not NOT1 (N3295, N3283);
not NOT1 (N3296, N3295);
nand NAND4 (N3297, N3289, N2688, N2882, N1461);
xor XOR2 (N3298, N3293, N1049);
not NOT1 (N3299, N3291);
nand NAND2 (N3300, N3299, N1796);
nor NOR3 (N3301, N3281, N2978, N1355);
xor XOR2 (N3302, N3296, N1616);
not NOT1 (N3303, N3292);
not NOT1 (N3304, N3300);
or OR3 (N3305, N3285, N2716, N1419);
nand NAND3 (N3306, N3303, N1964, N2384);
xor XOR2 (N3307, N3302, N2376);
xor XOR2 (N3308, N3298, N223);
nor NOR2 (N3309, N3290, N2087);
and AND3 (N3310, N3305, N2675, N3121);
xor XOR2 (N3311, N3307, N1788);
buf BUF1 (N3312, N3297);
and AND3 (N3313, N3301, N656, N157);
not NOT1 (N3314, N3311);
and AND3 (N3315, N3306, N2282, N811);
or OR2 (N3316, N3304, N1270);
not NOT1 (N3317, N3312);
or OR3 (N3318, N3313, N2613, N1308);
and AND2 (N3319, N3278, N1402);
nand NAND2 (N3320, N3309, N1536);
xor XOR2 (N3321, N3317, N2741);
xor XOR2 (N3322, N3320, N2230);
and AND4 (N3323, N3315, N605, N1193, N963);
xor XOR2 (N3324, N3294, N2537);
and AND2 (N3325, N3308, N947);
and AND2 (N3326, N3321, N354);
nand NAND2 (N3327, N3318, N1254);
or OR3 (N3328, N3325, N2890, N2360);
not NOT1 (N3329, N3323);
xor XOR2 (N3330, N3324, N729);
nor NOR4 (N3331, N3310, N3048, N2996, N2930);
buf BUF1 (N3332, N3322);
buf BUF1 (N3333, N3331);
not NOT1 (N3334, N3319);
not NOT1 (N3335, N3334);
xor XOR2 (N3336, N3330, N1040);
not NOT1 (N3337, N3326);
nand NAND4 (N3338, N3329, N3149, N974, N129);
or OR4 (N3339, N3336, N2477, N2433, N3275);
and AND2 (N3340, N3335, N1456);
xor XOR2 (N3341, N3339, N2567);
nor NOR3 (N3342, N3340, N2869, N966);
and AND3 (N3343, N3327, N3026, N3328);
buf BUF1 (N3344, N2137);
and AND4 (N3345, N3342, N2873, N2379, N1797);
or OR2 (N3346, N3337, N2474);
nor NOR4 (N3347, N3338, N2166, N1151, N924);
not NOT1 (N3348, N3343);
or OR3 (N3349, N3333, N482, N239);
nor NOR4 (N3350, N3344, N99, N2531, N821);
not NOT1 (N3351, N3316);
and AND3 (N3352, N3347, N2684, N2972);
and AND4 (N3353, N3346, N1681, N1316, N691);
xor XOR2 (N3354, N3351, N2341);
and AND2 (N3355, N3352, N1005);
nand NAND2 (N3356, N3354, N2425);
nand NAND3 (N3357, N3341, N3293, N238);
and AND4 (N3358, N3355, N2408, N2372, N544);
buf BUF1 (N3359, N3353);
not NOT1 (N3360, N3356);
nor NOR2 (N3361, N3345, N1428);
not NOT1 (N3362, N3360);
buf BUF1 (N3363, N3357);
or OR2 (N3364, N3359, N252);
nand NAND2 (N3365, N3349, N1877);
or OR2 (N3366, N3362, N2305);
and AND2 (N3367, N3365, N2721);
nor NOR4 (N3368, N3366, N2578, N1516, N3062);
xor XOR2 (N3369, N3332, N869);
nand NAND4 (N3370, N3358, N614, N1207, N235);
nor NOR4 (N3371, N3348, N534, N1519, N1559);
and AND2 (N3372, N3364, N523);
not NOT1 (N3373, N3363);
not NOT1 (N3374, N3373);
not NOT1 (N3375, N3350);
or OR4 (N3376, N3370, N2309, N715, N2118);
not NOT1 (N3377, N3361);
xor XOR2 (N3378, N3375, N46);
nand NAND4 (N3379, N3314, N587, N2856, N1742);
xor XOR2 (N3380, N3372, N1682);
nor NOR4 (N3381, N3377, N3000, N647, N2782);
not NOT1 (N3382, N3380);
buf BUF1 (N3383, N3367);
buf BUF1 (N3384, N3378);
and AND3 (N3385, N3369, N1640, N1871);
nand NAND3 (N3386, N3374, N341, N2064);
and AND2 (N3387, N3382, N1845);
nor NOR4 (N3388, N3386, N651, N1636, N541);
or OR3 (N3389, N3379, N2925, N151);
xor XOR2 (N3390, N3384, N1368);
xor XOR2 (N3391, N3381, N231);
buf BUF1 (N3392, N3388);
buf BUF1 (N3393, N3368);
nor NOR3 (N3394, N3389, N1922, N976);
nor NOR4 (N3395, N3371, N1775, N1866, N2749);
xor XOR2 (N3396, N3392, N1456);
not NOT1 (N3397, N3387);
xor XOR2 (N3398, N3385, N1147);
nand NAND3 (N3399, N3376, N2564, N659);
and AND3 (N3400, N3393, N1988, N2730);
nor NOR2 (N3401, N3394, N1849);
not NOT1 (N3402, N3396);
buf BUF1 (N3403, N3399);
or OR3 (N3404, N3397, N1579, N2786);
or OR3 (N3405, N3403, N1125, N3035);
xor XOR2 (N3406, N3402, N1639);
and AND2 (N3407, N3383, N1717);
not NOT1 (N3408, N3404);
or OR4 (N3409, N3406, N1762, N1249, N2307);
and AND3 (N3410, N3391, N1166, N3143);
and AND3 (N3411, N3390, N140, N794);
and AND2 (N3412, N3398, N870);
not NOT1 (N3413, N3401);
buf BUF1 (N3414, N3408);
buf BUF1 (N3415, N3405);
nor NOR2 (N3416, N3395, N220);
not NOT1 (N3417, N3413);
xor XOR2 (N3418, N3400, N2267);
and AND3 (N3419, N3410, N1310, N2570);
not NOT1 (N3420, N3414);
not NOT1 (N3421, N3419);
or OR4 (N3422, N3420, N2077, N2119, N1556);
buf BUF1 (N3423, N3418);
xor XOR2 (N3424, N3409, N2028);
nand NAND4 (N3425, N3422, N2602, N437, N515);
not NOT1 (N3426, N3417);
buf BUF1 (N3427, N3416);
and AND2 (N3428, N3423, N936);
nand NAND4 (N3429, N3407, N1907, N2905, N1017);
or OR4 (N3430, N3425, N449, N157, N2422);
not NOT1 (N3431, N3412);
not NOT1 (N3432, N3430);
nor NOR2 (N3433, N3411, N3113);
and AND2 (N3434, N3427, N2672);
nor NOR2 (N3435, N3434, N1681);
nor NOR2 (N3436, N3415, N777);
not NOT1 (N3437, N3426);
nor NOR3 (N3438, N3431, N3101, N821);
or OR3 (N3439, N3432, N2145, N3241);
buf BUF1 (N3440, N3433);
nor NOR2 (N3441, N3440, N2593);
and AND2 (N3442, N3436, N2019);
nand NAND2 (N3443, N3428, N2002);
xor XOR2 (N3444, N3435, N1838);
nand NAND4 (N3445, N3444, N180, N2966, N1032);
xor XOR2 (N3446, N3445, N815);
nand NAND4 (N3447, N3421, N2240, N3215, N2497);
or OR3 (N3448, N3439, N474, N858);
xor XOR2 (N3449, N3446, N1902);
xor XOR2 (N3450, N3437, N2927);
not NOT1 (N3451, N3442);
nor NOR2 (N3452, N3438, N227);
not NOT1 (N3453, N3441);
or OR4 (N3454, N3443, N1437, N3020, N196);
nand NAND2 (N3455, N3448, N341);
nand NAND2 (N3456, N3454, N2810);
buf BUF1 (N3457, N3451);
and AND3 (N3458, N3453, N2295, N2517);
not NOT1 (N3459, N3449);
or OR4 (N3460, N3456, N3278, N1717, N495);
xor XOR2 (N3461, N3447, N2198);
not NOT1 (N3462, N3461);
nand NAND4 (N3463, N3458, N621, N2359, N290);
nand NAND4 (N3464, N3459, N951, N2872, N130);
and AND3 (N3465, N3464, N1292, N2254);
not NOT1 (N3466, N3460);
and AND3 (N3467, N3455, N2768, N1089);
nor NOR3 (N3468, N3450, N716, N2546);
and AND3 (N3469, N3467, N208, N3366);
nand NAND2 (N3470, N3429, N3289);
or OR2 (N3471, N3469, N891);
or OR4 (N3472, N3463, N1388, N2176, N2476);
and AND4 (N3473, N3466, N1712, N763, N1194);
buf BUF1 (N3474, N3471);
buf BUF1 (N3475, N3468);
nor NOR2 (N3476, N3465, N1162);
not NOT1 (N3477, N3457);
or OR4 (N3478, N3475, N570, N1325, N481);
nand NAND2 (N3479, N3472, N2275);
buf BUF1 (N3480, N3470);
and AND3 (N3481, N3479, N270, N733);
nor NOR4 (N3482, N3462, N293, N3024, N308);
xor XOR2 (N3483, N3480, N1960);
xor XOR2 (N3484, N3477, N1224);
xor XOR2 (N3485, N3481, N897);
or OR4 (N3486, N3478, N180, N3088, N2370);
not NOT1 (N3487, N3424);
or OR4 (N3488, N3487, N63, N2816, N66);
xor XOR2 (N3489, N3474, N3242);
nor NOR4 (N3490, N3452, N2734, N2740, N1240);
nor NOR4 (N3491, N3488, N1587, N3119, N2828);
nand NAND3 (N3492, N3486, N1454, N659);
nor NOR2 (N3493, N3473, N2192);
buf BUF1 (N3494, N3492);
not NOT1 (N3495, N3493);
xor XOR2 (N3496, N3485, N2747);
and AND3 (N3497, N3490, N1997, N1632);
xor XOR2 (N3498, N3496, N240);
buf BUF1 (N3499, N3498);
nor NOR4 (N3500, N3484, N229, N622, N1300);
buf BUF1 (N3501, N3497);
nand NAND2 (N3502, N3494, N2062);
xor XOR2 (N3503, N3495, N2768);
not NOT1 (N3504, N3489);
and AND4 (N3505, N3503, N1294, N2344, N2611);
nand NAND2 (N3506, N3483, N487);
xor XOR2 (N3507, N3501, N2073);
buf BUF1 (N3508, N3504);
nand NAND2 (N3509, N3491, N2209);
not NOT1 (N3510, N3507);
and AND2 (N3511, N3500, N1752);
or OR4 (N3512, N3509, N2106, N2930, N1455);
or OR4 (N3513, N3510, N2354, N2551, N3339);
not NOT1 (N3514, N3482);
buf BUF1 (N3515, N3514);
and AND3 (N3516, N3502, N2773, N3265);
not NOT1 (N3517, N3499);
nand NAND4 (N3518, N3515, N456, N535, N1719);
not NOT1 (N3519, N3505);
not NOT1 (N3520, N3516);
or OR4 (N3521, N3517, N544, N1967, N1480);
xor XOR2 (N3522, N3511, N1707);
xor XOR2 (N3523, N3476, N1068);
buf BUF1 (N3524, N3521);
and AND3 (N3525, N3519, N3396, N3190);
nand NAND3 (N3526, N3524, N982, N1253);
not NOT1 (N3527, N3526);
not NOT1 (N3528, N3525);
and AND3 (N3529, N3522, N1824, N2530);
nor NOR4 (N3530, N3508, N1198, N632, N858);
nor NOR2 (N3531, N3527, N2270);
or OR4 (N3532, N3530, N1155, N865, N1911);
not NOT1 (N3533, N3532);
or OR3 (N3534, N3533, N2158, N702);
not NOT1 (N3535, N3534);
not NOT1 (N3536, N3523);
nor NOR4 (N3537, N3506, N890, N2544, N1545);
buf BUF1 (N3538, N3537);
not NOT1 (N3539, N3538);
buf BUF1 (N3540, N3518);
nor NOR4 (N3541, N3540, N1631, N1229, N517);
not NOT1 (N3542, N3520);
nor NOR3 (N3543, N3541, N3334, N1354);
and AND2 (N3544, N3529, N1083);
and AND4 (N3545, N3531, N903, N459, N3255);
nor NOR2 (N3546, N3528, N3209);
xor XOR2 (N3547, N3512, N816);
and AND2 (N3548, N3543, N2603);
and AND3 (N3549, N3548, N1198, N1173);
and AND3 (N3550, N3544, N2931, N2404);
nand NAND4 (N3551, N3550, N2180, N178, N1883);
nor NOR3 (N3552, N3547, N1270, N1047);
and AND4 (N3553, N3535, N704, N180, N610);
not NOT1 (N3554, N3513);
and AND3 (N3555, N3546, N919, N1930);
or OR4 (N3556, N3555, N1350, N549, N2233);
buf BUF1 (N3557, N3552);
and AND3 (N3558, N3557, N909, N1933);
xor XOR2 (N3559, N3545, N1477);
or OR2 (N3560, N3559, N3378);
nand NAND3 (N3561, N3539, N772, N1620);
nor NOR2 (N3562, N3560, N3327);
and AND2 (N3563, N3554, N594);
and AND2 (N3564, N3536, N3363);
xor XOR2 (N3565, N3564, N199);
and AND4 (N3566, N3549, N3490, N325, N177);
xor XOR2 (N3567, N3561, N1509);
xor XOR2 (N3568, N3565, N2257);
not NOT1 (N3569, N3567);
or OR2 (N3570, N3558, N2560);
and AND2 (N3571, N3568, N442);
or OR4 (N3572, N3569, N383, N1643, N3081);
not NOT1 (N3573, N3563);
buf BUF1 (N3574, N3553);
or OR3 (N3575, N3571, N3234, N1517);
xor XOR2 (N3576, N3574, N1296);
xor XOR2 (N3577, N3556, N3570);
and AND4 (N3578, N3158, N2038, N2752, N1157);
nor NOR4 (N3579, N3576, N358, N242, N3025);
nand NAND4 (N3580, N3572, N1938, N1603, N1417);
nor NOR3 (N3581, N3573, N2914, N975);
nor NOR4 (N3582, N3578, N2755, N1646, N560);
nand NAND3 (N3583, N3566, N287, N1799);
not NOT1 (N3584, N3575);
xor XOR2 (N3585, N3542, N3096);
or OR4 (N3586, N3585, N381, N2291, N1786);
not NOT1 (N3587, N3562);
nor NOR3 (N3588, N3583, N761, N3014);
or OR3 (N3589, N3581, N2101, N537);
buf BUF1 (N3590, N3587);
xor XOR2 (N3591, N3582, N1604);
buf BUF1 (N3592, N3584);
and AND3 (N3593, N3590, N680, N1461);
buf BUF1 (N3594, N3577);
nor NOR4 (N3595, N3588, N3072, N3513, N2176);
or OR3 (N3596, N3580, N1956, N3109);
or OR2 (N3597, N3579, N3107);
or OR3 (N3598, N3595, N246, N3010);
or OR4 (N3599, N3589, N2001, N3136, N2209);
nor NOR4 (N3600, N3599, N2586, N1443, N1944);
xor XOR2 (N3601, N3592, N946);
xor XOR2 (N3602, N3596, N1253);
not NOT1 (N3603, N3602);
nor NOR2 (N3604, N3601, N2642);
or OR2 (N3605, N3600, N1603);
or OR3 (N3606, N3605, N2815, N305);
xor XOR2 (N3607, N3551, N3537);
nand NAND2 (N3608, N3597, N1055);
nor NOR4 (N3609, N3604, N1822, N432, N2561);
buf BUF1 (N3610, N3603);
nand NAND4 (N3611, N3594, N1985, N835, N2189);
not NOT1 (N3612, N3609);
nor NOR2 (N3613, N3608, N2476);
xor XOR2 (N3614, N3607, N2725);
not NOT1 (N3615, N3598);
nor NOR2 (N3616, N3586, N1585);
or OR2 (N3617, N3612, N557);
xor XOR2 (N3618, N3614, N57);
buf BUF1 (N3619, N3613);
xor XOR2 (N3620, N3591, N1757);
nor NOR3 (N3621, N3620, N2287, N951);
nand NAND4 (N3622, N3615, N696, N1381, N3166);
or OR3 (N3623, N3618, N2463, N1986);
xor XOR2 (N3624, N3610, N2785);
nor NOR3 (N3625, N3623, N1141, N3288);
nand NAND2 (N3626, N3611, N2556);
not NOT1 (N3627, N3622);
nor NOR4 (N3628, N3606, N278, N841, N3215);
nor NOR4 (N3629, N3616, N2844, N553, N575);
and AND3 (N3630, N3617, N1093, N632);
or OR4 (N3631, N3621, N917, N2042, N684);
xor XOR2 (N3632, N3624, N2833);
and AND2 (N3633, N3630, N2068);
xor XOR2 (N3634, N3633, N2154);
or OR2 (N3635, N3629, N384);
xor XOR2 (N3636, N3635, N1530);
xor XOR2 (N3637, N3627, N1522);
buf BUF1 (N3638, N3626);
buf BUF1 (N3639, N3637);
buf BUF1 (N3640, N3639);
or OR4 (N3641, N3634, N1275, N1928, N2295);
nor NOR2 (N3642, N3625, N1688);
or OR3 (N3643, N3642, N269, N3461);
xor XOR2 (N3644, N3641, N1530);
nor NOR2 (N3645, N3628, N1446);
not NOT1 (N3646, N3644);
buf BUF1 (N3647, N3593);
buf BUF1 (N3648, N3636);
buf BUF1 (N3649, N3646);
nand NAND2 (N3650, N3649, N3554);
buf BUF1 (N3651, N3643);
or OR3 (N3652, N3638, N3221, N2080);
nand NAND2 (N3653, N3619, N340);
nand NAND2 (N3654, N3648, N1798);
or OR2 (N3655, N3653, N2327);
nor NOR3 (N3656, N3645, N2199, N1178);
nand NAND4 (N3657, N3632, N9, N562, N3505);
not NOT1 (N3658, N3652);
nor NOR3 (N3659, N3657, N3416, N325);
not NOT1 (N3660, N3659);
or OR4 (N3661, N3651, N1416, N748, N3068);
nor NOR2 (N3662, N3656, N3287);
not NOT1 (N3663, N3647);
nand NAND2 (N3664, N3660, N1950);
buf BUF1 (N3665, N3663);
or OR2 (N3666, N3650, N962);
buf BUF1 (N3667, N3662);
nor NOR2 (N3668, N3667, N937);
nand NAND2 (N3669, N3658, N3440);
buf BUF1 (N3670, N3640);
nor NOR3 (N3671, N3655, N1898, N270);
xor XOR2 (N3672, N3661, N1016);
nand NAND2 (N3673, N3665, N2942);
or OR3 (N3674, N3668, N1044, N2416);
and AND4 (N3675, N3631, N659, N1029, N2269);
or OR2 (N3676, N3673, N3428);
nor NOR3 (N3677, N3671, N1597, N3038);
nand NAND3 (N3678, N3675, N47, N2621);
xor XOR2 (N3679, N3672, N354);
not NOT1 (N3680, N3669);
xor XOR2 (N3681, N3679, N3488);
or OR2 (N3682, N3681, N2882);
and AND3 (N3683, N3677, N213, N3114);
or OR2 (N3684, N3683, N8);
nand NAND2 (N3685, N3684, N1297);
buf BUF1 (N3686, N3666);
nor NOR2 (N3687, N3676, N2946);
xor XOR2 (N3688, N3686, N213);
and AND2 (N3689, N3680, N354);
buf BUF1 (N3690, N3689);
or OR2 (N3691, N3690, N2157);
xor XOR2 (N3692, N3670, N3607);
nand NAND2 (N3693, N3682, N1049);
or OR2 (N3694, N3692, N3651);
xor XOR2 (N3695, N3694, N3551);
buf BUF1 (N3696, N3685);
and AND2 (N3697, N3664, N3549);
nor NOR2 (N3698, N3697, N1405);
xor XOR2 (N3699, N3674, N1900);
nand NAND3 (N3700, N3695, N1590, N2520);
nor NOR3 (N3701, N3698, N41, N3310);
and AND4 (N3702, N3678, N1988, N262, N1089);
or OR2 (N3703, N3699, N339);
buf BUF1 (N3704, N3693);
nor NOR3 (N3705, N3687, N1831, N3124);
not NOT1 (N3706, N3704);
xor XOR2 (N3707, N3654, N1659);
or OR3 (N3708, N3707, N1011, N3376);
and AND4 (N3709, N3700, N1510, N856, N1833);
xor XOR2 (N3710, N3703, N1073);
and AND2 (N3711, N3696, N3429);
not NOT1 (N3712, N3711);
and AND3 (N3713, N3705, N3704, N1296);
xor XOR2 (N3714, N3691, N18);
nand NAND4 (N3715, N3709, N2992, N3637, N219);
nor NOR4 (N3716, N3702, N852, N3274, N1244);
or OR4 (N3717, N3688, N1108, N3136, N3048);
nand NAND4 (N3718, N3708, N2084, N3053, N2977);
or OR3 (N3719, N3714, N1985, N2380);
xor XOR2 (N3720, N3713, N496);
nand NAND4 (N3721, N3715, N1368, N1527, N362);
nand NAND2 (N3722, N3721, N3108);
buf BUF1 (N3723, N3722);
and AND3 (N3724, N3706, N3122, N2697);
nand NAND4 (N3725, N3717, N3340, N3282, N891);
buf BUF1 (N3726, N3720);
or OR3 (N3727, N3726, N2139, N221);
nor NOR3 (N3728, N3725, N2805, N1134);
nand NAND3 (N3729, N3728, N2841, N2960);
xor XOR2 (N3730, N3701, N1887);
buf BUF1 (N3731, N3730);
buf BUF1 (N3732, N3712);
not NOT1 (N3733, N3731);
not NOT1 (N3734, N3724);
nand NAND4 (N3735, N3723, N2357, N1224, N3347);
nand NAND2 (N3736, N3732, N1821);
nand NAND2 (N3737, N3727, N1331);
nor NOR4 (N3738, N3729, N303, N2764, N1252);
xor XOR2 (N3739, N3718, N3302);
nand NAND3 (N3740, N3738, N50, N3234);
or OR2 (N3741, N3739, N2613);
buf BUF1 (N3742, N3736);
nand NAND3 (N3743, N3742, N700, N1429);
not NOT1 (N3744, N3716);
or OR2 (N3745, N3735, N649);
not NOT1 (N3746, N3740);
or OR2 (N3747, N3745, N131);
or OR4 (N3748, N3719, N55, N53, N786);
not NOT1 (N3749, N3737);
buf BUF1 (N3750, N3744);
and AND4 (N3751, N3746, N1685, N890, N1450);
nor NOR4 (N3752, N3748, N1029, N2530, N1307);
xor XOR2 (N3753, N3752, N519);
xor XOR2 (N3754, N3751, N983);
and AND2 (N3755, N3743, N835);
nand NAND3 (N3756, N3710, N3199, N3689);
or OR4 (N3757, N3756, N1909, N2180, N575);
not NOT1 (N3758, N3753);
and AND2 (N3759, N3733, N3571);
or OR2 (N3760, N3757, N3654);
or OR2 (N3761, N3754, N910);
nor NOR2 (N3762, N3747, N3050);
not NOT1 (N3763, N3762);
nor NOR4 (N3764, N3755, N2883, N1250, N3733);
nor NOR3 (N3765, N3758, N2358, N2480);
nand NAND3 (N3766, N3760, N1393, N3348);
nand NAND4 (N3767, N3750, N1389, N2707, N1737);
xor XOR2 (N3768, N3763, N3542);
not NOT1 (N3769, N3749);
not NOT1 (N3770, N3766);
nor NOR2 (N3771, N3768, N1198);
xor XOR2 (N3772, N3767, N3123);
buf BUF1 (N3773, N3764);
nand NAND2 (N3774, N3769, N3469);
not NOT1 (N3775, N3761);
and AND3 (N3776, N3771, N3231, N3657);
nand NAND4 (N3777, N3741, N741, N2008, N3174);
nor NOR4 (N3778, N3776, N2021, N3353, N1646);
or OR4 (N3779, N3759, N3323, N3375, N2082);
nand NAND3 (N3780, N3779, N217, N1822);
nor NOR4 (N3781, N3780, N1568, N2755, N3776);
nand NAND2 (N3782, N3775, N932);
not NOT1 (N3783, N3770);
xor XOR2 (N3784, N3734, N459);
nand NAND2 (N3785, N3784, N1418);
not NOT1 (N3786, N3774);
buf BUF1 (N3787, N3783);
not NOT1 (N3788, N3778);
xor XOR2 (N3789, N3782, N455);
buf BUF1 (N3790, N3781);
not NOT1 (N3791, N3790);
or OR3 (N3792, N3787, N1271, N3749);
not NOT1 (N3793, N3791);
buf BUF1 (N3794, N3786);
nand NAND4 (N3795, N3777, N326, N2965, N1769);
nand NAND4 (N3796, N3788, N3695, N839, N738);
buf BUF1 (N3797, N3772);
buf BUF1 (N3798, N3789);
nor NOR2 (N3799, N3795, N3601);
and AND2 (N3800, N3785, N1852);
buf BUF1 (N3801, N3798);
buf BUF1 (N3802, N3800);
not NOT1 (N3803, N3801);
nand NAND3 (N3804, N3802, N797, N986);
buf BUF1 (N3805, N3796);
and AND4 (N3806, N3792, N1283, N1720, N322);
nor NOR2 (N3807, N3803, N495);
nand NAND3 (N3808, N3794, N2529, N3274);
xor XOR2 (N3809, N3773, N1385);
or OR4 (N3810, N3809, N1542, N827, N909);
buf BUF1 (N3811, N3810);
and AND4 (N3812, N3797, N1688, N556, N3431);
buf BUF1 (N3813, N3808);
or OR2 (N3814, N3812, N247);
not NOT1 (N3815, N3814);
or OR4 (N3816, N3765, N445, N3547, N3299);
buf BUF1 (N3817, N3807);
nor NOR2 (N3818, N3811, N3117);
xor XOR2 (N3819, N3804, N2214);
or OR4 (N3820, N3818, N2383, N678, N1276);
and AND2 (N3821, N3817, N605);
or OR2 (N3822, N3806, N2443);
nand NAND4 (N3823, N3805, N908, N2548, N1891);
nand NAND3 (N3824, N3813, N3797, N2600);
and AND4 (N3825, N3821, N2366, N1496, N2936);
buf BUF1 (N3826, N3793);
xor XOR2 (N3827, N3825, N3634);
nand NAND2 (N3828, N3819, N2497);
nand NAND4 (N3829, N3823, N1416, N421, N942);
not NOT1 (N3830, N3829);
and AND4 (N3831, N3816, N1814, N945, N1660);
nor NOR2 (N3832, N3815, N2138);
xor XOR2 (N3833, N3830, N959);
nand NAND3 (N3834, N3826, N3056, N1600);
or OR4 (N3835, N3822, N2177, N197, N1788);
not NOT1 (N3836, N3828);
nand NAND2 (N3837, N3835, N2781);
not NOT1 (N3838, N3824);
nor NOR4 (N3839, N3827, N1844, N1495, N457);
and AND3 (N3840, N3836, N3487, N1854);
xor XOR2 (N3841, N3838, N2989);
nor NOR4 (N3842, N3837, N1538, N1675, N848);
or OR2 (N3843, N3834, N1103);
nor NOR4 (N3844, N3820, N1435, N3195, N1059);
and AND3 (N3845, N3832, N1783, N190);
nand NAND4 (N3846, N3841, N1498, N3700, N1041);
nand NAND3 (N3847, N3845, N3338, N1323);
or OR3 (N3848, N3843, N509, N581);
nand NAND4 (N3849, N3847, N13, N3290, N2068);
buf BUF1 (N3850, N3831);
or OR3 (N3851, N3839, N2658, N1783);
nand NAND2 (N3852, N3799, N1692);
and AND3 (N3853, N3844, N3646, N413);
and AND3 (N3854, N3851, N3624, N1754);
buf BUF1 (N3855, N3854);
and AND3 (N3856, N3849, N3617, N806);
nand NAND2 (N3857, N3850, N693);
xor XOR2 (N3858, N3853, N538);
not NOT1 (N3859, N3846);
buf BUF1 (N3860, N3859);
buf BUF1 (N3861, N3857);
not NOT1 (N3862, N3848);
or OR3 (N3863, N3852, N1229, N1619);
buf BUF1 (N3864, N3855);
or OR3 (N3865, N3860, N2465, N2342);
nor NOR4 (N3866, N3861, N3379, N721, N1494);
nor NOR3 (N3867, N3833, N33, N3794);
buf BUF1 (N3868, N3856);
and AND4 (N3869, N3867, N1407, N905, N249);
nand NAND4 (N3870, N3866, N1595, N3026, N748);
nand NAND2 (N3871, N3870, N3220);
and AND4 (N3872, N3864, N339, N1597, N2118);
nand NAND3 (N3873, N3869, N132, N1155);
buf BUF1 (N3874, N3868);
or OR4 (N3875, N3874, N334, N676, N951);
nor NOR3 (N3876, N3872, N2041, N1657);
not NOT1 (N3877, N3863);
buf BUF1 (N3878, N3858);
xor XOR2 (N3879, N3878, N2420);
nand NAND2 (N3880, N3873, N1746);
and AND3 (N3881, N3871, N735, N1619);
or OR4 (N3882, N3881, N621, N3263, N3645);
not NOT1 (N3883, N3865);
nand NAND3 (N3884, N3880, N3114, N1288);
not NOT1 (N3885, N3876);
buf BUF1 (N3886, N3882);
xor XOR2 (N3887, N3862, N615);
not NOT1 (N3888, N3887);
xor XOR2 (N3889, N3884, N1377);
nand NAND4 (N3890, N3879, N2065, N3791, N1100);
nor NOR4 (N3891, N3877, N754, N2894, N2442);
xor XOR2 (N3892, N3883, N2221);
or OR4 (N3893, N3840, N2446, N1071, N42);
nand NAND4 (N3894, N3886, N451, N3503, N3606);
buf BUF1 (N3895, N3842);
buf BUF1 (N3896, N3889);
buf BUF1 (N3897, N3891);
not NOT1 (N3898, N3893);
xor XOR2 (N3899, N3897, N81);
buf BUF1 (N3900, N3888);
xor XOR2 (N3901, N3875, N2512);
buf BUF1 (N3902, N3900);
not NOT1 (N3903, N3890);
or OR3 (N3904, N3902, N1532, N272);
or OR3 (N3905, N3904, N3271, N2133);
xor XOR2 (N3906, N3896, N1283);
xor XOR2 (N3907, N3903, N2815);
or OR3 (N3908, N3895, N2672, N1262);
or OR3 (N3909, N3908, N3840, N848);
xor XOR2 (N3910, N3906, N2354);
nor NOR4 (N3911, N3905, N627, N3746, N2128);
buf BUF1 (N3912, N3885);
not NOT1 (N3913, N3907);
nor NOR3 (N3914, N3910, N3767, N3258);
nand NAND2 (N3915, N3892, N24);
nor NOR3 (N3916, N3915, N1343, N932);
xor XOR2 (N3917, N3894, N106);
buf BUF1 (N3918, N3901);
or OR4 (N3919, N3899, N1476, N1368, N1570);
nand NAND3 (N3920, N3919, N2214, N3763);
nor NOR4 (N3921, N3911, N3830, N1364, N2851);
xor XOR2 (N3922, N3920, N3776);
buf BUF1 (N3923, N3917);
not NOT1 (N3924, N3922);
not NOT1 (N3925, N3924);
xor XOR2 (N3926, N3898, N1661);
and AND4 (N3927, N3921, N2234, N187, N3864);
nor NOR2 (N3928, N3916, N3664);
xor XOR2 (N3929, N3927, N151);
and AND4 (N3930, N3912, N1114, N580, N671);
or OR3 (N3931, N3930, N2531, N44);
nor NOR3 (N3932, N3913, N736, N2037);
nor NOR3 (N3933, N3914, N2090, N2529);
nor NOR4 (N3934, N3918, N3294, N1906, N1790);
and AND2 (N3935, N3929, N716);
buf BUF1 (N3936, N3923);
nor NOR3 (N3937, N3935, N3205, N26);
xor XOR2 (N3938, N3928, N3790);
buf BUF1 (N3939, N3931);
not NOT1 (N3940, N3937);
nor NOR2 (N3941, N3934, N304);
xor XOR2 (N3942, N3938, N1784);
or OR2 (N3943, N3941, N3085);
nand NAND3 (N3944, N3940, N2201, N2424);
nand NAND3 (N3945, N3943, N1495, N2524);
not NOT1 (N3946, N3942);
or OR3 (N3947, N3925, N2317, N3748);
or OR4 (N3948, N3939, N3137, N2505, N1711);
nand NAND2 (N3949, N3932, N455);
nor NOR3 (N3950, N3949, N1254, N1636);
buf BUF1 (N3951, N3945);
not NOT1 (N3952, N3951);
nor NOR4 (N3953, N3950, N1342, N2451, N2493);
or OR3 (N3954, N3944, N2218, N1801);
and AND4 (N3955, N3909, N2452, N3302, N653);
not NOT1 (N3956, N3926);
nor NOR4 (N3957, N3954, N3340, N3475, N108);
nand NAND4 (N3958, N3948, N3439, N2132, N484);
nor NOR2 (N3959, N3936, N2787);
nand NAND4 (N3960, N3947, N2437, N2829, N2777);
not NOT1 (N3961, N3933);
buf BUF1 (N3962, N3955);
or OR2 (N3963, N3956, N2859);
nand NAND4 (N3964, N3962, N3102, N2602, N1402);
not NOT1 (N3965, N3957);
xor XOR2 (N3966, N3960, N914);
nand NAND2 (N3967, N3953, N2422);
nand NAND3 (N3968, N3966, N3867, N3086);
and AND2 (N3969, N3958, N2840);
not NOT1 (N3970, N3964);
or OR2 (N3971, N3963, N3081);
xor XOR2 (N3972, N3961, N662);
nor NOR3 (N3973, N3946, N3937, N3361);
not NOT1 (N3974, N3952);
nor NOR3 (N3975, N3973, N565, N2487);
or OR2 (N3976, N3965, N203);
buf BUF1 (N3977, N3972);
nor NOR2 (N3978, N3959, N2415);
and AND4 (N3979, N3975, N2603, N3896, N955);
or OR2 (N3980, N3978, N3682);
nand NAND2 (N3981, N3969, N984);
nor NOR2 (N3982, N3981, N3241);
nor NOR4 (N3983, N3976, N1943, N1566, N3233);
and AND2 (N3984, N3977, N3514);
and AND3 (N3985, N3974, N1662, N1042);
buf BUF1 (N3986, N3979);
nor NOR2 (N3987, N3971, N538);
not NOT1 (N3988, N3986);
nor NOR4 (N3989, N3967, N3662, N863, N3356);
nand NAND3 (N3990, N3987, N192, N3238);
buf BUF1 (N3991, N3989);
or OR3 (N3992, N3990, N1592, N1202);
nand NAND3 (N3993, N3980, N915, N2413);
nor NOR3 (N3994, N3992, N2907, N3256);
nand NAND4 (N3995, N3991, N3934, N3506, N320);
or OR4 (N3996, N3993, N2103, N3556, N628);
not NOT1 (N3997, N3996);
or OR3 (N3998, N3984, N2634, N3189);
or OR3 (N3999, N3983, N174, N255);
nor NOR3 (N4000, N3994, N1400, N1550);
xor XOR2 (N4001, N4000, N1783);
not NOT1 (N4002, N4001);
xor XOR2 (N4003, N3968, N3663);
not NOT1 (N4004, N3982);
or OR3 (N4005, N3970, N2192, N2178);
nor NOR3 (N4006, N3995, N3821, N769);
nand NAND3 (N4007, N4006, N1564, N308);
xor XOR2 (N4008, N3998, N543);
xor XOR2 (N4009, N3988, N435);
nor NOR4 (N4010, N4003, N676, N613, N2203);
buf BUF1 (N4011, N4008);
or OR2 (N4012, N4011, N2173);
or OR3 (N4013, N4005, N3763, N349);
nor NOR4 (N4014, N3985, N3185, N1569, N2248);
buf BUF1 (N4015, N3997);
buf BUF1 (N4016, N4012);
buf BUF1 (N4017, N4013);
nor NOR3 (N4018, N4007, N3558, N2465);
nand NAND4 (N4019, N4002, N2325, N2425, N3485);
nand NAND4 (N4020, N4009, N1702, N1686, N228);
xor XOR2 (N4021, N4018, N105);
or OR3 (N4022, N4004, N4008, N3146);
xor XOR2 (N4023, N3999, N128);
not NOT1 (N4024, N4023);
and AND2 (N4025, N4021, N908);
xor XOR2 (N4026, N4020, N1731);
buf BUF1 (N4027, N4016);
nor NOR3 (N4028, N4025, N2466, N1411);
not NOT1 (N4029, N4015);
and AND3 (N4030, N4024, N1093, N1500);
nor NOR3 (N4031, N4030, N765, N172);
not NOT1 (N4032, N4029);
not NOT1 (N4033, N4017);
buf BUF1 (N4034, N4031);
buf BUF1 (N4035, N4014);
or OR3 (N4036, N4034, N2954, N1451);
nor NOR2 (N4037, N4036, N93);
and AND2 (N4038, N4010, N2704);
nand NAND3 (N4039, N4037, N2214, N386);
or OR3 (N4040, N4033, N3492, N848);
buf BUF1 (N4041, N4027);
buf BUF1 (N4042, N4028);
nor NOR2 (N4043, N4038, N1196);
buf BUF1 (N4044, N4022);
xor XOR2 (N4045, N4032, N3385);
xor XOR2 (N4046, N4041, N1427);
xor XOR2 (N4047, N4040, N2796);
buf BUF1 (N4048, N4019);
and AND4 (N4049, N4046, N657, N2289, N801);
not NOT1 (N4050, N4047);
nand NAND3 (N4051, N4050, N968, N3428);
buf BUF1 (N4052, N4048);
and AND3 (N4053, N4039, N2086, N2524);
nor NOR3 (N4054, N4051, N1437, N3010);
not NOT1 (N4055, N4054);
buf BUF1 (N4056, N4055);
or OR4 (N4057, N4026, N1317, N25, N2360);
nor NOR3 (N4058, N4056, N2038, N979);
nand NAND2 (N4059, N4058, N1501);
not NOT1 (N4060, N4043);
nand NAND2 (N4061, N4049, N3877);
buf BUF1 (N4062, N4060);
or OR3 (N4063, N4035, N341, N1961);
and AND2 (N4064, N4057, N2702);
not NOT1 (N4065, N4062);
nand NAND4 (N4066, N4063, N2945, N1489, N2096);
not NOT1 (N4067, N4045);
and AND4 (N4068, N4059, N3588, N2348, N3561);
xor XOR2 (N4069, N4044, N2125);
nor NOR3 (N4070, N4053, N3395, N1047);
xor XOR2 (N4071, N4067, N969);
buf BUF1 (N4072, N4070);
or OR4 (N4073, N4066, N2991, N1757, N1714);
and AND2 (N4074, N4042, N2949);
not NOT1 (N4075, N4052);
and AND3 (N4076, N4072, N1148, N793);
buf BUF1 (N4077, N4075);
xor XOR2 (N4078, N4076, N3761);
or OR2 (N4079, N4068, N1289);
buf BUF1 (N4080, N4064);
nand NAND2 (N4081, N4078, N2719);
nor NOR3 (N4082, N4065, N131, N1270);
nor NOR4 (N4083, N4061, N3651, N3344, N2844);
not NOT1 (N4084, N4079);
buf BUF1 (N4085, N4074);
xor XOR2 (N4086, N4071, N1173);
xor XOR2 (N4087, N4077, N3710);
or OR4 (N4088, N4087, N875, N2146, N2625);
and AND2 (N4089, N4084, N1684);
nand NAND2 (N4090, N4082, N3541);
xor XOR2 (N4091, N4081, N1781);
not NOT1 (N4092, N4091);
or OR3 (N4093, N4088, N2627, N14);
not NOT1 (N4094, N4092);
buf BUF1 (N4095, N4073);
not NOT1 (N4096, N4086);
and AND4 (N4097, N4095, N1593, N1933, N2780);
or OR2 (N4098, N4096, N190);
or OR3 (N4099, N4094, N3256, N2317);
not NOT1 (N4100, N4097);
not NOT1 (N4101, N4093);
nand NAND4 (N4102, N4083, N2661, N2062, N839);
and AND2 (N4103, N4085, N445);
nor NOR3 (N4104, N4069, N3401, N3410);
nand NAND2 (N4105, N4090, N438);
and AND3 (N4106, N4103, N3270, N1585);
not NOT1 (N4107, N4080);
nor NOR3 (N4108, N4100, N3992, N3394);
or OR4 (N4109, N4108, N2770, N2339, N50);
nand NAND4 (N4110, N4104, N206, N4006, N3298);
not NOT1 (N4111, N4109);
and AND3 (N4112, N4107, N1034, N2890);
nand NAND2 (N4113, N4110, N3916);
or OR3 (N4114, N4089, N3849, N3731);
and AND2 (N4115, N4111, N615);
not NOT1 (N4116, N4112);
nand NAND4 (N4117, N4098, N774, N2594, N1453);
nand NAND3 (N4118, N4099, N2592, N467);
and AND3 (N4119, N4101, N975, N3905);
buf BUF1 (N4120, N4117);
xor XOR2 (N4121, N4120, N1963);
or OR2 (N4122, N4121, N3454);
nor NOR3 (N4123, N4106, N1649, N3462);
or OR2 (N4124, N4113, N1306);
or OR2 (N4125, N4116, N2959);
buf BUF1 (N4126, N4123);
xor XOR2 (N4127, N4105, N1974);
buf BUF1 (N4128, N4122);
and AND2 (N4129, N4128, N1703);
and AND4 (N4130, N4119, N1033, N4117, N7);
xor XOR2 (N4131, N4129, N1890);
or OR3 (N4132, N4130, N2150, N3345);
or OR2 (N4133, N4132, N94);
xor XOR2 (N4134, N4133, N325);
buf BUF1 (N4135, N4134);
xor XOR2 (N4136, N4126, N4026);
nor NOR3 (N4137, N4135, N2859, N1988);
and AND2 (N4138, N4137, N1823);
nor NOR4 (N4139, N4136, N2694, N981, N2711);
buf BUF1 (N4140, N4118);
buf BUF1 (N4141, N4138);
not NOT1 (N4142, N4140);
buf BUF1 (N4143, N4127);
nor NOR3 (N4144, N4141, N3835, N2506);
or OR4 (N4145, N4144, N1158, N2948, N1973);
nand NAND2 (N4146, N4145, N2951);
nor NOR2 (N4147, N4139, N2453);
buf BUF1 (N4148, N4147);
buf BUF1 (N4149, N4143);
and AND4 (N4150, N4146, N3320, N1686, N815);
not NOT1 (N4151, N4102);
xor XOR2 (N4152, N4124, N519);
and AND2 (N4153, N4114, N3466);
and AND3 (N4154, N4152, N909, N2602);
xor XOR2 (N4155, N4150, N2214);
nand NAND4 (N4156, N4151, N739, N14, N2011);
xor XOR2 (N4157, N4153, N3625);
nor NOR2 (N4158, N4148, N528);
xor XOR2 (N4159, N4158, N4107);
xor XOR2 (N4160, N4125, N82);
nor NOR2 (N4161, N4160, N3381);
nor NOR2 (N4162, N4161, N3798);
or OR3 (N4163, N4131, N863, N2542);
xor XOR2 (N4164, N4162, N3403);
nand NAND2 (N4165, N4115, N3364);
or OR3 (N4166, N4163, N1410, N2386);
or OR2 (N4167, N4149, N2313);
xor XOR2 (N4168, N4164, N1236);
nand NAND2 (N4169, N4159, N3656);
xor XOR2 (N4170, N4155, N1245);
buf BUF1 (N4171, N4168);
not NOT1 (N4172, N4171);
and AND4 (N4173, N4166, N2372, N11, N370);
and AND2 (N4174, N4154, N3953);
xor XOR2 (N4175, N4157, N2081);
buf BUF1 (N4176, N4165);
and AND2 (N4177, N4174, N2391);
nor NOR4 (N4178, N4177, N3693, N2543, N1634);
nand NAND3 (N4179, N4167, N1298, N422);
xor XOR2 (N4180, N4169, N103);
xor XOR2 (N4181, N4179, N3341);
nor NOR4 (N4182, N4156, N3745, N416, N611);
buf BUF1 (N4183, N4172);
not NOT1 (N4184, N4175);
or OR2 (N4185, N4180, N1107);
xor XOR2 (N4186, N4185, N1122);
nor NOR2 (N4187, N4178, N952);
or OR3 (N4188, N4176, N605, N138);
nor NOR2 (N4189, N4182, N651);
and AND2 (N4190, N4189, N972);
not NOT1 (N4191, N4187);
nor NOR2 (N4192, N4186, N355);
not NOT1 (N4193, N4184);
nor NOR3 (N4194, N4173, N2724, N3867);
not NOT1 (N4195, N4188);
and AND4 (N4196, N4183, N962, N673, N984);
nand NAND3 (N4197, N4195, N1603, N3860);
xor XOR2 (N4198, N4142, N3021);
xor XOR2 (N4199, N4197, N1205);
nand NAND2 (N4200, N4198, N2844);
and AND2 (N4201, N4199, N1447);
and AND3 (N4202, N4192, N700, N2655);
and AND3 (N4203, N4202, N2992, N784);
buf BUF1 (N4204, N4181);
and AND3 (N4205, N4204, N1536, N2237);
not NOT1 (N4206, N4191);
nor NOR3 (N4207, N4196, N4057, N3757);
or OR3 (N4208, N4194, N2740, N431);
nor NOR3 (N4209, N4207, N2083, N1522);
not NOT1 (N4210, N4206);
nand NAND4 (N4211, N4200, N91, N4038, N109);
buf BUF1 (N4212, N4209);
buf BUF1 (N4213, N4201);
buf BUF1 (N4214, N4205);
xor XOR2 (N4215, N4193, N1650);
not NOT1 (N4216, N4211);
and AND2 (N4217, N4213, N3328);
not NOT1 (N4218, N4210);
and AND2 (N4219, N4190, N127);
xor XOR2 (N4220, N4203, N832);
buf BUF1 (N4221, N4215);
not NOT1 (N4222, N4221);
not NOT1 (N4223, N4218);
nand NAND2 (N4224, N4223, N2614);
buf BUF1 (N4225, N4170);
or OR2 (N4226, N4222, N3445);
and AND4 (N4227, N4214, N2460, N295, N2886);
nor NOR3 (N4228, N4224, N1741, N816);
nor NOR3 (N4229, N4227, N2020, N3523);
and AND3 (N4230, N4225, N2985, N1507);
nor NOR2 (N4231, N4226, N3355);
and AND2 (N4232, N4217, N1913);
xor XOR2 (N4233, N4216, N1814);
nand NAND3 (N4234, N4229, N3646, N2533);
buf BUF1 (N4235, N4230);
or OR4 (N4236, N4208, N1143, N349, N318);
xor XOR2 (N4237, N4232, N4001);
buf BUF1 (N4238, N4212);
buf BUF1 (N4239, N4219);
xor XOR2 (N4240, N4220, N2600);
nand NAND3 (N4241, N4240, N737, N2119);
and AND2 (N4242, N4239, N1050);
and AND2 (N4243, N4238, N2261);
not NOT1 (N4244, N4234);
or OR4 (N4245, N4243, N3467, N1920, N1321);
xor XOR2 (N4246, N4233, N3266);
and AND4 (N4247, N4246, N262, N959, N1047);
and AND4 (N4248, N4244, N39, N955, N1923);
and AND4 (N4249, N4228, N306, N697, N1509);
not NOT1 (N4250, N4247);
not NOT1 (N4251, N4242);
or OR4 (N4252, N4249, N2724, N1474, N1632);
xor XOR2 (N4253, N4235, N1017);
xor XOR2 (N4254, N4236, N3812);
xor XOR2 (N4255, N4237, N3565);
nor NOR4 (N4256, N4248, N241, N473, N1478);
and AND4 (N4257, N4250, N1071, N1062, N3297);
or OR2 (N4258, N4251, N2903);
or OR3 (N4259, N4256, N3824, N1330);
xor XOR2 (N4260, N4255, N1109);
xor XOR2 (N4261, N4241, N2994);
nand NAND2 (N4262, N4261, N4244);
xor XOR2 (N4263, N4254, N3374);
xor XOR2 (N4264, N4257, N1411);
not NOT1 (N4265, N4259);
or OR3 (N4266, N4252, N2232, N3913);
or OR4 (N4267, N4263, N2328, N3708, N2102);
nor NOR2 (N4268, N4260, N4140);
buf BUF1 (N4269, N4268);
not NOT1 (N4270, N4269);
and AND4 (N4271, N4266, N3797, N141, N2381);
and AND3 (N4272, N4264, N3606, N3277);
and AND4 (N4273, N4265, N2614, N3977, N680);
buf BUF1 (N4274, N4273);
nand NAND2 (N4275, N4274, N4014);
buf BUF1 (N4276, N4262);
nor NOR2 (N4277, N4253, N1893);
nor NOR4 (N4278, N4231, N1234, N3302, N1965);
xor XOR2 (N4279, N4267, N1144);
not NOT1 (N4280, N4276);
or OR3 (N4281, N4277, N3090, N195);
not NOT1 (N4282, N4278);
xor XOR2 (N4283, N4282, N1214);
and AND3 (N4284, N4258, N4225, N464);
nand NAND3 (N4285, N4281, N2567, N384);
and AND3 (N4286, N4245, N3816, N596);
not NOT1 (N4287, N4275);
nor NOR4 (N4288, N4286, N388, N3034, N1448);
nor NOR4 (N4289, N4279, N2652, N888, N3889);
buf BUF1 (N4290, N4288);
buf BUF1 (N4291, N4290);
buf BUF1 (N4292, N4284);
nor NOR4 (N4293, N4292, N284, N89, N2269);
and AND4 (N4294, N4291, N172, N1719, N3039);
and AND3 (N4295, N4294, N1611, N207);
and AND3 (N4296, N4285, N3867, N418);
nor NOR3 (N4297, N4270, N381, N1449);
nor NOR4 (N4298, N4280, N2461, N1600, N3682);
not NOT1 (N4299, N4296);
or OR3 (N4300, N4272, N1911, N963);
nor NOR2 (N4301, N4299, N2920);
or OR2 (N4302, N4295, N512);
xor XOR2 (N4303, N4289, N703);
buf BUF1 (N4304, N4302);
nand NAND3 (N4305, N4293, N1657, N2733);
and AND3 (N4306, N4304, N1435, N80);
not NOT1 (N4307, N4271);
or OR2 (N4308, N4300, N934);
buf BUF1 (N4309, N4283);
or OR4 (N4310, N4305, N1208, N1528, N2697);
or OR2 (N4311, N4301, N213);
and AND2 (N4312, N4307, N1125);
xor XOR2 (N4313, N4287, N3108);
nor NOR2 (N4314, N4303, N2637);
nand NAND2 (N4315, N4311, N3935);
buf BUF1 (N4316, N4315);
buf BUF1 (N4317, N4309);
or OR3 (N4318, N4317, N741, N3691);
nand NAND2 (N4319, N4306, N2829);
buf BUF1 (N4320, N4298);
and AND2 (N4321, N4319, N3039);
nor NOR2 (N4322, N4314, N2025);
nand NAND4 (N4323, N4318, N2291, N452, N3239);
not NOT1 (N4324, N4320);
xor XOR2 (N4325, N4308, N3592);
xor XOR2 (N4326, N4297, N1113);
buf BUF1 (N4327, N4321);
nor NOR3 (N4328, N4327, N2156, N2864);
or OR3 (N4329, N4326, N4068, N574);
and AND3 (N4330, N4329, N3361, N2093);
not NOT1 (N4331, N4325);
nand NAND2 (N4332, N4323, N3767);
buf BUF1 (N4333, N4331);
and AND2 (N4334, N4313, N2538);
nand NAND4 (N4335, N4333, N1596, N3360, N652);
and AND4 (N4336, N4328, N3136, N719, N2593);
not NOT1 (N4337, N4332);
nand NAND3 (N4338, N4322, N92, N451);
or OR3 (N4339, N4335, N3525, N381);
nor NOR2 (N4340, N4337, N3292);
and AND4 (N4341, N4310, N1375, N3412, N630);
nand NAND3 (N4342, N4324, N2035, N2429);
nand NAND2 (N4343, N4341, N3673);
nand NAND3 (N4344, N4340, N676, N2246);
buf BUF1 (N4345, N4344);
and AND4 (N4346, N4312, N1058, N144, N877);
buf BUF1 (N4347, N4342);
nand NAND3 (N4348, N4343, N3082, N885);
nand NAND2 (N4349, N4330, N2501);
xor XOR2 (N4350, N4345, N3037);
buf BUF1 (N4351, N4339);
buf BUF1 (N4352, N4334);
xor XOR2 (N4353, N4348, N2660);
nand NAND4 (N4354, N4349, N3671, N104, N1321);
nor NOR4 (N4355, N4347, N248, N3142, N757);
xor XOR2 (N4356, N4338, N2437);
nor NOR2 (N4357, N4346, N3977);
nor NOR2 (N4358, N4350, N4151);
not NOT1 (N4359, N4354);
nor NOR4 (N4360, N4353, N3248, N2109, N2007);
buf BUF1 (N4361, N4336);
or OR3 (N4362, N4352, N3639, N3127);
buf BUF1 (N4363, N4360);
not NOT1 (N4364, N4351);
or OR2 (N4365, N4362, N272);
nor NOR4 (N4366, N4355, N1209, N4244, N1619);
or OR2 (N4367, N4366, N1093);
or OR4 (N4368, N4363, N1584, N2167, N4068);
not NOT1 (N4369, N4361);
xor XOR2 (N4370, N4356, N1467);
not NOT1 (N4371, N4367);
nor NOR4 (N4372, N4368, N4041, N393, N192);
nor NOR2 (N4373, N4357, N1079);
nor NOR4 (N4374, N4364, N2283, N63, N3743);
or OR2 (N4375, N4370, N2226);
xor XOR2 (N4376, N4372, N2613);
and AND4 (N4377, N4369, N2618, N2532, N1106);
not NOT1 (N4378, N4365);
xor XOR2 (N4379, N4373, N1475);
buf BUF1 (N4380, N4376);
buf BUF1 (N4381, N4374);
not NOT1 (N4382, N4381);
nor NOR4 (N4383, N4375, N1549, N559, N4172);
not NOT1 (N4384, N4380);
xor XOR2 (N4385, N4383, N1844);
xor XOR2 (N4386, N4385, N3498);
and AND4 (N4387, N4358, N2011, N2676, N552);
nand NAND2 (N4388, N4316, N1045);
not NOT1 (N4389, N4387);
and AND4 (N4390, N4388, N52, N3650, N315);
not NOT1 (N4391, N4389);
buf BUF1 (N4392, N4379);
nand NAND3 (N4393, N4377, N3937, N3399);
buf BUF1 (N4394, N4371);
nand NAND4 (N4395, N4359, N3343, N2376, N3058);
not NOT1 (N4396, N4390);
nor NOR3 (N4397, N4394, N2787, N4300);
or OR2 (N4398, N4384, N1464);
xor XOR2 (N4399, N4395, N3847);
and AND4 (N4400, N4396, N2262, N2858, N3930);
or OR4 (N4401, N4386, N3407, N3048, N19);
nand NAND4 (N4402, N4382, N1276, N2792, N3670);
not NOT1 (N4403, N4399);
xor XOR2 (N4404, N4397, N3480);
buf BUF1 (N4405, N4404);
and AND4 (N4406, N4401, N778, N2765, N418);
or OR2 (N4407, N4378, N481);
or OR2 (N4408, N4392, N2149);
xor XOR2 (N4409, N4408, N676);
and AND3 (N4410, N4398, N1122, N1808);
or OR3 (N4411, N4407, N1737, N2742);
not NOT1 (N4412, N4400);
and AND3 (N4413, N4405, N633, N692);
xor XOR2 (N4414, N4413, N477);
nor NOR3 (N4415, N4403, N3777, N1383);
xor XOR2 (N4416, N4409, N3115);
xor XOR2 (N4417, N4402, N3460);
and AND3 (N4418, N4406, N899, N3033);
xor XOR2 (N4419, N4411, N4225);
buf BUF1 (N4420, N4416);
not NOT1 (N4421, N4393);
not NOT1 (N4422, N4419);
not NOT1 (N4423, N4418);
buf BUF1 (N4424, N4412);
and AND3 (N4425, N4414, N2917, N3375);
or OR3 (N4426, N4423, N292, N3551);
buf BUF1 (N4427, N4424);
and AND3 (N4428, N4421, N4255, N4062);
xor XOR2 (N4429, N4426, N2370);
buf BUF1 (N4430, N4422);
xor XOR2 (N4431, N4417, N4419);
nor NOR2 (N4432, N4430, N780);
nand NAND2 (N4433, N4427, N2710);
and AND2 (N4434, N4432, N594);
not NOT1 (N4435, N4434);
nand NAND2 (N4436, N4410, N2898);
nor NOR3 (N4437, N4431, N2622, N1325);
nand NAND3 (N4438, N4435, N782, N2845);
not NOT1 (N4439, N4429);
buf BUF1 (N4440, N4438);
not NOT1 (N4441, N4436);
not NOT1 (N4442, N4437);
or OR3 (N4443, N4440, N4372, N3083);
not NOT1 (N4444, N4425);
xor XOR2 (N4445, N4442, N697);
xor XOR2 (N4446, N4444, N1397);
nor NOR2 (N4447, N4433, N1167);
and AND4 (N4448, N4446, N1670, N791, N2308);
and AND2 (N4449, N4428, N3391);
and AND3 (N4450, N4391, N3100, N2197);
or OR3 (N4451, N4445, N550, N2703);
xor XOR2 (N4452, N4420, N2639);
and AND2 (N4453, N4441, N550);
xor XOR2 (N4454, N4452, N2573);
xor XOR2 (N4455, N4439, N2978);
and AND4 (N4456, N4450, N2887, N2928, N2901);
and AND4 (N4457, N4447, N1853, N1443, N4094);
buf BUF1 (N4458, N4443);
xor XOR2 (N4459, N4454, N4144);
not NOT1 (N4460, N4459);
xor XOR2 (N4461, N4455, N2518);
xor XOR2 (N4462, N4448, N3122);
or OR4 (N4463, N4415, N3510, N304, N4349);
and AND2 (N4464, N4453, N2762);
or OR4 (N4465, N4458, N4254, N1994, N54);
xor XOR2 (N4466, N4456, N4054);
and AND2 (N4467, N4451, N1556);
nor NOR2 (N4468, N4465, N1677);
nor NOR2 (N4469, N4461, N680);
or OR3 (N4470, N4468, N377, N4037);
not NOT1 (N4471, N4462);
and AND3 (N4472, N4466, N3951, N1466);
and AND4 (N4473, N4471, N4357, N146, N2843);
or OR4 (N4474, N4449, N3386, N1412, N2590);
buf BUF1 (N4475, N4473);
and AND2 (N4476, N4457, N3040);
and AND3 (N4477, N4469, N3977, N10);
and AND2 (N4478, N4475, N959);
xor XOR2 (N4479, N4460, N1008);
or OR4 (N4480, N4477, N4403, N433, N4058);
buf BUF1 (N4481, N4467);
nand NAND4 (N4482, N4464, N3289, N3399, N1171);
not NOT1 (N4483, N4482);
xor XOR2 (N4484, N4463, N406);
nor NOR2 (N4485, N4480, N3303);
xor XOR2 (N4486, N4472, N3458);
buf BUF1 (N4487, N4483);
xor XOR2 (N4488, N4481, N3653);
nor NOR4 (N4489, N4487, N597, N726, N1909);
buf BUF1 (N4490, N4476);
or OR4 (N4491, N4490, N2736, N4373, N3197);
nand NAND2 (N4492, N4478, N3875);
or OR3 (N4493, N4489, N4047, N2279);
and AND4 (N4494, N4486, N826, N3520, N1803);
nor NOR4 (N4495, N4474, N1406, N2469, N3427);
nor NOR2 (N4496, N4494, N3677);
or OR3 (N4497, N4491, N1722, N1278);
nor NOR4 (N4498, N4488, N4359, N98, N2276);
nand NAND3 (N4499, N4470, N1686, N3416);
or OR4 (N4500, N4484, N2559, N4016, N3284);
or OR3 (N4501, N4499, N2103, N888);
nor NOR3 (N4502, N4492, N3945, N2872);
nor NOR3 (N4503, N4479, N600, N4255);
buf BUF1 (N4504, N4503);
and AND3 (N4505, N4498, N3207, N4424);
xor XOR2 (N4506, N4493, N1031);
buf BUF1 (N4507, N4504);
or OR3 (N4508, N4497, N3629, N3536);
or OR2 (N4509, N4485, N3066);
or OR3 (N4510, N4496, N2770, N3561);
nor NOR4 (N4511, N4500, N1000, N2414, N572);
not NOT1 (N4512, N4508);
xor XOR2 (N4513, N4502, N1687);
nor NOR3 (N4514, N4505, N4003, N3603);
and AND3 (N4515, N4501, N639, N565);
and AND2 (N4516, N4514, N3279);
nor NOR2 (N4517, N4515, N2957);
or OR3 (N4518, N4513, N4116, N3087);
nor NOR2 (N4519, N4517, N1746);
nor NOR3 (N4520, N4509, N901, N2913);
xor XOR2 (N4521, N4520, N3492);
xor XOR2 (N4522, N4521, N3837);
xor XOR2 (N4523, N4519, N3617);
xor XOR2 (N4524, N4510, N788);
xor XOR2 (N4525, N4512, N4441);
buf BUF1 (N4526, N4524);
xor XOR2 (N4527, N4523, N2445);
buf BUF1 (N4528, N4527);
buf BUF1 (N4529, N4522);
buf BUF1 (N4530, N4511);
xor XOR2 (N4531, N4528, N3992);
or OR4 (N4532, N4507, N224, N3636, N234);
or OR3 (N4533, N4530, N1690, N313);
and AND3 (N4534, N4526, N3026, N4372);
buf BUF1 (N4535, N4533);
and AND3 (N4536, N4518, N1716, N3326);
not NOT1 (N4537, N4529);
buf BUF1 (N4538, N4537);
nand NAND4 (N4539, N4531, N3870, N1035, N435);
or OR3 (N4540, N4525, N3187, N3967);
buf BUF1 (N4541, N4536);
buf BUF1 (N4542, N4532);
not NOT1 (N4543, N4516);
nor NOR4 (N4544, N4535, N720, N2742, N1463);
xor XOR2 (N4545, N4542, N76);
buf BUF1 (N4546, N4539);
nor NOR3 (N4547, N4541, N2215, N2313);
not NOT1 (N4548, N4540);
buf BUF1 (N4549, N4534);
buf BUF1 (N4550, N4548);
and AND4 (N4551, N4506, N1354, N850, N1049);
nand NAND3 (N4552, N4551, N469, N1190);
or OR3 (N4553, N4544, N2086, N161);
nand NAND4 (N4554, N4546, N1178, N4271, N4200);
xor XOR2 (N4555, N4543, N4434);
or OR4 (N4556, N4552, N2037, N3885, N3759);
or OR4 (N4557, N4550, N609, N3085, N3091);
and AND3 (N4558, N4554, N804, N3826);
nor NOR2 (N4559, N4555, N2776);
and AND3 (N4560, N4545, N3248, N1912);
buf BUF1 (N4561, N4495);
nand NAND3 (N4562, N4549, N370, N1293);
buf BUF1 (N4563, N4559);
xor XOR2 (N4564, N4563, N2455);
nand NAND3 (N4565, N4557, N3649, N2053);
not NOT1 (N4566, N4561);
nor NOR2 (N4567, N4566, N199);
or OR2 (N4568, N4565, N1980);
buf BUF1 (N4569, N4568);
or OR2 (N4570, N4547, N3123);
buf BUF1 (N4571, N4569);
not NOT1 (N4572, N4556);
not NOT1 (N4573, N4564);
not NOT1 (N4574, N4560);
and AND3 (N4575, N4538, N487, N3839);
and AND3 (N4576, N4558, N4139, N2255);
buf BUF1 (N4577, N4574);
nor NOR4 (N4578, N4571, N1452, N3470, N3229);
xor XOR2 (N4579, N4567, N2814);
or OR4 (N4580, N4573, N2463, N683, N3220);
or OR3 (N4581, N4553, N3105, N1362);
and AND4 (N4582, N4579, N28, N2754, N1644);
and AND2 (N4583, N4577, N3547);
not NOT1 (N4584, N4576);
and AND4 (N4585, N4578, N3719, N1565, N271);
xor XOR2 (N4586, N4583, N2524);
nand NAND3 (N4587, N4575, N3992, N1503);
or OR4 (N4588, N4586, N4041, N1328, N1208);
nand NAND2 (N4589, N4572, N3818);
buf BUF1 (N4590, N4581);
nor NOR3 (N4591, N4570, N2492, N2971);
not NOT1 (N4592, N4580);
nor NOR4 (N4593, N4589, N4029, N304, N2594);
xor XOR2 (N4594, N4591, N2724);
not NOT1 (N4595, N4584);
not NOT1 (N4596, N4595);
xor XOR2 (N4597, N4562, N3147);
nand NAND2 (N4598, N4593, N1519);
nor NOR4 (N4599, N4596, N352, N2232, N2940);
not NOT1 (N4600, N4594);
nor NOR4 (N4601, N4597, N4445, N1119, N4151);
xor XOR2 (N4602, N4582, N4174);
buf BUF1 (N4603, N4588);
xor XOR2 (N4604, N4598, N4430);
and AND2 (N4605, N4602, N1104);
not NOT1 (N4606, N4600);
and AND3 (N4607, N4592, N3420, N214);
nand NAND2 (N4608, N4603, N4147);
or OR3 (N4609, N4601, N594, N4344);
and AND2 (N4610, N4585, N200);
nand NAND3 (N4611, N4607, N4295, N772);
or OR4 (N4612, N4608, N1542, N3455, N1073);
and AND2 (N4613, N4587, N3081);
xor XOR2 (N4614, N4605, N4347);
xor XOR2 (N4615, N4612, N173);
nor NOR2 (N4616, N4609, N4173);
and AND2 (N4617, N4599, N1798);
or OR4 (N4618, N4617, N2258, N3116, N732);
or OR2 (N4619, N4606, N4385);
nand NAND3 (N4620, N4613, N1757, N4003);
and AND4 (N4621, N4611, N298, N1368, N3059);
xor XOR2 (N4622, N4616, N2198);
or OR3 (N4623, N4614, N593, N2900);
not NOT1 (N4624, N4622);
nor NOR2 (N4625, N4624, N2648);
or OR3 (N4626, N4618, N309, N4463);
nand NAND4 (N4627, N4621, N4071, N1765, N4051);
nor NOR2 (N4628, N4620, N4069);
and AND3 (N4629, N4619, N3234, N2757);
xor XOR2 (N4630, N4610, N936);
not NOT1 (N4631, N4627);
or OR3 (N4632, N4626, N4032, N2337);
buf BUF1 (N4633, N4625);
and AND4 (N4634, N4633, N3530, N2146, N2195);
or OR3 (N4635, N4623, N2545, N951);
not NOT1 (N4636, N4629);
not NOT1 (N4637, N4634);
nor NOR2 (N4638, N4631, N358);
or OR4 (N4639, N4615, N3342, N2574, N2552);
xor XOR2 (N4640, N4590, N3709);
xor XOR2 (N4641, N4604, N4195);
not NOT1 (N4642, N4641);
not NOT1 (N4643, N4637);
or OR4 (N4644, N4643, N1541, N256, N3412);
buf BUF1 (N4645, N4632);
nor NOR3 (N4646, N4642, N2822, N2452);
buf BUF1 (N4647, N4644);
nor NOR3 (N4648, N4645, N4134, N2943);
nor NOR3 (N4649, N4646, N3261, N3860);
xor XOR2 (N4650, N4635, N2453);
nand NAND3 (N4651, N4640, N2121, N2360);
and AND2 (N4652, N4638, N1601);
nor NOR3 (N4653, N4649, N3435, N758);
not NOT1 (N4654, N4652);
nor NOR4 (N4655, N4630, N4094, N4464, N1777);
not NOT1 (N4656, N4636);
or OR4 (N4657, N4651, N2290, N95, N1053);
nand NAND4 (N4658, N4654, N1761, N2272, N925);
not NOT1 (N4659, N4650);
or OR4 (N4660, N4658, N298, N3910, N4243);
nor NOR2 (N4661, N4660, N2432);
nor NOR3 (N4662, N4639, N1991, N3909);
nand NAND4 (N4663, N4656, N1191, N4377, N1064);
and AND3 (N4664, N4662, N2921, N3789);
not NOT1 (N4665, N4661);
or OR2 (N4666, N4647, N1371);
not NOT1 (N4667, N4648);
not NOT1 (N4668, N4657);
buf BUF1 (N4669, N4664);
nand NAND2 (N4670, N4659, N2349);
and AND2 (N4671, N4667, N3492);
nor NOR4 (N4672, N4665, N4365, N2463, N1674);
nor NOR2 (N4673, N4670, N4413);
nand NAND2 (N4674, N4663, N664);
and AND2 (N4675, N4673, N4122);
nand NAND3 (N4676, N4675, N2994, N4150);
not NOT1 (N4677, N4674);
nor NOR2 (N4678, N4676, N3887);
buf BUF1 (N4679, N4653);
or OR2 (N4680, N4628, N2995);
xor XOR2 (N4681, N4680, N4520);
and AND4 (N4682, N4655, N1740, N2441, N841);
nor NOR3 (N4683, N4668, N1188, N2508);
nor NOR2 (N4684, N4677, N141);
not NOT1 (N4685, N4672);
or OR4 (N4686, N4681, N1396, N1014, N2192);
nor NOR3 (N4687, N4684, N3341, N160);
or OR4 (N4688, N4687, N1277, N1618, N51);
xor XOR2 (N4689, N4688, N3211);
xor XOR2 (N4690, N4689, N2643);
buf BUF1 (N4691, N4666);
xor XOR2 (N4692, N4671, N2042);
not NOT1 (N4693, N4683);
buf BUF1 (N4694, N4690);
nand NAND2 (N4695, N4686, N180);
xor XOR2 (N4696, N4682, N3101);
nor NOR3 (N4697, N4696, N1326, N2829);
nor NOR3 (N4698, N4679, N2301, N1514);
nor NOR3 (N4699, N4695, N49, N3237);
buf BUF1 (N4700, N4697);
buf BUF1 (N4701, N4692);
nand NAND4 (N4702, N4678, N4118, N1835, N3515);
xor XOR2 (N4703, N4669, N3453);
not NOT1 (N4704, N4685);
xor XOR2 (N4705, N4704, N2685);
buf BUF1 (N4706, N4694);
xor XOR2 (N4707, N4705, N3153);
and AND3 (N4708, N4701, N4059, N1640);
nand NAND2 (N4709, N4706, N1920);
buf BUF1 (N4710, N4709);
buf BUF1 (N4711, N4700);
and AND4 (N4712, N4710, N2156, N508, N817);
nor NOR2 (N4713, N4698, N2693);
buf BUF1 (N4714, N4708);
nor NOR3 (N4715, N4693, N822, N1425);
xor XOR2 (N4716, N4707, N2835);
buf BUF1 (N4717, N4716);
nand NAND2 (N4718, N4712, N3760);
nand NAND2 (N4719, N4717, N3605);
not NOT1 (N4720, N4703);
nand NAND2 (N4721, N4715, N2432);
xor XOR2 (N4722, N4718, N3997);
or OR4 (N4723, N4699, N1348, N1026, N3639);
not NOT1 (N4724, N4714);
nor NOR4 (N4725, N4702, N1147, N2082, N709);
nand NAND4 (N4726, N4720, N3343, N4175, N3191);
nand NAND4 (N4727, N4691, N2340, N1951, N3818);
xor XOR2 (N4728, N4723, N3422);
not NOT1 (N4729, N4726);
and AND2 (N4730, N4713, N3194);
nand NAND4 (N4731, N4729, N3161, N3505, N3338);
and AND2 (N4732, N4722, N4132);
xor XOR2 (N4733, N4721, N4730);
nand NAND2 (N4734, N1216, N9);
or OR3 (N4735, N4719, N4339, N1448);
not NOT1 (N4736, N4725);
nor NOR3 (N4737, N4732, N517, N1103);
buf BUF1 (N4738, N4736);
nor NOR2 (N4739, N4733, N2503);
nor NOR3 (N4740, N4734, N323, N4247);
xor XOR2 (N4741, N4739, N3903);
or OR2 (N4742, N4741, N3329);
buf BUF1 (N4743, N4742);
buf BUF1 (N4744, N4728);
xor XOR2 (N4745, N4744, N4212);
and AND4 (N4746, N4727, N1252, N3894, N3387);
and AND2 (N4747, N4731, N956);
not NOT1 (N4748, N4745);
not NOT1 (N4749, N4740);
nand NAND3 (N4750, N4749, N3112, N1564);
not NOT1 (N4751, N4743);
not NOT1 (N4752, N4738);
xor XOR2 (N4753, N4750, N3328);
or OR2 (N4754, N4724, N2300);
xor XOR2 (N4755, N4747, N436);
nor NOR4 (N4756, N4751, N4247, N2272, N38);
nor NOR3 (N4757, N4735, N759, N1031);
xor XOR2 (N4758, N4711, N4060);
nor NOR3 (N4759, N4754, N1415, N869);
nor NOR4 (N4760, N4753, N2110, N1782, N255);
xor XOR2 (N4761, N4760, N3560);
xor XOR2 (N4762, N4756, N1347);
and AND3 (N4763, N4761, N326, N693);
buf BUF1 (N4764, N4758);
buf BUF1 (N4765, N4762);
nor NOR3 (N4766, N4765, N3573, N4708);
xor XOR2 (N4767, N4757, N2755);
nand NAND2 (N4768, N4752, N4551);
and AND2 (N4769, N4737, N3323);
not NOT1 (N4770, N4767);
buf BUF1 (N4771, N4755);
nor NOR2 (N4772, N4748, N1447);
buf BUF1 (N4773, N4769);
not NOT1 (N4774, N4766);
or OR4 (N4775, N4771, N1506, N1357, N2507);
and AND3 (N4776, N4759, N4232, N4740);
and AND3 (N4777, N4768, N4185, N989);
or OR4 (N4778, N4775, N3852, N4152, N3967);
nor NOR4 (N4779, N4778, N4693, N2619, N3507);
not NOT1 (N4780, N4764);
or OR4 (N4781, N4774, N3253, N1364, N1950);
and AND4 (N4782, N4777, N3673, N3282, N3097);
not NOT1 (N4783, N4763);
or OR4 (N4784, N4780, N1221, N590, N3278);
not NOT1 (N4785, N4776);
xor XOR2 (N4786, N4784, N1403);
nand NAND3 (N4787, N4773, N2007, N1257);
xor XOR2 (N4788, N4779, N3598);
buf BUF1 (N4789, N4781);
not NOT1 (N4790, N4785);
or OR4 (N4791, N4746, N2133, N3035, N4608);
buf BUF1 (N4792, N4790);
and AND2 (N4793, N4789, N2768);
nand NAND3 (N4794, N4783, N2810, N2752);
buf BUF1 (N4795, N4770);
and AND4 (N4796, N4791, N4344, N2262, N1353);
nor NOR2 (N4797, N4782, N3850);
not NOT1 (N4798, N4796);
xor XOR2 (N4799, N4788, N2295);
nand NAND4 (N4800, N4792, N4421, N4566, N3348);
not NOT1 (N4801, N4800);
and AND2 (N4802, N4798, N4587);
nand NAND4 (N4803, N4787, N455, N3089, N2049);
and AND2 (N4804, N4795, N2989);
not NOT1 (N4805, N4794);
not NOT1 (N4806, N4786);
and AND4 (N4807, N4797, N2751, N96, N4677);
not NOT1 (N4808, N4807);
nor NOR4 (N4809, N4772, N1905, N2043, N2328);
or OR3 (N4810, N4805, N1073, N3875);
not NOT1 (N4811, N4808);
nand NAND3 (N4812, N4806, N3040, N2050);
nor NOR4 (N4813, N4793, N4415, N3160, N3592);
nand NAND2 (N4814, N4801, N506);
xor XOR2 (N4815, N4811, N4790);
nor NOR3 (N4816, N4804, N2771, N1415);
nor NOR3 (N4817, N4813, N902, N3797);
xor XOR2 (N4818, N4817, N2626);
buf BUF1 (N4819, N4816);
or OR4 (N4820, N4815, N4140, N3554, N1677);
not NOT1 (N4821, N4812);
buf BUF1 (N4822, N4821);
nor NOR2 (N4823, N4822, N3556);
not NOT1 (N4824, N4814);
or OR2 (N4825, N4810, N4635);
nor NOR2 (N4826, N4802, N879);
nor NOR4 (N4827, N4825, N4324, N2228, N3358);
buf BUF1 (N4828, N4823);
nor NOR4 (N4829, N4824, N4598, N2417, N213);
buf BUF1 (N4830, N4826);
nor NOR2 (N4831, N4828, N1707);
nand NAND2 (N4832, N4819, N17);
or OR3 (N4833, N4818, N2148, N3388);
xor XOR2 (N4834, N4833, N4562);
xor XOR2 (N4835, N4809, N1782);
or OR3 (N4836, N4835, N3142, N875);
not NOT1 (N4837, N4829);
xor XOR2 (N4838, N4836, N2701);
not NOT1 (N4839, N4799);
not NOT1 (N4840, N4827);
nand NAND2 (N4841, N4820, N25);
buf BUF1 (N4842, N4832);
or OR3 (N4843, N4830, N3345, N849);
and AND4 (N4844, N4843, N1283, N1508, N4296);
not NOT1 (N4845, N4831);
buf BUF1 (N4846, N4840);
nor NOR2 (N4847, N4841, N2320);
xor XOR2 (N4848, N4846, N3988);
not NOT1 (N4849, N4848);
and AND2 (N4850, N4839, N4829);
xor XOR2 (N4851, N4834, N2787);
nor NOR4 (N4852, N4837, N1433, N2329, N567);
nand NAND4 (N4853, N4847, N3564, N4536, N1352);
or OR3 (N4854, N4838, N3492, N757);
nand NAND3 (N4855, N4853, N4740, N1586);
and AND3 (N4856, N4854, N1073, N2110);
xor XOR2 (N4857, N4842, N4794);
xor XOR2 (N4858, N4857, N3398);
not NOT1 (N4859, N4850);
not NOT1 (N4860, N4859);
and AND2 (N4861, N4855, N1565);
not NOT1 (N4862, N4858);
nand NAND3 (N4863, N4844, N3510, N3270);
nand NAND4 (N4864, N4861, N1187, N130, N3041);
xor XOR2 (N4865, N4864, N2044);
nand NAND2 (N4866, N4849, N3331);
not NOT1 (N4867, N4860);
nand NAND3 (N4868, N4863, N4688, N1382);
and AND2 (N4869, N4868, N2686);
xor XOR2 (N4870, N4803, N4731);
buf BUF1 (N4871, N4852);
not NOT1 (N4872, N4851);
buf BUF1 (N4873, N4870);
buf BUF1 (N4874, N4871);
and AND3 (N4875, N4869, N2211, N4798);
not NOT1 (N4876, N4856);
and AND2 (N4877, N4874, N2161);
buf BUF1 (N4878, N4845);
nor NOR3 (N4879, N4876, N602, N137);
or OR3 (N4880, N4872, N4873, N3565);
and AND2 (N4881, N2072, N3210);
and AND2 (N4882, N4877, N3354);
or OR2 (N4883, N4881, N3162);
buf BUF1 (N4884, N4875);
nand NAND3 (N4885, N4866, N1350, N500);
and AND2 (N4886, N4880, N4158);
nor NOR4 (N4887, N4883, N443, N2308, N1040);
buf BUF1 (N4888, N4884);
and AND3 (N4889, N4865, N4066, N2934);
xor XOR2 (N4890, N4878, N1055);
buf BUF1 (N4891, N4889);
nor NOR4 (N4892, N4887, N265, N85, N3503);
or OR2 (N4893, N4891, N4644);
nor NOR3 (N4894, N4893, N2692, N4232);
nor NOR2 (N4895, N4867, N3570);
nor NOR2 (N4896, N4886, N15);
buf BUF1 (N4897, N4862);
buf BUF1 (N4898, N4896);
or OR4 (N4899, N4888, N4292, N3359, N3886);
buf BUF1 (N4900, N4898);
nor NOR3 (N4901, N4894, N4663, N619);
not NOT1 (N4902, N4879);
not NOT1 (N4903, N4897);
and AND3 (N4904, N4903, N2163, N4185);
not NOT1 (N4905, N4904);
and AND2 (N4906, N4900, N4053);
buf BUF1 (N4907, N4899);
nor NOR4 (N4908, N4906, N2163, N194, N1186);
nand NAND3 (N4909, N4902, N3837, N3965);
or OR4 (N4910, N4882, N1108, N3494, N2745);
xor XOR2 (N4911, N4905, N3533);
nor NOR3 (N4912, N4885, N802, N1757);
nand NAND3 (N4913, N4890, N930, N3889);
not NOT1 (N4914, N4909);
and AND3 (N4915, N4908, N834, N4214);
or OR2 (N4916, N4901, N1698);
xor XOR2 (N4917, N4907, N4641);
xor XOR2 (N4918, N4895, N3811);
xor XOR2 (N4919, N4892, N4865);
nand NAND4 (N4920, N4917, N1579, N854, N3148);
nor NOR3 (N4921, N4910, N637, N49);
and AND2 (N4922, N4911, N3310);
and AND4 (N4923, N4914, N633, N358, N711);
not NOT1 (N4924, N4920);
xor XOR2 (N4925, N4921, N1944);
not NOT1 (N4926, N4915);
nand NAND3 (N4927, N4918, N541, N3250);
and AND4 (N4928, N4922, N4804, N334, N300);
or OR4 (N4929, N4924, N4143, N2424, N1884);
nand NAND3 (N4930, N4919, N347, N542);
or OR3 (N4931, N4927, N2619, N648);
xor XOR2 (N4932, N4928, N3905);
and AND4 (N4933, N4923, N3996, N1384, N2233);
nand NAND2 (N4934, N4932, N3168);
buf BUF1 (N4935, N4931);
and AND4 (N4936, N4926, N4562, N2053, N2452);
nand NAND4 (N4937, N4916, N4167, N744, N4294);
or OR2 (N4938, N4935, N63);
and AND3 (N4939, N4938, N1259, N1716);
not NOT1 (N4940, N4939);
nand NAND2 (N4941, N4929, N712);
buf BUF1 (N4942, N4940);
nor NOR4 (N4943, N4936, N1817, N491, N510);
not NOT1 (N4944, N4943);
nand NAND2 (N4945, N4912, N733);
or OR2 (N4946, N4934, N3855);
xor XOR2 (N4947, N4944, N3427);
or OR2 (N4948, N4933, N4587);
nor NOR4 (N4949, N4945, N1955, N2995, N2019);
xor XOR2 (N4950, N4946, N1850);
and AND4 (N4951, N4937, N1357, N1195, N1092);
or OR3 (N4952, N4947, N2625, N816);
nor NOR4 (N4953, N4951, N3581, N4743, N3500);
or OR3 (N4954, N4925, N1752, N3443);
buf BUF1 (N4955, N4941);
buf BUF1 (N4956, N4955);
nor NOR4 (N4957, N4949, N2114, N4769, N2914);
or OR2 (N4958, N4954, N3068);
nand NAND4 (N4959, N4957, N4006, N200, N1458);
nand NAND2 (N4960, N4942, N994);
or OR4 (N4961, N4960, N3008, N449, N4073);
or OR4 (N4962, N4959, N1181, N567, N2575);
not NOT1 (N4963, N4958);
xor XOR2 (N4964, N4963, N4774);
xor XOR2 (N4965, N4950, N495);
xor XOR2 (N4966, N4953, N4772);
not NOT1 (N4967, N4948);
buf BUF1 (N4968, N4913);
not NOT1 (N4969, N4967);
not NOT1 (N4970, N4969);
not NOT1 (N4971, N4952);
nor NOR4 (N4972, N4966, N1448, N4679, N4380);
and AND3 (N4973, N4970, N1746, N1996);
or OR3 (N4974, N4930, N928, N1886);
nand NAND4 (N4975, N4968, N1170, N2087, N255);
xor XOR2 (N4976, N4975, N836);
not NOT1 (N4977, N4964);
xor XOR2 (N4978, N4965, N1283);
or OR2 (N4979, N4962, N3311);
or OR3 (N4980, N4961, N587, N3728);
nor NOR2 (N4981, N4956, N3485);
not NOT1 (N4982, N4981);
nor NOR3 (N4983, N4976, N1008, N3097);
nand NAND3 (N4984, N4977, N348, N3331);
nand NAND2 (N4985, N4984, N1686);
buf BUF1 (N4986, N4971);
nor NOR3 (N4987, N4974, N3900, N1574);
nand NAND3 (N4988, N4973, N1897, N3332);
and AND3 (N4989, N4982, N1117, N3611);
not NOT1 (N4990, N4978);
nor NOR4 (N4991, N4985, N790, N3311, N3752);
nor NOR3 (N4992, N4991, N4481, N618);
nand NAND2 (N4993, N4979, N2988);
buf BUF1 (N4994, N4993);
not NOT1 (N4995, N4989);
nor NOR4 (N4996, N4990, N4683, N1549, N4880);
not NOT1 (N4997, N4987);
or OR2 (N4998, N4992, N2772);
and AND2 (N4999, N4994, N3499);
xor XOR2 (N5000, N4998, N3428);
buf BUF1 (N5001, N4972);
nand NAND2 (N5002, N4980, N247);
xor XOR2 (N5003, N4999, N829);
buf BUF1 (N5004, N4996);
buf BUF1 (N5005, N4997);
xor XOR2 (N5006, N4983, N2140);
not NOT1 (N5007, N5004);
not NOT1 (N5008, N5001);
nand NAND3 (N5009, N4986, N725, N334);
or OR3 (N5010, N5002, N4373, N358);
nand NAND4 (N5011, N5005, N1595, N3706, N2518);
buf BUF1 (N5012, N5008);
not NOT1 (N5013, N5011);
or OR4 (N5014, N5006, N1004, N4935, N3829);
xor XOR2 (N5015, N5010, N1296);
or OR4 (N5016, N5000, N2354, N2739, N290);
not NOT1 (N5017, N5003);
buf BUF1 (N5018, N5013);
buf BUF1 (N5019, N5018);
buf BUF1 (N5020, N4995);
buf BUF1 (N5021, N5012);
xor XOR2 (N5022, N4988, N5004);
not NOT1 (N5023, N5017);
xor XOR2 (N5024, N5021, N2976);
not NOT1 (N5025, N5009);
buf BUF1 (N5026, N5022);
not NOT1 (N5027, N5020);
nor NOR4 (N5028, N5014, N2783, N4749, N2267);
not NOT1 (N5029, N5025);
nor NOR3 (N5030, N5019, N4800, N955);
and AND4 (N5031, N5029, N4040, N3519, N3853);
and AND4 (N5032, N5015, N3143, N4190, N4237);
nor NOR2 (N5033, N5030, N4082);
buf BUF1 (N5034, N5032);
or OR4 (N5035, N5007, N3772, N1799, N1848);
nand NAND4 (N5036, N5031, N414, N2702, N3326);
buf BUF1 (N5037, N5016);
buf BUF1 (N5038, N5033);
and AND3 (N5039, N5037, N186, N1014);
buf BUF1 (N5040, N5039);
or OR4 (N5041, N5023, N2792, N1737, N1772);
not NOT1 (N5042, N5040);
buf BUF1 (N5043, N5026);
not NOT1 (N5044, N5043);
nand NAND3 (N5045, N5042, N639, N2140);
nor NOR2 (N5046, N5045, N3963);
buf BUF1 (N5047, N5034);
nand NAND3 (N5048, N5041, N861, N2152);
buf BUF1 (N5049, N5038);
or OR4 (N5050, N5049, N96, N2413, N4182);
not NOT1 (N5051, N5048);
buf BUF1 (N5052, N5047);
or OR2 (N5053, N5052, N2186);
nand NAND2 (N5054, N5028, N1214);
nor NOR4 (N5055, N5024, N1856, N3813, N4034);
nor NOR4 (N5056, N5055, N3581, N3407, N4077);
not NOT1 (N5057, N5027);
nand NAND4 (N5058, N5035, N136, N2254, N4485);
nor NOR4 (N5059, N5046, N2039, N2897, N2413);
buf BUF1 (N5060, N5053);
and AND3 (N5061, N5054, N3946, N1402);
xor XOR2 (N5062, N5036, N4239);
buf BUF1 (N5063, N5056);
nand NAND4 (N5064, N5050, N3596, N4078, N4856);
buf BUF1 (N5065, N5057);
nand NAND2 (N5066, N5059, N4874);
xor XOR2 (N5067, N5064, N4465);
not NOT1 (N5068, N5065);
xor XOR2 (N5069, N5063, N1220);
buf BUF1 (N5070, N5062);
and AND3 (N5071, N5058, N716, N4531);
not NOT1 (N5072, N5060);
buf BUF1 (N5073, N5044);
buf BUF1 (N5074, N5067);
xor XOR2 (N5075, N5066, N4994);
nand NAND2 (N5076, N5051, N2697);
nor NOR2 (N5077, N5072, N2244);
nand NAND2 (N5078, N5076, N4378);
and AND3 (N5079, N5071, N2654, N3708);
nand NAND4 (N5080, N5079, N1338, N5029, N3441);
and AND2 (N5081, N5075, N4249);
xor XOR2 (N5082, N5080, N2385);
buf BUF1 (N5083, N5069);
or OR2 (N5084, N5083, N777);
buf BUF1 (N5085, N5068);
and AND3 (N5086, N5081, N4333, N1702);
buf BUF1 (N5087, N5070);
buf BUF1 (N5088, N5087);
and AND3 (N5089, N5077, N263, N2647);
nor NOR2 (N5090, N5085, N266);
nand NAND4 (N5091, N5090, N667, N1929, N4280);
nor NOR3 (N5092, N5082, N3341, N4574);
nor NOR2 (N5093, N5089, N2484);
xor XOR2 (N5094, N5084, N1340);
xor XOR2 (N5095, N5061, N2554);
nand NAND2 (N5096, N5074, N1409);
xor XOR2 (N5097, N5095, N3817);
nor NOR2 (N5098, N5094, N3711);
or OR2 (N5099, N5078, N4191);
not NOT1 (N5100, N5073);
nor NOR3 (N5101, N5093, N2328, N2508);
nor NOR4 (N5102, N5092, N4392, N469, N4421);
buf BUF1 (N5103, N5097);
buf BUF1 (N5104, N5098);
xor XOR2 (N5105, N5086, N2532);
not NOT1 (N5106, N5102);
or OR4 (N5107, N5103, N674, N1852, N3449);
nor NOR4 (N5108, N5088, N2384, N4505, N2618);
nor NOR2 (N5109, N5104, N804);
or OR3 (N5110, N5091, N1192, N1805);
nand NAND4 (N5111, N5106, N4472, N215, N1096);
nor NOR2 (N5112, N5111, N101);
nand NAND4 (N5113, N5112, N5087, N2265, N2361);
or OR3 (N5114, N5113, N424, N3425);
not NOT1 (N5115, N5101);
xor XOR2 (N5116, N5110, N1471);
nor NOR2 (N5117, N5109, N3546);
nor NOR4 (N5118, N5107, N4983, N1498, N607);
and AND3 (N5119, N5099, N3625, N762);
and AND3 (N5120, N5105, N4517, N201);
not NOT1 (N5121, N5116);
or OR2 (N5122, N5108, N3386);
not NOT1 (N5123, N5121);
xor XOR2 (N5124, N5118, N3941);
and AND4 (N5125, N5122, N1705, N1248, N1285);
xor XOR2 (N5126, N5123, N2831);
nor NOR2 (N5127, N5125, N3493);
buf BUF1 (N5128, N5127);
nor NOR3 (N5129, N5115, N1594, N2580);
not NOT1 (N5130, N5100);
and AND4 (N5131, N5124, N496, N1100, N2392);
xor XOR2 (N5132, N5126, N3041);
nand NAND4 (N5133, N5131, N1200, N2548, N4780);
not NOT1 (N5134, N5114);
not NOT1 (N5135, N5120);
xor XOR2 (N5136, N5132, N4486);
not NOT1 (N5137, N5136);
not NOT1 (N5138, N5137);
and AND2 (N5139, N5129, N4956);
and AND3 (N5140, N5130, N3319, N1039);
xor XOR2 (N5141, N5117, N4878);
and AND3 (N5142, N5141, N4044, N2528);
or OR3 (N5143, N5133, N2715, N3006);
or OR4 (N5144, N5134, N4103, N2348, N1264);
not NOT1 (N5145, N5138);
buf BUF1 (N5146, N5128);
and AND4 (N5147, N5142, N4007, N97, N4665);
or OR3 (N5148, N5140, N143, N2838);
buf BUF1 (N5149, N5139);
buf BUF1 (N5150, N5144);
nor NOR4 (N5151, N5146, N189, N185, N3707);
and AND4 (N5152, N5119, N1415, N500, N3828);
nand NAND2 (N5153, N5149, N2477);
or OR2 (N5154, N5152, N685);
nand NAND4 (N5155, N5150, N3964, N1658, N792);
buf BUF1 (N5156, N5096);
xor XOR2 (N5157, N5147, N3029);
nor NOR2 (N5158, N5154, N425);
or OR3 (N5159, N5148, N3285, N1260);
xor XOR2 (N5160, N5158, N37);
nor NOR3 (N5161, N5155, N2183, N4083);
not NOT1 (N5162, N5156);
and AND2 (N5163, N5160, N2058);
nand NAND3 (N5164, N5151, N4713, N4186);
xor XOR2 (N5165, N5153, N2575);
nand NAND4 (N5166, N5161, N4188, N276, N1801);
and AND3 (N5167, N5165, N2718, N2659);
not NOT1 (N5168, N5157);
or OR2 (N5169, N5145, N2930);
xor XOR2 (N5170, N5169, N871);
xor XOR2 (N5171, N5166, N4489);
or OR2 (N5172, N5170, N1207);
buf BUF1 (N5173, N5135);
not NOT1 (N5174, N5159);
xor XOR2 (N5175, N5143, N2086);
xor XOR2 (N5176, N5167, N1583);
not NOT1 (N5177, N5171);
xor XOR2 (N5178, N5163, N2752);
not NOT1 (N5179, N5164);
xor XOR2 (N5180, N5177, N1678);
or OR3 (N5181, N5176, N3660, N4061);
or OR3 (N5182, N5180, N1773, N4661);
nand NAND4 (N5183, N5162, N4875, N3152, N2578);
or OR4 (N5184, N5173, N5154, N2137, N1328);
not NOT1 (N5185, N5179);
buf BUF1 (N5186, N5185);
or OR3 (N5187, N5182, N233, N2403);
or OR3 (N5188, N5168, N3747, N3827);
nor NOR2 (N5189, N5184, N64);
buf BUF1 (N5190, N5175);
buf BUF1 (N5191, N5183);
or OR2 (N5192, N5186, N2175);
xor XOR2 (N5193, N5181, N4508);
and AND2 (N5194, N5191, N503);
xor XOR2 (N5195, N5178, N1283);
or OR4 (N5196, N5194, N2343, N2238, N1542);
buf BUF1 (N5197, N5174);
xor XOR2 (N5198, N5197, N3333);
xor XOR2 (N5199, N5188, N2495);
not NOT1 (N5200, N5192);
and AND4 (N5201, N5190, N3447, N3184, N770);
nand NAND2 (N5202, N5199, N3089);
or OR4 (N5203, N5172, N991, N242, N974);
and AND3 (N5204, N5203, N2601, N3974);
and AND2 (N5205, N5193, N5182);
nor NOR2 (N5206, N5205, N3478);
buf BUF1 (N5207, N5195);
not NOT1 (N5208, N5196);
buf BUF1 (N5209, N5187);
buf BUF1 (N5210, N5201);
not NOT1 (N5211, N5200);
or OR3 (N5212, N5198, N4230, N2);
buf BUF1 (N5213, N5206);
nand NAND4 (N5214, N5211, N4446, N2990, N1727);
not NOT1 (N5215, N5204);
nand NAND2 (N5216, N5202, N4229);
not NOT1 (N5217, N5209);
not NOT1 (N5218, N5213);
and AND2 (N5219, N5218, N5153);
or OR3 (N5220, N5214, N3383, N3581);
nor NOR4 (N5221, N5220, N2096, N2430, N3658);
xor XOR2 (N5222, N5215, N1479);
nand NAND3 (N5223, N5210, N747, N1098);
not NOT1 (N5224, N5219);
xor XOR2 (N5225, N5222, N4665);
and AND2 (N5226, N5221, N1543);
or OR3 (N5227, N5224, N3923, N2271);
nor NOR4 (N5228, N5226, N476, N4118, N3329);
or OR3 (N5229, N5217, N3783, N1220);
or OR2 (N5230, N5228, N4475);
nand NAND3 (N5231, N5230, N358, N2846);
nor NOR4 (N5232, N5208, N4463, N2525, N4086);
not NOT1 (N5233, N5223);
or OR4 (N5234, N5225, N842, N1432, N623);
or OR2 (N5235, N5212, N1117);
nand NAND4 (N5236, N5234, N2949, N2582, N2439);
xor XOR2 (N5237, N5229, N3498);
nand NAND2 (N5238, N5227, N2208);
not NOT1 (N5239, N5238);
xor XOR2 (N5240, N5235, N47);
buf BUF1 (N5241, N5231);
nor NOR2 (N5242, N5233, N2940);
not NOT1 (N5243, N5232);
buf BUF1 (N5244, N5207);
nor NOR4 (N5245, N5236, N1608, N2714, N2058);
nor NOR4 (N5246, N5244, N624, N3723, N674);
and AND3 (N5247, N5241, N1073, N3126);
or OR3 (N5248, N5189, N265, N4103);
xor XOR2 (N5249, N5248, N2424);
not NOT1 (N5250, N5242);
xor XOR2 (N5251, N5216, N1018);
nor NOR3 (N5252, N5246, N2612, N2636);
buf BUF1 (N5253, N5245);
or OR4 (N5254, N5243, N2028, N2484, N3580);
buf BUF1 (N5255, N5252);
nand NAND4 (N5256, N5251, N526, N1499, N3051);
nor NOR2 (N5257, N5247, N3664);
nand NAND2 (N5258, N5257, N4644);
xor XOR2 (N5259, N5254, N628);
xor XOR2 (N5260, N5256, N4327);
not NOT1 (N5261, N5258);
xor XOR2 (N5262, N5255, N2041);
xor XOR2 (N5263, N5240, N986);
or OR2 (N5264, N5239, N3977);
nor NOR2 (N5265, N5261, N2142);
nand NAND2 (N5266, N5237, N981);
nand NAND3 (N5267, N5250, N4318, N2224);
and AND4 (N5268, N5264, N498, N2148, N2721);
buf BUF1 (N5269, N5267);
buf BUF1 (N5270, N5265);
or OR4 (N5271, N5249, N2886, N1323, N4045);
nor NOR2 (N5272, N5271, N1269);
and AND4 (N5273, N5268, N3080, N3540, N3876);
not NOT1 (N5274, N5270);
xor XOR2 (N5275, N5272, N724);
buf BUF1 (N5276, N5274);
not NOT1 (N5277, N5260);
and AND4 (N5278, N5277, N955, N1004, N107);
buf BUF1 (N5279, N5278);
nand NAND4 (N5280, N5273, N3703, N1126, N2673);
nor NOR3 (N5281, N5263, N3912, N1466);
not NOT1 (N5282, N5276);
or OR2 (N5283, N5262, N4937);
nand NAND2 (N5284, N5259, N2032);
and AND4 (N5285, N5282, N1953, N513, N2379);
xor XOR2 (N5286, N5266, N1740);
xor XOR2 (N5287, N5286, N635);
nand NAND4 (N5288, N5281, N4412, N1776, N3754);
or OR2 (N5289, N5253, N3936);
not NOT1 (N5290, N5280);
nor NOR4 (N5291, N5289, N4124, N2686, N2904);
nor NOR4 (N5292, N5285, N3743, N3257, N2036);
and AND2 (N5293, N5279, N1082);
nor NOR4 (N5294, N5288, N2995, N3644, N3425);
nand NAND4 (N5295, N5290, N315, N4984, N3168);
nor NOR4 (N5296, N5287, N4752, N4226, N2762);
and AND4 (N5297, N5295, N3810, N3918, N373);
nor NOR3 (N5298, N5296, N4974, N626);
not NOT1 (N5299, N5284);
nor NOR4 (N5300, N5297, N1978, N3884, N2274);
buf BUF1 (N5301, N5291);
xor XOR2 (N5302, N5300, N4431);
xor XOR2 (N5303, N5301, N1416);
and AND3 (N5304, N5292, N2791, N2701);
and AND2 (N5305, N5275, N2482);
nor NOR3 (N5306, N5269, N4371, N110);
xor XOR2 (N5307, N5299, N3780);
nand NAND2 (N5308, N5293, N1306);
xor XOR2 (N5309, N5294, N3305);
nand NAND2 (N5310, N5309, N4003);
buf BUF1 (N5311, N5302);
not NOT1 (N5312, N5308);
buf BUF1 (N5313, N5298);
nand NAND4 (N5314, N5307, N4941, N1897, N2790);
or OR3 (N5315, N5311, N3552, N4151);
nand NAND3 (N5316, N5312, N2253, N2514);
nand NAND2 (N5317, N5310, N2388);
buf BUF1 (N5318, N5306);
or OR4 (N5319, N5304, N1025, N4361, N374);
not NOT1 (N5320, N5317);
buf BUF1 (N5321, N5283);
or OR2 (N5322, N5305, N4060);
and AND2 (N5323, N5303, N4476);
nand NAND4 (N5324, N5316, N2716, N565, N5019);
xor XOR2 (N5325, N5320, N3830);
nand NAND3 (N5326, N5325, N1314, N1859);
buf BUF1 (N5327, N5324);
or OR2 (N5328, N5313, N1809);
or OR2 (N5329, N5318, N636);
nand NAND2 (N5330, N5328, N3109);
xor XOR2 (N5331, N5323, N2541);
nor NOR2 (N5332, N5327, N1305);
buf BUF1 (N5333, N5332);
and AND3 (N5334, N5329, N3369, N4504);
and AND3 (N5335, N5319, N1046, N2413);
and AND4 (N5336, N5314, N2779, N3424, N1767);
buf BUF1 (N5337, N5333);
xor XOR2 (N5338, N5322, N406);
nand NAND3 (N5339, N5331, N4250, N1708);
buf BUF1 (N5340, N5335);
not NOT1 (N5341, N5336);
xor XOR2 (N5342, N5340, N5182);
and AND3 (N5343, N5337, N496, N1713);
not NOT1 (N5344, N5339);
or OR3 (N5345, N5338, N372, N3138);
nor NOR4 (N5346, N5326, N3130, N1996, N5086);
and AND3 (N5347, N5330, N1210, N1454);
and AND4 (N5348, N5341, N5209, N4729, N5256);
and AND4 (N5349, N5346, N4638, N1654, N1116);
or OR3 (N5350, N5347, N3746, N4493);
nor NOR3 (N5351, N5343, N35, N3946);
nor NOR2 (N5352, N5349, N4172);
or OR2 (N5353, N5351, N4010);
nor NOR4 (N5354, N5348, N641, N5004, N1221);
xor XOR2 (N5355, N5334, N477);
or OR3 (N5356, N5321, N2674, N4963);
and AND3 (N5357, N5355, N1433, N1234);
xor XOR2 (N5358, N5356, N4531);
nand NAND3 (N5359, N5315, N5033, N3922);
xor XOR2 (N5360, N5359, N5295);
or OR3 (N5361, N5360, N352, N2130);
not NOT1 (N5362, N5353);
and AND4 (N5363, N5352, N248, N3160, N3102);
and AND2 (N5364, N5361, N2780);
xor XOR2 (N5365, N5342, N5052);
nor NOR2 (N5366, N5364, N3795);
and AND3 (N5367, N5345, N4309, N2457);
xor XOR2 (N5368, N5367, N106);
not NOT1 (N5369, N5362);
xor XOR2 (N5370, N5368, N502);
or OR3 (N5371, N5354, N4664, N3805);
nand NAND3 (N5372, N5357, N5191, N2140);
xor XOR2 (N5373, N5370, N3653);
buf BUF1 (N5374, N5369);
nand NAND2 (N5375, N5371, N4511);
xor XOR2 (N5376, N5375, N875);
nand NAND2 (N5377, N5350, N3555);
buf BUF1 (N5378, N5374);
xor XOR2 (N5379, N5372, N386);
not NOT1 (N5380, N5378);
xor XOR2 (N5381, N5376, N2868);
nand NAND4 (N5382, N5363, N2502, N5375, N2772);
not NOT1 (N5383, N5344);
and AND4 (N5384, N5380, N637, N2589, N4358);
nor NOR3 (N5385, N5379, N3273, N2064);
or OR4 (N5386, N5373, N1113, N2818, N1434);
or OR3 (N5387, N5358, N1555, N3677);
and AND2 (N5388, N5365, N4860);
xor XOR2 (N5389, N5384, N4073);
not NOT1 (N5390, N5381);
or OR2 (N5391, N5377, N2931);
and AND3 (N5392, N5390, N3647, N851);
or OR3 (N5393, N5366, N2936, N5318);
not NOT1 (N5394, N5385);
nor NOR2 (N5395, N5394, N5146);
not NOT1 (N5396, N5388);
or OR2 (N5397, N5391, N5080);
not NOT1 (N5398, N5387);
and AND2 (N5399, N5389, N1836);
buf BUF1 (N5400, N5397);
buf BUF1 (N5401, N5383);
nor NOR2 (N5402, N5399, N2108);
xor XOR2 (N5403, N5395, N3750);
buf BUF1 (N5404, N5398);
or OR2 (N5405, N5400, N3167);
xor XOR2 (N5406, N5402, N3495);
not NOT1 (N5407, N5392);
nand NAND4 (N5408, N5396, N4213, N5137, N2600);
not NOT1 (N5409, N5405);
nand NAND3 (N5410, N5408, N542, N3875);
or OR3 (N5411, N5393, N3156, N698);
buf BUF1 (N5412, N5411);
not NOT1 (N5413, N5382);
nand NAND3 (N5414, N5404, N915, N5158);
not NOT1 (N5415, N5403);
xor XOR2 (N5416, N5410, N5305);
or OR2 (N5417, N5414, N1862);
or OR3 (N5418, N5386, N279, N5411);
xor XOR2 (N5419, N5401, N3533);
not NOT1 (N5420, N5409);
not NOT1 (N5421, N5417);
and AND2 (N5422, N5421, N4210);
not NOT1 (N5423, N5422);
buf BUF1 (N5424, N5412);
and AND2 (N5425, N5418, N3459);
xor XOR2 (N5426, N5425, N3411);
and AND4 (N5427, N5406, N1817, N2327, N3043);
nor NOR2 (N5428, N5424, N2934);
nor NOR4 (N5429, N5426, N2104, N2479, N2141);
or OR2 (N5430, N5413, N851);
not NOT1 (N5431, N5428);
nor NOR2 (N5432, N5431, N1322);
and AND2 (N5433, N5432, N1126);
buf BUF1 (N5434, N5433);
and AND3 (N5435, N5420, N4282, N5251);
nand NAND2 (N5436, N5429, N763);
xor XOR2 (N5437, N5435, N1342);
xor XOR2 (N5438, N5436, N1339);
not NOT1 (N5439, N5427);
or OR2 (N5440, N5419, N5386);
nand NAND4 (N5441, N5438, N3268, N2336, N2954);
nor NOR3 (N5442, N5415, N3329, N4830);
xor XOR2 (N5443, N5430, N3098);
nor NOR3 (N5444, N5423, N613, N4454);
nand NAND4 (N5445, N5434, N1863, N5428, N3800);
nor NOR3 (N5446, N5437, N3904, N4661);
xor XOR2 (N5447, N5441, N4870);
nor NOR4 (N5448, N5445, N340, N4431, N4387);
buf BUF1 (N5449, N5416);
nor NOR4 (N5450, N5444, N1683, N96, N293);
xor XOR2 (N5451, N5450, N4290);
buf BUF1 (N5452, N5443);
nor NOR2 (N5453, N5442, N4359);
nor NOR4 (N5454, N5439, N2668, N2885, N1023);
xor XOR2 (N5455, N5453, N350);
or OR2 (N5456, N5452, N1051);
and AND2 (N5457, N5446, N2593);
not NOT1 (N5458, N5451);
or OR4 (N5459, N5455, N1702, N4399, N5321);
or OR4 (N5460, N5407, N213, N4622, N1102);
not NOT1 (N5461, N5454);
not NOT1 (N5462, N5460);
nor NOR3 (N5463, N5458, N3979, N4152);
nor NOR3 (N5464, N5447, N4424, N3028);
nor NOR3 (N5465, N5461, N2791, N1398);
buf BUF1 (N5466, N5464);
xor XOR2 (N5467, N5465, N5352);
nand NAND4 (N5468, N5462, N21, N2130, N2065);
buf BUF1 (N5469, N5457);
xor XOR2 (N5470, N5449, N2065);
buf BUF1 (N5471, N5456);
and AND2 (N5472, N5466, N773);
xor XOR2 (N5473, N5459, N1096);
xor XOR2 (N5474, N5467, N1068);
buf BUF1 (N5475, N5473);
buf BUF1 (N5476, N5440);
buf BUF1 (N5477, N5476);
xor XOR2 (N5478, N5475, N2402);
xor XOR2 (N5479, N5470, N2775);
and AND3 (N5480, N5478, N3106, N3859);
and AND2 (N5481, N5463, N345);
or OR3 (N5482, N5480, N4619, N1485);
and AND3 (N5483, N5472, N403, N3399);
not NOT1 (N5484, N5474);
not NOT1 (N5485, N5477);
nand NAND4 (N5486, N5482, N1663, N5295, N1252);
nor NOR2 (N5487, N5479, N3987);
nand NAND4 (N5488, N5483, N4332, N282, N1717);
xor XOR2 (N5489, N5448, N1027);
and AND4 (N5490, N5486, N4715, N3300, N233);
or OR4 (N5491, N5490, N296, N3362, N5480);
not NOT1 (N5492, N5469);
not NOT1 (N5493, N5492);
buf BUF1 (N5494, N5481);
or OR2 (N5495, N5488, N3319);
not NOT1 (N5496, N5471);
and AND2 (N5497, N5484, N2172);
and AND2 (N5498, N5489, N1619);
not NOT1 (N5499, N5498);
not NOT1 (N5500, N5487);
nand NAND2 (N5501, N5491, N3085);
buf BUF1 (N5502, N5495);
and AND3 (N5503, N5499, N1652, N3391);
or OR2 (N5504, N5494, N992);
xor XOR2 (N5505, N5496, N1105);
or OR2 (N5506, N5468, N66);
xor XOR2 (N5507, N5500, N5492);
or OR2 (N5508, N5501, N972);
not NOT1 (N5509, N5502);
nor NOR3 (N5510, N5504, N4579, N1545);
or OR3 (N5511, N5507, N1952, N2155);
and AND4 (N5512, N5493, N4878, N1344, N4703);
or OR2 (N5513, N5505, N548);
xor XOR2 (N5514, N5508, N2891);
buf BUF1 (N5515, N5509);
xor XOR2 (N5516, N5515, N4705);
xor XOR2 (N5517, N5503, N832);
nand NAND4 (N5518, N5514, N1928, N4894, N4114);
nand NAND2 (N5519, N5512, N2948);
not NOT1 (N5520, N5510);
or OR2 (N5521, N5520, N4768);
not NOT1 (N5522, N5506);
or OR2 (N5523, N5516, N2288);
not NOT1 (N5524, N5497);
not NOT1 (N5525, N5511);
and AND4 (N5526, N5525, N2502, N4155, N3457);
nand NAND3 (N5527, N5517, N1958, N2041);
xor XOR2 (N5528, N5519, N2607);
not NOT1 (N5529, N5524);
nor NOR4 (N5530, N5522, N3510, N2090, N1267);
xor XOR2 (N5531, N5527, N4706);
or OR2 (N5532, N5513, N3443);
and AND3 (N5533, N5532, N4283, N1924);
or OR3 (N5534, N5485, N2397, N1545);
nand NAND4 (N5535, N5533, N3724, N4068, N266);
nand NAND4 (N5536, N5521, N1680, N2300, N5275);
buf BUF1 (N5537, N5536);
and AND3 (N5538, N5537, N1049, N4720);
nor NOR3 (N5539, N5530, N3280, N2748);
nand NAND2 (N5540, N5526, N443);
nor NOR3 (N5541, N5523, N1935, N365);
and AND4 (N5542, N5534, N5368, N4454, N800);
buf BUF1 (N5543, N5518);
nor NOR2 (N5544, N5531, N1874);
nand NAND4 (N5545, N5538, N1712, N2375, N2518);
nand NAND4 (N5546, N5539, N4725, N1893, N4116);
nor NOR4 (N5547, N5528, N15, N2208, N514);
or OR3 (N5548, N5535, N439, N5205);
not NOT1 (N5549, N5547);
or OR4 (N5550, N5529, N1914, N1195, N5274);
xor XOR2 (N5551, N5548, N4062);
buf BUF1 (N5552, N5544);
not NOT1 (N5553, N5551);
nand NAND4 (N5554, N5541, N406, N123, N2343);
or OR3 (N5555, N5543, N4512, N3495);
and AND3 (N5556, N5555, N3541, N1837);
xor XOR2 (N5557, N5549, N2438);
and AND2 (N5558, N5554, N4585);
nand NAND2 (N5559, N5545, N4223);
nand NAND2 (N5560, N5550, N2183);
buf BUF1 (N5561, N5560);
nor NOR3 (N5562, N5542, N2718, N1448);
and AND3 (N5563, N5558, N2124, N1410);
buf BUF1 (N5564, N5552);
nor NOR3 (N5565, N5553, N4913, N4313);
nor NOR3 (N5566, N5564, N5152, N1762);
not NOT1 (N5567, N5561);
buf BUF1 (N5568, N5557);
buf BUF1 (N5569, N5556);
nand NAND2 (N5570, N5566, N3611);
xor XOR2 (N5571, N5570, N4349);
xor XOR2 (N5572, N5569, N1532);
or OR2 (N5573, N5559, N5234);
buf BUF1 (N5574, N5573);
not NOT1 (N5575, N5563);
nand NAND2 (N5576, N5562, N4415);
nor NOR2 (N5577, N5540, N4659);
buf BUF1 (N5578, N5571);
not NOT1 (N5579, N5567);
and AND3 (N5580, N5578, N2348, N5209);
and AND4 (N5581, N5568, N4571, N134, N1469);
nor NOR4 (N5582, N5574, N1701, N187, N3738);
nand NAND4 (N5583, N5572, N1199, N621, N2344);
nand NAND4 (N5584, N5579, N1115, N4315, N5401);
not NOT1 (N5585, N5580);
xor XOR2 (N5586, N5546, N2950);
not NOT1 (N5587, N5581);
nor NOR4 (N5588, N5576, N3757, N742, N5528);
or OR4 (N5589, N5582, N3580, N4874, N4739);
buf BUF1 (N5590, N5588);
or OR2 (N5591, N5585, N955);
and AND4 (N5592, N5584, N1474, N1680, N4277);
xor XOR2 (N5593, N5577, N5507);
nor NOR4 (N5594, N5591, N308, N1545, N1335);
nor NOR2 (N5595, N5590, N4699);
not NOT1 (N5596, N5575);
buf BUF1 (N5597, N5587);
xor XOR2 (N5598, N5586, N1147);
and AND3 (N5599, N5595, N5090, N2085);
and AND4 (N5600, N5583, N1016, N2697, N4992);
buf BUF1 (N5601, N5593);
or OR4 (N5602, N5601, N1915, N968, N2250);
not NOT1 (N5603, N5596);
buf BUF1 (N5604, N5598);
not NOT1 (N5605, N5565);
and AND4 (N5606, N5602, N1303, N3326, N3086);
and AND4 (N5607, N5599, N4617, N1748, N2029);
not NOT1 (N5608, N5606);
xor XOR2 (N5609, N5608, N5153);
not NOT1 (N5610, N5600);
nor NOR2 (N5611, N5603, N1866);
nor NOR2 (N5612, N5611, N2440);
xor XOR2 (N5613, N5594, N4316);
nor NOR4 (N5614, N5605, N5353, N4615, N960);
and AND2 (N5615, N5609, N1991);
nor NOR3 (N5616, N5614, N600, N3910);
nor NOR4 (N5617, N5616, N909, N2843, N2939);
buf BUF1 (N5618, N5613);
xor XOR2 (N5619, N5615, N4535);
buf BUF1 (N5620, N5604);
nand NAND3 (N5621, N5592, N1515, N3847);
and AND2 (N5622, N5621, N3287);
nor NOR2 (N5623, N5619, N3215);
nand NAND3 (N5624, N5589, N1602, N3424);
and AND2 (N5625, N5620, N1938);
nor NOR2 (N5626, N5618, N1405);
buf BUF1 (N5627, N5622);
nand NAND2 (N5628, N5612, N640);
or OR3 (N5629, N5625, N5348, N5163);
nand NAND4 (N5630, N5623, N1326, N1260, N3248);
xor XOR2 (N5631, N5629, N729);
xor XOR2 (N5632, N5624, N2897);
buf BUF1 (N5633, N5617);
or OR2 (N5634, N5628, N309);
nor NOR3 (N5635, N5630, N5362, N2462);
nor NOR4 (N5636, N5632, N3654, N2655, N3612);
nand NAND2 (N5637, N5597, N1962);
nor NOR3 (N5638, N5631, N3822, N5444);
nand NAND4 (N5639, N5638, N228, N3635, N2611);
and AND2 (N5640, N5634, N358);
buf BUF1 (N5641, N5636);
and AND2 (N5642, N5641, N3364);
xor XOR2 (N5643, N5640, N2484);
nor NOR2 (N5644, N5627, N3117);
or OR4 (N5645, N5607, N4652, N975, N1103);
buf BUF1 (N5646, N5626);
not NOT1 (N5647, N5644);
buf BUF1 (N5648, N5633);
or OR2 (N5649, N5646, N5229);
xor XOR2 (N5650, N5643, N3102);
not NOT1 (N5651, N5647);
buf BUF1 (N5652, N5651);
xor XOR2 (N5653, N5637, N1280);
buf BUF1 (N5654, N5648);
buf BUF1 (N5655, N5639);
nand NAND3 (N5656, N5635, N937, N2793);
or OR4 (N5657, N5610, N1296, N5605, N2294);
xor XOR2 (N5658, N5657, N1350);
nand NAND2 (N5659, N5642, N5556);
and AND4 (N5660, N5649, N2902, N2755, N4685);
xor XOR2 (N5661, N5654, N4406);
buf BUF1 (N5662, N5650);
and AND3 (N5663, N5658, N1344, N5051);
nand NAND4 (N5664, N5662, N1539, N3561, N4638);
not NOT1 (N5665, N5659);
xor XOR2 (N5666, N5653, N4794);
nand NAND2 (N5667, N5663, N1342);
or OR4 (N5668, N5661, N809, N215, N4492);
nor NOR3 (N5669, N5668, N4171, N110);
xor XOR2 (N5670, N5652, N5160);
xor XOR2 (N5671, N5666, N448);
or OR2 (N5672, N5655, N3344);
or OR4 (N5673, N5667, N3317, N3118, N186);
or OR3 (N5674, N5665, N1569, N2976);
nand NAND3 (N5675, N5660, N593, N63);
or OR4 (N5676, N5671, N3009, N1143, N3964);
and AND3 (N5677, N5673, N1862, N4316);
or OR3 (N5678, N5669, N1112, N3463);
nand NAND4 (N5679, N5674, N1123, N2821, N3937);
nand NAND2 (N5680, N5645, N2287);
xor XOR2 (N5681, N5675, N2225);
buf BUF1 (N5682, N5679);
and AND2 (N5683, N5676, N3422);
nor NOR3 (N5684, N5682, N2419, N358);
buf BUF1 (N5685, N5656);
buf BUF1 (N5686, N5683);
buf BUF1 (N5687, N5681);
not NOT1 (N5688, N5678);
xor XOR2 (N5689, N5664, N2381);
and AND3 (N5690, N5680, N1822, N5667);
and AND2 (N5691, N5677, N4664);
xor XOR2 (N5692, N5690, N2952);
or OR4 (N5693, N5684, N4579, N4478, N4823);
nor NOR4 (N5694, N5693, N2735, N5059, N1392);
and AND4 (N5695, N5686, N1612, N1147, N5170);
and AND3 (N5696, N5691, N928, N3964);
and AND4 (N5697, N5696, N1347, N4742, N5343);
not NOT1 (N5698, N5694);
xor XOR2 (N5699, N5692, N5174);
nand NAND3 (N5700, N5672, N1367, N4426);
not NOT1 (N5701, N5670);
not NOT1 (N5702, N5688);
buf BUF1 (N5703, N5685);
and AND3 (N5704, N5700, N3517, N2900);
and AND4 (N5705, N5698, N2040, N2336, N1702);
not NOT1 (N5706, N5702);
nor NOR2 (N5707, N5689, N2879);
xor XOR2 (N5708, N5705, N1473);
xor XOR2 (N5709, N5707, N3231);
and AND4 (N5710, N5695, N1832, N3268, N33);
not NOT1 (N5711, N5710);
nand NAND2 (N5712, N5706, N954);
and AND2 (N5713, N5704, N1573);
nand NAND4 (N5714, N5701, N4536, N4879, N4522);
xor XOR2 (N5715, N5711, N870);
xor XOR2 (N5716, N5687, N660);
nand NAND3 (N5717, N5709, N4188, N1333);
and AND4 (N5718, N5712, N575, N1804, N1806);
or OR3 (N5719, N5716, N1357, N1173);
not NOT1 (N5720, N5719);
buf BUF1 (N5721, N5715);
buf BUF1 (N5722, N5721);
xor XOR2 (N5723, N5722, N2902);
or OR2 (N5724, N5714, N1605);
not NOT1 (N5725, N5708);
buf BUF1 (N5726, N5718);
and AND4 (N5727, N5697, N4548, N283, N105);
not NOT1 (N5728, N5713);
and AND2 (N5729, N5717, N208);
nand NAND3 (N5730, N5720, N3052, N3230);
xor XOR2 (N5731, N5730, N1758);
xor XOR2 (N5732, N5699, N829);
nand NAND4 (N5733, N5703, N3579, N2722, N798);
nand NAND2 (N5734, N5726, N4933);
or OR4 (N5735, N5727, N723, N3155, N1266);
and AND4 (N5736, N5734, N320, N4932, N3415);
nand NAND2 (N5737, N5735, N2920);
nand NAND4 (N5738, N5729, N4364, N3480, N4206);
and AND4 (N5739, N5738, N4322, N2163, N3667);
buf BUF1 (N5740, N5739);
or OR4 (N5741, N5731, N551, N1131, N1591);
nand NAND3 (N5742, N5737, N762, N4529);
xor XOR2 (N5743, N5742, N320);
and AND4 (N5744, N5732, N4236, N5370, N4331);
xor XOR2 (N5745, N5724, N1788);
or OR2 (N5746, N5740, N3999);
xor XOR2 (N5747, N5743, N2422);
and AND3 (N5748, N5744, N3477, N905);
nand NAND3 (N5749, N5736, N1833, N2317);
or OR3 (N5750, N5748, N4827, N2381);
xor XOR2 (N5751, N5747, N2207);
and AND4 (N5752, N5750, N1671, N4266, N4893);
buf BUF1 (N5753, N5728);
buf BUF1 (N5754, N5749);
nor NOR3 (N5755, N5754, N3841, N2674);
buf BUF1 (N5756, N5753);
nor NOR2 (N5757, N5752, N5506);
nor NOR4 (N5758, N5746, N197, N723, N4543);
xor XOR2 (N5759, N5741, N4738);
xor XOR2 (N5760, N5725, N2431);
buf BUF1 (N5761, N5745);
and AND3 (N5762, N5756, N2308, N3550);
nand NAND4 (N5763, N5733, N1751, N4002, N5749);
xor XOR2 (N5764, N5760, N4513);
not NOT1 (N5765, N5764);
nor NOR4 (N5766, N5762, N4337, N2650, N4916);
nor NOR4 (N5767, N5765, N5539, N4723, N3771);
buf BUF1 (N5768, N5763);
not NOT1 (N5769, N5759);
not NOT1 (N5770, N5723);
or OR4 (N5771, N5767, N484, N5714, N4639);
and AND2 (N5772, N5751, N4579);
or OR2 (N5773, N5757, N3121);
and AND4 (N5774, N5761, N1249, N1096, N3456);
xor XOR2 (N5775, N5772, N285);
nand NAND2 (N5776, N5769, N4956);
xor XOR2 (N5777, N5755, N5677);
nand NAND3 (N5778, N5768, N3637, N3531);
buf BUF1 (N5779, N5775);
nor NOR3 (N5780, N5778, N2506, N1278);
nand NAND4 (N5781, N5766, N3569, N3047, N3031);
nand NAND4 (N5782, N5781, N2535, N2050, N4154);
nor NOR3 (N5783, N5779, N2213, N3627);
buf BUF1 (N5784, N5783);
buf BUF1 (N5785, N5771);
not NOT1 (N5786, N5782);
or OR3 (N5787, N5784, N3667, N153);
not NOT1 (N5788, N5777);
not NOT1 (N5789, N5788);
or OR4 (N5790, N5785, N1641, N5192, N1312);
nor NOR2 (N5791, N5780, N2719);
not NOT1 (N5792, N5774);
nor NOR4 (N5793, N5790, N3557, N1384, N158);
or OR3 (N5794, N5787, N2928, N5091);
or OR2 (N5795, N5789, N3623);
and AND4 (N5796, N5776, N362, N129, N2745);
nand NAND4 (N5797, N5792, N54, N569, N2796);
not NOT1 (N5798, N5795);
or OR4 (N5799, N5773, N317, N1073, N5114);
not NOT1 (N5800, N5791);
nand NAND4 (N5801, N5800, N5697, N4072, N5056);
not NOT1 (N5802, N5796);
or OR4 (N5803, N5770, N4367, N944, N3898);
and AND4 (N5804, N5758, N4012, N2965, N3592);
xor XOR2 (N5805, N5801, N4108);
and AND2 (N5806, N5804, N3505);
or OR4 (N5807, N5786, N3224, N2036, N2373);
nand NAND3 (N5808, N5807, N5427, N3233);
buf BUF1 (N5809, N5806);
not NOT1 (N5810, N5809);
and AND3 (N5811, N5803, N5776, N478);
buf BUF1 (N5812, N5794);
nand NAND3 (N5813, N5797, N4954, N3187);
and AND3 (N5814, N5810, N2538, N1007);
not NOT1 (N5815, N5805);
xor XOR2 (N5816, N5811, N4016);
xor XOR2 (N5817, N5814, N4320);
not NOT1 (N5818, N5798);
nor NOR4 (N5819, N5813, N1383, N5209, N1494);
xor XOR2 (N5820, N5799, N3988);
nand NAND3 (N5821, N5812, N5784, N2291);
nor NOR4 (N5822, N5818, N5558, N2709, N1874);
not NOT1 (N5823, N5821);
nand NAND2 (N5824, N5816, N3630);
and AND2 (N5825, N5793, N1781);
nor NOR3 (N5826, N5817, N2179, N2052);
nand NAND2 (N5827, N5820, N3355);
not NOT1 (N5828, N5824);
buf BUF1 (N5829, N5819);
nor NOR3 (N5830, N5823, N3603, N2920);
and AND2 (N5831, N5828, N468);
nor NOR4 (N5832, N5826, N1675, N461, N3430);
not NOT1 (N5833, N5808);
buf BUF1 (N5834, N5825);
or OR3 (N5835, N5834, N1845, N1826);
not NOT1 (N5836, N5829);
and AND4 (N5837, N5836, N1752, N5684, N5597);
nor NOR3 (N5838, N5802, N5091, N1670);
buf BUF1 (N5839, N5835);
nor NOR4 (N5840, N5839, N4368, N2306, N877);
and AND4 (N5841, N5830, N891, N5493, N1984);
or OR3 (N5842, N5838, N4816, N3693);
or OR2 (N5843, N5842, N3526);
xor XOR2 (N5844, N5843, N579);
or OR2 (N5845, N5844, N4088);
and AND2 (N5846, N5815, N2649);
xor XOR2 (N5847, N5833, N4919);
xor XOR2 (N5848, N5841, N1694);
nand NAND2 (N5849, N5832, N3633);
buf BUF1 (N5850, N5840);
and AND3 (N5851, N5827, N2866, N4578);
buf BUF1 (N5852, N5845);
xor XOR2 (N5853, N5849, N3909);
xor XOR2 (N5854, N5853, N5650);
buf BUF1 (N5855, N5837);
and AND3 (N5856, N5855, N1042, N3742);
buf BUF1 (N5857, N5852);
nand NAND4 (N5858, N5822, N614, N2138, N4633);
xor XOR2 (N5859, N5856, N2723);
nor NOR4 (N5860, N5858, N5562, N746, N4283);
and AND4 (N5861, N5847, N2540, N4134, N3674);
buf BUF1 (N5862, N5857);
buf BUF1 (N5863, N5848);
or OR2 (N5864, N5850, N1886);
not NOT1 (N5865, N5854);
and AND3 (N5866, N5831, N740, N1276);
or OR2 (N5867, N5846, N2233);
or OR3 (N5868, N5863, N3805, N381);
not NOT1 (N5869, N5868);
buf BUF1 (N5870, N5860);
xor XOR2 (N5871, N5866, N3765);
nor NOR2 (N5872, N5859, N3788);
and AND2 (N5873, N5864, N4865);
or OR3 (N5874, N5851, N5646, N3534);
nand NAND2 (N5875, N5867, N279);
or OR3 (N5876, N5862, N5228, N1477);
nand NAND3 (N5877, N5876, N4271, N5787);
nor NOR2 (N5878, N5869, N323);
buf BUF1 (N5879, N5865);
xor XOR2 (N5880, N5878, N2206);
nand NAND3 (N5881, N5880, N1751, N3791);
nor NOR2 (N5882, N5871, N4923);
or OR3 (N5883, N5877, N4194, N5754);
not NOT1 (N5884, N5883);
xor XOR2 (N5885, N5873, N2591);
not NOT1 (N5886, N5872);
or OR3 (N5887, N5861, N2436, N1557);
nand NAND2 (N5888, N5875, N4133);
nor NOR4 (N5889, N5886, N4346, N3756, N4714);
nand NAND3 (N5890, N5884, N4366, N4872);
nor NOR2 (N5891, N5889, N3082);
not NOT1 (N5892, N5890);
or OR4 (N5893, N5882, N4384, N1487, N2839);
or OR4 (N5894, N5887, N572, N2720, N2789);
or OR2 (N5895, N5891, N2178);
nand NAND4 (N5896, N5870, N3500, N2134, N2420);
or OR4 (N5897, N5888, N1262, N4366, N3098);
nand NAND4 (N5898, N5885, N5380, N4305, N620);
nand NAND3 (N5899, N5898, N1087, N3464);
nand NAND4 (N5900, N5892, N3141, N3556, N4240);
nand NAND3 (N5901, N5895, N133, N1885);
and AND3 (N5902, N5894, N1786, N2654);
buf BUF1 (N5903, N5893);
and AND4 (N5904, N5901, N2422, N457, N2329);
or OR3 (N5905, N5897, N3656, N265);
or OR3 (N5906, N5879, N4847, N5547);
or OR3 (N5907, N5905, N2405, N4123);
xor XOR2 (N5908, N5900, N4533);
nand NAND3 (N5909, N5881, N3321, N4824);
xor XOR2 (N5910, N5896, N1248);
not NOT1 (N5911, N5904);
nand NAND4 (N5912, N5910, N1474, N4501, N4292);
nor NOR2 (N5913, N5912, N4540);
or OR4 (N5914, N5911, N4677, N697, N2432);
or OR2 (N5915, N5908, N2238);
and AND2 (N5916, N5902, N4321);
or OR4 (N5917, N5874, N3071, N470, N4146);
and AND2 (N5918, N5909, N1887);
nand NAND3 (N5919, N5915, N3832, N4353);
and AND4 (N5920, N5899, N2812, N3045, N1829);
not NOT1 (N5921, N5914);
not NOT1 (N5922, N5907);
or OR4 (N5923, N5903, N5733, N2385, N160);
or OR4 (N5924, N5918, N2476, N1538, N5694);
not NOT1 (N5925, N5919);
buf BUF1 (N5926, N5913);
not NOT1 (N5927, N5921);
and AND2 (N5928, N5926, N4382);
nor NOR4 (N5929, N5906, N43, N2285, N5200);
nand NAND4 (N5930, N5923, N4634, N4304, N5788);
nand NAND2 (N5931, N5930, N3665);
buf BUF1 (N5932, N5924);
nor NOR4 (N5933, N5922, N4141, N2187, N3420);
or OR4 (N5934, N5916, N3371, N1783, N3536);
or OR3 (N5935, N5934, N322, N3390);
nor NOR2 (N5936, N5925, N4314);
and AND3 (N5937, N5928, N5421, N5844);
and AND4 (N5938, N5932, N1135, N2182, N5640);
xor XOR2 (N5939, N5937, N5825);
buf BUF1 (N5940, N5936);
and AND3 (N5941, N5938, N4786, N3240);
or OR4 (N5942, N5931, N1108, N2194, N3464);
nor NOR2 (N5943, N5917, N5761);
buf BUF1 (N5944, N5939);
nand NAND3 (N5945, N5933, N4877, N5749);
xor XOR2 (N5946, N5920, N339);
buf BUF1 (N5947, N5944);
not NOT1 (N5948, N5942);
and AND4 (N5949, N5940, N2479, N70, N4570);
not NOT1 (N5950, N5945);
or OR2 (N5951, N5941, N4221);
xor XOR2 (N5952, N5935, N217);
not NOT1 (N5953, N5948);
xor XOR2 (N5954, N5950, N4199);
nor NOR4 (N5955, N5946, N2875, N3560, N4154);
xor XOR2 (N5956, N5949, N4964);
buf BUF1 (N5957, N5952);
and AND3 (N5958, N5943, N5854, N4586);
xor XOR2 (N5959, N5929, N889);
nand NAND3 (N5960, N5927, N979, N4969);
nand NAND2 (N5961, N5957, N4858);
or OR2 (N5962, N5954, N4452);
and AND4 (N5963, N5958, N5337, N4281, N525);
nand NAND4 (N5964, N5953, N772, N645, N960);
not NOT1 (N5965, N5956);
nor NOR3 (N5966, N5960, N3175, N3153);
buf BUF1 (N5967, N5955);
or OR2 (N5968, N5947, N1600);
xor XOR2 (N5969, N5966, N5009);
xor XOR2 (N5970, N5965, N4530);
buf BUF1 (N5971, N5963);
and AND3 (N5972, N5964, N3161, N1868);
nand NAND4 (N5973, N5961, N273, N772, N4569);
nor NOR4 (N5974, N5970, N3919, N1274, N1105);
nor NOR4 (N5975, N5959, N4257, N4758, N2231);
or OR4 (N5976, N5972, N1867, N1599, N4671);
or OR2 (N5977, N5962, N2210);
buf BUF1 (N5978, N5967);
xor XOR2 (N5979, N5974, N5070);
buf BUF1 (N5980, N5978);
buf BUF1 (N5981, N5976);
not NOT1 (N5982, N5975);
nand NAND4 (N5983, N5980, N3377, N2513, N2841);
nor NOR3 (N5984, N5969, N1820, N2294);
not NOT1 (N5985, N5984);
not NOT1 (N5986, N5968);
and AND2 (N5987, N5979, N4637);
and AND3 (N5988, N5982, N1147, N2664);
or OR4 (N5989, N5983, N3040, N5604, N3626);
or OR3 (N5990, N5951, N3753, N3858);
and AND3 (N5991, N5985, N4602, N2545);
nand NAND4 (N5992, N5971, N5150, N1567, N4434);
xor XOR2 (N5993, N5981, N4244);
or OR3 (N5994, N5990, N1909, N4848);
xor XOR2 (N5995, N5987, N5426);
not NOT1 (N5996, N5993);
nand NAND3 (N5997, N5988, N5547, N3852);
nand NAND2 (N5998, N5994, N5643);
nand NAND3 (N5999, N5977, N4064, N5314);
nor NOR2 (N6000, N5997, N3102);
xor XOR2 (N6001, N5986, N543);
not NOT1 (N6002, N5992);
or OR2 (N6003, N5996, N4006);
not NOT1 (N6004, N5989);
xor XOR2 (N6005, N6000, N789);
and AND4 (N6006, N6002, N2071, N3744, N429);
or OR2 (N6007, N6004, N4120);
xor XOR2 (N6008, N5999, N387);
not NOT1 (N6009, N6003);
nand NAND3 (N6010, N6008, N922, N3927);
or OR4 (N6011, N6005, N616, N2008, N4401);
buf BUF1 (N6012, N5991);
buf BUF1 (N6013, N5973);
nand NAND2 (N6014, N6010, N4614);
nor NOR4 (N6015, N6001, N585, N4820, N675);
not NOT1 (N6016, N6015);
or OR4 (N6017, N6007, N1070, N1497, N2476);
not NOT1 (N6018, N6006);
and AND4 (N6019, N5998, N4490, N2704, N1062);
xor XOR2 (N6020, N6017, N3743);
nand NAND3 (N6021, N6019, N5993, N3680);
xor XOR2 (N6022, N6014, N4497);
xor XOR2 (N6023, N6021, N1527);
not NOT1 (N6024, N6009);
nand NAND4 (N6025, N6020, N4771, N5540, N4961);
and AND2 (N6026, N6011, N1114);
xor XOR2 (N6027, N6016, N326);
not NOT1 (N6028, N6024);
not NOT1 (N6029, N6013);
nand NAND2 (N6030, N6025, N2167);
nand NAND4 (N6031, N6022, N1719, N1037, N2003);
not NOT1 (N6032, N6031);
nor NOR3 (N6033, N6029, N5157, N5362);
or OR4 (N6034, N6018, N3466, N2449, N537);
not NOT1 (N6035, N6023);
nand NAND3 (N6036, N6033, N979, N4893);
nand NAND3 (N6037, N6027, N1759, N4047);
or OR3 (N6038, N6032, N6018, N4666);
or OR2 (N6039, N6026, N2614);
xor XOR2 (N6040, N6035, N4129);
nor NOR4 (N6041, N6012, N2926, N5204, N5346);
nor NOR2 (N6042, N6034, N3537);
xor XOR2 (N6043, N6036, N2151);
not NOT1 (N6044, N6028);
nand NAND4 (N6045, N6043, N722, N1170, N4537);
buf BUF1 (N6046, N6030);
nor NOR4 (N6047, N6040, N5011, N1221, N2171);
or OR3 (N6048, N6044, N2803, N2580);
buf BUF1 (N6049, N6045);
buf BUF1 (N6050, N6042);
xor XOR2 (N6051, N6037, N1357);
or OR3 (N6052, N5995, N4827, N273);
buf BUF1 (N6053, N6051);
nor NOR3 (N6054, N6041, N4493, N2067);
not NOT1 (N6055, N6050);
nand NAND2 (N6056, N6054, N1152);
xor XOR2 (N6057, N6039, N2820);
nand NAND4 (N6058, N6055, N1929, N4096, N3334);
nor NOR2 (N6059, N6058, N5953);
not NOT1 (N6060, N6048);
and AND2 (N6061, N6046, N4366);
not NOT1 (N6062, N6038);
nor NOR2 (N6063, N6062, N1029);
and AND2 (N6064, N6056, N3478);
not NOT1 (N6065, N6052);
or OR2 (N6066, N6059, N1652);
or OR3 (N6067, N6049, N408, N578);
not NOT1 (N6068, N6067);
not NOT1 (N6069, N6065);
nor NOR3 (N6070, N6063, N2957, N4179);
buf BUF1 (N6071, N6070);
nand NAND4 (N6072, N6061, N5700, N4359, N3587);
nand NAND2 (N6073, N6069, N5345);
xor XOR2 (N6074, N6060, N1946);
xor XOR2 (N6075, N6071, N5021);
or OR3 (N6076, N6068, N3586, N4832);
nor NOR2 (N6077, N6057, N1082);
and AND2 (N6078, N6076, N1229);
and AND3 (N6079, N6066, N2288, N6045);
not NOT1 (N6080, N6077);
buf BUF1 (N6081, N6074);
not NOT1 (N6082, N6047);
buf BUF1 (N6083, N6072);
buf BUF1 (N6084, N6081);
nor NOR4 (N6085, N6080, N5291, N3490, N1443);
and AND3 (N6086, N6082, N3923, N3630);
not NOT1 (N6087, N6078);
buf BUF1 (N6088, N6086);
xor XOR2 (N6089, N6085, N5491);
xor XOR2 (N6090, N6053, N4266);
or OR3 (N6091, N6088, N3026, N4895);
nand NAND3 (N6092, N6089, N4335, N1584);
buf BUF1 (N6093, N6092);
nand NAND2 (N6094, N6079, N4668);
buf BUF1 (N6095, N6087);
nor NOR3 (N6096, N6093, N2875, N4590);
or OR2 (N6097, N6084, N4612);
buf BUF1 (N6098, N6073);
nand NAND3 (N6099, N6097, N4331, N4364);
buf BUF1 (N6100, N6098);
nand NAND3 (N6101, N6099, N3716, N1188);
nand NAND4 (N6102, N6100, N2798, N518, N5990);
xor XOR2 (N6103, N6101, N1359);
or OR4 (N6104, N6095, N659, N1290, N2037);
xor XOR2 (N6105, N6104, N3440);
nor NOR4 (N6106, N6064, N2561, N1672, N2010);
nor NOR3 (N6107, N6102, N83, N3578);
xor XOR2 (N6108, N6107, N4632);
buf BUF1 (N6109, N6091);
or OR2 (N6110, N6108, N994);
or OR4 (N6111, N6090, N242, N4602, N785);
nor NOR3 (N6112, N6110, N498, N5188);
and AND4 (N6113, N6096, N4923, N4179, N2472);
buf BUF1 (N6114, N6094);
not NOT1 (N6115, N6111);
nand NAND4 (N6116, N6109, N119, N997, N6111);
nor NOR2 (N6117, N6106, N1125);
or OR2 (N6118, N6113, N4512);
buf BUF1 (N6119, N6114);
nor NOR4 (N6120, N6112, N6075, N1236, N4683);
and AND4 (N6121, N1010, N720, N2339, N4060);
nand NAND4 (N6122, N6115, N3343, N3422, N1870);
buf BUF1 (N6123, N6105);
not NOT1 (N6124, N6116);
nor NOR4 (N6125, N6121, N5408, N4364, N842);
or OR3 (N6126, N6119, N3736, N5325);
buf BUF1 (N6127, N6125);
or OR4 (N6128, N6120, N5754, N5210, N695);
and AND2 (N6129, N6103, N4553);
buf BUF1 (N6130, N6126);
nand NAND4 (N6131, N6129, N5684, N3512, N5946);
buf BUF1 (N6132, N6123);
or OR4 (N6133, N6118, N5887, N3871, N1292);
and AND4 (N6134, N6131, N446, N4356, N1655);
not NOT1 (N6135, N6134);
not NOT1 (N6136, N6117);
and AND4 (N6137, N6124, N3069, N4291, N1622);
xor XOR2 (N6138, N6083, N2089);
xor XOR2 (N6139, N6138, N243);
xor XOR2 (N6140, N6135, N196);
xor XOR2 (N6141, N6136, N6030);
nor NOR4 (N6142, N6139, N4600, N1295, N1098);
buf BUF1 (N6143, N6127);
or OR2 (N6144, N6140, N3525);
and AND2 (N6145, N6144, N1393);
nand NAND3 (N6146, N6137, N3747, N3547);
xor XOR2 (N6147, N6145, N1385);
buf BUF1 (N6148, N6146);
xor XOR2 (N6149, N6128, N35);
or OR3 (N6150, N6132, N2979, N6065);
nand NAND4 (N6151, N6150, N244, N5365, N1232);
nand NAND2 (N6152, N6151, N5890);
not NOT1 (N6153, N6143);
nand NAND2 (N6154, N6152, N3794);
nor NOR2 (N6155, N6130, N2044);
buf BUF1 (N6156, N6133);
buf BUF1 (N6157, N6147);
nand NAND2 (N6158, N6148, N3344);
buf BUF1 (N6159, N6122);
xor XOR2 (N6160, N6156, N5910);
or OR3 (N6161, N6149, N1742, N2496);
or OR2 (N6162, N6141, N1659);
or OR4 (N6163, N6160, N3441, N4321, N3745);
xor XOR2 (N6164, N6158, N119);
not NOT1 (N6165, N6157);
xor XOR2 (N6166, N6153, N4022);
buf BUF1 (N6167, N6164);
xor XOR2 (N6168, N6165, N3099);
nor NOR4 (N6169, N6142, N812, N2555, N5753);
nor NOR2 (N6170, N6154, N6038);
not NOT1 (N6171, N6170);
xor XOR2 (N6172, N6166, N702);
or OR4 (N6173, N6155, N2081, N2285, N679);
xor XOR2 (N6174, N6163, N5863);
xor XOR2 (N6175, N6167, N3843);
xor XOR2 (N6176, N6161, N2988);
and AND3 (N6177, N6168, N5752, N5903);
and AND4 (N6178, N6175, N1604, N2396, N5771);
nand NAND3 (N6179, N6162, N4316, N4183);
not NOT1 (N6180, N6171);
not NOT1 (N6181, N6174);
buf BUF1 (N6182, N6180);
not NOT1 (N6183, N6173);
nor NOR2 (N6184, N6176, N2528);
xor XOR2 (N6185, N6183, N2736);
not NOT1 (N6186, N6181);
nand NAND3 (N6187, N6172, N5047, N5359);
or OR2 (N6188, N6186, N2851);
xor XOR2 (N6189, N6159, N1814);
buf BUF1 (N6190, N6169);
xor XOR2 (N6191, N6177, N6050);
nand NAND2 (N6192, N6191, N1128);
nor NOR4 (N6193, N6192, N3671, N607, N53);
nand NAND3 (N6194, N6185, N2783, N2078);
nor NOR3 (N6195, N6182, N5473, N3706);
or OR4 (N6196, N6193, N5407, N2158, N2499);
nand NAND2 (N6197, N6187, N4573);
nor NOR3 (N6198, N6189, N1511, N3703);
or OR3 (N6199, N6197, N3140, N5530);
nand NAND4 (N6200, N6179, N1964, N3239, N6194);
nor NOR4 (N6201, N639, N2486, N2335, N2843);
or OR3 (N6202, N6195, N6090, N3052);
buf BUF1 (N6203, N6202);
and AND3 (N6204, N6184, N5644, N3234);
not NOT1 (N6205, N6196);
nand NAND3 (N6206, N6188, N3691, N1381);
or OR3 (N6207, N6200, N1660, N2097);
or OR3 (N6208, N6190, N6172, N1613);
xor XOR2 (N6209, N6207, N1269);
nor NOR3 (N6210, N6178, N735, N4539);
xor XOR2 (N6211, N6201, N40);
or OR2 (N6212, N6206, N2956);
xor XOR2 (N6213, N6211, N4514);
xor XOR2 (N6214, N6205, N1246);
not NOT1 (N6215, N6212);
xor XOR2 (N6216, N6210, N2700);
buf BUF1 (N6217, N6215);
nor NOR2 (N6218, N6204, N69);
buf BUF1 (N6219, N6213);
xor XOR2 (N6220, N6209, N3110);
not NOT1 (N6221, N6214);
nor NOR2 (N6222, N6217, N2163);
not NOT1 (N6223, N6208);
or OR4 (N6224, N6223, N4720, N5257, N1039);
not NOT1 (N6225, N6219);
and AND3 (N6226, N6225, N5884, N50);
nand NAND3 (N6227, N6203, N436, N3481);
or OR4 (N6228, N6199, N1606, N5383, N4605);
or OR4 (N6229, N6227, N2855, N5006, N1596);
xor XOR2 (N6230, N6198, N4005);
not NOT1 (N6231, N6216);
nor NOR3 (N6232, N6224, N6022, N717);
buf BUF1 (N6233, N6229);
buf BUF1 (N6234, N6231);
not NOT1 (N6235, N6232);
or OR3 (N6236, N6233, N4679, N1364);
xor XOR2 (N6237, N6220, N857);
or OR3 (N6238, N6221, N2382, N2364);
buf BUF1 (N6239, N6230);
xor XOR2 (N6240, N6228, N4955);
nand NAND2 (N6241, N6222, N884);
xor XOR2 (N6242, N6234, N4802);
xor XOR2 (N6243, N6242, N3440);
nand NAND3 (N6244, N6236, N3235, N319);
not NOT1 (N6245, N6226);
nand NAND4 (N6246, N6241, N1675, N3087, N5405);
nor NOR3 (N6247, N6235, N6160, N4714);
nand NAND2 (N6248, N6238, N1393);
xor XOR2 (N6249, N6245, N3480);
nand NAND3 (N6250, N6247, N4705, N1858);
buf BUF1 (N6251, N6248);
xor XOR2 (N6252, N6246, N3184);
not NOT1 (N6253, N6249);
nor NOR4 (N6254, N6240, N245, N3577, N3867);
not NOT1 (N6255, N6251);
or OR2 (N6256, N6244, N6014);
buf BUF1 (N6257, N6252);
or OR2 (N6258, N6218, N4736);
not NOT1 (N6259, N6254);
and AND2 (N6260, N6250, N4840);
nor NOR4 (N6261, N6239, N2951, N4055, N1701);
nor NOR3 (N6262, N6257, N4159, N6045);
xor XOR2 (N6263, N6237, N1235);
or OR2 (N6264, N6253, N1863);
buf BUF1 (N6265, N6264);
buf BUF1 (N6266, N6256);
nand NAND3 (N6267, N6263, N735, N2945);
not NOT1 (N6268, N6265);
not NOT1 (N6269, N6260);
xor XOR2 (N6270, N6261, N4693);
xor XOR2 (N6271, N6269, N2638);
buf BUF1 (N6272, N6271);
nand NAND3 (N6273, N6255, N162, N5246);
nand NAND2 (N6274, N6259, N4450);
xor XOR2 (N6275, N6274, N6130);
nor NOR3 (N6276, N6266, N3046, N21);
nor NOR3 (N6277, N6273, N5969, N6250);
not NOT1 (N6278, N6267);
nor NOR4 (N6279, N6268, N6103, N4408, N3607);
xor XOR2 (N6280, N6272, N4879);
not NOT1 (N6281, N6276);
and AND4 (N6282, N6262, N929, N4843, N3322);
nor NOR2 (N6283, N6281, N5999);
buf BUF1 (N6284, N6279);
not NOT1 (N6285, N6277);
and AND4 (N6286, N6280, N5479, N6251, N1363);
buf BUF1 (N6287, N6284);
and AND3 (N6288, N6282, N710, N3300);
xor XOR2 (N6289, N6275, N1388);
nor NOR3 (N6290, N6287, N5516, N1099);
nand NAND4 (N6291, N6286, N885, N5889, N5364);
or OR2 (N6292, N6290, N5155);
nand NAND4 (N6293, N6258, N6290, N5230, N4732);
or OR4 (N6294, N6292, N1410, N579, N2958);
nand NAND3 (N6295, N6291, N1150, N5881);
nand NAND4 (N6296, N6295, N5002, N3323, N5005);
buf BUF1 (N6297, N6270);
and AND2 (N6298, N6288, N1733);
and AND4 (N6299, N6297, N766, N705, N4652);
nor NOR2 (N6300, N6285, N3029);
and AND3 (N6301, N6294, N5978, N2211);
nand NAND4 (N6302, N6298, N4578, N3512, N5575);
and AND4 (N6303, N6299, N2468, N3096, N2696);
xor XOR2 (N6304, N6283, N5644);
xor XOR2 (N6305, N6302, N2795);
xor XOR2 (N6306, N6304, N2148);
or OR3 (N6307, N6303, N5152, N4136);
xor XOR2 (N6308, N6301, N3879);
nand NAND3 (N6309, N6305, N4143, N270);
or OR4 (N6310, N6289, N3960, N3113, N4603);
nor NOR2 (N6311, N6307, N2751);
xor XOR2 (N6312, N6296, N3160);
nor NOR4 (N6313, N6310, N3307, N2126, N3508);
nor NOR4 (N6314, N6306, N5157, N1918, N3765);
xor XOR2 (N6315, N6243, N2158);
or OR2 (N6316, N6293, N4321);
xor XOR2 (N6317, N6311, N2497);
buf BUF1 (N6318, N6312);
not NOT1 (N6319, N6317);
nor NOR2 (N6320, N6316, N5160);
buf BUF1 (N6321, N6315);
and AND4 (N6322, N6278, N2524, N1888, N5502);
xor XOR2 (N6323, N6300, N4195);
xor XOR2 (N6324, N6309, N1049);
or OR3 (N6325, N6319, N870, N24);
and AND3 (N6326, N6314, N2102, N668);
xor XOR2 (N6327, N6308, N3837);
not NOT1 (N6328, N6327);
nand NAND4 (N6329, N6328, N1093, N1759, N3838);
xor XOR2 (N6330, N6323, N5243);
or OR4 (N6331, N6329, N5382, N304, N5379);
and AND3 (N6332, N6326, N1199, N2024);
buf BUF1 (N6333, N6325);
nand NAND2 (N6334, N6313, N3434);
xor XOR2 (N6335, N6321, N419);
buf BUF1 (N6336, N6324);
not NOT1 (N6337, N6318);
nor NOR2 (N6338, N6337, N3829);
buf BUF1 (N6339, N6332);
xor XOR2 (N6340, N6331, N4291);
and AND2 (N6341, N6322, N3785);
xor XOR2 (N6342, N6320, N3533);
not NOT1 (N6343, N6335);
or OR3 (N6344, N6338, N5931, N4677);
buf BUF1 (N6345, N6344);
buf BUF1 (N6346, N6340);
not NOT1 (N6347, N6336);
buf BUF1 (N6348, N6341);
not NOT1 (N6349, N6348);
or OR3 (N6350, N6339, N5877, N5459);
or OR2 (N6351, N6343, N5086);
nor NOR4 (N6352, N6330, N5673, N2633, N2139);
buf BUF1 (N6353, N6333);
or OR4 (N6354, N6345, N4397, N4057, N202);
xor XOR2 (N6355, N6334, N1169);
xor XOR2 (N6356, N6351, N5811);
not NOT1 (N6357, N6355);
not NOT1 (N6358, N6352);
nor NOR3 (N6359, N6342, N6281, N679);
nand NAND2 (N6360, N6358, N3897);
xor XOR2 (N6361, N6353, N222);
nor NOR3 (N6362, N6356, N426, N464);
or OR4 (N6363, N6361, N4144, N2606, N110);
xor XOR2 (N6364, N6346, N1946);
not NOT1 (N6365, N6364);
not NOT1 (N6366, N6365);
xor XOR2 (N6367, N6359, N5797);
or OR4 (N6368, N6366, N2702, N2840, N4425);
not NOT1 (N6369, N6350);
nand NAND3 (N6370, N6347, N1143, N2344);
xor XOR2 (N6371, N6367, N3005);
nand NAND3 (N6372, N6371, N727, N1913);
buf BUF1 (N6373, N6354);
or OR2 (N6374, N6349, N2439);
not NOT1 (N6375, N6372);
xor XOR2 (N6376, N6374, N3882);
or OR3 (N6377, N6360, N784, N2869);
or OR3 (N6378, N6369, N3223, N5974);
xor XOR2 (N6379, N6376, N5641);
not NOT1 (N6380, N6370);
buf BUF1 (N6381, N6379);
nor NOR4 (N6382, N6378, N4562, N6283, N3037);
nor NOR2 (N6383, N6362, N1186);
buf BUF1 (N6384, N6373);
nor NOR2 (N6385, N6377, N1715);
nor NOR4 (N6386, N6363, N4070, N4023, N3270);
nor NOR2 (N6387, N6384, N4150);
or OR2 (N6388, N6368, N3848);
and AND2 (N6389, N6387, N4139);
not NOT1 (N6390, N6383);
or OR3 (N6391, N6386, N6151, N1555);
nor NOR2 (N6392, N6382, N4670);
buf BUF1 (N6393, N6380);
nand NAND3 (N6394, N6357, N4491, N3695);
or OR4 (N6395, N6394, N6033, N2946, N5692);
not NOT1 (N6396, N6393);
nand NAND4 (N6397, N6385, N578, N5122, N409);
not NOT1 (N6398, N6389);
buf BUF1 (N6399, N6381);
xor XOR2 (N6400, N6398, N822);
nor NOR3 (N6401, N6375, N1395, N969);
and AND4 (N6402, N6395, N1069, N5879, N2318);
nor NOR3 (N6403, N6390, N3856, N2098);
xor XOR2 (N6404, N6401, N6360);
not NOT1 (N6405, N6399);
not NOT1 (N6406, N6397);
nor NOR4 (N6407, N6404, N5051, N4160, N6185);
or OR2 (N6408, N6406, N2521);
xor XOR2 (N6409, N6402, N876);
nor NOR4 (N6410, N6408, N5456, N345, N3097);
and AND2 (N6411, N6392, N5575);
nand NAND4 (N6412, N6388, N6100, N2524, N2228);
nor NOR2 (N6413, N6410, N1100);
and AND3 (N6414, N6391, N6290, N4064);
buf BUF1 (N6415, N6405);
xor XOR2 (N6416, N6396, N6181);
nand NAND4 (N6417, N6413, N5788, N4193, N3338);
and AND2 (N6418, N6400, N3364);
not NOT1 (N6419, N6412);
not NOT1 (N6420, N6414);
nand NAND2 (N6421, N6407, N5044);
buf BUF1 (N6422, N6411);
or OR3 (N6423, N6403, N504, N4827);
or OR3 (N6424, N6415, N2518, N605);
and AND2 (N6425, N6420, N6080);
nand NAND3 (N6426, N6424, N3572, N3732);
buf BUF1 (N6427, N6419);
nor NOR2 (N6428, N6409, N1709);
not NOT1 (N6429, N6423);
or OR3 (N6430, N6422, N1398, N3271);
nand NAND2 (N6431, N6421, N4680);
or OR4 (N6432, N6417, N3733, N2287, N3573);
and AND3 (N6433, N6432, N1143, N4283);
nand NAND2 (N6434, N6425, N1729);
xor XOR2 (N6435, N6433, N2477);
and AND2 (N6436, N6435, N6288);
or OR2 (N6437, N6428, N1317);
and AND4 (N6438, N6434, N1672, N3231, N282);
nand NAND2 (N6439, N6426, N4358);
nand NAND3 (N6440, N6431, N4485, N433);
nand NAND4 (N6441, N6437, N6119, N777, N2592);
not NOT1 (N6442, N6436);
not NOT1 (N6443, N6438);
buf BUF1 (N6444, N6440);
and AND4 (N6445, N6441, N970, N3143, N5446);
not NOT1 (N6446, N6429);
xor XOR2 (N6447, N6442, N2195);
xor XOR2 (N6448, N6445, N1911);
nor NOR2 (N6449, N6416, N5623);
nand NAND2 (N6450, N6427, N1903);
nand NAND3 (N6451, N6448, N1886, N725);
or OR2 (N6452, N6447, N3319);
or OR2 (N6453, N6451, N654);
xor XOR2 (N6454, N6449, N4730);
or OR3 (N6455, N6452, N2177, N1406);
buf BUF1 (N6456, N6444);
nand NAND4 (N6457, N6446, N4093, N521, N1463);
nand NAND3 (N6458, N6454, N5234, N4651);
buf BUF1 (N6459, N6457);
nor NOR4 (N6460, N6458, N2155, N715, N1363);
not NOT1 (N6461, N6443);
nand NAND3 (N6462, N6453, N3706, N829);
nor NOR4 (N6463, N6456, N3031, N6426, N2681);
or OR4 (N6464, N6439, N20, N1271, N5303);
xor XOR2 (N6465, N6462, N4624);
not NOT1 (N6466, N6463);
nor NOR4 (N6467, N6459, N907, N2237, N1038);
or OR4 (N6468, N6418, N1079, N1714, N5988);
or OR2 (N6469, N6465, N2927);
not NOT1 (N6470, N6464);
or OR3 (N6471, N6470, N4469, N697);
nor NOR2 (N6472, N6450, N5815);
xor XOR2 (N6473, N6460, N3684);
not NOT1 (N6474, N6467);
nand NAND4 (N6475, N6469, N5137, N447, N847);
xor XOR2 (N6476, N6475, N4226);
xor XOR2 (N6477, N6471, N1621);
or OR2 (N6478, N6461, N2243);
nor NOR4 (N6479, N6478, N1081, N3263, N855);
buf BUF1 (N6480, N6430);
and AND4 (N6481, N6473, N4213, N4030, N3132);
nand NAND2 (N6482, N6477, N28);
nand NAND4 (N6483, N6468, N6157, N3427, N3520);
not NOT1 (N6484, N6483);
buf BUF1 (N6485, N6472);
not NOT1 (N6486, N6482);
or OR3 (N6487, N6484, N1049, N4924);
or OR4 (N6488, N6487, N355, N3385, N6072);
xor XOR2 (N6489, N6466, N1900);
or OR3 (N6490, N6486, N5450, N3730);
nor NOR2 (N6491, N6474, N2901);
nor NOR3 (N6492, N6491, N6070, N5167);
not NOT1 (N6493, N6479);
nor NOR3 (N6494, N6490, N5695, N1042);
nor NOR2 (N6495, N6485, N4801);
buf BUF1 (N6496, N6489);
nand NAND3 (N6497, N6492, N1894, N6469);
nand NAND3 (N6498, N6455, N493, N4472);
buf BUF1 (N6499, N6493);
xor XOR2 (N6500, N6496, N1251);
and AND3 (N6501, N6494, N2479, N3494);
nor NOR4 (N6502, N6498, N5840, N3032, N654);
nor NOR3 (N6503, N6480, N6233, N5835);
nand NAND2 (N6504, N6495, N2005);
buf BUF1 (N6505, N6481);
buf BUF1 (N6506, N6502);
and AND2 (N6507, N6499, N4543);
nor NOR4 (N6508, N6507, N5449, N3677, N3192);
buf BUF1 (N6509, N6476);
or OR2 (N6510, N6497, N2339);
xor XOR2 (N6511, N6504, N5929);
nor NOR2 (N6512, N6500, N510);
nand NAND2 (N6513, N6503, N2037);
and AND3 (N6514, N6506, N5117, N5649);
buf BUF1 (N6515, N6514);
not NOT1 (N6516, N6505);
and AND4 (N6517, N6510, N1722, N2943, N4823);
not NOT1 (N6518, N6517);
nor NOR2 (N6519, N6518, N5);
xor XOR2 (N6520, N6519, N1580);
nor NOR3 (N6521, N6513, N1791, N1051);
nor NOR2 (N6522, N6512, N967);
buf BUF1 (N6523, N6515);
nor NOR3 (N6524, N6509, N5090, N1162);
and AND4 (N6525, N6508, N1810, N4010, N1234);
nor NOR4 (N6526, N6516, N125, N6273, N3573);
and AND4 (N6527, N6526, N3865, N1251, N4525);
xor XOR2 (N6528, N6522, N3649);
xor XOR2 (N6529, N6511, N2389);
or OR3 (N6530, N6525, N1393, N4172);
xor XOR2 (N6531, N6524, N1350);
not NOT1 (N6532, N6520);
xor XOR2 (N6533, N6529, N3184);
and AND3 (N6534, N6531, N4723, N2260);
nand NAND4 (N6535, N6534, N6306, N362, N4818);
xor XOR2 (N6536, N6521, N285);
nand NAND3 (N6537, N6535, N1335, N4712);
nand NAND3 (N6538, N6532, N3292, N5153);
nor NOR2 (N6539, N6538, N1293);
nand NAND3 (N6540, N6527, N444, N4440);
nand NAND4 (N6541, N6539, N6060, N6022, N2317);
and AND3 (N6542, N6541, N5468, N6459);
buf BUF1 (N6543, N6537);
nor NOR2 (N6544, N6501, N3602);
xor XOR2 (N6545, N6488, N6066);
buf BUF1 (N6546, N6540);
not NOT1 (N6547, N6542);
buf BUF1 (N6548, N6528);
nand NAND4 (N6549, N6547, N2070, N642, N2104);
nor NOR4 (N6550, N6546, N2965, N5537, N34);
not NOT1 (N6551, N6544);
xor XOR2 (N6552, N6543, N3206);
xor XOR2 (N6553, N6551, N5282);
or OR3 (N6554, N6550, N4263, N5734);
and AND3 (N6555, N6549, N2704, N4021);
buf BUF1 (N6556, N6523);
nor NOR2 (N6557, N6536, N3278);
buf BUF1 (N6558, N6554);
buf BUF1 (N6559, N6555);
buf BUF1 (N6560, N6530);
xor XOR2 (N6561, N6559, N5773);
nand NAND4 (N6562, N6557, N2424, N1573, N2997);
and AND2 (N6563, N6560, N5993);
buf BUF1 (N6564, N6556);
nor NOR4 (N6565, N6552, N5302, N1023, N1148);
nand NAND2 (N6566, N6565, N2014);
xor XOR2 (N6567, N6548, N1116);
and AND4 (N6568, N6561, N5066, N5004, N6474);
buf BUF1 (N6569, N6562);
nor NOR3 (N6570, N6563, N5426, N3018);
nor NOR4 (N6571, N6567, N4896, N4686, N6493);
and AND4 (N6572, N6570, N1745, N5025, N3203);
and AND3 (N6573, N6571, N1548, N4802);
buf BUF1 (N6574, N6573);
not NOT1 (N6575, N6572);
or OR3 (N6576, N6564, N5189, N3318);
and AND4 (N6577, N6575, N68, N3415, N3792);
buf BUF1 (N6578, N6569);
nor NOR3 (N6579, N6576, N730, N2963);
xor XOR2 (N6580, N6577, N2237);
nor NOR4 (N6581, N6533, N5784, N6475, N6024);
or OR4 (N6582, N6578, N5809, N2541, N2548);
nand NAND4 (N6583, N6545, N179, N2548, N1505);
nand NAND2 (N6584, N6583, N264);
nand NAND2 (N6585, N6579, N2142);
nand NAND2 (N6586, N6584, N6013);
and AND2 (N6587, N6585, N1421);
not NOT1 (N6588, N6581);
xor XOR2 (N6589, N6558, N1002);
nand NAND3 (N6590, N6582, N1966, N2732);
buf BUF1 (N6591, N6590);
xor XOR2 (N6592, N6591, N1364);
or OR4 (N6593, N6586, N4060, N6378, N5513);
buf BUF1 (N6594, N6587);
and AND3 (N6595, N6574, N4302, N4787);
nor NOR4 (N6596, N6580, N509, N5686, N6029);
and AND3 (N6597, N6588, N2555, N5455);
not NOT1 (N6598, N6593);
not NOT1 (N6599, N6598);
buf BUF1 (N6600, N6599);
nand NAND4 (N6601, N6553, N2996, N1571, N2779);
nand NAND2 (N6602, N6600, N2598);
not NOT1 (N6603, N6566);
nand NAND4 (N6604, N6597, N4896, N2126, N2667);
nor NOR2 (N6605, N6592, N4101);
nand NAND2 (N6606, N6589, N2194);
nor NOR4 (N6607, N6605, N4850, N1559, N2982);
and AND4 (N6608, N6568, N4152, N6456, N5055);
nor NOR4 (N6609, N6601, N6172, N6082, N994);
and AND4 (N6610, N6594, N4460, N5898, N5899);
not NOT1 (N6611, N6608);
nor NOR4 (N6612, N6611, N6479, N4772, N4546);
not NOT1 (N6613, N6612);
buf BUF1 (N6614, N6610);
and AND3 (N6615, N6602, N2667, N1959);
and AND2 (N6616, N6603, N2798);
and AND4 (N6617, N6614, N4409, N806, N1354);
or OR4 (N6618, N6604, N4961, N6343, N4509);
and AND4 (N6619, N6609, N4123, N5784, N3064);
nand NAND4 (N6620, N6617, N2999, N2733, N2968);
and AND4 (N6621, N6616, N3408, N3928, N2161);
nand NAND2 (N6622, N6613, N3224);
buf BUF1 (N6623, N6619);
nand NAND4 (N6624, N6607, N4056, N3282, N5361);
nand NAND2 (N6625, N6606, N3925);
and AND4 (N6626, N6618, N6057, N745, N1832);
xor XOR2 (N6627, N6624, N3756);
and AND2 (N6628, N6615, N2431);
xor XOR2 (N6629, N6625, N190);
or OR2 (N6630, N6628, N554);
xor XOR2 (N6631, N6629, N3601);
not NOT1 (N6632, N6626);
and AND4 (N6633, N6630, N2685, N2780, N4215);
nand NAND3 (N6634, N6633, N5806, N3179);
nor NOR2 (N6635, N6632, N2624);
xor XOR2 (N6636, N6627, N6371);
or OR3 (N6637, N6631, N1088, N3089);
and AND2 (N6638, N6596, N4691);
or OR2 (N6639, N6635, N5217);
and AND3 (N6640, N6637, N3926, N5463);
and AND2 (N6641, N6622, N2467);
and AND2 (N6642, N6623, N5094);
xor XOR2 (N6643, N6620, N5122);
not NOT1 (N6644, N6621);
and AND2 (N6645, N6643, N4269);
and AND3 (N6646, N6634, N3644, N1234);
nor NOR4 (N6647, N6644, N412, N3561, N2579);
nor NOR2 (N6648, N6641, N5691);
xor XOR2 (N6649, N6648, N486);
nand NAND4 (N6650, N6640, N2981, N2438, N2821);
or OR3 (N6651, N6638, N3340, N943);
and AND2 (N6652, N6639, N5446);
xor XOR2 (N6653, N6649, N2477);
and AND2 (N6654, N6646, N84);
buf BUF1 (N6655, N6652);
buf BUF1 (N6656, N6655);
nor NOR3 (N6657, N6595, N3500, N4438);
not NOT1 (N6658, N6636);
or OR3 (N6659, N6657, N4102, N6615);
and AND2 (N6660, N6658, N6274);
nor NOR4 (N6661, N6650, N731, N520, N3045);
nand NAND3 (N6662, N6660, N1524, N4142);
or OR4 (N6663, N6647, N4196, N1171, N1317);
nor NOR3 (N6664, N6642, N2849, N6283);
or OR2 (N6665, N6653, N3461);
xor XOR2 (N6666, N6651, N6323);
xor XOR2 (N6667, N6661, N1670);
and AND3 (N6668, N6659, N2002, N5152);
or OR3 (N6669, N6665, N3124, N2240);
and AND2 (N6670, N6656, N4949);
nand NAND2 (N6671, N6667, N3034);
and AND4 (N6672, N6670, N2521, N5198, N648);
nand NAND4 (N6673, N6669, N262, N4831, N6299);
buf BUF1 (N6674, N6671);
not NOT1 (N6675, N6666);
buf BUF1 (N6676, N6654);
not NOT1 (N6677, N6673);
and AND3 (N6678, N6674, N5439, N875);
buf BUF1 (N6679, N6664);
nor NOR4 (N6680, N6679, N3638, N6662, N661);
nand NAND3 (N6681, N1942, N6296, N1044);
not NOT1 (N6682, N6645);
nor NOR4 (N6683, N6672, N4451, N1266, N844);
or OR4 (N6684, N6675, N6267, N3789, N4904);
buf BUF1 (N6685, N6682);
buf BUF1 (N6686, N6683);
buf BUF1 (N6687, N6676);
xor XOR2 (N6688, N6677, N3805);
nand NAND3 (N6689, N6686, N3978, N1043);
xor XOR2 (N6690, N6668, N5986);
xor XOR2 (N6691, N6684, N6092);
or OR3 (N6692, N6687, N4216, N6557);
or OR3 (N6693, N6663, N2426, N446);
and AND2 (N6694, N6678, N4376);
xor XOR2 (N6695, N6691, N438);
nand NAND3 (N6696, N6693, N23, N6216);
nor NOR4 (N6697, N6694, N6343, N6164, N6463);
xor XOR2 (N6698, N6695, N2512);
not NOT1 (N6699, N6690);
and AND3 (N6700, N6697, N2579, N3281);
and AND3 (N6701, N6680, N4315, N6071);
buf BUF1 (N6702, N6681);
xor XOR2 (N6703, N6685, N6361);
nor NOR3 (N6704, N6701, N5649, N2354);
buf BUF1 (N6705, N6689);
not NOT1 (N6706, N6702);
and AND2 (N6707, N6705, N945);
and AND4 (N6708, N6699, N5951, N1341, N4205);
buf BUF1 (N6709, N6707);
buf BUF1 (N6710, N6692);
buf BUF1 (N6711, N6688);
or OR3 (N6712, N6711, N2006, N3865);
xor XOR2 (N6713, N6703, N5223);
xor XOR2 (N6714, N6704, N53);
and AND3 (N6715, N6710, N2896, N5394);
xor XOR2 (N6716, N6714, N4080);
buf BUF1 (N6717, N6709);
buf BUF1 (N6718, N6712);
nand NAND4 (N6719, N6696, N2951, N814, N417);
buf BUF1 (N6720, N6713);
not NOT1 (N6721, N6698);
not NOT1 (N6722, N6700);
nor NOR3 (N6723, N6720, N4043, N3286);
or OR3 (N6724, N6717, N4125, N6070);
nand NAND2 (N6725, N6721, N409);
buf BUF1 (N6726, N6718);
buf BUF1 (N6727, N6724);
and AND3 (N6728, N6716, N4412, N5341);
or OR3 (N6729, N6725, N6098, N6463);
buf BUF1 (N6730, N6723);
nand NAND4 (N6731, N6715, N4691, N1586, N3102);
nand NAND3 (N6732, N6722, N1747, N1451);
buf BUF1 (N6733, N6719);
nor NOR4 (N6734, N6729, N4535, N1353, N2553);
xor XOR2 (N6735, N6731, N6002);
and AND4 (N6736, N6727, N4150, N1492, N6377);
or OR4 (N6737, N6726, N2678, N5674, N42);
or OR2 (N6738, N6737, N885);
nor NOR2 (N6739, N6734, N1819);
nand NAND4 (N6740, N6730, N1869, N357, N2804);
nand NAND3 (N6741, N6732, N6630, N755);
or OR3 (N6742, N6741, N4289, N820);
nand NAND2 (N6743, N6708, N6724);
nand NAND4 (N6744, N6728, N4167, N5801, N4252);
or OR2 (N6745, N6743, N6004);
nor NOR2 (N6746, N6706, N2899);
and AND3 (N6747, N6746, N1191, N1319);
nor NOR3 (N6748, N6739, N6365, N5444);
nand NAND3 (N6749, N6735, N3931, N3147);
xor XOR2 (N6750, N6738, N279);
xor XOR2 (N6751, N6742, N5046);
not NOT1 (N6752, N6744);
nand NAND4 (N6753, N6749, N6436, N6351, N4757);
nor NOR4 (N6754, N6745, N5025, N5889, N2118);
not NOT1 (N6755, N6751);
or OR4 (N6756, N6753, N2514, N2611, N4437);
xor XOR2 (N6757, N6750, N885);
not NOT1 (N6758, N6754);
nand NAND3 (N6759, N6752, N2761, N4730);
nor NOR3 (N6760, N6755, N5004, N1959);
nor NOR2 (N6761, N6748, N6066);
or OR3 (N6762, N6747, N309, N6149);
xor XOR2 (N6763, N6762, N2749);
xor XOR2 (N6764, N6758, N869);
nor NOR2 (N6765, N6763, N4515);
nor NOR4 (N6766, N6756, N5962, N2447, N5804);
nor NOR2 (N6767, N6759, N247);
xor XOR2 (N6768, N6767, N6403);
not NOT1 (N6769, N6768);
nand NAND4 (N6770, N6736, N4415, N1994, N2540);
nand NAND3 (N6771, N6766, N546, N6280);
nor NOR2 (N6772, N6771, N3450);
or OR4 (N6773, N6765, N4856, N2882, N2154);
and AND2 (N6774, N6769, N2720);
buf BUF1 (N6775, N6770);
not NOT1 (N6776, N6757);
xor XOR2 (N6777, N6776, N2702);
nor NOR4 (N6778, N6733, N6710, N1960, N4467);
buf BUF1 (N6779, N6775);
nor NOR2 (N6780, N6761, N3190);
buf BUF1 (N6781, N6779);
buf BUF1 (N6782, N6772);
or OR3 (N6783, N6774, N4029, N5357);
nor NOR2 (N6784, N6780, N1439);
and AND2 (N6785, N6777, N2947);
xor XOR2 (N6786, N6782, N1551);
not NOT1 (N6787, N6783);
not NOT1 (N6788, N6778);
or OR2 (N6789, N6760, N1600);
nor NOR3 (N6790, N6787, N2782, N3237);
xor XOR2 (N6791, N6764, N35);
buf BUF1 (N6792, N6784);
not NOT1 (N6793, N6740);
or OR2 (N6794, N6792, N692);
xor XOR2 (N6795, N6786, N5569);
and AND4 (N6796, N6785, N1153, N985, N3432);
and AND4 (N6797, N6788, N4640, N3965, N4134);
and AND4 (N6798, N6794, N2637, N6022, N1012);
not NOT1 (N6799, N6773);
or OR4 (N6800, N6793, N1147, N2974, N750);
or OR3 (N6801, N6800, N4153, N6798);
nor NOR2 (N6802, N4099, N3677);
xor XOR2 (N6803, N6795, N758);
buf BUF1 (N6804, N6802);
buf BUF1 (N6805, N6804);
not NOT1 (N6806, N6781);
or OR4 (N6807, N6789, N6290, N3878, N3816);
and AND2 (N6808, N6805, N1547);
buf BUF1 (N6809, N6807);
and AND4 (N6810, N6808, N2243, N3878, N2945);
not NOT1 (N6811, N6803);
not NOT1 (N6812, N6799);
nand NAND4 (N6813, N6811, N1510, N1869, N6386);
not NOT1 (N6814, N6806);
and AND4 (N6815, N6790, N4499, N5259, N475);
nand NAND2 (N6816, N6809, N5371);
and AND3 (N6817, N6791, N2754, N5208);
xor XOR2 (N6818, N6814, N3143);
nand NAND3 (N6819, N6797, N6539, N3544);
or OR4 (N6820, N6810, N49, N3092, N2857);
nor NOR2 (N6821, N6812, N4914);
not NOT1 (N6822, N6815);
nor NOR2 (N6823, N6818, N3006);
and AND4 (N6824, N6823, N991, N3712, N2963);
not NOT1 (N6825, N6801);
not NOT1 (N6826, N6820);
buf BUF1 (N6827, N6826);
and AND3 (N6828, N6796, N5616, N6313);
xor XOR2 (N6829, N6825, N4976);
xor XOR2 (N6830, N6829, N4309);
nor NOR3 (N6831, N6827, N6556, N862);
nor NOR3 (N6832, N6813, N4194, N656);
not NOT1 (N6833, N6832);
or OR4 (N6834, N6822, N6381, N887, N5551);
nand NAND2 (N6835, N6830, N3226);
not NOT1 (N6836, N6835);
nand NAND2 (N6837, N6828, N4274);
buf BUF1 (N6838, N6819);
nand NAND4 (N6839, N6834, N1648, N3157, N1215);
buf BUF1 (N6840, N6839);
nand NAND3 (N6841, N6837, N3897, N4271);
or OR3 (N6842, N6821, N441, N6040);
not NOT1 (N6843, N6833);
and AND2 (N6844, N6816, N654);
nand NAND2 (N6845, N6817, N2060);
nor NOR4 (N6846, N6838, N2362, N2890, N6614);
and AND3 (N6847, N6843, N3411, N6615);
nand NAND2 (N6848, N6840, N1695);
or OR3 (N6849, N6848, N4288, N2193);
nor NOR2 (N6850, N6847, N3659);
nor NOR2 (N6851, N6841, N925);
xor XOR2 (N6852, N6836, N6343);
nand NAND3 (N6853, N6852, N2972, N1535);
buf BUF1 (N6854, N6853);
or OR3 (N6855, N6831, N928, N3203);
buf BUF1 (N6856, N6854);
nor NOR4 (N6857, N6856, N2158, N3044, N3660);
xor XOR2 (N6858, N6824, N6050);
nor NOR3 (N6859, N6844, N4607, N5157);
buf BUF1 (N6860, N6849);
and AND2 (N6861, N6857, N4616);
and AND3 (N6862, N6858, N4311, N4356);
nand NAND4 (N6863, N6861, N2865, N1047, N5582);
buf BUF1 (N6864, N6859);
and AND4 (N6865, N6864, N1870, N396, N4639);
and AND2 (N6866, N6862, N4158);
nand NAND3 (N6867, N6850, N3421, N2729);
not NOT1 (N6868, N6845);
nor NOR4 (N6869, N6868, N6378, N3659, N2174);
and AND2 (N6870, N6860, N4807);
not NOT1 (N6871, N6863);
and AND3 (N6872, N6870, N850, N1734);
and AND2 (N6873, N6871, N3561);
and AND3 (N6874, N6842, N2567, N2936);
nor NOR3 (N6875, N6869, N3510, N459);
xor XOR2 (N6876, N6865, N237);
buf BUF1 (N6877, N6876);
buf BUF1 (N6878, N6855);
not NOT1 (N6879, N6878);
xor XOR2 (N6880, N6873, N4886);
and AND2 (N6881, N6877, N2513);
xor XOR2 (N6882, N6866, N3926);
not NOT1 (N6883, N6872);
and AND2 (N6884, N6880, N6301);
nor NOR2 (N6885, N6881, N6224);
xor XOR2 (N6886, N6875, N5618);
or OR2 (N6887, N6874, N4411);
buf BUF1 (N6888, N6883);
not NOT1 (N6889, N6886);
xor XOR2 (N6890, N6887, N6747);
and AND2 (N6891, N6885, N4167);
xor XOR2 (N6892, N6846, N2423);
or OR4 (N6893, N6884, N815, N4287, N806);
or OR2 (N6894, N6893, N1392);
and AND2 (N6895, N6867, N3032);
and AND4 (N6896, N6892, N3361, N4324, N2538);
xor XOR2 (N6897, N6879, N4346);
buf BUF1 (N6898, N6882);
and AND4 (N6899, N6851, N3548, N5133, N5547);
nor NOR3 (N6900, N6889, N5461, N5125);
and AND3 (N6901, N6896, N2748, N2956);
nor NOR3 (N6902, N6888, N4021, N5446);
or OR3 (N6903, N6895, N3673, N6410);
nand NAND4 (N6904, N6894, N1950, N962, N2216);
or OR2 (N6905, N6891, N1934);
buf BUF1 (N6906, N6901);
not NOT1 (N6907, N6897);
xor XOR2 (N6908, N6899, N3829);
and AND2 (N6909, N6902, N4119);
buf BUF1 (N6910, N6908);
buf BUF1 (N6911, N6907);
or OR2 (N6912, N6890, N3319);
xor XOR2 (N6913, N6905, N4535);
xor XOR2 (N6914, N6913, N6463);
nand NAND3 (N6915, N6912, N2748, N4612);
not NOT1 (N6916, N6909);
nor NOR4 (N6917, N6900, N354, N1569, N240);
nor NOR4 (N6918, N6911, N4183, N3798, N5924);
nand NAND4 (N6919, N6914, N4210, N6239, N2877);
nor NOR2 (N6920, N6915, N6676);
nor NOR4 (N6921, N6917, N6246, N1055, N4703);
xor XOR2 (N6922, N6910, N6675);
or OR4 (N6923, N6919, N2758, N1938, N5036);
or OR4 (N6924, N6904, N2670, N2043, N2303);
or OR3 (N6925, N6921, N4403, N1613);
xor XOR2 (N6926, N6916, N2691);
xor XOR2 (N6927, N6906, N1814);
and AND2 (N6928, N6903, N4660);
and AND4 (N6929, N6928, N4328, N6610, N6659);
buf BUF1 (N6930, N6924);
nand NAND4 (N6931, N6927, N2991, N2073, N1224);
buf BUF1 (N6932, N6923);
or OR4 (N6933, N6922, N4062, N2082, N800);
and AND3 (N6934, N6926, N509, N1125);
nor NOR4 (N6935, N6932, N5359, N6508, N75);
or OR4 (N6936, N6925, N5005, N2076, N2012);
nand NAND2 (N6937, N6920, N3798);
or OR2 (N6938, N6937, N648);
and AND2 (N6939, N6929, N3354);
buf BUF1 (N6940, N6935);
nand NAND2 (N6941, N6936, N329);
not NOT1 (N6942, N6938);
or OR2 (N6943, N6931, N4718);
or OR3 (N6944, N6943, N1070, N5823);
nand NAND4 (N6945, N6930, N6158, N2299, N4749);
nand NAND3 (N6946, N6944, N3765, N3026);
not NOT1 (N6947, N6941);
or OR4 (N6948, N6947, N5348, N2238, N2328);
nand NAND2 (N6949, N6940, N1404);
and AND2 (N6950, N6948, N6855);
buf BUF1 (N6951, N6939);
buf BUF1 (N6952, N6933);
nor NOR4 (N6953, N6949, N367, N2726, N620);
nand NAND3 (N6954, N6942, N1533, N4691);
buf BUF1 (N6955, N6953);
or OR2 (N6956, N6955, N1237);
not NOT1 (N6957, N6945);
nand NAND2 (N6958, N6951, N6336);
nor NOR3 (N6959, N6956, N5266, N6002);
xor XOR2 (N6960, N6934, N2544);
nor NOR3 (N6961, N6958, N1193, N1888);
not NOT1 (N6962, N6954);
or OR2 (N6963, N6960, N4787);
buf BUF1 (N6964, N6946);
or OR2 (N6965, N6962, N2224);
or OR3 (N6966, N6961, N2317, N4310);
nand NAND4 (N6967, N6966, N2825, N1666, N1086);
xor XOR2 (N6968, N6952, N4162);
xor XOR2 (N6969, N6950, N5271);
or OR2 (N6970, N6968, N6148);
xor XOR2 (N6971, N6957, N5272);
and AND2 (N6972, N6970, N5105);
nand NAND3 (N6973, N6918, N2572, N4781);
not NOT1 (N6974, N6964);
and AND2 (N6975, N6973, N3404);
and AND4 (N6976, N6971, N3447, N6683, N3242);
or OR4 (N6977, N6975, N4817, N4573, N5032);
not NOT1 (N6978, N6977);
or OR3 (N6979, N6972, N255, N4239);
or OR4 (N6980, N6976, N670, N3009, N6222);
nand NAND3 (N6981, N6898, N4478, N3373);
xor XOR2 (N6982, N6974, N3562);
buf BUF1 (N6983, N6965);
nor NOR3 (N6984, N6959, N5234, N4288);
nor NOR4 (N6985, N6963, N2812, N5581, N1914);
nor NOR4 (N6986, N6980, N6315, N6650, N3133);
and AND2 (N6987, N6979, N4542);
not NOT1 (N6988, N6978);
buf BUF1 (N6989, N6988);
nand NAND3 (N6990, N6986, N2730, N4875);
nand NAND4 (N6991, N6981, N427, N4214, N5821);
nand NAND4 (N6992, N6987, N6537, N6131, N3253);
not NOT1 (N6993, N6967);
not NOT1 (N6994, N6983);
nand NAND3 (N6995, N6991, N1408, N684);
buf BUF1 (N6996, N6984);
nand NAND3 (N6997, N6989, N3500, N3742);
xor XOR2 (N6998, N6992, N4848);
xor XOR2 (N6999, N6969, N56);
nand NAND3 (N7000, N6999, N3039, N4220);
and AND3 (N7001, N6993, N4935, N5720);
or OR2 (N7002, N6990, N6925);
nand NAND4 (N7003, N6982, N6581, N4773, N3862);
xor XOR2 (N7004, N7001, N4361);
buf BUF1 (N7005, N7002);
or OR2 (N7006, N7000, N3047);
nand NAND2 (N7007, N6995, N2218);
not NOT1 (N7008, N7007);
xor XOR2 (N7009, N7004, N2721);
and AND3 (N7010, N7009, N3808, N5568);
or OR4 (N7011, N7003, N1372, N271, N5599);
nand NAND4 (N7012, N7006, N3780, N1124, N3865);
or OR3 (N7013, N6994, N5309, N6644);
buf BUF1 (N7014, N7005);
nor NOR2 (N7015, N6996, N5327);
xor XOR2 (N7016, N7008, N5170);
nand NAND2 (N7017, N7012, N1297);
xor XOR2 (N7018, N6985, N6801);
buf BUF1 (N7019, N7017);
and AND3 (N7020, N7015, N3446, N5947);
buf BUF1 (N7021, N7016);
not NOT1 (N7022, N7014);
buf BUF1 (N7023, N7021);
not NOT1 (N7024, N7022);
and AND2 (N7025, N7013, N2684);
nor NOR3 (N7026, N6998, N3967, N886);
not NOT1 (N7027, N7026);
and AND3 (N7028, N6997, N1377, N5406);
nor NOR2 (N7029, N7028, N3319);
xor XOR2 (N7030, N7023, N6072);
buf BUF1 (N7031, N7018);
nor NOR2 (N7032, N7029, N1703);
not NOT1 (N7033, N7024);
and AND3 (N7034, N7031, N1062, N5804);
or OR3 (N7035, N7019, N2886, N3685);
xor XOR2 (N7036, N7035, N5247);
xor XOR2 (N7037, N7025, N6029);
or OR3 (N7038, N7033, N5369, N246);
nand NAND3 (N7039, N7020, N6162, N3705);
and AND2 (N7040, N7011, N2987);
nor NOR4 (N7041, N7036, N6595, N5744, N3392);
not NOT1 (N7042, N7034);
nor NOR2 (N7043, N7042, N113);
buf BUF1 (N7044, N7030);
nor NOR3 (N7045, N7038, N2557, N2607);
or OR4 (N7046, N7040, N750, N1336, N6221);
xor XOR2 (N7047, N7027, N2428);
not NOT1 (N7048, N7047);
nand NAND2 (N7049, N7039, N1980);
or OR4 (N7050, N7046, N4330, N4363, N6143);
and AND2 (N7051, N7041, N2662);
nor NOR2 (N7052, N7037, N6863);
or OR3 (N7053, N7048, N5881, N4228);
not NOT1 (N7054, N7053);
nor NOR3 (N7055, N7045, N6913, N6356);
nand NAND4 (N7056, N7032, N353, N4290, N1714);
nor NOR2 (N7057, N7049, N3338);
buf BUF1 (N7058, N7044);
and AND3 (N7059, N7010, N2635, N3032);
xor XOR2 (N7060, N7054, N2052);
nand NAND4 (N7061, N7043, N480, N6328, N2570);
xor XOR2 (N7062, N7058, N3811);
or OR2 (N7063, N7050, N4440);
and AND2 (N7064, N7052, N3454);
or OR4 (N7065, N7061, N2414, N6411, N1322);
not NOT1 (N7066, N7064);
and AND2 (N7067, N7056, N5896);
nor NOR4 (N7068, N7065, N3508, N2680, N23);
buf BUF1 (N7069, N7060);
not NOT1 (N7070, N7051);
or OR2 (N7071, N7066, N2070);
buf BUF1 (N7072, N7063);
and AND4 (N7073, N7057, N5079, N4894, N5090);
not NOT1 (N7074, N7068);
buf BUF1 (N7075, N7074);
nand NAND2 (N7076, N7070, N4721);
and AND2 (N7077, N7072, N6246);
not NOT1 (N7078, N7077);
not NOT1 (N7079, N7076);
xor XOR2 (N7080, N7073, N1509);
and AND2 (N7081, N7067, N5028);
not NOT1 (N7082, N7079);
or OR3 (N7083, N7082, N3610, N5689);
or OR3 (N7084, N7081, N2315, N2086);
or OR4 (N7085, N7084, N4865, N6344, N2126);
buf BUF1 (N7086, N7085);
not NOT1 (N7087, N7086);
or OR3 (N7088, N7083, N1462, N4547);
or OR3 (N7089, N7062, N2818, N1454);
not NOT1 (N7090, N7087);
or OR4 (N7091, N7071, N4218, N854, N5318);
nor NOR3 (N7092, N7059, N6011, N2761);
xor XOR2 (N7093, N7080, N3974);
nor NOR2 (N7094, N7089, N2151);
or OR3 (N7095, N7055, N2780, N5178);
nand NAND2 (N7096, N7078, N1795);
or OR2 (N7097, N7069, N1585);
nand NAND2 (N7098, N7088, N3576);
or OR4 (N7099, N7095, N1522, N3131, N742);
not NOT1 (N7100, N7092);
not NOT1 (N7101, N7099);
not NOT1 (N7102, N7096);
not NOT1 (N7103, N7097);
or OR3 (N7104, N7100, N3061, N4719);
buf BUF1 (N7105, N7094);
not NOT1 (N7106, N7091);
not NOT1 (N7107, N7104);
nand NAND3 (N7108, N7075, N1307, N6878);
nand NAND4 (N7109, N7101, N2243, N5748, N935);
xor XOR2 (N7110, N7102, N3770);
buf BUF1 (N7111, N7090);
or OR4 (N7112, N7110, N4844, N559, N1145);
not NOT1 (N7113, N7098);
xor XOR2 (N7114, N7109, N2552);
and AND3 (N7115, N7107, N5245, N1933);
not NOT1 (N7116, N7114);
and AND4 (N7117, N7112, N6414, N17, N5549);
nor NOR4 (N7118, N7115, N3073, N2877, N1096);
xor XOR2 (N7119, N7108, N5378);
nand NAND4 (N7120, N7105, N504, N4039, N4337);
xor XOR2 (N7121, N7120, N1382);
nor NOR3 (N7122, N7111, N634, N2845);
nor NOR2 (N7123, N7106, N1643);
nand NAND2 (N7124, N7116, N1738);
or OR3 (N7125, N7103, N1602, N128);
buf BUF1 (N7126, N7121);
and AND4 (N7127, N7125, N1952, N5138, N3921);
xor XOR2 (N7128, N7117, N4453);
not NOT1 (N7129, N7119);
buf BUF1 (N7130, N7118);
not NOT1 (N7131, N7126);
and AND4 (N7132, N7131, N6848, N4085, N2109);
xor XOR2 (N7133, N7123, N269);
buf BUF1 (N7134, N7122);
nand NAND2 (N7135, N7124, N1160);
and AND3 (N7136, N7132, N6316, N6741);
nor NOR2 (N7137, N7129, N1919);
not NOT1 (N7138, N7134);
nand NAND3 (N7139, N7137, N5990, N3055);
nor NOR3 (N7140, N7128, N2264, N752);
or OR3 (N7141, N7127, N1115, N2353);
not NOT1 (N7142, N7093);
and AND2 (N7143, N7140, N6974);
not NOT1 (N7144, N7130);
or OR4 (N7145, N7143, N4153, N4778, N1946);
and AND3 (N7146, N7141, N1729, N591);
xor XOR2 (N7147, N7133, N1726);
or OR3 (N7148, N7142, N5836, N4970);
nor NOR4 (N7149, N7145, N1142, N699, N1657);
or OR4 (N7150, N7146, N4360, N287, N2498);
or OR3 (N7151, N7148, N319, N1660);
nor NOR3 (N7152, N7149, N6153, N6677);
nor NOR4 (N7153, N7144, N5717, N1328, N4734);
nor NOR4 (N7154, N7139, N6559, N5318, N4019);
nor NOR2 (N7155, N7136, N4041);
or OR4 (N7156, N7150, N4889, N817, N3904);
xor XOR2 (N7157, N7151, N6475);
or OR3 (N7158, N7155, N353, N4029);
buf BUF1 (N7159, N7152);
buf BUF1 (N7160, N7153);
nand NAND2 (N7161, N7160, N4877);
and AND2 (N7162, N7135, N4776);
xor XOR2 (N7163, N7138, N693);
and AND2 (N7164, N7154, N1961);
or OR3 (N7165, N7157, N3194, N2077);
nand NAND4 (N7166, N7161, N596, N2038, N2159);
nand NAND4 (N7167, N7162, N2377, N1265, N4338);
xor XOR2 (N7168, N7158, N3730);
buf BUF1 (N7169, N7164);
nand NAND3 (N7170, N7166, N6933, N322);
and AND2 (N7171, N7165, N5031);
or OR3 (N7172, N7169, N3692, N4627);
nand NAND3 (N7173, N7156, N1261, N6558);
buf BUF1 (N7174, N7113);
or OR4 (N7175, N7147, N4872, N2275, N853);
nand NAND3 (N7176, N7167, N3732, N1608);
buf BUF1 (N7177, N7173);
nand NAND4 (N7178, N7159, N4410, N4009, N2926);
or OR4 (N7179, N7163, N1223, N3189, N4455);
nand NAND2 (N7180, N7174, N2111);
nor NOR2 (N7181, N7172, N1245);
or OR2 (N7182, N7176, N1692);
or OR2 (N7183, N7170, N6413);
buf BUF1 (N7184, N7183);
or OR3 (N7185, N7180, N6552, N959);
and AND2 (N7186, N7177, N1256);
buf BUF1 (N7187, N7182);
not NOT1 (N7188, N7168);
xor XOR2 (N7189, N7188, N4158);
buf BUF1 (N7190, N7179);
nand NAND4 (N7191, N7184, N1046, N544, N3876);
nand NAND3 (N7192, N7171, N2882, N3573);
buf BUF1 (N7193, N7175);
nand NAND3 (N7194, N7189, N5152, N5410);
buf BUF1 (N7195, N7186);
and AND2 (N7196, N7191, N1885);
buf BUF1 (N7197, N7193);
xor XOR2 (N7198, N7192, N2292);
or OR4 (N7199, N7194, N4445, N2373, N987);
and AND3 (N7200, N7181, N5497, N9);
xor XOR2 (N7201, N7195, N4079);
buf BUF1 (N7202, N7200);
buf BUF1 (N7203, N7199);
or OR4 (N7204, N7185, N7001, N2033, N6148);
nor NOR2 (N7205, N7202, N2811);
not NOT1 (N7206, N7190);
nor NOR3 (N7207, N7198, N6360, N512);
xor XOR2 (N7208, N7187, N3690);
xor XOR2 (N7209, N7204, N5620);
not NOT1 (N7210, N7203);
or OR4 (N7211, N7205, N6315, N5624, N459);
and AND2 (N7212, N7196, N83);
and AND3 (N7213, N7178, N339, N3514);
not NOT1 (N7214, N7212);
xor XOR2 (N7215, N7201, N929);
buf BUF1 (N7216, N7211);
xor XOR2 (N7217, N7208, N6921);
buf BUF1 (N7218, N7217);
or OR4 (N7219, N7210, N4030, N2238, N6037);
and AND4 (N7220, N7206, N7197, N7004, N5963);
nor NOR3 (N7221, N6570, N2458, N4656);
nor NOR2 (N7222, N7220, N1101);
or OR4 (N7223, N7213, N1448, N540, N2503);
nor NOR3 (N7224, N7216, N4692, N6633);
or OR2 (N7225, N7222, N4191);
nor NOR4 (N7226, N7207, N833, N1187, N1202);
nand NAND2 (N7227, N7215, N1173);
nand NAND2 (N7228, N7219, N2285);
not NOT1 (N7229, N7221);
nor NOR3 (N7230, N7218, N1442, N52);
not NOT1 (N7231, N7226);
buf BUF1 (N7232, N7225);
and AND4 (N7233, N7230, N5475, N5906, N1486);
buf BUF1 (N7234, N7227);
and AND2 (N7235, N7231, N4589);
or OR2 (N7236, N7229, N7228);
nor NOR3 (N7237, N1052, N5227, N833);
nand NAND2 (N7238, N7214, N2531);
xor XOR2 (N7239, N7224, N4671);
xor XOR2 (N7240, N7223, N2038);
nor NOR2 (N7241, N7238, N4471);
nand NAND2 (N7242, N7240, N4314);
nand NAND4 (N7243, N7235, N4734, N6856, N2365);
xor XOR2 (N7244, N7209, N488);
not NOT1 (N7245, N7232);
buf BUF1 (N7246, N7242);
buf BUF1 (N7247, N7243);
not NOT1 (N7248, N7246);
xor XOR2 (N7249, N7247, N5174);
or OR3 (N7250, N7233, N5561, N6242);
not NOT1 (N7251, N7249);
and AND3 (N7252, N7237, N4805, N2211);
xor XOR2 (N7253, N7245, N2213);
buf BUF1 (N7254, N7251);
nor NOR3 (N7255, N7252, N6074, N4956);
or OR4 (N7256, N7234, N4174, N6530, N6728);
not NOT1 (N7257, N7250);
nor NOR4 (N7258, N7241, N4447, N4137, N1824);
and AND2 (N7259, N7244, N2150);
xor XOR2 (N7260, N7236, N529);
not NOT1 (N7261, N7258);
xor XOR2 (N7262, N7256, N1974);
or OR4 (N7263, N7262, N4545, N6373, N1578);
xor XOR2 (N7264, N7248, N6686);
or OR3 (N7265, N7261, N5934, N4820);
and AND4 (N7266, N7255, N6070, N1906, N4942);
nor NOR2 (N7267, N7259, N4838);
buf BUF1 (N7268, N7267);
not NOT1 (N7269, N7253);
not NOT1 (N7270, N7266);
and AND3 (N7271, N7269, N983, N383);
or OR2 (N7272, N7268, N5907);
xor XOR2 (N7273, N7270, N211);
nor NOR3 (N7274, N7273, N1474, N6156);
not NOT1 (N7275, N7263);
nor NOR3 (N7276, N7264, N3023, N958);
not NOT1 (N7277, N7254);
or OR4 (N7278, N7277, N4189, N1141, N4137);
or OR4 (N7279, N7275, N4446, N6038, N5381);
xor XOR2 (N7280, N7239, N4832);
and AND4 (N7281, N7260, N2186, N7033, N3691);
and AND3 (N7282, N7276, N7128, N1353);
nor NOR2 (N7283, N7257, N7184);
and AND4 (N7284, N7280, N491, N3963, N756);
buf BUF1 (N7285, N7271);
or OR2 (N7286, N7272, N6110);
buf BUF1 (N7287, N7265);
and AND3 (N7288, N7274, N6984, N255);
xor XOR2 (N7289, N7284, N2543);
nand NAND4 (N7290, N7288, N1823, N695, N6070);
xor XOR2 (N7291, N7283, N5428);
nor NOR4 (N7292, N7286, N5454, N3566, N1207);
and AND4 (N7293, N7285, N5264, N3064, N3915);
buf BUF1 (N7294, N7290);
xor XOR2 (N7295, N7292, N1199);
nor NOR4 (N7296, N7291, N1326, N2530, N3716);
xor XOR2 (N7297, N7287, N2050);
not NOT1 (N7298, N7296);
xor XOR2 (N7299, N7279, N3013);
or OR2 (N7300, N7281, N2767);
buf BUF1 (N7301, N7293);
buf BUF1 (N7302, N7301);
nor NOR2 (N7303, N7278, N3102);
not NOT1 (N7304, N7300);
and AND4 (N7305, N7299, N6140, N3199, N6179);
buf BUF1 (N7306, N7289);
xor XOR2 (N7307, N7298, N2048);
and AND2 (N7308, N7282, N4992);
not NOT1 (N7309, N7306);
xor XOR2 (N7310, N7295, N3118);
buf BUF1 (N7311, N7308);
and AND4 (N7312, N7307, N4949, N4590, N1020);
xor XOR2 (N7313, N7294, N4723);
buf BUF1 (N7314, N7309);
and AND3 (N7315, N7310, N3097, N6231);
xor XOR2 (N7316, N7313, N5342);
buf BUF1 (N7317, N7297);
and AND4 (N7318, N7314, N2434, N4114, N5903);
and AND4 (N7319, N7304, N627, N231, N2480);
nor NOR3 (N7320, N7315, N1262, N3954);
nor NOR2 (N7321, N7312, N6486);
nor NOR4 (N7322, N7319, N3121, N1567, N4717);
or OR4 (N7323, N7321, N2169, N3619, N5195);
xor XOR2 (N7324, N7323, N164);
nor NOR3 (N7325, N7320, N2799, N345);
nand NAND2 (N7326, N7302, N7317);
buf BUF1 (N7327, N3440);
not NOT1 (N7328, N7326);
nand NAND3 (N7329, N7303, N2972, N5869);
and AND4 (N7330, N7311, N4877, N2213, N4807);
or OR2 (N7331, N7316, N5730);
nand NAND3 (N7332, N7331, N6804, N810);
not NOT1 (N7333, N7318);
xor XOR2 (N7334, N7322, N4359);
and AND4 (N7335, N7334, N2573, N4122, N4226);
and AND2 (N7336, N7327, N1600);
nor NOR3 (N7337, N7305, N1470, N2858);
xor XOR2 (N7338, N7336, N5179);
and AND4 (N7339, N7335, N4312, N1010, N5303);
buf BUF1 (N7340, N7337);
xor XOR2 (N7341, N7333, N6529);
and AND2 (N7342, N7328, N5255);
or OR2 (N7343, N7332, N1728);
nand NAND4 (N7344, N7343, N4703, N915, N4535);
buf BUF1 (N7345, N7338);
xor XOR2 (N7346, N7325, N6235);
nor NOR2 (N7347, N7346, N3389);
not NOT1 (N7348, N7342);
xor XOR2 (N7349, N7347, N4529);
nor NOR2 (N7350, N7329, N4540);
nand NAND4 (N7351, N7330, N689, N6021, N3843);
xor XOR2 (N7352, N7340, N3173);
xor XOR2 (N7353, N7341, N5953);
nor NOR2 (N7354, N7349, N2903);
and AND3 (N7355, N7339, N4447, N2031);
buf BUF1 (N7356, N7353);
nor NOR3 (N7357, N7345, N6003, N6169);
nand NAND3 (N7358, N7355, N1534, N458);
and AND2 (N7359, N7348, N102);
or OR3 (N7360, N7358, N3416, N4509);
nand NAND3 (N7361, N7360, N5800, N479);
buf BUF1 (N7362, N7352);
not NOT1 (N7363, N7361);
and AND4 (N7364, N7362, N448, N2056, N460);
nor NOR2 (N7365, N7350, N6828);
nand NAND4 (N7366, N7359, N1212, N1056, N6397);
nor NOR3 (N7367, N7364, N2717, N148);
or OR4 (N7368, N7354, N7354, N3031, N1792);
and AND3 (N7369, N7366, N4299, N5956);
buf BUF1 (N7370, N7369);
and AND4 (N7371, N7370, N4735, N5666, N6968);
nor NOR4 (N7372, N7351, N4981, N5784, N7156);
and AND2 (N7373, N7367, N402);
nor NOR2 (N7374, N7357, N1703);
nor NOR4 (N7375, N7365, N6569, N5428, N6956);
not NOT1 (N7376, N7363);
nor NOR4 (N7377, N7344, N6785, N6713, N3502);
not NOT1 (N7378, N7376);
or OR2 (N7379, N7374, N2786);
or OR3 (N7380, N7377, N1993, N2798);
buf BUF1 (N7381, N7356);
buf BUF1 (N7382, N7380);
and AND3 (N7383, N7368, N6755, N5952);
buf BUF1 (N7384, N7381);
buf BUF1 (N7385, N7373);
buf BUF1 (N7386, N7382);
or OR2 (N7387, N7378, N3399);
nor NOR3 (N7388, N7324, N3662, N2275);
buf BUF1 (N7389, N7385);
and AND2 (N7390, N7383, N3659);
nand NAND4 (N7391, N7387, N315, N2375, N5463);
not NOT1 (N7392, N7384);
buf BUF1 (N7393, N7372);
nand NAND2 (N7394, N7393, N2541);
xor XOR2 (N7395, N7388, N2489);
buf BUF1 (N7396, N7391);
xor XOR2 (N7397, N7379, N946);
xor XOR2 (N7398, N7395, N537);
nand NAND2 (N7399, N7386, N2490);
xor XOR2 (N7400, N7396, N4080);
or OR2 (N7401, N7389, N2202);
xor XOR2 (N7402, N7390, N5340);
or OR2 (N7403, N7394, N2072);
or OR2 (N7404, N7403, N4092);
xor XOR2 (N7405, N7401, N285);
nand NAND4 (N7406, N7404, N6620, N6207, N1330);
nor NOR4 (N7407, N7402, N5553, N347, N3508);
or OR2 (N7408, N7398, N3333);
xor XOR2 (N7409, N7408, N3968);
buf BUF1 (N7410, N7409);
and AND3 (N7411, N7399, N1714, N5081);
nor NOR2 (N7412, N7397, N6871);
buf BUF1 (N7413, N7371);
not NOT1 (N7414, N7410);
nor NOR3 (N7415, N7375, N3402, N5961);
buf BUF1 (N7416, N7415);
not NOT1 (N7417, N7412);
xor XOR2 (N7418, N7392, N1504);
or OR3 (N7419, N7407, N4014, N45);
xor XOR2 (N7420, N7400, N1845);
nand NAND4 (N7421, N7411, N6013, N2132, N973);
not NOT1 (N7422, N7418);
buf BUF1 (N7423, N7419);
not NOT1 (N7424, N7417);
not NOT1 (N7425, N7413);
nor NOR3 (N7426, N7422, N6963, N6030);
nor NOR2 (N7427, N7426, N6863);
nor NOR3 (N7428, N7420, N3687, N3958);
buf BUF1 (N7429, N7414);
nand NAND2 (N7430, N7425, N1566);
not NOT1 (N7431, N7424);
nand NAND2 (N7432, N7428, N3853);
buf BUF1 (N7433, N7427);
buf BUF1 (N7434, N7406);
or OR4 (N7435, N7430, N1598, N5573, N6792);
or OR2 (N7436, N7416, N4900);
not NOT1 (N7437, N7423);
nor NOR4 (N7438, N7429, N79, N7061, N3944);
buf BUF1 (N7439, N7438);
or OR3 (N7440, N7439, N6499, N6640);
and AND2 (N7441, N7437, N2443);
xor XOR2 (N7442, N7432, N1521);
xor XOR2 (N7443, N7440, N7379);
buf BUF1 (N7444, N7434);
xor XOR2 (N7445, N7433, N683);
nor NOR4 (N7446, N7445, N3554, N750, N2705);
or OR3 (N7447, N7435, N4726, N3937);
nor NOR3 (N7448, N7442, N342, N5666);
xor XOR2 (N7449, N7444, N7165);
not NOT1 (N7450, N7436);
and AND3 (N7451, N7449, N7361, N7262);
not NOT1 (N7452, N7431);
or OR3 (N7453, N7446, N3680, N1537);
nand NAND4 (N7454, N7443, N3144, N5293, N2258);
not NOT1 (N7455, N7454);
xor XOR2 (N7456, N7448, N2509);
not NOT1 (N7457, N7455);
or OR4 (N7458, N7447, N3269, N5924, N2610);
nand NAND3 (N7459, N7453, N2801, N1634);
or OR2 (N7460, N7405, N6651);
and AND4 (N7461, N7458, N1100, N5463, N5648);
nand NAND2 (N7462, N7451, N1215);
nand NAND2 (N7463, N7456, N6302);
nor NOR2 (N7464, N7450, N2321);
not NOT1 (N7465, N7459);
xor XOR2 (N7466, N7460, N5273);
nand NAND4 (N7467, N7421, N1942, N5913, N2534);
buf BUF1 (N7468, N7467);
xor XOR2 (N7469, N7441, N1641);
buf BUF1 (N7470, N7464);
or OR4 (N7471, N7469, N6754, N2455, N4969);
and AND4 (N7472, N7462, N2969, N3540, N6026);
nand NAND2 (N7473, N7471, N3072);
buf BUF1 (N7474, N7457);
xor XOR2 (N7475, N7474, N4020);
or OR4 (N7476, N7470, N4122, N2219, N6573);
buf BUF1 (N7477, N7463);
nand NAND3 (N7478, N7477, N5614, N2708);
or OR2 (N7479, N7461, N5754);
or OR2 (N7480, N7466, N4136);
and AND2 (N7481, N7465, N6634);
not NOT1 (N7482, N7472);
or OR3 (N7483, N7480, N3213, N1010);
and AND2 (N7484, N7483, N1452);
buf BUF1 (N7485, N7481);
buf BUF1 (N7486, N7473);
and AND4 (N7487, N7486, N4542, N4948, N4450);
or OR4 (N7488, N7476, N5228, N6230, N5225);
not NOT1 (N7489, N7475);
buf BUF1 (N7490, N7452);
and AND2 (N7491, N7485, N7383);
nand NAND4 (N7492, N7489, N5550, N3513, N1385);
buf BUF1 (N7493, N7488);
nor NOR4 (N7494, N7492, N4002, N5524, N2300);
buf BUF1 (N7495, N7484);
buf BUF1 (N7496, N7468);
buf BUF1 (N7497, N7490);
buf BUF1 (N7498, N7495);
and AND4 (N7499, N7491, N2332, N7013, N1431);
buf BUF1 (N7500, N7496);
xor XOR2 (N7501, N7493, N3905);
buf BUF1 (N7502, N7499);
or OR3 (N7503, N7478, N58, N3886);
not NOT1 (N7504, N7502);
nand NAND3 (N7505, N7504, N470, N5401);
buf BUF1 (N7506, N7503);
nor NOR2 (N7507, N7482, N2309);
xor XOR2 (N7508, N7506, N746);
xor XOR2 (N7509, N7500, N6897);
not NOT1 (N7510, N7479);
nand NAND3 (N7511, N7487, N3800, N6181);
or OR3 (N7512, N7508, N1764, N4142);
xor XOR2 (N7513, N7497, N3672);
nand NAND3 (N7514, N7510, N346, N2001);
buf BUF1 (N7515, N7511);
nor NOR4 (N7516, N7509, N6590, N550, N6952);
xor XOR2 (N7517, N7516, N6015);
and AND2 (N7518, N7501, N3303);
buf BUF1 (N7519, N7507);
not NOT1 (N7520, N7518);
not NOT1 (N7521, N7517);
xor XOR2 (N7522, N7514, N6838);
nand NAND3 (N7523, N7519, N7311, N4323);
xor XOR2 (N7524, N7512, N2106);
nor NOR3 (N7525, N7505, N1453, N2811);
not NOT1 (N7526, N7522);
not NOT1 (N7527, N7515);
nor NOR3 (N7528, N7498, N1495, N340);
xor XOR2 (N7529, N7528, N6744);
nor NOR4 (N7530, N7521, N5879, N305, N1340);
nor NOR3 (N7531, N7529, N3733, N7252);
nand NAND2 (N7532, N7527, N1123);
or OR2 (N7533, N7494, N6679);
not NOT1 (N7534, N7513);
and AND2 (N7535, N7530, N3343);
or OR3 (N7536, N7535, N3220, N2048);
nor NOR3 (N7537, N7526, N1998, N5806);
buf BUF1 (N7538, N7536);
nor NOR3 (N7539, N7523, N4511, N7209);
and AND4 (N7540, N7538, N6503, N1191, N4291);
or OR4 (N7541, N7532, N4688, N6853, N402);
buf BUF1 (N7542, N7534);
nand NAND2 (N7543, N7533, N5898);
xor XOR2 (N7544, N7531, N4596);
xor XOR2 (N7545, N7520, N3736);
buf BUF1 (N7546, N7525);
xor XOR2 (N7547, N7537, N2721);
nor NOR4 (N7548, N7545, N2916, N988, N6430);
and AND4 (N7549, N7547, N6087, N1109, N6704);
nor NOR4 (N7550, N7544, N7386, N2850, N4012);
buf BUF1 (N7551, N7548);
nor NOR4 (N7552, N7543, N6817, N4708, N5440);
not NOT1 (N7553, N7542);
buf BUF1 (N7554, N7551);
xor XOR2 (N7555, N7553, N2770);
nand NAND3 (N7556, N7540, N6176, N5366);
xor XOR2 (N7557, N7524, N1509);
xor XOR2 (N7558, N7557, N896);
xor XOR2 (N7559, N7558, N1447);
buf BUF1 (N7560, N7539);
nor NOR2 (N7561, N7541, N2356);
not NOT1 (N7562, N7555);
and AND4 (N7563, N7552, N1106, N4434, N2695);
nand NAND3 (N7564, N7556, N1401, N5319);
not NOT1 (N7565, N7554);
and AND4 (N7566, N7564, N3692, N1878, N6410);
and AND2 (N7567, N7560, N3393);
and AND4 (N7568, N7562, N717, N4437, N5723);
buf BUF1 (N7569, N7567);
or OR2 (N7570, N7566, N1495);
xor XOR2 (N7571, N7565, N3605);
xor XOR2 (N7572, N7570, N1548);
or OR4 (N7573, N7572, N4166, N916, N374);
not NOT1 (N7574, N7561);
nor NOR3 (N7575, N7571, N2064, N2847);
xor XOR2 (N7576, N7573, N2727);
xor XOR2 (N7577, N7559, N1538);
nor NOR3 (N7578, N7576, N3958, N1511);
xor XOR2 (N7579, N7574, N1155);
and AND3 (N7580, N7579, N5286, N5935);
xor XOR2 (N7581, N7546, N6363);
nand NAND2 (N7582, N7581, N2687);
nor NOR4 (N7583, N7563, N7023, N1065, N2676);
not NOT1 (N7584, N7550);
xor XOR2 (N7585, N7583, N3320);
xor XOR2 (N7586, N7580, N5745);
xor XOR2 (N7587, N7577, N4657);
nand NAND3 (N7588, N7569, N4893, N3127);
nor NOR3 (N7589, N7587, N2163, N1995);
xor XOR2 (N7590, N7588, N141);
xor XOR2 (N7591, N7590, N6526);
and AND4 (N7592, N7584, N4617, N1160, N7518);
and AND4 (N7593, N7589, N3566, N3013, N6265);
xor XOR2 (N7594, N7591, N221);
xor XOR2 (N7595, N7592, N4309);
not NOT1 (N7596, N7585);
or OR2 (N7597, N7593, N6432);
xor XOR2 (N7598, N7582, N3627);
and AND3 (N7599, N7595, N3669, N4326);
nand NAND2 (N7600, N7578, N417);
or OR2 (N7601, N7599, N759);
nand NAND4 (N7602, N7575, N5178, N7232, N2007);
or OR4 (N7603, N7598, N2896, N2551, N7007);
nor NOR4 (N7604, N7603, N6299, N4942, N3018);
xor XOR2 (N7605, N7568, N501);
buf BUF1 (N7606, N7604);
xor XOR2 (N7607, N7600, N906);
xor XOR2 (N7608, N7605, N2349);
nor NOR3 (N7609, N7596, N2528, N7435);
or OR3 (N7610, N7602, N4077, N7246);
or OR4 (N7611, N7610, N2112, N6246, N4236);
nor NOR3 (N7612, N7606, N3270, N1320);
or OR3 (N7613, N7586, N394, N5124);
not NOT1 (N7614, N7594);
nand NAND2 (N7615, N7549, N3647);
xor XOR2 (N7616, N7615, N2299);
xor XOR2 (N7617, N7611, N5236);
not NOT1 (N7618, N7601);
xor XOR2 (N7619, N7612, N6524);
or OR2 (N7620, N7618, N66);
and AND3 (N7621, N7597, N5437, N3637);
not NOT1 (N7622, N7620);
not NOT1 (N7623, N7621);
or OR2 (N7624, N7617, N4683);
buf BUF1 (N7625, N7613);
or OR3 (N7626, N7623, N5007, N855);
or OR4 (N7627, N7622, N5772, N7466, N3868);
or OR4 (N7628, N7614, N6381, N2749, N7356);
nand NAND2 (N7629, N7619, N6160);
xor XOR2 (N7630, N7624, N2308);
not NOT1 (N7631, N7628);
buf BUF1 (N7632, N7608);
and AND4 (N7633, N7629, N3969, N6842, N1523);
not NOT1 (N7634, N7632);
or OR4 (N7635, N7607, N4873, N5370, N7155);
buf BUF1 (N7636, N7625);
nand NAND4 (N7637, N7630, N1746, N3858, N2988);
xor XOR2 (N7638, N7634, N2798);
buf BUF1 (N7639, N7635);
and AND3 (N7640, N7609, N4702, N4454);
and AND2 (N7641, N7633, N5341);
not NOT1 (N7642, N7631);
and AND3 (N7643, N7627, N3130, N1753);
nor NOR3 (N7644, N7639, N6221, N1834);
buf BUF1 (N7645, N7641);
and AND4 (N7646, N7645, N2085, N6415, N7134);
and AND3 (N7647, N7646, N826, N7359);
and AND2 (N7648, N7642, N5390);
nand NAND4 (N7649, N7648, N5272, N2844, N2715);
or OR2 (N7650, N7626, N3390);
xor XOR2 (N7651, N7636, N4150);
buf BUF1 (N7652, N7650);
nor NOR3 (N7653, N7638, N3655, N5770);
not NOT1 (N7654, N7649);
or OR4 (N7655, N7654, N6476, N6282, N626);
nand NAND4 (N7656, N7637, N2789, N7295, N4494);
nor NOR2 (N7657, N7653, N170);
buf BUF1 (N7658, N7657);
not NOT1 (N7659, N7656);
buf BUF1 (N7660, N7655);
buf BUF1 (N7661, N7643);
and AND3 (N7662, N7660, N1698, N2669);
or OR3 (N7663, N7647, N1243, N3105);
buf BUF1 (N7664, N7640);
nor NOR2 (N7665, N7652, N1828);
nand NAND2 (N7666, N7658, N5950);
or OR2 (N7667, N7644, N7376);
buf BUF1 (N7668, N7616);
nand NAND2 (N7669, N7663, N3340);
nor NOR4 (N7670, N7662, N4416, N4724, N7125);
buf BUF1 (N7671, N7667);
nor NOR3 (N7672, N7659, N1996, N6132);
not NOT1 (N7673, N7672);
nor NOR3 (N7674, N7668, N7396, N2801);
xor XOR2 (N7675, N7661, N6445);
nand NAND2 (N7676, N7674, N7594);
buf BUF1 (N7677, N7665);
or OR4 (N7678, N7677, N6840, N773, N2402);
not NOT1 (N7679, N7675);
and AND4 (N7680, N7678, N4804, N1363, N2746);
nand NAND2 (N7681, N7673, N4375);
not NOT1 (N7682, N7681);
xor XOR2 (N7683, N7682, N704);
nor NOR3 (N7684, N7671, N408, N2506);
and AND3 (N7685, N7679, N7139, N7373);
or OR4 (N7686, N7670, N24, N4269, N7098);
and AND3 (N7687, N7684, N6706, N5127);
or OR4 (N7688, N7683, N2703, N824, N799);
not NOT1 (N7689, N7676);
nor NOR2 (N7690, N7669, N5889);
and AND2 (N7691, N7689, N3971);
buf BUF1 (N7692, N7664);
xor XOR2 (N7693, N7651, N1311);
nor NOR3 (N7694, N7686, N539, N862);
and AND4 (N7695, N7690, N2120, N1613, N5629);
not NOT1 (N7696, N7692);
not NOT1 (N7697, N7695);
nor NOR4 (N7698, N7666, N5441, N2834, N1431);
nand NAND4 (N7699, N7697, N2861, N3645, N6781);
nor NOR2 (N7700, N7688, N3348);
buf BUF1 (N7701, N7694);
nand NAND3 (N7702, N7693, N4937, N7460);
or OR2 (N7703, N7702, N6404);
or OR2 (N7704, N7696, N2100);
nor NOR2 (N7705, N7680, N5333);
buf BUF1 (N7706, N7685);
buf BUF1 (N7707, N7699);
buf BUF1 (N7708, N7705);
buf BUF1 (N7709, N7701);
nor NOR3 (N7710, N7698, N6140, N3386);
not NOT1 (N7711, N7704);
nor NOR4 (N7712, N7709, N1213, N6111, N1452);
xor XOR2 (N7713, N7710, N871);
or OR4 (N7714, N7700, N4946, N5480, N1968);
buf BUF1 (N7715, N7707);
nand NAND2 (N7716, N7714, N3098);
nand NAND2 (N7717, N7703, N2686);
not NOT1 (N7718, N7708);
and AND2 (N7719, N7711, N2202);
not NOT1 (N7720, N7717);
or OR3 (N7721, N7720, N5683, N2652);
nor NOR3 (N7722, N7718, N6171, N3425);
not NOT1 (N7723, N7706);
xor XOR2 (N7724, N7719, N6804);
xor XOR2 (N7725, N7723, N3371);
not NOT1 (N7726, N7713);
nand NAND4 (N7727, N7725, N4592, N3154, N2108);
not NOT1 (N7728, N7724);
and AND4 (N7729, N7728, N4512, N578, N4060);
or OR3 (N7730, N7712, N3941, N5865);
xor XOR2 (N7731, N7715, N537);
nand NAND4 (N7732, N7730, N1513, N4549, N3155);
nand NAND3 (N7733, N7691, N4259, N2498);
or OR3 (N7734, N7727, N1148, N5480);
nor NOR3 (N7735, N7687, N3126, N1658);
or OR3 (N7736, N7731, N2718, N4957);
buf BUF1 (N7737, N7722);
nand NAND4 (N7738, N7736, N823, N3410, N6021);
nand NAND2 (N7739, N7734, N7548);
nor NOR2 (N7740, N7739, N4261);
xor XOR2 (N7741, N7735, N6011);
and AND2 (N7742, N7738, N7111);
nand NAND3 (N7743, N7729, N4337, N5954);
and AND3 (N7744, N7742, N398, N3275);
buf BUF1 (N7745, N7744);
nand NAND4 (N7746, N7743, N5148, N5311, N1328);
nand NAND4 (N7747, N7721, N1324, N4458, N6596);
nor NOR4 (N7748, N7733, N5535, N1023, N5997);
buf BUF1 (N7749, N7740);
not NOT1 (N7750, N7748);
not NOT1 (N7751, N7741);
and AND3 (N7752, N7732, N1141, N2074);
and AND3 (N7753, N7751, N2692, N1954);
not NOT1 (N7754, N7716);
and AND2 (N7755, N7753, N2719);
nor NOR3 (N7756, N7726, N3617, N2546);
not NOT1 (N7757, N7754);
xor XOR2 (N7758, N7745, N1426);
nor NOR2 (N7759, N7758, N5961);
and AND4 (N7760, N7750, N740, N7008, N3212);
not NOT1 (N7761, N7756);
nor NOR2 (N7762, N7737, N5804);
nor NOR2 (N7763, N7752, N2168);
xor XOR2 (N7764, N7760, N7537);
nand NAND4 (N7765, N7764, N3453, N7609, N3016);
buf BUF1 (N7766, N7747);
not NOT1 (N7767, N7759);
not NOT1 (N7768, N7767);
xor XOR2 (N7769, N7766, N5669);
nand NAND2 (N7770, N7762, N2022);
nor NOR2 (N7771, N7770, N4502);
buf BUF1 (N7772, N7761);
xor XOR2 (N7773, N7757, N4718);
or OR4 (N7774, N7765, N1961, N5154, N6650);
buf BUF1 (N7775, N7773);
or OR4 (N7776, N7769, N4450, N4729, N1704);
buf BUF1 (N7777, N7768);
not NOT1 (N7778, N7755);
not NOT1 (N7779, N7763);
nand NAND4 (N7780, N7746, N475, N64, N4858);
not NOT1 (N7781, N7780);
xor XOR2 (N7782, N7774, N2028);
xor XOR2 (N7783, N7775, N428);
xor XOR2 (N7784, N7749, N1725);
not NOT1 (N7785, N7778);
not NOT1 (N7786, N7784);
nand NAND2 (N7787, N7772, N5142);
xor XOR2 (N7788, N7779, N479);
buf BUF1 (N7789, N7786);
and AND4 (N7790, N7777, N523, N721, N3451);
not NOT1 (N7791, N7789);
and AND2 (N7792, N7782, N3709);
buf BUF1 (N7793, N7771);
buf BUF1 (N7794, N7787);
nand NAND4 (N7795, N7791, N3474, N6257, N3777);
nor NOR3 (N7796, N7794, N2896, N5088);
buf BUF1 (N7797, N7781);
or OR3 (N7798, N7796, N3133, N4455);
or OR4 (N7799, N7798, N7150, N6660, N3115);
and AND4 (N7800, N7788, N1323, N2758, N389);
nand NAND2 (N7801, N7797, N3951);
and AND3 (N7802, N7793, N1242, N4621);
nand NAND4 (N7803, N7795, N96, N3042, N6593);
and AND2 (N7804, N7776, N6638);
xor XOR2 (N7805, N7802, N2975);
buf BUF1 (N7806, N7792);
and AND2 (N7807, N7801, N3391);
buf BUF1 (N7808, N7806);
not NOT1 (N7809, N7805);
xor XOR2 (N7810, N7809, N2409);
or OR2 (N7811, N7800, N1310);
nand NAND4 (N7812, N7811, N1645, N1221, N2253);
not NOT1 (N7813, N7803);
nor NOR4 (N7814, N7804, N2229, N4250, N1470);
xor XOR2 (N7815, N7814, N1554);
not NOT1 (N7816, N7810);
xor XOR2 (N7817, N7812, N7327);
xor XOR2 (N7818, N7790, N2893);
nand NAND4 (N7819, N7785, N6257, N1127, N6706);
buf BUF1 (N7820, N7799);
and AND2 (N7821, N7808, N1347);
buf BUF1 (N7822, N7820);
not NOT1 (N7823, N7807);
buf BUF1 (N7824, N7823);
xor XOR2 (N7825, N7815, N7477);
xor XOR2 (N7826, N7819, N1918);
nand NAND4 (N7827, N7824, N4176, N789, N2865);
and AND4 (N7828, N7825, N5437, N1065, N3089);
buf BUF1 (N7829, N7817);
xor XOR2 (N7830, N7828, N4836);
not NOT1 (N7831, N7818);
nor NOR4 (N7832, N7826, N2318, N7551, N1115);
or OR4 (N7833, N7829, N2412, N2567, N7109);
not NOT1 (N7834, N7821);
not NOT1 (N7835, N7833);
not NOT1 (N7836, N7831);
nor NOR2 (N7837, N7827, N5333);
buf BUF1 (N7838, N7813);
buf BUF1 (N7839, N7832);
nor NOR4 (N7840, N7836, N6180, N7739, N2995);
buf BUF1 (N7841, N7835);
nor NOR3 (N7842, N7837, N5748, N7176);
or OR2 (N7843, N7830, N1507);
nor NOR2 (N7844, N7822, N7073);
or OR4 (N7845, N7816, N7738, N853, N4056);
or OR3 (N7846, N7841, N6182, N6506);
xor XOR2 (N7847, N7845, N5811);
or OR2 (N7848, N7842, N2446);
not NOT1 (N7849, N7838);
xor XOR2 (N7850, N7846, N6808);
or OR3 (N7851, N7840, N151, N6488);
and AND4 (N7852, N7849, N6032, N3438, N2624);
or OR4 (N7853, N7834, N2407, N2729, N4685);
nand NAND3 (N7854, N7843, N5322, N4506);
xor XOR2 (N7855, N7844, N3071);
xor XOR2 (N7856, N7783, N863);
nand NAND4 (N7857, N7855, N7741, N6438, N7081);
not NOT1 (N7858, N7856);
nand NAND4 (N7859, N7850, N6422, N2614, N1318);
xor XOR2 (N7860, N7857, N4167);
xor XOR2 (N7861, N7859, N5672);
not NOT1 (N7862, N7839);
nand NAND3 (N7863, N7853, N50, N370);
nand NAND2 (N7864, N7852, N6312);
xor XOR2 (N7865, N7860, N6488);
not NOT1 (N7866, N7854);
and AND2 (N7867, N7848, N769);
or OR2 (N7868, N7867, N1244);
nand NAND2 (N7869, N7864, N7483);
buf BUF1 (N7870, N7861);
not NOT1 (N7871, N7863);
not NOT1 (N7872, N7871);
xor XOR2 (N7873, N7858, N4277);
xor XOR2 (N7874, N7869, N6729);
nand NAND4 (N7875, N7851, N7216, N3853, N4286);
not NOT1 (N7876, N7866);
not NOT1 (N7877, N7876);
and AND2 (N7878, N7875, N758);
nand NAND4 (N7879, N7862, N1113, N3439, N4239);
buf BUF1 (N7880, N7847);
not NOT1 (N7881, N7872);
and AND2 (N7882, N7881, N4851);
nor NOR2 (N7883, N7874, N6664);
xor XOR2 (N7884, N7873, N1539);
buf BUF1 (N7885, N7870);
and AND4 (N7886, N7877, N2040, N355, N3211);
not NOT1 (N7887, N7882);
buf BUF1 (N7888, N7884);
not NOT1 (N7889, N7885);
and AND3 (N7890, N7880, N1537, N5414);
xor XOR2 (N7891, N7888, N1555);
or OR3 (N7892, N7886, N2992, N596);
buf BUF1 (N7893, N7879);
not NOT1 (N7894, N7891);
not NOT1 (N7895, N7892);
or OR3 (N7896, N7868, N1570, N5932);
nand NAND3 (N7897, N7878, N664, N6649);
nand NAND2 (N7898, N7893, N6793);
and AND2 (N7899, N7890, N6100);
buf BUF1 (N7900, N7898);
nand NAND3 (N7901, N7899, N3745, N6431);
buf BUF1 (N7902, N7889);
or OR2 (N7903, N7896, N608);
or OR4 (N7904, N7900, N2445, N5691, N7656);
not NOT1 (N7905, N7902);
or OR3 (N7906, N7904, N5372, N7789);
or OR2 (N7907, N7865, N6545);
nor NOR2 (N7908, N7903, N7290);
and AND2 (N7909, N7906, N2882);
or OR3 (N7910, N7897, N6202, N3740);
nand NAND2 (N7911, N7883, N792);
buf BUF1 (N7912, N7905);
or OR3 (N7913, N7909, N6190, N3994);
buf BUF1 (N7914, N7910);
buf BUF1 (N7915, N7894);
not NOT1 (N7916, N7912);
or OR4 (N7917, N7911, N3268, N5089, N6654);
nand NAND3 (N7918, N7917, N4637, N3780);
nor NOR3 (N7919, N7908, N6271, N6353);
buf BUF1 (N7920, N7914);
xor XOR2 (N7921, N7920, N7416);
or OR4 (N7922, N7921, N5993, N7747, N3858);
or OR4 (N7923, N7901, N2265, N6253, N837);
or OR4 (N7924, N7923, N2878, N1082, N7612);
xor XOR2 (N7925, N7887, N4734);
or OR2 (N7926, N7907, N6129);
xor XOR2 (N7927, N7924, N7449);
and AND3 (N7928, N7895, N1206, N6283);
buf BUF1 (N7929, N7919);
nor NOR3 (N7930, N7929, N2643, N426);
nand NAND4 (N7931, N7925, N3792, N7545, N4182);
buf BUF1 (N7932, N7926);
nand NAND2 (N7933, N7915, N3733);
and AND2 (N7934, N7930, N5617);
buf BUF1 (N7935, N7922);
buf BUF1 (N7936, N7927);
buf BUF1 (N7937, N7931);
nand NAND3 (N7938, N7937, N4133, N6399);
buf BUF1 (N7939, N7918);
not NOT1 (N7940, N7932);
or OR3 (N7941, N7933, N5615, N5784);
nor NOR3 (N7942, N7935, N2185, N5953);
and AND3 (N7943, N7941, N783, N1110);
nand NAND2 (N7944, N7939, N5358);
or OR4 (N7945, N7934, N6640, N6958, N3389);
xor XOR2 (N7946, N7938, N3916);
nand NAND4 (N7947, N7928, N4287, N5723, N3524);
nand NAND2 (N7948, N7916, N858);
or OR2 (N7949, N7936, N626);
and AND2 (N7950, N7943, N6107);
and AND3 (N7951, N7946, N3016, N4348);
nand NAND3 (N7952, N7947, N6404, N142);
and AND2 (N7953, N7944, N5311);
nand NAND3 (N7954, N7942, N2135, N7353);
xor XOR2 (N7955, N7952, N1736);
or OR4 (N7956, N7948, N286, N649, N1675);
or OR2 (N7957, N7955, N3779);
nand NAND4 (N7958, N7951, N5646, N5077, N135);
nand NAND2 (N7959, N7953, N6411);
or OR3 (N7960, N7956, N5238, N6388);
nor NOR4 (N7961, N7949, N1921, N6029, N4299);
or OR2 (N7962, N7945, N5189);
xor XOR2 (N7963, N7962, N6044);
buf BUF1 (N7964, N7940);
nor NOR2 (N7965, N7964, N5734);
nand NAND2 (N7966, N7960, N7534);
not NOT1 (N7967, N7966);
nand NAND2 (N7968, N7958, N4344);
nor NOR4 (N7969, N7950, N1881, N2878, N2312);
xor XOR2 (N7970, N7954, N6025);
nand NAND2 (N7971, N7959, N2615);
or OR4 (N7972, N7971, N6894, N5550, N1482);
or OR3 (N7973, N7957, N7880, N4804);
buf BUF1 (N7974, N7913);
xor XOR2 (N7975, N7974, N322);
not NOT1 (N7976, N7969);
nand NAND2 (N7977, N7975, N5562);
xor XOR2 (N7978, N7961, N3863);
nand NAND3 (N7979, N7967, N1939, N3486);
nand NAND2 (N7980, N7965, N3986);
nor NOR2 (N7981, N7970, N778);
nand NAND4 (N7982, N7973, N881, N2235, N588);
buf BUF1 (N7983, N7968);
or OR3 (N7984, N7980, N2993, N7352);
or OR4 (N7985, N7978, N1212, N6488, N1943);
xor XOR2 (N7986, N7982, N7277);
not NOT1 (N7987, N7981);
not NOT1 (N7988, N7976);
or OR4 (N7989, N7987, N5542, N2312, N6295);
not NOT1 (N7990, N7977);
not NOT1 (N7991, N7979);
xor XOR2 (N7992, N7972, N782);
nand NAND2 (N7993, N7990, N6500);
nand NAND4 (N7994, N7986, N719, N677, N5476);
buf BUF1 (N7995, N7963);
or OR4 (N7996, N7985, N6006, N6118, N1152);
nand NAND3 (N7997, N7993, N2375, N3470);
nand NAND2 (N7998, N7994, N5247);
not NOT1 (N7999, N7996);
and AND3 (N8000, N7991, N3322, N3216);
buf BUF1 (N8001, N7997);
not NOT1 (N8002, N7984);
buf BUF1 (N8003, N7983);
not NOT1 (N8004, N7989);
xor XOR2 (N8005, N8000, N6118);
and AND4 (N8006, N8005, N1701, N4225, N5817);
or OR4 (N8007, N7998, N6574, N7859, N6353);
buf BUF1 (N8008, N8004);
and AND3 (N8009, N8003, N6947, N7616);
nor NOR2 (N8010, N8006, N2952);
nor NOR4 (N8011, N7995, N2054, N7498, N5726);
nor NOR2 (N8012, N8001, N1274);
nor NOR2 (N8013, N8010, N6412);
not NOT1 (N8014, N8007);
xor XOR2 (N8015, N8014, N3478);
buf BUF1 (N8016, N7992);
xor XOR2 (N8017, N8012, N5029);
not NOT1 (N8018, N7988);
not NOT1 (N8019, N8017);
and AND2 (N8020, N8015, N1687);
not NOT1 (N8021, N7999);
nand NAND2 (N8022, N8013, N1258);
buf BUF1 (N8023, N8009);
or OR4 (N8024, N8021, N5240, N8002, N2139);
buf BUF1 (N8025, N1725);
buf BUF1 (N8026, N8024);
and AND3 (N8027, N8023, N531, N3162);
and AND2 (N8028, N8016, N4069);
nand NAND2 (N8029, N8026, N1640);
buf BUF1 (N8030, N8019);
buf BUF1 (N8031, N8028);
not NOT1 (N8032, N8018);
and AND4 (N8033, N8029, N5296, N4388, N1506);
not NOT1 (N8034, N8032);
and AND4 (N8035, N8033, N1322, N4293, N5262);
xor XOR2 (N8036, N8025, N754);
nor NOR4 (N8037, N8022, N1982, N3907, N1914);
not NOT1 (N8038, N8034);
or OR3 (N8039, N8030, N645, N2751);
buf BUF1 (N8040, N8035);
or OR3 (N8041, N8008, N5526, N6056);
nor NOR4 (N8042, N8020, N6971, N1142, N5633);
xor XOR2 (N8043, N8037, N6144);
or OR3 (N8044, N8041, N2492, N1734);
not NOT1 (N8045, N8031);
not NOT1 (N8046, N8040);
or OR3 (N8047, N8042, N2549, N1924);
not NOT1 (N8048, N8047);
and AND3 (N8049, N8039, N5079, N7164);
buf BUF1 (N8050, N8046);
nand NAND3 (N8051, N8050, N7127, N6531);
buf BUF1 (N8052, N8044);
or OR4 (N8053, N8048, N6614, N2345, N6416);
or OR3 (N8054, N8011, N3795, N4523);
xor XOR2 (N8055, N8053, N3939);
nor NOR4 (N8056, N8051, N7235, N599, N6884);
nor NOR3 (N8057, N8056, N6961, N3506);
or OR3 (N8058, N8043, N6348, N7167);
and AND4 (N8059, N8052, N4136, N7877, N3933);
xor XOR2 (N8060, N8058, N321);
buf BUF1 (N8061, N8054);
buf BUF1 (N8062, N8027);
nand NAND3 (N8063, N8045, N6467, N4889);
or OR4 (N8064, N8061, N1991, N2869, N628);
and AND4 (N8065, N8038, N2027, N4085, N122);
nor NOR2 (N8066, N8057, N3405);
or OR3 (N8067, N8059, N1391, N1970);
not NOT1 (N8068, N8062);
nor NOR2 (N8069, N8065, N5130);
buf BUF1 (N8070, N8068);
not NOT1 (N8071, N8064);
not NOT1 (N8072, N8070);
xor XOR2 (N8073, N8055, N5730);
xor XOR2 (N8074, N8069, N411);
buf BUF1 (N8075, N8067);
and AND4 (N8076, N8074, N2595, N5984, N2885);
xor XOR2 (N8077, N8076, N5893);
buf BUF1 (N8078, N8072);
xor XOR2 (N8079, N8036, N2924);
nand NAND4 (N8080, N8063, N6152, N3234, N2008);
buf BUF1 (N8081, N8078);
xor XOR2 (N8082, N8073, N2775);
and AND4 (N8083, N8080, N5840, N4296, N5742);
and AND4 (N8084, N8077, N1824, N408, N7452);
or OR2 (N8085, N8083, N3778);
nand NAND4 (N8086, N8060, N7406, N6416, N6989);
or OR2 (N8087, N8082, N7391);
buf BUF1 (N8088, N8081);
nand NAND3 (N8089, N8084, N664, N5024);
not NOT1 (N8090, N8049);
nor NOR4 (N8091, N8079, N2485, N7058, N5339);
and AND2 (N8092, N8086, N7848);
not NOT1 (N8093, N8066);
buf BUF1 (N8094, N8093);
buf BUF1 (N8095, N8087);
or OR2 (N8096, N8092, N1575);
not NOT1 (N8097, N8089);
not NOT1 (N8098, N8075);
and AND3 (N8099, N8096, N7372, N1563);
not NOT1 (N8100, N8085);
or OR4 (N8101, N8097, N3242, N5552, N4920);
or OR2 (N8102, N8101, N3101);
buf BUF1 (N8103, N8090);
not NOT1 (N8104, N8091);
or OR2 (N8105, N8094, N450);
or OR2 (N8106, N8104, N728);
not NOT1 (N8107, N8102);
nor NOR3 (N8108, N8100, N38, N2988);
nand NAND3 (N8109, N8088, N855, N8089);
not NOT1 (N8110, N8105);
nand NAND3 (N8111, N8108, N5602, N2803);
and AND4 (N8112, N8106, N4940, N7808, N3999);
xor XOR2 (N8113, N8107, N2539);
or OR2 (N8114, N8098, N6765);
not NOT1 (N8115, N8114);
nand NAND3 (N8116, N8112, N5757, N1468);
nand NAND3 (N8117, N8116, N1324, N5927);
xor XOR2 (N8118, N8110, N6879);
nor NOR3 (N8119, N8117, N2629, N3324);
xor XOR2 (N8120, N8115, N2289);
xor XOR2 (N8121, N8103, N3911);
or OR4 (N8122, N8121, N5358, N7458, N1443);
and AND2 (N8123, N8099, N2915);
and AND4 (N8124, N8111, N997, N4010, N904);
buf BUF1 (N8125, N8119);
nand NAND4 (N8126, N8120, N5031, N4771, N6541);
not NOT1 (N8127, N8095);
nand NAND4 (N8128, N8127, N6014, N7844, N6034);
buf BUF1 (N8129, N8125);
buf BUF1 (N8130, N8113);
not NOT1 (N8131, N8123);
or OR4 (N8132, N8118, N7078, N6544, N3966);
buf BUF1 (N8133, N8129);
not NOT1 (N8134, N8128);
not NOT1 (N8135, N8124);
or OR2 (N8136, N8071, N4169);
or OR3 (N8137, N8134, N8003, N5219);
and AND4 (N8138, N8135, N1624, N2208, N6221);
and AND2 (N8139, N8137, N5829);
or OR3 (N8140, N8122, N885, N4112);
nor NOR4 (N8141, N8140, N304, N4937, N6305);
not NOT1 (N8142, N8131);
nor NOR2 (N8143, N8139, N2982);
nor NOR3 (N8144, N8132, N4257, N1542);
nand NAND4 (N8145, N8130, N4169, N3414, N2149);
and AND3 (N8146, N8126, N2523, N3451);
nor NOR2 (N8147, N8141, N4251);
xor XOR2 (N8148, N8138, N4763);
not NOT1 (N8149, N8133);
xor XOR2 (N8150, N8136, N2070);
buf BUF1 (N8151, N8148);
xor XOR2 (N8152, N8143, N3336);
nand NAND3 (N8153, N8109, N4734, N557);
and AND3 (N8154, N8151, N3378, N2486);
buf BUF1 (N8155, N8149);
not NOT1 (N8156, N8154);
nor NOR4 (N8157, N8156, N5551, N3534, N738);
not NOT1 (N8158, N8150);
buf BUF1 (N8159, N8155);
buf BUF1 (N8160, N8159);
nand NAND4 (N8161, N8157, N5752, N5889, N6290);
and AND3 (N8162, N8146, N7161, N8027);
and AND4 (N8163, N8161, N7205, N1829, N940);
nor NOR4 (N8164, N8144, N1697, N2118, N2547);
or OR2 (N8165, N8163, N4598);
or OR3 (N8166, N8165, N521, N906);
or OR3 (N8167, N8152, N2281, N4868);
buf BUF1 (N8168, N8166);
or OR2 (N8169, N8145, N2849);
nor NOR2 (N8170, N8162, N7754);
or OR3 (N8171, N8142, N7238, N4805);
buf BUF1 (N8172, N8153);
nand NAND2 (N8173, N8169, N983);
buf BUF1 (N8174, N8171);
nor NOR2 (N8175, N8147, N6649);
nand NAND4 (N8176, N8175, N6051, N3595, N6845);
and AND3 (N8177, N8168, N407, N6827);
or OR2 (N8178, N8160, N252);
and AND3 (N8179, N8164, N2572, N3513);
or OR4 (N8180, N8179, N5689, N2716, N4836);
xor XOR2 (N8181, N8170, N5435);
nand NAND2 (N8182, N8176, N2188);
buf BUF1 (N8183, N8158);
or OR2 (N8184, N8174, N5089);
nor NOR2 (N8185, N8177, N1763);
or OR2 (N8186, N8183, N4105);
xor XOR2 (N8187, N8180, N5811);
not NOT1 (N8188, N8185);
nor NOR2 (N8189, N8181, N6938);
xor XOR2 (N8190, N8189, N3285);
buf BUF1 (N8191, N8178);
nor NOR2 (N8192, N8188, N1857);
xor XOR2 (N8193, N8184, N4927);
xor XOR2 (N8194, N8191, N4309);
not NOT1 (N8195, N8172);
buf BUF1 (N8196, N8187);
nor NOR4 (N8197, N8194, N3044, N1151, N727);
and AND3 (N8198, N8192, N36, N6330);
not NOT1 (N8199, N8198);
and AND2 (N8200, N8196, N2655);
xor XOR2 (N8201, N8195, N5915);
nand NAND4 (N8202, N8201, N1624, N4607, N834);
and AND3 (N8203, N8200, N4729, N1851);
and AND2 (N8204, N8199, N597);
buf BUF1 (N8205, N8186);
or OR4 (N8206, N8205, N7065, N2226, N2009);
or OR3 (N8207, N8203, N8166, N837);
not NOT1 (N8208, N8204);
not NOT1 (N8209, N8173);
buf BUF1 (N8210, N8193);
xor XOR2 (N8211, N8206, N6724);
buf BUF1 (N8212, N8209);
and AND2 (N8213, N8210, N1839);
xor XOR2 (N8214, N8208, N4704);
xor XOR2 (N8215, N8202, N3948);
not NOT1 (N8216, N8182);
not NOT1 (N8217, N8197);
and AND2 (N8218, N8215, N4345);
buf BUF1 (N8219, N8216);
or OR2 (N8220, N8211, N1835);
nor NOR2 (N8221, N8207, N7315);
nor NOR2 (N8222, N8213, N966);
xor XOR2 (N8223, N8219, N3818);
nor NOR3 (N8224, N8223, N4997, N1737);
buf BUF1 (N8225, N8190);
or OR4 (N8226, N8212, N1918, N7074, N3001);
buf BUF1 (N8227, N8167);
or OR4 (N8228, N8220, N4322, N4374, N4318);
buf BUF1 (N8229, N8225);
buf BUF1 (N8230, N8227);
nand NAND2 (N8231, N8229, N2322);
or OR4 (N8232, N8221, N765, N6702, N7250);
nor NOR4 (N8233, N8217, N6138, N10, N6063);
and AND3 (N8234, N8218, N6699, N441);
or OR4 (N8235, N8232, N3483, N3155, N1575);
and AND3 (N8236, N8222, N7601, N4816);
not NOT1 (N8237, N8233);
and AND2 (N8238, N8230, N4520);
and AND3 (N8239, N8228, N5854, N2283);
not NOT1 (N8240, N8238);
and AND2 (N8241, N8224, N4678);
buf BUF1 (N8242, N8226);
nand NAND4 (N8243, N8236, N6779, N6787, N6778);
not NOT1 (N8244, N8243);
and AND4 (N8245, N8241, N3285, N7949, N362);
or OR2 (N8246, N8239, N2744);
nor NOR3 (N8247, N8244, N7092, N1741);
buf BUF1 (N8248, N8235);
nor NOR4 (N8249, N8214, N4408, N8177, N7538);
or OR4 (N8250, N8231, N8220, N1700, N4561);
and AND2 (N8251, N8242, N7642);
not NOT1 (N8252, N8240);
buf BUF1 (N8253, N8245);
and AND2 (N8254, N8250, N7247);
nor NOR4 (N8255, N8234, N1183, N1564, N3891);
buf BUF1 (N8256, N8248);
and AND2 (N8257, N8252, N3185);
or OR4 (N8258, N8247, N4572, N2574, N1215);
not NOT1 (N8259, N8257);
buf BUF1 (N8260, N8254);
nand NAND4 (N8261, N8260, N7561, N3766, N5708);
not NOT1 (N8262, N8251);
xor XOR2 (N8263, N8261, N7758);
not NOT1 (N8264, N8237);
nand NAND3 (N8265, N8262, N5536, N682);
or OR2 (N8266, N8263, N3557);
xor XOR2 (N8267, N8246, N1393);
or OR2 (N8268, N8256, N7752);
nand NAND4 (N8269, N8267, N4446, N1881, N1442);
or OR3 (N8270, N8264, N4673, N4935);
not NOT1 (N8271, N8255);
nor NOR2 (N8272, N8270, N3582);
or OR3 (N8273, N8272, N2351, N3033);
xor XOR2 (N8274, N8249, N7054);
buf BUF1 (N8275, N8269);
xor XOR2 (N8276, N8266, N2007);
nor NOR4 (N8277, N8259, N807, N4486, N2968);
nor NOR4 (N8278, N8271, N4910, N7896, N3244);
buf BUF1 (N8279, N8258);
not NOT1 (N8280, N8274);
or OR2 (N8281, N8253, N602);
nand NAND4 (N8282, N8265, N8088, N4817, N5623);
nand NAND2 (N8283, N8281, N130);
nand NAND4 (N8284, N8283, N3424, N4813, N535);
nor NOR4 (N8285, N8275, N6317, N2129, N1029);
nor NOR2 (N8286, N8278, N6756);
buf BUF1 (N8287, N8276);
not NOT1 (N8288, N8282);
xor XOR2 (N8289, N8268, N904);
or OR4 (N8290, N8280, N2020, N4891, N4878);
not NOT1 (N8291, N8289);
buf BUF1 (N8292, N8273);
and AND2 (N8293, N8277, N2464);
not NOT1 (N8294, N8291);
or OR3 (N8295, N8286, N6801, N7180);
buf BUF1 (N8296, N8292);
nor NOR3 (N8297, N8285, N5433, N830);
nor NOR2 (N8298, N8288, N2573);
nor NOR3 (N8299, N8294, N419, N819);
or OR2 (N8300, N8295, N7482);
or OR4 (N8301, N8279, N2060, N1240, N591);
not NOT1 (N8302, N8296);
nand NAND3 (N8303, N8297, N2847, N6746);
xor XOR2 (N8304, N8293, N7205);
or OR2 (N8305, N8300, N1062);
not NOT1 (N8306, N8284);
or OR3 (N8307, N8302, N7672, N2819);
nand NAND2 (N8308, N8290, N2736);
xor XOR2 (N8309, N8304, N5038);
nand NAND3 (N8310, N8308, N5271, N3923);
not NOT1 (N8311, N8306);
xor XOR2 (N8312, N8310, N7829);
nor NOR2 (N8313, N8307, N1256);
nor NOR4 (N8314, N8312, N1749, N5295, N7938);
and AND2 (N8315, N8303, N3776);
or OR2 (N8316, N8299, N1994);
not NOT1 (N8317, N8309);
buf BUF1 (N8318, N8314);
nor NOR4 (N8319, N8298, N4792, N1252, N7458);
and AND4 (N8320, N8315, N6676, N4626, N4864);
not NOT1 (N8321, N8305);
xor XOR2 (N8322, N8287, N4799);
xor XOR2 (N8323, N8311, N690);
nand NAND3 (N8324, N8301, N4132, N2146);
buf BUF1 (N8325, N8324);
or OR2 (N8326, N8313, N873);
xor XOR2 (N8327, N8323, N662);
and AND2 (N8328, N8316, N6253);
and AND2 (N8329, N8319, N123);
nor NOR2 (N8330, N8325, N5309);
and AND4 (N8331, N8321, N4192, N5989, N828);
buf BUF1 (N8332, N8318);
not NOT1 (N8333, N8331);
and AND2 (N8334, N8317, N1211);
nand NAND3 (N8335, N8333, N5794, N3476);
or OR4 (N8336, N8328, N1515, N1807, N5427);
nor NOR3 (N8337, N8336, N7119, N4405);
nor NOR2 (N8338, N8320, N3183);
or OR2 (N8339, N8327, N2773);
and AND2 (N8340, N8337, N8260);
nand NAND2 (N8341, N8329, N8267);
buf BUF1 (N8342, N8332);
nor NOR4 (N8343, N8340, N5541, N1126, N1882);
or OR3 (N8344, N8334, N5948, N2684);
and AND4 (N8345, N8330, N7006, N1451, N1376);
xor XOR2 (N8346, N8326, N1579);
nand NAND4 (N8347, N8345, N5652, N8342, N825);
or OR2 (N8348, N5006, N3613);
and AND3 (N8349, N8343, N2618, N2249);
not NOT1 (N8350, N8322);
and AND3 (N8351, N8348, N4990, N832);
buf BUF1 (N8352, N8351);
or OR4 (N8353, N8335, N4766, N7968, N2116);
and AND2 (N8354, N8349, N4872);
nand NAND3 (N8355, N8346, N1781, N3651);
nand NAND3 (N8356, N8355, N4377, N8348);
or OR3 (N8357, N8341, N6535, N3052);
buf BUF1 (N8358, N8356);
buf BUF1 (N8359, N8344);
buf BUF1 (N8360, N8339);
nand NAND3 (N8361, N8353, N2652, N1383);
nor NOR4 (N8362, N8350, N6904, N5913, N5449);
and AND2 (N8363, N8361, N5517);
nand NAND3 (N8364, N8338, N5609, N218);
nand NAND2 (N8365, N8363, N2196);
xor XOR2 (N8366, N8358, N5927);
not NOT1 (N8367, N8352);
not NOT1 (N8368, N8367);
or OR4 (N8369, N8347, N6440, N5406, N8112);
xor XOR2 (N8370, N8359, N4996);
buf BUF1 (N8371, N8360);
buf BUF1 (N8372, N8371);
nor NOR3 (N8373, N8354, N6501, N4681);
buf BUF1 (N8374, N8366);
nand NAND3 (N8375, N8365, N3899, N7901);
nor NOR4 (N8376, N8362, N7163, N3117, N7279);
buf BUF1 (N8377, N8376);
xor XOR2 (N8378, N8374, N1906);
buf BUF1 (N8379, N8372);
and AND3 (N8380, N8369, N4459, N3594);
buf BUF1 (N8381, N8357);
nor NOR3 (N8382, N8379, N6362, N1063);
nand NAND2 (N8383, N8368, N7968);
and AND4 (N8384, N8381, N7583, N3590, N4508);
buf BUF1 (N8385, N8383);
xor XOR2 (N8386, N8373, N4631);
buf BUF1 (N8387, N8378);
nor NOR3 (N8388, N8364, N2570, N1416);
or OR2 (N8389, N8382, N5490);
or OR4 (N8390, N8384, N4636, N4770, N774);
and AND2 (N8391, N8386, N243);
nand NAND3 (N8392, N8377, N6341, N5432);
and AND3 (N8393, N8370, N7733, N889);
nor NOR2 (N8394, N8385, N5154);
nand NAND4 (N8395, N8392, N3670, N7028, N3449);
or OR4 (N8396, N8395, N5769, N3297, N8035);
xor XOR2 (N8397, N8391, N317);
xor XOR2 (N8398, N8387, N4796);
not NOT1 (N8399, N8398);
xor XOR2 (N8400, N8393, N1397);
or OR2 (N8401, N8380, N751);
nor NOR2 (N8402, N8400, N6855);
and AND2 (N8403, N8375, N1742);
nor NOR2 (N8404, N8401, N4371);
or OR4 (N8405, N8399, N1043, N5569, N2773);
nand NAND2 (N8406, N8405, N633);
xor XOR2 (N8407, N8389, N4358);
nor NOR4 (N8408, N8396, N3706, N1603, N1996);
buf BUF1 (N8409, N8390);
nor NOR4 (N8410, N8388, N5814, N4069, N4077);
or OR2 (N8411, N8407, N1206);
buf BUF1 (N8412, N8404);
and AND2 (N8413, N8406, N4947);
nand NAND2 (N8414, N8403, N4914);
not NOT1 (N8415, N8412);
not NOT1 (N8416, N8413);
xor XOR2 (N8417, N8414, N3277);
buf BUF1 (N8418, N8402);
nor NOR2 (N8419, N8408, N7045);
nor NOR3 (N8420, N8409, N3418, N5798);
not NOT1 (N8421, N8394);
and AND3 (N8422, N8420, N1418, N4251);
or OR3 (N8423, N8415, N3422, N2129);
nor NOR4 (N8424, N8422, N4084, N7981, N8193);
and AND3 (N8425, N8397, N7176, N5086);
not NOT1 (N8426, N8418);
not NOT1 (N8427, N8426);
nor NOR4 (N8428, N8421, N7928, N2242, N6453);
and AND4 (N8429, N8428, N5512, N2085, N5224);
and AND4 (N8430, N8427, N4495, N4367, N526);
xor XOR2 (N8431, N8419, N6000);
not NOT1 (N8432, N8411);
nor NOR3 (N8433, N8424, N2266, N6911);
not NOT1 (N8434, N8423);
nor NOR4 (N8435, N8430, N4449, N6962, N8335);
nor NOR4 (N8436, N8416, N496, N3499, N7736);
xor XOR2 (N8437, N8433, N1538);
buf BUF1 (N8438, N8436);
and AND4 (N8439, N8410, N2022, N5205, N3088);
or OR3 (N8440, N8438, N4619, N5891);
or OR3 (N8441, N8431, N4748, N3361);
or OR2 (N8442, N8437, N6123);
or OR3 (N8443, N8441, N5846, N6341);
nand NAND2 (N8444, N8443, N3862);
or OR3 (N8445, N8432, N3584, N96);
or OR4 (N8446, N8442, N7538, N1019, N6321);
not NOT1 (N8447, N8417);
nor NOR4 (N8448, N8435, N4956, N553, N3783);
nand NAND2 (N8449, N8429, N2315);
buf BUF1 (N8450, N8447);
xor XOR2 (N8451, N8444, N7265);
or OR4 (N8452, N8425, N2564, N145, N5808);
nand NAND2 (N8453, N8445, N8311);
buf BUF1 (N8454, N8451);
nand NAND3 (N8455, N8450, N5277, N1157);
nand NAND2 (N8456, N8448, N4534);
not NOT1 (N8457, N8456);
or OR2 (N8458, N8440, N1625);
and AND3 (N8459, N8452, N2632, N3417);
nand NAND2 (N8460, N8459, N3880);
and AND2 (N8461, N8460, N2204);
xor XOR2 (N8462, N8461, N3349);
or OR2 (N8463, N8449, N235);
or OR4 (N8464, N8457, N2165, N1445, N1204);
or OR3 (N8465, N8463, N1221, N5113);
nor NOR4 (N8466, N8455, N2547, N5250, N3598);
and AND4 (N8467, N8458, N4484, N8258, N7050);
xor XOR2 (N8468, N8453, N6037);
nand NAND3 (N8469, N8466, N512, N6144);
nand NAND4 (N8470, N8439, N523, N1245, N7190);
not NOT1 (N8471, N8465);
buf BUF1 (N8472, N8446);
nand NAND2 (N8473, N8471, N4946);
nor NOR4 (N8474, N8469, N6126, N4033, N4552);
and AND2 (N8475, N8470, N5594);
buf BUF1 (N8476, N8467);
and AND3 (N8477, N8473, N2312, N7078);
and AND4 (N8478, N8477, N1696, N5207, N2189);
or OR3 (N8479, N8468, N873, N7034);
nand NAND3 (N8480, N8464, N5666, N4948);
buf BUF1 (N8481, N8434);
xor XOR2 (N8482, N8476, N5758);
nand NAND4 (N8483, N8475, N5197, N6236, N8473);
or OR2 (N8484, N8478, N6343);
xor XOR2 (N8485, N8472, N1821);
buf BUF1 (N8486, N8484);
or OR4 (N8487, N8486, N2395, N4848, N5870);
buf BUF1 (N8488, N8482);
or OR2 (N8489, N8487, N2524);
or OR2 (N8490, N8485, N6342);
nand NAND2 (N8491, N8488, N341);
buf BUF1 (N8492, N8479);
xor XOR2 (N8493, N8480, N1491);
and AND3 (N8494, N8489, N186, N867);
xor XOR2 (N8495, N8483, N1210);
or OR2 (N8496, N8491, N7887);
nand NAND2 (N8497, N8496, N1479);
xor XOR2 (N8498, N8490, N6617);
and AND2 (N8499, N8497, N7293);
not NOT1 (N8500, N8481);
and AND4 (N8501, N8494, N6609, N807, N1236);
or OR2 (N8502, N8454, N2105);
nor NOR2 (N8503, N8498, N2204);
and AND2 (N8504, N8474, N4934);
xor XOR2 (N8505, N8462, N4203);
nand NAND3 (N8506, N8504, N6992, N6587);
buf BUF1 (N8507, N8503);
nand NAND2 (N8508, N8507, N2244);
or OR4 (N8509, N8505, N5464, N1747, N6071);
nand NAND2 (N8510, N8506, N670);
not NOT1 (N8511, N8502);
or OR2 (N8512, N8510, N997);
xor XOR2 (N8513, N8492, N8155);
nand NAND3 (N8514, N8511, N3745, N8385);
nor NOR2 (N8515, N8513, N3059);
or OR4 (N8516, N8512, N7601, N1871, N665);
nor NOR4 (N8517, N8493, N308, N6591, N1858);
xor XOR2 (N8518, N8517, N631);
xor XOR2 (N8519, N8516, N1767);
nor NOR4 (N8520, N8500, N1682, N434, N6169);
and AND2 (N8521, N8509, N3018);
xor XOR2 (N8522, N8501, N6718);
nor NOR3 (N8523, N8521, N5437, N5421);
nor NOR4 (N8524, N8508, N1138, N2702, N4192);
nor NOR3 (N8525, N8522, N4643, N2127);
buf BUF1 (N8526, N8514);
and AND4 (N8527, N8499, N7801, N7380, N3156);
buf BUF1 (N8528, N8520);
and AND2 (N8529, N8519, N2428);
nand NAND3 (N8530, N8523, N5260, N3758);
nand NAND3 (N8531, N8526, N1207, N1206);
buf BUF1 (N8532, N8495);
and AND2 (N8533, N8527, N1286);
nand NAND4 (N8534, N8532, N692, N4939, N7712);
and AND2 (N8535, N8528, N5559);
not NOT1 (N8536, N8535);
nand NAND3 (N8537, N8524, N7149, N6958);
not NOT1 (N8538, N8525);
and AND3 (N8539, N8534, N1686, N7759);
not NOT1 (N8540, N8533);
not NOT1 (N8541, N8536);
nor NOR2 (N8542, N8530, N2058);
or OR2 (N8543, N8518, N6780);
xor XOR2 (N8544, N8543, N6439);
and AND4 (N8545, N8540, N1423, N3628, N2185);
and AND3 (N8546, N8515, N1793, N879);
xor XOR2 (N8547, N8538, N276);
nor NOR2 (N8548, N8537, N7066);
buf BUF1 (N8549, N8542);
and AND3 (N8550, N8547, N4885, N8324);
buf BUF1 (N8551, N8548);
not NOT1 (N8552, N8545);
buf BUF1 (N8553, N8529);
buf BUF1 (N8554, N8544);
or OR3 (N8555, N8551, N8053, N7532);
buf BUF1 (N8556, N8554);
xor XOR2 (N8557, N8539, N1192);
and AND4 (N8558, N8531, N3513, N2301, N7405);
or OR4 (N8559, N8546, N6039, N5012, N4648);
and AND2 (N8560, N8555, N1662);
nor NOR3 (N8561, N8559, N8112, N6047);
xor XOR2 (N8562, N8561, N6987);
nand NAND2 (N8563, N8541, N6232);
and AND4 (N8564, N8550, N2587, N1958, N6018);
and AND4 (N8565, N8560, N3482, N6688, N7063);
buf BUF1 (N8566, N8558);
not NOT1 (N8567, N8563);
xor XOR2 (N8568, N8562, N4000);
not NOT1 (N8569, N8557);
nor NOR2 (N8570, N8567, N3461);
buf BUF1 (N8571, N8552);
nand NAND4 (N8572, N8570, N3755, N6093, N5672);
not NOT1 (N8573, N8568);
and AND3 (N8574, N8571, N3229, N4599);
or OR4 (N8575, N8569, N4533, N222, N6310);
and AND3 (N8576, N8575, N7377, N2115);
nor NOR3 (N8577, N8573, N4129, N3890);
and AND4 (N8578, N8572, N2168, N5647, N8223);
nor NOR3 (N8579, N8577, N1317, N6537);
not NOT1 (N8580, N8578);
or OR3 (N8581, N8576, N6808, N6428);
or OR4 (N8582, N8549, N4882, N1356, N6686);
or OR2 (N8583, N8581, N7770);
not NOT1 (N8584, N8566);
nor NOR2 (N8585, N8574, N5193);
nand NAND3 (N8586, N8565, N560, N5501);
or OR4 (N8587, N8584, N1120, N1483, N6627);
buf BUF1 (N8588, N8580);
nand NAND4 (N8589, N8553, N6139, N2909, N8017);
and AND2 (N8590, N8587, N729);
or OR4 (N8591, N8579, N3546, N1953, N604);
xor XOR2 (N8592, N8582, N8394);
nor NOR2 (N8593, N8586, N3659);
and AND4 (N8594, N8556, N5763, N7532, N4458);
or OR3 (N8595, N8593, N1856, N2304);
not NOT1 (N8596, N8595);
buf BUF1 (N8597, N8591);
buf BUF1 (N8598, N8590);
xor XOR2 (N8599, N8583, N3228);
not NOT1 (N8600, N8596);
or OR2 (N8601, N8599, N4751);
xor XOR2 (N8602, N8589, N6704);
nor NOR2 (N8603, N8588, N1172);
buf BUF1 (N8604, N8564);
xor XOR2 (N8605, N8597, N7162);
not NOT1 (N8606, N8604);
xor XOR2 (N8607, N8594, N7386);
nand NAND2 (N8608, N8601, N8236);
xor XOR2 (N8609, N8592, N3498);
nor NOR4 (N8610, N8600, N6853, N1135, N1082);
or OR4 (N8611, N8598, N2634, N3255, N1021);
nand NAND2 (N8612, N8602, N4885);
nand NAND4 (N8613, N8612, N712, N5814, N6895);
xor XOR2 (N8614, N8605, N1244);
not NOT1 (N8615, N8608);
nand NAND3 (N8616, N8611, N2101, N188);
nand NAND2 (N8617, N8613, N7957);
not NOT1 (N8618, N8617);
or OR2 (N8619, N8603, N1);
nor NOR2 (N8620, N8607, N3934);
buf BUF1 (N8621, N8618);
buf BUF1 (N8622, N8606);
nor NOR2 (N8623, N8620, N3218);
and AND2 (N8624, N8616, N7352);
buf BUF1 (N8625, N8621);
and AND3 (N8626, N8609, N1075, N8062);
or OR3 (N8627, N8623, N7338, N7740);
nand NAND3 (N8628, N8585, N6077, N6770);
buf BUF1 (N8629, N8626);
nor NOR4 (N8630, N8615, N8006, N2691, N7585);
not NOT1 (N8631, N8624);
and AND4 (N8632, N8628, N6766, N526, N5258);
buf BUF1 (N8633, N8614);
not NOT1 (N8634, N8633);
nand NAND2 (N8635, N8627, N3419);
xor XOR2 (N8636, N8622, N5874);
or OR3 (N8637, N8610, N489, N8302);
not NOT1 (N8638, N8630);
and AND3 (N8639, N8631, N49, N472);
and AND2 (N8640, N8638, N4299);
nor NOR4 (N8641, N8632, N190, N2442, N5219);
xor XOR2 (N8642, N8641, N1289);
not NOT1 (N8643, N8629);
and AND2 (N8644, N8640, N8401);
buf BUF1 (N8645, N8644);
nand NAND4 (N8646, N8637, N6206, N3614, N1994);
nor NOR4 (N8647, N8636, N328, N5560, N913);
or OR3 (N8648, N8625, N6956, N7956);
not NOT1 (N8649, N8634);
xor XOR2 (N8650, N8649, N1399);
nor NOR2 (N8651, N8639, N1558);
and AND4 (N8652, N8650, N8021, N7688, N6307);
and AND3 (N8653, N8647, N2042, N6279);
nand NAND4 (N8654, N8642, N5416, N2476, N3628);
nor NOR2 (N8655, N8648, N5265);
not NOT1 (N8656, N8645);
buf BUF1 (N8657, N8655);
or OR4 (N8658, N8656, N2590, N6500, N4022);
or OR4 (N8659, N8643, N6396, N5748, N8566);
xor XOR2 (N8660, N8652, N3771);
nand NAND3 (N8661, N8619, N2868, N8606);
and AND3 (N8662, N8653, N5782, N718);
not NOT1 (N8663, N8646);
xor XOR2 (N8664, N8663, N8363);
xor XOR2 (N8665, N8662, N2312);
or OR4 (N8666, N8657, N242, N2070, N649);
buf BUF1 (N8667, N8654);
buf BUF1 (N8668, N8665);
not NOT1 (N8669, N8661);
buf BUF1 (N8670, N8660);
not NOT1 (N8671, N8667);
not NOT1 (N8672, N8659);
xor XOR2 (N8673, N8671, N4964);
xor XOR2 (N8674, N8668, N6237);
and AND3 (N8675, N8674, N2566, N8412);
not NOT1 (N8676, N8664);
not NOT1 (N8677, N8635);
xor XOR2 (N8678, N8677, N3031);
or OR3 (N8679, N8678, N7605, N6092);
nor NOR3 (N8680, N8672, N8053, N3395);
xor XOR2 (N8681, N8680, N6402);
xor XOR2 (N8682, N8681, N2536);
or OR3 (N8683, N8675, N2956, N2603);
buf BUF1 (N8684, N8651);
not NOT1 (N8685, N8679);
and AND4 (N8686, N8685, N5269, N8335, N7450);
and AND4 (N8687, N8669, N7242, N5478, N941);
and AND3 (N8688, N8670, N8073, N7106);
not NOT1 (N8689, N8658);
and AND3 (N8690, N8689, N1878, N5536);
xor XOR2 (N8691, N8690, N7889);
buf BUF1 (N8692, N8684);
not NOT1 (N8693, N8683);
buf BUF1 (N8694, N8673);
xor XOR2 (N8695, N8691, N1381);
not NOT1 (N8696, N8666);
xor XOR2 (N8697, N8694, N183);
not NOT1 (N8698, N8676);
and AND4 (N8699, N8693, N3600, N4756, N7211);
or OR2 (N8700, N8696, N1906);
buf BUF1 (N8701, N8686);
xor XOR2 (N8702, N8699, N4603);
buf BUF1 (N8703, N8688);
not NOT1 (N8704, N8697);
nor NOR4 (N8705, N8682, N1069, N5430, N4417);
xor XOR2 (N8706, N8703, N5449);
nand NAND4 (N8707, N8695, N2339, N2995, N2270);
not NOT1 (N8708, N8706);
nor NOR3 (N8709, N8707, N787, N328);
and AND2 (N8710, N8704, N5238);
buf BUF1 (N8711, N8700);
not NOT1 (N8712, N8709);
buf BUF1 (N8713, N8698);
nor NOR3 (N8714, N8712, N8220, N5632);
and AND4 (N8715, N8708, N2918, N2330, N1032);
xor XOR2 (N8716, N8710, N3925);
nand NAND3 (N8717, N8715, N5424, N5605);
buf BUF1 (N8718, N8705);
nand NAND4 (N8719, N8717, N8678, N5642, N6129);
xor XOR2 (N8720, N8718, N8375);
and AND4 (N8721, N8714, N441, N2168, N3844);
xor XOR2 (N8722, N8701, N8169);
not NOT1 (N8723, N8719);
xor XOR2 (N8724, N8721, N5855);
xor XOR2 (N8725, N8724, N6758);
nor NOR2 (N8726, N8713, N8355);
nand NAND3 (N8727, N8725, N645, N3950);
not NOT1 (N8728, N8726);
or OR4 (N8729, N8702, N8235, N8518, N4509);
nand NAND3 (N8730, N8692, N4166, N1686);
and AND4 (N8731, N8716, N3468, N7039, N5892);
and AND4 (N8732, N8720, N8057, N2030, N1327);
or OR4 (N8733, N8727, N8205, N6488, N1216);
xor XOR2 (N8734, N8687, N2962);
buf BUF1 (N8735, N8729);
buf BUF1 (N8736, N8735);
or OR3 (N8737, N8730, N2756, N265);
or OR3 (N8738, N8732, N8442, N5418);
not NOT1 (N8739, N8723);
nand NAND3 (N8740, N8722, N3507, N11);
and AND3 (N8741, N8738, N4168, N5424);
or OR3 (N8742, N8740, N7353, N4828);
not NOT1 (N8743, N8737);
not NOT1 (N8744, N8734);
nor NOR4 (N8745, N8728, N5361, N597, N7478);
and AND2 (N8746, N8743, N5643);
or OR2 (N8747, N8736, N1556);
nor NOR3 (N8748, N8747, N3801, N5592);
buf BUF1 (N8749, N8731);
nor NOR3 (N8750, N8741, N5957, N1530);
nor NOR3 (N8751, N8711, N3670, N3858);
or OR3 (N8752, N8733, N379, N775);
buf BUF1 (N8753, N8752);
or OR4 (N8754, N8744, N1528, N7218, N752);
nor NOR3 (N8755, N8754, N3396, N1464);
or OR3 (N8756, N8746, N7729, N1383);
xor XOR2 (N8757, N8748, N219);
buf BUF1 (N8758, N8755);
xor XOR2 (N8759, N8751, N2179);
buf BUF1 (N8760, N8756);
xor XOR2 (N8761, N8745, N4429);
nor NOR3 (N8762, N8750, N1243, N841);
nand NAND3 (N8763, N8739, N2257, N7477);
xor XOR2 (N8764, N8760, N2891);
or OR4 (N8765, N8749, N3426, N2860, N4037);
nor NOR4 (N8766, N8759, N3423, N4387, N263);
not NOT1 (N8767, N8758);
nor NOR4 (N8768, N8763, N7813, N6124, N956);
and AND2 (N8769, N8764, N2077);
or OR2 (N8770, N8765, N6429);
not NOT1 (N8771, N8768);
not NOT1 (N8772, N8753);
nor NOR2 (N8773, N8769, N4009);
and AND4 (N8774, N8771, N1603, N3416, N2723);
nor NOR4 (N8775, N8757, N7115, N5359, N1652);
buf BUF1 (N8776, N8774);
or OR3 (N8777, N8776, N914, N3434);
xor XOR2 (N8778, N8777, N8621);
nor NOR4 (N8779, N8766, N5635, N4610, N1770);
nor NOR3 (N8780, N8762, N7008, N7822);
buf BUF1 (N8781, N8775);
xor XOR2 (N8782, N8742, N1126);
not NOT1 (N8783, N8778);
xor XOR2 (N8784, N8782, N8207);
nand NAND3 (N8785, N8784, N2583, N431);
xor XOR2 (N8786, N8783, N2013);
or OR4 (N8787, N8761, N3856, N8263, N5715);
and AND2 (N8788, N8770, N5568);
xor XOR2 (N8789, N8787, N4458);
buf BUF1 (N8790, N8772);
buf BUF1 (N8791, N8780);
nand NAND3 (N8792, N8781, N286, N7432);
nor NOR3 (N8793, N8786, N296, N2456);
xor XOR2 (N8794, N8789, N7325);
nand NAND3 (N8795, N8792, N6393, N1898);
nor NOR4 (N8796, N8795, N1301, N799, N5195);
xor XOR2 (N8797, N8785, N3752);
buf BUF1 (N8798, N8788);
nor NOR4 (N8799, N8793, N75, N2081, N7537);
and AND2 (N8800, N8773, N2902);
nand NAND4 (N8801, N8797, N2321, N184, N4073);
nand NAND2 (N8802, N8794, N2896);
nand NAND2 (N8803, N8796, N3619);
buf BUF1 (N8804, N8799);
nor NOR3 (N8805, N8801, N500, N5552);
xor XOR2 (N8806, N8804, N4548);
nor NOR3 (N8807, N8802, N4498, N1694);
buf BUF1 (N8808, N8807);
nand NAND3 (N8809, N8791, N2439, N3747);
buf BUF1 (N8810, N8767);
and AND4 (N8811, N8779, N3160, N6885, N2157);
or OR3 (N8812, N8810, N946, N7322);
nor NOR2 (N8813, N8808, N2591);
and AND2 (N8814, N8813, N5731);
or OR2 (N8815, N8811, N1491);
not NOT1 (N8816, N8803);
or OR3 (N8817, N8815, N2827, N7796);
or OR2 (N8818, N8817, N452);
nor NOR3 (N8819, N8805, N3835, N7272);
not NOT1 (N8820, N8798);
xor XOR2 (N8821, N8819, N6836);
not NOT1 (N8822, N8812);
nor NOR2 (N8823, N8790, N4757);
nand NAND4 (N8824, N8822, N8071, N7879, N6009);
nand NAND3 (N8825, N8820, N2930, N6972);
nor NOR2 (N8826, N8824, N7946);
not NOT1 (N8827, N8818);
xor XOR2 (N8828, N8825, N3178);
or OR4 (N8829, N8821, N908, N4819, N1824);
nand NAND4 (N8830, N8809, N5452, N4140, N8491);
nor NOR2 (N8831, N8806, N1871);
buf BUF1 (N8832, N8800);
or OR4 (N8833, N8828, N8248, N7392, N8180);
and AND4 (N8834, N8833, N4936, N4884, N1821);
xor XOR2 (N8835, N8814, N2530);
nor NOR3 (N8836, N8829, N8397, N4628);
and AND2 (N8837, N8816, N5158);
not NOT1 (N8838, N8826);
nand NAND3 (N8839, N8836, N1361, N318);
and AND4 (N8840, N8830, N1218, N7147, N3122);
buf BUF1 (N8841, N8832);
xor XOR2 (N8842, N8841, N5930);
or OR4 (N8843, N8834, N1897, N1764, N7331);
nand NAND4 (N8844, N8843, N57, N1222, N293);
not NOT1 (N8845, N8842);
or OR2 (N8846, N8827, N1916);
and AND3 (N8847, N8835, N3772, N1126);
buf BUF1 (N8848, N8823);
and AND3 (N8849, N8846, N3504, N8103);
buf BUF1 (N8850, N8838);
xor XOR2 (N8851, N8839, N3225);
and AND4 (N8852, N8848, N1318, N3201, N4607);
nand NAND4 (N8853, N8844, N6253, N6819, N2793);
nor NOR2 (N8854, N8850, N1657);
buf BUF1 (N8855, N8845);
not NOT1 (N8856, N8831);
xor XOR2 (N8857, N8855, N2423);
and AND4 (N8858, N8856, N8065, N6668, N644);
nand NAND4 (N8859, N8854, N2229, N2846, N6080);
or OR3 (N8860, N8837, N3976, N289);
nand NAND4 (N8861, N8840, N3112, N6117, N3962);
and AND4 (N8862, N8861, N8519, N8396, N786);
xor XOR2 (N8863, N8849, N1637);
and AND4 (N8864, N8863, N7561, N5549, N8157);
nor NOR3 (N8865, N8858, N3374, N3385);
buf BUF1 (N8866, N8851);
not NOT1 (N8867, N8865);
and AND3 (N8868, N8867, N5760, N7300);
xor XOR2 (N8869, N8864, N1637);
nand NAND3 (N8870, N8847, N7084, N1692);
not NOT1 (N8871, N8870);
or OR3 (N8872, N8853, N1080, N3759);
buf BUF1 (N8873, N8869);
not NOT1 (N8874, N8860);
or OR4 (N8875, N8873, N5301, N2125, N6068);
or OR2 (N8876, N8859, N4557);
nor NOR3 (N8877, N8866, N7166, N5158);
and AND4 (N8878, N8862, N3476, N256, N1641);
or OR3 (N8879, N8852, N1477, N1602);
buf BUF1 (N8880, N8874);
xor XOR2 (N8881, N8857, N1386);
buf BUF1 (N8882, N8868);
and AND2 (N8883, N8877, N3990);
or OR3 (N8884, N8878, N491, N1124);
xor XOR2 (N8885, N8875, N6401);
not NOT1 (N8886, N8883);
nor NOR2 (N8887, N8872, N4102);
xor XOR2 (N8888, N8880, N6750);
nor NOR3 (N8889, N8879, N3546, N3580);
buf BUF1 (N8890, N8886);
or OR2 (N8891, N8887, N7536);
nor NOR4 (N8892, N8884, N3045, N2528, N7291);
and AND2 (N8893, N8881, N2743);
and AND3 (N8894, N8893, N135, N4873);
nor NOR2 (N8895, N8876, N5691);
buf BUF1 (N8896, N8894);
xor XOR2 (N8897, N8891, N896);
buf BUF1 (N8898, N8897);
xor XOR2 (N8899, N8896, N3569);
or OR4 (N8900, N8882, N579, N2898, N5172);
and AND2 (N8901, N8889, N3233);
nand NAND2 (N8902, N8899, N7502);
xor XOR2 (N8903, N8901, N4284);
nor NOR3 (N8904, N8900, N5897, N4117);
or OR3 (N8905, N8898, N3890, N3309);
and AND3 (N8906, N8892, N5298, N3818);
and AND2 (N8907, N8903, N1954);
nor NOR2 (N8908, N8906, N132);
nor NOR3 (N8909, N8888, N544, N1804);
and AND4 (N8910, N8885, N4647, N3770, N1002);
and AND4 (N8911, N8907, N4772, N5719, N3433);
nand NAND4 (N8912, N8871, N5115, N1729, N4121);
xor XOR2 (N8913, N8912, N2);
nor NOR3 (N8914, N8908, N4601, N1046);
nand NAND2 (N8915, N8890, N4431);
not NOT1 (N8916, N8915);
xor XOR2 (N8917, N8895, N2794);
nand NAND4 (N8918, N8914, N6582, N6824, N6822);
nor NOR3 (N8919, N8911, N2924, N1831);
xor XOR2 (N8920, N8917, N1614);
not NOT1 (N8921, N8918);
nand NAND2 (N8922, N8904, N1449);
and AND4 (N8923, N8902, N1311, N972, N5801);
not NOT1 (N8924, N8920);
nand NAND3 (N8925, N8916, N3109, N654);
nand NAND3 (N8926, N8905, N954, N954);
and AND3 (N8927, N8921, N1943, N469);
and AND4 (N8928, N8923, N412, N7, N5093);
nor NOR2 (N8929, N8924, N1955);
xor XOR2 (N8930, N8925, N4621);
xor XOR2 (N8931, N8926, N7434);
nor NOR3 (N8932, N8913, N4472, N7363);
and AND3 (N8933, N8932, N5998, N5064);
or OR2 (N8934, N8922, N1358);
nor NOR4 (N8935, N8919, N1171, N1926, N4659);
or OR3 (N8936, N8931, N6172, N1400);
and AND2 (N8937, N8936, N430);
xor XOR2 (N8938, N8927, N5640);
nor NOR3 (N8939, N8929, N1864, N115);
or OR4 (N8940, N8930, N79, N1999, N3953);
nand NAND3 (N8941, N8939, N209, N771);
nor NOR3 (N8942, N8934, N4231, N2498);
nor NOR3 (N8943, N8910, N345, N2442);
nand NAND3 (N8944, N8933, N801, N4280);
nor NOR2 (N8945, N8944, N458);
not NOT1 (N8946, N8938);
xor XOR2 (N8947, N8937, N5382);
buf BUF1 (N8948, N8935);
nand NAND2 (N8949, N8941, N3249);
xor XOR2 (N8950, N8943, N7362);
or OR2 (N8951, N8945, N3541);
nand NAND4 (N8952, N8951, N1972, N8205, N7533);
not NOT1 (N8953, N8947);
and AND4 (N8954, N8948, N3010, N2801, N6990);
or OR3 (N8955, N8949, N5390, N2952);
nand NAND2 (N8956, N8952, N61);
and AND3 (N8957, N8950, N6582, N1590);
xor XOR2 (N8958, N8942, N1429);
buf BUF1 (N8959, N8940);
buf BUF1 (N8960, N8959);
nor NOR3 (N8961, N8928, N637, N4690);
nor NOR4 (N8962, N8953, N8700, N1539, N5484);
xor XOR2 (N8963, N8956, N3841);
nand NAND2 (N8964, N8962, N4804);
nor NOR2 (N8965, N8960, N5764);
nand NAND4 (N8966, N8946, N6927, N8428, N2539);
not NOT1 (N8967, N8955);
or OR4 (N8968, N8963, N2249, N8121, N1213);
nand NAND2 (N8969, N8961, N1014);
nor NOR4 (N8970, N8964, N3284, N6430, N5159);
buf BUF1 (N8971, N8968);
nor NOR2 (N8972, N8954, N4984);
and AND3 (N8973, N8966, N3243, N4029);
nor NOR4 (N8974, N8970, N2325, N2694, N4693);
not NOT1 (N8975, N8957);
nor NOR2 (N8976, N8965, N8111);
not NOT1 (N8977, N8969);
not NOT1 (N8978, N8974);
or OR4 (N8979, N8958, N6355, N5690, N892);
nor NOR2 (N8980, N8979, N930);
nor NOR4 (N8981, N8967, N6064, N6060, N6740);
nor NOR4 (N8982, N8980, N6560, N3422, N4970);
nor NOR2 (N8983, N8977, N870);
or OR3 (N8984, N8981, N2665, N8275);
nand NAND3 (N8985, N8983, N6397, N4090);
nor NOR2 (N8986, N8985, N8376);
nand NAND3 (N8987, N8986, N3775, N1995);
and AND3 (N8988, N8971, N5737, N4076);
or OR2 (N8989, N8973, N2967);
buf BUF1 (N8990, N8988);
not NOT1 (N8991, N8984);
or OR4 (N8992, N8972, N2597, N3363, N3832);
buf BUF1 (N8993, N8978);
and AND4 (N8994, N8975, N284, N1617, N678);
buf BUF1 (N8995, N8987);
or OR2 (N8996, N8982, N8764);
or OR3 (N8997, N8909, N3325, N6653);
and AND3 (N8998, N8976, N3478, N5809);
and AND4 (N8999, N8991, N8856, N1571, N1551);
nand NAND2 (N9000, N8996, N8808);
and AND4 (N9001, N9000, N4202, N7654, N2657);
and AND4 (N9002, N8995, N3879, N554, N122);
buf BUF1 (N9003, N8993);
or OR4 (N9004, N8999, N5045, N3590, N7110);
or OR2 (N9005, N8998, N6901);
xor XOR2 (N9006, N8992, N8571);
and AND2 (N9007, N8994, N7131);
not NOT1 (N9008, N9001);
buf BUF1 (N9009, N8989);
not NOT1 (N9010, N9002);
nand NAND4 (N9011, N8997, N2646, N6874, N6652);
or OR4 (N9012, N9009, N2016, N3166, N4629);
or OR2 (N9013, N9003, N4950);
not NOT1 (N9014, N8990);
buf BUF1 (N9015, N9014);
or OR2 (N9016, N9006, N1327);
or OR2 (N9017, N9016, N694);
xor XOR2 (N9018, N9008, N7126);
and AND2 (N9019, N9013, N7603);
xor XOR2 (N9020, N9004, N1224);
and AND3 (N9021, N9010, N2884, N6764);
nand NAND4 (N9022, N9020, N3062, N1595, N5839);
buf BUF1 (N9023, N9022);
buf BUF1 (N9024, N9017);
not NOT1 (N9025, N9021);
not NOT1 (N9026, N9007);
and AND4 (N9027, N9015, N7840, N8179, N1772);
and AND2 (N9028, N9023, N8740);
nand NAND4 (N9029, N9019, N7388, N6895, N6502);
nand NAND2 (N9030, N9024, N2576);
xor XOR2 (N9031, N9029, N2208);
nor NOR4 (N9032, N9018, N5851, N6318, N104);
nand NAND2 (N9033, N9031, N5940);
nand NAND2 (N9034, N9026, N8288);
not NOT1 (N9035, N9012);
buf BUF1 (N9036, N9005);
or OR3 (N9037, N9036, N2595, N2165);
nand NAND4 (N9038, N9028, N5825, N6290, N3626);
nand NAND4 (N9039, N9033, N4040, N2089, N3822);
xor XOR2 (N9040, N9011, N534);
and AND2 (N9041, N9027, N1202);
xor XOR2 (N9042, N9035, N1585);
xor XOR2 (N9043, N9041, N1555);
and AND2 (N9044, N9034, N3697);
buf BUF1 (N9045, N9043);
and AND4 (N9046, N9038, N7797, N1415, N4366);
or OR2 (N9047, N9025, N3132);
and AND2 (N9048, N9044, N8096);
buf BUF1 (N9049, N9048);
xor XOR2 (N9050, N9032, N7071);
and AND2 (N9051, N9040, N6195);
and AND4 (N9052, N9045, N4892, N5293, N6886);
or OR2 (N9053, N9051, N2905);
not NOT1 (N9054, N9039);
nor NOR3 (N9055, N9030, N4399, N8392);
xor XOR2 (N9056, N9055, N6566);
not NOT1 (N9057, N9053);
not NOT1 (N9058, N9056);
buf BUF1 (N9059, N9049);
xor XOR2 (N9060, N9042, N709);
xor XOR2 (N9061, N9058, N677);
buf BUF1 (N9062, N9037);
nor NOR4 (N9063, N9061, N4918, N8269, N1735);
nor NOR4 (N9064, N9047, N7208, N8908, N7056);
not NOT1 (N9065, N9057);
xor XOR2 (N9066, N9064, N1587);
xor XOR2 (N9067, N9060, N2672);
xor XOR2 (N9068, N9052, N5363);
nand NAND3 (N9069, N9067, N7171, N3759);
nor NOR4 (N9070, N9050, N3152, N2364, N3510);
xor XOR2 (N9071, N9059, N5142);
not NOT1 (N9072, N9065);
buf BUF1 (N9073, N9063);
and AND4 (N9074, N9068, N3302, N6042, N1783);
xor XOR2 (N9075, N9062, N2619);
and AND2 (N9076, N9066, N7564);
xor XOR2 (N9077, N9070, N8631);
xor XOR2 (N9078, N9075, N5748);
xor XOR2 (N9079, N9072, N3798);
or OR2 (N9080, N9054, N7205);
not NOT1 (N9081, N9078);
nand NAND2 (N9082, N9079, N5016);
buf BUF1 (N9083, N9080);
and AND2 (N9084, N9069, N2105);
not NOT1 (N9085, N9073);
and AND2 (N9086, N9084, N1079);
and AND3 (N9087, N9081, N7944, N2694);
not NOT1 (N9088, N9087);
or OR4 (N9089, N9046, N364, N1319, N6432);
not NOT1 (N9090, N9074);
buf BUF1 (N9091, N9076);
nand NAND4 (N9092, N9082, N7353, N7542, N8519);
xor XOR2 (N9093, N9085, N597);
not NOT1 (N9094, N9088);
not NOT1 (N9095, N9071);
or OR4 (N9096, N9091, N4104, N5263, N1547);
and AND3 (N9097, N9086, N5181, N2158);
xor XOR2 (N9098, N9093, N2937);
and AND2 (N9099, N9096, N3981);
and AND4 (N9100, N9083, N4228, N1294, N7973);
buf BUF1 (N9101, N9094);
not NOT1 (N9102, N9098);
buf BUF1 (N9103, N9097);
buf BUF1 (N9104, N9089);
not NOT1 (N9105, N9102);
or OR3 (N9106, N9077, N3884, N5207);
nor NOR2 (N9107, N9105, N929);
buf BUF1 (N9108, N9107);
and AND3 (N9109, N9099, N8845, N1102);
nor NOR2 (N9110, N9092, N4597);
nor NOR2 (N9111, N9100, N5992);
buf BUF1 (N9112, N9109);
and AND3 (N9113, N9103, N8186, N1301);
or OR2 (N9114, N9111, N3620);
and AND2 (N9115, N9108, N6264);
nand NAND4 (N9116, N9110, N5288, N2990, N1998);
nand NAND3 (N9117, N9101, N77, N6183);
and AND2 (N9118, N9104, N3570);
buf BUF1 (N9119, N9115);
not NOT1 (N9120, N9095);
nand NAND3 (N9121, N9116, N485, N7080);
not NOT1 (N9122, N9106);
nor NOR2 (N9123, N9119, N327);
and AND3 (N9124, N9114, N3554, N173);
not NOT1 (N9125, N9123);
and AND3 (N9126, N9125, N1839, N7674);
xor XOR2 (N9127, N9126, N832);
or OR4 (N9128, N9117, N6444, N2210, N1216);
and AND2 (N9129, N9113, N5287);
or OR3 (N9130, N9121, N7323, N1116);
nor NOR2 (N9131, N9122, N1398);
nor NOR4 (N9132, N9130, N72, N2559, N2240);
nor NOR4 (N9133, N9118, N6396, N3922, N6189);
nor NOR2 (N9134, N9124, N3673);
not NOT1 (N9135, N9134);
or OR3 (N9136, N9127, N8068, N8920);
nand NAND4 (N9137, N9112, N8759, N4630, N2800);
nand NAND4 (N9138, N9131, N6694, N279, N6726);
xor XOR2 (N9139, N9137, N5417);
xor XOR2 (N9140, N9139, N7095);
xor XOR2 (N9141, N9090, N1619);
or OR4 (N9142, N9140, N772, N398, N5740);
not NOT1 (N9143, N9135);
not NOT1 (N9144, N9128);
xor XOR2 (N9145, N9142, N2322);
xor XOR2 (N9146, N9129, N5477);
xor XOR2 (N9147, N9143, N4116);
nand NAND4 (N9148, N9120, N9019, N3196, N5261);
not NOT1 (N9149, N9145);
nand NAND2 (N9150, N9148, N1192);
buf BUF1 (N9151, N9147);
not NOT1 (N9152, N9138);
nor NOR3 (N9153, N9152, N6532, N8038);
buf BUF1 (N9154, N9153);
buf BUF1 (N9155, N9144);
or OR4 (N9156, N9136, N6141, N1458, N5960);
and AND2 (N9157, N9150, N4666);
or OR4 (N9158, N9141, N1069, N6509, N6638);
and AND2 (N9159, N9132, N5905);
and AND3 (N9160, N9133, N2125, N3753);
or OR3 (N9161, N9155, N6732, N6039);
nor NOR3 (N9162, N9161, N46, N4861);
buf BUF1 (N9163, N9160);
nor NOR2 (N9164, N9149, N112);
xor XOR2 (N9165, N9164, N4505);
and AND2 (N9166, N9154, N485);
or OR2 (N9167, N9157, N4401);
nand NAND3 (N9168, N9151, N3764, N1943);
nor NOR2 (N9169, N9168, N3581);
and AND2 (N9170, N9167, N4160);
not NOT1 (N9171, N9163);
nor NOR4 (N9172, N9165, N216, N133, N2721);
nand NAND2 (N9173, N9171, N7408);
or OR2 (N9174, N9159, N2515);
and AND2 (N9175, N9146, N8798);
nor NOR2 (N9176, N9170, N8086);
nand NAND3 (N9177, N9156, N2753, N5531);
not NOT1 (N9178, N9166);
xor XOR2 (N9179, N9173, N1231);
not NOT1 (N9180, N9175);
xor XOR2 (N9181, N9169, N3032);
nand NAND4 (N9182, N9180, N7397, N6931, N1212);
nor NOR2 (N9183, N9179, N5587);
and AND4 (N9184, N9183, N3828, N7274, N4495);
nand NAND3 (N9185, N9174, N978, N8746);
nand NAND4 (N9186, N9176, N3438, N3423, N3467);
not NOT1 (N9187, N9178);
or OR2 (N9188, N9184, N9140);
xor XOR2 (N9189, N9162, N792);
or OR4 (N9190, N9187, N1132, N4659, N5369);
not NOT1 (N9191, N9158);
buf BUF1 (N9192, N9186);
buf BUF1 (N9193, N9185);
and AND4 (N9194, N9192, N4876, N6547, N5193);
or OR4 (N9195, N9181, N8314, N6353, N1835);
and AND4 (N9196, N9190, N6808, N5486, N5622);
or OR3 (N9197, N9193, N2984, N91);
not NOT1 (N9198, N9194);
nand NAND3 (N9199, N9182, N8664, N765);
nand NAND3 (N9200, N9191, N5432, N3443);
nand NAND4 (N9201, N9172, N1471, N5841, N759);
and AND2 (N9202, N9199, N2522);
or OR2 (N9203, N9202, N4132);
buf BUF1 (N9204, N9203);
nor NOR3 (N9205, N9200, N3367, N2246);
not NOT1 (N9206, N9188);
nor NOR3 (N9207, N9177, N5644, N9198);
not NOT1 (N9208, N6194);
xor XOR2 (N9209, N9204, N1420);
or OR2 (N9210, N9207, N2565);
buf BUF1 (N9211, N9189);
nor NOR2 (N9212, N9209, N6274);
or OR3 (N9213, N9195, N1435, N5944);
and AND4 (N9214, N9213, N1386, N8928, N2719);
not NOT1 (N9215, N9196);
nor NOR3 (N9216, N9206, N3137, N1562);
xor XOR2 (N9217, N9197, N2923);
nand NAND3 (N9218, N9201, N7557, N6834);
xor XOR2 (N9219, N9217, N5097);
or OR2 (N9220, N9219, N6200);
buf BUF1 (N9221, N9216);
not NOT1 (N9222, N9212);
or OR3 (N9223, N9210, N5399, N6922);
or OR2 (N9224, N9211, N2806);
buf BUF1 (N9225, N9220);
and AND4 (N9226, N9223, N5401, N343, N9);
nand NAND3 (N9227, N9222, N1281, N8645);
and AND3 (N9228, N9218, N4689, N7899);
xor XOR2 (N9229, N9221, N8129);
xor XOR2 (N9230, N9214, N176);
buf BUF1 (N9231, N9224);
not NOT1 (N9232, N9227);
and AND2 (N9233, N9205, N4152);
nor NOR3 (N9234, N9230, N8693, N4517);
nor NOR4 (N9235, N9215, N1091, N3526, N2469);
not NOT1 (N9236, N9232);
nor NOR4 (N9237, N9208, N3010, N8801, N1860);
and AND2 (N9238, N9229, N5617);
not NOT1 (N9239, N9235);
nand NAND3 (N9240, N9233, N616, N8569);
not NOT1 (N9241, N9237);
buf BUF1 (N9242, N9239);
xor XOR2 (N9243, N9236, N550);
buf BUF1 (N9244, N9243);
not NOT1 (N9245, N9228);
nor NOR4 (N9246, N9241, N395, N5648, N3663);
not NOT1 (N9247, N9225);
or OR4 (N9248, N9231, N7376, N645, N9092);
and AND4 (N9249, N9244, N553, N7066, N3198);
and AND2 (N9250, N9248, N3517);
nor NOR3 (N9251, N9240, N3086, N6747);
or OR3 (N9252, N9250, N6753, N8385);
nor NOR4 (N9253, N9226, N3005, N212, N4809);
nand NAND2 (N9254, N9242, N978);
nor NOR4 (N9255, N9234, N3620, N4783, N261);
and AND4 (N9256, N9253, N5537, N3055, N5576);
xor XOR2 (N9257, N9247, N7211);
nand NAND4 (N9258, N9245, N8883, N361, N5205);
buf BUF1 (N9259, N9256);
xor XOR2 (N9260, N9246, N1195);
and AND2 (N9261, N9258, N1409);
nand NAND2 (N9262, N9249, N904);
and AND2 (N9263, N9262, N6571);
or OR2 (N9264, N9251, N8321);
or OR4 (N9265, N9257, N5589, N3197, N2928);
buf BUF1 (N9266, N9238);
and AND4 (N9267, N9259, N2043, N6700, N2551);
and AND4 (N9268, N9252, N5545, N4167, N1780);
xor XOR2 (N9269, N9255, N4418);
buf BUF1 (N9270, N9261);
and AND3 (N9271, N9264, N1812, N5306);
nand NAND3 (N9272, N9265, N2377, N8573);
xor XOR2 (N9273, N9268, N2431);
or OR2 (N9274, N9271, N1793);
not NOT1 (N9275, N9263);
or OR3 (N9276, N9274, N433, N5774);
not NOT1 (N9277, N9272);
xor XOR2 (N9278, N9267, N7218);
nand NAND3 (N9279, N9276, N8294, N2393);
or OR3 (N9280, N9277, N3123, N782);
not NOT1 (N9281, N9278);
buf BUF1 (N9282, N9281);
nand NAND3 (N9283, N9266, N3705, N8253);
not NOT1 (N9284, N9275);
or OR2 (N9285, N9273, N5564);
buf BUF1 (N9286, N9280);
or OR2 (N9287, N9279, N354);
buf BUF1 (N9288, N9285);
buf BUF1 (N9289, N9269);
nand NAND3 (N9290, N9284, N2715, N951);
xor XOR2 (N9291, N9270, N7554);
nor NOR2 (N9292, N9291, N5004);
xor XOR2 (N9293, N9288, N7552);
xor XOR2 (N9294, N9292, N2096);
nand NAND4 (N9295, N9294, N161, N6291, N7321);
nand NAND3 (N9296, N9283, N1324, N4747);
buf BUF1 (N9297, N9282);
buf BUF1 (N9298, N9286);
and AND4 (N9299, N9295, N6434, N8600, N1293);
or OR3 (N9300, N9254, N8152, N3498);
nor NOR3 (N9301, N9290, N8251, N4243);
or OR2 (N9302, N9296, N4726);
and AND4 (N9303, N9298, N5999, N4677, N2687);
not NOT1 (N9304, N9301);
and AND3 (N9305, N9287, N121, N8707);
nor NOR2 (N9306, N9293, N4149);
nor NOR2 (N9307, N9260, N4897);
nor NOR2 (N9308, N9304, N3476);
nor NOR2 (N9309, N9303, N2990);
nand NAND2 (N9310, N9299, N9122);
nor NOR4 (N9311, N9297, N176, N5373, N7686);
or OR4 (N9312, N9305, N1973, N7682, N3727);
nand NAND2 (N9313, N9312, N3188);
and AND3 (N9314, N9307, N408, N4486);
not NOT1 (N9315, N9310);
or OR4 (N9316, N9309, N2348, N4450, N677);
or OR3 (N9317, N9313, N4376, N2077);
buf BUF1 (N9318, N9317);
xor XOR2 (N9319, N9318, N3342);
xor XOR2 (N9320, N9289, N7977);
nor NOR4 (N9321, N9311, N2510, N2973, N4829);
or OR3 (N9322, N9308, N7145, N8801);
nor NOR4 (N9323, N9316, N4771, N5304, N2812);
xor XOR2 (N9324, N9322, N4616);
buf BUF1 (N9325, N9314);
nand NAND3 (N9326, N9300, N5676, N5525);
or OR4 (N9327, N9323, N1888, N1032, N805);
or OR3 (N9328, N9321, N5013, N965);
buf BUF1 (N9329, N9325);
or OR2 (N9330, N9319, N9146);
not NOT1 (N9331, N9315);
xor XOR2 (N9332, N9331, N1102);
or OR2 (N9333, N9306, N9228);
and AND2 (N9334, N9332, N8198);
xor XOR2 (N9335, N9302, N4004);
not NOT1 (N9336, N9333);
nand NAND3 (N9337, N9324, N4866, N5179);
and AND3 (N9338, N9336, N8557, N751);
nor NOR2 (N9339, N9337, N2988);
not NOT1 (N9340, N9326);
or OR3 (N9341, N9328, N7493, N5658);
or OR3 (N9342, N9339, N2302, N7257);
nand NAND4 (N9343, N9327, N8357, N30, N2293);
or OR4 (N9344, N9338, N5380, N803, N3336);
xor XOR2 (N9345, N9343, N4546);
nor NOR4 (N9346, N9342, N2715, N5973, N8448);
buf BUF1 (N9347, N9335);
xor XOR2 (N9348, N9334, N2921);
nor NOR4 (N9349, N9341, N8308, N7924, N4887);
nor NOR4 (N9350, N9329, N7564, N8307, N1693);
nor NOR4 (N9351, N9350, N5892, N6795, N7694);
or OR3 (N9352, N9330, N2195, N5618);
buf BUF1 (N9353, N9347);
xor XOR2 (N9354, N9351, N3120);
buf BUF1 (N9355, N9354);
and AND3 (N9356, N9352, N4677, N555);
not NOT1 (N9357, N9356);
nand NAND4 (N9358, N9348, N2119, N4945, N1751);
buf BUF1 (N9359, N9353);
not NOT1 (N9360, N9344);
nand NAND3 (N9361, N9358, N610, N8852);
buf BUF1 (N9362, N9340);
nand NAND4 (N9363, N9320, N91, N2527, N6012);
or OR4 (N9364, N9359, N3764, N8630, N1330);
not NOT1 (N9365, N9345);
and AND3 (N9366, N9363, N7016, N2596);
xor XOR2 (N9367, N9366, N64);
nor NOR2 (N9368, N9346, N8867);
buf BUF1 (N9369, N9367);
not NOT1 (N9370, N9349);
buf BUF1 (N9371, N9362);
not NOT1 (N9372, N9355);
nand NAND4 (N9373, N9364, N6909, N8434, N5698);
xor XOR2 (N9374, N9371, N6878);
or OR4 (N9375, N9372, N5950, N8381, N4292);
xor XOR2 (N9376, N9374, N7783);
nor NOR4 (N9377, N9361, N5333, N385, N8687);
and AND4 (N9378, N9370, N3865, N6813, N7920);
nand NAND4 (N9379, N9373, N2197, N8780, N3654);
xor XOR2 (N9380, N9379, N7592);
xor XOR2 (N9381, N9360, N4612);
buf BUF1 (N9382, N9376);
and AND3 (N9383, N9365, N1722, N7903);
buf BUF1 (N9384, N9368);
not NOT1 (N9385, N9375);
nand NAND2 (N9386, N9380, N8025);
buf BUF1 (N9387, N9385);
nand NAND3 (N9388, N9378, N1022, N2904);
or OR2 (N9389, N9357, N8270);
nor NOR3 (N9390, N9383, N641, N6733);
nand NAND4 (N9391, N9386, N672, N9135, N5417);
xor XOR2 (N9392, N9382, N9084);
xor XOR2 (N9393, N9384, N1532);
or OR4 (N9394, N9388, N5567, N312, N4831);
or OR3 (N9395, N9389, N9135, N6151);
buf BUF1 (N9396, N9395);
nand NAND2 (N9397, N9393, N145);
or OR2 (N9398, N9397, N5821);
xor XOR2 (N9399, N9381, N6189);
or OR2 (N9400, N9399, N2040);
and AND4 (N9401, N9369, N8900, N3468, N5179);
xor XOR2 (N9402, N9394, N2271);
xor XOR2 (N9403, N9398, N3802);
buf BUF1 (N9404, N9377);
nand NAND4 (N9405, N9387, N6926, N4139, N6299);
and AND4 (N9406, N9396, N2920, N3725, N4152);
nor NOR2 (N9407, N9402, N8243);
or OR2 (N9408, N9403, N7765);
or OR3 (N9409, N9391, N587, N9203);
nor NOR3 (N9410, N9404, N1676, N5331);
or OR4 (N9411, N9407, N5386, N7213, N4581);
nand NAND4 (N9412, N9405, N7201, N9404, N3562);
xor XOR2 (N9413, N9400, N1835);
and AND2 (N9414, N9401, N4347);
or OR2 (N9415, N9408, N3978);
nand NAND4 (N9416, N9409, N5252, N458, N1848);
and AND4 (N9417, N9414, N5740, N5590, N152);
buf BUF1 (N9418, N9406);
not NOT1 (N9419, N9410);
or OR3 (N9420, N9418, N2304, N114);
xor XOR2 (N9421, N9420, N2655);
not NOT1 (N9422, N9419);
buf BUF1 (N9423, N9422);
and AND2 (N9424, N9416, N1373);
or OR4 (N9425, N9415, N9019, N5022, N5975);
buf BUF1 (N9426, N9390);
buf BUF1 (N9427, N9412);
nand NAND4 (N9428, N9413, N6490, N1768, N3405);
buf BUF1 (N9429, N9392);
not NOT1 (N9430, N9421);
buf BUF1 (N9431, N9423);
nor NOR2 (N9432, N9427, N5396);
or OR2 (N9433, N9426, N1761);
nor NOR2 (N9434, N9429, N8594);
nor NOR4 (N9435, N9432, N6088, N6794, N9061);
buf BUF1 (N9436, N9435);
nand NAND2 (N9437, N9411, N6983);
not NOT1 (N9438, N9436);
or OR2 (N9439, N9438, N8057);
and AND2 (N9440, N9428, N2476);
not NOT1 (N9441, N9440);
nor NOR4 (N9442, N9433, N4534, N3694, N1633);
nor NOR3 (N9443, N9430, N3061, N301);
xor XOR2 (N9444, N9434, N4518);
xor XOR2 (N9445, N9444, N6628);
nor NOR2 (N9446, N9445, N3493);
xor XOR2 (N9447, N9439, N7657);
buf BUF1 (N9448, N9424);
nor NOR3 (N9449, N9437, N7861, N250);
nor NOR2 (N9450, N9449, N3345);
nor NOR4 (N9451, N9443, N2125, N768, N7937);
xor XOR2 (N9452, N9417, N1836);
nor NOR2 (N9453, N9441, N5011);
or OR2 (N9454, N9446, N7504);
nor NOR2 (N9455, N9451, N6431);
nor NOR2 (N9456, N9454, N6070);
not NOT1 (N9457, N9431);
and AND2 (N9458, N9425, N8063);
nand NAND2 (N9459, N9452, N6522);
or OR3 (N9460, N9458, N5538, N5185);
or OR4 (N9461, N9455, N3733, N1329, N5127);
and AND3 (N9462, N9450, N2076, N7246);
buf BUF1 (N9463, N9462);
not NOT1 (N9464, N9461);
buf BUF1 (N9465, N9460);
buf BUF1 (N9466, N9447);
nor NOR2 (N9467, N9459, N4989);
xor XOR2 (N9468, N9457, N5151);
nor NOR4 (N9469, N9464, N4397, N550, N7648);
buf BUF1 (N9470, N9456);
nor NOR3 (N9471, N9468, N2793, N436);
xor XOR2 (N9472, N9469, N7829);
xor XOR2 (N9473, N9465, N4451);
nor NOR4 (N9474, N9473, N3107, N611, N1797);
and AND2 (N9475, N9453, N9089);
xor XOR2 (N9476, N9467, N6617);
nand NAND4 (N9477, N9474, N7009, N8031, N3519);
and AND2 (N9478, N9463, N3844);
buf BUF1 (N9479, N9476);
nand NAND4 (N9480, N9466, N3794, N8115, N5715);
or OR3 (N9481, N9475, N7815, N2450);
and AND2 (N9482, N9471, N4388);
nand NAND2 (N9483, N9472, N8614);
buf BUF1 (N9484, N9448);
nor NOR2 (N9485, N9478, N2429);
buf BUF1 (N9486, N9481);
buf BUF1 (N9487, N9480);
buf BUF1 (N9488, N9482);
and AND3 (N9489, N9442, N5922, N435);
nand NAND4 (N9490, N9485, N1951, N5487, N692);
nor NOR3 (N9491, N9487, N1953, N2942);
not NOT1 (N9492, N9484);
xor XOR2 (N9493, N9486, N9174);
nand NAND3 (N9494, N9488, N8117, N1926);
buf BUF1 (N9495, N9470);
xor XOR2 (N9496, N9490, N7421);
xor XOR2 (N9497, N9496, N3993);
and AND3 (N9498, N9479, N790, N8820);
or OR4 (N9499, N9491, N3369, N92, N2163);
and AND4 (N9500, N9495, N9146, N3250, N6268);
xor XOR2 (N9501, N9497, N6935);
buf BUF1 (N9502, N9499);
nand NAND3 (N9503, N9493, N7562, N7506);
and AND4 (N9504, N9489, N3442, N1116, N3015);
nand NAND2 (N9505, N9477, N3297);
xor XOR2 (N9506, N9502, N1929);
xor XOR2 (N9507, N9500, N133);
nor NOR3 (N9508, N9501, N8442, N9243);
xor XOR2 (N9509, N9504, N4631);
buf BUF1 (N9510, N9498);
nor NOR4 (N9511, N9507, N1944, N8405, N8138);
buf BUF1 (N9512, N9508);
buf BUF1 (N9513, N9494);
and AND3 (N9514, N9503, N1543, N3806);
nor NOR3 (N9515, N9505, N6475, N5252);
nor NOR3 (N9516, N9511, N5416, N8365);
buf BUF1 (N9517, N9506);
nor NOR2 (N9518, N9515, N1629);
and AND3 (N9519, N9509, N1439, N8424);
not NOT1 (N9520, N9492);
nor NOR4 (N9521, N9520, N1933, N3552, N4109);
buf BUF1 (N9522, N9483);
nand NAND4 (N9523, N9522, N3764, N9440, N552);
nand NAND3 (N9524, N9516, N8083, N389);
nand NAND2 (N9525, N9521, N4776);
or OR2 (N9526, N9513, N32);
and AND3 (N9527, N9526, N2846, N6361);
and AND4 (N9528, N9517, N9447, N6462, N592);
nand NAND3 (N9529, N9512, N646, N555);
nor NOR4 (N9530, N9523, N4377, N8979, N5243);
nand NAND4 (N9531, N9529, N4274, N8969, N5969);
buf BUF1 (N9532, N9514);
and AND3 (N9533, N9531, N1010, N6134);
xor XOR2 (N9534, N9533, N7121);
not NOT1 (N9535, N9532);
and AND3 (N9536, N9518, N7694, N7012);
or OR2 (N9537, N9527, N154);
nor NOR3 (N9538, N9530, N8124, N3629);
xor XOR2 (N9539, N9519, N2848);
buf BUF1 (N9540, N9525);
nor NOR4 (N9541, N9535, N7780, N267, N6811);
xor XOR2 (N9542, N9537, N6278);
buf BUF1 (N9543, N9528);
buf BUF1 (N9544, N9538);
and AND4 (N9545, N9542, N6506, N1978, N5316);
buf BUF1 (N9546, N9510);
or OR4 (N9547, N9524, N4292, N7508, N2599);
nor NOR3 (N9548, N9545, N1727, N5547);
nor NOR4 (N9549, N9546, N8693, N1761, N3028);
nand NAND3 (N9550, N9548, N5828, N7994);
buf BUF1 (N9551, N9547);
nand NAND4 (N9552, N9543, N2873, N921, N6439);
xor XOR2 (N9553, N9549, N3917);
nor NOR3 (N9554, N9550, N4097, N1672);
and AND2 (N9555, N9541, N7868);
nand NAND3 (N9556, N9552, N3043, N4937);
nor NOR3 (N9557, N9556, N8673, N2236);
nor NOR3 (N9558, N9544, N1074, N1652);
xor XOR2 (N9559, N9540, N7230);
and AND4 (N9560, N9557, N7885, N5417, N4199);
buf BUF1 (N9561, N9554);
nand NAND3 (N9562, N9551, N7558, N4661);
nor NOR3 (N9563, N9560, N9126, N8254);
or OR3 (N9564, N9536, N577, N749);
and AND4 (N9565, N9553, N2629, N4708, N8539);
or OR2 (N9566, N9555, N8024);
xor XOR2 (N9567, N9563, N4490);
xor XOR2 (N9568, N9558, N4402);
buf BUF1 (N9569, N9565);
or OR4 (N9570, N9561, N8548, N7669, N1082);
xor XOR2 (N9571, N9562, N4246);
nor NOR3 (N9572, N9566, N5507, N6051);
xor XOR2 (N9573, N9539, N759);
or OR3 (N9574, N9534, N7720, N4412);
nor NOR4 (N9575, N9564, N5548, N714, N5276);
nand NAND4 (N9576, N9567, N3563, N6889, N2317);
or OR3 (N9577, N9559, N8336, N2559);
or OR4 (N9578, N9570, N5398, N7606, N1789);
not NOT1 (N9579, N9574);
nor NOR2 (N9580, N9575, N8542);
or OR2 (N9581, N9572, N7741);
buf BUF1 (N9582, N9571);
or OR4 (N9583, N9582, N4250, N995, N9341);
nand NAND4 (N9584, N9578, N8654, N2984, N2192);
not NOT1 (N9585, N9583);
nand NAND4 (N9586, N9573, N4805, N5446, N5311);
not NOT1 (N9587, N9585);
xor XOR2 (N9588, N9576, N9000);
and AND2 (N9589, N9586, N9033);
buf BUF1 (N9590, N9568);
and AND3 (N9591, N9590, N953, N2210);
and AND4 (N9592, N9589, N7709, N4114, N3163);
not NOT1 (N9593, N9584);
nand NAND4 (N9594, N9577, N571, N2485, N7423);
nand NAND2 (N9595, N9593, N4743);
nand NAND3 (N9596, N9592, N3961, N739);
nand NAND4 (N9597, N9579, N9447, N1198, N371);
and AND2 (N9598, N9594, N5509);
nand NAND2 (N9599, N9587, N6301);
and AND4 (N9600, N9595, N653, N6280, N5388);
buf BUF1 (N9601, N9591);
nor NOR4 (N9602, N9580, N500, N5415, N287);
xor XOR2 (N9603, N9588, N8556);
and AND2 (N9604, N9599, N1026);
and AND2 (N9605, N9604, N1118);
buf BUF1 (N9606, N9569);
not NOT1 (N9607, N9600);
xor XOR2 (N9608, N9601, N1916);
or OR4 (N9609, N9605, N6157, N2987, N4546);
nand NAND3 (N9610, N9609, N5296, N7167);
nand NAND4 (N9611, N9607, N3894, N761, N9190);
xor XOR2 (N9612, N9598, N5926);
xor XOR2 (N9613, N9602, N1743);
and AND4 (N9614, N9611, N6559, N7310, N4866);
and AND4 (N9615, N9603, N7706, N4636, N5817);
not NOT1 (N9616, N9615);
nor NOR2 (N9617, N9610, N4587);
nand NAND2 (N9618, N9617, N8858);
nand NAND3 (N9619, N9612, N5823, N3298);
xor XOR2 (N9620, N9606, N1048);
and AND3 (N9621, N9613, N5763, N4013);
nand NAND3 (N9622, N9616, N971, N2450);
or OR3 (N9623, N9614, N1127, N2956);
buf BUF1 (N9624, N9619);
and AND2 (N9625, N9623, N6751);
buf BUF1 (N9626, N9621);
nor NOR2 (N9627, N9620, N6901);
or OR3 (N9628, N9627, N8626, N9337);
or OR3 (N9629, N9622, N7873, N2425);
buf BUF1 (N9630, N9618);
xor XOR2 (N9631, N9597, N2325);
buf BUF1 (N9632, N9628);
nand NAND2 (N9633, N9632, N8636);
nand NAND3 (N9634, N9633, N9136, N7441);
buf BUF1 (N9635, N9634);
xor XOR2 (N9636, N9624, N4731);
xor XOR2 (N9637, N9581, N8300);
and AND2 (N9638, N9631, N5444);
and AND2 (N9639, N9626, N7619);
nor NOR4 (N9640, N9625, N7603, N328, N5598);
nor NOR3 (N9641, N9638, N2895, N5578);
and AND2 (N9642, N9640, N6679);
xor XOR2 (N9643, N9629, N6149);
nand NAND3 (N9644, N9608, N5494, N8932);
nand NAND3 (N9645, N9636, N7538, N7068);
or OR4 (N9646, N9635, N7525, N3172, N7896);
and AND4 (N9647, N9596, N8200, N2956, N6248);
nand NAND2 (N9648, N9642, N8955);
xor XOR2 (N9649, N9646, N1208);
buf BUF1 (N9650, N9645);
and AND2 (N9651, N9639, N3915);
and AND3 (N9652, N9637, N5118, N9358);
and AND4 (N9653, N9641, N7954, N1651, N1759);
nor NOR2 (N9654, N9653, N7253);
not NOT1 (N9655, N9650);
buf BUF1 (N9656, N9652);
nor NOR3 (N9657, N9655, N9230, N6251);
nor NOR2 (N9658, N9649, N7043);
buf BUF1 (N9659, N9657);
or OR2 (N9660, N9648, N7590);
buf BUF1 (N9661, N9659);
nor NOR3 (N9662, N9644, N1996, N8937);
not NOT1 (N9663, N9658);
and AND2 (N9664, N9647, N4710);
not NOT1 (N9665, N9654);
nor NOR4 (N9666, N9665, N2569, N7443, N9402);
buf BUF1 (N9667, N9643);
not NOT1 (N9668, N9656);
and AND3 (N9669, N9667, N1911, N991);
or OR2 (N9670, N9666, N1992);
xor XOR2 (N9671, N9630, N7524);
buf BUF1 (N9672, N9670);
or OR4 (N9673, N9664, N7050, N8884, N6923);
or OR2 (N9674, N9662, N606);
nor NOR3 (N9675, N9672, N4038, N5496);
nor NOR3 (N9676, N9671, N5947, N4191);
xor XOR2 (N9677, N9675, N4419);
buf BUF1 (N9678, N9661);
not NOT1 (N9679, N9677);
or OR2 (N9680, N9679, N9112);
xor XOR2 (N9681, N9663, N6348);
nor NOR3 (N9682, N9674, N9377, N2925);
not NOT1 (N9683, N9678);
nor NOR3 (N9684, N9669, N2521, N3021);
or OR2 (N9685, N9680, N4829);
not NOT1 (N9686, N9668);
and AND3 (N9687, N9682, N9234, N5667);
or OR3 (N9688, N9686, N1919, N1711);
nor NOR3 (N9689, N9685, N8817, N6058);
nand NAND2 (N9690, N9660, N678);
and AND4 (N9691, N9676, N1685, N2874, N3111);
or OR3 (N9692, N9683, N7742, N2981);
xor XOR2 (N9693, N9681, N1162);
and AND3 (N9694, N9687, N292, N5986);
nor NOR3 (N9695, N9693, N4260, N7408);
buf BUF1 (N9696, N9690);
nor NOR4 (N9697, N9689, N5575, N6019, N3321);
nor NOR2 (N9698, N9694, N6059);
buf BUF1 (N9699, N9695);
nand NAND2 (N9700, N9697, N5336);
buf BUF1 (N9701, N9673);
nand NAND2 (N9702, N9698, N342);
nor NOR3 (N9703, N9691, N4941, N9166);
nand NAND3 (N9704, N9692, N7874, N974);
and AND4 (N9705, N9651, N9461, N8319, N7545);
xor XOR2 (N9706, N9699, N8676);
nor NOR4 (N9707, N9684, N8366, N3975, N5054);
nor NOR3 (N9708, N9704, N4488, N1548);
nor NOR4 (N9709, N9700, N6372, N2230, N5092);
and AND3 (N9710, N9703, N3331, N5056);
or OR2 (N9711, N9709, N239);
or OR4 (N9712, N9710, N6614, N80, N3827);
xor XOR2 (N9713, N9708, N7906);
buf BUF1 (N9714, N9706);
nor NOR2 (N9715, N9714, N5700);
nand NAND2 (N9716, N9701, N1255);
nand NAND4 (N9717, N9712, N1486, N713, N4757);
nor NOR4 (N9718, N9715, N6778, N9110, N3795);
nand NAND3 (N9719, N9717, N7852, N2942);
xor XOR2 (N9720, N9713, N8488);
nand NAND2 (N9721, N9705, N1147);
or OR2 (N9722, N9721, N4741);
xor XOR2 (N9723, N9688, N7360);
buf BUF1 (N9724, N9707);
nor NOR2 (N9725, N9720, N3489);
not NOT1 (N9726, N9716);
nand NAND2 (N9727, N9711, N6926);
xor XOR2 (N9728, N9718, N2558);
nand NAND3 (N9729, N9724, N3132, N7408);
or OR3 (N9730, N9722, N6129, N3900);
or OR4 (N9731, N9725, N1803, N7491, N4526);
nor NOR2 (N9732, N9727, N7986);
or OR2 (N9733, N9719, N9423);
xor XOR2 (N9734, N9732, N3349);
xor XOR2 (N9735, N9730, N8118);
buf BUF1 (N9736, N9702);
nand NAND2 (N9737, N9731, N4333);
buf BUF1 (N9738, N9737);
or OR2 (N9739, N9738, N6055);
buf BUF1 (N9740, N9739);
nor NOR2 (N9741, N9728, N4729);
or OR4 (N9742, N9723, N6436, N1855, N5063);
buf BUF1 (N9743, N9735);
nor NOR3 (N9744, N9741, N2418, N2567);
or OR3 (N9745, N9734, N3809, N9586);
nor NOR4 (N9746, N9740, N8923, N2192, N4810);
buf BUF1 (N9747, N9726);
xor XOR2 (N9748, N9746, N9273);
nand NAND4 (N9749, N9729, N3031, N4106, N4850);
xor XOR2 (N9750, N9749, N4068);
or OR3 (N9751, N9696, N4202, N2575);
or OR4 (N9752, N9747, N3344, N7941, N5736);
xor XOR2 (N9753, N9743, N5330);
or OR2 (N9754, N9742, N1519);
and AND3 (N9755, N9748, N4746, N9386);
nor NOR2 (N9756, N9754, N3184);
xor XOR2 (N9757, N9733, N6897);
nor NOR2 (N9758, N9753, N418);
nor NOR4 (N9759, N9756, N3343, N724, N2589);
nand NAND3 (N9760, N9759, N91, N7135);
not NOT1 (N9761, N9752);
buf BUF1 (N9762, N9760);
buf BUF1 (N9763, N9757);
or OR3 (N9764, N9745, N6980, N5467);
and AND4 (N9765, N9764, N218, N3428, N4757);
nor NOR2 (N9766, N9765, N8005);
xor XOR2 (N9767, N9744, N3943);
nand NAND4 (N9768, N9750, N3212, N4119, N6404);
or OR4 (N9769, N9767, N9591, N7972, N2253);
or OR4 (N9770, N9758, N3760, N2424, N9522);
nor NOR4 (N9771, N9762, N7391, N767, N3406);
or OR3 (N9772, N9761, N1393, N1951);
and AND2 (N9773, N9769, N3515);
nor NOR4 (N9774, N9771, N1242, N3580, N2761);
nand NAND2 (N9775, N9773, N6860);
buf BUF1 (N9776, N9775);
nand NAND3 (N9777, N9774, N6813, N3186);
not NOT1 (N9778, N9751);
and AND3 (N9779, N9770, N9236, N3804);
nand NAND2 (N9780, N9763, N9488);
or OR2 (N9781, N9776, N3602);
buf BUF1 (N9782, N9779);
nor NOR4 (N9783, N9736, N5238, N4764, N1770);
and AND4 (N9784, N9781, N7309, N9461, N2380);
not NOT1 (N9785, N9766);
buf BUF1 (N9786, N9777);
or OR3 (N9787, N9755, N3821, N8587);
nand NAND3 (N9788, N9783, N6425, N8637);
xor XOR2 (N9789, N9782, N8454);
buf BUF1 (N9790, N9778);
and AND2 (N9791, N9790, N5791);
nor NOR3 (N9792, N9785, N6429, N3001);
xor XOR2 (N9793, N9789, N5520);
nand NAND4 (N9794, N9784, N1527, N4305, N5829);
and AND2 (N9795, N9794, N1433);
xor XOR2 (N9796, N9792, N5454);
nand NAND3 (N9797, N9780, N6183, N457);
xor XOR2 (N9798, N9797, N2272);
nand NAND4 (N9799, N9791, N1294, N1397, N3831);
or OR2 (N9800, N9788, N1925);
buf BUF1 (N9801, N9795);
nor NOR2 (N9802, N9787, N7561);
xor XOR2 (N9803, N9798, N9595);
buf BUF1 (N9804, N9802);
xor XOR2 (N9805, N9793, N4582);
not NOT1 (N9806, N9800);
and AND3 (N9807, N9804, N6732, N4091);
nor NOR2 (N9808, N9768, N1026);
nand NAND2 (N9809, N9801, N4033);
xor XOR2 (N9810, N9772, N7079);
buf BUF1 (N9811, N9786);
not NOT1 (N9812, N9799);
buf BUF1 (N9813, N9811);
xor XOR2 (N9814, N9812, N8761);
not NOT1 (N9815, N9808);
nor NOR3 (N9816, N9810, N4976, N7045);
or OR3 (N9817, N9813, N3402, N4673);
and AND2 (N9818, N9805, N7386);
nand NAND3 (N9819, N9809, N5412, N3664);
nand NAND4 (N9820, N9807, N5634, N4617, N175);
and AND4 (N9821, N9814, N6764, N9664, N3979);
nand NAND4 (N9822, N9817, N8858, N5114, N1506);
nor NOR3 (N9823, N9822, N7420, N8205);
nand NAND4 (N9824, N9806, N8065, N8175, N8072);
not NOT1 (N9825, N9815);
xor XOR2 (N9826, N9816, N6573);
not NOT1 (N9827, N9796);
not NOT1 (N9828, N9819);
not NOT1 (N9829, N9821);
and AND3 (N9830, N9824, N2285, N1319);
and AND2 (N9831, N9826, N6535);
xor XOR2 (N9832, N9827, N2377);
or OR4 (N9833, N9803, N357, N8191, N7133);
and AND4 (N9834, N9828, N1822, N1043, N3597);
or OR2 (N9835, N9833, N4625);
nand NAND3 (N9836, N9825, N2000, N1797);
nand NAND4 (N9837, N9823, N5285, N5147, N8494);
buf BUF1 (N9838, N9831);
buf BUF1 (N9839, N9832);
and AND2 (N9840, N9836, N9256);
nand NAND2 (N9841, N9838, N2271);
buf BUF1 (N9842, N9820);
xor XOR2 (N9843, N9839, N1132);
not NOT1 (N9844, N9818);
xor XOR2 (N9845, N9844, N8532);
not NOT1 (N9846, N9841);
nand NAND3 (N9847, N9845, N7074, N8984);
not NOT1 (N9848, N9846);
xor XOR2 (N9849, N9834, N503);
buf BUF1 (N9850, N9843);
nand NAND3 (N9851, N9835, N1185, N6853);
nor NOR3 (N9852, N9851, N9735, N2232);
and AND2 (N9853, N9837, N3422);
not NOT1 (N9854, N9849);
nor NOR2 (N9855, N9829, N7911);
nor NOR3 (N9856, N9850, N5046, N3779);
not NOT1 (N9857, N9853);
nor NOR2 (N9858, N9842, N853);
or OR3 (N9859, N9840, N9204, N8842);
and AND4 (N9860, N9852, N2866, N7723, N3792);
not NOT1 (N9861, N9855);
nand NAND2 (N9862, N9859, N916);
or OR2 (N9863, N9848, N33);
or OR2 (N9864, N9857, N49);
and AND2 (N9865, N9862, N2602);
and AND4 (N9866, N9830, N908, N6722, N388);
not NOT1 (N9867, N9856);
or OR2 (N9868, N9860, N2314);
and AND4 (N9869, N9866, N1339, N2187, N8018);
and AND2 (N9870, N9863, N3586);
or OR4 (N9871, N9865, N1699, N648, N5874);
nand NAND4 (N9872, N9854, N8156, N8516, N5494);
nor NOR4 (N9873, N9861, N7797, N7844, N472);
buf BUF1 (N9874, N9871);
buf BUF1 (N9875, N9872);
or OR2 (N9876, N9867, N4956);
and AND2 (N9877, N9858, N2236);
xor XOR2 (N9878, N9847, N940);
or OR3 (N9879, N9877, N2695, N5154);
buf BUF1 (N9880, N9879);
xor XOR2 (N9881, N9870, N1958);
not NOT1 (N9882, N9881);
or OR3 (N9883, N9864, N3161, N7399);
or OR3 (N9884, N9878, N1871, N5861);
buf BUF1 (N9885, N9884);
or OR2 (N9886, N9882, N7082);
not NOT1 (N9887, N9876);
nor NOR2 (N9888, N9874, N1438);
nor NOR3 (N9889, N9886, N8930, N1446);
xor XOR2 (N9890, N9885, N5022);
buf BUF1 (N9891, N9875);
nand NAND3 (N9892, N9883, N2516, N2055);
not NOT1 (N9893, N9891);
nor NOR4 (N9894, N9887, N6718, N8828, N2249);
and AND3 (N9895, N9893, N8415, N1084);
buf BUF1 (N9896, N9889);
or OR3 (N9897, N9892, N1355, N2372);
and AND3 (N9898, N9897, N6376, N1467);
buf BUF1 (N9899, N9880);
nand NAND2 (N9900, N9896, N7453);
not NOT1 (N9901, N9873);
or OR4 (N9902, N9900, N3256, N9729, N6464);
or OR3 (N9903, N9899, N5423, N2657);
and AND3 (N9904, N9894, N7371, N9219);
nand NAND3 (N9905, N9901, N5764, N7965);
not NOT1 (N9906, N9904);
not NOT1 (N9907, N9888);
buf BUF1 (N9908, N9905);
xor XOR2 (N9909, N9903, N2878);
and AND2 (N9910, N9908, N7904);
and AND3 (N9911, N9907, N6379, N731);
nor NOR2 (N9912, N9909, N7881);
buf BUF1 (N9913, N9868);
nand NAND2 (N9914, N9906, N6654);
buf BUF1 (N9915, N9911);
nand NAND4 (N9916, N9902, N2916, N9845, N8939);
xor XOR2 (N9917, N9910, N2216);
xor XOR2 (N9918, N9869, N7077);
nor NOR2 (N9919, N9895, N7865);
buf BUF1 (N9920, N9918);
nand NAND4 (N9921, N9919, N6671, N8222, N4909);
nor NOR4 (N9922, N9912, N5171, N8052, N5327);
and AND3 (N9923, N9913, N4872, N8571);
nor NOR2 (N9924, N9921, N7769);
and AND4 (N9925, N9916, N297, N2113, N7253);
nand NAND2 (N9926, N9898, N5049);
xor XOR2 (N9927, N9914, N1157);
nor NOR4 (N9928, N9926, N7657, N9553, N2632);
buf BUF1 (N9929, N9924);
or OR4 (N9930, N9929, N881, N9155, N4848);
nand NAND2 (N9931, N9917, N614);
or OR4 (N9932, N9925, N2361, N9169, N9138);
nand NAND3 (N9933, N9927, N4578, N3391);
nand NAND4 (N9934, N9920, N6046, N6843, N4570);
nor NOR2 (N9935, N9922, N1024);
xor XOR2 (N9936, N9935, N9349);
and AND2 (N9937, N9931, N1383);
and AND4 (N9938, N9934, N1212, N8210, N5464);
nor NOR3 (N9939, N9936, N958, N8311);
nand NAND4 (N9940, N9932, N5369, N3980, N4517);
or OR3 (N9941, N9937, N681, N2260);
nor NOR3 (N9942, N9915, N2779, N5147);
nand NAND4 (N9943, N9938, N7766, N4964, N7318);
and AND3 (N9944, N9930, N9133, N8865);
and AND4 (N9945, N9940, N732, N5771, N819);
nand NAND2 (N9946, N9939, N9878);
and AND3 (N9947, N9942, N7208, N2534);
nand NAND3 (N9948, N9944, N418, N7361);
nand NAND3 (N9949, N9923, N8633, N8859);
and AND3 (N9950, N9941, N7494, N2316);
xor XOR2 (N9951, N9945, N3483);
and AND2 (N9952, N9947, N2277);
or OR4 (N9953, N9949, N4883, N7744, N8621);
not NOT1 (N9954, N9948);
nand NAND2 (N9955, N9952, N4024);
or OR2 (N9956, N9955, N6398);
buf BUF1 (N9957, N9946);
or OR4 (N9958, N9950, N4558, N8270, N694);
nand NAND3 (N9959, N9943, N5040, N8007);
and AND2 (N9960, N9959, N9569);
nand NAND2 (N9961, N9951, N1909);
nand NAND4 (N9962, N9953, N8681, N3169, N4289);
nand NAND3 (N9963, N9957, N4479, N3011);
buf BUF1 (N9964, N9958);
not NOT1 (N9965, N9962);
xor XOR2 (N9966, N9960, N4010);
nand NAND4 (N9967, N9961, N77, N8416, N2563);
xor XOR2 (N9968, N9954, N6976);
xor XOR2 (N9969, N9928, N1553);
xor XOR2 (N9970, N9967, N3820);
not NOT1 (N9971, N9933);
nor NOR2 (N9972, N9966, N8962);
buf BUF1 (N9973, N9965);
or OR2 (N9974, N9890, N1935);
not NOT1 (N9975, N9969);
buf BUF1 (N9976, N9956);
nand NAND3 (N9977, N9970, N3638, N9303);
nor NOR2 (N9978, N9963, N7052);
nand NAND3 (N9979, N9973, N8395, N2829);
not NOT1 (N9980, N9971);
nand NAND2 (N9981, N9980, N6604);
and AND4 (N9982, N9972, N5106, N1166, N8196);
or OR3 (N9983, N9982, N2414, N2976);
nand NAND3 (N9984, N9981, N2989, N5353);
buf BUF1 (N9985, N9979);
nand NAND2 (N9986, N9976, N3872);
or OR4 (N9987, N9977, N5208, N8947, N2371);
or OR2 (N9988, N9985, N3716);
not NOT1 (N9989, N9984);
nand NAND3 (N9990, N9989, N6390, N7885);
buf BUF1 (N9991, N9983);
xor XOR2 (N9992, N9990, N1326);
xor XOR2 (N9993, N9987, N8806);
and AND4 (N9994, N9993, N4386, N3495, N9583);
buf BUF1 (N9995, N9991);
xor XOR2 (N9996, N9964, N8083);
not NOT1 (N9997, N9995);
nor NOR2 (N9998, N9992, N1007);
and AND4 (N9999, N9974, N7166, N8032, N2439);
and AND4 (N10000, N9997, N2042, N1969, N6430);
xor XOR2 (N10001, N9968, N2294);
xor XOR2 (N10002, N10001, N961);
or OR3 (N10003, N9998, N5709, N8367);
nor NOR4 (N10004, N10000, N6196, N1999, N1837);
buf BUF1 (N10005, N9986);
or OR2 (N10006, N9994, N7017);
not NOT1 (N10007, N10006);
or OR3 (N10008, N10007, N2202, N6819);
and AND2 (N10009, N9996, N5192);
nor NOR3 (N10010, N10004, N6835, N8215);
xor XOR2 (N10011, N9999, N6206);
xor XOR2 (N10012, N9988, N8993);
or OR3 (N10013, N9978, N3760, N6800);
nand NAND3 (N10014, N10003, N4017, N7477);
xor XOR2 (N10015, N10011, N4448);
nand NAND4 (N10016, N10012, N474, N4552, N1976);
and AND3 (N10017, N10008, N485, N1065);
buf BUF1 (N10018, N10005);
not NOT1 (N10019, N10013);
not NOT1 (N10020, N10016);
or OR4 (N10021, N10009, N9422, N6283, N5964);
buf BUF1 (N10022, N10018);
or OR2 (N10023, N10002, N8144);
xor XOR2 (N10024, N10014, N6787);
nand NAND4 (N10025, N10020, N4444, N4444, N1772);
nor NOR3 (N10026, N10017, N9593, N3692);
or OR3 (N10027, N10010, N9666, N5597);
not NOT1 (N10028, N9975);
xor XOR2 (N10029, N10024, N9536);
not NOT1 (N10030, N10028);
xor XOR2 (N10031, N10025, N7066);
nand NAND3 (N10032, N10029, N913, N1622);
nand NAND3 (N10033, N10032, N1043, N2221);
nand NAND4 (N10034, N10033, N4503, N8534, N4120);
not NOT1 (N10035, N10015);
and AND4 (N10036, N10026, N6303, N6477, N381);
buf BUF1 (N10037, N10022);
or OR2 (N10038, N10031, N5182);
and AND4 (N10039, N10035, N7925, N854, N4022);
or OR3 (N10040, N10037, N8145, N6160);
and AND3 (N10041, N10039, N7352, N4147);
nor NOR3 (N10042, N10040, N1877, N8224);
xor XOR2 (N10043, N10023, N4752);
xor XOR2 (N10044, N10021, N2647);
and AND4 (N10045, N10027, N8394, N2211, N3680);
xor XOR2 (N10046, N10019, N6724);
buf BUF1 (N10047, N10038);
and AND2 (N10048, N10046, N4794);
nor NOR4 (N10049, N10034, N8543, N14, N6838);
and AND4 (N10050, N10048, N78, N3558, N7342);
or OR4 (N10051, N10049, N7348, N1212, N6839);
nand NAND3 (N10052, N10036, N7383, N1957);
buf BUF1 (N10053, N10030);
and AND3 (N10054, N10051, N3530, N2249);
or OR2 (N10055, N10052, N3388);
or OR4 (N10056, N10042, N4584, N4568, N1687);
xor XOR2 (N10057, N10056, N2933);
xor XOR2 (N10058, N10043, N4114);
or OR3 (N10059, N10053, N6896, N6299);
or OR4 (N10060, N10047, N9927, N3276, N5145);
nor NOR2 (N10061, N10060, N2629);
xor XOR2 (N10062, N10058, N8459);
or OR2 (N10063, N10055, N5124);
not NOT1 (N10064, N10044);
buf BUF1 (N10065, N10063);
xor XOR2 (N10066, N10054, N5260);
nor NOR3 (N10067, N10062, N5104, N6379);
not NOT1 (N10068, N10064);
and AND3 (N10069, N10065, N7448, N5182);
buf BUF1 (N10070, N10050);
and AND2 (N10071, N10066, N8225);
and AND2 (N10072, N10061, N4499);
and AND2 (N10073, N10059, N6462);
not NOT1 (N10074, N10068);
not NOT1 (N10075, N10071);
and AND2 (N10076, N10070, N6529);
buf BUF1 (N10077, N10067);
nor NOR3 (N10078, N10076, N5991, N186);
not NOT1 (N10079, N10072);
not NOT1 (N10080, N10069);
buf BUF1 (N10081, N10074);
not NOT1 (N10082, N10041);
nand NAND2 (N10083, N10045, N2376);
xor XOR2 (N10084, N10082, N691);
and AND4 (N10085, N10081, N5945, N6725, N4966);
xor XOR2 (N10086, N10077, N4600);
not NOT1 (N10087, N10078);
not NOT1 (N10088, N10079);
and AND2 (N10089, N10085, N6685);
xor XOR2 (N10090, N10084, N505);
nand NAND3 (N10091, N10087, N708, N7304);
buf BUF1 (N10092, N10080);
xor XOR2 (N10093, N10090, N2569);
nand NAND4 (N10094, N10093, N9738, N3971, N8542);
xor XOR2 (N10095, N10083, N4526);
or OR4 (N10096, N10088, N7995, N8518, N6776);
and AND3 (N10097, N10091, N7238, N3244);
not NOT1 (N10098, N10092);
xor XOR2 (N10099, N10094, N7354);
nand NAND2 (N10100, N10089, N7681);
nor NOR3 (N10101, N10100, N6033, N9772);
not NOT1 (N10102, N10057);
nand NAND2 (N10103, N10097, N8670);
nand NAND3 (N10104, N10075, N5809, N5880);
buf BUF1 (N10105, N10073);
nor NOR4 (N10106, N10102, N353, N9372, N9030);
not NOT1 (N10107, N10106);
nor NOR2 (N10108, N10095, N4607);
nand NAND2 (N10109, N10103, N9405);
xor XOR2 (N10110, N10104, N6141);
nand NAND4 (N10111, N10098, N1837, N8310, N7203);
xor XOR2 (N10112, N10110, N3096);
and AND2 (N10113, N10109, N1589);
nand NAND4 (N10114, N10112, N3374, N1154, N3589);
and AND4 (N10115, N10113, N7811, N331, N7918);
not NOT1 (N10116, N10114);
nor NOR4 (N10117, N10108, N1, N6990, N4895);
not NOT1 (N10118, N10107);
nand NAND3 (N10119, N10086, N8019, N3662);
not NOT1 (N10120, N10115);
buf BUF1 (N10121, N10116);
or OR3 (N10122, N10120, N5960, N9519);
nand NAND4 (N10123, N10122, N990, N9808, N7482);
not NOT1 (N10124, N10105);
buf BUF1 (N10125, N10124);
not NOT1 (N10126, N10119);
xor XOR2 (N10127, N10125, N7075);
buf BUF1 (N10128, N10127);
nor NOR2 (N10129, N10128, N576);
xor XOR2 (N10130, N10096, N4660);
nor NOR3 (N10131, N10111, N7007, N289);
xor XOR2 (N10132, N10130, N1851);
nand NAND3 (N10133, N10099, N309, N1678);
and AND3 (N10134, N10133, N911, N5406);
or OR2 (N10135, N10134, N3280);
or OR2 (N10136, N10117, N4639);
xor XOR2 (N10137, N10132, N1638);
not NOT1 (N10138, N10136);
nor NOR2 (N10139, N10121, N1128);
nor NOR4 (N10140, N10118, N7729, N7986, N7239);
buf BUF1 (N10141, N10135);
nand NAND2 (N10142, N10101, N9879);
and AND4 (N10143, N10129, N7244, N5110, N6932);
buf BUF1 (N10144, N10141);
not NOT1 (N10145, N10143);
buf BUF1 (N10146, N10131);
not NOT1 (N10147, N10126);
nand NAND3 (N10148, N10144, N2786, N10072);
buf BUF1 (N10149, N10139);
nand NAND3 (N10150, N10138, N3515, N8605);
not NOT1 (N10151, N10148);
xor XOR2 (N10152, N10149, N4062);
not NOT1 (N10153, N10137);
and AND4 (N10154, N10145, N7286, N2345, N8537);
buf BUF1 (N10155, N10140);
buf BUF1 (N10156, N10151);
and AND3 (N10157, N10123, N664, N2866);
nor NOR4 (N10158, N10147, N10003, N4848, N6973);
buf BUF1 (N10159, N10155);
and AND2 (N10160, N10153, N266);
or OR2 (N10161, N10154, N4711);
or OR4 (N10162, N10158, N1221, N8560, N7794);
nor NOR3 (N10163, N10150, N8358, N6407);
buf BUF1 (N10164, N10156);
nand NAND3 (N10165, N10163, N1621, N6623);
nand NAND4 (N10166, N10164, N5508, N8808, N9291);
or OR4 (N10167, N10159, N4355, N5654, N2781);
nor NOR3 (N10168, N10157, N4595, N7431);
xor XOR2 (N10169, N10168, N6963);
nor NOR4 (N10170, N10142, N7781, N3616, N9242);
and AND3 (N10171, N10161, N5252, N3865);
not NOT1 (N10172, N10162);
and AND3 (N10173, N10146, N4796, N1196);
or OR2 (N10174, N10166, N3002);
nor NOR3 (N10175, N10160, N2720, N902);
nor NOR2 (N10176, N10152, N1176);
not NOT1 (N10177, N10170);
or OR2 (N10178, N10172, N5590);
and AND3 (N10179, N10174, N4865, N655);
and AND2 (N10180, N10179, N6049);
nor NOR4 (N10181, N10177, N9284, N7014, N2663);
not NOT1 (N10182, N10169);
nand NAND4 (N10183, N10171, N5412, N5856, N3242);
and AND4 (N10184, N10183, N8388, N9640, N1515);
or OR4 (N10185, N10182, N270, N1426, N2302);
nor NOR4 (N10186, N10167, N6343, N5518, N3418);
not NOT1 (N10187, N10178);
not NOT1 (N10188, N10181);
nor NOR2 (N10189, N10176, N4073);
nand NAND2 (N10190, N10165, N2785);
buf BUF1 (N10191, N10184);
nor NOR3 (N10192, N10175, N4663, N2435);
nand NAND4 (N10193, N10180, N2096, N9739, N5131);
not NOT1 (N10194, N10193);
and AND3 (N10195, N10188, N1410, N6167);
nand NAND2 (N10196, N10190, N8985);
buf BUF1 (N10197, N10187);
buf BUF1 (N10198, N10173);
buf BUF1 (N10199, N10196);
or OR3 (N10200, N10192, N5283, N671);
or OR4 (N10201, N10199, N2389, N7948, N1035);
nand NAND4 (N10202, N10191, N8124, N889, N6857);
or OR4 (N10203, N10186, N3167, N1392, N8251);
nor NOR4 (N10204, N10195, N6404, N3897, N160);
or OR4 (N10205, N10185, N2556, N4056, N1693);
and AND4 (N10206, N10194, N8595, N7545, N6708);
nor NOR3 (N10207, N10201, N8649, N5657);
nand NAND2 (N10208, N10202, N1850);
nand NAND2 (N10209, N10189, N216);
or OR4 (N10210, N10205, N6591, N8854, N9299);
buf BUF1 (N10211, N10198);
not NOT1 (N10212, N10207);
and AND2 (N10213, N10212, N8999);
and AND4 (N10214, N10206, N4909, N6614, N8260);
not NOT1 (N10215, N10214);
nand NAND3 (N10216, N10209, N2498, N9631);
nor NOR3 (N10217, N10211, N7659, N8084);
or OR2 (N10218, N10203, N2826);
or OR4 (N10219, N10217, N5746, N8888, N9838);
buf BUF1 (N10220, N10208);
not NOT1 (N10221, N10220);
xor XOR2 (N10222, N10221, N7997);
xor XOR2 (N10223, N10204, N7526);
nor NOR3 (N10224, N10222, N4489, N7766);
nand NAND2 (N10225, N10200, N4919);
nor NOR2 (N10226, N10223, N7858);
nand NAND2 (N10227, N10226, N3416);
nand NAND3 (N10228, N10210, N4964, N213);
nor NOR3 (N10229, N10228, N8487, N6863);
not NOT1 (N10230, N10229);
nor NOR3 (N10231, N10215, N8560, N1788);
and AND3 (N10232, N10225, N1784, N7758);
buf BUF1 (N10233, N10224);
not NOT1 (N10234, N10213);
and AND4 (N10235, N10218, N8138, N5281, N8617);
xor XOR2 (N10236, N10235, N8542);
buf BUF1 (N10237, N10219);
nand NAND4 (N10238, N10237, N4035, N4929, N5168);
or OR2 (N10239, N10231, N614);
xor XOR2 (N10240, N10239, N9982);
or OR4 (N10241, N10216, N4927, N9439, N724);
xor XOR2 (N10242, N10227, N5782);
or OR3 (N10243, N10230, N5111, N3933);
xor XOR2 (N10244, N10240, N6671);
buf BUF1 (N10245, N10244);
nor NOR2 (N10246, N10242, N362);
nand NAND3 (N10247, N10238, N5351, N1948);
and AND4 (N10248, N10246, N2160, N7991, N9155);
not NOT1 (N10249, N10243);
xor XOR2 (N10250, N10245, N227);
nor NOR2 (N10251, N10234, N4628);
nor NOR2 (N10252, N10232, N7515);
xor XOR2 (N10253, N10248, N1479);
nor NOR4 (N10254, N10249, N3722, N5069, N3602);
and AND3 (N10255, N10253, N6780, N5421);
or OR4 (N10256, N10251, N1901, N1768, N1300);
buf BUF1 (N10257, N10255);
not NOT1 (N10258, N10241);
and AND4 (N10259, N10247, N6009, N3576, N2740);
not NOT1 (N10260, N10236);
nor NOR2 (N10261, N10254, N9465);
xor XOR2 (N10262, N10252, N2826);
not NOT1 (N10263, N10258);
and AND3 (N10264, N10259, N8751, N9072);
and AND4 (N10265, N10260, N6709, N9428, N6063);
and AND3 (N10266, N10256, N714, N1909);
or OR4 (N10267, N10265, N4558, N6347, N6326);
not NOT1 (N10268, N10250);
buf BUF1 (N10269, N10257);
buf BUF1 (N10270, N10269);
nand NAND2 (N10271, N10261, N5926);
xor XOR2 (N10272, N10270, N4563);
and AND4 (N10273, N10262, N3313, N7372, N3949);
or OR2 (N10274, N10273, N4668);
buf BUF1 (N10275, N10268);
xor XOR2 (N10276, N10266, N2464);
nand NAND4 (N10277, N10233, N8642, N6896, N2135);
nor NOR2 (N10278, N10264, N8815);
nand NAND2 (N10279, N10278, N1948);
or OR3 (N10280, N10275, N4219, N3129);
or OR2 (N10281, N10274, N3474);
and AND3 (N10282, N10263, N115, N6068);
and AND3 (N10283, N10277, N1082, N2655);
xor XOR2 (N10284, N10271, N3477);
buf BUF1 (N10285, N10197);
buf BUF1 (N10286, N10282);
buf BUF1 (N10287, N10276);
nand NAND4 (N10288, N10279, N8078, N2245, N3453);
or OR4 (N10289, N10280, N2766, N2360, N4239);
buf BUF1 (N10290, N10267);
and AND3 (N10291, N10283, N5025, N2850);
nand NAND3 (N10292, N10287, N5889, N8934);
not NOT1 (N10293, N10285);
xor XOR2 (N10294, N10291, N9285);
nand NAND2 (N10295, N10289, N6110);
nand NAND3 (N10296, N10290, N3588, N971);
not NOT1 (N10297, N10286);
xor XOR2 (N10298, N10281, N3756);
or OR2 (N10299, N10296, N2623);
xor XOR2 (N10300, N10284, N1528);
or OR2 (N10301, N10295, N67);
nand NAND2 (N10302, N10298, N4675);
xor XOR2 (N10303, N10297, N8377);
or OR4 (N10304, N10272, N1190, N387, N1918);
buf BUF1 (N10305, N10301);
or OR3 (N10306, N10294, N8351, N3898);
and AND2 (N10307, N10293, N10128);
not NOT1 (N10308, N10305);
and AND4 (N10309, N10300, N5911, N2571, N6727);
nor NOR2 (N10310, N10299, N1934);
and AND3 (N10311, N10310, N5733, N1977);
and AND3 (N10312, N10306, N39, N3274);
and AND3 (N10313, N10302, N9431, N5208);
nor NOR4 (N10314, N10307, N986, N6304, N7495);
not NOT1 (N10315, N10308);
nor NOR4 (N10316, N10303, N7779, N2688, N8507);
or OR2 (N10317, N10304, N187);
and AND2 (N10318, N10312, N7727);
buf BUF1 (N10319, N10309);
not NOT1 (N10320, N10311);
not NOT1 (N10321, N10313);
not NOT1 (N10322, N10318);
buf BUF1 (N10323, N10321);
xor XOR2 (N10324, N10317, N3774);
buf BUF1 (N10325, N10288);
buf BUF1 (N10326, N10292);
buf BUF1 (N10327, N10324);
buf BUF1 (N10328, N10316);
not NOT1 (N10329, N10315);
buf BUF1 (N10330, N10326);
nand NAND2 (N10331, N10325, N2320);
buf BUF1 (N10332, N10328);
nand NAND3 (N10333, N10320, N9920, N7288);
nor NOR4 (N10334, N10314, N2076, N3509, N4262);
buf BUF1 (N10335, N10333);
and AND3 (N10336, N10322, N2532, N2412);
buf BUF1 (N10337, N10329);
buf BUF1 (N10338, N10330);
xor XOR2 (N10339, N10334, N787);
nor NOR2 (N10340, N10339, N8920);
nor NOR2 (N10341, N10332, N8613);
buf BUF1 (N10342, N10323);
and AND4 (N10343, N10337, N9942, N2447, N9402);
not NOT1 (N10344, N10331);
and AND4 (N10345, N10341, N3925, N2760, N9360);
and AND3 (N10346, N10345, N1911, N4281);
buf BUF1 (N10347, N10344);
not NOT1 (N10348, N10340);
and AND4 (N10349, N10346, N2461, N10260, N1688);
buf BUF1 (N10350, N10336);
and AND4 (N10351, N10349, N4482, N245, N4577);
buf BUF1 (N10352, N10351);
nand NAND2 (N10353, N10342, N2245);
or OR2 (N10354, N10343, N6245);
buf BUF1 (N10355, N10338);
buf BUF1 (N10356, N10353);
nor NOR2 (N10357, N10348, N525);
nor NOR2 (N10358, N10352, N4876);
or OR4 (N10359, N10319, N885, N867, N6342);
nand NAND3 (N10360, N10327, N478, N5489);
nand NAND3 (N10361, N10354, N2559, N1024);
or OR3 (N10362, N10357, N6046, N1218);
and AND3 (N10363, N10355, N9396, N1664);
xor XOR2 (N10364, N10363, N3156);
xor XOR2 (N10365, N10358, N1173);
buf BUF1 (N10366, N10360);
xor XOR2 (N10367, N10356, N1759);
nand NAND3 (N10368, N10359, N5043, N6248);
or OR4 (N10369, N10347, N6502, N9950, N5478);
not NOT1 (N10370, N10367);
and AND4 (N10371, N10364, N4249, N275, N1768);
or OR4 (N10372, N10368, N8446, N5747, N6497);
and AND2 (N10373, N10362, N3402);
not NOT1 (N10374, N10372);
nor NOR2 (N10375, N10335, N2065);
and AND4 (N10376, N10370, N1110, N2593, N5421);
buf BUF1 (N10377, N10374);
or OR2 (N10378, N10373, N8362);
not NOT1 (N10379, N10377);
or OR3 (N10380, N10369, N8144, N631);
nand NAND2 (N10381, N10350, N612);
nand NAND4 (N10382, N10365, N7213, N593, N1150);
or OR3 (N10383, N10366, N6539, N4275);
and AND4 (N10384, N10379, N9777, N420, N9263);
xor XOR2 (N10385, N10375, N2605);
buf BUF1 (N10386, N10376);
not NOT1 (N10387, N10382);
xor XOR2 (N10388, N10387, N478);
nor NOR2 (N10389, N10385, N4408);
xor XOR2 (N10390, N10384, N4555);
and AND4 (N10391, N10386, N5994, N8660, N5572);
and AND3 (N10392, N10390, N9436, N9153);
and AND3 (N10393, N10383, N9327, N9565);
xor XOR2 (N10394, N10392, N8216);
xor XOR2 (N10395, N10361, N5820);
nor NOR4 (N10396, N10393, N2060, N9733, N9009);
nand NAND4 (N10397, N10396, N10048, N2683, N5306);
and AND4 (N10398, N10395, N6605, N1179, N3940);
or OR2 (N10399, N10388, N4165);
or OR2 (N10400, N10381, N5778);
not NOT1 (N10401, N10399);
nor NOR2 (N10402, N10401, N8532);
nor NOR4 (N10403, N10371, N2455, N2219, N4695);
not NOT1 (N10404, N10398);
nand NAND2 (N10405, N10378, N8430);
xor XOR2 (N10406, N10397, N758);
or OR3 (N10407, N10380, N5351, N456);
and AND3 (N10408, N10389, N3647, N2803);
and AND3 (N10409, N10391, N9423, N2990);
and AND2 (N10410, N10404, N807);
buf BUF1 (N10411, N10405);
or OR4 (N10412, N10394, N6847, N4633, N1872);
not NOT1 (N10413, N10400);
not NOT1 (N10414, N10406);
or OR2 (N10415, N10411, N5080);
not NOT1 (N10416, N10402);
and AND4 (N10417, N10408, N5408, N342, N5421);
xor XOR2 (N10418, N10413, N9896);
or OR3 (N10419, N10409, N2874, N9378);
not NOT1 (N10420, N10418);
nor NOR4 (N10421, N10407, N4673, N7563, N111);
or OR3 (N10422, N10417, N1951, N5459);
or OR4 (N10423, N10419, N9638, N7894, N36);
nor NOR2 (N10424, N10423, N6026);
not NOT1 (N10425, N10403);
xor XOR2 (N10426, N10415, N9246);
buf BUF1 (N10427, N10410);
and AND2 (N10428, N10426, N7218);
nor NOR2 (N10429, N10420, N4485);
nor NOR4 (N10430, N10424, N10051, N1650, N8061);
buf BUF1 (N10431, N10430);
not NOT1 (N10432, N10429);
or OR4 (N10433, N10432, N2875, N5048, N9325);
or OR4 (N10434, N10427, N2935, N6362, N9866);
buf BUF1 (N10435, N10412);
and AND3 (N10436, N10431, N2530, N7856);
buf BUF1 (N10437, N10414);
xor XOR2 (N10438, N10437, N10322);
xor XOR2 (N10439, N10425, N983);
not NOT1 (N10440, N10438);
nand NAND4 (N10441, N10436, N5690, N1235, N10322);
or OR2 (N10442, N10428, N9020);
buf BUF1 (N10443, N10439);
xor XOR2 (N10444, N10442, N3824);
nor NOR4 (N10445, N10434, N6057, N7075, N392);
xor XOR2 (N10446, N10443, N8346);
or OR4 (N10447, N10444, N3386, N689, N7111);
nor NOR2 (N10448, N10416, N600);
not NOT1 (N10449, N10440);
and AND2 (N10450, N10446, N368);
and AND4 (N10451, N10449, N9035, N7501, N5151);
xor XOR2 (N10452, N10450, N6984);
xor XOR2 (N10453, N10452, N4259);
and AND3 (N10454, N10451, N2069, N2068);
not NOT1 (N10455, N10447);
nor NOR2 (N10456, N10421, N2810);
or OR2 (N10457, N10435, N1002);
nor NOR3 (N10458, N10422, N1734, N7518);
xor XOR2 (N10459, N10456, N5055);
nand NAND2 (N10460, N10454, N109);
nor NOR2 (N10461, N10445, N1052);
xor XOR2 (N10462, N10457, N4431);
buf BUF1 (N10463, N10448);
nor NOR2 (N10464, N10433, N5474);
nand NAND3 (N10465, N10453, N5066, N8524);
xor XOR2 (N10466, N10464, N7320);
nand NAND4 (N10467, N10458, N1182, N2749, N3455);
xor XOR2 (N10468, N10460, N7374);
or OR2 (N10469, N10441, N4121);
not NOT1 (N10470, N10463);
not NOT1 (N10471, N10455);
buf BUF1 (N10472, N10461);
xor XOR2 (N10473, N10465, N3777);
xor XOR2 (N10474, N10469, N4780);
not NOT1 (N10475, N10470);
not NOT1 (N10476, N10471);
and AND4 (N10477, N10468, N9117, N459, N7829);
nand NAND2 (N10478, N10472, N7257);
xor XOR2 (N10479, N10466, N3880);
buf BUF1 (N10480, N10478);
not NOT1 (N10481, N10473);
and AND2 (N10482, N10477, N6395);
and AND3 (N10483, N10482, N682, N7860);
buf BUF1 (N10484, N10481);
or OR4 (N10485, N10484, N93, N6387, N10295);
xor XOR2 (N10486, N10459, N10081);
xor XOR2 (N10487, N10476, N9248);
xor XOR2 (N10488, N10479, N378);
and AND4 (N10489, N10467, N136, N7259, N9417);
xor XOR2 (N10490, N10462, N61);
nor NOR3 (N10491, N10488, N1980, N7384);
and AND2 (N10492, N10489, N3521);
xor XOR2 (N10493, N10491, N4892);
nand NAND4 (N10494, N10474, N7620, N7334, N8524);
or OR2 (N10495, N10475, N7038);
not NOT1 (N10496, N10490);
xor XOR2 (N10497, N10492, N3723);
nand NAND4 (N10498, N10487, N296, N10098, N4610);
and AND2 (N10499, N10495, N9498);
nor NOR4 (N10500, N10480, N8993, N4671, N1514);
nand NAND2 (N10501, N10486, N6699);
not NOT1 (N10502, N10494);
not NOT1 (N10503, N10493);
xor XOR2 (N10504, N10483, N7037);
nor NOR4 (N10505, N10502, N6296, N4255, N3821);
or OR4 (N10506, N10496, N8249, N7675, N7885);
or OR4 (N10507, N10500, N3376, N5451, N4168);
buf BUF1 (N10508, N10501);
nor NOR4 (N10509, N10504, N143, N1282, N1952);
buf BUF1 (N10510, N10499);
not NOT1 (N10511, N10503);
or OR4 (N10512, N10497, N9957, N9702, N423);
nor NOR4 (N10513, N10506, N5262, N4301, N6000);
buf BUF1 (N10514, N10509);
xor XOR2 (N10515, N10507, N4111);
not NOT1 (N10516, N10508);
buf BUF1 (N10517, N10505);
buf BUF1 (N10518, N10515);
xor XOR2 (N10519, N10516, N1310);
nand NAND2 (N10520, N10514, N4737);
not NOT1 (N10521, N10512);
buf BUF1 (N10522, N10511);
xor XOR2 (N10523, N10518, N9009);
nand NAND2 (N10524, N10485, N7138);
buf BUF1 (N10525, N10523);
and AND2 (N10526, N10520, N7272);
or OR2 (N10527, N10517, N9576);
nand NAND2 (N10528, N10522, N10104);
or OR4 (N10529, N10527, N7402, N3695, N2012);
nor NOR3 (N10530, N10526, N3732, N8815);
nor NOR2 (N10531, N10525, N9139);
nand NAND2 (N10532, N10528, N5009);
or OR4 (N10533, N10519, N10299, N5736, N6452);
not NOT1 (N10534, N10529);
and AND3 (N10535, N10521, N6484, N8486);
or OR3 (N10536, N10510, N6339, N1877);
and AND4 (N10537, N10532, N6251, N5306, N976);
and AND2 (N10538, N10535, N4964);
nand NAND2 (N10539, N10537, N2482);
or OR2 (N10540, N10533, N2247);
and AND2 (N10541, N10498, N1354);
nand NAND3 (N10542, N10524, N7759, N7794);
nand NAND4 (N10543, N10538, N365, N227, N8100);
buf BUF1 (N10544, N10539);
nand NAND2 (N10545, N10542, N5227);
nor NOR2 (N10546, N10544, N6765);
or OR4 (N10547, N10541, N6804, N961, N1453);
nor NOR2 (N10548, N10545, N6197);
or OR4 (N10549, N10536, N8511, N4519, N2515);
buf BUF1 (N10550, N10543);
buf BUF1 (N10551, N10549);
not NOT1 (N10552, N10548);
buf BUF1 (N10553, N10540);
nand NAND2 (N10554, N10530, N894);
not NOT1 (N10555, N10534);
buf BUF1 (N10556, N10555);
nor NOR2 (N10557, N10513, N4501);
buf BUF1 (N10558, N10552);
and AND2 (N10559, N10550, N4339);
not NOT1 (N10560, N10557);
and AND3 (N10561, N10554, N1291, N2274);
not NOT1 (N10562, N10558);
nor NOR2 (N10563, N10556, N6012);
xor XOR2 (N10564, N10561, N1578);
and AND4 (N10565, N10546, N8279, N82, N10299);
buf BUF1 (N10566, N10547);
nand NAND4 (N10567, N10551, N942, N6522, N4238);
nand NAND4 (N10568, N10562, N10322, N8423, N861);
buf BUF1 (N10569, N10560);
nand NAND2 (N10570, N10531, N2475);
and AND4 (N10571, N10568, N9568, N8350, N930);
and AND4 (N10572, N10571, N4176, N8054, N6755);
buf BUF1 (N10573, N10566);
and AND3 (N10574, N10559, N7539, N1472);
or OR3 (N10575, N10563, N7979, N10063);
xor XOR2 (N10576, N10565, N3878);
not NOT1 (N10577, N10574);
not NOT1 (N10578, N10569);
nand NAND4 (N10579, N10572, N5849, N2412, N1777);
nand NAND2 (N10580, N10577, N1786);
or OR2 (N10581, N10576, N8336);
not NOT1 (N10582, N10579);
nor NOR4 (N10583, N10567, N8226, N8405, N9603);
xor XOR2 (N10584, N10581, N2087);
not NOT1 (N10585, N10582);
buf BUF1 (N10586, N10584);
or OR4 (N10587, N10586, N4369, N9246, N8287);
or OR4 (N10588, N10587, N3057, N5068, N4720);
nor NOR3 (N10589, N10588, N5240, N6764);
nand NAND3 (N10590, N10589, N51, N2219);
xor XOR2 (N10591, N10590, N6629);
nor NOR2 (N10592, N10580, N1291);
buf BUF1 (N10593, N10585);
xor XOR2 (N10594, N10573, N724);
nor NOR4 (N10595, N10583, N465, N6924, N8036);
and AND3 (N10596, N10575, N3967, N8058);
nand NAND2 (N10597, N10553, N8789);
not NOT1 (N10598, N10596);
not NOT1 (N10599, N10597);
nor NOR3 (N10600, N10593, N3204, N7463);
and AND2 (N10601, N10595, N6147);
buf BUF1 (N10602, N10564);
nor NOR3 (N10603, N10602, N5127, N5578);
nand NAND4 (N10604, N10598, N6325, N5517, N3884);
nor NOR3 (N10605, N10570, N9131, N4338);
buf BUF1 (N10606, N10605);
buf BUF1 (N10607, N10603);
xor XOR2 (N10608, N10601, N114);
nand NAND4 (N10609, N10600, N8502, N5081, N3519);
or OR4 (N10610, N10594, N10131, N5607, N7175);
nor NOR2 (N10611, N10608, N275);
nor NOR2 (N10612, N10610, N3521);
nor NOR4 (N10613, N10592, N3604, N3802, N5400);
not NOT1 (N10614, N10609);
not NOT1 (N10615, N10578);
nor NOR2 (N10616, N10607, N9554);
xor XOR2 (N10617, N10604, N8454);
nand NAND3 (N10618, N10606, N9033, N7350);
nor NOR2 (N10619, N10617, N2297);
not NOT1 (N10620, N10619);
and AND4 (N10621, N10612, N5264, N4063, N460);
xor XOR2 (N10622, N10613, N6963);
nand NAND3 (N10623, N10618, N9381, N2663);
xor XOR2 (N10624, N10591, N883);
nor NOR2 (N10625, N10616, N4046);
xor XOR2 (N10626, N10624, N10041);
xor XOR2 (N10627, N10614, N335);
nand NAND4 (N10628, N10599, N4259, N5721, N4768);
buf BUF1 (N10629, N10621);
nand NAND4 (N10630, N10628, N3952, N7694, N549);
xor XOR2 (N10631, N10611, N1304);
nand NAND3 (N10632, N10615, N8968, N7088);
nand NAND2 (N10633, N10626, N320);
nor NOR3 (N10634, N10633, N9869, N7378);
buf BUF1 (N10635, N10631);
xor XOR2 (N10636, N10623, N7669);
nor NOR2 (N10637, N10622, N2015);
buf BUF1 (N10638, N10634);
xor XOR2 (N10639, N10630, N4470);
or OR3 (N10640, N10637, N2141, N886);
buf BUF1 (N10641, N10627);
not NOT1 (N10642, N10632);
xor XOR2 (N10643, N10638, N4453);
not NOT1 (N10644, N10639);
nand NAND3 (N10645, N10644, N1989, N2541);
nor NOR4 (N10646, N10645, N1557, N478, N1660);
buf BUF1 (N10647, N10629);
nor NOR2 (N10648, N10636, N10091);
or OR3 (N10649, N10642, N3572, N2742);
and AND4 (N10650, N10647, N1153, N8787, N6607);
xor XOR2 (N10651, N10620, N4986);
not NOT1 (N10652, N10651);
nor NOR4 (N10653, N10649, N5517, N3811, N5629);
buf BUF1 (N10654, N10643);
xor XOR2 (N10655, N10653, N9907);
nor NOR4 (N10656, N10652, N9381, N7431, N7126);
not NOT1 (N10657, N10641);
not NOT1 (N10658, N10657);
or OR2 (N10659, N10646, N7511);
buf BUF1 (N10660, N10654);
or OR4 (N10661, N10625, N5592, N5779, N2328);
xor XOR2 (N10662, N10659, N819);
or OR4 (N10663, N10662, N723, N2393, N684);
not NOT1 (N10664, N10655);
nand NAND4 (N10665, N10640, N8353, N9979, N7371);
xor XOR2 (N10666, N10648, N91);
nor NOR4 (N10667, N10650, N9151, N1191, N6889);
and AND3 (N10668, N10667, N2539, N2510);
xor XOR2 (N10669, N10635, N654);
or OR3 (N10670, N10663, N3366, N8342);
or OR2 (N10671, N10661, N7496);
not NOT1 (N10672, N10664);
and AND4 (N10673, N10656, N5603, N7000, N6270);
and AND2 (N10674, N10669, N8639);
nor NOR4 (N10675, N10672, N690, N5056, N6482);
not NOT1 (N10676, N10668);
nand NAND2 (N10677, N10660, N10424);
and AND4 (N10678, N10677, N8150, N9523, N4050);
buf BUF1 (N10679, N10671);
nor NOR3 (N10680, N10666, N7500, N3857);
buf BUF1 (N10681, N10670);
not NOT1 (N10682, N10681);
not NOT1 (N10683, N10682);
or OR2 (N10684, N10676, N1347);
nand NAND2 (N10685, N10680, N6743);
or OR3 (N10686, N10678, N8359, N1107);
not NOT1 (N10687, N10674);
nor NOR4 (N10688, N10686, N8087, N5657, N10501);
nand NAND2 (N10689, N10688, N9683);
not NOT1 (N10690, N10679);
or OR2 (N10691, N10658, N810);
nand NAND2 (N10692, N10687, N10388);
or OR3 (N10693, N10685, N2190, N1891);
xor XOR2 (N10694, N10691, N8294);
and AND4 (N10695, N10690, N3964, N5667, N578);
nand NAND3 (N10696, N10695, N24, N4720);
xor XOR2 (N10697, N10673, N10217);
nand NAND2 (N10698, N10692, N696);
buf BUF1 (N10699, N10684);
or OR2 (N10700, N10694, N443);
not NOT1 (N10701, N10665);
xor XOR2 (N10702, N10701, N9898);
nor NOR4 (N10703, N10700, N10287, N1608, N9752);
or OR2 (N10704, N10683, N6033);
or OR4 (N10705, N10702, N8664, N4216, N4189);
nand NAND3 (N10706, N10705, N8154, N4011);
nand NAND2 (N10707, N10704, N7041);
and AND3 (N10708, N10706, N10648, N7234);
and AND4 (N10709, N10693, N5617, N7408, N2973);
or OR2 (N10710, N10709, N805);
xor XOR2 (N10711, N10697, N5231);
xor XOR2 (N10712, N10703, N8097);
and AND2 (N10713, N10689, N1011);
nand NAND3 (N10714, N10698, N3155, N8879);
buf BUF1 (N10715, N10713);
and AND2 (N10716, N10715, N461);
buf BUF1 (N10717, N10716);
and AND3 (N10718, N10675, N7637, N5654);
nand NAND3 (N10719, N10711, N234, N6411);
buf BUF1 (N10720, N10714);
or OR2 (N10721, N10712, N1359);
nand NAND4 (N10722, N10718, N4128, N5997, N1283);
xor XOR2 (N10723, N10722, N9662);
or OR4 (N10724, N10721, N7210, N5468, N9824);
buf BUF1 (N10725, N10723);
not NOT1 (N10726, N10707);
xor XOR2 (N10727, N10710, N4092);
or OR3 (N10728, N10699, N51, N840);
nor NOR3 (N10729, N10724, N6592, N9900);
and AND3 (N10730, N10725, N1528, N691);
buf BUF1 (N10731, N10727);
xor XOR2 (N10732, N10728, N848);
nand NAND4 (N10733, N10720, N6343, N6712, N9656);
not NOT1 (N10734, N10717);
buf BUF1 (N10735, N10708);
or OR3 (N10736, N10731, N8643, N7863);
not NOT1 (N10737, N10726);
nand NAND3 (N10738, N10696, N5839, N10525);
nor NOR2 (N10739, N10719, N610);
and AND3 (N10740, N10730, N147, N3934);
nor NOR4 (N10741, N10734, N3158, N2771, N157);
or OR4 (N10742, N10729, N9987, N339, N9987);
or OR3 (N10743, N10740, N6220, N7944);
xor XOR2 (N10744, N10741, N2782);
not NOT1 (N10745, N10743);
xor XOR2 (N10746, N10737, N9330);
nand NAND3 (N10747, N10745, N6112, N5926);
xor XOR2 (N10748, N10738, N10743);
nand NAND4 (N10749, N10733, N1606, N8432, N8146);
or OR2 (N10750, N10749, N9729);
xor XOR2 (N10751, N10744, N2960);
nor NOR4 (N10752, N10750, N10341, N8851, N2075);
or OR3 (N10753, N10752, N2377, N7136);
nand NAND2 (N10754, N10742, N1301);
buf BUF1 (N10755, N10735);
buf BUF1 (N10756, N10753);
buf BUF1 (N10757, N10754);
and AND3 (N10758, N10736, N2795, N10561);
and AND2 (N10759, N10755, N3186);
xor XOR2 (N10760, N10758, N10251);
xor XOR2 (N10761, N10748, N9878);
not NOT1 (N10762, N10757);
nand NAND4 (N10763, N10751, N7355, N7778, N2568);
xor XOR2 (N10764, N10746, N790);
and AND4 (N10765, N10747, N8229, N1991, N6703);
nand NAND2 (N10766, N10756, N5387);
or OR4 (N10767, N10766, N1334, N8903, N7438);
xor XOR2 (N10768, N10732, N6130);
nand NAND2 (N10769, N10768, N2542);
buf BUF1 (N10770, N10759);
nand NAND4 (N10771, N10763, N4662, N1897, N6110);
xor XOR2 (N10772, N10767, N2571);
nor NOR2 (N10773, N10772, N4050);
or OR3 (N10774, N10770, N9420, N4557);
or OR4 (N10775, N10765, N1559, N278, N4884);
and AND3 (N10776, N10760, N9028, N2687);
nor NOR3 (N10777, N10739, N4403, N6447);
nand NAND4 (N10778, N10774, N323, N9192, N5217);
not NOT1 (N10779, N10762);
not NOT1 (N10780, N10761);
nand NAND4 (N10781, N10778, N7687, N657, N3915);
xor XOR2 (N10782, N10781, N1129);
xor XOR2 (N10783, N10776, N4383);
nor NOR4 (N10784, N10769, N9749, N6940, N9510);
and AND4 (N10785, N10782, N4013, N5910, N5177);
buf BUF1 (N10786, N10775);
nand NAND4 (N10787, N10783, N2425, N1421, N4285);
not NOT1 (N10788, N10764);
or OR2 (N10789, N10771, N9350);
nor NOR4 (N10790, N10784, N10504, N1951, N6086);
xor XOR2 (N10791, N10788, N2917);
nand NAND4 (N10792, N10785, N5903, N7069, N3526);
not NOT1 (N10793, N10790);
not NOT1 (N10794, N10777);
nand NAND2 (N10795, N10780, N10709);
not NOT1 (N10796, N10789);
nor NOR3 (N10797, N10794, N10207, N3815);
buf BUF1 (N10798, N10787);
xor XOR2 (N10799, N10795, N2407);
nor NOR4 (N10800, N10796, N4490, N10198, N2746);
xor XOR2 (N10801, N10800, N6803);
buf BUF1 (N10802, N10799);
xor XOR2 (N10803, N10802, N6731);
or OR3 (N10804, N10786, N9794, N6651);
nand NAND3 (N10805, N10797, N5795, N9049);
buf BUF1 (N10806, N10801);
and AND2 (N10807, N10804, N3996);
or OR2 (N10808, N10805, N6330);
buf BUF1 (N10809, N10791);
not NOT1 (N10810, N10808);
xor XOR2 (N10811, N10810, N6194);
and AND2 (N10812, N10779, N5036);
buf BUF1 (N10813, N10792);
not NOT1 (N10814, N10809);
or OR4 (N10815, N10773, N566, N866, N8937);
xor XOR2 (N10816, N10803, N1249);
nor NOR2 (N10817, N10793, N915);
nand NAND2 (N10818, N10813, N5461);
xor XOR2 (N10819, N10815, N3951);
not NOT1 (N10820, N10814);
not NOT1 (N10821, N10798);
not NOT1 (N10822, N10806);
xor XOR2 (N10823, N10820, N8381);
and AND4 (N10824, N10817, N9036, N9824, N2743);
not NOT1 (N10825, N10824);
buf BUF1 (N10826, N10821);
xor XOR2 (N10827, N10819, N7585);
nor NOR4 (N10828, N10827, N7381, N8898, N5424);
and AND4 (N10829, N10818, N4952, N1347, N505);
xor XOR2 (N10830, N10811, N4152);
nor NOR3 (N10831, N10830, N1625, N2320);
or OR3 (N10832, N10829, N138, N2270);
or OR2 (N10833, N10812, N993);
xor XOR2 (N10834, N10825, N4904);
and AND2 (N10835, N10832, N5845);
buf BUF1 (N10836, N10823);
or OR4 (N10837, N10835, N4216, N2697, N228);
or OR4 (N10838, N10828, N1925, N8941, N8632);
buf BUF1 (N10839, N10833);
xor XOR2 (N10840, N10834, N5832);
not NOT1 (N10841, N10831);
and AND4 (N10842, N10840, N10032, N10631, N7590);
nor NOR3 (N10843, N10816, N10304, N4043);
xor XOR2 (N10844, N10807, N4124);
and AND2 (N10845, N10842, N3028);
nor NOR4 (N10846, N10826, N8880, N3378, N5354);
not NOT1 (N10847, N10844);
or OR3 (N10848, N10846, N10025, N1916);
buf BUF1 (N10849, N10847);
buf BUF1 (N10850, N10822);
not NOT1 (N10851, N10837);
or OR2 (N10852, N10850, N1774);
nor NOR2 (N10853, N10849, N10172);
nand NAND4 (N10854, N10843, N2743, N2268, N1337);
xor XOR2 (N10855, N10841, N5266);
nand NAND4 (N10856, N10848, N9206, N2337, N1320);
not NOT1 (N10857, N10851);
or OR4 (N10858, N10836, N3662, N8681, N7782);
buf BUF1 (N10859, N10858);
buf BUF1 (N10860, N10845);
and AND3 (N10861, N10854, N10571, N1788);
nand NAND3 (N10862, N10857, N9554, N4341);
nand NAND4 (N10863, N10859, N2169, N275, N10135);
nor NOR4 (N10864, N10861, N2905, N9399, N4300);
and AND4 (N10865, N10860, N7898, N8954, N261);
or OR2 (N10866, N10863, N10144);
and AND4 (N10867, N10866, N5067, N8544, N1842);
xor XOR2 (N10868, N10852, N10739);
or OR4 (N10869, N10868, N4740, N7689, N1392);
or OR4 (N10870, N10867, N3457, N10497, N7763);
or OR3 (N10871, N10865, N5420, N4196);
or OR4 (N10872, N10862, N3832, N9628, N2958);
not NOT1 (N10873, N10856);
nand NAND2 (N10874, N10855, N5819);
buf BUF1 (N10875, N10874);
or OR4 (N10876, N10864, N6540, N553, N1566);
nand NAND3 (N10877, N10838, N5913, N1795);
nor NOR3 (N10878, N10853, N8019, N9685);
not NOT1 (N10879, N10839);
nor NOR3 (N10880, N10871, N8559, N3683);
and AND2 (N10881, N10872, N10389);
nor NOR2 (N10882, N10876, N3520);
buf BUF1 (N10883, N10879);
or OR4 (N10884, N10875, N5342, N7448, N3684);
or OR3 (N10885, N10882, N3158, N1468);
buf BUF1 (N10886, N10885);
xor XOR2 (N10887, N10878, N10347);
or OR2 (N10888, N10873, N1994);
xor XOR2 (N10889, N10881, N6798);
or OR3 (N10890, N10880, N7391, N7157);
xor XOR2 (N10891, N10883, N4093);
and AND3 (N10892, N10884, N8298, N9845);
nand NAND3 (N10893, N10890, N10006, N1109);
buf BUF1 (N10894, N10892);
not NOT1 (N10895, N10894);
not NOT1 (N10896, N10870);
not NOT1 (N10897, N10877);
not NOT1 (N10898, N10886);
xor XOR2 (N10899, N10897, N1957);
nand NAND2 (N10900, N10889, N3149);
nand NAND2 (N10901, N10888, N4855);
or OR3 (N10902, N10891, N2998, N9905);
or OR2 (N10903, N10899, N8898);
nand NAND4 (N10904, N10895, N10147, N5988, N6896);
nand NAND4 (N10905, N10898, N7475, N8811, N1239);
buf BUF1 (N10906, N10869);
or OR4 (N10907, N10887, N6329, N8355, N1387);
not NOT1 (N10908, N10903);
nor NOR4 (N10909, N10900, N8439, N3641, N2747);
xor XOR2 (N10910, N10909, N8391);
xor XOR2 (N10911, N10906, N2152);
and AND3 (N10912, N10908, N8938, N8897);
buf BUF1 (N10913, N10910);
nor NOR4 (N10914, N10913, N5167, N728, N9198);
nor NOR3 (N10915, N10902, N2129, N10288);
xor XOR2 (N10916, N10914, N3636);
nor NOR2 (N10917, N10905, N8559);
buf BUF1 (N10918, N10917);
xor XOR2 (N10919, N10904, N5578);
buf BUF1 (N10920, N10915);
xor XOR2 (N10921, N10919, N1259);
xor XOR2 (N10922, N10896, N913);
nand NAND3 (N10923, N10916, N2026, N1472);
or OR3 (N10924, N10907, N9223, N1368);
and AND2 (N10925, N10920, N1804);
xor XOR2 (N10926, N10912, N224);
or OR3 (N10927, N10923, N10285, N8557);
not NOT1 (N10928, N10918);
nand NAND4 (N10929, N10926, N3834, N10295, N1037);
buf BUF1 (N10930, N10924);
xor XOR2 (N10931, N10922, N3000);
not NOT1 (N10932, N10927);
buf BUF1 (N10933, N10901);
xor XOR2 (N10934, N10931, N1417);
nand NAND3 (N10935, N10911, N5433, N8006);
not NOT1 (N10936, N10932);
and AND4 (N10937, N10928, N31, N5322, N2586);
nor NOR2 (N10938, N10929, N8477);
or OR3 (N10939, N10933, N7980, N1851);
xor XOR2 (N10940, N10937, N2427);
xor XOR2 (N10941, N10925, N8238);
nor NOR4 (N10942, N10939, N3087, N9415, N8518);
and AND3 (N10943, N10941, N5254, N7781);
nand NAND4 (N10944, N10942, N8919, N10227, N4828);
and AND3 (N10945, N10936, N2783, N4378);
nor NOR4 (N10946, N10944, N7283, N1229, N8613);
not NOT1 (N10947, N10945);
nor NOR3 (N10948, N10893, N2016, N9866);
nor NOR4 (N10949, N10935, N3552, N1063, N5335);
nand NAND4 (N10950, N10948, N4578, N802, N1838);
not NOT1 (N10951, N10938);
not NOT1 (N10952, N10950);
nor NOR3 (N10953, N10940, N5661, N3863);
buf BUF1 (N10954, N10930);
buf BUF1 (N10955, N10953);
not NOT1 (N10956, N10954);
nand NAND2 (N10957, N10943, N2873);
or OR3 (N10958, N10921, N4340, N5070);
nand NAND3 (N10959, N10952, N8986, N6874);
xor XOR2 (N10960, N10949, N7433);
buf BUF1 (N10961, N10958);
nand NAND3 (N10962, N10934, N5721, N6754);
or OR2 (N10963, N10959, N10096);
nor NOR4 (N10964, N10955, N5875, N3817, N5346);
buf BUF1 (N10965, N10961);
nand NAND3 (N10966, N10956, N5107, N2071);
not NOT1 (N10967, N10963);
not NOT1 (N10968, N10962);
and AND3 (N10969, N10968, N7799, N1450);
nand NAND4 (N10970, N10964, N1866, N2411, N2727);
nor NOR3 (N10971, N10969, N3502, N4464);
nand NAND2 (N10972, N10970, N1938);
xor XOR2 (N10973, N10966, N10110);
xor XOR2 (N10974, N10960, N7808);
not NOT1 (N10975, N10971);
xor XOR2 (N10976, N10974, N6468);
nor NOR2 (N10977, N10975, N2088);
buf BUF1 (N10978, N10965);
nor NOR2 (N10979, N10972, N6355);
or OR4 (N10980, N10976, N6129, N4519, N1630);
and AND4 (N10981, N10957, N2770, N336, N7288);
nand NAND2 (N10982, N10977, N10975);
nor NOR2 (N10983, N10980, N2008);
or OR2 (N10984, N10967, N7990);
or OR3 (N10985, N10984, N7999, N662);
nand NAND2 (N10986, N10982, N6257);
xor XOR2 (N10987, N10978, N4462);
buf BUF1 (N10988, N10979);
and AND4 (N10989, N10981, N1511, N1778, N9393);
nand NAND3 (N10990, N10951, N1185, N8194);
and AND2 (N10991, N10973, N914);
buf BUF1 (N10992, N10986);
buf BUF1 (N10993, N10990);
or OR3 (N10994, N10946, N7827, N1341);
or OR2 (N10995, N10985, N7290);
not NOT1 (N10996, N10987);
not NOT1 (N10997, N10989);
xor XOR2 (N10998, N10992, N8381);
or OR4 (N10999, N10997, N3247, N2531, N7716);
and AND4 (N11000, N10988, N8695, N7987, N6190);
or OR3 (N11001, N10995, N536, N2836);
not NOT1 (N11002, N10998);
and AND3 (N11003, N10994, N5778, N9699);
nand NAND2 (N11004, N11003, N3710);
or OR3 (N11005, N11004, N10187, N6463);
nand NAND3 (N11006, N10999, N103, N35);
nor NOR4 (N11007, N11006, N7058, N10767, N1347);
buf BUF1 (N11008, N10983);
or OR2 (N11009, N10993, N1038);
or OR3 (N11010, N11001, N7703, N10228);
xor XOR2 (N11011, N11000, N2039);
xor XOR2 (N11012, N11009, N8432);
buf BUF1 (N11013, N10991);
nand NAND3 (N11014, N10996, N9739, N5125);
not NOT1 (N11015, N11012);
or OR3 (N11016, N11005, N260, N4173);
nand NAND4 (N11017, N11015, N4490, N3660, N1298);
or OR2 (N11018, N11010, N6219);
nor NOR2 (N11019, N11017, N2521);
not NOT1 (N11020, N11013);
buf BUF1 (N11021, N11018);
buf BUF1 (N11022, N11020);
or OR3 (N11023, N11007, N7053, N9262);
not NOT1 (N11024, N11019);
xor XOR2 (N11025, N11023, N7190);
nand NAND2 (N11026, N10947, N8585);
nor NOR2 (N11027, N11026, N5131);
buf BUF1 (N11028, N11008);
not NOT1 (N11029, N11028);
xor XOR2 (N11030, N11014, N2287);
buf BUF1 (N11031, N11022);
not NOT1 (N11032, N11030);
or OR2 (N11033, N11032, N7027);
nand NAND4 (N11034, N11024, N7258, N2120, N5871);
not NOT1 (N11035, N11031);
nand NAND4 (N11036, N11034, N6035, N9672, N3037);
buf BUF1 (N11037, N11033);
or OR3 (N11038, N11011, N7777, N3681);
nand NAND4 (N11039, N11037, N4791, N9643, N3378);
xor XOR2 (N11040, N11016, N3173);
not NOT1 (N11041, N11027);
xor XOR2 (N11042, N11021, N231);
or OR2 (N11043, N11039, N6349);
not NOT1 (N11044, N11025);
xor XOR2 (N11045, N11042, N9505);
nor NOR3 (N11046, N11045, N8287, N2942);
not NOT1 (N11047, N11046);
or OR3 (N11048, N11040, N7678, N4685);
nand NAND4 (N11049, N11048, N7570, N868, N3794);
and AND3 (N11050, N11002, N10332, N8579);
nor NOR4 (N11051, N11041, N1995, N7503, N4308);
not NOT1 (N11052, N11049);
and AND2 (N11053, N11043, N3781);
buf BUF1 (N11054, N11051);
nor NOR3 (N11055, N11044, N9596, N4579);
xor XOR2 (N11056, N11054, N8933);
or OR2 (N11057, N11029, N4276);
nand NAND3 (N11058, N11052, N1140, N4181);
buf BUF1 (N11059, N11038);
xor XOR2 (N11060, N11055, N9774);
not NOT1 (N11061, N11057);
and AND2 (N11062, N11061, N6099);
and AND4 (N11063, N11056, N5702, N1909, N1372);
xor XOR2 (N11064, N11063, N10592);
nand NAND2 (N11065, N11060, N6236);
or OR3 (N11066, N11065, N4378, N10487);
or OR2 (N11067, N11062, N10240);
nand NAND2 (N11068, N11047, N8265);
nand NAND4 (N11069, N11067, N7264, N8216, N3863);
or OR3 (N11070, N11053, N7233, N10054);
not NOT1 (N11071, N11068);
or OR3 (N11072, N11070, N1618, N6033);
not NOT1 (N11073, N11066);
buf BUF1 (N11074, N11059);
nor NOR3 (N11075, N11050, N305, N5666);
and AND2 (N11076, N11071, N9939);
and AND2 (N11077, N11072, N7495);
nand NAND4 (N11078, N11074, N6113, N6852, N6817);
nand NAND2 (N11079, N11058, N1906);
and AND3 (N11080, N11035, N5862, N2335);
buf BUF1 (N11081, N11077);
buf BUF1 (N11082, N11079);
buf BUF1 (N11083, N11075);
or OR3 (N11084, N11081, N1671, N2953);
buf BUF1 (N11085, N11076);
not NOT1 (N11086, N11078);
buf BUF1 (N11087, N11082);
nor NOR4 (N11088, N11069, N7632, N9588, N2207);
xor XOR2 (N11089, N11073, N4857);
xor XOR2 (N11090, N11036, N5128);
xor XOR2 (N11091, N11083, N3832);
not NOT1 (N11092, N11086);
not NOT1 (N11093, N11089);
xor XOR2 (N11094, N11090, N7943);
xor XOR2 (N11095, N11084, N10702);
not NOT1 (N11096, N11093);
buf BUF1 (N11097, N11096);
nand NAND4 (N11098, N11088, N5629, N946, N7795);
not NOT1 (N11099, N11085);
nor NOR4 (N11100, N11080, N3689, N170, N1317);
nor NOR4 (N11101, N11097, N2346, N671, N2756);
nor NOR2 (N11102, N11095, N10218);
buf BUF1 (N11103, N11100);
not NOT1 (N11104, N11099);
buf BUF1 (N11105, N11092);
nor NOR4 (N11106, N11102, N8028, N4636, N5903);
xor XOR2 (N11107, N11101, N460);
xor XOR2 (N11108, N11105, N8026);
nor NOR3 (N11109, N11108, N2546, N8812);
and AND3 (N11110, N11091, N4518, N4184);
nand NAND4 (N11111, N11103, N3111, N6844, N5292);
nor NOR3 (N11112, N11098, N7276, N4295);
nand NAND4 (N11113, N11104, N8680, N1822, N4011);
nand NAND4 (N11114, N11064, N998, N6827, N1622);
nor NOR4 (N11115, N11106, N9539, N213, N1283);
not NOT1 (N11116, N11113);
xor XOR2 (N11117, N11111, N2699);
xor XOR2 (N11118, N11107, N8889);
not NOT1 (N11119, N11116);
not NOT1 (N11120, N11087);
buf BUF1 (N11121, N11110);
not NOT1 (N11122, N11094);
or OR2 (N11123, N11112, N3381);
or OR4 (N11124, N11115, N3075, N1297, N6148);
nor NOR3 (N11125, N11122, N6465, N3748);
nand NAND2 (N11126, N11117, N5468);
or OR2 (N11127, N11124, N2410);
xor XOR2 (N11128, N11121, N8765);
or OR3 (N11129, N11114, N3780, N5451);
nand NAND3 (N11130, N11109, N1917, N1783);
not NOT1 (N11131, N11125);
not NOT1 (N11132, N11128);
nor NOR2 (N11133, N11118, N2944);
buf BUF1 (N11134, N11126);
nor NOR4 (N11135, N11133, N1925, N10083, N7003);
not NOT1 (N11136, N11131);
not NOT1 (N11137, N11136);
or OR4 (N11138, N11120, N8276, N10575, N8869);
and AND2 (N11139, N11130, N8442);
nand NAND2 (N11140, N11139, N8786);
buf BUF1 (N11141, N11137);
and AND3 (N11142, N11129, N4107, N10976);
nor NOR2 (N11143, N11142, N8422);
buf BUF1 (N11144, N11127);
nor NOR3 (N11145, N11119, N6180, N8284);
buf BUF1 (N11146, N11132);
or OR3 (N11147, N11123, N3304, N5541);
buf BUF1 (N11148, N11141);
and AND4 (N11149, N11145, N9689, N7716, N7381);
buf BUF1 (N11150, N11138);
xor XOR2 (N11151, N11147, N7021);
nor NOR4 (N11152, N11150, N5723, N8941, N6060);
buf BUF1 (N11153, N11143);
buf BUF1 (N11154, N11151);
not NOT1 (N11155, N11148);
not NOT1 (N11156, N11152);
nand NAND3 (N11157, N11146, N4461, N9885);
not NOT1 (N11158, N11157);
xor XOR2 (N11159, N11153, N828);
nand NAND4 (N11160, N11134, N3153, N7985, N4511);
or OR3 (N11161, N11155, N2207, N5234);
xor XOR2 (N11162, N11156, N3844);
buf BUF1 (N11163, N11161);
xor XOR2 (N11164, N11149, N6428);
or OR4 (N11165, N11140, N9509, N4213, N10983);
xor XOR2 (N11166, N11135, N8514);
and AND4 (N11167, N11144, N10408, N510, N10421);
buf BUF1 (N11168, N11167);
nor NOR3 (N11169, N11159, N10447, N8373);
xor XOR2 (N11170, N11166, N7258);
not NOT1 (N11171, N11158);
xor XOR2 (N11172, N11170, N6216);
nor NOR3 (N11173, N11171, N10968, N1157);
nand NAND3 (N11174, N11160, N2904, N625);
not NOT1 (N11175, N11162);
buf BUF1 (N11176, N11173);
or OR2 (N11177, N11168, N8164);
nor NOR3 (N11178, N11154, N9559, N6642);
or OR3 (N11179, N11177, N2074, N9097);
or OR2 (N11180, N11172, N5301);
xor XOR2 (N11181, N11165, N10461);
xor XOR2 (N11182, N11174, N5191);
not NOT1 (N11183, N11176);
buf BUF1 (N11184, N11182);
and AND4 (N11185, N11179, N4054, N4680, N9012);
nand NAND3 (N11186, N11185, N10531, N1689);
nand NAND3 (N11187, N11178, N1636, N649);
nor NOR2 (N11188, N11180, N213);
and AND4 (N11189, N11186, N7766, N6329, N7373);
xor XOR2 (N11190, N11188, N1363);
or OR4 (N11191, N11163, N9914, N6173, N2239);
nand NAND3 (N11192, N11169, N3098, N369);
and AND4 (N11193, N11187, N7104, N3755, N9380);
or OR3 (N11194, N11175, N2448, N6016);
and AND4 (N11195, N11194, N11059, N4483, N3825);
or OR4 (N11196, N11164, N8117, N5481, N6592);
and AND3 (N11197, N11183, N7910, N6807);
nor NOR4 (N11198, N11191, N3124, N9898, N121);
buf BUF1 (N11199, N11189);
buf BUF1 (N11200, N11197);
not NOT1 (N11201, N11195);
nand NAND3 (N11202, N11192, N3696, N7488);
nor NOR3 (N11203, N11201, N10965, N8619);
not NOT1 (N11204, N11184);
not NOT1 (N11205, N11200);
not NOT1 (N11206, N11196);
and AND3 (N11207, N11202, N9723, N9139);
buf BUF1 (N11208, N11203);
buf BUF1 (N11209, N11207);
or OR3 (N11210, N11199, N5190, N10732);
nor NOR2 (N11211, N11208, N673);
xor XOR2 (N11212, N11204, N4935);
xor XOR2 (N11213, N11193, N4137);
nor NOR3 (N11214, N11213, N7774, N8934);
buf BUF1 (N11215, N11205);
nand NAND3 (N11216, N11210, N5592, N862);
and AND3 (N11217, N11206, N2148, N4691);
buf BUF1 (N11218, N11209);
xor XOR2 (N11219, N11212, N5497);
buf BUF1 (N11220, N11181);
nor NOR2 (N11221, N11218, N1917);
not NOT1 (N11222, N11215);
nand NAND4 (N11223, N11217, N10956, N5573, N6445);
xor XOR2 (N11224, N11221, N267);
and AND4 (N11225, N11223, N4837, N2377, N5215);
nor NOR3 (N11226, N11198, N3418, N1721);
nand NAND4 (N11227, N11190, N11191, N3926, N475);
buf BUF1 (N11228, N11211);
not NOT1 (N11229, N11225);
xor XOR2 (N11230, N11216, N2213);
nand NAND2 (N11231, N11227, N5379);
nand NAND2 (N11232, N11228, N10655);
nor NOR2 (N11233, N11232, N8563);
and AND3 (N11234, N11219, N6927, N5239);
nor NOR2 (N11235, N11230, N1786);
and AND2 (N11236, N11214, N1043);
or OR4 (N11237, N11234, N2703, N3520, N1753);
nor NOR2 (N11238, N11224, N8169);
nand NAND2 (N11239, N11220, N1680);
xor XOR2 (N11240, N11229, N7006);
or OR3 (N11241, N11240, N6693, N2860);
xor XOR2 (N11242, N11231, N2290);
xor XOR2 (N11243, N11233, N4800);
not NOT1 (N11244, N11222);
nor NOR2 (N11245, N11237, N8450);
not NOT1 (N11246, N11238);
nand NAND2 (N11247, N11244, N54);
or OR2 (N11248, N11239, N8195);
buf BUF1 (N11249, N11235);
or OR3 (N11250, N11226, N3069, N2571);
not NOT1 (N11251, N11249);
nor NOR4 (N11252, N11241, N5761, N6218, N3114);
xor XOR2 (N11253, N11245, N3212);
not NOT1 (N11254, N11236);
buf BUF1 (N11255, N11247);
not NOT1 (N11256, N11255);
nor NOR2 (N11257, N11250, N3846);
not NOT1 (N11258, N11243);
not NOT1 (N11259, N11258);
nand NAND2 (N11260, N11248, N9327);
nand NAND2 (N11261, N11251, N9167);
not NOT1 (N11262, N11253);
or OR2 (N11263, N11262, N3531);
or OR2 (N11264, N11256, N630);
and AND2 (N11265, N11242, N1924);
buf BUF1 (N11266, N11263);
xor XOR2 (N11267, N11266, N3073);
nor NOR2 (N11268, N11259, N4215);
not NOT1 (N11269, N11246);
and AND3 (N11270, N11260, N4511, N8916);
or OR2 (N11271, N11267, N181);
not NOT1 (N11272, N11264);
buf BUF1 (N11273, N11268);
and AND4 (N11274, N11271, N2805, N11150, N4224);
not NOT1 (N11275, N11270);
not NOT1 (N11276, N11269);
not NOT1 (N11277, N11273);
and AND3 (N11278, N11261, N1602, N9526);
not NOT1 (N11279, N11257);
and AND3 (N11280, N11265, N746, N5755);
nor NOR2 (N11281, N11274, N2831);
nand NAND3 (N11282, N11272, N5877, N1033);
xor XOR2 (N11283, N11277, N6357);
not NOT1 (N11284, N11282);
nor NOR4 (N11285, N11254, N5154, N10729, N8027);
not NOT1 (N11286, N11284);
or OR3 (N11287, N11286, N1862, N1827);
nand NAND2 (N11288, N11275, N3259);
buf BUF1 (N11289, N11279);
xor XOR2 (N11290, N11276, N7441);
nand NAND4 (N11291, N11290, N10289, N2524, N4220);
or OR4 (N11292, N11285, N3119, N5328, N9689);
nand NAND4 (N11293, N11287, N3078, N9572, N3730);
nand NAND4 (N11294, N11280, N1835, N385, N5154);
or OR4 (N11295, N11252, N6822, N7736, N6614);
not NOT1 (N11296, N11289);
xor XOR2 (N11297, N11283, N2437);
xor XOR2 (N11298, N11293, N10297);
and AND3 (N11299, N11288, N3826, N526);
buf BUF1 (N11300, N11297);
or OR2 (N11301, N11278, N3871);
xor XOR2 (N11302, N11294, N10847);
or OR4 (N11303, N11296, N7215, N6468, N9321);
xor XOR2 (N11304, N11298, N920);
nand NAND3 (N11305, N11291, N25, N2357);
xor XOR2 (N11306, N11295, N6058);
not NOT1 (N11307, N11299);
nand NAND4 (N11308, N11292, N4587, N2739, N4259);
nand NAND4 (N11309, N11303, N4607, N6273, N6437);
xor XOR2 (N11310, N11305, N1252);
or OR4 (N11311, N11304, N6369, N652, N6856);
and AND2 (N11312, N11306, N2821);
and AND3 (N11313, N11308, N7292, N3265);
buf BUF1 (N11314, N11309);
or OR2 (N11315, N11310, N10171);
or OR3 (N11316, N11315, N7257, N7464);
and AND2 (N11317, N11281, N7681);
nor NOR3 (N11318, N11301, N8210, N9864);
xor XOR2 (N11319, N11317, N7354);
and AND3 (N11320, N11313, N3264, N3829);
buf BUF1 (N11321, N11300);
buf BUF1 (N11322, N11311);
not NOT1 (N11323, N11314);
nand NAND4 (N11324, N11320, N7177, N9678, N2319);
nand NAND2 (N11325, N11322, N5239);
or OR3 (N11326, N11325, N1397, N9487);
not NOT1 (N11327, N11321);
or OR3 (N11328, N11312, N8408, N4609);
and AND2 (N11329, N11307, N5764);
nor NOR2 (N11330, N11323, N842);
not NOT1 (N11331, N11329);
or OR2 (N11332, N11326, N10801);
buf BUF1 (N11333, N11330);
nand NAND2 (N11334, N11318, N8689);
or OR2 (N11335, N11327, N6577);
xor XOR2 (N11336, N11316, N10689);
and AND4 (N11337, N11336, N4195, N2843, N6461);
nand NAND4 (N11338, N11328, N10226, N4618, N9120);
nor NOR2 (N11339, N11302, N4467);
and AND4 (N11340, N11333, N2225, N6369, N10);
nor NOR4 (N11341, N11338, N5343, N5166, N10477);
not NOT1 (N11342, N11337);
buf BUF1 (N11343, N11324);
and AND4 (N11344, N11341, N5322, N7689, N1178);
not NOT1 (N11345, N11339);
or OR2 (N11346, N11343, N7138);
xor XOR2 (N11347, N11334, N11251);
or OR4 (N11348, N11332, N1720, N2940, N11270);
buf BUF1 (N11349, N11342);
not NOT1 (N11350, N11348);
or OR2 (N11351, N11349, N7782);
and AND4 (N11352, N11319, N4057, N9863, N8811);
not NOT1 (N11353, N11352);
and AND4 (N11354, N11347, N689, N10013, N3420);
buf BUF1 (N11355, N11351);
buf BUF1 (N11356, N11355);
not NOT1 (N11357, N11345);
xor XOR2 (N11358, N11340, N6502);
buf BUF1 (N11359, N11350);
nor NOR2 (N11360, N11335, N8495);
or OR4 (N11361, N11360, N9891, N9247, N11032);
not NOT1 (N11362, N11359);
xor XOR2 (N11363, N11331, N1878);
not NOT1 (N11364, N11363);
not NOT1 (N11365, N11353);
or OR2 (N11366, N11362, N2544);
not NOT1 (N11367, N11358);
buf BUF1 (N11368, N11356);
buf BUF1 (N11369, N11357);
xor XOR2 (N11370, N11369, N2908);
and AND2 (N11371, N11370, N222);
nand NAND3 (N11372, N11368, N6012, N3811);
or OR3 (N11373, N11344, N6007, N6260);
nor NOR2 (N11374, N11354, N10943);
and AND3 (N11375, N11373, N1153, N4126);
not NOT1 (N11376, N11364);
nor NOR3 (N11377, N11371, N1794, N6799);
buf BUF1 (N11378, N11361);
not NOT1 (N11379, N11367);
buf BUF1 (N11380, N11379);
or OR2 (N11381, N11376, N6320);
not NOT1 (N11382, N11374);
nand NAND2 (N11383, N11366, N3622);
or OR3 (N11384, N11365, N2470, N8044);
nor NOR3 (N11385, N11346, N7465, N7018);
xor XOR2 (N11386, N11372, N1247);
nand NAND4 (N11387, N11384, N2466, N1362, N10841);
and AND4 (N11388, N11381, N3873, N9488, N10532);
nor NOR4 (N11389, N11383, N7378, N5727, N4094);
buf BUF1 (N11390, N11375);
xor XOR2 (N11391, N11378, N4961);
xor XOR2 (N11392, N11387, N8469);
xor XOR2 (N11393, N11377, N1821);
or OR3 (N11394, N11390, N7345, N2766);
not NOT1 (N11395, N11394);
or OR4 (N11396, N11385, N1947, N3496, N4077);
buf BUF1 (N11397, N11388);
buf BUF1 (N11398, N11382);
and AND4 (N11399, N11391, N1439, N802, N10777);
nor NOR3 (N11400, N11398, N10885, N3609);
nand NAND4 (N11401, N11395, N6119, N5395, N10050);
nor NOR4 (N11402, N11386, N6079, N1068, N4166);
nand NAND4 (N11403, N11392, N10468, N156, N7654);
or OR4 (N11404, N11400, N4534, N7315, N10619);
buf BUF1 (N11405, N11396);
nor NOR3 (N11406, N11401, N8676, N10987);
not NOT1 (N11407, N11380);
and AND4 (N11408, N11407, N11160, N6596, N8658);
nand NAND4 (N11409, N11399, N1783, N7570, N1708);
and AND2 (N11410, N11409, N9041);
and AND4 (N11411, N11408, N3473, N5631, N4967);
nor NOR3 (N11412, N11389, N1393, N10713);
not NOT1 (N11413, N11397);
not NOT1 (N11414, N11393);
buf BUF1 (N11415, N11412);
not NOT1 (N11416, N11406);
or OR3 (N11417, N11405, N1059, N10117);
not NOT1 (N11418, N11417);
nand NAND2 (N11419, N11418, N7993);
xor XOR2 (N11420, N11416, N7609);
xor XOR2 (N11421, N11411, N3535);
and AND3 (N11422, N11413, N5307, N9911);
and AND4 (N11423, N11421, N5424, N4624, N1789);
not NOT1 (N11424, N11414);
xor XOR2 (N11425, N11419, N2960);
or OR4 (N11426, N11402, N10161, N7896, N5903);
not NOT1 (N11427, N11415);
and AND2 (N11428, N11410, N3710);
or OR3 (N11429, N11424, N4655, N8439);
xor XOR2 (N11430, N11420, N5713);
nor NOR2 (N11431, N11429, N1924);
buf BUF1 (N11432, N11426);
nor NOR3 (N11433, N11430, N3924, N4693);
nor NOR4 (N11434, N11425, N8157, N10963, N1026);
xor XOR2 (N11435, N11422, N1222);
buf BUF1 (N11436, N11403);
xor XOR2 (N11437, N11434, N115);
or OR3 (N11438, N11427, N1886, N1646);
nand NAND4 (N11439, N11435, N6989, N6489, N8949);
nand NAND4 (N11440, N11439, N10921, N3172, N6507);
xor XOR2 (N11441, N11433, N3389);
buf BUF1 (N11442, N11441);
nor NOR2 (N11443, N11431, N6408);
not NOT1 (N11444, N11440);
nor NOR3 (N11445, N11436, N8995, N11310);
and AND3 (N11446, N11442, N3151, N5137);
nand NAND3 (N11447, N11428, N7094, N7572);
nor NOR2 (N11448, N11423, N2958);
nor NOR4 (N11449, N11445, N1476, N9529, N7023);
not NOT1 (N11450, N11446);
and AND3 (N11451, N11438, N8122, N8703);
not NOT1 (N11452, N11451);
and AND2 (N11453, N11450, N1488);
nor NOR3 (N11454, N11444, N8651, N2138);
xor XOR2 (N11455, N11452, N1525);
and AND4 (N11456, N11404, N5032, N5890, N9869);
buf BUF1 (N11457, N11456);
not NOT1 (N11458, N11454);
or OR4 (N11459, N11443, N3876, N3129, N9548);
not NOT1 (N11460, N11458);
not NOT1 (N11461, N11460);
nor NOR4 (N11462, N11432, N1793, N9628, N6060);
nand NAND4 (N11463, N11461, N5721, N7072, N84);
buf BUF1 (N11464, N11437);
or OR3 (N11465, N11448, N867, N5370);
nand NAND3 (N11466, N11459, N8213, N7401);
xor XOR2 (N11467, N11455, N6960);
nand NAND2 (N11468, N11457, N4772);
not NOT1 (N11469, N11468);
buf BUF1 (N11470, N11465);
not NOT1 (N11471, N11463);
and AND4 (N11472, N11466, N2690, N5626, N6836);
nand NAND2 (N11473, N11447, N8894);
nand NAND3 (N11474, N11462, N8963, N2758);
and AND2 (N11475, N11474, N9453);
and AND3 (N11476, N11453, N1451, N9596);
not NOT1 (N11477, N11469);
nor NOR4 (N11478, N11471, N7354, N2522, N2430);
not NOT1 (N11479, N11473);
or OR3 (N11480, N11476, N2199, N11042);
nand NAND2 (N11481, N11475, N9494);
and AND2 (N11482, N11479, N7909);
xor XOR2 (N11483, N11478, N11211);
or OR4 (N11484, N11449, N5960, N2836, N10519);
nand NAND3 (N11485, N11467, N964, N2960);
or OR3 (N11486, N11481, N7675, N2317);
nor NOR3 (N11487, N11484, N8574, N5555);
or OR3 (N11488, N11485, N3330, N8428);
not NOT1 (N11489, N11486);
and AND2 (N11490, N11487, N2316);
and AND3 (N11491, N11464, N9957, N6780);
xor XOR2 (N11492, N11488, N9408);
and AND4 (N11493, N11491, N11033, N1421, N2462);
nor NOR3 (N11494, N11493, N5469, N4805);
buf BUF1 (N11495, N11489);
not NOT1 (N11496, N11480);
or OR2 (N11497, N11490, N466);
nor NOR2 (N11498, N11470, N7639);
nor NOR2 (N11499, N11498, N6511);
or OR3 (N11500, N11499, N1602, N10567);
buf BUF1 (N11501, N11495);
or OR3 (N11502, N11482, N10560, N10880);
or OR2 (N11503, N11497, N1828);
or OR3 (N11504, N11492, N1424, N4204);
and AND3 (N11505, N11496, N8908, N5333);
and AND3 (N11506, N11472, N11074, N783);
xor XOR2 (N11507, N11494, N1297);
nand NAND4 (N11508, N11477, N930, N8300, N10964);
not NOT1 (N11509, N11504);
xor XOR2 (N11510, N11501, N4811);
buf BUF1 (N11511, N11508);
nor NOR2 (N11512, N11483, N4485);
nand NAND2 (N11513, N11506, N6152);
or OR3 (N11514, N11503, N206, N3049);
or OR4 (N11515, N11514, N10682, N5497, N2387);
buf BUF1 (N11516, N11505);
buf BUF1 (N11517, N11500);
nor NOR4 (N11518, N11515, N8793, N1543, N2710);
or OR3 (N11519, N11509, N9204, N2030);
buf BUF1 (N11520, N11512);
xor XOR2 (N11521, N11511, N6088);
not NOT1 (N11522, N11510);
nor NOR2 (N11523, N11520, N10914);
nand NAND4 (N11524, N11521, N9359, N9497, N9527);
not NOT1 (N11525, N11519);
buf BUF1 (N11526, N11522);
and AND3 (N11527, N11525, N2731, N4330);
nand NAND3 (N11528, N11513, N4036, N10611);
nand NAND3 (N11529, N11516, N3926, N2759);
nor NOR2 (N11530, N11518, N7576);
not NOT1 (N11531, N11529);
buf BUF1 (N11532, N11524);
xor XOR2 (N11533, N11502, N7351);
nand NAND3 (N11534, N11523, N5827, N8429);
nor NOR2 (N11535, N11534, N6439);
xor XOR2 (N11536, N11526, N906);
and AND2 (N11537, N11527, N7108);
xor XOR2 (N11538, N11535, N9229);
xor XOR2 (N11539, N11528, N2085);
not NOT1 (N11540, N11538);
nor NOR2 (N11541, N11531, N5091);
or OR4 (N11542, N11540, N4810, N9947, N5465);
xor XOR2 (N11543, N11507, N4557);
nand NAND4 (N11544, N11537, N514, N8481, N4055);
buf BUF1 (N11545, N11530);
xor XOR2 (N11546, N11544, N5173);
xor XOR2 (N11547, N11545, N176);
not NOT1 (N11548, N11547);
or OR2 (N11549, N11533, N6368);
not NOT1 (N11550, N11541);
buf BUF1 (N11551, N11536);
nor NOR3 (N11552, N11542, N3625, N7781);
xor XOR2 (N11553, N11543, N7355);
buf BUF1 (N11554, N11548);
nor NOR2 (N11555, N11517, N11117);
buf BUF1 (N11556, N11550);
buf BUF1 (N11557, N11556);
nor NOR2 (N11558, N11554, N665);
nand NAND2 (N11559, N11558, N1507);
nor NOR2 (N11560, N11551, N7205);
buf BUF1 (N11561, N11553);
xor XOR2 (N11562, N11532, N3210);
xor XOR2 (N11563, N11549, N1011);
not NOT1 (N11564, N11562);
and AND3 (N11565, N11559, N9732, N2670);
or OR3 (N11566, N11560, N11543, N10195);
nand NAND4 (N11567, N11561, N2548, N4357, N6440);
not NOT1 (N11568, N11539);
nand NAND4 (N11569, N11568, N7662, N4511, N10742);
buf BUF1 (N11570, N11569);
nand NAND2 (N11571, N11546, N4571);
and AND2 (N11572, N11552, N6666);
buf BUF1 (N11573, N11563);
nor NOR2 (N11574, N11566, N1755);
not NOT1 (N11575, N11573);
nor NOR4 (N11576, N11571, N7638, N832, N10830);
or OR4 (N11577, N11575, N346, N8899, N10478);
xor XOR2 (N11578, N11557, N8441);
or OR4 (N11579, N11572, N2901, N4099, N10042);
xor XOR2 (N11580, N11576, N11264);
not NOT1 (N11581, N11567);
buf BUF1 (N11582, N11565);
nor NOR3 (N11583, N11574, N11265, N9824);
nand NAND2 (N11584, N11570, N1728);
or OR2 (N11585, N11581, N6887);
or OR2 (N11586, N11555, N9700);
xor XOR2 (N11587, N11582, N1856);
not NOT1 (N11588, N11577);
buf BUF1 (N11589, N11583);
xor XOR2 (N11590, N11588, N7075);
and AND4 (N11591, N11589, N3502, N9596, N8082);
nor NOR2 (N11592, N11585, N786);
xor XOR2 (N11593, N11580, N8310);
nor NOR2 (N11594, N11592, N7703);
or OR4 (N11595, N11593, N499, N6089, N11566);
and AND2 (N11596, N11595, N2339);
nor NOR3 (N11597, N11587, N3558, N9363);
nand NAND4 (N11598, N11578, N9402, N216, N6705);
nor NOR4 (N11599, N11596, N748, N9075, N6933);
nand NAND4 (N11600, N11590, N476, N5712, N7091);
not NOT1 (N11601, N11598);
buf BUF1 (N11602, N11579);
nor NOR2 (N11603, N11599, N4900);
xor XOR2 (N11604, N11584, N7352);
and AND4 (N11605, N11600, N2864, N9482, N7996);
xor XOR2 (N11606, N11604, N6228);
or OR2 (N11607, N11601, N4989);
and AND2 (N11608, N11564, N10306);
and AND3 (N11609, N11605, N10667, N8470);
xor XOR2 (N11610, N11608, N2845);
nand NAND2 (N11611, N11602, N3329);
not NOT1 (N11612, N11610);
and AND3 (N11613, N11586, N8442, N3194);
nor NOR3 (N11614, N11607, N6601, N10502);
or OR2 (N11615, N11611, N10889);
nor NOR3 (N11616, N11613, N8886, N7481);
buf BUF1 (N11617, N11616);
xor XOR2 (N11618, N11591, N2393);
not NOT1 (N11619, N11614);
xor XOR2 (N11620, N11615, N445);
xor XOR2 (N11621, N11606, N7983);
nand NAND3 (N11622, N11620, N8708, N6106);
nor NOR3 (N11623, N11612, N10938, N3843);
not NOT1 (N11624, N11619);
xor XOR2 (N11625, N11618, N9707);
xor XOR2 (N11626, N11617, N8121);
and AND3 (N11627, N11594, N2139, N7611);
buf BUF1 (N11628, N11621);
not NOT1 (N11629, N11626);
or OR3 (N11630, N11627, N11333, N2090);
buf BUF1 (N11631, N11625);
nor NOR3 (N11632, N11629, N7314, N5876);
nand NAND3 (N11633, N11632, N11252, N8548);
not NOT1 (N11634, N11609);
and AND3 (N11635, N11624, N4809, N7449);
xor XOR2 (N11636, N11630, N4050);
and AND4 (N11637, N11635, N4729, N3969, N6898);
not NOT1 (N11638, N11636);
or OR4 (N11639, N11623, N4851, N9601, N9167);
and AND4 (N11640, N11631, N2424, N6897, N2638);
buf BUF1 (N11641, N11597);
nor NOR2 (N11642, N11641, N11149);
buf BUF1 (N11643, N11640);
nand NAND2 (N11644, N11638, N938);
xor XOR2 (N11645, N11603, N1910);
not NOT1 (N11646, N11643);
or OR2 (N11647, N11645, N1308);
or OR3 (N11648, N11642, N7806, N7245);
or OR4 (N11649, N11634, N2898, N718, N6376);
xor XOR2 (N11650, N11649, N7841);
nand NAND2 (N11651, N11650, N2264);
buf BUF1 (N11652, N11639);
buf BUF1 (N11653, N11647);
nor NOR4 (N11654, N11644, N3451, N9185, N8735);
or OR3 (N11655, N11648, N1720, N5514);
xor XOR2 (N11656, N11622, N1231);
nand NAND2 (N11657, N11637, N2500);
buf BUF1 (N11658, N11652);
xor XOR2 (N11659, N11651, N5463);
and AND4 (N11660, N11658, N8223, N6398, N9026);
and AND2 (N11661, N11660, N9140);
and AND3 (N11662, N11653, N9160, N2517);
not NOT1 (N11663, N11661);
and AND4 (N11664, N11646, N271, N502, N3194);
xor XOR2 (N11665, N11663, N608);
or OR4 (N11666, N11656, N6858, N11197, N8202);
buf BUF1 (N11667, N11662);
and AND2 (N11668, N11633, N3395);
nand NAND4 (N11669, N11654, N9581, N4289, N9188);
nor NOR4 (N11670, N11659, N8128, N7496, N9636);
or OR2 (N11671, N11664, N11307);
buf BUF1 (N11672, N11671);
buf BUF1 (N11673, N11657);
and AND2 (N11674, N11667, N1443);
buf BUF1 (N11675, N11668);
or OR4 (N11676, N11666, N6879, N3552, N8208);
not NOT1 (N11677, N11675);
or OR3 (N11678, N11670, N8871, N8209);
or OR3 (N11679, N11655, N954, N9474);
xor XOR2 (N11680, N11673, N9691);
nand NAND2 (N11681, N11665, N6354);
or OR4 (N11682, N11681, N4240, N4276, N10954);
nand NAND2 (N11683, N11674, N448);
not NOT1 (N11684, N11677);
and AND4 (N11685, N11683, N8831, N10786, N725);
not NOT1 (N11686, N11628);
and AND3 (N11687, N11672, N3254, N6710);
not NOT1 (N11688, N11684);
xor XOR2 (N11689, N11685, N4428);
nor NOR4 (N11690, N11689, N2466, N4079, N4154);
and AND3 (N11691, N11687, N2770, N8430);
buf BUF1 (N11692, N11682);
and AND4 (N11693, N11680, N5659, N5849, N2053);
nand NAND4 (N11694, N11686, N480, N11420, N5705);
buf BUF1 (N11695, N11676);
not NOT1 (N11696, N11678);
not NOT1 (N11697, N11695);
or OR4 (N11698, N11691, N2043, N6337, N9841);
nor NOR2 (N11699, N11697, N4871);
xor XOR2 (N11700, N11679, N9895);
buf BUF1 (N11701, N11694);
buf BUF1 (N11702, N11688);
xor XOR2 (N11703, N11700, N7376);
xor XOR2 (N11704, N11696, N2531);
and AND4 (N11705, N11690, N8898, N11054, N350);
and AND4 (N11706, N11702, N7005, N10647, N9116);
and AND2 (N11707, N11699, N10530);
nor NOR3 (N11708, N11698, N2464, N1154);
not NOT1 (N11709, N11708);
buf BUF1 (N11710, N11703);
or OR4 (N11711, N11707, N3246, N6588, N11298);
and AND4 (N11712, N11704, N7983, N4883, N3123);
xor XOR2 (N11713, N11701, N11416);
and AND3 (N11714, N11712, N819, N9331);
nor NOR2 (N11715, N11706, N1614);
nor NOR4 (N11716, N11705, N996, N4497, N1804);
or OR3 (N11717, N11693, N10441, N5341);
xor XOR2 (N11718, N11669, N10252);
xor XOR2 (N11719, N11692, N535);
nand NAND3 (N11720, N11711, N1312, N4289);
not NOT1 (N11721, N11720);
not NOT1 (N11722, N11715);
not NOT1 (N11723, N11709);
and AND3 (N11724, N11717, N9698, N5911);
xor XOR2 (N11725, N11721, N9579);
buf BUF1 (N11726, N11714);
nor NOR4 (N11727, N11710, N7475, N6799, N2094);
nor NOR4 (N11728, N11718, N5689, N10745, N8709);
xor XOR2 (N11729, N11719, N971);
nand NAND4 (N11730, N11724, N7634, N5795, N6851);
not NOT1 (N11731, N11727);
buf BUF1 (N11732, N11716);
nor NOR2 (N11733, N11732, N2886);
nand NAND3 (N11734, N11730, N92, N8155);
buf BUF1 (N11735, N11734);
nand NAND3 (N11736, N11728, N7714, N11653);
xor XOR2 (N11737, N11722, N3753);
nand NAND4 (N11738, N11731, N9935, N7754, N9887);
or OR3 (N11739, N11726, N4681, N6318);
xor XOR2 (N11740, N11735, N4160);
and AND3 (N11741, N11736, N11652, N7160);
buf BUF1 (N11742, N11740);
or OR4 (N11743, N11733, N4121, N353, N2672);
not NOT1 (N11744, N11743);
xor XOR2 (N11745, N11737, N10766);
xor XOR2 (N11746, N11739, N10671);
buf BUF1 (N11747, N11744);
xor XOR2 (N11748, N11713, N6149);
or OR3 (N11749, N11738, N9848, N190);
xor XOR2 (N11750, N11741, N8830);
or OR2 (N11751, N11725, N856);
or OR4 (N11752, N11749, N3367, N5297, N333);
and AND4 (N11753, N11746, N1398, N2762, N9200);
not NOT1 (N11754, N11745);
xor XOR2 (N11755, N11729, N93);
or OR3 (N11756, N11748, N10001, N11310);
xor XOR2 (N11757, N11750, N7007);
nor NOR3 (N11758, N11747, N4998, N5550);
nor NOR3 (N11759, N11723, N3726, N11192);
nand NAND3 (N11760, N11758, N1792, N7845);
xor XOR2 (N11761, N11752, N1527);
not NOT1 (N11762, N11761);
or OR2 (N11763, N11760, N3642);
nand NAND2 (N11764, N11754, N3147);
nand NAND3 (N11765, N11757, N1150, N9792);
or OR4 (N11766, N11742, N1307, N1327, N8721);
not NOT1 (N11767, N11759);
xor XOR2 (N11768, N11756, N6094);
buf BUF1 (N11769, N11764);
xor XOR2 (N11770, N11763, N3106);
not NOT1 (N11771, N11751);
nand NAND2 (N11772, N11765, N3756);
or OR2 (N11773, N11755, N7786);
nor NOR2 (N11774, N11767, N5194);
xor XOR2 (N11775, N11771, N3664);
or OR3 (N11776, N11770, N8962, N201);
nand NAND4 (N11777, N11772, N934, N11651, N10183);
and AND3 (N11778, N11768, N5043, N2010);
nand NAND2 (N11779, N11778, N11699);
nand NAND2 (N11780, N11753, N1594);
and AND2 (N11781, N11762, N4649);
and AND4 (N11782, N11766, N9959, N7616, N8336);
buf BUF1 (N11783, N11780);
or OR3 (N11784, N11769, N5231, N3738);
not NOT1 (N11785, N11777);
and AND3 (N11786, N11784, N6435, N8995);
not NOT1 (N11787, N11776);
and AND3 (N11788, N11785, N390, N11571);
nor NOR4 (N11789, N11788, N3086, N9500, N6103);
and AND4 (N11790, N11775, N192, N764, N11729);
and AND3 (N11791, N11779, N2149, N11483);
nor NOR4 (N11792, N11782, N2453, N3662, N805);
and AND2 (N11793, N11773, N1383);
nand NAND3 (N11794, N11793, N5248, N972);
xor XOR2 (N11795, N11783, N1607);
or OR3 (N11796, N11791, N11645, N5216);
buf BUF1 (N11797, N11790);
nand NAND3 (N11798, N11781, N3200, N7708);
xor XOR2 (N11799, N11795, N2801);
buf BUF1 (N11800, N11774);
nor NOR4 (N11801, N11789, N7102, N1815, N5410);
not NOT1 (N11802, N11797);
not NOT1 (N11803, N11796);
nand NAND4 (N11804, N11792, N5654, N5347, N11356);
nand NAND3 (N11805, N11803, N9240, N6337);
nand NAND2 (N11806, N11804, N11345);
xor XOR2 (N11807, N11806, N6042);
and AND3 (N11808, N11805, N8344, N4816);
or OR3 (N11809, N11787, N3934, N511);
xor XOR2 (N11810, N11809, N740);
nor NOR4 (N11811, N11808, N9318, N115, N3229);
and AND3 (N11812, N11802, N8704, N5557);
buf BUF1 (N11813, N11786);
nand NAND2 (N11814, N11813, N1064);
nor NOR4 (N11815, N11811, N565, N2640, N8177);
buf BUF1 (N11816, N11807);
or OR2 (N11817, N11798, N2522);
and AND2 (N11818, N11810, N9716);
xor XOR2 (N11819, N11801, N1687);
not NOT1 (N11820, N11816);
or OR4 (N11821, N11820, N6087, N6162, N745);
not NOT1 (N11822, N11815);
nor NOR2 (N11823, N11814, N7978);
nand NAND4 (N11824, N11819, N1897, N7706, N5182);
nor NOR4 (N11825, N11799, N2790, N7165, N8867);
xor XOR2 (N11826, N11823, N4827);
not NOT1 (N11827, N11822);
and AND2 (N11828, N11800, N8329);
not NOT1 (N11829, N11826);
and AND2 (N11830, N11794, N3862);
buf BUF1 (N11831, N11828);
buf BUF1 (N11832, N11824);
xor XOR2 (N11833, N11818, N10196);
buf BUF1 (N11834, N11829);
or OR3 (N11835, N11834, N2856, N5997);
buf BUF1 (N11836, N11832);
xor XOR2 (N11837, N11831, N10872);
buf BUF1 (N11838, N11817);
buf BUF1 (N11839, N11837);
xor XOR2 (N11840, N11839, N7073);
and AND2 (N11841, N11833, N2261);
xor XOR2 (N11842, N11838, N1746);
buf BUF1 (N11843, N11830);
buf BUF1 (N11844, N11821);
and AND2 (N11845, N11812, N3305);
buf BUF1 (N11846, N11841);
or OR4 (N11847, N11842, N769, N10501, N4890);
buf BUF1 (N11848, N11827);
nor NOR3 (N11849, N11840, N5362, N4126);
xor XOR2 (N11850, N11848, N2642);
and AND4 (N11851, N11850, N11736, N5440, N2034);
not NOT1 (N11852, N11825);
nor NOR3 (N11853, N11851, N5143, N10583);
xor XOR2 (N11854, N11852, N1825);
nand NAND3 (N11855, N11836, N11266, N9031);
buf BUF1 (N11856, N11835);
and AND2 (N11857, N11856, N3098);
nor NOR4 (N11858, N11849, N4612, N6364, N6724);
buf BUF1 (N11859, N11846);
nor NOR3 (N11860, N11843, N1170, N5748);
nand NAND2 (N11861, N11844, N10988);
nand NAND4 (N11862, N11861, N7016, N6283, N11041);
and AND2 (N11863, N11857, N2588);
buf BUF1 (N11864, N11863);
xor XOR2 (N11865, N11853, N7096);
and AND4 (N11866, N11858, N11243, N9666, N2546);
nand NAND2 (N11867, N11845, N4887);
not NOT1 (N11868, N11855);
nor NOR2 (N11869, N11854, N9723);
nor NOR3 (N11870, N11867, N3486, N6657);
or OR4 (N11871, N11866, N9656, N10222, N5023);
nor NOR4 (N11872, N11868, N9674, N6826, N3462);
or OR4 (N11873, N11872, N6979, N9182, N4259);
and AND3 (N11874, N11860, N10875, N10500);
not NOT1 (N11875, N11871);
nor NOR4 (N11876, N11874, N11523, N6190, N4958);
and AND2 (N11877, N11876, N11086);
and AND4 (N11878, N11875, N6038, N4897, N7905);
buf BUF1 (N11879, N11870);
and AND3 (N11880, N11865, N1312, N11060);
or OR4 (N11881, N11859, N2653, N4853, N7427);
not NOT1 (N11882, N11881);
buf BUF1 (N11883, N11847);
or OR4 (N11884, N11883, N6924, N418, N5612);
xor XOR2 (N11885, N11873, N8641);
and AND4 (N11886, N11862, N7829, N10864, N722);
nor NOR2 (N11887, N11884, N2537);
xor XOR2 (N11888, N11877, N938);
not NOT1 (N11889, N11880);
nor NOR4 (N11890, N11885, N4465, N8622, N2527);
and AND2 (N11891, N11878, N8473);
and AND4 (N11892, N11879, N3171, N3779, N86);
xor XOR2 (N11893, N11892, N1032);
buf BUF1 (N11894, N11890);
nor NOR2 (N11895, N11894, N4295);
nand NAND3 (N11896, N11882, N4931, N5796);
and AND3 (N11897, N11895, N4312, N3188);
nor NOR2 (N11898, N11887, N8557);
nor NOR3 (N11899, N11898, N1863, N11711);
xor XOR2 (N11900, N11869, N7688);
not NOT1 (N11901, N11899);
buf BUF1 (N11902, N11889);
buf BUF1 (N11903, N11900);
buf BUF1 (N11904, N11896);
and AND2 (N11905, N11902, N9209);
nor NOR4 (N11906, N11893, N7524, N6595, N8318);
nand NAND4 (N11907, N11903, N3118, N7102, N3050);
not NOT1 (N11908, N11891);
not NOT1 (N11909, N11901);
not NOT1 (N11910, N11909);
and AND4 (N11911, N11904, N11410, N2982, N11457);
not NOT1 (N11912, N11897);
nand NAND4 (N11913, N11864, N11754, N7052, N1690);
not NOT1 (N11914, N11908);
and AND2 (N11915, N11913, N9374);
nor NOR3 (N11916, N11914, N11002, N5401);
and AND4 (N11917, N11916, N8541, N10867, N6452);
and AND4 (N11918, N11912, N8347, N11017, N2144);
nand NAND4 (N11919, N11910, N7451, N9119, N8003);
and AND3 (N11920, N11915, N2051, N554);
xor XOR2 (N11921, N11919, N4337);
and AND4 (N11922, N11888, N2503, N805, N8361);
buf BUF1 (N11923, N11921);
and AND2 (N11924, N11886, N10102);
xor XOR2 (N11925, N11906, N7451);
nor NOR3 (N11926, N11905, N2215, N11084);
xor XOR2 (N11927, N11922, N2973);
nor NOR3 (N11928, N11926, N11737, N2029);
nor NOR4 (N11929, N11920, N9964, N545, N8143);
buf BUF1 (N11930, N11907);
xor XOR2 (N11931, N11930, N1621);
nand NAND2 (N11932, N11927, N4793);
and AND4 (N11933, N11911, N4780, N625, N5793);
nand NAND4 (N11934, N11923, N2570, N6687, N11797);
buf BUF1 (N11935, N11934);
not NOT1 (N11936, N11933);
or OR3 (N11937, N11918, N8347, N5203);
nor NOR3 (N11938, N11936, N11120, N248);
xor XOR2 (N11939, N11932, N970);
not NOT1 (N11940, N11931);
and AND3 (N11941, N11925, N6654, N10326);
buf BUF1 (N11942, N11928);
nand NAND4 (N11943, N11942, N1073, N6039, N494);
nor NOR3 (N11944, N11924, N6047, N9646);
and AND2 (N11945, N11929, N7353);
or OR3 (N11946, N11938, N11699, N7940);
and AND4 (N11947, N11935, N7893, N11548, N1558);
nor NOR2 (N11948, N11946, N4832);
or OR2 (N11949, N11939, N11526);
or OR3 (N11950, N11944, N3145, N6229);
nor NOR3 (N11951, N11945, N4516, N11782);
xor XOR2 (N11952, N11941, N4323);
nor NOR3 (N11953, N11937, N9054, N3360);
buf BUF1 (N11954, N11943);
or OR4 (N11955, N11951, N3394, N7310, N10207);
not NOT1 (N11956, N11949);
nor NOR4 (N11957, N11953, N1814, N7088, N6813);
nand NAND3 (N11958, N11957, N11187, N8909);
xor XOR2 (N11959, N11917, N3810);
not NOT1 (N11960, N11940);
xor XOR2 (N11961, N11950, N5028);
and AND3 (N11962, N11956, N4277, N4160);
nand NAND2 (N11963, N11952, N3934);
and AND4 (N11964, N11962, N10453, N1047, N2794);
and AND2 (N11965, N11947, N1541);
nor NOR4 (N11966, N11948, N1298, N2130, N1825);
nand NAND3 (N11967, N11961, N6526, N10178);
xor XOR2 (N11968, N11964, N5147);
buf BUF1 (N11969, N11963);
not NOT1 (N11970, N11968);
nand NAND3 (N11971, N11959, N1940, N6067);
or OR2 (N11972, N11971, N6454);
or OR4 (N11973, N11954, N8558, N2555, N9898);
buf BUF1 (N11974, N11970);
nor NOR3 (N11975, N11972, N10952, N8360);
xor XOR2 (N11976, N11955, N11154);
buf BUF1 (N11977, N11974);
and AND2 (N11978, N11977, N7285);
nand NAND2 (N11979, N11976, N7474);
or OR4 (N11980, N11975, N8955, N3301, N5580);
nand NAND2 (N11981, N11973, N9629);
nor NOR4 (N11982, N11967, N2527, N9515, N7249);
nor NOR3 (N11983, N11979, N2694, N6221);
buf BUF1 (N11984, N11969);
xor XOR2 (N11985, N11965, N1270);
or OR3 (N11986, N11980, N2218, N5223);
nor NOR3 (N11987, N11983, N4362, N8225);
nor NOR2 (N11988, N11960, N4677);
buf BUF1 (N11989, N11982);
not NOT1 (N11990, N11985);
buf BUF1 (N11991, N11990);
nand NAND4 (N11992, N11988, N7541, N2607, N5653);
buf BUF1 (N11993, N11984);
and AND3 (N11994, N11992, N2913, N2136);
or OR3 (N11995, N11981, N11949, N8597);
not NOT1 (N11996, N11978);
and AND3 (N11997, N11987, N6372, N7226);
nor NOR3 (N11998, N11995, N2035, N5633);
nand NAND2 (N11999, N11994, N1166);
or OR3 (N12000, N11996, N7392, N11749);
not NOT1 (N12001, N11986);
or OR2 (N12002, N11998, N9087);
and AND4 (N12003, N11989, N8768, N7048, N10531);
xor XOR2 (N12004, N12000, N1855);
and AND3 (N12005, N11999, N5046, N10110);
nand NAND3 (N12006, N12002, N9529, N7078);
not NOT1 (N12007, N11991);
xor XOR2 (N12008, N11997, N2222);
buf BUF1 (N12009, N12005);
nand NAND4 (N12010, N12008, N7348, N4222, N1350);
xor XOR2 (N12011, N12010, N3301);
or OR3 (N12012, N12003, N5254, N8767);
buf BUF1 (N12013, N12012);
or OR3 (N12014, N12011, N1633, N2131);
or OR2 (N12015, N12006, N7222);
buf BUF1 (N12016, N12009);
nand NAND2 (N12017, N12007, N1539);
and AND3 (N12018, N11958, N11111, N10140);
or OR2 (N12019, N12014, N9630);
not NOT1 (N12020, N12001);
nand NAND2 (N12021, N12018, N8533);
nor NOR3 (N12022, N12013, N8856, N6078);
buf BUF1 (N12023, N12022);
nand NAND2 (N12024, N12016, N6669);
xor XOR2 (N12025, N12021, N11390);
and AND3 (N12026, N12023, N4179, N11008);
nor NOR4 (N12027, N12020, N3686, N11317, N7510);
or OR3 (N12028, N12017, N9924, N10670);
nor NOR3 (N12029, N12026, N5934, N10809);
nand NAND3 (N12030, N12019, N766, N9630);
and AND4 (N12031, N12030, N4695, N5770, N2947);
nor NOR2 (N12032, N12024, N3107);
or OR4 (N12033, N12032, N10339, N8701, N4952);
nor NOR3 (N12034, N12029, N11552, N1547);
nand NAND2 (N12035, N12025, N3756);
and AND3 (N12036, N11966, N1589, N4696);
not NOT1 (N12037, N12033);
xor XOR2 (N12038, N11993, N39);
buf BUF1 (N12039, N12034);
nor NOR4 (N12040, N12015, N1084, N5339, N8650);
or OR4 (N12041, N12027, N11535, N6648, N5415);
or OR3 (N12042, N12036, N3886, N2493);
nand NAND3 (N12043, N12031, N3732, N10545);
nor NOR3 (N12044, N12038, N4963, N5329);
nand NAND4 (N12045, N12028, N6203, N8856, N3126);
not NOT1 (N12046, N12037);
buf BUF1 (N12047, N12035);
xor XOR2 (N12048, N12041, N936);
xor XOR2 (N12049, N12046, N6056);
nand NAND2 (N12050, N12040, N796);
and AND2 (N12051, N12042, N9794);
not NOT1 (N12052, N12051);
or OR4 (N12053, N12050, N4760, N44, N795);
xor XOR2 (N12054, N12039, N7815);
nand NAND3 (N12055, N12047, N9553, N9130);
not NOT1 (N12056, N12048);
nand NAND4 (N12057, N12043, N5095, N6591, N3913);
or OR3 (N12058, N12052, N10182, N6706);
xor XOR2 (N12059, N12055, N9017);
not NOT1 (N12060, N12049);
not NOT1 (N12061, N12045);
buf BUF1 (N12062, N12053);
or OR3 (N12063, N12059, N11128, N8210);
xor XOR2 (N12064, N12060, N8345);
xor XOR2 (N12065, N12044, N1013);
not NOT1 (N12066, N12057);
xor XOR2 (N12067, N12054, N9241);
not NOT1 (N12068, N12058);
xor XOR2 (N12069, N12062, N11683);
buf BUF1 (N12070, N12065);
nand NAND2 (N12071, N12064, N6364);
or OR3 (N12072, N12071, N6870, N6481);
buf BUF1 (N12073, N12061);
nor NOR3 (N12074, N12073, N1339, N7576);
buf BUF1 (N12075, N12068);
xor XOR2 (N12076, N12056, N3793);
not NOT1 (N12077, N12066);
and AND4 (N12078, N12069, N887, N6846, N8414);
nor NOR4 (N12079, N12063, N11027, N6767, N10325);
not NOT1 (N12080, N12076);
not NOT1 (N12081, N12075);
or OR3 (N12082, N12072, N11304, N2222);
nor NOR2 (N12083, N12079, N10649);
xor XOR2 (N12084, N12077, N985);
nor NOR4 (N12085, N12078, N9538, N11787, N7);
nor NOR2 (N12086, N12004, N2749);
and AND2 (N12087, N12081, N8621);
buf BUF1 (N12088, N12086);
nand NAND2 (N12089, N12088, N7402);
not NOT1 (N12090, N12087);
and AND3 (N12091, N12083, N2467, N1104);
and AND2 (N12092, N12089, N3599);
nor NOR2 (N12093, N12084, N1823);
or OR4 (N12094, N12090, N6894, N11219, N7258);
nand NAND2 (N12095, N12092, N7195);
or OR4 (N12096, N12093, N9592, N2681, N1088);
not NOT1 (N12097, N12067);
nor NOR2 (N12098, N12080, N2915);
buf BUF1 (N12099, N12096);
xor XOR2 (N12100, N12097, N430);
nand NAND4 (N12101, N12070, N10635, N837, N6880);
not NOT1 (N12102, N12091);
and AND3 (N12103, N12098, N4708, N5017);
nor NOR4 (N12104, N12103, N3750, N7150, N11952);
and AND2 (N12105, N12099, N5169);
xor XOR2 (N12106, N12094, N10923);
or OR2 (N12107, N12082, N10985);
nand NAND3 (N12108, N12100, N3587, N2780);
nand NAND4 (N12109, N12105, N6028, N10649, N8335);
xor XOR2 (N12110, N12095, N9479);
or OR4 (N12111, N12110, N2534, N5819, N11181);
buf BUF1 (N12112, N12085);
and AND4 (N12113, N12074, N1596, N10683, N11548);
and AND2 (N12114, N12104, N3493);
or OR3 (N12115, N12114, N2591, N1088);
xor XOR2 (N12116, N12115, N1476);
buf BUF1 (N12117, N12108);
not NOT1 (N12118, N12111);
not NOT1 (N12119, N12117);
buf BUF1 (N12120, N12102);
xor XOR2 (N12121, N12109, N5835);
and AND4 (N12122, N12120, N3188, N11776, N1186);
not NOT1 (N12123, N12121);
buf BUF1 (N12124, N12113);
buf BUF1 (N12125, N12118);
buf BUF1 (N12126, N12123);
not NOT1 (N12127, N12119);
nand NAND3 (N12128, N12124, N7467, N10704);
and AND3 (N12129, N12126, N10838, N2290);
buf BUF1 (N12130, N12116);
xor XOR2 (N12131, N12127, N3750);
buf BUF1 (N12132, N12122);
or OR2 (N12133, N12129, N2481);
xor XOR2 (N12134, N12131, N6114);
or OR2 (N12135, N12130, N8718);
or OR4 (N12136, N12112, N7119, N5633, N3383);
or OR2 (N12137, N12128, N7513);
and AND3 (N12138, N12132, N9849, N3934);
buf BUF1 (N12139, N12107);
not NOT1 (N12140, N12134);
nand NAND2 (N12141, N12139, N10755);
nor NOR4 (N12142, N12137, N9762, N9943, N8011);
buf BUF1 (N12143, N12138);
or OR2 (N12144, N12101, N9346);
nor NOR4 (N12145, N12136, N6663, N660, N965);
xor XOR2 (N12146, N12125, N11402);
xor XOR2 (N12147, N12135, N1018);
nand NAND4 (N12148, N12106, N3759, N12068, N6587);
nor NOR4 (N12149, N12143, N11096, N11769, N8661);
and AND3 (N12150, N12145, N8965, N9593);
nor NOR3 (N12151, N12133, N8247, N10358);
and AND3 (N12152, N12148, N1573, N1358);
buf BUF1 (N12153, N12142);
and AND3 (N12154, N12149, N1544, N4105);
nor NOR4 (N12155, N12140, N9635, N9764, N6107);
nand NAND3 (N12156, N12144, N4547, N5678);
not NOT1 (N12157, N12152);
nor NOR2 (N12158, N12147, N8875);
or OR2 (N12159, N12157, N2458);
nand NAND4 (N12160, N12150, N9346, N673, N79);
or OR3 (N12161, N12160, N6116, N1303);
and AND4 (N12162, N12158, N4948, N2275, N8455);
nand NAND2 (N12163, N12156, N3446);
and AND2 (N12164, N12163, N5207);
not NOT1 (N12165, N12159);
and AND3 (N12166, N12164, N11786, N2756);
xor XOR2 (N12167, N12166, N9219);
or OR2 (N12168, N12141, N2806);
nand NAND2 (N12169, N12165, N11021);
and AND2 (N12170, N12146, N10792);
nand NAND2 (N12171, N12169, N5220);
xor XOR2 (N12172, N12154, N6158);
not NOT1 (N12173, N12161);
buf BUF1 (N12174, N12168);
nand NAND2 (N12175, N12174, N1119);
buf BUF1 (N12176, N12173);
buf BUF1 (N12177, N12162);
nor NOR3 (N12178, N12177, N8014, N11836);
not NOT1 (N12179, N12172);
xor XOR2 (N12180, N12175, N8140);
buf BUF1 (N12181, N12153);
nor NOR4 (N12182, N12176, N495, N3579, N7713);
not NOT1 (N12183, N12178);
nand NAND3 (N12184, N12181, N11759, N11351);
not NOT1 (N12185, N12171);
not NOT1 (N12186, N12179);
not NOT1 (N12187, N12185);
nand NAND2 (N12188, N12187, N5085);
buf BUF1 (N12189, N12188);
nor NOR3 (N12190, N12155, N1392, N11154);
or OR4 (N12191, N12170, N6329, N7285, N1729);
buf BUF1 (N12192, N12151);
or OR2 (N12193, N12191, N11694);
nand NAND4 (N12194, N12193, N11811, N3284, N5807);
buf BUF1 (N12195, N12190);
nor NOR3 (N12196, N12194, N3392, N2062);
xor XOR2 (N12197, N12184, N7477);
and AND2 (N12198, N12182, N3588);
and AND2 (N12199, N12189, N766);
not NOT1 (N12200, N12198);
and AND2 (N12201, N12186, N2803);
nand NAND4 (N12202, N12167, N3005, N11969, N11968);
and AND4 (N12203, N12200, N7415, N3986, N8731);
xor XOR2 (N12204, N12199, N10248);
or OR2 (N12205, N12195, N8410);
xor XOR2 (N12206, N12204, N8005);
and AND2 (N12207, N12206, N5024);
and AND3 (N12208, N12183, N8838, N7721);
or OR3 (N12209, N12202, N3952, N559);
or OR4 (N12210, N12180, N3544, N10073, N6900);
not NOT1 (N12211, N12203);
and AND2 (N12212, N12197, N3446);
and AND2 (N12213, N12205, N2838);
nor NOR2 (N12214, N12207, N10033);
xor XOR2 (N12215, N12211, N7852);
xor XOR2 (N12216, N12214, N7125);
nor NOR2 (N12217, N12196, N8561);
and AND3 (N12218, N12216, N12086, N5356);
buf BUF1 (N12219, N12201);
not NOT1 (N12220, N12209);
not NOT1 (N12221, N12220);
not NOT1 (N12222, N12212);
or OR2 (N12223, N12213, N9675);
or OR4 (N12224, N12223, N3719, N5248, N9712);
and AND3 (N12225, N12208, N8405, N4158);
nand NAND3 (N12226, N12222, N10772, N870);
and AND3 (N12227, N12215, N4995, N6760);
or OR4 (N12228, N12226, N4909, N2705, N6515);
and AND4 (N12229, N12221, N7648, N3623, N6586);
buf BUF1 (N12230, N12225);
not NOT1 (N12231, N12227);
nand NAND4 (N12232, N12229, N8533, N3709, N8380);
not NOT1 (N12233, N12210);
nor NOR3 (N12234, N12230, N5079, N9560);
nor NOR4 (N12235, N12231, N9757, N12147, N8088);
not NOT1 (N12236, N12232);
not NOT1 (N12237, N12217);
not NOT1 (N12238, N12218);
and AND3 (N12239, N12236, N2637, N7851);
buf BUF1 (N12240, N12219);
or OR2 (N12241, N12224, N5744);
not NOT1 (N12242, N12234);
nand NAND3 (N12243, N12241, N2037, N9897);
nor NOR2 (N12244, N12238, N6530);
buf BUF1 (N12245, N12237);
and AND2 (N12246, N12240, N4626);
not NOT1 (N12247, N12235);
buf BUF1 (N12248, N12247);
and AND3 (N12249, N12246, N10301, N10544);
nand NAND2 (N12250, N12239, N791);
and AND2 (N12251, N12192, N8443);
not NOT1 (N12252, N12244);
or OR2 (N12253, N12252, N10513);
nand NAND2 (N12254, N12251, N8512);
or OR4 (N12255, N12242, N9331, N711, N9243);
not NOT1 (N12256, N12249);
or OR2 (N12257, N12228, N5454);
xor XOR2 (N12258, N12254, N2021);
not NOT1 (N12259, N12256);
nand NAND4 (N12260, N12233, N11763, N3149, N8130);
not NOT1 (N12261, N12253);
and AND3 (N12262, N12260, N1960, N2487);
and AND2 (N12263, N12248, N7275);
not NOT1 (N12264, N12245);
xor XOR2 (N12265, N12255, N3328);
nand NAND4 (N12266, N12261, N8040, N9293, N3059);
xor XOR2 (N12267, N12243, N7481);
and AND4 (N12268, N12250, N7875, N2775, N2037);
nor NOR3 (N12269, N12259, N5105, N5026);
xor XOR2 (N12270, N12258, N9400);
xor XOR2 (N12271, N12267, N9766);
nand NAND3 (N12272, N12265, N495, N10692);
not NOT1 (N12273, N12257);
not NOT1 (N12274, N12269);
and AND2 (N12275, N12273, N1685);
and AND2 (N12276, N12275, N6731);
not NOT1 (N12277, N12276);
nor NOR2 (N12278, N12272, N3473);
nor NOR2 (N12279, N12262, N184);
and AND2 (N12280, N12263, N4559);
not NOT1 (N12281, N12270);
and AND2 (N12282, N12266, N4255);
nand NAND2 (N12283, N12274, N10467);
xor XOR2 (N12284, N12271, N3862);
and AND3 (N12285, N12264, N3959, N7759);
buf BUF1 (N12286, N12277);
or OR4 (N12287, N12285, N5403, N4593, N1992);
nand NAND3 (N12288, N12281, N2294, N913);
and AND4 (N12289, N12282, N6770, N12093, N511);
not NOT1 (N12290, N12283);
or OR3 (N12291, N12288, N11160, N2313);
and AND3 (N12292, N12278, N11174, N8481);
and AND3 (N12293, N12280, N10773, N6473);
or OR4 (N12294, N12290, N9921, N5770, N1653);
buf BUF1 (N12295, N12268);
buf BUF1 (N12296, N12293);
xor XOR2 (N12297, N12286, N5148);
not NOT1 (N12298, N12295);
xor XOR2 (N12299, N12287, N6853);
not NOT1 (N12300, N12297);
nand NAND3 (N12301, N12299, N4777, N9027);
nand NAND2 (N12302, N12284, N7967);
nand NAND2 (N12303, N12291, N9736);
and AND4 (N12304, N12300, N9781, N3493, N129);
or OR4 (N12305, N12289, N10604, N10093, N3742);
nor NOR2 (N12306, N12292, N6247);
xor XOR2 (N12307, N12306, N9984);
xor XOR2 (N12308, N12303, N5474);
nor NOR3 (N12309, N12301, N3598, N2374);
or OR4 (N12310, N12298, N8891, N11399, N8989);
xor XOR2 (N12311, N12310, N4921);
and AND4 (N12312, N12311, N7095, N11877, N2132);
or OR3 (N12313, N12305, N8628, N9370);
not NOT1 (N12314, N12279);
not NOT1 (N12315, N12312);
nand NAND4 (N12316, N12304, N4740, N10175, N7434);
buf BUF1 (N12317, N12307);
and AND4 (N12318, N12296, N8722, N9233, N7871);
and AND4 (N12319, N12315, N2437, N759, N9594);
and AND3 (N12320, N12319, N946, N6497);
nand NAND4 (N12321, N12316, N9756, N7950, N7305);
buf BUF1 (N12322, N12313);
xor XOR2 (N12323, N12317, N9255);
and AND3 (N12324, N12322, N4882, N3742);
nand NAND2 (N12325, N12302, N12246);
and AND3 (N12326, N12323, N5807, N11890);
and AND4 (N12327, N12314, N11324, N10305, N9250);
not NOT1 (N12328, N12325);
not NOT1 (N12329, N12320);
buf BUF1 (N12330, N12309);
nand NAND4 (N12331, N12328, N8324, N10400, N12164);
nor NOR4 (N12332, N12330, N1488, N2757, N10323);
not NOT1 (N12333, N12318);
buf BUF1 (N12334, N12327);
buf BUF1 (N12335, N12331);
or OR2 (N12336, N12332, N11199);
xor XOR2 (N12337, N12324, N115);
nand NAND3 (N12338, N12294, N7088, N5220);
nand NAND3 (N12339, N12335, N2390, N9874);
nor NOR3 (N12340, N12329, N9291, N9181);
xor XOR2 (N12341, N12336, N2884);
nor NOR3 (N12342, N12341, N4652, N7664);
buf BUF1 (N12343, N12338);
not NOT1 (N12344, N12321);
and AND2 (N12345, N12344, N7201);
or OR3 (N12346, N12326, N10919, N1839);
and AND3 (N12347, N12334, N1101, N11329);
xor XOR2 (N12348, N12308, N4453);
nor NOR4 (N12349, N12343, N2808, N10530, N5995);
not NOT1 (N12350, N12337);
xor XOR2 (N12351, N12350, N11112);
or OR4 (N12352, N12345, N7275, N3771, N5193);
and AND4 (N12353, N12348, N2429, N6866, N4095);
buf BUF1 (N12354, N12340);
nand NAND3 (N12355, N12349, N5624, N10597);
or OR4 (N12356, N12339, N11499, N5247, N5091);
nand NAND4 (N12357, N12356, N4080, N3887, N5101);
nand NAND3 (N12358, N12347, N5687, N8104);
nand NAND4 (N12359, N12355, N1806, N7201, N1602);
not NOT1 (N12360, N12333);
not NOT1 (N12361, N12342);
xor XOR2 (N12362, N12353, N11618);
nor NOR4 (N12363, N12351, N6934, N3556, N3647);
and AND2 (N12364, N12363, N7097);
or OR2 (N12365, N12361, N10808);
and AND3 (N12366, N12357, N3365, N11480);
and AND2 (N12367, N12358, N11271);
not NOT1 (N12368, N12362);
buf BUF1 (N12369, N12366);
buf BUF1 (N12370, N12346);
buf BUF1 (N12371, N12359);
and AND4 (N12372, N12354, N776, N6542, N7511);
xor XOR2 (N12373, N12360, N2492);
buf BUF1 (N12374, N12369);
nor NOR3 (N12375, N12365, N9659, N3805);
not NOT1 (N12376, N12373);
nor NOR4 (N12377, N12364, N6891, N4125, N12204);
or OR4 (N12378, N12370, N9474, N3605, N1095);
xor XOR2 (N12379, N12352, N3535);
not NOT1 (N12380, N12367);
not NOT1 (N12381, N12379);
nand NAND2 (N12382, N12371, N10702);
and AND2 (N12383, N12376, N3797);
and AND4 (N12384, N12381, N4146, N8490, N5181);
not NOT1 (N12385, N12372);
buf BUF1 (N12386, N12380);
nand NAND3 (N12387, N12377, N11459, N4441);
nor NOR2 (N12388, N12368, N12348);
and AND4 (N12389, N12378, N11418, N7524, N183);
nor NOR4 (N12390, N12388, N4200, N11220, N8593);
and AND2 (N12391, N12390, N5729);
nor NOR3 (N12392, N12387, N3973, N99);
buf BUF1 (N12393, N12389);
nor NOR3 (N12394, N12385, N3007, N2787);
nor NOR2 (N12395, N12374, N4939);
and AND4 (N12396, N12391, N8628, N9011, N10203);
nor NOR2 (N12397, N12394, N10832);
buf BUF1 (N12398, N12392);
buf BUF1 (N12399, N12375);
buf BUF1 (N12400, N12386);
buf BUF1 (N12401, N12398);
and AND2 (N12402, N12400, N4983);
nor NOR3 (N12403, N12384, N7162, N1556);
and AND4 (N12404, N12383, N2831, N2203, N2043);
nand NAND2 (N12405, N12397, N1735);
or OR4 (N12406, N12405, N1623, N1752, N4405);
or OR2 (N12407, N12403, N356);
nand NAND3 (N12408, N12399, N11731, N11195);
and AND3 (N12409, N12406, N4093, N6604);
buf BUF1 (N12410, N12404);
nor NOR3 (N12411, N12396, N11601, N10923);
or OR2 (N12412, N12408, N6591);
or OR3 (N12413, N12395, N9751, N11974);
buf BUF1 (N12414, N12407);
xor XOR2 (N12415, N12413, N6652);
or OR2 (N12416, N12415, N7466);
nor NOR4 (N12417, N12412, N1675, N2054, N3174);
and AND3 (N12418, N12402, N211, N10422);
or OR2 (N12419, N12417, N178);
nor NOR4 (N12420, N12409, N9573, N700, N5628);
xor XOR2 (N12421, N12418, N5543);
buf BUF1 (N12422, N12410);
or OR2 (N12423, N12411, N6119);
nand NAND4 (N12424, N12421, N9634, N12105, N11201);
and AND3 (N12425, N12382, N3285, N5769);
nand NAND4 (N12426, N12393, N6426, N4865, N9692);
or OR2 (N12427, N12426, N10305);
nor NOR3 (N12428, N12401, N9889, N5594);
buf BUF1 (N12429, N12420);
xor XOR2 (N12430, N12419, N8782);
nand NAND3 (N12431, N12429, N539, N3331);
or OR3 (N12432, N12428, N3326, N12223);
buf BUF1 (N12433, N12427);
and AND3 (N12434, N12414, N402, N9535);
not NOT1 (N12435, N12416);
buf BUF1 (N12436, N12430);
buf BUF1 (N12437, N12431);
not NOT1 (N12438, N12424);
or OR4 (N12439, N12432, N626, N410, N6387);
buf BUF1 (N12440, N12423);
xor XOR2 (N12441, N12438, N1647);
xor XOR2 (N12442, N12435, N9947);
nand NAND3 (N12443, N12441, N5251, N8970);
buf BUF1 (N12444, N12425);
nand NAND3 (N12445, N12434, N6515, N91);
and AND4 (N12446, N12445, N849, N6610, N2286);
nand NAND3 (N12447, N12446, N2706, N8480);
nand NAND3 (N12448, N12447, N6753, N10845);
not NOT1 (N12449, N12448);
nor NOR3 (N12450, N12439, N10208, N10533);
and AND2 (N12451, N12436, N10305);
nand NAND2 (N12452, N12440, N11608);
not NOT1 (N12453, N12422);
not NOT1 (N12454, N12451);
nor NOR4 (N12455, N12444, N11418, N6534, N2278);
xor XOR2 (N12456, N12433, N525);
buf BUF1 (N12457, N12453);
and AND3 (N12458, N12449, N3538, N8139);
not NOT1 (N12459, N12457);
or OR4 (N12460, N12456, N1038, N6488, N4438);
not NOT1 (N12461, N12455);
not NOT1 (N12462, N12459);
xor XOR2 (N12463, N12461, N4992);
buf BUF1 (N12464, N12443);
or OR2 (N12465, N12437, N1992);
and AND4 (N12466, N12442, N1302, N11573, N10224);
buf BUF1 (N12467, N12460);
not NOT1 (N12468, N12450);
xor XOR2 (N12469, N12454, N2050);
xor XOR2 (N12470, N12467, N11532);
buf BUF1 (N12471, N12464);
or OR2 (N12472, N12469, N11537);
nor NOR4 (N12473, N12468, N2068, N4671, N6315);
not NOT1 (N12474, N12458);
and AND2 (N12475, N12452, N7855);
not NOT1 (N12476, N12471);
not NOT1 (N12477, N12470);
nand NAND3 (N12478, N12462, N4451, N1932);
buf BUF1 (N12479, N12465);
buf BUF1 (N12480, N12472);
xor XOR2 (N12481, N12479, N11943);
not NOT1 (N12482, N12475);
xor XOR2 (N12483, N12481, N12070);
xor XOR2 (N12484, N12483, N1349);
nor NOR3 (N12485, N12473, N9734, N9271);
xor XOR2 (N12486, N12463, N3671);
and AND2 (N12487, N12484, N4127);
not NOT1 (N12488, N12466);
xor XOR2 (N12489, N12478, N12245);
or OR2 (N12490, N12477, N8243);
and AND2 (N12491, N12474, N492);
nand NAND4 (N12492, N12487, N5130, N759, N2539);
nor NOR3 (N12493, N12491, N8480, N11648);
not NOT1 (N12494, N12488);
or OR4 (N12495, N12482, N194, N11836, N8623);
and AND4 (N12496, N12485, N8493, N8252, N9116);
xor XOR2 (N12497, N12480, N5792);
not NOT1 (N12498, N12497);
buf BUF1 (N12499, N12495);
nor NOR3 (N12500, N12498, N10599, N3364);
and AND2 (N12501, N12494, N6224);
and AND2 (N12502, N12492, N4560);
and AND2 (N12503, N12486, N316);
not NOT1 (N12504, N12493);
not NOT1 (N12505, N12502);
buf BUF1 (N12506, N12490);
or OR4 (N12507, N12501, N12400, N3277, N596);
or OR4 (N12508, N12476, N9004, N9695, N2715);
nand NAND4 (N12509, N12489, N12016, N9890, N1895);
not NOT1 (N12510, N12506);
not NOT1 (N12511, N12496);
or OR2 (N12512, N12510, N5369);
not NOT1 (N12513, N12505);
xor XOR2 (N12514, N12509, N3121);
or OR2 (N12515, N12508, N434);
buf BUF1 (N12516, N12500);
and AND4 (N12517, N12511, N12398, N11245, N5440);
xor XOR2 (N12518, N12499, N10767);
not NOT1 (N12519, N12518);
and AND4 (N12520, N12519, N11505, N8805, N1964);
or OR2 (N12521, N12512, N9560);
xor XOR2 (N12522, N12521, N9860);
buf BUF1 (N12523, N12513);
nor NOR4 (N12524, N12514, N3447, N9069, N6139);
or OR4 (N12525, N12503, N6616, N403, N4294);
nor NOR2 (N12526, N12516, N7934);
xor XOR2 (N12527, N12520, N545);
nand NAND4 (N12528, N12515, N8890, N3579, N2726);
xor XOR2 (N12529, N12527, N8260);
and AND3 (N12530, N12528, N3873, N10885);
xor XOR2 (N12531, N12529, N12394);
buf BUF1 (N12532, N12524);
xor XOR2 (N12533, N12531, N127);
nor NOR2 (N12534, N12533, N12264);
nor NOR3 (N12535, N12504, N7536, N9274);
not NOT1 (N12536, N12525);
or OR2 (N12537, N12522, N5720);
not NOT1 (N12538, N12536);
nand NAND4 (N12539, N12530, N11229, N6245, N4015);
nand NAND3 (N12540, N12535, N12006, N9531);
and AND4 (N12541, N12507, N8951, N782, N7647);
xor XOR2 (N12542, N12517, N3020);
nand NAND2 (N12543, N12538, N10409);
and AND2 (N12544, N12537, N4778);
nand NAND2 (N12545, N12526, N2461);
xor XOR2 (N12546, N12541, N197);
or OR3 (N12547, N12543, N12494, N11005);
or OR3 (N12548, N12534, N1734, N1714);
buf BUF1 (N12549, N12547);
not NOT1 (N12550, N12523);
xor XOR2 (N12551, N12540, N4159);
nor NOR2 (N12552, N12545, N10033);
nand NAND4 (N12553, N12552, N9573, N1305, N3282);
nand NAND3 (N12554, N12548, N961, N1425);
not NOT1 (N12555, N12549);
or OR3 (N12556, N12555, N11448, N825);
nor NOR2 (N12557, N12553, N46);
not NOT1 (N12558, N12542);
nand NAND4 (N12559, N12557, N378, N5132, N1276);
or OR4 (N12560, N12558, N7507, N3267, N8187);
buf BUF1 (N12561, N12560);
not NOT1 (N12562, N12561);
and AND4 (N12563, N12546, N1270, N12458, N9592);
nand NAND3 (N12564, N12551, N7724, N9047);
not NOT1 (N12565, N12550);
buf BUF1 (N12566, N12564);
and AND4 (N12567, N12554, N10344, N3252, N10106);
buf BUF1 (N12568, N12556);
nand NAND2 (N12569, N12539, N10817);
and AND3 (N12570, N12559, N1439, N4705);
not NOT1 (N12571, N12569);
buf BUF1 (N12572, N12562);
nor NOR3 (N12573, N12565, N3279, N2605);
nand NAND3 (N12574, N12563, N10065, N8934);
and AND4 (N12575, N12568, N9760, N5113, N1758);
not NOT1 (N12576, N12575);
nand NAND4 (N12577, N12571, N8637, N2207, N3772);
nand NAND2 (N12578, N12566, N7347);
nor NOR4 (N12579, N12578, N10184, N2625, N8319);
nand NAND4 (N12580, N12576, N2167, N11859, N11969);
or OR4 (N12581, N12567, N5767, N737, N10077);
nor NOR2 (N12582, N12577, N9427);
nor NOR3 (N12583, N12580, N8084, N5087);
nand NAND2 (N12584, N12581, N9147);
nor NOR2 (N12585, N12570, N8704);
buf BUF1 (N12586, N12573);
xor XOR2 (N12587, N12584, N4357);
and AND4 (N12588, N12574, N11804, N11069, N1162);
or OR4 (N12589, N12588, N6843, N156, N11362);
and AND3 (N12590, N12532, N5874, N2956);
nand NAND3 (N12591, N12579, N9703, N8490);
and AND2 (N12592, N12582, N9561);
and AND2 (N12593, N12590, N10433);
nand NAND4 (N12594, N12544, N4400, N1510, N4572);
or OR2 (N12595, N12593, N8179);
buf BUF1 (N12596, N12583);
not NOT1 (N12597, N12585);
not NOT1 (N12598, N12589);
buf BUF1 (N12599, N12591);
buf BUF1 (N12600, N12592);
not NOT1 (N12601, N12596);
buf BUF1 (N12602, N12594);
nand NAND2 (N12603, N12572, N5752);
nand NAND4 (N12604, N12599, N1423, N8930, N349);
nand NAND3 (N12605, N12597, N50, N6107);
xor XOR2 (N12606, N12586, N7688);
not NOT1 (N12607, N12587);
and AND2 (N12608, N12607, N12562);
buf BUF1 (N12609, N12601);
xor XOR2 (N12610, N12603, N11036);
or OR4 (N12611, N12598, N7111, N5517, N7011);
and AND3 (N12612, N12610, N8375, N11529);
or OR3 (N12613, N12612, N10881, N9327);
xor XOR2 (N12614, N12608, N918);
xor XOR2 (N12615, N12605, N9031);
or OR2 (N12616, N12613, N1685);
and AND3 (N12617, N12615, N11042, N6500);
buf BUF1 (N12618, N12609);
not NOT1 (N12619, N12600);
nor NOR2 (N12620, N12611, N3665);
buf BUF1 (N12621, N12616);
buf BUF1 (N12622, N12621);
not NOT1 (N12623, N12606);
not NOT1 (N12624, N12602);
nor NOR3 (N12625, N12604, N2536, N9618);
xor XOR2 (N12626, N12619, N12617);
nor NOR2 (N12627, N2474, N34);
or OR3 (N12628, N12620, N12399, N10299);
not NOT1 (N12629, N12627);
not NOT1 (N12630, N12614);
buf BUF1 (N12631, N12626);
and AND3 (N12632, N12618, N5062, N11135);
nand NAND2 (N12633, N12595, N1844);
and AND3 (N12634, N12631, N5855, N1732);
xor XOR2 (N12635, N12625, N7512);
nand NAND3 (N12636, N12634, N10860, N8737);
buf BUF1 (N12637, N12630);
buf BUF1 (N12638, N12633);
and AND3 (N12639, N12628, N3023, N7504);
or OR4 (N12640, N12636, N2968, N12342, N12222);
buf BUF1 (N12641, N12622);
xor XOR2 (N12642, N12632, N2607);
buf BUF1 (N12643, N12638);
nand NAND2 (N12644, N12641, N10612);
or OR3 (N12645, N12637, N7731, N3831);
not NOT1 (N12646, N12642);
not NOT1 (N12647, N12639);
xor XOR2 (N12648, N12647, N11687);
or OR3 (N12649, N12643, N3315, N3117);
nand NAND2 (N12650, N12623, N3279);
not NOT1 (N12651, N12644);
or OR3 (N12652, N12649, N12315, N5912);
buf BUF1 (N12653, N12629);
xor XOR2 (N12654, N12652, N2322);
and AND2 (N12655, N12635, N8394);
nor NOR4 (N12656, N12653, N918, N6949, N5864);
nand NAND2 (N12657, N12646, N3342);
buf BUF1 (N12658, N12650);
and AND3 (N12659, N12624, N11751, N1963);
or OR4 (N12660, N12651, N11681, N424, N8925);
not NOT1 (N12661, N12645);
not NOT1 (N12662, N12659);
buf BUF1 (N12663, N12657);
and AND4 (N12664, N12654, N6716, N2093, N9287);
nand NAND2 (N12665, N12648, N6770);
nor NOR4 (N12666, N12660, N7681, N3110, N11190);
or OR2 (N12667, N12666, N5076);
nor NOR3 (N12668, N12640, N6726, N1974);
nor NOR4 (N12669, N12663, N8, N11209, N5533);
not NOT1 (N12670, N12656);
xor XOR2 (N12671, N12669, N6340);
nand NAND3 (N12672, N12662, N11983, N3555);
and AND2 (N12673, N12655, N10935);
not NOT1 (N12674, N12664);
not NOT1 (N12675, N12671);
not NOT1 (N12676, N12668);
buf BUF1 (N12677, N12665);
xor XOR2 (N12678, N12675, N4192);
and AND4 (N12679, N12661, N11067, N6981, N4771);
nand NAND4 (N12680, N12676, N123, N8875, N9872);
xor XOR2 (N12681, N12667, N238);
and AND4 (N12682, N12681, N4549, N5332, N5913);
or OR3 (N12683, N12680, N8668, N9488);
nand NAND3 (N12684, N12683, N8601, N8152);
xor XOR2 (N12685, N12677, N1314);
buf BUF1 (N12686, N12685);
nand NAND2 (N12687, N12684, N10671);
nand NAND2 (N12688, N12673, N12413);
and AND4 (N12689, N12679, N2175, N4744, N11321);
and AND3 (N12690, N12682, N9724, N5381);
or OR3 (N12691, N12688, N8598, N688);
and AND4 (N12692, N12670, N1624, N7390, N8853);
nor NOR4 (N12693, N12674, N12536, N4493, N9878);
not NOT1 (N12694, N12658);
nor NOR3 (N12695, N12686, N3884, N3533);
not NOT1 (N12696, N12693);
xor XOR2 (N12697, N12678, N5512);
not NOT1 (N12698, N12691);
and AND4 (N12699, N12697, N1186, N9977, N2721);
xor XOR2 (N12700, N12698, N6320);
buf BUF1 (N12701, N12695);
buf BUF1 (N12702, N12694);
buf BUF1 (N12703, N12690);
nand NAND3 (N12704, N12703, N4962, N1459);
nand NAND4 (N12705, N12699, N12643, N3063, N6596);
nand NAND2 (N12706, N12696, N2342);
nor NOR4 (N12707, N12692, N5684, N11693, N10335);
xor XOR2 (N12708, N12689, N11258);
or OR4 (N12709, N12687, N3927, N7515, N6554);
buf BUF1 (N12710, N12707);
nand NAND2 (N12711, N12704, N12674);
or OR2 (N12712, N12709, N68);
or OR2 (N12713, N12672, N231);
or OR4 (N12714, N12705, N894, N6455, N6148);
buf BUF1 (N12715, N12714);
or OR3 (N12716, N12706, N7420, N2424);
not NOT1 (N12717, N12713);
nor NOR2 (N12718, N12717, N8603);
or OR2 (N12719, N12718, N2572);
xor XOR2 (N12720, N12711, N1285);
buf BUF1 (N12721, N12710);
xor XOR2 (N12722, N12708, N5454);
nor NOR2 (N12723, N12721, N6258);
xor XOR2 (N12724, N12712, N10644);
nand NAND4 (N12725, N12716, N11866, N5993, N8440);
xor XOR2 (N12726, N12702, N6405);
nand NAND4 (N12727, N12723, N2071, N8718, N1202);
nand NAND2 (N12728, N12726, N2870);
not NOT1 (N12729, N12722);
not NOT1 (N12730, N12700);
or OR4 (N12731, N12728, N7312, N6786, N3352);
xor XOR2 (N12732, N12727, N5817);
not NOT1 (N12733, N12719);
nand NAND3 (N12734, N12732, N8044, N9255);
or OR2 (N12735, N12720, N5148);
and AND3 (N12736, N12730, N10157, N12448);
xor XOR2 (N12737, N12731, N9254);
xor XOR2 (N12738, N12701, N8180);
not NOT1 (N12739, N12736);
buf BUF1 (N12740, N12733);
or OR3 (N12741, N12724, N4730, N3555);
xor XOR2 (N12742, N12740, N6515);
xor XOR2 (N12743, N12737, N9686);
buf BUF1 (N12744, N12734);
nor NOR3 (N12745, N12735, N8903, N10705);
nand NAND2 (N12746, N12743, N6090);
and AND3 (N12747, N12744, N8937, N5256);
nand NAND4 (N12748, N12741, N10282, N8912, N7665);
nand NAND4 (N12749, N12729, N1570, N1038, N12117);
buf BUF1 (N12750, N12745);
buf BUF1 (N12751, N12749);
buf BUF1 (N12752, N12739);
nand NAND3 (N12753, N12725, N2572, N8834);
nand NAND3 (N12754, N12748, N5618, N2396);
buf BUF1 (N12755, N12715);
and AND4 (N12756, N12750, N256, N9891, N3985);
nand NAND2 (N12757, N12738, N8607);
xor XOR2 (N12758, N12754, N6391);
buf BUF1 (N12759, N12755);
or OR4 (N12760, N12752, N1816, N8257, N471);
and AND4 (N12761, N12753, N9059, N12124, N7579);
xor XOR2 (N12762, N12746, N10334);
buf BUF1 (N12763, N12742);
buf BUF1 (N12764, N12747);
nor NOR4 (N12765, N12758, N4780, N333, N5237);
not NOT1 (N12766, N12762);
and AND3 (N12767, N12757, N6201, N10839);
xor XOR2 (N12768, N12765, N11199);
xor XOR2 (N12769, N12767, N8865);
nand NAND2 (N12770, N12759, N1321);
and AND2 (N12771, N12764, N3294);
buf BUF1 (N12772, N12771);
nor NOR3 (N12773, N12760, N11970, N2226);
buf BUF1 (N12774, N12751);
xor XOR2 (N12775, N12772, N2715);
xor XOR2 (N12776, N12766, N11905);
buf BUF1 (N12777, N12763);
not NOT1 (N12778, N12769);
and AND4 (N12779, N12773, N10648, N9026, N11047);
buf BUF1 (N12780, N12761);
buf BUF1 (N12781, N12770);
xor XOR2 (N12782, N12778, N11666);
xor XOR2 (N12783, N12756, N4198);
and AND3 (N12784, N12775, N4489, N6618);
or OR4 (N12785, N12784, N7724, N11116, N2085);
nor NOR3 (N12786, N12783, N7141, N2952);
xor XOR2 (N12787, N12785, N2784);
and AND2 (N12788, N12787, N431);
xor XOR2 (N12789, N12779, N10514);
nor NOR2 (N12790, N12768, N6841);
nand NAND2 (N12791, N12782, N10355);
nor NOR3 (N12792, N12789, N5600, N4951);
buf BUF1 (N12793, N12776);
or OR3 (N12794, N12780, N10858, N7160);
not NOT1 (N12795, N12790);
buf BUF1 (N12796, N12795);
and AND3 (N12797, N12774, N8581, N2282);
nor NOR2 (N12798, N12793, N2457);
nor NOR3 (N12799, N12796, N5243, N10738);
xor XOR2 (N12800, N12786, N1400);
or OR4 (N12801, N12794, N8617, N9660, N11696);
not NOT1 (N12802, N12800);
not NOT1 (N12803, N12791);
or OR3 (N12804, N12781, N8167, N8844);
xor XOR2 (N12805, N12792, N12113);
not NOT1 (N12806, N12777);
nor NOR4 (N12807, N12797, N11496, N12760, N7050);
or OR2 (N12808, N12806, N6162);
xor XOR2 (N12809, N12807, N11419);
buf BUF1 (N12810, N12805);
and AND4 (N12811, N12810, N3889, N6426, N8037);
nor NOR3 (N12812, N12798, N6325, N6181);
or OR3 (N12813, N12811, N8693, N9553);
nand NAND2 (N12814, N12788, N10715);
and AND4 (N12815, N12804, N8208, N9341, N2502);
xor XOR2 (N12816, N12814, N946);
nor NOR3 (N12817, N12816, N6118, N6855);
not NOT1 (N12818, N12813);
buf BUF1 (N12819, N12812);
or OR4 (N12820, N12803, N3354, N11140, N4008);
nor NOR2 (N12821, N12808, N4135);
nor NOR2 (N12822, N12818, N4679);
not NOT1 (N12823, N12815);
xor XOR2 (N12824, N12820, N1777);
nand NAND2 (N12825, N12817, N975);
buf BUF1 (N12826, N12825);
nand NAND3 (N12827, N12823, N9407, N4992);
xor XOR2 (N12828, N12799, N6410);
nor NOR2 (N12829, N12809, N10538);
buf BUF1 (N12830, N12826);
not NOT1 (N12831, N12801);
xor XOR2 (N12832, N12828, N1016);
nand NAND3 (N12833, N12832, N185, N3746);
and AND4 (N12834, N12822, N4611, N4692, N4483);
buf BUF1 (N12835, N12830);
or OR4 (N12836, N12835, N12675, N3086, N4554);
nor NOR3 (N12837, N12834, N2999, N12497);
and AND2 (N12838, N12837, N469);
nor NOR3 (N12839, N12831, N11075, N11504);
xor XOR2 (N12840, N12839, N11460);
buf BUF1 (N12841, N12827);
nand NAND4 (N12842, N12840, N4745, N7719, N10829);
or OR3 (N12843, N12819, N9519, N12077);
or OR3 (N12844, N12829, N10748, N3491);
nand NAND4 (N12845, N12844, N10278, N2794, N8488);
not NOT1 (N12846, N12821);
not NOT1 (N12847, N12841);
nand NAND4 (N12848, N12842, N8592, N11948, N2044);
or OR4 (N12849, N12847, N5692, N6990, N7324);
nand NAND2 (N12850, N12846, N11686);
nand NAND2 (N12851, N12848, N10834);
and AND2 (N12852, N12845, N10514);
nor NOR3 (N12853, N12851, N3876, N12529);
or OR4 (N12854, N12836, N9423, N10420, N3352);
xor XOR2 (N12855, N12824, N1866);
xor XOR2 (N12856, N12853, N12664);
nor NOR3 (N12857, N12855, N11971, N8235);
or OR4 (N12858, N12857, N5686, N10289, N7594);
xor XOR2 (N12859, N12852, N330);
nand NAND3 (N12860, N12843, N7252, N5190);
buf BUF1 (N12861, N12860);
xor XOR2 (N12862, N12833, N5841);
nand NAND4 (N12863, N12802, N4934, N10775, N5850);
not NOT1 (N12864, N12863);
not NOT1 (N12865, N12854);
buf BUF1 (N12866, N12865);
and AND4 (N12867, N12866, N10743, N10374, N2794);
nor NOR2 (N12868, N12867, N3544);
buf BUF1 (N12869, N12862);
and AND3 (N12870, N12856, N12688, N12462);
xor XOR2 (N12871, N12859, N8470);
buf BUF1 (N12872, N12871);
nand NAND2 (N12873, N12869, N10137);
xor XOR2 (N12874, N12868, N10203);
buf BUF1 (N12875, N12872);
xor XOR2 (N12876, N12838, N8474);
not NOT1 (N12877, N12864);
nor NOR3 (N12878, N12874, N6818, N4663);
or OR2 (N12879, N12875, N981);
nor NOR4 (N12880, N12858, N3043, N6802, N12577);
nor NOR4 (N12881, N12880, N1371, N2825, N487);
or OR4 (N12882, N12878, N1608, N4840, N85);
nand NAND2 (N12883, N12879, N10192);
buf BUF1 (N12884, N12883);
not NOT1 (N12885, N12876);
not NOT1 (N12886, N12884);
nor NOR2 (N12887, N12861, N2074);
nand NAND3 (N12888, N12882, N6477, N6561);
xor XOR2 (N12889, N12870, N5915);
not NOT1 (N12890, N12849);
nor NOR4 (N12891, N12850, N6070, N2083, N3816);
xor XOR2 (N12892, N12881, N8473);
xor XOR2 (N12893, N12873, N5147);
xor XOR2 (N12894, N12887, N677);
and AND4 (N12895, N12885, N8160, N6422, N10664);
nand NAND4 (N12896, N12890, N1667, N10395, N5002);
nand NAND3 (N12897, N12889, N8132, N6212);
nand NAND4 (N12898, N12897, N8205, N10764, N12078);
buf BUF1 (N12899, N12886);
buf BUF1 (N12900, N12898);
not NOT1 (N12901, N12896);
and AND2 (N12902, N12891, N12348);
nor NOR4 (N12903, N12895, N534, N5483, N3314);
xor XOR2 (N12904, N12877, N5473);
buf BUF1 (N12905, N12901);
nor NOR2 (N12906, N12894, N8663);
nor NOR4 (N12907, N12902, N11943, N3066, N11541);
and AND4 (N12908, N12899, N12103, N9324, N7048);
and AND4 (N12909, N12907, N4366, N6303, N316);
nor NOR3 (N12910, N12905, N11750, N4972);
and AND2 (N12911, N12893, N12893);
and AND4 (N12912, N12888, N3487, N2121, N5973);
buf BUF1 (N12913, N12910);
buf BUF1 (N12914, N12904);
or OR4 (N12915, N12911, N746, N10673, N12629);
and AND2 (N12916, N12900, N5578);
buf BUF1 (N12917, N12915);
not NOT1 (N12918, N12892);
or OR2 (N12919, N12918, N8594);
nor NOR2 (N12920, N12916, N1820);
or OR2 (N12921, N12913, N679);
not NOT1 (N12922, N12919);
xor XOR2 (N12923, N12903, N7368);
nand NAND4 (N12924, N12906, N6521, N12792, N3831);
and AND4 (N12925, N12914, N11377, N2539, N6841);
xor XOR2 (N12926, N12920, N7046);
or OR3 (N12927, N12924, N11839, N9839);
or OR2 (N12928, N12912, N1061);
or OR3 (N12929, N12926, N5907, N10730);
xor XOR2 (N12930, N12929, N5812);
nand NAND3 (N12931, N12917, N6718, N4894);
nand NAND3 (N12932, N12923, N5691, N10400);
nand NAND3 (N12933, N12921, N11455, N5400);
nand NAND4 (N12934, N12908, N11074, N270, N11419);
nand NAND2 (N12935, N12928, N7452);
and AND3 (N12936, N12935, N12789, N122);
buf BUF1 (N12937, N12927);
not NOT1 (N12938, N12932);
buf BUF1 (N12939, N12925);
nand NAND4 (N12940, N12939, N11056, N8329, N11468);
not NOT1 (N12941, N12931);
nand NAND2 (N12942, N12941, N4145);
buf BUF1 (N12943, N12909);
buf BUF1 (N12944, N12943);
xor XOR2 (N12945, N12942, N3239);
nand NAND3 (N12946, N12937, N10606, N6392);
xor XOR2 (N12947, N12940, N6784);
nor NOR3 (N12948, N12922, N4493, N5519);
buf BUF1 (N12949, N12930);
xor XOR2 (N12950, N12934, N8685);
or OR2 (N12951, N12944, N1814);
and AND4 (N12952, N12938, N5435, N8532, N7829);
nor NOR3 (N12953, N12950, N11500, N1427);
or OR3 (N12954, N12936, N6410, N10189);
buf BUF1 (N12955, N12949);
or OR4 (N12956, N12954, N5292, N3534, N9515);
nor NOR3 (N12957, N12947, N4022, N5468);
nand NAND4 (N12958, N12955, N6904, N10022, N3701);
or OR3 (N12959, N12945, N1005, N5430);
buf BUF1 (N12960, N12951);
buf BUF1 (N12961, N12960);
nand NAND3 (N12962, N12952, N8963, N4608);
nand NAND4 (N12963, N12946, N7578, N4381, N9068);
buf BUF1 (N12964, N12959);
nor NOR3 (N12965, N12958, N8566, N6847);
nand NAND4 (N12966, N12962, N6330, N4861, N4837);
xor XOR2 (N12967, N12963, N11151);
buf BUF1 (N12968, N12961);
not NOT1 (N12969, N12964);
and AND4 (N12970, N12956, N9365, N12869, N125);
buf BUF1 (N12971, N12969);
buf BUF1 (N12972, N12948);
nand NAND2 (N12973, N12968, N9809);
nand NAND2 (N12974, N12966, N12234);
xor XOR2 (N12975, N12957, N11472);
buf BUF1 (N12976, N12953);
or OR4 (N12977, N12967, N6759, N2106, N10878);
xor XOR2 (N12978, N12933, N1026);
nor NOR4 (N12979, N12971, N1004, N7991, N2043);
not NOT1 (N12980, N12972);
buf BUF1 (N12981, N12974);
not NOT1 (N12982, N12979);
and AND2 (N12983, N12977, N10350);
not NOT1 (N12984, N12975);
and AND4 (N12985, N12983, N1180, N1070, N6244);
buf BUF1 (N12986, N12980);
not NOT1 (N12987, N12965);
nor NOR2 (N12988, N12976, N7489);
nand NAND3 (N12989, N12970, N2691, N3688);
buf BUF1 (N12990, N12986);
xor XOR2 (N12991, N12989, N6689);
nor NOR2 (N12992, N12981, N7719);
buf BUF1 (N12993, N12973);
and AND2 (N12994, N12982, N1546);
or OR2 (N12995, N12993, N8569);
nand NAND2 (N12996, N12995, N7576);
or OR4 (N12997, N12991, N3684, N12643, N6513);
xor XOR2 (N12998, N12992, N7308);
xor XOR2 (N12999, N12978, N11036);
or OR2 (N13000, N12984, N11627);
or OR3 (N13001, N12994, N8148, N8665);
xor XOR2 (N13002, N12999, N3144);
or OR3 (N13003, N12996, N8702, N9700);
or OR2 (N13004, N12988, N1648);
or OR4 (N13005, N13000, N407, N8516, N2041);
not NOT1 (N13006, N13003);
nand NAND2 (N13007, N12998, N6977);
or OR2 (N13008, N12987, N460);
nand NAND4 (N13009, N13007, N6556, N7450, N3675);
not NOT1 (N13010, N12990);
or OR3 (N13011, N13006, N2121, N10051);
nand NAND2 (N13012, N13002, N2231);
nand NAND3 (N13013, N13005, N10310, N5119);
and AND2 (N13014, N13001, N10007);
and AND4 (N13015, N12985, N12825, N2875, N2501);
or OR3 (N13016, N13015, N2986, N7156);
nand NAND3 (N13017, N13013, N4299, N6454);
nor NOR4 (N13018, N12997, N5748, N2088, N1076);
buf BUF1 (N13019, N13009);
not NOT1 (N13020, N13004);
xor XOR2 (N13021, N13008, N11995);
nand NAND2 (N13022, N13011, N11599);
or OR3 (N13023, N13014, N1809, N3841);
buf BUF1 (N13024, N13022);
or OR3 (N13025, N13020, N12952, N4377);
nand NAND2 (N13026, N13019, N8455);
nor NOR4 (N13027, N13025, N2101, N861, N1766);
nor NOR3 (N13028, N13012, N10074, N8309);
not NOT1 (N13029, N13024);
or OR4 (N13030, N13016, N3556, N8763, N1745);
nand NAND2 (N13031, N13018, N5844);
xor XOR2 (N13032, N13030, N5199);
nor NOR3 (N13033, N13029, N3818, N1399);
buf BUF1 (N13034, N13021);
and AND4 (N13035, N13028, N11583, N6563, N5173);
or OR2 (N13036, N13033, N7080);
not NOT1 (N13037, N13010);
or OR2 (N13038, N13027, N5136);
xor XOR2 (N13039, N13031, N8416);
or OR2 (N13040, N13023, N7924);
nand NAND2 (N13041, N13017, N5);
buf BUF1 (N13042, N13026);
and AND4 (N13043, N13036, N2800, N5401, N8819);
and AND2 (N13044, N13039, N4202);
buf BUF1 (N13045, N13038);
and AND4 (N13046, N13032, N12395, N9513, N10736);
not NOT1 (N13047, N13034);
and AND2 (N13048, N13042, N4080);
buf BUF1 (N13049, N13044);
not NOT1 (N13050, N13035);
and AND2 (N13051, N13050, N2219);
buf BUF1 (N13052, N13037);
or OR3 (N13053, N13043, N2006, N10385);
or OR3 (N13054, N13040, N6989, N7924);
and AND3 (N13055, N13049, N5665, N5600);
and AND4 (N13056, N13041, N9863, N11549, N12761);
buf BUF1 (N13057, N13048);
not NOT1 (N13058, N13056);
nand NAND3 (N13059, N13057, N13034, N2898);
and AND4 (N13060, N13054, N5332, N355, N2206);
xor XOR2 (N13061, N13055, N12409);
xor XOR2 (N13062, N13052, N4676);
xor XOR2 (N13063, N13058, N8235);
buf BUF1 (N13064, N13060);
or OR3 (N13065, N13062, N7819, N880);
nor NOR4 (N13066, N13051, N2240, N5949, N3947);
nand NAND2 (N13067, N13045, N5962);
xor XOR2 (N13068, N13065, N8278);
or OR3 (N13069, N13067, N10707, N869);
nor NOR3 (N13070, N13069, N5298, N9324);
or OR4 (N13071, N13046, N2256, N9467, N8605);
nor NOR3 (N13072, N13064, N8846, N6807);
xor XOR2 (N13073, N13047, N2110);
or OR2 (N13074, N13053, N8442);
or OR2 (N13075, N13070, N11676);
nand NAND3 (N13076, N13074, N11857, N575);
or OR2 (N13077, N13063, N706);
nor NOR4 (N13078, N13075, N371, N7474, N4646);
nor NOR4 (N13079, N13078, N1102, N3741, N12087);
and AND2 (N13080, N13076, N10617);
nand NAND4 (N13081, N13059, N153, N7765, N5232);
or OR2 (N13082, N13066, N12445);
nor NOR2 (N13083, N13068, N8487);
xor XOR2 (N13084, N13061, N5339);
not NOT1 (N13085, N13080);
and AND2 (N13086, N13082, N10235);
nand NAND4 (N13087, N13079, N6014, N8790, N1544);
nand NAND4 (N13088, N13086, N9382, N11757, N7297);
nor NOR3 (N13089, N13083, N11681, N6142);
not NOT1 (N13090, N13089);
or OR2 (N13091, N13081, N699);
or OR3 (N13092, N13072, N9578, N3580);
buf BUF1 (N13093, N13087);
not NOT1 (N13094, N13084);
buf BUF1 (N13095, N13091);
or OR2 (N13096, N13095, N8639);
buf BUF1 (N13097, N13077);
nor NOR4 (N13098, N13096, N12046, N7527, N11207);
or OR2 (N13099, N13097, N1187);
nor NOR4 (N13100, N13090, N2769, N1756, N9252);
and AND3 (N13101, N13073, N748, N10294);
or OR4 (N13102, N13094, N1728, N12022, N11530);
not NOT1 (N13103, N13085);
or OR3 (N13104, N13099, N5267, N8665);
nand NAND2 (N13105, N13100, N5997);
or OR2 (N13106, N13101, N4606);
or OR3 (N13107, N13105, N1276, N11574);
nor NOR4 (N13108, N13103, N9661, N5730, N9664);
nand NAND4 (N13109, N13098, N10956, N2561, N1422);
buf BUF1 (N13110, N13108);
nor NOR3 (N13111, N13093, N3896, N1031);
nand NAND2 (N13112, N13111, N3341);
and AND4 (N13113, N13112, N4486, N4501, N869);
nor NOR3 (N13114, N13088, N11699, N12317);
nand NAND3 (N13115, N13102, N4109, N6560);
nor NOR3 (N13116, N13107, N12800, N10255);
nand NAND4 (N13117, N13106, N11812, N9858, N1363);
or OR3 (N13118, N13117, N3980, N4173);
buf BUF1 (N13119, N13114);
nand NAND3 (N13120, N13071, N959, N2189);
or OR2 (N13121, N13113, N1291);
buf BUF1 (N13122, N13119);
not NOT1 (N13123, N13120);
nand NAND2 (N13124, N13104, N8856);
or OR4 (N13125, N13092, N11929, N9233, N8486);
xor XOR2 (N13126, N13116, N12817);
buf BUF1 (N13127, N13115);
xor XOR2 (N13128, N13110, N11959);
nor NOR4 (N13129, N13118, N5509, N10165, N3498);
buf BUF1 (N13130, N13128);
nor NOR4 (N13131, N13129, N10605, N6637, N9636);
xor XOR2 (N13132, N13130, N7559);
or OR3 (N13133, N13109, N870, N5607);
nand NAND4 (N13134, N13123, N9153, N12180, N708);
nand NAND3 (N13135, N13134, N7455, N11803);
or OR4 (N13136, N13125, N9802, N11461, N9995);
xor XOR2 (N13137, N13135, N11814);
or OR4 (N13138, N13133, N12901, N9893, N4619);
not NOT1 (N13139, N13138);
nor NOR4 (N13140, N13136, N8655, N11846, N11620);
and AND4 (N13141, N13122, N2528, N12893, N1622);
and AND2 (N13142, N13140, N10149);
nor NOR2 (N13143, N13127, N580);
and AND3 (N13144, N13142, N9965, N10601);
nor NOR4 (N13145, N13141, N1437, N5688, N11318);
buf BUF1 (N13146, N13139);
xor XOR2 (N13147, N13126, N6136);
buf BUF1 (N13148, N13144);
xor XOR2 (N13149, N13148, N10645);
not NOT1 (N13150, N13124);
buf BUF1 (N13151, N13143);
not NOT1 (N13152, N13131);
or OR2 (N13153, N13137, N12004);
xor XOR2 (N13154, N13145, N11900);
nand NAND3 (N13155, N13121, N11901, N10943);
and AND4 (N13156, N13153, N435, N967, N7950);
not NOT1 (N13157, N13150);
or OR4 (N13158, N13151, N451, N9536, N9547);
nor NOR4 (N13159, N13156, N11305, N4304, N406);
not NOT1 (N13160, N13154);
nor NOR2 (N13161, N13160, N7525);
and AND4 (N13162, N13155, N11360, N6075, N10625);
xor XOR2 (N13163, N13161, N4437);
nor NOR3 (N13164, N13162, N6881, N2089);
xor XOR2 (N13165, N13158, N1996);
nor NOR3 (N13166, N13152, N4058, N12105);
not NOT1 (N13167, N13157);
not NOT1 (N13168, N13147);
not NOT1 (N13169, N13165);
xor XOR2 (N13170, N13167, N8633);
xor XOR2 (N13171, N13170, N10509);
xor XOR2 (N13172, N13171, N7394);
not NOT1 (N13173, N13166);
nor NOR2 (N13174, N13163, N7424);
and AND4 (N13175, N13164, N13167, N6046, N7817);
and AND4 (N13176, N13132, N11601, N6609, N3415);
or OR4 (N13177, N13174, N2106, N12725, N10331);
or OR4 (N13178, N13176, N6695, N6851, N2997);
nor NOR4 (N13179, N13149, N8097, N9009, N9895);
not NOT1 (N13180, N13168);
nor NOR4 (N13181, N13173, N1845, N3881, N7981);
nor NOR4 (N13182, N13172, N10523, N5778, N2730);
not NOT1 (N13183, N13175);
not NOT1 (N13184, N13183);
and AND2 (N13185, N13169, N10284);
nor NOR4 (N13186, N13185, N12985, N8645, N4698);
buf BUF1 (N13187, N13159);
buf BUF1 (N13188, N13184);
nor NOR2 (N13189, N13181, N5581);
nand NAND4 (N13190, N13182, N7613, N13120, N5350);
and AND2 (N13191, N13186, N6932);
xor XOR2 (N13192, N13187, N8285);
nand NAND2 (N13193, N13146, N1663);
or OR3 (N13194, N13179, N8186, N8074);
or OR3 (N13195, N13189, N2563, N1464);
xor XOR2 (N13196, N13192, N12187);
nand NAND3 (N13197, N13191, N9161, N6876);
buf BUF1 (N13198, N13188);
buf BUF1 (N13199, N13195);
xor XOR2 (N13200, N13180, N2471);
and AND3 (N13201, N13200, N8349, N7339);
and AND2 (N13202, N13198, N4559);
nand NAND2 (N13203, N13201, N12195);
buf BUF1 (N13204, N13203);
not NOT1 (N13205, N13177);
nor NOR2 (N13206, N13196, N8141);
or OR3 (N13207, N13206, N1408, N6008);
buf BUF1 (N13208, N13202);
nand NAND4 (N13209, N13207, N7525, N1386, N556);
and AND4 (N13210, N13204, N8021, N11943, N8245);
or OR3 (N13211, N13190, N3640, N11399);
and AND2 (N13212, N13209, N925);
nand NAND3 (N13213, N13205, N13144, N10684);
or OR4 (N13214, N13199, N7676, N12807, N10130);
buf BUF1 (N13215, N13193);
or OR4 (N13216, N13211, N4595, N8423, N9014);
nor NOR4 (N13217, N13210, N10090, N10120, N5555);
and AND2 (N13218, N13216, N6808);
and AND4 (N13219, N13213, N9861, N1213, N12431);
nor NOR3 (N13220, N13217, N2858, N3902);
buf BUF1 (N13221, N13208);
xor XOR2 (N13222, N13178, N850);
not NOT1 (N13223, N13219);
nor NOR3 (N13224, N13215, N5278, N3697);
buf BUF1 (N13225, N13194);
or OR2 (N13226, N13220, N3491);
or OR3 (N13227, N13218, N7112, N3549);
nand NAND4 (N13228, N13221, N11724, N10353, N8205);
xor XOR2 (N13229, N13197, N4442);
not NOT1 (N13230, N13214);
or OR4 (N13231, N13212, N4059, N7999, N5105);
buf BUF1 (N13232, N13230);
buf BUF1 (N13233, N13229);
not NOT1 (N13234, N13225);
xor XOR2 (N13235, N13228, N12438);
not NOT1 (N13236, N13231);
buf BUF1 (N13237, N13235);
or OR2 (N13238, N13236, N12454);
not NOT1 (N13239, N13226);
buf BUF1 (N13240, N13234);
xor XOR2 (N13241, N13227, N13148);
xor XOR2 (N13242, N13232, N7297);
nand NAND3 (N13243, N13233, N4687, N3136);
nand NAND3 (N13244, N13237, N8455, N12612);
xor XOR2 (N13245, N13238, N63);
nor NOR4 (N13246, N13243, N8011, N7759, N9265);
nor NOR4 (N13247, N13245, N5220, N12262, N12309);
nand NAND3 (N13248, N13222, N540, N1321);
buf BUF1 (N13249, N13239);
not NOT1 (N13250, N13241);
xor XOR2 (N13251, N13223, N4995);
not NOT1 (N13252, N13247);
xor XOR2 (N13253, N13242, N1841);
nand NAND4 (N13254, N13253, N10920, N13130, N9344);
and AND4 (N13255, N13249, N3564, N5952, N6372);
xor XOR2 (N13256, N13224, N4266);
not NOT1 (N13257, N13256);
nor NOR3 (N13258, N13244, N1456, N10814);
and AND3 (N13259, N13251, N2593, N4833);
and AND2 (N13260, N13240, N9971);
nand NAND4 (N13261, N13248, N6687, N10090, N1609);
not NOT1 (N13262, N13260);
and AND4 (N13263, N13255, N9084, N11279, N10891);
nand NAND3 (N13264, N13259, N5098, N8834);
and AND3 (N13265, N13261, N3695, N9743);
nor NOR4 (N13266, N13250, N12827, N2290, N6834);
buf BUF1 (N13267, N13254);
xor XOR2 (N13268, N13266, N4223);
and AND3 (N13269, N13264, N4311, N9366);
buf BUF1 (N13270, N13258);
nand NAND2 (N13271, N13270, N6200);
nand NAND2 (N13272, N13268, N8675);
nor NOR2 (N13273, N13262, N9072);
not NOT1 (N13274, N13265);
not NOT1 (N13275, N13273);
buf BUF1 (N13276, N13275);
xor XOR2 (N13277, N13274, N3060);
and AND4 (N13278, N13252, N12134, N10719, N13142);
nand NAND2 (N13279, N13276, N10852);
xor XOR2 (N13280, N13278, N9188);
xor XOR2 (N13281, N13280, N8831);
not NOT1 (N13282, N13263);
buf BUF1 (N13283, N13281);
not NOT1 (N13284, N13279);
not NOT1 (N13285, N13257);
or OR2 (N13286, N13283, N5046);
nor NOR3 (N13287, N13286, N3918, N4544);
and AND2 (N13288, N13284, N6404);
xor XOR2 (N13289, N13285, N8377);
and AND2 (N13290, N13269, N7633);
or OR4 (N13291, N13277, N1473, N4054, N12402);
xor XOR2 (N13292, N13246, N1031);
or OR3 (N13293, N13271, N12714, N7493);
not NOT1 (N13294, N13287);
not NOT1 (N13295, N13282);
nand NAND4 (N13296, N13293, N9765, N8673, N8215);
buf BUF1 (N13297, N13289);
buf BUF1 (N13298, N13288);
nand NAND3 (N13299, N13295, N8824, N1683);
or OR3 (N13300, N13299, N11761, N13185);
nor NOR3 (N13301, N13291, N7342, N4362);
xor XOR2 (N13302, N13297, N5827);
buf BUF1 (N13303, N13267);
nand NAND4 (N13304, N13292, N7629, N5501, N13203);
or OR4 (N13305, N13302, N12739, N3835, N5764);
buf BUF1 (N13306, N13303);
nand NAND2 (N13307, N13304, N1002);
xor XOR2 (N13308, N13298, N934);
xor XOR2 (N13309, N13296, N11291);
xor XOR2 (N13310, N13307, N5197);
xor XOR2 (N13311, N13305, N5309);
nor NOR4 (N13312, N13308, N7173, N9035, N2199);
not NOT1 (N13313, N13306);
and AND3 (N13314, N13311, N8411, N10714);
and AND3 (N13315, N13310, N10914, N2291);
nand NAND2 (N13316, N13313, N609);
buf BUF1 (N13317, N13314);
buf BUF1 (N13318, N13312);
not NOT1 (N13319, N13294);
buf BUF1 (N13320, N13318);
and AND2 (N13321, N13272, N10869);
not NOT1 (N13322, N13319);
or OR4 (N13323, N13320, N3958, N8623, N11686);
nand NAND2 (N13324, N13316, N3824);
xor XOR2 (N13325, N13301, N6243);
or OR3 (N13326, N13325, N7648, N3173);
nor NOR3 (N13327, N13300, N6328, N3623);
nand NAND2 (N13328, N13290, N649);
nor NOR2 (N13329, N13315, N185);
or OR4 (N13330, N13329, N847, N168, N6882);
buf BUF1 (N13331, N13326);
nor NOR2 (N13332, N13321, N9079);
or OR2 (N13333, N13330, N8050);
nor NOR4 (N13334, N13331, N610, N8214, N9210);
not NOT1 (N13335, N13333);
buf BUF1 (N13336, N13309);
nor NOR2 (N13337, N13335, N5702);
and AND2 (N13338, N13327, N9251);
not NOT1 (N13339, N13332);
nand NAND2 (N13340, N13328, N885);
nand NAND4 (N13341, N13334, N8254, N4349, N4734);
nand NAND2 (N13342, N13339, N361);
or OR4 (N13343, N13324, N3219, N3796, N7747);
or OR2 (N13344, N13337, N7913);
and AND4 (N13345, N13336, N10352, N3770, N4912);
xor XOR2 (N13346, N13342, N2823);
buf BUF1 (N13347, N13340);
or OR4 (N13348, N13346, N5976, N2048, N4521);
or OR3 (N13349, N13338, N8082, N8372);
buf BUF1 (N13350, N13349);
not NOT1 (N13351, N13317);
and AND3 (N13352, N13351, N11597, N10049);
not NOT1 (N13353, N13350);
or OR2 (N13354, N13343, N10360);
or OR3 (N13355, N13347, N12949, N8420);
buf BUF1 (N13356, N13341);
not NOT1 (N13357, N13352);
buf BUF1 (N13358, N13354);
nor NOR4 (N13359, N13345, N2207, N8853, N1288);
and AND3 (N13360, N13322, N1391, N2398);
not NOT1 (N13361, N13360);
nor NOR3 (N13362, N13353, N10982, N11060);
and AND2 (N13363, N13356, N4437);
or OR4 (N13364, N13357, N3223, N4060, N4136);
and AND3 (N13365, N13323, N4741, N7602);
nor NOR2 (N13366, N13359, N5751);
and AND4 (N13367, N13348, N7531, N7472, N1218);
not NOT1 (N13368, N13367);
not NOT1 (N13369, N13361);
nor NOR3 (N13370, N13358, N6870, N1438);
nand NAND4 (N13371, N13366, N10587, N8576, N4817);
not NOT1 (N13372, N13369);
and AND4 (N13373, N13363, N5206, N6462, N13193);
not NOT1 (N13374, N13373);
nor NOR4 (N13375, N13371, N2305, N8605, N3545);
xor XOR2 (N13376, N13374, N6567);
and AND4 (N13377, N13376, N2391, N569, N1291);
and AND3 (N13378, N13362, N11735, N10879);
and AND2 (N13379, N13370, N835);
not NOT1 (N13380, N13355);
and AND3 (N13381, N13380, N8433, N8102);
or OR3 (N13382, N13372, N5125, N10738);
xor XOR2 (N13383, N13364, N8588);
nor NOR4 (N13384, N13375, N8070, N286, N11008);
nand NAND2 (N13385, N13384, N1996);
nor NOR4 (N13386, N13379, N13271, N838, N3234);
and AND4 (N13387, N13382, N2153, N5601, N1432);
and AND3 (N13388, N13383, N7259, N9530);
xor XOR2 (N13389, N13388, N3635);
nor NOR4 (N13390, N13389, N3727, N12890, N10428);
or OR2 (N13391, N13381, N9325);
xor XOR2 (N13392, N13368, N11353);
nor NOR2 (N13393, N13390, N401);
xor XOR2 (N13394, N13391, N12154);
or OR4 (N13395, N13393, N6984, N5941, N9079);
or OR2 (N13396, N13377, N603);
or OR3 (N13397, N13392, N5490, N9715);
buf BUF1 (N13398, N13396);
xor XOR2 (N13399, N13365, N4376);
not NOT1 (N13400, N13387);
buf BUF1 (N13401, N13395);
and AND3 (N13402, N13397, N1077, N1507);
nand NAND3 (N13403, N13399, N2028, N8880);
nand NAND2 (N13404, N13385, N10225);
or OR4 (N13405, N13404, N8164, N983, N2335);
or OR4 (N13406, N13344, N3491, N9567, N9086);
xor XOR2 (N13407, N13405, N4392);
not NOT1 (N13408, N13406);
nand NAND2 (N13409, N13378, N7478);
not NOT1 (N13410, N13408);
and AND3 (N13411, N13386, N5287, N2787);
buf BUF1 (N13412, N13411);
nand NAND3 (N13413, N13394, N8582, N5411);
or OR4 (N13414, N13401, N11389, N2772, N6307);
or OR3 (N13415, N13403, N4967, N5758);
or OR3 (N13416, N13409, N11833, N1990);
not NOT1 (N13417, N13410);
or OR3 (N13418, N13398, N7441, N2007);
or OR2 (N13419, N13417, N12991);
not NOT1 (N13420, N13418);
nor NOR2 (N13421, N13412, N5587);
buf BUF1 (N13422, N13421);
not NOT1 (N13423, N13415);
and AND3 (N13424, N13416, N3028, N4275);
not NOT1 (N13425, N13402);
nor NOR3 (N13426, N13423, N3413, N10536);
buf BUF1 (N13427, N13424);
not NOT1 (N13428, N13419);
not NOT1 (N13429, N13413);
or OR2 (N13430, N13427, N2515);
and AND3 (N13431, N13426, N2059, N10168);
nor NOR3 (N13432, N13430, N5141, N8077);
nor NOR4 (N13433, N13432, N7894, N3540, N11519);
nor NOR4 (N13434, N13425, N12545, N9079, N4029);
nand NAND3 (N13435, N13422, N6640, N8618);
and AND3 (N13436, N13435, N240, N5352);
and AND2 (N13437, N13414, N9244);
nand NAND2 (N13438, N13428, N7246);
buf BUF1 (N13439, N13400);
nand NAND4 (N13440, N13436, N11244, N712, N9151);
or OR3 (N13441, N13439, N10623, N5055);
not NOT1 (N13442, N13437);
nor NOR4 (N13443, N13433, N13346, N337, N11502);
or OR4 (N13444, N13442, N4428, N6468, N8307);
nor NOR4 (N13445, N13434, N515, N13358, N10921);
not NOT1 (N13446, N13431);
and AND4 (N13447, N13420, N12177, N6826, N230);
xor XOR2 (N13448, N13447, N630);
and AND2 (N13449, N13440, N13335);
nand NAND3 (N13450, N13429, N2162, N3663);
not NOT1 (N13451, N13441);
and AND3 (N13452, N13438, N11663, N319);
or OR2 (N13453, N13448, N10292);
not NOT1 (N13454, N13449);
not NOT1 (N13455, N13444);
or OR4 (N13456, N13407, N7348, N4536, N1485);
or OR2 (N13457, N13445, N7320);
nand NAND2 (N13458, N13446, N6576);
buf BUF1 (N13459, N13457);
xor XOR2 (N13460, N13454, N2718);
not NOT1 (N13461, N13443);
nor NOR2 (N13462, N13456, N9006);
or OR4 (N13463, N13455, N5754, N1358, N8397);
or OR2 (N13464, N13463, N2925);
buf BUF1 (N13465, N13458);
xor XOR2 (N13466, N13461, N13038);
nand NAND4 (N13467, N13453, N8610, N2916, N3914);
and AND3 (N13468, N13452, N8719, N5545);
nand NAND2 (N13469, N13466, N1051);
nor NOR4 (N13470, N13459, N1901, N823, N2982);
xor XOR2 (N13471, N13465, N6221);
xor XOR2 (N13472, N13468, N8800);
nand NAND3 (N13473, N13462, N1636, N11914);
and AND2 (N13474, N13467, N6480);
xor XOR2 (N13475, N13451, N1417);
nand NAND3 (N13476, N13475, N12626, N789);
not NOT1 (N13477, N13464);
buf BUF1 (N13478, N13473);
nand NAND4 (N13479, N13469, N3488, N4895, N8795);
or OR4 (N13480, N13470, N10636, N2797, N7450);
not NOT1 (N13481, N13460);
xor XOR2 (N13482, N13478, N11701);
and AND2 (N13483, N13477, N12612);
or OR2 (N13484, N13482, N9982);
xor XOR2 (N13485, N13450, N3906);
not NOT1 (N13486, N13479);
buf BUF1 (N13487, N13474);
nand NAND3 (N13488, N13480, N4541, N6520);
nor NOR3 (N13489, N13471, N1462, N8319);
nand NAND3 (N13490, N13483, N4782, N8880);
buf BUF1 (N13491, N13476);
nand NAND4 (N13492, N13486, N1292, N12978, N6542);
not NOT1 (N13493, N13485);
and AND3 (N13494, N13492, N5249, N3522);
nand NAND2 (N13495, N13487, N4614);
and AND4 (N13496, N13493, N13128, N5577, N4015);
xor XOR2 (N13497, N13488, N1263);
and AND4 (N13498, N13494, N7, N4459, N2371);
xor XOR2 (N13499, N13495, N1466);
not NOT1 (N13500, N13490);
nand NAND3 (N13501, N13497, N10797, N5630);
and AND4 (N13502, N13484, N977, N7391, N2377);
not NOT1 (N13503, N13500);
xor XOR2 (N13504, N13489, N7613);
nor NOR3 (N13505, N13472, N8458, N11463);
nor NOR2 (N13506, N13496, N3);
buf BUF1 (N13507, N13491);
nor NOR4 (N13508, N13503, N7764, N13285, N11577);
buf BUF1 (N13509, N13506);
or OR4 (N13510, N13499, N89, N10944, N5977);
xor XOR2 (N13511, N13505, N2775);
xor XOR2 (N13512, N13507, N10587);
xor XOR2 (N13513, N13509, N10031);
and AND3 (N13514, N13498, N3460, N6737);
and AND2 (N13515, N13513, N6438);
nand NAND4 (N13516, N13501, N3374, N7598, N8158);
not NOT1 (N13517, N13514);
nand NAND4 (N13518, N13515, N2567, N184, N3888);
nand NAND2 (N13519, N13504, N12494);
xor XOR2 (N13520, N13518, N2511);
and AND4 (N13521, N13516, N5630, N7270, N9667);
and AND2 (N13522, N13502, N8578);
or OR3 (N13523, N13522, N4767, N9987);
nor NOR3 (N13524, N13517, N7273, N6412);
not NOT1 (N13525, N13508);
and AND3 (N13526, N13512, N2375, N4641);
nand NAND3 (N13527, N13481, N10048, N1255);
xor XOR2 (N13528, N13511, N7460);
xor XOR2 (N13529, N13528, N5051);
buf BUF1 (N13530, N13529);
buf BUF1 (N13531, N13524);
not NOT1 (N13532, N13523);
and AND2 (N13533, N13520, N9827);
and AND2 (N13534, N13526, N2012);
or OR3 (N13535, N13519, N9674, N10664);
xor XOR2 (N13536, N13525, N5369);
nor NOR2 (N13537, N13531, N7055);
not NOT1 (N13538, N13532);
buf BUF1 (N13539, N13534);
or OR4 (N13540, N13510, N11650, N3761, N984);
and AND2 (N13541, N13530, N3883);
nand NAND4 (N13542, N13538, N934, N7192, N3650);
nand NAND3 (N13543, N13539, N12617, N7173);
nand NAND2 (N13544, N13521, N7136);
or OR3 (N13545, N13541, N2718, N5607);
not NOT1 (N13546, N13543);
nand NAND3 (N13547, N13537, N11114, N6308);
or OR3 (N13548, N13544, N11786, N3146);
buf BUF1 (N13549, N13540);
nand NAND2 (N13550, N13533, N11596);
and AND3 (N13551, N13546, N743, N13349);
nor NOR4 (N13552, N13535, N7967, N7395, N11584);
not NOT1 (N13553, N13536);
nor NOR4 (N13554, N13553, N12829, N2268, N11485);
xor XOR2 (N13555, N13545, N4291);
not NOT1 (N13556, N13552);
buf BUF1 (N13557, N13527);
buf BUF1 (N13558, N13549);
nor NOR2 (N13559, N13554, N7690);
not NOT1 (N13560, N13555);
xor XOR2 (N13561, N13560, N607);
buf BUF1 (N13562, N13548);
not NOT1 (N13563, N13542);
or OR4 (N13564, N13556, N4111, N6938, N6423);
nand NAND2 (N13565, N13557, N3560);
or OR4 (N13566, N13551, N4706, N1910, N9971);
nand NAND4 (N13567, N13566, N5585, N2607, N4811);
nor NOR3 (N13568, N13561, N1582, N7053);
buf BUF1 (N13569, N13558);
or OR4 (N13570, N13564, N8927, N11268, N1938);
xor XOR2 (N13571, N13565, N9641);
nor NOR3 (N13572, N13569, N3810, N13539);
xor XOR2 (N13573, N13571, N10288);
nand NAND3 (N13574, N13572, N1533, N10160);
and AND3 (N13575, N13573, N6664, N1811);
and AND3 (N13576, N13562, N8256, N3314);
not NOT1 (N13577, N13550);
not NOT1 (N13578, N13577);
xor XOR2 (N13579, N13547, N9808);
buf BUF1 (N13580, N13567);
nand NAND4 (N13581, N13563, N7672, N2561, N9497);
or OR2 (N13582, N13568, N6999);
xor XOR2 (N13583, N13581, N6204);
xor XOR2 (N13584, N13580, N6337);
nor NOR4 (N13585, N13584, N3645, N3992, N11436);
nand NAND3 (N13586, N13559, N4023, N2139);
not NOT1 (N13587, N13583);
xor XOR2 (N13588, N13587, N7952);
xor XOR2 (N13589, N13576, N12218);
not NOT1 (N13590, N13575);
nand NAND4 (N13591, N13574, N4812, N8815, N1476);
nor NOR2 (N13592, N13582, N4964);
not NOT1 (N13593, N13585);
nor NOR3 (N13594, N13588, N6301, N11036);
nor NOR3 (N13595, N13592, N3993, N3147);
nor NOR4 (N13596, N13589, N3758, N7055, N1551);
and AND2 (N13597, N13578, N11648);
xor XOR2 (N13598, N13593, N3236);
nor NOR2 (N13599, N13598, N12099);
not NOT1 (N13600, N13570);
not NOT1 (N13601, N13594);
not NOT1 (N13602, N13595);
nand NAND3 (N13603, N13600, N6685, N7656);
nand NAND3 (N13604, N13599, N5067, N9211);
nor NOR4 (N13605, N13590, N4271, N8233, N4250);
or OR4 (N13606, N13602, N13323, N1243, N12218);
nand NAND4 (N13607, N13596, N878, N5982, N840);
and AND2 (N13608, N13597, N1727);
xor XOR2 (N13609, N13586, N7103);
buf BUF1 (N13610, N13604);
or OR4 (N13611, N13591, N7854, N10723, N4251);
not NOT1 (N13612, N13609);
and AND2 (N13613, N13606, N9523);
nor NOR2 (N13614, N13611, N8975);
or OR3 (N13615, N13605, N853, N2034);
buf BUF1 (N13616, N13613);
buf BUF1 (N13617, N13610);
nor NOR2 (N13618, N13608, N13184);
nor NOR3 (N13619, N13617, N1960, N5895);
not NOT1 (N13620, N13615);
nor NOR3 (N13621, N13579, N10745, N288);
nand NAND2 (N13622, N13619, N11754);
nand NAND3 (N13623, N13621, N9771, N13506);
nor NOR2 (N13624, N13618, N8757);
not NOT1 (N13625, N13620);
nor NOR2 (N13626, N13612, N9893);
and AND2 (N13627, N13603, N12178);
xor XOR2 (N13628, N13624, N12137);
and AND3 (N13629, N13622, N7958, N5027);
nand NAND4 (N13630, N13623, N2241, N5187, N7822);
nand NAND2 (N13631, N13616, N5417);
nand NAND2 (N13632, N13628, N11015);
not NOT1 (N13633, N13632);
buf BUF1 (N13634, N13630);
or OR4 (N13635, N13601, N8315, N10029, N12688);
buf BUF1 (N13636, N13614);
nor NOR2 (N13637, N13629, N8581);
buf BUF1 (N13638, N13607);
xor XOR2 (N13639, N13635, N6271);
nor NOR3 (N13640, N13639, N574, N8561);
and AND4 (N13641, N13636, N9054, N389, N6398);
and AND2 (N13642, N13626, N11576);
xor XOR2 (N13643, N13625, N4646);
or OR3 (N13644, N13641, N9039, N4129);
or OR2 (N13645, N13644, N8759);
buf BUF1 (N13646, N13645);
not NOT1 (N13647, N13633);
or OR2 (N13648, N13640, N9084);
or OR4 (N13649, N13638, N7408, N5120, N10465);
and AND3 (N13650, N13646, N7079, N8186);
nor NOR2 (N13651, N13634, N4334);
or OR3 (N13652, N13642, N10517, N6174);
not NOT1 (N13653, N13649);
xor XOR2 (N13654, N13637, N11687);
not NOT1 (N13655, N13643);
xor XOR2 (N13656, N13631, N4247);
and AND3 (N13657, N13627, N10807, N4575);
xor XOR2 (N13658, N13655, N3025);
nor NOR3 (N13659, N13657, N9608, N10506);
nor NOR3 (N13660, N13651, N6267, N8443);
xor XOR2 (N13661, N13652, N157);
nor NOR2 (N13662, N13654, N423);
xor XOR2 (N13663, N13656, N12680);
not NOT1 (N13664, N13658);
xor XOR2 (N13665, N13650, N8782);
nand NAND3 (N13666, N13647, N9650, N3087);
and AND3 (N13667, N13648, N5239, N10300);
xor XOR2 (N13668, N13663, N387);
or OR2 (N13669, N13659, N10465);
nand NAND4 (N13670, N13662, N2653, N12313, N858);
or OR3 (N13671, N13668, N6320, N4005);
nand NAND4 (N13672, N13664, N1609, N7771, N7283);
not NOT1 (N13673, N13667);
buf BUF1 (N13674, N13670);
nand NAND3 (N13675, N13653, N5976, N1198);
and AND4 (N13676, N13665, N12923, N8911, N9274);
or OR2 (N13677, N13675, N8879);
buf BUF1 (N13678, N13677);
not NOT1 (N13679, N13660);
and AND2 (N13680, N13678, N5945);
not NOT1 (N13681, N13671);
and AND2 (N13682, N13666, N7184);
or OR3 (N13683, N13679, N5929, N10114);
xor XOR2 (N13684, N13676, N12638);
buf BUF1 (N13685, N13681);
not NOT1 (N13686, N13661);
nand NAND3 (N13687, N13680, N748, N1572);
xor XOR2 (N13688, N13684, N2284);
not NOT1 (N13689, N13686);
buf BUF1 (N13690, N13687);
nor NOR4 (N13691, N13688, N6016, N12745, N2374);
not NOT1 (N13692, N13689);
xor XOR2 (N13693, N13682, N9600);
nor NOR2 (N13694, N13691, N13278);
xor XOR2 (N13695, N13674, N6904);
and AND4 (N13696, N13673, N837, N301, N5294);
xor XOR2 (N13697, N13695, N1876);
nor NOR4 (N13698, N13694, N7081, N11722, N1955);
xor XOR2 (N13699, N13690, N12451);
nor NOR3 (N13700, N13692, N8716, N2205);
not NOT1 (N13701, N13669);
not NOT1 (N13702, N13683);
or OR2 (N13703, N13672, N13019);
and AND4 (N13704, N13699, N8818, N11606, N1357);
or OR2 (N13705, N13702, N9616);
xor XOR2 (N13706, N13701, N8769);
buf BUF1 (N13707, N13698);
not NOT1 (N13708, N13705);
or OR4 (N13709, N13697, N1684, N12030, N670);
xor XOR2 (N13710, N13693, N9130);
or OR4 (N13711, N13700, N656, N1837, N30);
nand NAND2 (N13712, N13703, N7653);
and AND4 (N13713, N13712, N2821, N3172, N11553);
or OR3 (N13714, N13707, N13422, N6371);
not NOT1 (N13715, N13706);
xor XOR2 (N13716, N13713, N10136);
nor NOR3 (N13717, N13710, N10217, N13168);
buf BUF1 (N13718, N13717);
not NOT1 (N13719, N13711);
buf BUF1 (N13720, N13704);
nor NOR3 (N13721, N13718, N12032, N1854);
nor NOR2 (N13722, N13714, N10584);
and AND2 (N13723, N13709, N3177);
xor XOR2 (N13724, N13716, N10138);
buf BUF1 (N13725, N13696);
nor NOR3 (N13726, N13725, N6540, N5229);
not NOT1 (N13727, N13708);
not NOT1 (N13728, N13719);
and AND3 (N13729, N13728, N3559, N6670);
buf BUF1 (N13730, N13723);
and AND4 (N13731, N13727, N3096, N6914, N7892);
not NOT1 (N13732, N13685);
and AND3 (N13733, N13731, N9994, N3819);
and AND2 (N13734, N13732, N12988);
or OR4 (N13735, N13726, N414, N9106, N13167);
or OR2 (N13736, N13724, N9035);
xor XOR2 (N13737, N13734, N8567);
xor XOR2 (N13738, N13736, N1397);
not NOT1 (N13739, N13729);
and AND4 (N13740, N13738, N8852, N10972, N6997);
or OR3 (N13741, N13740, N4574, N6970);
or OR2 (N13742, N13721, N8422);
not NOT1 (N13743, N13742);
xor XOR2 (N13744, N13743, N3792);
buf BUF1 (N13745, N13715);
nor NOR4 (N13746, N13737, N7333, N2047, N2690);
nand NAND4 (N13747, N13720, N11885, N1096, N5926);
buf BUF1 (N13748, N13747);
nand NAND4 (N13749, N13730, N7093, N4792, N3597);
nand NAND4 (N13750, N13735, N4529, N8098, N3604);
nor NOR4 (N13751, N13749, N2360, N8917, N7958);
buf BUF1 (N13752, N13733);
nand NAND2 (N13753, N13748, N13044);
buf BUF1 (N13754, N13745);
buf BUF1 (N13755, N13744);
xor XOR2 (N13756, N13750, N11042);
xor XOR2 (N13757, N13754, N119);
and AND3 (N13758, N13756, N7690, N7600);
xor XOR2 (N13759, N13751, N10701);
and AND3 (N13760, N13758, N889, N11335);
nor NOR4 (N13761, N13755, N13738, N8322, N255);
and AND2 (N13762, N13746, N6261);
nand NAND2 (N13763, N13752, N12192);
and AND3 (N13764, N13722, N8716, N12567);
nor NOR2 (N13765, N13764, N10805);
nand NAND2 (N13766, N13762, N13603);
nand NAND3 (N13767, N13763, N5287, N8259);
nand NAND4 (N13768, N13739, N13015, N7866, N4293);
nor NOR3 (N13769, N13757, N9206, N7562);
buf BUF1 (N13770, N13768);
xor XOR2 (N13771, N13766, N12850);
xor XOR2 (N13772, N13769, N12803);
not NOT1 (N13773, N13772);
and AND3 (N13774, N13771, N6245, N1713);
nand NAND2 (N13775, N13741, N12156);
or OR2 (N13776, N13761, N1254);
not NOT1 (N13777, N13759);
and AND2 (N13778, N13765, N5919);
not NOT1 (N13779, N13776);
xor XOR2 (N13780, N13775, N10474);
buf BUF1 (N13781, N13760);
buf BUF1 (N13782, N13770);
buf BUF1 (N13783, N13767);
nand NAND2 (N13784, N13777, N8281);
xor XOR2 (N13785, N13784, N5099);
xor XOR2 (N13786, N13781, N10797);
or OR4 (N13787, N13753, N10752, N9384, N8951);
buf BUF1 (N13788, N13774);
and AND4 (N13789, N13786, N5369, N1931, N2701);
xor XOR2 (N13790, N13782, N4337);
xor XOR2 (N13791, N13790, N3599);
buf BUF1 (N13792, N13788);
buf BUF1 (N13793, N13791);
nand NAND3 (N13794, N13785, N539, N6920);
nor NOR3 (N13795, N13789, N10855, N12589);
or OR2 (N13796, N13783, N1250);
nor NOR4 (N13797, N13773, N6566, N915, N8666);
nor NOR3 (N13798, N13795, N1893, N13395);
buf BUF1 (N13799, N13797);
and AND4 (N13800, N13780, N5490, N6109, N9788);
or OR3 (N13801, N13794, N9752, N4491);
buf BUF1 (N13802, N13779);
nor NOR4 (N13803, N13800, N5456, N9063, N2525);
nand NAND3 (N13804, N13792, N7200, N11);
or OR2 (N13805, N13799, N10489);
nand NAND2 (N13806, N13803, N11876);
or OR3 (N13807, N13806, N8484, N630);
or OR4 (N13808, N13805, N5088, N1336, N12955);
not NOT1 (N13809, N13798);
not NOT1 (N13810, N13778);
buf BUF1 (N13811, N13810);
xor XOR2 (N13812, N13796, N11817);
xor XOR2 (N13813, N13804, N6712);
xor XOR2 (N13814, N13807, N7883);
nor NOR2 (N13815, N13811, N9307);
nand NAND3 (N13816, N13815, N3961, N11668);
nand NAND4 (N13817, N13812, N1941, N1639, N11852);
nand NAND4 (N13818, N13817, N4231, N10319, N9893);
not NOT1 (N13819, N13818);
buf BUF1 (N13820, N13802);
or OR2 (N13821, N13809, N7667);
nor NOR3 (N13822, N13808, N6196, N6523);
or OR3 (N13823, N13819, N2927, N10961);
nor NOR3 (N13824, N13787, N3146, N8069);
nor NOR4 (N13825, N13824, N10721, N6876, N9286);
buf BUF1 (N13826, N13820);
xor XOR2 (N13827, N13813, N6220);
nor NOR2 (N13828, N13823, N109);
nand NAND4 (N13829, N13826, N3796, N6395, N12050);
buf BUF1 (N13830, N13825);
xor XOR2 (N13831, N13814, N7714);
xor XOR2 (N13832, N13827, N2994);
or OR4 (N13833, N13832, N1256, N1383, N172);
xor XOR2 (N13834, N13829, N3813);
or OR2 (N13835, N13830, N3163);
nor NOR3 (N13836, N13822, N6890, N94);
not NOT1 (N13837, N13835);
not NOT1 (N13838, N13816);
or OR2 (N13839, N13836, N5579);
not NOT1 (N13840, N13837);
nor NOR2 (N13841, N13834, N2993);
nor NOR4 (N13842, N13801, N6162, N9138, N10436);
buf BUF1 (N13843, N13840);
xor XOR2 (N13844, N13821, N9188);
xor XOR2 (N13845, N13842, N11882);
xor XOR2 (N13846, N13831, N10152);
buf BUF1 (N13847, N13839);
not NOT1 (N13848, N13838);
buf BUF1 (N13849, N13844);
buf BUF1 (N13850, N13845);
xor XOR2 (N13851, N13846, N11281);
nor NOR2 (N13852, N13833, N6506);
xor XOR2 (N13853, N13841, N10191);
not NOT1 (N13854, N13851);
nor NOR4 (N13855, N13849, N10738, N7515, N12088);
not NOT1 (N13856, N13850);
not NOT1 (N13857, N13853);
xor XOR2 (N13858, N13847, N3902);
nor NOR4 (N13859, N13858, N5946, N3455, N12922);
nand NAND2 (N13860, N13852, N4575);
nor NOR3 (N13861, N13793, N8080, N3506);
xor XOR2 (N13862, N13859, N2217);
xor XOR2 (N13863, N13857, N11090);
and AND2 (N13864, N13854, N5200);
or OR4 (N13865, N13843, N11043, N4404, N38);
buf BUF1 (N13866, N13848);
buf BUF1 (N13867, N13860);
not NOT1 (N13868, N13864);
xor XOR2 (N13869, N13862, N574);
nor NOR3 (N13870, N13865, N2153, N8699);
not NOT1 (N13871, N13863);
xor XOR2 (N13872, N13868, N492);
xor XOR2 (N13873, N13872, N12021);
buf BUF1 (N13874, N13870);
or OR3 (N13875, N13861, N9273, N2558);
xor XOR2 (N13876, N13871, N11746);
nor NOR2 (N13877, N13869, N6119);
buf BUF1 (N13878, N13874);
xor XOR2 (N13879, N13876, N3225);
not NOT1 (N13880, N13873);
nand NAND2 (N13881, N13879, N9056);
not NOT1 (N13882, N13855);
or OR3 (N13883, N13866, N11672, N9042);
and AND2 (N13884, N13875, N5762);
xor XOR2 (N13885, N13880, N6072);
nand NAND4 (N13886, N13882, N4279, N10602, N3203);
xor XOR2 (N13887, N13878, N3877);
and AND3 (N13888, N13856, N11558, N1309);
nor NOR4 (N13889, N13887, N10156, N8074, N10400);
nand NAND4 (N13890, N13877, N12244, N10761, N11153);
xor XOR2 (N13891, N13885, N9619);
and AND2 (N13892, N13890, N5183);
buf BUF1 (N13893, N13891);
buf BUF1 (N13894, N13884);
nor NOR2 (N13895, N13883, N57);
nand NAND3 (N13896, N13889, N10661, N8213);
nand NAND4 (N13897, N13888, N3288, N12267, N330);
nor NOR4 (N13898, N13895, N6004, N9149, N13151);
and AND2 (N13899, N13893, N7216);
and AND2 (N13900, N13899, N6640);
not NOT1 (N13901, N13828);
nand NAND2 (N13902, N13886, N9929);
and AND2 (N13903, N13897, N12541);
xor XOR2 (N13904, N13903, N10896);
xor XOR2 (N13905, N13894, N9137);
nor NOR2 (N13906, N13881, N10703);
or OR2 (N13907, N13867, N12598);
not NOT1 (N13908, N13898);
buf BUF1 (N13909, N13906);
nor NOR4 (N13910, N13900, N6186, N11908, N13785);
xor XOR2 (N13911, N13901, N12975);
or OR2 (N13912, N13910, N2555);
and AND4 (N13913, N13912, N10240, N4350, N6331);
and AND3 (N13914, N13904, N2800, N148);
not NOT1 (N13915, N13905);
or OR2 (N13916, N13908, N2816);
not NOT1 (N13917, N13914);
buf BUF1 (N13918, N13916);
and AND3 (N13919, N13915, N290, N2267);
nand NAND2 (N13920, N13911, N1643);
xor XOR2 (N13921, N13913, N7598);
nand NAND3 (N13922, N13907, N6892, N1330);
nor NOR2 (N13923, N13922, N13539);
not NOT1 (N13924, N13921);
and AND3 (N13925, N13923, N1139, N1025);
nand NAND3 (N13926, N13924, N13490, N8261);
and AND3 (N13927, N13896, N8855, N5162);
nand NAND4 (N13928, N13927, N2876, N9376, N13816);
or OR2 (N13929, N13925, N11565);
not NOT1 (N13930, N13928);
nand NAND4 (N13931, N13920, N4046, N11474, N2548);
not NOT1 (N13932, N13929);
nand NAND4 (N13933, N13909, N4324, N3319, N4506);
or OR4 (N13934, N13902, N3446, N12545, N3318);
and AND3 (N13935, N13931, N7733, N859);
nand NAND2 (N13936, N13932, N8541);
and AND3 (N13937, N13936, N2305, N10562);
buf BUF1 (N13938, N13918);
not NOT1 (N13939, N13892);
or OR3 (N13940, N13930, N170, N4296);
nor NOR4 (N13941, N13934, N7863, N6533, N10828);
xor XOR2 (N13942, N13933, N8830);
and AND4 (N13943, N13919, N9806, N5693, N3200);
xor XOR2 (N13944, N13940, N1642);
nor NOR2 (N13945, N13943, N7988);
xor XOR2 (N13946, N13944, N313);
and AND4 (N13947, N13941, N147, N7159, N10015);
buf BUF1 (N13948, N13942);
or OR2 (N13949, N13935, N1519);
nor NOR4 (N13950, N13938, N3875, N8077, N10073);
buf BUF1 (N13951, N13939);
nor NOR3 (N13952, N13951, N6395, N9129);
buf BUF1 (N13953, N13947);
and AND2 (N13954, N13950, N12512);
or OR3 (N13955, N13937, N4717, N7061);
or OR2 (N13956, N13917, N8041);
nand NAND3 (N13957, N13953, N12338, N1190);
nor NOR4 (N13958, N13948, N4991, N13651, N12534);
xor XOR2 (N13959, N13946, N8879);
or OR4 (N13960, N13959, N164, N818, N12107);
or OR4 (N13961, N13960, N8444, N2055, N11444);
nor NOR4 (N13962, N13952, N12070, N6594, N777);
and AND4 (N13963, N13957, N3091, N56, N10843);
or OR4 (N13964, N13954, N8365, N8114, N4133);
not NOT1 (N13965, N13958);
nand NAND3 (N13966, N13963, N12413, N7205);
and AND2 (N13967, N13964, N8650);
buf BUF1 (N13968, N13966);
or OR4 (N13969, N13965, N2758, N10020, N306);
not NOT1 (N13970, N13949);
xor XOR2 (N13971, N13969, N2944);
nand NAND3 (N13972, N13961, N8145, N2470);
not NOT1 (N13973, N13967);
not NOT1 (N13974, N13945);
not NOT1 (N13975, N13973);
not NOT1 (N13976, N13962);
buf BUF1 (N13977, N13972);
not NOT1 (N13978, N13976);
xor XOR2 (N13979, N13926, N3503);
buf BUF1 (N13980, N13979);
buf BUF1 (N13981, N13978);
nor NOR4 (N13982, N13981, N1537, N1379, N13133);
and AND3 (N13983, N13955, N13089, N2229);
buf BUF1 (N13984, N13977);
and AND4 (N13985, N13956, N5294, N6755, N13389);
buf BUF1 (N13986, N13974);
xor XOR2 (N13987, N13971, N12046);
xor XOR2 (N13988, N13970, N10306);
nand NAND2 (N13989, N13985, N9644);
xor XOR2 (N13990, N13987, N2009);
not NOT1 (N13991, N13983);
xor XOR2 (N13992, N13982, N11404);
or OR2 (N13993, N13984, N10720);
nand NAND3 (N13994, N13993, N1371, N1966);
or OR2 (N13995, N13975, N3771);
and AND3 (N13996, N13988, N7797, N5767);
nand NAND2 (N13997, N13994, N5450);
not NOT1 (N13998, N13968);
not NOT1 (N13999, N13986);
or OR4 (N14000, N13989, N4137, N4049, N1307);
and AND4 (N14001, N13980, N774, N10716, N3405);
nor NOR3 (N14002, N13991, N6001, N12041);
and AND3 (N14003, N13998, N65, N7194);
or OR3 (N14004, N14001, N6106, N4900);
xor XOR2 (N14005, N13999, N1164);
xor XOR2 (N14006, N13990, N10768);
or OR2 (N14007, N14005, N6948);
and AND2 (N14008, N13997, N6889);
not NOT1 (N14009, N14007);
xor XOR2 (N14010, N13992, N12983);
nand NAND4 (N14011, N14008, N5550, N11105, N374);
buf BUF1 (N14012, N14010);
nand NAND4 (N14013, N14012, N8812, N7670, N7067);
nor NOR2 (N14014, N13996, N5774);
xor XOR2 (N14015, N14004, N2408);
nor NOR2 (N14016, N14013, N9021);
and AND3 (N14017, N14016, N4518, N13593);
or OR3 (N14018, N14003, N2176, N9950);
and AND3 (N14019, N14014, N8868, N2414);
and AND4 (N14020, N14015, N342, N2798, N13860);
buf BUF1 (N14021, N14018);
nand NAND3 (N14022, N14006, N10136, N12264);
nand NAND4 (N14023, N14017, N13481, N3700, N4596);
nand NAND4 (N14024, N14002, N10683, N7547, N3574);
nand NAND4 (N14025, N14019, N3823, N5464, N10653);
or OR2 (N14026, N14024, N9211);
and AND4 (N14027, N14000, N8998, N10482, N8357);
nor NOR2 (N14028, N14009, N3275);
nor NOR2 (N14029, N14028, N1563);
nor NOR4 (N14030, N14027, N10779, N3723, N1072);
or OR4 (N14031, N14022, N12607, N6199, N5165);
and AND3 (N14032, N14023, N7306, N11239);
xor XOR2 (N14033, N14021, N4507);
xor XOR2 (N14034, N14020, N9819);
xor XOR2 (N14035, N14033, N5304);
buf BUF1 (N14036, N14029);
nand NAND4 (N14037, N14026, N2751, N12924, N9233);
buf BUF1 (N14038, N14037);
nand NAND2 (N14039, N14036, N9503);
nand NAND3 (N14040, N14038, N10290, N7052);
xor XOR2 (N14041, N14032, N8907);
buf BUF1 (N14042, N14030);
xor XOR2 (N14043, N14040, N9296);
xor XOR2 (N14044, N14043, N233);
or OR4 (N14045, N14011, N10349, N4895, N7696);
nand NAND3 (N14046, N14031, N12842, N8477);
buf BUF1 (N14047, N14039);
or OR3 (N14048, N14035, N54, N6489);
not NOT1 (N14049, N13995);
and AND4 (N14050, N14044, N6579, N6345, N4714);
or OR4 (N14051, N14042, N457, N9599, N12936);
or OR4 (N14052, N14047, N5380, N13076, N3684);
buf BUF1 (N14053, N14052);
xor XOR2 (N14054, N14051, N365);
not NOT1 (N14055, N14045);
buf BUF1 (N14056, N14041);
buf BUF1 (N14057, N14048);
and AND3 (N14058, N14054, N5994, N2053);
nand NAND4 (N14059, N14025, N2364, N13456, N12243);
xor XOR2 (N14060, N14056, N4741);
buf BUF1 (N14061, N14034);
or OR3 (N14062, N14059, N6111, N13451);
and AND4 (N14063, N14058, N389, N12493, N9273);
nor NOR2 (N14064, N14057, N7849);
nor NOR3 (N14065, N14046, N8800, N10792);
or OR4 (N14066, N14049, N8230, N1082, N3066);
nand NAND2 (N14067, N14060, N4931);
nand NAND2 (N14068, N14066, N12843);
buf BUF1 (N14069, N14063);
nand NAND2 (N14070, N14062, N4406);
and AND4 (N14071, N14068, N836, N4784, N2687);
or OR3 (N14072, N14070, N8729, N8694);
or OR3 (N14073, N14050, N538, N7053);
xor XOR2 (N14074, N14072, N6090);
nor NOR4 (N14075, N14053, N12557, N2879, N119);
nor NOR2 (N14076, N14064, N11117);
nor NOR2 (N14077, N14075, N2802);
nand NAND4 (N14078, N14061, N310, N2580, N12645);
or OR4 (N14079, N14074, N13792, N2001, N6134);
nor NOR2 (N14080, N14077, N11582);
or OR3 (N14081, N14080, N2502, N8231);
and AND3 (N14082, N14073, N128, N10940);
xor XOR2 (N14083, N14071, N3096);
not NOT1 (N14084, N14076);
not NOT1 (N14085, N14084);
and AND3 (N14086, N14085, N4197, N6951);
or OR2 (N14087, N14055, N10044);
nor NOR2 (N14088, N14083, N2581);
nand NAND4 (N14089, N14081, N7554, N11974, N11054);
buf BUF1 (N14090, N14086);
buf BUF1 (N14091, N14087);
and AND4 (N14092, N14091, N3106, N6634, N13372);
nand NAND3 (N14093, N14065, N2894, N1031);
not NOT1 (N14094, N14090);
xor XOR2 (N14095, N14093, N11293);
xor XOR2 (N14096, N14094, N2159);
xor XOR2 (N14097, N14082, N9735);
nor NOR2 (N14098, N14088, N11940);
or OR3 (N14099, N14098, N5956, N2945);
xor XOR2 (N14100, N14078, N2971);
not NOT1 (N14101, N14097);
buf BUF1 (N14102, N14092);
or OR3 (N14103, N14100, N3482, N13568);
and AND2 (N14104, N14099, N13730);
or OR4 (N14105, N14096, N3993, N13463, N9680);
not NOT1 (N14106, N14105);
xor XOR2 (N14107, N14095, N4703);
buf BUF1 (N14108, N14069);
not NOT1 (N14109, N14067);
and AND4 (N14110, N14079, N5988, N3737, N9847);
buf BUF1 (N14111, N14102);
buf BUF1 (N14112, N14107);
not NOT1 (N14113, N14110);
and AND2 (N14114, N14112, N9419);
xor XOR2 (N14115, N14113, N9350);
and AND3 (N14116, N14104, N1496, N5427);
not NOT1 (N14117, N14114);
buf BUF1 (N14118, N14115);
not NOT1 (N14119, N14118);
buf BUF1 (N14120, N14119);
or OR2 (N14121, N14108, N13201);
buf BUF1 (N14122, N14117);
buf BUF1 (N14123, N14120);
or OR2 (N14124, N14122, N11857);
not NOT1 (N14125, N14101);
buf BUF1 (N14126, N14109);
and AND2 (N14127, N14126, N9844);
buf BUF1 (N14128, N14103);
xor XOR2 (N14129, N14128, N6884);
buf BUF1 (N14130, N14127);
buf BUF1 (N14131, N14111);
not NOT1 (N14132, N14123);
not NOT1 (N14133, N14106);
and AND4 (N14134, N14132, N1250, N8668, N11923);
buf BUF1 (N14135, N14125);
xor XOR2 (N14136, N14124, N7837);
nor NOR4 (N14137, N14131, N8227, N8753, N7683);
nand NAND4 (N14138, N14137, N7966, N7024, N6022);
nor NOR3 (N14139, N14136, N6816, N10901);
buf BUF1 (N14140, N14138);
not NOT1 (N14141, N14139);
or OR2 (N14142, N14133, N12828);
nand NAND3 (N14143, N14089, N4537, N12157);
or OR3 (N14144, N14121, N452, N4957);
or OR2 (N14145, N14116, N5026);
or OR3 (N14146, N14145, N12941, N12784);
or OR3 (N14147, N14143, N13431, N7053);
xor XOR2 (N14148, N14134, N3549);
and AND3 (N14149, N14130, N9085, N6108);
not NOT1 (N14150, N14148);
xor XOR2 (N14151, N14141, N7188);
and AND2 (N14152, N14129, N7102);
xor XOR2 (N14153, N14149, N7657);
xor XOR2 (N14154, N14152, N12840);
nor NOR3 (N14155, N14140, N5495, N624);
and AND3 (N14156, N14153, N4837, N13907);
nor NOR2 (N14157, N14154, N10846);
buf BUF1 (N14158, N14151);
buf BUF1 (N14159, N14150);
buf BUF1 (N14160, N14158);
xor XOR2 (N14161, N14155, N2155);
nand NAND4 (N14162, N14159, N4948, N397, N10515);
buf BUF1 (N14163, N14161);
not NOT1 (N14164, N14146);
nand NAND4 (N14165, N14156, N9593, N559, N12558);
xor XOR2 (N14166, N14165, N2228);
buf BUF1 (N14167, N14160);
nand NAND3 (N14168, N14167, N10862, N5097);
or OR4 (N14169, N14135, N12376, N10914, N6544);
or OR2 (N14170, N14157, N7608);
not NOT1 (N14171, N14142);
xor XOR2 (N14172, N14168, N7441);
nor NOR2 (N14173, N14147, N8123);
buf BUF1 (N14174, N14162);
nand NAND3 (N14175, N14170, N3264, N6000);
nor NOR4 (N14176, N14173, N10191, N12449, N12802);
nor NOR3 (N14177, N14171, N8927, N9767);
xor XOR2 (N14178, N14174, N9518);
xor XOR2 (N14179, N14175, N8004);
and AND2 (N14180, N14178, N7131);
nand NAND3 (N14181, N14163, N1879, N3886);
nor NOR3 (N14182, N14177, N7829, N13002);
nor NOR2 (N14183, N14169, N4076);
and AND4 (N14184, N14181, N10036, N11121, N11548);
not NOT1 (N14185, N14166);
nand NAND4 (N14186, N14172, N11795, N6990, N1891);
nand NAND4 (N14187, N14186, N12574, N11940, N6911);
xor XOR2 (N14188, N14179, N566);
and AND3 (N14189, N14144, N12504, N1491);
xor XOR2 (N14190, N14188, N13673);
or OR2 (N14191, N14183, N593);
xor XOR2 (N14192, N14164, N2064);
not NOT1 (N14193, N14176);
nor NOR3 (N14194, N14184, N6170, N8678);
nand NAND3 (N14195, N14182, N5419, N11282);
nand NAND2 (N14196, N14193, N9756);
buf BUF1 (N14197, N14190);
nand NAND4 (N14198, N14194, N13911, N11617, N5439);
and AND3 (N14199, N14180, N1017, N10601);
buf BUF1 (N14200, N14198);
or OR2 (N14201, N14192, N13060);
buf BUF1 (N14202, N14197);
nand NAND4 (N14203, N14200, N5946, N2210, N720);
buf BUF1 (N14204, N14199);
not NOT1 (N14205, N14203);
and AND4 (N14206, N14205, N12280, N1327, N3841);
buf BUF1 (N14207, N14202);
and AND2 (N14208, N14185, N10097);
nor NOR2 (N14209, N14187, N10912);
xor XOR2 (N14210, N14195, N8186);
and AND2 (N14211, N14191, N5588);
buf BUF1 (N14212, N14189);
nand NAND4 (N14213, N14208, N13864, N6957, N12294);
not NOT1 (N14214, N14196);
nand NAND2 (N14215, N14214, N3818);
not NOT1 (N14216, N14211);
nand NAND2 (N14217, N14210, N8041);
or OR2 (N14218, N14215, N9336);
nand NAND4 (N14219, N14209, N1766, N12306, N14037);
or OR3 (N14220, N14212, N3165, N4925);
or OR2 (N14221, N14207, N6118);
xor XOR2 (N14222, N14218, N8608);
not NOT1 (N14223, N14206);
not NOT1 (N14224, N14217);
not NOT1 (N14225, N14221);
buf BUF1 (N14226, N14201);
nor NOR3 (N14227, N14226, N1033, N13200);
or OR3 (N14228, N14216, N3505, N8754);
buf BUF1 (N14229, N14223);
or OR4 (N14230, N14220, N11416, N8230, N3333);
nand NAND4 (N14231, N14230, N14226, N8608, N13735);
or OR4 (N14232, N14219, N13273, N6535, N1281);
nor NOR2 (N14233, N14204, N14058);
nand NAND3 (N14234, N14224, N7696, N13703);
not NOT1 (N14235, N14229);
or OR3 (N14236, N14232, N11551, N1592);
not NOT1 (N14237, N14225);
nor NOR2 (N14238, N14233, N2121);
nand NAND2 (N14239, N14231, N7219);
and AND2 (N14240, N14235, N753);
xor XOR2 (N14241, N14228, N2608);
buf BUF1 (N14242, N14237);
not NOT1 (N14243, N14241);
and AND4 (N14244, N14242, N14171, N11318, N3107);
xor XOR2 (N14245, N14238, N3349);
xor XOR2 (N14246, N14234, N2819);
xor XOR2 (N14247, N14244, N10352);
nor NOR4 (N14248, N14236, N12168, N128, N10404);
nand NAND3 (N14249, N14248, N5287, N7743);
buf BUF1 (N14250, N14245);
buf BUF1 (N14251, N14240);
nor NOR2 (N14252, N14243, N2972);
xor XOR2 (N14253, N14251, N11975);
nor NOR3 (N14254, N14213, N11516, N3309);
nor NOR2 (N14255, N14247, N447);
buf BUF1 (N14256, N14222);
nor NOR2 (N14257, N14239, N5003);
nor NOR4 (N14258, N14246, N6987, N4230, N9296);
buf BUF1 (N14259, N14254);
xor XOR2 (N14260, N14256, N12790);
nand NAND2 (N14261, N14260, N9613);
and AND4 (N14262, N14258, N2760, N7442, N13007);
or OR4 (N14263, N14255, N2680, N9696, N4302);
not NOT1 (N14264, N14252);
buf BUF1 (N14265, N14261);
or OR4 (N14266, N14249, N709, N13585, N2566);
or OR4 (N14267, N14227, N1222, N7679, N8588);
buf BUF1 (N14268, N14266);
or OR4 (N14269, N14253, N7203, N8889, N557);
buf BUF1 (N14270, N14257);
xor XOR2 (N14271, N14269, N12445);
and AND2 (N14272, N14259, N8204);
and AND3 (N14273, N14270, N9514, N6963);
nand NAND2 (N14274, N14268, N5067);
not NOT1 (N14275, N14267);
xor XOR2 (N14276, N14275, N7651);
xor XOR2 (N14277, N14264, N2953);
nand NAND4 (N14278, N14271, N8962, N11473, N388);
and AND4 (N14279, N14274, N4020, N7760, N825);
or OR3 (N14280, N14276, N2089, N9106);
xor XOR2 (N14281, N14280, N1495);
buf BUF1 (N14282, N14281);
buf BUF1 (N14283, N14278);
not NOT1 (N14284, N14273);
xor XOR2 (N14285, N14283, N971);
buf BUF1 (N14286, N14262);
buf BUF1 (N14287, N14282);
nand NAND3 (N14288, N14277, N6181, N8168);
and AND2 (N14289, N14272, N5227);
buf BUF1 (N14290, N14285);
buf BUF1 (N14291, N14265);
nand NAND4 (N14292, N14263, N11243, N1504, N6683);
nand NAND4 (N14293, N14288, N120, N8460, N2234);
buf BUF1 (N14294, N14289);
xor XOR2 (N14295, N14250, N3929);
and AND2 (N14296, N14294, N8591);
and AND2 (N14297, N14295, N9158);
not NOT1 (N14298, N14290);
xor XOR2 (N14299, N14292, N9830);
buf BUF1 (N14300, N14284);
not NOT1 (N14301, N14287);
buf BUF1 (N14302, N14296);
nor NOR3 (N14303, N14286, N6633, N826);
nand NAND4 (N14304, N14301, N9747, N7608, N8507);
buf BUF1 (N14305, N14293);
buf BUF1 (N14306, N14300);
or OR2 (N14307, N14303, N646);
nand NAND4 (N14308, N14298, N8050, N11204, N9195);
buf BUF1 (N14309, N14297);
not NOT1 (N14310, N14304);
nand NAND2 (N14311, N14307, N3241);
and AND3 (N14312, N14311, N10380, N12056);
buf BUF1 (N14313, N14291);
not NOT1 (N14314, N14306);
not NOT1 (N14315, N14299);
nand NAND4 (N14316, N14308, N7857, N6488, N4969);
buf BUF1 (N14317, N14314);
not NOT1 (N14318, N14315);
not NOT1 (N14319, N14313);
buf BUF1 (N14320, N14302);
xor XOR2 (N14321, N14319, N9070);
or OR2 (N14322, N14309, N387);
and AND3 (N14323, N14279, N11551, N640);
buf BUF1 (N14324, N14322);
not NOT1 (N14325, N14317);
buf BUF1 (N14326, N14325);
nand NAND2 (N14327, N14324, N1213);
or OR3 (N14328, N14321, N11789, N6069);
and AND2 (N14329, N14318, N13458);
or OR2 (N14330, N14320, N6001);
and AND3 (N14331, N14330, N3146, N13030);
nand NAND3 (N14332, N14329, N1838, N8722);
and AND4 (N14333, N14305, N3616, N13413, N14022);
nand NAND3 (N14334, N14331, N9054, N4862);
buf BUF1 (N14335, N14310);
not NOT1 (N14336, N14327);
nor NOR4 (N14337, N14332, N13748, N2328, N6093);
nand NAND3 (N14338, N14337, N8463, N11109);
and AND3 (N14339, N14334, N4348, N3249);
and AND3 (N14340, N14312, N3252, N4072);
and AND3 (N14341, N14335, N11341, N3767);
buf BUF1 (N14342, N14338);
or OR3 (N14343, N14316, N12706, N7145);
nand NAND2 (N14344, N14342, N7469);
not NOT1 (N14345, N14344);
nor NOR3 (N14346, N14339, N769, N12266);
or OR3 (N14347, N14345, N9252, N8919);
not NOT1 (N14348, N14340);
nor NOR4 (N14349, N14323, N2804, N3220, N12276);
or OR2 (N14350, N14349, N12861);
and AND2 (N14351, N14350, N11877);
xor XOR2 (N14352, N14346, N480);
nor NOR4 (N14353, N14326, N7293, N7167, N1050);
nand NAND3 (N14354, N14347, N5615, N2610);
nor NOR2 (N14355, N14328, N1674);
and AND4 (N14356, N14341, N9090, N13942, N2821);
nand NAND4 (N14357, N14343, N9788, N3464, N5423);
buf BUF1 (N14358, N14352);
xor XOR2 (N14359, N14333, N3294);
nor NOR3 (N14360, N14351, N7393, N3731);
nor NOR2 (N14361, N14353, N14338);
nand NAND4 (N14362, N14359, N296, N7023, N2545);
xor XOR2 (N14363, N14360, N9922);
nand NAND2 (N14364, N14358, N5747);
not NOT1 (N14365, N14356);
and AND3 (N14366, N14361, N11254, N7144);
buf BUF1 (N14367, N14336);
not NOT1 (N14368, N14354);
nor NOR4 (N14369, N14363, N14140, N9682, N11591);
nand NAND2 (N14370, N14348, N11878);
nand NAND3 (N14371, N14357, N7655, N7524);
and AND3 (N14372, N14370, N7824, N10992);
nor NOR3 (N14373, N14368, N12813, N3623);
xor XOR2 (N14374, N14373, N255);
not NOT1 (N14375, N14365);
xor XOR2 (N14376, N14375, N8496);
not NOT1 (N14377, N14364);
buf BUF1 (N14378, N14355);
buf BUF1 (N14379, N14377);
nor NOR2 (N14380, N14376, N4856);
and AND4 (N14381, N14379, N7279, N9596, N2111);
buf BUF1 (N14382, N14366);
nor NOR2 (N14383, N14380, N5609);
or OR4 (N14384, N14369, N3403, N10956, N4116);
or OR2 (N14385, N14372, N13853);
xor XOR2 (N14386, N14371, N4472);
nor NOR2 (N14387, N14367, N12910);
and AND3 (N14388, N14386, N4442, N9232);
not NOT1 (N14389, N14383);
and AND3 (N14390, N14374, N3378, N2427);
nor NOR3 (N14391, N14384, N2865, N7531);
and AND2 (N14392, N14378, N542);
not NOT1 (N14393, N14391);
nand NAND2 (N14394, N14387, N10043);
and AND3 (N14395, N14390, N14061, N5683);
not NOT1 (N14396, N14381);
and AND2 (N14397, N14394, N2359);
nor NOR4 (N14398, N14392, N8592, N3417, N1635);
nor NOR4 (N14399, N14395, N7860, N11246, N2160);
nand NAND2 (N14400, N14382, N9821);
not NOT1 (N14401, N14397);
not NOT1 (N14402, N14399);
nor NOR3 (N14403, N14393, N14332, N8975);
or OR3 (N14404, N14398, N7479, N801);
buf BUF1 (N14405, N14389);
nand NAND3 (N14406, N14403, N8322, N8477);
nand NAND4 (N14407, N14396, N787, N3230, N2897);
xor XOR2 (N14408, N14362, N12679);
xor XOR2 (N14409, N14402, N2455);
buf BUF1 (N14410, N14405);
nand NAND4 (N14411, N14388, N5980, N11285, N10228);
or OR3 (N14412, N14407, N8848, N2275);
not NOT1 (N14413, N14408);
xor XOR2 (N14414, N14413, N10074);
nor NOR3 (N14415, N14414, N4183, N7957);
xor XOR2 (N14416, N14404, N1053);
or OR2 (N14417, N14410, N12158);
or OR3 (N14418, N14409, N13288, N6838);
buf BUF1 (N14419, N14416);
not NOT1 (N14420, N14400);
nand NAND2 (N14421, N14418, N10265);
buf BUF1 (N14422, N14401);
and AND4 (N14423, N14419, N9799, N11635, N1869);
and AND2 (N14424, N14406, N3540);
not NOT1 (N14425, N14420);
nand NAND3 (N14426, N14415, N8710, N7406);
nor NOR2 (N14427, N14424, N433);
and AND3 (N14428, N14425, N14219, N4783);
nand NAND2 (N14429, N14421, N982);
not NOT1 (N14430, N14417);
buf BUF1 (N14431, N14412);
nand NAND2 (N14432, N14429, N11007);
xor XOR2 (N14433, N14427, N13579);
nand NAND4 (N14434, N14430, N11604, N6615, N6004);
nor NOR4 (N14435, N14434, N2725, N6988, N9968);
xor XOR2 (N14436, N14423, N3805);
and AND3 (N14437, N14436, N3329, N5320);
not NOT1 (N14438, N14437);
buf BUF1 (N14439, N14426);
nand NAND4 (N14440, N14428, N10739, N10507, N3422);
nor NOR3 (N14441, N14432, N7607, N3677);
nor NOR3 (N14442, N14422, N13995, N697);
and AND3 (N14443, N14431, N1554, N12116);
or OR4 (N14444, N14385, N6649, N11379, N1253);
or OR3 (N14445, N14435, N3178, N1355);
buf BUF1 (N14446, N14439);
not NOT1 (N14447, N14442);
nand NAND4 (N14448, N14438, N5849, N493, N769);
and AND3 (N14449, N14445, N8203, N5128);
not NOT1 (N14450, N14444);
xor XOR2 (N14451, N14447, N3321);
not NOT1 (N14452, N14450);
and AND3 (N14453, N14451, N6298, N4491);
and AND2 (N14454, N14449, N9699);
or OR2 (N14455, N14448, N5526);
nor NOR2 (N14456, N14446, N10610);
buf BUF1 (N14457, N14455);
nand NAND3 (N14458, N14433, N7995, N10661);
or OR4 (N14459, N14411, N8023, N10566, N8209);
and AND4 (N14460, N14454, N7871, N8013, N11617);
nand NAND4 (N14461, N14459, N4743, N299, N3389);
buf BUF1 (N14462, N14456);
and AND4 (N14463, N14453, N448, N3468, N3116);
buf BUF1 (N14464, N14458);
and AND3 (N14465, N14463, N3634, N978);
buf BUF1 (N14466, N14452);
buf BUF1 (N14467, N14460);
nand NAND4 (N14468, N14461, N14146, N12500, N5115);
xor XOR2 (N14469, N14457, N13091);
or OR3 (N14470, N14464, N667, N8321);
buf BUF1 (N14471, N14441);
nor NOR2 (N14472, N14468, N14434);
nor NOR2 (N14473, N14443, N5228);
or OR3 (N14474, N14472, N11655, N5645);
and AND4 (N14475, N14469, N13628, N2045, N1284);
nand NAND4 (N14476, N14473, N12759, N1562, N8128);
xor XOR2 (N14477, N14466, N4986);
or OR3 (N14478, N14476, N11252, N13381);
buf BUF1 (N14479, N14474);
nand NAND2 (N14480, N14470, N5929);
not NOT1 (N14481, N14477);
nand NAND4 (N14482, N14462, N1347, N889, N3801);
buf BUF1 (N14483, N14482);
or OR2 (N14484, N14481, N12608);
not NOT1 (N14485, N14479);
nand NAND3 (N14486, N14475, N13980, N12102);
and AND2 (N14487, N14471, N9574);
or OR2 (N14488, N14483, N5108);
buf BUF1 (N14489, N14465);
nor NOR2 (N14490, N14485, N3696);
and AND3 (N14491, N14488, N4539, N1445);
xor XOR2 (N14492, N14491, N12045);
nor NOR2 (N14493, N14489, N8239);
nor NOR2 (N14494, N14467, N1897);
and AND2 (N14495, N14492, N3342);
xor XOR2 (N14496, N14484, N11188);
or OR4 (N14497, N14487, N4811, N13387, N8065);
nor NOR3 (N14498, N14496, N4287, N9385);
buf BUF1 (N14499, N14480);
and AND2 (N14500, N14478, N5180);
not NOT1 (N14501, N14490);
not NOT1 (N14502, N14494);
buf BUF1 (N14503, N14493);
buf BUF1 (N14504, N14500);
or OR4 (N14505, N14486, N6441, N10763, N4526);
not NOT1 (N14506, N14440);
or OR3 (N14507, N14504, N2329, N10528);
nand NAND2 (N14508, N14497, N330);
xor XOR2 (N14509, N14506, N8836);
or OR2 (N14510, N14495, N14119);
and AND2 (N14511, N14502, N10727);
buf BUF1 (N14512, N14509);
nand NAND2 (N14513, N14501, N2461);
or OR2 (N14514, N14503, N5553);
xor XOR2 (N14515, N14511, N3012);
and AND3 (N14516, N14512, N8666, N2432);
or OR4 (N14517, N14498, N13625, N2261, N137);
nand NAND2 (N14518, N14515, N6584);
nand NAND2 (N14519, N14505, N11054);
buf BUF1 (N14520, N14518);
or OR3 (N14521, N14517, N5398, N12155);
or OR2 (N14522, N14513, N12622);
or OR2 (N14523, N14510, N343);
xor XOR2 (N14524, N14523, N4812);
and AND3 (N14525, N14524, N2775, N6448);
nor NOR3 (N14526, N14508, N11363, N2789);
buf BUF1 (N14527, N14507);
and AND2 (N14528, N14514, N10944);
buf BUF1 (N14529, N14519);
and AND4 (N14530, N14520, N10332, N6949, N14339);
buf BUF1 (N14531, N14516);
nand NAND2 (N14532, N14528, N10161);
not NOT1 (N14533, N14532);
and AND2 (N14534, N14521, N4616);
and AND4 (N14535, N14529, N248, N5209, N3792);
not NOT1 (N14536, N14522);
buf BUF1 (N14537, N14531);
xor XOR2 (N14538, N14534, N5886);
not NOT1 (N14539, N14533);
nor NOR4 (N14540, N14530, N6222, N1984, N12266);
buf BUF1 (N14541, N14527);
or OR3 (N14542, N14499, N1699, N13924);
and AND3 (N14543, N14535, N10695, N8219);
not NOT1 (N14544, N14537);
not NOT1 (N14545, N14543);
not NOT1 (N14546, N14526);
and AND4 (N14547, N14542, N9980, N11582, N7827);
or OR4 (N14548, N14544, N10455, N12340, N11374);
or OR3 (N14549, N14525, N2004, N10737);
nand NAND2 (N14550, N14536, N10326);
xor XOR2 (N14551, N14550, N8458);
buf BUF1 (N14552, N14540);
nor NOR4 (N14553, N14538, N11157, N8675, N5455);
and AND3 (N14554, N14546, N2073, N14369);
buf BUF1 (N14555, N14539);
nor NOR2 (N14556, N14547, N7703);
xor XOR2 (N14557, N14545, N10894);
not NOT1 (N14558, N14553);
nand NAND3 (N14559, N14552, N4677, N4078);
buf BUF1 (N14560, N14551);
or OR3 (N14561, N14554, N5957, N952);
xor XOR2 (N14562, N14557, N10107);
nand NAND4 (N14563, N14556, N1898, N12249, N2320);
nand NAND4 (N14564, N14541, N11661, N8673, N7130);
and AND2 (N14565, N14558, N737);
and AND2 (N14566, N14559, N3430);
nand NAND3 (N14567, N14548, N12958, N1390);
or OR2 (N14568, N14560, N10847);
not NOT1 (N14569, N14568);
buf BUF1 (N14570, N14555);
or OR4 (N14571, N14569, N1032, N10640, N4101);
nor NOR2 (N14572, N14570, N11979);
xor XOR2 (N14573, N14571, N2836);
nand NAND3 (N14574, N14564, N9258, N3252);
nand NAND2 (N14575, N14567, N3808);
and AND3 (N14576, N14562, N2097, N4669);
xor XOR2 (N14577, N14563, N1031);
nand NAND4 (N14578, N14561, N2433, N10701, N3479);
or OR3 (N14579, N14574, N9975, N4486);
not NOT1 (N14580, N14549);
nor NOR3 (N14581, N14565, N6876, N3121);
not NOT1 (N14582, N14575);
and AND3 (N14583, N14582, N10773, N6601);
nand NAND4 (N14584, N14579, N10013, N7601, N13343);
buf BUF1 (N14585, N14578);
xor XOR2 (N14586, N14576, N1391);
buf BUF1 (N14587, N14572);
xor XOR2 (N14588, N14566, N13313);
buf BUF1 (N14589, N14584);
xor XOR2 (N14590, N14587, N6525);
nand NAND4 (N14591, N14585, N8190, N7708, N12169);
nand NAND3 (N14592, N14580, N5247, N13312);
xor XOR2 (N14593, N14586, N9216);
or OR3 (N14594, N14593, N3386, N798);
not NOT1 (N14595, N14573);
not NOT1 (N14596, N14595);
not NOT1 (N14597, N14592);
and AND2 (N14598, N14597, N10657);
xor XOR2 (N14599, N14581, N11402);
nor NOR4 (N14600, N14577, N4671, N2581, N7158);
not NOT1 (N14601, N14594);
or OR3 (N14602, N14599, N12319, N3301);
not NOT1 (N14603, N14596);
not NOT1 (N14604, N14598);
and AND2 (N14605, N14588, N8890);
not NOT1 (N14606, N14583);
not NOT1 (N14607, N14600);
or OR2 (N14608, N14589, N11541);
nand NAND2 (N14609, N14606, N11262);
nand NAND3 (N14610, N14601, N455, N8625);
not NOT1 (N14611, N14602);
not NOT1 (N14612, N14611);
nand NAND4 (N14613, N14605, N10038, N11624, N299);
or OR4 (N14614, N14607, N14584, N4097, N3502);
and AND2 (N14615, N14612, N1017);
nor NOR4 (N14616, N14610, N2667, N6094, N1067);
nand NAND2 (N14617, N14590, N4335);
and AND4 (N14618, N14613, N3041, N13535, N3459);
nor NOR2 (N14619, N14617, N12337);
buf BUF1 (N14620, N14608);
or OR2 (N14621, N14615, N9607);
not NOT1 (N14622, N14591);
or OR2 (N14623, N14618, N5976);
nor NOR2 (N14624, N14604, N9423);
and AND3 (N14625, N14619, N2235, N10143);
nor NOR3 (N14626, N14609, N4535, N10097);
or OR3 (N14627, N14622, N6009, N3479);
xor XOR2 (N14628, N14616, N9340);
not NOT1 (N14629, N14620);
or OR4 (N14630, N14624, N10280, N11768, N4846);
nor NOR2 (N14631, N14614, N7414);
nand NAND3 (N14632, N14631, N4236, N12134);
xor XOR2 (N14633, N14603, N6302);
buf BUF1 (N14634, N14630);
buf BUF1 (N14635, N14629);
or OR3 (N14636, N14633, N529, N5123);
and AND4 (N14637, N14628, N6147, N1094, N10770);
and AND4 (N14638, N14626, N3435, N5907, N505);
not NOT1 (N14639, N14632);
not NOT1 (N14640, N14623);
xor XOR2 (N14641, N14638, N13743);
buf BUF1 (N14642, N14621);
buf BUF1 (N14643, N14627);
buf BUF1 (N14644, N14625);
buf BUF1 (N14645, N14637);
and AND3 (N14646, N14645, N9885, N7219);
or OR4 (N14647, N14636, N7093, N1822, N9049);
not NOT1 (N14648, N14646);
nand NAND3 (N14649, N14643, N858, N3704);
buf BUF1 (N14650, N14635);
not NOT1 (N14651, N14639);
xor XOR2 (N14652, N14651, N13151);
nand NAND3 (N14653, N14649, N14344, N8965);
xor XOR2 (N14654, N14653, N14618);
and AND3 (N14655, N14644, N2707, N14394);
xor XOR2 (N14656, N14648, N8527);
and AND2 (N14657, N14642, N8824);
not NOT1 (N14658, N14652);
buf BUF1 (N14659, N14647);
or OR4 (N14660, N14640, N12717, N8716, N3569);
buf BUF1 (N14661, N14641);
not NOT1 (N14662, N14634);
xor XOR2 (N14663, N14654, N10614);
xor XOR2 (N14664, N14656, N10895);
nor NOR4 (N14665, N14659, N11093, N5898, N5045);
buf BUF1 (N14666, N14655);
not NOT1 (N14667, N14663);
and AND3 (N14668, N14665, N5124, N10724);
nand NAND4 (N14669, N14661, N7096, N4172, N1400);
buf BUF1 (N14670, N14650);
buf BUF1 (N14671, N14660);
xor XOR2 (N14672, N14667, N1540);
xor XOR2 (N14673, N14658, N3423);
and AND4 (N14674, N14666, N12683, N12054, N2911);
and AND2 (N14675, N14670, N6329);
nand NAND2 (N14676, N14657, N1159);
or OR2 (N14677, N14675, N14109);
nor NOR3 (N14678, N14674, N4833, N6248);
nand NAND2 (N14679, N14668, N9235);
and AND3 (N14680, N14662, N11524, N1928);
nor NOR4 (N14681, N14676, N11947, N8474, N4838);
not NOT1 (N14682, N14669);
nand NAND3 (N14683, N14678, N8751, N13286);
xor XOR2 (N14684, N14682, N13585);
and AND2 (N14685, N14673, N8528);
or OR2 (N14686, N14680, N10832);
buf BUF1 (N14687, N14685);
nor NOR3 (N14688, N14683, N14450, N4654);
nor NOR2 (N14689, N14671, N3901);
nor NOR3 (N14690, N14687, N5065, N5100);
not NOT1 (N14691, N14672);
nand NAND3 (N14692, N14681, N2940, N9735);
buf BUF1 (N14693, N14689);
or OR4 (N14694, N14664, N11536, N2250, N5915);
nand NAND3 (N14695, N14691, N10771, N13542);
or OR2 (N14696, N14692, N1674);
nor NOR4 (N14697, N14688, N6408, N4689, N6279);
xor XOR2 (N14698, N14679, N9356);
not NOT1 (N14699, N14696);
and AND3 (N14700, N14699, N11205, N8120);
nor NOR4 (N14701, N14698, N5688, N9879, N14530);
nor NOR2 (N14702, N14684, N9986);
and AND3 (N14703, N14690, N10731, N12323);
nand NAND4 (N14704, N14686, N9394, N1817, N12387);
and AND4 (N14705, N14695, N4420, N4293, N3950);
not NOT1 (N14706, N14703);
xor XOR2 (N14707, N14697, N11195);
nand NAND4 (N14708, N14706, N8027, N10113, N5209);
and AND4 (N14709, N14702, N2538, N14191, N6548);
not NOT1 (N14710, N14694);
and AND2 (N14711, N14705, N12720);
and AND2 (N14712, N14704, N625);
buf BUF1 (N14713, N14707);
buf BUF1 (N14714, N14693);
or OR3 (N14715, N14713, N11505, N6835);
and AND4 (N14716, N14714, N11656, N9146, N5050);
nand NAND4 (N14717, N14708, N13860, N3724, N10969);
not NOT1 (N14718, N14715);
xor XOR2 (N14719, N14712, N2317);
and AND2 (N14720, N14701, N5379);
or OR3 (N14721, N14718, N14180, N1136);
xor XOR2 (N14722, N14717, N8655);
or OR3 (N14723, N14721, N7638, N10778);
buf BUF1 (N14724, N14719);
nand NAND2 (N14725, N14723, N10198);
or OR2 (N14726, N14722, N2974);
not NOT1 (N14727, N14677);
xor XOR2 (N14728, N14725, N6689);
xor XOR2 (N14729, N14709, N4270);
not NOT1 (N14730, N14716);
nand NAND3 (N14731, N14728, N7435, N6069);
nand NAND2 (N14732, N14710, N8229);
buf BUF1 (N14733, N14700);
and AND3 (N14734, N14711, N7528, N13272);
nand NAND2 (N14735, N14733, N7043);
or OR2 (N14736, N14720, N6345);
nor NOR2 (N14737, N14727, N4653);
buf BUF1 (N14738, N14734);
nand NAND2 (N14739, N14738, N12066);
nand NAND2 (N14740, N14736, N11446);
or OR2 (N14741, N14732, N13665);
nor NOR4 (N14742, N14724, N12566, N8062, N1179);
or OR3 (N14743, N14735, N10592, N4026);
not NOT1 (N14744, N14743);
nand NAND4 (N14745, N14742, N1244, N5696, N75);
nor NOR3 (N14746, N14739, N14493, N12647);
nor NOR3 (N14747, N14741, N3265, N11145);
not NOT1 (N14748, N14737);
or OR3 (N14749, N14729, N10167, N13999);
not NOT1 (N14750, N14731);
not NOT1 (N14751, N14750);
or OR3 (N14752, N14740, N1393, N12132);
and AND4 (N14753, N14730, N8086, N6687, N9891);
xor XOR2 (N14754, N14745, N11199);
buf BUF1 (N14755, N14751);
or OR2 (N14756, N14755, N13545);
buf BUF1 (N14757, N14748);
buf BUF1 (N14758, N14726);
or OR3 (N14759, N14747, N3074, N1175);
or OR3 (N14760, N14756, N29, N181);
and AND3 (N14761, N14749, N10351, N4756);
or OR4 (N14762, N14754, N9897, N9854, N3332);
and AND3 (N14763, N14762, N2624, N7038);
not NOT1 (N14764, N14760);
nand NAND4 (N14765, N14744, N13565, N4317, N10074);
and AND3 (N14766, N14752, N13571, N4220);
nor NOR3 (N14767, N14765, N9699, N8767);
or OR3 (N14768, N14757, N11859, N4954);
nand NAND4 (N14769, N14764, N9202, N6739, N10487);
or OR2 (N14770, N14767, N4671);
nor NOR4 (N14771, N14761, N13401, N11703, N304);
xor XOR2 (N14772, N14753, N4385);
xor XOR2 (N14773, N14770, N1856);
nor NOR4 (N14774, N14758, N6546, N12110, N5129);
or OR4 (N14775, N14774, N10518, N12641, N12569);
or OR4 (N14776, N14773, N4458, N2938, N8290);
nor NOR2 (N14777, N14769, N14480);
buf BUF1 (N14778, N14772);
nor NOR4 (N14779, N14746, N13277, N5598, N1197);
and AND3 (N14780, N14777, N10665, N2790);
not NOT1 (N14781, N14775);
and AND4 (N14782, N14776, N5145, N8905, N3638);
not NOT1 (N14783, N14778);
nand NAND3 (N14784, N14759, N2064, N2353);
nand NAND4 (N14785, N14768, N13131, N12927, N13948);
nor NOR3 (N14786, N14782, N4654, N2788);
buf BUF1 (N14787, N14781);
xor XOR2 (N14788, N14771, N11653);
not NOT1 (N14789, N14785);
or OR3 (N14790, N14789, N10150, N8838);
and AND2 (N14791, N14763, N5300);
buf BUF1 (N14792, N14791);
or OR2 (N14793, N14779, N5443);
and AND3 (N14794, N14792, N11508, N8072);
and AND4 (N14795, N14794, N3668, N4553, N12333);
nor NOR4 (N14796, N14793, N10161, N8848, N1989);
or OR3 (N14797, N14784, N4413, N14794);
or OR3 (N14798, N14766, N4134, N14146);
nor NOR4 (N14799, N14780, N673, N5336, N4305);
or OR2 (N14800, N14787, N5335);
xor XOR2 (N14801, N14797, N9435);
nand NAND4 (N14802, N14799, N7718, N1305, N7851);
xor XOR2 (N14803, N14786, N6207);
xor XOR2 (N14804, N14803, N10306);
nor NOR2 (N14805, N14788, N12958);
nand NAND3 (N14806, N14783, N2469, N8411);
and AND4 (N14807, N14798, N2393, N11010, N11140);
nor NOR2 (N14808, N14800, N3379);
nor NOR2 (N14809, N14795, N7891);
or OR3 (N14810, N14802, N7607, N7208);
nand NAND3 (N14811, N14805, N14078, N6410);
xor XOR2 (N14812, N14807, N870);
nor NOR2 (N14813, N14811, N3554);
not NOT1 (N14814, N14804);
nor NOR4 (N14815, N14801, N6680, N5651, N5312);
nand NAND3 (N14816, N14806, N14259, N8524);
not NOT1 (N14817, N14790);
nand NAND3 (N14818, N14810, N12047, N12947);
nand NAND4 (N14819, N14809, N2390, N7640, N4414);
or OR2 (N14820, N14818, N3585);
buf BUF1 (N14821, N14813);
not NOT1 (N14822, N14817);
buf BUF1 (N14823, N14822);
not NOT1 (N14824, N14808);
xor XOR2 (N14825, N14824, N4800);
xor XOR2 (N14826, N14812, N12726);
nand NAND3 (N14827, N14796, N2651, N5674);
xor XOR2 (N14828, N14825, N10964);
not NOT1 (N14829, N14815);
nor NOR2 (N14830, N14828, N4500);
xor XOR2 (N14831, N14816, N1727);
not NOT1 (N14832, N14819);
buf BUF1 (N14833, N14830);
not NOT1 (N14834, N14826);
and AND3 (N14835, N14814, N13597, N13088);
nor NOR4 (N14836, N14835, N1195, N2580, N10549);
xor XOR2 (N14837, N14820, N3106);
not NOT1 (N14838, N14823);
not NOT1 (N14839, N14837);
and AND3 (N14840, N14832, N4860, N1272);
xor XOR2 (N14841, N14829, N382);
nand NAND3 (N14842, N14840, N11661, N382);
buf BUF1 (N14843, N14841);
nor NOR2 (N14844, N14843, N10649);
nand NAND4 (N14845, N14844, N2427, N8083, N4313);
xor XOR2 (N14846, N14836, N8690);
xor XOR2 (N14847, N14821, N11637);
nor NOR2 (N14848, N14845, N13660);
or OR3 (N14849, N14838, N14643, N5747);
and AND2 (N14850, N14834, N3761);
xor XOR2 (N14851, N14848, N6122);
nor NOR4 (N14852, N14839, N9718, N13663, N3165);
nor NOR4 (N14853, N14831, N5020, N5850, N14703);
buf BUF1 (N14854, N14827);
buf BUF1 (N14855, N14833);
and AND2 (N14856, N14846, N13053);
xor XOR2 (N14857, N14855, N10613);
buf BUF1 (N14858, N14857);
xor XOR2 (N14859, N14849, N3411);
xor XOR2 (N14860, N14852, N8233);
nand NAND4 (N14861, N14851, N4871, N503, N6384);
nand NAND3 (N14862, N14860, N13452, N14309);
and AND4 (N14863, N14853, N10058, N5251, N2961);
not NOT1 (N14864, N14854);
not NOT1 (N14865, N14842);
buf BUF1 (N14866, N14847);
nand NAND2 (N14867, N14866, N599);
nor NOR4 (N14868, N14858, N10610, N9738, N9264);
nor NOR4 (N14869, N14863, N3452, N5677, N541);
or OR2 (N14870, N14868, N229);
xor XOR2 (N14871, N14861, N654);
buf BUF1 (N14872, N14862);
xor XOR2 (N14873, N14859, N13690);
and AND4 (N14874, N14873, N7074, N14746, N12616);
buf BUF1 (N14875, N14872);
not NOT1 (N14876, N14856);
not NOT1 (N14877, N14871);
nor NOR3 (N14878, N14870, N2636, N10846);
nor NOR4 (N14879, N14878, N6035, N6860, N5443);
nand NAND2 (N14880, N14867, N5041);
nand NAND2 (N14881, N14877, N11223);
or OR2 (N14882, N14876, N14558);
not NOT1 (N14883, N14879);
or OR3 (N14884, N14850, N14570, N3286);
or OR4 (N14885, N14875, N9970, N14499, N2785);
nor NOR2 (N14886, N14882, N2058);
or OR3 (N14887, N14881, N754, N14444);
nor NOR4 (N14888, N14874, N12673, N3060, N313);
not NOT1 (N14889, N14869);
nor NOR4 (N14890, N14885, N2743, N6032, N13407);
nand NAND4 (N14891, N14890, N4470, N7590, N14340);
nor NOR3 (N14892, N14887, N9455, N1965);
buf BUF1 (N14893, N14880);
not NOT1 (N14894, N14889);
xor XOR2 (N14895, N14864, N11191);
xor XOR2 (N14896, N14893, N6525);
nor NOR4 (N14897, N14884, N13419, N5194, N11772);
and AND3 (N14898, N14865, N12449, N11688);
not NOT1 (N14899, N14896);
and AND3 (N14900, N14899, N6828, N8206);
or OR4 (N14901, N14888, N12975, N9117, N7181);
or OR3 (N14902, N14900, N12011, N9813);
nor NOR2 (N14903, N14894, N9027);
or OR4 (N14904, N14897, N10792, N10020, N5644);
and AND3 (N14905, N14891, N11766, N9752);
not NOT1 (N14906, N14901);
buf BUF1 (N14907, N14906);
and AND2 (N14908, N14903, N1257);
xor XOR2 (N14909, N14898, N13849);
nor NOR2 (N14910, N14907, N4097);
xor XOR2 (N14911, N14886, N7911);
or OR2 (N14912, N14911, N3739);
or OR4 (N14913, N14905, N14811, N11742, N4321);
nor NOR4 (N14914, N14908, N10106, N12891, N13763);
or OR2 (N14915, N14904, N359);
xor XOR2 (N14916, N14913, N2066);
buf BUF1 (N14917, N14892);
and AND4 (N14918, N14895, N11631, N13703, N13977);
xor XOR2 (N14919, N14902, N7126);
nor NOR2 (N14920, N14915, N2872);
not NOT1 (N14921, N14916);
nand NAND4 (N14922, N14921, N4936, N12990, N5635);
nand NAND2 (N14923, N14920, N5705);
xor XOR2 (N14924, N14923, N7104);
nor NOR4 (N14925, N14909, N4280, N9293, N11129);
xor XOR2 (N14926, N14883, N5639);
and AND3 (N14927, N14926, N9695, N7925);
buf BUF1 (N14928, N14919);
not NOT1 (N14929, N14912);
nand NAND2 (N14930, N14914, N7292);
or OR4 (N14931, N14927, N11782, N4244, N10485);
nor NOR4 (N14932, N14930, N13568, N5933, N12900);
buf BUF1 (N14933, N14922);
not NOT1 (N14934, N14929);
nand NAND4 (N14935, N14934, N5672, N3548, N6965);
xor XOR2 (N14936, N14917, N4637);
nor NOR2 (N14937, N14931, N5215);
nand NAND2 (N14938, N14937, N6899);
and AND3 (N14939, N14918, N11705, N10497);
nor NOR4 (N14940, N14932, N13637, N11448, N10188);
and AND4 (N14941, N14935, N9589, N11635, N4162);
or OR4 (N14942, N14928, N10788, N8713, N4144);
nor NOR4 (N14943, N14925, N7619, N13340, N9268);
nor NOR3 (N14944, N14924, N4677, N367);
nor NOR4 (N14945, N14944, N13780, N185, N3753);
and AND2 (N14946, N14943, N13345);
buf BUF1 (N14947, N14936);
not NOT1 (N14948, N14942);
or OR2 (N14949, N14941, N266);
or OR4 (N14950, N14933, N14664, N11329, N495);
nor NOR2 (N14951, N14938, N8815);
nor NOR3 (N14952, N14940, N8839, N5999);
not NOT1 (N14953, N14946);
and AND2 (N14954, N14910, N12425);
xor XOR2 (N14955, N14952, N9483);
xor XOR2 (N14956, N14954, N1933);
xor XOR2 (N14957, N14951, N2138);
nor NOR4 (N14958, N14950, N2704, N1058, N13073);
or OR4 (N14959, N14955, N6263, N4391, N13592);
xor XOR2 (N14960, N14947, N1673);
buf BUF1 (N14961, N14957);
nand NAND4 (N14962, N14948, N9175, N6464, N1019);
not NOT1 (N14963, N14961);
or OR4 (N14964, N14960, N12581, N8849, N3566);
xor XOR2 (N14965, N14956, N7551);
not NOT1 (N14966, N14945);
buf BUF1 (N14967, N14958);
nand NAND3 (N14968, N14964, N9672, N6857);
and AND4 (N14969, N14953, N8660, N6988, N9881);
not NOT1 (N14970, N14939);
nor NOR4 (N14971, N14967, N3107, N7340, N1284);
buf BUF1 (N14972, N14969);
buf BUF1 (N14973, N14949);
nor NOR4 (N14974, N14972, N8794, N13783, N8431);
xor XOR2 (N14975, N14971, N6711);
or OR4 (N14976, N14970, N1122, N577, N10237);
nor NOR2 (N14977, N14962, N10418);
or OR2 (N14978, N14974, N2901);
nor NOR4 (N14979, N14966, N7967, N6045, N425);
or OR4 (N14980, N14973, N2503, N7070, N2780);
xor XOR2 (N14981, N14978, N12748);
buf BUF1 (N14982, N14980);
nor NOR3 (N14983, N14981, N6913, N171);
nor NOR2 (N14984, N14977, N11321);
not NOT1 (N14985, N14984);
or OR4 (N14986, N14982, N2582, N14444, N9241);
nor NOR4 (N14987, N14965, N11189, N11566, N5117);
buf BUF1 (N14988, N14986);
and AND4 (N14989, N14985, N13401, N4107, N6981);
nand NAND2 (N14990, N14988, N14237);
and AND4 (N14991, N14959, N3698, N12171, N5706);
nor NOR4 (N14992, N14987, N8102, N12093, N8884);
nand NAND4 (N14993, N14991, N12868, N9154, N65);
nor NOR3 (N14994, N14983, N11636, N1601);
nor NOR3 (N14995, N14976, N8346, N8023);
not NOT1 (N14996, N14995);
not NOT1 (N14997, N14994);
buf BUF1 (N14998, N14992);
and AND4 (N14999, N14996, N7676, N11609, N6133);
not NOT1 (N15000, N14999);
or OR3 (N15001, N14968, N7554, N12560);
or OR4 (N15002, N14998, N6727, N10154, N11189);
nand NAND2 (N15003, N15000, N1721);
xor XOR2 (N15004, N14975, N8350);
not NOT1 (N15005, N15003);
buf BUF1 (N15006, N14979);
or OR4 (N15007, N15002, N14691, N1419, N13280);
not NOT1 (N15008, N14997);
xor XOR2 (N15009, N15007, N3193);
buf BUF1 (N15010, N14989);
not NOT1 (N15011, N15008);
nor NOR2 (N15012, N15010, N10069);
nand NAND2 (N15013, N15012, N12614);
nor NOR4 (N15014, N14993, N10461, N14132, N13810);
buf BUF1 (N15015, N15006);
or OR2 (N15016, N15009, N12074);
not NOT1 (N15017, N14963);
and AND3 (N15018, N15017, N8635, N1397);
and AND2 (N15019, N15004, N2042);
nand NAND4 (N15020, N15011, N7920, N3836, N7809);
and AND4 (N15021, N15016, N1952, N3088, N6190);
and AND4 (N15022, N15019, N2429, N7681, N13996);
not NOT1 (N15023, N14990);
or OR4 (N15024, N15013, N5472, N8451, N8914);
nor NOR4 (N15025, N15014, N693, N14503, N8266);
or OR3 (N15026, N15025, N431, N5427);
nand NAND2 (N15027, N15026, N9106);
buf BUF1 (N15028, N15001);
and AND4 (N15029, N15020, N10248, N1942, N1205);
or OR3 (N15030, N15023, N1369, N4665);
buf BUF1 (N15031, N15005);
xor XOR2 (N15032, N15030, N5729);
nand NAND2 (N15033, N15028, N11438);
xor XOR2 (N15034, N15027, N12869);
xor XOR2 (N15035, N15015, N12713);
and AND2 (N15036, N15033, N5651);
nand NAND3 (N15037, N15036, N10342, N10004);
buf BUF1 (N15038, N15032);
nand NAND2 (N15039, N15035, N13919);
not NOT1 (N15040, N15038);
nand NAND4 (N15041, N15040, N6149, N3408, N12728);
xor XOR2 (N15042, N15037, N6782);
buf BUF1 (N15043, N15024);
and AND4 (N15044, N15018, N2969, N9244, N1535);
or OR2 (N15045, N15034, N10796);
buf BUF1 (N15046, N15031);
or OR3 (N15047, N15044, N8490, N993);
and AND2 (N15048, N15042, N9698);
xor XOR2 (N15049, N15029, N4402);
nand NAND2 (N15050, N15046, N12647);
nor NOR4 (N15051, N15021, N4756, N5642, N2135);
nor NOR3 (N15052, N15039, N9683, N8652);
nand NAND3 (N15053, N15050, N10416, N13063);
nand NAND3 (N15054, N15045, N3249, N13950);
or OR4 (N15055, N15043, N968, N12073, N9102);
not NOT1 (N15056, N15055);
buf BUF1 (N15057, N15054);
not NOT1 (N15058, N15022);
nand NAND3 (N15059, N15057, N1192, N10368);
and AND2 (N15060, N15056, N1389);
not NOT1 (N15061, N15041);
and AND3 (N15062, N15058, N886, N7171);
nor NOR3 (N15063, N15053, N7947, N2794);
nor NOR3 (N15064, N15051, N4973, N6519);
nor NOR4 (N15065, N15059, N8252, N10870, N1882);
buf BUF1 (N15066, N15065);
and AND3 (N15067, N15061, N8412, N13165);
nand NAND2 (N15068, N15048, N2289);
nor NOR3 (N15069, N15067, N9066, N1411);
not NOT1 (N15070, N15068);
nor NOR3 (N15071, N15063, N13193, N12244);
or OR4 (N15072, N15052, N13817, N5587, N654);
and AND2 (N15073, N15069, N12595);
buf BUF1 (N15074, N15047);
and AND2 (N15075, N15064, N1107);
nor NOR4 (N15076, N15060, N14065, N10827, N9988);
or OR3 (N15077, N15074, N3258, N2574);
buf BUF1 (N15078, N15077);
xor XOR2 (N15079, N15075, N10904);
and AND4 (N15080, N15062, N6336, N1771, N7264);
and AND3 (N15081, N15078, N13814, N12746);
not NOT1 (N15082, N15071);
buf BUF1 (N15083, N15073);
nand NAND3 (N15084, N15076, N2354, N934);
and AND3 (N15085, N15049, N5936, N4432);
xor XOR2 (N15086, N15082, N14474);
nor NOR2 (N15087, N15066, N10767);
buf BUF1 (N15088, N15080);
or OR2 (N15089, N15087, N2647);
nand NAND2 (N15090, N15079, N11358);
nor NOR2 (N15091, N15084, N1487);
nor NOR4 (N15092, N15072, N3810, N11118, N10306);
and AND2 (N15093, N15090, N3826);
not NOT1 (N15094, N15081);
xor XOR2 (N15095, N15089, N7471);
not NOT1 (N15096, N15085);
nor NOR3 (N15097, N15091, N5238, N10468);
nor NOR3 (N15098, N15094, N7028, N2710);
not NOT1 (N15099, N15092);
nand NAND4 (N15100, N15099, N3998, N7595, N9293);
buf BUF1 (N15101, N15100);
xor XOR2 (N15102, N15097, N13616);
xor XOR2 (N15103, N15095, N7607);
nand NAND3 (N15104, N15098, N6284, N9875);
and AND2 (N15105, N15103, N2748);
not NOT1 (N15106, N15086);
and AND3 (N15107, N15093, N8142, N14801);
nand NAND4 (N15108, N15088, N11817, N11866, N9748);
nand NAND2 (N15109, N15105, N4158);
buf BUF1 (N15110, N15108);
xor XOR2 (N15111, N15106, N14821);
and AND4 (N15112, N15111, N9447, N13966, N3150);
not NOT1 (N15113, N15112);
nand NAND4 (N15114, N15101, N5605, N6610, N4587);
buf BUF1 (N15115, N15102);
xor XOR2 (N15116, N15070, N12202);
or OR4 (N15117, N15113, N11037, N3955, N5861);
or OR2 (N15118, N15096, N8663);
and AND3 (N15119, N15110, N2943, N10145);
buf BUF1 (N15120, N15114);
nor NOR4 (N15121, N15118, N798, N8258, N12536);
xor XOR2 (N15122, N15107, N13314);
or OR3 (N15123, N15116, N14388, N3467);
xor XOR2 (N15124, N15083, N5500);
nand NAND3 (N15125, N15121, N13692, N12009);
not NOT1 (N15126, N15124);
xor XOR2 (N15127, N15122, N14444);
and AND2 (N15128, N15109, N1035);
buf BUF1 (N15129, N15119);
nor NOR2 (N15130, N15127, N12789);
nor NOR4 (N15131, N15117, N4873, N6912, N7599);
or OR3 (N15132, N15104, N5599, N7293);
xor XOR2 (N15133, N15132, N8110);
xor XOR2 (N15134, N15115, N5000);
and AND2 (N15135, N15123, N3365);
and AND2 (N15136, N15130, N7310);
buf BUF1 (N15137, N15131);
and AND3 (N15138, N15125, N5732, N9133);
xor XOR2 (N15139, N15137, N8242);
not NOT1 (N15140, N15128);
or OR2 (N15141, N15139, N7090);
and AND2 (N15142, N15136, N4017);
not NOT1 (N15143, N15120);
or OR3 (N15144, N15138, N6921, N11557);
nor NOR2 (N15145, N15143, N10205);
nand NAND3 (N15146, N15133, N10166, N11416);
or OR2 (N15147, N15129, N6383);
and AND3 (N15148, N15134, N8207, N13233);
not NOT1 (N15149, N15135);
nand NAND3 (N15150, N15147, N12864, N13861);
or OR3 (N15151, N15142, N9017, N9903);
and AND4 (N15152, N15148, N13933, N10210, N10065);
not NOT1 (N15153, N15152);
nor NOR3 (N15154, N15126, N2468, N14585);
and AND2 (N15155, N15140, N13378);
buf BUF1 (N15156, N15144);
and AND3 (N15157, N15151, N8986, N7808);
not NOT1 (N15158, N15141);
nand NAND4 (N15159, N15153, N1598, N7557, N10185);
xor XOR2 (N15160, N15155, N9291);
nor NOR3 (N15161, N15158, N12395, N7635);
buf BUF1 (N15162, N15150);
buf BUF1 (N15163, N15149);
not NOT1 (N15164, N15157);
and AND4 (N15165, N15164, N5736, N1714, N14740);
nand NAND2 (N15166, N15159, N3615);
and AND2 (N15167, N15145, N12949);
or OR2 (N15168, N15156, N5966);
xor XOR2 (N15169, N15162, N4369);
nand NAND3 (N15170, N15163, N9299, N11784);
xor XOR2 (N15171, N15168, N7218);
not NOT1 (N15172, N15170);
nor NOR4 (N15173, N15169, N9506, N3310, N8882);
or OR2 (N15174, N15171, N4335);
or OR3 (N15175, N15146, N4913, N5439);
not NOT1 (N15176, N15154);
buf BUF1 (N15177, N15176);
nor NOR3 (N15178, N15165, N12201, N7574);
or OR4 (N15179, N15167, N6642, N9528, N5219);
or OR4 (N15180, N15166, N15126, N7529, N2294);
or OR2 (N15181, N15174, N1345);
and AND4 (N15182, N15181, N1844, N3727, N5649);
buf BUF1 (N15183, N15175);
not NOT1 (N15184, N15178);
buf BUF1 (N15185, N15161);
xor XOR2 (N15186, N15172, N9447);
nor NOR4 (N15187, N15186, N7877, N13373, N10112);
or OR2 (N15188, N15184, N9318);
nor NOR2 (N15189, N15173, N1044);
or OR3 (N15190, N15188, N4794, N3091);
buf BUF1 (N15191, N15179);
buf BUF1 (N15192, N15177);
nand NAND2 (N15193, N15183, N14409);
buf BUF1 (N15194, N15189);
xor XOR2 (N15195, N15182, N14143);
nand NAND3 (N15196, N15191, N6076, N11498);
xor XOR2 (N15197, N15196, N11526);
and AND3 (N15198, N15197, N13537, N15116);
not NOT1 (N15199, N15193);
not NOT1 (N15200, N15180);
buf BUF1 (N15201, N15160);
or OR3 (N15202, N15198, N15054, N8483);
xor XOR2 (N15203, N15194, N1473);
xor XOR2 (N15204, N15199, N3641);
buf BUF1 (N15205, N15185);
and AND2 (N15206, N15195, N8273);
nand NAND2 (N15207, N15206, N1328);
nor NOR3 (N15208, N15205, N13619, N7490);
and AND2 (N15209, N15190, N4597);
xor XOR2 (N15210, N15200, N14755);
or OR4 (N15211, N15209, N10199, N14881, N2617);
nand NAND3 (N15212, N15208, N10128, N6223);
nand NAND3 (N15213, N15204, N8254, N12500);
and AND4 (N15214, N15210, N8621, N11884, N10569);
xor XOR2 (N15215, N15192, N2653);
buf BUF1 (N15216, N15212);
and AND3 (N15217, N15215, N15165, N8086);
not NOT1 (N15218, N15187);
buf BUF1 (N15219, N15213);
nand NAND4 (N15220, N15207, N12389, N11429, N3590);
nor NOR2 (N15221, N15217, N10263);
or OR3 (N15222, N15203, N12222, N6376);
and AND4 (N15223, N15202, N10757, N5556, N10596);
nand NAND4 (N15224, N15214, N5334, N5612, N9677);
not NOT1 (N15225, N15218);
buf BUF1 (N15226, N15223);
or OR2 (N15227, N15226, N8223);
nand NAND2 (N15228, N15221, N1202);
nand NAND2 (N15229, N15211, N9104);
or OR2 (N15230, N15216, N14255);
not NOT1 (N15231, N15224);
and AND3 (N15232, N15220, N10915, N7334);
nand NAND2 (N15233, N15201, N9551);
nor NOR4 (N15234, N15219, N12346, N7526, N4354);
nand NAND3 (N15235, N15227, N5940, N13668);
or OR2 (N15236, N15233, N11215);
xor XOR2 (N15237, N15229, N10706);
nand NAND4 (N15238, N15222, N11464, N11657, N969);
and AND3 (N15239, N15234, N8226, N12313);
xor XOR2 (N15240, N15239, N5202);
and AND2 (N15241, N15232, N5302);
nor NOR4 (N15242, N15230, N8364, N10930, N625);
nand NAND2 (N15243, N15238, N5587);
buf BUF1 (N15244, N15231);
nor NOR2 (N15245, N15235, N5310);
and AND2 (N15246, N15243, N1343);
not NOT1 (N15247, N15237);
buf BUF1 (N15248, N15225);
nand NAND4 (N15249, N15245, N13479, N720, N5383);
xor XOR2 (N15250, N15240, N10241);
or OR4 (N15251, N15249, N12181, N3580, N10810);
not NOT1 (N15252, N15248);
or OR4 (N15253, N15250, N4032, N4206, N2981);
nand NAND3 (N15254, N15247, N1104, N14003);
not NOT1 (N15255, N15252);
not NOT1 (N15256, N15241);
xor XOR2 (N15257, N15251, N13309);
buf BUF1 (N15258, N15257);
buf BUF1 (N15259, N15228);
and AND4 (N15260, N15246, N707, N6853, N9838);
buf BUF1 (N15261, N15244);
and AND4 (N15262, N15258, N11540, N5842, N2447);
and AND2 (N15263, N15253, N567);
nand NAND4 (N15264, N15263, N14591, N8679, N6472);
nor NOR3 (N15265, N15256, N14931, N14175);
xor XOR2 (N15266, N15255, N6207);
and AND2 (N15267, N15254, N13292);
or OR3 (N15268, N15262, N8674, N2740);
and AND3 (N15269, N15266, N14831, N5215);
buf BUF1 (N15270, N15260);
not NOT1 (N15271, N15268);
and AND2 (N15272, N15236, N12734);
nor NOR2 (N15273, N15242, N9235);
nor NOR4 (N15274, N15271, N3552, N2113, N2824);
and AND3 (N15275, N15269, N13078, N3954);
or OR3 (N15276, N15264, N8388, N14442);
not NOT1 (N15277, N15272);
and AND3 (N15278, N15270, N14954, N11465);
and AND4 (N15279, N15275, N8646, N3948, N6542);
nand NAND2 (N15280, N15267, N14298);
not NOT1 (N15281, N15261);
nand NAND2 (N15282, N15265, N14512);
nor NOR4 (N15283, N15278, N2028, N4057, N4373);
or OR4 (N15284, N15274, N10582, N11999, N9177);
and AND4 (N15285, N15279, N13371, N3490, N2674);
buf BUF1 (N15286, N15277);
xor XOR2 (N15287, N15276, N9571);
nor NOR3 (N15288, N15285, N10227, N10262);
not NOT1 (N15289, N15282);
nor NOR2 (N15290, N15288, N14827);
not NOT1 (N15291, N15259);
nand NAND4 (N15292, N15289, N2422, N5071, N11073);
buf BUF1 (N15293, N15280);
or OR2 (N15294, N15287, N13757);
not NOT1 (N15295, N15292);
or OR4 (N15296, N15293, N13911, N5388, N12445);
or OR3 (N15297, N15273, N13319, N8530);
not NOT1 (N15298, N15284);
and AND3 (N15299, N15298, N5388, N7652);
nor NOR2 (N15300, N15281, N5832);
buf BUF1 (N15301, N15294);
not NOT1 (N15302, N15299);
and AND4 (N15303, N15283, N14218, N7701, N12397);
and AND2 (N15304, N15302, N14699);
xor XOR2 (N15305, N15301, N52);
xor XOR2 (N15306, N15291, N14306);
and AND2 (N15307, N15296, N8358);
and AND2 (N15308, N15305, N13482);
xor XOR2 (N15309, N15300, N8487);
xor XOR2 (N15310, N15306, N616);
nand NAND2 (N15311, N15286, N7328);
or OR4 (N15312, N15310, N10995, N1842, N8365);
buf BUF1 (N15313, N15290);
nand NAND3 (N15314, N15297, N12104, N5739);
nor NOR2 (N15315, N15307, N8688);
nand NAND4 (N15316, N15295, N2023, N9126, N4280);
buf BUF1 (N15317, N15313);
xor XOR2 (N15318, N15308, N9076);
not NOT1 (N15319, N15318);
nor NOR3 (N15320, N15304, N3760, N6021);
nor NOR2 (N15321, N15315, N325);
or OR4 (N15322, N15320, N13834, N9344, N2341);
nand NAND2 (N15323, N15314, N13);
or OR2 (N15324, N15323, N13107);
xor XOR2 (N15325, N15311, N5466);
nor NOR4 (N15326, N15324, N4619, N2123, N13317);
buf BUF1 (N15327, N15303);
nand NAND3 (N15328, N15312, N2201, N13196);
nor NOR3 (N15329, N15322, N7676, N6578);
nand NAND2 (N15330, N15326, N10721);
or OR3 (N15331, N15330, N5978, N9977);
nand NAND4 (N15332, N15329, N11696, N13557, N4047);
and AND3 (N15333, N15317, N6500, N2809);
and AND2 (N15334, N15333, N15152);
xor XOR2 (N15335, N15316, N11664);
nand NAND2 (N15336, N15327, N1136);
buf BUF1 (N15337, N15309);
and AND3 (N15338, N15328, N11790, N358);
or OR4 (N15339, N15334, N7450, N14066, N9350);
and AND4 (N15340, N15321, N12283, N5275, N340);
or OR2 (N15341, N15336, N9742);
buf BUF1 (N15342, N15335);
or OR4 (N15343, N15319, N10232, N4040, N9820);
and AND2 (N15344, N15337, N12964);
and AND4 (N15345, N15342, N1812, N6743, N8605);
nand NAND3 (N15346, N15338, N4666, N1705);
not NOT1 (N15347, N15341);
nor NOR3 (N15348, N15344, N10249, N13824);
nand NAND4 (N15349, N15332, N9096, N11068, N630);
not NOT1 (N15350, N15331);
nor NOR2 (N15351, N15325, N7409);
nand NAND4 (N15352, N15339, N2535, N7056, N9292);
xor XOR2 (N15353, N15348, N10812);
buf BUF1 (N15354, N15349);
not NOT1 (N15355, N15346);
buf BUF1 (N15356, N15347);
and AND3 (N15357, N15356, N14764, N3060);
buf BUF1 (N15358, N15345);
buf BUF1 (N15359, N15340);
nor NOR4 (N15360, N15353, N4481, N6812, N1580);
nand NAND4 (N15361, N15350, N3179, N10471, N15324);
nor NOR4 (N15362, N15361, N6522, N3380, N7200);
nor NOR2 (N15363, N15360, N12436);
nor NOR3 (N15364, N15351, N11881, N14630);
not NOT1 (N15365, N15357);
and AND3 (N15366, N15359, N3327, N5438);
xor XOR2 (N15367, N15364, N10900);
nor NOR3 (N15368, N15355, N793, N3494);
buf BUF1 (N15369, N15365);
buf BUF1 (N15370, N15369);
nand NAND4 (N15371, N15370, N2644, N3568, N3944);
not NOT1 (N15372, N15362);
or OR2 (N15373, N15372, N12416);
nand NAND2 (N15374, N15363, N12853);
buf BUF1 (N15375, N15371);
not NOT1 (N15376, N15358);
and AND2 (N15377, N15376, N1582);
nand NAND4 (N15378, N15375, N11099, N13242, N13903);
nand NAND2 (N15379, N15374, N14875);
nand NAND2 (N15380, N15367, N12354);
nor NOR4 (N15381, N15352, N9313, N3822, N3183);
buf BUF1 (N15382, N15366);
and AND2 (N15383, N15354, N13248);
buf BUF1 (N15384, N15373);
buf BUF1 (N15385, N15343);
and AND4 (N15386, N15379, N9058, N13344, N2326);
nand NAND4 (N15387, N15385, N3490, N10194, N14914);
buf BUF1 (N15388, N15384);
xor XOR2 (N15389, N15388, N14179);
xor XOR2 (N15390, N15378, N13089);
or OR3 (N15391, N15390, N6146, N5851);
and AND4 (N15392, N15382, N3024, N2762, N12804);
nor NOR2 (N15393, N15381, N5066);
buf BUF1 (N15394, N15393);
not NOT1 (N15395, N15392);
nand NAND2 (N15396, N15377, N10637);
nor NOR4 (N15397, N15368, N5706, N13146, N12338);
nand NAND4 (N15398, N15396, N70, N10050, N10078);
buf BUF1 (N15399, N15394);
buf BUF1 (N15400, N15391);
or OR3 (N15401, N15395, N7422, N3120);
and AND4 (N15402, N15387, N10681, N4726, N5409);
xor XOR2 (N15403, N15383, N15343);
buf BUF1 (N15404, N15402);
xor XOR2 (N15405, N15398, N4731);
not NOT1 (N15406, N15400);
and AND2 (N15407, N15404, N11639);
xor XOR2 (N15408, N15407, N8736);
nor NOR2 (N15409, N15386, N209);
xor XOR2 (N15410, N15401, N10289);
not NOT1 (N15411, N15408);
xor XOR2 (N15412, N15411, N12783);
nand NAND2 (N15413, N15405, N1202);
nand NAND3 (N15414, N15399, N6964, N11916);
and AND4 (N15415, N15410, N14537, N12729, N12422);
or OR2 (N15416, N15397, N4929);
buf BUF1 (N15417, N15413);
or OR3 (N15418, N15406, N10924, N10515);
and AND3 (N15419, N15380, N15037, N7629);
nor NOR3 (N15420, N15403, N5828, N2241);
xor XOR2 (N15421, N15418, N370);
buf BUF1 (N15422, N15414);
nor NOR2 (N15423, N15415, N5830);
nand NAND3 (N15424, N15389, N13882, N3692);
nand NAND3 (N15425, N15416, N12158, N4602);
not NOT1 (N15426, N15422);
and AND4 (N15427, N15424, N7391, N6686, N12910);
and AND3 (N15428, N15419, N7424, N7638);
buf BUF1 (N15429, N15425);
not NOT1 (N15430, N15421);
xor XOR2 (N15431, N15427, N3439);
not NOT1 (N15432, N15426);
or OR3 (N15433, N15409, N8781, N13166);
not NOT1 (N15434, N15428);
buf BUF1 (N15435, N15432);
buf BUF1 (N15436, N15431);
nand NAND2 (N15437, N15420, N4530);
nor NOR4 (N15438, N15429, N256, N2906, N5897);
or OR4 (N15439, N15430, N4681, N6236, N4061);
nor NOR4 (N15440, N15412, N1534, N5598, N14483);
xor XOR2 (N15441, N15439, N10450);
and AND3 (N15442, N15438, N5082, N14977);
or OR2 (N15443, N15434, N15280);
and AND4 (N15444, N15433, N15283, N12390, N13847);
not NOT1 (N15445, N15443);
and AND2 (N15446, N15437, N1411);
xor XOR2 (N15447, N15446, N9594);
nand NAND4 (N15448, N15417, N5842, N2731, N7465);
or OR4 (N15449, N15436, N5127, N10022, N14411);
buf BUF1 (N15450, N15423);
nor NOR2 (N15451, N15445, N4520);
or OR3 (N15452, N15450, N11025, N13592);
buf BUF1 (N15453, N15444);
nand NAND4 (N15454, N15435, N9586, N4166, N8718);
xor XOR2 (N15455, N15441, N9059);
buf BUF1 (N15456, N15454);
and AND3 (N15457, N15449, N1513, N2205);
not NOT1 (N15458, N15447);
nor NOR2 (N15459, N15455, N13230);
not NOT1 (N15460, N15457);
and AND4 (N15461, N15448, N775, N12683, N13562);
or OR2 (N15462, N15442, N3945);
and AND3 (N15463, N15452, N11137, N420);
nor NOR4 (N15464, N15453, N13088, N7254, N12998);
or OR3 (N15465, N15463, N4832, N12500);
nand NAND4 (N15466, N15462, N13314, N8579, N425);
buf BUF1 (N15467, N15458);
xor XOR2 (N15468, N15456, N10841);
xor XOR2 (N15469, N15451, N62);
nand NAND4 (N15470, N15461, N8762, N470, N2907);
or OR4 (N15471, N15459, N7084, N13690, N9635);
and AND4 (N15472, N15465, N7888, N13605, N4634);
and AND4 (N15473, N15471, N12207, N13397, N3341);
nand NAND3 (N15474, N15472, N9168, N5962);
buf BUF1 (N15475, N15474);
not NOT1 (N15476, N15466);
nand NAND4 (N15477, N15469, N15107, N4415, N11316);
nand NAND4 (N15478, N15475, N4080, N3005, N2409);
xor XOR2 (N15479, N15473, N13715);
xor XOR2 (N15480, N15478, N14626);
buf BUF1 (N15481, N15467);
nor NOR4 (N15482, N15480, N872, N8126, N9518);
or OR4 (N15483, N15470, N8016, N13454, N7288);
nor NOR2 (N15484, N15464, N12494);
or OR2 (N15485, N15440, N2277);
and AND4 (N15486, N15484, N6397, N9347, N7151);
and AND2 (N15487, N15477, N12287);
nor NOR2 (N15488, N15481, N472);
and AND4 (N15489, N15479, N1951, N3872, N1489);
xor XOR2 (N15490, N15460, N4713);
buf BUF1 (N15491, N15483);
xor XOR2 (N15492, N15482, N7143);
xor XOR2 (N15493, N15491, N7629);
nor NOR2 (N15494, N15489, N4993);
xor XOR2 (N15495, N15487, N12205);
and AND3 (N15496, N15490, N2527, N4463);
buf BUF1 (N15497, N15492);
xor XOR2 (N15498, N15497, N9324);
xor XOR2 (N15499, N15476, N1167);
nor NOR4 (N15500, N15486, N225, N14418, N1989);
or OR4 (N15501, N15495, N11355, N7815, N9720);
buf BUF1 (N15502, N15494);
or OR4 (N15503, N15501, N13595, N7774, N14282);
not NOT1 (N15504, N15488);
and AND4 (N15505, N15500, N5256, N10510, N9183);
and AND2 (N15506, N15505, N9466);
not NOT1 (N15507, N15506);
or OR4 (N15508, N15485, N2791, N13495, N3549);
not NOT1 (N15509, N15504);
or OR4 (N15510, N15499, N13137, N4290, N13906);
or OR4 (N15511, N15496, N4916, N4800, N4724);
xor XOR2 (N15512, N15509, N410);
or OR3 (N15513, N15503, N8250, N11461);
buf BUF1 (N15514, N15512);
or OR3 (N15515, N15514, N5489, N2335);
xor XOR2 (N15516, N15510, N5393);
xor XOR2 (N15517, N15516, N2198);
or OR3 (N15518, N15517, N14494, N10340);
or OR2 (N15519, N15507, N1787);
nor NOR2 (N15520, N15468, N3591);
buf BUF1 (N15521, N15513);
nor NOR2 (N15522, N15515, N3031);
nand NAND2 (N15523, N15508, N3858);
xor XOR2 (N15524, N15498, N14558);
nand NAND3 (N15525, N15511, N11699, N5975);
nor NOR2 (N15526, N15522, N76);
and AND4 (N15527, N15519, N6203, N7072, N8442);
and AND2 (N15528, N15524, N2106);
nand NAND3 (N15529, N15528, N2547, N4869);
nand NAND3 (N15530, N15525, N8268, N12886);
buf BUF1 (N15531, N15523);
buf BUF1 (N15532, N15531);
buf BUF1 (N15533, N15532);
nand NAND4 (N15534, N15520, N14212, N11456, N6632);
not NOT1 (N15535, N15493);
and AND4 (N15536, N15529, N968, N1353, N584);
xor XOR2 (N15537, N15535, N9269);
nor NOR2 (N15538, N15502, N12554);
xor XOR2 (N15539, N15518, N15284);
not NOT1 (N15540, N15538);
nor NOR2 (N15541, N15534, N12565);
nor NOR2 (N15542, N15521, N7167);
xor XOR2 (N15543, N15527, N13996);
and AND2 (N15544, N15543, N2849);
xor XOR2 (N15545, N15542, N6355);
nand NAND2 (N15546, N15537, N13670);
or OR2 (N15547, N15533, N13787);
or OR2 (N15548, N15544, N12876);
and AND3 (N15549, N15536, N5338, N7846);
and AND2 (N15550, N15541, N3329);
nand NAND4 (N15551, N15545, N13772, N10334, N11354);
nand NAND4 (N15552, N15526, N7861, N8576, N332);
nand NAND2 (N15553, N15540, N7094);
or OR4 (N15554, N15551, N7169, N8601, N9976);
or OR2 (N15555, N15554, N4087);
or OR4 (N15556, N15549, N5415, N13452, N6043);
buf BUF1 (N15557, N15530);
and AND4 (N15558, N15555, N10552, N11599, N15450);
and AND3 (N15559, N15539, N1832, N10873);
nand NAND2 (N15560, N15557, N2605);
buf BUF1 (N15561, N15546);
and AND2 (N15562, N15560, N12360);
xor XOR2 (N15563, N15548, N14914);
buf BUF1 (N15564, N15553);
not NOT1 (N15565, N15564);
xor XOR2 (N15566, N15562, N4135);
xor XOR2 (N15567, N15556, N11040);
xor XOR2 (N15568, N15563, N7284);
not NOT1 (N15569, N15568);
nand NAND4 (N15570, N15559, N8756, N14447, N6132);
or OR2 (N15571, N15547, N7310);
nand NAND2 (N15572, N15550, N6055);
and AND3 (N15573, N15569, N11779, N9659);
nand NAND2 (N15574, N15571, N3568);
and AND4 (N15575, N15567, N3999, N7685, N2250);
not NOT1 (N15576, N15552);
not NOT1 (N15577, N15573);
buf BUF1 (N15578, N15575);
xor XOR2 (N15579, N15578, N6737);
or OR3 (N15580, N15577, N10187, N4966);
or OR2 (N15581, N15579, N4072);
or OR2 (N15582, N15566, N9966);
and AND3 (N15583, N15558, N5573, N4666);
or OR3 (N15584, N15572, N6039, N6114);
nor NOR2 (N15585, N15574, N1657);
nor NOR4 (N15586, N15561, N3411, N2220, N3459);
xor XOR2 (N15587, N15565, N10220);
not NOT1 (N15588, N15583);
and AND3 (N15589, N15586, N8272, N4752);
or OR2 (N15590, N15584, N15032);
nand NAND3 (N15591, N15576, N14781, N12288);
not NOT1 (N15592, N15570);
and AND2 (N15593, N15582, N10898);
xor XOR2 (N15594, N15591, N15421);
buf BUF1 (N15595, N15587);
not NOT1 (N15596, N15594);
nor NOR3 (N15597, N15595, N4971, N13568);
not NOT1 (N15598, N15593);
xor XOR2 (N15599, N15581, N2915);
and AND4 (N15600, N15588, N5045, N7370, N11041);
nor NOR4 (N15601, N15590, N1963, N15459, N608);
buf BUF1 (N15602, N15600);
not NOT1 (N15603, N15589);
and AND4 (N15604, N15597, N2921, N4082, N10598);
or OR2 (N15605, N15602, N403);
nor NOR3 (N15606, N15604, N11032, N13911);
buf BUF1 (N15607, N15580);
not NOT1 (N15608, N15607);
xor XOR2 (N15609, N15605, N11964);
and AND2 (N15610, N15598, N9591);
and AND3 (N15611, N15606, N2707, N14498);
xor XOR2 (N15612, N15611, N8154);
nor NOR3 (N15613, N15610, N7964, N5855);
xor XOR2 (N15614, N15608, N3964);
not NOT1 (N15615, N15585);
buf BUF1 (N15616, N15603);
not NOT1 (N15617, N15614);
not NOT1 (N15618, N15599);
nor NOR4 (N15619, N15615, N12700, N2606, N8090);
nor NOR2 (N15620, N15601, N8205);
or OR3 (N15621, N15620, N1831, N5151);
xor XOR2 (N15622, N15621, N12041);
or OR2 (N15623, N15616, N677);
xor XOR2 (N15624, N15622, N7830);
nand NAND3 (N15625, N15596, N6549, N14171);
buf BUF1 (N15626, N15625);
not NOT1 (N15627, N15613);
nor NOR3 (N15628, N15592, N9525, N15002);
or OR2 (N15629, N15627, N12102);
buf BUF1 (N15630, N15628);
not NOT1 (N15631, N15609);
or OR3 (N15632, N15612, N4374, N8368);
not NOT1 (N15633, N15631);
buf BUF1 (N15634, N15626);
xor XOR2 (N15635, N15624, N1805);
and AND4 (N15636, N15617, N20, N10306, N13704);
nor NOR4 (N15637, N15618, N15229, N12362, N6624);
and AND4 (N15638, N15632, N8024, N12246, N4025);
and AND3 (N15639, N15619, N15174, N2574);
or OR2 (N15640, N15636, N4838);
xor XOR2 (N15641, N15633, N6011);
nand NAND4 (N15642, N15634, N14680, N3020, N7314);
nand NAND4 (N15643, N15629, N7934, N11044, N12956);
nor NOR3 (N15644, N15638, N8311, N4146);
or OR2 (N15645, N15630, N5201);
or OR4 (N15646, N15635, N1310, N14946, N13769);
buf BUF1 (N15647, N15623);
not NOT1 (N15648, N15639);
not NOT1 (N15649, N15637);
or OR4 (N15650, N15647, N15223, N5358, N13301);
or OR4 (N15651, N15646, N4955, N32, N1185);
and AND3 (N15652, N15642, N2486, N11180);
nor NOR4 (N15653, N15644, N596, N8883, N3158);
nand NAND4 (N15654, N15653, N9766, N123, N857);
and AND3 (N15655, N15654, N1566, N8978);
xor XOR2 (N15656, N15651, N15651);
and AND4 (N15657, N15640, N7696, N12570, N1669);
or OR3 (N15658, N15649, N4766, N1503);
xor XOR2 (N15659, N15655, N2043);
and AND2 (N15660, N15650, N134);
nand NAND2 (N15661, N15641, N2919);
nor NOR3 (N15662, N15660, N3411, N4157);
nand NAND3 (N15663, N15648, N6183, N11630);
not NOT1 (N15664, N15657);
not NOT1 (N15665, N15658);
nand NAND3 (N15666, N15662, N4458, N9017);
not NOT1 (N15667, N15643);
nand NAND3 (N15668, N15645, N6093, N4125);
xor XOR2 (N15669, N15666, N9607);
buf BUF1 (N15670, N15656);
nand NAND4 (N15671, N15670, N8653, N9560, N7636);
or OR4 (N15672, N15671, N9410, N11955, N8030);
nand NAND2 (N15673, N15672, N6460);
nand NAND4 (N15674, N15659, N9312, N11994, N3955);
nand NAND4 (N15675, N15673, N2424, N9430, N1276);
nor NOR3 (N15676, N15675, N5192, N11894);
not NOT1 (N15677, N15669);
nand NAND3 (N15678, N15664, N14193, N309);
and AND3 (N15679, N15678, N1842, N9344);
xor XOR2 (N15680, N15661, N14283);
nand NAND4 (N15681, N15676, N9849, N6632, N1497);
nand NAND2 (N15682, N15663, N4846);
xor XOR2 (N15683, N15679, N7445);
or OR2 (N15684, N15680, N4763);
or OR2 (N15685, N15674, N3209);
and AND3 (N15686, N15685, N1665, N117);
or OR4 (N15687, N15681, N8564, N3150, N3384);
not NOT1 (N15688, N15686);
or OR4 (N15689, N15683, N572, N11086, N12538);
not NOT1 (N15690, N15677);
buf BUF1 (N15691, N15690);
nand NAND3 (N15692, N15684, N10415, N11367);
not NOT1 (N15693, N15652);
or OR3 (N15694, N15667, N2759, N5072);
nor NOR2 (N15695, N15692, N12961);
buf BUF1 (N15696, N15691);
nand NAND2 (N15697, N15693, N418);
nand NAND3 (N15698, N15694, N11471, N10110);
xor XOR2 (N15699, N15689, N8667);
xor XOR2 (N15700, N15682, N2142);
nor NOR2 (N15701, N15700, N11210);
not NOT1 (N15702, N15687);
not NOT1 (N15703, N15702);
buf BUF1 (N15704, N15699);
not NOT1 (N15705, N15703);
nor NOR3 (N15706, N15701, N10833, N10632);
buf BUF1 (N15707, N15706);
not NOT1 (N15708, N15695);
nor NOR4 (N15709, N15665, N4122, N9553, N15590);
and AND4 (N15710, N15697, N8012, N1491, N9949);
buf BUF1 (N15711, N15707);
or OR3 (N15712, N15705, N13462, N1087);
not NOT1 (N15713, N15704);
and AND3 (N15714, N15698, N3463, N9224);
buf BUF1 (N15715, N15713);
and AND4 (N15716, N15696, N5916, N12619, N5343);
nand NAND4 (N15717, N15711, N7231, N15078, N3025);
nor NOR3 (N15718, N15710, N2587, N10444);
nor NOR2 (N15719, N15712, N14617);
nand NAND4 (N15720, N15709, N12492, N200, N3262);
not NOT1 (N15721, N15688);
nor NOR4 (N15722, N15721, N11181, N7544, N5865);
nand NAND2 (N15723, N15717, N10193);
buf BUF1 (N15724, N15715);
buf BUF1 (N15725, N15722);
and AND2 (N15726, N15668, N4237);
nand NAND3 (N15727, N15708, N12510, N33);
not NOT1 (N15728, N15718);
xor XOR2 (N15729, N15726, N13984);
buf BUF1 (N15730, N15725);
not NOT1 (N15731, N15716);
or OR3 (N15732, N15719, N5533, N3406);
and AND4 (N15733, N15724, N10076, N7012, N11244);
nor NOR4 (N15734, N15732, N7313, N4430, N2051);
nand NAND2 (N15735, N15730, N8472);
buf BUF1 (N15736, N15723);
nor NOR4 (N15737, N15734, N13759, N7368, N10217);
xor XOR2 (N15738, N15736, N8887);
nand NAND3 (N15739, N15720, N7098, N13768);
xor XOR2 (N15740, N15735, N12740);
buf BUF1 (N15741, N15738);
buf BUF1 (N15742, N15739);
or OR2 (N15743, N15740, N11346);
xor XOR2 (N15744, N15729, N10447);
buf BUF1 (N15745, N15744);
nand NAND3 (N15746, N15727, N8397, N5084);
not NOT1 (N15747, N15743);
and AND3 (N15748, N15745, N8343, N1427);
and AND2 (N15749, N15714, N2626);
and AND2 (N15750, N15741, N6298);
and AND2 (N15751, N15728, N4617);
nand NAND3 (N15752, N15749, N15522, N1537);
xor XOR2 (N15753, N15747, N7123);
nor NOR3 (N15754, N15753, N5627, N10034);
nand NAND4 (N15755, N15737, N13388, N5507, N6209);
nand NAND3 (N15756, N15751, N2210, N9058);
xor XOR2 (N15757, N15755, N7092);
xor XOR2 (N15758, N15746, N7663);
and AND2 (N15759, N15754, N6200);
nor NOR3 (N15760, N15756, N10243, N9986);
or OR3 (N15761, N15752, N13922, N14125);
and AND2 (N15762, N15759, N14852);
and AND2 (N15763, N15757, N9480);
or OR3 (N15764, N15760, N1090, N14051);
or OR4 (N15765, N15748, N13525, N4357, N6106);
and AND2 (N15766, N15763, N15750);
buf BUF1 (N15767, N7939);
not NOT1 (N15768, N15733);
or OR4 (N15769, N15731, N11466, N11701, N802);
nor NOR2 (N15770, N15758, N4431);
or OR4 (N15771, N15770, N13879, N15183, N6255);
or OR4 (N15772, N15742, N5781, N5654, N8923);
and AND4 (N15773, N15761, N14515, N9023, N14674);
xor XOR2 (N15774, N15767, N10994);
not NOT1 (N15775, N15771);
or OR3 (N15776, N15765, N11226, N7954);
nand NAND4 (N15777, N15764, N8680, N5211, N100);
xor XOR2 (N15778, N15774, N13079);
not NOT1 (N15779, N15768);
xor XOR2 (N15780, N15772, N1556);
nand NAND3 (N15781, N15775, N3718, N14486);
not NOT1 (N15782, N15773);
nor NOR4 (N15783, N15769, N5060, N3803, N1397);
or OR4 (N15784, N15781, N474, N8007, N11715);
and AND3 (N15785, N15776, N14366, N11849);
not NOT1 (N15786, N15784);
or OR3 (N15787, N15786, N7899, N5101);
xor XOR2 (N15788, N15787, N2764);
nand NAND3 (N15789, N15783, N96, N8648);
buf BUF1 (N15790, N15777);
and AND3 (N15791, N15790, N7284, N5715);
or OR2 (N15792, N15782, N12788);
buf BUF1 (N15793, N15778);
xor XOR2 (N15794, N15793, N12161);
or OR2 (N15795, N15789, N13516);
or OR2 (N15796, N15766, N13579);
nor NOR4 (N15797, N15762, N11518, N1956, N9938);
nor NOR3 (N15798, N15796, N3753, N1537);
xor XOR2 (N15799, N15779, N5784);
or OR2 (N15800, N15798, N5687);
not NOT1 (N15801, N15788);
or OR4 (N15802, N15791, N2305, N3987, N1101);
xor XOR2 (N15803, N15795, N6591);
and AND3 (N15804, N15792, N8577, N6802);
not NOT1 (N15805, N15803);
nand NAND4 (N15806, N15804, N10378, N12672, N15054);
not NOT1 (N15807, N15797);
buf BUF1 (N15808, N15785);
and AND2 (N15809, N15807, N2554);
or OR4 (N15810, N15808, N15385, N7982, N6645);
and AND2 (N15811, N15780, N9431);
buf BUF1 (N15812, N15811);
xor XOR2 (N15813, N15800, N15530);
and AND4 (N15814, N15799, N7653, N6378, N159);
and AND2 (N15815, N15809, N13770);
not NOT1 (N15816, N15814);
not NOT1 (N15817, N15802);
buf BUF1 (N15818, N15794);
and AND4 (N15819, N15806, N8605, N13060, N3982);
or OR3 (N15820, N15801, N14327, N6389);
not NOT1 (N15821, N15816);
or OR3 (N15822, N15810, N5836, N12873);
not NOT1 (N15823, N15819);
buf BUF1 (N15824, N15805);
nor NOR4 (N15825, N15822, N8544, N6230, N947);
or OR4 (N15826, N15824, N7174, N584, N9132);
nand NAND2 (N15827, N15815, N14717);
nand NAND4 (N15828, N15821, N15082, N15279, N6457);
not NOT1 (N15829, N15825);
xor XOR2 (N15830, N15820, N6475);
xor XOR2 (N15831, N15818, N11091);
or OR2 (N15832, N15830, N927);
xor XOR2 (N15833, N15827, N4396);
buf BUF1 (N15834, N15817);
or OR4 (N15835, N15833, N10769, N3309, N3754);
or OR3 (N15836, N15829, N6052, N4239);
or OR4 (N15837, N15835, N8409, N4790, N5140);
xor XOR2 (N15838, N15832, N9882);
nor NOR2 (N15839, N15837, N2832);
and AND2 (N15840, N15812, N775);
xor XOR2 (N15841, N15831, N2989);
xor XOR2 (N15842, N15834, N609);
not NOT1 (N15843, N15842);
nand NAND4 (N15844, N15828, N7301, N14208, N9012);
buf BUF1 (N15845, N15836);
nor NOR4 (N15846, N15845, N7529, N2174, N1556);
xor XOR2 (N15847, N15813, N13043);
buf BUF1 (N15848, N15847);
nor NOR4 (N15849, N15839, N11598, N13479, N14734);
and AND4 (N15850, N15841, N24, N6127, N1145);
and AND2 (N15851, N15843, N731);
not NOT1 (N15852, N15826);
xor XOR2 (N15853, N15849, N10916);
or OR3 (N15854, N15848, N8373, N7433);
not NOT1 (N15855, N15850);
buf BUF1 (N15856, N15853);
xor XOR2 (N15857, N15840, N14423);
not NOT1 (N15858, N15854);
nand NAND3 (N15859, N15851, N2470, N10292);
nand NAND2 (N15860, N15856, N13994);
buf BUF1 (N15861, N15855);
or OR4 (N15862, N15852, N2844, N2173, N10421);
buf BUF1 (N15863, N15858);
not NOT1 (N15864, N15861);
buf BUF1 (N15865, N15862);
nand NAND2 (N15866, N15857, N7555);
buf BUF1 (N15867, N15859);
and AND4 (N15868, N15846, N7730, N15268, N14700);
nor NOR2 (N15869, N15867, N9043);
xor XOR2 (N15870, N15863, N10617);
and AND2 (N15871, N15865, N12558);
nand NAND2 (N15872, N15870, N1942);
not NOT1 (N15873, N15860);
and AND3 (N15874, N15873, N5195, N5927);
and AND2 (N15875, N15866, N14488);
nor NOR3 (N15876, N15869, N13359, N8605);
buf BUF1 (N15877, N15844);
buf BUF1 (N15878, N15877);
nand NAND3 (N15879, N15872, N12093, N5305);
or OR4 (N15880, N15878, N2297, N14342, N13035);
nor NOR4 (N15881, N15876, N13729, N2615, N12616);
xor XOR2 (N15882, N15864, N6008);
xor XOR2 (N15883, N15879, N2300);
not NOT1 (N15884, N15874);
or OR4 (N15885, N15883, N10891, N6749, N14742);
nor NOR3 (N15886, N15871, N11032, N2704);
not NOT1 (N15887, N15881);
nor NOR2 (N15888, N15882, N7562);
nand NAND3 (N15889, N15880, N15409, N13063);
xor XOR2 (N15890, N15886, N16);
nor NOR4 (N15891, N15868, N9149, N4140, N14453);
buf BUF1 (N15892, N15838);
or OR3 (N15893, N15884, N7328, N12680);
xor XOR2 (N15894, N15823, N8165);
nor NOR2 (N15895, N15893, N4087);
nor NOR4 (N15896, N15895, N85, N6408, N628);
not NOT1 (N15897, N15890);
xor XOR2 (N15898, N15894, N9758);
or OR2 (N15899, N15887, N7177);
or OR3 (N15900, N15888, N14518, N4081);
buf BUF1 (N15901, N15889);
buf BUF1 (N15902, N15901);
nand NAND4 (N15903, N15897, N14907, N10654, N4440);
not NOT1 (N15904, N15885);
nand NAND4 (N15905, N15904, N15025, N10386, N14813);
not NOT1 (N15906, N15898);
xor XOR2 (N15907, N15896, N3132);
nor NOR2 (N15908, N15905, N15168);
or OR2 (N15909, N15903, N6647);
buf BUF1 (N15910, N15902);
or OR4 (N15911, N15892, N9770, N1717, N10099);
nand NAND4 (N15912, N15891, N5662, N14570, N9078);
nor NOR4 (N15913, N15910, N1884, N12871, N11416);
buf BUF1 (N15914, N15875);
buf BUF1 (N15915, N15900);
xor XOR2 (N15916, N15908, N8495);
buf BUF1 (N15917, N15912);
nor NOR2 (N15918, N15915, N2020);
nand NAND4 (N15919, N15906, N13156, N9200, N3728);
buf BUF1 (N15920, N15914);
xor XOR2 (N15921, N15907, N12392);
not NOT1 (N15922, N15911);
nand NAND4 (N15923, N15919, N5810, N11134, N12170);
nand NAND3 (N15924, N15922, N12872, N5446);
and AND4 (N15925, N15916, N2387, N11078, N7114);
xor XOR2 (N15926, N15909, N13330);
not NOT1 (N15927, N15921);
or OR3 (N15928, N15924, N4318, N5798);
xor XOR2 (N15929, N15927, N3016);
not NOT1 (N15930, N15920);
nand NAND4 (N15931, N15926, N13805, N12731, N2991);
and AND3 (N15932, N15929, N7306, N5863);
xor XOR2 (N15933, N15930, N13446);
xor XOR2 (N15934, N15925, N2019);
nor NOR2 (N15935, N15933, N40);
nor NOR3 (N15936, N15931, N2290, N12692);
not NOT1 (N15937, N15918);
or OR3 (N15938, N15934, N4550, N12718);
or OR4 (N15939, N15917, N13226, N1794, N2659);
xor XOR2 (N15940, N15923, N1005);
nand NAND2 (N15941, N15938, N998);
buf BUF1 (N15942, N15913);
nor NOR4 (N15943, N15941, N15622, N15898, N1883);
and AND4 (N15944, N15937, N6548, N3377, N10359);
xor XOR2 (N15945, N15936, N3719);
and AND4 (N15946, N15944, N4910, N13281, N6268);
and AND3 (N15947, N15928, N4759, N308);
nor NOR2 (N15948, N15899, N12006);
and AND2 (N15949, N15947, N8643);
and AND2 (N15950, N15946, N11241);
nor NOR3 (N15951, N15940, N7782, N7856);
nand NAND4 (N15952, N15943, N13113, N10170, N9502);
buf BUF1 (N15953, N15945);
xor XOR2 (N15954, N15942, N401);
nand NAND4 (N15955, N15949, N11222, N11131, N6629);
xor XOR2 (N15956, N15952, N2373);
and AND3 (N15957, N15954, N5888, N5711);
nor NOR4 (N15958, N15932, N4315, N2649, N5399);
nand NAND4 (N15959, N15935, N8750, N2077, N6688);
nor NOR2 (N15960, N15956, N18);
or OR2 (N15961, N15959, N2866);
buf BUF1 (N15962, N15961);
and AND4 (N15963, N15955, N1970, N14531, N12301);
not NOT1 (N15964, N15957);
xor XOR2 (N15965, N15951, N15273);
nand NAND2 (N15966, N15953, N12479);
nor NOR3 (N15967, N15966, N6872, N7147);
nand NAND4 (N15968, N15962, N3932, N485, N7458);
or OR3 (N15969, N15963, N6996, N4246);
nand NAND2 (N15970, N15960, N12320);
and AND4 (N15971, N15969, N8061, N1600, N6363);
buf BUF1 (N15972, N15965);
xor XOR2 (N15973, N15968, N14782);
nand NAND2 (N15974, N15948, N7133);
or OR3 (N15975, N15974, N1733, N8997);
or OR3 (N15976, N15970, N4916, N15926);
xor XOR2 (N15977, N15964, N1833);
buf BUF1 (N15978, N15958);
buf BUF1 (N15979, N15977);
nor NOR4 (N15980, N15972, N12617, N2206, N6015);
or OR2 (N15981, N15973, N13953);
nor NOR4 (N15982, N15978, N8066, N7479, N15425);
and AND2 (N15983, N15980, N6856);
buf BUF1 (N15984, N15981);
or OR3 (N15985, N15982, N8299, N11618);
or OR3 (N15986, N15967, N2116, N6811);
and AND3 (N15987, N15979, N14398, N7888);
buf BUF1 (N15988, N15985);
xor XOR2 (N15989, N15984, N10153);
not NOT1 (N15990, N15989);
buf BUF1 (N15991, N15971);
not NOT1 (N15992, N15975);
nor NOR2 (N15993, N15986, N7751);
or OR2 (N15994, N15950, N11233);
buf BUF1 (N15995, N15976);
not NOT1 (N15996, N15991);
and AND2 (N15997, N15992, N11956);
and AND4 (N15998, N15993, N14842, N7194, N10046);
or OR2 (N15999, N15983, N10723);
nor NOR3 (N16000, N15990, N173, N7974);
xor XOR2 (N16001, N15987, N13268);
and AND2 (N16002, N15998, N9675);
and AND2 (N16003, N15988, N8572);
buf BUF1 (N16004, N15997);
xor XOR2 (N16005, N16003, N5870);
and AND3 (N16006, N16005, N150, N15606);
not NOT1 (N16007, N16006);
nand NAND2 (N16008, N16004, N8420);
or OR2 (N16009, N16001, N6617);
buf BUF1 (N16010, N15996);
and AND2 (N16011, N15999, N12176);
xor XOR2 (N16012, N16002, N3392);
nand NAND2 (N16013, N16008, N3311);
nor NOR4 (N16014, N16011, N7276, N13735, N13089);
or OR2 (N16015, N15995, N10738);
nor NOR4 (N16016, N16014, N8138, N7550, N9647);
and AND2 (N16017, N16013, N15500);
and AND2 (N16018, N15994, N13216);
xor XOR2 (N16019, N16009, N4285);
endmodule