// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N109,N114,N101,N112,N116,N117,N108,N115,N110,N118;

xor XOR2 (N19, N16, N1);
or OR3 (N20, N10, N12, N12);
not NOT1 (N21, N20);
buf BUF1 (N22, N11);
xor XOR2 (N23, N19, N17);
xor XOR2 (N24, N17, N2);
nand NAND4 (N25, N10, N4, N7, N13);
nor NOR3 (N26, N2, N8, N17);
or OR3 (N27, N8, N14, N24);
buf BUF1 (N28, N26);
or OR4 (N29, N11, N8, N21, N24);
xor XOR2 (N30, N7, N19);
and AND3 (N31, N30, N18, N21);
nand NAND4 (N32, N20, N28, N30, N10);
xor XOR2 (N33, N7, N26);
xor XOR2 (N34, N15, N4);
not NOT1 (N35, N12);
xor XOR2 (N36, N27, N19);
nand NAND3 (N37, N35, N12, N21);
and AND3 (N38, N32, N34, N30);
xor XOR2 (N39, N32, N28);
nand NAND2 (N40, N38, N24);
nor NOR2 (N41, N23, N32);
nor NOR2 (N42, N25, N40);
nand NAND3 (N43, N3, N42, N20);
buf BUF1 (N44, N6);
and AND4 (N45, N44, N14, N3, N18);
or OR3 (N46, N33, N21, N22);
xor XOR2 (N47, N17, N6);
not NOT1 (N48, N37);
nand NAND2 (N49, N41, N12);
not NOT1 (N50, N48);
not NOT1 (N51, N39);
not NOT1 (N52, N43);
xor XOR2 (N53, N31, N34);
buf BUF1 (N54, N45);
nor NOR4 (N55, N29, N51, N24, N36);
buf BUF1 (N56, N2);
xor XOR2 (N57, N51, N40);
buf BUF1 (N58, N54);
buf BUF1 (N59, N52);
nor NOR4 (N60, N50, N37, N3, N49);
not NOT1 (N61, N38);
or OR4 (N62, N46, N46, N46, N1);
or OR2 (N63, N58, N53);
or OR4 (N64, N49, N5, N47, N49);
buf BUF1 (N65, N40);
and AND4 (N66, N57, N40, N17, N35);
or OR2 (N67, N63, N49);
and AND4 (N68, N65, N49, N15, N12);
nor NOR3 (N69, N67, N26, N50);
xor XOR2 (N70, N61, N8);
and AND3 (N71, N60, N64, N29);
nor NOR3 (N72, N58, N69, N19);
or OR2 (N73, N18, N9);
nor NOR2 (N74, N56, N3);
nor NOR4 (N75, N68, N59, N52, N35);
nand NAND4 (N76, N61, N48, N41, N59);
or OR2 (N77, N73, N69);
or OR2 (N78, N77, N50);
not NOT1 (N79, N76);
or OR3 (N80, N66, N52, N79);
buf BUF1 (N81, N50);
nand NAND2 (N82, N75, N45);
nor NOR2 (N83, N71, N19);
or OR4 (N84, N82, N57, N4, N60);
xor XOR2 (N85, N83, N43);
buf BUF1 (N86, N74);
nand NAND3 (N87, N84, N77, N46);
and AND3 (N88, N86, N83, N3);
nor NOR2 (N89, N78, N43);
nand NAND3 (N90, N55, N53, N73);
xor XOR2 (N91, N85, N38);
nand NAND2 (N92, N81, N30);
buf BUF1 (N93, N70);
or OR2 (N94, N90, N6);
not NOT1 (N95, N62);
nor NOR3 (N96, N88, N26, N46);
xor XOR2 (N97, N94, N66);
xor XOR2 (N98, N72, N87);
buf BUF1 (N99, N38);
and AND4 (N100, N89, N3, N48, N42);
or OR4 (N101, N92, N89, N14, N7);
buf BUF1 (N102, N99);
xor XOR2 (N103, N97, N75);
xor XOR2 (N104, N93, N45);
nor NOR4 (N105, N103, N82, N2, N90);
nand NAND4 (N106, N102, N43, N6, N25);
not NOT1 (N107, N91);
buf BUF1 (N108, N106);
xor XOR2 (N109, N98, N38);
and AND3 (N110, N95, N19, N71);
nand NAND3 (N111, N107, N107, N53);
and AND4 (N112, N100, N64, N18, N11);
nand NAND4 (N113, N104, N51, N63, N9);
or OR4 (N114, N105, N53, N50, N9);
xor XOR2 (N115, N80, N11);
xor XOR2 (N116, N96, N46);
or OR4 (N117, N111, N72, N94, N61);
buf BUF1 (N118, N113);
endmodule