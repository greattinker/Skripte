// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N203,N196,N189,N207,N202,N206,N199,N209,N197,N210;

buf BUF1 (N11, N9);
buf BUF1 (N12, N10);
and AND3 (N13, N5, N10, N11);
xor XOR2 (N14, N9, N13);
nor NOR4 (N15, N6, N6, N8, N10);
not NOT1 (N16, N1);
xor XOR2 (N17, N1, N7);
nor NOR4 (N18, N4, N4, N5, N7);
buf BUF1 (N19, N14);
xor XOR2 (N20, N1, N12);
nor NOR2 (N21, N7, N4);
nand NAND3 (N22, N2, N6, N18);
xor XOR2 (N23, N4, N13);
xor XOR2 (N24, N19, N2);
nand NAND3 (N25, N21, N14, N6);
xor XOR2 (N26, N3, N24);
and AND3 (N27, N10, N24, N18);
nand NAND3 (N28, N11, N9, N6);
nor NOR4 (N29, N16, N16, N3, N7);
buf BUF1 (N30, N28);
nand NAND3 (N31, N30, N21, N5);
and AND2 (N32, N25, N20);
buf BUF1 (N33, N1);
or OR3 (N34, N15, N9, N25);
not NOT1 (N35, N22);
nand NAND3 (N36, N33, N9, N14);
nor NOR3 (N37, N26, N7, N7);
nand NAND2 (N38, N32, N28);
xor XOR2 (N39, N35, N34);
nand NAND3 (N40, N13, N20, N19);
not NOT1 (N41, N36);
buf BUF1 (N42, N40);
nor NOR4 (N43, N39, N38, N4, N2);
nand NAND4 (N44, N20, N1, N27, N19);
not NOT1 (N45, N28);
nand NAND2 (N46, N42, N42);
buf BUF1 (N47, N37);
or OR3 (N48, N46, N36, N36);
buf BUF1 (N49, N43);
nand NAND4 (N50, N44, N4, N44, N12);
xor XOR2 (N51, N47, N1);
buf BUF1 (N52, N31);
nor NOR4 (N53, N50, N4, N5, N33);
buf BUF1 (N54, N49);
buf BUF1 (N55, N23);
nor NOR2 (N56, N54, N45);
xor XOR2 (N57, N3, N7);
xor XOR2 (N58, N57, N34);
xor XOR2 (N59, N48, N35);
buf BUF1 (N60, N59);
and AND4 (N61, N52, N59, N56, N29);
buf BUF1 (N62, N24);
xor XOR2 (N63, N42, N31);
xor XOR2 (N64, N62, N62);
nand NAND3 (N65, N64, N54, N21);
buf BUF1 (N66, N65);
nor NOR2 (N67, N53, N20);
buf BUF1 (N68, N55);
not NOT1 (N69, N17);
nand NAND4 (N70, N61, N68, N22, N55);
nor NOR2 (N71, N6, N29);
or OR2 (N72, N60, N29);
buf BUF1 (N73, N72);
nand NAND2 (N74, N51, N60);
and AND2 (N75, N63, N26);
nand NAND4 (N76, N70, N26, N12, N70);
nor NOR3 (N77, N71, N70, N18);
xor XOR2 (N78, N76, N32);
and AND4 (N79, N67, N78, N35, N37);
xor XOR2 (N80, N11, N76);
or OR2 (N81, N77, N23);
and AND4 (N82, N79, N64, N18, N55);
or OR2 (N83, N69, N72);
xor XOR2 (N84, N83, N4);
not NOT1 (N85, N58);
nor NOR3 (N86, N41, N41, N51);
not NOT1 (N87, N74);
nor NOR2 (N88, N82, N65);
nand NAND2 (N89, N87, N52);
nand NAND4 (N90, N80, N62, N89, N42);
or OR2 (N91, N56, N58);
and AND2 (N92, N90, N86);
or OR3 (N93, N87, N66, N82);
not NOT1 (N94, N68);
nand NAND2 (N95, N92, N51);
buf BUF1 (N96, N91);
nand NAND3 (N97, N88, N63, N75);
or OR4 (N98, N66, N55, N82, N15);
buf BUF1 (N99, N96);
nor NOR2 (N100, N95, N29);
or OR4 (N101, N84, N79, N84, N51);
nor NOR2 (N102, N73, N11);
nand NAND4 (N103, N94, N71, N92, N24);
nor NOR2 (N104, N98, N65);
buf BUF1 (N105, N103);
not NOT1 (N106, N100);
nor NOR2 (N107, N102, N11);
or OR4 (N108, N101, N22, N17, N101);
not NOT1 (N109, N85);
nand NAND4 (N110, N99, N89, N44, N65);
nand NAND3 (N111, N97, N85, N29);
and AND3 (N112, N107, N9, N43);
nand NAND3 (N113, N111, N29, N31);
nand NAND3 (N114, N109, N81, N112);
buf BUF1 (N115, N34);
nand NAND3 (N116, N84, N82, N32);
not NOT1 (N117, N105);
nor NOR2 (N118, N108, N18);
and AND2 (N119, N115, N17);
nand NAND2 (N120, N110, N37);
nor NOR3 (N121, N117, N104, N56);
nor NOR3 (N122, N92, N14, N109);
nand NAND4 (N123, N119, N4, N112, N46);
nor NOR4 (N124, N93, N38, N54, N18);
or OR2 (N125, N118, N67);
and AND2 (N126, N116, N24);
xor XOR2 (N127, N120, N85);
and AND2 (N128, N123, N23);
nor NOR3 (N129, N127, N85, N99);
xor XOR2 (N130, N124, N39);
buf BUF1 (N131, N121);
nand NAND4 (N132, N126, N69, N103, N11);
nor NOR2 (N133, N132, N131);
or OR3 (N134, N36, N88, N34);
buf BUF1 (N135, N129);
nand NAND4 (N136, N135, N78, N122, N86);
nand NAND2 (N137, N106, N87);
not NOT1 (N138, N114);
nand NAND3 (N139, N70, N82, N79);
and AND3 (N140, N138, N17, N64);
not NOT1 (N141, N137);
nor NOR2 (N142, N136, N28);
or OR4 (N143, N140, N77, N14, N110);
buf BUF1 (N144, N142);
xor XOR2 (N145, N134, N60);
buf BUF1 (N146, N141);
not NOT1 (N147, N145);
not NOT1 (N148, N146);
or OR4 (N149, N139, N18, N42, N37);
xor XOR2 (N150, N113, N34);
xor XOR2 (N151, N149, N75);
xor XOR2 (N152, N133, N133);
xor XOR2 (N153, N152, N44);
not NOT1 (N154, N153);
and AND4 (N155, N151, N146, N39, N69);
not NOT1 (N156, N154);
nor NOR4 (N157, N128, N77, N100, N118);
xor XOR2 (N158, N150, N66);
buf BUF1 (N159, N158);
or OR2 (N160, N147, N64);
and AND4 (N161, N148, N42, N93, N2);
and AND3 (N162, N160, N95, N3);
nor NOR3 (N163, N155, N151, N71);
not NOT1 (N164, N143);
xor XOR2 (N165, N125, N41);
buf BUF1 (N166, N161);
not NOT1 (N167, N159);
or OR4 (N168, N144, N153, N52, N35);
buf BUF1 (N169, N167);
or OR3 (N170, N169, N85, N47);
or OR3 (N171, N163, N116, N92);
nand NAND2 (N172, N162, N76);
nor NOR3 (N173, N165, N98, N58);
buf BUF1 (N174, N168);
nand NAND4 (N175, N156, N124, N158, N11);
not NOT1 (N176, N130);
or OR2 (N177, N172, N120);
nand NAND2 (N178, N157, N50);
nor NOR3 (N179, N170, N159, N110);
buf BUF1 (N180, N171);
not NOT1 (N181, N180);
not NOT1 (N182, N166);
nor NOR4 (N183, N182, N118, N133, N69);
buf BUF1 (N184, N175);
or OR4 (N185, N183, N53, N143, N92);
buf BUF1 (N186, N173);
buf BUF1 (N187, N178);
and AND2 (N188, N164, N122);
nor NOR4 (N189, N174, N142, N30, N83);
xor XOR2 (N190, N176, N23);
nand NAND4 (N191, N188, N49, N32, N108);
not NOT1 (N192, N177);
or OR2 (N193, N184, N26);
or OR4 (N194, N185, N29, N107, N15);
xor XOR2 (N195, N191, N59);
and AND4 (N196, N179, N54, N127, N132);
not NOT1 (N197, N187);
nand NAND2 (N198, N193, N93);
xor XOR2 (N199, N190, N58);
not NOT1 (N200, N186);
or OR3 (N201, N200, N82, N25);
xor XOR2 (N202, N198, N136);
or OR3 (N203, N201, N73, N66);
not NOT1 (N204, N194);
not NOT1 (N205, N181);
or OR4 (N206, N195, N29, N87, N108);
nor NOR4 (N207, N192, N137, N126, N115);
not NOT1 (N208, N204);
and AND4 (N209, N205, N195, N81, N74);
or OR4 (N210, N208, N5, N93, N143);
endmodule