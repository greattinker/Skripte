// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N3507,N3510,N3498,N3500,N3486,N3499,N3509,N3505,N3511,N3515;

not NOT1 (N16, N2);
not NOT1 (N17, N2);
xor XOR2 (N18, N12, N5);
nand NAND4 (N19, N2, N17, N16, N8);
nor NOR2 (N20, N16, N5);
or OR2 (N21, N12, N5);
buf BUF1 (N22, N13);
not NOT1 (N23, N1);
nand NAND4 (N24, N7, N6, N7, N14);
xor XOR2 (N25, N10, N11);
nand NAND4 (N26, N10, N13, N19, N6);
buf BUF1 (N27, N21);
not NOT1 (N28, N25);
nand NAND4 (N29, N22, N26, N1, N18);
and AND4 (N30, N27, N19, N17, N20);
nand NAND4 (N31, N3, N11, N2, N28);
not NOT1 (N32, N23);
or OR2 (N33, N30, N28);
xor XOR2 (N34, N10, N28);
nand NAND2 (N35, N29, N1);
and AND2 (N36, N26, N20);
buf BUF1 (N37, N3);
nor NOR2 (N38, N35, N17);
xor XOR2 (N39, N1, N20);
or OR4 (N40, N4, N5, N14, N17);
nand NAND3 (N41, N38, N27, N23);
not NOT1 (N42, N31);
not NOT1 (N43, N42);
not NOT1 (N44, N33);
nor NOR2 (N45, N39, N24);
nor NOR4 (N46, N20, N45, N42, N12);
or OR3 (N47, N18, N25, N9);
xor XOR2 (N48, N37, N33);
and AND2 (N49, N46, N11);
nor NOR2 (N50, N47, N23);
not NOT1 (N51, N50);
nor NOR4 (N52, N51, N9, N19, N15);
buf BUF1 (N53, N41);
xor XOR2 (N54, N34, N2);
or OR3 (N55, N52, N39, N27);
nand NAND4 (N56, N54, N28, N3, N26);
or OR3 (N57, N32, N54, N10);
buf BUF1 (N58, N53);
xor XOR2 (N59, N48, N49);
xor XOR2 (N60, N50, N18);
nand NAND4 (N61, N59, N48, N12, N27);
and AND2 (N62, N56, N44);
nand NAND3 (N63, N8, N30, N8);
nor NOR4 (N64, N62, N16, N50, N27);
or OR3 (N65, N60, N55, N8);
xor XOR2 (N66, N17, N37);
and AND2 (N67, N40, N51);
or OR4 (N68, N64, N43, N28, N42);
buf BUF1 (N69, N48);
buf BUF1 (N70, N65);
not NOT1 (N71, N61);
nor NOR3 (N72, N57, N38, N60);
nor NOR3 (N73, N63, N37, N43);
buf BUF1 (N74, N71);
nand NAND4 (N75, N74, N17, N61, N52);
not NOT1 (N76, N68);
or OR2 (N77, N70, N23);
nor NOR3 (N78, N72, N76, N69);
not NOT1 (N79, N36);
buf BUF1 (N80, N12);
and AND2 (N81, N78, N32);
not NOT1 (N82, N70);
and AND3 (N83, N67, N21, N62);
or OR3 (N84, N81, N79, N3);
and AND2 (N85, N33, N71);
xor XOR2 (N86, N77, N22);
xor XOR2 (N87, N75, N2);
nand NAND4 (N88, N83, N67, N64, N10);
nor NOR3 (N89, N84, N14, N63);
not NOT1 (N90, N73);
xor XOR2 (N91, N89, N34);
not NOT1 (N92, N58);
xor XOR2 (N93, N80, N80);
and AND2 (N94, N92, N91);
nor NOR4 (N95, N33, N17, N3, N73);
or OR4 (N96, N85, N33, N33, N56);
nand NAND4 (N97, N87, N90, N91, N36);
and AND4 (N98, N31, N34, N67, N11);
nor NOR2 (N99, N98, N37);
nand NAND3 (N100, N95, N36, N21);
nor NOR4 (N101, N86, N78, N51, N83);
not NOT1 (N102, N96);
buf BUF1 (N103, N97);
nand NAND4 (N104, N101, N8, N67, N57);
xor XOR2 (N105, N82, N4);
not NOT1 (N106, N102);
nor NOR2 (N107, N100, N61);
nand NAND3 (N108, N94, N78, N51);
or OR3 (N109, N103, N36, N105);
and AND4 (N110, N10, N68, N80, N90);
not NOT1 (N111, N99);
and AND3 (N112, N108, N33, N50);
nor NOR4 (N113, N112, N92, N63, N112);
nor NOR4 (N114, N106, N10, N110, N26);
xor XOR2 (N115, N107, N23);
or OR3 (N116, N86, N15, N87);
nor NOR2 (N117, N66, N74);
or OR4 (N118, N104, N106, N34, N58);
or OR2 (N119, N113, N52);
or OR3 (N120, N119, N113, N30);
not NOT1 (N121, N116);
xor XOR2 (N122, N93, N19);
and AND3 (N123, N109, N76, N86);
and AND2 (N124, N111, N118);
not NOT1 (N125, N94);
not NOT1 (N126, N122);
buf BUF1 (N127, N124);
xor XOR2 (N128, N120, N54);
nand NAND4 (N129, N125, N13, N34, N32);
nand NAND2 (N130, N114, N75);
nand NAND3 (N131, N123, N29, N114);
nand NAND4 (N132, N130, N59, N46, N3);
and AND3 (N133, N131, N116, N31);
xor XOR2 (N134, N88, N105);
xor XOR2 (N135, N134, N102);
or OR3 (N136, N128, N37, N33);
buf BUF1 (N137, N132);
or OR3 (N138, N129, N42, N26);
nand NAND3 (N139, N127, N61, N47);
xor XOR2 (N140, N126, N105);
or OR3 (N141, N115, N83, N87);
buf BUF1 (N142, N121);
nor NOR3 (N143, N136, N44, N106);
and AND2 (N144, N140, N125);
or OR4 (N145, N144, N111, N97, N95);
xor XOR2 (N146, N142, N73);
or OR3 (N147, N137, N127, N94);
or OR2 (N148, N133, N131);
not NOT1 (N149, N146);
nor NOR4 (N150, N141, N51, N54, N45);
nor NOR3 (N151, N117, N7, N16);
xor XOR2 (N152, N143, N66);
buf BUF1 (N153, N151);
buf BUF1 (N154, N148);
nor NOR4 (N155, N139, N65, N83, N31);
nand NAND2 (N156, N145, N81);
nand NAND3 (N157, N138, N150, N54);
nor NOR3 (N158, N95, N73, N30);
xor XOR2 (N159, N149, N117);
xor XOR2 (N160, N156, N46);
and AND4 (N161, N155, N25, N121, N49);
not NOT1 (N162, N152);
or OR2 (N163, N161, N155);
and AND4 (N164, N154, N121, N161, N91);
buf BUF1 (N165, N163);
nand NAND4 (N166, N157, N151, N71, N163);
xor XOR2 (N167, N158, N163);
not NOT1 (N168, N167);
nand NAND3 (N169, N166, N123, N53);
and AND2 (N170, N147, N43);
or OR3 (N171, N170, N142, N150);
buf BUF1 (N172, N160);
xor XOR2 (N173, N169, N48);
nand NAND4 (N174, N153, N1, N171, N2);
and AND3 (N175, N43, N41, N59);
nand NAND4 (N176, N165, N68, N27, N69);
buf BUF1 (N177, N173);
nor NOR3 (N178, N172, N47, N53);
and AND4 (N179, N162, N14, N137, N156);
and AND3 (N180, N135, N64, N130);
nor NOR4 (N181, N159, N32, N176, N10);
not NOT1 (N182, N141);
not NOT1 (N183, N179);
buf BUF1 (N184, N177);
or OR4 (N185, N182, N109, N134, N4);
xor XOR2 (N186, N180, N152);
not NOT1 (N187, N164);
not NOT1 (N188, N174);
not NOT1 (N189, N181);
nor NOR4 (N190, N186, N34, N86, N28);
nand NAND2 (N191, N190, N147);
not NOT1 (N192, N189);
xor XOR2 (N193, N175, N40);
xor XOR2 (N194, N188, N134);
buf BUF1 (N195, N183);
buf BUF1 (N196, N187);
or OR3 (N197, N184, N139, N161);
or OR2 (N198, N194, N156);
xor XOR2 (N199, N168, N114);
nor NOR2 (N200, N185, N176);
and AND2 (N201, N197, N182);
xor XOR2 (N202, N199, N30);
xor XOR2 (N203, N191, N162);
or OR2 (N204, N195, N93);
or OR2 (N205, N192, N109);
buf BUF1 (N206, N198);
nand NAND4 (N207, N178, N197, N185, N40);
not NOT1 (N208, N205);
or OR2 (N209, N206, N57);
nand NAND4 (N210, N196, N18, N44, N48);
xor XOR2 (N211, N200, N156);
xor XOR2 (N212, N211, N38);
nor NOR3 (N213, N210, N53, N119);
buf BUF1 (N214, N209);
not NOT1 (N215, N204);
not NOT1 (N216, N207);
buf BUF1 (N217, N216);
nor NOR4 (N218, N208, N33, N35, N134);
and AND2 (N219, N201, N172);
xor XOR2 (N220, N203, N78);
nand NAND2 (N221, N218, N13);
buf BUF1 (N222, N213);
xor XOR2 (N223, N214, N180);
and AND3 (N224, N212, N101, N62);
not NOT1 (N225, N202);
not NOT1 (N226, N193);
and AND3 (N227, N225, N19, N156);
nand NAND3 (N228, N215, N193, N202);
buf BUF1 (N229, N227);
nand NAND4 (N230, N220, N63, N222, N68);
nor NOR4 (N231, N11, N102, N84, N125);
buf BUF1 (N232, N229);
nand NAND4 (N233, N231, N134, N123, N225);
not NOT1 (N234, N233);
or OR3 (N235, N230, N26, N1);
and AND3 (N236, N219, N70, N13);
not NOT1 (N237, N235);
buf BUF1 (N238, N234);
not NOT1 (N239, N237);
not NOT1 (N240, N217);
nand NAND3 (N241, N221, N97, N63);
or OR4 (N242, N236, N92, N170, N52);
xor XOR2 (N243, N226, N40);
not NOT1 (N244, N242);
buf BUF1 (N245, N243);
nand NAND2 (N246, N245, N4);
not NOT1 (N247, N238);
and AND3 (N248, N241, N175, N70);
buf BUF1 (N249, N244);
nor NOR4 (N250, N232, N217, N57, N183);
not NOT1 (N251, N224);
not NOT1 (N252, N250);
not NOT1 (N253, N240);
nor NOR4 (N254, N249, N82, N240, N209);
not NOT1 (N255, N228);
nor NOR3 (N256, N248, N204, N132);
or OR2 (N257, N239, N40);
or OR4 (N258, N246, N27, N242, N73);
buf BUF1 (N259, N254);
nor NOR2 (N260, N251, N206);
buf BUF1 (N261, N258);
nand NAND4 (N262, N247, N52, N165, N110);
and AND3 (N263, N255, N139, N192);
not NOT1 (N264, N256);
nor NOR4 (N265, N260, N241, N81, N119);
and AND4 (N266, N265, N122, N259, N98);
and AND2 (N267, N78, N236);
or OR3 (N268, N262, N234, N195);
nor NOR4 (N269, N263, N172, N25, N28);
or OR3 (N270, N267, N228, N65);
not NOT1 (N271, N268);
nand NAND3 (N272, N264, N94, N224);
and AND3 (N273, N271, N71, N124);
nor NOR4 (N274, N269, N132, N190, N70);
xor XOR2 (N275, N257, N140);
xor XOR2 (N276, N273, N101);
not NOT1 (N277, N270);
not NOT1 (N278, N276);
or OR3 (N279, N275, N84, N16);
nor NOR4 (N280, N278, N269, N51, N217);
nor NOR3 (N281, N253, N15, N222);
or OR3 (N282, N266, N192, N115);
or OR3 (N283, N282, N251, N15);
or OR4 (N284, N280, N169, N50, N163);
nor NOR2 (N285, N284, N61);
nand NAND3 (N286, N277, N256, N197);
buf BUF1 (N287, N281);
nor NOR3 (N288, N287, N120, N165);
not NOT1 (N289, N283);
or OR3 (N290, N288, N112, N82);
or OR2 (N291, N223, N159);
buf BUF1 (N292, N285);
or OR3 (N293, N274, N167, N54);
nand NAND2 (N294, N272, N155);
not NOT1 (N295, N292);
buf BUF1 (N296, N293);
nand NAND3 (N297, N290, N8, N182);
or OR3 (N298, N295, N270, N27);
xor XOR2 (N299, N297, N84);
nor NOR3 (N300, N279, N288, N23);
nor NOR3 (N301, N289, N98, N248);
xor XOR2 (N302, N299, N77);
xor XOR2 (N303, N252, N74);
and AND4 (N304, N301, N203, N222, N237);
and AND4 (N305, N300, N153, N246, N104);
not NOT1 (N306, N286);
and AND3 (N307, N261, N78, N69);
nand NAND2 (N308, N306, N16);
and AND2 (N309, N298, N155);
nand NAND3 (N310, N296, N187, N174);
buf BUF1 (N311, N304);
nor NOR3 (N312, N310, N153, N223);
and AND3 (N313, N302, N305, N291);
or OR4 (N314, N116, N80, N209, N16);
nand NAND2 (N315, N107, N312);
and AND4 (N316, N120, N234, N312, N222);
and AND3 (N317, N308, N291, N13);
and AND3 (N318, N315, N255, N20);
or OR4 (N319, N316, N263, N62, N175);
and AND4 (N320, N311, N195, N306, N241);
not NOT1 (N321, N318);
xor XOR2 (N322, N294, N298);
nand NAND4 (N323, N320, N132, N5, N46);
nor NOR3 (N324, N313, N209, N107);
nand NAND3 (N325, N323, N64, N278);
not NOT1 (N326, N325);
xor XOR2 (N327, N321, N174);
or OR4 (N328, N303, N34, N69, N113);
not NOT1 (N329, N324);
not NOT1 (N330, N326);
nand NAND4 (N331, N330, N323, N305, N215);
nand NAND2 (N332, N328, N85);
xor XOR2 (N333, N332, N272);
xor XOR2 (N334, N327, N327);
nand NAND2 (N335, N322, N255);
or OR2 (N336, N329, N112);
xor XOR2 (N337, N331, N233);
not NOT1 (N338, N314);
nor NOR4 (N339, N337, N161, N54, N129);
buf BUF1 (N340, N317);
xor XOR2 (N341, N334, N245);
buf BUF1 (N342, N333);
nor NOR3 (N343, N309, N102, N58);
nand NAND2 (N344, N336, N289);
nor NOR2 (N345, N343, N177);
nor NOR4 (N346, N342, N27, N341, N174);
xor XOR2 (N347, N231, N297);
and AND3 (N348, N340, N197, N202);
nand NAND3 (N349, N338, N312, N64);
and AND2 (N350, N344, N227);
not NOT1 (N351, N339);
not NOT1 (N352, N351);
xor XOR2 (N353, N319, N235);
and AND4 (N354, N349, N168, N74, N77);
not NOT1 (N355, N353);
nor NOR2 (N356, N335, N21);
nand NAND4 (N357, N352, N217, N68, N191);
nor NOR4 (N358, N347, N23, N53, N226);
or OR4 (N359, N307, N355, N32, N49);
and AND4 (N360, N266, N181, N105, N339);
or OR3 (N361, N356, N79, N35);
nor NOR3 (N362, N359, N314, N263);
buf BUF1 (N363, N361);
xor XOR2 (N364, N357, N250);
not NOT1 (N365, N345);
xor XOR2 (N366, N364, N259);
buf BUF1 (N367, N366);
or OR4 (N368, N358, N327, N132, N18);
or OR3 (N369, N350, N335, N210);
nor NOR3 (N370, N354, N110, N154);
buf BUF1 (N371, N360);
nor NOR2 (N372, N346, N128);
buf BUF1 (N373, N369);
buf BUF1 (N374, N372);
or OR3 (N375, N371, N244, N213);
and AND2 (N376, N348, N106);
xor XOR2 (N377, N365, N64);
and AND4 (N378, N363, N119, N355, N210);
and AND2 (N379, N373, N277);
nor NOR2 (N380, N370, N41);
or OR4 (N381, N378, N284, N52, N47);
buf BUF1 (N382, N380);
and AND4 (N383, N362, N45, N91, N315);
xor XOR2 (N384, N374, N177);
xor XOR2 (N385, N382, N191);
nand NAND2 (N386, N376, N152);
nor NOR2 (N387, N384, N105);
and AND3 (N388, N381, N207, N254);
nand NAND4 (N389, N385, N320, N50, N30);
or OR4 (N390, N389, N61, N230, N58);
nor NOR4 (N391, N383, N122, N312, N175);
and AND2 (N392, N377, N285);
xor XOR2 (N393, N379, N243);
and AND4 (N394, N388, N223, N172, N48);
and AND3 (N395, N375, N305, N261);
xor XOR2 (N396, N394, N52);
or OR3 (N397, N395, N81, N253);
and AND3 (N398, N396, N159, N233);
or OR4 (N399, N391, N346, N389, N324);
nor NOR4 (N400, N367, N329, N392, N69);
or OR4 (N401, N232, N214, N269, N309);
xor XOR2 (N402, N390, N259);
xor XOR2 (N403, N402, N313);
buf BUF1 (N404, N386);
nand NAND3 (N405, N393, N222, N108);
or OR3 (N406, N397, N269, N370);
not NOT1 (N407, N398);
xor XOR2 (N408, N406, N124);
or OR3 (N409, N408, N207, N6);
or OR2 (N410, N409, N366);
nand NAND4 (N411, N368, N340, N182, N390);
nor NOR4 (N412, N400, N17, N196, N233);
and AND2 (N413, N399, N317);
or OR4 (N414, N405, N39, N20, N68);
or OR4 (N415, N401, N156, N143, N179);
and AND3 (N416, N412, N126, N413);
or OR2 (N417, N160, N33);
nand NAND2 (N418, N411, N279);
nor NOR4 (N419, N414, N59, N121, N165);
not NOT1 (N420, N416);
nor NOR2 (N421, N403, N59);
nand NAND2 (N422, N410, N273);
buf BUF1 (N423, N417);
not NOT1 (N424, N415);
not NOT1 (N425, N424);
and AND4 (N426, N420, N68, N336, N318);
not NOT1 (N427, N426);
not NOT1 (N428, N407);
not NOT1 (N429, N428);
nand NAND3 (N430, N423, N336, N69);
xor XOR2 (N431, N425, N232);
and AND4 (N432, N418, N126, N265, N173);
nand NAND3 (N433, N430, N139, N263);
nand NAND3 (N434, N422, N80, N23);
and AND4 (N435, N432, N145, N108, N159);
or OR3 (N436, N433, N232, N198);
xor XOR2 (N437, N429, N283);
nand NAND2 (N438, N436, N176);
nand NAND4 (N439, N434, N374, N338, N359);
not NOT1 (N440, N387);
and AND4 (N441, N431, N299, N87, N26);
buf BUF1 (N442, N435);
and AND3 (N443, N441, N91, N44);
and AND2 (N444, N404, N355);
buf BUF1 (N445, N421);
xor XOR2 (N446, N438, N120);
nor NOR3 (N447, N427, N230, N243);
or OR3 (N448, N419, N100, N401);
buf BUF1 (N449, N440);
nand NAND2 (N450, N442, N28);
not NOT1 (N451, N447);
or OR4 (N452, N444, N6, N225, N234);
not NOT1 (N453, N450);
and AND2 (N454, N452, N8);
not NOT1 (N455, N445);
buf BUF1 (N456, N453);
buf BUF1 (N457, N456);
not NOT1 (N458, N437);
not NOT1 (N459, N454);
not NOT1 (N460, N459);
or OR4 (N461, N460, N253, N73, N50);
xor XOR2 (N462, N457, N67);
or OR3 (N463, N462, N419, N244);
nor NOR3 (N464, N461, N456, N164);
or OR3 (N465, N455, N203, N271);
nand NAND4 (N466, N465, N213, N382, N144);
nor NOR3 (N467, N451, N373, N348);
not NOT1 (N468, N449);
nor NOR2 (N469, N463, N142);
or OR2 (N470, N466, N457);
and AND4 (N471, N468, N185, N361, N128);
and AND3 (N472, N443, N155, N154);
xor XOR2 (N473, N469, N153);
nor NOR2 (N474, N448, N255);
and AND4 (N475, N471, N132, N189, N379);
xor XOR2 (N476, N464, N336);
not NOT1 (N477, N472);
or OR2 (N478, N473, N341);
or OR3 (N479, N475, N38, N35);
not NOT1 (N480, N477);
xor XOR2 (N481, N474, N248);
not NOT1 (N482, N478);
not NOT1 (N483, N481);
nor NOR4 (N484, N470, N391, N404, N461);
or OR3 (N485, N439, N369, N323);
not NOT1 (N486, N479);
nand NAND4 (N487, N458, N183, N323, N155);
or OR4 (N488, N483, N275, N47, N286);
buf BUF1 (N489, N484);
or OR3 (N490, N476, N406, N208);
xor XOR2 (N491, N467, N20);
or OR3 (N492, N485, N144, N82);
buf BUF1 (N493, N488);
nor NOR2 (N494, N489, N74);
nor NOR2 (N495, N487, N369);
buf BUF1 (N496, N494);
and AND4 (N497, N480, N381, N289, N24);
not NOT1 (N498, N486);
or OR2 (N499, N495, N10);
buf BUF1 (N500, N496);
buf BUF1 (N501, N446);
xor XOR2 (N502, N497, N267);
buf BUF1 (N503, N500);
or OR2 (N504, N490, N306);
nor NOR4 (N505, N498, N177, N432, N424);
buf BUF1 (N506, N503);
xor XOR2 (N507, N502, N254);
nor NOR4 (N508, N499, N179, N114, N372);
and AND4 (N509, N482, N450, N331, N124);
nand NAND3 (N510, N507, N137, N354);
buf BUF1 (N511, N506);
not NOT1 (N512, N509);
and AND4 (N513, N491, N364, N492, N480);
and AND4 (N514, N9, N244, N471, N270);
nand NAND3 (N515, N493, N49, N464);
nand NAND2 (N516, N505, N44);
buf BUF1 (N517, N508);
not NOT1 (N518, N515);
or OR3 (N519, N516, N406, N396);
not NOT1 (N520, N513);
buf BUF1 (N521, N519);
nand NAND2 (N522, N514, N179);
not NOT1 (N523, N501);
nand NAND2 (N524, N510, N96);
buf BUF1 (N525, N522);
nor NOR4 (N526, N520, N340, N75, N271);
and AND2 (N527, N525, N64);
buf BUF1 (N528, N512);
xor XOR2 (N529, N528, N33);
or OR3 (N530, N527, N191, N429);
nand NAND2 (N531, N517, N342);
or OR2 (N532, N523, N218);
nand NAND3 (N533, N521, N74, N428);
xor XOR2 (N534, N518, N122);
buf BUF1 (N535, N532);
not NOT1 (N536, N530);
or OR2 (N537, N526, N138);
nor NOR3 (N538, N534, N68, N359);
or OR4 (N539, N537, N55, N414, N235);
nor NOR2 (N540, N533, N232);
or OR4 (N541, N536, N116, N24, N13);
buf BUF1 (N542, N529);
or OR4 (N543, N539, N146, N246, N407);
or OR4 (N544, N540, N185, N405, N397);
and AND4 (N545, N538, N195, N403, N310);
buf BUF1 (N546, N531);
buf BUF1 (N547, N542);
not NOT1 (N548, N511);
xor XOR2 (N549, N546, N439);
nand NAND3 (N550, N504, N46, N58);
nand NAND4 (N551, N550, N419, N52, N7);
nand NAND2 (N552, N545, N165);
buf BUF1 (N553, N535);
not NOT1 (N554, N548);
or OR4 (N555, N554, N425, N537, N438);
not NOT1 (N556, N543);
xor XOR2 (N557, N556, N247);
and AND3 (N558, N524, N86, N59);
and AND2 (N559, N555, N295);
nand NAND3 (N560, N558, N506, N196);
xor XOR2 (N561, N551, N4);
buf BUF1 (N562, N557);
or OR3 (N563, N547, N246, N121);
buf BUF1 (N564, N559);
and AND4 (N565, N541, N214, N92, N315);
buf BUF1 (N566, N563);
or OR4 (N567, N565, N213, N75, N364);
nor NOR4 (N568, N564, N308, N490, N49);
nand NAND3 (N569, N562, N264, N472);
buf BUF1 (N570, N569);
not NOT1 (N571, N544);
or OR2 (N572, N553, N346);
nand NAND2 (N573, N571, N267);
nor NOR4 (N574, N566, N164, N362, N441);
or OR3 (N575, N560, N67, N535);
nand NAND3 (N576, N572, N483, N274);
nor NOR2 (N577, N568, N156);
or OR3 (N578, N549, N115, N531);
nor NOR2 (N579, N574, N466);
xor XOR2 (N580, N578, N259);
and AND3 (N581, N575, N53, N518);
and AND3 (N582, N573, N238, N278);
nand NAND3 (N583, N577, N434, N156);
and AND4 (N584, N570, N189, N479, N31);
and AND4 (N585, N583, N164, N343, N404);
nor NOR2 (N586, N580, N275);
nor NOR3 (N587, N582, N130, N234);
not NOT1 (N588, N552);
not NOT1 (N589, N581);
nand NAND3 (N590, N589, N406, N518);
not NOT1 (N591, N586);
or OR2 (N592, N585, N480);
nand NAND2 (N593, N584, N26);
or OR2 (N594, N591, N556);
nand NAND3 (N595, N594, N496, N83);
nand NAND2 (N596, N592, N283);
buf BUF1 (N597, N596);
or OR4 (N598, N593, N348, N464, N74);
nand NAND2 (N599, N561, N174);
and AND2 (N600, N590, N452);
nand NAND2 (N601, N595, N227);
or OR3 (N602, N567, N483, N548);
nor NOR3 (N603, N599, N139, N121);
nor NOR4 (N604, N576, N225, N380, N560);
nand NAND4 (N605, N579, N333, N257, N14);
nand NAND3 (N606, N600, N101, N234);
buf BUF1 (N607, N587);
nand NAND2 (N608, N607, N567);
not NOT1 (N609, N604);
buf BUF1 (N610, N603);
not NOT1 (N611, N598);
not NOT1 (N612, N597);
nand NAND3 (N613, N605, N356, N568);
buf BUF1 (N614, N611);
not NOT1 (N615, N608);
nand NAND4 (N616, N614, N193, N510, N455);
or OR3 (N617, N606, N68, N548);
and AND4 (N618, N615, N3, N113, N56);
nand NAND4 (N619, N612, N287, N309, N92);
and AND3 (N620, N588, N262, N310);
or OR4 (N621, N601, N211, N184, N463);
or OR3 (N622, N610, N192, N60);
and AND2 (N623, N616, N539);
and AND4 (N624, N619, N337, N297, N374);
or OR2 (N625, N618, N546);
or OR3 (N626, N602, N141, N31);
xor XOR2 (N627, N621, N302);
xor XOR2 (N628, N626, N596);
nand NAND4 (N629, N623, N52, N302, N198);
xor XOR2 (N630, N617, N321);
or OR2 (N631, N609, N287);
nor NOR3 (N632, N630, N577, N622);
nand NAND4 (N633, N33, N434, N234, N375);
or OR3 (N634, N633, N441, N605);
nor NOR4 (N635, N631, N517, N306, N585);
and AND4 (N636, N629, N255, N88, N69);
nand NAND3 (N637, N613, N486, N426);
nor NOR4 (N638, N628, N518, N604, N535);
buf BUF1 (N639, N636);
or OR2 (N640, N625, N608);
nand NAND4 (N641, N624, N198, N58, N299);
nor NOR4 (N642, N632, N300, N22, N628);
and AND4 (N643, N639, N361, N166, N147);
or OR4 (N644, N620, N411, N216, N200);
nand NAND2 (N645, N640, N631);
buf BUF1 (N646, N634);
nand NAND4 (N647, N627, N319, N427, N220);
nand NAND2 (N648, N646, N53);
not NOT1 (N649, N638);
xor XOR2 (N650, N643, N622);
not NOT1 (N651, N637);
nand NAND2 (N652, N648, N253);
and AND3 (N653, N644, N643, N507);
nor NOR4 (N654, N635, N342, N458, N428);
xor XOR2 (N655, N647, N615);
nand NAND2 (N656, N650, N102);
buf BUF1 (N657, N653);
xor XOR2 (N658, N654, N357);
not NOT1 (N659, N645);
not NOT1 (N660, N651);
not NOT1 (N661, N656);
nand NAND4 (N662, N658, N403, N478, N134);
buf BUF1 (N663, N652);
xor XOR2 (N664, N660, N62);
not NOT1 (N665, N657);
and AND4 (N666, N661, N484, N73, N588);
or OR3 (N667, N649, N46, N597);
xor XOR2 (N668, N655, N156);
and AND3 (N669, N664, N171, N539);
nor NOR4 (N670, N669, N598, N192, N453);
nor NOR4 (N671, N666, N616, N340, N537);
xor XOR2 (N672, N667, N356);
not NOT1 (N673, N659);
nor NOR4 (N674, N670, N606, N649, N553);
xor XOR2 (N675, N673, N196);
not NOT1 (N676, N665);
or OR3 (N677, N672, N442, N200);
or OR3 (N678, N677, N210, N166);
nand NAND2 (N679, N675, N430);
nand NAND3 (N680, N668, N412, N584);
xor XOR2 (N681, N674, N501);
nor NOR4 (N682, N679, N411, N393, N529);
and AND4 (N683, N662, N326, N493, N456);
xor XOR2 (N684, N681, N487);
and AND3 (N685, N676, N508, N218);
buf BUF1 (N686, N682);
or OR3 (N687, N678, N114, N142);
xor XOR2 (N688, N687, N686);
nand NAND3 (N689, N214, N487, N215);
nand NAND4 (N690, N680, N609, N556, N307);
buf BUF1 (N691, N671);
buf BUF1 (N692, N688);
not NOT1 (N693, N641);
buf BUF1 (N694, N642);
or OR4 (N695, N683, N3, N387, N387);
buf BUF1 (N696, N689);
or OR4 (N697, N690, N2, N332, N149);
nor NOR4 (N698, N692, N369, N139, N273);
nor NOR2 (N699, N663, N174);
nor NOR3 (N700, N685, N21, N643);
nor NOR4 (N701, N700, N566, N202, N209);
buf BUF1 (N702, N699);
and AND2 (N703, N684, N244);
not NOT1 (N704, N703);
and AND2 (N705, N693, N593);
and AND3 (N706, N694, N46, N555);
not NOT1 (N707, N701);
buf BUF1 (N708, N706);
not NOT1 (N709, N708);
or OR4 (N710, N696, N336, N302, N623);
nor NOR4 (N711, N702, N507, N204, N641);
nor NOR4 (N712, N697, N16, N565, N484);
or OR4 (N713, N695, N15, N146, N522);
xor XOR2 (N714, N691, N523);
nor NOR4 (N715, N704, N672, N592, N97);
nand NAND3 (N716, N712, N564, N439);
xor XOR2 (N717, N707, N135);
nand NAND4 (N718, N716, N498, N59, N530);
xor XOR2 (N719, N713, N572);
nor NOR3 (N720, N698, N173, N540);
nor NOR2 (N721, N720, N467);
nand NAND3 (N722, N710, N282, N225);
and AND4 (N723, N714, N334, N291, N718);
nand NAND3 (N724, N291, N40, N399);
or OR3 (N725, N719, N487, N28);
xor XOR2 (N726, N717, N30);
nor NOR2 (N727, N723, N711);
nor NOR4 (N728, N578, N400, N682, N409);
or OR4 (N729, N721, N340, N58, N118);
and AND4 (N730, N705, N237, N637, N655);
not NOT1 (N731, N729);
or OR2 (N732, N725, N624);
buf BUF1 (N733, N732);
nor NOR3 (N734, N731, N561, N461);
buf BUF1 (N735, N726);
nand NAND3 (N736, N709, N407, N271);
not NOT1 (N737, N727);
nand NAND2 (N738, N724, N149);
and AND4 (N739, N730, N360, N203, N412);
not NOT1 (N740, N722);
buf BUF1 (N741, N734);
xor XOR2 (N742, N740, N157);
and AND2 (N743, N715, N27);
not NOT1 (N744, N741);
or OR2 (N745, N733, N420);
buf BUF1 (N746, N728);
xor XOR2 (N747, N735, N615);
or OR3 (N748, N746, N49, N374);
nand NAND3 (N749, N738, N620, N208);
nand NAND4 (N750, N743, N504, N678, N480);
xor XOR2 (N751, N742, N663);
nand NAND2 (N752, N739, N135);
and AND2 (N753, N747, N530);
or OR4 (N754, N752, N512, N660, N363);
nand NAND3 (N755, N754, N738, N421);
xor XOR2 (N756, N744, N187);
nor NOR2 (N757, N745, N435);
buf BUF1 (N758, N753);
or OR3 (N759, N748, N661, N285);
nor NOR4 (N760, N757, N203, N137, N53);
xor XOR2 (N761, N749, N750);
buf BUF1 (N762, N175);
nor NOR2 (N763, N758, N409);
and AND2 (N764, N756, N725);
or OR2 (N765, N764, N631);
nand NAND3 (N766, N751, N542, N73);
xor XOR2 (N767, N755, N144);
or OR4 (N768, N767, N244, N215, N322);
and AND2 (N769, N760, N224);
not NOT1 (N770, N765);
not NOT1 (N771, N737);
not NOT1 (N772, N736);
or OR4 (N773, N770, N112, N276, N736);
nand NAND2 (N774, N763, N634);
buf BUF1 (N775, N774);
or OR3 (N776, N773, N125, N409);
nand NAND4 (N777, N768, N329, N485, N758);
nor NOR3 (N778, N762, N523, N445);
and AND4 (N779, N771, N548, N318, N340);
not NOT1 (N780, N779);
or OR3 (N781, N769, N474, N457);
buf BUF1 (N782, N759);
not NOT1 (N783, N766);
and AND4 (N784, N776, N383, N89, N463);
nor NOR4 (N785, N783, N621, N650, N605);
nand NAND4 (N786, N782, N330, N572, N533);
nand NAND2 (N787, N775, N106);
nand NAND2 (N788, N778, N282);
xor XOR2 (N789, N787, N373);
not NOT1 (N790, N784);
nand NAND2 (N791, N790, N701);
or OR2 (N792, N777, N196);
buf BUF1 (N793, N786);
xor XOR2 (N794, N791, N598);
xor XOR2 (N795, N794, N319);
and AND3 (N796, N761, N105, N781);
nand NAND2 (N797, N614, N239);
nor NOR2 (N798, N792, N130);
and AND4 (N799, N788, N178, N58, N83);
nand NAND3 (N800, N797, N157, N592);
and AND4 (N801, N800, N249, N329, N219);
not NOT1 (N802, N801);
and AND4 (N803, N795, N209, N45, N330);
nand NAND4 (N804, N799, N548, N384, N478);
xor XOR2 (N805, N804, N557);
nor NOR2 (N806, N789, N345);
and AND4 (N807, N802, N101, N693, N460);
and AND2 (N808, N803, N16);
xor XOR2 (N809, N772, N360);
buf BUF1 (N810, N806);
or OR3 (N811, N807, N39, N142);
nand NAND4 (N812, N811, N169, N301, N276);
or OR2 (N813, N809, N211);
or OR4 (N814, N805, N629, N71, N788);
xor XOR2 (N815, N796, N284);
buf BUF1 (N816, N812);
nor NOR4 (N817, N815, N250, N503, N100);
or OR3 (N818, N817, N139, N454);
nand NAND2 (N819, N816, N793);
nand NAND3 (N820, N494, N281, N233);
not NOT1 (N821, N785);
xor XOR2 (N822, N821, N799);
not NOT1 (N823, N780);
nand NAND2 (N824, N814, N792);
or OR4 (N825, N808, N710, N219, N60);
xor XOR2 (N826, N820, N806);
xor XOR2 (N827, N819, N369);
and AND3 (N828, N826, N226, N239);
nand NAND2 (N829, N798, N733);
nand NAND3 (N830, N825, N124, N485);
not NOT1 (N831, N810);
nor NOR4 (N832, N829, N264, N167, N756);
not NOT1 (N833, N813);
nor NOR3 (N834, N831, N266, N599);
nand NAND3 (N835, N832, N93, N567);
or OR4 (N836, N835, N441, N680, N576);
buf BUF1 (N837, N822);
or OR4 (N838, N830, N140, N335, N203);
and AND2 (N839, N834, N201);
nor NOR4 (N840, N838, N501, N800, N515);
or OR4 (N841, N839, N191, N57, N209);
and AND2 (N842, N836, N403);
and AND4 (N843, N827, N201, N795, N32);
buf BUF1 (N844, N843);
buf BUF1 (N845, N818);
not NOT1 (N846, N842);
nor NOR4 (N847, N828, N141, N192, N806);
buf BUF1 (N848, N833);
nor NOR3 (N849, N844, N269, N415);
or OR4 (N850, N845, N50, N796, N788);
or OR2 (N851, N824, N497);
nand NAND2 (N852, N841, N594);
or OR2 (N853, N823, N289);
buf BUF1 (N854, N853);
nor NOR2 (N855, N846, N812);
xor XOR2 (N856, N855, N157);
xor XOR2 (N857, N847, N355);
nand NAND3 (N858, N857, N564, N413);
and AND2 (N859, N852, N194);
nor NOR4 (N860, N848, N400, N608, N329);
xor XOR2 (N861, N856, N475);
buf BUF1 (N862, N860);
not NOT1 (N863, N840);
not NOT1 (N864, N858);
not NOT1 (N865, N849);
nor NOR2 (N866, N861, N252);
buf BUF1 (N867, N865);
not NOT1 (N868, N859);
or OR4 (N869, N868, N265, N67, N13);
or OR2 (N870, N851, N24);
not NOT1 (N871, N854);
not NOT1 (N872, N837);
and AND4 (N873, N867, N201, N863, N819);
xor XOR2 (N874, N667, N487);
nand NAND3 (N875, N850, N191, N379);
nor NOR3 (N876, N872, N407, N191);
nand NAND4 (N877, N871, N255, N232, N191);
and AND4 (N878, N866, N468, N181, N622);
nand NAND2 (N879, N877, N152);
xor XOR2 (N880, N878, N380);
or OR3 (N881, N880, N54, N585);
buf BUF1 (N882, N864);
not NOT1 (N883, N879);
xor XOR2 (N884, N862, N815);
and AND4 (N885, N870, N349, N436, N129);
xor XOR2 (N886, N876, N422);
or OR2 (N887, N869, N678);
or OR4 (N888, N873, N159, N789, N624);
nor NOR2 (N889, N888, N12);
not NOT1 (N890, N874);
and AND2 (N891, N886, N631);
not NOT1 (N892, N884);
and AND4 (N893, N889, N315, N588, N730);
or OR2 (N894, N891, N86);
and AND3 (N895, N875, N2, N30);
not NOT1 (N896, N894);
and AND2 (N897, N895, N721);
buf BUF1 (N898, N890);
nand NAND3 (N899, N896, N703, N597);
not NOT1 (N900, N892);
and AND3 (N901, N900, N746, N785);
and AND4 (N902, N881, N432, N493, N630);
not NOT1 (N903, N882);
nor NOR3 (N904, N899, N389, N870);
buf BUF1 (N905, N901);
and AND2 (N906, N893, N904);
not NOT1 (N907, N71);
nor NOR3 (N908, N898, N173, N903);
nor NOR2 (N909, N374, N424);
and AND4 (N910, N909, N401, N667, N29);
not NOT1 (N911, N887);
not NOT1 (N912, N906);
xor XOR2 (N913, N912, N750);
nor NOR4 (N914, N911, N272, N136, N577);
and AND4 (N915, N908, N810, N864, N735);
xor XOR2 (N916, N907, N93);
not NOT1 (N917, N910);
nor NOR3 (N918, N897, N92, N704);
not NOT1 (N919, N916);
nand NAND4 (N920, N883, N728, N533, N913);
xor XOR2 (N921, N559, N23);
nor NOR3 (N922, N917, N443, N628);
or OR2 (N923, N919, N771);
xor XOR2 (N924, N905, N797);
nand NAND3 (N925, N920, N682, N195);
xor XOR2 (N926, N925, N254);
and AND2 (N927, N885, N292);
or OR3 (N928, N914, N650, N924);
and AND3 (N929, N912, N415, N547);
buf BUF1 (N930, N923);
buf BUF1 (N931, N930);
nor NOR3 (N932, N926, N361, N68);
or OR3 (N933, N927, N177, N186);
xor XOR2 (N934, N933, N285);
not NOT1 (N935, N932);
nor NOR2 (N936, N915, N681);
not NOT1 (N937, N931);
nor NOR4 (N938, N936, N323, N147, N470);
xor XOR2 (N939, N928, N884);
nor NOR4 (N940, N938, N246, N449, N483);
not NOT1 (N941, N918);
nor NOR4 (N942, N929, N334, N654, N21);
and AND4 (N943, N921, N749, N514, N742);
buf BUF1 (N944, N943);
nor NOR2 (N945, N937, N711);
nor NOR3 (N946, N934, N294, N724);
xor XOR2 (N947, N939, N657);
and AND4 (N948, N942, N199, N249, N459);
nor NOR4 (N949, N945, N207, N524, N860);
and AND2 (N950, N922, N533);
nor NOR2 (N951, N902, N566);
or OR2 (N952, N951, N188);
nand NAND4 (N953, N952, N780, N922, N237);
nand NAND2 (N954, N949, N522);
not NOT1 (N955, N953);
nor NOR4 (N956, N950, N189, N653, N460);
and AND3 (N957, N947, N205, N173);
and AND3 (N958, N957, N554, N746);
not NOT1 (N959, N944);
nand NAND4 (N960, N940, N569, N876, N896);
nor NOR4 (N961, N941, N308, N115, N532);
not NOT1 (N962, N959);
xor XOR2 (N963, N955, N872);
and AND3 (N964, N958, N723, N564);
xor XOR2 (N965, N954, N196);
not NOT1 (N966, N963);
nor NOR2 (N967, N935, N827);
or OR3 (N968, N967, N711, N635);
not NOT1 (N969, N964);
xor XOR2 (N970, N962, N405);
nand NAND4 (N971, N946, N606, N653, N529);
nor NOR3 (N972, N969, N180, N953);
nand NAND3 (N973, N966, N298, N674);
and AND2 (N974, N968, N50);
and AND3 (N975, N965, N399, N931);
nor NOR4 (N976, N971, N530, N498, N424);
not NOT1 (N977, N972);
nor NOR3 (N978, N975, N883, N926);
not NOT1 (N979, N956);
and AND3 (N980, N948, N545, N896);
and AND2 (N981, N973, N403);
buf BUF1 (N982, N970);
or OR4 (N983, N976, N72, N269, N731);
xor XOR2 (N984, N982, N527);
nor NOR2 (N985, N977, N675);
or OR3 (N986, N984, N55, N105);
buf BUF1 (N987, N981);
or OR3 (N988, N980, N879, N815);
xor XOR2 (N989, N985, N236);
buf BUF1 (N990, N974);
xor XOR2 (N991, N987, N244);
or OR3 (N992, N988, N750, N541);
nor NOR3 (N993, N986, N442, N413);
not NOT1 (N994, N961);
or OR2 (N995, N993, N194);
xor XOR2 (N996, N990, N623);
nor NOR4 (N997, N991, N101, N727, N717);
buf BUF1 (N998, N995);
and AND3 (N999, N994, N904, N23);
buf BUF1 (N1000, N999);
buf BUF1 (N1001, N960);
not NOT1 (N1002, N978);
not NOT1 (N1003, N979);
not NOT1 (N1004, N1003);
nor NOR3 (N1005, N989, N980, N75);
xor XOR2 (N1006, N1004, N328);
buf BUF1 (N1007, N983);
xor XOR2 (N1008, N1007, N239);
xor XOR2 (N1009, N1000, N768);
and AND4 (N1010, N1005, N437, N539, N903);
not NOT1 (N1011, N997);
nor NOR3 (N1012, N998, N616, N224);
buf BUF1 (N1013, N1002);
nand NAND2 (N1014, N1010, N157);
buf BUF1 (N1015, N1009);
or OR2 (N1016, N1001, N793);
xor XOR2 (N1017, N992, N99);
buf BUF1 (N1018, N1008);
not NOT1 (N1019, N1012);
or OR2 (N1020, N996, N568);
or OR4 (N1021, N1020, N420, N137, N883);
nor NOR3 (N1022, N1013, N550, N80);
not NOT1 (N1023, N1022);
not NOT1 (N1024, N1018);
nor NOR3 (N1025, N1024, N716, N375);
not NOT1 (N1026, N1023);
and AND2 (N1027, N1015, N804);
buf BUF1 (N1028, N1017);
xor XOR2 (N1029, N1011, N225);
and AND2 (N1030, N1025, N421);
or OR2 (N1031, N1029, N343);
not NOT1 (N1032, N1014);
buf BUF1 (N1033, N1027);
and AND2 (N1034, N1021, N819);
buf BUF1 (N1035, N1032);
or OR4 (N1036, N1031, N56, N437, N951);
or OR2 (N1037, N1036, N802);
and AND2 (N1038, N1026, N207);
and AND4 (N1039, N1033, N224, N438, N1023);
and AND4 (N1040, N1030, N499, N890, N593);
xor XOR2 (N1041, N1019, N664);
nor NOR2 (N1042, N1006, N609);
nor NOR2 (N1043, N1035, N888);
xor XOR2 (N1044, N1041, N701);
nor NOR3 (N1045, N1044, N785, N446);
xor XOR2 (N1046, N1037, N999);
not NOT1 (N1047, N1028);
nor NOR3 (N1048, N1046, N166, N150);
xor XOR2 (N1049, N1045, N728);
and AND4 (N1050, N1049, N875, N129, N933);
and AND3 (N1051, N1040, N446, N776);
or OR4 (N1052, N1042, N566, N665, N120);
xor XOR2 (N1053, N1016, N270);
nor NOR4 (N1054, N1052, N141, N462, N163);
and AND4 (N1055, N1048, N728, N1049, N826);
or OR2 (N1056, N1053, N386);
nor NOR4 (N1057, N1038, N687, N411, N827);
nand NAND2 (N1058, N1047, N249);
or OR4 (N1059, N1057, N220, N585, N820);
nor NOR4 (N1060, N1043, N306, N878, N849);
xor XOR2 (N1061, N1050, N968);
and AND2 (N1062, N1059, N189);
nor NOR4 (N1063, N1058, N128, N397, N740);
and AND3 (N1064, N1061, N364, N1022);
and AND4 (N1065, N1056, N517, N762, N567);
or OR4 (N1066, N1064, N193, N361, N127);
and AND4 (N1067, N1063, N401, N729, N391);
or OR4 (N1068, N1065, N675, N418, N667);
nor NOR4 (N1069, N1055, N514, N806, N4);
xor XOR2 (N1070, N1068, N355);
and AND2 (N1071, N1060, N564);
nand NAND4 (N1072, N1039, N991, N18, N1070);
nor NOR3 (N1073, N522, N903, N188);
xor XOR2 (N1074, N1054, N80);
nand NAND4 (N1075, N1051, N272, N927, N119);
xor XOR2 (N1076, N1067, N1);
buf BUF1 (N1077, N1072);
or OR2 (N1078, N1076, N622);
and AND4 (N1079, N1071, N63, N365, N635);
xor XOR2 (N1080, N1077, N165);
xor XOR2 (N1081, N1062, N106);
buf BUF1 (N1082, N1080);
xor XOR2 (N1083, N1081, N110);
or OR3 (N1084, N1078, N231, N1080);
nor NOR4 (N1085, N1079, N211, N882, N1055);
buf BUF1 (N1086, N1069);
and AND4 (N1087, N1066, N380, N322, N768);
or OR4 (N1088, N1075, N75, N1022, N63);
or OR2 (N1089, N1086, N706);
xor XOR2 (N1090, N1084, N754);
or OR4 (N1091, N1087, N151, N99, N926);
nor NOR2 (N1092, N1090, N318);
or OR2 (N1093, N1088, N400);
xor XOR2 (N1094, N1085, N427);
nor NOR2 (N1095, N1094, N165);
and AND3 (N1096, N1095, N838, N431);
not NOT1 (N1097, N1092);
or OR4 (N1098, N1082, N238, N234, N387);
nand NAND2 (N1099, N1073, N346);
not NOT1 (N1100, N1099);
nand NAND3 (N1101, N1034, N916, N375);
nor NOR2 (N1102, N1074, N701);
nand NAND4 (N1103, N1098, N118, N788, N597);
or OR4 (N1104, N1093, N984, N572, N96);
buf BUF1 (N1105, N1103);
and AND2 (N1106, N1104, N629);
not NOT1 (N1107, N1096);
nand NAND3 (N1108, N1089, N903, N361);
nand NAND4 (N1109, N1108, N542, N1108, N780);
not NOT1 (N1110, N1091);
nand NAND2 (N1111, N1100, N395);
nand NAND4 (N1112, N1102, N832, N1024, N260);
xor XOR2 (N1113, N1111, N1068);
or OR4 (N1114, N1107, N720, N717, N938);
nand NAND4 (N1115, N1101, N816, N458, N58);
buf BUF1 (N1116, N1105);
and AND2 (N1117, N1097, N1108);
nand NAND2 (N1118, N1106, N153);
xor XOR2 (N1119, N1112, N597);
or OR2 (N1120, N1083, N213);
and AND4 (N1121, N1119, N267, N61, N122);
buf BUF1 (N1122, N1115);
nor NOR2 (N1123, N1116, N289);
buf BUF1 (N1124, N1122);
not NOT1 (N1125, N1114);
and AND2 (N1126, N1113, N347);
xor XOR2 (N1127, N1120, N481);
nor NOR2 (N1128, N1127, N410);
nor NOR3 (N1129, N1118, N737, N1068);
nor NOR3 (N1130, N1124, N660, N760);
xor XOR2 (N1131, N1123, N128);
nand NAND2 (N1132, N1121, N970);
nand NAND3 (N1133, N1125, N510, N439);
and AND2 (N1134, N1126, N442);
and AND4 (N1135, N1132, N428, N430, N110);
nor NOR2 (N1136, N1109, N1130);
xor XOR2 (N1137, N610, N487);
not NOT1 (N1138, N1131);
nand NAND4 (N1139, N1129, N885, N861, N305);
nor NOR3 (N1140, N1128, N935, N325);
or OR4 (N1141, N1136, N811, N397, N139);
nand NAND4 (N1142, N1139, N319, N977, N637);
not NOT1 (N1143, N1138);
not NOT1 (N1144, N1143);
or OR4 (N1145, N1140, N424, N913, N412);
or OR2 (N1146, N1137, N1144);
nand NAND2 (N1147, N413, N28);
not NOT1 (N1148, N1133);
not NOT1 (N1149, N1148);
not NOT1 (N1150, N1147);
nor NOR4 (N1151, N1135, N505, N622, N669);
not NOT1 (N1152, N1117);
nand NAND2 (N1153, N1152, N586);
nor NOR4 (N1154, N1134, N527, N1034, N1124);
xor XOR2 (N1155, N1150, N21);
nand NAND3 (N1156, N1149, N1142, N712);
xor XOR2 (N1157, N1043, N1126);
xor XOR2 (N1158, N1141, N6);
nor NOR4 (N1159, N1157, N1029, N919, N727);
nor NOR2 (N1160, N1159, N252);
or OR4 (N1161, N1151, N125, N123, N460);
or OR4 (N1162, N1161, N856, N584, N453);
not NOT1 (N1163, N1158);
and AND2 (N1164, N1110, N480);
or OR4 (N1165, N1156, N8, N413, N877);
and AND4 (N1166, N1165, N538, N40, N641);
buf BUF1 (N1167, N1164);
buf BUF1 (N1168, N1155);
nand NAND3 (N1169, N1154, N392, N340);
nor NOR4 (N1170, N1153, N289, N1099, N287);
not NOT1 (N1171, N1162);
nand NAND2 (N1172, N1166, N482);
not NOT1 (N1173, N1146);
nor NOR3 (N1174, N1160, N199, N926);
nand NAND2 (N1175, N1169, N121);
xor XOR2 (N1176, N1173, N278);
or OR3 (N1177, N1168, N668, N292);
nand NAND2 (N1178, N1170, N1051);
nor NOR2 (N1179, N1167, N118);
xor XOR2 (N1180, N1179, N1093);
and AND2 (N1181, N1178, N1131);
not NOT1 (N1182, N1176);
xor XOR2 (N1183, N1180, N1074);
buf BUF1 (N1184, N1171);
nand NAND3 (N1185, N1184, N170, N76);
buf BUF1 (N1186, N1183);
xor XOR2 (N1187, N1186, N263);
xor XOR2 (N1188, N1182, N924);
nor NOR4 (N1189, N1185, N803, N70, N355);
buf BUF1 (N1190, N1188);
xor XOR2 (N1191, N1190, N181);
buf BUF1 (N1192, N1174);
xor XOR2 (N1193, N1192, N1116);
not NOT1 (N1194, N1177);
not NOT1 (N1195, N1194);
nand NAND2 (N1196, N1175, N698);
nand NAND3 (N1197, N1172, N390, N411);
and AND2 (N1198, N1163, N654);
and AND3 (N1199, N1187, N284, N538);
xor XOR2 (N1200, N1193, N140);
or OR3 (N1201, N1181, N36, N55);
not NOT1 (N1202, N1198);
nor NOR4 (N1203, N1197, N553, N141, N591);
nor NOR4 (N1204, N1196, N940, N905, N440);
not NOT1 (N1205, N1199);
or OR3 (N1206, N1191, N794, N469);
xor XOR2 (N1207, N1204, N1045);
buf BUF1 (N1208, N1205);
buf BUF1 (N1209, N1200);
or OR3 (N1210, N1189, N575, N1189);
not NOT1 (N1211, N1201);
not NOT1 (N1212, N1211);
xor XOR2 (N1213, N1208, N827);
nor NOR2 (N1214, N1195, N1208);
not NOT1 (N1215, N1209);
xor XOR2 (N1216, N1210, N275);
xor XOR2 (N1217, N1145, N1001);
buf BUF1 (N1218, N1217);
not NOT1 (N1219, N1213);
nand NAND3 (N1220, N1203, N578, N104);
nor NOR3 (N1221, N1206, N18, N1003);
xor XOR2 (N1222, N1221, N290);
or OR3 (N1223, N1219, N1209, N614);
and AND3 (N1224, N1216, N14, N1121);
xor XOR2 (N1225, N1202, N313);
nand NAND2 (N1226, N1214, N1166);
not NOT1 (N1227, N1212);
or OR4 (N1228, N1226, N605, N1056, N678);
buf BUF1 (N1229, N1224);
and AND2 (N1230, N1207, N485);
xor XOR2 (N1231, N1228, N269);
xor XOR2 (N1232, N1229, N1149);
xor XOR2 (N1233, N1230, N279);
nor NOR3 (N1234, N1218, N1146, N997);
or OR2 (N1235, N1227, N856);
or OR4 (N1236, N1231, N479, N387, N359);
nand NAND2 (N1237, N1222, N552);
xor XOR2 (N1238, N1237, N587);
nand NAND3 (N1239, N1225, N1148, N484);
not NOT1 (N1240, N1235);
not NOT1 (N1241, N1238);
nand NAND2 (N1242, N1240, N890);
or OR4 (N1243, N1239, N234, N1053, N575);
and AND3 (N1244, N1220, N85, N590);
and AND3 (N1245, N1233, N746, N1010);
not NOT1 (N1246, N1241);
xor XOR2 (N1247, N1234, N1110);
xor XOR2 (N1248, N1244, N1170);
nand NAND3 (N1249, N1248, N254, N354);
xor XOR2 (N1250, N1223, N176);
or OR4 (N1251, N1232, N711, N1117, N596);
and AND3 (N1252, N1245, N686, N785);
not NOT1 (N1253, N1249);
nand NAND2 (N1254, N1253, N1035);
nor NOR2 (N1255, N1251, N146);
nand NAND2 (N1256, N1246, N1081);
xor XOR2 (N1257, N1247, N943);
not NOT1 (N1258, N1236);
buf BUF1 (N1259, N1215);
not NOT1 (N1260, N1242);
and AND4 (N1261, N1257, N473, N445, N4);
nor NOR2 (N1262, N1260, N367);
nor NOR2 (N1263, N1262, N925);
xor XOR2 (N1264, N1243, N387);
nor NOR3 (N1265, N1252, N662, N673);
xor XOR2 (N1266, N1261, N72);
nand NAND4 (N1267, N1254, N256, N963, N943);
not NOT1 (N1268, N1266);
nor NOR2 (N1269, N1256, N646);
and AND3 (N1270, N1265, N647, N1025);
nand NAND3 (N1271, N1270, N1155, N328);
nor NOR4 (N1272, N1255, N797, N51, N143);
and AND4 (N1273, N1258, N654, N754, N1052);
or OR3 (N1274, N1264, N74, N179);
or OR4 (N1275, N1259, N62, N751, N672);
not NOT1 (N1276, N1274);
nand NAND2 (N1277, N1271, N350);
or OR2 (N1278, N1263, N929);
not NOT1 (N1279, N1269);
and AND4 (N1280, N1278, N1000, N743, N989);
nor NOR2 (N1281, N1267, N294);
not NOT1 (N1282, N1277);
or OR2 (N1283, N1281, N523);
or OR2 (N1284, N1282, N1160);
xor XOR2 (N1285, N1279, N1001);
xor XOR2 (N1286, N1284, N261);
nand NAND3 (N1287, N1275, N940, N1229);
xor XOR2 (N1288, N1276, N607);
and AND2 (N1289, N1283, N1185);
xor XOR2 (N1290, N1250, N493);
nor NOR4 (N1291, N1288, N597, N804, N1062);
nand NAND2 (N1292, N1289, N1155);
nor NOR3 (N1293, N1287, N296, N329);
nor NOR4 (N1294, N1291, N398, N1087, N1261);
buf BUF1 (N1295, N1286);
nor NOR2 (N1296, N1290, N612);
nor NOR4 (N1297, N1272, N968, N366, N77);
not NOT1 (N1298, N1280);
or OR3 (N1299, N1268, N1033, N158);
nand NAND4 (N1300, N1285, N204, N1281, N1040);
not NOT1 (N1301, N1293);
nor NOR4 (N1302, N1300, N118, N1043, N788);
not NOT1 (N1303, N1294);
buf BUF1 (N1304, N1302);
not NOT1 (N1305, N1301);
xor XOR2 (N1306, N1273, N249);
xor XOR2 (N1307, N1306, N7);
or OR4 (N1308, N1297, N1158, N1229, N702);
nor NOR3 (N1309, N1292, N851, N279);
nand NAND3 (N1310, N1299, N806, N169);
not NOT1 (N1311, N1310);
not NOT1 (N1312, N1305);
nand NAND2 (N1313, N1308, N978);
or OR3 (N1314, N1303, N531, N162);
nand NAND2 (N1315, N1307, N768);
nand NAND3 (N1316, N1312, N1203, N344);
or OR4 (N1317, N1313, N973, N172, N701);
xor XOR2 (N1318, N1317, N799);
and AND2 (N1319, N1314, N274);
xor XOR2 (N1320, N1298, N554);
xor XOR2 (N1321, N1309, N1316);
buf BUF1 (N1322, N923);
and AND2 (N1323, N1321, N39);
or OR2 (N1324, N1295, N1152);
nand NAND4 (N1325, N1311, N140, N846, N887);
or OR3 (N1326, N1324, N172, N297);
nand NAND4 (N1327, N1322, N193, N393, N371);
buf BUF1 (N1328, N1304);
xor XOR2 (N1329, N1296, N4);
buf BUF1 (N1330, N1320);
buf BUF1 (N1331, N1325);
nor NOR3 (N1332, N1328, N1162, N1052);
buf BUF1 (N1333, N1329);
or OR4 (N1334, N1332, N601, N1018, N153);
nand NAND4 (N1335, N1331, N556, N126, N1098);
xor XOR2 (N1336, N1318, N188);
and AND3 (N1337, N1327, N855, N277);
or OR2 (N1338, N1336, N1171);
buf BUF1 (N1339, N1330);
or OR3 (N1340, N1334, N1040, N54);
nor NOR4 (N1341, N1335, N1026, N668, N13);
xor XOR2 (N1342, N1323, N477);
or OR4 (N1343, N1341, N981, N71, N1227);
nand NAND3 (N1344, N1340, N451, N1077);
not NOT1 (N1345, N1344);
xor XOR2 (N1346, N1333, N1209);
and AND2 (N1347, N1346, N1002);
nor NOR4 (N1348, N1338, N217, N640, N1192);
or OR4 (N1349, N1339, N249, N772, N618);
xor XOR2 (N1350, N1343, N415);
nand NAND2 (N1351, N1348, N58);
nor NOR3 (N1352, N1326, N233, N982);
nor NOR2 (N1353, N1342, N973);
nor NOR3 (N1354, N1319, N1107, N95);
nand NAND3 (N1355, N1351, N235, N508);
nor NOR3 (N1356, N1353, N1298, N1325);
not NOT1 (N1357, N1356);
or OR2 (N1358, N1350, N72);
not NOT1 (N1359, N1354);
nand NAND2 (N1360, N1357, N1293);
nor NOR3 (N1361, N1359, N727, N14);
buf BUF1 (N1362, N1352);
not NOT1 (N1363, N1360);
nor NOR3 (N1364, N1349, N356, N1154);
or OR3 (N1365, N1347, N922, N1081);
xor XOR2 (N1366, N1315, N957);
xor XOR2 (N1367, N1345, N428);
xor XOR2 (N1368, N1362, N75);
buf BUF1 (N1369, N1367);
nand NAND3 (N1370, N1369, N932, N561);
nand NAND4 (N1371, N1370, N381, N726, N42);
and AND2 (N1372, N1368, N901);
buf BUF1 (N1373, N1355);
not NOT1 (N1374, N1358);
or OR3 (N1375, N1361, N581, N785);
xor XOR2 (N1376, N1372, N516);
buf BUF1 (N1377, N1337);
not NOT1 (N1378, N1374);
xor XOR2 (N1379, N1376, N1275);
or OR3 (N1380, N1363, N1299, N1325);
buf BUF1 (N1381, N1366);
or OR2 (N1382, N1365, N1194);
or OR4 (N1383, N1379, N1353, N1265, N496);
buf BUF1 (N1384, N1383);
xor XOR2 (N1385, N1373, N1094);
buf BUF1 (N1386, N1381);
nor NOR3 (N1387, N1386, N674, N546);
buf BUF1 (N1388, N1387);
nor NOR4 (N1389, N1377, N620, N1214, N599);
xor XOR2 (N1390, N1389, N553);
xor XOR2 (N1391, N1371, N1037);
or OR2 (N1392, N1375, N1076);
or OR4 (N1393, N1382, N894, N284, N825);
xor XOR2 (N1394, N1391, N610);
buf BUF1 (N1395, N1392);
or OR4 (N1396, N1380, N857, N727, N526);
nand NAND2 (N1397, N1385, N897);
not NOT1 (N1398, N1390);
nor NOR4 (N1399, N1396, N1048, N95, N873);
xor XOR2 (N1400, N1398, N696);
buf BUF1 (N1401, N1400);
and AND2 (N1402, N1395, N236);
xor XOR2 (N1403, N1397, N993);
nand NAND3 (N1404, N1378, N379, N609);
nor NOR3 (N1405, N1384, N829, N1014);
nor NOR3 (N1406, N1403, N705, N1298);
or OR2 (N1407, N1399, N1196);
and AND2 (N1408, N1405, N472);
xor XOR2 (N1409, N1402, N856);
buf BUF1 (N1410, N1401);
or OR3 (N1411, N1394, N574, N1243);
or OR3 (N1412, N1408, N1063, N1224);
and AND4 (N1413, N1404, N397, N1388, N1144);
and AND4 (N1414, N864, N667, N1041, N1312);
not NOT1 (N1415, N1412);
buf BUF1 (N1416, N1364);
and AND4 (N1417, N1415, N365, N172, N184);
or OR2 (N1418, N1410, N325);
or OR2 (N1419, N1414, N1272);
or OR4 (N1420, N1418, N986, N486, N571);
or OR3 (N1421, N1393, N149, N948);
and AND4 (N1422, N1421, N933, N783, N1063);
or OR4 (N1423, N1420, N720, N102, N887);
nand NAND3 (N1424, N1419, N2, N346);
buf BUF1 (N1425, N1407);
or OR3 (N1426, N1413, N1343, N908);
xor XOR2 (N1427, N1422, N3);
and AND2 (N1428, N1416, N1252);
xor XOR2 (N1429, N1423, N777);
and AND2 (N1430, N1426, N1333);
not NOT1 (N1431, N1424);
buf BUF1 (N1432, N1409);
or OR4 (N1433, N1427, N137, N736, N263);
buf BUF1 (N1434, N1430);
and AND4 (N1435, N1434, N1433, N907, N195);
nor NOR4 (N1436, N1048, N739, N939, N863);
nand NAND3 (N1437, N1417, N214, N733);
or OR2 (N1438, N1435, N50);
and AND2 (N1439, N1438, N1145);
or OR4 (N1440, N1431, N835, N1257, N18);
nor NOR2 (N1441, N1425, N266);
or OR4 (N1442, N1406, N710, N198, N41);
nor NOR3 (N1443, N1428, N126, N199);
nor NOR4 (N1444, N1442, N708, N638, N863);
not NOT1 (N1445, N1411);
not NOT1 (N1446, N1444);
nor NOR4 (N1447, N1429, N238, N379, N504);
or OR3 (N1448, N1445, N1193, N1437);
not NOT1 (N1449, N245);
and AND4 (N1450, N1441, N1287, N1273, N675);
nand NAND3 (N1451, N1447, N373, N1131);
nand NAND4 (N1452, N1451, N190, N36, N450);
nand NAND2 (N1453, N1443, N772);
not NOT1 (N1454, N1450);
and AND2 (N1455, N1432, N848);
and AND3 (N1456, N1449, N1428, N1412);
not NOT1 (N1457, N1439);
nor NOR2 (N1458, N1440, N1011);
or OR2 (N1459, N1453, N420);
nand NAND2 (N1460, N1458, N1162);
nand NAND3 (N1461, N1452, N413, N932);
and AND2 (N1462, N1459, N100);
and AND2 (N1463, N1454, N539);
xor XOR2 (N1464, N1461, N1146);
nand NAND3 (N1465, N1446, N534, N127);
nor NOR3 (N1466, N1448, N1119, N975);
buf BUF1 (N1467, N1465);
or OR3 (N1468, N1460, N517, N1325);
nand NAND4 (N1469, N1462, N465, N1325, N210);
xor XOR2 (N1470, N1466, N441);
not NOT1 (N1471, N1436);
and AND3 (N1472, N1456, N575, N519);
and AND4 (N1473, N1457, N463, N479, N1144);
and AND4 (N1474, N1463, N207, N497, N1337);
and AND2 (N1475, N1473, N865);
and AND4 (N1476, N1470, N505, N1047, N364);
nand NAND2 (N1477, N1471, N452);
nand NAND3 (N1478, N1476, N649, N735);
nand NAND4 (N1479, N1478, N178, N76, N769);
and AND3 (N1480, N1468, N1273, N15);
nand NAND2 (N1481, N1475, N518);
not NOT1 (N1482, N1477);
xor XOR2 (N1483, N1479, N1367);
buf BUF1 (N1484, N1455);
and AND3 (N1485, N1467, N273, N1153);
nor NOR3 (N1486, N1483, N176, N641);
nand NAND4 (N1487, N1472, N982, N831, N1273);
xor XOR2 (N1488, N1482, N287);
and AND4 (N1489, N1481, N491, N267, N440);
nand NAND4 (N1490, N1488, N1170, N443, N1225);
nand NAND3 (N1491, N1486, N539, N1215);
and AND2 (N1492, N1485, N760);
buf BUF1 (N1493, N1464);
or OR2 (N1494, N1490, N627);
or OR3 (N1495, N1487, N541, N1320);
xor XOR2 (N1496, N1474, N883);
xor XOR2 (N1497, N1489, N1164);
buf BUF1 (N1498, N1480);
buf BUF1 (N1499, N1469);
xor XOR2 (N1500, N1497, N1479);
nor NOR3 (N1501, N1491, N671, N1294);
and AND2 (N1502, N1492, N1250);
buf BUF1 (N1503, N1494);
xor XOR2 (N1504, N1493, N603);
not NOT1 (N1505, N1504);
and AND4 (N1506, N1484, N978, N147, N432);
nand NAND3 (N1507, N1502, N1061, N40);
buf BUF1 (N1508, N1498);
and AND2 (N1509, N1506, N550);
not NOT1 (N1510, N1503);
nand NAND4 (N1511, N1500, N965, N528, N285);
nor NOR3 (N1512, N1511, N1399, N1468);
xor XOR2 (N1513, N1510, N1161);
nand NAND4 (N1514, N1495, N19, N63, N261);
buf BUF1 (N1515, N1508);
nand NAND3 (N1516, N1509, N1418, N1509);
buf BUF1 (N1517, N1514);
nor NOR3 (N1518, N1499, N451, N479);
and AND4 (N1519, N1512, N255, N1242, N582);
buf BUF1 (N1520, N1501);
and AND4 (N1521, N1513, N413, N250, N1463);
buf BUF1 (N1522, N1505);
xor XOR2 (N1523, N1515, N478);
and AND3 (N1524, N1496, N391, N313);
nor NOR2 (N1525, N1523, N925);
nand NAND4 (N1526, N1516, N1187, N1402, N124);
xor XOR2 (N1527, N1522, N145);
nand NAND4 (N1528, N1517, N221, N196, N1442);
not NOT1 (N1529, N1519);
xor XOR2 (N1530, N1526, N248);
buf BUF1 (N1531, N1524);
and AND3 (N1532, N1528, N900, N99);
xor XOR2 (N1533, N1518, N1311);
buf BUF1 (N1534, N1521);
not NOT1 (N1535, N1520);
not NOT1 (N1536, N1533);
and AND2 (N1537, N1525, N1063);
and AND4 (N1538, N1527, N1409, N709, N1346);
nor NOR3 (N1539, N1537, N884, N1461);
nand NAND2 (N1540, N1534, N333);
buf BUF1 (N1541, N1532);
nand NAND4 (N1542, N1538, N1253, N1151, N911);
nor NOR2 (N1543, N1540, N1019);
xor XOR2 (N1544, N1536, N1111);
xor XOR2 (N1545, N1541, N840);
or OR3 (N1546, N1535, N915, N343);
not NOT1 (N1547, N1546);
nor NOR3 (N1548, N1530, N1344, N959);
nand NAND3 (N1549, N1507, N774, N1379);
xor XOR2 (N1550, N1544, N778);
nand NAND3 (N1551, N1543, N983, N1037);
nor NOR3 (N1552, N1531, N54, N1504);
nand NAND3 (N1553, N1549, N1521, N284);
or OR3 (N1554, N1542, N1248, N680);
and AND2 (N1555, N1547, N949);
or OR4 (N1556, N1545, N673, N1043, N1409);
or OR3 (N1557, N1556, N807, N1105);
nand NAND3 (N1558, N1548, N32, N1133);
and AND2 (N1559, N1539, N1548);
nor NOR3 (N1560, N1555, N241, N352);
and AND2 (N1561, N1551, N1147);
not NOT1 (N1562, N1554);
buf BUF1 (N1563, N1561);
and AND4 (N1564, N1558, N789, N527, N1529);
nor NOR2 (N1565, N1540, N1177);
not NOT1 (N1566, N1563);
not NOT1 (N1567, N1557);
and AND2 (N1568, N1564, N298);
nand NAND4 (N1569, N1560, N864, N1278, N1416);
or OR2 (N1570, N1567, N1535);
nand NAND2 (N1571, N1552, N1346);
xor XOR2 (N1572, N1562, N1425);
nor NOR3 (N1573, N1565, N368, N501);
nor NOR3 (N1574, N1550, N724, N864);
xor XOR2 (N1575, N1569, N182);
not NOT1 (N1576, N1553);
and AND2 (N1577, N1559, N869);
or OR4 (N1578, N1575, N1037, N954, N975);
xor XOR2 (N1579, N1573, N10);
nand NAND2 (N1580, N1572, N1576);
buf BUF1 (N1581, N1010);
and AND2 (N1582, N1578, N687);
and AND3 (N1583, N1566, N1483, N629);
not NOT1 (N1584, N1570);
xor XOR2 (N1585, N1577, N756);
not NOT1 (N1586, N1568);
buf BUF1 (N1587, N1579);
nand NAND3 (N1588, N1574, N1276, N741);
and AND2 (N1589, N1584, N728);
xor XOR2 (N1590, N1581, N1206);
or OR2 (N1591, N1571, N87);
not NOT1 (N1592, N1586);
nand NAND4 (N1593, N1589, N1544, N906, N662);
buf BUF1 (N1594, N1585);
and AND2 (N1595, N1583, N1100);
or OR4 (N1596, N1594, N1218, N1412, N267);
and AND4 (N1597, N1592, N773, N1072, N1221);
nor NOR4 (N1598, N1580, N1317, N1220, N9);
and AND4 (N1599, N1595, N39, N1330, N354);
nand NAND4 (N1600, N1591, N901, N1477, N214);
buf BUF1 (N1601, N1588);
and AND3 (N1602, N1601, N33, N788);
buf BUF1 (N1603, N1600);
buf BUF1 (N1604, N1596);
not NOT1 (N1605, N1593);
not NOT1 (N1606, N1603);
or OR2 (N1607, N1605, N158);
nand NAND3 (N1608, N1607, N889, N34);
nand NAND2 (N1609, N1598, N1494);
or OR4 (N1610, N1606, N439, N262, N845);
not NOT1 (N1611, N1608);
xor XOR2 (N1612, N1587, N1464);
and AND2 (N1613, N1597, N1453);
nand NAND3 (N1614, N1609, N1021, N179);
or OR4 (N1615, N1614, N651, N1132, N356);
and AND3 (N1616, N1602, N651, N414);
or OR3 (N1617, N1599, N1303, N1086);
not NOT1 (N1618, N1615);
xor XOR2 (N1619, N1611, N645);
xor XOR2 (N1620, N1613, N28);
buf BUF1 (N1621, N1612);
nand NAND4 (N1622, N1604, N1115, N469, N861);
not NOT1 (N1623, N1610);
not NOT1 (N1624, N1616);
buf BUF1 (N1625, N1623);
buf BUF1 (N1626, N1590);
not NOT1 (N1627, N1620);
and AND3 (N1628, N1625, N1501, N765);
or OR3 (N1629, N1626, N120, N1432);
not NOT1 (N1630, N1582);
buf BUF1 (N1631, N1618);
buf BUF1 (N1632, N1619);
nor NOR2 (N1633, N1631, N127);
xor XOR2 (N1634, N1622, N846);
nand NAND4 (N1635, N1630, N1460, N215, N1294);
nor NOR4 (N1636, N1635, N1443, N112, N771);
not NOT1 (N1637, N1629);
and AND3 (N1638, N1621, N1162, N1222);
xor XOR2 (N1639, N1632, N1445);
buf BUF1 (N1640, N1627);
xor XOR2 (N1641, N1636, N1302);
not NOT1 (N1642, N1639);
xor XOR2 (N1643, N1637, N943);
nor NOR3 (N1644, N1633, N495, N591);
nor NOR4 (N1645, N1644, N1236, N536, N1144);
or OR2 (N1646, N1643, N113);
xor XOR2 (N1647, N1628, N120);
and AND2 (N1648, N1641, N678);
not NOT1 (N1649, N1634);
not NOT1 (N1650, N1647);
xor XOR2 (N1651, N1640, N402);
and AND4 (N1652, N1646, N1409, N368, N48);
nor NOR2 (N1653, N1624, N1518);
buf BUF1 (N1654, N1653);
not NOT1 (N1655, N1617);
buf BUF1 (N1656, N1638);
nor NOR2 (N1657, N1650, N50);
and AND3 (N1658, N1645, N561, N566);
or OR2 (N1659, N1657, N29);
not NOT1 (N1660, N1649);
not NOT1 (N1661, N1659);
nand NAND2 (N1662, N1661, N1621);
not NOT1 (N1663, N1656);
nor NOR3 (N1664, N1662, N147, N1301);
or OR2 (N1665, N1655, N871);
not NOT1 (N1666, N1651);
buf BUF1 (N1667, N1658);
buf BUF1 (N1668, N1648);
buf BUF1 (N1669, N1660);
buf BUF1 (N1670, N1663);
nor NOR4 (N1671, N1654, N653, N875, N1553);
nor NOR4 (N1672, N1671, N1417, N1598, N344);
xor XOR2 (N1673, N1669, N1546);
and AND4 (N1674, N1652, N1237, N150, N1451);
nand NAND2 (N1675, N1672, N488);
nand NAND4 (N1676, N1667, N702, N843, N1537);
and AND3 (N1677, N1675, N901, N140);
and AND2 (N1678, N1670, N724);
not NOT1 (N1679, N1665);
xor XOR2 (N1680, N1677, N61);
or OR2 (N1681, N1680, N1349);
buf BUF1 (N1682, N1668);
xor XOR2 (N1683, N1673, N1611);
and AND3 (N1684, N1683, N108, N1339);
or OR3 (N1685, N1681, N1110, N864);
nand NAND2 (N1686, N1679, N75);
xor XOR2 (N1687, N1686, N297);
or OR2 (N1688, N1674, N1119);
not NOT1 (N1689, N1682);
buf BUF1 (N1690, N1688);
xor XOR2 (N1691, N1664, N1663);
not NOT1 (N1692, N1691);
and AND2 (N1693, N1684, N1691);
xor XOR2 (N1694, N1685, N615);
nor NOR4 (N1695, N1694, N1133, N577, N1402);
xor XOR2 (N1696, N1666, N1661);
nand NAND3 (N1697, N1696, N822, N532);
xor XOR2 (N1698, N1695, N717);
and AND3 (N1699, N1689, N168, N366);
nor NOR4 (N1700, N1690, N224, N1144, N1499);
buf BUF1 (N1701, N1676);
nor NOR4 (N1702, N1678, N1006, N1593, N730);
not NOT1 (N1703, N1698);
nand NAND3 (N1704, N1692, N924, N519);
nand NAND4 (N1705, N1697, N1064, N402, N811);
nand NAND4 (N1706, N1705, N725, N1207, N1036);
xor XOR2 (N1707, N1642, N1283);
buf BUF1 (N1708, N1693);
xor XOR2 (N1709, N1706, N1636);
buf BUF1 (N1710, N1704);
nor NOR2 (N1711, N1702, N491);
buf BUF1 (N1712, N1708);
nor NOR4 (N1713, N1710, N816, N74, N88);
nand NAND4 (N1714, N1711, N1456, N1671, N1586);
not NOT1 (N1715, N1714);
xor XOR2 (N1716, N1707, N624);
or OR4 (N1717, N1716, N573, N248, N1283);
and AND2 (N1718, N1713, N1660);
nand NAND4 (N1719, N1715, N166, N1137, N1484);
buf BUF1 (N1720, N1719);
nand NAND4 (N1721, N1717, N276, N1720, N1692);
buf BUF1 (N1722, N1715);
xor XOR2 (N1723, N1701, N500);
not NOT1 (N1724, N1687);
not NOT1 (N1725, N1721);
nand NAND3 (N1726, N1709, N463, N1531);
nor NOR4 (N1727, N1722, N240, N728, N1545);
or OR4 (N1728, N1712, N798, N833, N1019);
or OR2 (N1729, N1725, N1712);
not NOT1 (N1730, N1727);
or OR2 (N1731, N1700, N1327);
xor XOR2 (N1732, N1703, N145);
nor NOR4 (N1733, N1728, N968, N185, N383);
or OR4 (N1734, N1724, N777, N1265, N550);
not NOT1 (N1735, N1734);
nor NOR3 (N1736, N1726, N506, N496);
nor NOR4 (N1737, N1735, N230, N794, N1287);
nand NAND4 (N1738, N1733, N880, N175, N1524);
xor XOR2 (N1739, N1732, N591);
not NOT1 (N1740, N1738);
buf BUF1 (N1741, N1699);
xor XOR2 (N1742, N1731, N199);
buf BUF1 (N1743, N1718);
or OR3 (N1744, N1741, N1240, N1582);
not NOT1 (N1745, N1736);
not NOT1 (N1746, N1742);
nor NOR4 (N1747, N1730, N1380, N1295, N572);
xor XOR2 (N1748, N1743, N995);
nor NOR2 (N1749, N1723, N1263);
and AND2 (N1750, N1729, N804);
buf BUF1 (N1751, N1749);
not NOT1 (N1752, N1747);
or OR4 (N1753, N1739, N1136, N289, N1380);
xor XOR2 (N1754, N1744, N254);
xor XOR2 (N1755, N1753, N794);
buf BUF1 (N1756, N1751);
nand NAND3 (N1757, N1752, N754, N1678);
and AND4 (N1758, N1748, N441, N886, N13);
or OR2 (N1759, N1740, N1316);
buf BUF1 (N1760, N1745);
not NOT1 (N1761, N1756);
nor NOR2 (N1762, N1746, N1570);
and AND2 (N1763, N1737, N407);
buf BUF1 (N1764, N1761);
not NOT1 (N1765, N1762);
buf BUF1 (N1766, N1760);
and AND4 (N1767, N1759, N1483, N1500, N422);
nor NOR2 (N1768, N1764, N164);
xor XOR2 (N1769, N1757, N15);
nand NAND2 (N1770, N1750, N341);
or OR3 (N1771, N1767, N1703, N1534);
buf BUF1 (N1772, N1758);
nor NOR2 (N1773, N1763, N651);
buf BUF1 (N1774, N1754);
nand NAND2 (N1775, N1768, N1122);
not NOT1 (N1776, N1765);
and AND2 (N1777, N1775, N1724);
nor NOR4 (N1778, N1777, N1683, N343, N506);
nor NOR3 (N1779, N1770, N1677, N890);
not NOT1 (N1780, N1776);
and AND2 (N1781, N1773, N1252);
not NOT1 (N1782, N1771);
or OR4 (N1783, N1778, N1148, N859, N179);
nand NAND4 (N1784, N1779, N1288, N358, N1570);
nor NOR3 (N1785, N1781, N662, N140);
or OR4 (N1786, N1780, N1666, N638, N832);
buf BUF1 (N1787, N1784);
or OR4 (N1788, N1783, N791, N1217, N637);
and AND4 (N1789, N1782, N980, N1411, N1609);
or OR3 (N1790, N1774, N137, N879);
nand NAND3 (N1791, N1787, N446, N665);
nor NOR2 (N1792, N1788, N390);
buf BUF1 (N1793, N1789);
xor XOR2 (N1794, N1769, N366);
nand NAND2 (N1795, N1786, N727);
nor NOR3 (N1796, N1755, N1108, N1538);
and AND3 (N1797, N1772, N1724, N1170);
and AND4 (N1798, N1797, N1343, N301, N610);
buf BUF1 (N1799, N1766);
or OR3 (N1800, N1796, N1705, N1451);
or OR2 (N1801, N1793, N860);
and AND3 (N1802, N1790, N803, N874);
and AND3 (N1803, N1792, N120, N949);
xor XOR2 (N1804, N1794, N1361);
or OR2 (N1805, N1798, N1588);
not NOT1 (N1806, N1804);
or OR3 (N1807, N1785, N955, N109);
xor XOR2 (N1808, N1802, N1697);
and AND2 (N1809, N1800, N359);
nor NOR3 (N1810, N1799, N1784, N60);
nor NOR2 (N1811, N1801, N1343);
nand NAND2 (N1812, N1809, N1328);
nand NAND2 (N1813, N1803, N854);
nor NOR4 (N1814, N1810, N967, N1389, N1147);
buf BUF1 (N1815, N1806);
or OR3 (N1816, N1805, N18, N770);
or OR3 (N1817, N1813, N1257, N1583);
xor XOR2 (N1818, N1795, N1521);
buf BUF1 (N1819, N1816);
nor NOR2 (N1820, N1791, N1215);
not NOT1 (N1821, N1811);
not NOT1 (N1822, N1812);
buf BUF1 (N1823, N1820);
or OR4 (N1824, N1821, N210, N961, N13);
nand NAND4 (N1825, N1824, N195, N666, N1142);
or OR4 (N1826, N1823, N1222, N244, N325);
nand NAND4 (N1827, N1815, N1583, N151, N230);
not NOT1 (N1828, N1817);
not NOT1 (N1829, N1818);
nand NAND2 (N1830, N1822, N237);
nand NAND3 (N1831, N1825, N173, N1221);
not NOT1 (N1832, N1814);
xor XOR2 (N1833, N1808, N747);
nand NAND2 (N1834, N1826, N746);
buf BUF1 (N1835, N1832);
xor XOR2 (N1836, N1827, N362);
nor NOR3 (N1837, N1831, N843, N848);
not NOT1 (N1838, N1835);
buf BUF1 (N1839, N1836);
or OR3 (N1840, N1834, N1393, N1581);
nand NAND3 (N1841, N1829, N108, N62);
xor XOR2 (N1842, N1819, N611);
buf BUF1 (N1843, N1807);
not NOT1 (N1844, N1838);
or OR2 (N1845, N1841, N773);
buf BUF1 (N1846, N1844);
nor NOR4 (N1847, N1839, N1443, N758, N1821);
nor NOR3 (N1848, N1828, N483, N428);
or OR3 (N1849, N1848, N1584, N803);
buf BUF1 (N1850, N1837);
xor XOR2 (N1851, N1830, N1545);
and AND4 (N1852, N1843, N977, N907, N1775);
nor NOR3 (N1853, N1846, N348, N180);
nand NAND2 (N1854, N1842, N1427);
nand NAND2 (N1855, N1852, N408);
and AND2 (N1856, N1840, N466);
xor XOR2 (N1857, N1845, N450);
nor NOR3 (N1858, N1850, N371, N534);
buf BUF1 (N1859, N1854);
not NOT1 (N1860, N1855);
buf BUF1 (N1861, N1853);
or OR2 (N1862, N1849, N1363);
nor NOR2 (N1863, N1859, N1156);
nand NAND3 (N1864, N1856, N1234, N1173);
xor XOR2 (N1865, N1862, N1347);
not NOT1 (N1866, N1865);
and AND4 (N1867, N1866, N1636, N1732, N84);
nor NOR4 (N1868, N1863, N1830, N664, N1403);
xor XOR2 (N1869, N1867, N1828);
and AND2 (N1870, N1869, N1433);
not NOT1 (N1871, N1857);
buf BUF1 (N1872, N1864);
nand NAND2 (N1873, N1833, N797);
not NOT1 (N1874, N1847);
nand NAND4 (N1875, N1851, N762, N1097, N1761);
xor XOR2 (N1876, N1872, N1612);
or OR2 (N1877, N1874, N1786);
nor NOR4 (N1878, N1860, N1011, N793, N1818);
xor XOR2 (N1879, N1870, N1779);
nor NOR3 (N1880, N1871, N1441, N461);
and AND3 (N1881, N1876, N797, N1344);
nand NAND4 (N1882, N1878, N1071, N632, N699);
nand NAND3 (N1883, N1875, N237, N1698);
nand NAND2 (N1884, N1868, N545);
nand NAND4 (N1885, N1879, N1432, N231, N1458);
xor XOR2 (N1886, N1880, N138);
xor XOR2 (N1887, N1877, N1462);
or OR2 (N1888, N1887, N1532);
nor NOR3 (N1889, N1858, N97, N595);
or OR2 (N1890, N1885, N735);
nor NOR2 (N1891, N1888, N149);
not NOT1 (N1892, N1886);
or OR4 (N1893, N1861, N1781, N1314, N188);
nand NAND2 (N1894, N1892, N797);
buf BUF1 (N1895, N1882);
and AND4 (N1896, N1893, N291, N3, N1165);
xor XOR2 (N1897, N1896, N141);
not NOT1 (N1898, N1897);
not NOT1 (N1899, N1881);
xor XOR2 (N1900, N1884, N193);
nand NAND2 (N1901, N1883, N829);
and AND2 (N1902, N1895, N243);
nor NOR4 (N1903, N1894, N1056, N1382, N136);
not NOT1 (N1904, N1901);
nand NAND4 (N1905, N1891, N576, N750, N974);
not NOT1 (N1906, N1905);
nand NAND4 (N1907, N1900, N25, N381, N738);
or OR3 (N1908, N1898, N52, N1157);
and AND4 (N1909, N1907, N1631, N419, N23);
buf BUF1 (N1910, N1903);
or OR2 (N1911, N1899, N1484);
not NOT1 (N1912, N1911);
not NOT1 (N1913, N1906);
buf BUF1 (N1914, N1904);
and AND2 (N1915, N1909, N1772);
nor NOR3 (N1916, N1915, N259, N787);
nor NOR2 (N1917, N1902, N101);
nor NOR4 (N1918, N1910, N725, N180, N1086);
nor NOR4 (N1919, N1873, N630, N1034, N1200);
and AND3 (N1920, N1913, N1138, N189);
xor XOR2 (N1921, N1912, N838);
or OR2 (N1922, N1890, N1707);
and AND2 (N1923, N1908, N828);
xor XOR2 (N1924, N1916, N1434);
not NOT1 (N1925, N1921);
and AND2 (N1926, N1919, N285);
nor NOR3 (N1927, N1924, N149, N1452);
not NOT1 (N1928, N1926);
nor NOR3 (N1929, N1917, N1084, N1635);
or OR4 (N1930, N1920, N1308, N543, N21);
not NOT1 (N1931, N1927);
nor NOR2 (N1932, N1930, N1656);
nor NOR4 (N1933, N1925, N661, N54, N1036);
xor XOR2 (N1934, N1922, N450);
or OR2 (N1935, N1931, N1107);
xor XOR2 (N1936, N1923, N611);
and AND2 (N1937, N1889, N374);
not NOT1 (N1938, N1937);
not NOT1 (N1939, N1918);
xor XOR2 (N1940, N1938, N796);
nand NAND3 (N1941, N1928, N1048, N1927);
and AND2 (N1942, N1929, N764);
and AND2 (N1943, N1935, N551);
nor NOR3 (N1944, N1914, N1099, N151);
or OR4 (N1945, N1933, N159, N808, N764);
nand NAND2 (N1946, N1940, N1379);
nand NAND3 (N1947, N1941, N1239, N964);
nand NAND2 (N1948, N1945, N1911);
nor NOR2 (N1949, N1939, N1677);
buf BUF1 (N1950, N1932);
nand NAND2 (N1951, N1934, N590);
and AND4 (N1952, N1946, N1693, N1316, N1818);
and AND4 (N1953, N1944, N1792, N1735, N1241);
or OR2 (N1954, N1950, N432);
and AND3 (N1955, N1948, N513, N279);
nor NOR2 (N1956, N1942, N76);
buf BUF1 (N1957, N1955);
nand NAND2 (N1958, N1951, N1802);
or OR2 (N1959, N1956, N1166);
xor XOR2 (N1960, N1954, N901);
buf BUF1 (N1961, N1936);
and AND3 (N1962, N1961, N594, N930);
and AND3 (N1963, N1953, N1453, N1245);
nor NOR4 (N1964, N1947, N113, N1244, N1485);
nand NAND4 (N1965, N1964, N379, N1845, N1021);
buf BUF1 (N1966, N1957);
nand NAND3 (N1967, N1952, N250, N1702);
or OR2 (N1968, N1965, N171);
and AND3 (N1969, N1966, N1661, N1855);
not NOT1 (N1970, N1949);
xor XOR2 (N1971, N1958, N1893);
and AND4 (N1972, N1969, N1052, N1288, N586);
or OR2 (N1973, N1970, N1050);
nor NOR3 (N1974, N1943, N1051, N1655);
and AND2 (N1975, N1959, N1033);
and AND2 (N1976, N1972, N795);
xor XOR2 (N1977, N1960, N1246);
or OR4 (N1978, N1971, N515, N1231, N196);
not NOT1 (N1979, N1978);
or OR2 (N1980, N1975, N997);
not NOT1 (N1981, N1967);
not NOT1 (N1982, N1963);
buf BUF1 (N1983, N1980);
and AND2 (N1984, N1976, N747);
not NOT1 (N1985, N1984);
xor XOR2 (N1986, N1981, N687);
and AND4 (N1987, N1977, N43, N1313, N1398);
nand NAND3 (N1988, N1962, N913, N43);
not NOT1 (N1989, N1986);
not NOT1 (N1990, N1973);
and AND3 (N1991, N1989, N619, N945);
not NOT1 (N1992, N1985);
nor NOR4 (N1993, N1968, N485, N1116, N1240);
nor NOR2 (N1994, N1988, N1748);
and AND4 (N1995, N1990, N1090, N1467, N1507);
xor XOR2 (N1996, N1983, N1741);
not NOT1 (N1997, N1987);
nand NAND3 (N1998, N1993, N1716, N484);
xor XOR2 (N1999, N1998, N211);
xor XOR2 (N2000, N1982, N1676);
buf BUF1 (N2001, N1974);
not NOT1 (N2002, N1979);
buf BUF1 (N2003, N1992);
and AND3 (N2004, N1997, N1181, N622);
or OR2 (N2005, N1996, N1752);
xor XOR2 (N2006, N1991, N939);
nor NOR3 (N2007, N2003, N103, N1072);
not NOT1 (N2008, N1999);
nor NOR3 (N2009, N1994, N1532, N1881);
not NOT1 (N2010, N2009);
and AND2 (N2011, N2010, N1047);
nor NOR3 (N2012, N2005, N1578, N806);
and AND3 (N2013, N2012, N1973, N1256);
and AND4 (N2014, N2001, N31, N1348, N1502);
or OR4 (N2015, N2011, N9, N1002, N47);
or OR3 (N2016, N2015, N1644, N234);
or OR4 (N2017, N2004, N1974, N1347, N163);
buf BUF1 (N2018, N2013);
nor NOR2 (N2019, N2018, N135);
and AND3 (N2020, N2008, N1484, N199);
and AND2 (N2021, N2000, N329);
not NOT1 (N2022, N2021);
buf BUF1 (N2023, N2022);
and AND4 (N2024, N1995, N680, N1297, N1285);
nand NAND2 (N2025, N2024, N104);
not NOT1 (N2026, N2016);
nor NOR2 (N2027, N2023, N44);
or OR2 (N2028, N2020, N462);
not NOT1 (N2029, N2028);
not NOT1 (N2030, N2017);
nor NOR2 (N2031, N2029, N406);
and AND2 (N2032, N2014, N806);
xor XOR2 (N2033, N2032, N1860);
xor XOR2 (N2034, N2031, N421);
buf BUF1 (N2035, N2033);
xor XOR2 (N2036, N2002, N1668);
nor NOR2 (N2037, N2007, N650);
not NOT1 (N2038, N2037);
not NOT1 (N2039, N2019);
xor XOR2 (N2040, N2025, N1691);
nand NAND4 (N2041, N2026, N562, N1666, N1588);
or OR2 (N2042, N2006, N1266);
xor XOR2 (N2043, N2027, N700);
buf BUF1 (N2044, N2042);
nand NAND3 (N2045, N2030, N284, N249);
and AND2 (N2046, N2041, N648);
or OR3 (N2047, N2044, N362, N1778);
or OR4 (N2048, N2038, N1688, N1101, N1536);
nor NOR3 (N2049, N2048, N882, N73);
nand NAND3 (N2050, N2045, N1973, N1333);
and AND4 (N2051, N2046, N733, N260, N665);
nand NAND4 (N2052, N2035, N215, N1442, N1883);
not NOT1 (N2053, N2040);
not NOT1 (N2054, N2050);
buf BUF1 (N2055, N2047);
buf BUF1 (N2056, N2036);
buf BUF1 (N2057, N2053);
or OR3 (N2058, N2034, N936, N1303);
nand NAND2 (N2059, N2049, N1135);
buf BUF1 (N2060, N2056);
nand NAND4 (N2061, N2043, N385, N492, N1576);
nand NAND2 (N2062, N2061, N1556);
nor NOR4 (N2063, N2060, N1389, N467, N115);
xor XOR2 (N2064, N2051, N772);
and AND3 (N2065, N2054, N1707, N1916);
not NOT1 (N2066, N2059);
or OR2 (N2067, N2063, N1857);
or OR2 (N2068, N2052, N534);
nand NAND3 (N2069, N2055, N1083, N1848);
buf BUF1 (N2070, N2039);
nor NOR3 (N2071, N2069, N263, N720);
or OR2 (N2072, N2058, N1949);
xor XOR2 (N2073, N2067, N468);
nor NOR3 (N2074, N2072, N420, N807);
buf BUF1 (N2075, N2074);
and AND2 (N2076, N2073, N1686);
and AND4 (N2077, N2076, N273, N1130, N1795);
not NOT1 (N2078, N2062);
not NOT1 (N2079, N2065);
or OR3 (N2080, N2078, N801, N1204);
nand NAND2 (N2081, N2064, N1286);
xor XOR2 (N2082, N2081, N1136);
buf BUF1 (N2083, N2080);
buf BUF1 (N2084, N2068);
xor XOR2 (N2085, N2070, N1168);
and AND4 (N2086, N2075, N1924, N860, N993);
not NOT1 (N2087, N2083);
xor XOR2 (N2088, N2077, N545);
or OR3 (N2089, N2057, N5, N1958);
not NOT1 (N2090, N2066);
xor XOR2 (N2091, N2090, N431);
or OR2 (N2092, N2082, N1318);
and AND2 (N2093, N2092, N1290);
or OR3 (N2094, N2088, N952, N1587);
xor XOR2 (N2095, N2071, N1491);
xor XOR2 (N2096, N2093, N1226);
nor NOR4 (N2097, N2095, N1852, N146, N502);
nor NOR3 (N2098, N2084, N443, N2072);
or OR2 (N2099, N2091, N886);
buf BUF1 (N2100, N2099);
not NOT1 (N2101, N2079);
not NOT1 (N2102, N2085);
and AND2 (N2103, N2094, N424);
buf BUF1 (N2104, N2101);
and AND4 (N2105, N2100, N1567, N1414, N511);
xor XOR2 (N2106, N2105, N2083);
buf BUF1 (N2107, N2089);
nand NAND2 (N2108, N2097, N1136);
xor XOR2 (N2109, N2103, N436);
and AND4 (N2110, N2087, N1240, N2099, N556);
or OR3 (N2111, N2107, N1347, N1607);
nor NOR4 (N2112, N2096, N1950, N1880, N772);
nor NOR3 (N2113, N2098, N940, N980);
not NOT1 (N2114, N2086);
nand NAND3 (N2115, N2112, N453, N722);
nand NAND2 (N2116, N2113, N683);
not NOT1 (N2117, N2108);
xor XOR2 (N2118, N2110, N538);
not NOT1 (N2119, N2118);
nand NAND4 (N2120, N2106, N580, N142, N1260);
nor NOR4 (N2121, N2104, N674, N582, N447);
xor XOR2 (N2122, N2121, N1641);
nand NAND3 (N2123, N2102, N1494, N2073);
nand NAND3 (N2124, N2116, N185, N1815);
nor NOR2 (N2125, N2123, N608);
not NOT1 (N2126, N2119);
and AND3 (N2127, N2111, N271, N1320);
buf BUF1 (N2128, N2109);
buf BUF1 (N2129, N2120);
nor NOR4 (N2130, N2117, N709, N1755, N2073);
or OR2 (N2131, N2125, N2098);
not NOT1 (N2132, N2124);
not NOT1 (N2133, N2122);
and AND2 (N2134, N2130, N297);
nor NOR2 (N2135, N2127, N175);
xor XOR2 (N2136, N2115, N781);
not NOT1 (N2137, N2129);
or OR2 (N2138, N2134, N1315);
xor XOR2 (N2139, N2128, N1102);
buf BUF1 (N2140, N2138);
and AND4 (N2141, N2137, N1318, N1211, N1227);
buf BUF1 (N2142, N2141);
xor XOR2 (N2143, N2142, N581);
xor XOR2 (N2144, N2143, N1384);
nand NAND4 (N2145, N2133, N744, N1234, N527);
or OR3 (N2146, N2140, N1343, N977);
nand NAND3 (N2147, N2146, N1249, N420);
or OR2 (N2148, N2126, N803);
nor NOR2 (N2149, N2139, N1928);
buf BUF1 (N2150, N2114);
or OR3 (N2151, N2148, N872, N2129);
nor NOR2 (N2152, N2147, N489);
or OR4 (N2153, N2150, N1930, N1744, N741);
or OR4 (N2154, N2135, N852, N1788, N2129);
nand NAND2 (N2155, N2149, N768);
and AND3 (N2156, N2155, N1359, N136);
xor XOR2 (N2157, N2156, N5);
nor NOR3 (N2158, N2132, N1034, N1690);
buf BUF1 (N2159, N2152);
and AND3 (N2160, N2157, N108, N1871);
nor NOR4 (N2161, N2131, N49, N1809, N2144);
or OR3 (N2162, N1258, N1884, N1511);
and AND3 (N2163, N2158, N109, N1478);
nor NOR4 (N2164, N2163, N1642, N288, N2117);
not NOT1 (N2165, N2159);
buf BUF1 (N2166, N2160);
xor XOR2 (N2167, N2161, N2086);
and AND2 (N2168, N2151, N332);
or OR2 (N2169, N2167, N1907);
or OR4 (N2170, N2165, N1281, N778, N948);
buf BUF1 (N2171, N2162);
nand NAND2 (N2172, N2145, N133);
nand NAND3 (N2173, N2169, N464, N1874);
buf BUF1 (N2174, N2171);
or OR2 (N2175, N2164, N2033);
and AND3 (N2176, N2136, N1951, N1891);
or OR2 (N2177, N2166, N1509);
and AND3 (N2178, N2176, N163, N1847);
or OR4 (N2179, N2172, N703, N2038, N231);
not NOT1 (N2180, N2170);
buf BUF1 (N2181, N2154);
and AND2 (N2182, N2178, N668);
xor XOR2 (N2183, N2153, N1937);
nand NAND4 (N2184, N2175, N1394, N1340, N971);
xor XOR2 (N2185, N2168, N715);
nor NOR2 (N2186, N2174, N1088);
buf BUF1 (N2187, N2181);
or OR2 (N2188, N2187, N1389);
and AND3 (N2189, N2179, N1971, N1787);
buf BUF1 (N2190, N2185);
and AND3 (N2191, N2177, N28, N802);
nor NOR3 (N2192, N2182, N1327, N1155);
or OR2 (N2193, N2186, N87);
nand NAND4 (N2194, N2184, N2099, N309, N848);
xor XOR2 (N2195, N2190, N1234);
xor XOR2 (N2196, N2173, N2042);
and AND4 (N2197, N2191, N334, N1392, N1305);
nor NOR2 (N2198, N2196, N2132);
not NOT1 (N2199, N2194);
and AND3 (N2200, N2189, N704, N548);
xor XOR2 (N2201, N2180, N1323);
and AND4 (N2202, N2199, N771, N2172, N1980);
buf BUF1 (N2203, N2183);
buf BUF1 (N2204, N2201);
xor XOR2 (N2205, N2192, N513);
and AND4 (N2206, N2198, N234, N1393, N2155);
nor NOR2 (N2207, N2202, N667);
xor XOR2 (N2208, N2204, N648);
or OR3 (N2209, N2203, N1779, N1283);
buf BUF1 (N2210, N2207);
nand NAND2 (N2211, N2206, N648);
not NOT1 (N2212, N2195);
buf BUF1 (N2213, N2208);
or OR3 (N2214, N2197, N325, N397);
or OR4 (N2215, N2188, N593, N397, N168);
buf BUF1 (N2216, N2215);
buf BUF1 (N2217, N2200);
nor NOR3 (N2218, N2216, N692, N927);
nand NAND4 (N2219, N2211, N658, N97, N1364);
nor NOR4 (N2220, N2219, N2029, N1192, N75);
nor NOR3 (N2221, N2193, N1707, N1823);
or OR4 (N2222, N2214, N388, N1025, N174);
and AND3 (N2223, N2220, N182, N761);
xor XOR2 (N2224, N2212, N966);
not NOT1 (N2225, N2217);
or OR4 (N2226, N2213, N2055, N842, N505);
nor NOR2 (N2227, N2225, N89);
and AND4 (N2228, N2221, N1630, N2058, N906);
nand NAND3 (N2229, N2227, N50, N79);
xor XOR2 (N2230, N2222, N1434);
or OR4 (N2231, N2226, N506, N2042, N1449);
nor NOR3 (N2232, N2205, N619, N1762);
or OR2 (N2233, N2229, N1879);
buf BUF1 (N2234, N2210);
nor NOR3 (N2235, N2224, N1402, N507);
not NOT1 (N2236, N2218);
nor NOR4 (N2237, N2232, N901, N1177, N347);
or OR3 (N2238, N2231, N392, N482);
nor NOR3 (N2239, N2238, N2191, N1598);
or OR3 (N2240, N2236, N1671, N925);
or OR3 (N2241, N2230, N575, N1063);
nand NAND2 (N2242, N2233, N705);
buf BUF1 (N2243, N2235);
xor XOR2 (N2244, N2228, N926);
and AND2 (N2245, N2242, N357);
nand NAND2 (N2246, N2240, N1850);
buf BUF1 (N2247, N2246);
buf BUF1 (N2248, N2234);
nand NAND3 (N2249, N2247, N1195, N2147);
not NOT1 (N2250, N2209);
nand NAND2 (N2251, N2249, N1856);
buf BUF1 (N2252, N2243);
buf BUF1 (N2253, N2252);
xor XOR2 (N2254, N2244, N527);
nand NAND2 (N2255, N2245, N1642);
buf BUF1 (N2256, N2241);
or OR2 (N2257, N2223, N660);
not NOT1 (N2258, N2251);
xor XOR2 (N2259, N2248, N322);
not NOT1 (N2260, N2258);
not NOT1 (N2261, N2255);
buf BUF1 (N2262, N2257);
not NOT1 (N2263, N2259);
buf BUF1 (N2264, N2250);
not NOT1 (N2265, N2256);
xor XOR2 (N2266, N2262, N930);
or OR3 (N2267, N2239, N1080, N1549);
xor XOR2 (N2268, N2265, N882);
nor NOR4 (N2269, N2264, N1199, N1646, N703);
nor NOR4 (N2270, N2269, N1113, N1191, N1985);
nand NAND4 (N2271, N2261, N177, N786, N1177);
buf BUF1 (N2272, N2270);
not NOT1 (N2273, N2272);
not NOT1 (N2274, N2260);
buf BUF1 (N2275, N2273);
and AND3 (N2276, N2267, N2251, N504);
xor XOR2 (N2277, N2275, N368);
nand NAND2 (N2278, N2276, N257);
buf BUF1 (N2279, N2237);
nand NAND3 (N2280, N2266, N1732, N407);
and AND3 (N2281, N2278, N389, N1902);
buf BUF1 (N2282, N2268);
nand NAND4 (N2283, N2271, N987, N1304, N1166);
and AND4 (N2284, N2254, N1357, N1397, N1535);
buf BUF1 (N2285, N2284);
nor NOR3 (N2286, N2283, N101, N1838);
buf BUF1 (N2287, N2285);
or OR2 (N2288, N2279, N765);
nor NOR2 (N2289, N2286, N1549);
buf BUF1 (N2290, N2289);
xor XOR2 (N2291, N2288, N16);
or OR2 (N2292, N2277, N874);
buf BUF1 (N2293, N2281);
xor XOR2 (N2294, N2253, N1620);
buf BUF1 (N2295, N2293);
not NOT1 (N2296, N2280);
xor XOR2 (N2297, N2263, N733);
nand NAND4 (N2298, N2292, N507, N277, N1195);
buf BUF1 (N2299, N2287);
nand NAND2 (N2300, N2294, N361);
not NOT1 (N2301, N2282);
buf BUF1 (N2302, N2300);
and AND3 (N2303, N2301, N606, N332);
or OR2 (N2304, N2274, N44);
not NOT1 (N2305, N2297);
and AND3 (N2306, N2304, N27, N1573);
nand NAND4 (N2307, N2291, N238, N834, N835);
and AND4 (N2308, N2299, N17, N1012, N1203);
or OR4 (N2309, N2302, N1075, N131, N2154);
nand NAND2 (N2310, N2303, N1632);
or OR2 (N2311, N2305, N1735);
or OR2 (N2312, N2306, N759);
and AND4 (N2313, N2309, N1124, N1395, N546);
xor XOR2 (N2314, N2290, N1551);
or OR2 (N2315, N2308, N662);
or OR4 (N2316, N2307, N373, N1111, N1343);
nand NAND2 (N2317, N2315, N447);
or OR4 (N2318, N2311, N2222, N1249, N498);
or OR2 (N2319, N2317, N1462);
and AND4 (N2320, N2295, N1669, N1577, N1132);
nand NAND2 (N2321, N2313, N798);
not NOT1 (N2322, N2319);
and AND2 (N2323, N2321, N99);
buf BUF1 (N2324, N2298);
or OR2 (N2325, N2314, N174);
and AND2 (N2326, N2325, N431);
not NOT1 (N2327, N2324);
not NOT1 (N2328, N2310);
nor NOR2 (N2329, N2320, N2106);
and AND4 (N2330, N2312, N1326, N1383, N231);
xor XOR2 (N2331, N2328, N549);
buf BUF1 (N2332, N2322);
and AND3 (N2333, N2318, N156, N725);
buf BUF1 (N2334, N2296);
and AND2 (N2335, N2323, N1412);
and AND4 (N2336, N2330, N1725, N1695, N313);
xor XOR2 (N2337, N2334, N1054);
and AND4 (N2338, N2331, N698, N1070, N939);
not NOT1 (N2339, N2329);
or OR4 (N2340, N2332, N2123, N1541, N763);
not NOT1 (N2341, N2333);
nor NOR3 (N2342, N2341, N2140, N1697);
xor XOR2 (N2343, N2327, N1107);
not NOT1 (N2344, N2340);
or OR4 (N2345, N2338, N300, N1367, N593);
nand NAND3 (N2346, N2326, N1551, N303);
buf BUF1 (N2347, N2343);
nand NAND3 (N2348, N2344, N2341, N984);
xor XOR2 (N2349, N2337, N2301);
nand NAND3 (N2350, N2339, N1068, N1508);
nand NAND3 (N2351, N2346, N334, N1233);
nor NOR3 (N2352, N2347, N1226, N188);
xor XOR2 (N2353, N2348, N1401);
and AND4 (N2354, N2316, N1303, N1743, N592);
buf BUF1 (N2355, N2352);
nand NAND2 (N2356, N2336, N2007);
buf BUF1 (N2357, N2355);
not NOT1 (N2358, N2335);
or OR2 (N2359, N2349, N1149);
nand NAND3 (N2360, N2354, N2164, N1989);
xor XOR2 (N2361, N2345, N94);
or OR3 (N2362, N2350, N1712, N1183);
or OR4 (N2363, N2360, N1080, N1802, N506);
nor NOR4 (N2364, N2362, N2119, N1254, N182);
xor XOR2 (N2365, N2356, N511);
and AND3 (N2366, N2363, N573, N1838);
xor XOR2 (N2367, N2364, N1409);
nor NOR3 (N2368, N2366, N1231, N56);
buf BUF1 (N2369, N2357);
xor XOR2 (N2370, N2359, N1984);
buf BUF1 (N2371, N2351);
and AND2 (N2372, N2353, N612);
and AND2 (N2373, N2365, N2003);
buf BUF1 (N2374, N2372);
not NOT1 (N2375, N2367);
buf BUF1 (N2376, N2361);
and AND3 (N2377, N2342, N1609, N1655);
xor XOR2 (N2378, N2371, N1888);
not NOT1 (N2379, N2358);
nand NAND3 (N2380, N2370, N844, N1393);
not NOT1 (N2381, N2374);
not NOT1 (N2382, N2375);
buf BUF1 (N2383, N2380);
xor XOR2 (N2384, N2369, N1281);
nor NOR4 (N2385, N2377, N540, N983, N650);
or OR3 (N2386, N2381, N2062, N1407);
nor NOR4 (N2387, N2386, N456, N212, N451);
and AND2 (N2388, N2368, N1371);
and AND2 (N2389, N2373, N304);
nor NOR3 (N2390, N2383, N1635, N1605);
or OR4 (N2391, N2385, N1140, N304, N1919);
nor NOR4 (N2392, N2388, N1571, N1797, N1281);
nor NOR2 (N2393, N2378, N1656);
xor XOR2 (N2394, N2384, N613);
buf BUF1 (N2395, N2376);
or OR4 (N2396, N2382, N642, N1391, N1288);
not NOT1 (N2397, N2390);
not NOT1 (N2398, N2395);
nand NAND4 (N2399, N2391, N1395, N277, N2260);
nand NAND3 (N2400, N2397, N316, N793);
nor NOR3 (N2401, N2394, N379, N2362);
nand NAND4 (N2402, N2401, N1416, N1911, N1732);
buf BUF1 (N2403, N2392);
buf BUF1 (N2404, N2402);
not NOT1 (N2405, N2400);
not NOT1 (N2406, N2405);
nand NAND3 (N2407, N2396, N1609, N1848);
and AND2 (N2408, N2398, N1750);
not NOT1 (N2409, N2404);
nand NAND4 (N2410, N2408, N1007, N1385, N881);
not NOT1 (N2411, N2410);
nand NAND2 (N2412, N2403, N1932);
and AND3 (N2413, N2379, N258, N98);
nand NAND4 (N2414, N2399, N456, N1641, N666);
or OR4 (N2415, N2409, N67, N1303, N47);
or OR4 (N2416, N2415, N807, N2377, N340);
and AND3 (N2417, N2406, N2178, N428);
not NOT1 (N2418, N2393);
buf BUF1 (N2419, N2389);
or OR3 (N2420, N2387, N2016, N1091);
not NOT1 (N2421, N2407);
nand NAND4 (N2422, N2419, N1924, N387, N2280);
or OR3 (N2423, N2413, N240, N1190);
not NOT1 (N2424, N2418);
buf BUF1 (N2425, N2411);
not NOT1 (N2426, N2423);
buf BUF1 (N2427, N2417);
xor XOR2 (N2428, N2421, N418);
xor XOR2 (N2429, N2428, N1827);
buf BUF1 (N2430, N2424);
or OR2 (N2431, N2420, N1601);
or OR3 (N2432, N2430, N772, N2362);
nor NOR3 (N2433, N2416, N1053, N835);
buf BUF1 (N2434, N2433);
nand NAND3 (N2435, N2427, N2027, N691);
or OR2 (N2436, N2435, N1737);
nand NAND2 (N2437, N2434, N1433);
or OR2 (N2438, N2412, N2388);
xor XOR2 (N2439, N2425, N609);
or OR3 (N2440, N2437, N318, N489);
or OR3 (N2441, N2439, N864, N334);
nor NOR3 (N2442, N2438, N161, N1998);
xor XOR2 (N2443, N2414, N889);
or OR2 (N2444, N2429, N1047);
and AND2 (N2445, N2443, N1237);
buf BUF1 (N2446, N2440);
or OR3 (N2447, N2446, N1572, N1473);
not NOT1 (N2448, N2441);
xor XOR2 (N2449, N2432, N192);
and AND4 (N2450, N2449, N641, N2334, N1752);
or OR4 (N2451, N2445, N1571, N1321, N1250);
nand NAND2 (N2452, N2442, N146);
or OR2 (N2453, N2422, N153);
or OR2 (N2454, N2448, N510);
nand NAND4 (N2455, N2426, N30, N365, N728);
buf BUF1 (N2456, N2453);
or OR4 (N2457, N2451, N1522, N527, N2132);
and AND3 (N2458, N2450, N963, N1540);
xor XOR2 (N2459, N2431, N880);
or OR2 (N2460, N2452, N1983);
or OR2 (N2461, N2444, N2255);
buf BUF1 (N2462, N2461);
or OR4 (N2463, N2454, N1643, N2413, N2359);
nor NOR4 (N2464, N2458, N753, N168, N1861);
nand NAND3 (N2465, N2457, N1588, N91);
nor NOR2 (N2466, N2459, N2408);
buf BUF1 (N2467, N2456);
xor XOR2 (N2468, N2464, N1091);
nand NAND4 (N2469, N2447, N2050, N823, N744);
nor NOR3 (N2470, N2463, N641, N618);
nand NAND2 (N2471, N2455, N790);
nand NAND3 (N2472, N2471, N493, N1987);
and AND2 (N2473, N2460, N2449);
or OR2 (N2474, N2472, N1250);
buf BUF1 (N2475, N2462);
or OR3 (N2476, N2468, N418, N1629);
nor NOR2 (N2477, N2467, N1986);
nand NAND3 (N2478, N2469, N995, N375);
or OR3 (N2479, N2475, N697, N1657);
and AND3 (N2480, N2478, N540, N1029);
and AND3 (N2481, N2470, N2296, N1208);
nor NOR3 (N2482, N2481, N81, N1092);
nor NOR3 (N2483, N2474, N2161, N1738);
nor NOR2 (N2484, N2473, N266);
or OR2 (N2485, N2482, N1817);
nor NOR4 (N2486, N2484, N1427, N1763, N984);
xor XOR2 (N2487, N2476, N1199);
and AND3 (N2488, N2480, N781, N192);
xor XOR2 (N2489, N2487, N959);
nor NOR4 (N2490, N2436, N2249, N815, N110);
and AND4 (N2491, N2488, N2363, N1972, N618);
not NOT1 (N2492, N2486);
not NOT1 (N2493, N2485);
nand NAND4 (N2494, N2492, N735, N700, N6);
or OR4 (N2495, N2494, N2262, N1627, N1332);
and AND3 (N2496, N2465, N565, N1258);
xor XOR2 (N2497, N2483, N2436);
or OR2 (N2498, N2497, N848);
nand NAND4 (N2499, N2466, N1776, N377, N1663);
xor XOR2 (N2500, N2495, N963);
or OR3 (N2501, N2477, N81, N1255);
or OR3 (N2502, N2501, N2158, N2190);
buf BUF1 (N2503, N2502);
or OR3 (N2504, N2498, N1918, N978);
or OR3 (N2505, N2504, N1789, N345);
not NOT1 (N2506, N2491);
buf BUF1 (N2507, N2506);
buf BUF1 (N2508, N2496);
and AND3 (N2509, N2490, N2177, N415);
nand NAND4 (N2510, N2489, N2156, N858, N1861);
and AND3 (N2511, N2499, N232, N965);
nand NAND3 (N2512, N2505, N1733, N813);
not NOT1 (N2513, N2503);
xor XOR2 (N2514, N2508, N1110);
and AND2 (N2515, N2513, N1241);
buf BUF1 (N2516, N2507);
xor XOR2 (N2517, N2479, N740);
xor XOR2 (N2518, N2517, N1949);
or OR2 (N2519, N2514, N884);
nor NOR3 (N2520, N2519, N369, N1011);
or OR4 (N2521, N2515, N466, N293, N483);
nand NAND4 (N2522, N2521, N921, N2120, N1371);
or OR3 (N2523, N2522, N2129, N908);
and AND2 (N2524, N2523, N919);
and AND4 (N2525, N2524, N2227, N2010, N1391);
buf BUF1 (N2526, N2525);
not NOT1 (N2527, N2500);
xor XOR2 (N2528, N2520, N913);
nor NOR4 (N2529, N2528, N2254, N1533, N158);
buf BUF1 (N2530, N2511);
nand NAND4 (N2531, N2518, N1003, N1604, N1512);
or OR2 (N2532, N2512, N1346);
nand NAND2 (N2533, N2530, N530);
nand NAND2 (N2534, N2533, N1948);
and AND3 (N2535, N2493, N1329, N2285);
nor NOR2 (N2536, N2535, N2461);
nor NOR2 (N2537, N2510, N277);
and AND2 (N2538, N2537, N1573);
or OR2 (N2539, N2516, N2170);
not NOT1 (N2540, N2529);
and AND2 (N2541, N2539, N2206);
xor XOR2 (N2542, N2540, N2354);
xor XOR2 (N2543, N2542, N2454);
or OR2 (N2544, N2509, N1537);
buf BUF1 (N2545, N2544);
buf BUF1 (N2546, N2543);
nand NAND4 (N2547, N2532, N1016, N1509, N640);
not NOT1 (N2548, N2546);
and AND3 (N2549, N2526, N848, N1283);
buf BUF1 (N2550, N2538);
nor NOR4 (N2551, N2536, N154, N564, N2454);
nand NAND2 (N2552, N2541, N179);
xor XOR2 (N2553, N2552, N740);
buf BUF1 (N2554, N2550);
and AND4 (N2555, N2553, N1215, N336, N555);
or OR3 (N2556, N2554, N1869, N1485);
xor XOR2 (N2557, N2555, N1899);
nor NOR3 (N2558, N2557, N1250, N2325);
nand NAND3 (N2559, N2548, N2006, N1622);
buf BUF1 (N2560, N2527);
xor XOR2 (N2561, N2558, N1746);
xor XOR2 (N2562, N2556, N2390);
nand NAND2 (N2563, N2545, N2274);
xor XOR2 (N2564, N2547, N618);
not NOT1 (N2565, N2531);
nand NAND4 (N2566, N2560, N916, N1616, N1470);
xor XOR2 (N2567, N2534, N54);
xor XOR2 (N2568, N2567, N2156);
not NOT1 (N2569, N2562);
xor XOR2 (N2570, N2568, N593);
buf BUF1 (N2571, N2559);
not NOT1 (N2572, N2549);
not NOT1 (N2573, N2570);
buf BUF1 (N2574, N2569);
nor NOR2 (N2575, N2572, N2441);
buf BUF1 (N2576, N2551);
buf BUF1 (N2577, N2574);
and AND4 (N2578, N2566, N242, N49, N1283);
buf BUF1 (N2579, N2571);
xor XOR2 (N2580, N2563, N928);
and AND4 (N2581, N2561, N1696, N1098, N2239);
xor XOR2 (N2582, N2576, N1843);
not NOT1 (N2583, N2564);
xor XOR2 (N2584, N2579, N2169);
nor NOR4 (N2585, N2573, N513, N698, N711);
or OR2 (N2586, N2582, N900);
buf BUF1 (N2587, N2586);
xor XOR2 (N2588, N2583, N1088);
buf BUF1 (N2589, N2575);
buf BUF1 (N2590, N2587);
nor NOR4 (N2591, N2585, N788, N1076, N729);
xor XOR2 (N2592, N2578, N1988);
or OR3 (N2593, N2581, N1555, N782);
nand NAND3 (N2594, N2580, N860, N1035);
nand NAND3 (N2595, N2591, N458, N615);
and AND2 (N2596, N2589, N2277);
nor NOR3 (N2597, N2594, N367, N371);
nand NAND2 (N2598, N2592, N1316);
not NOT1 (N2599, N2590);
not NOT1 (N2600, N2598);
nor NOR2 (N2601, N2577, N231);
nor NOR3 (N2602, N2584, N1486, N234);
and AND4 (N2603, N2599, N760, N27, N1540);
nor NOR4 (N2604, N2602, N2392, N57, N886);
or OR2 (N2605, N2600, N159);
and AND2 (N2606, N2597, N1417);
not NOT1 (N2607, N2606);
nor NOR2 (N2608, N2607, N31);
not NOT1 (N2609, N2603);
not NOT1 (N2610, N2608);
not NOT1 (N2611, N2588);
buf BUF1 (N2612, N2611);
nor NOR4 (N2613, N2610, N1296, N663, N1020);
and AND2 (N2614, N2595, N277);
nand NAND3 (N2615, N2612, N2346, N320);
nand NAND3 (N2616, N2613, N2577, N1079);
buf BUF1 (N2617, N2601);
nor NOR2 (N2618, N2565, N338);
not NOT1 (N2619, N2605);
buf BUF1 (N2620, N2596);
nor NOR4 (N2621, N2615, N780, N1709, N2002);
xor XOR2 (N2622, N2604, N2063);
buf BUF1 (N2623, N2621);
nor NOR4 (N2624, N2622, N738, N136, N1328);
not NOT1 (N2625, N2619);
not NOT1 (N2626, N2620);
nor NOR2 (N2627, N2616, N1127);
xor XOR2 (N2628, N2626, N1067);
nor NOR3 (N2629, N2628, N344, N1057);
not NOT1 (N2630, N2627);
nor NOR4 (N2631, N2614, N275, N277, N2153);
nor NOR2 (N2632, N2625, N934);
nor NOR4 (N2633, N2618, N235, N1320, N1722);
nand NAND2 (N2634, N2632, N232);
nor NOR4 (N2635, N2633, N2264, N1585, N2508);
and AND4 (N2636, N2624, N57, N130, N421);
or OR4 (N2637, N2630, N96, N607, N1037);
buf BUF1 (N2638, N2609);
or OR4 (N2639, N2593, N840, N1442, N1973);
and AND2 (N2640, N2638, N1162);
not NOT1 (N2641, N2635);
buf BUF1 (N2642, N2617);
xor XOR2 (N2643, N2640, N2009);
or OR4 (N2644, N2637, N1514, N656, N1562);
not NOT1 (N2645, N2634);
or OR4 (N2646, N2644, N1568, N916, N967);
or OR2 (N2647, N2623, N2438);
nand NAND2 (N2648, N2629, N566);
nand NAND2 (N2649, N2647, N993);
nand NAND4 (N2650, N2645, N2556, N850, N128);
xor XOR2 (N2651, N2649, N2301);
and AND2 (N2652, N2641, N1181);
buf BUF1 (N2653, N2639);
and AND3 (N2654, N2643, N2632, N981);
not NOT1 (N2655, N2642);
nor NOR4 (N2656, N2650, N461, N1582, N1730);
not NOT1 (N2657, N2656);
nand NAND3 (N2658, N2646, N2272, N2188);
buf BUF1 (N2659, N2657);
nand NAND2 (N2660, N2653, N737);
and AND2 (N2661, N2648, N186);
and AND2 (N2662, N2659, N480);
and AND4 (N2663, N2655, N2150, N2409, N983);
buf BUF1 (N2664, N2631);
and AND4 (N2665, N2636, N1470, N921, N248);
not NOT1 (N2666, N2665);
nor NOR2 (N2667, N2652, N447);
buf BUF1 (N2668, N2660);
not NOT1 (N2669, N2664);
nand NAND2 (N2670, N2669, N1073);
or OR3 (N2671, N2663, N1279, N2553);
nor NOR3 (N2672, N2668, N536, N1344);
or OR4 (N2673, N2658, N1067, N2559, N2601);
nand NAND2 (N2674, N2671, N2388);
nand NAND3 (N2675, N2651, N2334, N1002);
not NOT1 (N2676, N2654);
nand NAND4 (N2677, N2666, N352, N2578, N1688);
and AND4 (N2678, N2675, N931, N32, N543);
or OR4 (N2679, N2667, N1124, N2531, N2339);
or OR2 (N2680, N2678, N2026);
or OR2 (N2681, N2680, N751);
or OR4 (N2682, N2681, N1737, N446, N985);
not NOT1 (N2683, N2676);
nand NAND4 (N2684, N2670, N2355, N1018, N2570);
buf BUF1 (N2685, N2683);
and AND4 (N2686, N2685, N516, N2512, N2034);
nand NAND2 (N2687, N2686, N1621);
and AND2 (N2688, N2687, N778);
and AND3 (N2689, N2661, N1682, N395);
nor NOR3 (N2690, N2684, N375, N741);
xor XOR2 (N2691, N2688, N2074);
buf BUF1 (N2692, N2672);
buf BUF1 (N2693, N2691);
and AND2 (N2694, N2674, N2584);
not NOT1 (N2695, N2692);
xor XOR2 (N2696, N2694, N1019);
nand NAND4 (N2697, N2682, N598, N2192, N564);
xor XOR2 (N2698, N2677, N1878);
not NOT1 (N2699, N2690);
not NOT1 (N2700, N2673);
and AND3 (N2701, N2699, N1134, N125);
nor NOR4 (N2702, N2695, N2618, N1592, N3);
nand NAND2 (N2703, N2701, N2429);
not NOT1 (N2704, N2679);
not NOT1 (N2705, N2702);
nand NAND3 (N2706, N2698, N1554, N2134);
buf BUF1 (N2707, N2704);
and AND2 (N2708, N2707, N372);
not NOT1 (N2709, N2696);
nand NAND2 (N2710, N2697, N1987);
xor XOR2 (N2711, N2709, N769);
buf BUF1 (N2712, N2706);
nor NOR2 (N2713, N2712, N2231);
and AND3 (N2714, N2662, N1895, N2485);
and AND3 (N2715, N2693, N2352, N1220);
or OR4 (N2716, N2714, N2231, N1973, N559);
and AND4 (N2717, N2713, N1677, N1802, N2051);
buf BUF1 (N2718, N2711);
buf BUF1 (N2719, N2718);
or OR3 (N2720, N2719, N103, N999);
or OR2 (N2721, N2710, N2130);
nor NOR2 (N2722, N2716, N2086);
or OR3 (N2723, N2717, N1374, N2456);
or OR3 (N2724, N2720, N1986, N2521);
nand NAND4 (N2725, N2715, N1942, N1997, N167);
not NOT1 (N2726, N2705);
xor XOR2 (N2727, N2708, N575);
nand NAND2 (N2728, N2725, N1062);
and AND3 (N2729, N2700, N1488, N284);
not NOT1 (N2730, N2689);
nand NAND3 (N2731, N2724, N281, N1326);
nor NOR2 (N2732, N2726, N997);
and AND4 (N2733, N2722, N2524, N2379, N1305);
or OR4 (N2734, N2727, N209, N334, N1536);
buf BUF1 (N2735, N2732);
xor XOR2 (N2736, N2729, N2454);
or OR2 (N2737, N2730, N750);
nor NOR4 (N2738, N2736, N1462, N1138, N847);
xor XOR2 (N2739, N2737, N1316);
nand NAND2 (N2740, N2738, N1256);
buf BUF1 (N2741, N2733);
xor XOR2 (N2742, N2741, N423);
buf BUF1 (N2743, N2734);
and AND3 (N2744, N2740, N1048, N2681);
buf BUF1 (N2745, N2739);
xor XOR2 (N2746, N2723, N2740);
or OR4 (N2747, N2721, N1417, N126, N250);
xor XOR2 (N2748, N2746, N254);
not NOT1 (N2749, N2703);
nand NAND2 (N2750, N2748, N2530);
and AND4 (N2751, N2749, N1601, N627, N742);
and AND2 (N2752, N2731, N2538);
nand NAND4 (N2753, N2745, N1143, N1985, N703);
and AND4 (N2754, N2728, N1830, N1562, N2074);
buf BUF1 (N2755, N2747);
not NOT1 (N2756, N2742);
nand NAND4 (N2757, N2750, N2469, N2740, N1053);
or OR2 (N2758, N2752, N226);
or OR3 (N2759, N2751, N832, N1221);
not NOT1 (N2760, N2753);
xor XOR2 (N2761, N2754, N582);
and AND4 (N2762, N2761, N273, N246, N1240);
or OR4 (N2763, N2762, N1490, N2400, N852);
or OR3 (N2764, N2757, N1375, N1242);
nor NOR3 (N2765, N2735, N1863, N483);
or OR3 (N2766, N2744, N1000, N487);
nor NOR2 (N2767, N2755, N895);
and AND3 (N2768, N2764, N648, N1653);
xor XOR2 (N2769, N2760, N1604);
nor NOR3 (N2770, N2768, N2167, N1816);
not NOT1 (N2771, N2743);
and AND2 (N2772, N2756, N823);
or OR2 (N2773, N2759, N841);
and AND2 (N2774, N2763, N590);
nand NAND3 (N2775, N2765, N702, N2154);
buf BUF1 (N2776, N2770);
xor XOR2 (N2777, N2773, N112);
buf BUF1 (N2778, N2772);
nor NOR3 (N2779, N2771, N652, N130);
buf BUF1 (N2780, N2774);
xor XOR2 (N2781, N2777, N1468);
nand NAND2 (N2782, N2776, N2400);
nor NOR3 (N2783, N2758, N2509, N68);
nand NAND3 (N2784, N2783, N2305, N2071);
and AND2 (N2785, N2769, N1015);
not NOT1 (N2786, N2784);
buf BUF1 (N2787, N2778);
not NOT1 (N2788, N2780);
and AND3 (N2789, N2779, N796, N1812);
not NOT1 (N2790, N2767);
nand NAND4 (N2791, N2789, N2289, N2053, N1252);
xor XOR2 (N2792, N2782, N944);
nor NOR3 (N2793, N2786, N607, N2597);
and AND2 (N2794, N2787, N1298);
nand NAND3 (N2795, N2794, N315, N2525);
xor XOR2 (N2796, N2791, N362);
nand NAND3 (N2797, N2788, N2305, N2620);
xor XOR2 (N2798, N2797, N1061);
nand NAND3 (N2799, N2793, N1114, N1032);
and AND4 (N2800, N2781, N1055, N2356, N476);
buf BUF1 (N2801, N2799);
xor XOR2 (N2802, N2801, N1387);
buf BUF1 (N2803, N2800);
not NOT1 (N2804, N2796);
not NOT1 (N2805, N2775);
buf BUF1 (N2806, N2804);
nor NOR3 (N2807, N2802, N1794, N95);
and AND3 (N2808, N2798, N1830, N925);
not NOT1 (N2809, N2803);
buf BUF1 (N2810, N2805);
or OR2 (N2811, N2810, N1460);
or OR2 (N2812, N2766, N2420);
nor NOR3 (N2813, N2807, N2178, N2768);
nand NAND3 (N2814, N2812, N1576, N9);
nand NAND3 (N2815, N2792, N1366, N2300);
or OR3 (N2816, N2809, N806, N1495);
and AND4 (N2817, N2808, N2167, N2639, N479);
xor XOR2 (N2818, N2815, N59);
xor XOR2 (N2819, N2790, N83);
nor NOR2 (N2820, N2813, N1968);
or OR3 (N2821, N2819, N2307, N307);
nor NOR4 (N2822, N2816, N1103, N2488, N931);
nand NAND3 (N2823, N2822, N1596, N306);
buf BUF1 (N2824, N2795);
or OR2 (N2825, N2824, N1789);
nand NAND4 (N2826, N2818, N238, N1316, N526);
xor XOR2 (N2827, N2825, N1201);
not NOT1 (N2828, N2820);
nand NAND4 (N2829, N2806, N844, N241, N1967);
and AND4 (N2830, N2814, N659, N1015, N2412);
nand NAND2 (N2831, N2829, N2720);
buf BUF1 (N2832, N2811);
not NOT1 (N2833, N2830);
not NOT1 (N2834, N2832);
xor XOR2 (N2835, N2821, N859);
nand NAND4 (N2836, N2834, N1877, N819, N2777);
and AND2 (N2837, N2828, N1661);
or OR4 (N2838, N2835, N2095, N797, N2639);
xor XOR2 (N2839, N2826, N977);
nor NOR2 (N2840, N2833, N1580);
or OR2 (N2841, N2785, N2767);
or OR2 (N2842, N2838, N1208);
nand NAND4 (N2843, N2817, N162, N2314, N336);
nor NOR3 (N2844, N2841, N993, N2396);
not NOT1 (N2845, N2839);
not NOT1 (N2846, N2840);
or OR2 (N2847, N2823, N2609);
nand NAND2 (N2848, N2847, N1845);
or OR4 (N2849, N2842, N2679, N2819, N466);
buf BUF1 (N2850, N2827);
or OR3 (N2851, N2850, N2046, N1233);
not NOT1 (N2852, N2843);
buf BUF1 (N2853, N2849);
xor XOR2 (N2854, N2836, N973);
buf BUF1 (N2855, N2846);
xor XOR2 (N2856, N2831, N2007);
xor XOR2 (N2857, N2837, N271);
nand NAND4 (N2858, N2852, N1700, N2564, N67);
not NOT1 (N2859, N2855);
xor XOR2 (N2860, N2857, N755);
not NOT1 (N2861, N2845);
nand NAND4 (N2862, N2860, N2569, N1344, N312);
xor XOR2 (N2863, N2844, N1253);
buf BUF1 (N2864, N2862);
nor NOR3 (N2865, N2848, N2307, N2448);
xor XOR2 (N2866, N2861, N1180);
xor XOR2 (N2867, N2853, N1561);
nand NAND4 (N2868, N2854, N2319, N2350, N2602);
buf BUF1 (N2869, N2856);
buf BUF1 (N2870, N2868);
not NOT1 (N2871, N2863);
and AND2 (N2872, N2851, N1192);
xor XOR2 (N2873, N2872, N972);
not NOT1 (N2874, N2867);
xor XOR2 (N2875, N2874, N615);
not NOT1 (N2876, N2870);
nor NOR2 (N2877, N2859, N2772);
xor XOR2 (N2878, N2858, N979);
nand NAND3 (N2879, N2866, N2133, N2747);
not NOT1 (N2880, N2873);
xor XOR2 (N2881, N2865, N1005);
nor NOR2 (N2882, N2869, N420);
buf BUF1 (N2883, N2875);
and AND2 (N2884, N2877, N2864);
nor NOR2 (N2885, N2028, N1049);
buf BUF1 (N2886, N2879);
xor XOR2 (N2887, N2876, N401);
and AND4 (N2888, N2880, N2067, N628, N398);
nand NAND4 (N2889, N2885, N429, N2465, N935);
nor NOR2 (N2890, N2888, N2348);
xor XOR2 (N2891, N2884, N912);
nor NOR3 (N2892, N2889, N475, N2386);
and AND4 (N2893, N2881, N703, N1172, N2469);
not NOT1 (N2894, N2886);
nor NOR4 (N2895, N2892, N419, N2405, N2587);
nor NOR3 (N2896, N2882, N2069, N1655);
xor XOR2 (N2897, N2891, N613);
buf BUF1 (N2898, N2896);
and AND3 (N2899, N2878, N617, N654);
xor XOR2 (N2900, N2890, N331);
nor NOR2 (N2901, N2887, N2071);
nor NOR4 (N2902, N2898, N1583, N505, N312);
buf BUF1 (N2903, N2894);
buf BUF1 (N2904, N2897);
nand NAND4 (N2905, N2883, N1806, N1272, N1036);
or OR4 (N2906, N2871, N87, N785, N561);
and AND4 (N2907, N2905, N2283, N1001, N1367);
buf BUF1 (N2908, N2902);
buf BUF1 (N2909, N2900);
nor NOR3 (N2910, N2904, N92, N445);
or OR2 (N2911, N2903, N716);
xor XOR2 (N2912, N2899, N687);
and AND4 (N2913, N2911, N770, N690, N2536);
nor NOR3 (N2914, N2907, N212, N1737);
and AND2 (N2915, N2912, N684);
or OR2 (N2916, N2909, N413);
and AND2 (N2917, N2908, N1764);
xor XOR2 (N2918, N2901, N1465);
nand NAND2 (N2919, N2895, N1492);
not NOT1 (N2920, N2918);
or OR2 (N2921, N2906, N2480);
or OR3 (N2922, N2917, N135, N2118);
not NOT1 (N2923, N2910);
and AND4 (N2924, N2923, N1060, N2820, N1048);
not NOT1 (N2925, N2914);
nand NAND2 (N2926, N2921, N2027);
and AND4 (N2927, N2919, N477, N2030, N2570);
or OR3 (N2928, N2913, N487, N1562);
or OR2 (N2929, N2927, N596);
not NOT1 (N2930, N2920);
nand NAND2 (N2931, N2930, N2100);
or OR4 (N2932, N2931, N2251, N1666, N174);
xor XOR2 (N2933, N2932, N155);
buf BUF1 (N2934, N2928);
nand NAND4 (N2935, N2893, N2697, N1718, N1434);
and AND3 (N2936, N2924, N2398, N1911);
buf BUF1 (N2937, N2916);
and AND4 (N2938, N2934, N2156, N697, N98);
or OR3 (N2939, N2937, N1668, N1996);
nor NOR4 (N2940, N2939, N2030, N1713, N310);
buf BUF1 (N2941, N2933);
nor NOR2 (N2942, N2941, N1262);
nand NAND2 (N2943, N2926, N1221);
or OR2 (N2944, N2940, N2631);
nor NOR2 (N2945, N2944, N2467);
or OR4 (N2946, N2943, N510, N2306, N284);
buf BUF1 (N2947, N2945);
nand NAND3 (N2948, N2936, N2127, N2580);
nand NAND3 (N2949, N2925, N2916, N2925);
nand NAND4 (N2950, N2948, N628, N202, N2353);
nand NAND3 (N2951, N2946, N2881, N1012);
buf BUF1 (N2952, N2950);
nand NAND3 (N2953, N2935, N777, N77);
buf BUF1 (N2954, N2929);
nor NOR2 (N2955, N2952, N1359);
nor NOR3 (N2956, N2915, N1586, N738);
nor NOR4 (N2957, N2947, N2649, N11, N139);
buf BUF1 (N2958, N2949);
and AND3 (N2959, N2951, N1765, N1973);
nand NAND3 (N2960, N2942, N1654, N785);
not NOT1 (N2961, N2957);
or OR3 (N2962, N2954, N555, N1270);
buf BUF1 (N2963, N2953);
xor XOR2 (N2964, N2961, N2217);
and AND4 (N2965, N2964, N2934, N2823, N1904);
nand NAND2 (N2966, N2962, N1264);
or OR3 (N2967, N2958, N100, N387);
and AND3 (N2968, N2963, N2310, N1794);
or OR2 (N2969, N2938, N639);
nand NAND2 (N2970, N2967, N2813);
nand NAND2 (N2971, N2968, N372);
and AND2 (N2972, N2922, N645);
and AND2 (N2973, N2965, N2804);
buf BUF1 (N2974, N2973);
buf BUF1 (N2975, N2972);
nand NAND2 (N2976, N2966, N2439);
xor XOR2 (N2977, N2970, N662);
buf BUF1 (N2978, N2971);
or OR2 (N2979, N2974, N786);
buf BUF1 (N2980, N2977);
xor XOR2 (N2981, N2978, N1287);
nor NOR4 (N2982, N2955, N2423, N1723, N1006);
nor NOR3 (N2983, N2976, N2601, N1254);
or OR4 (N2984, N2979, N45, N1571, N162);
buf BUF1 (N2985, N2983);
not NOT1 (N2986, N2959);
not NOT1 (N2987, N2969);
nor NOR4 (N2988, N2986, N1062, N503, N1991);
nand NAND3 (N2989, N2988, N1875, N933);
and AND3 (N2990, N2985, N2184, N797);
or OR3 (N2991, N2987, N2051, N1729);
xor XOR2 (N2992, N2975, N2894);
or OR4 (N2993, N2981, N443, N2326, N668);
nand NAND4 (N2994, N2956, N2007, N2566, N1176);
buf BUF1 (N2995, N2989);
nor NOR3 (N2996, N2984, N2150, N2451);
nor NOR3 (N2997, N2982, N2667, N1173);
and AND3 (N2998, N2994, N2219, N1098);
nand NAND2 (N2999, N2995, N1726);
nand NAND3 (N3000, N2997, N1096, N1949);
nor NOR2 (N3001, N2993, N1128);
buf BUF1 (N3002, N3000);
xor XOR2 (N3003, N3001, N2000);
and AND3 (N3004, N2991, N1594, N2956);
buf BUF1 (N3005, N2980);
buf BUF1 (N3006, N2998);
buf BUF1 (N3007, N3003);
or OR4 (N3008, N3004, N581, N2869, N2714);
or OR3 (N3009, N2990, N2146, N2203);
or OR2 (N3010, N2960, N966);
buf BUF1 (N3011, N2996);
buf BUF1 (N3012, N2999);
nor NOR2 (N3013, N3008, N1492);
buf BUF1 (N3014, N3012);
and AND2 (N3015, N3002, N1184);
buf BUF1 (N3016, N3009);
and AND2 (N3017, N3006, N1172);
nand NAND4 (N3018, N3015, N2689, N2819, N194);
not NOT1 (N3019, N3017);
nor NOR4 (N3020, N3013, N1179, N2346, N972);
xor XOR2 (N3021, N3010, N2035);
buf BUF1 (N3022, N3020);
or OR3 (N3023, N3019, N478, N1372);
xor XOR2 (N3024, N3021, N1798);
buf BUF1 (N3025, N3016);
buf BUF1 (N3026, N3014);
xor XOR2 (N3027, N2992, N816);
or OR4 (N3028, N3018, N2899, N1359, N1943);
nand NAND3 (N3029, N3026, N1606, N1290);
nor NOR2 (N3030, N3025, N1656);
and AND4 (N3031, N3023, N1592, N533, N1913);
nand NAND2 (N3032, N3030, N670);
xor XOR2 (N3033, N3032, N2200);
or OR3 (N3034, N3022, N1807, N1175);
xor XOR2 (N3035, N3034, N621);
nor NOR2 (N3036, N3031, N1960);
buf BUF1 (N3037, N3024);
or OR3 (N3038, N3037, N2257, N206);
not NOT1 (N3039, N3029);
or OR3 (N3040, N3035, N644, N1221);
nand NAND4 (N3041, N3028, N207, N2142, N179);
and AND4 (N3042, N3027, N600, N2463, N1107);
not NOT1 (N3043, N3039);
not NOT1 (N3044, N3042);
buf BUF1 (N3045, N3007);
and AND4 (N3046, N3043, N1406, N2962, N2401);
not NOT1 (N3047, N3033);
or OR4 (N3048, N3041, N2186, N370, N2542);
xor XOR2 (N3049, N3036, N1638);
or OR3 (N3050, N3046, N2462, N2290);
and AND2 (N3051, N3011, N488);
buf BUF1 (N3052, N3040);
and AND4 (N3053, N3048, N1386, N2637, N1162);
and AND4 (N3054, N3051, N2671, N2710, N2192);
nor NOR4 (N3055, N3044, N1246, N1034, N2699);
and AND4 (N3056, N3055, N95, N1458, N2267);
and AND4 (N3057, N3049, N1361, N872, N122);
buf BUF1 (N3058, N3038);
and AND4 (N3059, N3005, N399, N3008, N278);
xor XOR2 (N3060, N3057, N537);
nand NAND2 (N3061, N3052, N1441);
buf BUF1 (N3062, N3059);
or OR3 (N3063, N3062, N1578, N149);
not NOT1 (N3064, N3045);
not NOT1 (N3065, N3058);
buf BUF1 (N3066, N3063);
buf BUF1 (N3067, N3053);
nor NOR3 (N3068, N3065, N2928, N64);
not NOT1 (N3069, N3068);
or OR2 (N3070, N3047, N123);
not NOT1 (N3071, N3067);
nand NAND4 (N3072, N3056, N737, N2238, N606);
buf BUF1 (N3073, N3054);
nand NAND4 (N3074, N3064, N343, N1682, N2833);
or OR2 (N3075, N3060, N1668);
nor NOR4 (N3076, N3075, N2898, N2091, N550);
nor NOR2 (N3077, N3076, N39);
or OR3 (N3078, N3050, N1254, N1407);
buf BUF1 (N3079, N3066);
nor NOR4 (N3080, N3061, N2247, N1248, N1330);
nand NAND2 (N3081, N3073, N2159);
nand NAND3 (N3082, N3079, N820, N2053);
not NOT1 (N3083, N3070);
xor XOR2 (N3084, N3071, N1894);
nor NOR2 (N3085, N3084, N224);
nor NOR3 (N3086, N3082, N2716, N2291);
not NOT1 (N3087, N3085);
not NOT1 (N3088, N3077);
or OR2 (N3089, N3087, N1320);
nand NAND4 (N3090, N3069, N2978, N936, N2227);
xor XOR2 (N3091, N3086, N781);
nand NAND4 (N3092, N3089, N580, N808, N683);
not NOT1 (N3093, N3081);
nor NOR4 (N3094, N3093, N2244, N2536, N564);
or OR4 (N3095, N3074, N1839, N1098, N2417);
xor XOR2 (N3096, N3092, N1386);
or OR4 (N3097, N3090, N1648, N1480, N1058);
xor XOR2 (N3098, N3091, N67);
or OR4 (N3099, N3080, N1120, N2454, N1310);
or OR3 (N3100, N3095, N2028, N1099);
nor NOR4 (N3101, N3083, N1246, N1375, N935);
nand NAND3 (N3102, N3101, N2859, N2647);
nor NOR2 (N3103, N3097, N618);
buf BUF1 (N3104, N3098);
or OR3 (N3105, N3102, N1166, N2286);
nor NOR4 (N3106, N3103, N1579, N2349, N2766);
and AND2 (N3107, N3096, N2041);
and AND2 (N3108, N3106, N123);
not NOT1 (N3109, N3107);
and AND4 (N3110, N3108, N2662, N2515, N2555);
or OR2 (N3111, N3110, N1416);
or OR2 (N3112, N3105, N1887);
nand NAND4 (N3113, N3078, N2870, N1377, N721);
nor NOR3 (N3114, N3072, N1254, N2892);
and AND3 (N3115, N3111, N663, N1435);
or OR2 (N3116, N3109, N1207);
not NOT1 (N3117, N3113);
xor XOR2 (N3118, N3117, N964);
nor NOR3 (N3119, N3088, N1675, N2552);
xor XOR2 (N3120, N3119, N733);
not NOT1 (N3121, N3115);
nand NAND4 (N3122, N3114, N113, N980, N907);
xor XOR2 (N3123, N3112, N808);
xor XOR2 (N3124, N3104, N658);
nor NOR2 (N3125, N3099, N2308);
nor NOR4 (N3126, N3094, N818, N2678, N2934);
not NOT1 (N3127, N3121);
buf BUF1 (N3128, N3126);
buf BUF1 (N3129, N3127);
not NOT1 (N3130, N3125);
or OR2 (N3131, N3118, N506);
buf BUF1 (N3132, N3124);
or OR4 (N3133, N3131, N1562, N22, N537);
not NOT1 (N3134, N3132);
not NOT1 (N3135, N3128);
xor XOR2 (N3136, N3129, N1286);
nor NOR3 (N3137, N3134, N1309, N2549);
or OR3 (N3138, N3120, N202, N2623);
nor NOR2 (N3139, N3116, N928);
not NOT1 (N3140, N3100);
or OR2 (N3141, N3137, N2560);
and AND4 (N3142, N3136, N2485, N2439, N26);
and AND3 (N3143, N3142, N1649, N553);
and AND3 (N3144, N3133, N1298, N2815);
or OR4 (N3145, N3130, N1627, N887, N2597);
not NOT1 (N3146, N3123);
not NOT1 (N3147, N3146);
nand NAND2 (N3148, N3138, N208);
nor NOR3 (N3149, N3140, N337, N1260);
nand NAND3 (N3150, N3145, N2391, N91);
and AND3 (N3151, N3148, N3048, N1379);
xor XOR2 (N3152, N3143, N589);
and AND2 (N3153, N3135, N1565);
xor XOR2 (N3154, N3151, N1929);
nand NAND2 (N3155, N3153, N3);
buf BUF1 (N3156, N3155);
buf BUF1 (N3157, N3156);
buf BUF1 (N3158, N3154);
xor XOR2 (N3159, N3147, N967);
xor XOR2 (N3160, N3152, N2198);
and AND2 (N3161, N3158, N2453);
nand NAND3 (N3162, N3141, N15, N2941);
nand NAND2 (N3163, N3161, N3060);
and AND4 (N3164, N3144, N358, N691, N2208);
nand NAND4 (N3165, N3163, N2980, N1872, N1251);
or OR2 (N3166, N3159, N179);
and AND4 (N3167, N3122, N403, N2347, N3100);
not NOT1 (N3168, N3167);
nand NAND2 (N3169, N3157, N860);
and AND2 (N3170, N3166, N1411);
or OR3 (N3171, N3168, N29, N1983);
not NOT1 (N3172, N3160);
or OR2 (N3173, N3149, N83);
buf BUF1 (N3174, N3139);
nor NOR2 (N3175, N3169, N3045);
nand NAND4 (N3176, N3174, N2431, N1433, N1333);
or OR2 (N3177, N3150, N2467);
nor NOR2 (N3178, N3162, N2343);
and AND3 (N3179, N3177, N1240, N757);
xor XOR2 (N3180, N3173, N2343);
or OR4 (N3181, N3165, N1228, N2768, N2989);
buf BUF1 (N3182, N3164);
or OR4 (N3183, N3179, N1278, N1917, N1486);
nor NOR3 (N3184, N3178, N395, N443);
or OR4 (N3185, N3170, N1800, N1468, N2294);
buf BUF1 (N3186, N3183);
and AND3 (N3187, N3172, N3118, N2374);
nand NAND4 (N3188, N3180, N257, N1226, N2027);
xor XOR2 (N3189, N3175, N1598);
nor NOR3 (N3190, N3188, N573, N229);
nor NOR3 (N3191, N3181, N3059, N2051);
not NOT1 (N3192, N3190);
buf BUF1 (N3193, N3187);
and AND4 (N3194, N3176, N31, N1206, N1200);
nand NAND4 (N3195, N3182, N3005, N3021, N2274);
not NOT1 (N3196, N3195);
nor NOR4 (N3197, N3192, N716, N348, N2986);
and AND4 (N3198, N3197, N2287, N26, N1592);
and AND2 (N3199, N3194, N2346);
xor XOR2 (N3200, N3198, N514);
nand NAND2 (N3201, N3189, N1970);
and AND4 (N3202, N3185, N245, N1150, N1110);
nand NAND2 (N3203, N3186, N987);
nand NAND4 (N3204, N3201, N417, N1167, N3095);
and AND4 (N3205, N3191, N825, N6, N3180);
or OR4 (N3206, N3203, N443, N1305, N2628);
not NOT1 (N3207, N3202);
and AND3 (N3208, N3171, N2370, N1657);
nand NAND4 (N3209, N3204, N2122, N2683, N864);
buf BUF1 (N3210, N3200);
and AND4 (N3211, N3207, N1324, N2533, N3078);
nor NOR3 (N3212, N3205, N1903, N1864);
buf BUF1 (N3213, N3211);
nand NAND4 (N3214, N3184, N2990, N1485, N2539);
nor NOR2 (N3215, N3206, N2318);
or OR3 (N3216, N3210, N1672, N581);
and AND4 (N3217, N3196, N1954, N2527, N1408);
nand NAND2 (N3218, N3215, N841);
not NOT1 (N3219, N3212);
nand NAND3 (N3220, N3208, N1632, N434);
nor NOR3 (N3221, N3209, N2608, N2394);
buf BUF1 (N3222, N3213);
xor XOR2 (N3223, N3220, N1122);
or OR4 (N3224, N3199, N2878, N2681, N2895);
nand NAND3 (N3225, N3218, N1198, N2774);
buf BUF1 (N3226, N3221);
nand NAND3 (N3227, N3214, N407, N83);
nand NAND3 (N3228, N3219, N2351, N2896);
not NOT1 (N3229, N3227);
buf BUF1 (N3230, N3226);
xor XOR2 (N3231, N3230, N85);
not NOT1 (N3232, N3228);
nor NOR4 (N3233, N3223, N2532, N2559, N1692);
or OR3 (N3234, N3233, N1988, N790);
buf BUF1 (N3235, N3222);
not NOT1 (N3236, N3193);
not NOT1 (N3237, N3231);
buf BUF1 (N3238, N3225);
nor NOR4 (N3239, N3224, N2112, N337, N1921);
and AND4 (N3240, N3238, N2426, N934, N2461);
or OR4 (N3241, N3240, N21, N2258, N2742);
or OR4 (N3242, N3241, N2103, N2885, N2589);
or OR4 (N3243, N3217, N362, N2201, N1196);
xor XOR2 (N3244, N3236, N253);
and AND3 (N3245, N3235, N2499, N1088);
xor XOR2 (N3246, N3237, N2673);
nand NAND2 (N3247, N3242, N1636);
nor NOR2 (N3248, N3246, N2746);
or OR3 (N3249, N3229, N1544, N332);
nand NAND2 (N3250, N3216, N2224);
nor NOR3 (N3251, N3243, N504, N1597);
xor XOR2 (N3252, N3245, N562);
or OR2 (N3253, N3249, N93);
buf BUF1 (N3254, N3244);
or OR3 (N3255, N3232, N268, N2202);
buf BUF1 (N3256, N3234);
buf BUF1 (N3257, N3254);
nor NOR3 (N3258, N3252, N2683, N1850);
buf BUF1 (N3259, N3247);
nor NOR2 (N3260, N3257, N1528);
nand NAND3 (N3261, N3251, N390, N2145);
nand NAND3 (N3262, N3258, N1289, N543);
not NOT1 (N3263, N3260);
or OR3 (N3264, N3256, N1605, N815);
xor XOR2 (N3265, N3248, N1994);
not NOT1 (N3266, N3255);
or OR4 (N3267, N3266, N1035, N2867, N1490);
xor XOR2 (N3268, N3263, N2146);
not NOT1 (N3269, N3267);
or OR2 (N3270, N3265, N2802);
not NOT1 (N3271, N3239);
and AND4 (N3272, N3259, N2475, N3056, N1573);
nand NAND3 (N3273, N3264, N814, N1218);
and AND2 (N3274, N3272, N2803);
and AND4 (N3275, N3269, N2447, N1434, N1955);
buf BUF1 (N3276, N3270);
and AND4 (N3277, N3271, N2113, N87, N1648);
or OR4 (N3278, N3277, N1093, N273, N279);
nor NOR2 (N3279, N3276, N2119);
nor NOR2 (N3280, N3273, N3241);
or OR3 (N3281, N3250, N2798, N777);
xor XOR2 (N3282, N3281, N426);
nor NOR3 (N3283, N3268, N2320, N752);
nand NAND3 (N3284, N3279, N291, N925);
or OR4 (N3285, N3284, N2379, N734, N2842);
buf BUF1 (N3286, N3262);
and AND4 (N3287, N3261, N18, N514, N3279);
nand NAND2 (N3288, N3274, N3092);
not NOT1 (N3289, N3280);
nor NOR2 (N3290, N3282, N2712);
or OR3 (N3291, N3253, N1721, N1735);
nor NOR4 (N3292, N3278, N1175, N321, N2586);
and AND3 (N3293, N3289, N1527, N2813);
xor XOR2 (N3294, N3292, N2997);
xor XOR2 (N3295, N3288, N2896);
and AND3 (N3296, N3294, N2034, N1156);
buf BUF1 (N3297, N3283);
xor XOR2 (N3298, N3285, N370);
not NOT1 (N3299, N3298);
and AND2 (N3300, N3286, N168);
nand NAND2 (N3301, N3299, N1497);
not NOT1 (N3302, N3297);
and AND2 (N3303, N3301, N524);
nor NOR4 (N3304, N3295, N2761, N2259, N114);
or OR4 (N3305, N3293, N2639, N2824, N145);
buf BUF1 (N3306, N3291);
or OR2 (N3307, N3287, N1954);
not NOT1 (N3308, N3302);
or OR2 (N3309, N3290, N2720);
nand NAND4 (N3310, N3303, N3173, N756, N723);
and AND4 (N3311, N3307, N1153, N122, N869);
nand NAND2 (N3312, N3296, N193);
and AND3 (N3313, N3305, N348, N1284);
and AND3 (N3314, N3311, N2172, N2279);
and AND3 (N3315, N3308, N172, N3223);
nand NAND3 (N3316, N3300, N1372, N2484);
nand NAND4 (N3317, N3316, N728, N764, N1106);
not NOT1 (N3318, N3313);
and AND4 (N3319, N3314, N1989, N10, N2471);
and AND3 (N3320, N3310, N3001, N3142);
xor XOR2 (N3321, N3317, N2342);
not NOT1 (N3322, N3318);
not NOT1 (N3323, N3275);
nand NAND2 (N3324, N3306, N1316);
not NOT1 (N3325, N3323);
or OR3 (N3326, N3309, N511, N67);
and AND2 (N3327, N3324, N740);
buf BUF1 (N3328, N3322);
nor NOR4 (N3329, N3312, N3203, N2644, N1103);
not NOT1 (N3330, N3327);
and AND2 (N3331, N3320, N1164);
buf BUF1 (N3332, N3328);
xor XOR2 (N3333, N3330, N294);
xor XOR2 (N3334, N3315, N1282);
nand NAND2 (N3335, N3334, N1779);
not NOT1 (N3336, N3332);
not NOT1 (N3337, N3333);
buf BUF1 (N3338, N3335);
nor NOR4 (N3339, N3304, N3287, N1774, N3154);
nor NOR3 (N3340, N3329, N1443, N997);
or OR4 (N3341, N3337, N2226, N472, N3185);
and AND2 (N3342, N3338, N68);
and AND3 (N3343, N3336, N2169, N3258);
or OR4 (N3344, N3331, N950, N2879, N2186);
nand NAND4 (N3345, N3325, N1616, N1948, N2756);
not NOT1 (N3346, N3340);
nor NOR3 (N3347, N3343, N2710, N2749);
not NOT1 (N3348, N3326);
and AND3 (N3349, N3339, N2114, N2781);
or OR2 (N3350, N3348, N1933);
not NOT1 (N3351, N3350);
buf BUF1 (N3352, N3342);
nand NAND4 (N3353, N3352, N2956, N2765, N1749);
not NOT1 (N3354, N3345);
not NOT1 (N3355, N3347);
or OR2 (N3356, N3353, N577);
buf BUF1 (N3357, N3321);
and AND3 (N3358, N3356, N2679, N2912);
xor XOR2 (N3359, N3358, N3032);
not NOT1 (N3360, N3351);
buf BUF1 (N3361, N3354);
xor XOR2 (N3362, N3349, N2899);
not NOT1 (N3363, N3361);
not NOT1 (N3364, N3357);
buf BUF1 (N3365, N3364);
or OR4 (N3366, N3355, N3002, N1050, N284);
nor NOR2 (N3367, N3365, N3255);
xor XOR2 (N3368, N3359, N510);
xor XOR2 (N3369, N3319, N2781);
nor NOR2 (N3370, N3346, N891);
or OR4 (N3371, N3344, N2932, N1281, N3307);
not NOT1 (N3372, N3369);
not NOT1 (N3373, N3368);
buf BUF1 (N3374, N3367);
xor XOR2 (N3375, N3371, N1829);
nor NOR3 (N3376, N3360, N877, N2145);
nor NOR4 (N3377, N3362, N2557, N1672, N3211);
nand NAND2 (N3378, N3373, N3365);
nand NAND3 (N3379, N3370, N2305, N2824);
nand NAND2 (N3380, N3375, N3043);
buf BUF1 (N3381, N3372);
buf BUF1 (N3382, N3381);
and AND4 (N3383, N3374, N1804, N1445, N2549);
nand NAND2 (N3384, N3341, N2616);
nand NAND2 (N3385, N3383, N1889);
nand NAND3 (N3386, N3376, N2066, N2477);
nand NAND2 (N3387, N3363, N454);
xor XOR2 (N3388, N3380, N2911);
nand NAND4 (N3389, N3387, N1606, N353, N1061);
xor XOR2 (N3390, N3385, N1378);
buf BUF1 (N3391, N3384);
and AND3 (N3392, N3389, N2576, N1705);
buf BUF1 (N3393, N3366);
nand NAND4 (N3394, N3379, N1033, N1881, N228);
or OR4 (N3395, N3391, N1760, N628, N3201);
or OR4 (N3396, N3386, N29, N3025, N2548);
buf BUF1 (N3397, N3382);
xor XOR2 (N3398, N3393, N2407);
nor NOR3 (N3399, N3394, N3068, N2942);
nand NAND3 (N3400, N3395, N2518, N1461);
and AND4 (N3401, N3378, N1049, N1589, N757);
xor XOR2 (N3402, N3397, N846);
not NOT1 (N3403, N3398);
or OR4 (N3404, N3399, N2857, N589, N656);
xor XOR2 (N3405, N3390, N538);
nand NAND4 (N3406, N3404, N1172, N3388, N434);
nand NAND3 (N3407, N2823, N830, N646);
and AND3 (N3408, N3396, N712, N2517);
buf BUF1 (N3409, N3405);
or OR3 (N3410, N3406, N2238, N3321);
buf BUF1 (N3411, N3409);
and AND2 (N3412, N3403, N1679);
nor NOR3 (N3413, N3411, N2266, N1096);
buf BUF1 (N3414, N3401);
xor XOR2 (N3415, N3414, N1355);
or OR3 (N3416, N3408, N1059, N3117);
and AND4 (N3417, N3377, N3123, N1172, N827);
or OR2 (N3418, N3412, N1881);
and AND3 (N3419, N3417, N2267, N3379);
nand NAND2 (N3420, N3418, N611);
xor XOR2 (N3421, N3413, N1263);
or OR4 (N3422, N3392, N1528, N841, N328);
and AND4 (N3423, N3410, N2105, N2188, N1325);
buf BUF1 (N3424, N3415);
nand NAND4 (N3425, N3419, N1715, N50, N3071);
nor NOR3 (N3426, N3420, N618, N2747);
and AND4 (N3427, N3402, N270, N1833, N1390);
xor XOR2 (N3428, N3427, N1054);
or OR4 (N3429, N3426, N2563, N3227, N2782);
nor NOR2 (N3430, N3424, N12);
or OR4 (N3431, N3400, N2976, N258, N3224);
buf BUF1 (N3432, N3425);
xor XOR2 (N3433, N3429, N575);
nand NAND4 (N3434, N3422, N1129, N2917, N849);
and AND4 (N3435, N3421, N90, N1452, N304);
xor XOR2 (N3436, N3432, N1941);
and AND4 (N3437, N3407, N2801, N1120, N2256);
buf BUF1 (N3438, N3431);
and AND4 (N3439, N3437, N239, N2856, N2493);
nor NOR4 (N3440, N3435, N2483, N1356, N2025);
or OR4 (N3441, N3428, N2328, N2544, N1863);
buf BUF1 (N3442, N3433);
and AND2 (N3443, N3442, N1369);
buf BUF1 (N3444, N3439);
xor XOR2 (N3445, N3423, N524);
not NOT1 (N3446, N3434);
buf BUF1 (N3447, N3416);
nand NAND4 (N3448, N3436, N3039, N343, N1265);
xor XOR2 (N3449, N3430, N1128);
and AND2 (N3450, N3448, N19);
not NOT1 (N3451, N3446);
buf BUF1 (N3452, N3443);
and AND3 (N3453, N3452, N3325, N286);
xor XOR2 (N3454, N3445, N3281);
not NOT1 (N3455, N3453);
xor XOR2 (N3456, N3444, N1597);
buf BUF1 (N3457, N3447);
and AND4 (N3458, N3451, N514, N2516, N3042);
nor NOR3 (N3459, N3458, N2250, N1258);
or OR2 (N3460, N3438, N2552);
nor NOR4 (N3461, N3441, N2645, N743, N347);
buf BUF1 (N3462, N3461);
not NOT1 (N3463, N3462);
buf BUF1 (N3464, N3457);
nand NAND3 (N3465, N3464, N1022, N3165);
xor XOR2 (N3466, N3459, N2821);
buf BUF1 (N3467, N3450);
and AND3 (N3468, N3454, N893, N2373);
buf BUF1 (N3469, N3465);
buf BUF1 (N3470, N3463);
and AND2 (N3471, N3460, N1567);
xor XOR2 (N3472, N3440, N2151);
nand NAND4 (N3473, N3449, N740, N2373, N1952);
nand NAND4 (N3474, N3471, N1350, N1499, N1482);
and AND3 (N3475, N3455, N485, N249);
nor NOR2 (N3476, N3466, N140);
or OR4 (N3477, N3476, N612, N2448, N1417);
xor XOR2 (N3478, N3468, N3080);
nand NAND4 (N3479, N3470, N165, N1858, N790);
and AND4 (N3480, N3469, N2110, N2285, N273);
buf BUF1 (N3481, N3472);
or OR3 (N3482, N3475, N1823, N3356);
xor XOR2 (N3483, N3480, N247);
or OR2 (N3484, N3477, N2173);
or OR4 (N3485, N3473, N705, N1654, N556);
xor XOR2 (N3486, N3482, N2270);
and AND4 (N3487, N3478, N3069, N802, N1191);
and AND4 (N3488, N3481, N2889, N2867, N511);
not NOT1 (N3489, N3485);
xor XOR2 (N3490, N3487, N1135);
not NOT1 (N3491, N3490);
nand NAND2 (N3492, N3484, N357);
and AND4 (N3493, N3483, N185, N3027, N164);
not NOT1 (N3494, N3474);
or OR3 (N3495, N3479, N2548, N1133);
xor XOR2 (N3496, N3493, N702);
buf BUF1 (N3497, N3491);
not NOT1 (N3498, N3488);
or OR3 (N3499, N3456, N1863, N1881);
or OR3 (N3500, N3497, N718, N3138);
and AND3 (N3501, N3495, N3342, N2017);
or OR4 (N3502, N3492, N2535, N2823, N964);
not NOT1 (N3503, N3467);
xor XOR2 (N3504, N3494, N157);
not NOT1 (N3505, N3501);
nand NAND3 (N3506, N3504, N2356, N376);
or OR3 (N3507, N3503, N1617, N2317);
not NOT1 (N3508, N3506);
nor NOR4 (N3509, N3496, N3384, N3406, N1946);
not NOT1 (N3510, N3508);
and AND2 (N3511, N3502, N746);
nand NAND2 (N3512, N3489, N3021);
and AND3 (N3513, N3512, N1415, N468);
buf BUF1 (N3514, N3513);
not NOT1 (N3515, N3514);
endmodule