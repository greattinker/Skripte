// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N411,N391,N381,N413,N409,N396,N387,N404,N414,N415;

nor NOR2 (N16, N4, N1);
and AND2 (N17, N9, N11);
and AND4 (N18, N4, N8, N9, N16);
nor NOR4 (N19, N7, N16, N8, N11);
not NOT1 (N20, N1);
nand NAND3 (N21, N18, N19, N15);
or OR3 (N22, N19, N11, N4);
and AND4 (N23, N4, N1, N22, N7);
xor XOR2 (N24, N19, N16);
nand NAND4 (N25, N11, N18, N4, N15);
xor XOR2 (N26, N19, N20);
xor XOR2 (N27, N16, N21);
nand NAND4 (N28, N7, N21, N3, N10);
not NOT1 (N29, N24);
not NOT1 (N30, N25);
xor XOR2 (N31, N1, N13);
buf BUF1 (N32, N27);
nand NAND4 (N33, N23, N6, N22, N5);
and AND3 (N34, N30, N3, N7);
or OR4 (N35, N23, N16, N31, N28);
not NOT1 (N36, N5);
nand NAND3 (N37, N15, N32, N20);
and AND4 (N38, N1, N12, N29, N16);
and AND4 (N39, N31, N36, N35, N9);
nor NOR3 (N40, N5, N19, N25);
buf BUF1 (N41, N4);
xor XOR2 (N42, N17, N11);
and AND2 (N43, N7, N39);
buf BUF1 (N44, N24);
not NOT1 (N45, N38);
and AND2 (N46, N41, N30);
nor NOR4 (N47, N44, N2, N3, N38);
or OR3 (N48, N42, N6, N4);
nand NAND3 (N49, N46, N45, N44);
xor XOR2 (N50, N13, N34);
nand NAND4 (N51, N47, N16, N24, N31);
and AND4 (N52, N9, N45, N9, N31);
nand NAND2 (N53, N37, N3);
xor XOR2 (N54, N50, N50);
and AND4 (N55, N43, N17, N7, N16);
and AND2 (N56, N26, N1);
xor XOR2 (N57, N33, N47);
not NOT1 (N58, N56);
nor NOR4 (N59, N58, N1, N56, N58);
xor XOR2 (N60, N54, N51);
nor NOR3 (N61, N8, N37, N1);
not NOT1 (N62, N59);
not NOT1 (N63, N60);
nor NOR4 (N64, N53, N32, N50, N14);
nor NOR3 (N65, N57, N36, N39);
nor NOR2 (N66, N52, N12);
xor XOR2 (N67, N61, N64);
xor XOR2 (N68, N8, N14);
or OR4 (N69, N62, N16, N60, N32);
xor XOR2 (N70, N49, N18);
buf BUF1 (N71, N70);
xor XOR2 (N72, N67, N48);
not NOT1 (N73, N41);
not NOT1 (N74, N71);
and AND2 (N75, N40, N32);
xor XOR2 (N76, N63, N20);
or OR2 (N77, N75, N63);
or OR4 (N78, N68, N20, N74, N28);
not NOT1 (N79, N33);
and AND4 (N80, N65, N18, N46, N47);
or OR3 (N81, N76, N34, N24);
buf BUF1 (N82, N79);
xor XOR2 (N83, N81, N2);
nor NOR4 (N84, N66, N13, N45, N72);
nor NOR3 (N85, N52, N37, N47);
not NOT1 (N86, N80);
buf BUF1 (N87, N86);
and AND2 (N88, N84, N22);
xor XOR2 (N89, N69, N2);
and AND2 (N90, N87, N26);
nand NAND2 (N91, N82, N62);
buf BUF1 (N92, N73);
or OR4 (N93, N91, N36, N58, N22);
nand NAND4 (N94, N55, N9, N77, N43);
and AND3 (N95, N4, N57, N18);
or OR3 (N96, N92, N38, N7);
xor XOR2 (N97, N96, N83);
and AND3 (N98, N84, N27, N22);
xor XOR2 (N99, N85, N41);
or OR4 (N100, N88, N74, N71, N22);
or OR3 (N101, N90, N91, N57);
xor XOR2 (N102, N98, N32);
nand NAND3 (N103, N100, N74, N54);
or OR3 (N104, N101, N73, N32);
and AND2 (N105, N102, N57);
xor XOR2 (N106, N89, N58);
not NOT1 (N107, N105);
nor NOR2 (N108, N94, N74);
nor NOR2 (N109, N104, N70);
nor NOR3 (N110, N93, N8, N76);
nand NAND4 (N111, N108, N108, N71, N54);
not NOT1 (N112, N106);
and AND3 (N113, N103, N95, N85);
or OR4 (N114, N93, N41, N68, N18);
nor NOR4 (N115, N112, N52, N105, N102);
xor XOR2 (N116, N110, N76);
buf BUF1 (N117, N111);
nand NAND2 (N118, N97, N101);
and AND4 (N119, N115, N51, N85, N114);
xor XOR2 (N120, N101, N91);
xor XOR2 (N121, N78, N64);
nand NAND2 (N122, N113, N108);
nand NAND4 (N123, N109, N86, N48, N59);
not NOT1 (N124, N99);
nand NAND3 (N125, N116, N62, N32);
xor XOR2 (N126, N119, N2);
buf BUF1 (N127, N123);
and AND4 (N128, N125, N33, N46, N58);
and AND4 (N129, N117, N91, N39, N112);
nand NAND4 (N130, N126, N43, N78, N74);
or OR4 (N131, N122, N32, N24, N67);
nand NAND2 (N132, N121, N106);
or OR3 (N133, N128, N69, N87);
nand NAND3 (N134, N131, N80, N60);
xor XOR2 (N135, N107, N44);
and AND4 (N136, N129, N69, N109, N18);
xor XOR2 (N137, N133, N44);
or OR3 (N138, N118, N18, N131);
and AND2 (N139, N134, N22);
not NOT1 (N140, N132);
nor NOR2 (N141, N139, N118);
buf BUF1 (N142, N141);
nor NOR3 (N143, N142, N135, N63);
or OR2 (N144, N87, N42);
not NOT1 (N145, N137);
nand NAND4 (N146, N130, N141, N130, N68);
buf BUF1 (N147, N143);
xor XOR2 (N148, N138, N132);
nor NOR2 (N149, N140, N112);
and AND4 (N150, N136, N129, N116, N106);
nand NAND3 (N151, N149, N37, N95);
buf BUF1 (N152, N120);
nand NAND2 (N153, N124, N49);
buf BUF1 (N154, N145);
and AND4 (N155, N148, N33, N116, N127);
or OR2 (N156, N131, N128);
buf BUF1 (N157, N152);
not NOT1 (N158, N157);
nor NOR4 (N159, N150, N69, N51, N10);
xor XOR2 (N160, N151, N109);
and AND4 (N161, N155, N88, N158, N53);
nor NOR2 (N162, N32, N65);
nor NOR4 (N163, N162, N17, N77, N67);
buf BUF1 (N164, N159);
buf BUF1 (N165, N161);
not NOT1 (N166, N153);
nand NAND4 (N167, N154, N121, N125, N108);
nand NAND4 (N168, N164, N142, N103, N31);
xor XOR2 (N169, N165, N43);
buf BUF1 (N170, N166);
and AND4 (N171, N156, N142, N137, N138);
buf BUF1 (N172, N160);
nor NOR2 (N173, N146, N90);
or OR3 (N174, N167, N1, N6);
nor NOR4 (N175, N173, N10, N30, N45);
and AND4 (N176, N174, N120, N131, N93);
not NOT1 (N177, N147);
or OR3 (N178, N176, N164, N123);
nand NAND3 (N179, N144, N52, N99);
xor XOR2 (N180, N172, N173);
nand NAND2 (N181, N170, N45);
and AND3 (N182, N178, N111, N177);
nand NAND4 (N183, N171, N85, N37, N106);
buf BUF1 (N184, N9);
nand NAND2 (N185, N175, N147);
buf BUF1 (N186, N179);
xor XOR2 (N187, N180, N107);
and AND4 (N188, N187, N179, N127, N8);
nand NAND2 (N189, N168, N80);
not NOT1 (N190, N185);
xor XOR2 (N191, N163, N167);
not NOT1 (N192, N186);
nand NAND3 (N193, N192, N155, N26);
and AND2 (N194, N188, N118);
and AND4 (N195, N191, N88, N13, N115);
and AND3 (N196, N183, N97, N87);
or OR4 (N197, N193, N20, N44, N193);
xor XOR2 (N198, N182, N107);
and AND4 (N199, N184, N100, N153, N147);
and AND2 (N200, N197, N52);
nor NOR3 (N201, N181, N54, N68);
and AND2 (N202, N196, N18);
and AND3 (N203, N190, N132, N4);
and AND3 (N204, N194, N36, N172);
and AND3 (N205, N198, N24, N51);
and AND4 (N206, N203, N18, N17, N1);
nand NAND2 (N207, N195, N105);
not NOT1 (N208, N169);
nand NAND3 (N209, N204, N120, N83);
nor NOR3 (N210, N199, N20, N175);
buf BUF1 (N211, N205);
and AND2 (N212, N208, N31);
and AND2 (N213, N206, N90);
and AND4 (N214, N210, N65, N75, N202);
or OR4 (N215, N209, N204, N69, N57);
and AND2 (N216, N123, N98);
or OR2 (N217, N201, N97);
buf BUF1 (N218, N214);
xor XOR2 (N219, N216, N5);
nor NOR2 (N220, N218, N54);
xor XOR2 (N221, N211, N5);
nor NOR2 (N222, N213, N46);
nand NAND4 (N223, N200, N111, N98, N49);
and AND3 (N224, N215, N3, N7);
xor XOR2 (N225, N221, N125);
and AND4 (N226, N225, N19, N105, N23);
xor XOR2 (N227, N217, N109);
or OR3 (N228, N219, N92, N201);
nor NOR4 (N229, N228, N114, N166, N201);
nand NAND2 (N230, N220, N4);
nor NOR2 (N231, N207, N97);
or OR4 (N232, N189, N209, N54, N85);
not NOT1 (N233, N222);
and AND4 (N234, N233, N204, N105, N201);
nand NAND4 (N235, N232, N111, N194, N198);
not NOT1 (N236, N224);
and AND4 (N237, N235, N224, N24, N218);
or OR3 (N238, N231, N112, N163);
nor NOR2 (N239, N236, N4);
nor NOR2 (N240, N237, N38);
nand NAND3 (N241, N239, N239, N133);
nand NAND3 (N242, N240, N85, N181);
nand NAND2 (N243, N223, N203);
and AND2 (N244, N229, N195);
nand NAND4 (N245, N212, N54, N33, N239);
nand NAND3 (N246, N238, N1, N60);
nand NAND2 (N247, N234, N151);
xor XOR2 (N248, N245, N144);
or OR4 (N249, N226, N103, N92, N234);
not NOT1 (N250, N248);
xor XOR2 (N251, N249, N57);
nor NOR2 (N252, N243, N202);
nor NOR2 (N253, N251, N127);
and AND4 (N254, N244, N244, N84, N236);
xor XOR2 (N255, N230, N118);
nor NOR3 (N256, N241, N217, N85);
buf BUF1 (N257, N255);
xor XOR2 (N258, N253, N51);
or OR2 (N259, N256, N239);
or OR3 (N260, N250, N59, N23);
nor NOR4 (N261, N247, N124, N198, N12);
or OR3 (N262, N246, N227, N147);
nand NAND2 (N263, N179, N173);
nand NAND2 (N264, N259, N6);
or OR2 (N265, N252, N204);
nor NOR2 (N266, N258, N228);
or OR3 (N267, N262, N196, N204);
or OR2 (N268, N242, N19);
nand NAND2 (N269, N263, N105);
and AND4 (N270, N266, N218, N43, N47);
nor NOR2 (N271, N265, N164);
not NOT1 (N272, N260);
xor XOR2 (N273, N261, N211);
buf BUF1 (N274, N264);
and AND2 (N275, N269, N137);
nor NOR3 (N276, N257, N37, N142);
xor XOR2 (N277, N270, N44);
not NOT1 (N278, N277);
not NOT1 (N279, N275);
not NOT1 (N280, N271);
xor XOR2 (N281, N267, N260);
not NOT1 (N282, N276);
xor XOR2 (N283, N268, N51);
xor XOR2 (N284, N283, N230);
not NOT1 (N285, N273);
buf BUF1 (N286, N272);
not NOT1 (N287, N284);
or OR4 (N288, N285, N287, N49, N122);
buf BUF1 (N289, N41);
or OR3 (N290, N274, N50, N65);
and AND2 (N291, N289, N173);
not NOT1 (N292, N288);
buf BUF1 (N293, N290);
xor XOR2 (N294, N286, N21);
or OR4 (N295, N278, N210, N150, N128);
not NOT1 (N296, N281);
xor XOR2 (N297, N292, N185);
xor XOR2 (N298, N282, N34);
buf BUF1 (N299, N296);
and AND4 (N300, N291, N188, N241, N139);
nor NOR4 (N301, N254, N298, N243, N1);
nand NAND2 (N302, N66, N297);
and AND3 (N303, N72, N82, N112);
nor NOR2 (N304, N279, N124);
or OR2 (N305, N303, N103);
not NOT1 (N306, N293);
and AND3 (N307, N299, N119, N129);
and AND2 (N308, N305, N307);
nand NAND4 (N309, N27, N25, N13, N28);
xor XOR2 (N310, N309, N59);
or OR4 (N311, N306, N66, N217, N130);
or OR2 (N312, N300, N103);
buf BUF1 (N313, N280);
xor XOR2 (N314, N310, N102);
buf BUF1 (N315, N302);
and AND3 (N316, N294, N7, N273);
or OR2 (N317, N313, N302);
not NOT1 (N318, N311);
xor XOR2 (N319, N295, N133);
xor XOR2 (N320, N314, N153);
and AND2 (N321, N312, N154);
or OR4 (N322, N321, N200, N220, N262);
nor NOR2 (N323, N308, N250);
buf BUF1 (N324, N316);
and AND3 (N325, N319, N165, N154);
and AND2 (N326, N324, N75);
nand NAND4 (N327, N323, N285, N71, N113);
or OR4 (N328, N325, N163, N185, N120);
and AND2 (N329, N320, N310);
not NOT1 (N330, N322);
xor XOR2 (N331, N301, N115);
or OR2 (N332, N318, N50);
xor XOR2 (N333, N315, N98);
and AND4 (N334, N328, N249, N35, N33);
or OR4 (N335, N329, N105, N287, N15);
or OR2 (N336, N330, N39);
nand NAND2 (N337, N333, N45);
nor NOR4 (N338, N326, N7, N204, N59);
and AND4 (N339, N332, N207, N68, N20);
buf BUF1 (N340, N317);
nor NOR2 (N341, N336, N231);
nand NAND4 (N342, N340, N167, N114, N54);
and AND3 (N343, N304, N129, N334);
buf BUF1 (N344, N261);
nor NOR2 (N345, N335, N255);
xor XOR2 (N346, N345, N316);
nand NAND4 (N347, N341, N124, N133, N183);
nor NOR2 (N348, N331, N262);
and AND4 (N349, N342, N117, N191, N158);
buf BUF1 (N350, N338);
or OR3 (N351, N350, N39, N168);
nand NAND4 (N352, N339, N244, N2, N72);
not NOT1 (N353, N343);
nor NOR2 (N354, N347, N261);
nand NAND2 (N355, N353, N89);
buf BUF1 (N356, N354);
buf BUF1 (N357, N327);
buf BUF1 (N358, N357);
not NOT1 (N359, N358);
and AND2 (N360, N355, N137);
nand NAND3 (N361, N348, N260, N310);
and AND4 (N362, N349, N277, N79, N344);
or OR2 (N363, N71, N342);
and AND4 (N364, N337, N175, N89, N276);
and AND4 (N365, N359, N292, N16, N260);
buf BUF1 (N366, N352);
buf BUF1 (N367, N365);
nand NAND3 (N368, N367, N137, N348);
buf BUF1 (N369, N346);
nor NOR3 (N370, N364, N261, N368);
nor NOR2 (N371, N237, N49);
or OR4 (N372, N361, N263, N32, N74);
buf BUF1 (N373, N362);
xor XOR2 (N374, N363, N258);
not NOT1 (N375, N373);
or OR2 (N376, N351, N280);
buf BUF1 (N377, N375);
not NOT1 (N378, N370);
nand NAND3 (N379, N376, N186, N73);
nor NOR3 (N380, N379, N152, N330);
not NOT1 (N381, N372);
not NOT1 (N382, N369);
or OR4 (N383, N356, N247, N67, N91);
or OR3 (N384, N382, N315, N17);
buf BUF1 (N385, N380);
not NOT1 (N386, N374);
buf BUF1 (N387, N378);
not NOT1 (N388, N386);
buf BUF1 (N389, N377);
not NOT1 (N390, N383);
or OR2 (N391, N366, N138);
and AND3 (N392, N389, N312, N232);
not NOT1 (N393, N388);
nor NOR3 (N394, N390, N221, N28);
nand NAND3 (N395, N385, N238, N337);
xor XOR2 (N396, N371, N118);
nand NAND4 (N397, N393, N57, N216, N142);
xor XOR2 (N398, N392, N301);
buf BUF1 (N399, N395);
and AND3 (N400, N360, N110, N383);
not NOT1 (N401, N394);
nor NOR4 (N402, N397, N284, N2, N172);
not NOT1 (N403, N402);
nor NOR4 (N404, N403, N87, N147, N83);
not NOT1 (N405, N400);
nor NOR3 (N406, N405, N83, N314);
xor XOR2 (N407, N398, N322);
nand NAND4 (N408, N407, N103, N375, N171);
xor XOR2 (N409, N406, N358);
nand NAND4 (N410, N384, N223, N21, N136);
buf BUF1 (N411, N408);
buf BUF1 (N412, N401);
nand NAND2 (N413, N399, N206);
nand NAND2 (N414, N412, N249);
buf BUF1 (N415, N410);
endmodule