// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N411,N421,N419,N407,N414,N404,N416,N401,N420,N422;

nand NAND3 (N23, N7, N2, N10);
and AND2 (N24, N11, N5);
nor NOR4 (N25, N12, N7, N7, N22);
nor NOR4 (N26, N19, N10, N21, N4);
not NOT1 (N27, N21);
buf BUF1 (N28, N7);
nand NAND3 (N29, N5, N2, N15);
not NOT1 (N30, N27);
buf BUF1 (N31, N5);
xor XOR2 (N32, N29, N27);
not NOT1 (N33, N13);
xor XOR2 (N34, N28, N20);
nand NAND2 (N35, N24, N20);
and AND3 (N36, N31, N3, N2);
xor XOR2 (N37, N20, N15);
nor NOR4 (N38, N37, N14, N9, N5);
nand NAND4 (N39, N35, N33, N23, N10);
buf BUF1 (N40, N14);
not NOT1 (N41, N21);
nand NAND3 (N42, N25, N40, N34);
xor XOR2 (N43, N37, N24);
xor XOR2 (N44, N27, N26);
buf BUF1 (N45, N21);
and AND4 (N46, N43, N23, N41, N27);
and AND2 (N47, N18, N23);
nor NOR4 (N48, N46, N13, N25, N47);
xor XOR2 (N49, N35, N32);
nor NOR4 (N50, N43, N25, N13, N46);
xor XOR2 (N51, N38, N28);
buf BUF1 (N52, N30);
not NOT1 (N53, N36);
not NOT1 (N54, N39);
nand NAND2 (N55, N54, N44);
nand NAND3 (N56, N44, N49, N24);
or OR4 (N57, N45, N17, N25, N39);
nand NAND3 (N58, N56, N29, N44);
not NOT1 (N59, N26);
nand NAND4 (N60, N58, N29, N46, N20);
nand NAND2 (N61, N51, N42);
nand NAND3 (N62, N6, N50, N32);
or OR4 (N63, N17, N28, N27, N21);
nor NOR2 (N64, N62, N6);
not NOT1 (N65, N52);
nor NOR3 (N66, N65, N20, N46);
nor NOR3 (N67, N59, N9, N51);
nand NAND4 (N68, N53, N31, N43, N66);
and AND4 (N69, N36, N14, N32, N6);
xor XOR2 (N70, N60, N38);
not NOT1 (N71, N64);
xor XOR2 (N72, N67, N13);
nor NOR3 (N73, N69, N16, N55);
xor XOR2 (N74, N16, N25);
nand NAND2 (N75, N68, N56);
and AND3 (N76, N63, N29, N32);
xor XOR2 (N77, N72, N33);
nor NOR3 (N78, N74, N51, N30);
xor XOR2 (N79, N77, N10);
nand NAND3 (N80, N70, N9, N73);
buf BUF1 (N81, N74);
or OR2 (N82, N75, N19);
not NOT1 (N83, N57);
buf BUF1 (N84, N82);
nor NOR4 (N85, N81, N75, N61, N33);
xor XOR2 (N86, N49, N49);
xor XOR2 (N87, N48, N74);
or OR2 (N88, N80, N81);
not NOT1 (N89, N84);
xor XOR2 (N90, N87, N89);
xor XOR2 (N91, N33, N62);
nand NAND4 (N92, N76, N86, N76, N62);
nand NAND3 (N93, N82, N39, N78);
nor NOR3 (N94, N13, N24, N91);
not NOT1 (N95, N79);
nor NOR2 (N96, N81, N3);
nor NOR3 (N97, N96, N29, N44);
and AND2 (N98, N94, N50);
not NOT1 (N99, N97);
nor NOR2 (N100, N85, N84);
buf BUF1 (N101, N71);
not NOT1 (N102, N95);
buf BUF1 (N103, N93);
not NOT1 (N104, N99);
and AND2 (N105, N102, N58);
buf BUF1 (N106, N90);
or OR2 (N107, N100, N46);
xor XOR2 (N108, N103, N49);
xor XOR2 (N109, N106, N69);
and AND4 (N110, N88, N14, N101, N39);
nand NAND2 (N111, N27, N36);
nor NOR2 (N112, N107, N84);
xor XOR2 (N113, N108, N80);
xor XOR2 (N114, N111, N63);
nor NOR3 (N115, N105, N114, N41);
or OR3 (N116, N60, N73, N57);
buf BUF1 (N117, N104);
and AND4 (N118, N115, N68, N76, N54);
nor NOR4 (N119, N116, N113, N102, N82);
nor NOR4 (N120, N104, N10, N17, N13);
nand NAND4 (N121, N119, N85, N35, N77);
nand NAND3 (N122, N83, N27, N15);
xor XOR2 (N123, N112, N65);
xor XOR2 (N124, N110, N57);
nor NOR2 (N125, N117, N97);
not NOT1 (N126, N118);
buf BUF1 (N127, N126);
nor NOR4 (N128, N120, N89, N110, N43);
nor NOR3 (N129, N122, N118, N107);
or OR2 (N130, N123, N79);
buf BUF1 (N131, N127);
nor NOR4 (N132, N124, N94, N51, N42);
and AND2 (N133, N130, N128);
or OR3 (N134, N129, N26, N20);
or OR2 (N135, N116, N39);
nand NAND2 (N136, N135, N35);
buf BUF1 (N137, N134);
or OR4 (N138, N131, N34, N31, N134);
buf BUF1 (N139, N136);
not NOT1 (N140, N121);
xor XOR2 (N141, N125, N27);
and AND4 (N142, N132, N30, N107, N81);
or OR3 (N143, N98, N123, N73);
and AND2 (N144, N139, N128);
xor XOR2 (N145, N143, N20);
xor XOR2 (N146, N144, N116);
nand NAND3 (N147, N137, N118, N7);
not NOT1 (N148, N146);
not NOT1 (N149, N148);
xor XOR2 (N150, N138, N118);
xor XOR2 (N151, N142, N135);
xor XOR2 (N152, N151, N143);
nand NAND3 (N153, N152, N26, N106);
nor NOR2 (N154, N140, N126);
nand NAND3 (N155, N150, N154, N33);
xor XOR2 (N156, N102, N49);
buf BUF1 (N157, N145);
nor NOR4 (N158, N153, N111, N12, N32);
buf BUF1 (N159, N158);
nor NOR3 (N160, N157, N95, N106);
and AND3 (N161, N109, N115, N154);
xor XOR2 (N162, N141, N126);
nor NOR3 (N163, N147, N29, N56);
buf BUF1 (N164, N156);
nor NOR2 (N165, N161, N93);
nor NOR3 (N166, N149, N17, N3);
and AND4 (N167, N163, N107, N30, N137);
xor XOR2 (N168, N159, N57);
not NOT1 (N169, N166);
nand NAND4 (N170, N162, N44, N153, N80);
and AND3 (N171, N169, N113, N108);
and AND3 (N172, N165, N37, N64);
xor XOR2 (N173, N164, N121);
not NOT1 (N174, N172);
or OR2 (N175, N155, N31);
not NOT1 (N176, N167);
buf BUF1 (N177, N174);
and AND3 (N178, N160, N167, N96);
or OR2 (N179, N168, N30);
and AND3 (N180, N178, N66, N22);
not NOT1 (N181, N173);
nor NOR4 (N182, N92, N56, N138, N114);
and AND4 (N183, N182, N161, N1, N96);
or OR4 (N184, N181, N117, N99, N164);
xor XOR2 (N185, N171, N145);
and AND4 (N186, N170, N176, N83, N35);
xor XOR2 (N187, N120, N127);
xor XOR2 (N188, N133, N125);
buf BUF1 (N189, N186);
and AND2 (N190, N187, N174);
nor NOR4 (N191, N179, N113, N17, N66);
xor XOR2 (N192, N183, N8);
nor NOR4 (N193, N177, N97, N89, N8);
buf BUF1 (N194, N190);
nor NOR3 (N195, N191, N39, N66);
and AND2 (N196, N188, N146);
and AND2 (N197, N189, N88);
nor NOR3 (N198, N184, N69, N179);
not NOT1 (N199, N195);
nor NOR3 (N200, N199, N18, N193);
nor NOR3 (N201, N36, N101, N86);
nor NOR3 (N202, N192, N47, N102);
nand NAND4 (N203, N185, N155, N53, N57);
buf BUF1 (N204, N175);
or OR4 (N205, N196, N114, N11, N24);
or OR4 (N206, N197, N188, N118, N172);
not NOT1 (N207, N202);
or OR2 (N208, N201, N186);
or OR4 (N209, N204, N201, N137, N171);
nand NAND3 (N210, N208, N179, N76);
nand NAND2 (N211, N209, N55);
xor XOR2 (N212, N205, N20);
and AND4 (N213, N180, N7, N138, N125);
not NOT1 (N214, N210);
buf BUF1 (N215, N203);
buf BUF1 (N216, N206);
and AND4 (N217, N216, N20, N63, N157);
xor XOR2 (N218, N211, N119);
not NOT1 (N219, N213);
buf BUF1 (N220, N214);
and AND2 (N221, N220, N217);
or OR3 (N222, N57, N25, N31);
or OR2 (N223, N198, N176);
and AND3 (N224, N207, N50, N134);
nor NOR2 (N225, N215, N197);
not NOT1 (N226, N224);
or OR2 (N227, N221, N154);
and AND3 (N228, N222, N192, N115);
not NOT1 (N229, N219);
and AND2 (N230, N200, N94);
nor NOR2 (N231, N225, N67);
and AND3 (N232, N231, N49, N124);
nor NOR4 (N233, N223, N194, N166, N106);
buf BUF1 (N234, N64);
and AND2 (N235, N227, N110);
buf BUF1 (N236, N212);
buf BUF1 (N237, N232);
or OR2 (N238, N228, N207);
or OR4 (N239, N229, N27, N20, N21);
and AND4 (N240, N226, N81, N218, N4);
nand NAND3 (N241, N69, N121, N96);
or OR4 (N242, N235, N42, N198, N80);
nand NAND4 (N243, N237, N208, N212, N65);
nand NAND2 (N244, N233, N162);
nor NOR2 (N245, N236, N37);
xor XOR2 (N246, N239, N200);
buf BUF1 (N247, N242);
not NOT1 (N248, N240);
or OR3 (N249, N243, N65, N177);
nand NAND2 (N250, N249, N110);
nor NOR4 (N251, N246, N63, N241, N94);
nor NOR4 (N252, N135, N193, N228, N27);
nand NAND3 (N253, N238, N201, N251);
not NOT1 (N254, N52);
not NOT1 (N255, N252);
nor NOR4 (N256, N248, N46, N160, N94);
and AND2 (N257, N250, N238);
nand NAND4 (N258, N253, N195, N236, N21);
nor NOR4 (N259, N255, N25, N141, N217);
buf BUF1 (N260, N259);
not NOT1 (N261, N244);
xor XOR2 (N262, N247, N56);
and AND2 (N263, N230, N120);
not NOT1 (N264, N260);
and AND2 (N265, N245, N53);
and AND3 (N266, N234, N158, N112);
xor XOR2 (N267, N266, N259);
and AND3 (N268, N264, N106, N185);
or OR4 (N269, N267, N186, N80, N144);
nand NAND4 (N270, N265, N38, N227, N265);
nor NOR3 (N271, N268, N142, N191);
nand NAND4 (N272, N263, N71, N185, N218);
nand NAND2 (N273, N272, N182);
nor NOR3 (N274, N254, N26, N238);
nor NOR4 (N275, N256, N67, N133, N243);
buf BUF1 (N276, N258);
nand NAND3 (N277, N271, N174, N211);
not NOT1 (N278, N261);
not NOT1 (N279, N275);
nand NAND3 (N280, N276, N191, N83);
buf BUF1 (N281, N280);
not NOT1 (N282, N270);
or OR2 (N283, N277, N113);
nor NOR2 (N284, N273, N236);
xor XOR2 (N285, N283, N247);
not NOT1 (N286, N257);
or OR3 (N287, N274, N83, N50);
not NOT1 (N288, N269);
or OR3 (N289, N278, N147, N180);
and AND3 (N290, N289, N112, N171);
not NOT1 (N291, N290);
nand NAND3 (N292, N287, N232, N234);
or OR4 (N293, N282, N144, N130, N153);
not NOT1 (N294, N288);
xor XOR2 (N295, N279, N188);
and AND3 (N296, N281, N60, N150);
or OR3 (N297, N296, N271, N17);
nand NAND4 (N298, N285, N5, N195, N276);
or OR3 (N299, N284, N131, N214);
not NOT1 (N300, N286);
buf BUF1 (N301, N293);
buf BUF1 (N302, N291);
xor XOR2 (N303, N300, N151);
buf BUF1 (N304, N295);
nand NAND4 (N305, N301, N46, N232, N280);
buf BUF1 (N306, N292);
nand NAND3 (N307, N262, N178, N272);
nand NAND2 (N308, N297, N303);
nand NAND3 (N309, N155, N221, N243);
not NOT1 (N310, N306);
nand NAND3 (N311, N304, N238, N154);
or OR4 (N312, N307, N141, N213, N12);
not NOT1 (N313, N305);
buf BUF1 (N314, N302);
nand NAND3 (N315, N312, N308, N256);
or OR3 (N316, N86, N42, N249);
xor XOR2 (N317, N309, N28);
xor XOR2 (N318, N314, N274);
not NOT1 (N319, N310);
buf BUF1 (N320, N294);
xor XOR2 (N321, N316, N36);
buf BUF1 (N322, N298);
nand NAND3 (N323, N317, N141, N3);
xor XOR2 (N324, N299, N131);
buf BUF1 (N325, N313);
nand NAND3 (N326, N319, N322, N149);
not NOT1 (N327, N315);
buf BUF1 (N328, N265);
xor XOR2 (N329, N326, N284);
buf BUF1 (N330, N329);
buf BUF1 (N331, N328);
and AND3 (N332, N311, N241, N205);
xor XOR2 (N333, N327, N44);
nor NOR4 (N334, N332, N165, N241, N280);
xor XOR2 (N335, N320, N54);
buf BUF1 (N336, N330);
not NOT1 (N337, N324);
not NOT1 (N338, N325);
nand NAND2 (N339, N323, N234);
or OR4 (N340, N318, N53, N175, N333);
and AND2 (N341, N180, N83);
not NOT1 (N342, N339);
and AND2 (N343, N321, N3);
xor XOR2 (N344, N331, N166);
and AND2 (N345, N341, N20);
or OR2 (N346, N345, N133);
xor XOR2 (N347, N334, N210);
xor XOR2 (N348, N338, N5);
or OR2 (N349, N335, N142);
or OR3 (N350, N349, N291, N127);
and AND4 (N351, N346, N273, N322, N104);
or OR2 (N352, N343, N18);
and AND3 (N353, N347, N200, N250);
not NOT1 (N354, N340);
and AND3 (N355, N342, N23, N84);
and AND4 (N356, N352, N236, N114, N110);
xor XOR2 (N357, N353, N160);
buf BUF1 (N358, N351);
nor NOR4 (N359, N354, N176, N86, N215);
not NOT1 (N360, N359);
and AND3 (N361, N357, N157, N14);
and AND2 (N362, N360, N316);
and AND4 (N363, N355, N246, N152, N247);
nor NOR2 (N364, N350, N109);
or OR3 (N365, N363, N246, N257);
nor NOR4 (N366, N336, N51, N313, N7);
buf BUF1 (N367, N337);
and AND2 (N368, N358, N315);
buf BUF1 (N369, N366);
or OR4 (N370, N356, N27, N184, N74);
or OR2 (N371, N368, N361);
or OR3 (N372, N249, N114, N2);
nand NAND4 (N373, N364, N46, N71, N38);
nand NAND2 (N374, N362, N262);
nand NAND4 (N375, N365, N111, N84, N11);
not NOT1 (N376, N370);
or OR3 (N377, N348, N25, N350);
and AND3 (N378, N377, N85, N121);
and AND4 (N379, N376, N230, N124, N166);
not NOT1 (N380, N375);
nand NAND4 (N381, N373, N10, N191, N87);
not NOT1 (N382, N378);
nand NAND3 (N383, N380, N122, N308);
nand NAND3 (N384, N367, N203, N188);
nor NOR4 (N385, N379, N51, N133, N273);
nor NOR3 (N386, N344, N223, N297);
not NOT1 (N387, N386);
or OR4 (N388, N383, N30, N148, N121);
xor XOR2 (N389, N381, N377);
or OR2 (N390, N387, N269);
and AND3 (N391, N372, N248, N262);
or OR4 (N392, N374, N330, N289, N175);
buf BUF1 (N393, N369);
xor XOR2 (N394, N389, N105);
and AND3 (N395, N385, N117, N274);
not NOT1 (N396, N391);
or OR4 (N397, N371, N19, N331, N313);
nor NOR3 (N398, N384, N129, N195);
and AND4 (N399, N393, N27, N303, N112);
nor NOR2 (N400, N398, N386);
and AND2 (N401, N399, N237);
xor XOR2 (N402, N388, N343);
nand NAND3 (N403, N394, N337, N220);
buf BUF1 (N404, N396);
nor NOR2 (N405, N397, N299);
or OR3 (N406, N382, N26, N8);
or OR4 (N407, N403, N28, N253, N245);
nand NAND4 (N408, N402, N163, N262, N201);
xor XOR2 (N409, N408, N23);
buf BUF1 (N410, N406);
not NOT1 (N411, N392);
nor NOR3 (N412, N395, N296, N227);
buf BUF1 (N413, N390);
not NOT1 (N414, N409);
xor XOR2 (N415, N400, N406);
buf BUF1 (N416, N412);
nand NAND4 (N417, N410, N348, N403, N355);
and AND3 (N418, N417, N181, N56);
and AND4 (N419, N418, N87, N357, N219);
and AND2 (N420, N413, N92);
or OR2 (N421, N405, N113);
not NOT1 (N422, N415);
endmodule