// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N618,N616,N612,N604,N603,N613,N585,N617,N598,N619;

xor XOR2 (N20, N14, N8);
nand NAND4 (N21, N19, N5, N4, N20);
not NOT1 (N22, N20);
nor NOR2 (N23, N12, N5);
buf BUF1 (N24, N2);
xor XOR2 (N25, N10, N16);
and AND4 (N26, N17, N12, N18, N18);
not NOT1 (N27, N19);
not NOT1 (N28, N2);
nand NAND2 (N29, N7, N23);
or OR4 (N30, N2, N23, N27, N26);
buf BUF1 (N31, N28);
and AND3 (N32, N25, N16, N21);
and AND2 (N33, N19, N32);
nand NAND4 (N34, N26, N14, N5, N1);
or OR3 (N35, N18, N25, N24);
or OR3 (N36, N24, N10, N34);
buf BUF1 (N37, N34);
nor NOR2 (N38, N26, N4);
xor XOR2 (N39, N29, N18);
buf BUF1 (N40, N16);
xor XOR2 (N41, N30, N8);
not NOT1 (N42, N41);
nor NOR3 (N43, N40, N39, N28);
or OR2 (N44, N41, N11);
nand NAND2 (N45, N22, N28);
not NOT1 (N46, N37);
and AND2 (N47, N31, N2);
or OR4 (N48, N38, N38, N20, N33);
nand NAND3 (N49, N43, N46, N6);
or OR4 (N50, N44, N34, N7, N44);
and AND3 (N51, N50, N22, N28);
or OR4 (N52, N50, N25, N34, N16);
buf BUF1 (N53, N18);
or OR4 (N54, N52, N36, N31, N39);
not NOT1 (N55, N3);
xor XOR2 (N56, N35, N41);
nor NOR3 (N57, N51, N28, N55);
not NOT1 (N58, N25);
nand NAND3 (N59, N45, N37, N24);
nor NOR4 (N60, N58, N25, N49, N6);
or OR3 (N61, N18, N44, N57);
xor XOR2 (N62, N45, N12);
not NOT1 (N63, N56);
and AND4 (N64, N54, N35, N17, N12);
not NOT1 (N65, N48);
buf BUF1 (N66, N42);
nor NOR2 (N67, N60, N14);
not NOT1 (N68, N53);
not NOT1 (N69, N63);
xor XOR2 (N70, N64, N49);
not NOT1 (N71, N68);
and AND3 (N72, N66, N24, N16);
and AND4 (N73, N62, N36, N27, N8);
buf BUF1 (N74, N47);
buf BUF1 (N75, N61);
xor XOR2 (N76, N75, N8);
nor NOR2 (N77, N67, N24);
and AND3 (N78, N73, N70, N2);
nand NAND4 (N79, N30, N18, N70, N69);
xor XOR2 (N80, N79, N60);
xor XOR2 (N81, N42, N59);
and AND3 (N82, N67, N73, N46);
not NOT1 (N83, N78);
nor NOR4 (N84, N77, N42, N48, N8);
or OR2 (N85, N80, N3);
or OR3 (N86, N84, N85, N72);
or OR4 (N87, N56, N85, N42, N57);
nand NAND4 (N88, N33, N83, N49, N42);
not NOT1 (N89, N39);
buf BUF1 (N90, N81);
or OR3 (N91, N74, N38, N90);
nand NAND2 (N92, N80, N40);
and AND3 (N93, N91, N37, N59);
or OR4 (N94, N86, N60, N22, N66);
buf BUF1 (N95, N89);
not NOT1 (N96, N87);
or OR2 (N97, N95, N42);
nand NAND4 (N98, N76, N12, N60, N20);
buf BUF1 (N99, N92);
or OR2 (N100, N65, N46);
buf BUF1 (N101, N82);
buf BUF1 (N102, N96);
not NOT1 (N103, N93);
and AND4 (N104, N99, N4, N30, N84);
not NOT1 (N105, N102);
nand NAND4 (N106, N71, N51, N90, N47);
and AND4 (N107, N88, N83, N52, N33);
buf BUF1 (N108, N94);
nand NAND2 (N109, N106, N22);
nand NAND3 (N110, N105, N71, N98);
nand NAND3 (N111, N32, N105, N57);
or OR3 (N112, N104, N109, N77);
buf BUF1 (N113, N83);
or OR3 (N114, N103, N57, N57);
nor NOR4 (N115, N113, N78, N83, N87);
buf BUF1 (N116, N100);
and AND2 (N117, N112, N114);
or OR3 (N118, N106, N24, N41);
and AND4 (N119, N110, N61, N71, N78);
nor NOR4 (N120, N107, N115, N68, N105);
buf BUF1 (N121, N72);
nand NAND2 (N122, N101, N103);
nand NAND3 (N123, N118, N27, N77);
xor XOR2 (N124, N97, N60);
or OR2 (N125, N123, N44);
or OR2 (N126, N117, N67);
xor XOR2 (N127, N116, N114);
or OR4 (N128, N126, N125, N60, N5);
xor XOR2 (N129, N121, N60);
not NOT1 (N130, N49);
buf BUF1 (N131, N129);
and AND3 (N132, N131, N25, N88);
nand NAND4 (N133, N132, N114, N71, N10);
buf BUF1 (N134, N133);
not NOT1 (N135, N130);
buf BUF1 (N136, N134);
buf BUF1 (N137, N135);
or OR4 (N138, N137, N89, N129, N98);
buf BUF1 (N139, N119);
buf BUF1 (N140, N136);
and AND3 (N141, N124, N105, N50);
or OR3 (N142, N122, N86, N75);
nand NAND4 (N143, N108, N64, N109, N35);
nand NAND4 (N144, N142, N141, N75, N105);
not NOT1 (N145, N18);
nor NOR2 (N146, N120, N76);
not NOT1 (N147, N127);
nand NAND4 (N148, N140, N134, N139, N18);
buf BUF1 (N149, N148);
not NOT1 (N150, N12);
nand NAND2 (N151, N145, N97);
buf BUF1 (N152, N138);
xor XOR2 (N153, N152, N135);
nand NAND2 (N154, N149, N86);
not NOT1 (N155, N153);
nand NAND4 (N156, N150, N70, N79, N132);
not NOT1 (N157, N128);
and AND3 (N158, N147, N147, N143);
nor NOR2 (N159, N55, N120);
and AND4 (N160, N155, N7, N148, N25);
not NOT1 (N161, N160);
and AND3 (N162, N154, N156, N113);
or OR4 (N163, N80, N19, N18, N105);
buf BUF1 (N164, N144);
and AND4 (N165, N162, N96, N8, N88);
or OR4 (N166, N146, N138, N1, N50);
xor XOR2 (N167, N158, N126);
or OR4 (N168, N165, N88, N84, N122);
buf BUF1 (N169, N151);
xor XOR2 (N170, N164, N148);
or OR2 (N171, N163, N30);
xor XOR2 (N172, N168, N85);
nand NAND3 (N173, N111, N133, N32);
and AND4 (N174, N166, N85, N85, N12);
or OR3 (N175, N172, N110, N150);
nor NOR3 (N176, N173, N59, N12);
buf BUF1 (N177, N157);
and AND2 (N178, N170, N147);
and AND2 (N179, N161, N110);
not NOT1 (N180, N179);
xor XOR2 (N181, N180, N65);
nor NOR2 (N182, N181, N158);
nand NAND2 (N183, N176, N83);
buf BUF1 (N184, N174);
nand NAND2 (N185, N178, N66);
nand NAND2 (N186, N171, N162);
nor NOR4 (N187, N177, N159, N32, N75);
nand NAND4 (N188, N28, N182, N128, N148);
and AND2 (N189, N141, N94);
not NOT1 (N190, N167);
or OR2 (N191, N188, N186);
nand NAND4 (N192, N55, N44, N7, N148);
buf BUF1 (N193, N175);
and AND4 (N194, N193, N105, N76, N147);
xor XOR2 (N195, N184, N78);
xor XOR2 (N196, N191, N61);
nand NAND3 (N197, N187, N176, N104);
nor NOR2 (N198, N196, N63);
nor NOR2 (N199, N169, N154);
xor XOR2 (N200, N197, N168);
nor NOR3 (N201, N195, N131, N186);
or OR4 (N202, N199, N146, N192, N87);
buf BUF1 (N203, N65);
nor NOR3 (N204, N185, N126, N128);
buf BUF1 (N205, N203);
and AND3 (N206, N204, N129, N166);
or OR2 (N207, N190, N66);
xor XOR2 (N208, N198, N81);
nor NOR4 (N209, N207, N188, N181, N141);
or OR4 (N210, N201, N182, N127, N114);
nand NAND2 (N211, N183, N146);
nor NOR3 (N212, N208, N179, N184);
nand NAND3 (N213, N206, N141, N203);
buf BUF1 (N214, N211);
buf BUF1 (N215, N212);
nand NAND3 (N216, N214, N53, N57);
not NOT1 (N217, N216);
or OR2 (N218, N189, N135);
not NOT1 (N219, N202);
and AND3 (N220, N215, N165, N53);
nor NOR2 (N221, N217, N112);
nor NOR3 (N222, N194, N56, N21);
not NOT1 (N223, N221);
nand NAND4 (N224, N205, N59, N70, N8);
nor NOR3 (N225, N213, N162, N219);
nor NOR4 (N226, N196, N29, N4, N198);
not NOT1 (N227, N218);
or OR2 (N228, N225, N114);
xor XOR2 (N229, N226, N176);
nor NOR2 (N230, N222, N192);
and AND3 (N231, N229, N41, N82);
or OR4 (N232, N200, N222, N45, N71);
buf BUF1 (N233, N209);
nand NAND4 (N234, N228, N200, N205, N76);
or OR2 (N235, N232, N136);
and AND2 (N236, N233, N75);
xor XOR2 (N237, N220, N127);
nand NAND3 (N238, N210, N162, N228);
and AND3 (N239, N230, N82, N211);
or OR4 (N240, N224, N30, N103, N119);
nand NAND4 (N241, N239, N112, N230, N185);
and AND3 (N242, N238, N19, N208);
nand NAND3 (N243, N242, N83, N241);
nor NOR2 (N244, N225, N201);
buf BUF1 (N245, N237);
xor XOR2 (N246, N244, N38);
xor XOR2 (N247, N236, N117);
nor NOR2 (N248, N227, N154);
not NOT1 (N249, N240);
buf BUF1 (N250, N223);
not NOT1 (N251, N249);
xor XOR2 (N252, N243, N90);
nand NAND4 (N253, N251, N173, N183, N25);
or OR2 (N254, N248, N180);
buf BUF1 (N255, N254);
not NOT1 (N256, N231);
nand NAND3 (N257, N252, N61, N158);
xor XOR2 (N258, N246, N170);
xor XOR2 (N259, N245, N138);
not NOT1 (N260, N250);
and AND4 (N261, N260, N39, N64, N19);
not NOT1 (N262, N255);
buf BUF1 (N263, N261);
or OR2 (N264, N235, N32);
nand NAND3 (N265, N262, N127, N182);
nor NOR2 (N266, N265, N70);
nand NAND3 (N267, N247, N166, N121);
or OR2 (N268, N266, N115);
and AND3 (N269, N256, N129, N104);
or OR2 (N270, N234, N83);
or OR3 (N271, N263, N62, N93);
or OR3 (N272, N253, N51, N94);
not NOT1 (N273, N271);
nand NAND3 (N274, N272, N8, N45);
nor NOR4 (N275, N258, N211, N162, N146);
buf BUF1 (N276, N273);
nor NOR4 (N277, N268, N176, N269, N74);
nor NOR4 (N278, N258, N186, N24, N5);
not NOT1 (N279, N270);
nand NAND4 (N280, N274, N163, N207, N54);
buf BUF1 (N281, N267);
nor NOR4 (N282, N259, N255, N158, N189);
nand NAND4 (N283, N278, N213, N18, N230);
xor XOR2 (N284, N281, N10);
nand NAND4 (N285, N283, N7, N206, N283);
nand NAND3 (N286, N285, N165, N116);
nor NOR4 (N287, N286, N156, N210, N282);
xor XOR2 (N288, N45, N76);
buf BUF1 (N289, N257);
not NOT1 (N290, N289);
not NOT1 (N291, N284);
xor XOR2 (N292, N287, N205);
or OR2 (N293, N276, N56);
and AND2 (N294, N264, N148);
not NOT1 (N295, N275);
not NOT1 (N296, N280);
xor XOR2 (N297, N279, N26);
buf BUF1 (N298, N291);
and AND3 (N299, N296, N127, N179);
buf BUF1 (N300, N299);
not NOT1 (N301, N293);
nand NAND2 (N302, N301, N60);
buf BUF1 (N303, N292);
nand NAND2 (N304, N302, N239);
or OR3 (N305, N300, N278, N118);
nor NOR3 (N306, N295, N237, N285);
xor XOR2 (N307, N297, N79);
xor XOR2 (N308, N288, N262);
and AND2 (N309, N307, N265);
buf BUF1 (N310, N309);
nand NAND4 (N311, N304, N87, N191, N48);
xor XOR2 (N312, N294, N268);
not NOT1 (N313, N306);
xor XOR2 (N314, N305, N6);
buf BUF1 (N315, N311);
or OR3 (N316, N310, N214, N10);
not NOT1 (N317, N298);
not NOT1 (N318, N303);
and AND3 (N319, N308, N236, N223);
nor NOR4 (N320, N277, N58, N111, N297);
not NOT1 (N321, N314);
nand NAND4 (N322, N315, N282, N207, N274);
or OR3 (N323, N320, N127, N24);
not NOT1 (N324, N322);
nor NOR4 (N325, N316, N237, N82, N293);
and AND3 (N326, N312, N37, N63);
xor XOR2 (N327, N324, N223);
xor XOR2 (N328, N290, N249);
xor XOR2 (N329, N313, N203);
xor XOR2 (N330, N317, N115);
nand NAND4 (N331, N321, N196, N283, N48);
or OR4 (N332, N323, N47, N266, N268);
nor NOR2 (N333, N327, N30);
nand NAND2 (N334, N331, N283);
not NOT1 (N335, N326);
nand NAND4 (N336, N325, N177, N30, N274);
nor NOR2 (N337, N334, N19);
nand NAND4 (N338, N333, N232, N71, N39);
buf BUF1 (N339, N335);
xor XOR2 (N340, N339, N103);
xor XOR2 (N341, N336, N229);
and AND2 (N342, N337, N13);
nand NAND3 (N343, N329, N29, N328);
or OR4 (N344, N207, N281, N21, N21);
xor XOR2 (N345, N332, N329);
nand NAND3 (N346, N344, N82, N131);
or OR4 (N347, N345, N169, N236, N93);
and AND2 (N348, N346, N56);
xor XOR2 (N349, N341, N280);
or OR2 (N350, N343, N349);
buf BUF1 (N351, N124);
buf BUF1 (N352, N342);
or OR2 (N353, N347, N29);
and AND4 (N354, N338, N99, N75, N335);
xor XOR2 (N355, N354, N84);
and AND2 (N356, N340, N316);
and AND4 (N357, N351, N293, N194, N271);
buf BUF1 (N358, N353);
or OR4 (N359, N355, N276, N236, N80);
buf BUF1 (N360, N348);
xor XOR2 (N361, N319, N315);
buf BUF1 (N362, N357);
nor NOR4 (N363, N358, N166, N41, N32);
nor NOR4 (N364, N360, N215, N348, N212);
not NOT1 (N365, N356);
buf BUF1 (N366, N364);
nor NOR4 (N367, N330, N324, N211, N97);
nor NOR4 (N368, N350, N273, N174, N90);
not NOT1 (N369, N359);
nor NOR2 (N370, N367, N249);
nor NOR3 (N371, N363, N352, N83);
buf BUF1 (N372, N348);
and AND2 (N373, N362, N180);
buf BUF1 (N374, N366);
not NOT1 (N375, N369);
or OR4 (N376, N375, N343, N226, N59);
or OR2 (N377, N374, N296);
not NOT1 (N378, N368);
nand NAND4 (N379, N373, N322, N31, N225);
buf BUF1 (N380, N377);
or OR2 (N381, N379, N376);
not NOT1 (N382, N156);
buf BUF1 (N383, N381);
buf BUF1 (N384, N371);
buf BUF1 (N385, N372);
or OR2 (N386, N384, N271);
xor XOR2 (N387, N370, N112);
nor NOR2 (N388, N361, N219);
buf BUF1 (N389, N318);
or OR3 (N390, N365, N42, N236);
and AND2 (N391, N389, N311);
xor XOR2 (N392, N382, N303);
or OR4 (N393, N391, N9, N4, N257);
or OR3 (N394, N392, N252, N241);
nor NOR2 (N395, N387, N147);
buf BUF1 (N396, N390);
nor NOR4 (N397, N380, N367, N331, N358);
not NOT1 (N398, N378);
buf BUF1 (N399, N395);
buf BUF1 (N400, N393);
and AND3 (N401, N400, N316, N334);
buf BUF1 (N402, N383);
xor XOR2 (N403, N394, N367);
xor XOR2 (N404, N398, N16);
xor XOR2 (N405, N404, N54);
buf BUF1 (N406, N402);
nand NAND2 (N407, N403, N38);
xor XOR2 (N408, N399, N202);
nor NOR4 (N409, N386, N375, N12, N127);
nor NOR2 (N410, N397, N90);
or OR4 (N411, N388, N132, N93, N124);
nand NAND2 (N412, N409, N19);
xor XOR2 (N413, N407, N33);
nand NAND2 (N414, N413, N191);
xor XOR2 (N415, N411, N139);
not NOT1 (N416, N414);
nand NAND2 (N417, N412, N105);
xor XOR2 (N418, N401, N65);
not NOT1 (N419, N417);
or OR4 (N420, N416, N365, N297, N27);
and AND3 (N421, N418, N364, N138);
nand NAND4 (N422, N405, N243, N9, N245);
xor XOR2 (N423, N408, N74);
xor XOR2 (N424, N410, N76);
and AND4 (N425, N423, N201, N344, N383);
nand NAND2 (N426, N421, N64);
nand NAND4 (N427, N426, N248, N366, N274);
not NOT1 (N428, N406);
buf BUF1 (N429, N428);
nor NOR3 (N430, N425, N58, N164);
and AND3 (N431, N424, N372, N362);
and AND2 (N432, N427, N272);
buf BUF1 (N433, N422);
not NOT1 (N434, N430);
xor XOR2 (N435, N420, N273);
or OR2 (N436, N385, N340);
not NOT1 (N437, N429);
and AND2 (N438, N415, N284);
or OR3 (N439, N433, N245, N169);
xor XOR2 (N440, N436, N429);
xor XOR2 (N441, N437, N44);
and AND3 (N442, N435, N203, N341);
buf BUF1 (N443, N438);
buf BUF1 (N444, N442);
xor XOR2 (N445, N431, N120);
buf BUF1 (N446, N434);
nand NAND3 (N447, N441, N439, N26);
and AND4 (N448, N150, N109, N413, N414);
and AND2 (N449, N440, N79);
not NOT1 (N450, N432);
xor XOR2 (N451, N448, N71);
xor XOR2 (N452, N450, N85);
or OR3 (N453, N396, N133, N312);
buf BUF1 (N454, N453);
nor NOR2 (N455, N447, N386);
nand NAND3 (N456, N454, N26, N365);
xor XOR2 (N457, N443, N284);
or OR3 (N458, N446, N203, N84);
buf BUF1 (N459, N458);
or OR4 (N460, N457, N6, N133, N417);
nor NOR3 (N461, N455, N91, N413);
nor NOR4 (N462, N449, N55, N15, N372);
nor NOR3 (N463, N444, N294, N114);
or OR3 (N464, N445, N292, N262);
nor NOR2 (N465, N419, N249);
nand NAND2 (N466, N451, N290);
nor NOR4 (N467, N464, N49, N348, N275);
nand NAND2 (N468, N462, N325);
and AND2 (N469, N468, N410);
nor NOR4 (N470, N469, N284, N194, N320);
or OR4 (N471, N470, N174, N463, N61);
buf BUF1 (N472, N274);
nor NOR3 (N473, N467, N37, N80);
and AND2 (N474, N472, N229);
not NOT1 (N475, N459);
buf BUF1 (N476, N460);
buf BUF1 (N477, N474);
and AND4 (N478, N465, N86, N34, N129);
nor NOR3 (N479, N475, N15, N97);
not NOT1 (N480, N473);
xor XOR2 (N481, N456, N475);
not NOT1 (N482, N477);
xor XOR2 (N483, N478, N85);
xor XOR2 (N484, N482, N230);
or OR3 (N485, N471, N154, N235);
xor XOR2 (N486, N476, N360);
nor NOR4 (N487, N484, N185, N84, N165);
and AND2 (N488, N483, N265);
buf BUF1 (N489, N487);
nand NAND4 (N490, N481, N224, N401, N49);
nor NOR4 (N491, N488, N160, N403, N50);
and AND2 (N492, N461, N153);
nand NAND3 (N493, N466, N270, N95);
or OR2 (N494, N490, N440);
and AND4 (N495, N492, N284, N205, N202);
and AND4 (N496, N489, N490, N239, N458);
xor XOR2 (N497, N485, N200);
nand NAND4 (N498, N493, N99, N359, N314);
nor NOR3 (N499, N491, N244, N202);
or OR4 (N500, N452, N443, N54, N18);
nor NOR4 (N501, N495, N161, N436, N314);
and AND3 (N502, N496, N110, N209);
or OR3 (N503, N501, N362, N30);
not NOT1 (N504, N500);
not NOT1 (N505, N479);
xor XOR2 (N506, N480, N72);
xor XOR2 (N507, N502, N389);
xor XOR2 (N508, N507, N465);
nor NOR4 (N509, N497, N79, N270, N157);
buf BUF1 (N510, N499);
and AND4 (N511, N510, N284, N110, N234);
nor NOR3 (N512, N509, N487, N379);
not NOT1 (N513, N512);
and AND3 (N514, N503, N48, N254);
and AND4 (N515, N514, N448, N13, N352);
nor NOR4 (N516, N486, N300, N395, N1);
buf BUF1 (N517, N506);
nand NAND4 (N518, N513, N470, N215, N455);
xor XOR2 (N519, N494, N330);
not NOT1 (N520, N504);
or OR3 (N521, N505, N187, N53);
and AND2 (N522, N515, N98);
nand NAND3 (N523, N519, N347, N79);
nand NAND3 (N524, N522, N112, N495);
or OR3 (N525, N523, N382, N107);
nand NAND2 (N526, N498, N421);
nand NAND2 (N527, N518, N133);
nand NAND2 (N528, N516, N317);
buf BUF1 (N529, N525);
nand NAND3 (N530, N520, N350, N4);
or OR2 (N531, N517, N167);
xor XOR2 (N532, N529, N337);
nor NOR4 (N533, N521, N298, N92, N22);
nand NAND3 (N534, N508, N368, N346);
buf BUF1 (N535, N526);
nor NOR4 (N536, N524, N151, N191, N475);
and AND2 (N537, N530, N257);
and AND2 (N538, N534, N400);
and AND3 (N539, N535, N228, N308);
or OR4 (N540, N527, N299, N365, N223);
and AND2 (N541, N511, N220);
or OR2 (N542, N538, N391);
not NOT1 (N543, N531);
or OR4 (N544, N543, N281, N82, N118);
or OR2 (N545, N541, N66);
xor XOR2 (N546, N537, N346);
or OR3 (N547, N542, N19, N390);
and AND3 (N548, N528, N121, N163);
and AND4 (N549, N533, N52, N526, N422);
and AND3 (N550, N547, N50, N133);
or OR3 (N551, N546, N51, N453);
buf BUF1 (N552, N550);
or OR4 (N553, N549, N213, N333, N214);
not NOT1 (N554, N552);
and AND2 (N555, N553, N115);
not NOT1 (N556, N544);
buf BUF1 (N557, N536);
not NOT1 (N558, N557);
buf BUF1 (N559, N532);
buf BUF1 (N560, N559);
buf BUF1 (N561, N545);
xor XOR2 (N562, N540, N365);
not NOT1 (N563, N560);
nand NAND2 (N564, N561, N146);
nand NAND2 (N565, N563, N159);
nor NOR3 (N566, N548, N407, N309);
and AND3 (N567, N556, N560, N413);
xor XOR2 (N568, N551, N13);
or OR3 (N569, N565, N113, N308);
or OR2 (N570, N539, N27);
nand NAND3 (N571, N554, N388, N480);
not NOT1 (N572, N566);
buf BUF1 (N573, N571);
not NOT1 (N574, N567);
or OR4 (N575, N555, N81, N210, N428);
or OR4 (N576, N572, N327, N415, N529);
buf BUF1 (N577, N573);
buf BUF1 (N578, N558);
nand NAND3 (N579, N569, N70, N423);
nand NAND4 (N580, N574, N340, N58, N560);
nor NOR4 (N581, N579, N440, N255, N541);
not NOT1 (N582, N576);
and AND4 (N583, N580, N69, N244, N565);
or OR2 (N584, N581, N165);
not NOT1 (N585, N575);
nand NAND2 (N586, N562, N242);
or OR2 (N587, N583, N537);
and AND2 (N588, N564, N314);
and AND3 (N589, N582, N310, N3);
xor XOR2 (N590, N588, N212);
nand NAND2 (N591, N568, N300);
or OR2 (N592, N570, N112);
nor NOR2 (N593, N586, N50);
and AND2 (N594, N584, N250);
nor NOR3 (N595, N590, N388, N192);
not NOT1 (N596, N589);
not NOT1 (N597, N592);
nor NOR4 (N598, N593, N124, N22, N349);
buf BUF1 (N599, N578);
xor XOR2 (N600, N591, N472);
and AND4 (N601, N600, N431, N415, N281);
nand NAND3 (N602, N594, N442, N516);
xor XOR2 (N603, N595, N341);
nand NAND3 (N604, N601, N321, N164);
nand NAND3 (N605, N597, N89, N470);
xor XOR2 (N606, N599, N491);
nor NOR2 (N607, N587, N324);
buf BUF1 (N608, N602);
nor NOR3 (N609, N577, N154, N118);
or OR4 (N610, N606, N3, N386, N125);
or OR2 (N611, N608, N117);
and AND4 (N612, N610, N410, N117, N362);
buf BUF1 (N613, N596);
nand NAND2 (N614, N605, N534);
nand NAND3 (N615, N611, N89, N232);
xor XOR2 (N616, N614, N52);
xor XOR2 (N617, N609, N60);
nor NOR4 (N618, N607, N119, N463, N445);
xor XOR2 (N619, N615, N509);
endmodule