// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N3018,N2995,N2999,N3017,N3011,N3001,N3016,N3014,N3020,N3022;

buf BUF1 (N23, N19);
nor NOR2 (N24, N13, N2);
not NOT1 (N25, N2);
or OR3 (N26, N18, N22, N20);
nor NOR4 (N27, N5, N12, N24, N26);
nand NAND4 (N28, N17, N16, N18, N1);
nor NOR4 (N29, N13, N9, N6, N20);
nor NOR3 (N30, N12, N20, N11);
nand NAND4 (N31, N17, N25, N19, N21);
and AND4 (N32, N3, N2, N14, N26);
xor XOR2 (N33, N16, N24);
nor NOR2 (N34, N5, N3);
and AND3 (N35, N30, N12, N2);
or OR3 (N36, N21, N24, N31);
not NOT1 (N37, N36);
or OR4 (N38, N17, N33, N32, N24);
nand NAND4 (N39, N27, N15, N24, N33);
or OR3 (N40, N35, N30, N29);
or OR4 (N41, N30, N38, N13, N4);
and AND2 (N42, N22, N9);
and AND4 (N43, N29, N36, N3, N2);
buf BUF1 (N44, N19);
nand NAND3 (N45, N34, N10, N34);
not NOT1 (N46, N28);
buf BUF1 (N47, N44);
buf BUF1 (N48, N47);
or OR2 (N49, N39, N31);
buf BUF1 (N50, N45);
nor NOR3 (N51, N41, N36, N24);
buf BUF1 (N52, N23);
nand NAND2 (N53, N42, N45);
and AND2 (N54, N53, N35);
not NOT1 (N55, N50);
buf BUF1 (N56, N54);
nor NOR3 (N57, N49, N38, N6);
buf BUF1 (N58, N57);
nand NAND4 (N59, N46, N7, N15, N28);
and AND2 (N60, N52, N49);
and AND3 (N61, N55, N14, N24);
and AND3 (N62, N58, N33, N60);
and AND2 (N63, N15, N39);
or OR2 (N64, N40, N21);
xor XOR2 (N65, N62, N36);
buf BUF1 (N66, N64);
not NOT1 (N67, N59);
or OR2 (N68, N63, N52);
and AND2 (N69, N66, N7);
not NOT1 (N70, N56);
nor NOR2 (N71, N68, N5);
and AND2 (N72, N65, N47);
or OR3 (N73, N72, N69, N32);
and AND2 (N74, N20, N60);
nor NOR3 (N75, N74, N23, N52);
nor NOR3 (N76, N71, N17, N58);
not NOT1 (N77, N67);
nand NAND4 (N78, N43, N17, N14, N9);
nand NAND3 (N79, N61, N37, N48);
nand NAND4 (N80, N51, N44, N17, N71);
or OR2 (N81, N42, N42);
nand NAND4 (N82, N29, N16, N17, N74);
xor XOR2 (N83, N73, N34);
not NOT1 (N84, N78);
or OR2 (N85, N81, N82);
or OR4 (N86, N20, N39, N4, N1);
buf BUF1 (N87, N76);
or OR3 (N88, N85, N6, N14);
buf BUF1 (N89, N79);
not NOT1 (N90, N75);
xor XOR2 (N91, N77, N90);
or OR3 (N92, N57, N36, N37);
nor NOR4 (N93, N84, N53, N26, N52);
or OR3 (N94, N92, N72, N30);
xor XOR2 (N95, N83, N60);
buf BUF1 (N96, N87);
buf BUF1 (N97, N88);
nand NAND3 (N98, N95, N78, N73);
nor NOR3 (N99, N89, N16, N7);
buf BUF1 (N100, N86);
nor NOR2 (N101, N80, N80);
nor NOR4 (N102, N70, N46, N83, N57);
or OR2 (N103, N94, N64);
and AND3 (N104, N102, N73, N1);
xor XOR2 (N105, N93, N101);
buf BUF1 (N106, N67);
buf BUF1 (N107, N98);
not NOT1 (N108, N97);
nor NOR2 (N109, N107, N3);
xor XOR2 (N110, N99, N86);
xor XOR2 (N111, N109, N86);
nand NAND3 (N112, N106, N97, N5);
nand NAND4 (N113, N110, N39, N112, N11);
nand NAND2 (N114, N109, N36);
buf BUF1 (N115, N100);
not NOT1 (N116, N104);
buf BUF1 (N117, N116);
nor NOR3 (N118, N111, N113, N57);
buf BUF1 (N119, N3);
and AND3 (N120, N103, N7, N36);
nand NAND4 (N121, N117, N43, N106, N56);
not NOT1 (N122, N91);
nor NOR3 (N123, N118, N26, N114);
nand NAND4 (N124, N35, N29, N68, N1);
not NOT1 (N125, N108);
nand NAND2 (N126, N96, N88);
nand NAND4 (N127, N126, N41, N29, N29);
and AND4 (N128, N123, N66, N72, N2);
xor XOR2 (N129, N105, N78);
xor XOR2 (N130, N129, N117);
not NOT1 (N131, N124);
nor NOR3 (N132, N128, N48, N54);
or OR4 (N133, N125, N107, N128, N97);
buf BUF1 (N134, N115);
or OR4 (N135, N122, N94, N91, N9);
xor XOR2 (N136, N130, N1);
not NOT1 (N137, N135);
nand NAND2 (N138, N133, N41);
and AND2 (N139, N131, N124);
and AND3 (N140, N120, N30, N17);
nand NAND4 (N141, N119, N67, N85, N39);
nor NOR3 (N142, N140, N93, N99);
nor NOR2 (N143, N139, N127);
and AND4 (N144, N44, N27, N107, N59);
and AND3 (N145, N138, N25, N84);
nor NOR2 (N146, N121, N111);
xor XOR2 (N147, N132, N35);
xor XOR2 (N148, N144, N106);
or OR4 (N149, N134, N96, N108, N74);
nand NAND3 (N150, N143, N129, N141);
buf BUF1 (N151, N149);
and AND3 (N152, N131, N93, N78);
not NOT1 (N153, N150);
nand NAND4 (N154, N148, N89, N31, N105);
nand NAND4 (N155, N153, N38, N61, N117);
xor XOR2 (N156, N146, N9);
xor XOR2 (N157, N145, N56);
buf BUF1 (N158, N155);
and AND3 (N159, N156, N78, N110);
nand NAND3 (N160, N136, N32, N16);
nor NOR2 (N161, N152, N130);
nand NAND2 (N162, N157, N30);
xor XOR2 (N163, N161, N34);
nand NAND2 (N164, N162, N45);
buf BUF1 (N165, N160);
and AND4 (N166, N147, N164, N115, N52);
nand NAND3 (N167, N37, N19, N99);
nor NOR3 (N168, N165, N130, N30);
nor NOR3 (N169, N168, N32, N160);
xor XOR2 (N170, N169, N133);
not NOT1 (N171, N151);
nand NAND3 (N172, N142, N85, N97);
buf BUF1 (N173, N159);
xor XOR2 (N174, N173, N77);
or OR3 (N175, N154, N21, N173);
and AND4 (N176, N174, N89, N116, N96);
buf BUF1 (N177, N163);
nand NAND4 (N178, N175, N158, N165, N24);
buf BUF1 (N179, N98);
or OR3 (N180, N171, N37, N28);
xor XOR2 (N181, N166, N75);
and AND4 (N182, N179, N118, N83, N136);
nor NOR3 (N183, N177, N162, N48);
buf BUF1 (N184, N181);
or OR2 (N185, N182, N128);
buf BUF1 (N186, N180);
or OR3 (N187, N184, N135, N74);
buf BUF1 (N188, N137);
nor NOR4 (N189, N178, N115, N140, N46);
or OR3 (N190, N187, N15, N179);
xor XOR2 (N191, N188, N43);
buf BUF1 (N192, N189);
or OR3 (N193, N185, N167, N190);
not NOT1 (N194, N189);
xor XOR2 (N195, N35, N122);
xor XOR2 (N196, N194, N92);
or OR3 (N197, N172, N181, N82);
buf BUF1 (N198, N193);
or OR4 (N199, N198, N145, N5, N106);
nor NOR2 (N200, N186, N131);
nand NAND2 (N201, N170, N200);
or OR4 (N202, N83, N97, N46, N166);
or OR4 (N203, N191, N64, N171, N39);
xor XOR2 (N204, N202, N186);
nor NOR2 (N205, N196, N200);
and AND3 (N206, N176, N39, N152);
nor NOR2 (N207, N201, N147);
nand NAND4 (N208, N195, N56, N206, N13);
nor NOR2 (N209, N151, N114);
nor NOR2 (N210, N209, N106);
and AND4 (N211, N199, N195, N151, N14);
or OR3 (N212, N211, N34, N135);
and AND2 (N213, N210, N75);
and AND4 (N214, N207, N42, N20, N202);
nand NAND3 (N215, N212, N212, N151);
not NOT1 (N216, N192);
xor XOR2 (N217, N204, N163);
and AND2 (N218, N214, N138);
nand NAND4 (N219, N218, N141, N8, N26);
buf BUF1 (N220, N216);
or OR4 (N221, N203, N23, N86, N135);
buf BUF1 (N222, N221);
buf BUF1 (N223, N222);
not NOT1 (N224, N220);
nor NOR3 (N225, N205, N179, N187);
nand NAND4 (N226, N215, N153, N189, N197);
buf BUF1 (N227, N157);
and AND4 (N228, N224, N180, N183, N206);
nor NOR2 (N229, N51, N82);
not NOT1 (N230, N223);
xor XOR2 (N231, N213, N36);
nor NOR3 (N232, N219, N141, N9);
and AND3 (N233, N230, N133, N63);
nand NAND2 (N234, N226, N33);
nor NOR2 (N235, N228, N31);
not NOT1 (N236, N229);
nor NOR4 (N237, N233, N85, N118, N218);
nor NOR2 (N238, N217, N59);
and AND4 (N239, N234, N68, N160, N22);
nor NOR2 (N240, N235, N42);
xor XOR2 (N241, N231, N170);
buf BUF1 (N242, N227);
buf BUF1 (N243, N241);
nand NAND2 (N244, N239, N142);
nand NAND2 (N245, N244, N22);
not NOT1 (N246, N243);
or OR4 (N247, N225, N16, N84, N128);
nor NOR2 (N248, N245, N189);
buf BUF1 (N249, N236);
nor NOR3 (N250, N247, N242, N91);
not NOT1 (N251, N106);
not NOT1 (N252, N237);
nand NAND2 (N253, N238, N43);
and AND2 (N254, N248, N249);
buf BUF1 (N255, N159);
nor NOR4 (N256, N246, N120, N196, N132);
and AND2 (N257, N240, N202);
buf BUF1 (N258, N256);
not NOT1 (N259, N253);
and AND3 (N260, N254, N230, N136);
nor NOR3 (N261, N252, N132, N86);
xor XOR2 (N262, N251, N203);
not NOT1 (N263, N260);
xor XOR2 (N264, N208, N38);
nor NOR2 (N265, N259, N179);
not NOT1 (N266, N261);
buf BUF1 (N267, N258);
xor XOR2 (N268, N257, N265);
or OR2 (N269, N158, N69);
buf BUF1 (N270, N262);
not NOT1 (N271, N270);
xor XOR2 (N272, N269, N65);
and AND4 (N273, N272, N87, N89, N20);
nor NOR2 (N274, N263, N19);
xor XOR2 (N275, N271, N124);
xor XOR2 (N276, N273, N44);
buf BUF1 (N277, N250);
nand NAND3 (N278, N268, N188, N216);
buf BUF1 (N279, N275);
nor NOR3 (N280, N277, N246, N86);
or OR3 (N281, N266, N69, N17);
nor NOR4 (N282, N232, N50, N70, N134);
or OR4 (N283, N280, N2, N6, N56);
nand NAND2 (N284, N278, N274);
buf BUF1 (N285, N58);
and AND4 (N286, N284, N183, N7, N99);
nand NAND3 (N287, N255, N271, N175);
not NOT1 (N288, N267);
buf BUF1 (N289, N283);
or OR4 (N290, N286, N67, N289, N160);
not NOT1 (N291, N25);
not NOT1 (N292, N290);
or OR3 (N293, N291, N186, N198);
nand NAND4 (N294, N285, N223, N101, N82);
xor XOR2 (N295, N287, N268);
nand NAND4 (N296, N281, N154, N132, N35);
not NOT1 (N297, N276);
and AND4 (N298, N282, N90, N84, N192);
and AND3 (N299, N294, N9, N291);
and AND3 (N300, N288, N93, N267);
nor NOR4 (N301, N295, N61, N210, N176);
nand NAND3 (N302, N279, N48, N126);
buf BUF1 (N303, N300);
and AND2 (N304, N299, N61);
nand NAND3 (N305, N296, N227, N203);
nand NAND4 (N306, N297, N142, N32, N295);
and AND4 (N307, N298, N227, N71, N181);
not NOT1 (N308, N302);
not NOT1 (N309, N292);
nand NAND2 (N310, N304, N278);
not NOT1 (N311, N306);
and AND4 (N312, N264, N141, N252, N308);
or OR3 (N313, N189, N235, N49);
nand NAND3 (N314, N293, N198, N241);
buf BUF1 (N315, N314);
not NOT1 (N316, N310);
and AND2 (N317, N309, N127);
buf BUF1 (N318, N315);
nand NAND4 (N319, N316, N191, N71, N33);
and AND3 (N320, N305, N209, N160);
and AND2 (N321, N313, N107);
xor XOR2 (N322, N318, N266);
nand NAND2 (N323, N312, N27);
xor XOR2 (N324, N303, N274);
nor NOR3 (N325, N324, N81, N148);
or OR4 (N326, N322, N298, N119, N97);
not NOT1 (N327, N319);
nand NAND4 (N328, N320, N210, N245, N295);
xor XOR2 (N329, N307, N30);
xor XOR2 (N330, N311, N329);
and AND3 (N331, N146, N37, N285);
or OR3 (N332, N317, N21, N207);
or OR4 (N333, N325, N43, N176, N188);
or OR4 (N334, N326, N82, N242, N252);
and AND3 (N335, N331, N242, N225);
nand NAND3 (N336, N332, N164, N134);
and AND3 (N337, N334, N140, N189);
and AND2 (N338, N301, N15);
nand NAND4 (N339, N330, N169, N314, N321);
nor NOR2 (N340, N190, N155);
buf BUF1 (N341, N333);
buf BUF1 (N342, N336);
buf BUF1 (N343, N323);
not NOT1 (N344, N340);
nor NOR2 (N345, N344, N7);
xor XOR2 (N346, N343, N102);
xor XOR2 (N347, N335, N196);
nand NAND2 (N348, N341, N220);
nor NOR4 (N349, N342, N151, N8, N291);
buf BUF1 (N350, N327);
nor NOR2 (N351, N328, N101);
nand NAND3 (N352, N346, N249, N315);
xor XOR2 (N353, N348, N285);
xor XOR2 (N354, N352, N234);
not NOT1 (N355, N338);
xor XOR2 (N356, N347, N157);
nor NOR3 (N357, N345, N311, N230);
not NOT1 (N358, N351);
xor XOR2 (N359, N357, N184);
or OR3 (N360, N353, N262, N19);
not NOT1 (N361, N356);
and AND2 (N362, N349, N212);
and AND4 (N363, N362, N176, N123, N330);
nand NAND3 (N364, N358, N71, N350);
nand NAND2 (N365, N283, N222);
buf BUF1 (N366, N354);
or OR4 (N367, N337, N208, N7, N362);
nand NAND4 (N368, N367, N246, N128, N88);
nor NOR2 (N369, N355, N312);
nor NOR3 (N370, N364, N253, N89);
buf BUF1 (N371, N339);
not NOT1 (N372, N366);
nand NAND4 (N373, N363, N26, N13, N271);
xor XOR2 (N374, N370, N54);
not NOT1 (N375, N374);
or OR3 (N376, N369, N121, N209);
and AND4 (N377, N371, N186, N296, N358);
nand NAND2 (N378, N368, N207);
and AND2 (N379, N365, N154);
xor XOR2 (N380, N372, N322);
or OR4 (N381, N378, N83, N21, N260);
or OR4 (N382, N359, N94, N34, N346);
nor NOR2 (N383, N360, N189);
not NOT1 (N384, N377);
nand NAND2 (N385, N384, N3);
nor NOR4 (N386, N361, N343, N301, N27);
or OR2 (N387, N386, N89);
or OR3 (N388, N383, N243, N336);
nand NAND4 (N389, N379, N230, N359, N123);
nand NAND2 (N390, N375, N24);
not NOT1 (N391, N382);
xor XOR2 (N392, N381, N114);
xor XOR2 (N393, N380, N183);
not NOT1 (N394, N390);
buf BUF1 (N395, N392);
nor NOR3 (N396, N387, N312, N165);
or OR4 (N397, N376, N62, N377, N63);
and AND2 (N398, N385, N52);
xor XOR2 (N399, N393, N220);
and AND4 (N400, N397, N346, N17, N229);
nor NOR2 (N401, N399, N282);
or OR4 (N402, N396, N57, N364, N350);
nor NOR3 (N403, N394, N136, N154);
buf BUF1 (N404, N398);
and AND2 (N405, N401, N270);
nand NAND4 (N406, N404, N152, N158, N95);
not NOT1 (N407, N400);
nand NAND3 (N408, N406, N48, N347);
xor XOR2 (N409, N402, N29);
not NOT1 (N410, N388);
not NOT1 (N411, N403);
xor XOR2 (N412, N409, N207);
buf BUF1 (N413, N389);
nand NAND2 (N414, N410, N53);
xor XOR2 (N415, N373, N78);
or OR4 (N416, N413, N157, N26, N200);
buf BUF1 (N417, N405);
nor NOR2 (N418, N416, N181);
nand NAND4 (N419, N408, N387, N308, N237);
xor XOR2 (N420, N407, N337);
nand NAND2 (N421, N419, N144);
nor NOR4 (N422, N412, N372, N192, N180);
and AND3 (N423, N422, N205, N89);
nor NOR3 (N424, N415, N208, N117);
and AND4 (N425, N391, N302, N239, N339);
buf BUF1 (N426, N423);
and AND4 (N427, N425, N6, N75, N234);
nand NAND3 (N428, N424, N335, N208);
nor NOR4 (N429, N417, N153, N231, N381);
xor XOR2 (N430, N395, N357);
not NOT1 (N431, N426);
nand NAND2 (N432, N430, N45);
nand NAND4 (N433, N411, N121, N255, N367);
xor XOR2 (N434, N428, N149);
buf BUF1 (N435, N434);
nor NOR3 (N436, N420, N392, N326);
or OR2 (N437, N427, N63);
and AND4 (N438, N421, N423, N41, N268);
nand NAND2 (N439, N429, N415);
nor NOR2 (N440, N438, N60);
nand NAND3 (N441, N414, N391, N316);
or OR4 (N442, N431, N120, N101, N362);
nor NOR3 (N443, N440, N232, N10);
or OR2 (N444, N439, N408);
nor NOR3 (N445, N418, N422, N128);
buf BUF1 (N446, N441);
not NOT1 (N447, N436);
nor NOR4 (N448, N447, N74, N100, N338);
and AND4 (N449, N443, N104, N223, N362);
nand NAND3 (N450, N444, N11, N428);
xor XOR2 (N451, N445, N318);
not NOT1 (N452, N448);
or OR3 (N453, N451, N214, N192);
nand NAND4 (N454, N446, N154, N323, N141);
and AND3 (N455, N433, N331, N240);
xor XOR2 (N456, N450, N445);
and AND4 (N457, N435, N258, N316, N332);
nand NAND2 (N458, N452, N415);
nor NOR2 (N459, N453, N139);
and AND4 (N460, N432, N345, N414, N291);
nor NOR2 (N461, N455, N399);
or OR4 (N462, N437, N67, N300, N397);
and AND4 (N463, N458, N170, N38, N102);
nor NOR4 (N464, N460, N57, N23, N138);
xor XOR2 (N465, N461, N373);
xor XOR2 (N466, N464, N9);
nor NOR4 (N467, N449, N209, N425, N294);
and AND2 (N468, N467, N353);
nand NAND2 (N469, N442, N35);
xor XOR2 (N470, N456, N78);
nor NOR3 (N471, N454, N389, N433);
or OR3 (N472, N471, N420, N240);
nor NOR4 (N473, N470, N228, N203, N18);
not NOT1 (N474, N466);
not NOT1 (N475, N457);
not NOT1 (N476, N463);
or OR4 (N477, N462, N182, N373, N474);
and AND4 (N478, N284, N390, N8, N91);
nor NOR4 (N479, N475, N348, N40, N299);
nand NAND2 (N480, N459, N364);
buf BUF1 (N481, N472);
or OR3 (N482, N479, N17, N276);
xor XOR2 (N483, N477, N158);
nand NAND4 (N484, N469, N81, N403, N370);
not NOT1 (N485, N480);
not NOT1 (N486, N476);
and AND2 (N487, N481, N228);
buf BUF1 (N488, N478);
or OR4 (N489, N482, N244, N452, N78);
nor NOR4 (N490, N488, N407, N49, N271);
nor NOR4 (N491, N490, N335, N283, N141);
not NOT1 (N492, N468);
or OR2 (N493, N487, N106);
not NOT1 (N494, N492);
or OR2 (N495, N489, N210);
or OR4 (N496, N483, N356, N494, N187);
nor NOR2 (N497, N439, N431);
and AND2 (N498, N497, N158);
or OR3 (N499, N485, N222, N280);
buf BUF1 (N500, N496);
buf BUF1 (N501, N486);
buf BUF1 (N502, N495);
or OR3 (N503, N493, N288, N44);
not NOT1 (N504, N503);
xor XOR2 (N505, N499, N7);
or OR3 (N506, N505, N299, N159);
or OR2 (N507, N498, N439);
not NOT1 (N508, N507);
not NOT1 (N509, N504);
xor XOR2 (N510, N502, N41);
nand NAND3 (N511, N465, N400, N264);
not NOT1 (N512, N501);
nand NAND3 (N513, N511, N280, N257);
and AND3 (N514, N513, N167, N47);
nor NOR3 (N515, N514, N124, N192);
not NOT1 (N516, N500);
and AND4 (N517, N512, N176, N325, N448);
or OR2 (N518, N517, N147);
not NOT1 (N519, N516);
nor NOR3 (N520, N473, N207, N477);
nand NAND4 (N521, N518, N271, N87, N393);
nand NAND3 (N522, N509, N456, N448);
or OR4 (N523, N506, N407, N400, N278);
and AND4 (N524, N508, N261, N140, N240);
or OR3 (N525, N510, N421, N236);
buf BUF1 (N526, N515);
not NOT1 (N527, N521);
nor NOR4 (N528, N523, N438, N156, N258);
buf BUF1 (N529, N484);
nor NOR2 (N530, N529, N159);
nor NOR4 (N531, N520, N191, N266, N161);
buf BUF1 (N532, N522);
nor NOR3 (N533, N491, N113, N237);
nor NOR4 (N534, N527, N192, N170, N120);
buf BUF1 (N535, N534);
nand NAND3 (N536, N535, N227, N329);
buf BUF1 (N537, N528);
buf BUF1 (N538, N531);
nor NOR4 (N539, N537, N271, N510, N111);
or OR3 (N540, N525, N411, N268);
and AND4 (N541, N539, N34, N108, N167);
buf BUF1 (N542, N526);
and AND2 (N543, N530, N196);
xor XOR2 (N544, N519, N52);
xor XOR2 (N545, N538, N78);
buf BUF1 (N546, N533);
nand NAND4 (N547, N545, N488, N329, N148);
and AND2 (N548, N546, N258);
xor XOR2 (N549, N524, N334);
xor XOR2 (N550, N542, N397);
nand NAND4 (N551, N544, N203, N80, N506);
nor NOR3 (N552, N543, N253, N218);
and AND3 (N553, N552, N398, N477);
and AND3 (N554, N532, N106, N442);
buf BUF1 (N555, N549);
or OR3 (N556, N555, N379, N496);
nor NOR3 (N557, N551, N118, N316);
and AND4 (N558, N540, N485, N484, N172);
or OR4 (N559, N548, N423, N337, N377);
not NOT1 (N560, N554);
nand NAND2 (N561, N557, N440);
buf BUF1 (N562, N556);
buf BUF1 (N563, N547);
or OR3 (N564, N541, N130, N497);
nor NOR2 (N565, N536, N346);
nor NOR2 (N566, N559, N428);
nor NOR4 (N567, N565, N214, N459, N46);
not NOT1 (N568, N560);
xor XOR2 (N569, N550, N292);
xor XOR2 (N570, N553, N277);
nor NOR3 (N571, N562, N531, N250);
and AND2 (N572, N561, N265);
nor NOR3 (N573, N564, N75, N289);
nor NOR2 (N574, N572, N456);
not NOT1 (N575, N558);
not NOT1 (N576, N569);
xor XOR2 (N577, N563, N538);
nand NAND3 (N578, N576, N267, N446);
nor NOR3 (N579, N567, N550, N426);
buf BUF1 (N580, N571);
nor NOR3 (N581, N574, N347, N103);
buf BUF1 (N582, N579);
nand NAND2 (N583, N573, N212);
nor NOR2 (N584, N580, N406);
and AND2 (N585, N581, N88);
nand NAND4 (N586, N584, N476, N345, N405);
and AND2 (N587, N583, N348);
and AND3 (N588, N582, N392, N199);
nor NOR4 (N589, N570, N45, N487, N509);
and AND4 (N590, N578, N375, N468, N302);
or OR2 (N591, N587, N345);
and AND3 (N592, N591, N466, N207);
xor XOR2 (N593, N590, N399);
xor XOR2 (N594, N585, N109);
xor XOR2 (N595, N592, N363);
and AND2 (N596, N586, N264);
buf BUF1 (N597, N566);
nor NOR3 (N598, N568, N86, N135);
xor XOR2 (N599, N596, N316);
not NOT1 (N600, N595);
or OR2 (N601, N588, N414);
nor NOR2 (N602, N601, N479);
and AND2 (N603, N594, N325);
and AND3 (N604, N598, N543, N240);
buf BUF1 (N605, N593);
and AND4 (N606, N605, N530, N192, N204);
and AND2 (N607, N603, N37);
buf BUF1 (N608, N577);
nand NAND4 (N609, N589, N401, N37, N243);
nor NOR4 (N610, N575, N479, N436, N206);
buf BUF1 (N611, N609);
nor NOR2 (N612, N602, N365);
not NOT1 (N613, N608);
and AND2 (N614, N611, N445);
and AND2 (N615, N614, N248);
not NOT1 (N616, N599);
buf BUF1 (N617, N615);
buf BUF1 (N618, N610);
nor NOR3 (N619, N617, N15, N324);
nor NOR4 (N620, N613, N24, N430, N585);
and AND2 (N621, N616, N352);
nand NAND4 (N622, N604, N338, N154, N80);
nor NOR3 (N623, N607, N506, N385);
xor XOR2 (N624, N612, N101);
or OR2 (N625, N597, N96);
and AND4 (N626, N606, N558, N97, N346);
nand NAND2 (N627, N623, N94);
nand NAND4 (N628, N626, N286, N434, N239);
not NOT1 (N629, N621);
or OR3 (N630, N624, N109, N344);
xor XOR2 (N631, N628, N520);
or OR3 (N632, N620, N384, N239);
buf BUF1 (N633, N627);
or OR2 (N634, N633, N319);
or OR4 (N635, N630, N522, N337, N252);
not NOT1 (N636, N625);
not NOT1 (N637, N631);
not NOT1 (N638, N629);
buf BUF1 (N639, N636);
or OR3 (N640, N632, N404, N42);
nor NOR2 (N641, N637, N126);
nand NAND3 (N642, N638, N74, N42);
nor NOR3 (N643, N642, N224, N548);
nand NAND3 (N644, N634, N212, N568);
xor XOR2 (N645, N639, N521);
xor XOR2 (N646, N641, N39);
xor XOR2 (N647, N619, N551);
nor NOR4 (N648, N645, N151, N335, N512);
nand NAND4 (N649, N646, N202, N525, N334);
and AND3 (N650, N618, N582, N135);
and AND4 (N651, N649, N285, N403, N505);
and AND4 (N652, N650, N94, N285, N635);
buf BUF1 (N653, N26);
xor XOR2 (N654, N647, N227);
not NOT1 (N655, N643);
or OR4 (N656, N654, N213, N279, N549);
or OR4 (N657, N622, N516, N207, N280);
xor XOR2 (N658, N640, N309);
nor NOR3 (N659, N651, N83, N344);
not NOT1 (N660, N653);
or OR3 (N661, N600, N276, N511);
nor NOR2 (N662, N652, N48);
or OR2 (N663, N659, N531);
and AND2 (N664, N644, N94);
nand NAND2 (N665, N658, N265);
nand NAND4 (N666, N662, N299, N304, N78);
and AND4 (N667, N664, N477, N441, N574);
and AND2 (N668, N665, N644);
and AND4 (N669, N648, N403, N205, N530);
and AND3 (N670, N661, N340, N60);
or OR3 (N671, N667, N278, N472);
xor XOR2 (N672, N655, N405);
xor XOR2 (N673, N669, N256);
buf BUF1 (N674, N672);
not NOT1 (N675, N660);
xor XOR2 (N676, N671, N120);
not NOT1 (N677, N674);
or OR2 (N678, N663, N634);
nor NOR4 (N679, N668, N510, N253, N147);
and AND4 (N680, N666, N564, N404, N190);
and AND3 (N681, N677, N92, N535);
nor NOR3 (N682, N676, N179, N462);
not NOT1 (N683, N673);
or OR3 (N684, N656, N210, N658);
nor NOR4 (N685, N680, N83, N513, N185);
nand NAND3 (N686, N657, N546, N237);
nor NOR2 (N687, N686, N238);
buf BUF1 (N688, N670);
and AND3 (N689, N684, N527, N522);
buf BUF1 (N690, N685);
nor NOR3 (N691, N678, N215, N85);
nand NAND3 (N692, N682, N511, N54);
not NOT1 (N693, N691);
xor XOR2 (N694, N693, N204);
buf BUF1 (N695, N675);
not NOT1 (N696, N695);
nand NAND4 (N697, N689, N501, N484, N149);
nand NAND3 (N698, N679, N380, N692);
nand NAND2 (N699, N644, N347);
buf BUF1 (N700, N690);
buf BUF1 (N701, N683);
not NOT1 (N702, N699);
and AND3 (N703, N688, N563, N256);
and AND4 (N704, N702, N396, N619, N174);
and AND3 (N705, N704, N388, N383);
nand NAND2 (N706, N705, N118);
not NOT1 (N707, N697);
and AND4 (N708, N703, N145, N156, N636);
buf BUF1 (N709, N700);
not NOT1 (N710, N696);
or OR4 (N711, N681, N170, N322, N128);
buf BUF1 (N712, N710);
buf BUF1 (N713, N698);
nor NOR4 (N714, N707, N613, N14, N433);
and AND3 (N715, N713, N647, N547);
buf BUF1 (N716, N715);
not NOT1 (N717, N687);
or OR4 (N718, N706, N70, N31, N109);
not NOT1 (N719, N717);
nor NOR3 (N720, N712, N532, N569);
or OR4 (N721, N711, N672, N192, N96);
xor XOR2 (N722, N714, N193);
nor NOR3 (N723, N701, N525, N206);
and AND3 (N724, N708, N3, N61);
buf BUF1 (N725, N720);
xor XOR2 (N726, N723, N546);
xor XOR2 (N727, N721, N271);
and AND4 (N728, N727, N157, N29, N403);
not NOT1 (N729, N709);
xor XOR2 (N730, N728, N183);
nand NAND3 (N731, N694, N335, N646);
or OR4 (N732, N729, N669, N271, N492);
nand NAND4 (N733, N725, N420, N554, N360);
nor NOR2 (N734, N718, N201);
not NOT1 (N735, N733);
buf BUF1 (N736, N724);
xor XOR2 (N737, N722, N106);
nor NOR4 (N738, N734, N304, N414, N710);
nand NAND2 (N739, N716, N157);
buf BUF1 (N740, N726);
not NOT1 (N741, N735);
xor XOR2 (N742, N738, N451);
not NOT1 (N743, N719);
or OR4 (N744, N742, N98, N38, N311);
and AND3 (N745, N737, N246, N657);
and AND4 (N746, N740, N658, N652, N569);
xor XOR2 (N747, N731, N444);
nor NOR2 (N748, N745, N580);
and AND3 (N749, N741, N215, N543);
or OR3 (N750, N748, N573, N350);
buf BUF1 (N751, N743);
xor XOR2 (N752, N730, N66);
nor NOR3 (N753, N744, N311, N428);
xor XOR2 (N754, N750, N317);
not NOT1 (N755, N751);
nand NAND4 (N756, N739, N745, N42, N242);
buf BUF1 (N757, N752);
and AND4 (N758, N749, N621, N296, N104);
nor NOR3 (N759, N758, N556, N728);
xor XOR2 (N760, N736, N20);
and AND3 (N761, N747, N685, N540);
xor XOR2 (N762, N761, N596);
not NOT1 (N763, N754);
xor XOR2 (N764, N760, N633);
or OR4 (N765, N755, N447, N187, N2);
nand NAND3 (N766, N757, N547, N270);
buf BUF1 (N767, N766);
not NOT1 (N768, N732);
nand NAND2 (N769, N759, N410);
not NOT1 (N770, N767);
and AND2 (N771, N769, N281);
nand NAND4 (N772, N753, N298, N543, N349);
nor NOR3 (N773, N764, N147, N129);
buf BUF1 (N774, N765);
or OR3 (N775, N770, N387, N453);
buf BUF1 (N776, N746);
buf BUF1 (N777, N775);
nor NOR4 (N778, N756, N175, N84, N698);
or OR3 (N779, N771, N667, N582);
nor NOR3 (N780, N776, N396, N166);
nand NAND3 (N781, N777, N516, N604);
buf BUF1 (N782, N763);
buf BUF1 (N783, N778);
xor XOR2 (N784, N762, N749);
or OR4 (N785, N784, N366, N562, N519);
or OR4 (N786, N768, N436, N742, N179);
xor XOR2 (N787, N780, N616);
buf BUF1 (N788, N786);
or OR2 (N789, N788, N214);
xor XOR2 (N790, N781, N240);
and AND4 (N791, N773, N756, N671, N558);
nand NAND2 (N792, N785, N516);
nor NOR4 (N793, N774, N267, N355, N766);
nor NOR4 (N794, N791, N540, N640, N48);
buf BUF1 (N795, N793);
or OR2 (N796, N790, N567);
or OR4 (N797, N796, N109, N370, N356);
buf BUF1 (N798, N794);
not NOT1 (N799, N772);
and AND3 (N800, N797, N458, N680);
or OR4 (N801, N792, N8, N494, N577);
nor NOR3 (N802, N783, N354, N247);
and AND2 (N803, N801, N623);
nand NAND4 (N804, N795, N585, N28, N797);
nand NAND2 (N805, N789, N503);
and AND4 (N806, N802, N638, N165, N673);
nand NAND3 (N807, N805, N763, N96);
nor NOR4 (N808, N804, N161, N750, N578);
or OR3 (N809, N807, N492, N59);
and AND2 (N810, N809, N614);
buf BUF1 (N811, N799);
buf BUF1 (N812, N798);
buf BUF1 (N813, N811);
nand NAND4 (N814, N800, N201, N413, N289);
nor NOR2 (N815, N803, N273);
not NOT1 (N816, N813);
not NOT1 (N817, N808);
and AND2 (N818, N779, N582);
not NOT1 (N819, N782);
not NOT1 (N820, N787);
not NOT1 (N821, N819);
and AND2 (N822, N821, N640);
xor XOR2 (N823, N822, N235);
nor NOR2 (N824, N806, N400);
xor XOR2 (N825, N815, N560);
nor NOR3 (N826, N825, N761, N11);
nor NOR4 (N827, N818, N131, N778, N491);
not NOT1 (N828, N812);
nand NAND3 (N829, N823, N735, N271);
xor XOR2 (N830, N820, N526);
xor XOR2 (N831, N810, N162);
not NOT1 (N832, N828);
xor XOR2 (N833, N824, N770);
nand NAND2 (N834, N814, N686);
and AND2 (N835, N834, N273);
or OR4 (N836, N831, N142, N763, N697);
nand NAND4 (N837, N829, N550, N748, N64);
nand NAND2 (N838, N816, N490);
nand NAND4 (N839, N832, N26, N81, N335);
and AND2 (N840, N839, N364);
nand NAND2 (N841, N837, N692);
or OR4 (N842, N840, N67, N458, N539);
nor NOR2 (N843, N836, N551);
buf BUF1 (N844, N835);
buf BUF1 (N845, N844);
buf BUF1 (N846, N826);
not NOT1 (N847, N846);
nand NAND3 (N848, N843, N680, N151);
xor XOR2 (N849, N848, N690);
not NOT1 (N850, N833);
xor XOR2 (N851, N841, N505);
and AND2 (N852, N845, N119);
nor NOR3 (N853, N838, N564, N655);
and AND3 (N854, N827, N352, N423);
and AND4 (N855, N830, N86, N92, N580);
xor XOR2 (N856, N849, N684);
or OR2 (N857, N852, N137);
not NOT1 (N858, N857);
and AND2 (N859, N851, N121);
nor NOR4 (N860, N850, N489, N154, N483);
not NOT1 (N861, N855);
nand NAND2 (N862, N853, N22);
not NOT1 (N863, N861);
not NOT1 (N864, N847);
xor XOR2 (N865, N859, N733);
nand NAND3 (N866, N862, N475, N362);
or OR3 (N867, N842, N150, N635);
buf BUF1 (N868, N860);
or OR2 (N869, N854, N243);
nand NAND2 (N870, N865, N280);
buf BUF1 (N871, N864);
or OR4 (N872, N868, N602, N517, N225);
buf BUF1 (N873, N867);
xor XOR2 (N874, N817, N774);
buf BUF1 (N875, N869);
or OR2 (N876, N863, N771);
nor NOR3 (N877, N858, N189, N246);
not NOT1 (N878, N876);
or OR3 (N879, N872, N628, N709);
and AND4 (N880, N874, N376, N814, N244);
xor XOR2 (N881, N878, N824);
xor XOR2 (N882, N877, N375);
or OR3 (N883, N881, N696, N537);
and AND3 (N884, N880, N53, N146);
or OR3 (N885, N866, N661, N551);
nand NAND3 (N886, N882, N103, N66);
nor NOR2 (N887, N885, N151);
xor XOR2 (N888, N875, N819);
or OR2 (N889, N873, N858);
or OR3 (N890, N883, N556, N325);
and AND3 (N891, N871, N348, N521);
not NOT1 (N892, N889);
buf BUF1 (N893, N884);
not NOT1 (N894, N891);
buf BUF1 (N895, N893);
nand NAND2 (N896, N890, N571);
or OR2 (N897, N870, N169);
nor NOR4 (N898, N879, N654, N763, N559);
and AND2 (N899, N896, N196);
or OR2 (N900, N898, N340);
xor XOR2 (N901, N897, N747);
buf BUF1 (N902, N900);
and AND3 (N903, N886, N629, N240);
not NOT1 (N904, N888);
nand NAND3 (N905, N899, N739, N92);
nand NAND4 (N906, N856, N5, N206, N160);
xor XOR2 (N907, N892, N238);
not NOT1 (N908, N905);
nor NOR4 (N909, N895, N103, N129, N836);
and AND4 (N910, N906, N179, N20, N664);
or OR2 (N911, N909, N652);
and AND4 (N912, N910, N284, N177, N843);
and AND3 (N913, N911, N190, N480);
nor NOR3 (N914, N887, N878, N109);
and AND3 (N915, N894, N197, N588);
not NOT1 (N916, N912);
buf BUF1 (N917, N915);
nor NOR3 (N918, N917, N292, N708);
buf BUF1 (N919, N901);
nand NAND2 (N920, N902, N399);
xor XOR2 (N921, N919, N486);
not NOT1 (N922, N920);
not NOT1 (N923, N922);
and AND3 (N924, N923, N246, N313);
nor NOR2 (N925, N916, N696);
or OR3 (N926, N913, N924, N162);
and AND4 (N927, N466, N499, N762, N625);
and AND3 (N928, N907, N342, N681);
xor XOR2 (N929, N925, N346);
buf BUF1 (N930, N903);
and AND2 (N931, N904, N667);
nand NAND4 (N932, N931, N689, N589, N645);
and AND2 (N933, N918, N162);
and AND2 (N934, N914, N741);
nand NAND2 (N935, N927, N386);
nand NAND3 (N936, N934, N31, N625);
or OR3 (N937, N926, N609, N763);
buf BUF1 (N938, N932);
and AND4 (N939, N933, N728, N858, N883);
not NOT1 (N940, N936);
nor NOR4 (N941, N940, N21, N47, N106);
buf BUF1 (N942, N921);
and AND2 (N943, N930, N662);
nor NOR4 (N944, N939, N559, N29, N874);
buf BUF1 (N945, N943);
and AND2 (N946, N928, N845);
xor XOR2 (N947, N937, N177);
xor XOR2 (N948, N941, N430);
xor XOR2 (N949, N947, N324);
nor NOR2 (N950, N935, N18);
nor NOR2 (N951, N938, N607);
nand NAND3 (N952, N908, N33, N536);
and AND2 (N953, N946, N881);
nand NAND3 (N954, N951, N822, N310);
xor XOR2 (N955, N952, N935);
or OR4 (N956, N945, N587, N188, N286);
buf BUF1 (N957, N942);
nor NOR3 (N958, N929, N533, N612);
and AND4 (N959, N954, N691, N137, N62);
not NOT1 (N960, N950);
or OR3 (N961, N955, N676, N505);
not NOT1 (N962, N948);
not NOT1 (N963, N957);
nor NOR4 (N964, N963, N501, N171, N85);
and AND2 (N965, N958, N488);
buf BUF1 (N966, N964);
nand NAND4 (N967, N956, N345, N36, N91);
or OR4 (N968, N960, N734, N732, N494);
and AND4 (N969, N967, N368, N9, N573);
buf BUF1 (N970, N961);
and AND4 (N971, N965, N356, N325, N920);
and AND2 (N972, N959, N947);
buf BUF1 (N973, N944);
buf BUF1 (N974, N970);
and AND4 (N975, N968, N974, N351, N10);
nor NOR2 (N976, N3, N68);
not NOT1 (N977, N975);
xor XOR2 (N978, N969, N860);
or OR3 (N979, N977, N946, N834);
nand NAND4 (N980, N979, N671, N459, N752);
nor NOR3 (N981, N980, N146, N663);
nand NAND2 (N982, N962, N445);
nand NAND3 (N983, N972, N892, N950);
nand NAND4 (N984, N983, N765, N725, N252);
or OR3 (N985, N981, N755, N786);
and AND3 (N986, N976, N769, N704);
and AND3 (N987, N978, N676, N510);
not NOT1 (N988, N953);
buf BUF1 (N989, N985);
xor XOR2 (N990, N989, N248);
not NOT1 (N991, N987);
nor NOR2 (N992, N982, N971);
or OR3 (N993, N883, N429, N401);
nand NAND2 (N994, N984, N281);
buf BUF1 (N995, N993);
xor XOR2 (N996, N990, N775);
xor XOR2 (N997, N988, N913);
and AND4 (N998, N997, N946, N471, N316);
buf BUF1 (N999, N996);
buf BUF1 (N1000, N995);
and AND4 (N1001, N994, N1000, N932, N569);
xor XOR2 (N1002, N557, N372);
not NOT1 (N1003, N998);
or OR3 (N1004, N966, N711, N866);
xor XOR2 (N1005, N991, N603);
buf BUF1 (N1006, N973);
nor NOR4 (N1007, N1003, N509, N773, N567);
nor NOR3 (N1008, N1004, N1, N100);
buf BUF1 (N1009, N999);
nor NOR2 (N1010, N1009, N744);
xor XOR2 (N1011, N949, N530);
or OR2 (N1012, N1006, N654);
buf BUF1 (N1013, N1011);
not NOT1 (N1014, N1012);
xor XOR2 (N1015, N1010, N425);
buf BUF1 (N1016, N1014);
buf BUF1 (N1017, N1013);
or OR4 (N1018, N1001, N826, N322, N241);
or OR2 (N1019, N1002, N139);
and AND2 (N1020, N1007, N126);
nand NAND3 (N1021, N1008, N32, N373);
and AND2 (N1022, N1017, N73);
buf BUF1 (N1023, N1020);
or OR3 (N1024, N1023, N740, N574);
xor XOR2 (N1025, N986, N539);
nand NAND2 (N1026, N1016, N760);
and AND2 (N1027, N1019, N1011);
or OR4 (N1028, N1027, N593, N710, N979);
and AND2 (N1029, N1022, N756);
nor NOR4 (N1030, N1028, N787, N286, N616);
nand NAND4 (N1031, N1018, N926, N453, N275);
xor XOR2 (N1032, N1024, N709);
buf BUF1 (N1033, N1005);
buf BUF1 (N1034, N1025);
nand NAND4 (N1035, N1021, N853, N158, N543);
nand NAND2 (N1036, N1033, N722);
or OR3 (N1037, N1029, N792, N954);
nor NOR2 (N1038, N1032, N1028);
or OR4 (N1039, N1030, N704, N750, N696);
nand NAND2 (N1040, N1037, N559);
xor XOR2 (N1041, N1015, N128);
nand NAND3 (N1042, N1031, N500, N273);
and AND4 (N1043, N1040, N298, N682, N426);
or OR2 (N1044, N1042, N231);
or OR3 (N1045, N992, N717, N229);
buf BUF1 (N1046, N1045);
xor XOR2 (N1047, N1026, N234);
buf BUF1 (N1048, N1047);
nand NAND2 (N1049, N1039, N721);
buf BUF1 (N1050, N1038);
nor NOR2 (N1051, N1043, N438);
not NOT1 (N1052, N1051);
and AND4 (N1053, N1035, N10, N760, N887);
and AND3 (N1054, N1053, N244, N541);
nand NAND3 (N1055, N1052, N861, N11);
nor NOR4 (N1056, N1048, N114, N72, N370);
nor NOR4 (N1057, N1041, N716, N862, N152);
buf BUF1 (N1058, N1036);
nor NOR2 (N1059, N1049, N251);
nor NOR3 (N1060, N1054, N23, N778);
xor XOR2 (N1061, N1058, N927);
xor XOR2 (N1062, N1050, N145);
nand NAND3 (N1063, N1061, N844, N340);
nor NOR3 (N1064, N1062, N831, N639);
and AND4 (N1065, N1055, N642, N320, N457);
and AND3 (N1066, N1044, N960, N730);
not NOT1 (N1067, N1057);
xor XOR2 (N1068, N1060, N208);
nor NOR3 (N1069, N1046, N912, N672);
buf BUF1 (N1070, N1059);
nand NAND2 (N1071, N1070, N58);
nor NOR3 (N1072, N1063, N233, N246);
or OR2 (N1073, N1069, N553);
buf BUF1 (N1074, N1072);
xor XOR2 (N1075, N1065, N545);
xor XOR2 (N1076, N1066, N542);
xor XOR2 (N1077, N1074, N615);
nand NAND3 (N1078, N1075, N456, N332);
buf BUF1 (N1079, N1073);
nor NOR4 (N1080, N1077, N385, N397, N241);
xor XOR2 (N1081, N1080, N291);
or OR3 (N1082, N1064, N857, N582);
not NOT1 (N1083, N1068);
and AND2 (N1084, N1056, N784);
not NOT1 (N1085, N1034);
nor NOR2 (N1086, N1085, N635);
buf BUF1 (N1087, N1084);
nor NOR3 (N1088, N1086, N855, N121);
nor NOR2 (N1089, N1083, N310);
or OR3 (N1090, N1071, N225, N728);
nand NAND4 (N1091, N1082, N623, N631, N819);
or OR2 (N1092, N1089, N932);
xor XOR2 (N1093, N1087, N112);
or OR2 (N1094, N1092, N694);
buf BUF1 (N1095, N1090);
and AND2 (N1096, N1067, N701);
nor NOR3 (N1097, N1091, N651, N14);
buf BUF1 (N1098, N1095);
not NOT1 (N1099, N1088);
and AND4 (N1100, N1098, N7, N482, N1043);
and AND3 (N1101, N1078, N896, N615);
nand NAND3 (N1102, N1100, N129, N580);
or OR3 (N1103, N1093, N793, N896);
xor XOR2 (N1104, N1103, N297);
nand NAND4 (N1105, N1096, N39, N106, N127);
or OR2 (N1106, N1094, N790);
not NOT1 (N1107, N1101);
and AND3 (N1108, N1104, N1022, N692);
buf BUF1 (N1109, N1108);
buf BUF1 (N1110, N1109);
not NOT1 (N1111, N1097);
not NOT1 (N1112, N1079);
or OR3 (N1113, N1081, N55, N1065);
not NOT1 (N1114, N1102);
xor XOR2 (N1115, N1113, N77);
and AND2 (N1116, N1111, N858);
nand NAND3 (N1117, N1115, N302, N106);
or OR3 (N1118, N1116, N477, N1043);
xor XOR2 (N1119, N1099, N722);
nand NAND3 (N1120, N1118, N900, N1033);
nor NOR4 (N1121, N1076, N204, N648, N769);
buf BUF1 (N1122, N1121);
xor XOR2 (N1123, N1122, N10);
xor XOR2 (N1124, N1106, N372);
xor XOR2 (N1125, N1119, N448);
nand NAND2 (N1126, N1107, N743);
nor NOR2 (N1127, N1124, N317);
or OR4 (N1128, N1123, N836, N76, N844);
buf BUF1 (N1129, N1127);
buf BUF1 (N1130, N1125);
or OR4 (N1131, N1110, N492, N386, N1075);
xor XOR2 (N1132, N1130, N240);
nand NAND4 (N1133, N1105, N1076, N107, N251);
nor NOR2 (N1134, N1117, N353);
or OR4 (N1135, N1133, N1087, N1088, N948);
xor XOR2 (N1136, N1134, N1033);
or OR4 (N1137, N1129, N977, N822, N921);
not NOT1 (N1138, N1137);
nand NAND3 (N1139, N1128, N246, N225);
buf BUF1 (N1140, N1132);
or OR3 (N1141, N1114, N1127, N769);
buf BUF1 (N1142, N1141);
nor NOR4 (N1143, N1126, N237, N130, N877);
nor NOR3 (N1144, N1112, N401, N809);
nor NOR2 (N1145, N1131, N1015);
or OR3 (N1146, N1120, N216, N826);
not NOT1 (N1147, N1135);
not NOT1 (N1148, N1143);
buf BUF1 (N1149, N1138);
nand NAND3 (N1150, N1146, N425, N500);
xor XOR2 (N1151, N1148, N118);
and AND3 (N1152, N1145, N16, N1034);
nand NAND3 (N1153, N1144, N326, N772);
and AND3 (N1154, N1136, N493, N127);
nand NAND3 (N1155, N1140, N93, N474);
nand NAND3 (N1156, N1151, N734, N130);
nand NAND3 (N1157, N1139, N480, N997);
or OR3 (N1158, N1149, N536, N248);
nand NAND2 (N1159, N1147, N463);
and AND4 (N1160, N1158, N577, N422, N707);
nand NAND2 (N1161, N1150, N414);
buf BUF1 (N1162, N1155);
nand NAND2 (N1163, N1142, N745);
not NOT1 (N1164, N1163);
not NOT1 (N1165, N1157);
xor XOR2 (N1166, N1154, N1030);
not NOT1 (N1167, N1162);
not NOT1 (N1168, N1164);
not NOT1 (N1169, N1168);
not NOT1 (N1170, N1160);
xor XOR2 (N1171, N1153, N873);
nand NAND2 (N1172, N1152, N899);
nor NOR4 (N1173, N1172, N25, N893, N20);
nand NAND3 (N1174, N1161, N288, N410);
nand NAND3 (N1175, N1173, N643, N256);
or OR3 (N1176, N1170, N949, N402);
nand NAND4 (N1177, N1156, N1097, N139, N905);
xor XOR2 (N1178, N1174, N1065);
nand NAND4 (N1179, N1169, N931, N1043, N510);
buf BUF1 (N1180, N1179);
and AND3 (N1181, N1165, N498, N684);
nand NAND4 (N1182, N1181, N28, N162, N245);
nor NOR3 (N1183, N1167, N215, N374);
nor NOR2 (N1184, N1180, N957);
nor NOR4 (N1185, N1166, N246, N30, N954);
buf BUF1 (N1186, N1159);
or OR3 (N1187, N1182, N512, N623);
xor XOR2 (N1188, N1178, N650);
xor XOR2 (N1189, N1171, N365);
or OR4 (N1190, N1187, N451, N261, N768);
or OR3 (N1191, N1185, N49, N694);
or OR2 (N1192, N1186, N1079);
xor XOR2 (N1193, N1175, N203);
nor NOR2 (N1194, N1183, N284);
xor XOR2 (N1195, N1190, N1003);
nor NOR3 (N1196, N1192, N1058, N805);
not NOT1 (N1197, N1191);
and AND2 (N1198, N1195, N145);
nand NAND2 (N1199, N1184, N358);
and AND3 (N1200, N1197, N85, N579);
xor XOR2 (N1201, N1194, N991);
xor XOR2 (N1202, N1189, N624);
not NOT1 (N1203, N1200);
or OR2 (N1204, N1203, N233);
buf BUF1 (N1205, N1193);
and AND4 (N1206, N1205, N569, N998, N922);
nand NAND2 (N1207, N1204, N1063);
nand NAND2 (N1208, N1196, N935);
nor NOR3 (N1209, N1206, N1153, N816);
buf BUF1 (N1210, N1201);
or OR3 (N1211, N1209, N701, N635);
xor XOR2 (N1212, N1211, N469);
nand NAND2 (N1213, N1176, N1007);
nor NOR4 (N1214, N1212, N717, N1125, N431);
nand NAND2 (N1215, N1188, N32);
buf BUF1 (N1216, N1210);
xor XOR2 (N1217, N1177, N875);
and AND3 (N1218, N1208, N930, N384);
and AND4 (N1219, N1215, N810, N695, N769);
nor NOR4 (N1220, N1214, N38, N1190, N1082);
buf BUF1 (N1221, N1213);
buf BUF1 (N1222, N1198);
nand NAND4 (N1223, N1217, N573, N435, N225);
or OR3 (N1224, N1220, N801, N598);
xor XOR2 (N1225, N1223, N33);
or OR2 (N1226, N1221, N1150);
buf BUF1 (N1227, N1224);
and AND2 (N1228, N1216, N86);
or OR2 (N1229, N1225, N1102);
not NOT1 (N1230, N1218);
not NOT1 (N1231, N1228);
nand NAND2 (N1232, N1199, N403);
nor NOR2 (N1233, N1222, N668);
xor XOR2 (N1234, N1232, N812);
buf BUF1 (N1235, N1207);
buf BUF1 (N1236, N1233);
not NOT1 (N1237, N1235);
and AND4 (N1238, N1219, N453, N907, N171);
xor XOR2 (N1239, N1202, N1123);
xor XOR2 (N1240, N1237, N720);
nor NOR4 (N1241, N1226, N769, N220, N71);
xor XOR2 (N1242, N1239, N76);
not NOT1 (N1243, N1242);
and AND4 (N1244, N1241, N299, N113, N866);
xor XOR2 (N1245, N1229, N573);
and AND2 (N1246, N1245, N601);
xor XOR2 (N1247, N1246, N1242);
xor XOR2 (N1248, N1244, N1196);
not NOT1 (N1249, N1236);
buf BUF1 (N1250, N1248);
xor XOR2 (N1251, N1240, N687);
not NOT1 (N1252, N1251);
not NOT1 (N1253, N1227);
nand NAND3 (N1254, N1252, N686, N685);
nand NAND2 (N1255, N1243, N35);
xor XOR2 (N1256, N1250, N92);
and AND4 (N1257, N1234, N526, N831, N723);
or OR2 (N1258, N1254, N433);
buf BUF1 (N1259, N1253);
nand NAND4 (N1260, N1255, N13, N1097, N596);
nand NAND2 (N1261, N1247, N1250);
or OR3 (N1262, N1256, N1025, N205);
buf BUF1 (N1263, N1238);
nand NAND2 (N1264, N1258, N546);
and AND4 (N1265, N1262, N1204, N826, N988);
and AND2 (N1266, N1261, N309);
and AND4 (N1267, N1249, N843, N224, N195);
not NOT1 (N1268, N1267);
xor XOR2 (N1269, N1257, N624);
xor XOR2 (N1270, N1268, N1044);
buf BUF1 (N1271, N1269);
xor XOR2 (N1272, N1259, N612);
or OR3 (N1273, N1271, N948, N536);
xor XOR2 (N1274, N1230, N96);
nand NAND2 (N1275, N1260, N611);
xor XOR2 (N1276, N1265, N1023);
xor XOR2 (N1277, N1272, N866);
buf BUF1 (N1278, N1273);
and AND3 (N1279, N1278, N1012, N394);
xor XOR2 (N1280, N1274, N1259);
xor XOR2 (N1281, N1266, N1062);
nand NAND4 (N1282, N1231, N377, N1069, N541);
xor XOR2 (N1283, N1270, N1241);
nand NAND2 (N1284, N1276, N45);
nand NAND4 (N1285, N1275, N272, N1177, N402);
xor XOR2 (N1286, N1263, N507);
and AND4 (N1287, N1279, N313, N885, N657);
nor NOR4 (N1288, N1286, N439, N648, N605);
buf BUF1 (N1289, N1277);
xor XOR2 (N1290, N1280, N1216);
nor NOR3 (N1291, N1281, N892, N787);
xor XOR2 (N1292, N1283, N509);
nor NOR3 (N1293, N1287, N1173, N862);
nor NOR3 (N1294, N1285, N767, N703);
and AND2 (N1295, N1294, N408);
nand NAND4 (N1296, N1295, N640, N524, N793);
and AND3 (N1297, N1296, N724, N1007);
buf BUF1 (N1298, N1291);
or OR2 (N1299, N1284, N918);
or OR4 (N1300, N1293, N1259, N937, N1146);
and AND2 (N1301, N1299, N944);
xor XOR2 (N1302, N1282, N995);
not NOT1 (N1303, N1300);
or OR2 (N1304, N1301, N557);
xor XOR2 (N1305, N1292, N10);
xor XOR2 (N1306, N1302, N1175);
buf BUF1 (N1307, N1304);
xor XOR2 (N1308, N1290, N1254);
not NOT1 (N1309, N1303);
nor NOR2 (N1310, N1297, N333);
and AND3 (N1311, N1310, N1172, N438);
buf BUF1 (N1312, N1311);
nand NAND4 (N1313, N1309, N868, N989, N1029);
and AND3 (N1314, N1288, N803, N786);
or OR2 (N1315, N1313, N577);
nand NAND3 (N1316, N1315, N480, N1166);
buf BUF1 (N1317, N1312);
or OR4 (N1318, N1316, N14, N988, N754);
nor NOR2 (N1319, N1308, N78);
nand NAND2 (N1320, N1307, N775);
nand NAND3 (N1321, N1264, N36, N986);
buf BUF1 (N1322, N1320);
nor NOR3 (N1323, N1314, N952, N213);
nand NAND4 (N1324, N1305, N706, N490, N997);
and AND2 (N1325, N1324, N769);
not NOT1 (N1326, N1298);
or OR3 (N1327, N1317, N701, N564);
not NOT1 (N1328, N1321);
and AND4 (N1329, N1319, N265, N1016, N1263);
or OR4 (N1330, N1329, N1075, N1233, N18);
not NOT1 (N1331, N1318);
and AND4 (N1332, N1331, N1075, N199, N1131);
and AND3 (N1333, N1326, N808, N762);
not NOT1 (N1334, N1322);
nor NOR3 (N1335, N1333, N121, N714);
nor NOR3 (N1336, N1335, N1197, N993);
buf BUF1 (N1337, N1328);
nor NOR3 (N1338, N1330, N101, N203);
nand NAND4 (N1339, N1334, N718, N731, N897);
buf BUF1 (N1340, N1338);
xor XOR2 (N1341, N1332, N669);
buf BUF1 (N1342, N1340);
nand NAND2 (N1343, N1327, N1110);
or OR3 (N1344, N1306, N497, N436);
nor NOR2 (N1345, N1344, N826);
or OR3 (N1346, N1323, N183, N293);
nor NOR3 (N1347, N1341, N1053, N198);
and AND4 (N1348, N1289, N674, N1122, N428);
not NOT1 (N1349, N1347);
and AND2 (N1350, N1339, N1134);
nand NAND3 (N1351, N1337, N1131, N667);
xor XOR2 (N1352, N1349, N427);
and AND2 (N1353, N1325, N369);
nor NOR4 (N1354, N1343, N857, N1248, N432);
or OR2 (N1355, N1348, N593);
xor XOR2 (N1356, N1345, N1048);
xor XOR2 (N1357, N1336, N649);
nor NOR4 (N1358, N1355, N384, N815, N627);
buf BUF1 (N1359, N1346);
nor NOR4 (N1360, N1356, N18, N1330, N898);
nand NAND4 (N1361, N1358, N1360, N139, N496);
and AND3 (N1362, N633, N75, N34);
not NOT1 (N1363, N1353);
not NOT1 (N1364, N1350);
nand NAND2 (N1365, N1342, N229);
not NOT1 (N1366, N1362);
nand NAND3 (N1367, N1351, N414, N1108);
or OR4 (N1368, N1354, N1289, N808, N1124);
xor XOR2 (N1369, N1368, N895);
xor XOR2 (N1370, N1361, N866);
xor XOR2 (N1371, N1369, N1060);
and AND4 (N1372, N1352, N820, N670, N198);
not NOT1 (N1373, N1364);
and AND2 (N1374, N1359, N1234);
buf BUF1 (N1375, N1363);
nor NOR4 (N1376, N1365, N450, N777, N172);
and AND3 (N1377, N1374, N1233, N916);
not NOT1 (N1378, N1376);
buf BUF1 (N1379, N1366);
buf BUF1 (N1380, N1379);
nand NAND2 (N1381, N1377, N629);
nand NAND3 (N1382, N1367, N301, N846);
buf BUF1 (N1383, N1378);
buf BUF1 (N1384, N1375);
xor XOR2 (N1385, N1373, N961);
buf BUF1 (N1386, N1383);
and AND2 (N1387, N1382, N1236);
nor NOR3 (N1388, N1385, N1067, N828);
not NOT1 (N1389, N1357);
and AND3 (N1390, N1389, N566, N1111);
xor XOR2 (N1391, N1380, N572);
buf BUF1 (N1392, N1381);
nand NAND4 (N1393, N1371, N632, N821, N1172);
buf BUF1 (N1394, N1388);
nor NOR3 (N1395, N1391, N1220, N335);
nand NAND4 (N1396, N1393, N147, N984, N137);
xor XOR2 (N1397, N1394, N1156);
nand NAND2 (N1398, N1384, N619);
not NOT1 (N1399, N1392);
or OR2 (N1400, N1390, N639);
nor NOR4 (N1401, N1397, N745, N904, N179);
xor XOR2 (N1402, N1370, N712);
not NOT1 (N1403, N1402);
not NOT1 (N1404, N1387);
or OR4 (N1405, N1404, N1142, N187, N780);
xor XOR2 (N1406, N1399, N1369);
or OR4 (N1407, N1401, N121, N483, N981);
and AND2 (N1408, N1405, N618);
xor XOR2 (N1409, N1372, N620);
nand NAND4 (N1410, N1403, N400, N867, N929);
xor XOR2 (N1411, N1410, N697);
buf BUF1 (N1412, N1406);
buf BUF1 (N1413, N1398);
xor XOR2 (N1414, N1407, N1387);
xor XOR2 (N1415, N1414, N992);
buf BUF1 (N1416, N1400);
nand NAND4 (N1417, N1413, N368, N1035, N303);
buf BUF1 (N1418, N1411);
xor XOR2 (N1419, N1408, N749);
nor NOR4 (N1420, N1386, N122, N716, N206);
nand NAND4 (N1421, N1417, N24, N358, N702);
or OR2 (N1422, N1419, N1042);
nor NOR4 (N1423, N1396, N473, N543, N1164);
nor NOR4 (N1424, N1422, N526, N1337, N904);
xor XOR2 (N1425, N1423, N779);
nand NAND4 (N1426, N1421, N1075, N1165, N1266);
nand NAND4 (N1427, N1412, N469, N1049, N542);
nor NOR3 (N1428, N1420, N1224, N1164);
buf BUF1 (N1429, N1427);
and AND3 (N1430, N1428, N1174, N83);
buf BUF1 (N1431, N1415);
nand NAND3 (N1432, N1424, N1171, N675);
nor NOR2 (N1433, N1426, N424);
xor XOR2 (N1434, N1430, N227);
buf BUF1 (N1435, N1425);
and AND4 (N1436, N1433, N337, N1196, N248);
and AND4 (N1437, N1432, N876, N1366, N877);
and AND3 (N1438, N1429, N1155, N403);
xor XOR2 (N1439, N1418, N957);
and AND4 (N1440, N1409, N1164, N115, N1240);
not NOT1 (N1441, N1416);
xor XOR2 (N1442, N1395, N447);
xor XOR2 (N1443, N1441, N1380);
or OR2 (N1444, N1442, N953);
xor XOR2 (N1445, N1439, N1404);
and AND4 (N1446, N1431, N527, N458, N684);
buf BUF1 (N1447, N1445);
buf BUF1 (N1448, N1444);
or OR2 (N1449, N1447, N96);
and AND4 (N1450, N1435, N722, N975, N791);
not NOT1 (N1451, N1446);
nor NOR2 (N1452, N1440, N236);
xor XOR2 (N1453, N1437, N660);
not NOT1 (N1454, N1453);
nor NOR3 (N1455, N1452, N405, N692);
or OR4 (N1456, N1455, N952, N1033, N1120);
not NOT1 (N1457, N1454);
nand NAND4 (N1458, N1436, N1097, N882, N345);
and AND2 (N1459, N1434, N385);
not NOT1 (N1460, N1456);
xor XOR2 (N1461, N1460, N132);
xor XOR2 (N1462, N1461, N411);
nand NAND3 (N1463, N1451, N40, N1204);
not NOT1 (N1464, N1458);
xor XOR2 (N1465, N1449, N459);
nor NOR4 (N1466, N1438, N230, N369, N1196);
not NOT1 (N1467, N1450);
and AND3 (N1468, N1463, N653, N855);
not NOT1 (N1469, N1466);
or OR2 (N1470, N1459, N88);
and AND3 (N1471, N1469, N1282, N1240);
not NOT1 (N1472, N1467);
not NOT1 (N1473, N1472);
xor XOR2 (N1474, N1471, N1253);
nand NAND2 (N1475, N1457, N1130);
or OR2 (N1476, N1465, N1170);
nand NAND3 (N1477, N1448, N595, N203);
nand NAND3 (N1478, N1475, N1461, N99);
buf BUF1 (N1479, N1468);
or OR2 (N1480, N1462, N542);
not NOT1 (N1481, N1479);
and AND4 (N1482, N1477, N1368, N731, N1012);
not NOT1 (N1483, N1473);
buf BUF1 (N1484, N1470);
nor NOR3 (N1485, N1443, N833, N347);
xor XOR2 (N1486, N1481, N1272);
buf BUF1 (N1487, N1484);
or OR2 (N1488, N1485, N1462);
nand NAND4 (N1489, N1478, N1069, N1416, N1327);
nand NAND4 (N1490, N1482, N1209, N1142, N517);
not NOT1 (N1491, N1488);
nor NOR4 (N1492, N1490, N1278, N1198, N1214);
or OR2 (N1493, N1483, N855);
not NOT1 (N1494, N1476);
and AND3 (N1495, N1487, N715, N508);
and AND4 (N1496, N1480, N1082, N1228, N181);
nand NAND4 (N1497, N1492, N467, N108, N24);
not NOT1 (N1498, N1497);
nor NOR4 (N1499, N1491, N682, N75, N1190);
and AND4 (N1500, N1499, N960, N1145, N464);
not NOT1 (N1501, N1498);
nor NOR4 (N1502, N1501, N1051, N340, N807);
nand NAND2 (N1503, N1495, N623);
buf BUF1 (N1504, N1502);
not NOT1 (N1505, N1464);
buf BUF1 (N1506, N1503);
buf BUF1 (N1507, N1506);
xor XOR2 (N1508, N1504, N1268);
and AND3 (N1509, N1507, N76, N1163);
not NOT1 (N1510, N1474);
not NOT1 (N1511, N1500);
nor NOR2 (N1512, N1496, N1378);
not NOT1 (N1513, N1511);
nor NOR3 (N1514, N1512, N181, N839);
or OR3 (N1515, N1489, N60, N457);
and AND3 (N1516, N1515, N1228, N1193);
xor XOR2 (N1517, N1516, N1046);
and AND3 (N1518, N1513, N1140, N1318);
xor XOR2 (N1519, N1493, N874);
and AND3 (N1520, N1505, N164, N1304);
not NOT1 (N1521, N1519);
nor NOR3 (N1522, N1486, N1470, N700);
not NOT1 (N1523, N1508);
nor NOR2 (N1524, N1521, N294);
not NOT1 (N1525, N1522);
not NOT1 (N1526, N1510);
not NOT1 (N1527, N1517);
or OR2 (N1528, N1520, N527);
nor NOR2 (N1529, N1518, N806);
nand NAND2 (N1530, N1523, N271);
nand NAND4 (N1531, N1525, N881, N312, N788);
nand NAND3 (N1532, N1524, N1515, N507);
or OR4 (N1533, N1528, N1256, N85, N1165);
and AND3 (N1534, N1527, N1203, N694);
or OR4 (N1535, N1532, N911, N357, N1070);
not NOT1 (N1536, N1533);
xor XOR2 (N1537, N1535, N1107);
nor NOR3 (N1538, N1494, N69, N103);
nand NAND4 (N1539, N1531, N296, N160, N709);
buf BUF1 (N1540, N1514);
not NOT1 (N1541, N1534);
not NOT1 (N1542, N1537);
xor XOR2 (N1543, N1529, N211);
nand NAND3 (N1544, N1541, N383, N620);
not NOT1 (N1545, N1538);
or OR4 (N1546, N1544, N808, N870, N568);
not NOT1 (N1547, N1539);
and AND3 (N1548, N1509, N248, N128);
nand NAND2 (N1549, N1543, N1162);
buf BUF1 (N1550, N1546);
buf BUF1 (N1551, N1548);
buf BUF1 (N1552, N1540);
not NOT1 (N1553, N1530);
and AND3 (N1554, N1526, N10, N1414);
nor NOR2 (N1555, N1542, N294);
buf BUF1 (N1556, N1550);
nor NOR4 (N1557, N1547, N335, N445, N316);
and AND3 (N1558, N1556, N426, N268);
buf BUF1 (N1559, N1558);
and AND3 (N1560, N1559, N1114, N603);
buf BUF1 (N1561, N1557);
buf BUF1 (N1562, N1551);
buf BUF1 (N1563, N1553);
nor NOR4 (N1564, N1552, N467, N727, N795);
and AND4 (N1565, N1554, N749, N1485, N206);
buf BUF1 (N1566, N1545);
nand NAND3 (N1567, N1566, N199, N561);
or OR2 (N1568, N1549, N667);
nor NOR2 (N1569, N1560, N821);
nand NAND2 (N1570, N1536, N897);
and AND4 (N1571, N1567, N1341, N1026, N2);
xor XOR2 (N1572, N1570, N833);
and AND3 (N1573, N1563, N1373, N1346);
nor NOR3 (N1574, N1562, N717, N1049);
nor NOR3 (N1575, N1573, N945, N571);
nor NOR3 (N1576, N1569, N503, N1039);
buf BUF1 (N1577, N1561);
buf BUF1 (N1578, N1555);
or OR2 (N1579, N1568, N1000);
nor NOR4 (N1580, N1578, N402, N337, N658);
not NOT1 (N1581, N1579);
nand NAND3 (N1582, N1565, N887, N740);
and AND2 (N1583, N1575, N389);
nor NOR3 (N1584, N1581, N1396, N509);
xor XOR2 (N1585, N1574, N1396);
or OR4 (N1586, N1580, N223, N1358, N760);
xor XOR2 (N1587, N1571, N1580);
and AND4 (N1588, N1582, N1190, N445, N783);
xor XOR2 (N1589, N1588, N1339);
or OR4 (N1590, N1585, N113, N53, N1438);
and AND3 (N1591, N1587, N798, N1485);
nand NAND3 (N1592, N1586, N1457, N751);
xor XOR2 (N1593, N1572, N832);
nand NAND2 (N1594, N1564, N1289);
and AND2 (N1595, N1594, N82);
xor XOR2 (N1596, N1576, N1011);
nor NOR4 (N1597, N1593, N715, N328, N127);
xor XOR2 (N1598, N1597, N395);
buf BUF1 (N1599, N1598);
nor NOR3 (N1600, N1590, N942, N931);
nand NAND2 (N1601, N1577, N1583);
and AND2 (N1602, N830, N729);
nand NAND2 (N1603, N1595, N1427);
nor NOR2 (N1604, N1599, N1302);
not NOT1 (N1605, N1600);
nor NOR4 (N1606, N1601, N1263, N422, N1204);
or OR4 (N1607, N1602, N1567, N560, N823);
and AND4 (N1608, N1604, N433, N98, N608);
nor NOR3 (N1609, N1607, N838, N1237);
nand NAND4 (N1610, N1589, N384, N1325, N501);
buf BUF1 (N1611, N1606);
xor XOR2 (N1612, N1609, N379);
buf BUF1 (N1613, N1603);
xor XOR2 (N1614, N1612, N216);
or OR4 (N1615, N1596, N376, N737, N336);
or OR4 (N1616, N1591, N376, N1296, N1447);
nand NAND4 (N1617, N1584, N701, N1373, N1085);
or OR2 (N1618, N1616, N115);
xor XOR2 (N1619, N1610, N1182);
or OR3 (N1620, N1615, N959, N1227);
nand NAND2 (N1621, N1592, N1143);
buf BUF1 (N1622, N1618);
or OR4 (N1623, N1619, N720, N1044, N314);
buf BUF1 (N1624, N1621);
buf BUF1 (N1625, N1624);
xor XOR2 (N1626, N1613, N102);
buf BUF1 (N1627, N1623);
and AND2 (N1628, N1605, N899);
nand NAND4 (N1629, N1620, N535, N1307, N966);
and AND3 (N1630, N1627, N1076, N216);
xor XOR2 (N1631, N1630, N961);
xor XOR2 (N1632, N1629, N695);
buf BUF1 (N1633, N1632);
buf BUF1 (N1634, N1608);
not NOT1 (N1635, N1628);
nor NOR2 (N1636, N1622, N535);
not NOT1 (N1637, N1634);
or OR4 (N1638, N1625, N1301, N1153, N1337);
xor XOR2 (N1639, N1626, N193);
buf BUF1 (N1640, N1637);
xor XOR2 (N1641, N1631, N1179);
or OR3 (N1642, N1611, N1117, N1622);
xor XOR2 (N1643, N1641, N1642);
nand NAND2 (N1644, N1419, N49);
nor NOR4 (N1645, N1643, N686, N768, N1071);
nor NOR3 (N1646, N1638, N532, N1472);
xor XOR2 (N1647, N1645, N597);
or OR4 (N1648, N1647, N1027, N459, N1088);
nand NAND4 (N1649, N1644, N241, N1130, N832);
nand NAND3 (N1650, N1640, N331, N1437);
nor NOR4 (N1651, N1646, N715, N219, N1540);
xor XOR2 (N1652, N1649, N1501);
xor XOR2 (N1653, N1650, N479);
buf BUF1 (N1654, N1636);
or OR4 (N1655, N1648, N784, N888, N1008);
nand NAND3 (N1656, N1633, N1189, N805);
and AND3 (N1657, N1639, N1401, N503);
and AND3 (N1658, N1653, N1486, N1470);
buf BUF1 (N1659, N1617);
buf BUF1 (N1660, N1652);
nand NAND4 (N1661, N1656, N1193, N1208, N874);
and AND3 (N1662, N1657, N860, N588);
or OR4 (N1663, N1651, N665, N90, N349);
or OR4 (N1664, N1660, N1067, N1645, N179);
not NOT1 (N1665, N1635);
nor NOR2 (N1666, N1665, N1374);
and AND2 (N1667, N1614, N888);
nor NOR3 (N1668, N1662, N256, N340);
xor XOR2 (N1669, N1664, N468);
nand NAND2 (N1670, N1661, N801);
and AND2 (N1671, N1666, N572);
xor XOR2 (N1672, N1671, N250);
not NOT1 (N1673, N1672);
and AND4 (N1674, N1655, N663, N398, N1487);
nand NAND2 (N1675, N1674, N839);
nand NAND2 (N1676, N1670, N1574);
buf BUF1 (N1677, N1673);
nand NAND2 (N1678, N1659, N1586);
and AND2 (N1679, N1667, N1484);
and AND2 (N1680, N1663, N1607);
xor XOR2 (N1681, N1675, N395);
buf BUF1 (N1682, N1680);
nand NAND2 (N1683, N1676, N431);
nand NAND4 (N1684, N1683, N183, N1669, N1248);
nor NOR4 (N1685, N1251, N887, N483, N1455);
xor XOR2 (N1686, N1681, N1030);
not NOT1 (N1687, N1685);
xor XOR2 (N1688, N1687, N1296);
nand NAND2 (N1689, N1688, N1266);
not NOT1 (N1690, N1682);
or OR2 (N1691, N1678, N175);
buf BUF1 (N1692, N1689);
nand NAND2 (N1693, N1658, N418);
xor XOR2 (N1694, N1679, N902);
or OR4 (N1695, N1654, N977, N513, N1642);
and AND3 (N1696, N1668, N421, N1164);
or OR2 (N1697, N1690, N992);
xor XOR2 (N1698, N1686, N198);
buf BUF1 (N1699, N1677);
xor XOR2 (N1700, N1695, N923);
nor NOR4 (N1701, N1697, N553, N677, N1378);
xor XOR2 (N1702, N1699, N398);
not NOT1 (N1703, N1692);
buf BUF1 (N1704, N1693);
not NOT1 (N1705, N1701);
not NOT1 (N1706, N1691);
or OR2 (N1707, N1698, N1250);
and AND4 (N1708, N1704, N265, N832, N1161);
xor XOR2 (N1709, N1702, N987);
not NOT1 (N1710, N1705);
xor XOR2 (N1711, N1703, N1346);
nand NAND2 (N1712, N1684, N1365);
not NOT1 (N1713, N1712);
nor NOR3 (N1714, N1700, N701, N1631);
and AND2 (N1715, N1709, N1034);
or OR2 (N1716, N1715, N321);
nor NOR4 (N1717, N1713, N914, N1623, N553);
nand NAND2 (N1718, N1711, N97);
nor NOR3 (N1719, N1716, N1153, N1178);
buf BUF1 (N1720, N1694);
and AND4 (N1721, N1708, N115, N1077, N484);
xor XOR2 (N1722, N1717, N384);
not NOT1 (N1723, N1722);
nand NAND2 (N1724, N1706, N483);
nor NOR3 (N1725, N1718, N1096, N360);
nor NOR3 (N1726, N1725, N354, N16);
buf BUF1 (N1727, N1714);
xor XOR2 (N1728, N1721, N117);
xor XOR2 (N1729, N1726, N1039);
xor XOR2 (N1730, N1696, N502);
and AND4 (N1731, N1710, N177, N668, N721);
or OR2 (N1732, N1724, N761);
or OR4 (N1733, N1729, N377, N1086, N1558);
not NOT1 (N1734, N1723);
not NOT1 (N1735, N1730);
nand NAND2 (N1736, N1732, N742);
not NOT1 (N1737, N1735);
buf BUF1 (N1738, N1734);
or OR3 (N1739, N1719, N1302, N151);
and AND2 (N1740, N1707, N849);
or OR2 (N1741, N1728, N191);
and AND2 (N1742, N1727, N138);
buf BUF1 (N1743, N1736);
buf BUF1 (N1744, N1740);
not NOT1 (N1745, N1738);
nand NAND3 (N1746, N1733, N178, N1558);
buf BUF1 (N1747, N1741);
nand NAND3 (N1748, N1745, N313, N1500);
nand NAND2 (N1749, N1743, N1079);
or OR4 (N1750, N1748, N210, N1327, N1218);
buf BUF1 (N1751, N1737);
or OR2 (N1752, N1749, N1141);
buf BUF1 (N1753, N1720);
xor XOR2 (N1754, N1739, N525);
nor NOR3 (N1755, N1742, N1505, N145);
nor NOR3 (N1756, N1752, N1039, N1718);
nor NOR4 (N1757, N1731, N1604, N1290, N517);
buf BUF1 (N1758, N1750);
not NOT1 (N1759, N1757);
and AND4 (N1760, N1751, N247, N772, N1181);
nor NOR2 (N1761, N1759, N269);
xor XOR2 (N1762, N1746, N1706);
nand NAND2 (N1763, N1758, N1013);
xor XOR2 (N1764, N1754, N1708);
not NOT1 (N1765, N1762);
nand NAND2 (N1766, N1744, N1115);
not NOT1 (N1767, N1761);
or OR3 (N1768, N1766, N490, N940);
nor NOR3 (N1769, N1747, N45, N530);
buf BUF1 (N1770, N1764);
xor XOR2 (N1771, N1765, N320);
nand NAND4 (N1772, N1770, N1649, N657, N316);
and AND2 (N1773, N1771, N667);
and AND3 (N1774, N1753, N857, N1642);
nor NOR2 (N1775, N1756, N537);
xor XOR2 (N1776, N1775, N1500);
not NOT1 (N1777, N1773);
or OR3 (N1778, N1755, N15, N1321);
xor XOR2 (N1779, N1768, N524);
nand NAND3 (N1780, N1774, N532, N1551);
nor NOR4 (N1781, N1763, N1688, N1044, N851);
xor XOR2 (N1782, N1772, N614);
xor XOR2 (N1783, N1776, N794);
xor XOR2 (N1784, N1780, N300);
xor XOR2 (N1785, N1769, N1371);
nor NOR4 (N1786, N1778, N1775, N398, N1322);
or OR4 (N1787, N1784, N878, N1641, N12);
nand NAND2 (N1788, N1779, N193);
xor XOR2 (N1789, N1777, N1446);
xor XOR2 (N1790, N1785, N699);
xor XOR2 (N1791, N1786, N35);
nor NOR4 (N1792, N1782, N1320, N191, N1098);
nand NAND2 (N1793, N1792, N1260);
or OR4 (N1794, N1788, N501, N606, N336);
or OR3 (N1795, N1794, N1212, N938);
xor XOR2 (N1796, N1781, N1721);
not NOT1 (N1797, N1793);
and AND2 (N1798, N1787, N1745);
xor XOR2 (N1799, N1796, N322);
xor XOR2 (N1800, N1797, N679);
not NOT1 (N1801, N1783);
or OR2 (N1802, N1801, N1413);
nor NOR3 (N1803, N1795, N191, N1264);
and AND4 (N1804, N1790, N1666, N234, N1276);
nand NAND2 (N1805, N1803, N536);
not NOT1 (N1806, N1767);
and AND2 (N1807, N1802, N1532);
buf BUF1 (N1808, N1807);
xor XOR2 (N1809, N1804, N49);
and AND3 (N1810, N1800, N36, N518);
not NOT1 (N1811, N1810);
nor NOR4 (N1812, N1805, N109, N1231, N1639);
xor XOR2 (N1813, N1812, N847);
or OR2 (N1814, N1789, N393);
nand NAND3 (N1815, N1809, N733, N1799);
xor XOR2 (N1816, N395, N742);
nor NOR4 (N1817, N1816, N1655, N232, N1381);
nor NOR4 (N1818, N1813, N1801, N982, N1456);
xor XOR2 (N1819, N1811, N89);
nor NOR2 (N1820, N1760, N265);
or OR3 (N1821, N1819, N985, N701);
or OR4 (N1822, N1814, N455, N444, N141);
and AND3 (N1823, N1820, N9, N591);
or OR2 (N1824, N1806, N1365);
xor XOR2 (N1825, N1815, N769);
or OR2 (N1826, N1821, N757);
not NOT1 (N1827, N1823);
and AND4 (N1828, N1827, N1729, N1599, N607);
or OR4 (N1829, N1798, N260, N163, N110);
buf BUF1 (N1830, N1828);
xor XOR2 (N1831, N1824, N746);
nand NAND4 (N1832, N1825, N158, N1012, N1814);
nand NAND2 (N1833, N1822, N1773);
buf BUF1 (N1834, N1831);
and AND4 (N1835, N1833, N374, N246, N1012);
nand NAND2 (N1836, N1817, N1247);
nand NAND3 (N1837, N1832, N1497, N384);
nor NOR4 (N1838, N1836, N160, N60, N704);
buf BUF1 (N1839, N1834);
nand NAND4 (N1840, N1808, N349, N1200, N1839);
nor NOR3 (N1841, N603, N938, N260);
xor XOR2 (N1842, N1837, N1165);
and AND4 (N1843, N1826, N1076, N585, N914);
nand NAND4 (N1844, N1838, N1577, N975, N27);
nor NOR2 (N1845, N1841, N196);
and AND3 (N1846, N1829, N1834, N111);
and AND4 (N1847, N1844, N1651, N1336, N730);
not NOT1 (N1848, N1842);
and AND2 (N1849, N1848, N680);
or OR2 (N1850, N1835, N407);
buf BUF1 (N1851, N1846);
buf BUF1 (N1852, N1847);
not NOT1 (N1853, N1791);
nand NAND4 (N1854, N1818, N964, N1552, N1383);
and AND3 (N1855, N1853, N904, N450);
xor XOR2 (N1856, N1840, N725);
and AND3 (N1857, N1855, N746, N1112);
or OR2 (N1858, N1857, N1190);
nor NOR4 (N1859, N1845, N1459, N1367, N217);
nor NOR3 (N1860, N1854, N488, N919);
and AND2 (N1861, N1849, N364);
xor XOR2 (N1862, N1860, N1568);
not NOT1 (N1863, N1851);
xor XOR2 (N1864, N1863, N1748);
and AND2 (N1865, N1852, N1249);
buf BUF1 (N1866, N1843);
or OR3 (N1867, N1858, N682, N815);
and AND2 (N1868, N1866, N1287);
xor XOR2 (N1869, N1856, N84);
xor XOR2 (N1870, N1865, N1043);
nand NAND3 (N1871, N1830, N1257, N519);
xor XOR2 (N1872, N1868, N1004);
not NOT1 (N1873, N1862);
and AND4 (N1874, N1872, N1864, N1245, N1343);
nand NAND3 (N1875, N1168, N1333, N1247);
nor NOR2 (N1876, N1859, N1561);
xor XOR2 (N1877, N1874, N1394);
not NOT1 (N1878, N1876);
nor NOR3 (N1879, N1867, N1798, N1122);
not NOT1 (N1880, N1875);
nand NAND4 (N1881, N1869, N1152, N615, N430);
nand NAND3 (N1882, N1878, N1113, N1271);
buf BUF1 (N1883, N1877);
not NOT1 (N1884, N1850);
or OR2 (N1885, N1871, N214);
not NOT1 (N1886, N1885);
buf BUF1 (N1887, N1883);
nand NAND2 (N1888, N1887, N1312);
buf BUF1 (N1889, N1886);
nor NOR4 (N1890, N1879, N1026, N356, N476);
and AND3 (N1891, N1861, N1437, N193);
nor NOR3 (N1892, N1889, N119, N1793);
xor XOR2 (N1893, N1882, N332);
buf BUF1 (N1894, N1888);
or OR3 (N1895, N1892, N1028, N158);
nand NAND4 (N1896, N1870, N53, N600, N641);
not NOT1 (N1897, N1884);
nand NAND2 (N1898, N1896, N918);
xor XOR2 (N1899, N1898, N1427);
xor XOR2 (N1900, N1895, N1564);
and AND4 (N1901, N1890, N1674, N255, N1704);
and AND3 (N1902, N1893, N71, N873);
xor XOR2 (N1903, N1897, N374);
or OR2 (N1904, N1899, N59);
nand NAND2 (N1905, N1900, N432);
nor NOR3 (N1906, N1891, N1723, N409);
and AND4 (N1907, N1906, N1555, N352, N691);
not NOT1 (N1908, N1894);
and AND3 (N1909, N1903, N1355, N680);
and AND2 (N1910, N1908, N77);
nand NAND3 (N1911, N1901, N102, N450);
not NOT1 (N1912, N1880);
and AND3 (N1913, N1873, N36, N688);
or OR4 (N1914, N1905, N145, N1503, N464);
or OR4 (N1915, N1912, N690, N1813, N1059);
not NOT1 (N1916, N1911);
not NOT1 (N1917, N1910);
buf BUF1 (N1918, N1907);
nor NOR3 (N1919, N1902, N786, N1398);
not NOT1 (N1920, N1881);
nand NAND4 (N1921, N1913, N1803, N1083, N975);
nand NAND2 (N1922, N1917, N1787);
buf BUF1 (N1923, N1918);
not NOT1 (N1924, N1921);
nor NOR2 (N1925, N1916, N554);
or OR3 (N1926, N1914, N1708, N31);
nor NOR2 (N1927, N1909, N1290);
nand NAND2 (N1928, N1924, N1842);
nand NAND3 (N1929, N1922, N1423, N844);
and AND4 (N1930, N1923, N750, N1737, N1083);
not NOT1 (N1931, N1927);
and AND3 (N1932, N1930, N672, N1696);
xor XOR2 (N1933, N1929, N45);
or OR2 (N1934, N1904, N264);
buf BUF1 (N1935, N1915);
or OR2 (N1936, N1931, N17);
nor NOR4 (N1937, N1928, N1662, N1522, N1294);
nor NOR2 (N1938, N1925, N872);
and AND2 (N1939, N1936, N1297);
not NOT1 (N1940, N1935);
not NOT1 (N1941, N1939);
nor NOR3 (N1942, N1926, N1774, N141);
nand NAND2 (N1943, N1919, N883);
not NOT1 (N1944, N1942);
or OR4 (N1945, N1932, N684, N860, N238);
nand NAND2 (N1946, N1933, N1921);
nand NAND2 (N1947, N1941, N1506);
nor NOR2 (N1948, N1940, N1803);
nor NOR4 (N1949, N1947, N115, N1412, N316);
buf BUF1 (N1950, N1944);
nand NAND2 (N1951, N1943, N1933);
or OR4 (N1952, N1948, N227, N1874, N1893);
xor XOR2 (N1953, N1949, N667);
xor XOR2 (N1954, N1920, N422);
nor NOR4 (N1955, N1952, N1226, N782, N1947);
buf BUF1 (N1956, N1945);
nor NOR4 (N1957, N1937, N1260, N963, N644);
buf BUF1 (N1958, N1954);
and AND3 (N1959, N1950, N1864, N658);
xor XOR2 (N1960, N1956, N1137);
not NOT1 (N1961, N1951);
nor NOR3 (N1962, N1961, N1794, N573);
not NOT1 (N1963, N1938);
not NOT1 (N1964, N1934);
and AND2 (N1965, N1955, N1068);
not NOT1 (N1966, N1957);
and AND2 (N1967, N1959, N1419);
xor XOR2 (N1968, N1960, N1699);
or OR3 (N1969, N1962, N1911, N506);
not NOT1 (N1970, N1964);
or OR2 (N1971, N1963, N1381);
buf BUF1 (N1972, N1967);
xor XOR2 (N1973, N1970, N285);
nor NOR4 (N1974, N1969, N1930, N1381, N498);
nor NOR2 (N1975, N1972, N912);
xor XOR2 (N1976, N1974, N234);
or OR2 (N1977, N1946, N1158);
and AND2 (N1978, N1973, N1358);
nor NOR2 (N1979, N1976, N1329);
or OR3 (N1980, N1978, N406, N687);
buf BUF1 (N1981, N1966);
buf BUF1 (N1982, N1953);
nand NAND3 (N1983, N1979, N1014, N1156);
xor XOR2 (N1984, N1977, N1148);
or OR4 (N1985, N1981, N527, N847, N261);
nor NOR2 (N1986, N1983, N394);
nor NOR4 (N1987, N1980, N197, N1755, N850);
nand NAND3 (N1988, N1965, N1203, N1677);
or OR2 (N1989, N1982, N1171);
nand NAND2 (N1990, N1971, N1730);
xor XOR2 (N1991, N1986, N998);
or OR3 (N1992, N1987, N67, N160);
and AND3 (N1993, N1991, N333, N1043);
nor NOR2 (N1994, N1993, N1938);
not NOT1 (N1995, N1984);
buf BUF1 (N1996, N1988);
xor XOR2 (N1997, N1996, N1436);
buf BUF1 (N1998, N1985);
not NOT1 (N1999, N1975);
nor NOR4 (N2000, N1958, N1575, N869, N1629);
nor NOR3 (N2001, N1994, N1594, N628);
not NOT1 (N2002, N1992);
xor XOR2 (N2003, N1989, N469);
buf BUF1 (N2004, N2003);
not NOT1 (N2005, N2001);
buf BUF1 (N2006, N1997);
nor NOR3 (N2007, N2000, N215, N506);
xor XOR2 (N2008, N1998, N820);
nor NOR3 (N2009, N2002, N654, N191);
xor XOR2 (N2010, N2008, N589);
or OR3 (N2011, N2009, N1969, N1052);
nor NOR2 (N2012, N2005, N708);
or OR2 (N2013, N1999, N1624);
not NOT1 (N2014, N2010);
nand NAND3 (N2015, N2011, N70, N1756);
xor XOR2 (N2016, N2004, N67);
nor NOR4 (N2017, N2013, N1494, N1826, N908);
nand NAND2 (N2018, N2017, N855);
or OR2 (N2019, N2015, N478);
nor NOR4 (N2020, N1995, N934, N947, N536);
or OR2 (N2021, N2014, N1603);
or OR3 (N2022, N2016, N1396, N1918);
nand NAND4 (N2023, N1990, N875, N295, N1104);
buf BUF1 (N2024, N2019);
or OR3 (N2025, N2022, N1067, N242);
xor XOR2 (N2026, N2021, N2012);
not NOT1 (N2027, N1825);
nor NOR4 (N2028, N1968, N57, N445, N1450);
buf BUF1 (N2029, N2007);
xor XOR2 (N2030, N2023, N1652);
xor XOR2 (N2031, N2025, N1143);
buf BUF1 (N2032, N2030);
xor XOR2 (N2033, N2031, N1459);
buf BUF1 (N2034, N2028);
and AND4 (N2035, N2018, N915, N1493, N1095);
not NOT1 (N2036, N2027);
and AND4 (N2037, N2020, N950, N2005, N562);
buf BUF1 (N2038, N2036);
nor NOR4 (N2039, N2034, N173, N1398, N1105);
nor NOR3 (N2040, N2006, N1529, N1486);
nand NAND3 (N2041, N2035, N1406, N1803);
xor XOR2 (N2042, N2037, N1583);
not NOT1 (N2043, N2033);
not NOT1 (N2044, N2032);
or OR4 (N2045, N2042, N697, N1853, N141);
xor XOR2 (N2046, N2039, N323);
and AND4 (N2047, N2026, N1004, N24, N310);
not NOT1 (N2048, N2040);
nor NOR4 (N2049, N2041, N1692, N567, N211);
nor NOR2 (N2050, N2048, N1928);
buf BUF1 (N2051, N2045);
and AND2 (N2052, N2046, N554);
xor XOR2 (N2053, N2047, N1072);
buf BUF1 (N2054, N2043);
not NOT1 (N2055, N2038);
xor XOR2 (N2056, N2055, N967);
not NOT1 (N2057, N2050);
nor NOR3 (N2058, N2044, N440, N925);
or OR3 (N2059, N2054, N552, N740);
or OR3 (N2060, N2057, N1946, N102);
xor XOR2 (N2061, N2056, N247);
xor XOR2 (N2062, N2029, N2059);
and AND2 (N2063, N1624, N199);
or OR3 (N2064, N2060, N1311, N683);
or OR3 (N2065, N2049, N1626, N1226);
xor XOR2 (N2066, N2063, N1926);
nor NOR4 (N2067, N2064, N296, N1429, N933);
xor XOR2 (N2068, N2061, N1077);
nand NAND3 (N2069, N2068, N1139, N460);
xor XOR2 (N2070, N2062, N1818);
buf BUF1 (N2071, N2070);
or OR2 (N2072, N2066, N171);
nand NAND3 (N2073, N2065, N916, N657);
and AND2 (N2074, N2024, N30);
nor NOR2 (N2075, N2072, N949);
nand NAND3 (N2076, N2074, N1953, N845);
buf BUF1 (N2077, N2075);
or OR2 (N2078, N2051, N2008);
not NOT1 (N2079, N2073);
not NOT1 (N2080, N2053);
nor NOR3 (N2081, N2071, N790, N1944);
not NOT1 (N2082, N2079);
nor NOR4 (N2083, N2052, N1501, N316, N161);
xor XOR2 (N2084, N2067, N1437);
and AND4 (N2085, N2058, N1180, N307, N1814);
nand NAND3 (N2086, N2081, N1719, N1092);
and AND2 (N2087, N2083, N858);
xor XOR2 (N2088, N2086, N2083);
buf BUF1 (N2089, N2076);
not NOT1 (N2090, N2082);
not NOT1 (N2091, N2078);
nor NOR2 (N2092, N2091, N650);
or OR3 (N2093, N2080, N1933, N1223);
or OR3 (N2094, N2087, N171, N1069);
and AND2 (N2095, N2092, N1783);
xor XOR2 (N2096, N2077, N881);
xor XOR2 (N2097, N2084, N1422);
nor NOR4 (N2098, N2093, N1604, N1815, N603);
nor NOR3 (N2099, N2085, N567, N1165);
buf BUF1 (N2100, N2096);
nor NOR2 (N2101, N2097, N1609);
xor XOR2 (N2102, N2098, N1938);
xor XOR2 (N2103, N2095, N288);
not NOT1 (N2104, N2099);
and AND4 (N2105, N2101, N1881, N249, N974);
nor NOR2 (N2106, N2090, N1043);
nor NOR2 (N2107, N2089, N639);
nand NAND4 (N2108, N2100, N1197, N874, N1633);
nor NOR2 (N2109, N2108, N1853);
not NOT1 (N2110, N2094);
and AND2 (N2111, N2109, N693);
xor XOR2 (N2112, N2106, N516);
not NOT1 (N2113, N2107);
buf BUF1 (N2114, N2102);
and AND3 (N2115, N2113, N806, N1729);
buf BUF1 (N2116, N2105);
xor XOR2 (N2117, N2114, N2109);
and AND3 (N2118, N2069, N478, N1232);
buf BUF1 (N2119, N2117);
nor NOR3 (N2120, N2115, N188, N665);
not NOT1 (N2121, N2119);
xor XOR2 (N2122, N2111, N1363);
nand NAND2 (N2123, N2122, N110);
and AND3 (N2124, N2110, N1526, N1882);
nand NAND4 (N2125, N2121, N489, N298, N2040);
or OR3 (N2126, N2088, N964, N1092);
buf BUF1 (N2127, N2104);
and AND3 (N2128, N2120, N2089, N946);
and AND2 (N2129, N2128, N495);
xor XOR2 (N2130, N2123, N74);
or OR4 (N2131, N2126, N268, N1505, N17);
nand NAND2 (N2132, N2129, N1755);
xor XOR2 (N2133, N2103, N1214);
nand NAND4 (N2134, N2125, N215, N260, N986);
or OR2 (N2135, N2112, N228);
buf BUF1 (N2136, N2118);
not NOT1 (N2137, N2127);
buf BUF1 (N2138, N2133);
nor NOR2 (N2139, N2134, N1736);
xor XOR2 (N2140, N2138, N569);
and AND3 (N2141, N2140, N1576, N1413);
xor XOR2 (N2142, N2130, N1012);
not NOT1 (N2143, N2137);
xor XOR2 (N2144, N2131, N989);
and AND3 (N2145, N2144, N99, N1145);
not NOT1 (N2146, N2135);
or OR3 (N2147, N2136, N1417, N798);
or OR2 (N2148, N2139, N459);
xor XOR2 (N2149, N2146, N1393);
nand NAND4 (N2150, N2142, N1833, N1655, N1694);
xor XOR2 (N2151, N2150, N1787);
nand NAND3 (N2152, N2124, N281, N392);
nor NOR3 (N2153, N2145, N1975, N1809);
or OR4 (N2154, N2143, N474, N428, N753);
buf BUF1 (N2155, N2154);
nor NOR4 (N2156, N2132, N1784, N1444, N616);
or OR2 (N2157, N2147, N1348);
nor NOR3 (N2158, N2152, N331, N2155);
or OR2 (N2159, N2076, N1265);
and AND4 (N2160, N2149, N1903, N1992, N1512);
xor XOR2 (N2161, N2151, N1855);
not NOT1 (N2162, N2161);
nand NAND2 (N2163, N2116, N1004);
or OR4 (N2164, N2156, N2, N420, N2046);
or OR2 (N2165, N2159, N1464);
xor XOR2 (N2166, N2153, N2088);
or OR2 (N2167, N2160, N1746);
buf BUF1 (N2168, N2167);
not NOT1 (N2169, N2164);
xor XOR2 (N2170, N2148, N1022);
nor NOR4 (N2171, N2166, N1360, N2050, N853);
nor NOR2 (N2172, N2163, N67);
nand NAND2 (N2173, N2171, N696);
and AND2 (N2174, N2170, N1414);
buf BUF1 (N2175, N2158);
not NOT1 (N2176, N2172);
or OR4 (N2177, N2169, N297, N931, N426);
nand NAND4 (N2178, N2177, N576, N876, N1773);
and AND3 (N2179, N2168, N1148, N261);
xor XOR2 (N2180, N2174, N786);
buf BUF1 (N2181, N2179);
or OR4 (N2182, N2180, N350, N1161, N1414);
nor NOR3 (N2183, N2175, N610, N122);
not NOT1 (N2184, N2183);
xor XOR2 (N2185, N2141, N82);
nand NAND3 (N2186, N2165, N764, N1398);
buf BUF1 (N2187, N2157);
nand NAND3 (N2188, N2185, N199, N1428);
nand NAND3 (N2189, N2186, N1249, N167);
or OR2 (N2190, N2178, N36);
nand NAND4 (N2191, N2189, N1949, N397, N84);
nand NAND4 (N2192, N2173, N284, N1989, N1878);
not NOT1 (N2193, N2192);
not NOT1 (N2194, N2190);
nor NOR3 (N2195, N2176, N484, N1973);
buf BUF1 (N2196, N2191);
buf BUF1 (N2197, N2196);
or OR2 (N2198, N2181, N1469);
xor XOR2 (N2199, N2184, N1274);
xor XOR2 (N2200, N2182, N235);
not NOT1 (N2201, N2197);
buf BUF1 (N2202, N2193);
nand NAND4 (N2203, N2202, N953, N682, N1321);
nor NOR3 (N2204, N2194, N496, N915);
nor NOR4 (N2205, N2199, N1273, N1530, N1027);
and AND3 (N2206, N2204, N1960, N1886);
xor XOR2 (N2207, N2187, N1554);
xor XOR2 (N2208, N2205, N122);
xor XOR2 (N2209, N2203, N32);
xor XOR2 (N2210, N2198, N1611);
or OR3 (N2211, N2210, N2029, N119);
nor NOR3 (N2212, N2211, N1375, N1384);
nand NAND4 (N2213, N2206, N464, N1011, N498);
xor XOR2 (N2214, N2188, N532);
nor NOR2 (N2215, N2213, N2121);
xor XOR2 (N2216, N2214, N223);
and AND4 (N2217, N2195, N1443, N2105, N886);
nand NAND3 (N2218, N2162, N1931, N802);
buf BUF1 (N2219, N2216);
not NOT1 (N2220, N2208);
and AND2 (N2221, N2201, N1438);
nor NOR2 (N2222, N2221, N754);
nor NOR2 (N2223, N2217, N1826);
buf BUF1 (N2224, N2200);
nand NAND3 (N2225, N2224, N315, N54);
or OR3 (N2226, N2225, N601, N804);
nand NAND4 (N2227, N2222, N916, N1726, N1666);
or OR4 (N2228, N2220, N1733, N45, N490);
nand NAND2 (N2229, N2218, N1459);
buf BUF1 (N2230, N2228);
buf BUF1 (N2231, N2230);
or OR4 (N2232, N2212, N2168, N1581, N1032);
xor XOR2 (N2233, N2229, N560);
xor XOR2 (N2234, N2233, N1667);
not NOT1 (N2235, N2227);
nor NOR2 (N2236, N2223, N632);
nor NOR2 (N2237, N2219, N593);
and AND2 (N2238, N2234, N155);
nor NOR4 (N2239, N2215, N324, N1887, N2049);
not NOT1 (N2240, N2226);
buf BUF1 (N2241, N2231);
not NOT1 (N2242, N2232);
and AND2 (N2243, N2242, N489);
xor XOR2 (N2244, N2207, N960);
nand NAND2 (N2245, N2239, N1268);
nor NOR3 (N2246, N2244, N909, N1172);
nand NAND2 (N2247, N2243, N929);
nor NOR4 (N2248, N2237, N1273, N1732, N2037);
and AND2 (N2249, N2246, N14);
xor XOR2 (N2250, N2247, N1977);
nor NOR4 (N2251, N2248, N841, N2091, N1866);
not NOT1 (N2252, N2235);
xor XOR2 (N2253, N2240, N358);
and AND4 (N2254, N2209, N1126, N1788, N170);
buf BUF1 (N2255, N2254);
not NOT1 (N2256, N2253);
and AND3 (N2257, N2245, N1150, N1218);
buf BUF1 (N2258, N2241);
not NOT1 (N2259, N2255);
buf BUF1 (N2260, N2249);
nor NOR2 (N2261, N2250, N2249);
and AND2 (N2262, N2261, N2021);
and AND3 (N2263, N2259, N780, N929);
and AND4 (N2264, N2260, N1332, N628, N2216);
nand NAND4 (N2265, N2264, N1708, N2014, N1167);
buf BUF1 (N2266, N2256);
not NOT1 (N2267, N2266);
nand NAND3 (N2268, N2251, N1970, N214);
or OR4 (N2269, N2265, N1232, N817, N973);
nor NOR3 (N2270, N2252, N524, N2128);
xor XOR2 (N2271, N2268, N1705);
nand NAND4 (N2272, N2238, N173, N920, N1445);
nand NAND2 (N2273, N2272, N303);
and AND3 (N2274, N2262, N1570, N1372);
buf BUF1 (N2275, N2273);
and AND2 (N2276, N2258, N474);
nand NAND3 (N2277, N2270, N201, N1125);
buf BUF1 (N2278, N2257);
and AND2 (N2279, N2274, N117);
not NOT1 (N2280, N2271);
not NOT1 (N2281, N2277);
nor NOR3 (N2282, N2263, N1608, N1819);
nand NAND2 (N2283, N2279, N1640);
or OR4 (N2284, N2282, N1079, N2071, N2105);
nand NAND2 (N2285, N2236, N379);
buf BUF1 (N2286, N2267);
not NOT1 (N2287, N2278);
not NOT1 (N2288, N2283);
nand NAND4 (N2289, N2286, N1493, N2075, N1994);
xor XOR2 (N2290, N2289, N1391);
not NOT1 (N2291, N2290);
or OR4 (N2292, N2269, N1606, N990, N1282);
and AND3 (N2293, N2284, N2129, N1427);
nand NAND3 (N2294, N2276, N2192, N1515);
nand NAND2 (N2295, N2285, N1);
nor NOR3 (N2296, N2295, N1061, N1196);
not NOT1 (N2297, N2292);
xor XOR2 (N2298, N2280, N1575);
and AND2 (N2299, N2288, N584);
nand NAND2 (N2300, N2296, N596);
or OR3 (N2301, N2299, N534, N628);
xor XOR2 (N2302, N2281, N1165);
buf BUF1 (N2303, N2298);
nor NOR3 (N2304, N2294, N2090, N1462);
not NOT1 (N2305, N2275);
nand NAND3 (N2306, N2302, N2018, N2167);
and AND3 (N2307, N2287, N512, N322);
and AND4 (N2308, N2306, N651, N1286, N1224);
not NOT1 (N2309, N2308);
not NOT1 (N2310, N2309);
not NOT1 (N2311, N2300);
xor XOR2 (N2312, N2304, N441);
xor XOR2 (N2313, N2293, N646);
or OR2 (N2314, N2303, N206);
nor NOR3 (N2315, N2301, N1929, N56);
and AND3 (N2316, N2291, N269, N1762);
buf BUF1 (N2317, N2297);
xor XOR2 (N2318, N2310, N1471);
not NOT1 (N2319, N2318);
nor NOR3 (N2320, N2311, N1877, N1539);
buf BUF1 (N2321, N2307);
xor XOR2 (N2322, N2313, N1744);
not NOT1 (N2323, N2316);
xor XOR2 (N2324, N2319, N884);
nand NAND3 (N2325, N2320, N550, N1454);
or OR3 (N2326, N2321, N110, N2300);
xor XOR2 (N2327, N2326, N1514);
nor NOR3 (N2328, N2305, N1583, N1420);
xor XOR2 (N2329, N2312, N188);
buf BUF1 (N2330, N2324);
nor NOR3 (N2331, N2317, N1082, N367);
and AND4 (N2332, N2329, N841, N692, N99);
and AND2 (N2333, N2314, N1163);
xor XOR2 (N2334, N2323, N1809);
and AND2 (N2335, N2328, N2087);
or OR4 (N2336, N2325, N1171, N2132, N512);
nand NAND4 (N2337, N2330, N2057, N2101, N1832);
buf BUF1 (N2338, N2334);
not NOT1 (N2339, N2322);
buf BUF1 (N2340, N2335);
and AND3 (N2341, N2315, N596, N1903);
not NOT1 (N2342, N2338);
not NOT1 (N2343, N2340);
nor NOR4 (N2344, N2336, N733, N1223, N1374);
xor XOR2 (N2345, N2341, N1751);
nor NOR4 (N2346, N2344, N1113, N961, N1161);
xor XOR2 (N2347, N2346, N397);
nand NAND3 (N2348, N2332, N1352, N1907);
or OR4 (N2349, N2339, N1231, N32, N1283);
buf BUF1 (N2350, N2345);
or OR2 (N2351, N2337, N259);
xor XOR2 (N2352, N2343, N1070);
nand NAND2 (N2353, N2327, N498);
and AND3 (N2354, N2351, N137, N875);
buf BUF1 (N2355, N2349);
nor NOR3 (N2356, N2352, N1741, N1795);
and AND4 (N2357, N2348, N1792, N2203, N817);
and AND3 (N2358, N2354, N2159, N1156);
nand NAND4 (N2359, N2333, N470, N490, N1100);
buf BUF1 (N2360, N2353);
nor NOR2 (N2361, N2350, N343);
and AND3 (N2362, N2358, N1021, N1055);
or OR2 (N2363, N2361, N2038);
buf BUF1 (N2364, N2359);
and AND2 (N2365, N2342, N1878);
nand NAND3 (N2366, N2355, N1794, N2309);
nand NAND2 (N2367, N2331, N773);
nor NOR4 (N2368, N2357, N470, N1803, N505);
xor XOR2 (N2369, N2356, N1265);
buf BUF1 (N2370, N2369);
xor XOR2 (N2371, N2364, N1926);
not NOT1 (N2372, N2360);
buf BUF1 (N2373, N2372);
nand NAND4 (N2374, N2371, N95, N727, N1382);
nor NOR2 (N2375, N2374, N1405);
or OR3 (N2376, N2362, N425, N1634);
or OR3 (N2377, N2366, N1783, N1520);
not NOT1 (N2378, N2377);
nand NAND3 (N2379, N2365, N1654, N588);
xor XOR2 (N2380, N2370, N762);
or OR3 (N2381, N2347, N1631, N2345);
or OR2 (N2382, N2378, N261);
and AND3 (N2383, N2381, N1258, N705);
not NOT1 (N2384, N2380);
nand NAND2 (N2385, N2368, N1376);
buf BUF1 (N2386, N2375);
buf BUF1 (N2387, N2367);
nand NAND3 (N2388, N2376, N602, N695);
not NOT1 (N2389, N2379);
xor XOR2 (N2390, N2373, N1952);
xor XOR2 (N2391, N2389, N744);
xor XOR2 (N2392, N2391, N1693);
nand NAND4 (N2393, N2382, N1958, N36, N307);
not NOT1 (N2394, N2393);
nor NOR3 (N2395, N2394, N198, N2201);
not NOT1 (N2396, N2387);
not NOT1 (N2397, N2392);
not NOT1 (N2398, N2363);
xor XOR2 (N2399, N2383, N2004);
nor NOR2 (N2400, N2385, N937);
not NOT1 (N2401, N2396);
buf BUF1 (N2402, N2401);
not NOT1 (N2403, N2390);
nand NAND4 (N2404, N2397, N986, N2120, N876);
and AND2 (N2405, N2388, N1902);
not NOT1 (N2406, N2404);
xor XOR2 (N2407, N2386, N1618);
nor NOR2 (N2408, N2402, N1768);
not NOT1 (N2409, N2395);
not NOT1 (N2410, N2406);
or OR2 (N2411, N2384, N559);
nand NAND3 (N2412, N2400, N2284, N178);
nor NOR2 (N2413, N2408, N377);
not NOT1 (N2414, N2399);
or OR4 (N2415, N2405, N179, N1726, N2145);
nand NAND3 (N2416, N2410, N1257, N306);
or OR4 (N2417, N2416, N123, N2001, N1309);
not NOT1 (N2418, N2398);
or OR4 (N2419, N2413, N85, N1215, N1134);
nor NOR2 (N2420, N2418, N1611);
or OR4 (N2421, N2403, N431, N1771, N574);
buf BUF1 (N2422, N2421);
nand NAND2 (N2423, N2420, N1428);
nor NOR3 (N2424, N2414, N1520, N2271);
nand NAND2 (N2425, N2415, N1562);
nor NOR2 (N2426, N2419, N1377);
nor NOR3 (N2427, N2407, N2199, N1924);
not NOT1 (N2428, N2409);
not NOT1 (N2429, N2427);
or OR2 (N2430, N2429, N1538);
and AND2 (N2431, N2425, N1174);
and AND3 (N2432, N2423, N1981, N56);
buf BUF1 (N2433, N2428);
nor NOR2 (N2434, N2432, N156);
xor XOR2 (N2435, N2430, N435);
xor XOR2 (N2436, N2411, N1192);
nor NOR2 (N2437, N2435, N631);
buf BUF1 (N2438, N2417);
buf BUF1 (N2439, N2438);
or OR2 (N2440, N2436, N939);
or OR2 (N2441, N2437, N1166);
not NOT1 (N2442, N2431);
and AND2 (N2443, N2440, N43);
not NOT1 (N2444, N2439);
nor NOR4 (N2445, N2444, N645, N219, N745);
and AND2 (N2446, N2441, N247);
nand NAND4 (N2447, N2412, N1418, N2340, N178);
buf BUF1 (N2448, N2445);
xor XOR2 (N2449, N2433, N1617);
nand NAND3 (N2450, N2434, N150, N603);
or OR3 (N2451, N2448, N2327, N2009);
or OR4 (N2452, N2451, N2277, N754, N712);
nand NAND2 (N2453, N2443, N92);
and AND2 (N2454, N2426, N1839);
nor NOR2 (N2455, N2452, N455);
not NOT1 (N2456, N2422);
xor XOR2 (N2457, N2450, N1749);
or OR2 (N2458, N2442, N1793);
and AND2 (N2459, N2424, N1403);
or OR3 (N2460, N2457, N2357, N1243);
buf BUF1 (N2461, N2447);
or OR2 (N2462, N2454, N464);
or OR2 (N2463, N2460, N1980);
xor XOR2 (N2464, N2453, N114);
not NOT1 (N2465, N2462);
not NOT1 (N2466, N2464);
buf BUF1 (N2467, N2463);
or OR2 (N2468, N2449, N1344);
nand NAND2 (N2469, N2446, N1104);
and AND4 (N2470, N2466, N617, N2450, N858);
xor XOR2 (N2471, N2470, N1919);
and AND4 (N2472, N2467, N1056, N244, N192);
buf BUF1 (N2473, N2459);
not NOT1 (N2474, N2469);
nor NOR2 (N2475, N2472, N1441);
or OR4 (N2476, N2465, N2468, N1268, N1725);
nor NOR3 (N2477, N2351, N1541, N974);
buf BUF1 (N2478, N2475);
nand NAND4 (N2479, N2474, N367, N1361, N962);
buf BUF1 (N2480, N2476);
not NOT1 (N2481, N2455);
buf BUF1 (N2482, N2461);
buf BUF1 (N2483, N2480);
and AND3 (N2484, N2481, N2042, N1568);
buf BUF1 (N2485, N2478);
or OR2 (N2486, N2485, N1064);
or OR2 (N2487, N2456, N1563);
xor XOR2 (N2488, N2483, N505);
or OR4 (N2489, N2486, N1515, N2416, N301);
not NOT1 (N2490, N2484);
or OR3 (N2491, N2479, N1006, N126);
nand NAND3 (N2492, N2482, N2184, N1558);
not NOT1 (N2493, N2489);
not NOT1 (N2494, N2491);
nor NOR2 (N2495, N2493, N301);
nand NAND4 (N2496, N2471, N1420, N211, N163);
or OR4 (N2497, N2492, N438, N951, N1037);
xor XOR2 (N2498, N2487, N1448);
not NOT1 (N2499, N2495);
not NOT1 (N2500, N2490);
and AND3 (N2501, N2473, N1040, N2136);
not NOT1 (N2502, N2501);
nor NOR2 (N2503, N2496, N1739);
nor NOR3 (N2504, N2500, N790, N856);
nor NOR4 (N2505, N2488, N2447, N1616, N2060);
xor XOR2 (N2506, N2504, N1463);
buf BUF1 (N2507, N2497);
nor NOR4 (N2508, N2502, N2182, N171, N554);
not NOT1 (N2509, N2507);
xor XOR2 (N2510, N2506, N2286);
xor XOR2 (N2511, N2499, N78);
nand NAND4 (N2512, N2508, N2444, N322, N962);
and AND4 (N2513, N2477, N2381, N1775, N49);
and AND4 (N2514, N2505, N1345, N2103, N253);
nor NOR4 (N2515, N2513, N2238, N1015, N1933);
and AND4 (N2516, N2510, N1929, N1536, N1147);
nor NOR4 (N2517, N2511, N157, N2172, N1985);
and AND3 (N2518, N2458, N1390, N2233);
nand NAND3 (N2519, N2515, N2025, N1125);
buf BUF1 (N2520, N2517);
nand NAND4 (N2521, N2516, N1738, N1724, N2180);
not NOT1 (N2522, N2503);
and AND4 (N2523, N2498, N2306, N1417, N2221);
nor NOR3 (N2524, N2520, N1546, N1866);
and AND4 (N2525, N2523, N1058, N1440, N714);
nand NAND3 (N2526, N2524, N7, N1633);
nand NAND4 (N2527, N2519, N2326, N1820, N1202);
buf BUF1 (N2528, N2509);
not NOT1 (N2529, N2526);
and AND2 (N2530, N2512, N817);
or OR4 (N2531, N2525, N712, N1244, N1517);
nand NAND4 (N2532, N2531, N206, N607, N1829);
or OR4 (N2533, N2514, N2392, N1147, N1127);
nand NAND2 (N2534, N2532, N1204);
not NOT1 (N2535, N2522);
not NOT1 (N2536, N2527);
nand NAND3 (N2537, N2528, N2269, N27);
xor XOR2 (N2538, N2529, N78);
nor NOR3 (N2539, N2521, N504, N78);
or OR2 (N2540, N2536, N125);
xor XOR2 (N2541, N2494, N330);
xor XOR2 (N2542, N2537, N512);
xor XOR2 (N2543, N2530, N1939);
nor NOR3 (N2544, N2539, N1564, N1073);
buf BUF1 (N2545, N2541);
buf BUF1 (N2546, N2543);
nor NOR3 (N2547, N2518, N1063, N1888);
nand NAND4 (N2548, N2546, N174, N747, N1726);
xor XOR2 (N2549, N2540, N1709);
or OR4 (N2550, N2535, N698, N1500, N2021);
and AND4 (N2551, N2533, N1482, N2261, N2507);
buf BUF1 (N2552, N2545);
or OR2 (N2553, N2534, N887);
and AND4 (N2554, N2552, N1008, N949, N403);
not NOT1 (N2555, N2538);
nand NAND4 (N2556, N2549, N480, N331, N1879);
nand NAND4 (N2557, N2551, N173, N2422, N1384);
or OR3 (N2558, N2553, N1855, N1675);
and AND4 (N2559, N2550, N1896, N2398, N2004);
xor XOR2 (N2560, N2544, N830);
nand NAND4 (N2561, N2548, N1358, N1118, N942);
buf BUF1 (N2562, N2554);
and AND3 (N2563, N2562, N2250, N758);
nand NAND2 (N2564, N2561, N520);
nor NOR2 (N2565, N2555, N129);
nand NAND4 (N2566, N2563, N1458, N499, N1699);
nand NAND4 (N2567, N2560, N358, N684, N859);
and AND2 (N2568, N2557, N2114);
nor NOR2 (N2569, N2547, N219);
buf BUF1 (N2570, N2566);
not NOT1 (N2571, N2556);
or OR2 (N2572, N2558, N1843);
or OR3 (N2573, N2572, N987, N1789);
nor NOR2 (N2574, N2568, N2329);
buf BUF1 (N2575, N2542);
buf BUF1 (N2576, N2565);
and AND3 (N2577, N2575, N940, N777);
buf BUF1 (N2578, N2567);
xor XOR2 (N2579, N2564, N365);
xor XOR2 (N2580, N2571, N517);
buf BUF1 (N2581, N2570);
nand NAND2 (N2582, N2581, N1873);
nand NAND3 (N2583, N2559, N1162, N2123);
and AND4 (N2584, N2574, N2029, N683, N1941);
nand NAND4 (N2585, N2576, N1826, N163, N2252);
xor XOR2 (N2586, N2583, N1197);
nand NAND3 (N2587, N2579, N2066, N762);
xor XOR2 (N2588, N2569, N2100);
buf BUF1 (N2589, N2578);
xor XOR2 (N2590, N2585, N2494);
buf BUF1 (N2591, N2586);
or OR2 (N2592, N2580, N733);
nor NOR2 (N2593, N2573, N187);
nor NOR3 (N2594, N2587, N978, N443);
and AND4 (N2595, N2594, N1078, N2020, N693);
nand NAND2 (N2596, N2593, N351);
and AND3 (N2597, N2590, N821, N2229);
and AND4 (N2598, N2597, N1473, N149, N1683);
xor XOR2 (N2599, N2591, N169);
and AND3 (N2600, N2592, N401, N2444);
buf BUF1 (N2601, N2582);
or OR3 (N2602, N2595, N476, N1304);
buf BUF1 (N2603, N2600);
nor NOR2 (N2604, N2577, N1616);
and AND3 (N2605, N2602, N1587, N1715);
buf BUF1 (N2606, N2603);
buf BUF1 (N2607, N2601);
nor NOR2 (N2608, N2598, N816);
or OR2 (N2609, N2605, N1712);
not NOT1 (N2610, N2604);
nor NOR4 (N2611, N2584, N459, N2423, N2490);
buf BUF1 (N2612, N2607);
xor XOR2 (N2613, N2610, N560);
and AND3 (N2614, N2613, N156, N1065);
nand NAND2 (N2615, N2588, N2337);
not NOT1 (N2616, N2612);
and AND4 (N2617, N2615, N2289, N2541, N1998);
not NOT1 (N2618, N2608);
nand NAND3 (N2619, N2606, N1591, N1729);
nand NAND4 (N2620, N2589, N1479, N819, N1870);
and AND4 (N2621, N2599, N294, N2595, N1428);
nor NOR4 (N2622, N2620, N581, N813, N834);
buf BUF1 (N2623, N2614);
buf BUF1 (N2624, N2621);
or OR3 (N2625, N2623, N183, N1945);
nor NOR2 (N2626, N2622, N2180);
nand NAND3 (N2627, N2611, N2588, N647);
xor XOR2 (N2628, N2609, N2596);
nand NAND4 (N2629, N856, N743, N2131, N34);
and AND4 (N2630, N2616, N2283, N474, N601);
buf BUF1 (N2631, N2630);
not NOT1 (N2632, N2628);
and AND2 (N2633, N2627, N1309);
and AND4 (N2634, N2617, N615, N1094, N2625);
not NOT1 (N2635, N2056);
xor XOR2 (N2636, N2629, N2453);
buf BUF1 (N2637, N2635);
nor NOR4 (N2638, N2632, N234, N262, N898);
not NOT1 (N2639, N2631);
nor NOR2 (N2640, N2626, N363);
nand NAND3 (N2641, N2637, N399, N416);
buf BUF1 (N2642, N2640);
and AND2 (N2643, N2618, N1046);
buf BUF1 (N2644, N2642);
not NOT1 (N2645, N2636);
xor XOR2 (N2646, N2624, N563);
nand NAND4 (N2647, N2619, N1805, N628, N302);
or OR4 (N2648, N2638, N2337, N2160, N1604);
buf BUF1 (N2649, N2645);
or OR2 (N2650, N2648, N1587);
buf BUF1 (N2651, N2643);
nand NAND2 (N2652, N2633, N6);
and AND3 (N2653, N2651, N503, N2328);
xor XOR2 (N2654, N2650, N1078);
nand NAND4 (N2655, N2646, N1336, N2140, N33);
nor NOR3 (N2656, N2653, N526, N553);
nand NAND2 (N2657, N2656, N1909);
and AND2 (N2658, N2644, N936);
buf BUF1 (N2659, N2639);
or OR3 (N2660, N2649, N451, N2036);
nor NOR3 (N2661, N2655, N270, N538);
nand NAND3 (N2662, N2641, N221, N943);
xor XOR2 (N2663, N2661, N1939);
or OR2 (N2664, N2634, N408);
buf BUF1 (N2665, N2654);
not NOT1 (N2666, N2647);
nand NAND4 (N2667, N2657, N207, N310, N864);
not NOT1 (N2668, N2664);
nand NAND3 (N2669, N2659, N2236, N2360);
not NOT1 (N2670, N2668);
buf BUF1 (N2671, N2667);
xor XOR2 (N2672, N2652, N2571);
nand NAND3 (N2673, N2662, N463, N257);
nor NOR2 (N2674, N2666, N1628);
not NOT1 (N2675, N2672);
or OR2 (N2676, N2673, N1633);
xor XOR2 (N2677, N2676, N2615);
not NOT1 (N2678, N2670);
buf BUF1 (N2679, N2658);
or OR4 (N2680, N2675, N1115, N1261, N2293);
buf BUF1 (N2681, N2680);
and AND4 (N2682, N2671, N313, N1241, N506);
or OR4 (N2683, N2663, N1873, N2088, N2285);
and AND3 (N2684, N2683, N1787, N1482);
nor NOR4 (N2685, N2684, N2328, N2517, N1451);
or OR4 (N2686, N2685, N565, N1246, N1946);
and AND3 (N2687, N2686, N788, N2128);
not NOT1 (N2688, N2682);
buf BUF1 (N2689, N2665);
not NOT1 (N2690, N2689);
and AND3 (N2691, N2687, N2589, N434);
nor NOR3 (N2692, N2669, N2478, N871);
xor XOR2 (N2693, N2688, N1513);
or OR2 (N2694, N2677, N901);
nor NOR4 (N2695, N2694, N573, N2192, N1266);
nand NAND4 (N2696, N2690, N2154, N437, N2623);
not NOT1 (N2697, N2660);
or OR2 (N2698, N2691, N2409);
xor XOR2 (N2699, N2679, N613);
nor NOR2 (N2700, N2695, N177);
and AND2 (N2701, N2699, N2014);
or OR2 (N2702, N2692, N978);
or OR3 (N2703, N2678, N2109, N2313);
buf BUF1 (N2704, N2703);
xor XOR2 (N2705, N2702, N2074);
xor XOR2 (N2706, N2696, N2045);
not NOT1 (N2707, N2700);
buf BUF1 (N2708, N2705);
nor NOR3 (N2709, N2697, N1933, N2288);
xor XOR2 (N2710, N2698, N866);
buf BUF1 (N2711, N2710);
or OR2 (N2712, N2681, N1842);
or OR4 (N2713, N2707, N1574, N228, N2138);
nor NOR3 (N2714, N2708, N57, N1012);
nor NOR3 (N2715, N2712, N406, N1167);
or OR2 (N2716, N2709, N1589);
xor XOR2 (N2717, N2711, N1747);
nor NOR2 (N2718, N2704, N522);
nor NOR4 (N2719, N2713, N77, N2292, N27);
buf BUF1 (N2720, N2693);
buf BUF1 (N2721, N2674);
nand NAND2 (N2722, N2716, N1902);
not NOT1 (N2723, N2706);
nand NAND3 (N2724, N2719, N2118, N1049);
not NOT1 (N2725, N2701);
nor NOR2 (N2726, N2714, N914);
nand NAND4 (N2727, N2725, N2098, N1158, N2407);
and AND3 (N2728, N2726, N2677, N1614);
and AND2 (N2729, N2715, N1093);
and AND3 (N2730, N2724, N149, N2305);
not NOT1 (N2731, N2727);
nand NAND4 (N2732, N2720, N2201, N1499, N2114);
not NOT1 (N2733, N2729);
or OR3 (N2734, N2732, N2722, N2102);
xor XOR2 (N2735, N526, N2085);
not NOT1 (N2736, N2730);
not NOT1 (N2737, N2723);
not NOT1 (N2738, N2728);
not NOT1 (N2739, N2721);
nand NAND2 (N2740, N2718, N325);
or OR3 (N2741, N2731, N1710, N311);
and AND4 (N2742, N2717, N2494, N365, N2628);
nor NOR4 (N2743, N2736, N2702, N1215, N1442);
not NOT1 (N2744, N2737);
xor XOR2 (N2745, N2739, N109);
and AND3 (N2746, N2744, N2261, N127);
and AND2 (N2747, N2746, N125);
nor NOR2 (N2748, N2740, N348);
nand NAND3 (N2749, N2733, N257, N983);
buf BUF1 (N2750, N2747);
and AND3 (N2751, N2749, N463, N1570);
buf BUF1 (N2752, N2734);
nor NOR2 (N2753, N2750, N664);
or OR3 (N2754, N2741, N1344, N2694);
nand NAND2 (N2755, N2753, N1030);
not NOT1 (N2756, N2743);
and AND2 (N2757, N2751, N2336);
nor NOR2 (N2758, N2745, N1464);
xor XOR2 (N2759, N2754, N1318);
not NOT1 (N2760, N2759);
nor NOR2 (N2761, N2742, N979);
nand NAND4 (N2762, N2735, N1551, N400, N2192);
nor NOR3 (N2763, N2761, N2366, N728);
buf BUF1 (N2764, N2738);
xor XOR2 (N2765, N2757, N1439);
xor XOR2 (N2766, N2758, N1232);
and AND2 (N2767, N2765, N2413);
xor XOR2 (N2768, N2748, N1453);
or OR3 (N2769, N2756, N599, N2097);
xor XOR2 (N2770, N2767, N1517);
or OR2 (N2771, N2762, N2209);
xor XOR2 (N2772, N2771, N488);
or OR4 (N2773, N2764, N379, N1582, N913);
or OR3 (N2774, N2770, N140, N214);
nor NOR4 (N2775, N2772, N1153, N126, N2511);
nand NAND3 (N2776, N2768, N1348, N1913);
xor XOR2 (N2777, N2773, N1671);
or OR4 (N2778, N2775, N2741, N1659, N2342);
and AND4 (N2779, N2752, N58, N2173, N612);
xor XOR2 (N2780, N2777, N846);
buf BUF1 (N2781, N2776);
nor NOR3 (N2782, N2769, N1579, N2759);
not NOT1 (N2783, N2763);
and AND4 (N2784, N2755, N1444, N1433, N2140);
buf BUF1 (N2785, N2782);
or OR4 (N2786, N2780, N1935, N994, N1945);
xor XOR2 (N2787, N2778, N1049);
and AND3 (N2788, N2785, N1948, N597);
xor XOR2 (N2789, N2784, N518);
and AND3 (N2790, N2783, N1806, N1639);
not NOT1 (N2791, N2788);
and AND2 (N2792, N2789, N820);
nor NOR3 (N2793, N2774, N956, N1766);
not NOT1 (N2794, N2779);
xor XOR2 (N2795, N2781, N2057);
nor NOR3 (N2796, N2795, N829, N1351);
nor NOR3 (N2797, N2790, N520, N1344);
nor NOR2 (N2798, N2792, N1067);
not NOT1 (N2799, N2791);
nand NAND4 (N2800, N2793, N1368, N172, N1038);
nor NOR2 (N2801, N2787, N558);
buf BUF1 (N2802, N2801);
buf BUF1 (N2803, N2760);
nor NOR4 (N2804, N2798, N1648, N555, N1444);
and AND2 (N2805, N2786, N604);
and AND4 (N2806, N2794, N652, N157, N2528);
nand NAND4 (N2807, N2796, N569, N988, N2143);
buf BUF1 (N2808, N2807);
nor NOR3 (N2809, N2803, N641, N346);
and AND3 (N2810, N2799, N2031, N280);
buf BUF1 (N2811, N2766);
or OR2 (N2812, N2810, N329);
not NOT1 (N2813, N2797);
nor NOR3 (N2814, N2813, N2693, N2188);
not NOT1 (N2815, N2811);
or OR3 (N2816, N2802, N2360, N2298);
nand NAND4 (N2817, N2808, N1085, N174, N590);
nand NAND4 (N2818, N2816, N824, N1211, N1370);
nand NAND3 (N2819, N2814, N194, N2061);
nand NAND2 (N2820, N2805, N675);
nor NOR4 (N2821, N2819, N1864, N501, N2218);
nor NOR2 (N2822, N2821, N2437);
nor NOR3 (N2823, N2822, N2069, N1897);
or OR4 (N2824, N2809, N2097, N1264, N405);
buf BUF1 (N2825, N2800);
nor NOR2 (N2826, N2806, N1893);
buf BUF1 (N2827, N2826);
and AND2 (N2828, N2804, N1283);
xor XOR2 (N2829, N2828, N2426);
and AND3 (N2830, N2827, N1148, N815);
nor NOR4 (N2831, N2830, N23, N1943, N2611);
and AND4 (N2832, N2831, N37, N2795, N2322);
xor XOR2 (N2833, N2829, N387);
nand NAND4 (N2834, N2815, N1752, N2215, N87);
nor NOR3 (N2835, N2825, N1032, N2826);
nor NOR3 (N2836, N2835, N2762, N1288);
xor XOR2 (N2837, N2833, N2624);
or OR2 (N2838, N2832, N2262);
nand NAND4 (N2839, N2820, N518, N2190, N2456);
not NOT1 (N2840, N2838);
nor NOR4 (N2841, N2834, N183, N1257, N2374);
xor XOR2 (N2842, N2836, N1175);
not NOT1 (N2843, N2817);
or OR3 (N2844, N2842, N1929, N1839);
xor XOR2 (N2845, N2840, N1963);
nor NOR4 (N2846, N2839, N2109, N950, N2118);
nand NAND3 (N2847, N2823, N2055, N1446);
nor NOR3 (N2848, N2818, N1412, N1769);
buf BUF1 (N2849, N2837);
xor XOR2 (N2850, N2812, N262);
not NOT1 (N2851, N2849);
not NOT1 (N2852, N2851);
or OR2 (N2853, N2850, N2248);
or OR3 (N2854, N2852, N206, N445);
or OR3 (N2855, N2824, N270, N1538);
xor XOR2 (N2856, N2843, N350);
nor NOR2 (N2857, N2853, N450);
not NOT1 (N2858, N2844);
nor NOR2 (N2859, N2854, N2508);
xor XOR2 (N2860, N2855, N359);
nor NOR3 (N2861, N2848, N1908, N281);
not NOT1 (N2862, N2847);
and AND3 (N2863, N2861, N2414, N1749);
nor NOR4 (N2864, N2858, N952, N2214, N2257);
xor XOR2 (N2865, N2864, N225);
nor NOR4 (N2866, N2862, N1711, N1267, N2641);
or OR4 (N2867, N2865, N848, N1747, N985);
nor NOR2 (N2868, N2856, N2527);
or OR2 (N2869, N2841, N1897);
not NOT1 (N2870, N2868);
or OR3 (N2871, N2859, N2606, N2166);
and AND4 (N2872, N2857, N2197, N1986, N2026);
nand NAND2 (N2873, N2870, N2131);
or OR3 (N2874, N2866, N1471, N890);
not NOT1 (N2875, N2869);
and AND2 (N2876, N2871, N2026);
buf BUF1 (N2877, N2875);
nor NOR2 (N2878, N2877, N807);
nand NAND3 (N2879, N2878, N2506, N2456);
or OR2 (N2880, N2860, N1970);
not NOT1 (N2881, N2880);
and AND2 (N2882, N2872, N76);
or OR2 (N2883, N2876, N2333);
nand NAND4 (N2884, N2863, N1903, N77, N1793);
or OR2 (N2885, N2882, N1113);
and AND3 (N2886, N2885, N80, N166);
buf BUF1 (N2887, N2884);
nor NOR3 (N2888, N2887, N261, N2543);
or OR2 (N2889, N2881, N712);
not NOT1 (N2890, N2883);
and AND4 (N2891, N2845, N1584, N459, N1277);
buf BUF1 (N2892, N2888);
xor XOR2 (N2893, N2873, N2386);
or OR2 (N2894, N2867, N1057);
or OR4 (N2895, N2894, N1243, N2728, N501);
xor XOR2 (N2896, N2893, N1013);
nand NAND3 (N2897, N2889, N792, N1215);
nand NAND4 (N2898, N2895, N1066, N1437, N1620);
xor XOR2 (N2899, N2896, N2753);
xor XOR2 (N2900, N2898, N1917);
nand NAND3 (N2901, N2892, N97, N800);
not NOT1 (N2902, N2901);
buf BUF1 (N2903, N2879);
nor NOR2 (N2904, N2900, N1904);
not NOT1 (N2905, N2891);
nor NOR4 (N2906, N2886, N2336, N2394, N1416);
buf BUF1 (N2907, N2902);
or OR2 (N2908, N2899, N1847);
nor NOR2 (N2909, N2890, N2901);
or OR4 (N2910, N2909, N2875, N2195, N1324);
and AND2 (N2911, N2908, N1806);
buf BUF1 (N2912, N2910);
not NOT1 (N2913, N2905);
or OR3 (N2914, N2912, N239, N410);
buf BUF1 (N2915, N2874);
nand NAND2 (N2916, N2911, N2372);
not NOT1 (N2917, N2916);
not NOT1 (N2918, N2914);
and AND2 (N2919, N2917, N2868);
buf BUF1 (N2920, N2897);
nor NOR4 (N2921, N2904, N2315, N1349, N1020);
nand NAND2 (N2922, N2906, N442);
xor XOR2 (N2923, N2846, N616);
nand NAND2 (N2924, N2919, N892);
xor XOR2 (N2925, N2913, N435);
nand NAND2 (N2926, N2923, N399);
nand NAND2 (N2927, N2924, N1712);
buf BUF1 (N2928, N2927);
and AND2 (N2929, N2918, N1379);
and AND2 (N2930, N2928, N1742);
buf BUF1 (N2931, N2907);
buf BUF1 (N2932, N2922);
or OR3 (N2933, N2932, N669, N640);
not NOT1 (N2934, N2920);
or OR3 (N2935, N2921, N823, N1439);
xor XOR2 (N2936, N2925, N1152);
and AND4 (N2937, N2936, N1616, N2477, N2028);
nor NOR3 (N2938, N2937, N2534, N115);
nor NOR3 (N2939, N2931, N1583, N2568);
nor NOR2 (N2940, N2915, N2376);
buf BUF1 (N2941, N2930);
and AND3 (N2942, N2939, N1931, N1589);
not NOT1 (N2943, N2942);
buf BUF1 (N2944, N2933);
not NOT1 (N2945, N2941);
nand NAND2 (N2946, N2926, N2664);
and AND3 (N2947, N2938, N609, N2385);
buf BUF1 (N2948, N2935);
buf BUF1 (N2949, N2940);
not NOT1 (N2950, N2948);
xor XOR2 (N2951, N2929, N413);
not NOT1 (N2952, N2945);
not NOT1 (N2953, N2952);
xor XOR2 (N2954, N2944, N2217);
not NOT1 (N2955, N2934);
and AND3 (N2956, N2946, N2415, N1632);
nand NAND3 (N2957, N2943, N796, N240);
and AND4 (N2958, N2957, N422, N1194, N198);
xor XOR2 (N2959, N2949, N2246);
and AND3 (N2960, N2903, N965, N2141);
not NOT1 (N2961, N2951);
buf BUF1 (N2962, N2956);
xor XOR2 (N2963, N2955, N286);
buf BUF1 (N2964, N2963);
or OR3 (N2965, N2954, N509, N161);
nand NAND3 (N2966, N2959, N1805, N2411);
or OR3 (N2967, N2962, N1535, N1430);
not NOT1 (N2968, N2966);
nor NOR2 (N2969, N2968, N620);
nand NAND3 (N2970, N2960, N2122, N2285);
not NOT1 (N2971, N2953);
buf BUF1 (N2972, N2965);
or OR3 (N2973, N2971, N1315, N2195);
and AND2 (N2974, N2964, N2874);
xor XOR2 (N2975, N2967, N1651);
and AND3 (N2976, N2974, N2872, N1581);
nand NAND4 (N2977, N2969, N1264, N1965, N2013);
and AND4 (N2978, N2970, N1393, N2051, N501);
and AND2 (N2979, N2958, N1613);
xor XOR2 (N2980, N2977, N1401);
not NOT1 (N2981, N2950);
xor XOR2 (N2982, N2978, N166);
and AND4 (N2983, N2961, N1604, N2268, N122);
not NOT1 (N2984, N2981);
xor XOR2 (N2985, N2983, N1814);
xor XOR2 (N2986, N2984, N778);
and AND2 (N2987, N2975, N1199);
or OR3 (N2988, N2980, N2101, N2047);
nand NAND3 (N2989, N2985, N2752, N2149);
not NOT1 (N2990, N2986);
or OR3 (N2991, N2947, N1235, N376);
and AND2 (N2992, N2972, N1298);
not NOT1 (N2993, N2988);
nor NOR3 (N2994, N2989, N392, N789);
not NOT1 (N2995, N2991);
buf BUF1 (N2996, N2990);
and AND2 (N2997, N2993, N1925);
buf BUF1 (N2998, N2992);
xor XOR2 (N2999, N2987, N1366);
buf BUF1 (N3000, N2998);
or OR3 (N3001, N2994, N669, N2054);
nor NOR2 (N3002, N2997, N2590);
nor NOR3 (N3003, N3000, N1247, N1309);
nand NAND3 (N3004, N3003, N961, N55);
and AND2 (N3005, N2996, N2870);
xor XOR2 (N3006, N3004, N436);
buf BUF1 (N3007, N2973);
nand NAND4 (N3008, N2982, N1200, N1210, N900);
and AND3 (N3009, N3007, N2259, N33);
nor NOR2 (N3010, N3005, N2196);
xor XOR2 (N3011, N3002, N2276);
or OR4 (N3012, N3008, N1352, N557, N1439);
buf BUF1 (N3013, N3012);
and AND4 (N3014, N3013, N926, N1905, N969);
not NOT1 (N3015, N3006);
xor XOR2 (N3016, N2976, N1285);
not NOT1 (N3017, N3009);
and AND2 (N3018, N2979, N1749);
nand NAND4 (N3019, N3015, N1528, N1074, N450);
nor NOR2 (N3020, N3019, N900);
not NOT1 (N3021, N3010);
xor XOR2 (N3022, N3021, N2856);
endmodule