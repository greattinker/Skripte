// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N2006,N2013,N2011,N2016,N1992,N2017,N1998,N2002,N2015,N2018;

nor NOR4 (N19, N12, N4, N1, N16);
nor NOR3 (N20, N9, N15, N12);
buf BUF1 (N21, N12);
xor XOR2 (N22, N16, N4);
or OR3 (N23, N19, N16, N11);
or OR3 (N24, N6, N2, N18);
buf BUF1 (N25, N13);
xor XOR2 (N26, N24, N3);
nor NOR3 (N27, N6, N3, N25);
buf BUF1 (N28, N25);
nand NAND3 (N29, N25, N2, N18);
not NOT1 (N30, N1);
buf BUF1 (N31, N26);
and AND4 (N32, N14, N13, N26, N18);
or OR2 (N33, N28, N3);
buf BUF1 (N34, N30);
nor NOR3 (N35, N20, N6, N19);
xor XOR2 (N36, N27, N25);
buf BUF1 (N37, N35);
nor NOR4 (N38, N29, N14, N27, N12);
and AND2 (N39, N37, N12);
nand NAND3 (N40, N21, N13, N14);
and AND3 (N41, N33, N16, N14);
and AND2 (N42, N34, N26);
or OR3 (N43, N41, N21, N23);
not NOT1 (N44, N43);
and AND3 (N45, N4, N31, N24);
not NOT1 (N46, N2);
xor XOR2 (N47, N46, N14);
not NOT1 (N48, N39);
or OR3 (N49, N42, N20, N34);
buf BUF1 (N50, N36);
not NOT1 (N51, N50);
and AND3 (N52, N40, N13, N51);
and AND2 (N53, N49, N21);
nand NAND2 (N54, N34, N53);
not NOT1 (N55, N36);
or OR2 (N56, N22, N5);
buf BUF1 (N57, N32);
nand NAND3 (N58, N57, N57, N17);
or OR4 (N59, N48, N57, N32, N39);
not NOT1 (N60, N59);
or OR2 (N61, N55, N45);
xor XOR2 (N62, N19, N15);
nor NOR4 (N63, N38, N5, N41, N40);
nand NAND2 (N64, N44, N49);
xor XOR2 (N65, N58, N33);
and AND2 (N66, N47, N46);
or OR4 (N67, N56, N38, N53, N8);
buf BUF1 (N68, N64);
not NOT1 (N69, N67);
xor XOR2 (N70, N60, N69);
and AND3 (N71, N38, N66, N42);
or OR2 (N72, N27, N15);
nor NOR4 (N73, N54, N2, N30, N50);
xor XOR2 (N74, N73, N11);
nand NAND3 (N75, N62, N52, N40);
not NOT1 (N76, N28);
xor XOR2 (N77, N61, N63);
and AND3 (N78, N48, N23, N31);
nor NOR3 (N79, N65, N39, N10);
xor XOR2 (N80, N74, N33);
or OR4 (N81, N77, N77, N13, N6);
or OR2 (N82, N75, N20);
nor NOR3 (N83, N76, N63, N9);
xor XOR2 (N84, N83, N6);
nor NOR4 (N85, N78, N23, N16, N23);
not NOT1 (N86, N81);
nand NAND2 (N87, N82, N11);
or OR3 (N88, N86, N46, N65);
nand NAND4 (N89, N80, N39, N63, N22);
xor XOR2 (N90, N84, N88);
buf BUF1 (N91, N9);
not NOT1 (N92, N91);
nand NAND4 (N93, N71, N10, N65, N34);
and AND2 (N94, N87, N87);
and AND4 (N95, N93, N39, N70, N84);
nand NAND2 (N96, N67, N95);
nor NOR4 (N97, N86, N47, N35, N65);
buf BUF1 (N98, N89);
nor NOR4 (N99, N97, N47, N64, N42);
nor NOR3 (N100, N92, N83, N3);
not NOT1 (N101, N99);
not NOT1 (N102, N96);
or OR3 (N103, N72, N34, N38);
or OR4 (N104, N102, N76, N77, N94);
and AND4 (N105, N5, N61, N98, N12);
nor NOR2 (N106, N74, N35);
not NOT1 (N107, N103);
nor NOR2 (N108, N105, N94);
nand NAND3 (N109, N68, N96, N107);
nand NAND2 (N110, N84, N107);
nand NAND2 (N111, N104, N53);
buf BUF1 (N112, N108);
or OR2 (N113, N110, N48);
nand NAND3 (N114, N100, N12, N46);
buf BUF1 (N115, N112);
nor NOR3 (N116, N113, N103, N92);
and AND3 (N117, N101, N78, N28);
or OR3 (N118, N90, N20, N104);
not NOT1 (N119, N118);
and AND4 (N120, N119, N45, N62, N114);
not NOT1 (N121, N116);
buf BUF1 (N122, N81);
and AND2 (N123, N109, N5);
not NOT1 (N124, N120);
buf BUF1 (N125, N123);
buf BUF1 (N126, N125);
buf BUF1 (N127, N122);
and AND3 (N128, N126, N37, N127);
nand NAND2 (N129, N107, N115);
or OR2 (N130, N70, N28);
xor XOR2 (N131, N128, N25);
buf BUF1 (N132, N111);
not NOT1 (N133, N79);
not NOT1 (N134, N106);
xor XOR2 (N135, N132, N96);
xor XOR2 (N136, N133, N48);
or OR3 (N137, N85, N49, N94);
buf BUF1 (N138, N130);
not NOT1 (N139, N138);
nand NAND2 (N140, N134, N130);
nand NAND4 (N141, N139, N4, N80, N57);
or OR3 (N142, N140, N1, N86);
xor XOR2 (N143, N142, N20);
not NOT1 (N144, N131);
buf BUF1 (N145, N136);
nand NAND3 (N146, N145, N124, N133);
buf BUF1 (N147, N61);
xor XOR2 (N148, N146, N145);
and AND2 (N149, N129, N41);
nand NAND3 (N150, N143, N57, N16);
nor NOR2 (N151, N149, N149);
not NOT1 (N152, N117);
not NOT1 (N153, N147);
xor XOR2 (N154, N141, N80);
not NOT1 (N155, N151);
nor NOR3 (N156, N137, N25, N122);
and AND2 (N157, N148, N121);
not NOT1 (N158, N122);
not NOT1 (N159, N153);
xor XOR2 (N160, N159, N2);
buf BUF1 (N161, N150);
and AND3 (N162, N156, N2, N27);
xor XOR2 (N163, N157, N77);
or OR2 (N164, N161, N43);
not NOT1 (N165, N158);
and AND3 (N166, N162, N120, N140);
buf BUF1 (N167, N166);
not NOT1 (N168, N164);
or OR2 (N169, N163, N39);
nor NOR3 (N170, N152, N44, N61);
nor NOR2 (N171, N167, N47);
nor NOR2 (N172, N144, N102);
and AND2 (N173, N171, N134);
nor NOR3 (N174, N172, N37, N67);
and AND4 (N175, N154, N151, N149, N46);
buf BUF1 (N176, N170);
nand NAND3 (N177, N169, N158, N46);
buf BUF1 (N178, N177);
nor NOR2 (N179, N135, N174);
nand NAND3 (N180, N57, N172, N160);
xor XOR2 (N181, N94, N96);
buf BUF1 (N182, N178);
not NOT1 (N183, N181);
nand NAND2 (N184, N155, N5);
nand NAND4 (N185, N173, N32, N69, N35);
not NOT1 (N186, N180);
nor NOR2 (N187, N186, N133);
buf BUF1 (N188, N182);
or OR4 (N189, N165, N184, N41, N181);
or OR3 (N190, N52, N147, N11);
not NOT1 (N191, N179);
xor XOR2 (N192, N190, N127);
nand NAND3 (N193, N175, N42, N66);
not NOT1 (N194, N183);
nor NOR3 (N195, N193, N155, N70);
nand NAND3 (N196, N195, N156, N34);
xor XOR2 (N197, N168, N83);
or OR4 (N198, N189, N137, N70, N143);
or OR4 (N199, N187, N188, N131, N191);
and AND2 (N200, N109, N65);
or OR2 (N201, N148, N200);
and AND4 (N202, N85, N89, N176, N111);
not NOT1 (N203, N72);
and AND3 (N204, N185, N65, N35);
nand NAND4 (N205, N198, N187, N83, N165);
nor NOR2 (N206, N196, N116);
and AND3 (N207, N197, N43, N5);
nand NAND3 (N208, N194, N115, N173);
or OR2 (N209, N204, N205);
not NOT1 (N210, N165);
nor NOR3 (N211, N192, N82, N176);
xor XOR2 (N212, N206, N126);
or OR2 (N213, N208, N47);
and AND4 (N214, N199, N171, N179, N204);
and AND4 (N215, N213, N122, N142, N127);
or OR4 (N216, N212, N49, N29, N20);
and AND3 (N217, N209, N36, N178);
xor XOR2 (N218, N211, N51);
or OR2 (N219, N202, N193);
nand NAND4 (N220, N203, N125, N94, N38);
nand NAND2 (N221, N207, N45);
buf BUF1 (N222, N218);
xor XOR2 (N223, N201, N111);
nor NOR2 (N224, N216, N124);
nor NOR4 (N225, N215, N59, N153, N49);
not NOT1 (N226, N221);
xor XOR2 (N227, N219, N66);
and AND2 (N228, N214, N179);
and AND3 (N229, N224, N99, N223);
not NOT1 (N230, N167);
or OR4 (N231, N230, N150, N142, N116);
and AND2 (N232, N231, N180);
nand NAND4 (N233, N232, N130, N142, N29);
and AND4 (N234, N210, N89, N49, N64);
nor NOR2 (N235, N220, N164);
and AND2 (N236, N234, N227);
or OR2 (N237, N22, N85);
not NOT1 (N238, N226);
nor NOR3 (N239, N229, N84, N24);
nor NOR2 (N240, N217, N230);
and AND3 (N241, N238, N234, N115);
not NOT1 (N242, N240);
not NOT1 (N243, N222);
nor NOR2 (N244, N233, N64);
not NOT1 (N245, N225);
and AND3 (N246, N241, N220, N87);
xor XOR2 (N247, N239, N208);
xor XOR2 (N248, N242, N226);
buf BUF1 (N249, N228);
xor XOR2 (N250, N247, N190);
nand NAND4 (N251, N250, N4, N121, N190);
or OR2 (N252, N248, N207);
nor NOR2 (N253, N246, N236);
and AND2 (N254, N70, N8);
nand NAND2 (N255, N253, N12);
or OR4 (N256, N255, N224, N203, N240);
buf BUF1 (N257, N244);
and AND4 (N258, N252, N136, N240, N253);
or OR2 (N259, N235, N76);
xor XOR2 (N260, N243, N71);
xor XOR2 (N261, N254, N152);
or OR4 (N262, N249, N149, N232, N254);
buf BUF1 (N263, N251);
xor XOR2 (N264, N259, N189);
not NOT1 (N265, N256);
or OR4 (N266, N260, N102, N236, N239);
or OR4 (N267, N258, N228, N195, N81);
buf BUF1 (N268, N266);
nand NAND2 (N269, N268, N99);
or OR2 (N270, N269, N9);
nand NAND4 (N271, N237, N185, N265, N27);
xor XOR2 (N272, N59, N11);
buf BUF1 (N273, N263);
nor NOR2 (N274, N271, N68);
and AND4 (N275, N264, N253, N115, N49);
nor NOR3 (N276, N272, N115, N47);
buf BUF1 (N277, N257);
buf BUF1 (N278, N273);
nor NOR3 (N279, N274, N219, N250);
and AND3 (N280, N262, N70, N150);
xor XOR2 (N281, N275, N111);
buf BUF1 (N282, N261);
nor NOR3 (N283, N277, N60, N46);
or OR3 (N284, N245, N12, N53);
nand NAND3 (N285, N282, N130, N83);
nor NOR3 (N286, N281, N224, N161);
buf BUF1 (N287, N283);
not NOT1 (N288, N278);
nor NOR2 (N289, N284, N127);
or OR3 (N290, N280, N7, N248);
nor NOR2 (N291, N276, N156);
or OR4 (N292, N285, N20, N187, N153);
buf BUF1 (N293, N287);
and AND4 (N294, N286, N102, N193, N109);
xor XOR2 (N295, N267, N35);
or OR4 (N296, N288, N202, N130, N262);
not NOT1 (N297, N291);
not NOT1 (N298, N293);
buf BUF1 (N299, N294);
nand NAND2 (N300, N279, N286);
nand NAND3 (N301, N295, N106, N74);
xor XOR2 (N302, N290, N46);
or OR2 (N303, N296, N173);
or OR3 (N304, N297, N295, N22);
and AND3 (N305, N302, N202, N162);
buf BUF1 (N306, N300);
nor NOR3 (N307, N299, N31, N69);
nand NAND2 (N308, N289, N44);
or OR4 (N309, N307, N56, N80, N53);
xor XOR2 (N310, N292, N165);
nor NOR3 (N311, N305, N269, N114);
not NOT1 (N312, N303);
nor NOR2 (N313, N306, N76);
nand NAND3 (N314, N308, N284, N131);
nor NOR2 (N315, N313, N188);
nand NAND2 (N316, N270, N165);
nand NAND3 (N317, N298, N113, N270);
buf BUF1 (N318, N310);
not NOT1 (N319, N314);
not NOT1 (N320, N315);
buf BUF1 (N321, N304);
nor NOR2 (N322, N318, N11);
buf BUF1 (N323, N321);
and AND4 (N324, N312, N298, N104, N121);
nor NOR4 (N325, N316, N227, N151, N149);
or OR3 (N326, N301, N94, N171);
and AND3 (N327, N323, N194, N62);
and AND4 (N328, N324, N124, N159, N146);
not NOT1 (N329, N328);
or OR3 (N330, N326, N304, N226);
buf BUF1 (N331, N319);
nor NOR4 (N332, N330, N321, N296, N178);
or OR2 (N333, N325, N157);
xor XOR2 (N334, N309, N107);
or OR4 (N335, N334, N242, N248, N107);
buf BUF1 (N336, N320);
nand NAND3 (N337, N332, N291, N71);
buf BUF1 (N338, N311);
not NOT1 (N339, N327);
xor XOR2 (N340, N337, N55);
and AND2 (N341, N331, N247);
buf BUF1 (N342, N336);
nand NAND2 (N343, N338, N320);
buf BUF1 (N344, N339);
nor NOR3 (N345, N342, N3, N105);
not NOT1 (N346, N322);
xor XOR2 (N347, N343, N184);
xor XOR2 (N348, N347, N295);
or OR4 (N349, N341, N236, N130, N297);
buf BUF1 (N350, N335);
or OR3 (N351, N340, N77, N39);
not NOT1 (N352, N351);
or OR2 (N353, N333, N186);
or OR2 (N354, N329, N328);
not NOT1 (N355, N346);
and AND4 (N356, N317, N177, N265, N291);
and AND2 (N357, N354, N163);
and AND3 (N358, N345, N215, N339);
and AND2 (N359, N355, N76);
not NOT1 (N360, N358);
and AND2 (N361, N350, N194);
nand NAND2 (N362, N344, N132);
nand NAND3 (N363, N361, N252, N90);
and AND2 (N364, N362, N311);
buf BUF1 (N365, N364);
nor NOR4 (N366, N360, N339, N193, N331);
not NOT1 (N367, N349);
nor NOR2 (N368, N357, N60);
or OR3 (N369, N356, N36, N239);
not NOT1 (N370, N352);
not NOT1 (N371, N369);
not NOT1 (N372, N366);
not NOT1 (N373, N363);
nand NAND4 (N374, N367, N363, N287, N72);
buf BUF1 (N375, N353);
nor NOR3 (N376, N348, N32, N129);
nand NAND2 (N377, N376, N47);
not NOT1 (N378, N365);
nor NOR3 (N379, N368, N348, N24);
and AND4 (N380, N379, N126, N309, N331);
nand NAND2 (N381, N373, N33);
xor XOR2 (N382, N381, N279);
not NOT1 (N383, N370);
or OR2 (N384, N383, N202);
not NOT1 (N385, N384);
nand NAND4 (N386, N382, N349, N19, N161);
xor XOR2 (N387, N372, N223);
or OR4 (N388, N359, N380, N26, N47);
nor NOR3 (N389, N74, N364, N124);
not NOT1 (N390, N389);
buf BUF1 (N391, N386);
and AND2 (N392, N375, N165);
and AND3 (N393, N377, N59, N122);
nand NAND4 (N394, N390, N89, N352, N224);
buf BUF1 (N395, N392);
nand NAND4 (N396, N395, N315, N54, N99);
xor XOR2 (N397, N374, N23);
buf BUF1 (N398, N378);
or OR2 (N399, N391, N100);
or OR4 (N400, N371, N174, N315, N18);
nand NAND2 (N401, N396, N233);
not NOT1 (N402, N387);
or OR3 (N403, N399, N384, N100);
nand NAND4 (N404, N403, N50, N97, N190);
or OR4 (N405, N385, N214, N275, N301);
and AND3 (N406, N400, N166, N67);
not NOT1 (N407, N405);
nor NOR4 (N408, N393, N260, N371, N212);
not NOT1 (N409, N388);
and AND4 (N410, N401, N66, N204, N142);
nor NOR2 (N411, N397, N219);
nor NOR4 (N412, N402, N18, N138, N187);
xor XOR2 (N413, N412, N402);
or OR4 (N414, N406, N278, N281, N101);
buf BUF1 (N415, N407);
and AND4 (N416, N413, N384, N229, N178);
nand NAND4 (N417, N410, N313, N365, N414);
nand NAND2 (N418, N57, N53);
or OR3 (N419, N404, N171, N131);
buf BUF1 (N420, N408);
nand NAND4 (N421, N418, N207, N160, N167);
not NOT1 (N422, N394);
nand NAND3 (N423, N419, N78, N18);
nand NAND4 (N424, N411, N326, N69, N335);
or OR2 (N425, N424, N266);
buf BUF1 (N426, N416);
buf BUF1 (N427, N398);
or OR3 (N428, N409, N62, N417);
nor NOR4 (N429, N335, N193, N403, N374);
xor XOR2 (N430, N429, N85);
and AND2 (N431, N427, N260);
not NOT1 (N432, N430);
xor XOR2 (N433, N426, N257);
nor NOR4 (N434, N431, N208, N327, N394);
and AND3 (N435, N425, N273, N137);
buf BUF1 (N436, N415);
nor NOR2 (N437, N432, N114);
buf BUF1 (N438, N433);
and AND2 (N439, N438, N173);
not NOT1 (N440, N428);
nand NAND4 (N441, N436, N328, N210, N29);
or OR4 (N442, N441, N418, N247, N124);
or OR2 (N443, N420, N136);
buf BUF1 (N444, N421);
xor XOR2 (N445, N444, N324);
buf BUF1 (N446, N440);
not NOT1 (N447, N439);
xor XOR2 (N448, N437, N141);
buf BUF1 (N449, N445);
or OR3 (N450, N435, N343, N85);
xor XOR2 (N451, N448, N78);
nor NOR3 (N452, N434, N154, N124);
nand NAND4 (N453, N446, N259, N417, N323);
not NOT1 (N454, N452);
xor XOR2 (N455, N442, N192);
nand NAND4 (N456, N453, N254, N268, N310);
xor XOR2 (N457, N451, N137);
xor XOR2 (N458, N454, N149);
not NOT1 (N459, N447);
xor XOR2 (N460, N423, N313);
xor XOR2 (N461, N456, N187);
or OR3 (N462, N449, N203, N374);
or OR4 (N463, N461, N54, N394, N203);
or OR2 (N464, N458, N305);
buf BUF1 (N465, N462);
nor NOR4 (N466, N464, N330, N142, N260);
or OR4 (N467, N455, N93, N40, N67);
or OR2 (N468, N457, N102);
not NOT1 (N469, N467);
nand NAND4 (N470, N465, N128, N276, N222);
not NOT1 (N471, N450);
or OR4 (N472, N422, N212, N280, N179);
and AND3 (N473, N472, N273, N216);
nor NOR4 (N474, N468, N256, N38, N188);
or OR4 (N475, N463, N451, N468, N445);
not NOT1 (N476, N443);
or OR2 (N477, N460, N350);
xor XOR2 (N478, N473, N129);
not NOT1 (N479, N474);
and AND2 (N480, N476, N356);
and AND4 (N481, N480, N140, N429, N312);
nand NAND3 (N482, N475, N292, N124);
not NOT1 (N483, N479);
not NOT1 (N484, N470);
and AND3 (N485, N483, N241, N147);
buf BUF1 (N486, N484);
not NOT1 (N487, N469);
not NOT1 (N488, N485);
nor NOR3 (N489, N466, N266, N98);
not NOT1 (N490, N486);
not NOT1 (N491, N478);
not NOT1 (N492, N489);
not NOT1 (N493, N488);
nor NOR3 (N494, N459, N75, N243);
nor NOR2 (N495, N482, N444);
and AND4 (N496, N492, N349, N347, N451);
buf BUF1 (N497, N477);
not NOT1 (N498, N497);
nand NAND3 (N499, N490, N467, N297);
not NOT1 (N500, N495);
buf BUF1 (N501, N496);
or OR3 (N502, N499, N264, N234);
nand NAND4 (N503, N500, N322, N374, N495);
nor NOR4 (N504, N493, N254, N348, N450);
not NOT1 (N505, N494);
not NOT1 (N506, N487);
buf BUF1 (N507, N504);
or OR4 (N508, N481, N313, N79, N289);
buf BUF1 (N509, N502);
nor NOR4 (N510, N491, N103, N52, N299);
or OR2 (N511, N506, N210);
and AND3 (N512, N503, N210, N498);
buf BUF1 (N513, N478);
not NOT1 (N514, N512);
or OR4 (N515, N507, N35, N255, N138);
xor XOR2 (N516, N505, N15);
xor XOR2 (N517, N515, N201);
not NOT1 (N518, N513);
xor XOR2 (N519, N471, N443);
nor NOR2 (N520, N510, N344);
xor XOR2 (N521, N518, N139);
or OR3 (N522, N519, N59, N483);
not NOT1 (N523, N522);
nor NOR3 (N524, N508, N332, N314);
nand NAND3 (N525, N509, N366, N503);
buf BUF1 (N526, N517);
nand NAND2 (N527, N514, N220);
xor XOR2 (N528, N520, N277);
xor XOR2 (N529, N527, N78);
buf BUF1 (N530, N523);
nor NOR4 (N531, N525, N472, N344, N408);
not NOT1 (N532, N516);
nor NOR3 (N533, N532, N202, N137);
buf BUF1 (N534, N529);
buf BUF1 (N535, N524);
not NOT1 (N536, N530);
or OR2 (N537, N501, N309);
not NOT1 (N538, N531);
not NOT1 (N539, N536);
or OR2 (N540, N526, N455);
and AND4 (N541, N535, N238, N339, N439);
buf BUF1 (N542, N537);
nor NOR4 (N543, N538, N423, N526, N313);
buf BUF1 (N544, N533);
xor XOR2 (N545, N542, N463);
and AND4 (N546, N511, N2, N24, N221);
and AND4 (N547, N521, N492, N296, N322);
xor XOR2 (N548, N540, N380);
and AND4 (N549, N546, N170, N441, N183);
nand NAND3 (N550, N547, N476, N45);
or OR3 (N551, N539, N446, N334);
and AND3 (N552, N543, N138, N160);
and AND2 (N553, N528, N238);
nand NAND3 (N554, N549, N307, N527);
nor NOR2 (N555, N541, N230);
buf BUF1 (N556, N545);
nand NAND3 (N557, N551, N515, N427);
nand NAND3 (N558, N552, N342, N229);
nor NOR3 (N559, N548, N205, N28);
not NOT1 (N560, N557);
or OR2 (N561, N550, N544);
nor NOR4 (N562, N71, N47, N440, N476);
xor XOR2 (N563, N555, N452);
or OR4 (N564, N563, N345, N236, N76);
nand NAND4 (N565, N534, N295, N537, N469);
nand NAND3 (N566, N565, N119, N489);
and AND2 (N567, N561, N201);
nand NAND3 (N568, N566, N178, N4);
or OR2 (N569, N567, N73);
buf BUF1 (N570, N562);
buf BUF1 (N571, N570);
buf BUF1 (N572, N556);
buf BUF1 (N573, N572);
nor NOR4 (N574, N569, N206, N543, N16);
nand NAND2 (N575, N574, N123);
nor NOR3 (N576, N573, N182, N398);
not NOT1 (N577, N554);
and AND3 (N578, N558, N357, N185);
nor NOR3 (N579, N575, N329, N331);
buf BUF1 (N580, N579);
buf BUF1 (N581, N568);
and AND4 (N582, N560, N200, N217, N562);
and AND3 (N583, N553, N33, N183);
not NOT1 (N584, N576);
buf BUF1 (N585, N578);
and AND4 (N586, N559, N253, N146, N449);
or OR2 (N587, N577, N551);
and AND3 (N588, N564, N249, N60);
not NOT1 (N589, N585);
or OR2 (N590, N589, N377);
nor NOR3 (N591, N588, N372, N114);
and AND4 (N592, N591, N485, N192, N381);
or OR2 (N593, N587, N4);
nand NAND2 (N594, N581, N160);
nand NAND3 (N595, N584, N144, N466);
or OR2 (N596, N595, N58);
nand NAND2 (N597, N592, N517);
xor XOR2 (N598, N590, N162);
nand NAND2 (N599, N597, N119);
nor NOR3 (N600, N583, N278, N82);
nand NAND3 (N601, N600, N430, N113);
xor XOR2 (N602, N599, N293);
nand NAND4 (N603, N594, N181, N528, N256);
nand NAND4 (N604, N593, N419, N317, N132);
nand NAND4 (N605, N598, N109, N213, N72);
and AND3 (N606, N601, N244, N96);
nor NOR2 (N607, N603, N155);
buf BUF1 (N608, N605);
nand NAND2 (N609, N602, N508);
not NOT1 (N610, N604);
nand NAND2 (N611, N609, N50);
nor NOR2 (N612, N596, N463);
buf BUF1 (N613, N571);
xor XOR2 (N614, N608, N556);
buf BUF1 (N615, N607);
xor XOR2 (N616, N613, N56);
xor XOR2 (N617, N606, N555);
nor NOR2 (N618, N612, N615);
nand NAND4 (N619, N323, N111, N29, N507);
and AND4 (N620, N619, N375, N190, N305);
buf BUF1 (N621, N616);
or OR2 (N622, N610, N208);
not NOT1 (N623, N620);
and AND2 (N624, N618, N145);
nand NAND2 (N625, N614, N364);
not NOT1 (N626, N611);
xor XOR2 (N627, N625, N56);
or OR4 (N628, N580, N54, N9, N157);
nand NAND3 (N629, N626, N535, N126);
buf BUF1 (N630, N627);
and AND3 (N631, N621, N6, N279);
xor XOR2 (N632, N622, N340);
and AND3 (N633, N629, N304, N443);
nand NAND2 (N634, N631, N384);
and AND4 (N635, N632, N141, N239, N378);
buf BUF1 (N636, N628);
nand NAND2 (N637, N634, N350);
or OR2 (N638, N582, N111);
nand NAND4 (N639, N623, N446, N352, N426);
nand NAND4 (N640, N636, N100, N166, N3);
nand NAND3 (N641, N624, N58, N82);
buf BUF1 (N642, N617);
not NOT1 (N643, N633);
or OR3 (N644, N643, N221, N51);
not NOT1 (N645, N642);
nand NAND2 (N646, N644, N343);
buf BUF1 (N647, N630);
nand NAND2 (N648, N639, N469);
and AND4 (N649, N640, N382, N617, N117);
buf BUF1 (N650, N647);
nand NAND3 (N651, N648, N185, N68);
not NOT1 (N652, N649);
nand NAND4 (N653, N635, N96, N189, N502);
nand NAND3 (N654, N638, N88, N448);
and AND3 (N655, N645, N364, N29);
nand NAND3 (N656, N652, N325, N43);
buf BUF1 (N657, N656);
nand NAND2 (N658, N657, N643);
buf BUF1 (N659, N658);
not NOT1 (N660, N637);
nand NAND2 (N661, N651, N346);
nor NOR2 (N662, N659, N489);
nor NOR3 (N663, N660, N284, N162);
and AND4 (N664, N661, N455, N394, N20);
or OR2 (N665, N586, N195);
xor XOR2 (N666, N664, N309);
nor NOR3 (N667, N662, N297, N298);
buf BUF1 (N668, N646);
nor NOR4 (N669, N666, N200, N424, N459);
nand NAND4 (N670, N663, N427, N243, N147);
nor NOR4 (N671, N655, N310, N168, N154);
xor XOR2 (N672, N665, N592);
and AND3 (N673, N654, N503, N319);
or OR3 (N674, N650, N136, N248);
xor XOR2 (N675, N641, N100);
nor NOR2 (N676, N668, N12);
xor XOR2 (N677, N675, N490);
buf BUF1 (N678, N669);
xor XOR2 (N679, N678, N346);
buf BUF1 (N680, N672);
nor NOR2 (N681, N679, N562);
buf BUF1 (N682, N680);
and AND3 (N683, N681, N99, N70);
buf BUF1 (N684, N667);
nor NOR4 (N685, N677, N68, N155, N281);
nand NAND4 (N686, N682, N398, N87, N216);
or OR3 (N687, N674, N532, N502);
nand NAND4 (N688, N687, N498, N109, N132);
not NOT1 (N689, N686);
buf BUF1 (N690, N676);
or OR2 (N691, N688, N143);
buf BUF1 (N692, N683);
or OR3 (N693, N690, N530, N309);
not NOT1 (N694, N673);
nand NAND2 (N695, N653, N231);
and AND2 (N696, N671, N147);
xor XOR2 (N697, N692, N510);
xor XOR2 (N698, N691, N238);
xor XOR2 (N699, N696, N132);
nand NAND4 (N700, N685, N332, N383, N658);
not NOT1 (N701, N699);
not NOT1 (N702, N697);
nand NAND2 (N703, N695, N59);
nand NAND4 (N704, N693, N685, N150, N579);
buf BUF1 (N705, N684);
xor XOR2 (N706, N702, N595);
nor NOR3 (N707, N705, N629, N297);
not NOT1 (N708, N694);
not NOT1 (N709, N707);
buf BUF1 (N710, N706);
and AND3 (N711, N701, N229, N183);
buf BUF1 (N712, N689);
buf BUF1 (N713, N709);
and AND3 (N714, N700, N145, N53);
nor NOR2 (N715, N712, N72);
xor XOR2 (N716, N704, N672);
and AND2 (N717, N716, N216);
or OR3 (N718, N714, N243, N239);
or OR3 (N719, N703, N310, N718);
xor XOR2 (N720, N271, N36);
not NOT1 (N721, N698);
and AND4 (N722, N715, N29, N132, N121);
buf BUF1 (N723, N670);
buf BUF1 (N724, N710);
not NOT1 (N725, N722);
not NOT1 (N726, N719);
and AND4 (N727, N720, N485, N129, N448);
nor NOR2 (N728, N711, N179);
buf BUF1 (N729, N724);
not NOT1 (N730, N729);
or OR3 (N731, N726, N496, N206);
nor NOR2 (N732, N727, N501);
nor NOR3 (N733, N721, N313, N251);
xor XOR2 (N734, N723, N357);
or OR4 (N735, N731, N205, N494, N363);
and AND2 (N736, N725, N605);
buf BUF1 (N737, N717);
nor NOR2 (N738, N733, N178);
xor XOR2 (N739, N735, N478);
or OR4 (N740, N732, N541, N437, N464);
not NOT1 (N741, N737);
nor NOR4 (N742, N728, N2, N258, N415);
not NOT1 (N743, N730);
xor XOR2 (N744, N741, N34);
xor XOR2 (N745, N738, N389);
or OR3 (N746, N708, N47, N541);
xor XOR2 (N747, N739, N171);
xor XOR2 (N748, N736, N203);
or OR4 (N749, N743, N302, N126, N95);
not NOT1 (N750, N748);
buf BUF1 (N751, N740);
nand NAND3 (N752, N745, N350, N473);
xor XOR2 (N753, N734, N144);
nand NAND2 (N754, N749, N608);
nand NAND4 (N755, N746, N727, N675, N104);
not NOT1 (N756, N742);
nor NOR3 (N757, N754, N735, N690);
buf BUF1 (N758, N756);
nor NOR2 (N759, N755, N228);
xor XOR2 (N760, N747, N60);
not NOT1 (N761, N759);
not NOT1 (N762, N752);
nand NAND3 (N763, N758, N721, N20);
not NOT1 (N764, N750);
nand NAND4 (N765, N762, N423, N308, N446);
not NOT1 (N766, N763);
nor NOR4 (N767, N766, N463, N734, N199);
nor NOR2 (N768, N760, N623);
not NOT1 (N769, N757);
xor XOR2 (N770, N744, N146);
nor NOR4 (N771, N765, N565, N206, N565);
buf BUF1 (N772, N768);
nor NOR2 (N773, N771, N546);
buf BUF1 (N774, N753);
nor NOR3 (N775, N774, N305, N71);
nor NOR4 (N776, N751, N328, N1, N362);
nand NAND2 (N777, N764, N487);
nor NOR3 (N778, N773, N152, N358);
nand NAND2 (N779, N713, N181);
xor XOR2 (N780, N772, N143);
nand NAND3 (N781, N778, N605, N208);
nor NOR2 (N782, N777, N576);
and AND2 (N783, N767, N538);
or OR2 (N784, N781, N82);
or OR2 (N785, N775, N11);
not NOT1 (N786, N780);
buf BUF1 (N787, N783);
or OR2 (N788, N779, N594);
and AND3 (N789, N782, N97, N515);
and AND4 (N790, N787, N51, N56, N694);
nor NOR4 (N791, N790, N703, N358, N507);
xor XOR2 (N792, N784, N534);
or OR4 (N793, N785, N612, N478, N596);
or OR3 (N794, N770, N210, N111);
nor NOR4 (N795, N761, N364, N371, N183);
and AND2 (N796, N786, N422);
or OR3 (N797, N791, N167, N497);
nor NOR3 (N798, N794, N662, N791);
nand NAND4 (N799, N769, N118, N260, N387);
nand NAND2 (N800, N796, N624);
not NOT1 (N801, N799);
xor XOR2 (N802, N776, N758);
buf BUF1 (N803, N801);
nand NAND4 (N804, N797, N15, N153, N528);
and AND2 (N805, N792, N436);
not NOT1 (N806, N788);
buf BUF1 (N807, N802);
not NOT1 (N808, N798);
nor NOR2 (N809, N806, N462);
not NOT1 (N810, N803);
or OR2 (N811, N789, N193);
xor XOR2 (N812, N795, N781);
nor NOR3 (N813, N810, N567, N579);
xor XOR2 (N814, N800, N14);
nand NAND3 (N815, N811, N147, N617);
xor XOR2 (N816, N807, N402);
nand NAND3 (N817, N804, N403, N390);
or OR2 (N818, N812, N747);
not NOT1 (N819, N814);
xor XOR2 (N820, N815, N513);
xor XOR2 (N821, N808, N389);
nor NOR3 (N822, N793, N709, N239);
and AND3 (N823, N805, N399, N52);
nor NOR2 (N824, N817, N442);
buf BUF1 (N825, N809);
or OR4 (N826, N816, N420, N385, N200);
nand NAND3 (N827, N826, N478, N381);
and AND4 (N828, N825, N762, N330, N618);
not NOT1 (N829, N819);
not NOT1 (N830, N821);
xor XOR2 (N831, N820, N515);
and AND2 (N832, N824, N476);
not NOT1 (N833, N831);
not NOT1 (N834, N813);
and AND4 (N835, N822, N176, N773, N732);
nor NOR2 (N836, N830, N30);
xor XOR2 (N837, N827, N715);
or OR4 (N838, N836, N569, N665, N134);
or OR4 (N839, N832, N466, N282, N68);
buf BUF1 (N840, N818);
or OR2 (N841, N835, N582);
not NOT1 (N842, N841);
buf BUF1 (N843, N828);
not NOT1 (N844, N842);
nor NOR3 (N845, N829, N783, N178);
xor XOR2 (N846, N833, N548);
not NOT1 (N847, N839);
buf BUF1 (N848, N838);
buf BUF1 (N849, N844);
or OR2 (N850, N843, N413);
xor XOR2 (N851, N849, N637);
nand NAND4 (N852, N840, N377, N519, N38);
not NOT1 (N853, N851);
nand NAND4 (N854, N846, N562, N623, N688);
and AND4 (N855, N854, N728, N228, N351);
nor NOR2 (N856, N852, N402);
not NOT1 (N857, N856);
or OR2 (N858, N850, N368);
buf BUF1 (N859, N823);
nor NOR2 (N860, N837, N296);
not NOT1 (N861, N834);
buf BUF1 (N862, N845);
nor NOR4 (N863, N861, N522, N709, N830);
and AND2 (N864, N857, N465);
buf BUF1 (N865, N862);
or OR2 (N866, N863, N11);
nor NOR3 (N867, N858, N200, N142);
or OR3 (N868, N853, N680, N641);
xor XOR2 (N869, N859, N687);
not NOT1 (N870, N847);
and AND2 (N871, N864, N13);
buf BUF1 (N872, N871);
xor XOR2 (N873, N867, N112);
nor NOR3 (N874, N860, N494, N839);
buf BUF1 (N875, N868);
or OR4 (N876, N873, N214, N683, N401);
nor NOR4 (N877, N872, N239, N349, N83);
and AND2 (N878, N865, N159);
not NOT1 (N879, N878);
xor XOR2 (N880, N866, N361);
and AND2 (N881, N877, N724);
nand NAND2 (N882, N879, N89);
buf BUF1 (N883, N875);
nand NAND4 (N884, N869, N631, N847, N430);
xor XOR2 (N885, N876, N360);
nand NAND4 (N886, N881, N348, N339, N310);
xor XOR2 (N887, N882, N150);
and AND3 (N888, N870, N154, N51);
nor NOR3 (N889, N848, N783, N657);
nand NAND2 (N890, N884, N732);
and AND2 (N891, N889, N545);
not NOT1 (N892, N891);
and AND4 (N893, N890, N291, N832, N461);
nor NOR2 (N894, N855, N149);
and AND4 (N895, N887, N512, N793, N787);
buf BUF1 (N896, N892);
nand NAND2 (N897, N886, N328);
buf BUF1 (N898, N897);
nor NOR2 (N899, N895, N624);
nor NOR3 (N900, N888, N59, N806);
or OR4 (N901, N883, N629, N736, N146);
nor NOR4 (N902, N880, N351, N127, N658);
buf BUF1 (N903, N893);
not NOT1 (N904, N902);
and AND2 (N905, N900, N409);
not NOT1 (N906, N905);
nor NOR3 (N907, N874, N620, N7);
nand NAND2 (N908, N906, N316);
and AND4 (N909, N903, N242, N487, N366);
not NOT1 (N910, N896);
nand NAND3 (N911, N899, N252, N652);
and AND3 (N912, N901, N582, N891);
or OR2 (N913, N894, N910);
xor XOR2 (N914, N565, N36);
nor NOR2 (N915, N913, N25);
nand NAND3 (N916, N914, N466, N589);
nor NOR2 (N917, N909, N13);
buf BUF1 (N918, N916);
nand NAND2 (N919, N904, N608);
nand NAND3 (N920, N915, N420, N505);
buf BUF1 (N921, N907);
not NOT1 (N922, N919);
not NOT1 (N923, N898);
nor NOR2 (N924, N922, N788);
or OR2 (N925, N918, N144);
not NOT1 (N926, N920);
xor XOR2 (N927, N912, N20);
or OR3 (N928, N923, N916, N585);
xor XOR2 (N929, N921, N69);
buf BUF1 (N930, N928);
buf BUF1 (N931, N927);
xor XOR2 (N932, N885, N857);
or OR2 (N933, N911, N699);
or OR4 (N934, N931, N918, N723, N573);
or OR3 (N935, N926, N624, N604);
xor XOR2 (N936, N925, N222);
or OR4 (N937, N930, N109, N316, N72);
xor XOR2 (N938, N929, N821);
nor NOR2 (N939, N924, N123);
nand NAND2 (N940, N938, N656);
or OR4 (N941, N932, N380, N724, N249);
or OR2 (N942, N937, N888);
nor NOR4 (N943, N940, N937, N860, N928);
not NOT1 (N944, N943);
or OR2 (N945, N935, N157);
and AND2 (N946, N933, N271);
nand NAND3 (N947, N945, N735, N838);
or OR4 (N948, N941, N941, N579, N648);
not NOT1 (N949, N936);
nor NOR4 (N950, N917, N163, N149, N559);
xor XOR2 (N951, N942, N694);
buf BUF1 (N952, N951);
or OR2 (N953, N950, N385);
nor NOR3 (N954, N952, N926, N541);
and AND4 (N955, N947, N343, N178, N1);
not NOT1 (N956, N953);
not NOT1 (N957, N949);
nand NAND2 (N958, N954, N25);
nand NAND4 (N959, N946, N530, N935, N707);
nor NOR3 (N960, N958, N295, N460);
and AND2 (N961, N957, N109);
not NOT1 (N962, N908);
xor XOR2 (N963, N959, N531);
xor XOR2 (N964, N956, N647);
buf BUF1 (N965, N963);
buf BUF1 (N966, N960);
or OR3 (N967, N962, N137, N165);
and AND4 (N968, N934, N374, N813, N481);
not NOT1 (N969, N966);
or OR3 (N970, N939, N74, N450);
buf BUF1 (N971, N948);
or OR2 (N972, N968, N382);
not NOT1 (N973, N971);
and AND2 (N974, N961, N194);
buf BUF1 (N975, N964);
buf BUF1 (N976, N955);
or OR3 (N977, N944, N461, N876);
nand NAND3 (N978, N976, N566, N676);
and AND4 (N979, N977, N888, N316, N794);
buf BUF1 (N980, N973);
nand NAND4 (N981, N970, N744, N864, N188);
nand NAND2 (N982, N978, N490);
not NOT1 (N983, N980);
nand NAND4 (N984, N983, N851, N865, N861);
or OR4 (N985, N982, N815, N656, N825);
nor NOR2 (N986, N979, N826);
not NOT1 (N987, N974);
not NOT1 (N988, N981);
nand NAND2 (N989, N969, N602);
nor NOR4 (N990, N972, N506, N404, N240);
and AND2 (N991, N987, N544);
or OR3 (N992, N986, N959, N232);
not NOT1 (N993, N991);
not NOT1 (N994, N985);
nor NOR4 (N995, N984, N130, N273, N740);
and AND4 (N996, N975, N339, N207, N35);
nand NAND3 (N997, N990, N770, N931);
nor NOR2 (N998, N992, N614);
not NOT1 (N999, N997);
xor XOR2 (N1000, N998, N161);
or OR4 (N1001, N994, N392, N890, N107);
and AND4 (N1002, N988, N331, N118, N481);
nor NOR4 (N1003, N989, N294, N119, N906);
xor XOR2 (N1004, N1002, N302);
not NOT1 (N1005, N996);
nand NAND3 (N1006, N1003, N721, N330);
buf BUF1 (N1007, N1004);
buf BUF1 (N1008, N965);
or OR3 (N1009, N1008, N797, N324);
not NOT1 (N1010, N999);
nor NOR3 (N1011, N1001, N225, N366);
and AND2 (N1012, N1000, N563);
not NOT1 (N1013, N967);
and AND2 (N1014, N1013, N979);
and AND4 (N1015, N1006, N308, N120, N284);
and AND4 (N1016, N995, N147, N863, N497);
nor NOR4 (N1017, N993, N731, N908, N332);
buf BUF1 (N1018, N1007);
and AND2 (N1019, N1017, N480);
and AND3 (N1020, N1012, N158, N443);
and AND3 (N1021, N1011, N608, N908);
nor NOR4 (N1022, N1016, N957, N652, N704);
or OR4 (N1023, N1019, N634, N248, N842);
not NOT1 (N1024, N1021);
xor XOR2 (N1025, N1009, N315);
nor NOR2 (N1026, N1015, N880);
nand NAND3 (N1027, N1005, N162, N622);
not NOT1 (N1028, N1020);
buf BUF1 (N1029, N1022);
buf BUF1 (N1030, N1023);
nor NOR4 (N1031, N1027, N650, N588, N795);
xor XOR2 (N1032, N1029, N372);
or OR3 (N1033, N1024, N348, N546);
and AND2 (N1034, N1014, N39);
or OR4 (N1035, N1028, N855, N88, N124);
nand NAND4 (N1036, N1033, N271, N288, N605);
not NOT1 (N1037, N1035);
nor NOR3 (N1038, N1037, N167, N710);
and AND2 (N1039, N1010, N711);
nor NOR2 (N1040, N1038, N45);
xor XOR2 (N1041, N1039, N895);
nand NAND4 (N1042, N1018, N986, N368, N938);
or OR2 (N1043, N1042, N506);
xor XOR2 (N1044, N1041, N544);
nand NAND2 (N1045, N1043, N355);
and AND3 (N1046, N1034, N705, N59);
nor NOR2 (N1047, N1036, N312);
buf BUF1 (N1048, N1032);
or OR4 (N1049, N1040, N315, N460, N814);
buf BUF1 (N1050, N1031);
not NOT1 (N1051, N1049);
nand NAND3 (N1052, N1046, N818, N732);
and AND2 (N1053, N1030, N343);
nor NOR3 (N1054, N1025, N307, N1019);
buf BUF1 (N1055, N1054);
nor NOR4 (N1056, N1052, N367, N626, N700);
nand NAND3 (N1057, N1048, N189, N612);
or OR2 (N1058, N1056, N445);
buf BUF1 (N1059, N1053);
and AND3 (N1060, N1045, N971, N457);
and AND4 (N1061, N1059, N240, N547, N1020);
buf BUF1 (N1062, N1026);
not NOT1 (N1063, N1044);
or OR4 (N1064, N1060, N191, N328, N270);
and AND4 (N1065, N1047, N175, N818, N484);
and AND3 (N1066, N1064, N462, N1045);
nand NAND3 (N1067, N1055, N524, N619);
or OR4 (N1068, N1050, N432, N710, N973);
buf BUF1 (N1069, N1065);
nor NOR3 (N1070, N1057, N554, N135);
xor XOR2 (N1071, N1070, N115);
buf BUF1 (N1072, N1061);
xor XOR2 (N1073, N1051, N164);
not NOT1 (N1074, N1062);
not NOT1 (N1075, N1067);
nand NAND2 (N1076, N1071, N479);
or OR2 (N1077, N1069, N807);
or OR4 (N1078, N1075, N145, N275, N1070);
or OR4 (N1079, N1076, N440, N680, N815);
xor XOR2 (N1080, N1058, N433);
or OR3 (N1081, N1063, N131, N14);
nor NOR4 (N1082, N1080, N392, N208, N568);
not NOT1 (N1083, N1072);
and AND3 (N1084, N1082, N16, N79);
not NOT1 (N1085, N1077);
or OR2 (N1086, N1078, N315);
not NOT1 (N1087, N1068);
nand NAND3 (N1088, N1084, N207, N232);
xor XOR2 (N1089, N1073, N778);
nand NAND3 (N1090, N1088, N347, N464);
xor XOR2 (N1091, N1083, N131);
buf BUF1 (N1092, N1085);
nor NOR4 (N1093, N1087, N389, N1049, N1040);
and AND3 (N1094, N1086, N539, N297);
and AND4 (N1095, N1093, N787, N705, N572);
or OR4 (N1096, N1079, N594, N824, N892);
or OR2 (N1097, N1066, N170);
nand NAND4 (N1098, N1096, N165, N629, N391);
or OR3 (N1099, N1098, N13, N594);
buf BUF1 (N1100, N1081);
nor NOR2 (N1101, N1094, N185);
nand NAND2 (N1102, N1101, N19);
or OR3 (N1103, N1097, N1037, N597);
or OR3 (N1104, N1102, N64, N726);
buf BUF1 (N1105, N1090);
nor NOR3 (N1106, N1100, N779, N1098);
buf BUF1 (N1107, N1104);
xor XOR2 (N1108, N1091, N153);
nor NOR3 (N1109, N1074, N394, N775);
and AND4 (N1110, N1089, N344, N75, N323);
or OR3 (N1111, N1095, N301, N459);
not NOT1 (N1112, N1107);
nor NOR3 (N1113, N1105, N1028, N811);
xor XOR2 (N1114, N1099, N368);
nand NAND3 (N1115, N1110, N770, N100);
xor XOR2 (N1116, N1112, N332);
buf BUF1 (N1117, N1109);
nand NAND3 (N1118, N1108, N500, N1066);
nor NOR3 (N1119, N1111, N759, N1087);
and AND3 (N1120, N1115, N768, N799);
nor NOR4 (N1121, N1119, N725, N725, N505);
nand NAND3 (N1122, N1121, N954, N40);
buf BUF1 (N1123, N1117);
buf BUF1 (N1124, N1116);
buf BUF1 (N1125, N1120);
xor XOR2 (N1126, N1106, N285);
nand NAND4 (N1127, N1118, N1112, N676, N151);
nand NAND2 (N1128, N1123, N174);
or OR3 (N1129, N1103, N1043, N831);
or OR2 (N1130, N1124, N693);
or OR2 (N1131, N1127, N299);
nand NAND4 (N1132, N1092, N11, N5, N582);
buf BUF1 (N1133, N1132);
not NOT1 (N1134, N1125);
nand NAND4 (N1135, N1133, N318, N303, N51);
buf BUF1 (N1136, N1128);
nand NAND3 (N1137, N1122, N745, N1062);
xor XOR2 (N1138, N1129, N175);
xor XOR2 (N1139, N1136, N726);
or OR3 (N1140, N1131, N774, N375);
buf BUF1 (N1141, N1126);
nor NOR3 (N1142, N1137, N772, N833);
buf BUF1 (N1143, N1141);
buf BUF1 (N1144, N1135);
nand NAND3 (N1145, N1113, N775, N356);
nand NAND3 (N1146, N1139, N31, N709);
nand NAND4 (N1147, N1145, N254, N533, N206);
buf BUF1 (N1148, N1130);
not NOT1 (N1149, N1146);
buf BUF1 (N1150, N1143);
nor NOR4 (N1151, N1150, N299, N1082, N829);
not NOT1 (N1152, N1142);
not NOT1 (N1153, N1114);
xor XOR2 (N1154, N1151, N1146);
nor NOR2 (N1155, N1138, N79);
and AND3 (N1156, N1140, N807, N334);
not NOT1 (N1157, N1144);
not NOT1 (N1158, N1155);
or OR2 (N1159, N1153, N535);
and AND2 (N1160, N1152, N492);
and AND2 (N1161, N1154, N95);
not NOT1 (N1162, N1158);
not NOT1 (N1163, N1160);
and AND3 (N1164, N1157, N234, N231);
buf BUF1 (N1165, N1134);
not NOT1 (N1166, N1163);
or OR2 (N1167, N1147, N2);
not NOT1 (N1168, N1159);
nand NAND4 (N1169, N1167, N808, N291, N63);
not NOT1 (N1170, N1166);
and AND2 (N1171, N1164, N94);
nor NOR2 (N1172, N1171, N130);
not NOT1 (N1173, N1162);
nand NAND3 (N1174, N1173, N880, N367);
not NOT1 (N1175, N1165);
buf BUF1 (N1176, N1174);
or OR3 (N1177, N1156, N381, N126);
nand NAND4 (N1178, N1169, N828, N570, N232);
xor XOR2 (N1179, N1175, N751);
and AND4 (N1180, N1177, N278, N120, N223);
not NOT1 (N1181, N1178);
nand NAND2 (N1182, N1179, N854);
or OR4 (N1183, N1170, N14, N1023, N320);
nor NOR4 (N1184, N1172, N935, N890, N160);
buf BUF1 (N1185, N1180);
buf BUF1 (N1186, N1183);
buf BUF1 (N1187, N1185);
or OR2 (N1188, N1161, N961);
not NOT1 (N1189, N1181);
nand NAND3 (N1190, N1176, N205, N449);
nand NAND4 (N1191, N1190, N223, N761, N428);
and AND4 (N1192, N1168, N279, N554, N796);
or OR3 (N1193, N1189, N1170, N9);
or OR2 (N1194, N1187, N444);
or OR3 (N1195, N1193, N229, N1007);
xor XOR2 (N1196, N1149, N1021);
not NOT1 (N1197, N1195);
and AND4 (N1198, N1191, N492, N741, N580);
not NOT1 (N1199, N1194);
and AND3 (N1200, N1182, N515, N620);
xor XOR2 (N1201, N1148, N97);
not NOT1 (N1202, N1198);
and AND2 (N1203, N1197, N890);
nand NAND3 (N1204, N1203, N1169, N1021);
not NOT1 (N1205, N1196);
xor XOR2 (N1206, N1201, N672);
xor XOR2 (N1207, N1206, N421);
not NOT1 (N1208, N1202);
buf BUF1 (N1209, N1188);
and AND3 (N1210, N1205, N356, N668);
or OR3 (N1211, N1207, N791, N590);
not NOT1 (N1212, N1186);
buf BUF1 (N1213, N1210);
or OR3 (N1214, N1192, N761, N1171);
buf BUF1 (N1215, N1211);
or OR2 (N1216, N1184, N60);
and AND3 (N1217, N1200, N401, N670);
not NOT1 (N1218, N1204);
nand NAND4 (N1219, N1208, N516, N355, N33);
xor XOR2 (N1220, N1209, N300);
xor XOR2 (N1221, N1199, N393);
nand NAND2 (N1222, N1218, N602);
nand NAND3 (N1223, N1220, N957, N831);
buf BUF1 (N1224, N1223);
buf BUF1 (N1225, N1216);
or OR4 (N1226, N1225, N35, N207, N646);
and AND3 (N1227, N1224, N1031, N583);
buf BUF1 (N1228, N1213);
xor XOR2 (N1229, N1228, N971);
xor XOR2 (N1230, N1212, N35);
or OR2 (N1231, N1215, N831);
buf BUF1 (N1232, N1217);
nor NOR3 (N1233, N1214, N793, N870);
buf BUF1 (N1234, N1232);
buf BUF1 (N1235, N1219);
or OR4 (N1236, N1222, N743, N1228, N531);
not NOT1 (N1237, N1226);
xor XOR2 (N1238, N1236, N907);
and AND4 (N1239, N1235, N420, N827, N1027);
not NOT1 (N1240, N1238);
not NOT1 (N1241, N1237);
or OR3 (N1242, N1240, N648, N1048);
xor XOR2 (N1243, N1231, N596);
nand NAND3 (N1244, N1230, N1042, N319);
or OR3 (N1245, N1242, N518, N1070);
xor XOR2 (N1246, N1227, N489);
nand NAND4 (N1247, N1239, N361, N575, N788);
not NOT1 (N1248, N1246);
and AND4 (N1249, N1234, N211, N1144, N1167);
not NOT1 (N1250, N1247);
buf BUF1 (N1251, N1221);
not NOT1 (N1252, N1243);
xor XOR2 (N1253, N1251, N156);
nor NOR3 (N1254, N1250, N649, N782);
nor NOR3 (N1255, N1233, N611, N753);
nor NOR3 (N1256, N1244, N64, N228);
nand NAND3 (N1257, N1253, N1255, N404);
nor NOR4 (N1258, N217, N849, N1176, N538);
not NOT1 (N1259, N1241);
nand NAND3 (N1260, N1249, N1184, N136);
not NOT1 (N1261, N1257);
and AND3 (N1262, N1245, N138, N801);
or OR2 (N1263, N1259, N1022);
buf BUF1 (N1264, N1254);
or OR3 (N1265, N1261, N848, N667);
and AND2 (N1266, N1248, N454);
or OR4 (N1267, N1252, N1223, N1029, N1236);
buf BUF1 (N1268, N1260);
nand NAND4 (N1269, N1264, N837, N1215, N1004);
or OR3 (N1270, N1268, N321, N347);
and AND3 (N1271, N1269, N159, N207);
or OR2 (N1272, N1229, N764);
nor NOR2 (N1273, N1270, N994);
xor XOR2 (N1274, N1258, N1166);
xor XOR2 (N1275, N1274, N1184);
and AND3 (N1276, N1262, N555, N695);
or OR3 (N1277, N1275, N972, N328);
not NOT1 (N1278, N1267);
nor NOR4 (N1279, N1273, N61, N1101, N878);
nor NOR4 (N1280, N1265, N1240, N853, N806);
buf BUF1 (N1281, N1266);
xor XOR2 (N1282, N1277, N546);
buf BUF1 (N1283, N1279);
or OR2 (N1284, N1283, N630);
or OR4 (N1285, N1284, N564, N388, N412);
or OR4 (N1286, N1282, N416, N911, N963);
and AND4 (N1287, N1271, N448, N1269, N606);
not NOT1 (N1288, N1286);
buf BUF1 (N1289, N1276);
and AND4 (N1290, N1263, N3, N295, N1001);
buf BUF1 (N1291, N1287);
nand NAND3 (N1292, N1290, N1157, N1263);
xor XOR2 (N1293, N1289, N759);
or OR2 (N1294, N1280, N528);
or OR3 (N1295, N1281, N1146, N878);
buf BUF1 (N1296, N1293);
buf BUF1 (N1297, N1296);
not NOT1 (N1298, N1256);
not NOT1 (N1299, N1285);
and AND4 (N1300, N1288, N632, N212, N101);
and AND4 (N1301, N1278, N161, N1000, N955);
or OR2 (N1302, N1292, N455);
nor NOR3 (N1303, N1301, N958, N36);
nor NOR4 (N1304, N1291, N1297, N131, N992);
not NOT1 (N1305, N89);
buf BUF1 (N1306, N1294);
or OR4 (N1307, N1295, N988, N1041, N513);
buf BUF1 (N1308, N1298);
buf BUF1 (N1309, N1302);
not NOT1 (N1310, N1309);
or OR3 (N1311, N1300, N793, N603);
xor XOR2 (N1312, N1311, N520);
nor NOR2 (N1313, N1304, N1194);
nand NAND4 (N1314, N1306, N1011, N105, N598);
nand NAND4 (N1315, N1312, N49, N904, N294);
buf BUF1 (N1316, N1314);
nor NOR2 (N1317, N1315, N1109);
buf BUF1 (N1318, N1308);
nand NAND2 (N1319, N1307, N97);
nor NOR3 (N1320, N1316, N1241, N583);
xor XOR2 (N1321, N1299, N395);
not NOT1 (N1322, N1310);
and AND2 (N1323, N1321, N777);
buf BUF1 (N1324, N1313);
buf BUF1 (N1325, N1319);
nor NOR4 (N1326, N1317, N239, N589, N457);
xor XOR2 (N1327, N1322, N632);
and AND4 (N1328, N1323, N311, N1095, N434);
and AND2 (N1329, N1320, N677);
nor NOR3 (N1330, N1272, N335, N980);
buf BUF1 (N1331, N1318);
or OR4 (N1332, N1330, N76, N437, N360);
nor NOR4 (N1333, N1325, N1150, N909, N102);
buf BUF1 (N1334, N1303);
not NOT1 (N1335, N1334);
and AND4 (N1336, N1331, N158, N706, N1139);
nand NAND2 (N1337, N1326, N1097);
not NOT1 (N1338, N1329);
nand NAND3 (N1339, N1324, N165, N220);
nand NAND3 (N1340, N1332, N677, N824);
nor NOR3 (N1341, N1333, N1315, N751);
and AND2 (N1342, N1338, N1230);
xor XOR2 (N1343, N1305, N978);
buf BUF1 (N1344, N1327);
or OR3 (N1345, N1328, N1026, N1015);
and AND4 (N1346, N1337, N629, N6, N989);
not NOT1 (N1347, N1345);
or OR4 (N1348, N1347, N1070, N108, N114);
buf BUF1 (N1349, N1341);
nor NOR4 (N1350, N1348, N401, N1009, N614);
xor XOR2 (N1351, N1343, N274);
nor NOR2 (N1352, N1350, N447);
nand NAND3 (N1353, N1344, N542, N1174);
and AND3 (N1354, N1346, N801, N1339);
nand NAND3 (N1355, N908, N595, N525);
nor NOR2 (N1356, N1335, N1262);
or OR3 (N1357, N1356, N994, N1160);
not NOT1 (N1358, N1354);
xor XOR2 (N1359, N1355, N1055);
nand NAND2 (N1360, N1353, N701);
not NOT1 (N1361, N1360);
not NOT1 (N1362, N1361);
not NOT1 (N1363, N1352);
xor XOR2 (N1364, N1342, N1353);
nor NOR4 (N1365, N1364, N1343, N717, N1185);
nand NAND2 (N1366, N1363, N309);
not NOT1 (N1367, N1366);
nor NOR3 (N1368, N1365, N219, N634);
and AND2 (N1369, N1357, N632);
nand NAND2 (N1370, N1340, N182);
and AND3 (N1371, N1368, N927, N312);
nand NAND4 (N1372, N1359, N1337, N1146, N254);
nor NOR2 (N1373, N1370, N898);
and AND4 (N1374, N1336, N54, N771, N1369);
not NOT1 (N1375, N792);
buf BUF1 (N1376, N1358);
nor NOR2 (N1377, N1371, N1083);
xor XOR2 (N1378, N1377, N553);
nand NAND3 (N1379, N1378, N736, N323);
nand NAND3 (N1380, N1376, N1377, N55);
xor XOR2 (N1381, N1349, N742);
not NOT1 (N1382, N1381);
xor XOR2 (N1383, N1375, N1180);
buf BUF1 (N1384, N1379);
nand NAND2 (N1385, N1382, N604);
nor NOR3 (N1386, N1362, N1216, N935);
buf BUF1 (N1387, N1374);
and AND2 (N1388, N1383, N891);
nand NAND3 (N1389, N1388, N26, N354);
nor NOR4 (N1390, N1387, N718, N1146, N611);
xor XOR2 (N1391, N1389, N980);
nor NOR4 (N1392, N1384, N1274, N20, N901);
nand NAND2 (N1393, N1392, N1361);
or OR2 (N1394, N1351, N191);
not NOT1 (N1395, N1393);
nor NOR2 (N1396, N1390, N111);
nand NAND2 (N1397, N1396, N606);
and AND4 (N1398, N1385, N750, N514, N148);
and AND2 (N1399, N1372, N797);
and AND4 (N1400, N1394, N658, N1169, N203);
nand NAND4 (N1401, N1397, N1142, N743, N1138);
nand NAND4 (N1402, N1400, N1165, N741, N556);
nor NOR3 (N1403, N1395, N909, N206);
buf BUF1 (N1404, N1367);
and AND2 (N1405, N1386, N670);
nor NOR3 (N1406, N1373, N426, N685);
not NOT1 (N1407, N1391);
and AND3 (N1408, N1407, N945, N661);
or OR2 (N1409, N1405, N127);
nor NOR2 (N1410, N1402, N616);
nor NOR3 (N1411, N1408, N95, N1236);
nor NOR4 (N1412, N1409, N126, N1275, N142);
nor NOR3 (N1413, N1411, N1249, N1297);
nand NAND3 (N1414, N1398, N642, N255);
nand NAND3 (N1415, N1414, N169, N1194);
nor NOR3 (N1416, N1403, N1281, N1406);
or OR4 (N1417, N974, N682, N702, N556);
xor XOR2 (N1418, N1416, N24);
and AND2 (N1419, N1415, N458);
or OR2 (N1420, N1419, N1320);
xor XOR2 (N1421, N1417, N1141);
nand NAND2 (N1422, N1410, N963);
buf BUF1 (N1423, N1399);
buf BUF1 (N1424, N1422);
or OR3 (N1425, N1423, N181, N138);
or OR2 (N1426, N1401, N282);
buf BUF1 (N1427, N1421);
buf BUF1 (N1428, N1425);
xor XOR2 (N1429, N1418, N346);
or OR2 (N1430, N1413, N650);
not NOT1 (N1431, N1412);
xor XOR2 (N1432, N1380, N1049);
or OR3 (N1433, N1424, N1090, N1346);
nand NAND4 (N1434, N1426, N631, N1409, N962);
nor NOR4 (N1435, N1420, N779, N727, N120);
and AND3 (N1436, N1427, N1105, N440);
not NOT1 (N1437, N1404);
nor NOR2 (N1438, N1434, N1101);
and AND4 (N1439, N1432, N733, N53, N576);
xor XOR2 (N1440, N1428, N619);
nand NAND2 (N1441, N1429, N973);
xor XOR2 (N1442, N1439, N950);
or OR2 (N1443, N1442, N1069);
buf BUF1 (N1444, N1433);
not NOT1 (N1445, N1435);
buf BUF1 (N1446, N1438);
nor NOR4 (N1447, N1444, N36, N1117, N1192);
xor XOR2 (N1448, N1437, N1231);
not NOT1 (N1449, N1448);
nor NOR4 (N1450, N1431, N139, N820, N669);
or OR3 (N1451, N1447, N1073, N1162);
buf BUF1 (N1452, N1441);
nor NOR4 (N1453, N1430, N486, N268, N1195);
nor NOR4 (N1454, N1446, N1392, N1058, N432);
or OR3 (N1455, N1445, N1390, N1032);
buf BUF1 (N1456, N1455);
nand NAND4 (N1457, N1453, N477, N1426, N458);
nor NOR4 (N1458, N1443, N925, N788, N904);
and AND2 (N1459, N1449, N1145);
and AND3 (N1460, N1454, N683, N173);
nor NOR2 (N1461, N1460, N385);
not NOT1 (N1462, N1450);
not NOT1 (N1463, N1461);
buf BUF1 (N1464, N1462);
nor NOR4 (N1465, N1440, N65, N1154, N851);
and AND4 (N1466, N1465, N269, N1227, N547);
nand NAND2 (N1467, N1463, N1046);
and AND3 (N1468, N1436, N1419, N314);
or OR4 (N1469, N1467, N1143, N1426, N1266);
and AND4 (N1470, N1469, N485, N747, N1149);
buf BUF1 (N1471, N1466);
and AND3 (N1472, N1459, N1022, N1232);
not NOT1 (N1473, N1451);
or OR2 (N1474, N1468, N1324);
not NOT1 (N1475, N1464);
xor XOR2 (N1476, N1458, N1009);
or OR3 (N1477, N1473, N1020, N1414);
xor XOR2 (N1478, N1457, N1317);
nand NAND3 (N1479, N1477, N1237, N936);
xor XOR2 (N1480, N1474, N674);
nand NAND4 (N1481, N1475, N382, N666, N226);
and AND4 (N1482, N1470, N942, N540, N19);
xor XOR2 (N1483, N1478, N1406);
or OR2 (N1484, N1476, N131);
xor XOR2 (N1485, N1480, N1197);
or OR2 (N1486, N1483, N544);
or OR2 (N1487, N1484, N547);
and AND4 (N1488, N1471, N1347, N759, N1054);
or OR4 (N1489, N1482, N42, N7, N389);
and AND3 (N1490, N1452, N1414, N8);
nor NOR4 (N1491, N1489, N25, N1031, N11);
xor XOR2 (N1492, N1488, N408);
nor NOR4 (N1493, N1481, N1307, N1279, N70);
or OR2 (N1494, N1486, N150);
not NOT1 (N1495, N1494);
buf BUF1 (N1496, N1493);
not NOT1 (N1497, N1490);
and AND3 (N1498, N1496, N662, N1229);
buf BUF1 (N1499, N1492);
xor XOR2 (N1500, N1456, N287);
nor NOR3 (N1501, N1485, N495, N553);
or OR3 (N1502, N1495, N163, N18);
xor XOR2 (N1503, N1479, N960);
nor NOR4 (N1504, N1487, N1007, N59, N481);
nand NAND4 (N1505, N1504, N1087, N976, N58);
not NOT1 (N1506, N1499);
nor NOR4 (N1507, N1491, N419, N923, N718);
and AND3 (N1508, N1497, N82, N1498);
buf BUF1 (N1509, N1321);
and AND4 (N1510, N1503, N420, N1309, N1143);
or OR2 (N1511, N1510, N565);
buf BUF1 (N1512, N1502);
not NOT1 (N1513, N1472);
or OR2 (N1514, N1509, N1367);
nor NOR3 (N1515, N1501, N1382, N996);
nand NAND2 (N1516, N1513, N41);
nor NOR4 (N1517, N1505, N934, N1210, N1081);
buf BUF1 (N1518, N1514);
xor XOR2 (N1519, N1515, N1136);
buf BUF1 (N1520, N1500);
not NOT1 (N1521, N1519);
nand NAND4 (N1522, N1518, N115, N1403, N640);
nor NOR3 (N1523, N1506, N1185, N1205);
nor NOR3 (N1524, N1511, N217, N760);
buf BUF1 (N1525, N1512);
and AND3 (N1526, N1508, N823, N229);
not NOT1 (N1527, N1523);
nand NAND4 (N1528, N1527, N1414, N676, N226);
xor XOR2 (N1529, N1517, N797);
or OR2 (N1530, N1516, N574);
nor NOR2 (N1531, N1525, N1008);
nor NOR4 (N1532, N1521, N628, N619, N416);
or OR2 (N1533, N1522, N1420);
not NOT1 (N1534, N1529);
not NOT1 (N1535, N1507);
nor NOR4 (N1536, N1532, N524, N699, N1371);
or OR2 (N1537, N1536, N779);
nor NOR3 (N1538, N1524, N473, N17);
not NOT1 (N1539, N1535);
buf BUF1 (N1540, N1520);
xor XOR2 (N1541, N1538, N13);
buf BUF1 (N1542, N1530);
not NOT1 (N1543, N1541);
buf BUF1 (N1544, N1531);
nor NOR4 (N1545, N1534, N16, N584, N264);
or OR3 (N1546, N1539, N682, N846);
not NOT1 (N1547, N1542);
xor XOR2 (N1548, N1545, N72);
xor XOR2 (N1549, N1544, N622);
and AND4 (N1550, N1546, N302, N822, N1394);
nand NAND3 (N1551, N1547, N1474, N232);
nor NOR4 (N1552, N1550, N544, N1539, N335);
nand NAND2 (N1553, N1540, N185);
nand NAND4 (N1554, N1528, N216, N1267, N813);
or OR4 (N1555, N1533, N1090, N1088, N630);
buf BUF1 (N1556, N1554);
xor XOR2 (N1557, N1548, N97);
and AND4 (N1558, N1555, N922, N1127, N368);
nor NOR2 (N1559, N1552, N1106);
xor XOR2 (N1560, N1558, N715);
or OR4 (N1561, N1557, N651, N1043, N767);
buf BUF1 (N1562, N1556);
or OR4 (N1563, N1537, N157, N701, N856);
not NOT1 (N1564, N1553);
not NOT1 (N1565, N1562);
and AND2 (N1566, N1564, N40);
not NOT1 (N1567, N1559);
nor NOR4 (N1568, N1563, N1366, N1390, N944);
buf BUF1 (N1569, N1566);
xor XOR2 (N1570, N1561, N848);
nand NAND3 (N1571, N1560, N760, N92);
xor XOR2 (N1572, N1551, N735);
or OR4 (N1573, N1565, N270, N1440, N1526);
xor XOR2 (N1574, N370, N650);
or OR2 (N1575, N1570, N793);
nor NOR4 (N1576, N1567, N865, N425, N209);
or OR2 (N1577, N1574, N286);
nor NOR3 (N1578, N1572, N690, N888);
not NOT1 (N1579, N1576);
or OR4 (N1580, N1549, N1502, N86, N132);
xor XOR2 (N1581, N1577, N1128);
not NOT1 (N1582, N1579);
not NOT1 (N1583, N1575);
or OR3 (N1584, N1581, N22, N630);
xor XOR2 (N1585, N1571, N1150);
nand NAND4 (N1586, N1569, N1405, N253, N1465);
nor NOR2 (N1587, N1580, N674);
nor NOR4 (N1588, N1587, N285, N390, N617);
nand NAND4 (N1589, N1584, N1461, N146, N143);
and AND3 (N1590, N1573, N1181, N709);
buf BUF1 (N1591, N1568);
and AND2 (N1592, N1582, N238);
nor NOR2 (N1593, N1589, N1358);
buf BUF1 (N1594, N1585);
nor NOR3 (N1595, N1592, N993, N930);
nand NAND2 (N1596, N1586, N583);
not NOT1 (N1597, N1596);
buf BUF1 (N1598, N1583);
nand NAND3 (N1599, N1593, N484, N663);
not NOT1 (N1600, N1591);
and AND2 (N1601, N1543, N302);
xor XOR2 (N1602, N1578, N476);
nor NOR2 (N1603, N1590, N1380);
and AND3 (N1604, N1594, N785, N965);
nand NAND4 (N1605, N1597, N787, N772, N88);
buf BUF1 (N1606, N1602);
or OR3 (N1607, N1603, N6, N1373);
xor XOR2 (N1608, N1599, N2);
and AND2 (N1609, N1598, N156);
not NOT1 (N1610, N1588);
not NOT1 (N1611, N1610);
nand NAND3 (N1612, N1604, N1278, N777);
and AND2 (N1613, N1601, N467);
nand NAND2 (N1614, N1609, N564);
buf BUF1 (N1615, N1612);
nand NAND4 (N1616, N1611, N795, N222, N572);
or OR3 (N1617, N1613, N629, N317);
nor NOR3 (N1618, N1616, N360, N1446);
nand NAND2 (N1619, N1595, N668);
xor XOR2 (N1620, N1600, N105);
nand NAND3 (N1621, N1617, N409, N1033);
buf BUF1 (N1622, N1621);
buf BUF1 (N1623, N1622);
not NOT1 (N1624, N1614);
and AND2 (N1625, N1618, N1558);
xor XOR2 (N1626, N1620, N708);
xor XOR2 (N1627, N1625, N888);
and AND3 (N1628, N1615, N1326, N495);
xor XOR2 (N1629, N1624, N834);
buf BUF1 (N1630, N1623);
xor XOR2 (N1631, N1605, N278);
buf BUF1 (N1632, N1629);
or OR3 (N1633, N1607, N1515, N700);
and AND3 (N1634, N1633, N242, N1351);
nor NOR4 (N1635, N1626, N454, N1420, N1428);
nand NAND3 (N1636, N1628, N641, N205);
nand NAND2 (N1637, N1608, N958);
not NOT1 (N1638, N1627);
not NOT1 (N1639, N1637);
nor NOR4 (N1640, N1635, N348, N790, N590);
and AND4 (N1641, N1634, N709, N794, N1035);
buf BUF1 (N1642, N1606);
not NOT1 (N1643, N1636);
nand NAND3 (N1644, N1619, N456, N1484);
or OR2 (N1645, N1632, N516);
not NOT1 (N1646, N1630);
and AND3 (N1647, N1641, N1600, N536);
buf BUF1 (N1648, N1640);
or OR2 (N1649, N1638, N215);
not NOT1 (N1650, N1639);
buf BUF1 (N1651, N1650);
nand NAND2 (N1652, N1642, N1462);
not NOT1 (N1653, N1631);
xor XOR2 (N1654, N1651, N916);
nor NOR3 (N1655, N1648, N349, N1519);
buf BUF1 (N1656, N1654);
xor XOR2 (N1657, N1655, N433);
xor XOR2 (N1658, N1657, N1403);
buf BUF1 (N1659, N1658);
not NOT1 (N1660, N1649);
nor NOR3 (N1661, N1646, N1044, N1070);
buf BUF1 (N1662, N1660);
or OR3 (N1663, N1644, N922, N868);
nor NOR4 (N1664, N1643, N888, N1051, N291);
nand NAND3 (N1665, N1656, N795, N1265);
xor XOR2 (N1666, N1659, N1621);
nand NAND2 (N1667, N1652, N770);
buf BUF1 (N1668, N1647);
xor XOR2 (N1669, N1666, N1662);
nand NAND3 (N1670, N1073, N752, N1231);
or OR4 (N1671, N1661, N581, N554, N258);
buf BUF1 (N1672, N1664);
and AND2 (N1673, N1645, N399);
or OR2 (N1674, N1667, N964);
not NOT1 (N1675, N1653);
xor XOR2 (N1676, N1675, N373);
buf BUF1 (N1677, N1665);
buf BUF1 (N1678, N1663);
nand NAND3 (N1679, N1668, N1586, N1444);
and AND2 (N1680, N1669, N299);
or OR4 (N1681, N1676, N330, N589, N1370);
buf BUF1 (N1682, N1671);
or OR3 (N1683, N1673, N1409, N410);
buf BUF1 (N1684, N1677);
xor XOR2 (N1685, N1684, N936);
not NOT1 (N1686, N1683);
not NOT1 (N1687, N1682);
xor XOR2 (N1688, N1678, N967);
or OR4 (N1689, N1686, N976, N1249, N376);
buf BUF1 (N1690, N1688);
and AND3 (N1691, N1681, N268, N151);
xor XOR2 (N1692, N1685, N1296);
nand NAND2 (N1693, N1679, N927);
nor NOR3 (N1694, N1670, N1356, N978);
xor XOR2 (N1695, N1674, N1177);
nor NOR4 (N1696, N1695, N689, N451, N863);
nor NOR2 (N1697, N1692, N711);
nor NOR2 (N1698, N1697, N1190);
nand NAND4 (N1699, N1690, N720, N806, N1407);
nand NAND4 (N1700, N1693, N1399, N175, N867);
or OR4 (N1701, N1672, N1359, N1307, N927);
xor XOR2 (N1702, N1699, N316);
and AND3 (N1703, N1696, N607, N1228);
buf BUF1 (N1704, N1691);
or OR4 (N1705, N1694, N864, N1147, N1125);
and AND4 (N1706, N1698, N812, N466, N1333);
and AND2 (N1707, N1689, N1174);
xor XOR2 (N1708, N1687, N305);
xor XOR2 (N1709, N1703, N1583);
or OR3 (N1710, N1701, N58, N853);
or OR2 (N1711, N1700, N907);
nor NOR2 (N1712, N1707, N668);
nand NAND4 (N1713, N1709, N1152, N343, N446);
nand NAND3 (N1714, N1705, N496, N532);
nand NAND3 (N1715, N1706, N1259, N622);
not NOT1 (N1716, N1680);
not NOT1 (N1717, N1704);
or OR2 (N1718, N1716, N743);
buf BUF1 (N1719, N1711);
xor XOR2 (N1720, N1713, N1264);
not NOT1 (N1721, N1718);
not NOT1 (N1722, N1717);
and AND3 (N1723, N1714, N1438, N1455);
or OR4 (N1724, N1723, N198, N1140, N290);
or OR4 (N1725, N1724, N659, N1158, N1616);
nor NOR3 (N1726, N1720, N1303, N117);
xor XOR2 (N1727, N1719, N209);
xor XOR2 (N1728, N1722, N1304);
and AND2 (N1729, N1708, N351);
nand NAND3 (N1730, N1725, N469, N1570);
or OR4 (N1731, N1702, N1300, N345, N546);
buf BUF1 (N1732, N1710);
xor XOR2 (N1733, N1721, N1622);
buf BUF1 (N1734, N1727);
xor XOR2 (N1735, N1733, N236);
nand NAND3 (N1736, N1712, N220, N1106);
buf BUF1 (N1737, N1726);
not NOT1 (N1738, N1736);
nand NAND4 (N1739, N1731, N603, N849, N1000);
nor NOR3 (N1740, N1739, N978, N1399);
xor XOR2 (N1741, N1738, N598);
nor NOR2 (N1742, N1735, N1716);
nand NAND4 (N1743, N1741, N1196, N1367, N342);
or OR3 (N1744, N1729, N162, N793);
buf BUF1 (N1745, N1743);
nand NAND2 (N1746, N1744, N1485);
nand NAND4 (N1747, N1745, N503, N660, N1315);
buf BUF1 (N1748, N1728);
xor XOR2 (N1749, N1747, N345);
not NOT1 (N1750, N1734);
xor XOR2 (N1751, N1715, N353);
or OR4 (N1752, N1751, N654, N1421, N1742);
and AND2 (N1753, N136, N461);
or OR4 (N1754, N1746, N1066, N1152, N1185);
or OR2 (N1755, N1740, N1399);
and AND3 (N1756, N1750, N114, N1526);
not NOT1 (N1757, N1752);
xor XOR2 (N1758, N1730, N967);
buf BUF1 (N1759, N1754);
buf BUF1 (N1760, N1755);
or OR3 (N1761, N1753, N381, N412);
and AND3 (N1762, N1761, N1737, N183);
xor XOR2 (N1763, N140, N1476);
and AND2 (N1764, N1763, N177);
or OR4 (N1765, N1756, N1286, N549, N892);
nand NAND2 (N1766, N1757, N327);
or OR2 (N1767, N1766, N1577);
or OR2 (N1768, N1748, N686);
and AND4 (N1769, N1768, N943, N1119, N1743);
nor NOR3 (N1770, N1760, N1263, N1447);
nand NAND3 (N1771, N1758, N1516, N454);
or OR2 (N1772, N1765, N1289);
xor XOR2 (N1773, N1771, N1604);
or OR3 (N1774, N1773, N1404, N559);
not NOT1 (N1775, N1774);
nand NAND4 (N1776, N1775, N526, N1662, N1759);
nand NAND4 (N1777, N690, N1098, N866, N1251);
not NOT1 (N1778, N1732);
nand NAND2 (N1779, N1764, N484);
nand NAND4 (N1780, N1762, N1680, N1418, N490);
nand NAND2 (N1781, N1770, N44);
buf BUF1 (N1782, N1781);
nor NOR3 (N1783, N1769, N1335, N860);
or OR2 (N1784, N1767, N44);
nor NOR3 (N1785, N1749, N1146, N1701);
and AND4 (N1786, N1777, N1753, N875, N47);
or OR3 (N1787, N1780, N414, N1607);
nand NAND2 (N1788, N1787, N1334);
or OR3 (N1789, N1779, N608, N865);
nand NAND4 (N1790, N1776, N385, N636, N349);
and AND3 (N1791, N1790, N855, N398);
and AND3 (N1792, N1786, N1233, N399);
nand NAND2 (N1793, N1784, N495);
and AND2 (N1794, N1778, N541);
and AND4 (N1795, N1791, N837, N49, N1153);
buf BUF1 (N1796, N1795);
or OR2 (N1797, N1782, N811);
xor XOR2 (N1798, N1783, N712);
nor NOR4 (N1799, N1789, N805, N1062, N1590);
or OR2 (N1800, N1797, N649);
not NOT1 (N1801, N1796);
nor NOR4 (N1802, N1801, N282, N918, N361);
nand NAND3 (N1803, N1799, N1451, N212);
buf BUF1 (N1804, N1794);
and AND2 (N1805, N1798, N519);
or OR3 (N1806, N1803, N850, N1719);
nor NOR3 (N1807, N1804, N1266, N574);
not NOT1 (N1808, N1792);
buf BUF1 (N1809, N1805);
buf BUF1 (N1810, N1793);
nor NOR3 (N1811, N1772, N1079, N1570);
xor XOR2 (N1812, N1811, N1180);
nor NOR3 (N1813, N1812, N1707, N631);
xor XOR2 (N1814, N1802, N1711);
nand NAND2 (N1815, N1807, N1472);
buf BUF1 (N1816, N1800);
and AND3 (N1817, N1788, N1756, N1449);
buf BUF1 (N1818, N1785);
xor XOR2 (N1819, N1818, N1395);
not NOT1 (N1820, N1817);
not NOT1 (N1821, N1815);
buf BUF1 (N1822, N1819);
and AND2 (N1823, N1813, N1325);
and AND2 (N1824, N1814, N1463);
nand NAND2 (N1825, N1821, N1601);
xor XOR2 (N1826, N1809, N1780);
not NOT1 (N1827, N1822);
buf BUF1 (N1828, N1808);
not NOT1 (N1829, N1820);
nor NOR3 (N1830, N1825, N314, N1687);
nor NOR3 (N1831, N1830, N1401, N932);
xor XOR2 (N1832, N1826, N615);
nand NAND3 (N1833, N1831, N866, N822);
nor NOR3 (N1834, N1824, N1597, N305);
and AND4 (N1835, N1806, N1610, N1759, N1407);
xor XOR2 (N1836, N1835, N766);
or OR3 (N1837, N1834, N279, N1551);
not NOT1 (N1838, N1828);
not NOT1 (N1839, N1829);
buf BUF1 (N1840, N1839);
not NOT1 (N1841, N1840);
xor XOR2 (N1842, N1832, N1121);
and AND4 (N1843, N1816, N401, N1511, N26);
xor XOR2 (N1844, N1833, N1279);
or OR2 (N1845, N1837, N1597);
and AND4 (N1846, N1844, N551, N1048, N1455);
nand NAND2 (N1847, N1838, N182);
nand NAND3 (N1848, N1846, N1399, N1615);
or OR4 (N1849, N1843, N1193, N364, N1330);
nor NOR3 (N1850, N1836, N727, N1829);
or OR3 (N1851, N1848, N1561, N1346);
nor NOR2 (N1852, N1823, N1334);
not NOT1 (N1853, N1810);
not NOT1 (N1854, N1849);
or OR2 (N1855, N1841, N137);
nor NOR2 (N1856, N1854, N1341);
nor NOR3 (N1857, N1842, N450, N552);
xor XOR2 (N1858, N1827, N1658);
not NOT1 (N1859, N1856);
nor NOR4 (N1860, N1847, N1730, N698, N1754);
not NOT1 (N1861, N1850);
buf BUF1 (N1862, N1858);
buf BUF1 (N1863, N1860);
not NOT1 (N1864, N1852);
not NOT1 (N1865, N1864);
not NOT1 (N1866, N1853);
nor NOR3 (N1867, N1859, N410, N827);
buf BUF1 (N1868, N1855);
or OR3 (N1869, N1845, N299, N292);
nand NAND3 (N1870, N1851, N271, N281);
nor NOR2 (N1871, N1867, N1673);
buf BUF1 (N1872, N1865);
and AND2 (N1873, N1862, N684);
buf BUF1 (N1874, N1863);
nand NAND2 (N1875, N1861, N528);
xor XOR2 (N1876, N1872, N604);
nor NOR3 (N1877, N1866, N1181, N699);
xor XOR2 (N1878, N1873, N714);
nor NOR2 (N1879, N1876, N1019);
buf BUF1 (N1880, N1877);
nand NAND4 (N1881, N1878, N1329, N208, N171);
buf BUF1 (N1882, N1880);
nor NOR3 (N1883, N1868, N1664, N424);
xor XOR2 (N1884, N1870, N1605);
xor XOR2 (N1885, N1882, N232);
xor XOR2 (N1886, N1884, N1311);
buf BUF1 (N1887, N1875);
not NOT1 (N1888, N1879);
buf BUF1 (N1889, N1869);
and AND4 (N1890, N1886, N1841, N1654, N1107);
xor XOR2 (N1891, N1883, N612);
buf BUF1 (N1892, N1881);
xor XOR2 (N1893, N1890, N959);
nor NOR3 (N1894, N1893, N383, N275);
not NOT1 (N1895, N1891);
xor XOR2 (N1896, N1892, N1131);
or OR2 (N1897, N1871, N1414);
nand NAND2 (N1898, N1894, N457);
or OR4 (N1899, N1857, N368, N1894, N768);
and AND2 (N1900, N1874, N1388);
or OR2 (N1901, N1888, N79);
or OR4 (N1902, N1899, N1381, N863, N1352);
or OR3 (N1903, N1897, N164, N1756);
xor XOR2 (N1904, N1889, N1191);
buf BUF1 (N1905, N1901);
buf BUF1 (N1906, N1904);
buf BUF1 (N1907, N1902);
and AND3 (N1908, N1900, N699, N1101);
and AND2 (N1909, N1908, N210);
buf BUF1 (N1910, N1898);
and AND4 (N1911, N1895, N1034, N1476, N887);
nand NAND2 (N1912, N1896, N62);
nor NOR2 (N1913, N1885, N1023);
and AND4 (N1914, N1912, N1810, N1905, N1147);
xor XOR2 (N1915, N1552, N946);
nor NOR4 (N1916, N1887, N495, N337, N1264);
xor XOR2 (N1917, N1916, N83);
nand NAND2 (N1918, N1917, N1156);
and AND3 (N1919, N1909, N1551, N753);
nor NOR4 (N1920, N1907, N1574, N174, N742);
nand NAND4 (N1921, N1915, N108, N164, N1298);
xor XOR2 (N1922, N1918, N1519);
xor XOR2 (N1923, N1914, N704);
nor NOR4 (N1924, N1906, N1699, N994, N136);
nand NAND3 (N1925, N1920, N1751, N1192);
and AND2 (N1926, N1923, N1080);
or OR3 (N1927, N1926, N1635, N914);
nor NOR4 (N1928, N1911, N1656, N415, N1617);
or OR2 (N1929, N1924, N246);
and AND2 (N1930, N1910, N462);
nand NAND2 (N1931, N1929, N1423);
xor XOR2 (N1932, N1928, N866);
and AND3 (N1933, N1919, N1516, N379);
xor XOR2 (N1934, N1927, N1190);
xor XOR2 (N1935, N1921, N1758);
or OR3 (N1936, N1903, N1399, N800);
xor XOR2 (N1937, N1936, N1360);
xor XOR2 (N1938, N1933, N991);
nor NOR4 (N1939, N1938, N1386, N1252, N205);
not NOT1 (N1940, N1939);
buf BUF1 (N1941, N1931);
or OR4 (N1942, N1925, N497, N1037, N391);
nand NAND4 (N1943, N1932, N285, N1705, N1864);
or OR4 (N1944, N1934, N1699, N425, N352);
buf BUF1 (N1945, N1941);
buf BUF1 (N1946, N1942);
and AND4 (N1947, N1946, N1622, N1796, N1751);
not NOT1 (N1948, N1913);
xor XOR2 (N1949, N1945, N1138);
and AND3 (N1950, N1943, N1939, N915);
xor XOR2 (N1951, N1944, N1767);
not NOT1 (N1952, N1940);
or OR2 (N1953, N1951, N370);
buf BUF1 (N1954, N1949);
xor XOR2 (N1955, N1952, N1679);
and AND3 (N1956, N1954, N917, N239);
nor NOR2 (N1957, N1955, N598);
or OR4 (N1958, N1948, N1674, N338, N953);
or OR2 (N1959, N1947, N654);
nor NOR4 (N1960, N1958, N1479, N517, N1905);
nor NOR2 (N1961, N1953, N1267);
and AND2 (N1962, N1957, N453);
nor NOR2 (N1963, N1959, N1421);
and AND3 (N1964, N1962, N516, N313);
nor NOR3 (N1965, N1963, N435, N1512);
nor NOR4 (N1966, N1961, N79, N539, N1641);
buf BUF1 (N1967, N1956);
or OR3 (N1968, N1950, N1623, N713);
or OR2 (N1969, N1937, N1035);
buf BUF1 (N1970, N1930);
or OR3 (N1971, N1960, N182, N1127);
buf BUF1 (N1972, N1964);
buf BUF1 (N1973, N1966);
or OR4 (N1974, N1970, N775, N1653, N71);
or OR2 (N1975, N1974, N1221);
xor XOR2 (N1976, N1935, N958);
or OR4 (N1977, N1922, N340, N1032, N12);
or OR3 (N1978, N1972, N605, N1659);
nand NAND4 (N1979, N1975, N1945, N1511, N1440);
and AND3 (N1980, N1976, N1217, N1445);
and AND2 (N1981, N1967, N1210);
nor NOR4 (N1982, N1965, N1036, N1409, N1506);
nor NOR3 (N1983, N1969, N1578, N404);
and AND2 (N1984, N1980, N1432);
xor XOR2 (N1985, N1978, N975);
xor XOR2 (N1986, N1977, N613);
xor XOR2 (N1987, N1981, N412);
not NOT1 (N1988, N1979);
buf BUF1 (N1989, N1984);
nor NOR3 (N1990, N1989, N1837, N25);
nand NAND3 (N1991, N1986, N1148, N1647);
and AND3 (N1992, N1988, N885, N1303);
and AND2 (N1993, N1971, N37);
and AND2 (N1994, N1987, N884);
nand NAND2 (N1995, N1983, N1367);
buf BUF1 (N1996, N1973);
and AND2 (N1997, N1993, N1425);
not NOT1 (N1998, N1982);
and AND4 (N1999, N1994, N1791, N152, N124);
not NOT1 (N2000, N1999);
xor XOR2 (N2001, N1997, N1053);
buf BUF1 (N2002, N2000);
xor XOR2 (N2003, N1985, N1397);
and AND2 (N2004, N1990, N374);
and AND3 (N2005, N1991, N736, N16);
or OR2 (N2006, N1968, N1092);
xor XOR2 (N2007, N2003, N1118);
not NOT1 (N2008, N2001);
and AND3 (N2009, N2004, N245, N286);
buf BUF1 (N2010, N2007);
and AND4 (N2011, N2009, N719, N512, N579);
and AND4 (N2012, N2005, N1036, N1460, N685);
nor NOR2 (N2013, N1996, N351);
not NOT1 (N2014, N2012);
xor XOR2 (N2015, N2014, N1351);
or OR2 (N2016, N2010, N279);
buf BUF1 (N2017, N1995);
buf BUF1 (N2018, N2008);
endmodule