// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N2008,N1982,N2013,N2015,N2014,N1986,N2012,N2016,N2018,N2019;

or OR4 (N20, N15, N15, N17, N1);
nand NAND2 (N21, N1, N19);
xor XOR2 (N22, N3, N9);
not NOT1 (N23, N8);
or OR4 (N24, N5, N14, N19, N18);
and AND2 (N25, N7, N5);
and AND3 (N26, N11, N25, N17);
buf BUF1 (N27, N26);
nor NOR4 (N28, N19, N14, N4, N10);
xor XOR2 (N29, N19, N7);
buf BUF1 (N30, N17);
buf BUF1 (N31, N10);
buf BUF1 (N32, N28);
nand NAND3 (N33, N22, N3, N18);
xor XOR2 (N34, N24, N24);
and AND4 (N35, N23, N2, N5, N22);
or OR3 (N36, N33, N5, N11);
and AND4 (N37, N31, N7, N32, N12);
nor NOR2 (N38, N7, N27);
buf BUF1 (N39, N30);
nand NAND4 (N40, N27, N8, N10, N3);
xor XOR2 (N41, N38, N8);
nor NOR3 (N42, N29, N15, N14);
xor XOR2 (N43, N21, N23);
or OR2 (N44, N37, N32);
nor NOR4 (N45, N35, N18, N2, N31);
nand NAND4 (N46, N40, N35, N27, N31);
or OR3 (N47, N45, N32, N17);
not NOT1 (N48, N47);
not NOT1 (N49, N46);
nor NOR3 (N50, N42, N4, N12);
not NOT1 (N51, N39);
buf BUF1 (N52, N41);
and AND4 (N53, N51, N45, N14, N20);
and AND4 (N54, N3, N38, N7, N4);
buf BUF1 (N55, N36);
buf BUF1 (N56, N49);
nor NOR4 (N57, N44, N35, N31, N4);
or OR3 (N58, N34, N38, N36);
and AND3 (N59, N54, N34, N37);
xor XOR2 (N60, N53, N29);
nand NAND4 (N61, N52, N43, N50, N13);
buf BUF1 (N62, N41);
nand NAND4 (N63, N21, N24, N13, N13);
not NOT1 (N64, N48);
nand NAND2 (N65, N61, N31);
buf BUF1 (N66, N56);
nand NAND3 (N67, N65, N48, N39);
or OR4 (N68, N58, N46, N57, N26);
or OR2 (N69, N41, N66);
or OR3 (N70, N16, N19, N27);
and AND3 (N71, N62, N56, N49);
nand NAND3 (N72, N69, N13, N49);
xor XOR2 (N73, N59, N66);
or OR3 (N74, N70, N27, N48);
and AND2 (N75, N64, N56);
buf BUF1 (N76, N55);
nand NAND4 (N77, N74, N70, N46, N61);
or OR3 (N78, N73, N18, N18);
not NOT1 (N79, N75);
xor XOR2 (N80, N77, N39);
and AND4 (N81, N60, N78, N68, N29);
nand NAND4 (N82, N40, N63, N72, N26);
nor NOR2 (N83, N48, N17);
and AND4 (N84, N17, N66, N76, N43);
not NOT1 (N85, N73);
or OR3 (N86, N82, N42, N67);
nor NOR2 (N87, N62, N29);
or OR2 (N88, N75, N83);
xor XOR2 (N89, N39, N17);
not NOT1 (N90, N80);
nand NAND4 (N91, N71, N73, N11, N8);
and AND2 (N92, N86, N14);
nand NAND2 (N93, N87, N56);
and AND4 (N94, N85, N78, N8, N83);
not NOT1 (N95, N88);
nand NAND4 (N96, N93, N87, N7, N62);
buf BUF1 (N97, N90);
buf BUF1 (N98, N97);
not NOT1 (N99, N84);
buf BUF1 (N100, N91);
nand NAND2 (N101, N89, N22);
buf BUF1 (N102, N101);
not NOT1 (N103, N94);
or OR3 (N104, N95, N43, N98);
xor XOR2 (N105, N24, N25);
nor NOR3 (N106, N92, N68, N90);
buf BUF1 (N107, N104);
nor NOR3 (N108, N103, N44, N30);
nor NOR2 (N109, N108, N84);
not NOT1 (N110, N109);
nor NOR4 (N111, N106, N48, N63, N81);
nand NAND2 (N112, N60, N65);
or OR4 (N113, N96, N54, N60, N40);
nor NOR2 (N114, N107, N12);
not NOT1 (N115, N110);
nand NAND3 (N116, N105, N85, N52);
buf BUF1 (N117, N111);
and AND4 (N118, N113, N63, N117, N49);
buf BUF1 (N119, N61);
and AND3 (N120, N102, N20, N39);
buf BUF1 (N121, N118);
and AND4 (N122, N79, N53, N24, N112);
and AND2 (N123, N34, N27);
xor XOR2 (N124, N122, N85);
and AND4 (N125, N116, N18, N95, N24);
xor XOR2 (N126, N121, N18);
not NOT1 (N127, N120);
not NOT1 (N128, N114);
nor NOR4 (N129, N99, N5, N89, N27);
buf BUF1 (N130, N123);
nand NAND3 (N131, N100, N106, N77);
or OR4 (N132, N127, N27, N79, N44);
nand NAND3 (N133, N126, N45, N41);
nand NAND2 (N134, N130, N5);
nor NOR3 (N135, N125, N95, N15);
not NOT1 (N136, N132);
nor NOR2 (N137, N129, N84);
not NOT1 (N138, N136);
not NOT1 (N139, N131);
not NOT1 (N140, N128);
nand NAND4 (N141, N134, N23, N64, N45);
xor XOR2 (N142, N124, N96);
not NOT1 (N143, N139);
nand NAND3 (N144, N119, N19, N76);
nor NOR2 (N145, N133, N97);
nor NOR4 (N146, N135, N75, N24, N77);
and AND3 (N147, N142, N51, N26);
nor NOR3 (N148, N115, N63, N4);
and AND2 (N149, N138, N48);
xor XOR2 (N150, N140, N92);
nand NAND4 (N151, N144, N10, N4, N133);
xor XOR2 (N152, N151, N9);
and AND2 (N153, N146, N39);
and AND4 (N154, N153, N19, N52, N54);
nor NOR2 (N155, N148, N90);
buf BUF1 (N156, N154);
not NOT1 (N157, N143);
nor NOR4 (N158, N150, N105, N16, N94);
xor XOR2 (N159, N155, N146);
not NOT1 (N160, N157);
nand NAND3 (N161, N158, N74, N67);
and AND2 (N162, N141, N86);
or OR3 (N163, N137, N154, N53);
not NOT1 (N164, N162);
and AND4 (N165, N161, N61, N21, N61);
nand NAND2 (N166, N165, N149);
or OR2 (N167, N82, N20);
xor XOR2 (N168, N164, N118);
buf BUF1 (N169, N166);
not NOT1 (N170, N152);
nand NAND3 (N171, N169, N24, N26);
nand NAND4 (N172, N168, N21, N29, N45);
and AND3 (N173, N145, N92, N162);
or OR2 (N174, N171, N124);
nand NAND4 (N175, N167, N95, N140, N84);
or OR2 (N176, N172, N41);
xor XOR2 (N177, N159, N3);
buf BUF1 (N178, N163);
nand NAND4 (N179, N173, N105, N53, N58);
not NOT1 (N180, N156);
xor XOR2 (N181, N174, N22);
buf BUF1 (N182, N177);
or OR4 (N183, N181, N64, N69, N98);
and AND3 (N184, N160, N165, N28);
nand NAND3 (N185, N182, N84, N85);
nand NAND4 (N186, N184, N154, N127, N153);
nand NAND4 (N187, N176, N63, N35, N42);
buf BUF1 (N188, N186);
not NOT1 (N189, N183);
xor XOR2 (N190, N187, N66);
xor XOR2 (N191, N190, N60);
or OR2 (N192, N180, N121);
nand NAND3 (N193, N192, N50, N63);
buf BUF1 (N194, N189);
xor XOR2 (N195, N188, N126);
not NOT1 (N196, N185);
not NOT1 (N197, N147);
not NOT1 (N198, N178);
xor XOR2 (N199, N193, N169);
buf BUF1 (N200, N175);
nor NOR4 (N201, N195, N113, N104, N108);
and AND2 (N202, N191, N124);
and AND2 (N203, N170, N76);
not NOT1 (N204, N199);
or OR3 (N205, N198, N156, N112);
or OR2 (N206, N194, N121);
nor NOR4 (N207, N205, N107, N181, N38);
nand NAND3 (N208, N200, N159, N100);
or OR4 (N209, N197, N68, N203, N60);
and AND2 (N210, N104, N61);
not NOT1 (N211, N196);
not NOT1 (N212, N201);
xor XOR2 (N213, N211, N100);
nor NOR2 (N214, N213, N168);
nand NAND2 (N215, N214, N92);
xor XOR2 (N216, N212, N7);
buf BUF1 (N217, N209);
xor XOR2 (N218, N210, N6);
xor XOR2 (N219, N216, N212);
buf BUF1 (N220, N218);
or OR2 (N221, N217, N154);
nand NAND4 (N222, N215, N56, N119, N178);
buf BUF1 (N223, N219);
nand NAND4 (N224, N179, N182, N18, N45);
and AND3 (N225, N220, N174, N13);
nor NOR3 (N226, N225, N149, N128);
xor XOR2 (N227, N221, N185);
nor NOR2 (N228, N226, N225);
buf BUF1 (N229, N202);
and AND4 (N230, N206, N205, N159, N88);
buf BUF1 (N231, N223);
and AND2 (N232, N224, N208);
and AND3 (N233, N31, N13, N71);
nand NAND4 (N234, N230, N97, N114, N231);
xor XOR2 (N235, N50, N90);
or OR2 (N236, N204, N210);
nor NOR3 (N237, N233, N230, N53);
nor NOR2 (N238, N222, N131);
or OR3 (N239, N234, N63, N182);
or OR2 (N240, N207, N25);
nor NOR4 (N241, N235, N176, N218, N5);
nand NAND3 (N242, N228, N40, N79);
and AND4 (N243, N241, N164, N54, N146);
xor XOR2 (N244, N242, N25);
xor XOR2 (N245, N240, N117);
and AND3 (N246, N237, N7, N174);
not NOT1 (N247, N229);
nor NOR3 (N248, N246, N43, N111);
and AND4 (N249, N227, N6, N81, N24);
nand NAND4 (N250, N232, N43, N217, N232);
not NOT1 (N251, N238);
and AND4 (N252, N236, N107, N146, N182);
nand NAND3 (N253, N245, N132, N152);
nand NAND2 (N254, N244, N101);
and AND4 (N255, N251, N12, N37, N175);
or OR2 (N256, N255, N203);
buf BUF1 (N257, N256);
and AND3 (N258, N253, N141, N193);
buf BUF1 (N259, N250);
or OR4 (N260, N254, N218, N206, N149);
not NOT1 (N261, N258);
or OR2 (N262, N252, N163);
and AND2 (N263, N249, N5);
nor NOR2 (N264, N262, N160);
buf BUF1 (N265, N239);
xor XOR2 (N266, N243, N176);
not NOT1 (N267, N261);
nor NOR3 (N268, N265, N144, N24);
xor XOR2 (N269, N263, N28);
or OR3 (N270, N247, N120, N74);
nor NOR4 (N271, N248, N129, N1, N110);
xor XOR2 (N272, N270, N124);
or OR3 (N273, N264, N61, N118);
buf BUF1 (N274, N259);
or OR3 (N275, N268, N125, N61);
or OR4 (N276, N274, N122, N129, N54);
xor XOR2 (N277, N271, N46);
nor NOR3 (N278, N276, N266, N27);
or OR3 (N279, N56, N275, N272);
nand NAND2 (N280, N33, N5);
buf BUF1 (N281, N7);
not NOT1 (N282, N277);
xor XOR2 (N283, N273, N80);
or OR3 (N284, N283, N154, N170);
xor XOR2 (N285, N260, N208);
and AND2 (N286, N269, N183);
xor XOR2 (N287, N280, N85);
or OR2 (N288, N287, N125);
not NOT1 (N289, N282);
buf BUF1 (N290, N285);
buf BUF1 (N291, N286);
xor XOR2 (N292, N289, N40);
not NOT1 (N293, N288);
xor XOR2 (N294, N267, N209);
nand NAND3 (N295, N292, N98, N183);
xor XOR2 (N296, N281, N241);
buf BUF1 (N297, N293);
buf BUF1 (N298, N279);
buf BUF1 (N299, N298);
xor XOR2 (N300, N257, N253);
not NOT1 (N301, N295);
nor NOR2 (N302, N290, N272);
not NOT1 (N303, N301);
nor NOR3 (N304, N278, N127, N253);
not NOT1 (N305, N291);
and AND4 (N306, N296, N142, N63, N149);
not NOT1 (N307, N304);
or OR3 (N308, N300, N78, N120);
and AND3 (N309, N297, N64, N140);
nand NAND3 (N310, N302, N212, N255);
nand NAND2 (N311, N284, N82);
or OR4 (N312, N311, N14, N41, N233);
xor XOR2 (N313, N308, N12);
nor NOR4 (N314, N310, N171, N77, N200);
and AND2 (N315, N307, N293);
nand NAND3 (N316, N309, N17, N40);
nor NOR2 (N317, N313, N97);
buf BUF1 (N318, N315);
buf BUF1 (N319, N294);
or OR2 (N320, N316, N104);
or OR3 (N321, N306, N169, N320);
not NOT1 (N322, N255);
and AND4 (N323, N299, N67, N110, N240);
nor NOR3 (N324, N321, N215, N212);
and AND2 (N325, N319, N62);
or OR4 (N326, N323, N81, N305, N303);
buf BUF1 (N327, N119);
buf BUF1 (N328, N84);
or OR3 (N329, N322, N236, N171);
xor XOR2 (N330, N314, N70);
and AND3 (N331, N326, N46, N162);
xor XOR2 (N332, N317, N151);
nor NOR4 (N333, N329, N95, N71, N28);
nor NOR3 (N334, N327, N36, N59);
not NOT1 (N335, N328);
not NOT1 (N336, N334);
xor XOR2 (N337, N325, N279);
buf BUF1 (N338, N318);
nor NOR2 (N339, N335, N171);
or OR3 (N340, N339, N137, N179);
or OR2 (N341, N324, N322);
or OR2 (N342, N332, N232);
or OR3 (N343, N333, N80, N82);
nand NAND3 (N344, N343, N53, N29);
not NOT1 (N345, N340);
nand NAND4 (N346, N341, N326, N9, N266);
nor NOR2 (N347, N336, N188);
nand NAND3 (N348, N346, N194, N344);
or OR4 (N349, N211, N195, N240, N52);
nand NAND4 (N350, N312, N271, N308, N190);
xor XOR2 (N351, N331, N102);
or OR4 (N352, N337, N16, N43, N42);
nand NAND3 (N353, N349, N129, N349);
xor XOR2 (N354, N352, N229);
nor NOR2 (N355, N348, N185);
and AND2 (N356, N355, N71);
and AND4 (N357, N342, N337, N168, N128);
not NOT1 (N358, N351);
nand NAND2 (N359, N353, N4);
xor XOR2 (N360, N354, N162);
xor XOR2 (N361, N338, N145);
nand NAND2 (N362, N359, N292);
buf BUF1 (N363, N347);
nand NAND3 (N364, N330, N21, N179);
or OR3 (N365, N362, N58, N241);
and AND3 (N366, N350, N114, N285);
or OR4 (N367, N363, N118, N19, N64);
not NOT1 (N368, N364);
buf BUF1 (N369, N367);
and AND2 (N370, N369, N222);
or OR4 (N371, N370, N240, N317, N23);
not NOT1 (N372, N357);
or OR4 (N373, N371, N9, N123, N69);
not NOT1 (N374, N361);
xor XOR2 (N375, N372, N58);
buf BUF1 (N376, N356);
not NOT1 (N377, N376);
not NOT1 (N378, N345);
xor XOR2 (N379, N375, N346);
xor XOR2 (N380, N368, N51);
xor XOR2 (N381, N380, N155);
or OR3 (N382, N366, N257, N378);
nor NOR2 (N383, N382, N235);
nand NAND4 (N384, N300, N182, N342, N243);
and AND2 (N385, N383, N108);
nand NAND3 (N386, N374, N153, N151);
or OR3 (N387, N384, N15, N83);
nand NAND3 (N388, N373, N219, N207);
buf BUF1 (N389, N386);
xor XOR2 (N390, N358, N51);
buf BUF1 (N391, N377);
and AND2 (N392, N390, N349);
xor XOR2 (N393, N381, N368);
buf BUF1 (N394, N379);
not NOT1 (N395, N391);
and AND3 (N396, N395, N54, N29);
or OR2 (N397, N360, N122);
xor XOR2 (N398, N396, N85);
or OR4 (N399, N398, N204, N55, N106);
not NOT1 (N400, N365);
or OR3 (N401, N397, N37, N21);
not NOT1 (N402, N388);
nand NAND3 (N403, N399, N205, N266);
or OR3 (N404, N392, N364, N258);
or OR2 (N405, N389, N25);
and AND3 (N406, N400, N204, N63);
and AND2 (N407, N387, N315);
xor XOR2 (N408, N393, N387);
nor NOR2 (N409, N385, N292);
nor NOR3 (N410, N404, N360, N288);
not NOT1 (N411, N394);
nor NOR2 (N412, N410, N43);
not NOT1 (N413, N405);
xor XOR2 (N414, N409, N240);
and AND4 (N415, N401, N267, N126, N410);
xor XOR2 (N416, N407, N347);
buf BUF1 (N417, N413);
and AND4 (N418, N403, N163, N46, N140);
xor XOR2 (N419, N411, N237);
xor XOR2 (N420, N415, N57);
xor XOR2 (N421, N402, N357);
xor XOR2 (N422, N406, N103);
and AND4 (N423, N418, N188, N184, N83);
and AND4 (N424, N422, N290, N167, N59);
xor XOR2 (N425, N412, N109);
buf BUF1 (N426, N416);
and AND3 (N427, N419, N96, N123);
nand NAND4 (N428, N414, N257, N237, N314);
and AND2 (N429, N421, N14);
not NOT1 (N430, N427);
xor XOR2 (N431, N424, N346);
nor NOR2 (N432, N429, N75);
or OR2 (N433, N420, N159);
not NOT1 (N434, N428);
nor NOR4 (N435, N433, N399, N240, N121);
nand NAND3 (N436, N432, N102, N67);
buf BUF1 (N437, N436);
xor XOR2 (N438, N426, N272);
not NOT1 (N439, N417);
or OR4 (N440, N408, N93, N281, N338);
and AND3 (N441, N423, N81, N426);
buf BUF1 (N442, N434);
not NOT1 (N443, N435);
not NOT1 (N444, N443);
nand NAND3 (N445, N441, N149, N162);
buf BUF1 (N446, N445);
not NOT1 (N447, N430);
buf BUF1 (N448, N438);
nor NOR3 (N449, N440, N102, N353);
nor NOR3 (N450, N442, N20, N376);
nor NOR2 (N451, N425, N105);
nor NOR2 (N452, N437, N438);
nand NAND2 (N453, N447, N71);
not NOT1 (N454, N449);
and AND3 (N455, N431, N74, N76);
not NOT1 (N456, N439);
buf BUF1 (N457, N450);
nor NOR4 (N458, N454, N33, N324, N406);
xor XOR2 (N459, N446, N31);
and AND4 (N460, N444, N20, N238, N429);
buf BUF1 (N461, N451);
or OR2 (N462, N448, N196);
xor XOR2 (N463, N452, N368);
or OR3 (N464, N457, N422, N377);
xor XOR2 (N465, N460, N115);
buf BUF1 (N466, N453);
xor XOR2 (N467, N456, N183);
nor NOR2 (N468, N462, N451);
or OR4 (N469, N459, N404, N125, N13);
nor NOR4 (N470, N461, N328, N267, N359);
nor NOR3 (N471, N466, N298, N94);
nand NAND2 (N472, N467, N113);
nand NAND3 (N473, N464, N174, N81);
and AND4 (N474, N470, N126, N285, N459);
not NOT1 (N475, N463);
nor NOR4 (N476, N469, N315, N160, N225);
nor NOR2 (N477, N465, N63);
or OR2 (N478, N477, N325);
nor NOR2 (N479, N473, N329);
nor NOR2 (N480, N474, N428);
not NOT1 (N481, N471);
buf BUF1 (N482, N476);
nand NAND3 (N483, N480, N468, N245);
nand NAND4 (N484, N406, N304, N285, N303);
not NOT1 (N485, N455);
buf BUF1 (N486, N479);
not NOT1 (N487, N484);
not NOT1 (N488, N486);
or OR3 (N489, N483, N114, N30);
and AND2 (N490, N489, N437);
not NOT1 (N491, N485);
not NOT1 (N492, N458);
and AND4 (N493, N487, N117, N103, N273);
xor XOR2 (N494, N472, N100);
and AND3 (N495, N490, N493, N287);
nor NOR4 (N496, N7, N317, N487, N205);
buf BUF1 (N497, N492);
and AND4 (N498, N494, N448, N59, N96);
nand NAND4 (N499, N495, N293, N122, N75);
nand NAND4 (N500, N478, N99, N179, N225);
buf BUF1 (N501, N475);
xor XOR2 (N502, N501, N400);
xor XOR2 (N503, N491, N362);
not NOT1 (N504, N482);
or OR4 (N505, N504, N243, N116, N436);
nor NOR2 (N506, N503, N304);
buf BUF1 (N507, N496);
or OR3 (N508, N499, N295, N64);
and AND3 (N509, N500, N21, N327);
buf BUF1 (N510, N481);
xor XOR2 (N511, N505, N393);
not NOT1 (N512, N498);
nand NAND3 (N513, N497, N340, N511);
xor XOR2 (N514, N437, N264);
nor NOR3 (N515, N502, N54, N496);
buf BUF1 (N516, N507);
xor XOR2 (N517, N512, N495);
and AND3 (N518, N508, N340, N85);
buf BUF1 (N519, N488);
not NOT1 (N520, N519);
and AND4 (N521, N509, N295, N148, N395);
not NOT1 (N522, N520);
or OR3 (N523, N514, N352, N301);
nor NOR3 (N524, N513, N277, N2);
xor XOR2 (N525, N524, N414);
nand NAND3 (N526, N516, N165, N426);
not NOT1 (N527, N517);
xor XOR2 (N528, N515, N153);
buf BUF1 (N529, N521);
nand NAND2 (N530, N522, N17);
or OR4 (N531, N518, N116, N235, N448);
not NOT1 (N532, N523);
or OR4 (N533, N531, N41, N251, N512);
nand NAND2 (N534, N526, N447);
or OR3 (N535, N532, N200, N376);
not NOT1 (N536, N506);
nor NOR2 (N537, N528, N75);
not NOT1 (N538, N535);
xor XOR2 (N539, N529, N173);
and AND2 (N540, N533, N212);
nor NOR2 (N541, N540, N408);
nor NOR4 (N542, N534, N496, N386, N348);
nand NAND3 (N543, N527, N241, N202);
xor XOR2 (N544, N538, N118);
and AND4 (N545, N542, N263, N133, N218);
buf BUF1 (N546, N544);
nor NOR4 (N547, N539, N216, N46, N274);
and AND2 (N548, N510, N458);
nand NAND2 (N549, N541, N156);
and AND2 (N550, N548, N260);
or OR2 (N551, N547, N388);
nand NAND3 (N552, N543, N216, N421);
or OR2 (N553, N550, N61);
nor NOR3 (N554, N530, N26, N169);
buf BUF1 (N555, N545);
xor XOR2 (N556, N552, N207);
or OR2 (N557, N549, N185);
and AND2 (N558, N557, N82);
nand NAND3 (N559, N546, N478, N342);
nand NAND2 (N560, N536, N145);
xor XOR2 (N561, N558, N514);
buf BUF1 (N562, N551);
not NOT1 (N563, N561);
nand NAND3 (N564, N554, N13, N81);
nand NAND3 (N565, N556, N508, N266);
nor NOR2 (N566, N565, N16);
buf BUF1 (N567, N559);
and AND4 (N568, N562, N196, N371, N29);
and AND3 (N569, N560, N470, N386);
buf BUF1 (N570, N525);
xor XOR2 (N571, N570, N122);
nor NOR3 (N572, N567, N494, N491);
not NOT1 (N573, N537);
xor XOR2 (N574, N564, N310);
buf BUF1 (N575, N571);
buf BUF1 (N576, N569);
buf BUF1 (N577, N573);
xor XOR2 (N578, N575, N133);
not NOT1 (N579, N555);
xor XOR2 (N580, N566, N16);
xor XOR2 (N581, N577, N83);
or OR3 (N582, N574, N370, N352);
nand NAND4 (N583, N582, N210, N240, N560);
and AND2 (N584, N568, N165);
xor XOR2 (N585, N581, N193);
nor NOR4 (N586, N572, N321, N347, N55);
nand NAND4 (N587, N580, N364, N90, N230);
xor XOR2 (N588, N587, N254);
nand NAND3 (N589, N576, N64, N116);
nand NAND4 (N590, N563, N283, N211, N422);
xor XOR2 (N591, N588, N494);
nor NOR4 (N592, N586, N526, N358, N549);
nand NAND3 (N593, N553, N300, N73);
or OR2 (N594, N590, N440);
nand NAND3 (N595, N593, N330, N514);
or OR3 (N596, N585, N411, N207);
buf BUF1 (N597, N594);
not NOT1 (N598, N584);
buf BUF1 (N599, N597);
xor XOR2 (N600, N595, N4);
not NOT1 (N601, N600);
buf BUF1 (N602, N583);
not NOT1 (N603, N592);
or OR2 (N604, N591, N513);
nand NAND4 (N605, N602, N234, N158, N177);
and AND3 (N606, N596, N584, N208);
and AND3 (N607, N579, N420, N97);
or OR2 (N608, N603, N532);
not NOT1 (N609, N604);
buf BUF1 (N610, N607);
xor XOR2 (N611, N601, N253);
or OR3 (N612, N598, N597, N461);
nor NOR4 (N613, N578, N319, N602, N284);
or OR2 (N614, N606, N483);
nor NOR4 (N615, N610, N97, N383, N513);
or OR4 (N616, N611, N423, N15, N469);
nor NOR3 (N617, N613, N12, N561);
buf BUF1 (N618, N599);
not NOT1 (N619, N615);
and AND3 (N620, N619, N161, N329);
buf BUF1 (N621, N617);
nor NOR2 (N622, N621, N565);
nor NOR4 (N623, N608, N80, N134, N617);
nand NAND4 (N624, N612, N401, N181, N83);
nor NOR4 (N625, N624, N344, N171, N163);
not NOT1 (N626, N625);
xor XOR2 (N627, N614, N329);
buf BUF1 (N628, N609);
not NOT1 (N629, N620);
or OR2 (N630, N589, N405);
not NOT1 (N631, N616);
nor NOR2 (N632, N623, N78);
nor NOR2 (N633, N632, N536);
or OR3 (N634, N631, N219, N48);
nor NOR2 (N635, N605, N36);
nand NAND3 (N636, N635, N565, N6);
or OR3 (N637, N629, N64, N340);
or OR3 (N638, N634, N369, N167);
or OR3 (N639, N626, N497, N91);
buf BUF1 (N640, N628);
nand NAND3 (N641, N630, N141, N429);
not NOT1 (N642, N636);
not NOT1 (N643, N633);
not NOT1 (N644, N622);
not NOT1 (N645, N637);
and AND3 (N646, N642, N431, N170);
buf BUF1 (N647, N639);
xor XOR2 (N648, N638, N468);
and AND3 (N649, N647, N356, N460);
buf BUF1 (N650, N641);
buf BUF1 (N651, N646);
or OR4 (N652, N640, N499, N445, N164);
or OR4 (N653, N643, N236, N84, N295);
and AND2 (N654, N650, N510);
buf BUF1 (N655, N653);
and AND3 (N656, N618, N326, N289);
or OR2 (N657, N655, N401);
and AND2 (N658, N657, N208);
not NOT1 (N659, N654);
xor XOR2 (N660, N644, N205);
nor NOR4 (N661, N659, N611, N88, N343);
nor NOR4 (N662, N656, N581, N451, N451);
nor NOR2 (N663, N648, N302);
and AND4 (N664, N649, N618, N654, N594);
or OR4 (N665, N660, N316, N476, N238);
not NOT1 (N666, N663);
nand NAND3 (N667, N627, N433, N443);
or OR2 (N668, N658, N155);
buf BUF1 (N669, N661);
or OR4 (N670, N668, N642, N89, N550);
or OR3 (N671, N670, N409, N393);
buf BUF1 (N672, N665);
xor XOR2 (N673, N671, N76);
and AND3 (N674, N673, N430, N223);
not NOT1 (N675, N669);
not NOT1 (N676, N674);
xor XOR2 (N677, N667, N251);
or OR3 (N678, N651, N410, N289);
nor NOR3 (N679, N664, N343, N288);
or OR3 (N680, N677, N614, N144);
and AND4 (N681, N676, N390, N95, N374);
buf BUF1 (N682, N645);
not NOT1 (N683, N682);
xor XOR2 (N684, N672, N70);
or OR2 (N685, N679, N565);
and AND4 (N686, N684, N376, N667, N541);
not NOT1 (N687, N683);
buf BUF1 (N688, N685);
or OR4 (N689, N680, N686, N93, N656);
xor XOR2 (N690, N465, N165);
and AND2 (N691, N662, N65);
and AND4 (N692, N681, N597, N297, N286);
buf BUF1 (N693, N687);
and AND3 (N694, N690, N173, N552);
buf BUF1 (N695, N675);
nand NAND3 (N696, N688, N173, N264);
and AND2 (N697, N696, N292);
nand NAND3 (N698, N666, N445, N683);
and AND4 (N699, N694, N161, N473, N49);
buf BUF1 (N700, N695);
xor XOR2 (N701, N698, N108);
buf BUF1 (N702, N701);
not NOT1 (N703, N691);
nand NAND4 (N704, N689, N347, N644, N288);
and AND4 (N705, N693, N44, N445, N594);
or OR3 (N706, N702, N126, N175);
nand NAND3 (N707, N697, N259, N607);
xor XOR2 (N708, N692, N44);
not NOT1 (N709, N706);
nor NOR3 (N710, N652, N98, N385);
nor NOR2 (N711, N700, N82);
and AND4 (N712, N710, N641, N551, N41);
or OR3 (N713, N712, N637, N223);
not NOT1 (N714, N711);
nor NOR2 (N715, N713, N236);
nand NAND3 (N716, N708, N102, N623);
xor XOR2 (N717, N705, N69);
buf BUF1 (N718, N707);
buf BUF1 (N719, N715);
not NOT1 (N720, N709);
xor XOR2 (N721, N714, N138);
nand NAND4 (N722, N716, N402, N292, N578);
and AND4 (N723, N718, N243, N306, N20);
nand NAND4 (N724, N719, N68, N205, N232);
or OR3 (N725, N703, N501, N522);
xor XOR2 (N726, N678, N134);
xor XOR2 (N727, N704, N609);
and AND3 (N728, N723, N198, N303);
not NOT1 (N729, N725);
nor NOR2 (N730, N699, N509);
nand NAND3 (N731, N730, N120, N495);
not NOT1 (N732, N731);
buf BUF1 (N733, N728);
or OR4 (N734, N724, N206, N220, N506);
buf BUF1 (N735, N734);
buf BUF1 (N736, N735);
nor NOR4 (N737, N732, N170, N229, N211);
nand NAND3 (N738, N737, N137, N241);
buf BUF1 (N739, N733);
or OR3 (N740, N739, N458, N258);
and AND4 (N741, N721, N635, N80, N337);
nand NAND3 (N742, N740, N193, N737);
and AND2 (N743, N727, N154);
nand NAND2 (N744, N742, N559);
buf BUF1 (N745, N741);
nand NAND4 (N746, N717, N170, N682, N506);
and AND4 (N747, N743, N614, N413, N301);
and AND4 (N748, N736, N401, N281, N552);
nor NOR4 (N749, N745, N566, N458, N93);
and AND2 (N750, N726, N574);
or OR4 (N751, N749, N473, N359, N457);
nand NAND4 (N752, N748, N29, N252, N210);
or OR4 (N753, N722, N89, N646, N284);
not NOT1 (N754, N738);
not NOT1 (N755, N751);
and AND3 (N756, N753, N29, N355);
and AND4 (N757, N754, N218, N273, N238);
or OR2 (N758, N752, N415);
and AND4 (N759, N744, N495, N309, N353);
buf BUF1 (N760, N756);
or OR4 (N761, N758, N659, N269, N244);
xor XOR2 (N762, N760, N702);
nor NOR2 (N763, N729, N233);
or OR4 (N764, N746, N129, N238, N528);
nor NOR3 (N765, N720, N739, N472);
not NOT1 (N766, N750);
xor XOR2 (N767, N763, N660);
buf BUF1 (N768, N764);
nand NAND3 (N769, N766, N544, N263);
not NOT1 (N770, N747);
buf BUF1 (N771, N761);
nand NAND3 (N772, N757, N274, N176);
nand NAND2 (N773, N770, N590);
xor XOR2 (N774, N765, N675);
buf BUF1 (N775, N755);
nand NAND4 (N776, N762, N620, N8, N698);
nor NOR4 (N777, N775, N59, N515, N355);
or OR3 (N778, N771, N410, N237);
not NOT1 (N779, N772);
nand NAND4 (N780, N769, N367, N341, N130);
xor XOR2 (N781, N767, N634);
nand NAND3 (N782, N779, N334, N150);
xor XOR2 (N783, N781, N296);
xor XOR2 (N784, N776, N267);
buf BUF1 (N785, N777);
nor NOR3 (N786, N782, N63, N245);
nor NOR4 (N787, N785, N679, N93, N741);
nand NAND2 (N788, N774, N359);
xor XOR2 (N789, N780, N485);
nand NAND4 (N790, N788, N630, N249, N264);
or OR3 (N791, N787, N120, N155);
and AND4 (N792, N773, N662, N724, N272);
nor NOR3 (N793, N783, N762, N709);
nand NAND4 (N794, N792, N693, N135, N401);
and AND3 (N795, N789, N222, N385);
not NOT1 (N796, N784);
or OR3 (N797, N791, N435, N6);
xor XOR2 (N798, N797, N571);
buf BUF1 (N799, N768);
and AND4 (N800, N778, N153, N95, N6);
nor NOR2 (N801, N800, N418);
nor NOR3 (N802, N759, N118, N182);
not NOT1 (N803, N801);
or OR4 (N804, N793, N767, N486, N385);
not NOT1 (N805, N802);
and AND4 (N806, N798, N394, N617, N492);
nand NAND2 (N807, N796, N794);
and AND4 (N808, N466, N20, N448, N642);
or OR3 (N809, N799, N759, N653);
nand NAND2 (N810, N805, N739);
buf BUF1 (N811, N804);
nand NAND3 (N812, N790, N538, N538);
not NOT1 (N813, N807);
or OR2 (N814, N806, N256);
not NOT1 (N815, N808);
nand NAND4 (N816, N795, N521, N677, N21);
buf BUF1 (N817, N810);
and AND3 (N818, N786, N352, N679);
and AND2 (N819, N818, N401);
buf BUF1 (N820, N809);
nand NAND4 (N821, N819, N573, N701, N392);
xor XOR2 (N822, N821, N78);
nand NAND4 (N823, N811, N483, N172, N467);
and AND3 (N824, N814, N454, N599);
and AND2 (N825, N803, N716);
buf BUF1 (N826, N820);
nor NOR4 (N827, N817, N592, N570, N362);
not NOT1 (N828, N812);
buf BUF1 (N829, N826);
nand NAND3 (N830, N824, N116, N414);
not NOT1 (N831, N829);
nor NOR4 (N832, N815, N492, N160, N268);
nor NOR4 (N833, N830, N417, N109, N184);
xor XOR2 (N834, N822, N670);
xor XOR2 (N835, N816, N559);
or OR4 (N836, N834, N500, N741, N555);
xor XOR2 (N837, N835, N80);
nor NOR2 (N838, N827, N521);
or OR3 (N839, N838, N524, N656);
not NOT1 (N840, N825);
and AND4 (N841, N833, N147, N814, N451);
and AND4 (N842, N831, N786, N451, N72);
and AND2 (N843, N813, N606);
or OR2 (N844, N839, N43);
nand NAND3 (N845, N836, N200, N146);
and AND4 (N846, N844, N721, N127, N449);
nor NOR4 (N847, N837, N313, N335, N571);
nand NAND2 (N848, N841, N613);
nand NAND4 (N849, N840, N629, N388, N22);
nand NAND4 (N850, N843, N638, N782, N587);
buf BUF1 (N851, N847);
buf BUF1 (N852, N851);
and AND2 (N853, N823, N411);
and AND3 (N854, N849, N737, N486);
not NOT1 (N855, N853);
xor XOR2 (N856, N854, N766);
nor NOR3 (N857, N856, N58, N643);
not NOT1 (N858, N832);
nor NOR2 (N859, N852, N55);
nor NOR3 (N860, N846, N239, N432);
nor NOR4 (N861, N858, N478, N37, N620);
or OR4 (N862, N859, N405, N540, N34);
not NOT1 (N863, N855);
buf BUF1 (N864, N848);
xor XOR2 (N865, N850, N592);
and AND3 (N866, N845, N134, N117);
not NOT1 (N867, N860);
or OR4 (N868, N863, N271, N705, N745);
or OR3 (N869, N865, N400, N261);
or OR4 (N870, N861, N645, N570, N8);
xor XOR2 (N871, N842, N207);
xor XOR2 (N872, N870, N113);
or OR4 (N873, N871, N173, N552, N81);
nor NOR4 (N874, N867, N429, N405, N63);
buf BUF1 (N875, N874);
or OR3 (N876, N866, N549, N838);
and AND2 (N877, N868, N646);
buf BUF1 (N878, N876);
and AND2 (N879, N875, N448);
nor NOR3 (N880, N872, N222, N790);
nor NOR2 (N881, N877, N359);
not NOT1 (N882, N862);
xor XOR2 (N883, N878, N237);
buf BUF1 (N884, N879);
buf BUF1 (N885, N882);
nor NOR4 (N886, N828, N207, N141, N624);
nand NAND2 (N887, N881, N264);
nand NAND2 (N888, N887, N542);
nor NOR3 (N889, N888, N707, N148);
xor XOR2 (N890, N873, N119);
nand NAND2 (N891, N890, N213);
and AND3 (N892, N886, N417, N787);
or OR2 (N893, N889, N345);
or OR2 (N894, N884, N105);
and AND3 (N895, N893, N331, N457);
buf BUF1 (N896, N894);
xor XOR2 (N897, N895, N525);
or OR4 (N898, N885, N803, N886, N893);
and AND4 (N899, N857, N306, N357, N57);
or OR2 (N900, N883, N68);
nor NOR3 (N901, N869, N716, N396);
nand NAND2 (N902, N892, N801);
xor XOR2 (N903, N864, N507);
and AND2 (N904, N897, N292);
and AND3 (N905, N899, N564, N148);
nand NAND3 (N906, N905, N275, N335);
and AND4 (N907, N896, N250, N742, N178);
not NOT1 (N908, N900);
xor XOR2 (N909, N898, N392);
nand NAND4 (N910, N880, N190, N137, N639);
nor NOR2 (N911, N909, N567);
nor NOR3 (N912, N906, N601, N614);
nor NOR2 (N913, N907, N46);
buf BUF1 (N914, N903);
buf BUF1 (N915, N902);
buf BUF1 (N916, N901);
or OR4 (N917, N913, N394, N894, N23);
nand NAND4 (N918, N915, N856, N406, N735);
not NOT1 (N919, N908);
xor XOR2 (N920, N918, N785);
nand NAND3 (N921, N920, N314, N735);
xor XOR2 (N922, N904, N26);
buf BUF1 (N923, N917);
and AND2 (N924, N916, N226);
not NOT1 (N925, N911);
or OR3 (N926, N923, N396, N858);
buf BUF1 (N927, N891);
nor NOR2 (N928, N924, N863);
nand NAND2 (N929, N925, N673);
xor XOR2 (N930, N922, N157);
not NOT1 (N931, N910);
nand NAND3 (N932, N928, N827, N200);
not NOT1 (N933, N914);
xor XOR2 (N934, N931, N873);
xor XOR2 (N935, N912, N162);
xor XOR2 (N936, N930, N35);
or OR4 (N937, N933, N392, N275, N348);
nand NAND2 (N938, N934, N796);
or OR2 (N939, N927, N747);
nor NOR2 (N940, N926, N740);
nor NOR4 (N941, N929, N636, N676, N524);
not NOT1 (N942, N938);
nor NOR2 (N943, N939, N420);
nand NAND3 (N944, N942, N807, N568);
buf BUF1 (N945, N943);
nand NAND4 (N946, N936, N591, N483, N35);
not NOT1 (N947, N946);
or OR3 (N948, N947, N933, N404);
or OR3 (N949, N940, N875, N815);
not NOT1 (N950, N921);
xor XOR2 (N951, N941, N882);
buf BUF1 (N952, N937);
and AND4 (N953, N945, N565, N7, N896);
and AND2 (N954, N932, N762);
nand NAND2 (N955, N919, N629);
xor XOR2 (N956, N951, N443);
buf BUF1 (N957, N952);
and AND4 (N958, N955, N275, N608, N795);
nand NAND3 (N959, N935, N36, N734);
and AND2 (N960, N944, N872);
xor XOR2 (N961, N950, N171);
buf BUF1 (N962, N957);
and AND2 (N963, N956, N633);
or OR2 (N964, N960, N274);
and AND3 (N965, N949, N738, N571);
and AND4 (N966, N965, N138, N80, N611);
or OR3 (N967, N953, N542, N142);
nor NOR4 (N968, N966, N657, N159, N870);
or OR3 (N969, N968, N85, N8);
xor XOR2 (N970, N969, N447);
not NOT1 (N971, N959);
nor NOR4 (N972, N948, N637, N213, N942);
buf BUF1 (N973, N963);
buf BUF1 (N974, N964);
nand NAND4 (N975, N967, N768, N352, N364);
nor NOR2 (N976, N970, N252);
and AND4 (N977, N954, N494, N687, N259);
not NOT1 (N978, N973);
not NOT1 (N979, N974);
buf BUF1 (N980, N972);
nor NOR2 (N981, N961, N917);
not NOT1 (N982, N979);
or OR2 (N983, N982, N625);
xor XOR2 (N984, N983, N870);
buf BUF1 (N985, N984);
nand NAND4 (N986, N978, N763, N598, N729);
and AND4 (N987, N981, N69, N305, N653);
or OR3 (N988, N976, N909, N374);
xor XOR2 (N989, N988, N532);
xor XOR2 (N990, N962, N974);
or OR4 (N991, N980, N574, N786, N84);
nand NAND3 (N992, N985, N468, N225);
buf BUF1 (N993, N971);
not NOT1 (N994, N975);
or OR4 (N995, N987, N484, N959, N372);
xor XOR2 (N996, N977, N778);
not NOT1 (N997, N991);
buf BUF1 (N998, N995);
or OR2 (N999, N993, N755);
not NOT1 (N1000, N986);
and AND3 (N1001, N999, N133, N189);
nor NOR4 (N1002, N997, N420, N877, N254);
xor XOR2 (N1003, N1001, N666);
xor XOR2 (N1004, N992, N542);
not NOT1 (N1005, N1004);
nor NOR3 (N1006, N990, N146, N26);
or OR4 (N1007, N958, N741, N871, N1002);
buf BUF1 (N1008, N287);
or OR4 (N1009, N996, N692, N794, N947);
nand NAND2 (N1010, N1005, N386);
or OR3 (N1011, N1000, N928, N185);
or OR2 (N1012, N1008, N40);
and AND3 (N1013, N1006, N959, N949);
or OR4 (N1014, N1012, N52, N465, N751);
not NOT1 (N1015, N998);
or OR2 (N1016, N989, N129);
or OR3 (N1017, N1015, N507, N358);
or OR4 (N1018, N1014, N501, N51, N994);
and AND2 (N1019, N157, N22);
not NOT1 (N1020, N1007);
and AND4 (N1021, N1013, N332, N823, N913);
or OR4 (N1022, N1018, N907, N497, N910);
not NOT1 (N1023, N1017);
nor NOR4 (N1024, N1022, N840, N134, N63);
nor NOR4 (N1025, N1024, N746, N364, N296);
or OR4 (N1026, N1011, N230, N452, N276);
nor NOR4 (N1027, N1026, N286, N659, N948);
and AND4 (N1028, N1016, N826, N59, N869);
xor XOR2 (N1029, N1027, N3);
nand NAND4 (N1030, N1003, N95, N224, N141);
nor NOR3 (N1031, N1010, N69, N791);
or OR2 (N1032, N1019, N363);
or OR3 (N1033, N1028, N4, N405);
xor XOR2 (N1034, N1023, N459);
and AND4 (N1035, N1031, N481, N979, N67);
buf BUF1 (N1036, N1021);
nor NOR2 (N1037, N1020, N575);
and AND2 (N1038, N1009, N588);
not NOT1 (N1039, N1025);
nor NOR3 (N1040, N1036, N797, N204);
nor NOR4 (N1041, N1040, N468, N485, N476);
and AND4 (N1042, N1033, N849, N796, N1011);
nand NAND2 (N1043, N1034, N176);
nand NAND4 (N1044, N1038, N24, N791, N776);
buf BUF1 (N1045, N1039);
buf BUF1 (N1046, N1041);
nor NOR2 (N1047, N1037, N386);
nor NOR2 (N1048, N1047, N453);
buf BUF1 (N1049, N1032);
or OR4 (N1050, N1030, N629, N900, N1025);
nand NAND3 (N1051, N1048, N985, N287);
and AND3 (N1052, N1050, N772, N763);
or OR2 (N1053, N1035, N795);
xor XOR2 (N1054, N1045, N620);
xor XOR2 (N1055, N1054, N564);
or OR3 (N1056, N1055, N600, N127);
nor NOR2 (N1057, N1046, N138);
xor XOR2 (N1058, N1053, N1048);
nor NOR3 (N1059, N1056, N595, N342);
buf BUF1 (N1060, N1058);
xor XOR2 (N1061, N1049, N339);
buf BUF1 (N1062, N1042);
and AND2 (N1063, N1029, N583);
nand NAND2 (N1064, N1059, N426);
buf BUF1 (N1065, N1043);
buf BUF1 (N1066, N1063);
and AND4 (N1067, N1064, N254, N957, N1034);
xor XOR2 (N1068, N1066, N449);
and AND3 (N1069, N1051, N982, N753);
buf BUF1 (N1070, N1069);
or OR2 (N1071, N1052, N260);
not NOT1 (N1072, N1065);
nor NOR2 (N1073, N1070, N597);
not NOT1 (N1074, N1044);
nor NOR4 (N1075, N1060, N727, N526, N998);
nor NOR3 (N1076, N1074, N485, N662);
and AND4 (N1077, N1076, N558, N729, N1029);
not NOT1 (N1078, N1071);
buf BUF1 (N1079, N1057);
or OR2 (N1080, N1067, N231);
and AND3 (N1081, N1068, N781, N811);
and AND4 (N1082, N1062, N527, N771, N341);
or OR4 (N1083, N1077, N843, N548, N584);
and AND3 (N1084, N1080, N1042, N59);
or OR2 (N1085, N1072, N236);
not NOT1 (N1086, N1075);
nand NAND3 (N1087, N1079, N621, N957);
not NOT1 (N1088, N1086);
nand NAND2 (N1089, N1083, N262);
nor NOR3 (N1090, N1088, N306, N852);
nand NAND4 (N1091, N1087, N417, N743, N515);
nor NOR3 (N1092, N1084, N842, N250);
not NOT1 (N1093, N1089);
nor NOR2 (N1094, N1093, N345);
nor NOR4 (N1095, N1082, N978, N365, N658);
or OR4 (N1096, N1090, N311, N311, N1065);
buf BUF1 (N1097, N1085);
xor XOR2 (N1098, N1095, N554);
nand NAND4 (N1099, N1094, N156, N1058, N902);
and AND2 (N1100, N1081, N374);
not NOT1 (N1101, N1100);
xor XOR2 (N1102, N1091, N962);
xor XOR2 (N1103, N1102, N444);
and AND4 (N1104, N1098, N480, N464, N433);
nor NOR2 (N1105, N1097, N771);
buf BUF1 (N1106, N1105);
xor XOR2 (N1107, N1101, N667);
buf BUF1 (N1108, N1103);
or OR4 (N1109, N1078, N1040, N889, N1062);
nor NOR2 (N1110, N1061, N1088);
nand NAND2 (N1111, N1096, N1017);
xor XOR2 (N1112, N1092, N1006);
nand NAND3 (N1113, N1109, N1090, N117);
nor NOR2 (N1114, N1073, N674);
buf BUF1 (N1115, N1106);
and AND3 (N1116, N1112, N127, N629);
buf BUF1 (N1117, N1099);
xor XOR2 (N1118, N1111, N781);
xor XOR2 (N1119, N1104, N583);
xor XOR2 (N1120, N1108, N163);
nor NOR3 (N1121, N1113, N442, N912);
xor XOR2 (N1122, N1120, N29);
nand NAND3 (N1123, N1114, N192, N825);
or OR4 (N1124, N1117, N382, N652, N333);
nand NAND3 (N1125, N1110, N313, N811);
buf BUF1 (N1126, N1119);
not NOT1 (N1127, N1126);
not NOT1 (N1128, N1121);
xor XOR2 (N1129, N1116, N112);
buf BUF1 (N1130, N1118);
or OR3 (N1131, N1128, N195, N485);
buf BUF1 (N1132, N1129);
not NOT1 (N1133, N1127);
nand NAND4 (N1134, N1107, N943, N808, N403);
xor XOR2 (N1135, N1123, N495);
xor XOR2 (N1136, N1125, N330);
or OR3 (N1137, N1122, N665, N644);
buf BUF1 (N1138, N1124);
nand NAND4 (N1139, N1133, N110, N634, N301);
not NOT1 (N1140, N1139);
buf BUF1 (N1141, N1132);
nor NOR3 (N1142, N1134, N323, N93);
or OR2 (N1143, N1135, N135);
nor NOR2 (N1144, N1143, N539);
or OR3 (N1145, N1140, N8, N107);
or OR2 (N1146, N1141, N242);
or OR4 (N1147, N1138, N757, N68, N50);
or OR4 (N1148, N1137, N101, N917, N621);
buf BUF1 (N1149, N1130);
nand NAND4 (N1150, N1115, N594, N31, N178);
nand NAND2 (N1151, N1142, N689);
and AND2 (N1152, N1144, N1019);
and AND4 (N1153, N1149, N576, N9, N553);
nand NAND2 (N1154, N1146, N34);
and AND2 (N1155, N1151, N1033);
buf BUF1 (N1156, N1147);
or OR2 (N1157, N1131, N125);
not NOT1 (N1158, N1155);
and AND3 (N1159, N1152, N267, N1059);
and AND4 (N1160, N1159, N587, N447, N278);
buf BUF1 (N1161, N1145);
buf BUF1 (N1162, N1156);
xor XOR2 (N1163, N1150, N390);
and AND3 (N1164, N1148, N1104, N822);
not NOT1 (N1165, N1160);
buf BUF1 (N1166, N1154);
nand NAND4 (N1167, N1158, N226, N655, N1050);
nor NOR2 (N1168, N1157, N615);
xor XOR2 (N1169, N1136, N549);
not NOT1 (N1170, N1166);
nor NOR3 (N1171, N1163, N970, N938);
nor NOR2 (N1172, N1162, N270);
nor NOR2 (N1173, N1164, N205);
buf BUF1 (N1174, N1167);
xor XOR2 (N1175, N1173, N75);
or OR2 (N1176, N1174, N290);
and AND3 (N1177, N1176, N795, N876);
or OR2 (N1178, N1161, N509);
nand NAND2 (N1179, N1171, N918);
nor NOR3 (N1180, N1165, N933, N884);
nand NAND4 (N1181, N1177, N65, N617, N169);
nor NOR4 (N1182, N1180, N1132, N1148, N732);
nand NAND4 (N1183, N1153, N773, N300, N481);
xor XOR2 (N1184, N1170, N857);
not NOT1 (N1185, N1175);
xor XOR2 (N1186, N1184, N390);
xor XOR2 (N1187, N1182, N1027);
buf BUF1 (N1188, N1178);
nor NOR3 (N1189, N1185, N735, N717);
nor NOR2 (N1190, N1187, N1040);
and AND2 (N1191, N1188, N563);
nand NAND4 (N1192, N1172, N764, N955, N639);
or OR2 (N1193, N1192, N956);
xor XOR2 (N1194, N1190, N399);
nand NAND4 (N1195, N1169, N153, N368, N1086);
nor NOR4 (N1196, N1183, N744, N504, N519);
nand NAND4 (N1197, N1186, N801, N688, N119);
nand NAND2 (N1198, N1193, N292);
or OR3 (N1199, N1191, N224, N1100);
nand NAND3 (N1200, N1195, N306, N106);
or OR2 (N1201, N1181, N1162);
xor XOR2 (N1202, N1197, N853);
not NOT1 (N1203, N1196);
nor NOR4 (N1204, N1168, N1158, N566, N605);
xor XOR2 (N1205, N1202, N435);
not NOT1 (N1206, N1198);
nor NOR2 (N1207, N1205, N266);
not NOT1 (N1208, N1179);
buf BUF1 (N1209, N1208);
not NOT1 (N1210, N1201);
nor NOR2 (N1211, N1194, N669);
nor NOR2 (N1212, N1206, N1148);
buf BUF1 (N1213, N1203);
buf BUF1 (N1214, N1204);
not NOT1 (N1215, N1209);
buf BUF1 (N1216, N1199);
buf BUF1 (N1217, N1211);
and AND3 (N1218, N1212, N472, N249);
nand NAND4 (N1219, N1189, N932, N422, N416);
nand NAND2 (N1220, N1219, N472);
xor XOR2 (N1221, N1214, N265);
or OR3 (N1222, N1217, N421, N903);
nor NOR2 (N1223, N1210, N1005);
and AND3 (N1224, N1221, N58, N933);
or OR2 (N1225, N1200, N988);
not NOT1 (N1226, N1224);
nand NAND2 (N1227, N1225, N1170);
and AND2 (N1228, N1220, N527);
nor NOR4 (N1229, N1227, N306, N326, N96);
or OR2 (N1230, N1216, N343);
xor XOR2 (N1231, N1226, N165);
buf BUF1 (N1232, N1218);
xor XOR2 (N1233, N1215, N229);
not NOT1 (N1234, N1213);
buf BUF1 (N1235, N1234);
xor XOR2 (N1236, N1222, N891);
not NOT1 (N1237, N1231);
or OR4 (N1238, N1223, N129, N426, N387);
xor XOR2 (N1239, N1207, N940);
nand NAND4 (N1240, N1239, N1239, N732, N1050);
buf BUF1 (N1241, N1235);
or OR3 (N1242, N1230, N754, N207);
xor XOR2 (N1243, N1236, N727);
buf BUF1 (N1244, N1240);
and AND4 (N1245, N1232, N178, N159, N45);
nor NOR3 (N1246, N1245, N568, N811);
or OR2 (N1247, N1241, N87);
or OR4 (N1248, N1238, N177, N819, N1214);
and AND3 (N1249, N1246, N11, N1049);
nand NAND4 (N1250, N1244, N851, N751, N448);
buf BUF1 (N1251, N1249);
not NOT1 (N1252, N1233);
and AND4 (N1253, N1248, N61, N311, N502);
xor XOR2 (N1254, N1243, N578);
nand NAND3 (N1255, N1228, N1218, N531);
and AND2 (N1256, N1250, N1023);
nor NOR2 (N1257, N1229, N1045);
buf BUF1 (N1258, N1257);
and AND3 (N1259, N1254, N883, N44);
nand NAND3 (N1260, N1259, N265, N872);
nand NAND4 (N1261, N1251, N380, N352, N493);
xor XOR2 (N1262, N1255, N1215);
buf BUF1 (N1263, N1260);
and AND3 (N1264, N1252, N965, N737);
and AND2 (N1265, N1263, N417);
nand NAND2 (N1266, N1247, N1118);
buf BUF1 (N1267, N1258);
buf BUF1 (N1268, N1253);
nor NOR2 (N1269, N1264, N293);
xor XOR2 (N1270, N1268, N1217);
and AND4 (N1271, N1261, N1003, N327, N767);
nor NOR2 (N1272, N1269, N378);
not NOT1 (N1273, N1242);
buf BUF1 (N1274, N1262);
and AND4 (N1275, N1237, N769, N1212, N623);
xor XOR2 (N1276, N1270, N422);
not NOT1 (N1277, N1274);
xor XOR2 (N1278, N1271, N790);
xor XOR2 (N1279, N1267, N369);
and AND3 (N1280, N1277, N153, N121);
not NOT1 (N1281, N1275);
buf BUF1 (N1282, N1265);
and AND2 (N1283, N1278, N372);
buf BUF1 (N1284, N1273);
xor XOR2 (N1285, N1281, N1236);
not NOT1 (N1286, N1280);
buf BUF1 (N1287, N1286);
nor NOR2 (N1288, N1283, N275);
and AND3 (N1289, N1288, N531, N743);
nor NOR3 (N1290, N1279, N204, N338);
xor XOR2 (N1291, N1289, N1184);
and AND4 (N1292, N1284, N1214, N519, N587);
not NOT1 (N1293, N1290);
nor NOR3 (N1294, N1272, N228, N902);
or OR3 (N1295, N1291, N1140, N216);
or OR3 (N1296, N1294, N1227, N994);
nor NOR2 (N1297, N1256, N1135);
nand NAND3 (N1298, N1295, N414, N556);
nand NAND2 (N1299, N1266, N840);
not NOT1 (N1300, N1299);
buf BUF1 (N1301, N1282);
and AND4 (N1302, N1297, N620, N42, N766);
nor NOR4 (N1303, N1285, N725, N839, N704);
not NOT1 (N1304, N1298);
not NOT1 (N1305, N1276);
buf BUF1 (N1306, N1302);
xor XOR2 (N1307, N1305, N257);
or OR3 (N1308, N1307, N1210, N386);
or OR3 (N1309, N1287, N712, N1079);
nand NAND4 (N1310, N1304, N1294, N687, N1176);
buf BUF1 (N1311, N1306);
nand NAND3 (N1312, N1310, N146, N421);
or OR3 (N1313, N1308, N616, N661);
or OR3 (N1314, N1313, N153, N690);
or OR2 (N1315, N1314, N1197);
and AND4 (N1316, N1300, N1087, N291, N1104);
not NOT1 (N1317, N1315);
not NOT1 (N1318, N1292);
not NOT1 (N1319, N1303);
or OR4 (N1320, N1318, N554, N1183, N1106);
and AND2 (N1321, N1296, N1280);
xor XOR2 (N1322, N1311, N591);
and AND3 (N1323, N1312, N289, N835);
and AND3 (N1324, N1322, N1196, N1268);
not NOT1 (N1325, N1323);
not NOT1 (N1326, N1316);
xor XOR2 (N1327, N1320, N1017);
and AND2 (N1328, N1319, N153);
nor NOR4 (N1329, N1301, N640, N848, N308);
not NOT1 (N1330, N1328);
buf BUF1 (N1331, N1326);
or OR3 (N1332, N1324, N530, N1307);
nand NAND3 (N1333, N1325, N863, N80);
buf BUF1 (N1334, N1327);
or OR3 (N1335, N1333, N843, N989);
xor XOR2 (N1336, N1317, N269);
buf BUF1 (N1337, N1335);
buf BUF1 (N1338, N1337);
buf BUF1 (N1339, N1329);
not NOT1 (N1340, N1339);
and AND4 (N1341, N1309, N505, N1264, N142);
not NOT1 (N1342, N1331);
xor XOR2 (N1343, N1330, N272);
or OR2 (N1344, N1321, N1270);
nor NOR4 (N1345, N1344, N186, N859, N994);
not NOT1 (N1346, N1342);
xor XOR2 (N1347, N1341, N207);
nor NOR4 (N1348, N1336, N996, N663, N615);
nand NAND3 (N1349, N1347, N13, N498);
nor NOR3 (N1350, N1338, N1326, N238);
xor XOR2 (N1351, N1343, N142);
buf BUF1 (N1352, N1334);
nor NOR4 (N1353, N1349, N1161, N801, N1272);
not NOT1 (N1354, N1332);
not NOT1 (N1355, N1346);
buf BUF1 (N1356, N1354);
and AND4 (N1357, N1345, N181, N1262, N119);
not NOT1 (N1358, N1356);
or OR2 (N1359, N1352, N266);
buf BUF1 (N1360, N1357);
or OR3 (N1361, N1358, N1312, N961);
and AND4 (N1362, N1361, N1165, N257, N1036);
nor NOR2 (N1363, N1340, N656);
or OR3 (N1364, N1359, N652, N51);
and AND3 (N1365, N1364, N1068, N206);
nor NOR2 (N1366, N1362, N725);
xor XOR2 (N1367, N1355, N1352);
nor NOR3 (N1368, N1366, N911, N1108);
nor NOR3 (N1369, N1353, N15, N1338);
xor XOR2 (N1370, N1363, N971);
and AND2 (N1371, N1365, N5);
not NOT1 (N1372, N1371);
and AND2 (N1373, N1367, N1347);
or OR4 (N1374, N1293, N405, N350, N1288);
or OR2 (N1375, N1351, N1047);
xor XOR2 (N1376, N1374, N158);
nand NAND2 (N1377, N1348, N326);
nor NOR2 (N1378, N1376, N246);
nor NOR4 (N1379, N1370, N319, N874, N939);
buf BUF1 (N1380, N1375);
nand NAND4 (N1381, N1379, N262, N1080, N456);
or OR3 (N1382, N1372, N309, N240);
or OR3 (N1383, N1350, N160, N42);
nor NOR3 (N1384, N1383, N677, N541);
or OR2 (N1385, N1378, N207);
or OR4 (N1386, N1369, N1157, N618, N590);
buf BUF1 (N1387, N1381);
and AND2 (N1388, N1368, N375);
buf BUF1 (N1389, N1382);
not NOT1 (N1390, N1377);
xor XOR2 (N1391, N1373, N467);
not NOT1 (N1392, N1360);
nor NOR3 (N1393, N1384, N966, N480);
nand NAND4 (N1394, N1393, N1216, N1297, N25);
nor NOR3 (N1395, N1385, N799, N216);
buf BUF1 (N1396, N1395);
nand NAND4 (N1397, N1387, N1335, N399, N452);
nor NOR3 (N1398, N1392, N1207, N762);
not NOT1 (N1399, N1396);
or OR4 (N1400, N1389, N1068, N151, N1216);
and AND2 (N1401, N1390, N52);
xor XOR2 (N1402, N1386, N485);
and AND4 (N1403, N1402, N296, N679, N829);
not NOT1 (N1404, N1397);
nor NOR4 (N1405, N1398, N955, N754, N534);
and AND4 (N1406, N1391, N1300, N474, N894);
nand NAND4 (N1407, N1399, N1160, N836, N1154);
nor NOR2 (N1408, N1403, N372);
buf BUF1 (N1409, N1407);
and AND3 (N1410, N1408, N1281, N182);
buf BUF1 (N1411, N1406);
not NOT1 (N1412, N1405);
xor XOR2 (N1413, N1380, N318);
not NOT1 (N1414, N1394);
nand NAND2 (N1415, N1412, N564);
buf BUF1 (N1416, N1415);
nor NOR4 (N1417, N1401, N1278, N675, N533);
buf BUF1 (N1418, N1404);
and AND4 (N1419, N1400, N659, N1316, N845);
xor XOR2 (N1420, N1411, N905);
or OR4 (N1421, N1416, N165, N218, N842);
nand NAND3 (N1422, N1414, N1314, N297);
nor NOR2 (N1423, N1388, N350);
not NOT1 (N1424, N1419);
or OR4 (N1425, N1418, N653, N715, N1120);
and AND3 (N1426, N1420, N122, N1345);
nand NAND4 (N1427, N1426, N456, N633, N725);
buf BUF1 (N1428, N1417);
or OR2 (N1429, N1409, N341);
nand NAND2 (N1430, N1421, N24);
not NOT1 (N1431, N1410);
nor NOR4 (N1432, N1430, N1132, N246, N12);
nand NAND3 (N1433, N1422, N361, N1421);
or OR4 (N1434, N1423, N508, N386, N978);
nand NAND3 (N1435, N1431, N856, N1117);
nor NOR3 (N1436, N1435, N718, N840);
nor NOR3 (N1437, N1429, N815, N1274);
not NOT1 (N1438, N1413);
buf BUF1 (N1439, N1432);
nand NAND2 (N1440, N1425, N1132);
and AND3 (N1441, N1424, N365, N528);
nor NOR2 (N1442, N1427, N1048);
or OR4 (N1443, N1434, N1216, N941, N575);
or OR3 (N1444, N1438, N48, N121);
or OR2 (N1445, N1436, N837);
nand NAND4 (N1446, N1433, N21, N1161, N1353);
xor XOR2 (N1447, N1440, N265);
or OR3 (N1448, N1441, N744, N1214);
nand NAND2 (N1449, N1439, N335);
not NOT1 (N1450, N1445);
nor NOR4 (N1451, N1446, N112, N209, N87);
and AND4 (N1452, N1442, N1393, N58, N1065);
or OR4 (N1453, N1449, N134, N1187, N1356);
and AND3 (N1454, N1428, N127, N1227);
xor XOR2 (N1455, N1451, N547);
buf BUF1 (N1456, N1455);
or OR4 (N1457, N1448, N1323, N44, N1241);
nand NAND2 (N1458, N1452, N1117);
not NOT1 (N1459, N1454);
not NOT1 (N1460, N1437);
or OR2 (N1461, N1453, N64);
nand NAND3 (N1462, N1459, N1312, N863);
buf BUF1 (N1463, N1458);
nor NOR3 (N1464, N1456, N1166, N417);
not NOT1 (N1465, N1461);
xor XOR2 (N1466, N1460, N450);
not NOT1 (N1467, N1464);
and AND2 (N1468, N1443, N197);
nand NAND4 (N1469, N1466, N215, N277, N782);
and AND3 (N1470, N1462, N1398, N1351);
nor NOR4 (N1471, N1467, N1235, N1340, N643);
and AND2 (N1472, N1465, N1245);
nor NOR2 (N1473, N1463, N936);
or OR4 (N1474, N1457, N223, N347, N478);
nor NOR2 (N1475, N1472, N573);
or OR2 (N1476, N1468, N717);
not NOT1 (N1477, N1444);
and AND3 (N1478, N1470, N408, N937);
nand NAND4 (N1479, N1476, N1404, N1256, N1268);
or OR2 (N1480, N1475, N883);
not NOT1 (N1481, N1477);
nand NAND3 (N1482, N1469, N1019, N1326);
nor NOR3 (N1483, N1479, N285, N1434);
nand NAND4 (N1484, N1450, N47, N1054, N1074);
or OR2 (N1485, N1478, N1395);
nor NOR4 (N1486, N1473, N792, N472, N675);
buf BUF1 (N1487, N1486);
not NOT1 (N1488, N1474);
nand NAND4 (N1489, N1485, N1190, N876, N992);
nor NOR3 (N1490, N1487, N1016, N757);
or OR3 (N1491, N1483, N137, N334);
xor XOR2 (N1492, N1471, N270);
not NOT1 (N1493, N1490);
buf BUF1 (N1494, N1447);
nand NAND2 (N1495, N1493, N39);
not NOT1 (N1496, N1491);
nor NOR2 (N1497, N1492, N482);
or OR3 (N1498, N1488, N93, N444);
and AND2 (N1499, N1494, N462);
not NOT1 (N1500, N1480);
nor NOR4 (N1501, N1498, N513, N760, N761);
xor XOR2 (N1502, N1482, N232);
buf BUF1 (N1503, N1495);
nand NAND4 (N1504, N1496, N948, N603, N1484);
xor XOR2 (N1505, N1235, N161);
and AND4 (N1506, N1505, N755, N386, N1448);
buf BUF1 (N1507, N1501);
and AND4 (N1508, N1504, N1060, N341, N1187);
not NOT1 (N1509, N1481);
nand NAND3 (N1510, N1506, N1262, N495);
xor XOR2 (N1511, N1508, N203);
nor NOR4 (N1512, N1500, N332, N118, N646);
and AND2 (N1513, N1510, N782);
nor NOR2 (N1514, N1511, N714);
and AND3 (N1515, N1514, N1400, N156);
buf BUF1 (N1516, N1499);
buf BUF1 (N1517, N1516);
not NOT1 (N1518, N1502);
and AND4 (N1519, N1513, N760, N1191, N726);
nor NOR2 (N1520, N1497, N225);
not NOT1 (N1521, N1489);
or OR4 (N1522, N1521, N1320, N454, N559);
or OR2 (N1523, N1515, N465);
xor XOR2 (N1524, N1519, N1520);
not NOT1 (N1525, N608);
buf BUF1 (N1526, N1517);
xor XOR2 (N1527, N1522, N210);
nor NOR4 (N1528, N1507, N1487, N1034, N1316);
not NOT1 (N1529, N1523);
nand NAND4 (N1530, N1518, N1439, N1048, N1280);
and AND2 (N1531, N1512, N864);
not NOT1 (N1532, N1525);
buf BUF1 (N1533, N1529);
nand NAND2 (N1534, N1528, N320);
and AND4 (N1535, N1530, N978, N560, N596);
not NOT1 (N1536, N1532);
and AND2 (N1537, N1531, N180);
nand NAND2 (N1538, N1527, N895);
nor NOR4 (N1539, N1534, N24, N1201, N236);
nand NAND3 (N1540, N1533, N690, N459);
buf BUF1 (N1541, N1536);
and AND3 (N1542, N1540, N41, N495);
not NOT1 (N1543, N1526);
nor NOR3 (N1544, N1503, N1151, N1528);
buf BUF1 (N1545, N1539);
xor XOR2 (N1546, N1538, N898);
or OR2 (N1547, N1542, N61);
nand NAND4 (N1548, N1545, N312, N1278, N1044);
not NOT1 (N1549, N1541);
nand NAND4 (N1550, N1535, N567, N895, N1205);
not NOT1 (N1551, N1509);
or OR3 (N1552, N1551, N1534, N521);
not NOT1 (N1553, N1544);
not NOT1 (N1554, N1546);
nand NAND4 (N1555, N1554, N1096, N1199, N816);
buf BUF1 (N1556, N1553);
and AND3 (N1557, N1556, N644, N326);
nor NOR4 (N1558, N1550, N1403, N1513, N1249);
buf BUF1 (N1559, N1557);
nand NAND2 (N1560, N1549, N730);
and AND2 (N1561, N1558, N748);
buf BUF1 (N1562, N1561);
and AND3 (N1563, N1548, N712, N1173);
xor XOR2 (N1564, N1563, N218);
xor XOR2 (N1565, N1524, N39);
or OR4 (N1566, N1543, N1223, N1053, N1285);
not NOT1 (N1567, N1560);
buf BUF1 (N1568, N1562);
nor NOR2 (N1569, N1552, N780);
nor NOR3 (N1570, N1567, N321, N1139);
or OR4 (N1571, N1564, N582, N1130, N593);
not NOT1 (N1572, N1571);
xor XOR2 (N1573, N1565, N133);
nor NOR3 (N1574, N1570, N751, N469);
nor NOR3 (N1575, N1566, N527, N1350);
and AND3 (N1576, N1559, N1301, N469);
buf BUF1 (N1577, N1575);
or OR2 (N1578, N1555, N803);
and AND4 (N1579, N1569, N1143, N1569, N242);
not NOT1 (N1580, N1572);
nor NOR4 (N1581, N1568, N261, N385, N237);
buf BUF1 (N1582, N1580);
nand NAND2 (N1583, N1537, N306);
nor NOR2 (N1584, N1579, N761);
or OR3 (N1585, N1581, N458, N126);
and AND3 (N1586, N1578, N1380, N64);
xor XOR2 (N1587, N1547, N433);
xor XOR2 (N1588, N1582, N1245);
nor NOR2 (N1589, N1573, N1320);
and AND4 (N1590, N1583, N364, N77, N733);
nand NAND3 (N1591, N1588, N1370, N1357);
nor NOR4 (N1592, N1590, N291, N790, N863);
and AND3 (N1593, N1577, N865, N12);
or OR3 (N1594, N1574, N904, N757);
and AND4 (N1595, N1594, N1498, N1474, N271);
nor NOR2 (N1596, N1595, N472);
nand NAND3 (N1597, N1586, N266, N358);
buf BUF1 (N1598, N1587);
not NOT1 (N1599, N1592);
nor NOR3 (N1600, N1597, N1376, N432);
buf BUF1 (N1601, N1600);
buf BUF1 (N1602, N1589);
or OR3 (N1603, N1593, N1037, N1419);
nor NOR2 (N1604, N1596, N475);
not NOT1 (N1605, N1585);
or OR4 (N1606, N1602, N368, N45, N823);
and AND3 (N1607, N1598, N292, N784);
and AND3 (N1608, N1576, N1331, N119);
and AND2 (N1609, N1584, N592);
and AND2 (N1610, N1609, N824);
nor NOR3 (N1611, N1603, N711, N1539);
nor NOR4 (N1612, N1604, N1130, N963, N479);
xor XOR2 (N1613, N1605, N854);
xor XOR2 (N1614, N1606, N1269);
not NOT1 (N1615, N1591);
nor NOR3 (N1616, N1611, N1167, N449);
xor XOR2 (N1617, N1610, N1033);
buf BUF1 (N1618, N1608);
nor NOR3 (N1619, N1616, N573, N1132);
nand NAND4 (N1620, N1599, N643, N291, N876);
not NOT1 (N1621, N1614);
buf BUF1 (N1622, N1619);
or OR2 (N1623, N1617, N144);
not NOT1 (N1624, N1621);
not NOT1 (N1625, N1615);
buf BUF1 (N1626, N1620);
buf BUF1 (N1627, N1607);
or OR4 (N1628, N1601, N1369, N305, N134);
and AND2 (N1629, N1622, N32);
buf BUF1 (N1630, N1627);
nor NOR2 (N1631, N1629, N855);
nor NOR2 (N1632, N1623, N1617);
nor NOR4 (N1633, N1626, N1291, N498, N1387);
nor NOR2 (N1634, N1624, N1067);
not NOT1 (N1635, N1634);
and AND4 (N1636, N1632, N1225, N1018, N1181);
not NOT1 (N1637, N1625);
and AND3 (N1638, N1635, N1236, N774);
xor XOR2 (N1639, N1633, N1002);
and AND3 (N1640, N1630, N1227, N1128);
or OR2 (N1641, N1618, N593);
not NOT1 (N1642, N1638);
or OR4 (N1643, N1612, N874, N1230, N741);
buf BUF1 (N1644, N1641);
xor XOR2 (N1645, N1631, N1098);
or OR3 (N1646, N1639, N506, N1469);
or OR4 (N1647, N1646, N126, N219, N1462);
or OR3 (N1648, N1640, N176, N612);
nor NOR4 (N1649, N1644, N6, N1285, N134);
xor XOR2 (N1650, N1648, N456);
not NOT1 (N1651, N1649);
nand NAND4 (N1652, N1613, N1005, N605, N125);
and AND3 (N1653, N1637, N173, N801);
or OR4 (N1654, N1647, N404, N122, N133);
buf BUF1 (N1655, N1645);
xor XOR2 (N1656, N1653, N691);
nor NOR4 (N1657, N1656, N730, N82, N865);
not NOT1 (N1658, N1657);
xor XOR2 (N1659, N1643, N1455);
nand NAND4 (N1660, N1650, N1442, N835, N1300);
nand NAND4 (N1661, N1660, N137, N1356, N1640);
or OR3 (N1662, N1642, N1423, N183);
nor NOR4 (N1663, N1661, N279, N299, N1322);
or OR2 (N1664, N1628, N606);
buf BUF1 (N1665, N1654);
buf BUF1 (N1666, N1659);
nand NAND2 (N1667, N1664, N46);
buf BUF1 (N1668, N1667);
or OR4 (N1669, N1663, N589, N1081, N1152);
xor XOR2 (N1670, N1655, N470);
and AND4 (N1671, N1669, N1075, N1088, N26);
buf BUF1 (N1672, N1666);
and AND3 (N1673, N1658, N1054, N846);
xor XOR2 (N1674, N1665, N1062);
nand NAND2 (N1675, N1671, N357);
and AND2 (N1676, N1675, N105);
xor XOR2 (N1677, N1670, N970);
or OR3 (N1678, N1636, N1631, N411);
not NOT1 (N1679, N1652);
not NOT1 (N1680, N1673);
nor NOR4 (N1681, N1668, N977, N350, N275);
and AND3 (N1682, N1651, N677, N913);
buf BUF1 (N1683, N1679);
buf BUF1 (N1684, N1676);
and AND3 (N1685, N1672, N630, N1558);
not NOT1 (N1686, N1680);
buf BUF1 (N1687, N1678);
not NOT1 (N1688, N1662);
or OR2 (N1689, N1682, N939);
nand NAND4 (N1690, N1685, N398, N237, N1584);
or OR3 (N1691, N1686, N214, N304);
not NOT1 (N1692, N1687);
buf BUF1 (N1693, N1681);
xor XOR2 (N1694, N1690, N405);
nand NAND4 (N1695, N1688, N1589, N799, N9);
and AND3 (N1696, N1695, N1410, N1330);
nand NAND2 (N1697, N1674, N384);
not NOT1 (N1698, N1683);
not NOT1 (N1699, N1694);
buf BUF1 (N1700, N1693);
xor XOR2 (N1701, N1697, N1111);
buf BUF1 (N1702, N1696);
nor NOR4 (N1703, N1684, N1673, N227, N710);
not NOT1 (N1704, N1701);
buf BUF1 (N1705, N1689);
or OR2 (N1706, N1699, N93);
buf BUF1 (N1707, N1703);
and AND2 (N1708, N1704, N994);
not NOT1 (N1709, N1700);
not NOT1 (N1710, N1692);
xor XOR2 (N1711, N1677, N105);
nor NOR3 (N1712, N1691, N1017, N1696);
nor NOR3 (N1713, N1706, N1460, N1061);
and AND4 (N1714, N1709, N907, N160, N1666);
buf BUF1 (N1715, N1711);
nor NOR2 (N1716, N1698, N463);
and AND2 (N1717, N1714, N1529);
nand NAND2 (N1718, N1716, N983);
buf BUF1 (N1719, N1712);
or OR3 (N1720, N1710, N1047, N292);
xor XOR2 (N1721, N1713, N1273);
nand NAND3 (N1722, N1715, N192, N623);
or OR4 (N1723, N1721, N634, N285, N1121);
not NOT1 (N1724, N1708);
or OR4 (N1725, N1720, N1366, N641, N533);
nand NAND3 (N1726, N1724, N545, N930);
nand NAND3 (N1727, N1705, N38, N631);
xor XOR2 (N1728, N1726, N551);
and AND4 (N1729, N1718, N1627, N1196, N1352);
and AND2 (N1730, N1707, N832);
not NOT1 (N1731, N1725);
not NOT1 (N1732, N1702);
nand NAND4 (N1733, N1722, N664, N1693, N180);
xor XOR2 (N1734, N1719, N642);
and AND4 (N1735, N1717, N475, N380, N1365);
xor XOR2 (N1736, N1733, N894);
not NOT1 (N1737, N1723);
nor NOR3 (N1738, N1737, N287, N1305);
buf BUF1 (N1739, N1730);
nand NAND4 (N1740, N1731, N649, N1236, N596);
xor XOR2 (N1741, N1728, N335);
not NOT1 (N1742, N1732);
xor XOR2 (N1743, N1727, N1263);
and AND2 (N1744, N1739, N411);
and AND3 (N1745, N1743, N798, N1215);
buf BUF1 (N1746, N1734);
nor NOR3 (N1747, N1744, N851, N1476);
xor XOR2 (N1748, N1747, N1014);
and AND2 (N1749, N1729, N876);
and AND4 (N1750, N1736, N1336, N123, N1308);
xor XOR2 (N1751, N1742, N1002);
xor XOR2 (N1752, N1741, N312);
xor XOR2 (N1753, N1746, N129);
buf BUF1 (N1754, N1740);
and AND4 (N1755, N1749, N1663, N1031, N1729);
and AND3 (N1756, N1748, N1598, N1404);
nor NOR2 (N1757, N1753, N1555);
not NOT1 (N1758, N1750);
xor XOR2 (N1759, N1751, N1085);
not NOT1 (N1760, N1758);
xor XOR2 (N1761, N1759, N713);
and AND3 (N1762, N1752, N1343, N565);
or OR4 (N1763, N1761, N1595, N314, N90);
nand NAND3 (N1764, N1754, N1643, N502);
not NOT1 (N1765, N1763);
nor NOR3 (N1766, N1738, N901, N878);
buf BUF1 (N1767, N1735);
not NOT1 (N1768, N1764);
buf BUF1 (N1769, N1762);
and AND4 (N1770, N1755, N261, N1608, N863);
nand NAND4 (N1771, N1770, N590, N1477, N81);
xor XOR2 (N1772, N1768, N1454);
and AND4 (N1773, N1765, N1102, N1252, N588);
xor XOR2 (N1774, N1756, N537);
xor XOR2 (N1775, N1769, N294);
not NOT1 (N1776, N1772);
or OR4 (N1777, N1776, N691, N1035, N941);
xor XOR2 (N1778, N1775, N526);
or OR2 (N1779, N1745, N234);
or OR4 (N1780, N1766, N882, N1220, N1115);
and AND2 (N1781, N1767, N1065);
nand NAND3 (N1782, N1757, N1471, N352);
xor XOR2 (N1783, N1782, N1070);
nand NAND4 (N1784, N1774, N1641, N728, N740);
buf BUF1 (N1785, N1778);
nand NAND2 (N1786, N1785, N635);
nor NOR4 (N1787, N1777, N1209, N713, N1628);
xor XOR2 (N1788, N1773, N1340);
buf BUF1 (N1789, N1784);
not NOT1 (N1790, N1787);
nor NOR3 (N1791, N1789, N1170, N98);
buf BUF1 (N1792, N1780);
nor NOR3 (N1793, N1788, N1691, N454);
or OR2 (N1794, N1779, N1417);
nand NAND3 (N1795, N1786, N4, N1077);
not NOT1 (N1796, N1793);
buf BUF1 (N1797, N1794);
or OR4 (N1798, N1797, N31, N1754, N1457);
nand NAND4 (N1799, N1760, N1502, N1662, N1768);
xor XOR2 (N1800, N1783, N982);
not NOT1 (N1801, N1795);
nand NAND3 (N1802, N1771, N922, N734);
nor NOR3 (N1803, N1792, N532, N1417);
xor XOR2 (N1804, N1802, N358);
not NOT1 (N1805, N1791);
not NOT1 (N1806, N1800);
buf BUF1 (N1807, N1798);
buf BUF1 (N1808, N1790);
nand NAND3 (N1809, N1803, N614, N1233);
or OR4 (N1810, N1801, N113, N1045, N832);
or OR2 (N1811, N1810, N674);
not NOT1 (N1812, N1796);
and AND4 (N1813, N1806, N965, N1464, N1520);
and AND3 (N1814, N1799, N1505, N1351);
or OR4 (N1815, N1805, N482, N829, N1282);
or OR3 (N1816, N1808, N1364, N1403);
not NOT1 (N1817, N1816);
nor NOR3 (N1818, N1814, N598, N1487);
and AND2 (N1819, N1815, N998);
and AND4 (N1820, N1818, N1392, N958, N852);
or OR4 (N1821, N1781, N1391, N1301, N199);
or OR2 (N1822, N1817, N176);
buf BUF1 (N1823, N1819);
not NOT1 (N1824, N1812);
or OR3 (N1825, N1823, N12, N427);
xor XOR2 (N1826, N1820, N1254);
buf BUF1 (N1827, N1811);
xor XOR2 (N1828, N1807, N1751);
buf BUF1 (N1829, N1804);
and AND4 (N1830, N1824, N100, N623, N65);
or OR3 (N1831, N1809, N713, N749);
buf BUF1 (N1832, N1828);
or OR3 (N1833, N1827, N774, N971);
buf BUF1 (N1834, N1831);
or OR2 (N1835, N1832, N1803);
or OR2 (N1836, N1825, N1162);
and AND3 (N1837, N1834, N969, N1219);
xor XOR2 (N1838, N1829, N927);
or OR4 (N1839, N1813, N24, N164, N1168);
buf BUF1 (N1840, N1830);
buf BUF1 (N1841, N1833);
nand NAND4 (N1842, N1826, N53, N597, N686);
xor XOR2 (N1843, N1839, N155);
xor XOR2 (N1844, N1822, N88);
buf BUF1 (N1845, N1844);
buf BUF1 (N1846, N1821);
nand NAND3 (N1847, N1837, N824, N31);
nor NOR4 (N1848, N1843, N1489, N219, N625);
xor XOR2 (N1849, N1845, N695);
not NOT1 (N1850, N1849);
or OR2 (N1851, N1850, N342);
xor XOR2 (N1852, N1848, N1491);
not NOT1 (N1853, N1838);
not NOT1 (N1854, N1853);
and AND3 (N1855, N1842, N625, N1015);
not NOT1 (N1856, N1851);
not NOT1 (N1857, N1852);
nand NAND3 (N1858, N1855, N930, N1455);
and AND4 (N1859, N1856, N999, N1009, N398);
or OR3 (N1860, N1846, N823, N1158);
and AND2 (N1861, N1847, N964);
nand NAND2 (N1862, N1840, N225);
nor NOR2 (N1863, N1859, N1848);
xor XOR2 (N1864, N1854, N1448);
or OR2 (N1865, N1860, N118);
buf BUF1 (N1866, N1863);
and AND2 (N1867, N1864, N1532);
nor NOR2 (N1868, N1866, N543);
and AND3 (N1869, N1862, N984, N668);
xor XOR2 (N1870, N1868, N1058);
nor NOR4 (N1871, N1841, N1649, N1505, N293);
nor NOR3 (N1872, N1869, N699, N832);
and AND3 (N1873, N1836, N120, N1219);
and AND3 (N1874, N1858, N1626, N1560);
buf BUF1 (N1875, N1873);
or OR2 (N1876, N1874, N907);
buf BUF1 (N1877, N1867);
not NOT1 (N1878, N1835);
nor NOR3 (N1879, N1876, N710, N1267);
not NOT1 (N1880, N1879);
or OR4 (N1881, N1871, N1558, N167, N720);
xor XOR2 (N1882, N1880, N744);
buf BUF1 (N1883, N1870);
xor XOR2 (N1884, N1881, N999);
buf BUF1 (N1885, N1872);
not NOT1 (N1886, N1882);
and AND3 (N1887, N1877, N347, N173);
or OR3 (N1888, N1878, N1159, N1813);
nand NAND2 (N1889, N1887, N1590);
and AND2 (N1890, N1888, N596);
or OR4 (N1891, N1889, N1367, N1030, N557);
not NOT1 (N1892, N1884);
and AND4 (N1893, N1890, N66, N512, N603);
nand NAND4 (N1894, N1892, N1024, N1059, N1774);
or OR4 (N1895, N1885, N1415, N908, N1204);
and AND4 (N1896, N1893, N1848, N321, N498);
not NOT1 (N1897, N1891);
xor XOR2 (N1898, N1857, N524);
nand NAND3 (N1899, N1897, N300, N424);
nand NAND4 (N1900, N1865, N1361, N1463, N794);
nor NOR3 (N1901, N1883, N385, N1410);
nor NOR4 (N1902, N1895, N1761, N18, N1659);
nand NAND3 (N1903, N1886, N1666, N528);
and AND4 (N1904, N1898, N188, N948, N119);
nand NAND3 (N1905, N1899, N1052, N1745);
xor XOR2 (N1906, N1903, N1110);
or OR4 (N1907, N1875, N501, N1268, N308);
nand NAND4 (N1908, N1861, N1791, N1527, N160);
buf BUF1 (N1909, N1900);
not NOT1 (N1910, N1896);
buf BUF1 (N1911, N1902);
nor NOR2 (N1912, N1905, N1043);
nand NAND3 (N1913, N1912, N146, N1279);
or OR3 (N1914, N1913, N692, N328);
nor NOR3 (N1915, N1906, N1221, N332);
nor NOR4 (N1916, N1907, N1351, N672, N568);
buf BUF1 (N1917, N1901);
nand NAND3 (N1918, N1904, N1445, N187);
buf BUF1 (N1919, N1915);
nor NOR3 (N1920, N1918, N35, N1569);
nor NOR4 (N1921, N1911, N142, N459, N1462);
buf BUF1 (N1922, N1908);
or OR4 (N1923, N1916, N1004, N1281, N1526);
and AND2 (N1924, N1894, N593);
or OR2 (N1925, N1923, N1585);
nor NOR3 (N1926, N1924, N937, N1456);
not NOT1 (N1927, N1910);
and AND2 (N1928, N1917, N1524);
nor NOR4 (N1929, N1909, N1112, N1000, N1880);
and AND3 (N1930, N1929, N141, N205);
nand NAND3 (N1931, N1919, N721, N1512);
or OR2 (N1932, N1926, N711);
or OR2 (N1933, N1920, N465);
and AND2 (N1934, N1914, N1782);
and AND4 (N1935, N1930, N466, N282, N40);
not NOT1 (N1936, N1928);
not NOT1 (N1937, N1925);
nor NOR2 (N1938, N1931, N410);
not NOT1 (N1939, N1938);
nor NOR2 (N1940, N1936, N1776);
or OR2 (N1941, N1921, N837);
xor XOR2 (N1942, N1922, N1636);
and AND3 (N1943, N1939, N746, N225);
and AND4 (N1944, N1943, N937, N11, N339);
or OR2 (N1945, N1941, N1868);
not NOT1 (N1946, N1932);
or OR2 (N1947, N1937, N860);
or OR3 (N1948, N1935, N1342, N1456);
nor NOR4 (N1949, N1944, N471, N994, N38);
xor XOR2 (N1950, N1949, N1247);
buf BUF1 (N1951, N1948);
or OR4 (N1952, N1942, N151, N1497, N235);
and AND4 (N1953, N1950, N716, N1116, N572);
buf BUF1 (N1954, N1934);
and AND2 (N1955, N1953, N1467);
xor XOR2 (N1956, N1951, N885);
and AND2 (N1957, N1927, N352);
xor XOR2 (N1958, N1956, N1141);
not NOT1 (N1959, N1946);
xor XOR2 (N1960, N1954, N1037);
not NOT1 (N1961, N1945);
nor NOR3 (N1962, N1958, N1251, N903);
not NOT1 (N1963, N1940);
nand NAND3 (N1964, N1952, N537, N1470);
xor XOR2 (N1965, N1959, N1249);
buf BUF1 (N1966, N1964);
nor NOR2 (N1967, N1966, N1053);
not NOT1 (N1968, N1967);
nand NAND4 (N1969, N1968, N807, N472, N875);
buf BUF1 (N1970, N1965);
and AND4 (N1971, N1961, N665, N94, N1190);
and AND4 (N1972, N1970, N538, N620, N644);
nand NAND4 (N1973, N1957, N418, N675, N1315);
and AND4 (N1974, N1955, N146, N1389, N208);
buf BUF1 (N1975, N1972);
not NOT1 (N1976, N1963);
or OR2 (N1977, N1971, N266);
buf BUF1 (N1978, N1962);
xor XOR2 (N1979, N1977, N1851);
and AND3 (N1980, N1973, N7, N1320);
and AND4 (N1981, N1960, N1085, N1332, N846);
or OR3 (N1982, N1978, N1553, N1165);
xor XOR2 (N1983, N1947, N1141);
not NOT1 (N1984, N1974);
nor NOR4 (N1985, N1979, N168, N283, N1078);
not NOT1 (N1986, N1969);
nand NAND2 (N1987, N1980, N1640);
nand NAND2 (N1988, N1985, N299);
nand NAND2 (N1989, N1981, N19);
xor XOR2 (N1990, N1983, N1817);
xor XOR2 (N1991, N1988, N800);
nand NAND4 (N1992, N1990, N1881, N693, N931);
not NOT1 (N1993, N1984);
and AND3 (N1994, N1993, N294, N660);
xor XOR2 (N1995, N1994, N542);
nand NAND2 (N1996, N1991, N1790);
xor XOR2 (N1997, N1975, N1456);
not NOT1 (N1998, N1976);
nor NOR2 (N1999, N1998, N1329);
buf BUF1 (N2000, N1997);
and AND2 (N2001, N1933, N194);
and AND4 (N2002, N2001, N1739, N1265, N1474);
and AND4 (N2003, N1992, N701, N863, N538);
buf BUF1 (N2004, N2002);
xor XOR2 (N2005, N2003, N62);
and AND3 (N2006, N1996, N713, N1837);
nand NAND3 (N2007, N2000, N1803, N1378);
nand NAND2 (N2008, N2006, N559);
nand NAND2 (N2009, N2007, N1948);
not NOT1 (N2010, N2009);
xor XOR2 (N2011, N2005, N1278);
not NOT1 (N2012, N2010);
or OR3 (N2013, N1995, N974, N1411);
and AND4 (N2014, N1987, N107, N147, N1003);
nand NAND2 (N2015, N2004, N1010);
nor NOR4 (N2016, N2011, N1311, N386, N38);
not NOT1 (N2017, N1999);
xor XOR2 (N2018, N1989, N2006);
and AND4 (N2019, N2017, N118, N698, N777);
endmodule