// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N796,N813,N808,N806,N818,N817,N815,N811,N814,N819;

buf BUF1 (N20, N5);
and AND4 (N21, N19, N4, N5, N1);
nand NAND3 (N22, N10, N18, N7);
nand NAND4 (N23, N7, N6, N18, N22);
xor XOR2 (N24, N10, N3);
nand NAND4 (N25, N13, N19, N5, N20);
nand NAND4 (N26, N5, N22, N25, N12);
not NOT1 (N27, N4);
xor XOR2 (N28, N12, N18);
nor NOR2 (N29, N15, N23);
xor XOR2 (N30, N11, N1);
or OR3 (N31, N19, N2, N16);
and AND2 (N32, N20, N11);
nand NAND3 (N33, N13, N15, N5);
and AND3 (N34, N32, N10, N25);
nor NOR2 (N35, N28, N11);
and AND4 (N36, N33, N15, N10, N10);
nor NOR2 (N37, N34, N35);
nand NAND2 (N38, N21, N21);
not NOT1 (N39, N12);
nor NOR3 (N40, N29, N34, N37);
xor XOR2 (N41, N8, N12);
not NOT1 (N42, N26);
xor XOR2 (N43, N40, N12);
buf BUF1 (N44, N31);
not NOT1 (N45, N39);
nand NAND2 (N46, N24, N9);
not NOT1 (N47, N38);
buf BUF1 (N48, N41);
not NOT1 (N49, N46);
xor XOR2 (N50, N49, N6);
or OR2 (N51, N44, N30);
buf BUF1 (N52, N23);
or OR4 (N53, N52, N21, N21, N22);
nand NAND3 (N54, N43, N42, N17);
nand NAND4 (N55, N41, N40, N49, N51);
not NOT1 (N56, N37);
xor XOR2 (N57, N55, N8);
nand NAND2 (N58, N53, N31);
not NOT1 (N59, N58);
buf BUF1 (N60, N45);
not NOT1 (N61, N48);
and AND2 (N62, N60, N57);
nand NAND3 (N63, N12, N49, N39);
xor XOR2 (N64, N61, N21);
xor XOR2 (N65, N63, N16);
nand NAND4 (N66, N50, N65, N57, N35);
or OR4 (N67, N44, N59, N17, N56);
buf BUF1 (N68, N48);
nand NAND4 (N69, N64, N9, N46, N37);
and AND3 (N70, N38, N69, N19);
not NOT1 (N71, N55);
buf BUF1 (N72, N68);
and AND4 (N73, N71, N70, N9, N20);
and AND4 (N74, N55, N66, N40, N58);
not NOT1 (N75, N27);
and AND3 (N76, N61, N51, N41);
nand NAND3 (N77, N62, N31, N35);
and AND3 (N78, N36, N9, N22);
nand NAND2 (N79, N73, N9);
nor NOR3 (N80, N77, N12, N18);
nand NAND4 (N81, N67, N20, N70, N46);
xor XOR2 (N82, N76, N16);
and AND3 (N83, N79, N67, N4);
nor NOR3 (N84, N80, N48, N38);
or OR3 (N85, N75, N71, N62);
or OR4 (N86, N83, N18, N78, N81);
not NOT1 (N87, N86);
buf BUF1 (N88, N44);
buf BUF1 (N89, N39);
nand NAND2 (N90, N85, N14);
or OR3 (N91, N54, N70, N63);
not NOT1 (N92, N91);
xor XOR2 (N93, N84, N48);
and AND2 (N94, N93, N7);
buf BUF1 (N95, N94);
nand NAND4 (N96, N88, N62, N20, N36);
nand NAND4 (N97, N90, N30, N31, N12);
xor XOR2 (N98, N82, N15);
not NOT1 (N99, N72);
not NOT1 (N100, N99);
xor XOR2 (N101, N100, N61);
xor XOR2 (N102, N95, N99);
and AND3 (N103, N96, N46, N97);
nand NAND2 (N104, N51, N5);
and AND4 (N105, N92, N60, N58, N86);
nand NAND2 (N106, N74, N45);
xor XOR2 (N107, N89, N82);
nand NAND3 (N108, N87, N40, N76);
or OR4 (N109, N98, N15, N12, N54);
buf BUF1 (N110, N102);
and AND2 (N111, N105, N37);
and AND4 (N112, N108, N6, N27, N111);
nand NAND3 (N113, N67, N65, N63);
and AND2 (N114, N110, N3);
and AND3 (N115, N101, N106, N111);
nand NAND4 (N116, N22, N91, N92, N93);
or OR4 (N117, N107, N64, N82, N69);
or OR3 (N118, N103, N90, N87);
or OR4 (N119, N117, N52, N12, N49);
nor NOR3 (N120, N104, N55, N13);
nor NOR4 (N121, N116, N18, N114, N53);
xor XOR2 (N122, N49, N28);
and AND2 (N123, N121, N23);
nor NOR4 (N124, N115, N64, N74, N21);
or OR2 (N125, N118, N88);
or OR2 (N126, N47, N50);
nor NOR2 (N127, N109, N126);
not NOT1 (N128, N118);
nor NOR2 (N129, N112, N91);
and AND2 (N130, N120, N27);
xor XOR2 (N131, N124, N104);
nor NOR3 (N132, N119, N38, N98);
nand NAND2 (N133, N127, N55);
not NOT1 (N134, N123);
not NOT1 (N135, N113);
nor NOR4 (N136, N130, N36, N10, N43);
buf BUF1 (N137, N125);
nand NAND4 (N138, N132, N132, N102, N47);
buf BUF1 (N139, N136);
not NOT1 (N140, N134);
nand NAND2 (N141, N137, N83);
nor NOR4 (N142, N141, N73, N73, N18);
and AND3 (N143, N135, N55, N33);
nor NOR4 (N144, N139, N51, N44, N32);
or OR4 (N145, N133, N139, N76, N2);
xor XOR2 (N146, N128, N135);
or OR4 (N147, N131, N144, N139, N15);
buf BUF1 (N148, N76);
or OR2 (N149, N142, N49);
nor NOR3 (N150, N146, N41, N59);
nor NOR4 (N151, N145, N46, N89, N116);
and AND2 (N152, N140, N112);
and AND2 (N153, N147, N4);
buf BUF1 (N154, N149);
nand NAND3 (N155, N143, N95, N29);
buf BUF1 (N156, N138);
nand NAND3 (N157, N151, N14, N124);
or OR3 (N158, N153, N45, N51);
buf BUF1 (N159, N155);
and AND4 (N160, N148, N72, N43, N36);
nand NAND4 (N161, N154, N36, N79, N94);
xor XOR2 (N162, N160, N128);
nor NOR2 (N163, N152, N101);
not NOT1 (N164, N158);
buf BUF1 (N165, N129);
not NOT1 (N166, N163);
xor XOR2 (N167, N162, N131);
not NOT1 (N168, N122);
buf BUF1 (N169, N159);
buf BUF1 (N170, N165);
xor XOR2 (N171, N168, N78);
xor XOR2 (N172, N157, N47);
buf BUF1 (N173, N166);
not NOT1 (N174, N173);
and AND2 (N175, N174, N24);
or OR4 (N176, N167, N86, N166, N60);
not NOT1 (N177, N170);
nand NAND2 (N178, N169, N34);
xor XOR2 (N179, N177, N124);
xor XOR2 (N180, N171, N111);
not NOT1 (N181, N178);
and AND4 (N182, N161, N64, N181, N152);
not NOT1 (N183, N179);
not NOT1 (N184, N146);
and AND2 (N185, N176, N46);
xor XOR2 (N186, N164, N155);
or OR4 (N187, N172, N50, N148, N75);
xor XOR2 (N188, N175, N182);
or OR4 (N189, N183, N78, N63, N106);
not NOT1 (N190, N101);
nand NAND2 (N191, N188, N101);
nand NAND2 (N192, N186, N31);
xor XOR2 (N193, N184, N134);
and AND3 (N194, N192, N114, N2);
nand NAND2 (N195, N156, N174);
not NOT1 (N196, N189);
buf BUF1 (N197, N193);
and AND2 (N198, N194, N40);
buf BUF1 (N199, N185);
or OR4 (N200, N197, N138, N195, N18);
and AND3 (N201, N16, N23, N105);
nand NAND2 (N202, N198, N126);
not NOT1 (N203, N201);
and AND4 (N204, N202, N2, N123, N155);
nor NOR4 (N205, N180, N35, N63, N73);
or OR4 (N206, N191, N124, N170, N9);
not NOT1 (N207, N200);
buf BUF1 (N208, N187);
and AND2 (N209, N204, N74);
and AND4 (N210, N207, N183, N9, N138);
buf BUF1 (N211, N199);
not NOT1 (N212, N203);
nand NAND2 (N213, N210, N22);
xor XOR2 (N214, N212, N73);
nand NAND2 (N215, N211, N176);
not NOT1 (N216, N209);
xor XOR2 (N217, N190, N149);
xor XOR2 (N218, N206, N77);
xor XOR2 (N219, N217, N161);
nor NOR4 (N220, N215, N69, N140, N210);
or OR2 (N221, N213, N107);
buf BUF1 (N222, N205);
nand NAND3 (N223, N220, N36, N162);
and AND3 (N224, N218, N170, N214);
and AND2 (N225, N190, N133);
not NOT1 (N226, N224);
nand NAND3 (N227, N221, N127, N81);
xor XOR2 (N228, N219, N226);
and AND2 (N229, N12, N198);
buf BUF1 (N230, N227);
nand NAND3 (N231, N150, N119, N25);
nand NAND4 (N232, N196, N156, N90, N20);
not NOT1 (N233, N229);
nand NAND2 (N234, N231, N184);
nor NOR4 (N235, N234, N46, N19, N214);
nor NOR2 (N236, N228, N94);
or OR3 (N237, N223, N107, N188);
and AND3 (N238, N235, N189, N33);
xor XOR2 (N239, N225, N157);
not NOT1 (N240, N208);
and AND4 (N241, N230, N22, N197, N182);
or OR4 (N242, N238, N78, N87, N219);
nor NOR4 (N243, N236, N223, N242, N25);
nor NOR3 (N244, N118, N50, N59);
not NOT1 (N245, N233);
buf BUF1 (N246, N222);
nand NAND2 (N247, N232, N38);
nor NOR2 (N248, N244, N9);
nor NOR4 (N249, N248, N196, N144, N94);
and AND3 (N250, N243, N173, N184);
nor NOR4 (N251, N245, N168, N176, N224);
nand NAND2 (N252, N246, N219);
or OR2 (N253, N237, N200);
xor XOR2 (N254, N252, N28);
not NOT1 (N255, N216);
buf BUF1 (N256, N254);
nand NAND4 (N257, N253, N229, N118, N18);
nor NOR2 (N258, N255, N164);
or OR2 (N259, N241, N20);
not NOT1 (N260, N249);
xor XOR2 (N261, N240, N145);
not NOT1 (N262, N260);
nor NOR2 (N263, N262, N159);
xor XOR2 (N264, N251, N247);
buf BUF1 (N265, N215);
or OR4 (N266, N258, N242, N179, N152);
and AND3 (N267, N239, N197, N39);
not NOT1 (N268, N259);
nand NAND3 (N269, N263, N56, N79);
not NOT1 (N270, N268);
not NOT1 (N271, N250);
xor XOR2 (N272, N256, N245);
nor NOR3 (N273, N269, N257, N270);
xor XOR2 (N274, N214, N213);
or OR3 (N275, N175, N130, N131);
buf BUF1 (N276, N265);
and AND3 (N277, N266, N136, N129);
xor XOR2 (N278, N274, N250);
nand NAND4 (N279, N271, N260, N230, N150);
nand NAND3 (N280, N275, N31, N14);
xor XOR2 (N281, N280, N252);
buf BUF1 (N282, N279);
and AND3 (N283, N267, N259, N143);
buf BUF1 (N284, N264);
xor XOR2 (N285, N261, N50);
and AND3 (N286, N285, N69, N5);
nand NAND2 (N287, N273, N121);
xor XOR2 (N288, N286, N37);
nand NAND4 (N289, N287, N104, N272, N84);
and AND3 (N290, N274, N97, N288);
nor NOR4 (N291, N33, N120, N60, N117);
and AND4 (N292, N276, N290, N261, N96);
not NOT1 (N293, N39);
nor NOR4 (N294, N278, N85, N80, N184);
buf BUF1 (N295, N283);
or OR4 (N296, N289, N62, N220, N269);
nor NOR2 (N297, N293, N212);
xor XOR2 (N298, N291, N246);
not NOT1 (N299, N277);
or OR2 (N300, N298, N118);
not NOT1 (N301, N281);
and AND2 (N302, N282, N125);
nand NAND3 (N303, N299, N280, N155);
nor NOR3 (N304, N301, N67, N32);
xor XOR2 (N305, N302, N14);
xor XOR2 (N306, N304, N255);
nor NOR3 (N307, N296, N84, N212);
nor NOR4 (N308, N305, N303, N267, N12);
buf BUF1 (N309, N158);
nor NOR4 (N310, N292, N172, N81, N242);
nand NAND4 (N311, N310, N100, N150, N208);
nor NOR4 (N312, N294, N22, N2, N207);
xor XOR2 (N313, N284, N17);
not NOT1 (N314, N313);
nand NAND2 (N315, N297, N238);
not NOT1 (N316, N311);
not NOT1 (N317, N315);
and AND3 (N318, N317, N269, N15);
nand NAND4 (N319, N307, N107, N156, N172);
nor NOR4 (N320, N312, N236, N33, N256);
not NOT1 (N321, N306);
and AND4 (N322, N308, N303, N247, N269);
nor NOR4 (N323, N300, N298, N65, N207);
or OR4 (N324, N295, N56, N22, N192);
or OR4 (N325, N324, N175, N77, N258);
and AND4 (N326, N318, N233, N314, N33);
not NOT1 (N327, N164);
nor NOR4 (N328, N309, N157, N72, N141);
buf BUF1 (N329, N327);
nor NOR3 (N330, N326, N157, N327);
not NOT1 (N331, N328);
buf BUF1 (N332, N330);
xor XOR2 (N333, N322, N286);
buf BUF1 (N334, N316);
nand NAND2 (N335, N334, N141);
nand NAND4 (N336, N331, N39, N293, N92);
buf BUF1 (N337, N336);
not NOT1 (N338, N333);
nand NAND4 (N339, N325, N94, N50, N221);
or OR4 (N340, N320, N183, N338, N67);
and AND3 (N341, N61, N64, N22);
or OR2 (N342, N340, N149);
and AND3 (N343, N342, N265, N79);
nor NOR4 (N344, N339, N318, N27, N322);
xor XOR2 (N345, N344, N60);
xor XOR2 (N346, N343, N189);
xor XOR2 (N347, N335, N12);
nand NAND4 (N348, N321, N54, N10, N118);
not NOT1 (N349, N337);
or OR3 (N350, N323, N93, N197);
or OR3 (N351, N332, N50, N113);
and AND2 (N352, N347, N169);
buf BUF1 (N353, N349);
buf BUF1 (N354, N345);
nor NOR2 (N355, N354, N21);
nand NAND4 (N356, N350, N8, N332, N204);
buf BUF1 (N357, N355);
and AND2 (N358, N319, N138);
and AND4 (N359, N358, N132, N48, N250);
nand NAND2 (N360, N353, N111);
buf BUF1 (N361, N359);
buf BUF1 (N362, N329);
nor NOR2 (N363, N361, N50);
xor XOR2 (N364, N348, N26);
xor XOR2 (N365, N357, N288);
not NOT1 (N366, N351);
or OR3 (N367, N366, N193, N306);
and AND3 (N368, N365, N283, N29);
nor NOR4 (N369, N341, N324, N167, N92);
nor NOR3 (N370, N352, N9, N324);
nor NOR3 (N371, N362, N216, N45);
and AND4 (N372, N369, N317, N306, N194);
buf BUF1 (N373, N363);
nor NOR3 (N374, N367, N152, N36);
xor XOR2 (N375, N373, N34);
nor NOR2 (N376, N364, N204);
nor NOR3 (N377, N375, N47, N278);
and AND2 (N378, N374, N24);
xor XOR2 (N379, N346, N160);
xor XOR2 (N380, N368, N232);
not NOT1 (N381, N371);
nand NAND3 (N382, N360, N215, N321);
buf BUF1 (N383, N370);
nand NAND2 (N384, N378, N364);
nor NOR4 (N385, N383, N5, N123, N132);
or OR4 (N386, N356, N267, N384, N52);
nand NAND4 (N387, N386, N280, N179, N207);
nor NOR2 (N388, N112, N277);
nand NAND4 (N389, N381, N306, N307, N319);
not NOT1 (N390, N379);
xor XOR2 (N391, N372, N82);
not NOT1 (N392, N385);
not NOT1 (N393, N391);
xor XOR2 (N394, N388, N383);
buf BUF1 (N395, N377);
or OR2 (N396, N389, N154);
and AND4 (N397, N393, N100, N168, N300);
not NOT1 (N398, N397);
and AND3 (N399, N390, N217, N86);
nor NOR3 (N400, N395, N293, N361);
nor NOR4 (N401, N399, N193, N141, N211);
and AND4 (N402, N401, N13, N235, N277);
nand NAND4 (N403, N380, N145, N311, N265);
nand NAND2 (N404, N394, N122);
xor XOR2 (N405, N387, N361);
xor XOR2 (N406, N402, N290);
nor NOR2 (N407, N405, N16);
buf BUF1 (N408, N382);
nor NOR3 (N409, N400, N334, N254);
nand NAND3 (N410, N403, N44, N86);
xor XOR2 (N411, N406, N26);
and AND3 (N412, N409, N305, N406);
nand NAND3 (N413, N410, N300, N398);
nor NOR4 (N414, N161, N38, N318, N221);
nor NOR4 (N415, N413, N402, N81, N149);
nand NAND2 (N416, N408, N195);
nor NOR4 (N417, N415, N284, N273, N155);
and AND4 (N418, N407, N74, N294, N73);
xor XOR2 (N419, N392, N99);
xor XOR2 (N420, N376, N34);
not NOT1 (N421, N412);
buf BUF1 (N422, N404);
nor NOR4 (N423, N396, N141, N67, N308);
not NOT1 (N424, N421);
nand NAND2 (N425, N417, N233);
not NOT1 (N426, N419);
and AND3 (N427, N414, N66, N86);
buf BUF1 (N428, N420);
or OR4 (N429, N416, N421, N334, N43);
not NOT1 (N430, N428);
nor NOR2 (N431, N411, N423);
xor XOR2 (N432, N295, N34);
buf BUF1 (N433, N418);
not NOT1 (N434, N431);
and AND2 (N435, N425, N133);
nand NAND2 (N436, N426, N251);
xor XOR2 (N437, N422, N360);
or OR2 (N438, N424, N216);
xor XOR2 (N439, N437, N262);
xor XOR2 (N440, N434, N385);
xor XOR2 (N441, N427, N423);
xor XOR2 (N442, N432, N52);
not NOT1 (N443, N433);
or OR3 (N444, N435, N371, N436);
buf BUF1 (N445, N61);
and AND3 (N446, N444, N119, N337);
xor XOR2 (N447, N442, N81);
xor XOR2 (N448, N429, N157);
buf BUF1 (N449, N441);
or OR2 (N450, N446, N432);
nor NOR4 (N451, N449, N332, N156, N293);
buf BUF1 (N452, N443);
nand NAND4 (N453, N440, N316, N65, N152);
nor NOR4 (N454, N453, N82, N298, N22);
nand NAND2 (N455, N451, N321);
or OR2 (N456, N452, N391);
nand NAND4 (N457, N439, N347, N71, N326);
buf BUF1 (N458, N430);
buf BUF1 (N459, N458);
xor XOR2 (N460, N448, N11);
xor XOR2 (N461, N450, N418);
nand NAND4 (N462, N457, N410, N99, N123);
buf BUF1 (N463, N445);
xor XOR2 (N464, N456, N117);
not NOT1 (N465, N460);
nor NOR3 (N466, N465, N2, N331);
not NOT1 (N467, N438);
buf BUF1 (N468, N463);
nor NOR2 (N469, N467, N184);
and AND2 (N470, N466, N339);
xor XOR2 (N471, N459, N124);
buf BUF1 (N472, N469);
nor NOR2 (N473, N464, N24);
or OR3 (N474, N461, N452, N416);
or OR4 (N475, N473, N303, N128, N346);
xor XOR2 (N476, N462, N5);
nor NOR2 (N477, N447, N125);
nand NAND4 (N478, N476, N79, N266, N157);
and AND4 (N479, N474, N120, N350, N346);
and AND2 (N480, N477, N310);
or OR2 (N481, N455, N51);
nand NAND3 (N482, N481, N218, N236);
nor NOR2 (N483, N468, N471);
nand NAND3 (N484, N111, N169, N379);
or OR2 (N485, N484, N332);
not NOT1 (N486, N478);
xor XOR2 (N487, N454, N321);
nand NAND3 (N488, N479, N202, N315);
buf BUF1 (N489, N488);
nand NAND4 (N490, N485, N47, N92, N469);
nand NAND3 (N491, N480, N123, N280);
buf BUF1 (N492, N489);
not NOT1 (N493, N487);
not NOT1 (N494, N492);
buf BUF1 (N495, N482);
xor XOR2 (N496, N475, N266);
not NOT1 (N497, N490);
nor NOR4 (N498, N493, N253, N274, N112);
xor XOR2 (N499, N494, N376);
and AND4 (N500, N486, N410, N443, N414);
nand NAND4 (N501, N495, N186, N452, N119);
nor NOR3 (N502, N500, N117, N307);
buf BUF1 (N503, N498);
xor XOR2 (N504, N501, N89);
or OR3 (N505, N491, N50, N467);
not NOT1 (N506, N483);
or OR4 (N507, N503, N65, N243, N192);
buf BUF1 (N508, N506);
or OR2 (N509, N497, N171);
buf BUF1 (N510, N509);
buf BUF1 (N511, N472);
nand NAND4 (N512, N504, N263, N366, N17);
and AND2 (N513, N499, N454);
nand NAND2 (N514, N511, N110);
nand NAND4 (N515, N470, N183, N375, N247);
nand NAND2 (N516, N507, N271);
nand NAND3 (N517, N515, N99, N14);
or OR2 (N518, N517, N453);
or OR3 (N519, N505, N340, N399);
buf BUF1 (N520, N508);
nand NAND3 (N521, N520, N235, N208);
xor XOR2 (N522, N513, N139);
xor XOR2 (N523, N512, N195);
or OR2 (N524, N496, N331);
buf BUF1 (N525, N502);
buf BUF1 (N526, N524);
not NOT1 (N527, N514);
nand NAND2 (N528, N525, N213);
not NOT1 (N529, N527);
nand NAND4 (N530, N519, N252, N492, N94);
nand NAND3 (N531, N523, N517, N433);
xor XOR2 (N532, N516, N304);
not NOT1 (N533, N528);
and AND2 (N534, N531, N153);
nor NOR4 (N535, N522, N66, N332, N18);
or OR2 (N536, N534, N470);
or OR4 (N537, N533, N423, N355, N48);
xor XOR2 (N538, N530, N87);
not NOT1 (N539, N510);
nor NOR3 (N540, N538, N531, N525);
xor XOR2 (N541, N536, N241);
nor NOR2 (N542, N532, N286);
and AND4 (N543, N542, N27, N256, N231);
or OR4 (N544, N541, N286, N167, N247);
nor NOR3 (N545, N543, N205, N30);
and AND2 (N546, N539, N376);
nand NAND3 (N547, N535, N541, N281);
buf BUF1 (N548, N518);
or OR3 (N549, N521, N6, N157);
nor NOR4 (N550, N529, N242, N220, N402);
xor XOR2 (N551, N526, N59);
nor NOR2 (N552, N545, N472);
nand NAND4 (N553, N552, N125, N133, N448);
not NOT1 (N554, N550);
nand NAND3 (N555, N553, N433, N508);
nor NOR4 (N556, N544, N439, N385, N62);
buf BUF1 (N557, N551);
not NOT1 (N558, N554);
buf BUF1 (N559, N547);
xor XOR2 (N560, N556, N176);
or OR3 (N561, N558, N319, N368);
nor NOR4 (N562, N537, N462, N110, N542);
nand NAND4 (N563, N562, N323, N329, N74);
xor XOR2 (N564, N559, N250);
and AND2 (N565, N555, N118);
and AND2 (N566, N563, N359);
or OR3 (N567, N560, N339, N60);
nor NOR2 (N568, N557, N130);
not NOT1 (N569, N564);
and AND4 (N570, N565, N239, N280, N363);
not NOT1 (N571, N548);
buf BUF1 (N572, N561);
or OR3 (N573, N572, N329, N413);
not NOT1 (N574, N573);
or OR4 (N575, N540, N195, N275, N28);
buf BUF1 (N576, N571);
xor XOR2 (N577, N566, N174);
not NOT1 (N578, N568);
xor XOR2 (N579, N549, N315);
and AND4 (N580, N570, N70, N280, N289);
nand NAND3 (N581, N567, N3, N170);
not NOT1 (N582, N577);
nand NAND3 (N583, N574, N526, N560);
nand NAND3 (N584, N583, N382, N422);
nand NAND4 (N585, N546, N386, N424, N217);
nand NAND3 (N586, N584, N561, N470);
nand NAND4 (N587, N586, N512, N25, N414);
and AND3 (N588, N582, N401, N273);
or OR3 (N589, N585, N131, N550);
or OR4 (N590, N569, N85, N556, N192);
buf BUF1 (N591, N580);
buf BUF1 (N592, N578);
xor XOR2 (N593, N587, N363);
or OR2 (N594, N593, N104);
nor NOR2 (N595, N592, N577);
not NOT1 (N596, N589);
not NOT1 (N597, N575);
not NOT1 (N598, N597);
xor XOR2 (N599, N590, N554);
or OR2 (N600, N579, N63);
or OR4 (N601, N591, N445, N67, N506);
xor XOR2 (N602, N596, N13);
xor XOR2 (N603, N595, N305);
not NOT1 (N604, N603);
nor NOR4 (N605, N600, N358, N309, N279);
nand NAND3 (N606, N598, N569, N531);
not NOT1 (N607, N605);
not NOT1 (N608, N594);
not NOT1 (N609, N606);
xor XOR2 (N610, N604, N558);
not NOT1 (N611, N599);
nand NAND2 (N612, N576, N409);
or OR2 (N613, N602, N388);
buf BUF1 (N614, N609);
buf BUF1 (N615, N613);
buf BUF1 (N616, N611);
and AND4 (N617, N601, N539, N403, N536);
nor NOR2 (N618, N607, N469);
and AND3 (N619, N588, N284, N213);
xor XOR2 (N620, N618, N211);
or OR2 (N621, N619, N562);
and AND4 (N622, N612, N379, N437, N219);
and AND2 (N623, N620, N19);
or OR2 (N624, N581, N386);
and AND2 (N625, N624, N169);
nand NAND3 (N626, N616, N531, N394);
nand NAND3 (N627, N615, N500, N209);
xor XOR2 (N628, N608, N532);
buf BUF1 (N629, N621);
and AND4 (N630, N626, N305, N378, N10);
nand NAND3 (N631, N628, N308, N117);
buf BUF1 (N632, N623);
not NOT1 (N633, N625);
nand NAND3 (N634, N629, N230, N64);
and AND2 (N635, N634, N491);
not NOT1 (N636, N610);
buf BUF1 (N637, N622);
buf BUF1 (N638, N633);
nand NAND2 (N639, N637, N329);
and AND2 (N640, N635, N114);
nor NOR4 (N641, N627, N264, N341, N351);
buf BUF1 (N642, N631);
or OR3 (N643, N617, N164, N143);
buf BUF1 (N644, N639);
and AND4 (N645, N630, N68, N609, N305);
buf BUF1 (N646, N644);
buf BUF1 (N647, N638);
buf BUF1 (N648, N646);
or OR3 (N649, N640, N61, N227);
xor XOR2 (N650, N645, N36);
xor XOR2 (N651, N647, N617);
not NOT1 (N652, N651);
buf BUF1 (N653, N642);
buf BUF1 (N654, N632);
nand NAND2 (N655, N649, N329);
buf BUF1 (N656, N636);
nor NOR2 (N657, N643, N288);
nor NOR2 (N658, N654, N465);
nor NOR2 (N659, N658, N395);
xor XOR2 (N660, N614, N629);
xor XOR2 (N661, N660, N228);
nor NOR2 (N662, N657, N238);
not NOT1 (N663, N662);
nand NAND2 (N664, N652, N477);
and AND2 (N665, N653, N370);
not NOT1 (N666, N641);
not NOT1 (N667, N656);
nand NAND3 (N668, N663, N121, N103);
or OR4 (N669, N661, N455, N28, N375);
buf BUF1 (N670, N659);
not NOT1 (N671, N655);
not NOT1 (N672, N667);
xor XOR2 (N673, N669, N654);
and AND3 (N674, N672, N18, N348);
or OR4 (N675, N674, N246, N155, N506);
nor NOR2 (N676, N675, N333);
not NOT1 (N677, N666);
nand NAND3 (N678, N650, N380, N471);
nand NAND3 (N679, N676, N310, N331);
nor NOR3 (N680, N665, N52, N90);
buf BUF1 (N681, N671);
or OR4 (N682, N648, N517, N677, N459);
not NOT1 (N683, N341);
not NOT1 (N684, N670);
nor NOR3 (N685, N664, N121, N238);
nor NOR3 (N686, N684, N384, N489);
or OR4 (N687, N683, N114, N249, N558);
and AND4 (N688, N678, N251, N345, N251);
or OR4 (N689, N688, N514, N520, N473);
nand NAND4 (N690, N682, N627, N674, N165);
or OR3 (N691, N690, N273, N648);
buf BUF1 (N692, N673);
buf BUF1 (N693, N687);
not NOT1 (N694, N685);
nand NAND2 (N695, N689, N501);
or OR4 (N696, N691, N115, N363, N164);
not NOT1 (N697, N668);
xor XOR2 (N698, N680, N642);
not NOT1 (N699, N679);
nand NAND2 (N700, N695, N116);
nor NOR2 (N701, N696, N399);
not NOT1 (N702, N697);
nand NAND2 (N703, N700, N416);
nor NOR3 (N704, N693, N60, N501);
not NOT1 (N705, N699);
or OR4 (N706, N702, N175, N181, N311);
buf BUF1 (N707, N704);
nand NAND2 (N708, N705, N499);
not NOT1 (N709, N706);
or OR3 (N710, N698, N419, N583);
nand NAND3 (N711, N694, N4, N604);
xor XOR2 (N712, N707, N465);
nor NOR2 (N713, N708, N503);
and AND2 (N714, N713, N508);
xor XOR2 (N715, N692, N637);
or OR3 (N716, N709, N194, N499);
and AND2 (N717, N703, N86);
not NOT1 (N718, N710);
nand NAND3 (N719, N686, N58, N642);
not NOT1 (N720, N716);
buf BUF1 (N721, N714);
nor NOR4 (N722, N712, N461, N386, N105);
xor XOR2 (N723, N719, N19);
and AND4 (N724, N718, N210, N281, N576);
or OR4 (N725, N681, N89, N535, N353);
xor XOR2 (N726, N717, N110);
nand NAND2 (N727, N725, N397);
xor XOR2 (N728, N724, N90);
not NOT1 (N729, N720);
nand NAND4 (N730, N723, N584, N122, N92);
nor NOR3 (N731, N701, N715, N655);
or OR4 (N732, N69, N628, N339, N580);
not NOT1 (N733, N722);
nor NOR4 (N734, N733, N258, N499, N219);
and AND2 (N735, N734, N221);
nor NOR2 (N736, N728, N171);
and AND3 (N737, N711, N524, N648);
xor XOR2 (N738, N735, N143);
xor XOR2 (N739, N721, N537);
not NOT1 (N740, N737);
not NOT1 (N741, N727);
not NOT1 (N742, N736);
xor XOR2 (N743, N732, N685);
nand NAND2 (N744, N726, N424);
xor XOR2 (N745, N743, N619);
nor NOR3 (N746, N730, N409, N312);
nor NOR2 (N747, N731, N39);
and AND3 (N748, N729, N199, N12);
or OR3 (N749, N742, N173, N148);
nor NOR2 (N750, N745, N127);
buf BUF1 (N751, N750);
and AND3 (N752, N740, N222, N701);
or OR3 (N753, N747, N337, N264);
not NOT1 (N754, N752);
buf BUF1 (N755, N744);
nor NOR4 (N756, N749, N285, N538, N538);
nand NAND4 (N757, N738, N601, N330, N512);
xor XOR2 (N758, N755, N346);
xor XOR2 (N759, N748, N514);
buf BUF1 (N760, N753);
or OR2 (N761, N746, N155);
xor XOR2 (N762, N741, N519);
buf BUF1 (N763, N759);
nand NAND2 (N764, N760, N361);
or OR4 (N765, N756, N446, N620, N55);
xor XOR2 (N766, N763, N622);
nand NAND3 (N767, N765, N482, N356);
nor NOR4 (N768, N764, N394, N142, N527);
xor XOR2 (N769, N758, N747);
nor NOR2 (N770, N769, N150);
or OR2 (N771, N766, N424);
buf BUF1 (N772, N739);
buf BUF1 (N773, N770);
and AND3 (N774, N772, N320, N453);
or OR2 (N775, N761, N4);
xor XOR2 (N776, N762, N570);
and AND4 (N777, N754, N716, N160, N32);
not NOT1 (N778, N776);
nand NAND4 (N779, N757, N648, N400, N414);
and AND2 (N780, N751, N436);
not NOT1 (N781, N768);
and AND2 (N782, N779, N273);
nand NAND3 (N783, N774, N195, N371);
or OR2 (N784, N775, N166);
nand NAND2 (N785, N784, N733);
and AND2 (N786, N767, N479);
buf BUF1 (N787, N777);
buf BUF1 (N788, N781);
buf BUF1 (N789, N786);
and AND4 (N790, N771, N785, N560, N340);
nand NAND4 (N791, N528, N263, N747, N497);
xor XOR2 (N792, N788, N612);
buf BUF1 (N793, N791);
xor XOR2 (N794, N793, N563);
xor XOR2 (N795, N780, N389);
not NOT1 (N796, N790);
or OR4 (N797, N783, N390, N168, N319);
buf BUF1 (N798, N794);
buf BUF1 (N799, N778);
nand NAND4 (N800, N795, N776, N595, N306);
not NOT1 (N801, N789);
nor NOR3 (N802, N799, N140, N159);
xor XOR2 (N803, N802, N258);
or OR3 (N804, N782, N325, N433);
buf BUF1 (N805, N792);
buf BUF1 (N806, N787);
or OR4 (N807, N801, N661, N391, N140);
buf BUF1 (N808, N797);
nand NAND4 (N809, N807, N120, N281, N748);
and AND2 (N810, N805, N702);
nor NOR4 (N811, N800, N663, N602, N661);
nor NOR2 (N812, N798, N748);
buf BUF1 (N813, N803);
and AND4 (N814, N809, N372, N9, N380);
and AND4 (N815, N804, N567, N344, N607);
and AND2 (N816, N773, N444);
not NOT1 (N817, N812);
nand NAND4 (N818, N810, N573, N782, N339);
and AND3 (N819, N816, N735, N535);
endmodule