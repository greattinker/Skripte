// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N4018,N4011,N4006,N4014,N3994,N4019,N4017,N4009,N4010,N4021;

or OR3 (N22, N7, N4, N13);
not NOT1 (N23, N9);
nor NOR2 (N24, N13, N15);
or OR4 (N25, N20, N2, N11, N24);
xor XOR2 (N26, N17, N8);
nor NOR3 (N27, N26, N2, N3);
and AND3 (N28, N12, N27, N12);
nor NOR3 (N29, N25, N26, N14);
buf BUF1 (N30, N22);
buf BUF1 (N31, N4);
xor XOR2 (N32, N5, N9);
not NOT1 (N33, N18);
xor XOR2 (N34, N19, N1);
xor XOR2 (N35, N20, N19);
nand NAND2 (N36, N12, N24);
nor NOR3 (N37, N34, N30, N1);
nor NOR3 (N38, N32, N3, N37);
or OR4 (N39, N36, N28, N12, N21);
nand NAND4 (N40, N20, N11, N3, N13);
and AND3 (N41, N2, N23, N36);
and AND3 (N42, N25, N10, N4);
or OR3 (N43, N33, N10, N9);
or OR4 (N44, N1, N25, N22, N34);
buf BUF1 (N45, N31);
and AND4 (N46, N44, N3, N26, N15);
buf BUF1 (N47, N42);
xor XOR2 (N48, N47, N39);
and AND3 (N49, N6, N26, N9);
and AND4 (N50, N46, N31, N31, N20);
or OR2 (N51, N40, N26);
nand NAND3 (N52, N38, N17, N39);
or OR2 (N53, N45, N36);
and AND3 (N54, N52, N17, N53);
or OR3 (N55, N22, N2, N49);
nand NAND3 (N56, N10, N47, N35);
or OR2 (N57, N36, N19);
nor NOR3 (N58, N50, N56, N21);
not NOT1 (N59, N40);
not NOT1 (N60, N55);
nand NAND3 (N61, N59, N53, N40);
buf BUF1 (N62, N48);
not NOT1 (N63, N51);
not NOT1 (N64, N63);
not NOT1 (N65, N54);
nand NAND4 (N66, N57, N23, N18, N38);
buf BUF1 (N67, N41);
not NOT1 (N68, N64);
not NOT1 (N69, N60);
not NOT1 (N70, N61);
buf BUF1 (N71, N29);
nand NAND2 (N72, N65, N52);
not NOT1 (N73, N62);
nand NAND2 (N74, N73, N33);
nor NOR3 (N75, N43, N73, N53);
nand NAND4 (N76, N75, N27, N34, N45);
or OR4 (N77, N72, N58, N8, N56);
xor XOR2 (N78, N51, N6);
nor NOR4 (N79, N70, N42, N49, N3);
and AND4 (N80, N74, N47, N42, N5);
nor NOR2 (N81, N78, N24);
nand NAND2 (N82, N66, N50);
nand NAND2 (N83, N68, N6);
nand NAND3 (N84, N76, N60, N18);
or OR4 (N85, N79, N77, N2, N27);
nand NAND4 (N86, N57, N9, N73, N78);
nand NAND4 (N87, N81, N51, N35, N78);
nor NOR3 (N88, N84, N42, N37);
xor XOR2 (N89, N88, N69);
not NOT1 (N90, N73);
buf BUF1 (N91, N82);
nand NAND4 (N92, N86, N77, N77, N17);
xor XOR2 (N93, N90, N6);
buf BUF1 (N94, N71);
xor XOR2 (N95, N87, N39);
or OR2 (N96, N92, N20);
or OR3 (N97, N80, N42, N58);
not NOT1 (N98, N97);
xor XOR2 (N99, N98, N52);
not NOT1 (N100, N94);
nand NAND3 (N101, N96, N100, N96);
or OR2 (N102, N91, N55);
or OR3 (N103, N34, N100, N76);
nor NOR2 (N104, N103, N95);
and AND3 (N105, N81, N86, N88);
and AND3 (N106, N83, N37, N70);
and AND3 (N107, N67, N50, N19);
and AND2 (N108, N85, N50);
buf BUF1 (N109, N93);
not NOT1 (N110, N99);
nand NAND3 (N111, N102, N77, N94);
or OR2 (N112, N104, N75);
not NOT1 (N113, N101);
and AND3 (N114, N111, N93, N52);
nand NAND3 (N115, N105, N73, N87);
nor NOR4 (N116, N109, N84, N62, N12);
and AND4 (N117, N114, N75, N28, N37);
not NOT1 (N118, N117);
nand NAND3 (N119, N118, N90, N24);
nor NOR2 (N120, N106, N34);
nor NOR3 (N121, N112, N112, N108);
xor XOR2 (N122, N38, N16);
and AND2 (N123, N120, N14);
nand NAND3 (N124, N121, N52, N48);
and AND4 (N125, N123, N60, N70, N34);
buf BUF1 (N126, N125);
nor NOR4 (N127, N89, N33, N101, N105);
or OR3 (N128, N124, N66, N106);
xor XOR2 (N129, N110, N85);
xor XOR2 (N130, N128, N45);
xor XOR2 (N131, N127, N85);
buf BUF1 (N132, N115);
nor NOR4 (N133, N129, N107, N62, N14);
buf BUF1 (N134, N32);
xor XOR2 (N135, N113, N127);
or OR3 (N136, N131, N43, N58);
and AND3 (N137, N136, N87, N114);
or OR3 (N138, N126, N114, N123);
not NOT1 (N139, N132);
buf BUF1 (N140, N122);
not NOT1 (N141, N140);
buf BUF1 (N142, N138);
nor NOR4 (N143, N134, N20, N62, N95);
and AND3 (N144, N130, N98, N111);
buf BUF1 (N145, N142);
nand NAND2 (N146, N145, N2);
xor XOR2 (N147, N116, N90);
nand NAND4 (N148, N133, N27, N147, N34);
not NOT1 (N149, N28);
nand NAND3 (N150, N137, N85, N43);
xor XOR2 (N151, N146, N11);
nor NOR3 (N152, N150, N8, N96);
xor XOR2 (N153, N151, N119);
not NOT1 (N154, N63);
or OR3 (N155, N139, N77, N10);
nor NOR4 (N156, N152, N1, N88, N121);
buf BUF1 (N157, N155);
buf BUF1 (N158, N144);
not NOT1 (N159, N135);
buf BUF1 (N160, N141);
buf BUF1 (N161, N160);
buf BUF1 (N162, N154);
buf BUF1 (N163, N159);
buf BUF1 (N164, N157);
xor XOR2 (N165, N156, N161);
xor XOR2 (N166, N91, N70);
or OR3 (N167, N158, N53, N108);
buf BUF1 (N168, N153);
and AND3 (N169, N164, N41, N146);
nand NAND2 (N170, N168, N60);
xor XOR2 (N171, N167, N24);
buf BUF1 (N172, N149);
xor XOR2 (N173, N162, N100);
and AND2 (N174, N166, N17);
or OR4 (N175, N174, N2, N152, N85);
nand NAND4 (N176, N165, N156, N145, N159);
nor NOR4 (N177, N172, N71, N21, N57);
nor NOR4 (N178, N163, N161, N26, N24);
or OR4 (N179, N175, N8, N153, N27);
or OR3 (N180, N143, N178, N96);
nor NOR2 (N181, N131, N161);
or OR4 (N182, N176, N81, N156, N29);
nor NOR4 (N183, N169, N142, N45, N38);
not NOT1 (N184, N181);
nand NAND2 (N185, N180, N168);
or OR4 (N186, N148, N144, N97, N97);
nand NAND4 (N187, N182, N144, N68, N27);
or OR2 (N188, N173, N41);
or OR2 (N189, N179, N34);
xor XOR2 (N190, N188, N165);
buf BUF1 (N191, N190);
nand NAND4 (N192, N187, N24, N62, N55);
not NOT1 (N193, N191);
xor XOR2 (N194, N171, N99);
buf BUF1 (N195, N185);
buf BUF1 (N196, N186);
not NOT1 (N197, N184);
not NOT1 (N198, N197);
nand NAND4 (N199, N198, N175, N70, N145);
buf BUF1 (N200, N170);
nor NOR3 (N201, N194, N136, N149);
nand NAND4 (N202, N201, N19, N163, N128);
and AND3 (N203, N200, N65, N66);
or OR3 (N204, N199, N26, N10);
and AND3 (N205, N203, N104, N151);
and AND2 (N206, N177, N53);
not NOT1 (N207, N204);
or OR2 (N208, N195, N18);
or OR4 (N209, N205, N8, N63, N8);
nor NOR4 (N210, N189, N148, N21, N161);
nor NOR2 (N211, N183, N75);
nor NOR4 (N212, N208, N139, N50, N27);
and AND3 (N213, N196, N21, N184);
or OR2 (N214, N211, N156);
xor XOR2 (N215, N193, N207);
not NOT1 (N216, N49);
buf BUF1 (N217, N216);
not NOT1 (N218, N206);
and AND3 (N219, N218, N176, N166);
not NOT1 (N220, N213);
xor XOR2 (N221, N219, N216);
or OR2 (N222, N215, N109);
nand NAND2 (N223, N221, N35);
buf BUF1 (N224, N214);
and AND4 (N225, N202, N201, N118, N53);
and AND4 (N226, N212, N177, N94, N10);
xor XOR2 (N227, N217, N129);
buf BUF1 (N228, N222);
nand NAND3 (N229, N228, N59, N111);
nor NOR4 (N230, N224, N228, N142, N133);
nor NOR3 (N231, N220, N107, N136);
buf BUF1 (N232, N226);
nor NOR4 (N233, N210, N7, N4, N111);
and AND2 (N234, N225, N185);
nand NAND2 (N235, N229, N210);
nor NOR4 (N236, N234, N208, N136, N157);
not NOT1 (N237, N227);
xor XOR2 (N238, N230, N104);
nand NAND3 (N239, N237, N106, N237);
nor NOR4 (N240, N235, N210, N121, N223);
buf BUF1 (N241, N185);
and AND4 (N242, N192, N124, N159, N119);
xor XOR2 (N243, N236, N198);
buf BUF1 (N244, N239);
or OR3 (N245, N238, N177, N4);
nand NAND3 (N246, N231, N95, N64);
or OR2 (N247, N232, N130);
buf BUF1 (N248, N244);
buf BUF1 (N249, N243);
nand NAND2 (N250, N240, N132);
xor XOR2 (N251, N249, N48);
not NOT1 (N252, N241);
xor XOR2 (N253, N250, N80);
nand NAND2 (N254, N252, N169);
buf BUF1 (N255, N254);
or OR3 (N256, N251, N115, N49);
buf BUF1 (N257, N248);
nand NAND2 (N258, N245, N69);
or OR4 (N259, N246, N121, N240, N22);
xor XOR2 (N260, N258, N161);
or OR3 (N261, N257, N27, N115);
xor XOR2 (N262, N261, N227);
nor NOR4 (N263, N255, N148, N216, N13);
nor NOR2 (N264, N209, N1);
and AND2 (N265, N263, N92);
or OR4 (N266, N233, N168, N125, N194);
not NOT1 (N267, N265);
xor XOR2 (N268, N264, N1);
or OR4 (N269, N268, N54, N25, N35);
nand NAND2 (N270, N262, N189);
nor NOR2 (N271, N266, N129);
and AND3 (N272, N253, N64, N14);
or OR2 (N273, N242, N130);
nand NAND2 (N274, N271, N103);
or OR3 (N275, N269, N122, N218);
nor NOR4 (N276, N259, N112, N61, N25);
buf BUF1 (N277, N247);
nand NAND3 (N278, N275, N145, N78);
not NOT1 (N279, N256);
nor NOR2 (N280, N270, N124);
nor NOR3 (N281, N278, N220, N251);
and AND3 (N282, N279, N73, N259);
or OR4 (N283, N281, N153, N229, N143);
not NOT1 (N284, N260);
or OR4 (N285, N272, N230, N126, N176);
xor XOR2 (N286, N285, N128);
not NOT1 (N287, N277);
buf BUF1 (N288, N286);
nor NOR2 (N289, N273, N72);
nand NAND4 (N290, N283, N256, N208, N158);
nor NOR3 (N291, N287, N127, N224);
not NOT1 (N292, N291);
not NOT1 (N293, N267);
buf BUF1 (N294, N289);
and AND3 (N295, N284, N281, N244);
and AND2 (N296, N295, N127);
nand NAND3 (N297, N290, N12, N203);
xor XOR2 (N298, N280, N6);
not NOT1 (N299, N297);
nor NOR3 (N300, N282, N127, N130);
nor NOR4 (N301, N293, N164, N246, N171);
nor NOR2 (N302, N276, N7);
and AND3 (N303, N300, N261, N243);
nand NAND3 (N304, N274, N231, N214);
and AND2 (N305, N288, N245);
not NOT1 (N306, N303);
buf BUF1 (N307, N301);
not NOT1 (N308, N306);
nand NAND4 (N309, N307, N234, N260, N88);
nor NOR2 (N310, N305, N39);
or OR3 (N311, N298, N78, N65);
buf BUF1 (N312, N309);
nand NAND4 (N313, N310, N49, N23, N35);
xor XOR2 (N314, N311, N120);
or OR4 (N315, N292, N244, N270, N78);
and AND2 (N316, N312, N247);
not NOT1 (N317, N314);
or OR3 (N318, N296, N213, N300);
nor NOR4 (N319, N318, N89, N246, N90);
nand NAND3 (N320, N316, N155, N314);
or OR4 (N321, N315, N31, N300, N192);
not NOT1 (N322, N317);
not NOT1 (N323, N299);
not NOT1 (N324, N321);
nand NAND4 (N325, N313, N260, N237, N249);
nor NOR3 (N326, N304, N24, N223);
and AND3 (N327, N326, N46, N263);
nand NAND3 (N328, N319, N164, N41);
or OR3 (N329, N328, N312, N282);
and AND4 (N330, N322, N273, N105, N251);
not NOT1 (N331, N308);
not NOT1 (N332, N330);
or OR4 (N333, N327, N320, N125, N16);
xor XOR2 (N334, N132, N40);
nor NOR4 (N335, N302, N37, N17, N147);
not NOT1 (N336, N334);
and AND4 (N337, N325, N108, N66, N274);
xor XOR2 (N338, N331, N81);
nor NOR4 (N339, N294, N66, N234, N107);
buf BUF1 (N340, N338);
or OR3 (N341, N323, N154, N321);
buf BUF1 (N342, N332);
nor NOR3 (N343, N341, N246, N157);
and AND3 (N344, N336, N179, N121);
nand NAND3 (N345, N340, N37, N214);
and AND3 (N346, N324, N307, N192);
nor NOR4 (N347, N343, N66, N325, N110);
xor XOR2 (N348, N342, N229);
xor XOR2 (N349, N329, N217);
buf BUF1 (N350, N339);
nor NOR3 (N351, N346, N95, N285);
nor NOR3 (N352, N348, N99, N126);
nor NOR3 (N353, N347, N57, N241);
nand NAND2 (N354, N352, N67);
not NOT1 (N355, N337);
or OR4 (N356, N335, N302, N210, N187);
and AND4 (N357, N345, N2, N286, N293);
or OR2 (N358, N333, N102);
not NOT1 (N359, N344);
and AND3 (N360, N359, N172, N112);
xor XOR2 (N361, N357, N64);
xor XOR2 (N362, N353, N239);
nand NAND4 (N363, N355, N131, N153, N139);
buf BUF1 (N364, N358);
xor XOR2 (N365, N356, N53);
xor XOR2 (N366, N351, N104);
or OR3 (N367, N360, N99, N22);
nor NOR4 (N368, N366, N278, N93, N152);
buf BUF1 (N369, N367);
not NOT1 (N370, N364);
xor XOR2 (N371, N370, N144);
nor NOR2 (N372, N362, N138);
nor NOR3 (N373, N349, N112, N191);
xor XOR2 (N374, N354, N126);
nand NAND3 (N375, N373, N353, N231);
and AND2 (N376, N350, N300);
or OR4 (N377, N363, N112, N171, N51);
nand NAND2 (N378, N376, N262);
or OR3 (N379, N361, N135, N271);
or OR3 (N380, N374, N122, N63);
nor NOR3 (N381, N379, N76, N325);
buf BUF1 (N382, N381);
not NOT1 (N383, N368);
nand NAND2 (N384, N372, N56);
and AND3 (N385, N382, N135, N209);
buf BUF1 (N386, N365);
xor XOR2 (N387, N380, N126);
or OR2 (N388, N383, N117);
or OR2 (N389, N377, N234);
xor XOR2 (N390, N375, N1);
nor NOR2 (N391, N371, N129);
and AND2 (N392, N385, N30);
nor NOR4 (N393, N391, N382, N220, N219);
not NOT1 (N394, N388);
not NOT1 (N395, N386);
nand NAND3 (N396, N387, N88, N15);
xor XOR2 (N397, N396, N354);
xor XOR2 (N398, N369, N159);
or OR2 (N399, N392, N279);
nor NOR2 (N400, N393, N146);
buf BUF1 (N401, N399);
nor NOR4 (N402, N378, N181, N211, N396);
xor XOR2 (N403, N402, N114);
buf BUF1 (N404, N397);
xor XOR2 (N405, N404, N2);
not NOT1 (N406, N395);
nor NOR3 (N407, N405, N393, N238);
buf BUF1 (N408, N398);
xor XOR2 (N409, N403, N67);
nand NAND2 (N410, N400, N344);
and AND4 (N411, N408, N90, N276, N4);
buf BUF1 (N412, N409);
nand NAND4 (N413, N410, N282, N50, N273);
or OR4 (N414, N389, N218, N294, N260);
or OR3 (N415, N411, N207, N109);
xor XOR2 (N416, N413, N359);
xor XOR2 (N417, N406, N371);
not NOT1 (N418, N390);
not NOT1 (N419, N407);
nor NOR2 (N420, N415, N408);
nand NAND2 (N421, N418, N320);
nand NAND3 (N422, N412, N216, N18);
and AND3 (N423, N414, N229, N211);
not NOT1 (N424, N394);
and AND3 (N425, N416, N273, N132);
nand NAND2 (N426, N424, N183);
not NOT1 (N427, N421);
and AND4 (N428, N417, N279, N334, N71);
or OR3 (N429, N420, N334, N256);
not NOT1 (N430, N419);
buf BUF1 (N431, N425);
and AND4 (N432, N384, N287, N342, N19);
nand NAND4 (N433, N432, N265, N24, N70);
not NOT1 (N434, N401);
or OR2 (N435, N422, N102);
buf BUF1 (N436, N426);
nor NOR3 (N437, N423, N53, N358);
nor NOR4 (N438, N437, N1, N201, N298);
and AND2 (N439, N434, N392);
buf BUF1 (N440, N436);
not NOT1 (N441, N440);
xor XOR2 (N442, N427, N268);
nor NOR2 (N443, N442, N89);
xor XOR2 (N444, N429, N380);
not NOT1 (N445, N438);
nor NOR3 (N446, N443, N360, N259);
nor NOR2 (N447, N441, N172);
not NOT1 (N448, N447);
xor XOR2 (N449, N439, N367);
or OR4 (N450, N428, N32, N119, N361);
or OR4 (N451, N445, N289, N3, N12);
nand NAND2 (N452, N448, N231);
xor XOR2 (N453, N431, N311);
nand NAND4 (N454, N453, N11, N158, N336);
nor NOR3 (N455, N449, N325, N413);
not NOT1 (N456, N454);
buf BUF1 (N457, N451);
not NOT1 (N458, N435);
buf BUF1 (N459, N446);
xor XOR2 (N460, N457, N260);
and AND3 (N461, N430, N85, N27);
nor NOR4 (N462, N461, N217, N135, N329);
not NOT1 (N463, N452);
and AND3 (N464, N459, N23, N273);
not NOT1 (N465, N450);
and AND4 (N466, N464, N359, N249, N251);
and AND4 (N467, N456, N335, N374, N219);
not NOT1 (N468, N467);
xor XOR2 (N469, N433, N92);
not NOT1 (N470, N460);
not NOT1 (N471, N470);
and AND4 (N472, N463, N37, N329, N147);
nand NAND3 (N473, N444, N82, N341);
or OR3 (N474, N469, N434, N120);
buf BUF1 (N475, N473);
buf BUF1 (N476, N468);
xor XOR2 (N477, N462, N53);
nand NAND3 (N478, N472, N262, N136);
and AND3 (N479, N477, N349, N375);
not NOT1 (N480, N476);
xor XOR2 (N481, N465, N470);
or OR2 (N482, N474, N78);
nor NOR3 (N483, N455, N333, N196);
and AND2 (N484, N482, N39);
not NOT1 (N485, N458);
buf BUF1 (N486, N485);
nor NOR2 (N487, N480, N359);
xor XOR2 (N488, N479, N48);
not NOT1 (N489, N481);
xor XOR2 (N490, N489, N141);
buf BUF1 (N491, N471);
nand NAND2 (N492, N484, N282);
and AND2 (N493, N490, N363);
nand NAND3 (N494, N486, N379, N345);
or OR4 (N495, N483, N265, N74, N268);
nand NAND2 (N496, N494, N222);
or OR3 (N497, N495, N317, N307);
buf BUF1 (N498, N488);
nand NAND2 (N499, N466, N79);
buf BUF1 (N500, N491);
nand NAND3 (N501, N497, N333, N475);
buf BUF1 (N502, N135);
buf BUF1 (N503, N496);
nor NOR4 (N504, N493, N460, N96, N172);
nor NOR3 (N505, N501, N68, N493);
not NOT1 (N506, N500);
not NOT1 (N507, N499);
nand NAND4 (N508, N504, N125, N344, N348);
buf BUF1 (N509, N502);
buf BUF1 (N510, N487);
not NOT1 (N511, N510);
and AND2 (N512, N498, N484);
and AND3 (N513, N512, N481, N286);
buf BUF1 (N514, N507);
nor NOR4 (N515, N513, N341, N492, N245);
not NOT1 (N516, N330);
or OR4 (N517, N514, N337, N372, N103);
xor XOR2 (N518, N509, N235);
nor NOR3 (N519, N508, N95, N44);
or OR3 (N520, N516, N45, N336);
and AND3 (N521, N520, N203, N32);
or OR4 (N522, N478, N521, N133, N156);
nand NAND3 (N523, N183, N324, N466);
buf BUF1 (N524, N506);
or OR2 (N525, N519, N174);
not NOT1 (N526, N503);
or OR3 (N527, N511, N34, N35);
nor NOR2 (N528, N515, N247);
buf BUF1 (N529, N522);
or OR3 (N530, N527, N272, N164);
xor XOR2 (N531, N517, N251);
nand NAND4 (N532, N529, N210, N306, N492);
not NOT1 (N533, N526);
buf BUF1 (N534, N518);
buf BUF1 (N535, N532);
nand NAND4 (N536, N533, N13, N423, N336);
nand NAND4 (N537, N534, N234, N80, N401);
nand NAND2 (N538, N530, N267);
or OR2 (N539, N525, N25);
buf BUF1 (N540, N535);
buf BUF1 (N541, N538);
not NOT1 (N542, N537);
not NOT1 (N543, N539);
nand NAND2 (N544, N536, N176);
xor XOR2 (N545, N543, N104);
or OR2 (N546, N540, N481);
or OR3 (N547, N544, N313, N334);
nor NOR4 (N548, N541, N99, N77, N371);
xor XOR2 (N549, N548, N337);
or OR4 (N550, N505, N399, N242, N485);
or OR2 (N551, N531, N428);
and AND3 (N552, N547, N332, N254);
or OR2 (N553, N528, N254);
buf BUF1 (N554, N550);
nor NOR4 (N555, N523, N107, N68, N124);
nor NOR2 (N556, N546, N155);
and AND2 (N557, N556, N332);
not NOT1 (N558, N524);
nand NAND4 (N559, N549, N245, N142, N469);
not NOT1 (N560, N551);
nor NOR4 (N561, N553, N42, N142, N353);
and AND2 (N562, N554, N484);
xor XOR2 (N563, N561, N444);
buf BUF1 (N564, N563);
and AND3 (N565, N545, N423, N4);
nand NAND3 (N566, N560, N134, N263);
or OR2 (N567, N562, N273);
buf BUF1 (N568, N552);
or OR2 (N569, N566, N279);
buf BUF1 (N570, N558);
and AND2 (N571, N564, N472);
buf BUF1 (N572, N557);
or OR2 (N573, N555, N223);
buf BUF1 (N574, N573);
buf BUF1 (N575, N565);
and AND4 (N576, N571, N568, N11, N261);
nand NAND2 (N577, N361, N8);
xor XOR2 (N578, N574, N137);
buf BUF1 (N579, N542);
not NOT1 (N580, N577);
nor NOR4 (N581, N575, N274, N533, N120);
xor XOR2 (N582, N578, N528);
nand NAND3 (N583, N581, N376, N237);
xor XOR2 (N584, N567, N273);
xor XOR2 (N585, N570, N348);
xor XOR2 (N586, N584, N499);
xor XOR2 (N587, N572, N256);
nor NOR2 (N588, N586, N585);
xor XOR2 (N589, N28, N432);
and AND4 (N590, N559, N219, N360, N263);
or OR3 (N591, N579, N554, N323);
and AND3 (N592, N580, N262, N408);
nor NOR2 (N593, N569, N154);
not NOT1 (N594, N587);
not NOT1 (N595, N591);
or OR3 (N596, N583, N92, N333);
or OR4 (N597, N588, N6, N338, N289);
xor XOR2 (N598, N592, N457);
or OR2 (N599, N593, N397);
and AND2 (N600, N590, N553);
xor XOR2 (N601, N596, N34);
xor XOR2 (N602, N595, N340);
xor XOR2 (N603, N594, N65);
buf BUF1 (N604, N582);
buf BUF1 (N605, N597);
nor NOR2 (N606, N589, N587);
nand NAND2 (N607, N602, N185);
buf BUF1 (N608, N603);
buf BUF1 (N609, N605);
xor XOR2 (N610, N604, N75);
buf BUF1 (N611, N609);
nand NAND2 (N612, N611, N374);
not NOT1 (N613, N598);
buf BUF1 (N614, N576);
buf BUF1 (N615, N607);
nor NOR3 (N616, N608, N201, N354);
not NOT1 (N617, N613);
nor NOR2 (N618, N606, N49);
buf BUF1 (N619, N615);
nand NAND2 (N620, N612, N422);
and AND2 (N621, N601, N375);
nor NOR2 (N622, N619, N284);
buf BUF1 (N623, N600);
and AND3 (N624, N610, N93, N394);
nand NAND4 (N625, N621, N385, N259, N100);
not NOT1 (N626, N625);
not NOT1 (N627, N622);
or OR3 (N628, N627, N627, N15);
buf BUF1 (N629, N618);
xor XOR2 (N630, N626, N145);
or OR4 (N631, N617, N424, N142, N276);
nand NAND3 (N632, N624, N587, N442);
not NOT1 (N633, N620);
or OR2 (N634, N628, N95);
nor NOR4 (N635, N629, N451, N150, N213);
xor XOR2 (N636, N623, N611);
nor NOR2 (N637, N631, N507);
or OR3 (N638, N632, N32, N499);
nor NOR4 (N639, N634, N145, N401, N366);
not NOT1 (N640, N630);
not NOT1 (N641, N638);
xor XOR2 (N642, N616, N400);
or OR2 (N643, N639, N372);
or OR4 (N644, N643, N164, N394, N129);
and AND3 (N645, N641, N559, N228);
nor NOR2 (N646, N635, N352);
and AND2 (N647, N645, N189);
nor NOR4 (N648, N642, N81, N337, N561);
xor XOR2 (N649, N647, N350);
not NOT1 (N650, N649);
buf BUF1 (N651, N636);
or OR3 (N652, N646, N356, N342);
nand NAND3 (N653, N637, N54, N569);
or OR2 (N654, N648, N98);
xor XOR2 (N655, N652, N551);
not NOT1 (N656, N654);
buf BUF1 (N657, N640);
xor XOR2 (N658, N657, N119);
nand NAND3 (N659, N658, N17, N321);
buf BUF1 (N660, N633);
not NOT1 (N661, N651);
nand NAND3 (N662, N655, N540, N490);
nor NOR4 (N663, N644, N210, N193, N546);
nand NAND3 (N664, N661, N293, N144);
buf BUF1 (N665, N662);
nor NOR4 (N666, N614, N61, N315, N54);
and AND2 (N667, N665, N99);
and AND4 (N668, N664, N495, N263, N486);
xor XOR2 (N669, N663, N182);
nor NOR4 (N670, N660, N409, N113, N481);
nor NOR2 (N671, N668, N436);
xor XOR2 (N672, N670, N26);
xor XOR2 (N673, N667, N266);
not NOT1 (N674, N669);
and AND4 (N675, N666, N33, N408, N37);
nor NOR4 (N676, N650, N646, N512, N15);
or OR4 (N677, N675, N122, N195, N645);
xor XOR2 (N678, N653, N33);
or OR2 (N679, N674, N636);
buf BUF1 (N680, N677);
nand NAND3 (N681, N672, N645, N47);
xor XOR2 (N682, N673, N561);
nor NOR4 (N683, N671, N241, N527, N236);
buf BUF1 (N684, N681);
not NOT1 (N685, N683);
xor XOR2 (N686, N676, N377);
or OR3 (N687, N659, N642, N176);
nor NOR3 (N688, N687, N207, N628);
buf BUF1 (N689, N599);
not NOT1 (N690, N684);
not NOT1 (N691, N689);
buf BUF1 (N692, N686);
buf BUF1 (N693, N691);
or OR4 (N694, N656, N445, N377, N410);
nand NAND3 (N695, N694, N54, N381);
buf BUF1 (N696, N682);
nor NOR4 (N697, N688, N456, N442, N101);
nand NAND3 (N698, N678, N291, N334);
nor NOR3 (N699, N685, N652, N365);
nor NOR4 (N700, N696, N619, N437, N578);
nor NOR3 (N701, N698, N73, N80);
nand NAND3 (N702, N680, N4, N385);
and AND2 (N703, N695, N698);
xor XOR2 (N704, N702, N433);
buf BUF1 (N705, N703);
or OR2 (N706, N697, N496);
nor NOR3 (N707, N693, N245, N325);
and AND4 (N708, N705, N627, N219, N216);
nand NAND4 (N709, N700, N63, N194, N73);
not NOT1 (N710, N699);
or OR4 (N711, N704, N579, N536, N466);
xor XOR2 (N712, N707, N455);
xor XOR2 (N713, N710, N563);
nand NAND2 (N714, N679, N659);
nor NOR4 (N715, N714, N539, N141, N356);
not NOT1 (N716, N712);
buf BUF1 (N717, N709);
and AND3 (N718, N701, N300, N554);
and AND3 (N719, N692, N247, N97);
not NOT1 (N720, N708);
or OR4 (N721, N716, N682, N103, N29);
buf BUF1 (N722, N706);
buf BUF1 (N723, N721);
nand NAND4 (N724, N690, N320, N212, N133);
not NOT1 (N725, N724);
not NOT1 (N726, N711);
buf BUF1 (N727, N726);
xor XOR2 (N728, N720, N167);
xor XOR2 (N729, N727, N548);
nor NOR3 (N730, N717, N104, N649);
and AND3 (N731, N713, N142, N32);
not NOT1 (N732, N718);
nand NAND3 (N733, N730, N629, N582);
nand NAND3 (N734, N725, N586, N201);
nor NOR3 (N735, N719, N41, N95);
nor NOR3 (N736, N734, N117, N316);
not NOT1 (N737, N715);
xor XOR2 (N738, N736, N612);
buf BUF1 (N739, N735);
nand NAND3 (N740, N732, N317, N647);
nor NOR4 (N741, N739, N5, N394, N652);
or OR4 (N742, N728, N400, N513, N524);
nor NOR2 (N743, N729, N224);
and AND2 (N744, N722, N13);
and AND4 (N745, N743, N239, N161, N132);
nor NOR2 (N746, N738, N523);
xor XOR2 (N747, N745, N161);
buf BUF1 (N748, N746);
buf BUF1 (N749, N733);
or OR4 (N750, N741, N592, N613, N709);
nor NOR3 (N751, N742, N344, N659);
and AND2 (N752, N744, N323);
or OR2 (N753, N748, N2);
xor XOR2 (N754, N747, N680);
and AND4 (N755, N723, N107, N177, N153);
nand NAND4 (N756, N755, N533, N383, N218);
buf BUF1 (N757, N750);
xor XOR2 (N758, N737, N646);
nand NAND3 (N759, N753, N46, N396);
buf BUF1 (N760, N754);
and AND3 (N761, N759, N555, N624);
not NOT1 (N762, N731);
buf BUF1 (N763, N756);
xor XOR2 (N764, N760, N619);
nand NAND4 (N765, N752, N10, N260, N267);
xor XOR2 (N766, N761, N439);
or OR4 (N767, N757, N626, N521, N591);
or OR4 (N768, N758, N375, N280, N382);
nand NAND4 (N769, N768, N563, N150, N739);
buf BUF1 (N770, N740);
buf BUF1 (N771, N769);
and AND2 (N772, N762, N33);
nand NAND3 (N773, N749, N535, N191);
not NOT1 (N774, N764);
or OR4 (N775, N765, N146, N360, N283);
buf BUF1 (N776, N772);
buf BUF1 (N777, N767);
buf BUF1 (N778, N777);
nor NOR3 (N779, N766, N670, N647);
nand NAND2 (N780, N775, N665);
or OR4 (N781, N774, N187, N729, N187);
not NOT1 (N782, N780);
nor NOR4 (N783, N771, N768, N118, N673);
or OR2 (N784, N776, N492);
nand NAND2 (N785, N781, N678);
or OR4 (N786, N784, N110, N302, N458);
nor NOR4 (N787, N782, N588, N678, N658);
or OR3 (N788, N783, N238, N775);
buf BUF1 (N789, N786);
xor XOR2 (N790, N773, N301);
and AND4 (N791, N785, N103, N348, N93);
not NOT1 (N792, N763);
buf BUF1 (N793, N751);
not NOT1 (N794, N779);
nor NOR3 (N795, N788, N716, N2);
nor NOR4 (N796, N792, N272, N131, N477);
xor XOR2 (N797, N794, N542);
nand NAND3 (N798, N787, N675, N549);
not NOT1 (N799, N770);
xor XOR2 (N800, N799, N432);
not NOT1 (N801, N791);
buf BUF1 (N802, N790);
not NOT1 (N803, N795);
and AND4 (N804, N789, N436, N759, N732);
nor NOR3 (N805, N803, N607, N628);
and AND3 (N806, N800, N18, N53);
and AND4 (N807, N796, N64, N56, N74);
or OR2 (N808, N806, N647);
nand NAND4 (N809, N808, N688, N21, N548);
not NOT1 (N810, N805);
not NOT1 (N811, N797);
and AND2 (N812, N807, N666);
or OR3 (N813, N778, N767, N462);
not NOT1 (N814, N801);
buf BUF1 (N815, N812);
nand NAND3 (N816, N802, N793, N135);
or OR2 (N817, N629, N459);
not NOT1 (N818, N815);
and AND4 (N819, N813, N426, N116, N163);
buf BUF1 (N820, N798);
nor NOR3 (N821, N804, N104, N784);
or OR4 (N822, N811, N582, N414, N639);
or OR3 (N823, N817, N397, N209);
buf BUF1 (N824, N809);
nor NOR3 (N825, N818, N294, N58);
nor NOR3 (N826, N814, N793, N177);
buf BUF1 (N827, N825);
xor XOR2 (N828, N821, N214);
xor XOR2 (N829, N826, N179);
nor NOR4 (N830, N820, N105, N448, N644);
nand NAND3 (N831, N824, N117, N645);
xor XOR2 (N832, N829, N72);
nand NAND2 (N833, N819, N665);
buf BUF1 (N834, N810);
not NOT1 (N835, N831);
not NOT1 (N836, N827);
nor NOR4 (N837, N835, N201, N202, N763);
nand NAND4 (N838, N834, N75, N86, N611);
not NOT1 (N839, N833);
and AND2 (N840, N837, N538);
xor XOR2 (N841, N830, N528);
and AND3 (N842, N841, N389, N578);
nor NOR2 (N843, N816, N293);
buf BUF1 (N844, N822);
nand NAND2 (N845, N832, N782);
buf BUF1 (N846, N836);
or OR2 (N847, N839, N20);
nor NOR4 (N848, N842, N616, N225, N47);
xor XOR2 (N849, N847, N629);
and AND4 (N850, N845, N230, N157, N706);
or OR3 (N851, N846, N78, N305);
buf BUF1 (N852, N851);
not NOT1 (N853, N848);
and AND2 (N854, N853, N75);
not NOT1 (N855, N850);
or OR4 (N856, N828, N333, N493, N490);
or OR2 (N857, N852, N88);
nand NAND3 (N858, N855, N697, N648);
not NOT1 (N859, N840);
nor NOR3 (N860, N823, N41, N493);
not NOT1 (N861, N857);
nand NAND3 (N862, N859, N295, N476);
buf BUF1 (N863, N854);
not NOT1 (N864, N860);
xor XOR2 (N865, N861, N629);
or OR2 (N866, N843, N12);
buf BUF1 (N867, N844);
or OR3 (N868, N856, N36, N836);
nor NOR2 (N869, N849, N485);
not NOT1 (N870, N858);
nand NAND2 (N871, N865, N91);
and AND2 (N872, N866, N7);
or OR4 (N873, N838, N218, N572, N12);
nor NOR4 (N874, N868, N465, N394, N613);
xor XOR2 (N875, N869, N477);
not NOT1 (N876, N871);
or OR3 (N877, N874, N555, N448);
nand NAND3 (N878, N875, N773, N795);
nor NOR4 (N879, N872, N594, N876, N582);
not NOT1 (N880, N821);
buf BUF1 (N881, N873);
not NOT1 (N882, N878);
or OR3 (N883, N877, N507, N866);
nor NOR3 (N884, N864, N177, N859);
or OR4 (N885, N870, N406, N774, N205);
and AND3 (N886, N881, N512, N858);
and AND2 (N887, N886, N511);
not NOT1 (N888, N880);
nor NOR4 (N889, N884, N373, N813, N645);
nor NOR2 (N890, N885, N492);
nand NAND4 (N891, N889, N35, N837, N81);
nor NOR4 (N892, N867, N82, N868, N146);
xor XOR2 (N893, N890, N854);
buf BUF1 (N894, N883);
and AND4 (N895, N891, N566, N794, N138);
nand NAND2 (N896, N879, N88);
nor NOR4 (N897, N896, N413, N337, N103);
buf BUF1 (N898, N893);
or OR4 (N899, N862, N136, N708, N345);
nor NOR3 (N900, N895, N897, N878);
not NOT1 (N901, N666);
not NOT1 (N902, N901);
not NOT1 (N903, N894);
not NOT1 (N904, N899);
xor XOR2 (N905, N863, N189);
not NOT1 (N906, N882);
xor XOR2 (N907, N888, N132);
not NOT1 (N908, N906);
buf BUF1 (N909, N904);
not NOT1 (N910, N908);
xor XOR2 (N911, N900, N27);
nor NOR4 (N912, N898, N364, N834, N848);
nor NOR4 (N913, N903, N559, N873, N833);
or OR3 (N914, N905, N735, N723);
xor XOR2 (N915, N909, N95);
nor NOR2 (N916, N907, N324);
nand NAND3 (N917, N914, N903, N51);
nand NAND3 (N918, N902, N390, N903);
nor NOR3 (N919, N887, N708, N355);
xor XOR2 (N920, N913, N158);
or OR2 (N921, N918, N756);
or OR2 (N922, N915, N338);
nand NAND4 (N923, N920, N167, N6, N306);
and AND4 (N924, N921, N139, N613, N678);
buf BUF1 (N925, N911);
buf BUF1 (N926, N922);
buf BUF1 (N927, N919);
nor NOR4 (N928, N916, N795, N652, N840);
xor XOR2 (N929, N892, N836);
buf BUF1 (N930, N926);
nor NOR2 (N931, N923, N766);
nor NOR2 (N932, N930, N713);
xor XOR2 (N933, N929, N842);
and AND3 (N934, N932, N901, N368);
xor XOR2 (N935, N925, N798);
nand NAND2 (N936, N933, N136);
buf BUF1 (N937, N910);
and AND2 (N938, N936, N303);
nand NAND4 (N939, N931, N379, N466, N555);
nor NOR4 (N940, N938, N431, N204, N201);
not NOT1 (N941, N917);
nor NOR2 (N942, N928, N372);
or OR3 (N943, N940, N520, N358);
nor NOR3 (N944, N939, N57, N14);
buf BUF1 (N945, N943);
nand NAND2 (N946, N924, N515);
xor XOR2 (N947, N942, N43);
not NOT1 (N948, N946);
not NOT1 (N949, N947);
buf BUF1 (N950, N934);
not NOT1 (N951, N950);
buf BUF1 (N952, N937);
not NOT1 (N953, N952);
or OR2 (N954, N945, N94);
and AND4 (N955, N927, N536, N329, N936);
nor NOR3 (N956, N954, N934, N715);
nand NAND4 (N957, N951, N62, N205, N747);
not NOT1 (N958, N949);
nand NAND2 (N959, N957, N579);
not NOT1 (N960, N941);
nand NAND2 (N961, N956, N894);
or OR3 (N962, N958, N146, N382);
or OR4 (N963, N944, N744, N501, N623);
and AND3 (N964, N962, N334, N895);
xor XOR2 (N965, N935, N380);
or OR4 (N966, N960, N885, N168, N203);
buf BUF1 (N967, N963);
buf BUF1 (N968, N964);
or OR4 (N969, N967, N169, N810, N268);
not NOT1 (N970, N966);
xor XOR2 (N971, N912, N174);
not NOT1 (N972, N969);
nand NAND2 (N973, N961, N845);
and AND2 (N974, N970, N874);
buf BUF1 (N975, N973);
xor XOR2 (N976, N959, N889);
nand NAND4 (N977, N965, N964, N96, N344);
and AND4 (N978, N971, N301, N534, N779);
nor NOR3 (N979, N968, N537, N192);
xor XOR2 (N980, N978, N595);
not NOT1 (N981, N955);
or OR3 (N982, N977, N548, N619);
or OR3 (N983, N976, N597, N385);
or OR2 (N984, N983, N720);
xor XOR2 (N985, N979, N719);
or OR3 (N986, N985, N864, N789);
nand NAND3 (N987, N975, N701, N866);
not NOT1 (N988, N984);
not NOT1 (N989, N972);
or OR4 (N990, N974, N707, N948, N817);
nand NAND2 (N991, N518, N532);
not NOT1 (N992, N990);
not NOT1 (N993, N953);
nor NOR2 (N994, N988, N842);
nor NOR4 (N995, N991, N708, N567, N60);
nor NOR4 (N996, N987, N876, N698, N985);
not NOT1 (N997, N995);
not NOT1 (N998, N992);
not NOT1 (N999, N980);
buf BUF1 (N1000, N994);
and AND3 (N1001, N981, N826, N476);
xor XOR2 (N1002, N1000, N388);
nand NAND4 (N1003, N1002, N822, N462, N768);
not NOT1 (N1004, N997);
nand NAND2 (N1005, N989, N434);
xor XOR2 (N1006, N1003, N699);
xor XOR2 (N1007, N996, N234);
buf BUF1 (N1008, N993);
xor XOR2 (N1009, N986, N670);
and AND4 (N1010, N998, N6, N460, N772);
or OR3 (N1011, N1007, N395, N357);
buf BUF1 (N1012, N1001);
nand NAND4 (N1013, N1005, N319, N791, N623);
and AND3 (N1014, N1004, N742, N916);
nand NAND2 (N1015, N1011, N646);
buf BUF1 (N1016, N1013);
and AND2 (N1017, N1008, N355);
nand NAND4 (N1018, N1012, N752, N995, N383);
and AND4 (N1019, N999, N174, N840, N291);
xor XOR2 (N1020, N982, N757);
xor XOR2 (N1021, N1017, N810);
nor NOR3 (N1022, N1010, N64, N99);
or OR3 (N1023, N1021, N821, N901);
or OR2 (N1024, N1020, N144);
buf BUF1 (N1025, N1019);
not NOT1 (N1026, N1016);
xor XOR2 (N1027, N1026, N715);
xor XOR2 (N1028, N1018, N881);
nand NAND4 (N1029, N1015, N133, N142, N634);
not NOT1 (N1030, N1023);
nand NAND4 (N1031, N1014, N843, N118, N818);
buf BUF1 (N1032, N1028);
nand NAND4 (N1033, N1006, N727, N351, N591);
xor XOR2 (N1034, N1009, N676);
nand NAND2 (N1035, N1030, N543);
or OR4 (N1036, N1032, N250, N697, N850);
nand NAND2 (N1037, N1034, N28);
not NOT1 (N1038, N1031);
xor XOR2 (N1039, N1027, N282);
buf BUF1 (N1040, N1038);
or OR3 (N1041, N1036, N491, N329);
nand NAND4 (N1042, N1040, N799, N504, N491);
nor NOR2 (N1043, N1037, N872);
or OR2 (N1044, N1033, N1012);
or OR2 (N1045, N1022, N969);
or OR2 (N1046, N1042, N1037);
xor XOR2 (N1047, N1029, N741);
and AND2 (N1048, N1045, N767);
xor XOR2 (N1049, N1035, N73);
xor XOR2 (N1050, N1048, N242);
buf BUF1 (N1051, N1046);
nor NOR2 (N1052, N1051, N574);
xor XOR2 (N1053, N1024, N415);
buf BUF1 (N1054, N1052);
buf BUF1 (N1055, N1041);
not NOT1 (N1056, N1044);
nor NOR4 (N1057, N1055, N114, N557, N330);
and AND4 (N1058, N1039, N507, N892, N577);
nand NAND4 (N1059, N1054, N85, N309, N385);
xor XOR2 (N1060, N1058, N861);
nand NAND2 (N1061, N1025, N251);
or OR2 (N1062, N1056, N1037);
not NOT1 (N1063, N1050);
nand NAND3 (N1064, N1049, N1052, N213);
xor XOR2 (N1065, N1059, N207);
nand NAND3 (N1066, N1063, N592, N622);
and AND2 (N1067, N1053, N484);
not NOT1 (N1068, N1064);
xor XOR2 (N1069, N1065, N601);
or OR3 (N1070, N1067, N363, N788);
xor XOR2 (N1071, N1069, N806);
or OR2 (N1072, N1068, N140);
nor NOR4 (N1073, N1043, N1017, N85, N21);
xor XOR2 (N1074, N1057, N472);
or OR2 (N1075, N1074, N724);
buf BUF1 (N1076, N1061);
not NOT1 (N1077, N1062);
not NOT1 (N1078, N1066);
nor NOR4 (N1079, N1070, N594, N606, N875);
buf BUF1 (N1080, N1072);
nand NAND4 (N1081, N1047, N15, N567, N52);
and AND3 (N1082, N1081, N733, N1035);
nor NOR3 (N1083, N1077, N929, N710);
nand NAND2 (N1084, N1078, N11);
nand NAND4 (N1085, N1071, N1016, N1045, N501);
nand NAND4 (N1086, N1075, N905, N903, N303);
not NOT1 (N1087, N1080);
and AND4 (N1088, N1073, N447, N576, N1048);
xor XOR2 (N1089, N1085, N1044);
buf BUF1 (N1090, N1086);
and AND3 (N1091, N1083, N367, N615);
and AND2 (N1092, N1089, N577);
nand NAND2 (N1093, N1079, N978);
buf BUF1 (N1094, N1076);
xor XOR2 (N1095, N1094, N335);
nand NAND2 (N1096, N1093, N683);
or OR3 (N1097, N1088, N827, N1034);
nand NAND3 (N1098, N1087, N586, N434);
xor XOR2 (N1099, N1096, N539);
and AND2 (N1100, N1098, N347);
buf BUF1 (N1101, N1082);
not NOT1 (N1102, N1060);
or OR3 (N1103, N1101, N909, N626);
buf BUF1 (N1104, N1102);
xor XOR2 (N1105, N1084, N324);
buf BUF1 (N1106, N1105);
not NOT1 (N1107, N1100);
and AND2 (N1108, N1090, N740);
or OR4 (N1109, N1103, N55, N418, N870);
xor XOR2 (N1110, N1107, N430);
xor XOR2 (N1111, N1106, N881);
nand NAND4 (N1112, N1097, N700, N818, N253);
buf BUF1 (N1113, N1104);
nand NAND2 (N1114, N1092, N648);
or OR2 (N1115, N1095, N325);
xor XOR2 (N1116, N1111, N862);
and AND3 (N1117, N1116, N859, N765);
xor XOR2 (N1118, N1115, N378);
not NOT1 (N1119, N1108);
xor XOR2 (N1120, N1119, N1084);
xor XOR2 (N1121, N1109, N615);
xor XOR2 (N1122, N1112, N1042);
or OR3 (N1123, N1099, N388, N172);
xor XOR2 (N1124, N1110, N334);
buf BUF1 (N1125, N1113);
not NOT1 (N1126, N1117);
buf BUF1 (N1127, N1091);
buf BUF1 (N1128, N1124);
xor XOR2 (N1129, N1121, N89);
not NOT1 (N1130, N1129);
buf BUF1 (N1131, N1120);
nand NAND3 (N1132, N1122, N1039, N553);
buf BUF1 (N1133, N1130);
buf BUF1 (N1134, N1132);
nor NOR3 (N1135, N1118, N1015, N767);
or OR4 (N1136, N1127, N765, N499, N811);
nor NOR4 (N1137, N1126, N1095, N832, N1060);
nand NAND2 (N1138, N1131, N743);
or OR3 (N1139, N1136, N249, N135);
nor NOR3 (N1140, N1134, N673, N939);
nand NAND2 (N1141, N1125, N524);
or OR3 (N1142, N1141, N274, N864);
or OR2 (N1143, N1142, N36);
nand NAND4 (N1144, N1143, N1060, N138, N1058);
buf BUF1 (N1145, N1138);
xor XOR2 (N1146, N1140, N562);
nand NAND2 (N1147, N1137, N581);
not NOT1 (N1148, N1135);
or OR3 (N1149, N1133, N854, N86);
xor XOR2 (N1150, N1149, N541);
nor NOR4 (N1151, N1150, N24, N354, N167);
and AND3 (N1152, N1148, N178, N525);
nor NOR2 (N1153, N1145, N667);
nand NAND3 (N1154, N1153, N867, N731);
buf BUF1 (N1155, N1139);
buf BUF1 (N1156, N1154);
or OR3 (N1157, N1156, N327, N77);
xor XOR2 (N1158, N1144, N1110);
buf BUF1 (N1159, N1123);
and AND3 (N1160, N1146, N810, N1020);
xor XOR2 (N1161, N1147, N563);
xor XOR2 (N1162, N1159, N321);
nand NAND3 (N1163, N1155, N1041, N1115);
buf BUF1 (N1164, N1162);
buf BUF1 (N1165, N1164);
buf BUF1 (N1166, N1114);
not NOT1 (N1167, N1166);
nor NOR4 (N1168, N1161, N469, N550, N320);
or OR4 (N1169, N1157, N434, N149, N723);
not NOT1 (N1170, N1167);
not NOT1 (N1171, N1169);
and AND4 (N1172, N1168, N240, N574, N135);
nor NOR4 (N1173, N1163, N266, N876, N513);
nor NOR2 (N1174, N1160, N193);
and AND4 (N1175, N1165, N715, N835, N434);
nand NAND2 (N1176, N1128, N525);
buf BUF1 (N1177, N1151);
nand NAND4 (N1178, N1152, N506, N619, N1120);
buf BUF1 (N1179, N1178);
xor XOR2 (N1180, N1179, N364);
or OR3 (N1181, N1175, N51, N1132);
nor NOR4 (N1182, N1158, N426, N788, N138);
nand NAND3 (N1183, N1182, N888, N878);
and AND3 (N1184, N1181, N357, N550);
nand NAND2 (N1185, N1180, N10);
nand NAND4 (N1186, N1183, N4, N20, N431);
nand NAND2 (N1187, N1185, N427);
and AND2 (N1188, N1184, N649);
buf BUF1 (N1189, N1176);
or OR3 (N1190, N1170, N811, N142);
or OR3 (N1191, N1172, N509, N480);
nand NAND3 (N1192, N1174, N13, N179);
buf BUF1 (N1193, N1187);
nand NAND2 (N1194, N1192, N257);
xor XOR2 (N1195, N1191, N203);
not NOT1 (N1196, N1189);
nor NOR3 (N1197, N1177, N548, N895);
xor XOR2 (N1198, N1186, N741);
not NOT1 (N1199, N1197);
nand NAND4 (N1200, N1196, N705, N387, N651);
buf BUF1 (N1201, N1195);
and AND3 (N1202, N1198, N626, N80);
nand NAND2 (N1203, N1200, N114);
xor XOR2 (N1204, N1193, N636);
and AND2 (N1205, N1199, N326);
and AND2 (N1206, N1205, N517);
nand NAND2 (N1207, N1173, N315);
nand NAND4 (N1208, N1188, N598, N4, N415);
or OR2 (N1209, N1171, N51);
nor NOR4 (N1210, N1207, N597, N940, N386);
nand NAND4 (N1211, N1194, N1054, N210, N307);
buf BUF1 (N1212, N1204);
xor XOR2 (N1213, N1208, N986);
nand NAND3 (N1214, N1211, N702, N204);
not NOT1 (N1215, N1203);
nor NOR2 (N1216, N1190, N795);
xor XOR2 (N1217, N1212, N197);
nor NOR4 (N1218, N1215, N371, N1071, N43);
and AND3 (N1219, N1210, N889, N89);
xor XOR2 (N1220, N1206, N1142);
not NOT1 (N1221, N1217);
nor NOR4 (N1222, N1201, N642, N1038, N47);
nand NAND2 (N1223, N1221, N409);
nand NAND2 (N1224, N1216, N419);
xor XOR2 (N1225, N1222, N56);
xor XOR2 (N1226, N1220, N12);
or OR4 (N1227, N1209, N266, N31, N531);
xor XOR2 (N1228, N1225, N616);
buf BUF1 (N1229, N1213);
buf BUF1 (N1230, N1223);
and AND3 (N1231, N1218, N1114, N647);
xor XOR2 (N1232, N1227, N38);
buf BUF1 (N1233, N1228);
xor XOR2 (N1234, N1231, N511);
or OR3 (N1235, N1230, N822, N790);
nor NOR3 (N1236, N1234, N1126, N659);
and AND4 (N1237, N1214, N564, N267, N3);
and AND4 (N1238, N1232, N991, N231, N1117);
xor XOR2 (N1239, N1233, N409);
nor NOR2 (N1240, N1236, N1133);
not NOT1 (N1241, N1235);
and AND4 (N1242, N1241, N1047, N810, N911);
nor NOR3 (N1243, N1226, N439, N160);
and AND2 (N1244, N1224, N952);
xor XOR2 (N1245, N1240, N964);
and AND3 (N1246, N1202, N754, N292);
nand NAND2 (N1247, N1246, N1201);
and AND2 (N1248, N1245, N324);
or OR3 (N1249, N1247, N1016, N421);
or OR4 (N1250, N1229, N248, N165, N434);
nand NAND3 (N1251, N1250, N736, N761);
or OR2 (N1252, N1242, N437);
xor XOR2 (N1253, N1244, N2);
nor NOR2 (N1254, N1253, N775);
nor NOR4 (N1255, N1252, N138, N720, N1070);
xor XOR2 (N1256, N1238, N710);
nand NAND2 (N1257, N1248, N5);
buf BUF1 (N1258, N1239);
and AND2 (N1259, N1237, N661);
xor XOR2 (N1260, N1243, N1165);
xor XOR2 (N1261, N1254, N1227);
nor NOR3 (N1262, N1260, N817, N1105);
and AND4 (N1263, N1261, N485, N613, N1197);
xor XOR2 (N1264, N1256, N486);
nor NOR4 (N1265, N1255, N1182, N592, N1206);
not NOT1 (N1266, N1249);
and AND2 (N1267, N1258, N1100);
xor XOR2 (N1268, N1265, N1069);
nand NAND4 (N1269, N1251, N47, N221, N8);
not NOT1 (N1270, N1259);
nand NAND2 (N1271, N1257, N616);
or OR3 (N1272, N1268, N306, N632);
nor NOR2 (N1273, N1271, N290);
nand NAND2 (N1274, N1219, N179);
buf BUF1 (N1275, N1273);
or OR2 (N1276, N1263, N328);
or OR4 (N1277, N1274, N1006, N274, N136);
xor XOR2 (N1278, N1272, N905);
and AND3 (N1279, N1276, N1252, N1229);
or OR4 (N1280, N1267, N1040, N811, N340);
xor XOR2 (N1281, N1270, N62);
not NOT1 (N1282, N1278);
xor XOR2 (N1283, N1280, N218);
xor XOR2 (N1284, N1277, N420);
xor XOR2 (N1285, N1281, N135);
not NOT1 (N1286, N1262);
buf BUF1 (N1287, N1283);
nor NOR4 (N1288, N1269, N981, N756, N11);
or OR3 (N1289, N1266, N1235, N207);
nor NOR3 (N1290, N1286, N453, N835);
xor XOR2 (N1291, N1275, N264);
nor NOR2 (N1292, N1282, N5);
xor XOR2 (N1293, N1289, N114);
not NOT1 (N1294, N1290);
not NOT1 (N1295, N1293);
nor NOR3 (N1296, N1284, N344, N142);
or OR4 (N1297, N1292, N211, N643, N752);
and AND3 (N1298, N1295, N709, N892);
xor XOR2 (N1299, N1296, N752);
not NOT1 (N1300, N1299);
buf BUF1 (N1301, N1300);
and AND2 (N1302, N1279, N824);
not NOT1 (N1303, N1285);
not NOT1 (N1304, N1298);
not NOT1 (N1305, N1288);
nand NAND3 (N1306, N1291, N603, N857);
nor NOR2 (N1307, N1294, N32);
buf BUF1 (N1308, N1297);
and AND3 (N1309, N1305, N1191, N669);
xor XOR2 (N1310, N1302, N193);
nand NAND2 (N1311, N1303, N979);
not NOT1 (N1312, N1287);
or OR2 (N1313, N1311, N1217);
and AND4 (N1314, N1304, N840, N244, N1128);
and AND4 (N1315, N1309, N504, N239, N498);
nand NAND2 (N1316, N1307, N49);
and AND3 (N1317, N1316, N1192, N14);
and AND3 (N1318, N1264, N928, N133);
and AND3 (N1319, N1318, N44, N504);
buf BUF1 (N1320, N1306);
not NOT1 (N1321, N1308);
nor NOR4 (N1322, N1312, N1217, N571, N1247);
nor NOR2 (N1323, N1301, N823);
not NOT1 (N1324, N1313);
or OR2 (N1325, N1317, N838);
not NOT1 (N1326, N1315);
nand NAND3 (N1327, N1319, N338, N578);
or OR3 (N1328, N1322, N27, N698);
nand NAND4 (N1329, N1321, N120, N1179, N147);
buf BUF1 (N1330, N1320);
buf BUF1 (N1331, N1330);
nor NOR4 (N1332, N1329, N956, N961, N875);
not NOT1 (N1333, N1323);
or OR4 (N1334, N1310, N739, N621, N1277);
and AND3 (N1335, N1332, N346, N765);
and AND4 (N1336, N1325, N1282, N718, N272);
and AND3 (N1337, N1324, N298, N314);
nand NAND4 (N1338, N1331, N971, N1256, N426);
nand NAND3 (N1339, N1334, N1289, N1229);
or OR4 (N1340, N1314, N889, N869, N1002);
and AND4 (N1341, N1336, N787, N804, N683);
nand NAND4 (N1342, N1339, N879, N326, N1316);
nand NAND2 (N1343, N1327, N902);
buf BUF1 (N1344, N1342);
buf BUF1 (N1345, N1333);
xor XOR2 (N1346, N1344, N1042);
nor NOR4 (N1347, N1328, N1185, N575, N791);
and AND3 (N1348, N1347, N847, N142);
nor NOR3 (N1349, N1340, N570, N100);
and AND4 (N1350, N1337, N501, N1063, N596);
and AND2 (N1351, N1341, N869);
not NOT1 (N1352, N1349);
or OR3 (N1353, N1335, N995, N485);
and AND3 (N1354, N1345, N620, N328);
nor NOR4 (N1355, N1343, N403, N254, N858);
not NOT1 (N1356, N1348);
nand NAND4 (N1357, N1354, N1169, N653, N536);
not NOT1 (N1358, N1338);
nor NOR2 (N1359, N1352, N89);
buf BUF1 (N1360, N1357);
not NOT1 (N1361, N1326);
nor NOR3 (N1362, N1361, N476, N375);
buf BUF1 (N1363, N1346);
and AND3 (N1364, N1363, N629, N550);
nor NOR3 (N1365, N1360, N585, N848);
and AND4 (N1366, N1365, N1237, N910, N12);
not NOT1 (N1367, N1358);
buf BUF1 (N1368, N1359);
nand NAND4 (N1369, N1368, N605, N1269, N1217);
and AND4 (N1370, N1355, N818, N1184, N59);
nand NAND4 (N1371, N1362, N860, N1131, N260);
not NOT1 (N1372, N1369);
nor NOR3 (N1373, N1353, N539, N755);
or OR2 (N1374, N1356, N846);
and AND3 (N1375, N1370, N1337, N333);
nand NAND3 (N1376, N1364, N122, N91);
nor NOR3 (N1377, N1367, N500, N943);
buf BUF1 (N1378, N1350);
nor NOR4 (N1379, N1378, N1225, N837, N120);
buf BUF1 (N1380, N1373);
buf BUF1 (N1381, N1375);
nand NAND2 (N1382, N1351, N1269);
nand NAND4 (N1383, N1372, N778, N1131, N1349);
not NOT1 (N1384, N1371);
or OR4 (N1385, N1377, N182, N1357, N164);
xor XOR2 (N1386, N1366, N1286);
nand NAND2 (N1387, N1380, N1125);
or OR4 (N1388, N1381, N848, N713, N279);
buf BUF1 (N1389, N1388);
nor NOR4 (N1390, N1382, N1047, N964, N280);
nand NAND3 (N1391, N1384, N990, N567);
not NOT1 (N1392, N1390);
nor NOR4 (N1393, N1389, N316, N22, N817);
not NOT1 (N1394, N1392);
nand NAND4 (N1395, N1374, N868, N28, N563);
xor XOR2 (N1396, N1385, N44);
nor NOR3 (N1397, N1387, N404, N503);
not NOT1 (N1398, N1394);
buf BUF1 (N1399, N1395);
not NOT1 (N1400, N1379);
buf BUF1 (N1401, N1386);
xor XOR2 (N1402, N1401, N334);
xor XOR2 (N1403, N1391, N611);
not NOT1 (N1404, N1397);
or OR4 (N1405, N1393, N148, N412, N459);
nor NOR4 (N1406, N1398, N511, N28, N1380);
or OR4 (N1407, N1383, N766, N1253, N86);
nand NAND4 (N1408, N1405, N201, N615, N790);
xor XOR2 (N1409, N1376, N930);
buf BUF1 (N1410, N1406);
and AND4 (N1411, N1407, N468, N1047, N900);
xor XOR2 (N1412, N1411, N100);
xor XOR2 (N1413, N1410, N680);
nand NAND3 (N1414, N1396, N1297, N317);
nand NAND2 (N1415, N1412, N630);
or OR3 (N1416, N1409, N979, N1273);
or OR2 (N1417, N1402, N89);
nor NOR3 (N1418, N1408, N505, N254);
nor NOR2 (N1419, N1416, N856);
buf BUF1 (N1420, N1404);
or OR2 (N1421, N1419, N1336);
xor XOR2 (N1422, N1420, N846);
not NOT1 (N1423, N1413);
buf BUF1 (N1424, N1421);
xor XOR2 (N1425, N1423, N238);
xor XOR2 (N1426, N1399, N790);
or OR3 (N1427, N1422, N185, N260);
or OR4 (N1428, N1424, N873, N393, N705);
and AND2 (N1429, N1428, N960);
nand NAND4 (N1430, N1427, N1276, N1333, N967);
buf BUF1 (N1431, N1418);
and AND3 (N1432, N1426, N977, N348);
xor XOR2 (N1433, N1403, N343);
buf BUF1 (N1434, N1433);
xor XOR2 (N1435, N1432, N469);
xor XOR2 (N1436, N1430, N880);
buf BUF1 (N1437, N1434);
buf BUF1 (N1438, N1429);
or OR3 (N1439, N1400, N119, N715);
nor NOR2 (N1440, N1437, N1285);
not NOT1 (N1441, N1435);
nor NOR3 (N1442, N1439, N899, N619);
or OR3 (N1443, N1414, N881, N395);
buf BUF1 (N1444, N1431);
and AND2 (N1445, N1440, N1042);
not NOT1 (N1446, N1442);
or OR2 (N1447, N1441, N218);
nor NOR3 (N1448, N1438, N870, N565);
or OR4 (N1449, N1446, N1356, N39, N922);
nor NOR4 (N1450, N1449, N706, N1275, N1210);
and AND3 (N1451, N1450, N543, N990);
and AND3 (N1452, N1425, N850, N1016);
and AND2 (N1453, N1443, N1025);
buf BUF1 (N1454, N1445);
buf BUF1 (N1455, N1415);
not NOT1 (N1456, N1452);
or OR2 (N1457, N1455, N1091);
buf BUF1 (N1458, N1451);
nand NAND2 (N1459, N1448, N803);
or OR3 (N1460, N1459, N1171, N841);
not NOT1 (N1461, N1460);
or OR3 (N1462, N1444, N265, N1008);
not NOT1 (N1463, N1454);
nand NAND4 (N1464, N1417, N653, N1129, N303);
nor NOR3 (N1465, N1453, N469, N907);
nand NAND4 (N1466, N1463, N1302, N281, N630);
and AND2 (N1467, N1465, N478);
buf BUF1 (N1468, N1456);
buf BUF1 (N1469, N1462);
buf BUF1 (N1470, N1447);
nor NOR3 (N1471, N1466, N194, N395);
xor XOR2 (N1472, N1469, N869);
xor XOR2 (N1473, N1472, N1357);
or OR4 (N1474, N1461, N902, N1186, N1233);
and AND4 (N1475, N1468, N1119, N622, N1032);
nand NAND2 (N1476, N1471, N788);
or OR2 (N1477, N1467, N1293);
buf BUF1 (N1478, N1436);
or OR3 (N1479, N1475, N488, N320);
nor NOR2 (N1480, N1470, N541);
and AND2 (N1481, N1478, N1219);
and AND2 (N1482, N1458, N921);
buf BUF1 (N1483, N1464);
nor NOR2 (N1484, N1473, N697);
buf BUF1 (N1485, N1479);
not NOT1 (N1486, N1482);
buf BUF1 (N1487, N1484);
xor XOR2 (N1488, N1474, N1345);
buf BUF1 (N1489, N1476);
buf BUF1 (N1490, N1481);
not NOT1 (N1491, N1480);
not NOT1 (N1492, N1489);
and AND3 (N1493, N1487, N116, N89);
xor XOR2 (N1494, N1485, N371);
xor XOR2 (N1495, N1486, N902);
xor XOR2 (N1496, N1483, N455);
and AND4 (N1497, N1493, N235, N1275, N877);
nor NOR2 (N1498, N1477, N444);
not NOT1 (N1499, N1490);
not NOT1 (N1500, N1498);
and AND2 (N1501, N1457, N269);
and AND4 (N1502, N1500, N1397, N325, N725);
or OR4 (N1503, N1497, N1190, N986, N783);
nand NAND2 (N1504, N1503, N1052);
buf BUF1 (N1505, N1491);
or OR3 (N1506, N1494, N683, N1405);
not NOT1 (N1507, N1499);
xor XOR2 (N1508, N1496, N648);
and AND2 (N1509, N1492, N1000);
buf BUF1 (N1510, N1488);
and AND2 (N1511, N1508, N185);
xor XOR2 (N1512, N1502, N1262);
xor XOR2 (N1513, N1512, N1449);
buf BUF1 (N1514, N1501);
nor NOR4 (N1515, N1506, N698, N1508, N284);
and AND2 (N1516, N1509, N688);
buf BUF1 (N1517, N1510);
buf BUF1 (N1518, N1504);
nand NAND2 (N1519, N1505, N240);
or OR4 (N1520, N1513, N743, N124, N356);
nor NOR4 (N1521, N1515, N1477, N482, N291);
nor NOR3 (N1522, N1507, N810, N1515);
nor NOR2 (N1523, N1517, N1207);
xor XOR2 (N1524, N1516, N89);
nand NAND2 (N1525, N1495, N138);
xor XOR2 (N1526, N1518, N498);
and AND3 (N1527, N1522, N433, N142);
xor XOR2 (N1528, N1520, N999);
nor NOR4 (N1529, N1525, N130, N417, N1399);
nand NAND3 (N1530, N1521, N845, N1065);
and AND2 (N1531, N1527, N31);
buf BUF1 (N1532, N1511);
nor NOR3 (N1533, N1519, N1093, N721);
and AND3 (N1534, N1524, N1505, N1244);
nor NOR2 (N1535, N1532, N1428);
or OR3 (N1536, N1526, N237, N13);
buf BUF1 (N1537, N1535);
not NOT1 (N1538, N1533);
buf BUF1 (N1539, N1530);
or OR2 (N1540, N1534, N918);
nor NOR3 (N1541, N1537, N61, N720);
nand NAND3 (N1542, N1529, N450, N1066);
buf BUF1 (N1543, N1536);
buf BUF1 (N1544, N1528);
xor XOR2 (N1545, N1538, N950);
and AND3 (N1546, N1545, N1159, N104);
buf BUF1 (N1547, N1540);
xor XOR2 (N1548, N1543, N69);
xor XOR2 (N1549, N1539, N1489);
and AND4 (N1550, N1549, N745, N655, N1262);
not NOT1 (N1551, N1547);
not NOT1 (N1552, N1542);
or OR4 (N1553, N1551, N361, N583, N718);
and AND3 (N1554, N1523, N682, N1537);
buf BUF1 (N1555, N1541);
nor NOR3 (N1556, N1550, N410, N1371);
buf BUF1 (N1557, N1514);
not NOT1 (N1558, N1548);
xor XOR2 (N1559, N1553, N1165);
and AND4 (N1560, N1558, N1495, N802, N721);
buf BUF1 (N1561, N1546);
nand NAND2 (N1562, N1552, N606);
nand NAND4 (N1563, N1531, N548, N835, N307);
nor NOR4 (N1564, N1544, N895, N356, N1198);
or OR2 (N1565, N1562, N343);
and AND2 (N1566, N1565, N662);
xor XOR2 (N1567, N1559, N764);
nor NOR3 (N1568, N1560, N91, N165);
nand NAND3 (N1569, N1563, N1327, N505);
nand NAND2 (N1570, N1564, N1313);
xor XOR2 (N1571, N1568, N1006);
and AND4 (N1572, N1554, N375, N1211, N788);
or OR2 (N1573, N1557, N511);
nor NOR4 (N1574, N1570, N156, N252, N780);
not NOT1 (N1575, N1573);
buf BUF1 (N1576, N1561);
and AND4 (N1577, N1574, N1292, N1536, N1565);
or OR4 (N1578, N1577, N1388, N1194, N225);
not NOT1 (N1579, N1569);
or OR2 (N1580, N1576, N12);
xor XOR2 (N1581, N1579, N1046);
xor XOR2 (N1582, N1572, N69);
buf BUF1 (N1583, N1571);
or OR4 (N1584, N1580, N1040, N1391, N30);
and AND4 (N1585, N1578, N1050, N1196, N1399);
not NOT1 (N1586, N1566);
nor NOR3 (N1587, N1586, N808, N104);
or OR3 (N1588, N1583, N1247, N1091);
nor NOR3 (N1589, N1556, N320, N774);
and AND2 (N1590, N1588, N300);
and AND3 (N1591, N1567, N1179, N881);
or OR2 (N1592, N1582, N998);
and AND4 (N1593, N1584, N1071, N938, N525);
or OR3 (N1594, N1592, N157, N587);
and AND4 (N1595, N1590, N1159, N1567, N1174);
not NOT1 (N1596, N1589);
nand NAND3 (N1597, N1585, N1444, N846);
not NOT1 (N1598, N1587);
or OR2 (N1599, N1596, N296);
or OR4 (N1600, N1595, N387, N508, N742);
or OR2 (N1601, N1598, N1382);
buf BUF1 (N1602, N1600);
xor XOR2 (N1603, N1593, N1444);
not NOT1 (N1604, N1601);
buf BUF1 (N1605, N1602);
and AND2 (N1606, N1605, N441);
nor NOR4 (N1607, N1597, N556, N458, N72);
or OR3 (N1608, N1581, N173, N724);
xor XOR2 (N1609, N1575, N762);
buf BUF1 (N1610, N1607);
xor XOR2 (N1611, N1610, N1156);
and AND4 (N1612, N1603, N1010, N178, N949);
nand NAND4 (N1613, N1606, N1121, N1126, N511);
nand NAND3 (N1614, N1604, N480, N353);
nor NOR4 (N1615, N1608, N233, N792, N1606);
and AND4 (N1616, N1615, N1176, N1131, N241);
xor XOR2 (N1617, N1611, N1530);
xor XOR2 (N1618, N1614, N1547);
not NOT1 (N1619, N1591);
not NOT1 (N1620, N1619);
and AND2 (N1621, N1599, N1057);
nor NOR3 (N1622, N1616, N151, N1315);
xor XOR2 (N1623, N1613, N1486);
xor XOR2 (N1624, N1612, N1216);
nor NOR2 (N1625, N1620, N1080);
nor NOR3 (N1626, N1623, N1433, N1469);
buf BUF1 (N1627, N1594);
and AND4 (N1628, N1609, N34, N572, N190);
not NOT1 (N1629, N1625);
not NOT1 (N1630, N1626);
or OR3 (N1631, N1627, N1448, N1610);
nor NOR3 (N1632, N1631, N394, N1081);
nand NAND3 (N1633, N1624, N542, N1233);
nand NAND2 (N1634, N1622, N306);
nand NAND2 (N1635, N1618, N611);
xor XOR2 (N1636, N1632, N1599);
not NOT1 (N1637, N1635);
nand NAND3 (N1638, N1637, N1415, N826);
and AND2 (N1639, N1638, N40);
not NOT1 (N1640, N1617);
not NOT1 (N1641, N1633);
nand NAND2 (N1642, N1641, N898);
nand NAND3 (N1643, N1621, N1161, N444);
nor NOR4 (N1644, N1629, N1361, N1292, N789);
nor NOR4 (N1645, N1630, N1286, N178, N670);
nand NAND2 (N1646, N1636, N104);
not NOT1 (N1647, N1639);
xor XOR2 (N1648, N1643, N1515);
or OR3 (N1649, N1634, N1112, N1530);
not NOT1 (N1650, N1628);
xor XOR2 (N1651, N1646, N1236);
not NOT1 (N1652, N1649);
buf BUF1 (N1653, N1644);
and AND2 (N1654, N1652, N742);
not NOT1 (N1655, N1555);
or OR4 (N1656, N1648, N314, N413, N1434);
nor NOR4 (N1657, N1645, N887, N515, N1077);
nand NAND3 (N1658, N1654, N338, N828);
nand NAND4 (N1659, N1653, N1325, N239, N745);
or OR4 (N1660, N1656, N1472, N1044, N1539);
or OR4 (N1661, N1650, N532, N616, N578);
or OR4 (N1662, N1642, N691, N227, N241);
or OR2 (N1663, N1659, N1456);
or OR2 (N1664, N1640, N195);
and AND4 (N1665, N1662, N1340, N378, N948);
and AND2 (N1666, N1664, N666);
or OR2 (N1667, N1663, N1382);
buf BUF1 (N1668, N1666);
buf BUF1 (N1669, N1658);
xor XOR2 (N1670, N1657, N784);
nor NOR3 (N1671, N1665, N1036, N724);
and AND3 (N1672, N1660, N321, N620);
or OR4 (N1673, N1671, N936, N865, N748);
nand NAND3 (N1674, N1655, N1180, N1434);
nor NOR3 (N1675, N1669, N1386, N1526);
nand NAND4 (N1676, N1661, N444, N1013, N536);
or OR2 (N1677, N1651, N730);
and AND2 (N1678, N1675, N280);
xor XOR2 (N1679, N1670, N624);
nand NAND4 (N1680, N1672, N1274, N264, N1679);
nor NOR3 (N1681, N887, N1471, N1598);
buf BUF1 (N1682, N1680);
or OR2 (N1683, N1682, N632);
xor XOR2 (N1684, N1676, N1563);
nand NAND3 (N1685, N1683, N19, N1501);
or OR3 (N1686, N1667, N1452, N1378);
xor XOR2 (N1687, N1681, N672);
nor NOR3 (N1688, N1684, N1412, N1373);
xor XOR2 (N1689, N1673, N846);
nor NOR2 (N1690, N1687, N357);
or OR3 (N1691, N1674, N523, N200);
not NOT1 (N1692, N1688);
and AND3 (N1693, N1692, N103, N433);
and AND4 (N1694, N1691, N1045, N550, N1538);
buf BUF1 (N1695, N1677);
or OR4 (N1696, N1694, N1273, N1262, N921);
not NOT1 (N1697, N1668);
buf BUF1 (N1698, N1678);
xor XOR2 (N1699, N1686, N1326);
buf BUF1 (N1700, N1697);
or OR3 (N1701, N1698, N1140, N162);
buf BUF1 (N1702, N1699);
not NOT1 (N1703, N1647);
nand NAND3 (N1704, N1703, N9, N1029);
buf BUF1 (N1705, N1689);
or OR4 (N1706, N1695, N1516, N1429, N1334);
and AND3 (N1707, N1705, N1443, N1304);
xor XOR2 (N1708, N1702, N1151);
nand NAND3 (N1709, N1704, N854, N1334);
nand NAND4 (N1710, N1709, N1069, N911, N274);
buf BUF1 (N1711, N1701);
not NOT1 (N1712, N1707);
nand NAND2 (N1713, N1708, N170);
nand NAND3 (N1714, N1693, N48, N106);
xor XOR2 (N1715, N1714, N1659);
buf BUF1 (N1716, N1700);
and AND2 (N1717, N1690, N275);
or OR3 (N1718, N1713, N861, N1194);
buf BUF1 (N1719, N1717);
not NOT1 (N1720, N1718);
and AND2 (N1721, N1696, N1244);
not NOT1 (N1722, N1721);
or OR2 (N1723, N1716, N1069);
and AND2 (N1724, N1722, N763);
xor XOR2 (N1725, N1723, N497);
nand NAND2 (N1726, N1710, N1448);
or OR4 (N1727, N1720, N368, N1130, N55);
not NOT1 (N1728, N1706);
or OR2 (N1729, N1715, N546);
buf BUF1 (N1730, N1727);
nand NAND2 (N1731, N1726, N1634);
and AND4 (N1732, N1712, N13, N1334, N998);
not NOT1 (N1733, N1730);
xor XOR2 (N1734, N1685, N94);
buf BUF1 (N1735, N1711);
nand NAND3 (N1736, N1719, N670, N705);
xor XOR2 (N1737, N1734, N1164);
and AND3 (N1738, N1736, N255, N612);
buf BUF1 (N1739, N1724);
not NOT1 (N1740, N1739);
not NOT1 (N1741, N1740);
nand NAND2 (N1742, N1732, N735);
or OR4 (N1743, N1733, N205, N1120, N356);
not NOT1 (N1744, N1728);
or OR3 (N1745, N1741, N1487, N1166);
and AND2 (N1746, N1737, N1559);
nor NOR4 (N1747, N1744, N960, N1294, N718);
nand NAND4 (N1748, N1742, N1584, N890, N1200);
nand NAND4 (N1749, N1725, N902, N743, N812);
or OR3 (N1750, N1743, N1519, N70);
not NOT1 (N1751, N1729);
nor NOR3 (N1752, N1745, N696, N1239);
buf BUF1 (N1753, N1751);
nor NOR3 (N1754, N1747, N413, N30);
or OR3 (N1755, N1754, N1693, N1174);
nor NOR3 (N1756, N1731, N1076, N1131);
buf BUF1 (N1757, N1748);
buf BUF1 (N1758, N1757);
buf BUF1 (N1759, N1758);
nand NAND2 (N1760, N1753, N1607);
or OR2 (N1761, N1756, N1399);
or OR4 (N1762, N1746, N368, N1549, N46);
xor XOR2 (N1763, N1759, N1728);
xor XOR2 (N1764, N1738, N1412);
nor NOR2 (N1765, N1735, N823);
and AND3 (N1766, N1761, N933, N1634);
xor XOR2 (N1767, N1763, N48);
or OR3 (N1768, N1750, N968, N1472);
and AND3 (N1769, N1764, N54, N645);
nor NOR4 (N1770, N1749, N90, N1224, N416);
xor XOR2 (N1771, N1770, N1388);
nor NOR3 (N1772, N1771, N289, N329);
not NOT1 (N1773, N1769);
not NOT1 (N1774, N1765);
nand NAND3 (N1775, N1768, N441, N1565);
not NOT1 (N1776, N1775);
not NOT1 (N1777, N1755);
and AND3 (N1778, N1774, N204, N346);
not NOT1 (N1779, N1777);
buf BUF1 (N1780, N1773);
nor NOR2 (N1781, N1779, N401);
buf BUF1 (N1782, N1781);
xor XOR2 (N1783, N1760, N1620);
and AND3 (N1784, N1752, N1175, N916);
not NOT1 (N1785, N1762);
nand NAND3 (N1786, N1782, N554, N156);
nand NAND3 (N1787, N1780, N898, N446);
or OR3 (N1788, N1787, N184, N306);
and AND3 (N1789, N1772, N900, N1658);
or OR4 (N1790, N1767, N1315, N37, N627);
and AND2 (N1791, N1783, N735);
xor XOR2 (N1792, N1789, N485);
buf BUF1 (N1793, N1790);
and AND3 (N1794, N1792, N495, N738);
or OR3 (N1795, N1785, N1092, N1600);
or OR4 (N1796, N1794, N567, N1222, N955);
not NOT1 (N1797, N1766);
xor XOR2 (N1798, N1791, N1699);
buf BUF1 (N1799, N1793);
or OR4 (N1800, N1784, N949, N463, N45);
or OR3 (N1801, N1778, N1316, N1649);
buf BUF1 (N1802, N1795);
nand NAND3 (N1803, N1797, N1548, N1405);
and AND4 (N1804, N1776, N967, N1638, N1284);
buf BUF1 (N1805, N1802);
or OR4 (N1806, N1805, N786, N957, N1103);
or OR4 (N1807, N1788, N1777, N1783, N1614);
or OR2 (N1808, N1801, N1423);
buf BUF1 (N1809, N1808);
xor XOR2 (N1810, N1786, N425);
nand NAND2 (N1811, N1804, N419);
or OR3 (N1812, N1809, N1069, N1710);
nand NAND3 (N1813, N1807, N876, N860);
not NOT1 (N1814, N1806);
not NOT1 (N1815, N1799);
nor NOR4 (N1816, N1813, N522, N394, N1527);
nor NOR3 (N1817, N1811, N359, N1613);
and AND4 (N1818, N1817, N703, N774, N1035);
nand NAND2 (N1819, N1810, N1280);
xor XOR2 (N1820, N1819, N1669);
nand NAND4 (N1821, N1820, N862, N782, N1527);
buf BUF1 (N1822, N1796);
xor XOR2 (N1823, N1814, N1807);
or OR3 (N1824, N1803, N1179, N223);
buf BUF1 (N1825, N1816);
and AND4 (N1826, N1823, N858, N1623, N1005);
xor XOR2 (N1827, N1821, N155);
nor NOR4 (N1828, N1815, N368, N1154, N1063);
and AND2 (N1829, N1825, N762);
not NOT1 (N1830, N1818);
nor NOR3 (N1831, N1812, N1407, N1218);
not NOT1 (N1832, N1829);
or OR3 (N1833, N1827, N1592, N1234);
nand NAND2 (N1834, N1800, N280);
nand NAND2 (N1835, N1798, N1140);
nor NOR4 (N1836, N1830, N116, N540, N607);
nor NOR3 (N1837, N1833, N952, N368);
nand NAND4 (N1838, N1836, N1757, N580, N393);
and AND2 (N1839, N1834, N399);
and AND3 (N1840, N1826, N1639, N45);
buf BUF1 (N1841, N1840);
xor XOR2 (N1842, N1837, N225);
nor NOR4 (N1843, N1841, N342, N436, N253);
not NOT1 (N1844, N1842);
nor NOR3 (N1845, N1824, N332, N1676);
nand NAND4 (N1846, N1828, N1444, N786, N1571);
not NOT1 (N1847, N1838);
buf BUF1 (N1848, N1832);
nor NOR2 (N1849, N1831, N588);
xor XOR2 (N1850, N1848, N351);
or OR4 (N1851, N1839, N52, N1327, N930);
not NOT1 (N1852, N1845);
not NOT1 (N1853, N1850);
or OR3 (N1854, N1847, N509, N355);
not NOT1 (N1855, N1854);
buf BUF1 (N1856, N1843);
buf BUF1 (N1857, N1822);
nor NOR2 (N1858, N1856, N410);
and AND4 (N1859, N1853, N462, N92, N1237);
nand NAND2 (N1860, N1851, N1308);
buf BUF1 (N1861, N1859);
or OR2 (N1862, N1844, N1229);
nor NOR4 (N1863, N1858, N1085, N1341, N364);
not NOT1 (N1864, N1861);
not NOT1 (N1865, N1852);
not NOT1 (N1866, N1835);
nand NAND3 (N1867, N1855, N576, N638);
xor XOR2 (N1868, N1865, N1080);
xor XOR2 (N1869, N1857, N1225);
xor XOR2 (N1870, N1866, N557);
nand NAND2 (N1871, N1868, N901);
nand NAND3 (N1872, N1867, N1726, N679);
nor NOR4 (N1873, N1849, N1235, N193, N690);
buf BUF1 (N1874, N1872);
and AND4 (N1875, N1871, N1583, N281, N456);
or OR3 (N1876, N1875, N821, N43);
buf BUF1 (N1877, N1873);
buf BUF1 (N1878, N1860);
xor XOR2 (N1879, N1869, N21);
buf BUF1 (N1880, N1876);
xor XOR2 (N1881, N1880, N1033);
nand NAND3 (N1882, N1874, N1484, N837);
or OR2 (N1883, N1881, N1832);
not NOT1 (N1884, N1878);
buf BUF1 (N1885, N1864);
or OR2 (N1886, N1877, N1036);
and AND3 (N1887, N1879, N1158, N1289);
xor XOR2 (N1888, N1885, N1388);
and AND4 (N1889, N1886, N784, N79, N1457);
not NOT1 (N1890, N1887);
buf BUF1 (N1891, N1883);
nand NAND4 (N1892, N1870, N268, N1081, N1810);
nor NOR2 (N1893, N1884, N758);
not NOT1 (N1894, N1890);
or OR4 (N1895, N1893, N1568, N1530, N35);
buf BUF1 (N1896, N1895);
not NOT1 (N1897, N1846);
not NOT1 (N1898, N1889);
or OR3 (N1899, N1862, N1011, N235);
xor XOR2 (N1900, N1863, N411);
not NOT1 (N1901, N1882);
and AND4 (N1902, N1901, N50, N166, N1460);
xor XOR2 (N1903, N1891, N374);
nor NOR2 (N1904, N1899, N81);
buf BUF1 (N1905, N1897);
or OR2 (N1906, N1900, N1507);
xor XOR2 (N1907, N1896, N1046);
or OR4 (N1908, N1904, N22, N602, N546);
and AND2 (N1909, N1905, N254);
nor NOR4 (N1910, N1909, N961, N1709, N1000);
xor XOR2 (N1911, N1908, N1548);
or OR3 (N1912, N1910, N1700, N1550);
buf BUF1 (N1913, N1907);
or OR3 (N1914, N1888, N1283, N24);
nor NOR2 (N1915, N1906, N1277);
not NOT1 (N1916, N1898);
and AND3 (N1917, N1915, N435, N1024);
not NOT1 (N1918, N1912);
not NOT1 (N1919, N1917);
buf BUF1 (N1920, N1894);
buf BUF1 (N1921, N1918);
or OR4 (N1922, N1913, N1681, N435, N923);
buf BUF1 (N1923, N1921);
xor XOR2 (N1924, N1903, N1779);
not NOT1 (N1925, N1911);
xor XOR2 (N1926, N1920, N1014);
nor NOR4 (N1927, N1914, N370, N1192, N773);
buf BUF1 (N1928, N1923);
and AND3 (N1929, N1924, N1403, N829);
xor XOR2 (N1930, N1927, N753);
and AND4 (N1931, N1922, N1238, N249, N1254);
nand NAND3 (N1932, N1931, N247, N1428);
nor NOR4 (N1933, N1930, N792, N612, N627);
nand NAND3 (N1934, N1928, N1658, N1839);
not NOT1 (N1935, N1902);
nor NOR2 (N1936, N1932, N313);
buf BUF1 (N1937, N1936);
or OR2 (N1938, N1935, N265);
and AND2 (N1939, N1925, N533);
not NOT1 (N1940, N1939);
nand NAND3 (N1941, N1929, N1693, N444);
xor XOR2 (N1942, N1892, N1924);
not NOT1 (N1943, N1926);
nand NAND4 (N1944, N1937, N210, N1011, N1578);
and AND2 (N1945, N1941, N1490);
buf BUF1 (N1946, N1942);
nand NAND2 (N1947, N1916, N1299);
nand NAND4 (N1948, N1933, N1080, N429, N1561);
nor NOR4 (N1949, N1944, N622, N1268, N176);
not NOT1 (N1950, N1934);
xor XOR2 (N1951, N1943, N1835);
and AND3 (N1952, N1938, N268, N480);
nand NAND2 (N1953, N1949, N591);
and AND2 (N1954, N1946, N1335);
nand NAND4 (N1955, N1947, N974, N970, N414);
nand NAND2 (N1956, N1953, N1047);
not NOT1 (N1957, N1951);
not NOT1 (N1958, N1948);
nand NAND2 (N1959, N1919, N738);
or OR3 (N1960, N1945, N1816, N424);
xor XOR2 (N1961, N1959, N1908);
or OR3 (N1962, N1955, N1798, N1380);
buf BUF1 (N1963, N1940);
xor XOR2 (N1964, N1960, N1368);
nand NAND4 (N1965, N1964, N196, N1415, N1835);
not NOT1 (N1966, N1957);
buf BUF1 (N1967, N1958);
or OR4 (N1968, N1965, N1182, N382, N1230);
nor NOR4 (N1969, N1956, N1158, N1473, N829);
nor NOR2 (N1970, N1968, N1585);
xor XOR2 (N1971, N1967, N223);
nand NAND4 (N1972, N1966, N1578, N1048, N850);
or OR4 (N1973, N1970, N1477, N1103, N1403);
nor NOR4 (N1974, N1963, N465, N837, N1960);
and AND4 (N1975, N1973, N311, N482, N1166);
not NOT1 (N1976, N1969);
not NOT1 (N1977, N1975);
or OR2 (N1978, N1974, N1815);
xor XOR2 (N1979, N1971, N1636);
buf BUF1 (N1980, N1962);
and AND3 (N1981, N1952, N1190, N664);
buf BUF1 (N1982, N1961);
nand NAND4 (N1983, N1980, N573, N183, N1782);
xor XOR2 (N1984, N1979, N976);
nor NOR4 (N1985, N1954, N240, N342, N712);
not NOT1 (N1986, N1981);
or OR3 (N1987, N1984, N1242, N1945);
and AND4 (N1988, N1976, N1407, N466, N1661);
nand NAND4 (N1989, N1983, N367, N1133, N836);
buf BUF1 (N1990, N1977);
or OR3 (N1991, N1987, N858, N30);
xor XOR2 (N1992, N1985, N1857);
not NOT1 (N1993, N1992);
nand NAND3 (N1994, N1972, N152, N930);
buf BUF1 (N1995, N1991);
nor NOR2 (N1996, N1994, N520);
xor XOR2 (N1997, N1986, N1475);
buf BUF1 (N1998, N1988);
and AND3 (N1999, N1950, N391, N1879);
and AND4 (N2000, N1998, N1519, N773, N1223);
nor NOR3 (N2001, N1989, N255, N953);
buf BUF1 (N2002, N1978);
and AND3 (N2003, N2002, N1101, N1339);
xor XOR2 (N2004, N1990, N1053);
xor XOR2 (N2005, N2001, N1633);
nand NAND3 (N2006, N2004, N1424, N756);
or OR2 (N2007, N1982, N1600);
nor NOR2 (N2008, N2003, N1563);
nor NOR4 (N2009, N1993, N442, N1587, N1071);
nand NAND4 (N2010, N1995, N248, N1791, N1008);
not NOT1 (N2011, N2007);
buf BUF1 (N2012, N1999);
nor NOR4 (N2013, N2011, N1691, N800, N971);
or OR2 (N2014, N2009, N1391);
buf BUF1 (N2015, N2012);
buf BUF1 (N2016, N2015);
nand NAND2 (N2017, N2008, N975);
and AND3 (N2018, N2010, N1017, N1806);
nand NAND3 (N2019, N2018, N1328, N334);
and AND3 (N2020, N2014, N1511, N965);
nand NAND4 (N2021, N2016, N400, N1123, N1325);
not NOT1 (N2022, N1996);
nor NOR3 (N2023, N2020, N1552, N1059);
and AND2 (N2024, N2021, N1534);
xor XOR2 (N2025, N2024, N1596);
buf BUF1 (N2026, N2025);
buf BUF1 (N2027, N2019);
or OR3 (N2028, N2023, N433, N22);
nor NOR4 (N2029, N2017, N706, N16, N279);
not NOT1 (N2030, N2022);
xor XOR2 (N2031, N2006, N1615);
not NOT1 (N2032, N1997);
nor NOR4 (N2033, N2005, N2022, N593, N1115);
not NOT1 (N2034, N2028);
nand NAND4 (N2035, N2029, N129, N918, N1803);
and AND2 (N2036, N2030, N388);
buf BUF1 (N2037, N2033);
xor XOR2 (N2038, N2034, N1450);
or OR4 (N2039, N2000, N1317, N1254, N678);
not NOT1 (N2040, N2037);
and AND4 (N2041, N2013, N781, N1536, N588);
and AND3 (N2042, N2040, N466, N1370);
nor NOR4 (N2043, N2038, N71, N1637, N300);
or OR2 (N2044, N2032, N533);
nand NAND4 (N2045, N2042, N1267, N890, N1385);
and AND4 (N2046, N2026, N1126, N779, N419);
buf BUF1 (N2047, N2031);
buf BUF1 (N2048, N2039);
nand NAND4 (N2049, N2048, N1252, N1038, N267);
or OR4 (N2050, N2041, N787, N1186, N1174);
xor XOR2 (N2051, N2050, N938);
buf BUF1 (N2052, N2036);
buf BUF1 (N2053, N2045);
or OR4 (N2054, N2043, N700, N111, N145);
not NOT1 (N2055, N2052);
buf BUF1 (N2056, N2044);
or OR4 (N2057, N2056, N1621, N839, N1525);
and AND2 (N2058, N2057, N416);
or OR3 (N2059, N2053, N792, N743);
and AND2 (N2060, N2051, N1328);
nand NAND2 (N2061, N2054, N1154);
buf BUF1 (N2062, N2046);
buf BUF1 (N2063, N2062);
xor XOR2 (N2064, N2060, N959);
or OR3 (N2065, N2063, N1427, N1107);
nand NAND4 (N2066, N2055, N1259, N84, N1146);
nand NAND3 (N2067, N2049, N562, N249);
buf BUF1 (N2068, N2067);
not NOT1 (N2069, N2061);
and AND2 (N2070, N2058, N207);
and AND4 (N2071, N2035, N408, N1016, N694);
nor NOR2 (N2072, N2047, N2036);
not NOT1 (N2073, N2065);
xor XOR2 (N2074, N2073, N7);
or OR3 (N2075, N2059, N837, N1899);
not NOT1 (N2076, N2071);
or OR3 (N2077, N2074, N332, N51);
nand NAND2 (N2078, N2070, N357);
buf BUF1 (N2079, N2078);
buf BUF1 (N2080, N2027);
nand NAND2 (N2081, N2064, N1358);
nor NOR4 (N2082, N2079, N1911, N1304, N1566);
nand NAND3 (N2083, N2081, N338, N1164);
nand NAND3 (N2084, N2076, N2048, N727);
or OR3 (N2085, N2077, N1397, N1341);
nand NAND2 (N2086, N2082, N1672);
nand NAND3 (N2087, N2066, N1716, N925);
and AND2 (N2088, N2084, N71);
not NOT1 (N2089, N2068);
buf BUF1 (N2090, N2089);
and AND3 (N2091, N2090, N882, N1578);
xor XOR2 (N2092, N2080, N1772);
or OR3 (N2093, N2087, N1682, N467);
and AND3 (N2094, N2069, N1419, N1397);
buf BUF1 (N2095, N2092);
xor XOR2 (N2096, N2088, N803);
buf BUF1 (N2097, N2094);
buf BUF1 (N2098, N2072);
nor NOR4 (N2099, N2091, N870, N1105, N1718);
and AND4 (N2100, N2083, N945, N269, N629);
or OR4 (N2101, N2093, N2066, N1815, N305);
buf BUF1 (N2102, N2085);
not NOT1 (N2103, N2075);
nor NOR4 (N2104, N2096, N1205, N1334, N1408);
and AND3 (N2105, N2095, N1845, N1095);
or OR4 (N2106, N2098, N933, N697, N304);
nor NOR4 (N2107, N2101, N508, N953, N1672);
xor XOR2 (N2108, N2105, N905);
xor XOR2 (N2109, N2097, N250);
or OR2 (N2110, N2107, N916);
nor NOR2 (N2111, N2109, N122);
xor XOR2 (N2112, N2110, N1960);
xor XOR2 (N2113, N2112, N995);
or OR3 (N2114, N2106, N1232, N525);
xor XOR2 (N2115, N2111, N2063);
nand NAND2 (N2116, N2115, N119);
buf BUF1 (N2117, N2108);
or OR3 (N2118, N2100, N814, N1165);
or OR3 (N2119, N2114, N645, N137);
and AND4 (N2120, N2116, N2039, N2005, N1921);
xor XOR2 (N2121, N2120, N919);
xor XOR2 (N2122, N2099, N109);
and AND2 (N2123, N2102, N1891);
nor NOR4 (N2124, N2117, N1157, N738, N1459);
nand NAND4 (N2125, N2104, N714, N315, N1706);
nand NAND3 (N2126, N2086, N2087, N661);
or OR3 (N2127, N2103, N1517, N682);
not NOT1 (N2128, N2123);
nand NAND2 (N2129, N2118, N323);
and AND3 (N2130, N2119, N1458, N933);
or OR4 (N2131, N2121, N1479, N1693, N1682);
and AND3 (N2132, N2131, N324, N1771);
nand NAND2 (N2133, N2113, N2002);
or OR3 (N2134, N2129, N759, N1911);
buf BUF1 (N2135, N2126);
not NOT1 (N2136, N2130);
xor XOR2 (N2137, N2125, N1899);
and AND3 (N2138, N2127, N1624, N1480);
nor NOR4 (N2139, N2133, N1352, N1205, N640);
nand NAND2 (N2140, N2138, N1735);
or OR4 (N2141, N2132, N1178, N744, N408);
xor XOR2 (N2142, N2124, N251);
or OR2 (N2143, N2140, N1441);
and AND3 (N2144, N2141, N606, N1828);
not NOT1 (N2145, N2143);
nand NAND2 (N2146, N2135, N830);
xor XOR2 (N2147, N2144, N1202);
nand NAND2 (N2148, N2142, N1501);
nor NOR3 (N2149, N2147, N1505, N1461);
buf BUF1 (N2150, N2128);
and AND2 (N2151, N2145, N1989);
nor NOR3 (N2152, N2148, N82, N1130);
xor XOR2 (N2153, N2151, N46);
nand NAND4 (N2154, N2146, N1018, N1930, N2012);
buf BUF1 (N2155, N2139);
and AND2 (N2156, N2153, N546);
xor XOR2 (N2157, N2134, N897);
and AND4 (N2158, N2122, N1391, N1800, N1960);
xor XOR2 (N2159, N2137, N995);
nor NOR4 (N2160, N2152, N925, N52, N1086);
buf BUF1 (N2161, N2160);
nor NOR3 (N2162, N2150, N1100, N864);
buf BUF1 (N2163, N2149);
nand NAND2 (N2164, N2159, N1594);
not NOT1 (N2165, N2163);
nand NAND4 (N2166, N2136, N104, N269, N893);
buf BUF1 (N2167, N2165);
not NOT1 (N2168, N2154);
or OR4 (N2169, N2164, N369, N915, N1250);
xor XOR2 (N2170, N2158, N29);
and AND3 (N2171, N2156, N1285, N236);
or OR3 (N2172, N2162, N1135, N1743);
or OR3 (N2173, N2167, N1206, N1617);
nor NOR3 (N2174, N2169, N1343, N2093);
buf BUF1 (N2175, N2170);
xor XOR2 (N2176, N2171, N415);
buf BUF1 (N2177, N2155);
and AND3 (N2178, N2176, N1324, N1789);
nand NAND4 (N2179, N2161, N80, N1346, N569);
nor NOR2 (N2180, N2157, N547);
or OR3 (N2181, N2178, N453, N1590);
nand NAND4 (N2182, N2179, N1086, N1734, N2042);
nor NOR2 (N2183, N2175, N289);
or OR2 (N2184, N2181, N162);
and AND2 (N2185, N2183, N617);
or OR4 (N2186, N2177, N133, N437, N4);
or OR4 (N2187, N2172, N1917, N265, N1617);
nor NOR2 (N2188, N2168, N390);
nand NAND2 (N2189, N2188, N1425);
or OR3 (N2190, N2166, N635, N1152);
not NOT1 (N2191, N2185);
not NOT1 (N2192, N2189);
or OR2 (N2193, N2186, N612);
nand NAND4 (N2194, N2173, N626, N1343, N1777);
nor NOR4 (N2195, N2184, N2192, N754, N1443);
xor XOR2 (N2196, N1449, N1429);
not NOT1 (N2197, N2191);
xor XOR2 (N2198, N2174, N1780);
or OR3 (N2199, N2194, N420, N2186);
xor XOR2 (N2200, N2195, N993);
nand NAND2 (N2201, N2197, N1636);
not NOT1 (N2202, N2182);
xor XOR2 (N2203, N2201, N475);
not NOT1 (N2204, N2202);
not NOT1 (N2205, N2187);
buf BUF1 (N2206, N2196);
nand NAND3 (N2207, N2199, N1107, N519);
nor NOR3 (N2208, N2180, N1043, N2114);
buf BUF1 (N2209, N2204);
or OR4 (N2210, N2208, N621, N1415, N1174);
buf BUF1 (N2211, N2206);
buf BUF1 (N2212, N2211);
or OR4 (N2213, N2198, N1636, N1675, N318);
nand NAND4 (N2214, N2210, N94, N73, N1221);
buf BUF1 (N2215, N2193);
or OR3 (N2216, N2200, N2034, N689);
buf BUF1 (N2217, N2209);
nor NOR3 (N2218, N2216, N1885, N2195);
or OR4 (N2219, N2205, N24, N1, N1773);
buf BUF1 (N2220, N2219);
not NOT1 (N2221, N2207);
not NOT1 (N2222, N2214);
and AND2 (N2223, N2217, N751);
xor XOR2 (N2224, N2203, N2157);
not NOT1 (N2225, N2212);
buf BUF1 (N2226, N2223);
xor XOR2 (N2227, N2218, N2139);
or OR3 (N2228, N2220, N795, N1728);
or OR2 (N2229, N2222, N1559);
xor XOR2 (N2230, N2227, N1476);
nor NOR2 (N2231, N2213, N684);
buf BUF1 (N2232, N2230);
buf BUF1 (N2233, N2225);
buf BUF1 (N2234, N2215);
nand NAND4 (N2235, N2234, N813, N1143, N1496);
xor XOR2 (N2236, N2229, N651);
xor XOR2 (N2237, N2232, N1174);
buf BUF1 (N2238, N2237);
not NOT1 (N2239, N2235);
and AND2 (N2240, N2238, N899);
xor XOR2 (N2241, N2236, N1831);
nand NAND4 (N2242, N2224, N2061, N229, N54);
nor NOR4 (N2243, N2242, N1844, N194, N1564);
buf BUF1 (N2244, N2233);
xor XOR2 (N2245, N2239, N1679);
nand NAND3 (N2246, N2190, N758, N1131);
nor NOR3 (N2247, N2244, N972, N1808);
and AND3 (N2248, N2228, N710, N237);
not NOT1 (N2249, N2245);
xor XOR2 (N2250, N2246, N1861);
xor XOR2 (N2251, N2249, N1307);
not NOT1 (N2252, N2241);
nor NOR4 (N2253, N2243, N1553, N497, N136);
nand NAND2 (N2254, N2250, N941);
nand NAND3 (N2255, N2253, N837, N1319);
not NOT1 (N2256, N2231);
xor XOR2 (N2257, N2247, N1330);
not NOT1 (N2258, N2226);
or OR2 (N2259, N2252, N1165);
not NOT1 (N2260, N2258);
nand NAND2 (N2261, N2240, N797);
xor XOR2 (N2262, N2260, N1255);
not NOT1 (N2263, N2251);
or OR3 (N2264, N2262, N2029, N1298);
nor NOR2 (N2265, N2259, N505);
nand NAND4 (N2266, N2265, N2100, N551, N1339);
or OR2 (N2267, N2264, N135);
and AND4 (N2268, N2261, N570, N2168, N1567);
xor XOR2 (N2269, N2248, N614);
nor NOR2 (N2270, N2268, N92);
nand NAND4 (N2271, N2269, N175, N792, N1575);
and AND4 (N2272, N2254, N2129, N1056, N1071);
xor XOR2 (N2273, N2266, N257);
not NOT1 (N2274, N2256);
xor XOR2 (N2275, N2272, N1912);
nor NOR3 (N2276, N2221, N692, N1221);
or OR4 (N2277, N2257, N706, N1218, N122);
buf BUF1 (N2278, N2263);
and AND3 (N2279, N2276, N1686, N1566);
nand NAND4 (N2280, N2271, N559, N306, N2203);
or OR2 (N2281, N2267, N887);
buf BUF1 (N2282, N2273);
or OR3 (N2283, N2274, N1744, N261);
and AND3 (N2284, N2275, N536, N322);
not NOT1 (N2285, N2280);
and AND2 (N2286, N2283, N1872);
nand NAND2 (N2287, N2277, N2093);
buf BUF1 (N2288, N2255);
nand NAND4 (N2289, N2285, N1435, N723, N1245);
and AND2 (N2290, N2288, N1866);
buf BUF1 (N2291, N2286);
nor NOR4 (N2292, N2284, N977, N1182, N1048);
or OR2 (N2293, N2282, N1993);
xor XOR2 (N2294, N2292, N2088);
buf BUF1 (N2295, N2293);
buf BUF1 (N2296, N2279);
not NOT1 (N2297, N2281);
nand NAND2 (N2298, N2278, N48);
xor XOR2 (N2299, N2295, N1528);
nand NAND4 (N2300, N2297, N1232, N1291, N1707);
and AND4 (N2301, N2270, N657, N1245, N745);
or OR4 (N2302, N2300, N857, N954, N230);
or OR3 (N2303, N2294, N921, N1074);
nand NAND3 (N2304, N2291, N252, N1167);
buf BUF1 (N2305, N2289);
or OR2 (N2306, N2287, N1949);
and AND4 (N2307, N2305, N262, N1125, N2153);
nor NOR3 (N2308, N2296, N1013, N346);
not NOT1 (N2309, N2306);
or OR4 (N2310, N2298, N2129, N1481, N166);
and AND3 (N2311, N2301, N2069, N1172);
or OR3 (N2312, N2309, N1857, N110);
and AND4 (N2313, N2310, N67, N1081, N1152);
buf BUF1 (N2314, N2312);
nor NOR2 (N2315, N2313, N2238);
nor NOR3 (N2316, N2303, N1981, N178);
xor XOR2 (N2317, N2290, N1112);
not NOT1 (N2318, N2314);
xor XOR2 (N2319, N2302, N447);
nor NOR3 (N2320, N2319, N636, N1773);
nand NAND2 (N2321, N2299, N355);
or OR2 (N2322, N2311, N2308);
xor XOR2 (N2323, N2173, N1363);
not NOT1 (N2324, N2321);
and AND4 (N2325, N2315, N1503, N467, N1394);
nand NAND3 (N2326, N2324, N1227, N908);
xor XOR2 (N2327, N2325, N1495);
or OR3 (N2328, N2307, N1660, N1365);
xor XOR2 (N2329, N2323, N239);
nor NOR2 (N2330, N2317, N2093);
xor XOR2 (N2331, N2328, N1629);
buf BUF1 (N2332, N2320);
buf BUF1 (N2333, N2330);
and AND2 (N2334, N2326, N1291);
and AND4 (N2335, N2316, N940, N647, N830);
nor NOR2 (N2336, N2322, N2309);
buf BUF1 (N2337, N2336);
xor XOR2 (N2338, N2337, N39);
xor XOR2 (N2339, N2332, N49);
nand NAND2 (N2340, N2335, N1961);
nor NOR2 (N2341, N2318, N2283);
nand NAND2 (N2342, N2331, N1586);
buf BUF1 (N2343, N2333);
nor NOR4 (N2344, N2342, N2238, N225, N1002);
not NOT1 (N2345, N2344);
xor XOR2 (N2346, N2345, N1806);
xor XOR2 (N2347, N2304, N2015);
nor NOR3 (N2348, N2346, N172, N1352);
nor NOR3 (N2349, N2341, N227, N1174);
xor XOR2 (N2350, N2340, N2151);
xor XOR2 (N2351, N2338, N1477);
nand NAND2 (N2352, N2350, N2051);
xor XOR2 (N2353, N2343, N1671);
and AND4 (N2354, N2327, N1958, N1847, N683);
and AND2 (N2355, N2351, N981);
buf BUF1 (N2356, N2339);
buf BUF1 (N2357, N2356);
nand NAND4 (N2358, N2329, N670, N2033, N405);
not NOT1 (N2359, N2347);
or OR4 (N2360, N2359, N1833, N2316, N885);
nor NOR4 (N2361, N2357, N945, N1086, N1116);
or OR2 (N2362, N2361, N68);
nor NOR2 (N2363, N2353, N2261);
buf BUF1 (N2364, N2358);
nand NAND4 (N2365, N2363, N283, N1974, N1631);
xor XOR2 (N2366, N2360, N460);
buf BUF1 (N2367, N2348);
buf BUF1 (N2368, N2367);
and AND3 (N2369, N2352, N1469, N1679);
buf BUF1 (N2370, N2362);
buf BUF1 (N2371, N2368);
buf BUF1 (N2372, N2365);
nor NOR4 (N2373, N2370, N1072, N1905, N2019);
and AND2 (N2374, N2369, N458);
nand NAND4 (N2375, N2372, N652, N2194, N1776);
and AND3 (N2376, N2334, N1812, N189);
xor XOR2 (N2377, N2364, N397);
xor XOR2 (N2378, N2373, N1146);
nand NAND4 (N2379, N2376, N1275, N1633, N1997);
or OR2 (N2380, N2378, N811);
buf BUF1 (N2381, N2355);
or OR4 (N2382, N2380, N1796, N1453, N1884);
xor XOR2 (N2383, N2374, N1364);
nand NAND3 (N2384, N2375, N970, N2319);
nor NOR4 (N2385, N2384, N1824, N914, N1620);
buf BUF1 (N2386, N2383);
or OR2 (N2387, N2366, N979);
and AND2 (N2388, N2379, N857);
xor XOR2 (N2389, N2349, N905);
and AND3 (N2390, N2388, N2278, N685);
nor NOR4 (N2391, N2382, N429, N184, N2320);
nand NAND3 (N2392, N2354, N1654, N2173);
and AND4 (N2393, N2377, N1945, N1035, N2069);
nand NAND2 (N2394, N2392, N617);
buf BUF1 (N2395, N2385);
buf BUF1 (N2396, N2395);
buf BUF1 (N2397, N2387);
xor XOR2 (N2398, N2389, N662);
buf BUF1 (N2399, N2394);
or OR2 (N2400, N2391, N2327);
buf BUF1 (N2401, N2397);
xor XOR2 (N2402, N2400, N2362);
nand NAND2 (N2403, N2386, N639);
and AND4 (N2404, N2403, N1152, N207, N1512);
xor XOR2 (N2405, N2402, N2154);
buf BUF1 (N2406, N2396);
buf BUF1 (N2407, N2381);
xor XOR2 (N2408, N2405, N1908);
buf BUF1 (N2409, N2399);
buf BUF1 (N2410, N2390);
or OR2 (N2411, N2410, N1289);
and AND2 (N2412, N2401, N1971);
not NOT1 (N2413, N2407);
nand NAND4 (N2414, N2398, N471, N676, N926);
or OR3 (N2415, N2404, N2279, N1538);
or OR3 (N2416, N2413, N1512, N1975);
or OR3 (N2417, N2415, N1303, N239);
or OR3 (N2418, N2393, N709, N1339);
and AND2 (N2419, N2416, N2090);
or OR2 (N2420, N2412, N5);
not NOT1 (N2421, N2411);
or OR2 (N2422, N2420, N872);
not NOT1 (N2423, N2414);
nor NOR4 (N2424, N2406, N614, N159, N577);
or OR4 (N2425, N2417, N1240, N1462, N434);
buf BUF1 (N2426, N2408);
nor NOR3 (N2427, N2419, N180, N764);
xor XOR2 (N2428, N2421, N812);
nand NAND4 (N2429, N2425, N1165, N2294, N2381);
buf BUF1 (N2430, N2423);
nand NAND4 (N2431, N2409, N1533, N2344, N1541);
nand NAND4 (N2432, N2430, N2077, N1954, N332);
or OR4 (N2433, N2422, N2413, N2186, N841);
buf BUF1 (N2434, N2433);
nor NOR2 (N2435, N2426, N1373);
and AND3 (N2436, N2428, N2086, N1324);
nor NOR2 (N2437, N2432, N819);
or OR2 (N2438, N2431, N1180);
not NOT1 (N2439, N2424);
nand NAND3 (N2440, N2429, N332, N448);
and AND3 (N2441, N2436, N124, N2056);
nand NAND2 (N2442, N2371, N240);
buf BUF1 (N2443, N2438);
buf BUF1 (N2444, N2427);
or OR3 (N2445, N2439, N1068, N20);
nand NAND4 (N2446, N2435, N2266, N390, N1405);
xor XOR2 (N2447, N2444, N2084);
and AND2 (N2448, N2418, N1304);
xor XOR2 (N2449, N2440, N518);
buf BUF1 (N2450, N2434);
and AND2 (N2451, N2447, N2070);
xor XOR2 (N2452, N2445, N68);
xor XOR2 (N2453, N2437, N1714);
not NOT1 (N2454, N2442);
nand NAND2 (N2455, N2451, N2073);
or OR2 (N2456, N2449, N295);
nand NAND4 (N2457, N2441, N54, N567, N1070);
buf BUF1 (N2458, N2455);
or OR2 (N2459, N2446, N2092);
or OR4 (N2460, N2448, N2458, N2272, N707);
xor XOR2 (N2461, N1514, N1016);
or OR3 (N2462, N2454, N283, N271);
or OR4 (N2463, N2457, N1087, N1047, N1612);
nand NAND4 (N2464, N2462, N2023, N2114, N745);
or OR3 (N2465, N2450, N1376, N1089);
not NOT1 (N2466, N2459);
buf BUF1 (N2467, N2443);
or OR2 (N2468, N2461, N1411);
and AND4 (N2469, N2467, N1644, N1040, N199);
buf BUF1 (N2470, N2456);
buf BUF1 (N2471, N2460);
or OR2 (N2472, N2469, N2448);
and AND2 (N2473, N2470, N2117);
and AND2 (N2474, N2465, N2073);
or OR4 (N2475, N2464, N1096, N1057, N1991);
not NOT1 (N2476, N2468);
buf BUF1 (N2477, N2475);
xor XOR2 (N2478, N2472, N2230);
nand NAND3 (N2479, N2452, N391, N161);
xor XOR2 (N2480, N2479, N215);
or OR2 (N2481, N2474, N276);
xor XOR2 (N2482, N2471, N2433);
xor XOR2 (N2483, N2480, N1176);
and AND2 (N2484, N2463, N503);
nor NOR4 (N2485, N2473, N610, N933, N1129);
nand NAND4 (N2486, N2477, N2083, N1309, N1738);
or OR4 (N2487, N2453, N2042, N1979, N2139);
or OR3 (N2488, N2486, N269, N511);
nor NOR2 (N2489, N2487, N1199);
and AND2 (N2490, N2489, N1617);
or OR3 (N2491, N2488, N1243, N2276);
nand NAND3 (N2492, N2481, N1570, N611);
xor XOR2 (N2493, N2478, N1165);
not NOT1 (N2494, N2492);
nand NAND3 (N2495, N2466, N214, N1323);
and AND4 (N2496, N2476, N118, N1553, N1252);
or OR3 (N2497, N2490, N1264, N46);
or OR4 (N2498, N2497, N951, N777, N470);
buf BUF1 (N2499, N2496);
nand NAND3 (N2500, N2485, N275, N1484);
not NOT1 (N2501, N2494);
or OR3 (N2502, N2491, N1737, N367);
nand NAND3 (N2503, N2482, N1539, N1001);
buf BUF1 (N2504, N2495);
nor NOR4 (N2505, N2503, N145, N2166, N1219);
xor XOR2 (N2506, N2484, N2214);
nand NAND4 (N2507, N2493, N1362, N1480, N2118);
not NOT1 (N2508, N2501);
nor NOR3 (N2509, N2498, N839, N726);
nand NAND3 (N2510, N2506, N383, N1143);
buf BUF1 (N2511, N2505);
nor NOR2 (N2512, N2502, N1817);
nor NOR4 (N2513, N2504, N986, N152, N11);
nand NAND2 (N2514, N2507, N2132);
nand NAND2 (N2515, N2510, N433);
and AND3 (N2516, N2511, N1943, N1071);
buf BUF1 (N2517, N2509);
nor NOR4 (N2518, N2516, N1744, N1934, N173);
and AND2 (N2519, N2518, N301);
buf BUF1 (N2520, N2514);
xor XOR2 (N2521, N2519, N2462);
nor NOR3 (N2522, N2517, N970, N717);
xor XOR2 (N2523, N2513, N1930);
and AND4 (N2524, N2512, N1407, N1066, N1315);
nand NAND2 (N2525, N2500, N2243);
and AND3 (N2526, N2523, N368, N1308);
xor XOR2 (N2527, N2524, N859);
nor NOR3 (N2528, N2515, N1451, N780);
nand NAND4 (N2529, N2483, N746, N960, N1925);
xor XOR2 (N2530, N2499, N1718);
and AND2 (N2531, N2530, N463);
and AND2 (N2532, N2528, N682);
xor XOR2 (N2533, N2531, N1426);
nor NOR2 (N2534, N2520, N1586);
nor NOR4 (N2535, N2529, N474, N1924, N2227);
or OR3 (N2536, N2526, N2365, N2461);
nand NAND2 (N2537, N2535, N1763);
nand NAND4 (N2538, N2508, N2355, N2001, N2351);
nor NOR2 (N2539, N2537, N89);
or OR3 (N2540, N2525, N2405, N400);
and AND4 (N2541, N2540, N1996, N2208, N2136);
nand NAND2 (N2542, N2539, N1854);
buf BUF1 (N2543, N2538);
not NOT1 (N2544, N2534);
nor NOR3 (N2545, N2533, N838, N2028);
nor NOR3 (N2546, N2541, N2535, N1570);
or OR3 (N2547, N2521, N2297, N51);
not NOT1 (N2548, N2532);
not NOT1 (N2549, N2522);
buf BUF1 (N2550, N2547);
not NOT1 (N2551, N2543);
or OR3 (N2552, N2546, N687, N2313);
or OR2 (N2553, N2551, N986);
nand NAND3 (N2554, N2548, N365, N1923);
xor XOR2 (N2555, N2544, N1418);
buf BUF1 (N2556, N2536);
nand NAND2 (N2557, N2545, N2314);
not NOT1 (N2558, N2556);
xor XOR2 (N2559, N2550, N44);
not NOT1 (N2560, N2559);
buf BUF1 (N2561, N2558);
and AND3 (N2562, N2560, N495, N96);
buf BUF1 (N2563, N2554);
not NOT1 (N2564, N2563);
or OR4 (N2565, N2553, N674, N862, N1476);
buf BUF1 (N2566, N2552);
not NOT1 (N2567, N2564);
nor NOR3 (N2568, N2567, N709, N1661);
nor NOR3 (N2569, N2549, N607, N407);
xor XOR2 (N2570, N2542, N420);
nand NAND4 (N2571, N2565, N2260, N1280, N2120);
and AND3 (N2572, N2561, N1318, N780);
xor XOR2 (N2573, N2527, N2370);
xor XOR2 (N2574, N2562, N1283);
not NOT1 (N2575, N2566);
and AND3 (N2576, N2570, N2419, N2365);
nand NAND2 (N2577, N2572, N1249);
buf BUF1 (N2578, N2568);
xor XOR2 (N2579, N2575, N124);
or OR4 (N2580, N2557, N1210, N2290, N634);
nand NAND2 (N2581, N2576, N518);
xor XOR2 (N2582, N2581, N858);
buf BUF1 (N2583, N2579);
xor XOR2 (N2584, N2578, N300);
nor NOR2 (N2585, N2577, N1128);
xor XOR2 (N2586, N2584, N160);
nor NOR4 (N2587, N2582, N892, N1746, N25);
nor NOR3 (N2588, N2580, N1114, N568);
or OR3 (N2589, N2569, N185, N912);
nor NOR4 (N2590, N2571, N443, N1941, N828);
xor XOR2 (N2591, N2573, N126);
not NOT1 (N2592, N2589);
not NOT1 (N2593, N2587);
nand NAND2 (N2594, N2592, N1812);
buf BUF1 (N2595, N2586);
or OR4 (N2596, N2594, N223, N736, N2456);
and AND2 (N2597, N2588, N69);
xor XOR2 (N2598, N2591, N2088);
and AND3 (N2599, N2583, N216, N376);
buf BUF1 (N2600, N2597);
not NOT1 (N2601, N2598);
nand NAND4 (N2602, N2601, N700, N439, N434);
buf BUF1 (N2603, N2590);
and AND4 (N2604, N2555, N2235, N100, N1812);
nand NAND3 (N2605, N2603, N46, N118);
xor XOR2 (N2606, N2599, N2001);
buf BUF1 (N2607, N2602);
nor NOR4 (N2608, N2596, N1112, N2598, N1600);
not NOT1 (N2609, N2585);
and AND3 (N2610, N2608, N902, N2399);
xor XOR2 (N2611, N2595, N1887);
nand NAND4 (N2612, N2611, N1430, N558, N1706);
not NOT1 (N2613, N2605);
xor XOR2 (N2614, N2610, N892);
xor XOR2 (N2615, N2593, N1682);
or OR3 (N2616, N2612, N822, N1531);
buf BUF1 (N2617, N2604);
not NOT1 (N2618, N2609);
xor XOR2 (N2619, N2617, N1876);
nor NOR4 (N2620, N2615, N930, N1956, N1402);
not NOT1 (N2621, N2616);
and AND2 (N2622, N2600, N1229);
xor XOR2 (N2623, N2574, N853);
not NOT1 (N2624, N2619);
xor XOR2 (N2625, N2620, N1833);
and AND3 (N2626, N2613, N1488, N2370);
xor XOR2 (N2627, N2622, N1209);
buf BUF1 (N2628, N2626);
xor XOR2 (N2629, N2621, N995);
and AND2 (N2630, N2618, N1749);
not NOT1 (N2631, N2628);
nand NAND2 (N2632, N2627, N696);
nand NAND3 (N2633, N2631, N1669, N1803);
buf BUF1 (N2634, N2607);
and AND4 (N2635, N2606, N2195, N1597, N2114);
buf BUF1 (N2636, N2633);
nor NOR4 (N2637, N2614, N2486, N2437, N1244);
and AND4 (N2638, N2632, N806, N1176, N1609);
not NOT1 (N2639, N2638);
xor XOR2 (N2640, N2636, N1877);
xor XOR2 (N2641, N2640, N215);
and AND3 (N2642, N2634, N1902, N2428);
xor XOR2 (N2643, N2637, N1745);
nand NAND2 (N2644, N2625, N1042);
nor NOR3 (N2645, N2639, N1383, N2637);
and AND2 (N2646, N2645, N2118);
xor XOR2 (N2647, N2643, N1889);
and AND4 (N2648, N2624, N2434, N1310, N2314);
and AND2 (N2649, N2629, N456);
not NOT1 (N2650, N2648);
xor XOR2 (N2651, N2641, N1719);
nor NOR2 (N2652, N2642, N408);
or OR2 (N2653, N2650, N2135);
buf BUF1 (N2654, N2647);
not NOT1 (N2655, N2646);
buf BUF1 (N2656, N2653);
nand NAND3 (N2657, N2652, N1966, N11);
not NOT1 (N2658, N2644);
buf BUF1 (N2659, N2651);
buf BUF1 (N2660, N2623);
or OR4 (N2661, N2659, N2620, N317, N358);
nand NAND3 (N2662, N2654, N1646, N1860);
not NOT1 (N2663, N2655);
or OR2 (N2664, N2656, N648);
buf BUF1 (N2665, N2657);
or OR3 (N2666, N2630, N1853, N467);
buf BUF1 (N2667, N2649);
xor XOR2 (N2668, N2666, N1406);
or OR2 (N2669, N2661, N2276);
xor XOR2 (N2670, N2635, N2556);
buf BUF1 (N2671, N2660);
buf BUF1 (N2672, N2662);
and AND3 (N2673, N2672, N254, N258);
nand NAND4 (N2674, N2667, N1986, N2310, N1394);
nor NOR2 (N2675, N2670, N2022);
nand NAND2 (N2676, N2675, N2368);
not NOT1 (N2677, N2658);
nor NOR3 (N2678, N2674, N709, N1783);
nor NOR4 (N2679, N2669, N75, N1294, N2397);
xor XOR2 (N2680, N2679, N1158);
xor XOR2 (N2681, N2664, N2204);
xor XOR2 (N2682, N2676, N1165);
not NOT1 (N2683, N2665);
or OR2 (N2684, N2683, N624);
or OR4 (N2685, N2663, N1014, N1165, N2472);
and AND2 (N2686, N2678, N1667);
and AND4 (N2687, N2668, N88, N1497, N1640);
not NOT1 (N2688, N2681);
nand NAND3 (N2689, N2682, N1405, N1353);
nand NAND3 (N2690, N2684, N1902, N123);
nand NAND4 (N2691, N2680, N1841, N1511, N1532);
or OR3 (N2692, N2677, N466, N51);
xor XOR2 (N2693, N2692, N1329);
or OR3 (N2694, N2690, N668, N2083);
nand NAND2 (N2695, N2685, N395);
and AND3 (N2696, N2689, N2503, N2208);
not NOT1 (N2697, N2673);
nand NAND2 (N2698, N2693, N227);
nand NAND2 (N2699, N2687, N1250);
and AND2 (N2700, N2694, N2334);
or OR3 (N2701, N2688, N714, N2362);
not NOT1 (N2702, N2700);
nand NAND4 (N2703, N2698, N2444, N2453, N2293);
or OR2 (N2704, N2696, N2665);
nor NOR4 (N2705, N2691, N2405, N2254, N325);
or OR3 (N2706, N2705, N2593, N1871);
buf BUF1 (N2707, N2702);
not NOT1 (N2708, N2707);
nand NAND4 (N2709, N2703, N437, N343, N1637);
nor NOR4 (N2710, N2709, N2011, N1541, N229);
xor XOR2 (N2711, N2699, N2196);
nor NOR3 (N2712, N2697, N1294, N606);
not NOT1 (N2713, N2710);
xor XOR2 (N2714, N2686, N1855);
and AND3 (N2715, N2701, N773, N1200);
buf BUF1 (N2716, N2704);
buf BUF1 (N2717, N2714);
or OR4 (N2718, N2711, N1190, N777, N521);
buf BUF1 (N2719, N2671);
xor XOR2 (N2720, N2706, N1869);
or OR2 (N2721, N2715, N2201);
nand NAND4 (N2722, N2718, N846, N1287, N687);
nand NAND2 (N2723, N2716, N1066);
not NOT1 (N2724, N2721);
xor XOR2 (N2725, N2717, N570);
or OR3 (N2726, N2722, N881, N2125);
or OR3 (N2727, N2712, N290, N1449);
nand NAND3 (N2728, N2726, N146, N2372);
or OR2 (N2729, N2724, N1573);
nand NAND4 (N2730, N2727, N1097, N414, N1037);
buf BUF1 (N2731, N2695);
nand NAND4 (N2732, N2729, N2484, N414, N2477);
xor XOR2 (N2733, N2708, N894);
buf BUF1 (N2734, N2725);
not NOT1 (N2735, N2728);
xor XOR2 (N2736, N2734, N1489);
buf BUF1 (N2737, N2719);
xor XOR2 (N2738, N2730, N746);
buf BUF1 (N2739, N2713);
nand NAND2 (N2740, N2720, N1088);
or OR3 (N2741, N2739, N2728, N2273);
not NOT1 (N2742, N2741);
nand NAND3 (N2743, N2731, N1696, N436);
nor NOR2 (N2744, N2737, N1399);
not NOT1 (N2745, N2744);
xor XOR2 (N2746, N2742, N22);
and AND3 (N2747, N2733, N1959, N941);
or OR2 (N2748, N2735, N392);
xor XOR2 (N2749, N2738, N947);
nor NOR3 (N2750, N2749, N258, N2430);
buf BUF1 (N2751, N2745);
or OR3 (N2752, N2723, N666, N749);
buf BUF1 (N2753, N2732);
and AND3 (N2754, N2740, N2282, N1597);
and AND4 (N2755, N2754, N489, N1663, N685);
and AND3 (N2756, N2750, N1756, N1446);
or OR4 (N2757, N2736, N2507, N1294, N817);
and AND4 (N2758, N2743, N1507, N337, N802);
nor NOR4 (N2759, N2757, N1051, N2305, N1626);
nand NAND2 (N2760, N2759, N2570);
or OR2 (N2761, N2756, N1859);
not NOT1 (N2762, N2751);
and AND2 (N2763, N2755, N1929);
nor NOR3 (N2764, N2746, N393, N2300);
xor XOR2 (N2765, N2758, N2117);
and AND3 (N2766, N2747, N348, N1843);
or OR2 (N2767, N2766, N2093);
and AND3 (N2768, N2748, N2466, N1535);
xor XOR2 (N2769, N2762, N417);
buf BUF1 (N2770, N2765);
xor XOR2 (N2771, N2752, N2496);
xor XOR2 (N2772, N2771, N2700);
or OR3 (N2773, N2753, N2753, N1988);
nand NAND4 (N2774, N2769, N2323, N1814, N2569);
buf BUF1 (N2775, N2768);
and AND2 (N2776, N2761, N385);
xor XOR2 (N2777, N2775, N835);
nand NAND3 (N2778, N2763, N2244, N741);
or OR3 (N2779, N2774, N2368, N2431);
nor NOR3 (N2780, N2779, N2654, N1960);
not NOT1 (N2781, N2778);
and AND4 (N2782, N2781, N2441, N361, N358);
not NOT1 (N2783, N2782);
and AND2 (N2784, N2776, N443);
or OR4 (N2785, N2773, N1900, N2699, N1990);
or OR4 (N2786, N2785, N308, N1880, N395);
not NOT1 (N2787, N2770);
and AND3 (N2788, N2772, N473, N376);
or OR4 (N2789, N2786, N402, N2255, N803);
not NOT1 (N2790, N2780);
not NOT1 (N2791, N2777);
nand NAND2 (N2792, N2760, N1492);
xor XOR2 (N2793, N2788, N1878);
and AND4 (N2794, N2783, N1205, N1701, N2522);
and AND2 (N2795, N2787, N908);
xor XOR2 (N2796, N2794, N2077);
nor NOR2 (N2797, N2795, N980);
nand NAND4 (N2798, N2790, N756, N882, N1307);
not NOT1 (N2799, N2798);
not NOT1 (N2800, N2799);
and AND4 (N2801, N2784, N2626, N2383, N997);
nand NAND2 (N2802, N2792, N405);
buf BUF1 (N2803, N2789);
xor XOR2 (N2804, N2791, N2062);
not NOT1 (N2805, N2796);
buf BUF1 (N2806, N2764);
nor NOR2 (N2807, N2803, N89);
not NOT1 (N2808, N2800);
buf BUF1 (N2809, N2806);
xor XOR2 (N2810, N2804, N389);
nand NAND4 (N2811, N2767, N940, N834, N271);
buf BUF1 (N2812, N2793);
nand NAND3 (N2813, N2805, N2216, N394);
nand NAND2 (N2814, N2811, N431);
buf BUF1 (N2815, N2802);
nor NOR3 (N2816, N2801, N1571, N1846);
and AND4 (N2817, N2815, N1196, N2288, N898);
xor XOR2 (N2818, N2810, N53);
not NOT1 (N2819, N2812);
and AND2 (N2820, N2819, N2475);
and AND4 (N2821, N2813, N1405, N1958, N1479);
buf BUF1 (N2822, N2797);
not NOT1 (N2823, N2817);
not NOT1 (N2824, N2821);
or OR3 (N2825, N2820, N871, N1324);
nor NOR2 (N2826, N2809, N893);
nand NAND2 (N2827, N2823, N2740);
not NOT1 (N2828, N2816);
buf BUF1 (N2829, N2826);
not NOT1 (N2830, N2818);
or OR4 (N2831, N2822, N210, N1703, N1298);
nor NOR3 (N2832, N2827, N1870, N319);
xor XOR2 (N2833, N2808, N1823);
or OR3 (N2834, N2828, N612, N910);
nand NAND4 (N2835, N2814, N674, N201, N2461);
not NOT1 (N2836, N2835);
xor XOR2 (N2837, N2830, N2626);
or OR3 (N2838, N2831, N662, N862);
nand NAND4 (N2839, N2824, N497, N2791, N2449);
xor XOR2 (N2840, N2834, N603);
and AND3 (N2841, N2829, N2243, N2071);
xor XOR2 (N2842, N2807, N2409);
xor XOR2 (N2843, N2836, N948);
or OR4 (N2844, N2842, N1670, N1933, N844);
or OR3 (N2845, N2837, N2299, N1691);
xor XOR2 (N2846, N2845, N1141);
xor XOR2 (N2847, N2844, N38);
not NOT1 (N2848, N2841);
xor XOR2 (N2849, N2840, N2250);
or OR4 (N2850, N2843, N2227, N2003, N19);
and AND3 (N2851, N2850, N1699, N1479);
nor NOR2 (N2852, N2847, N2448);
or OR3 (N2853, N2851, N1478, N300);
xor XOR2 (N2854, N2833, N1877);
buf BUF1 (N2855, N2839);
xor XOR2 (N2856, N2852, N2421);
not NOT1 (N2857, N2832);
buf BUF1 (N2858, N2848);
and AND3 (N2859, N2854, N2196, N2689);
xor XOR2 (N2860, N2838, N2294);
buf BUF1 (N2861, N2825);
buf BUF1 (N2862, N2858);
nand NAND4 (N2863, N2862, N2136, N427, N1198);
nand NAND3 (N2864, N2863, N287, N1606);
nand NAND4 (N2865, N2856, N1355, N2025, N661);
buf BUF1 (N2866, N2865);
or OR3 (N2867, N2860, N697, N2846);
xor XOR2 (N2868, N2775, N1342);
or OR4 (N2869, N2857, N671, N1035, N1905);
xor XOR2 (N2870, N2869, N125);
xor XOR2 (N2871, N2849, N503);
or OR4 (N2872, N2870, N1958, N2441, N986);
and AND2 (N2873, N2864, N1936);
buf BUF1 (N2874, N2868);
not NOT1 (N2875, N2874);
nand NAND2 (N2876, N2871, N181);
and AND4 (N2877, N2867, N459, N1687, N1739);
or OR3 (N2878, N2853, N2408, N2651);
nand NAND2 (N2879, N2855, N1245);
buf BUF1 (N2880, N2878);
xor XOR2 (N2881, N2876, N712);
not NOT1 (N2882, N2879);
and AND4 (N2883, N2866, N2265, N204, N337);
nor NOR4 (N2884, N2872, N1591, N2763, N472);
or OR3 (N2885, N2883, N1776, N1447);
buf BUF1 (N2886, N2880);
or OR4 (N2887, N2875, N569, N2514, N953);
nand NAND2 (N2888, N2861, N1881);
nor NOR4 (N2889, N2885, N2433, N1943, N256);
not NOT1 (N2890, N2888);
or OR4 (N2891, N2884, N903, N419, N1402);
xor XOR2 (N2892, N2882, N1119);
xor XOR2 (N2893, N2886, N1681);
nor NOR4 (N2894, N2877, N2582, N140, N52);
buf BUF1 (N2895, N2889);
or OR4 (N2896, N2895, N1281, N568, N1460);
or OR3 (N2897, N2859, N851, N690);
and AND3 (N2898, N2873, N2063, N1397);
nor NOR2 (N2899, N2898, N2512);
nor NOR4 (N2900, N2891, N824, N147, N173);
or OR3 (N2901, N2899, N675, N2879);
nor NOR3 (N2902, N2896, N1802, N170);
xor XOR2 (N2903, N2902, N2069);
nand NAND3 (N2904, N2894, N1387, N1722);
buf BUF1 (N2905, N2900);
or OR4 (N2906, N2887, N2085, N157, N2516);
nand NAND4 (N2907, N2901, N1681, N486, N1542);
and AND2 (N2908, N2907, N208);
or OR4 (N2909, N2892, N571, N1145, N2409);
and AND2 (N2910, N2890, N969);
or OR3 (N2911, N2908, N654, N1942);
nor NOR3 (N2912, N2910, N2038, N2281);
not NOT1 (N2913, N2903);
not NOT1 (N2914, N2905);
and AND4 (N2915, N2912, N1741, N2791, N1795);
nand NAND2 (N2916, N2913, N2752);
nand NAND2 (N2917, N2909, N1440);
and AND2 (N2918, N2917, N765);
and AND3 (N2919, N2911, N2680, N835);
not NOT1 (N2920, N2906);
buf BUF1 (N2921, N2916);
not NOT1 (N2922, N2881);
xor XOR2 (N2923, N2921, N1732);
nor NOR4 (N2924, N2919, N2915, N2386, N2377);
xor XOR2 (N2925, N68, N1155);
buf BUF1 (N2926, N2924);
xor XOR2 (N2927, N2897, N1786);
nand NAND3 (N2928, N2922, N2491, N100);
nor NOR2 (N2929, N2918, N1027);
and AND2 (N2930, N2893, N1439);
and AND3 (N2931, N2926, N2537, N1183);
nand NAND4 (N2932, N2931, N1840, N760, N2587);
nand NAND2 (N2933, N2904, N2058);
not NOT1 (N2934, N2914);
buf BUF1 (N2935, N2930);
and AND4 (N2936, N2928, N787, N725, N2550);
buf BUF1 (N2937, N2936);
or OR2 (N2938, N2937, N1092);
or OR3 (N2939, N2925, N2736, N2801);
buf BUF1 (N2940, N2923);
and AND3 (N2941, N2938, N2358, N741);
nor NOR4 (N2942, N2935, N1501, N2212, N897);
nand NAND4 (N2943, N2932, N835, N2552, N504);
nand NAND3 (N2944, N2941, N893, N813);
nor NOR3 (N2945, N2942, N2316, N2114);
or OR2 (N2946, N2920, N1363);
or OR3 (N2947, N2943, N1942, N403);
not NOT1 (N2948, N2945);
and AND2 (N2949, N2947, N1556);
not NOT1 (N2950, N2940);
not NOT1 (N2951, N2933);
and AND2 (N2952, N2944, N2634);
or OR2 (N2953, N2948, N2264);
nor NOR4 (N2954, N2953, N1882, N2775, N2274);
not NOT1 (N2955, N2950);
nand NAND4 (N2956, N2934, N2128, N510, N948);
xor XOR2 (N2957, N2929, N1523);
nand NAND3 (N2958, N2927, N1335, N369);
nor NOR4 (N2959, N2952, N2169, N1602, N2021);
xor XOR2 (N2960, N2939, N2238);
not NOT1 (N2961, N2954);
or OR3 (N2962, N2949, N555, N927);
xor XOR2 (N2963, N2962, N88);
nor NOR2 (N2964, N2958, N2274);
buf BUF1 (N2965, N2957);
buf BUF1 (N2966, N2960);
xor XOR2 (N2967, N2965, N650);
buf BUF1 (N2968, N2966);
xor XOR2 (N2969, N2968, N1217);
nor NOR4 (N2970, N2969, N758, N1295, N1610);
nor NOR2 (N2971, N2956, N1528);
nor NOR3 (N2972, N2961, N1846, N956);
nor NOR3 (N2973, N2951, N1543, N2913);
nor NOR2 (N2974, N2955, N2904);
nor NOR3 (N2975, N2964, N455, N1167);
and AND3 (N2976, N2975, N758, N1623);
xor XOR2 (N2977, N2976, N2351);
or OR3 (N2978, N2959, N2051, N173);
nor NOR4 (N2979, N2970, N1971, N1186, N2225);
and AND3 (N2980, N2978, N883, N93);
nor NOR4 (N2981, N2979, N2925, N1018, N620);
and AND4 (N2982, N2972, N1445, N2190, N2220);
nand NAND4 (N2983, N2982, N2401, N1670, N275);
buf BUF1 (N2984, N2971);
or OR2 (N2985, N2980, N78);
or OR4 (N2986, N2981, N2912, N1239, N1013);
and AND4 (N2987, N2985, N320, N1528, N2663);
and AND2 (N2988, N2963, N219);
nor NOR2 (N2989, N2946, N440);
or OR3 (N2990, N2986, N2038, N1999);
buf BUF1 (N2991, N2989);
nand NAND2 (N2992, N2988, N676);
xor XOR2 (N2993, N2983, N1713);
nor NOR3 (N2994, N2977, N576, N1039);
xor XOR2 (N2995, N2984, N2311);
or OR2 (N2996, N2994, N2928);
xor XOR2 (N2997, N2996, N213);
and AND2 (N2998, N2995, N1203);
xor XOR2 (N2999, N2987, N2448);
nand NAND4 (N3000, N2967, N417, N1418, N11);
nand NAND2 (N3001, N2997, N793);
nor NOR3 (N3002, N3000, N999, N81);
nor NOR3 (N3003, N2990, N1638, N971);
not NOT1 (N3004, N2993);
buf BUF1 (N3005, N2991);
buf BUF1 (N3006, N2999);
nor NOR4 (N3007, N2992, N815, N680, N2838);
or OR4 (N3008, N3007, N664, N2260, N1109);
buf BUF1 (N3009, N3006);
buf BUF1 (N3010, N3002);
buf BUF1 (N3011, N2973);
nand NAND2 (N3012, N3011, N2452);
nor NOR3 (N3013, N3001, N1546, N339);
nand NAND3 (N3014, N3005, N1250, N2731);
or OR2 (N3015, N3008, N1324);
xor XOR2 (N3016, N3009, N2155);
nor NOR2 (N3017, N2998, N2754);
nor NOR3 (N3018, N3012, N2673, N1617);
and AND4 (N3019, N3018, N1220, N1098, N893);
buf BUF1 (N3020, N3010);
xor XOR2 (N3021, N3004, N1739);
nand NAND4 (N3022, N3013, N190, N1960, N1477);
xor XOR2 (N3023, N3022, N2580);
xor XOR2 (N3024, N3023, N1546);
xor XOR2 (N3025, N3019, N1603);
nand NAND2 (N3026, N3003, N2292);
not NOT1 (N3027, N3014);
nor NOR4 (N3028, N3017, N1399, N2257, N1068);
nand NAND2 (N3029, N3021, N1843);
buf BUF1 (N3030, N3024);
buf BUF1 (N3031, N3028);
nor NOR3 (N3032, N3020, N644, N1304);
xor XOR2 (N3033, N3032, N2247);
or OR2 (N3034, N3026, N2213);
and AND2 (N3035, N3025, N2306);
nand NAND4 (N3036, N3027, N727, N2654, N1662);
nand NAND3 (N3037, N3035, N1332, N1227);
nor NOR4 (N3038, N3015, N2987, N2086, N367);
nand NAND4 (N3039, N3036, N2660, N1455, N1636);
xor XOR2 (N3040, N3031, N1772);
or OR2 (N3041, N3039, N645);
nand NAND4 (N3042, N3034, N261, N2725, N1189);
buf BUF1 (N3043, N3041);
nor NOR4 (N3044, N3042, N848, N2458, N942);
and AND3 (N3045, N3029, N1221, N2635);
or OR4 (N3046, N2974, N2879, N1580, N370);
buf BUF1 (N3047, N3045);
or OR4 (N3048, N3037, N439, N1126, N2359);
nor NOR3 (N3049, N3046, N2872, N694);
and AND3 (N3050, N3030, N1548, N2702);
not NOT1 (N3051, N3044);
nand NAND3 (N3052, N3049, N722, N1269);
buf BUF1 (N3053, N3052);
or OR3 (N3054, N3038, N323, N2293);
or OR2 (N3055, N3033, N2210);
nor NOR3 (N3056, N3053, N2411, N974);
nand NAND3 (N3057, N3043, N1085, N2125);
not NOT1 (N3058, N3048);
buf BUF1 (N3059, N3016);
nand NAND3 (N3060, N3051, N316, N1068);
nand NAND2 (N3061, N3054, N2072);
not NOT1 (N3062, N3055);
or OR3 (N3063, N3057, N2987, N2988);
nand NAND4 (N3064, N3050, N1011, N487, N2857);
buf BUF1 (N3065, N3063);
and AND3 (N3066, N3065, N1231, N1347);
not NOT1 (N3067, N3056);
nor NOR3 (N3068, N3064, N2668, N1729);
not NOT1 (N3069, N3068);
or OR4 (N3070, N3066, N1658, N1353, N90);
nand NAND4 (N3071, N3040, N2396, N2710, N2996);
buf BUF1 (N3072, N3067);
xor XOR2 (N3073, N3071, N835);
buf BUF1 (N3074, N3072);
nor NOR4 (N3075, N3069, N1739, N2993, N2095);
and AND2 (N3076, N3062, N1132);
nand NAND2 (N3077, N3075, N1642);
not NOT1 (N3078, N3076);
or OR3 (N3079, N3059, N2594, N2858);
nor NOR4 (N3080, N3079, N1326, N2763, N2584);
and AND3 (N3081, N3074, N995, N2482);
nand NAND2 (N3082, N3060, N477);
xor XOR2 (N3083, N3058, N2539);
nand NAND3 (N3084, N3083, N537, N1023);
xor XOR2 (N3085, N3082, N484);
nor NOR3 (N3086, N3078, N339, N1470);
nor NOR3 (N3087, N3070, N643, N1608);
nor NOR3 (N3088, N3061, N91, N2525);
buf BUF1 (N3089, N3081);
xor XOR2 (N3090, N3089, N2364);
nor NOR2 (N3091, N3073, N2307);
xor XOR2 (N3092, N3084, N3000);
not NOT1 (N3093, N3085);
nand NAND3 (N3094, N3090, N683, N25);
buf BUF1 (N3095, N3086);
xor XOR2 (N3096, N3080, N92);
or OR4 (N3097, N3093, N2338, N149, N679);
xor XOR2 (N3098, N3092, N2687);
or OR3 (N3099, N3047, N2040, N577);
nand NAND4 (N3100, N3098, N1150, N2845, N1593);
nand NAND2 (N3101, N3100, N78);
and AND2 (N3102, N3088, N1871);
nand NAND4 (N3103, N3102, N3056, N1541, N995);
nand NAND4 (N3104, N3077, N2156, N2959, N1220);
buf BUF1 (N3105, N3094);
xor XOR2 (N3106, N3105, N3008);
or OR2 (N3107, N3087, N216);
or OR4 (N3108, N3099, N2551, N1148, N2729);
not NOT1 (N3109, N3101);
nor NOR2 (N3110, N3109, N557);
and AND2 (N3111, N3106, N669);
and AND4 (N3112, N3104, N803, N1559, N1572);
nand NAND3 (N3113, N3103, N302, N6);
or OR3 (N3114, N3108, N2736, N2943);
not NOT1 (N3115, N3095);
or OR2 (N3116, N3114, N2107);
nor NOR4 (N3117, N3097, N1800, N1549, N936);
or OR3 (N3118, N3096, N2251, N1684);
or OR3 (N3119, N3113, N149, N1989);
and AND4 (N3120, N3115, N2765, N1680, N1757);
buf BUF1 (N3121, N3116);
and AND4 (N3122, N3118, N462, N2665, N1887);
nor NOR3 (N3123, N3111, N1173, N712);
not NOT1 (N3124, N3107);
and AND2 (N3125, N3122, N396);
and AND4 (N3126, N3117, N2567, N949, N863);
or OR3 (N3127, N3126, N948, N2440);
buf BUF1 (N3128, N3127);
not NOT1 (N3129, N3128);
and AND4 (N3130, N3120, N2072, N2739, N213);
nor NOR3 (N3131, N3130, N1671, N793);
nor NOR3 (N3132, N3125, N2672, N401);
nor NOR3 (N3133, N3119, N346, N659);
xor XOR2 (N3134, N3091, N2947);
nand NAND4 (N3135, N3129, N1567, N2226, N620);
xor XOR2 (N3136, N3121, N562);
nor NOR4 (N3137, N3124, N2541, N1659, N2413);
xor XOR2 (N3138, N3123, N2497);
and AND3 (N3139, N3136, N2565, N802);
or OR3 (N3140, N3137, N2059, N97);
xor XOR2 (N3141, N3139, N314);
and AND4 (N3142, N3138, N1072, N1284, N649);
not NOT1 (N3143, N3140);
and AND4 (N3144, N3112, N776, N2514, N1474);
not NOT1 (N3145, N3135);
xor XOR2 (N3146, N3143, N985);
nor NOR3 (N3147, N3110, N2483, N2490);
buf BUF1 (N3148, N3142);
not NOT1 (N3149, N3148);
not NOT1 (N3150, N3149);
or OR4 (N3151, N3145, N1968, N1176, N1189);
not NOT1 (N3152, N3147);
not NOT1 (N3153, N3144);
or OR4 (N3154, N3134, N2372, N497, N3048);
not NOT1 (N3155, N3131);
and AND2 (N3156, N3133, N1517);
nand NAND2 (N3157, N3155, N2473);
buf BUF1 (N3158, N3132);
or OR4 (N3159, N3141, N1158, N2991, N2667);
and AND2 (N3160, N3156, N966);
nand NAND3 (N3161, N3151, N889, N1663);
not NOT1 (N3162, N3152);
or OR4 (N3163, N3150, N542, N1559, N316);
not NOT1 (N3164, N3160);
buf BUF1 (N3165, N3164);
buf BUF1 (N3166, N3153);
and AND2 (N3167, N3158, N2293);
nor NOR4 (N3168, N3163, N2192, N2310, N1868);
nor NOR3 (N3169, N3157, N2238, N2391);
and AND3 (N3170, N3161, N604, N152);
xor XOR2 (N3171, N3166, N2923);
nor NOR4 (N3172, N3171, N1545, N2491, N1319);
nand NAND4 (N3173, N3170, N223, N174, N2384);
xor XOR2 (N3174, N3162, N597);
nor NOR4 (N3175, N3173, N2636, N1363, N2827);
and AND4 (N3176, N3169, N2649, N131, N1922);
nand NAND2 (N3177, N3146, N35);
xor XOR2 (N3178, N3174, N2322);
nand NAND4 (N3179, N3176, N3081, N2921, N446);
nand NAND4 (N3180, N3154, N1121, N2764, N665);
buf BUF1 (N3181, N3159);
or OR4 (N3182, N3181, N394, N120, N33);
xor XOR2 (N3183, N3167, N662);
or OR2 (N3184, N3179, N457);
xor XOR2 (N3185, N3182, N2934);
not NOT1 (N3186, N3185);
nand NAND3 (N3187, N3175, N2528, N2959);
not NOT1 (N3188, N3172);
buf BUF1 (N3189, N3178);
nor NOR4 (N3190, N3168, N1433, N168, N1216);
not NOT1 (N3191, N3190);
not NOT1 (N3192, N3189);
not NOT1 (N3193, N3180);
xor XOR2 (N3194, N3177, N1258);
not NOT1 (N3195, N3194);
and AND3 (N3196, N3192, N2994, N2717);
nor NOR3 (N3197, N3183, N2250, N2021);
not NOT1 (N3198, N3193);
or OR4 (N3199, N3188, N948, N1042, N2395);
nor NOR3 (N3200, N3187, N823, N2313);
nor NOR2 (N3201, N3165, N1820);
nor NOR4 (N3202, N3184, N227, N14, N2371);
nor NOR4 (N3203, N3200, N2103, N754, N1580);
nor NOR2 (N3204, N3198, N2985);
buf BUF1 (N3205, N3203);
not NOT1 (N3206, N3199);
or OR3 (N3207, N3204, N3035, N1960);
not NOT1 (N3208, N3196);
nand NAND2 (N3209, N3206, N2985);
xor XOR2 (N3210, N3207, N1432);
xor XOR2 (N3211, N3205, N1348);
buf BUF1 (N3212, N3201);
nand NAND2 (N3213, N3211, N860);
nor NOR3 (N3214, N3202, N2262, N3130);
nor NOR2 (N3215, N3209, N307);
buf BUF1 (N3216, N3197);
buf BUF1 (N3217, N3215);
or OR2 (N3218, N3210, N2205);
nand NAND3 (N3219, N3214, N2555, N978);
and AND3 (N3220, N3213, N1139, N1936);
not NOT1 (N3221, N3212);
not NOT1 (N3222, N3208);
or OR4 (N3223, N3216, N238, N2987, N2064);
xor XOR2 (N3224, N3195, N838);
xor XOR2 (N3225, N3219, N1832);
nor NOR2 (N3226, N3218, N1627);
and AND2 (N3227, N3191, N1009);
xor XOR2 (N3228, N3217, N119);
not NOT1 (N3229, N3223);
buf BUF1 (N3230, N3220);
buf BUF1 (N3231, N3221);
or OR3 (N3232, N3186, N2185, N3158);
and AND2 (N3233, N3227, N617);
nor NOR2 (N3234, N3222, N332);
or OR3 (N3235, N3232, N1048, N1319);
nor NOR2 (N3236, N3226, N3166);
nand NAND4 (N3237, N3225, N931, N2910, N1377);
and AND3 (N3238, N3230, N1115, N1179);
nor NOR4 (N3239, N3236, N1319, N2653, N95);
nor NOR2 (N3240, N3235, N740);
and AND3 (N3241, N3239, N402, N528);
or OR3 (N3242, N3224, N710, N2416);
or OR3 (N3243, N3242, N1662, N1364);
xor XOR2 (N3244, N3228, N1513);
or OR4 (N3245, N3233, N1857, N1487, N2086);
nand NAND3 (N3246, N3229, N159, N965);
buf BUF1 (N3247, N3234);
buf BUF1 (N3248, N3247);
not NOT1 (N3249, N3240);
and AND2 (N3250, N3246, N574);
buf BUF1 (N3251, N3238);
nor NOR3 (N3252, N3248, N3163, N1075);
or OR4 (N3253, N3252, N1120, N2541, N1223);
not NOT1 (N3254, N3231);
not NOT1 (N3255, N3249);
or OR3 (N3256, N3250, N840, N2177);
nand NAND2 (N3257, N3251, N1380);
nor NOR2 (N3258, N3243, N1623);
and AND4 (N3259, N3257, N952, N2940, N637);
not NOT1 (N3260, N3258);
buf BUF1 (N3261, N3241);
or OR4 (N3262, N3244, N1675, N2097, N1380);
or OR4 (N3263, N3260, N1617, N1262, N1901);
not NOT1 (N3264, N3253);
and AND2 (N3265, N3263, N2249);
buf BUF1 (N3266, N3261);
buf BUF1 (N3267, N3254);
and AND2 (N3268, N3245, N772);
buf BUF1 (N3269, N3256);
and AND2 (N3270, N3255, N1090);
and AND2 (N3271, N3264, N1751);
buf BUF1 (N3272, N3259);
xor XOR2 (N3273, N3270, N720);
and AND3 (N3274, N3268, N2537, N149);
xor XOR2 (N3275, N3272, N1133);
or OR4 (N3276, N3266, N2999, N2966, N542);
buf BUF1 (N3277, N3265);
xor XOR2 (N3278, N3237, N503);
or OR2 (N3279, N3262, N2565);
not NOT1 (N3280, N3269);
not NOT1 (N3281, N3278);
nand NAND2 (N3282, N3273, N1120);
buf BUF1 (N3283, N3277);
nor NOR3 (N3284, N3267, N2336, N2613);
not NOT1 (N3285, N3271);
nor NOR2 (N3286, N3281, N2141);
nor NOR2 (N3287, N3274, N308);
xor XOR2 (N3288, N3284, N62);
or OR4 (N3289, N3276, N1563, N1924, N1107);
or OR3 (N3290, N3283, N348, N680);
buf BUF1 (N3291, N3286);
not NOT1 (N3292, N3285);
nor NOR3 (N3293, N3289, N521, N232);
or OR3 (N3294, N3282, N1550, N2349);
or OR2 (N3295, N3275, N1290);
or OR3 (N3296, N3291, N2774, N2522);
xor XOR2 (N3297, N3295, N2427);
or OR4 (N3298, N3280, N1405, N1562, N1494);
xor XOR2 (N3299, N3288, N1493);
xor XOR2 (N3300, N3296, N259);
and AND3 (N3301, N3279, N2496, N800);
and AND2 (N3302, N3294, N2502);
not NOT1 (N3303, N3298);
xor XOR2 (N3304, N3297, N2611);
xor XOR2 (N3305, N3300, N1361);
nand NAND3 (N3306, N3287, N1185, N420);
nand NAND3 (N3307, N3301, N2723, N624);
nor NOR3 (N3308, N3305, N1410, N1096);
xor XOR2 (N3309, N3293, N2936);
and AND4 (N3310, N3308, N303, N1686, N651);
not NOT1 (N3311, N3290);
or OR3 (N3312, N3302, N2716, N2596);
and AND3 (N3313, N3309, N2151, N853);
nand NAND3 (N3314, N3307, N503, N37);
buf BUF1 (N3315, N3306);
xor XOR2 (N3316, N3313, N1845);
nor NOR3 (N3317, N3310, N2813, N118);
buf BUF1 (N3318, N3312);
and AND3 (N3319, N3304, N1579, N1424);
and AND3 (N3320, N3311, N16, N2814);
xor XOR2 (N3321, N3299, N121);
buf BUF1 (N3322, N3303);
not NOT1 (N3323, N3322);
nand NAND3 (N3324, N3316, N3193, N577);
or OR4 (N3325, N3317, N157, N3231, N2480);
and AND4 (N3326, N3325, N88, N302, N3012);
or OR3 (N3327, N3292, N1943, N2672);
and AND4 (N3328, N3318, N733, N2761, N347);
nand NAND2 (N3329, N3324, N2102);
nor NOR2 (N3330, N3327, N1108);
nor NOR2 (N3331, N3329, N3180);
nand NAND3 (N3332, N3323, N1197, N1219);
nor NOR2 (N3333, N3326, N826);
buf BUF1 (N3334, N3320);
or OR3 (N3335, N3334, N2824, N2222);
and AND2 (N3336, N3321, N289);
nand NAND2 (N3337, N3332, N672);
nand NAND4 (N3338, N3328, N2684, N2204, N300);
xor XOR2 (N3339, N3333, N821);
and AND3 (N3340, N3338, N1967, N1684);
not NOT1 (N3341, N3337);
and AND2 (N3342, N3339, N3154);
xor XOR2 (N3343, N3335, N2134);
buf BUF1 (N3344, N3330);
nor NOR3 (N3345, N3343, N2187, N1984);
nor NOR3 (N3346, N3342, N754, N2230);
not NOT1 (N3347, N3340);
xor XOR2 (N3348, N3341, N993);
nor NOR3 (N3349, N3347, N1723, N2126);
nor NOR4 (N3350, N3344, N465, N1354, N1857);
or OR3 (N3351, N3346, N3232, N1865);
nand NAND2 (N3352, N3348, N1431);
xor XOR2 (N3353, N3350, N3299);
nand NAND2 (N3354, N3315, N1264);
buf BUF1 (N3355, N3351);
not NOT1 (N3356, N3354);
xor XOR2 (N3357, N3356, N1228);
not NOT1 (N3358, N3352);
xor XOR2 (N3359, N3314, N2719);
not NOT1 (N3360, N3353);
and AND4 (N3361, N3349, N2269, N2232, N703);
and AND2 (N3362, N3355, N808);
or OR2 (N3363, N3357, N2355);
buf BUF1 (N3364, N3363);
xor XOR2 (N3365, N3336, N227);
buf BUF1 (N3366, N3319);
not NOT1 (N3367, N3331);
not NOT1 (N3368, N3366);
buf BUF1 (N3369, N3361);
xor XOR2 (N3370, N3368, N713);
buf BUF1 (N3371, N3369);
not NOT1 (N3372, N3345);
nand NAND4 (N3373, N3360, N2807, N148, N3228);
nand NAND3 (N3374, N3370, N449, N2641);
buf BUF1 (N3375, N3373);
nor NOR2 (N3376, N3372, N2507);
and AND3 (N3377, N3358, N1978, N1908);
and AND4 (N3378, N3359, N2155, N329, N2917);
xor XOR2 (N3379, N3377, N2618);
xor XOR2 (N3380, N3364, N2736);
or OR4 (N3381, N3362, N306, N2931, N177);
or OR3 (N3382, N3381, N1311, N1552);
nand NAND3 (N3383, N3376, N1017, N2966);
or OR4 (N3384, N3365, N2349, N2822, N2394);
buf BUF1 (N3385, N3379);
buf BUF1 (N3386, N3385);
nand NAND4 (N3387, N3384, N3122, N291, N1208);
not NOT1 (N3388, N3374);
not NOT1 (N3389, N3375);
and AND2 (N3390, N3371, N1921);
not NOT1 (N3391, N3386);
buf BUF1 (N3392, N3390);
not NOT1 (N3393, N3389);
buf BUF1 (N3394, N3367);
and AND2 (N3395, N3378, N2014);
nor NOR2 (N3396, N3388, N3311);
and AND3 (N3397, N3394, N242, N714);
not NOT1 (N3398, N3380);
nand NAND3 (N3399, N3382, N235, N1341);
not NOT1 (N3400, N3387);
nor NOR4 (N3401, N3400, N2127, N365, N53);
xor XOR2 (N3402, N3399, N1353);
or OR4 (N3403, N3397, N2690, N932, N3059);
xor XOR2 (N3404, N3403, N2231);
not NOT1 (N3405, N3398);
or OR4 (N3406, N3393, N2514, N558, N2770);
not NOT1 (N3407, N3392);
and AND3 (N3408, N3401, N2775, N598);
or OR3 (N3409, N3402, N2832, N1439);
nand NAND3 (N3410, N3391, N1220, N1049);
not NOT1 (N3411, N3383);
nor NOR4 (N3412, N3410, N3369, N298, N687);
not NOT1 (N3413, N3405);
nand NAND2 (N3414, N3409, N461);
xor XOR2 (N3415, N3411, N3292);
or OR4 (N3416, N3404, N1825, N2921, N661);
or OR4 (N3417, N3415, N1221, N2603, N1641);
nand NAND4 (N3418, N3416, N500, N2565, N2566);
buf BUF1 (N3419, N3408);
nor NOR3 (N3420, N3406, N1947, N584);
nor NOR3 (N3421, N3414, N1549, N1585);
buf BUF1 (N3422, N3418);
nor NOR3 (N3423, N3396, N1629, N1537);
nor NOR2 (N3424, N3421, N425);
buf BUF1 (N3425, N3420);
nand NAND3 (N3426, N3425, N699, N1631);
and AND3 (N3427, N3422, N1435, N830);
buf BUF1 (N3428, N3413);
nor NOR3 (N3429, N3407, N1568, N1995);
xor XOR2 (N3430, N3428, N2657);
not NOT1 (N3431, N3423);
and AND2 (N3432, N3395, N3338);
xor XOR2 (N3433, N3417, N459);
nand NAND4 (N3434, N3432, N617, N610, N420);
or OR4 (N3435, N3434, N2215, N2728, N2207);
xor XOR2 (N3436, N3427, N240);
or OR3 (N3437, N3424, N485, N2084);
xor XOR2 (N3438, N3436, N1688);
nor NOR2 (N3439, N3435, N2419);
not NOT1 (N3440, N3426);
xor XOR2 (N3441, N3437, N1127);
not NOT1 (N3442, N3429);
xor XOR2 (N3443, N3433, N1779);
xor XOR2 (N3444, N3442, N2576);
nor NOR2 (N3445, N3412, N2134);
or OR3 (N3446, N3443, N2562, N2477);
xor XOR2 (N3447, N3446, N1359);
not NOT1 (N3448, N3438);
nand NAND4 (N3449, N3440, N63, N1000, N2894);
nand NAND3 (N3450, N3448, N929, N17);
or OR4 (N3451, N3441, N1180, N219, N2643);
nand NAND3 (N3452, N3451, N3026, N2034);
buf BUF1 (N3453, N3447);
not NOT1 (N3454, N3445);
buf BUF1 (N3455, N3452);
and AND2 (N3456, N3430, N2005);
or OR4 (N3457, N3455, N2415, N2035, N2172);
xor XOR2 (N3458, N3419, N1925);
buf BUF1 (N3459, N3431);
buf BUF1 (N3460, N3439);
buf BUF1 (N3461, N3456);
not NOT1 (N3462, N3453);
nand NAND3 (N3463, N3457, N2155, N2751);
nor NOR2 (N3464, N3450, N3233);
not NOT1 (N3465, N3464);
and AND2 (N3466, N3449, N1122);
xor XOR2 (N3467, N3463, N3077);
and AND4 (N3468, N3444, N2205, N1871, N2104);
xor XOR2 (N3469, N3467, N1239);
nand NAND3 (N3470, N3460, N2431, N179);
nor NOR2 (N3471, N3459, N1028);
nor NOR2 (N3472, N3462, N199);
or OR2 (N3473, N3472, N604);
xor XOR2 (N3474, N3470, N3161);
or OR2 (N3475, N3458, N991);
and AND2 (N3476, N3465, N3223);
nand NAND3 (N3477, N3474, N1664, N944);
not NOT1 (N3478, N3476);
or OR2 (N3479, N3475, N2611);
or OR2 (N3480, N3461, N1663);
not NOT1 (N3481, N3473);
xor XOR2 (N3482, N3480, N3341);
nor NOR3 (N3483, N3471, N3408, N627);
nor NOR4 (N3484, N3477, N1751, N2897, N2670);
not NOT1 (N3485, N3482);
or OR2 (N3486, N3466, N2350);
not NOT1 (N3487, N3481);
or OR2 (N3488, N3469, N3246);
nor NOR2 (N3489, N3468, N683);
buf BUF1 (N3490, N3485);
not NOT1 (N3491, N3484);
and AND2 (N3492, N3488, N2507);
and AND3 (N3493, N3479, N3328, N424);
not NOT1 (N3494, N3487);
nand NAND2 (N3495, N3489, N1618);
or OR3 (N3496, N3491, N2242, N3384);
and AND3 (N3497, N3492, N295, N1844);
not NOT1 (N3498, N3496);
nor NOR3 (N3499, N3495, N3107, N2453);
xor XOR2 (N3500, N3478, N2358);
nand NAND3 (N3501, N3454, N2150, N1115);
or OR4 (N3502, N3486, N899, N2106, N718);
buf BUF1 (N3503, N3490);
or OR2 (N3504, N3500, N1724);
nor NOR4 (N3505, N3501, N749, N1128, N401);
buf BUF1 (N3506, N3503);
and AND4 (N3507, N3483, N1358, N167, N313);
nor NOR3 (N3508, N3507, N224, N2273);
nand NAND2 (N3509, N3504, N1065);
xor XOR2 (N3510, N3509, N2721);
or OR4 (N3511, N3497, N2133, N1425, N784);
xor XOR2 (N3512, N3506, N1679);
buf BUF1 (N3513, N3510);
buf BUF1 (N3514, N3513);
nor NOR3 (N3515, N3493, N1988, N3034);
not NOT1 (N3516, N3494);
not NOT1 (N3517, N3511);
buf BUF1 (N3518, N3498);
or OR3 (N3519, N3518, N2896, N655);
nand NAND3 (N3520, N3502, N3219, N3128);
nand NAND2 (N3521, N3516, N2585);
buf BUF1 (N3522, N3512);
not NOT1 (N3523, N3517);
and AND2 (N3524, N3520, N2026);
nand NAND4 (N3525, N3515, N565, N2677, N1410);
and AND3 (N3526, N3519, N3007, N1984);
xor XOR2 (N3527, N3523, N2765);
nor NOR3 (N3528, N3526, N1298, N1873);
not NOT1 (N3529, N3521);
or OR2 (N3530, N3514, N2298);
buf BUF1 (N3531, N3499);
nand NAND2 (N3532, N3528, N1612);
and AND2 (N3533, N3532, N678);
and AND3 (N3534, N3530, N108, N1908);
buf BUF1 (N3535, N3527);
buf BUF1 (N3536, N3524);
and AND2 (N3537, N3531, N2688);
buf BUF1 (N3538, N3505);
and AND2 (N3539, N3538, N2444);
or OR4 (N3540, N3508, N652, N2467, N2149);
buf BUF1 (N3541, N3535);
nand NAND2 (N3542, N3537, N2624);
or OR2 (N3543, N3539, N199);
nand NAND2 (N3544, N3522, N504);
nand NAND2 (N3545, N3542, N307);
buf BUF1 (N3546, N3541);
not NOT1 (N3547, N3546);
and AND3 (N3548, N3533, N354, N567);
and AND2 (N3549, N3525, N2402);
or OR4 (N3550, N3549, N2822, N1445, N380);
xor XOR2 (N3551, N3540, N3150);
nand NAND2 (N3552, N3543, N696);
nand NAND4 (N3553, N3545, N1227, N1814, N1421);
xor XOR2 (N3554, N3548, N2323);
xor XOR2 (N3555, N3551, N3437);
xor XOR2 (N3556, N3547, N1476);
or OR2 (N3557, N3550, N1393);
and AND3 (N3558, N3557, N808, N1221);
or OR2 (N3559, N3552, N2477);
or OR2 (N3560, N3559, N1451);
not NOT1 (N3561, N3558);
xor XOR2 (N3562, N3553, N1087);
and AND2 (N3563, N3554, N1300);
buf BUF1 (N3564, N3563);
or OR2 (N3565, N3536, N2793);
buf BUF1 (N3566, N3556);
xor XOR2 (N3567, N3564, N1379);
and AND3 (N3568, N3555, N2346, N491);
nor NOR2 (N3569, N3566, N656);
buf BUF1 (N3570, N3569);
nor NOR3 (N3571, N3544, N721, N630);
and AND3 (N3572, N3534, N1802, N1941);
xor XOR2 (N3573, N3570, N3493);
nor NOR4 (N3574, N3560, N1827, N768, N67);
and AND4 (N3575, N3574, N3405, N3218, N309);
xor XOR2 (N3576, N3572, N89);
or OR2 (N3577, N3567, N2312);
nor NOR3 (N3578, N3562, N2189, N3030);
buf BUF1 (N3579, N3575);
xor XOR2 (N3580, N3579, N1717);
xor XOR2 (N3581, N3573, N386);
nand NAND2 (N3582, N3568, N3105);
and AND3 (N3583, N3565, N968, N378);
or OR3 (N3584, N3529, N472, N473);
buf BUF1 (N3585, N3583);
or OR4 (N3586, N3584, N3225, N3527, N74);
buf BUF1 (N3587, N3561);
nor NOR2 (N3588, N3582, N1861);
or OR2 (N3589, N3571, N238);
nor NOR4 (N3590, N3581, N3073, N1694, N2605);
or OR2 (N3591, N3589, N518);
buf BUF1 (N3592, N3585);
buf BUF1 (N3593, N3577);
nand NAND3 (N3594, N3588, N518, N797);
and AND3 (N3595, N3594, N2278, N1970);
or OR3 (N3596, N3593, N1295, N548);
nor NOR3 (N3597, N3578, N3497, N2692);
or OR4 (N3598, N3576, N1692, N333, N2444);
or OR3 (N3599, N3591, N2810, N868);
or OR4 (N3600, N3597, N724, N1286, N150);
not NOT1 (N3601, N3599);
not NOT1 (N3602, N3587);
not NOT1 (N3603, N3598);
nand NAND3 (N3604, N3592, N711, N3029);
buf BUF1 (N3605, N3590);
nand NAND3 (N3606, N3596, N3462, N2666);
nor NOR3 (N3607, N3601, N1405, N1456);
nor NOR2 (N3608, N3586, N1777);
buf BUF1 (N3609, N3600);
or OR4 (N3610, N3609, N785, N2533, N1983);
xor XOR2 (N3611, N3595, N520);
xor XOR2 (N3612, N3604, N449);
or OR4 (N3613, N3605, N1300, N2330, N2448);
not NOT1 (N3614, N3603);
xor XOR2 (N3615, N3611, N2902);
nor NOR3 (N3616, N3602, N130, N1738);
nand NAND2 (N3617, N3610, N2246);
or OR3 (N3618, N3613, N2098, N3230);
and AND2 (N3619, N3606, N2512);
buf BUF1 (N3620, N3607);
nand NAND4 (N3621, N3617, N1953, N2888, N118);
not NOT1 (N3622, N3619);
not NOT1 (N3623, N3608);
nand NAND2 (N3624, N3623, N3303);
or OR2 (N3625, N3580, N1948);
buf BUF1 (N3626, N3622);
and AND2 (N3627, N3612, N337);
nor NOR2 (N3628, N3625, N1956);
buf BUF1 (N3629, N3616);
nand NAND3 (N3630, N3624, N1428, N1056);
or OR4 (N3631, N3628, N1849, N1895, N2278);
xor XOR2 (N3632, N3614, N423);
buf BUF1 (N3633, N3627);
or OR3 (N3634, N3633, N2335, N153);
nand NAND2 (N3635, N3629, N1647);
xor XOR2 (N3636, N3634, N2240);
and AND2 (N3637, N3626, N2126);
nand NAND2 (N3638, N3635, N3596);
or OR2 (N3639, N3618, N2741);
buf BUF1 (N3640, N3639);
nand NAND2 (N3641, N3621, N1275);
buf BUF1 (N3642, N3641);
or OR4 (N3643, N3640, N3461, N3448, N2784);
buf BUF1 (N3644, N3638);
buf BUF1 (N3645, N3620);
buf BUF1 (N3646, N3632);
buf BUF1 (N3647, N3644);
buf BUF1 (N3648, N3631);
nor NOR2 (N3649, N3637, N3061);
or OR2 (N3650, N3649, N2542);
buf BUF1 (N3651, N3636);
not NOT1 (N3652, N3647);
and AND2 (N3653, N3646, N595);
xor XOR2 (N3654, N3650, N3118);
or OR4 (N3655, N3651, N3632, N3481, N1162);
and AND4 (N3656, N3655, N462, N3080, N147);
buf BUF1 (N3657, N3656);
buf BUF1 (N3658, N3648);
and AND4 (N3659, N3653, N2953, N1442, N2700);
nor NOR3 (N3660, N3643, N1366, N2018);
not NOT1 (N3661, N3645);
nor NOR2 (N3662, N3661, N2586);
nand NAND2 (N3663, N3658, N508);
buf BUF1 (N3664, N3657);
nand NAND3 (N3665, N3654, N171, N485);
or OR2 (N3666, N3660, N1800);
buf BUF1 (N3667, N3662);
nand NAND2 (N3668, N3667, N2355);
or OR2 (N3669, N3664, N1700);
not NOT1 (N3670, N3642);
nor NOR3 (N3671, N3663, N72, N879);
and AND3 (N3672, N3669, N2532, N1377);
xor XOR2 (N3673, N3630, N3158);
not NOT1 (N3674, N3672);
or OR4 (N3675, N3670, N1647, N2924, N17);
xor XOR2 (N3676, N3673, N2408);
and AND4 (N3677, N3659, N294, N188, N3628);
or OR2 (N3678, N3615, N1869);
xor XOR2 (N3679, N3677, N2484);
and AND2 (N3680, N3666, N3241);
buf BUF1 (N3681, N3674);
nor NOR2 (N3682, N3671, N1906);
not NOT1 (N3683, N3681);
xor XOR2 (N3684, N3679, N1278);
not NOT1 (N3685, N3675);
buf BUF1 (N3686, N3678);
buf BUF1 (N3687, N3684);
or OR2 (N3688, N3683, N88);
and AND3 (N3689, N3676, N3059, N1171);
xor XOR2 (N3690, N3682, N409);
or OR2 (N3691, N3690, N3644);
xor XOR2 (N3692, N3665, N557);
xor XOR2 (N3693, N3686, N708);
nor NOR2 (N3694, N3668, N563);
and AND3 (N3695, N3687, N1148, N2904);
or OR4 (N3696, N3688, N700, N27, N2492);
or OR2 (N3697, N3692, N485);
buf BUF1 (N3698, N3685);
nand NAND4 (N3699, N3652, N2180, N2629, N2354);
xor XOR2 (N3700, N3693, N1138);
and AND3 (N3701, N3694, N1225, N1143);
not NOT1 (N3702, N3700);
nor NOR2 (N3703, N3698, N9);
buf BUF1 (N3704, N3703);
buf BUF1 (N3705, N3680);
buf BUF1 (N3706, N3696);
xor XOR2 (N3707, N3706, N3178);
and AND2 (N3708, N3702, N475);
or OR4 (N3709, N3707, N3099, N2328, N2225);
buf BUF1 (N3710, N3699);
xor XOR2 (N3711, N3701, N11);
nand NAND4 (N3712, N3691, N1563, N127, N107);
or OR4 (N3713, N3705, N1552, N961, N2405);
not NOT1 (N3714, N3709);
or OR2 (N3715, N3713, N225);
not NOT1 (N3716, N3712);
xor XOR2 (N3717, N3711, N2682);
nor NOR2 (N3718, N3715, N1220);
or OR3 (N3719, N3716, N2348, N1365);
not NOT1 (N3720, N3717);
xor XOR2 (N3721, N3708, N919);
xor XOR2 (N3722, N3714, N2175);
nor NOR4 (N3723, N3720, N2612, N750, N1084);
nand NAND3 (N3724, N3723, N3094, N2922);
and AND3 (N3725, N3722, N1664, N955);
nand NAND4 (N3726, N3704, N1101, N1984, N744);
xor XOR2 (N3727, N3689, N3674);
xor XOR2 (N3728, N3726, N3633);
and AND4 (N3729, N3727, N3715, N63, N641);
nand NAND2 (N3730, N3725, N2206);
nand NAND4 (N3731, N3724, N1704, N336, N1111);
nor NOR3 (N3732, N3718, N1053, N2749);
nor NOR3 (N3733, N3731, N275, N2683);
not NOT1 (N3734, N3710);
or OR4 (N3735, N3734, N3345, N459, N3362);
and AND3 (N3736, N3733, N237, N2779);
not NOT1 (N3737, N3730);
xor XOR2 (N3738, N3719, N1653);
xor XOR2 (N3739, N3738, N1465);
and AND4 (N3740, N3732, N1894, N1299, N988);
buf BUF1 (N3741, N3721);
nor NOR3 (N3742, N3737, N2231, N1801);
or OR4 (N3743, N3736, N233, N3589, N2753);
buf BUF1 (N3744, N3695);
xor XOR2 (N3745, N3735, N2863);
xor XOR2 (N3746, N3697, N725);
or OR4 (N3747, N3729, N752, N2076, N163);
nor NOR3 (N3748, N3744, N500, N3729);
or OR2 (N3749, N3739, N2813);
nand NAND4 (N3750, N3741, N2585, N352, N1693);
xor XOR2 (N3751, N3750, N3597);
nand NAND3 (N3752, N3740, N669, N845);
xor XOR2 (N3753, N3748, N1535);
buf BUF1 (N3754, N3749);
or OR2 (N3755, N3754, N1188);
and AND3 (N3756, N3745, N29, N2936);
buf BUF1 (N3757, N3753);
buf BUF1 (N3758, N3743);
xor XOR2 (N3759, N3742, N1879);
xor XOR2 (N3760, N3757, N3626);
not NOT1 (N3761, N3751);
nor NOR2 (N3762, N3746, N2523);
not NOT1 (N3763, N3762);
or OR3 (N3764, N3756, N974, N1820);
buf BUF1 (N3765, N3728);
not NOT1 (N3766, N3760);
nand NAND2 (N3767, N3766, N1228);
or OR4 (N3768, N3765, N3745, N987, N1445);
xor XOR2 (N3769, N3755, N2583);
buf BUF1 (N3770, N3747);
nand NAND3 (N3771, N3767, N1877, N1842);
nor NOR2 (N3772, N3763, N864);
or OR3 (N3773, N3758, N908, N1553);
buf BUF1 (N3774, N3771);
buf BUF1 (N3775, N3768);
nor NOR3 (N3776, N3772, N2508, N1222);
nor NOR2 (N3777, N3769, N1696);
or OR2 (N3778, N3776, N328);
or OR2 (N3779, N3774, N2772);
buf BUF1 (N3780, N3777);
not NOT1 (N3781, N3773);
xor XOR2 (N3782, N3778, N1926);
nor NOR2 (N3783, N3775, N2883);
buf BUF1 (N3784, N3752);
or OR4 (N3785, N3783, N1513, N2431, N1097);
and AND3 (N3786, N3782, N1710, N1598);
and AND3 (N3787, N3786, N785, N2017);
buf BUF1 (N3788, N3764);
xor XOR2 (N3789, N3761, N330);
not NOT1 (N3790, N3770);
xor XOR2 (N3791, N3789, N3520);
nor NOR3 (N3792, N3787, N2929, N2520);
buf BUF1 (N3793, N3784);
buf BUF1 (N3794, N3792);
nand NAND4 (N3795, N3794, N3608, N938, N1910);
not NOT1 (N3796, N3795);
or OR2 (N3797, N3780, N2552);
nand NAND4 (N3798, N3790, N586, N1701, N3582);
nand NAND2 (N3799, N3796, N1443);
buf BUF1 (N3800, N3785);
not NOT1 (N3801, N3797);
xor XOR2 (N3802, N3798, N1377);
nand NAND3 (N3803, N3793, N452, N2573);
xor XOR2 (N3804, N3788, N3096);
nor NOR3 (N3805, N3759, N747, N3593);
buf BUF1 (N3806, N3799);
and AND3 (N3807, N3801, N1723, N463);
nor NOR3 (N3808, N3804, N1386, N111);
or OR4 (N3809, N3803, N860, N342, N3012);
buf BUF1 (N3810, N3802);
not NOT1 (N3811, N3809);
buf BUF1 (N3812, N3791);
xor XOR2 (N3813, N3810, N3498);
xor XOR2 (N3814, N3808, N1767);
buf BUF1 (N3815, N3779);
not NOT1 (N3816, N3781);
buf BUF1 (N3817, N3812);
nor NOR3 (N3818, N3800, N1822, N2153);
buf BUF1 (N3819, N3805);
and AND2 (N3820, N3806, N1285);
nand NAND3 (N3821, N3817, N3067, N2197);
xor XOR2 (N3822, N3821, N1296);
xor XOR2 (N3823, N3814, N1819);
nand NAND2 (N3824, N3819, N2112);
not NOT1 (N3825, N3820);
buf BUF1 (N3826, N3815);
buf BUF1 (N3827, N3813);
or OR3 (N3828, N3825, N1000, N620);
and AND4 (N3829, N3828, N455, N2795, N3171);
or OR3 (N3830, N3807, N1336, N1333);
xor XOR2 (N3831, N3822, N2205);
xor XOR2 (N3832, N3826, N3476);
buf BUF1 (N3833, N3811);
nor NOR4 (N3834, N3823, N1368, N2855, N3771);
nand NAND3 (N3835, N3830, N1846, N782);
nor NOR3 (N3836, N3829, N541, N634);
nand NAND2 (N3837, N3834, N2085);
or OR4 (N3838, N3832, N3683, N1989, N2531);
buf BUF1 (N3839, N3837);
not NOT1 (N3840, N3827);
nand NAND3 (N3841, N3824, N2887, N3800);
xor XOR2 (N3842, N3841, N80);
not NOT1 (N3843, N3842);
nand NAND4 (N3844, N3836, N56, N1561, N1963);
not NOT1 (N3845, N3816);
xor XOR2 (N3846, N3835, N801);
or OR4 (N3847, N3840, N711, N3129, N1486);
xor XOR2 (N3848, N3839, N2333);
or OR3 (N3849, N3844, N533, N2187);
nor NOR3 (N3850, N3849, N427, N1878);
xor XOR2 (N3851, N3848, N49);
and AND2 (N3852, N3845, N1517);
nand NAND3 (N3853, N3847, N7, N273);
nor NOR4 (N3854, N3851, N2413, N1575, N543);
nand NAND4 (N3855, N3818, N1660, N2088, N2029);
xor XOR2 (N3856, N3855, N2600);
buf BUF1 (N3857, N3843);
nor NOR4 (N3858, N3857, N734, N1678, N2173);
not NOT1 (N3859, N3846);
and AND3 (N3860, N3859, N1878, N1036);
and AND3 (N3861, N3850, N1008, N218);
and AND3 (N3862, N3853, N2997, N97);
and AND4 (N3863, N3861, N2711, N3518, N151);
not NOT1 (N3864, N3863);
or OR3 (N3865, N3864, N977, N2410);
buf BUF1 (N3866, N3858);
and AND3 (N3867, N3866, N2761, N157);
nor NOR4 (N3868, N3831, N955, N108, N2795);
xor XOR2 (N3869, N3865, N1830);
nand NAND2 (N3870, N3852, N2310);
or OR3 (N3871, N3838, N1291, N2304);
not NOT1 (N3872, N3854);
not NOT1 (N3873, N3860);
buf BUF1 (N3874, N3862);
xor XOR2 (N3875, N3856, N2356);
nor NOR4 (N3876, N3833, N218, N2790, N1089);
nor NOR2 (N3877, N3868, N2813);
not NOT1 (N3878, N3875);
nand NAND3 (N3879, N3871, N2646, N825);
not NOT1 (N3880, N3878);
nand NAND3 (N3881, N3867, N1791, N1258);
xor XOR2 (N3882, N3881, N3488);
and AND4 (N3883, N3869, N3683, N130, N3780);
nor NOR2 (N3884, N3873, N2663);
and AND3 (N3885, N3884, N1854, N3744);
nand NAND3 (N3886, N3880, N3073, N2740);
buf BUF1 (N3887, N3883);
and AND2 (N3888, N3876, N496);
not NOT1 (N3889, N3885);
nand NAND3 (N3890, N3886, N2272, N3660);
nor NOR2 (N3891, N3882, N1346);
or OR2 (N3892, N3891, N2954);
buf BUF1 (N3893, N3889);
buf BUF1 (N3894, N3887);
buf BUF1 (N3895, N3874);
nand NAND4 (N3896, N3895, N3024, N139, N948);
nor NOR3 (N3897, N3870, N3417, N1066);
nand NAND2 (N3898, N3896, N3190);
not NOT1 (N3899, N3890);
xor XOR2 (N3900, N3888, N2631);
xor XOR2 (N3901, N3892, N2198);
or OR3 (N3902, N3872, N2688, N3619);
not NOT1 (N3903, N3893);
not NOT1 (N3904, N3897);
or OR2 (N3905, N3899, N1080);
not NOT1 (N3906, N3879);
nand NAND2 (N3907, N3904, N1049);
nand NAND3 (N3908, N3898, N1376, N2240);
nand NAND2 (N3909, N3894, N2629);
not NOT1 (N3910, N3907);
nor NOR4 (N3911, N3900, N30, N3284, N2971);
or OR2 (N3912, N3909, N3140);
not NOT1 (N3913, N3912);
nand NAND4 (N3914, N3906, N3338, N469, N2693);
xor XOR2 (N3915, N3903, N3033);
not NOT1 (N3916, N3905);
or OR2 (N3917, N3916, N3696);
nand NAND2 (N3918, N3902, N1526);
xor XOR2 (N3919, N3877, N2087);
nor NOR4 (N3920, N3919, N1652, N3136, N3900);
buf BUF1 (N3921, N3920);
not NOT1 (N3922, N3915);
nor NOR4 (N3923, N3914, N941, N185, N3651);
nor NOR2 (N3924, N3908, N3314);
nand NAND2 (N3925, N3901, N666);
not NOT1 (N3926, N3910);
or OR3 (N3927, N3924, N2314, N1336);
xor XOR2 (N3928, N3927, N895);
not NOT1 (N3929, N3926);
and AND3 (N3930, N3922, N951, N424);
or OR2 (N3931, N3928, N1854);
nor NOR2 (N3932, N3931, N2469);
or OR2 (N3933, N3929, N2805);
not NOT1 (N3934, N3933);
xor XOR2 (N3935, N3911, N2662);
and AND3 (N3936, N3921, N3079, N2194);
or OR4 (N3937, N3936, N1006, N33, N3701);
nand NAND2 (N3938, N3935, N2914);
and AND4 (N3939, N3932, N3794, N2523, N822);
or OR4 (N3940, N3937, N3812, N479, N3351);
nor NOR2 (N3941, N3925, N2589);
and AND3 (N3942, N3940, N2434, N832);
not NOT1 (N3943, N3918);
xor XOR2 (N3944, N3941, N3420);
nand NAND4 (N3945, N3934, N2111, N1972, N2468);
nor NOR4 (N3946, N3944, N3915, N2808, N1029);
or OR3 (N3947, N3923, N930, N497);
or OR3 (N3948, N3947, N3083, N2802);
and AND2 (N3949, N3942, N2267);
and AND2 (N3950, N3913, N1059);
or OR3 (N3951, N3943, N1359, N1997);
buf BUF1 (N3952, N3945);
buf BUF1 (N3953, N3949);
or OR4 (N3954, N3950, N3373, N1506, N773);
and AND2 (N3955, N3917, N115);
buf BUF1 (N3956, N3939);
not NOT1 (N3957, N3952);
nand NAND2 (N3958, N3957, N3693);
and AND4 (N3959, N3948, N2832, N3708, N2982);
xor XOR2 (N3960, N3938, N1269);
nor NOR3 (N3961, N3958, N974, N3730);
xor XOR2 (N3962, N3961, N2780);
buf BUF1 (N3963, N3960);
xor XOR2 (N3964, N3955, N2770);
nor NOR2 (N3965, N3954, N1633);
nand NAND2 (N3966, N3964, N2779);
not NOT1 (N3967, N3951);
or OR3 (N3968, N3956, N2103, N3467);
buf BUF1 (N3969, N3963);
not NOT1 (N3970, N3966);
or OR4 (N3971, N3967, N3534, N1977, N712);
or OR2 (N3972, N3968, N3837);
and AND3 (N3973, N3970, N1725, N2952);
or OR3 (N3974, N3953, N3878, N3442);
nor NOR4 (N3975, N3962, N1709, N227, N272);
buf BUF1 (N3976, N3973);
nand NAND2 (N3977, N3965, N1050);
nor NOR4 (N3978, N3974, N2530, N420, N3060);
xor XOR2 (N3979, N3976, N2769);
or OR4 (N3980, N3946, N1536, N1589, N929);
nor NOR4 (N3981, N3930, N315, N3454, N1056);
nand NAND2 (N3982, N3959, N3585);
buf BUF1 (N3983, N3978);
or OR3 (N3984, N3972, N3848, N3682);
not NOT1 (N3985, N3982);
buf BUF1 (N3986, N3975);
or OR2 (N3987, N3969, N3759);
or OR3 (N3988, N3971, N2852, N1467);
or OR3 (N3989, N3988, N2236, N2800);
nor NOR2 (N3990, N3987, N2643);
or OR2 (N3991, N3980, N464);
and AND2 (N3992, N3985, N998);
nor NOR3 (N3993, N3989, N1894, N3250);
nor NOR3 (N3994, N3984, N2751, N1162);
nand NAND3 (N3995, N3986, N3191, N2331);
xor XOR2 (N3996, N3992, N1754);
and AND3 (N3997, N3981, N2601, N714);
and AND4 (N3998, N3991, N1716, N2429, N3691);
and AND4 (N3999, N3990, N3485, N1207, N605);
xor XOR2 (N4000, N3979, N2839);
buf BUF1 (N4001, N3995);
nand NAND4 (N4002, N4000, N3427, N2308, N3760);
buf BUF1 (N4003, N3998);
nor NOR3 (N4004, N3977, N2490, N1721);
buf BUF1 (N4005, N3983);
not NOT1 (N4006, N4004);
not NOT1 (N4007, N4001);
not NOT1 (N4008, N3993);
xor XOR2 (N4009, N3997, N3150);
or OR4 (N4010, N4005, N1852, N825, N866);
buf BUF1 (N4011, N4008);
and AND4 (N4012, N4002, N1381, N2327, N3658);
xor XOR2 (N4013, N4012, N2476);
not NOT1 (N4014, N4007);
nor NOR4 (N4015, N4003, N1491, N3597, N2553);
xor XOR2 (N4016, N4015, N1662);
nor NOR3 (N4017, N3996, N997, N1230);
and AND4 (N4018, N4016, N1493, N621, N2465);
and AND3 (N4019, N4013, N3199, N3677);
xor XOR2 (N4020, N3999, N1928);
or OR4 (N4021, N4020, N1601, N134, N1527);
endmodule