// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N3008,N2988,N3005,N2993,N3011,N3007,N3010,N2995,N2982,N3012;

not NOT1 (N13, N11);
or OR2 (N14, N9, N4);
nand NAND2 (N15, N9, N8);
buf BUF1 (N16, N14);
nand NAND4 (N17, N8, N12, N8, N13);
not NOT1 (N18, N6);
and AND4 (N19, N13, N15, N15, N7);
buf BUF1 (N20, N7);
not NOT1 (N21, N16);
nand NAND4 (N22, N17, N16, N7, N17);
or OR4 (N23, N14, N5, N9, N15);
and AND3 (N24, N2, N2, N17);
buf BUF1 (N25, N23);
buf BUF1 (N26, N23);
or OR3 (N27, N14, N16, N7);
nand NAND2 (N28, N10, N23);
or OR4 (N29, N28, N4, N26, N24);
buf BUF1 (N30, N7);
or OR4 (N31, N18, N26, N15, N17);
xor XOR2 (N32, N10, N25);
buf BUF1 (N33, N7);
or OR4 (N34, N33, N22, N8, N28);
xor XOR2 (N35, N34, N27);
xor XOR2 (N36, N2, N33);
nand NAND2 (N37, N36, N36);
buf BUF1 (N38, N36);
xor XOR2 (N39, N32, N24);
nor NOR3 (N40, N30, N2, N13);
and AND3 (N41, N31, N10, N8);
not NOT1 (N42, N35);
buf BUF1 (N43, N41);
nand NAND2 (N44, N20, N2);
buf BUF1 (N45, N29);
xor XOR2 (N46, N44, N21);
nor NOR2 (N47, N7, N32);
and AND4 (N48, N19, N15, N19, N15);
buf BUF1 (N49, N48);
or OR2 (N50, N45, N9);
and AND4 (N51, N47, N10, N24, N3);
not NOT1 (N52, N51);
not NOT1 (N53, N42);
and AND2 (N54, N53, N47);
xor XOR2 (N55, N50, N44);
or OR2 (N56, N54, N39);
buf BUF1 (N57, N7);
or OR4 (N58, N43, N14, N4, N27);
nand NAND3 (N59, N49, N30, N20);
not NOT1 (N60, N52);
nor NOR3 (N61, N38, N10, N41);
not NOT1 (N62, N46);
xor XOR2 (N63, N62, N52);
or OR4 (N64, N37, N30, N25, N63);
buf BUF1 (N65, N41);
and AND3 (N66, N65, N53, N27);
and AND4 (N67, N55, N54, N12, N17);
not NOT1 (N68, N66);
nand NAND4 (N69, N59, N7, N61, N66);
buf BUF1 (N70, N33);
and AND3 (N71, N69, N58, N38);
buf BUF1 (N72, N64);
and AND4 (N73, N62, N11, N3, N25);
not NOT1 (N74, N70);
or OR4 (N75, N72, N6, N68, N61);
nand NAND4 (N76, N21, N62, N62, N10);
nand NAND2 (N77, N60, N38);
xor XOR2 (N78, N73, N32);
xor XOR2 (N79, N56, N20);
not NOT1 (N80, N76);
nand NAND4 (N81, N75, N24, N13, N72);
or OR4 (N82, N80, N35, N55, N2);
and AND4 (N83, N40, N68, N42, N82);
or OR3 (N84, N76, N25, N82);
nor NOR4 (N85, N84, N59, N80, N40);
buf BUF1 (N86, N77);
xor XOR2 (N87, N83, N36);
or OR3 (N88, N85, N83, N12);
not NOT1 (N89, N67);
buf BUF1 (N90, N71);
nand NAND4 (N91, N86, N86, N57, N11);
xor XOR2 (N92, N77, N23);
not NOT1 (N93, N78);
buf BUF1 (N94, N91);
nor NOR2 (N95, N93, N77);
not NOT1 (N96, N95);
xor XOR2 (N97, N94, N77);
and AND2 (N98, N97, N40);
buf BUF1 (N99, N88);
not NOT1 (N100, N96);
buf BUF1 (N101, N89);
nand NAND4 (N102, N99, N7, N4, N72);
buf BUF1 (N103, N79);
buf BUF1 (N104, N103);
nand NAND4 (N105, N104, N44, N51, N27);
xor XOR2 (N106, N101, N100);
buf BUF1 (N107, N1);
nor NOR2 (N108, N107, N48);
buf BUF1 (N109, N105);
nand NAND2 (N110, N106, N20);
not NOT1 (N111, N110);
and AND4 (N112, N108, N62, N69, N105);
or OR3 (N113, N74, N87, N73);
nand NAND2 (N114, N52, N15);
nand NAND3 (N115, N81, N98, N31);
nand NAND2 (N116, N7, N79);
nor NOR4 (N117, N90, N80, N43, N17);
or OR4 (N118, N114, N95, N109, N93);
or OR4 (N119, N94, N30, N107, N81);
and AND4 (N120, N116, N102, N44, N13);
not NOT1 (N121, N21);
or OR2 (N122, N111, N9);
nand NAND4 (N123, N115, N7, N48, N83);
or OR4 (N124, N113, N19, N20, N62);
not NOT1 (N125, N92);
buf BUF1 (N126, N125);
nand NAND3 (N127, N122, N51, N51);
buf BUF1 (N128, N119);
nand NAND2 (N129, N112, N28);
or OR4 (N130, N129, N109, N59, N46);
buf BUF1 (N131, N121);
nand NAND4 (N132, N120, N37, N4, N31);
xor XOR2 (N133, N126, N74);
not NOT1 (N134, N133);
or OR4 (N135, N124, N5, N6, N5);
xor XOR2 (N136, N135, N5);
or OR4 (N137, N136, N72, N30, N24);
buf BUF1 (N138, N137);
buf BUF1 (N139, N128);
or OR3 (N140, N117, N112, N97);
buf BUF1 (N141, N130);
and AND3 (N142, N138, N107, N96);
buf BUF1 (N143, N127);
nor NOR4 (N144, N132, N113, N94, N9);
xor XOR2 (N145, N141, N48);
nand NAND4 (N146, N140, N55, N46, N105);
xor XOR2 (N147, N123, N45);
or OR3 (N148, N142, N40, N127);
buf BUF1 (N149, N145);
xor XOR2 (N150, N149, N118);
nand NAND4 (N151, N149, N6, N88, N144);
or OR2 (N152, N63, N128);
not NOT1 (N153, N131);
buf BUF1 (N154, N147);
and AND2 (N155, N146, N68);
and AND2 (N156, N151, N75);
not NOT1 (N157, N154);
nor NOR4 (N158, N153, N111, N120, N140);
xor XOR2 (N159, N139, N90);
and AND2 (N160, N159, N70);
buf BUF1 (N161, N152);
nor NOR4 (N162, N150, N141, N53, N1);
and AND3 (N163, N158, N16, N47);
nor NOR4 (N164, N162, N21, N160, N141);
xor XOR2 (N165, N153, N25);
or OR4 (N166, N163, N32, N23, N102);
buf BUF1 (N167, N166);
xor XOR2 (N168, N155, N65);
xor XOR2 (N169, N156, N69);
nor NOR3 (N170, N148, N131, N78);
buf BUF1 (N171, N165);
buf BUF1 (N172, N161);
and AND2 (N173, N164, N119);
buf BUF1 (N174, N171);
buf BUF1 (N175, N172);
nor NOR4 (N176, N169, N15, N91, N83);
buf BUF1 (N177, N167);
not NOT1 (N178, N170);
or OR2 (N179, N134, N160);
and AND3 (N180, N157, N78, N20);
nor NOR2 (N181, N168, N172);
buf BUF1 (N182, N173);
not NOT1 (N183, N178);
and AND2 (N184, N174, N79);
not NOT1 (N185, N175);
buf BUF1 (N186, N177);
or OR2 (N187, N176, N161);
buf BUF1 (N188, N184);
nand NAND4 (N189, N185, N163, N107, N179);
buf BUF1 (N190, N185);
xor XOR2 (N191, N183, N164);
or OR3 (N192, N182, N118, N170);
buf BUF1 (N193, N187);
and AND4 (N194, N181, N3, N37, N58);
nor NOR3 (N195, N188, N15, N134);
or OR4 (N196, N195, N8, N48, N186);
nor NOR2 (N197, N29, N74);
or OR3 (N198, N189, N183, N75);
and AND3 (N199, N180, N145, N198);
nor NOR2 (N200, N124, N124);
nor NOR4 (N201, N193, N163, N7, N26);
not NOT1 (N202, N190);
nor NOR4 (N203, N202, N55, N70, N157);
or OR4 (N204, N196, N15, N45, N143);
and AND4 (N205, N34, N5, N142, N130);
and AND2 (N206, N204, N149);
or OR2 (N207, N200, N22);
nor NOR2 (N208, N191, N93);
not NOT1 (N209, N203);
buf BUF1 (N210, N209);
nand NAND3 (N211, N201, N110, N95);
nand NAND4 (N212, N197, N113, N183, N109);
nand NAND3 (N213, N211, N173, N27);
or OR2 (N214, N192, N34);
not NOT1 (N215, N207);
not NOT1 (N216, N205);
or OR2 (N217, N194, N69);
not NOT1 (N218, N210);
not NOT1 (N219, N214);
not NOT1 (N220, N212);
xor XOR2 (N221, N217, N219);
nand NAND2 (N222, N61, N38);
not NOT1 (N223, N218);
nand NAND2 (N224, N220, N207);
nor NOR4 (N225, N208, N81, N164, N97);
and AND2 (N226, N225, N96);
nor NOR2 (N227, N206, N17);
or OR4 (N228, N222, N217, N220, N163);
and AND3 (N229, N224, N170, N186);
xor XOR2 (N230, N215, N147);
xor XOR2 (N231, N229, N207);
or OR4 (N232, N226, N68, N170, N145);
and AND4 (N233, N199, N113, N57, N96);
xor XOR2 (N234, N233, N157);
buf BUF1 (N235, N232);
nor NOR4 (N236, N221, N188, N52, N58);
and AND2 (N237, N234, N128);
or OR2 (N238, N216, N197);
nand NAND2 (N239, N213, N155);
xor XOR2 (N240, N239, N140);
nand NAND4 (N241, N240, N188, N156, N163);
and AND3 (N242, N235, N4, N146);
buf BUF1 (N243, N230);
xor XOR2 (N244, N223, N232);
buf BUF1 (N245, N238);
nor NOR4 (N246, N237, N204, N139, N230);
not NOT1 (N247, N227);
and AND3 (N248, N236, N21, N231);
xor XOR2 (N249, N32, N101);
not NOT1 (N250, N241);
nor NOR4 (N251, N246, N231, N16, N68);
xor XOR2 (N252, N242, N250);
buf BUF1 (N253, N76);
nand NAND2 (N254, N252, N133);
nand NAND2 (N255, N243, N100);
nand NAND3 (N256, N249, N171, N181);
xor XOR2 (N257, N256, N141);
buf BUF1 (N258, N247);
nand NAND4 (N259, N245, N184, N214, N206);
nor NOR3 (N260, N258, N84, N102);
nor NOR2 (N261, N257, N242);
buf BUF1 (N262, N228);
buf BUF1 (N263, N244);
xor XOR2 (N264, N260, N165);
nand NAND3 (N265, N263, N256, N240);
not NOT1 (N266, N262);
and AND3 (N267, N253, N148, N58);
and AND4 (N268, N265, N96, N146, N146);
or OR2 (N269, N261, N203);
nand NAND3 (N270, N248, N151, N33);
or OR3 (N271, N255, N186, N42);
and AND3 (N272, N270, N258, N6);
nand NAND4 (N273, N259, N90, N227, N242);
or OR2 (N274, N268, N68);
xor XOR2 (N275, N251, N250);
and AND3 (N276, N275, N222, N150);
not NOT1 (N277, N269);
not NOT1 (N278, N274);
nand NAND4 (N279, N254, N48, N66, N189);
nor NOR4 (N280, N273, N192, N3, N121);
or OR3 (N281, N277, N210, N21);
xor XOR2 (N282, N279, N150);
and AND3 (N283, N264, N127, N132);
xor XOR2 (N284, N282, N263);
buf BUF1 (N285, N267);
xor XOR2 (N286, N280, N145);
buf BUF1 (N287, N276);
not NOT1 (N288, N284);
xor XOR2 (N289, N285, N92);
not NOT1 (N290, N281);
and AND3 (N291, N289, N190, N37);
nand NAND2 (N292, N291, N269);
nor NOR3 (N293, N283, N216, N216);
not NOT1 (N294, N271);
nand NAND2 (N295, N294, N205);
nor NOR3 (N296, N292, N167, N78);
nand NAND4 (N297, N278, N207, N212, N92);
nor NOR4 (N298, N297, N159, N138, N132);
not NOT1 (N299, N288);
or OR2 (N300, N293, N85);
xor XOR2 (N301, N295, N223);
and AND3 (N302, N272, N183, N124);
buf BUF1 (N303, N299);
xor XOR2 (N304, N290, N161);
or OR4 (N305, N298, N108, N285, N89);
not NOT1 (N306, N286);
and AND3 (N307, N266, N166, N10);
or OR4 (N308, N306, N43, N273, N203);
buf BUF1 (N309, N304);
not NOT1 (N310, N308);
nor NOR2 (N311, N305, N244);
or OR3 (N312, N300, N217, N270);
or OR4 (N313, N287, N244, N140, N94);
xor XOR2 (N314, N310, N91);
nand NAND4 (N315, N302, N247, N30, N221);
nand NAND2 (N316, N309, N233);
and AND3 (N317, N314, N303, N258);
or OR2 (N318, N74, N258);
or OR3 (N319, N311, N75, N262);
and AND2 (N320, N317, N98);
buf BUF1 (N321, N316);
nand NAND4 (N322, N321, N135, N168, N238);
or OR2 (N323, N319, N24);
not NOT1 (N324, N323);
nor NOR3 (N325, N318, N164, N42);
buf BUF1 (N326, N307);
and AND3 (N327, N301, N123, N279);
and AND3 (N328, N296, N166, N248);
nor NOR4 (N329, N320, N26, N103, N243);
xor XOR2 (N330, N324, N5);
and AND2 (N331, N327, N29);
xor XOR2 (N332, N328, N322);
nor NOR4 (N333, N55, N332, N307, N163);
nand NAND4 (N334, N333, N119, N127, N181);
not NOT1 (N335, N233);
nor NOR4 (N336, N325, N80, N189, N319);
nand NAND2 (N337, N335, N149);
and AND2 (N338, N331, N213);
nor NOR4 (N339, N336, N325, N198, N44);
nor NOR3 (N340, N334, N105, N248);
nand NAND3 (N341, N329, N107, N80);
buf BUF1 (N342, N313);
and AND2 (N343, N338, N206);
buf BUF1 (N344, N312);
buf BUF1 (N345, N330);
and AND3 (N346, N326, N85, N206);
nor NOR3 (N347, N344, N144, N112);
not NOT1 (N348, N343);
or OR3 (N349, N337, N182, N106);
not NOT1 (N350, N315);
and AND4 (N351, N345, N172, N329, N77);
or OR2 (N352, N347, N47);
not NOT1 (N353, N350);
nor NOR3 (N354, N340, N171, N165);
xor XOR2 (N355, N342, N287);
nand NAND2 (N356, N349, N232);
and AND2 (N357, N353, N93);
and AND4 (N358, N351, N195, N238, N178);
or OR3 (N359, N346, N255, N191);
and AND4 (N360, N339, N95, N110, N13);
nor NOR3 (N361, N348, N126, N325);
nand NAND4 (N362, N357, N208, N76, N271);
or OR3 (N363, N341, N63, N312);
xor XOR2 (N364, N363, N217);
nand NAND3 (N365, N355, N169, N79);
nand NAND3 (N366, N358, N266, N193);
and AND4 (N367, N366, N244, N279, N348);
xor XOR2 (N368, N356, N184);
or OR2 (N369, N365, N124);
and AND2 (N370, N360, N182);
not NOT1 (N371, N370);
and AND4 (N372, N369, N259, N88, N192);
nand NAND3 (N373, N354, N318, N50);
not NOT1 (N374, N359);
xor XOR2 (N375, N352, N324);
nand NAND2 (N376, N367, N303);
and AND4 (N377, N376, N317, N228, N133);
xor XOR2 (N378, N361, N121);
not NOT1 (N379, N375);
and AND2 (N380, N373, N56);
buf BUF1 (N381, N380);
xor XOR2 (N382, N362, N366);
or OR4 (N383, N364, N357, N321, N35);
not NOT1 (N384, N379);
xor XOR2 (N385, N378, N323);
nand NAND4 (N386, N371, N364, N116, N273);
nand NAND4 (N387, N377, N97, N168, N239);
xor XOR2 (N388, N384, N223);
xor XOR2 (N389, N385, N339);
and AND2 (N390, N383, N39);
not NOT1 (N391, N387);
buf BUF1 (N392, N372);
nand NAND2 (N393, N374, N357);
nand NAND3 (N394, N368, N393, N273);
buf BUF1 (N395, N163);
nor NOR3 (N396, N388, N23, N76);
or OR3 (N397, N389, N59, N128);
xor XOR2 (N398, N390, N44);
and AND3 (N399, N381, N266, N387);
nand NAND4 (N400, N392, N2, N268, N302);
nor NOR3 (N401, N398, N281, N271);
xor XOR2 (N402, N401, N257);
nor NOR4 (N403, N382, N253, N311, N258);
xor XOR2 (N404, N402, N275);
xor XOR2 (N405, N399, N245);
or OR2 (N406, N403, N132);
and AND4 (N407, N391, N78, N348, N66);
nand NAND3 (N408, N394, N383, N129);
buf BUF1 (N409, N397);
or OR2 (N410, N404, N276);
or OR3 (N411, N407, N242, N369);
or OR4 (N412, N411, N316, N335, N111);
xor XOR2 (N413, N405, N292);
buf BUF1 (N414, N409);
nand NAND2 (N415, N395, N231);
or OR4 (N416, N406, N249, N163, N138);
and AND2 (N417, N408, N7);
buf BUF1 (N418, N416);
buf BUF1 (N419, N396);
nor NOR2 (N420, N417, N109);
and AND3 (N421, N412, N110, N321);
xor XOR2 (N422, N410, N7);
buf BUF1 (N423, N422);
nand NAND3 (N424, N400, N228, N217);
nor NOR3 (N425, N386, N237, N365);
xor XOR2 (N426, N420, N79);
and AND2 (N427, N425, N5);
nand NAND3 (N428, N419, N68, N189);
nor NOR4 (N429, N424, N340, N34, N415);
buf BUF1 (N430, N276);
xor XOR2 (N431, N421, N10);
not NOT1 (N432, N414);
and AND4 (N433, N432, N203, N403, N14);
xor XOR2 (N434, N427, N261);
buf BUF1 (N435, N418);
not NOT1 (N436, N413);
buf BUF1 (N437, N430);
and AND2 (N438, N423, N54);
nand NAND2 (N439, N426, N306);
xor XOR2 (N440, N431, N345);
xor XOR2 (N441, N429, N137);
not NOT1 (N442, N436);
buf BUF1 (N443, N435);
or OR3 (N444, N428, N8, N412);
xor XOR2 (N445, N442, N100);
xor XOR2 (N446, N441, N344);
not NOT1 (N447, N445);
not NOT1 (N448, N447);
not NOT1 (N449, N438);
not NOT1 (N450, N449);
buf BUF1 (N451, N446);
not NOT1 (N452, N450);
and AND3 (N453, N437, N190, N299);
buf BUF1 (N454, N434);
or OR3 (N455, N452, N33, N301);
not NOT1 (N456, N451);
or OR4 (N457, N444, N104, N250, N259);
xor XOR2 (N458, N439, N394);
buf BUF1 (N459, N456);
xor XOR2 (N460, N443, N371);
buf BUF1 (N461, N457);
xor XOR2 (N462, N461, N157);
nor NOR3 (N463, N453, N98, N199);
buf BUF1 (N464, N459);
nor NOR3 (N465, N455, N26, N194);
nor NOR4 (N466, N463, N369, N75, N188);
not NOT1 (N467, N466);
and AND2 (N468, N448, N229);
xor XOR2 (N469, N460, N159);
not NOT1 (N470, N440);
or OR3 (N471, N462, N204, N252);
nor NOR2 (N472, N465, N328);
or OR3 (N473, N468, N142, N118);
or OR4 (N474, N454, N23, N15, N196);
and AND3 (N475, N473, N397, N8);
or OR4 (N476, N472, N402, N391, N128);
not NOT1 (N477, N475);
not NOT1 (N478, N477);
nand NAND2 (N479, N458, N133);
nand NAND2 (N480, N469, N22);
not NOT1 (N481, N479);
not NOT1 (N482, N478);
and AND2 (N483, N476, N282);
and AND3 (N484, N480, N226, N15);
not NOT1 (N485, N483);
and AND3 (N486, N471, N45, N153);
or OR4 (N487, N482, N403, N227, N444);
or OR2 (N488, N467, N74);
and AND3 (N489, N481, N409, N331);
buf BUF1 (N490, N464);
nand NAND4 (N491, N488, N270, N475, N370);
and AND4 (N492, N491, N183, N181, N288);
and AND3 (N493, N474, N16, N80);
xor XOR2 (N494, N489, N424);
not NOT1 (N495, N486);
or OR4 (N496, N490, N282, N390, N87);
or OR4 (N497, N470, N77, N168, N240);
xor XOR2 (N498, N496, N378);
nand NAND2 (N499, N494, N149);
and AND3 (N500, N485, N248, N357);
xor XOR2 (N501, N497, N485);
not NOT1 (N502, N433);
or OR4 (N503, N499, N10, N294, N341);
buf BUF1 (N504, N503);
nor NOR3 (N505, N498, N140, N123);
or OR3 (N506, N504, N484, N372);
nor NOR4 (N507, N498, N168, N221, N427);
not NOT1 (N508, N487);
nor NOR3 (N509, N505, N366, N456);
or OR3 (N510, N501, N257, N343);
buf BUF1 (N511, N495);
or OR2 (N512, N492, N129);
and AND3 (N513, N509, N179, N501);
not NOT1 (N514, N508);
and AND2 (N515, N512, N280);
buf BUF1 (N516, N507);
nand NAND4 (N517, N500, N393, N354, N360);
not NOT1 (N518, N493);
nand NAND3 (N519, N516, N448, N410);
and AND2 (N520, N515, N247);
nor NOR2 (N521, N518, N433);
and AND4 (N522, N506, N410, N29, N278);
xor XOR2 (N523, N520, N166);
nand NAND2 (N524, N513, N365);
not NOT1 (N525, N514);
not NOT1 (N526, N524);
or OR2 (N527, N510, N248);
nor NOR2 (N528, N523, N181);
buf BUF1 (N529, N525);
nand NAND4 (N530, N528, N400, N289, N17);
not NOT1 (N531, N522);
not NOT1 (N532, N511);
xor XOR2 (N533, N517, N147);
xor XOR2 (N534, N521, N427);
xor XOR2 (N535, N530, N303);
not NOT1 (N536, N526);
xor XOR2 (N537, N502, N501);
nand NAND4 (N538, N529, N417, N341, N485);
not NOT1 (N539, N532);
or OR4 (N540, N527, N295, N249, N112);
or OR4 (N541, N537, N290, N56, N102);
buf BUF1 (N542, N533);
nand NAND3 (N543, N536, N434, N374);
nand NAND4 (N544, N519, N486, N509, N100);
not NOT1 (N545, N534);
nor NOR2 (N546, N545, N481);
and AND4 (N547, N531, N92, N515, N62);
not NOT1 (N548, N543);
or OR3 (N549, N544, N161, N214);
buf BUF1 (N550, N540);
not NOT1 (N551, N539);
xor XOR2 (N552, N541, N115);
buf BUF1 (N553, N552);
not NOT1 (N554, N538);
or OR3 (N555, N546, N100, N34);
not NOT1 (N556, N542);
not NOT1 (N557, N556);
nor NOR4 (N558, N548, N374, N506, N276);
nor NOR2 (N559, N557, N360);
not NOT1 (N560, N551);
nand NAND3 (N561, N550, N31, N486);
or OR2 (N562, N560, N506);
xor XOR2 (N563, N549, N123);
xor XOR2 (N564, N561, N374);
and AND4 (N565, N558, N277, N193, N248);
nand NAND3 (N566, N559, N515, N51);
buf BUF1 (N567, N564);
or OR3 (N568, N562, N411, N518);
not NOT1 (N569, N554);
buf BUF1 (N570, N569);
xor XOR2 (N571, N563, N147);
xor XOR2 (N572, N565, N161);
not NOT1 (N573, N566);
xor XOR2 (N574, N568, N222);
nand NAND3 (N575, N553, N287, N309);
not NOT1 (N576, N574);
nor NOR2 (N577, N547, N168);
nor NOR4 (N578, N575, N217, N80, N461);
nand NAND3 (N579, N535, N156, N305);
xor XOR2 (N580, N578, N451);
not NOT1 (N581, N555);
and AND2 (N582, N579, N231);
nand NAND4 (N583, N572, N155, N456, N268);
nand NAND3 (N584, N583, N540, N516);
xor XOR2 (N585, N573, N229);
xor XOR2 (N586, N567, N490);
and AND3 (N587, N581, N343, N401);
not NOT1 (N588, N576);
not NOT1 (N589, N587);
xor XOR2 (N590, N586, N325);
nand NAND3 (N591, N577, N427, N541);
buf BUF1 (N592, N584);
nand NAND2 (N593, N585, N64);
and AND3 (N594, N571, N344, N289);
buf BUF1 (N595, N588);
buf BUF1 (N596, N594);
not NOT1 (N597, N580);
or OR4 (N598, N591, N389, N353, N1);
not NOT1 (N599, N582);
and AND3 (N600, N598, N518, N153);
or OR4 (N601, N600, N99, N18, N271);
and AND4 (N602, N599, N114, N111, N160);
or OR4 (N603, N602, N498, N53, N226);
or OR4 (N604, N589, N557, N466, N586);
not NOT1 (N605, N601);
and AND2 (N606, N596, N212);
not NOT1 (N607, N595);
not NOT1 (N608, N593);
or OR2 (N609, N597, N38);
not NOT1 (N610, N607);
nor NOR4 (N611, N592, N208, N108, N536);
nand NAND2 (N612, N570, N275);
not NOT1 (N613, N603);
not NOT1 (N614, N611);
nand NAND4 (N615, N604, N386, N368, N398);
not NOT1 (N616, N608);
or OR4 (N617, N612, N515, N229, N172);
and AND4 (N618, N590, N460, N6, N366);
not NOT1 (N619, N605);
nand NAND3 (N620, N615, N159, N496);
or OR4 (N621, N618, N238, N98, N86);
xor XOR2 (N622, N613, N114);
not NOT1 (N623, N621);
xor XOR2 (N624, N617, N282);
nor NOR4 (N625, N622, N289, N399, N22);
nand NAND3 (N626, N609, N125, N218);
not NOT1 (N627, N610);
nand NAND4 (N628, N625, N562, N425, N379);
or OR2 (N629, N624, N587);
buf BUF1 (N630, N620);
nor NOR4 (N631, N626, N560, N406, N451);
and AND3 (N632, N614, N384, N34);
buf BUF1 (N633, N623);
nor NOR3 (N634, N632, N519, N341);
nor NOR2 (N635, N630, N105);
nand NAND4 (N636, N627, N612, N297, N289);
nand NAND4 (N637, N631, N601, N166, N170);
nand NAND3 (N638, N633, N226, N70);
nand NAND3 (N639, N635, N549, N616);
not NOT1 (N640, N182);
nand NAND4 (N641, N639, N95, N294, N585);
not NOT1 (N642, N637);
buf BUF1 (N643, N634);
not NOT1 (N644, N636);
and AND2 (N645, N644, N75);
buf BUF1 (N646, N629);
xor XOR2 (N647, N640, N587);
not NOT1 (N648, N628);
or OR3 (N649, N606, N141, N489);
not NOT1 (N650, N648);
buf BUF1 (N651, N650);
nor NOR4 (N652, N619, N280, N36, N528);
buf BUF1 (N653, N647);
not NOT1 (N654, N642);
nor NOR3 (N655, N651, N76, N643);
and AND2 (N656, N497, N440);
buf BUF1 (N657, N654);
not NOT1 (N658, N653);
nor NOR3 (N659, N655, N379, N315);
xor XOR2 (N660, N638, N564);
buf BUF1 (N661, N649);
nand NAND3 (N662, N645, N572, N316);
nor NOR2 (N663, N658, N449);
nand NAND3 (N664, N657, N651, N218);
nor NOR3 (N665, N652, N88, N171);
nor NOR4 (N666, N661, N181, N422, N499);
xor XOR2 (N667, N656, N482);
xor XOR2 (N668, N641, N229);
and AND3 (N669, N668, N560, N411);
xor XOR2 (N670, N664, N342);
not NOT1 (N671, N667);
nand NAND2 (N672, N666, N19);
nor NOR4 (N673, N669, N179, N269, N132);
not NOT1 (N674, N672);
nor NOR3 (N675, N674, N353, N407);
nor NOR3 (N676, N663, N358, N520);
buf BUF1 (N677, N675);
xor XOR2 (N678, N676, N513);
nor NOR2 (N679, N659, N4);
or OR4 (N680, N665, N211, N467, N319);
and AND3 (N681, N670, N607, N315);
or OR4 (N682, N677, N669, N235, N52);
buf BUF1 (N683, N682);
nor NOR3 (N684, N679, N615, N35);
xor XOR2 (N685, N646, N170);
buf BUF1 (N686, N681);
nand NAND3 (N687, N673, N326, N46);
nor NOR2 (N688, N686, N112);
nor NOR3 (N689, N660, N626, N560);
buf BUF1 (N690, N662);
or OR3 (N691, N685, N426, N324);
or OR2 (N692, N691, N155);
or OR2 (N693, N684, N470);
xor XOR2 (N694, N671, N149);
and AND4 (N695, N693, N533, N607, N559);
and AND3 (N696, N695, N191, N497);
not NOT1 (N697, N694);
nand NAND2 (N698, N697, N337);
nand NAND2 (N699, N687, N643);
nor NOR3 (N700, N688, N502, N278);
not NOT1 (N701, N699);
or OR4 (N702, N689, N124, N293, N77);
nand NAND4 (N703, N702, N429, N225, N669);
and AND3 (N704, N700, N179, N692);
or OR3 (N705, N365, N462, N536);
xor XOR2 (N706, N701, N466);
or OR3 (N707, N690, N478, N664);
nor NOR4 (N708, N707, N583, N295, N464);
xor XOR2 (N709, N703, N5);
not NOT1 (N710, N683);
or OR4 (N711, N678, N513, N574, N188);
buf BUF1 (N712, N698);
nor NOR3 (N713, N710, N309, N409);
xor XOR2 (N714, N705, N36);
nand NAND4 (N715, N704, N614, N188, N404);
buf BUF1 (N716, N709);
and AND4 (N717, N715, N220, N128, N334);
nor NOR4 (N718, N716, N500, N392, N605);
and AND4 (N719, N717, N410, N176, N599);
xor XOR2 (N720, N706, N535);
xor XOR2 (N721, N713, N32);
xor XOR2 (N722, N712, N445);
not NOT1 (N723, N708);
and AND2 (N724, N723, N490);
nor NOR3 (N725, N721, N229, N18);
nor NOR4 (N726, N720, N461, N351, N254);
and AND3 (N727, N725, N195, N322);
buf BUF1 (N728, N719);
not NOT1 (N729, N722);
and AND4 (N730, N724, N664, N51, N571);
buf BUF1 (N731, N728);
buf BUF1 (N732, N711);
and AND3 (N733, N680, N340, N572);
not NOT1 (N734, N729);
buf BUF1 (N735, N727);
xor XOR2 (N736, N696, N114);
nor NOR3 (N737, N733, N11, N647);
nor NOR4 (N738, N737, N238, N146, N226);
nand NAND3 (N739, N731, N255, N659);
or OR3 (N740, N718, N267, N685);
and AND3 (N741, N738, N103, N236);
not NOT1 (N742, N741);
nand NAND4 (N743, N726, N385, N420, N446);
nand NAND3 (N744, N732, N144, N209);
nor NOR3 (N745, N742, N93, N619);
nand NAND4 (N746, N736, N572, N63, N605);
and AND3 (N747, N746, N227, N25);
nand NAND4 (N748, N735, N45, N104, N106);
or OR3 (N749, N748, N747, N588);
and AND2 (N750, N227, N95);
nor NOR2 (N751, N750, N510);
nand NAND2 (N752, N739, N11);
xor XOR2 (N753, N745, N521);
nand NAND4 (N754, N751, N205, N417, N653);
nand NAND4 (N755, N714, N190, N125, N27);
and AND3 (N756, N740, N57, N283);
nor NOR4 (N757, N754, N279, N219, N394);
not NOT1 (N758, N730);
nor NOR4 (N759, N756, N383, N67, N552);
not NOT1 (N760, N734);
not NOT1 (N761, N759);
nand NAND4 (N762, N752, N362, N58, N23);
nand NAND3 (N763, N757, N365, N11);
nor NOR4 (N764, N758, N473, N168, N58);
nand NAND3 (N765, N749, N495, N733);
xor XOR2 (N766, N743, N131);
buf BUF1 (N767, N761);
not NOT1 (N768, N767);
nor NOR3 (N769, N744, N548, N469);
or OR3 (N770, N762, N616, N343);
and AND4 (N771, N765, N721, N196, N525);
or OR3 (N772, N760, N594, N375);
nand NAND4 (N773, N764, N519, N379, N163);
and AND3 (N774, N763, N474, N715);
nor NOR3 (N775, N766, N464, N90);
or OR3 (N776, N772, N292, N443);
or OR4 (N777, N773, N98, N111, N748);
not NOT1 (N778, N775);
xor XOR2 (N779, N771, N673);
nor NOR3 (N780, N769, N725, N360);
and AND2 (N781, N770, N65);
buf BUF1 (N782, N755);
xor XOR2 (N783, N774, N294);
xor XOR2 (N784, N776, N197);
and AND2 (N785, N784, N69);
xor XOR2 (N786, N780, N315);
nand NAND4 (N787, N768, N227, N84, N739);
buf BUF1 (N788, N778);
nor NOR2 (N789, N783, N700);
or OR2 (N790, N785, N543);
or OR4 (N791, N789, N674, N537, N591);
or OR3 (N792, N753, N726, N97);
xor XOR2 (N793, N777, N202);
buf BUF1 (N794, N791);
nor NOR3 (N795, N782, N89, N707);
buf BUF1 (N796, N788);
or OR4 (N797, N790, N388, N62, N168);
or OR3 (N798, N779, N672, N161);
buf BUF1 (N799, N797);
and AND2 (N800, N796, N555);
and AND2 (N801, N799, N500);
xor XOR2 (N802, N794, N700);
nand NAND3 (N803, N787, N787, N34);
buf BUF1 (N804, N793);
and AND4 (N805, N798, N531, N166, N728);
buf BUF1 (N806, N805);
not NOT1 (N807, N802);
nor NOR3 (N808, N806, N445, N699);
nand NAND4 (N809, N781, N745, N16, N504);
and AND3 (N810, N807, N694, N170);
nand NAND4 (N811, N809, N675, N107, N100);
nor NOR3 (N812, N786, N762, N609);
and AND3 (N813, N810, N781, N299);
nand NAND3 (N814, N812, N61, N31);
and AND2 (N815, N808, N254);
nand NAND4 (N816, N804, N87, N469, N523);
or OR2 (N817, N795, N199);
not NOT1 (N818, N815);
not NOT1 (N819, N817);
or OR4 (N820, N818, N214, N800, N67);
nor NOR4 (N821, N258, N19, N282, N592);
not NOT1 (N822, N813);
nor NOR3 (N823, N811, N31, N228);
or OR3 (N824, N801, N285, N125);
nor NOR4 (N825, N822, N419, N522, N529);
or OR3 (N826, N825, N118, N793);
nand NAND4 (N827, N820, N535, N454, N770);
buf BUF1 (N828, N821);
buf BUF1 (N829, N827);
buf BUF1 (N830, N816);
buf BUF1 (N831, N819);
nand NAND3 (N832, N829, N716, N265);
or OR3 (N833, N803, N377, N645);
nand NAND2 (N834, N833, N18);
xor XOR2 (N835, N831, N92);
nor NOR2 (N836, N824, N294);
not NOT1 (N837, N834);
nor NOR3 (N838, N828, N499, N287);
buf BUF1 (N839, N823);
xor XOR2 (N840, N814, N757);
buf BUF1 (N841, N838);
or OR2 (N842, N839, N649);
nor NOR3 (N843, N835, N385, N226);
or OR2 (N844, N826, N647);
nor NOR3 (N845, N830, N558, N781);
xor XOR2 (N846, N844, N180);
or OR3 (N847, N846, N497, N353);
nand NAND3 (N848, N792, N310, N520);
nand NAND2 (N849, N836, N97);
buf BUF1 (N850, N845);
not NOT1 (N851, N843);
nor NOR4 (N852, N851, N170, N43, N767);
or OR2 (N853, N832, N760);
or OR4 (N854, N848, N608, N279, N851);
not NOT1 (N855, N850);
buf BUF1 (N856, N852);
not NOT1 (N857, N837);
or OR2 (N858, N847, N462);
xor XOR2 (N859, N855, N505);
or OR3 (N860, N841, N763, N245);
buf BUF1 (N861, N853);
not NOT1 (N862, N861);
nand NAND2 (N863, N857, N149);
nor NOR3 (N864, N862, N825, N567);
and AND4 (N865, N859, N184, N285, N519);
and AND2 (N866, N840, N140);
and AND2 (N867, N858, N758);
and AND2 (N868, N865, N362);
and AND3 (N869, N867, N405, N432);
nor NOR3 (N870, N842, N868, N21);
xor XOR2 (N871, N43, N77);
xor XOR2 (N872, N864, N564);
nand NAND3 (N873, N870, N426, N281);
not NOT1 (N874, N869);
not NOT1 (N875, N866);
buf BUF1 (N876, N872);
not NOT1 (N877, N860);
nand NAND4 (N878, N863, N226, N622, N90);
nor NOR2 (N879, N856, N424);
not NOT1 (N880, N875);
nand NAND2 (N881, N854, N299);
or OR4 (N882, N878, N462, N799, N195);
or OR4 (N883, N881, N627, N841, N44);
not NOT1 (N884, N880);
or OR3 (N885, N871, N704, N492);
xor XOR2 (N886, N849, N256);
or OR2 (N887, N882, N751);
xor XOR2 (N888, N873, N153);
nand NAND2 (N889, N885, N155);
nand NAND2 (N890, N888, N571);
buf BUF1 (N891, N890);
not NOT1 (N892, N879);
or OR2 (N893, N884, N352);
and AND2 (N894, N891, N220);
xor XOR2 (N895, N894, N809);
nand NAND2 (N896, N886, N349);
and AND2 (N897, N876, N327);
xor XOR2 (N898, N897, N507);
buf BUF1 (N899, N877);
nor NOR4 (N900, N896, N352, N804, N108);
not NOT1 (N901, N892);
or OR2 (N902, N895, N477);
xor XOR2 (N903, N902, N491);
not NOT1 (N904, N893);
nand NAND2 (N905, N900, N555);
and AND4 (N906, N889, N744, N453, N567);
buf BUF1 (N907, N899);
not NOT1 (N908, N906);
buf BUF1 (N909, N907);
nand NAND4 (N910, N909, N211, N9, N841);
and AND3 (N911, N903, N596, N559);
nand NAND3 (N912, N904, N332, N96);
xor XOR2 (N913, N883, N134);
and AND4 (N914, N908, N629, N218, N435);
xor XOR2 (N915, N912, N837);
and AND3 (N916, N911, N209, N294);
not NOT1 (N917, N916);
buf BUF1 (N918, N913);
not NOT1 (N919, N901);
or OR2 (N920, N905, N584);
buf BUF1 (N921, N917);
not NOT1 (N922, N898);
nand NAND4 (N923, N919, N867, N194, N260);
buf BUF1 (N924, N920);
or OR3 (N925, N874, N329, N102);
not NOT1 (N926, N925);
not NOT1 (N927, N910);
not NOT1 (N928, N921);
xor XOR2 (N929, N927, N677);
or OR2 (N930, N929, N605);
buf BUF1 (N931, N887);
buf BUF1 (N932, N914);
not NOT1 (N933, N924);
buf BUF1 (N934, N930);
nor NOR2 (N935, N934, N153);
or OR2 (N936, N926, N305);
not NOT1 (N937, N931);
buf BUF1 (N938, N935);
or OR4 (N939, N922, N937, N423, N185);
and AND3 (N940, N47, N432, N342);
and AND2 (N941, N918, N719);
or OR3 (N942, N932, N619, N241);
nand NAND3 (N943, N941, N182, N893);
nand NAND3 (N944, N933, N436, N332);
buf BUF1 (N945, N939);
not NOT1 (N946, N915);
and AND3 (N947, N944, N734, N744);
not NOT1 (N948, N943);
and AND3 (N949, N938, N850, N183);
nand NAND2 (N950, N923, N770);
or OR4 (N951, N942, N813, N741, N575);
buf BUF1 (N952, N946);
xor XOR2 (N953, N949, N735);
nor NOR3 (N954, N950, N875, N474);
nand NAND4 (N955, N948, N209, N551, N232);
nor NOR4 (N956, N928, N884, N385, N293);
not NOT1 (N957, N936);
nand NAND4 (N958, N956, N900, N135, N519);
xor XOR2 (N959, N955, N590);
xor XOR2 (N960, N951, N176);
xor XOR2 (N961, N940, N893);
or OR2 (N962, N953, N859);
nor NOR2 (N963, N945, N111);
xor XOR2 (N964, N959, N471);
nor NOR2 (N965, N963, N17);
or OR4 (N966, N964, N158, N540, N646);
or OR4 (N967, N954, N807, N586, N265);
buf BUF1 (N968, N966);
not NOT1 (N969, N947);
xor XOR2 (N970, N969, N422);
or OR3 (N971, N957, N829, N745);
xor XOR2 (N972, N952, N592);
xor XOR2 (N973, N962, N179);
xor XOR2 (N974, N960, N865);
buf BUF1 (N975, N972);
or OR2 (N976, N975, N545);
or OR2 (N977, N958, N397);
or OR3 (N978, N971, N460, N869);
or OR4 (N979, N961, N404, N556, N172);
nand NAND4 (N980, N970, N94, N257, N371);
not NOT1 (N981, N967);
xor XOR2 (N982, N976, N896);
not NOT1 (N983, N979);
not NOT1 (N984, N974);
or OR2 (N985, N973, N691);
xor XOR2 (N986, N965, N470);
nor NOR2 (N987, N977, N31);
nor NOR4 (N988, N983, N718, N799, N725);
not NOT1 (N989, N968);
not NOT1 (N990, N981);
and AND4 (N991, N985, N825, N263, N327);
and AND4 (N992, N987, N140, N791, N453);
and AND3 (N993, N988, N854, N521);
and AND3 (N994, N991, N57, N228);
or OR3 (N995, N994, N220, N40);
not NOT1 (N996, N992);
or OR4 (N997, N993, N599, N94, N252);
buf BUF1 (N998, N982);
nor NOR2 (N999, N980, N542);
and AND3 (N1000, N996, N951, N707);
nor NOR2 (N1001, N1000, N341);
not NOT1 (N1002, N998);
and AND3 (N1003, N986, N636, N420);
buf BUF1 (N1004, N990);
xor XOR2 (N1005, N984, N241);
nor NOR4 (N1006, N997, N895, N57, N20);
not NOT1 (N1007, N978);
or OR3 (N1008, N1001, N859, N351);
buf BUF1 (N1009, N999);
not NOT1 (N1010, N1003);
buf BUF1 (N1011, N1006);
buf BUF1 (N1012, N1007);
nor NOR2 (N1013, N1008, N806);
buf BUF1 (N1014, N1004);
buf BUF1 (N1015, N989);
nor NOR3 (N1016, N1012, N63, N968);
nand NAND3 (N1017, N1010, N699, N334);
and AND3 (N1018, N1013, N128, N117);
nor NOR2 (N1019, N1011, N59);
nor NOR2 (N1020, N1019, N359);
and AND2 (N1021, N1015, N852);
xor XOR2 (N1022, N1020, N514);
buf BUF1 (N1023, N1017);
and AND3 (N1024, N1021, N485, N120);
nor NOR4 (N1025, N1022, N363, N853, N841);
nand NAND4 (N1026, N1009, N33, N285, N343);
or OR2 (N1027, N1025, N145);
buf BUF1 (N1028, N1002);
nand NAND2 (N1029, N1024, N747);
xor XOR2 (N1030, N1016, N60);
nor NOR2 (N1031, N1030, N218);
xor XOR2 (N1032, N1014, N122);
or OR2 (N1033, N1023, N24);
and AND3 (N1034, N995, N775, N652);
not NOT1 (N1035, N1026);
xor XOR2 (N1036, N1029, N392);
buf BUF1 (N1037, N1033);
nor NOR2 (N1038, N1005, N795);
nor NOR2 (N1039, N1018, N747);
nand NAND3 (N1040, N1037, N505, N362);
not NOT1 (N1041, N1034);
or OR3 (N1042, N1035, N273, N928);
not NOT1 (N1043, N1027);
and AND2 (N1044, N1031, N54);
nor NOR3 (N1045, N1043, N362, N32);
nor NOR3 (N1046, N1036, N900, N757);
nor NOR3 (N1047, N1038, N385, N583);
and AND2 (N1048, N1044, N850);
and AND3 (N1049, N1039, N232, N652);
xor XOR2 (N1050, N1032, N835);
nor NOR2 (N1051, N1050, N646);
not NOT1 (N1052, N1045);
or OR3 (N1053, N1051, N420, N1034);
nand NAND4 (N1054, N1046, N226, N259, N1037);
or OR2 (N1055, N1052, N6);
or OR2 (N1056, N1047, N510);
not NOT1 (N1057, N1054);
nor NOR3 (N1058, N1055, N411, N551);
or OR3 (N1059, N1042, N730, N262);
nor NOR4 (N1060, N1053, N188, N285, N483);
buf BUF1 (N1061, N1059);
nor NOR2 (N1062, N1049, N767);
nor NOR3 (N1063, N1062, N817, N625);
nand NAND3 (N1064, N1061, N692, N1046);
or OR4 (N1065, N1056, N739, N437, N721);
nor NOR3 (N1066, N1064, N548, N892);
xor XOR2 (N1067, N1057, N169);
xor XOR2 (N1068, N1065, N313);
and AND3 (N1069, N1028, N553, N930);
and AND4 (N1070, N1041, N731, N524, N733);
buf BUF1 (N1071, N1069);
nor NOR4 (N1072, N1063, N751, N756, N659);
or OR3 (N1073, N1048, N1011, N1055);
nor NOR3 (N1074, N1067, N1043, N878);
nand NAND2 (N1075, N1073, N599);
nor NOR3 (N1076, N1060, N717, N727);
nand NAND4 (N1077, N1071, N130, N1041, N1072);
nand NAND2 (N1078, N725, N664);
nand NAND2 (N1079, N1058, N703);
nand NAND2 (N1080, N1078, N1001);
or OR3 (N1081, N1077, N766, N757);
not NOT1 (N1082, N1076);
xor XOR2 (N1083, N1068, N92);
and AND4 (N1084, N1083, N973, N455, N937);
xor XOR2 (N1085, N1084, N43);
buf BUF1 (N1086, N1070);
xor XOR2 (N1087, N1080, N310);
nor NOR3 (N1088, N1082, N127, N219);
xor XOR2 (N1089, N1079, N828);
buf BUF1 (N1090, N1074);
xor XOR2 (N1091, N1085, N102);
xor XOR2 (N1092, N1090, N1040);
xor XOR2 (N1093, N705, N268);
nor NOR3 (N1094, N1093, N306, N765);
nand NAND4 (N1095, N1081, N257, N239, N800);
nor NOR2 (N1096, N1066, N461);
nand NAND3 (N1097, N1092, N949, N50);
and AND2 (N1098, N1089, N24);
not NOT1 (N1099, N1097);
and AND2 (N1100, N1099, N713);
xor XOR2 (N1101, N1075, N1021);
buf BUF1 (N1102, N1087);
buf BUF1 (N1103, N1086);
xor XOR2 (N1104, N1096, N753);
nand NAND3 (N1105, N1098, N258, N1040);
nand NAND2 (N1106, N1102, N737);
or OR3 (N1107, N1101, N360, N577);
not NOT1 (N1108, N1091);
or OR4 (N1109, N1106, N590, N22, N1065);
buf BUF1 (N1110, N1108);
nor NOR4 (N1111, N1110, N690, N393, N881);
and AND4 (N1112, N1105, N618, N981, N869);
nand NAND4 (N1113, N1112, N991, N59, N370);
nand NAND3 (N1114, N1109, N330, N715);
nand NAND4 (N1115, N1113, N132, N548, N697);
not NOT1 (N1116, N1115);
and AND4 (N1117, N1103, N956, N208, N222);
and AND4 (N1118, N1114, N743, N458, N74);
buf BUF1 (N1119, N1107);
not NOT1 (N1120, N1116);
and AND4 (N1121, N1095, N353, N13, N1039);
buf BUF1 (N1122, N1111);
and AND2 (N1123, N1122, N598);
or OR2 (N1124, N1100, N442);
nor NOR4 (N1125, N1124, N779, N223, N573);
or OR2 (N1126, N1118, N408);
not NOT1 (N1127, N1125);
buf BUF1 (N1128, N1120);
nor NOR3 (N1129, N1117, N873, N208);
nand NAND4 (N1130, N1104, N77, N853, N251);
not NOT1 (N1131, N1130);
not NOT1 (N1132, N1123);
nand NAND3 (N1133, N1129, N891, N322);
nor NOR4 (N1134, N1088, N792, N380, N931);
xor XOR2 (N1135, N1126, N169);
nor NOR4 (N1136, N1134, N229, N706, N345);
and AND2 (N1137, N1127, N963);
buf BUF1 (N1138, N1119);
buf BUF1 (N1139, N1132);
and AND3 (N1140, N1137, N892, N1137);
nand NAND4 (N1141, N1131, N66, N30, N590);
nor NOR2 (N1142, N1121, N21);
not NOT1 (N1143, N1140);
not NOT1 (N1144, N1143);
not NOT1 (N1145, N1135);
nor NOR3 (N1146, N1139, N76, N849);
or OR3 (N1147, N1128, N1000, N915);
and AND2 (N1148, N1144, N890);
and AND4 (N1149, N1146, N12, N987, N29);
not NOT1 (N1150, N1149);
not NOT1 (N1151, N1147);
not NOT1 (N1152, N1142);
not NOT1 (N1153, N1152);
xor XOR2 (N1154, N1138, N607);
xor XOR2 (N1155, N1153, N985);
buf BUF1 (N1156, N1150);
or OR3 (N1157, N1133, N929, N650);
and AND3 (N1158, N1145, N553, N585);
and AND3 (N1159, N1156, N1111, N303);
nor NOR3 (N1160, N1157, N568, N304);
or OR4 (N1161, N1148, N572, N194, N772);
buf BUF1 (N1162, N1160);
nand NAND4 (N1163, N1159, N397, N476, N540);
xor XOR2 (N1164, N1162, N715);
not NOT1 (N1165, N1164);
not NOT1 (N1166, N1155);
nand NAND3 (N1167, N1166, N40, N518);
xor XOR2 (N1168, N1167, N889);
or OR4 (N1169, N1163, N974, N624, N617);
buf BUF1 (N1170, N1161);
xor XOR2 (N1171, N1169, N457);
nor NOR3 (N1172, N1168, N255, N803);
nor NOR3 (N1173, N1165, N24, N38);
nand NAND3 (N1174, N1094, N1068, N773);
nor NOR4 (N1175, N1173, N259, N419, N1087);
not NOT1 (N1176, N1136);
nor NOR2 (N1177, N1141, N196);
or OR4 (N1178, N1174, N151, N692, N1027);
or OR4 (N1179, N1154, N45, N487, N635);
nor NOR2 (N1180, N1151, N1066);
nor NOR4 (N1181, N1172, N410, N974, N945);
buf BUF1 (N1182, N1179);
buf BUF1 (N1183, N1178);
xor XOR2 (N1184, N1183, N794);
nor NOR3 (N1185, N1171, N427, N1054);
buf BUF1 (N1186, N1176);
and AND4 (N1187, N1177, N1079, N231, N457);
and AND2 (N1188, N1186, N217);
nand NAND4 (N1189, N1180, N985, N717, N1058);
nor NOR3 (N1190, N1184, N1030, N1113);
buf BUF1 (N1191, N1188);
buf BUF1 (N1192, N1187);
and AND3 (N1193, N1185, N177, N668);
nand NAND2 (N1194, N1182, N1023);
nand NAND3 (N1195, N1193, N759, N620);
nand NAND2 (N1196, N1190, N165);
or OR4 (N1197, N1192, N1011, N1077, N1016);
nor NOR2 (N1198, N1191, N669);
and AND3 (N1199, N1181, N544, N382);
and AND4 (N1200, N1158, N425, N940, N847);
nand NAND3 (N1201, N1195, N39, N413);
xor XOR2 (N1202, N1194, N167);
nor NOR2 (N1203, N1202, N1178);
nor NOR3 (N1204, N1175, N690, N1153);
buf BUF1 (N1205, N1203);
xor XOR2 (N1206, N1201, N117);
buf BUF1 (N1207, N1198);
or OR3 (N1208, N1197, N567, N1191);
not NOT1 (N1209, N1196);
nor NOR4 (N1210, N1207, N171, N482, N141);
buf BUF1 (N1211, N1200);
or OR4 (N1212, N1209, N728, N353, N153);
buf BUF1 (N1213, N1199);
buf BUF1 (N1214, N1206);
xor XOR2 (N1215, N1170, N829);
nand NAND3 (N1216, N1210, N1005, N341);
buf BUF1 (N1217, N1213);
not NOT1 (N1218, N1214);
nand NAND4 (N1219, N1208, N1109, N569, N341);
nand NAND4 (N1220, N1212, N659, N1120, N1115);
nor NOR4 (N1221, N1217, N609, N537, N386);
nand NAND4 (N1222, N1216, N1114, N473, N522);
nor NOR4 (N1223, N1204, N649, N527, N562);
and AND2 (N1224, N1219, N1220);
buf BUF1 (N1225, N366);
not NOT1 (N1226, N1189);
nor NOR4 (N1227, N1224, N748, N76, N504);
or OR3 (N1228, N1211, N1197, N920);
or OR3 (N1229, N1218, N163, N461);
xor XOR2 (N1230, N1228, N943);
nor NOR4 (N1231, N1221, N813, N181, N955);
xor XOR2 (N1232, N1225, N755);
or OR2 (N1233, N1232, N112);
or OR4 (N1234, N1222, N266, N503, N922);
and AND3 (N1235, N1223, N1113, N145);
nor NOR3 (N1236, N1233, N1026, N461);
or OR2 (N1237, N1226, N246);
not NOT1 (N1238, N1230);
nand NAND2 (N1239, N1227, N832);
nor NOR3 (N1240, N1236, N440, N361);
xor XOR2 (N1241, N1235, N970);
nor NOR3 (N1242, N1231, N7, N650);
nor NOR3 (N1243, N1229, N76, N547);
buf BUF1 (N1244, N1239);
buf BUF1 (N1245, N1215);
or OR4 (N1246, N1240, N218, N400, N232);
nand NAND2 (N1247, N1237, N1237);
nand NAND4 (N1248, N1241, N113, N1133, N534);
nor NOR4 (N1249, N1238, N101, N245, N34);
and AND3 (N1250, N1243, N596, N238);
nand NAND3 (N1251, N1234, N280, N1139);
or OR2 (N1252, N1246, N13);
nand NAND4 (N1253, N1248, N993, N1093, N279);
and AND2 (N1254, N1253, N951);
and AND2 (N1255, N1254, N1204);
nand NAND3 (N1256, N1250, N1244, N931);
nand NAND3 (N1257, N951, N1163, N851);
xor XOR2 (N1258, N1255, N1240);
xor XOR2 (N1259, N1205, N359);
nor NOR2 (N1260, N1249, N492);
buf BUF1 (N1261, N1251);
xor XOR2 (N1262, N1259, N510);
buf BUF1 (N1263, N1260);
nand NAND4 (N1264, N1261, N682, N255, N826);
not NOT1 (N1265, N1252);
xor XOR2 (N1266, N1262, N460);
nand NAND2 (N1267, N1257, N624);
or OR4 (N1268, N1242, N666, N798, N277);
not NOT1 (N1269, N1247);
nand NAND3 (N1270, N1269, N565, N1135);
not NOT1 (N1271, N1268);
nand NAND2 (N1272, N1267, N1203);
nand NAND4 (N1273, N1266, N270, N576, N826);
not NOT1 (N1274, N1258);
and AND3 (N1275, N1256, N1093, N914);
xor XOR2 (N1276, N1245, N1054);
or OR2 (N1277, N1264, N118);
buf BUF1 (N1278, N1271);
nor NOR4 (N1279, N1270, N93, N1226, N525);
not NOT1 (N1280, N1265);
buf BUF1 (N1281, N1273);
buf BUF1 (N1282, N1278);
nand NAND4 (N1283, N1275, N1158, N839, N256);
xor XOR2 (N1284, N1272, N880);
and AND2 (N1285, N1274, N1199);
not NOT1 (N1286, N1281);
buf BUF1 (N1287, N1285);
nand NAND3 (N1288, N1279, N481, N914);
and AND2 (N1289, N1282, N1063);
buf BUF1 (N1290, N1280);
xor XOR2 (N1291, N1288, N9);
xor XOR2 (N1292, N1291, N1045);
xor XOR2 (N1293, N1283, N926);
and AND2 (N1294, N1289, N1237);
xor XOR2 (N1295, N1292, N747);
not NOT1 (N1296, N1284);
buf BUF1 (N1297, N1290);
xor XOR2 (N1298, N1293, N669);
xor XOR2 (N1299, N1298, N385);
not NOT1 (N1300, N1299);
buf BUF1 (N1301, N1296);
not NOT1 (N1302, N1295);
xor XOR2 (N1303, N1277, N136);
xor XOR2 (N1304, N1263, N688);
nand NAND3 (N1305, N1294, N959, N703);
or OR4 (N1306, N1303, N1260, N738, N1136);
nand NAND4 (N1307, N1301, N465, N569, N505);
xor XOR2 (N1308, N1305, N839);
not NOT1 (N1309, N1276);
buf BUF1 (N1310, N1297);
not NOT1 (N1311, N1310);
nor NOR2 (N1312, N1307, N1240);
xor XOR2 (N1313, N1309, N90);
not NOT1 (N1314, N1286);
buf BUF1 (N1315, N1304);
xor XOR2 (N1316, N1306, N631);
buf BUF1 (N1317, N1302);
or OR2 (N1318, N1287, N321);
and AND4 (N1319, N1314, N1006, N959, N656);
not NOT1 (N1320, N1318);
buf BUF1 (N1321, N1320);
not NOT1 (N1322, N1317);
not NOT1 (N1323, N1322);
nor NOR2 (N1324, N1312, N1114);
nand NAND2 (N1325, N1308, N329);
buf BUF1 (N1326, N1315);
not NOT1 (N1327, N1313);
xor XOR2 (N1328, N1324, N134);
nand NAND3 (N1329, N1323, N503, N121);
or OR4 (N1330, N1326, N433, N741, N664);
xor XOR2 (N1331, N1311, N70);
nor NOR4 (N1332, N1300, N868, N413, N644);
or OR3 (N1333, N1330, N419, N109);
nand NAND4 (N1334, N1316, N848, N590, N985);
xor XOR2 (N1335, N1321, N138);
nor NOR2 (N1336, N1328, N878);
and AND2 (N1337, N1332, N1239);
not NOT1 (N1338, N1337);
buf BUF1 (N1339, N1335);
or OR4 (N1340, N1336, N1004, N1317, N983);
and AND4 (N1341, N1333, N168, N1270, N343);
xor XOR2 (N1342, N1334, N548);
xor XOR2 (N1343, N1342, N348);
nor NOR4 (N1344, N1340, N941, N458, N754);
nand NAND2 (N1345, N1339, N642);
nor NOR3 (N1346, N1331, N920, N1238);
nand NAND4 (N1347, N1344, N273, N674, N993);
xor XOR2 (N1348, N1341, N47);
or OR3 (N1349, N1348, N892, N475);
buf BUF1 (N1350, N1319);
or OR4 (N1351, N1346, N764, N1154, N896);
nor NOR3 (N1352, N1351, N950, N164);
and AND2 (N1353, N1349, N400);
or OR3 (N1354, N1352, N452, N151);
xor XOR2 (N1355, N1327, N774);
not NOT1 (N1356, N1350);
buf BUF1 (N1357, N1355);
nand NAND3 (N1358, N1329, N502, N1326);
and AND3 (N1359, N1345, N415, N603);
xor XOR2 (N1360, N1358, N363);
nor NOR3 (N1361, N1343, N1276, N792);
xor XOR2 (N1362, N1359, N958);
nor NOR3 (N1363, N1356, N1227, N996);
buf BUF1 (N1364, N1338);
not NOT1 (N1365, N1353);
nor NOR2 (N1366, N1360, N769);
and AND2 (N1367, N1357, N1100);
xor XOR2 (N1368, N1365, N482);
or OR3 (N1369, N1367, N259, N148);
nor NOR4 (N1370, N1361, N1262, N1270, N360);
nor NOR4 (N1371, N1363, N1297, N77, N618);
or OR4 (N1372, N1371, N691, N727, N1318);
xor XOR2 (N1373, N1364, N840);
nand NAND4 (N1374, N1366, N182, N534, N1132);
and AND4 (N1375, N1369, N36, N455, N852);
buf BUF1 (N1376, N1370);
xor XOR2 (N1377, N1375, N331);
or OR2 (N1378, N1325, N47);
and AND3 (N1379, N1372, N725, N758);
nand NAND4 (N1380, N1374, N403, N357, N809);
xor XOR2 (N1381, N1373, N369);
nor NOR4 (N1382, N1354, N1039, N136, N1342);
xor XOR2 (N1383, N1382, N692);
buf BUF1 (N1384, N1347);
or OR3 (N1385, N1377, N1081, N868);
not NOT1 (N1386, N1379);
and AND4 (N1387, N1383, N825, N87, N430);
buf BUF1 (N1388, N1362);
not NOT1 (N1389, N1388);
or OR3 (N1390, N1380, N763, N1263);
xor XOR2 (N1391, N1384, N365);
and AND2 (N1392, N1387, N23);
nand NAND4 (N1393, N1390, N822, N1310, N15);
xor XOR2 (N1394, N1378, N578);
nor NOR4 (N1395, N1389, N630, N920, N203);
xor XOR2 (N1396, N1391, N1067);
buf BUF1 (N1397, N1386);
not NOT1 (N1398, N1376);
or OR4 (N1399, N1398, N95, N1063, N992);
nor NOR2 (N1400, N1396, N1302);
nor NOR4 (N1401, N1392, N806, N949, N1384);
nor NOR2 (N1402, N1381, N242);
xor XOR2 (N1403, N1368, N636);
nand NAND4 (N1404, N1397, N441, N1350, N811);
not NOT1 (N1405, N1400);
and AND3 (N1406, N1393, N1227, N1399);
not NOT1 (N1407, N77);
and AND2 (N1408, N1401, N395);
and AND3 (N1409, N1407, N634, N213);
nor NOR4 (N1410, N1403, N843, N897, N131);
xor XOR2 (N1411, N1410, N906);
nor NOR3 (N1412, N1395, N1125, N654);
xor XOR2 (N1413, N1411, N347);
xor XOR2 (N1414, N1402, N1262);
xor XOR2 (N1415, N1412, N24);
nor NOR3 (N1416, N1414, N362, N1093);
and AND3 (N1417, N1408, N1082, N553);
buf BUF1 (N1418, N1385);
and AND4 (N1419, N1406, N652, N869, N838);
and AND3 (N1420, N1415, N1348, N487);
and AND2 (N1421, N1417, N425);
nand NAND2 (N1422, N1418, N268);
xor XOR2 (N1423, N1419, N674);
xor XOR2 (N1424, N1409, N696);
or OR2 (N1425, N1421, N631);
xor XOR2 (N1426, N1424, N232);
buf BUF1 (N1427, N1416);
nor NOR2 (N1428, N1422, N306);
nor NOR3 (N1429, N1428, N1360, N517);
or OR4 (N1430, N1420, N779, N713, N1080);
buf BUF1 (N1431, N1426);
and AND3 (N1432, N1394, N1358, N480);
or OR2 (N1433, N1413, N1155);
nand NAND2 (N1434, N1404, N1284);
nor NOR3 (N1435, N1430, N375, N1003);
nand NAND4 (N1436, N1435, N1318, N720, N318);
nand NAND3 (N1437, N1425, N1124, N379);
and AND2 (N1438, N1434, N516);
nand NAND3 (N1439, N1438, N705, N1043);
xor XOR2 (N1440, N1436, N1282);
and AND4 (N1441, N1440, N574, N1084, N686);
and AND3 (N1442, N1441, N138, N444);
xor XOR2 (N1443, N1427, N615);
not NOT1 (N1444, N1432);
xor XOR2 (N1445, N1429, N146);
buf BUF1 (N1446, N1443);
buf BUF1 (N1447, N1446);
not NOT1 (N1448, N1445);
or OR2 (N1449, N1431, N1178);
nand NAND4 (N1450, N1448, N829, N657, N633);
or OR2 (N1451, N1447, N1078);
buf BUF1 (N1452, N1449);
or OR3 (N1453, N1437, N707, N858);
or OR3 (N1454, N1444, N1251, N160);
not NOT1 (N1455, N1450);
xor XOR2 (N1456, N1451, N812);
not NOT1 (N1457, N1455);
buf BUF1 (N1458, N1457);
xor XOR2 (N1459, N1433, N261);
buf BUF1 (N1460, N1405);
buf BUF1 (N1461, N1456);
nand NAND4 (N1462, N1461, N201, N1340, N39);
not NOT1 (N1463, N1462);
not NOT1 (N1464, N1442);
or OR4 (N1465, N1463, N1353, N1395, N206);
not NOT1 (N1466, N1452);
nand NAND2 (N1467, N1464, N493);
or OR4 (N1468, N1465, N754, N1422, N505);
buf BUF1 (N1469, N1467);
and AND3 (N1470, N1423, N906, N168);
xor XOR2 (N1471, N1453, N785);
nor NOR4 (N1472, N1469, N558, N12, N951);
nand NAND2 (N1473, N1460, N1468);
xor XOR2 (N1474, N1256, N1358);
and AND2 (N1475, N1458, N1169);
or OR2 (N1476, N1439, N232);
and AND4 (N1477, N1476, N1457, N361, N388);
xor XOR2 (N1478, N1477, N1359);
or OR2 (N1479, N1478, N51);
or OR2 (N1480, N1473, N463);
nand NAND4 (N1481, N1479, N304, N167, N104);
buf BUF1 (N1482, N1454);
buf BUF1 (N1483, N1466);
not NOT1 (N1484, N1474);
nand NAND2 (N1485, N1480, N72);
xor XOR2 (N1486, N1471, N7);
and AND4 (N1487, N1482, N887, N1268, N440);
and AND3 (N1488, N1472, N503, N209);
xor XOR2 (N1489, N1488, N650);
xor XOR2 (N1490, N1481, N268);
or OR2 (N1491, N1489, N780);
not NOT1 (N1492, N1484);
xor XOR2 (N1493, N1491, N1471);
nand NAND3 (N1494, N1470, N982, N546);
nor NOR4 (N1495, N1475, N1237, N1263, N1182);
nor NOR4 (N1496, N1490, N458, N361, N842);
or OR3 (N1497, N1483, N1384, N1488);
or OR2 (N1498, N1494, N1347);
nand NAND4 (N1499, N1486, N566, N207, N898);
and AND3 (N1500, N1459, N287, N1281);
nand NAND2 (N1501, N1493, N655);
xor XOR2 (N1502, N1485, N522);
nor NOR2 (N1503, N1496, N192);
not NOT1 (N1504, N1497);
or OR4 (N1505, N1503, N1007, N871, N658);
or OR3 (N1506, N1502, N580, N1457);
buf BUF1 (N1507, N1505);
or OR3 (N1508, N1495, N521, N72);
buf BUF1 (N1509, N1499);
and AND2 (N1510, N1492, N158);
nand NAND2 (N1511, N1504, N926);
not NOT1 (N1512, N1509);
nand NAND2 (N1513, N1501, N607);
xor XOR2 (N1514, N1500, N1500);
nor NOR4 (N1515, N1507, N379, N829, N1349);
buf BUF1 (N1516, N1487);
not NOT1 (N1517, N1508);
not NOT1 (N1518, N1498);
xor XOR2 (N1519, N1516, N257);
and AND3 (N1520, N1518, N719, N612);
not NOT1 (N1521, N1515);
nand NAND2 (N1522, N1521, N1017);
or OR3 (N1523, N1514, N1104, N398);
not NOT1 (N1524, N1519);
and AND4 (N1525, N1520, N887, N1234, N546);
and AND3 (N1526, N1513, N165, N953);
nor NOR3 (N1527, N1526, N738, N495);
not NOT1 (N1528, N1524);
and AND4 (N1529, N1523, N1159, N916, N1407);
nand NAND2 (N1530, N1510, N100);
or OR3 (N1531, N1529, N163, N1214);
or OR2 (N1532, N1531, N871);
nor NOR4 (N1533, N1532, N230, N1400, N130);
xor XOR2 (N1534, N1517, N1373);
or OR2 (N1535, N1525, N1432);
or OR3 (N1536, N1530, N1176, N434);
and AND3 (N1537, N1528, N1388, N758);
nor NOR2 (N1538, N1522, N1454);
xor XOR2 (N1539, N1533, N593);
nand NAND2 (N1540, N1534, N744);
nand NAND3 (N1541, N1539, N1227, N593);
nand NAND2 (N1542, N1536, N1112);
nand NAND4 (N1543, N1506, N93, N64, N818);
not NOT1 (N1544, N1540);
xor XOR2 (N1545, N1527, N1317);
xor XOR2 (N1546, N1545, N44);
or OR2 (N1547, N1546, N1302);
and AND2 (N1548, N1547, N1005);
or OR3 (N1549, N1537, N969, N9);
or OR2 (N1550, N1511, N902);
nand NAND4 (N1551, N1550, N159, N1063, N969);
and AND2 (N1552, N1541, N777);
nand NAND4 (N1553, N1535, N1072, N823, N123);
buf BUF1 (N1554, N1549);
and AND3 (N1555, N1553, N560, N450);
and AND3 (N1556, N1543, N952, N1120);
nand NAND3 (N1557, N1552, N1187, N759);
nand NAND2 (N1558, N1551, N509);
buf BUF1 (N1559, N1556);
nor NOR2 (N1560, N1548, N1413);
buf BUF1 (N1561, N1558);
or OR2 (N1562, N1560, N63);
nor NOR2 (N1563, N1559, N1446);
and AND4 (N1564, N1562, N1532, N638, N218);
nor NOR4 (N1565, N1564, N1057, N1188, N721);
or OR3 (N1566, N1512, N1011, N1084);
nand NAND4 (N1567, N1555, N972, N605, N783);
xor XOR2 (N1568, N1566, N609);
buf BUF1 (N1569, N1544);
buf BUF1 (N1570, N1568);
not NOT1 (N1571, N1565);
buf BUF1 (N1572, N1570);
nor NOR2 (N1573, N1557, N625);
or OR3 (N1574, N1572, N167, N115);
buf BUF1 (N1575, N1569);
and AND2 (N1576, N1563, N669);
or OR2 (N1577, N1561, N290);
buf BUF1 (N1578, N1573);
buf BUF1 (N1579, N1578);
xor XOR2 (N1580, N1542, N1002);
nor NOR4 (N1581, N1574, N676, N1040, N1442);
xor XOR2 (N1582, N1581, N972);
buf BUF1 (N1583, N1567);
or OR4 (N1584, N1538, N417, N1, N74);
or OR2 (N1585, N1580, N1018);
nand NAND3 (N1586, N1582, N950, N1011);
xor XOR2 (N1587, N1571, N548);
or OR4 (N1588, N1587, N154, N487, N859);
xor XOR2 (N1589, N1575, N969);
or OR3 (N1590, N1585, N1153, N1068);
buf BUF1 (N1591, N1579);
or OR2 (N1592, N1577, N1118);
or OR2 (N1593, N1592, N1370);
and AND3 (N1594, N1590, N1230, N974);
nand NAND2 (N1595, N1589, N16);
nand NAND4 (N1596, N1588, N1005, N1426, N718);
buf BUF1 (N1597, N1583);
nand NAND2 (N1598, N1586, N580);
not NOT1 (N1599, N1584);
nand NAND4 (N1600, N1599, N220, N930, N78);
nand NAND4 (N1601, N1576, N1088, N1187, N1065);
xor XOR2 (N1602, N1600, N1322);
xor XOR2 (N1603, N1554, N345);
xor XOR2 (N1604, N1602, N312);
xor XOR2 (N1605, N1596, N1307);
nand NAND3 (N1606, N1595, N1177, N275);
buf BUF1 (N1607, N1605);
not NOT1 (N1608, N1597);
not NOT1 (N1609, N1591);
buf BUF1 (N1610, N1593);
not NOT1 (N1611, N1594);
nor NOR3 (N1612, N1611, N1458, N1610);
or OR4 (N1613, N833, N229, N1031, N1506);
or OR4 (N1614, N1606, N1328, N472, N800);
nand NAND2 (N1615, N1603, N562);
not NOT1 (N1616, N1609);
buf BUF1 (N1617, N1604);
nand NAND4 (N1618, N1613, N710, N308, N1506);
buf BUF1 (N1619, N1601);
and AND2 (N1620, N1618, N250);
not NOT1 (N1621, N1617);
and AND3 (N1622, N1607, N1453, N897);
and AND2 (N1623, N1598, N387);
and AND3 (N1624, N1619, N292, N448);
buf BUF1 (N1625, N1608);
nand NAND3 (N1626, N1622, N159, N1021);
xor XOR2 (N1627, N1621, N1027);
buf BUF1 (N1628, N1623);
buf BUF1 (N1629, N1616);
nand NAND2 (N1630, N1626, N1434);
xor XOR2 (N1631, N1614, N901);
not NOT1 (N1632, N1629);
buf BUF1 (N1633, N1632);
nand NAND2 (N1634, N1615, N911);
xor XOR2 (N1635, N1634, N105);
buf BUF1 (N1636, N1627);
xor XOR2 (N1637, N1633, N850);
buf BUF1 (N1638, N1637);
and AND3 (N1639, N1636, N299, N281);
or OR2 (N1640, N1620, N995);
xor XOR2 (N1641, N1612, N341);
nand NAND2 (N1642, N1630, N584);
nor NOR3 (N1643, N1639, N120, N1081);
nor NOR3 (N1644, N1643, N784, N219);
nor NOR4 (N1645, N1635, N966, N545, N1217);
nand NAND4 (N1646, N1625, N282, N926, N196);
xor XOR2 (N1647, N1641, N541);
buf BUF1 (N1648, N1646);
xor XOR2 (N1649, N1644, N117);
not NOT1 (N1650, N1631);
buf BUF1 (N1651, N1649);
not NOT1 (N1652, N1648);
not NOT1 (N1653, N1642);
not NOT1 (N1654, N1638);
nand NAND4 (N1655, N1624, N829, N1652, N1644);
nand NAND3 (N1656, N914, N952, N107);
nand NAND4 (N1657, N1656, N1437, N921, N1294);
xor XOR2 (N1658, N1655, N1359);
and AND4 (N1659, N1628, N1586, N1430, N486);
nand NAND2 (N1660, N1640, N1477);
nor NOR2 (N1661, N1647, N971);
and AND2 (N1662, N1653, N310);
nor NOR3 (N1663, N1662, N1013, N976);
or OR4 (N1664, N1654, N996, N1310, N1147);
buf BUF1 (N1665, N1650);
and AND3 (N1666, N1659, N466, N704);
or OR3 (N1667, N1660, N228, N1003);
not NOT1 (N1668, N1661);
or OR2 (N1669, N1665, N1575);
buf BUF1 (N1670, N1651);
and AND2 (N1671, N1664, N1486);
xor XOR2 (N1672, N1670, N844);
and AND3 (N1673, N1671, N616, N132);
nor NOR4 (N1674, N1669, N107, N1555, N874);
or OR3 (N1675, N1673, N1346, N1208);
or OR3 (N1676, N1657, N1056, N970);
and AND4 (N1677, N1675, N982, N781, N1560);
nand NAND4 (N1678, N1677, N775, N802, N887);
xor XOR2 (N1679, N1658, N141);
or OR2 (N1680, N1676, N458);
not NOT1 (N1681, N1674);
and AND2 (N1682, N1681, N948);
xor XOR2 (N1683, N1667, N980);
nand NAND2 (N1684, N1666, N1252);
or OR3 (N1685, N1683, N1250, N801);
nand NAND2 (N1686, N1668, N1458);
not NOT1 (N1687, N1679);
xor XOR2 (N1688, N1672, N236);
and AND3 (N1689, N1680, N339, N752);
and AND2 (N1690, N1645, N1025);
buf BUF1 (N1691, N1688);
buf BUF1 (N1692, N1687);
nand NAND3 (N1693, N1685, N11, N535);
and AND3 (N1694, N1686, N930, N1010);
nor NOR4 (N1695, N1663, N756, N1372, N765);
or OR3 (N1696, N1694, N1151, N837);
buf BUF1 (N1697, N1695);
buf BUF1 (N1698, N1689);
not NOT1 (N1699, N1698);
or OR4 (N1700, N1678, N1482, N1022, N289);
xor XOR2 (N1701, N1697, N1564);
not NOT1 (N1702, N1691);
and AND4 (N1703, N1692, N659, N937, N754);
and AND2 (N1704, N1682, N1375);
buf BUF1 (N1705, N1696);
nor NOR4 (N1706, N1705, N667, N1691, N1656);
and AND2 (N1707, N1699, N1584);
nand NAND3 (N1708, N1684, N1087, N1324);
not NOT1 (N1709, N1690);
buf BUF1 (N1710, N1693);
buf BUF1 (N1711, N1702);
and AND2 (N1712, N1709, N653);
nand NAND4 (N1713, N1700, N1069, N175, N1548);
nand NAND2 (N1714, N1712, N1504);
or OR4 (N1715, N1714, N183, N91, N79);
or OR2 (N1716, N1706, N595);
nand NAND4 (N1717, N1707, N1367, N396, N544);
xor XOR2 (N1718, N1717, N798);
or OR3 (N1719, N1701, N1221, N5);
xor XOR2 (N1720, N1719, N160);
not NOT1 (N1721, N1716);
xor XOR2 (N1722, N1710, N864);
nor NOR3 (N1723, N1703, N1329, N1216);
and AND4 (N1724, N1708, N451, N427, N411);
and AND3 (N1725, N1722, N1576, N1065);
nor NOR3 (N1726, N1704, N1242, N337);
and AND4 (N1727, N1721, N1054, N204, N728);
and AND3 (N1728, N1718, N140, N54);
xor XOR2 (N1729, N1725, N906);
nor NOR3 (N1730, N1728, N492, N596);
xor XOR2 (N1731, N1726, N1431);
nor NOR4 (N1732, N1727, N696, N738, N760);
buf BUF1 (N1733, N1730);
or OR3 (N1734, N1715, N729, N1143);
nand NAND3 (N1735, N1729, N350, N1035);
nand NAND4 (N1736, N1711, N338, N314, N1677);
buf BUF1 (N1737, N1733);
or OR2 (N1738, N1735, N1371);
and AND2 (N1739, N1734, N35);
buf BUF1 (N1740, N1731);
nor NOR4 (N1741, N1737, N876, N1695, N489);
nand NAND4 (N1742, N1736, N675, N529, N30);
or OR4 (N1743, N1739, N786, N230, N1298);
buf BUF1 (N1744, N1732);
or OR2 (N1745, N1724, N1355);
buf BUF1 (N1746, N1742);
buf BUF1 (N1747, N1743);
buf BUF1 (N1748, N1745);
or OR3 (N1749, N1723, N465, N933);
and AND3 (N1750, N1713, N808, N1678);
nor NOR4 (N1751, N1749, N553, N71, N1659);
and AND3 (N1752, N1740, N91, N1686);
not NOT1 (N1753, N1747);
nor NOR3 (N1754, N1746, N1105, N1044);
buf BUF1 (N1755, N1744);
buf BUF1 (N1756, N1753);
nor NOR2 (N1757, N1751, N809);
or OR4 (N1758, N1755, N846, N397, N55);
not NOT1 (N1759, N1752);
and AND3 (N1760, N1748, N28, N1649);
and AND4 (N1761, N1760, N548, N1405, N1065);
nand NAND3 (N1762, N1750, N1484, N319);
and AND4 (N1763, N1761, N945, N31, N1623);
nand NAND3 (N1764, N1762, N1314, N1670);
nand NAND2 (N1765, N1741, N165);
and AND4 (N1766, N1765, N1222, N513, N296);
or OR4 (N1767, N1756, N1446, N443, N66);
not NOT1 (N1768, N1738);
not NOT1 (N1769, N1720);
buf BUF1 (N1770, N1757);
or OR2 (N1771, N1759, N1095);
xor XOR2 (N1772, N1770, N1754);
nor NOR2 (N1773, N1614, N469);
and AND4 (N1774, N1773, N140, N541, N935);
and AND2 (N1775, N1771, N957);
buf BUF1 (N1776, N1764);
not NOT1 (N1777, N1776);
xor XOR2 (N1778, N1775, N265);
or OR4 (N1779, N1774, N407, N223, N538);
and AND4 (N1780, N1772, N1018, N1338, N566);
nand NAND4 (N1781, N1780, N293, N1367, N180);
nor NOR2 (N1782, N1768, N951);
nand NAND4 (N1783, N1766, N463, N511, N1067);
buf BUF1 (N1784, N1781);
not NOT1 (N1785, N1769);
xor XOR2 (N1786, N1758, N1168);
buf BUF1 (N1787, N1784);
and AND3 (N1788, N1783, N1701, N100);
xor XOR2 (N1789, N1779, N886);
xor XOR2 (N1790, N1785, N1288);
nor NOR3 (N1791, N1786, N618, N1756);
nand NAND2 (N1792, N1790, N9);
and AND4 (N1793, N1791, N1383, N1056, N1757);
buf BUF1 (N1794, N1787);
buf BUF1 (N1795, N1794);
xor XOR2 (N1796, N1792, N999);
or OR3 (N1797, N1793, N717, N636);
xor XOR2 (N1798, N1777, N619);
buf BUF1 (N1799, N1782);
buf BUF1 (N1800, N1789);
xor XOR2 (N1801, N1778, N1605);
and AND2 (N1802, N1763, N1510);
not NOT1 (N1803, N1800);
not NOT1 (N1804, N1802);
or OR3 (N1805, N1797, N1246, N1374);
xor XOR2 (N1806, N1795, N717);
or OR2 (N1807, N1806, N1441);
and AND4 (N1808, N1796, N261, N378, N1101);
or OR3 (N1809, N1801, N1677, N742);
and AND4 (N1810, N1788, N365, N206, N853);
nand NAND4 (N1811, N1798, N788, N942, N1772);
buf BUF1 (N1812, N1811);
not NOT1 (N1813, N1810);
or OR3 (N1814, N1799, N447, N518);
xor XOR2 (N1815, N1807, N1054);
nor NOR2 (N1816, N1805, N272);
or OR4 (N1817, N1814, N435, N1421, N1264);
not NOT1 (N1818, N1809);
and AND2 (N1819, N1767, N1607);
buf BUF1 (N1820, N1803);
nor NOR3 (N1821, N1818, N206, N944);
or OR4 (N1822, N1821, N479, N766, N1235);
and AND3 (N1823, N1808, N799, N1);
not NOT1 (N1824, N1822);
and AND3 (N1825, N1824, N1424, N189);
xor XOR2 (N1826, N1820, N71);
nand NAND2 (N1827, N1817, N111);
or OR3 (N1828, N1812, N1797, N1247);
and AND3 (N1829, N1823, N536, N333);
buf BUF1 (N1830, N1816);
buf BUF1 (N1831, N1813);
or OR4 (N1832, N1825, N904, N724, N1142);
nand NAND4 (N1833, N1832, N796, N471, N1148);
nor NOR3 (N1834, N1815, N1335, N1771);
nor NOR4 (N1835, N1826, N1553, N1630, N702);
buf BUF1 (N1836, N1831);
not NOT1 (N1837, N1828);
nor NOR2 (N1838, N1827, N1341);
nor NOR3 (N1839, N1829, N339, N1615);
nand NAND4 (N1840, N1833, N1134, N1595, N218);
or OR4 (N1841, N1837, N270, N473, N611);
not NOT1 (N1842, N1835);
xor XOR2 (N1843, N1838, N544);
nand NAND4 (N1844, N1840, N909, N10, N1116);
buf BUF1 (N1845, N1843);
or OR2 (N1846, N1841, N377);
or OR3 (N1847, N1819, N709, N1472);
nand NAND2 (N1848, N1846, N1002);
nor NOR3 (N1849, N1848, N1203, N1631);
nand NAND3 (N1850, N1845, N1555, N869);
and AND2 (N1851, N1847, N1173);
nor NOR4 (N1852, N1849, N1100, N739, N1336);
not NOT1 (N1853, N1852);
buf BUF1 (N1854, N1836);
or OR4 (N1855, N1853, N508, N135, N934);
buf BUF1 (N1856, N1839);
buf BUF1 (N1857, N1804);
nand NAND3 (N1858, N1857, N1561, N1391);
xor XOR2 (N1859, N1842, N119);
or OR4 (N1860, N1834, N1267, N1716, N1528);
xor XOR2 (N1861, N1850, N591);
xor XOR2 (N1862, N1858, N1283);
not NOT1 (N1863, N1851);
buf BUF1 (N1864, N1844);
or OR4 (N1865, N1862, N1132, N1388, N649);
or OR4 (N1866, N1864, N1357, N197, N1343);
xor XOR2 (N1867, N1866, N858);
not NOT1 (N1868, N1856);
nor NOR4 (N1869, N1868, N950, N528, N811);
nand NAND4 (N1870, N1869, N932, N1699, N905);
not NOT1 (N1871, N1863);
nor NOR2 (N1872, N1855, N1189);
buf BUF1 (N1873, N1867);
xor XOR2 (N1874, N1859, N869);
xor XOR2 (N1875, N1860, N620);
nand NAND3 (N1876, N1865, N1690, N308);
nor NOR4 (N1877, N1870, N1285, N1334, N1671);
and AND2 (N1878, N1874, N1222);
xor XOR2 (N1879, N1878, N1307);
nand NAND3 (N1880, N1861, N1529, N60);
nand NAND4 (N1881, N1877, N594, N1091, N1397);
nor NOR4 (N1882, N1875, N959, N52, N56);
nand NAND3 (N1883, N1854, N1355, N1021);
nand NAND3 (N1884, N1872, N1457, N992);
buf BUF1 (N1885, N1876);
not NOT1 (N1886, N1883);
xor XOR2 (N1887, N1880, N1018);
nand NAND2 (N1888, N1879, N1692);
buf BUF1 (N1889, N1886);
or OR4 (N1890, N1881, N920, N220, N606);
not NOT1 (N1891, N1882);
and AND2 (N1892, N1889, N298);
or OR3 (N1893, N1887, N1232, N22);
or OR4 (N1894, N1890, N1866, N1234, N1315);
or OR2 (N1895, N1888, N1611);
xor XOR2 (N1896, N1873, N923);
and AND4 (N1897, N1884, N1050, N942, N1209);
buf BUF1 (N1898, N1895);
and AND3 (N1899, N1893, N1560, N1187);
and AND2 (N1900, N1885, N722);
nor NOR3 (N1901, N1899, N1179, N559);
nor NOR2 (N1902, N1896, N1343);
nor NOR3 (N1903, N1891, N276, N1258);
buf BUF1 (N1904, N1902);
nor NOR3 (N1905, N1871, N1035, N57);
xor XOR2 (N1906, N1830, N371);
not NOT1 (N1907, N1904);
not NOT1 (N1908, N1903);
not NOT1 (N1909, N1892);
not NOT1 (N1910, N1900);
nor NOR2 (N1911, N1910, N1670);
nor NOR3 (N1912, N1908, N677, N1499);
not NOT1 (N1913, N1907);
nand NAND2 (N1914, N1906, N1203);
xor XOR2 (N1915, N1901, N1760);
buf BUF1 (N1916, N1915);
nand NAND4 (N1917, N1905, N1233, N887, N1042);
xor XOR2 (N1918, N1898, N1001);
buf BUF1 (N1919, N1894);
nand NAND2 (N1920, N1909, N960);
buf BUF1 (N1921, N1897);
and AND2 (N1922, N1916, N965);
nand NAND3 (N1923, N1921, N35, N275);
not NOT1 (N1924, N1917);
or OR3 (N1925, N1912, N1, N9);
nor NOR4 (N1926, N1920, N870, N644, N962);
nor NOR3 (N1927, N1926, N1006, N1276);
nor NOR4 (N1928, N1919, N1229, N1669, N79);
xor XOR2 (N1929, N1928, N674);
xor XOR2 (N1930, N1922, N482);
nor NOR4 (N1931, N1927, N1205, N1184, N1153);
nand NAND3 (N1932, N1913, N357, N1059);
and AND3 (N1933, N1932, N1331, N1495);
nand NAND2 (N1934, N1925, N457);
xor XOR2 (N1935, N1934, N1548);
or OR3 (N1936, N1933, N1348, N33);
nand NAND2 (N1937, N1911, N1504);
xor XOR2 (N1938, N1937, N926);
not NOT1 (N1939, N1938);
nand NAND2 (N1940, N1923, N1169);
or OR3 (N1941, N1935, N1025, N306);
nand NAND3 (N1942, N1931, N1865, N1836);
or OR3 (N1943, N1941, N1089, N1580);
nor NOR4 (N1944, N1942, N617, N1248, N1459);
not NOT1 (N1945, N1943);
buf BUF1 (N1946, N1945);
buf BUF1 (N1947, N1944);
not NOT1 (N1948, N1924);
xor XOR2 (N1949, N1914, N1107);
not NOT1 (N1950, N1930);
buf BUF1 (N1951, N1950);
nor NOR3 (N1952, N1918, N670, N1437);
not NOT1 (N1953, N1940);
buf BUF1 (N1954, N1946);
nor NOR4 (N1955, N1952, N94, N717, N1054);
nor NOR4 (N1956, N1948, N821, N1191, N573);
not NOT1 (N1957, N1953);
buf BUF1 (N1958, N1947);
not NOT1 (N1959, N1955);
not NOT1 (N1960, N1939);
nand NAND4 (N1961, N1958, N1905, N1756, N998);
xor XOR2 (N1962, N1959, N1932);
not NOT1 (N1963, N1951);
and AND4 (N1964, N1957, N1297, N1361, N1178);
buf BUF1 (N1965, N1962);
nor NOR3 (N1966, N1964, N1479, N310);
nor NOR4 (N1967, N1954, N1392, N725, N878);
not NOT1 (N1968, N1963);
or OR3 (N1969, N1966, N342, N1322);
xor XOR2 (N1970, N1929, N544);
nand NAND3 (N1971, N1949, N1733, N816);
and AND4 (N1972, N1971, N594, N1373, N1620);
buf BUF1 (N1973, N1956);
xor XOR2 (N1974, N1970, N1578);
nor NOR2 (N1975, N1967, N321);
or OR4 (N1976, N1972, N1322, N294, N1430);
nor NOR3 (N1977, N1965, N1318, N725);
nand NAND4 (N1978, N1973, N1691, N1473, N1851);
buf BUF1 (N1979, N1976);
buf BUF1 (N1980, N1974);
and AND4 (N1981, N1936, N682, N763, N1798);
or OR3 (N1982, N1979, N622, N842);
nand NAND2 (N1983, N1969, N1567);
nand NAND3 (N1984, N1975, N1804, N393);
not NOT1 (N1985, N1983);
nand NAND4 (N1986, N1980, N297, N1959, N1789);
xor XOR2 (N1987, N1977, N1454);
or OR2 (N1988, N1968, N508);
xor XOR2 (N1989, N1987, N478);
and AND2 (N1990, N1989, N1727);
not NOT1 (N1991, N1982);
nor NOR3 (N1992, N1991, N1550, N1775);
xor XOR2 (N1993, N1981, N1024);
and AND2 (N1994, N1993, N1963);
xor XOR2 (N1995, N1992, N711);
buf BUF1 (N1996, N1986);
xor XOR2 (N1997, N1978, N236);
or OR4 (N1998, N1990, N836, N1879, N779);
nor NOR3 (N1999, N1960, N1740, N1754);
or OR4 (N2000, N1996, N1813, N1285, N1318);
buf BUF1 (N2001, N1961);
buf BUF1 (N2002, N2001);
buf BUF1 (N2003, N1988);
or OR3 (N2004, N2003, N1755, N513);
nand NAND4 (N2005, N2000, N1583, N501, N1983);
and AND3 (N2006, N2002, N1254, N145);
or OR3 (N2007, N1997, N679, N637);
xor XOR2 (N2008, N1985, N1622);
or OR4 (N2009, N1994, N485, N1756, N767);
or OR2 (N2010, N2004, N1070);
xor XOR2 (N2011, N1995, N1036);
and AND3 (N2012, N1984, N1976, N108);
or OR2 (N2013, N2006, N1884);
or OR2 (N2014, N2007, N1803);
nor NOR2 (N2015, N2012, N1931);
nor NOR3 (N2016, N2015, N230, N812);
not NOT1 (N2017, N1998);
nand NAND4 (N2018, N2011, N1625, N785, N238);
buf BUF1 (N2019, N2016);
nand NAND4 (N2020, N2005, N887, N1304, N1222);
nor NOR4 (N2021, N2017, N632, N1827, N391);
xor XOR2 (N2022, N2021, N802);
and AND2 (N2023, N2019, N683);
buf BUF1 (N2024, N1999);
xor XOR2 (N2025, N2022, N1597);
nor NOR3 (N2026, N2008, N405, N1607);
xor XOR2 (N2027, N2024, N465);
and AND4 (N2028, N2009, N963, N1925, N1326);
nor NOR2 (N2029, N2028, N143);
xor XOR2 (N2030, N2018, N1093);
nor NOR4 (N2031, N2030, N165, N927, N1571);
nand NAND2 (N2032, N2014, N446);
nand NAND3 (N2033, N2025, N378, N584);
xor XOR2 (N2034, N2033, N1939);
nor NOR4 (N2035, N2023, N937, N598, N1707);
xor XOR2 (N2036, N2020, N1146);
or OR2 (N2037, N2034, N1049);
not NOT1 (N2038, N2037);
not NOT1 (N2039, N2027);
or OR4 (N2040, N2039, N171, N538, N1230);
nor NOR2 (N2041, N2031, N842);
nand NAND3 (N2042, N2026, N1110, N1428);
nor NOR4 (N2043, N2038, N1725, N568, N955);
nor NOR3 (N2044, N2032, N123, N1791);
xor XOR2 (N2045, N2013, N1674);
nor NOR2 (N2046, N2040, N1905);
not NOT1 (N2047, N2036);
nand NAND4 (N2048, N2044, N169, N1609, N677);
xor XOR2 (N2049, N2046, N1584);
buf BUF1 (N2050, N2045);
nor NOR4 (N2051, N2029, N1070, N1630, N1737);
nor NOR3 (N2052, N2043, N1467, N981);
nor NOR4 (N2053, N2048, N1075, N1595, N293);
buf BUF1 (N2054, N2050);
nand NAND3 (N2055, N2053, N870, N476);
xor XOR2 (N2056, N2035, N82);
or OR4 (N2057, N2054, N1184, N1787, N295);
or OR4 (N2058, N2057, N448, N432, N886);
nand NAND3 (N2059, N2056, N1846, N1180);
xor XOR2 (N2060, N2051, N1110);
buf BUF1 (N2061, N2042);
and AND3 (N2062, N2010, N1697, N1237);
not NOT1 (N2063, N2062);
or OR4 (N2064, N2041, N2013, N454, N1512);
nand NAND4 (N2065, N2059, N1177, N900, N1508);
or OR4 (N2066, N2052, N1263, N532, N194);
buf BUF1 (N2067, N2055);
xor XOR2 (N2068, N2067, N338);
nand NAND2 (N2069, N2064, N440);
not NOT1 (N2070, N2068);
buf BUF1 (N2071, N2061);
nand NAND3 (N2072, N2071, N1383, N201);
or OR2 (N2073, N2047, N189);
nand NAND2 (N2074, N2073, N802);
buf BUF1 (N2075, N2069);
buf BUF1 (N2076, N2058);
buf BUF1 (N2077, N2065);
or OR2 (N2078, N2049, N1025);
buf BUF1 (N2079, N2075);
buf BUF1 (N2080, N2079);
and AND3 (N2081, N2070, N1468, N211);
nor NOR3 (N2082, N2066, N557, N1897);
or OR3 (N2083, N2076, N1130, N185);
not NOT1 (N2084, N2063);
buf BUF1 (N2085, N2072);
xor XOR2 (N2086, N2082, N480);
nor NOR2 (N2087, N2077, N528);
nor NOR4 (N2088, N2084, N1505, N787, N951);
nand NAND4 (N2089, N2080, N1575, N1021, N368);
buf BUF1 (N2090, N2088);
not NOT1 (N2091, N2060);
not NOT1 (N2092, N2089);
xor XOR2 (N2093, N2078, N744);
nand NAND4 (N2094, N2083, N1312, N1938, N1191);
or OR4 (N2095, N2091, N1374, N275, N326);
or OR4 (N2096, N2095, N1103, N2094, N1100);
and AND2 (N2097, N1274, N1900);
buf BUF1 (N2098, N2074);
or OR2 (N2099, N2086, N1307);
nor NOR4 (N2100, N2092, N1647, N911, N1663);
nor NOR2 (N2101, N2099, N156);
and AND4 (N2102, N2098, N1805, N870, N1897);
nand NAND2 (N2103, N2102, N1189);
or OR3 (N2104, N2100, N1540, N1350);
nor NOR3 (N2105, N2093, N1397, N1158);
nor NOR2 (N2106, N2085, N1809);
buf BUF1 (N2107, N2103);
xor XOR2 (N2108, N2107, N1057);
buf BUF1 (N2109, N2101);
or OR4 (N2110, N2081, N1476, N1091, N1479);
not NOT1 (N2111, N2096);
nand NAND2 (N2112, N2106, N1308);
nor NOR2 (N2113, N2112, N1650);
nor NOR4 (N2114, N2113, N1465, N887, N1005);
nor NOR4 (N2115, N2090, N1687, N1630, N1276);
nand NAND2 (N2116, N2097, N812);
not NOT1 (N2117, N2110);
not NOT1 (N2118, N2104);
and AND3 (N2119, N2111, N79, N1226);
not NOT1 (N2120, N2118);
and AND3 (N2121, N2114, N1150, N1458);
or OR4 (N2122, N2120, N1884, N908, N1410);
nor NOR3 (N2123, N2109, N1541, N837);
nand NAND4 (N2124, N2116, N266, N716, N156);
and AND2 (N2125, N2122, N1582);
not NOT1 (N2126, N2121);
xor XOR2 (N2127, N2125, N451);
nand NAND4 (N2128, N2108, N2093, N96, N2067);
buf BUF1 (N2129, N2117);
buf BUF1 (N2130, N2129);
or OR4 (N2131, N2087, N1960, N1499, N406);
buf BUF1 (N2132, N2128);
nand NAND2 (N2133, N2126, N320);
nor NOR4 (N2134, N2130, N1847, N682, N871);
xor XOR2 (N2135, N2115, N136);
xor XOR2 (N2136, N2134, N134);
nor NOR3 (N2137, N2133, N1348, N1799);
or OR4 (N2138, N2135, N742, N685, N585);
nand NAND4 (N2139, N2124, N1380, N1373, N770);
not NOT1 (N2140, N2132);
xor XOR2 (N2141, N2105, N697);
nand NAND4 (N2142, N2119, N1476, N373, N1681);
xor XOR2 (N2143, N2142, N560);
nor NOR4 (N2144, N2141, N1330, N1382, N528);
nor NOR3 (N2145, N2136, N763, N762);
nand NAND4 (N2146, N2143, N577, N1143, N2013);
or OR3 (N2147, N2139, N775, N221);
or OR2 (N2148, N2131, N618);
nand NAND4 (N2149, N2147, N568, N1830, N1858);
nand NAND3 (N2150, N2137, N1777, N514);
not NOT1 (N2151, N2150);
or OR3 (N2152, N2144, N744, N18);
nor NOR2 (N2153, N2149, N1593);
buf BUF1 (N2154, N2153);
nor NOR4 (N2155, N2151, N1431, N856, N1603);
not NOT1 (N2156, N2138);
nand NAND4 (N2157, N2156, N1455, N1537, N515);
buf BUF1 (N2158, N2123);
nand NAND4 (N2159, N2140, N2100, N553, N678);
nand NAND2 (N2160, N2152, N1322);
nor NOR4 (N2161, N2127, N69, N597, N1423);
buf BUF1 (N2162, N2158);
nor NOR4 (N2163, N2162, N1687, N809, N700);
or OR3 (N2164, N2154, N954, N214);
buf BUF1 (N2165, N2164);
nor NOR3 (N2166, N2146, N513, N1132);
xor XOR2 (N2167, N2148, N2114);
or OR3 (N2168, N2157, N1513, N2138);
xor XOR2 (N2169, N2167, N740);
and AND3 (N2170, N2165, N1395, N1899);
nor NOR4 (N2171, N2163, N1293, N1960, N1159);
buf BUF1 (N2172, N2161);
xor XOR2 (N2173, N2169, N1109);
buf BUF1 (N2174, N2172);
and AND3 (N2175, N2160, N207, N444);
or OR2 (N2176, N2170, N1195);
buf BUF1 (N2177, N2166);
not NOT1 (N2178, N2175);
xor XOR2 (N2179, N2145, N636);
nor NOR4 (N2180, N2177, N1687, N702, N1447);
and AND4 (N2181, N2171, N1063, N1270, N2070);
xor XOR2 (N2182, N2168, N1034);
not NOT1 (N2183, N2181);
nor NOR2 (N2184, N2178, N1011);
xor XOR2 (N2185, N2174, N1227);
buf BUF1 (N2186, N2159);
and AND4 (N2187, N2185, N810, N40, N1626);
nor NOR2 (N2188, N2155, N1876);
xor XOR2 (N2189, N2176, N1299);
nor NOR4 (N2190, N2186, N630, N1396, N1141);
or OR4 (N2191, N2184, N464, N1424, N1579);
nand NAND2 (N2192, N2191, N1030);
or OR4 (N2193, N2188, N667, N1432, N2022);
not NOT1 (N2194, N2183);
not NOT1 (N2195, N2182);
nand NAND3 (N2196, N2173, N2165, N424);
nand NAND4 (N2197, N2195, N703, N1967, N1904);
or OR3 (N2198, N2190, N206, N234);
and AND4 (N2199, N2179, N215, N1695, N1660);
and AND3 (N2200, N2197, N1072, N14);
buf BUF1 (N2201, N2198);
and AND3 (N2202, N2196, N1190, N659);
or OR2 (N2203, N2189, N287);
and AND4 (N2204, N2194, N925, N513, N1904);
or OR4 (N2205, N2202, N82, N1325, N2181);
nand NAND2 (N2206, N2203, N585);
nor NOR2 (N2207, N2201, N2034);
buf BUF1 (N2208, N2180);
buf BUF1 (N2209, N2205);
or OR4 (N2210, N2209, N178, N1298, N1430);
buf BUF1 (N2211, N2199);
nor NOR2 (N2212, N2204, N1901);
nand NAND4 (N2213, N2211, N1179, N1732, N1970);
xor XOR2 (N2214, N2213, N1886);
or OR2 (N2215, N2214, N217);
nand NAND3 (N2216, N2187, N206, N360);
buf BUF1 (N2217, N2208);
not NOT1 (N2218, N2212);
buf BUF1 (N2219, N2192);
xor XOR2 (N2220, N2216, N1646);
buf BUF1 (N2221, N2210);
and AND2 (N2222, N2215, N659);
buf BUF1 (N2223, N2220);
nor NOR4 (N2224, N2222, N109, N569, N221);
buf BUF1 (N2225, N2223);
xor XOR2 (N2226, N2193, N233);
nand NAND3 (N2227, N2221, N472, N50);
or OR2 (N2228, N2225, N1638);
buf BUF1 (N2229, N2200);
xor XOR2 (N2230, N2227, N1116);
xor XOR2 (N2231, N2228, N769);
nor NOR3 (N2232, N2230, N913, N23);
nor NOR2 (N2233, N2206, N1806);
buf BUF1 (N2234, N2224);
buf BUF1 (N2235, N2233);
nand NAND2 (N2236, N2219, N965);
xor XOR2 (N2237, N2226, N2003);
xor XOR2 (N2238, N2232, N534);
buf BUF1 (N2239, N2236);
nor NOR4 (N2240, N2229, N97, N463, N1834);
and AND2 (N2241, N2207, N1163);
not NOT1 (N2242, N2241);
nand NAND3 (N2243, N2235, N1735, N922);
or OR4 (N2244, N2234, N1134, N1021, N2185);
nor NOR2 (N2245, N2231, N1556);
nor NOR4 (N2246, N2217, N2067, N1387, N1887);
not NOT1 (N2247, N2238);
nand NAND4 (N2248, N2244, N166, N812, N2024);
xor XOR2 (N2249, N2248, N2104);
nor NOR2 (N2250, N2247, N2139);
not NOT1 (N2251, N2246);
nor NOR2 (N2252, N2250, N905);
or OR2 (N2253, N2239, N930);
not NOT1 (N2254, N2242);
nand NAND4 (N2255, N2243, N540, N1739, N2191);
buf BUF1 (N2256, N2240);
nor NOR2 (N2257, N2256, N242);
nor NOR2 (N2258, N2245, N2056);
nor NOR2 (N2259, N2252, N27);
not NOT1 (N2260, N2253);
xor XOR2 (N2261, N2259, N1452);
not NOT1 (N2262, N2249);
or OR4 (N2263, N2218, N970, N1321, N216);
not NOT1 (N2264, N2254);
or OR4 (N2265, N2258, N728, N2211, N1632);
nand NAND4 (N2266, N2260, N1247, N1328, N2020);
xor XOR2 (N2267, N2255, N467);
or OR4 (N2268, N2264, N487, N1167, N597);
buf BUF1 (N2269, N2265);
nor NOR2 (N2270, N2269, N795);
nand NAND4 (N2271, N2262, N992, N1703, N826);
nand NAND2 (N2272, N2257, N2109);
or OR3 (N2273, N2267, N2202, N1758);
or OR3 (N2274, N2261, N871, N888);
buf BUF1 (N2275, N2251);
or OR2 (N2276, N2273, N510);
or OR4 (N2277, N2271, N1648, N689, N353);
xor XOR2 (N2278, N2277, N2099);
buf BUF1 (N2279, N2270);
buf BUF1 (N2280, N2272);
nand NAND3 (N2281, N2278, N1356, N2192);
nor NOR3 (N2282, N2280, N1683, N907);
or OR3 (N2283, N2276, N1424, N1522);
not NOT1 (N2284, N2282);
nand NAND2 (N2285, N2274, N272);
xor XOR2 (N2286, N2275, N1276);
not NOT1 (N2287, N2266);
nor NOR3 (N2288, N2281, N749, N2057);
or OR4 (N2289, N2285, N530, N1250, N1613);
and AND4 (N2290, N2289, N1067, N987, N1481);
buf BUF1 (N2291, N2283);
not NOT1 (N2292, N2279);
nand NAND3 (N2293, N2291, N2257, N1869);
not NOT1 (N2294, N2286);
and AND4 (N2295, N2292, N1943, N662, N2264);
not NOT1 (N2296, N2288);
xor XOR2 (N2297, N2263, N1135);
and AND4 (N2298, N2284, N389, N125, N841);
xor XOR2 (N2299, N2296, N926);
and AND3 (N2300, N2290, N734, N1899);
xor XOR2 (N2301, N2237, N478);
buf BUF1 (N2302, N2298);
nand NAND4 (N2303, N2300, N1082, N1315, N205);
nand NAND3 (N2304, N2302, N1891, N1268);
nand NAND3 (N2305, N2299, N1205, N1855);
not NOT1 (N2306, N2295);
buf BUF1 (N2307, N2304);
xor XOR2 (N2308, N2301, N895);
xor XOR2 (N2309, N2287, N1184);
nor NOR2 (N2310, N2306, N1198);
and AND4 (N2311, N2303, N1590, N2017, N267);
and AND2 (N2312, N2305, N2156);
nand NAND3 (N2313, N2268, N852, N490);
buf BUF1 (N2314, N2293);
buf BUF1 (N2315, N2307);
buf BUF1 (N2316, N2315);
not NOT1 (N2317, N2309);
buf BUF1 (N2318, N2316);
or OR2 (N2319, N2317, N1323);
xor XOR2 (N2320, N2297, N1889);
buf BUF1 (N2321, N2318);
and AND4 (N2322, N2321, N551, N790, N2090);
or OR4 (N2323, N2310, N1069, N1953, N2130);
not NOT1 (N2324, N2314);
nand NAND3 (N2325, N2294, N835, N1642);
or OR2 (N2326, N2311, N502);
and AND3 (N2327, N2313, N1218, N1090);
xor XOR2 (N2328, N2320, N2206);
xor XOR2 (N2329, N2312, N1299);
and AND2 (N2330, N2319, N1398);
and AND4 (N2331, N2324, N332, N133, N1520);
nor NOR2 (N2332, N2308, N1085);
buf BUF1 (N2333, N2325);
not NOT1 (N2334, N2333);
nor NOR3 (N2335, N2332, N224, N42);
nor NOR3 (N2336, N2322, N2012, N1589);
and AND3 (N2337, N2336, N1890, N2171);
buf BUF1 (N2338, N2334);
nand NAND3 (N2339, N2323, N1887, N575);
buf BUF1 (N2340, N2327);
not NOT1 (N2341, N2329);
and AND3 (N2342, N2340, N1131, N1175);
or OR3 (N2343, N2331, N1711, N2035);
buf BUF1 (N2344, N2328);
nor NOR3 (N2345, N2343, N144, N905);
xor XOR2 (N2346, N2338, N2063);
nor NOR4 (N2347, N2344, N2291, N532, N232);
xor XOR2 (N2348, N2339, N68);
nor NOR3 (N2349, N2341, N1525, N687);
or OR4 (N2350, N2335, N218, N462, N1547);
or OR3 (N2351, N2326, N1389, N195);
xor XOR2 (N2352, N2348, N438);
nor NOR4 (N2353, N2347, N474, N147, N2074);
buf BUF1 (N2354, N2353);
not NOT1 (N2355, N2352);
or OR3 (N2356, N2350, N904, N867);
or OR3 (N2357, N2354, N1048, N2104);
nand NAND4 (N2358, N2345, N1134, N1014, N1528);
xor XOR2 (N2359, N2342, N350);
xor XOR2 (N2360, N2346, N981);
not NOT1 (N2361, N2349);
and AND3 (N2362, N2361, N2257, N743);
or OR4 (N2363, N2362, N717, N1165, N1312);
nand NAND3 (N2364, N2360, N1379, N1388);
not NOT1 (N2365, N2355);
and AND4 (N2366, N2351, N2085, N235, N1795);
buf BUF1 (N2367, N2364);
and AND3 (N2368, N2359, N1873, N433);
nor NOR2 (N2369, N2357, N2271);
and AND4 (N2370, N2363, N1301, N271, N2268);
buf BUF1 (N2371, N2366);
xor XOR2 (N2372, N2365, N2293);
not NOT1 (N2373, N2367);
nand NAND4 (N2374, N2358, N359, N1567, N2042);
and AND4 (N2375, N2374, N588, N2132, N577);
xor XOR2 (N2376, N2373, N1754);
nand NAND2 (N2377, N2375, N1982);
buf BUF1 (N2378, N2377);
nor NOR4 (N2379, N2330, N1664, N722, N492);
not NOT1 (N2380, N2376);
not NOT1 (N2381, N2368);
xor XOR2 (N2382, N2356, N1742);
nand NAND2 (N2383, N2370, N1585);
and AND4 (N2384, N2379, N1862, N1257, N1170);
and AND3 (N2385, N2383, N1109, N847);
buf BUF1 (N2386, N2372);
or OR2 (N2387, N2337, N2381);
xor XOR2 (N2388, N853, N883);
not NOT1 (N2389, N2378);
nand NAND2 (N2390, N2369, N1996);
and AND2 (N2391, N2384, N261);
nor NOR2 (N2392, N2380, N1011);
nand NAND2 (N2393, N2390, N487);
nor NOR3 (N2394, N2385, N1201, N2126);
buf BUF1 (N2395, N2382);
and AND2 (N2396, N2394, N2389);
nand NAND3 (N2397, N132, N1531, N2349);
or OR4 (N2398, N2392, N239, N2340, N982);
and AND2 (N2399, N2397, N280);
nand NAND3 (N2400, N2387, N1433, N1549);
nand NAND2 (N2401, N2398, N2357);
and AND3 (N2402, N2400, N1408, N316);
buf BUF1 (N2403, N2393);
and AND4 (N2404, N2371, N1528, N136, N1648);
nand NAND3 (N2405, N2402, N979, N2098);
not NOT1 (N2406, N2395);
xor XOR2 (N2407, N2391, N2258);
and AND4 (N2408, N2388, N722, N273, N1481);
or OR2 (N2409, N2401, N1212);
or OR3 (N2410, N2408, N133, N1185);
nor NOR4 (N2411, N2405, N662, N1138, N129);
or OR2 (N2412, N2399, N693);
nor NOR2 (N2413, N2406, N23);
buf BUF1 (N2414, N2404);
nand NAND4 (N2415, N2412, N1699, N1426, N2210);
nand NAND4 (N2416, N2410, N2403, N1587, N1637);
xor XOR2 (N2417, N624, N2073);
not NOT1 (N2418, N2415);
xor XOR2 (N2419, N2418, N1636);
or OR2 (N2420, N2386, N2300);
nor NOR2 (N2421, N2420, N941);
nand NAND3 (N2422, N2409, N402, N729);
and AND4 (N2423, N2416, N1348, N1373, N160);
and AND3 (N2424, N2417, N468, N289);
nor NOR2 (N2425, N2424, N1019);
or OR3 (N2426, N2421, N213, N855);
buf BUF1 (N2427, N2425);
nand NAND2 (N2428, N2427, N2086);
nor NOR3 (N2429, N2414, N746, N1241);
xor XOR2 (N2430, N2429, N1124);
xor XOR2 (N2431, N2430, N2395);
buf BUF1 (N2432, N2423);
xor XOR2 (N2433, N2422, N1335);
not NOT1 (N2434, N2426);
nor NOR2 (N2435, N2428, N1650);
buf BUF1 (N2436, N2407);
buf BUF1 (N2437, N2419);
nand NAND4 (N2438, N2432, N1315, N991, N516);
nand NAND4 (N2439, N2435, N1868, N1942, N2213);
buf BUF1 (N2440, N2436);
nor NOR2 (N2441, N2438, N2213);
xor XOR2 (N2442, N2437, N1474);
not NOT1 (N2443, N2431);
buf BUF1 (N2444, N2442);
nand NAND3 (N2445, N2411, N676, N1378);
not NOT1 (N2446, N2396);
xor XOR2 (N2447, N2439, N2307);
or OR2 (N2448, N2433, N1605);
not NOT1 (N2449, N2441);
buf BUF1 (N2450, N2447);
and AND2 (N2451, N2413, N2394);
not NOT1 (N2452, N2440);
xor XOR2 (N2453, N2448, N1653);
xor XOR2 (N2454, N2451, N729);
or OR4 (N2455, N2450, N1004, N775, N660);
and AND2 (N2456, N2454, N277);
or OR2 (N2457, N2434, N2127);
buf BUF1 (N2458, N2452);
nand NAND2 (N2459, N2453, N1641);
nand NAND4 (N2460, N2459, N1339, N973, N1768);
xor XOR2 (N2461, N2456, N1937);
buf BUF1 (N2462, N2445);
not NOT1 (N2463, N2462);
xor XOR2 (N2464, N2460, N1375);
nand NAND2 (N2465, N2457, N464);
not NOT1 (N2466, N2446);
nor NOR3 (N2467, N2463, N159, N1012);
buf BUF1 (N2468, N2466);
or OR2 (N2469, N2461, N1135);
buf BUF1 (N2470, N2464);
nand NAND3 (N2471, N2465, N79, N902);
xor XOR2 (N2472, N2458, N2409);
not NOT1 (N2473, N2468);
and AND3 (N2474, N2470, N2042, N2462);
and AND3 (N2475, N2472, N2110, N1044);
xor XOR2 (N2476, N2467, N2471);
not NOT1 (N2477, N2435);
buf BUF1 (N2478, N2449);
nand NAND2 (N2479, N2478, N233);
nand NAND4 (N2480, N2443, N182, N1782, N788);
buf BUF1 (N2481, N2480);
not NOT1 (N2482, N2476);
nor NOR4 (N2483, N2469, N2076, N2461, N40);
and AND2 (N2484, N2483, N1823);
not NOT1 (N2485, N2444);
or OR2 (N2486, N2481, N1462);
buf BUF1 (N2487, N2482);
nor NOR4 (N2488, N2477, N2156, N2429, N1904);
nor NOR4 (N2489, N2479, N498, N1566, N673);
buf BUF1 (N2490, N2485);
xor XOR2 (N2491, N2489, N2078);
xor XOR2 (N2492, N2455, N2223);
xor XOR2 (N2493, N2486, N1999);
nand NAND4 (N2494, N2474, N2219, N892, N390);
nor NOR2 (N2495, N2493, N2448);
and AND3 (N2496, N2487, N1143, N1625);
nor NOR3 (N2497, N2491, N1300, N426);
or OR2 (N2498, N2494, N350);
buf BUF1 (N2499, N2475);
not NOT1 (N2500, N2495);
not NOT1 (N2501, N2497);
and AND3 (N2502, N2473, N669, N838);
and AND4 (N2503, N2501, N286, N267, N1205);
nand NAND3 (N2504, N2492, N2090, N1620);
and AND2 (N2505, N2490, N1031);
nand NAND4 (N2506, N2499, N1503, N1333, N397);
buf BUF1 (N2507, N2488);
nand NAND3 (N2508, N2506, N69, N2265);
buf BUF1 (N2509, N2505);
nand NAND4 (N2510, N2508, N1670, N1736, N2408);
nor NOR3 (N2511, N2504, N1056, N2429);
not NOT1 (N2512, N2509);
xor XOR2 (N2513, N2498, N25);
not NOT1 (N2514, N2511);
nor NOR4 (N2515, N2513, N416, N1066, N1546);
or OR2 (N2516, N2510, N1965);
nand NAND2 (N2517, N2507, N1961);
and AND2 (N2518, N2502, N609);
and AND3 (N2519, N2484, N1758, N285);
xor XOR2 (N2520, N2512, N2005);
buf BUF1 (N2521, N2520);
not NOT1 (N2522, N2500);
or OR3 (N2523, N2517, N1003, N694);
nor NOR4 (N2524, N2522, N763, N306, N1384);
and AND4 (N2525, N2524, N1003, N73, N1279);
xor XOR2 (N2526, N2523, N383);
not NOT1 (N2527, N2521);
nor NOR2 (N2528, N2526, N1446);
or OR2 (N2529, N2503, N651);
and AND4 (N2530, N2527, N1186, N977, N2255);
xor XOR2 (N2531, N2525, N227);
not NOT1 (N2532, N2496);
not NOT1 (N2533, N2532);
not NOT1 (N2534, N2514);
or OR4 (N2535, N2519, N830, N913, N1937);
or OR3 (N2536, N2528, N284, N1191);
buf BUF1 (N2537, N2515);
xor XOR2 (N2538, N2518, N2386);
buf BUF1 (N2539, N2535);
nor NOR2 (N2540, N2533, N713);
or OR4 (N2541, N2531, N936, N960, N2344);
and AND3 (N2542, N2530, N837, N2061);
not NOT1 (N2543, N2536);
xor XOR2 (N2544, N2538, N2201);
not NOT1 (N2545, N2543);
or OR2 (N2546, N2529, N1027);
not NOT1 (N2547, N2544);
not NOT1 (N2548, N2542);
nand NAND2 (N2549, N2534, N2092);
and AND2 (N2550, N2540, N943);
xor XOR2 (N2551, N2545, N1236);
xor XOR2 (N2552, N2547, N67);
xor XOR2 (N2553, N2549, N483);
nor NOR3 (N2554, N2516, N2363, N350);
buf BUF1 (N2555, N2551);
xor XOR2 (N2556, N2550, N2489);
buf BUF1 (N2557, N2554);
and AND2 (N2558, N2537, N1223);
or OR4 (N2559, N2548, N167, N1563, N2001);
xor XOR2 (N2560, N2556, N448);
nor NOR2 (N2561, N2555, N2290);
xor XOR2 (N2562, N2558, N554);
or OR2 (N2563, N2562, N637);
buf BUF1 (N2564, N2552);
and AND2 (N2565, N2539, N2035);
nor NOR4 (N2566, N2565, N1938, N2457, N2433);
xor XOR2 (N2567, N2546, N140);
or OR2 (N2568, N2559, N2133);
nand NAND2 (N2569, N2564, N2525);
and AND4 (N2570, N2553, N1533, N559, N1187);
nor NOR4 (N2571, N2560, N2111, N1744, N1996);
buf BUF1 (N2572, N2563);
buf BUF1 (N2573, N2570);
or OR4 (N2574, N2567, N1947, N2365, N369);
not NOT1 (N2575, N2571);
nor NOR4 (N2576, N2561, N1971, N907, N1494);
xor XOR2 (N2577, N2566, N917);
and AND3 (N2578, N2573, N2020, N1252);
or OR3 (N2579, N2574, N1585, N2451);
buf BUF1 (N2580, N2572);
not NOT1 (N2581, N2575);
not NOT1 (N2582, N2577);
and AND2 (N2583, N2576, N131);
nor NOR4 (N2584, N2557, N1869, N1106, N323);
not NOT1 (N2585, N2578);
nand NAND2 (N2586, N2584, N1407);
buf BUF1 (N2587, N2583);
nor NOR2 (N2588, N2585, N1968);
or OR4 (N2589, N2541, N1948, N732, N1802);
nand NAND4 (N2590, N2579, N144, N1441, N150);
not NOT1 (N2591, N2587);
buf BUF1 (N2592, N2580);
nor NOR4 (N2593, N2582, N566, N2043, N1955);
nor NOR3 (N2594, N2593, N2320, N691);
xor XOR2 (N2595, N2592, N2280);
buf BUF1 (N2596, N2591);
nor NOR2 (N2597, N2569, N1110);
nand NAND3 (N2598, N2568, N2095, N2278);
buf BUF1 (N2599, N2595);
xor XOR2 (N2600, N2596, N1043);
not NOT1 (N2601, N2599);
or OR3 (N2602, N2590, N269, N180);
buf BUF1 (N2603, N2597);
xor XOR2 (N2604, N2602, N163);
not NOT1 (N2605, N2598);
and AND2 (N2606, N2594, N1711);
nand NAND2 (N2607, N2604, N2514);
or OR3 (N2608, N2588, N1905, N1625);
nand NAND4 (N2609, N2607, N1247, N1239, N2555);
not NOT1 (N2610, N2606);
xor XOR2 (N2611, N2586, N1033);
nand NAND2 (N2612, N2608, N2479);
nand NAND3 (N2613, N2609, N2081, N1759);
xor XOR2 (N2614, N2612, N1054);
xor XOR2 (N2615, N2613, N553);
or OR2 (N2616, N2603, N2614);
not NOT1 (N2617, N639);
buf BUF1 (N2618, N2610);
nand NAND4 (N2619, N2601, N2508, N1882, N1777);
nand NAND4 (N2620, N2618, N88, N309, N2537);
nand NAND3 (N2621, N2611, N1442, N699);
buf BUF1 (N2622, N2621);
xor XOR2 (N2623, N2622, N1795);
and AND2 (N2624, N2617, N275);
buf BUF1 (N2625, N2581);
and AND3 (N2626, N2616, N1528, N313);
or OR2 (N2627, N2624, N1442);
or OR3 (N2628, N2600, N771, N1308);
buf BUF1 (N2629, N2628);
xor XOR2 (N2630, N2625, N1391);
not NOT1 (N2631, N2589);
and AND2 (N2632, N2623, N388);
not NOT1 (N2633, N2619);
not NOT1 (N2634, N2627);
or OR4 (N2635, N2633, N749, N2406, N2091);
nand NAND2 (N2636, N2634, N889);
not NOT1 (N2637, N2632);
xor XOR2 (N2638, N2631, N1903);
not NOT1 (N2639, N2630);
nand NAND3 (N2640, N2635, N2377, N1960);
or OR2 (N2641, N2626, N1447);
buf BUF1 (N2642, N2637);
buf BUF1 (N2643, N2641);
and AND2 (N2644, N2643, N1919);
or OR4 (N2645, N2640, N1340, N1440, N246);
buf BUF1 (N2646, N2639);
nand NAND3 (N2647, N2636, N2544, N118);
nand NAND4 (N2648, N2647, N254, N405, N2066);
and AND2 (N2649, N2646, N776);
xor XOR2 (N2650, N2620, N538);
or OR2 (N2651, N2629, N1946);
and AND2 (N2652, N2605, N1852);
and AND4 (N2653, N2651, N889, N1159, N670);
not NOT1 (N2654, N2638);
or OR3 (N2655, N2653, N485, N1820);
buf BUF1 (N2656, N2650);
and AND2 (N2657, N2655, N999);
nor NOR2 (N2658, N2654, N7);
nand NAND4 (N2659, N2648, N97, N1413, N2520);
xor XOR2 (N2660, N2644, N2294);
buf BUF1 (N2661, N2659);
xor XOR2 (N2662, N2652, N1500);
buf BUF1 (N2663, N2657);
and AND2 (N2664, N2662, N2280);
or OR3 (N2665, N2661, N2002, N939);
not NOT1 (N2666, N2649);
and AND2 (N2667, N2666, N2573);
or OR3 (N2668, N2667, N994, N1048);
or OR4 (N2669, N2658, N1482, N2474, N2216);
xor XOR2 (N2670, N2669, N143);
buf BUF1 (N2671, N2660);
buf BUF1 (N2672, N2645);
buf BUF1 (N2673, N2642);
nand NAND4 (N2674, N2670, N1471, N2044, N341);
not NOT1 (N2675, N2674);
or OR2 (N2676, N2675, N589);
not NOT1 (N2677, N2671);
xor XOR2 (N2678, N2673, N2578);
nor NOR4 (N2679, N2665, N53, N2179, N1065);
or OR4 (N2680, N2679, N1825, N925, N481);
xor XOR2 (N2681, N2676, N2471);
nor NOR2 (N2682, N2664, N2119);
buf BUF1 (N2683, N2682);
not NOT1 (N2684, N2672);
nand NAND4 (N2685, N2678, N1266, N2013, N461);
nand NAND3 (N2686, N2615, N1113, N335);
and AND4 (N2687, N2656, N1241, N370, N2095);
and AND4 (N2688, N2677, N1378, N588, N921);
nor NOR3 (N2689, N2687, N2362, N1405);
nor NOR3 (N2690, N2663, N128, N2122);
not NOT1 (N2691, N2680);
not NOT1 (N2692, N2685);
nand NAND2 (N2693, N2692, N1283);
xor XOR2 (N2694, N2690, N2264);
or OR4 (N2695, N2689, N2382, N1153, N1302);
and AND2 (N2696, N2691, N2425);
and AND3 (N2697, N2695, N687, N480);
nor NOR3 (N2698, N2697, N1148, N945);
not NOT1 (N2699, N2698);
nor NOR4 (N2700, N2684, N1894, N212, N1178);
buf BUF1 (N2701, N2693);
buf BUF1 (N2702, N2683);
or OR2 (N2703, N2688, N1766);
xor XOR2 (N2704, N2686, N510);
nand NAND4 (N2705, N2703, N1736, N351, N1768);
nand NAND2 (N2706, N2668, N2334);
not NOT1 (N2707, N2681);
not NOT1 (N2708, N2694);
not NOT1 (N2709, N2707);
not NOT1 (N2710, N2708);
or OR2 (N2711, N2702, N2105);
nor NOR2 (N2712, N2709, N1616);
nor NOR3 (N2713, N2711, N823, N390);
buf BUF1 (N2714, N2700);
xor XOR2 (N2715, N2710, N2698);
nand NAND2 (N2716, N2715, N235);
buf BUF1 (N2717, N2716);
buf BUF1 (N2718, N2705);
and AND4 (N2719, N2718, N2347, N1201, N1192);
xor XOR2 (N2720, N2701, N516);
not NOT1 (N2721, N2714);
xor XOR2 (N2722, N2704, N1084);
xor XOR2 (N2723, N2706, N2558);
and AND2 (N2724, N2717, N1150);
or OR3 (N2725, N2696, N2599, N708);
not NOT1 (N2726, N2713);
xor XOR2 (N2727, N2699, N152);
nor NOR4 (N2728, N2720, N2408, N1589, N1151);
xor XOR2 (N2729, N2723, N379);
nand NAND4 (N2730, N2729, N1763, N970, N1853);
nor NOR2 (N2731, N2722, N1975);
nor NOR3 (N2732, N2724, N2703, N2560);
and AND4 (N2733, N2728, N509, N764, N2251);
not NOT1 (N2734, N2727);
and AND4 (N2735, N2725, N2207, N1520, N2139);
xor XOR2 (N2736, N2731, N2494);
nand NAND2 (N2737, N2719, N210);
nand NAND2 (N2738, N2721, N926);
not NOT1 (N2739, N2734);
not NOT1 (N2740, N2739);
xor XOR2 (N2741, N2737, N1095);
nor NOR4 (N2742, N2732, N1574, N836, N2220);
xor XOR2 (N2743, N2726, N422);
nor NOR4 (N2744, N2736, N2134, N947, N111);
nor NOR4 (N2745, N2738, N941, N1436, N1645);
nor NOR2 (N2746, N2745, N1848);
buf BUF1 (N2747, N2730);
not NOT1 (N2748, N2741);
not NOT1 (N2749, N2744);
and AND3 (N2750, N2740, N1367, N2457);
buf BUF1 (N2751, N2750);
nor NOR4 (N2752, N2743, N2309, N1384, N2340);
and AND4 (N2753, N2747, N1797, N1384, N69);
or OR3 (N2754, N2748, N749, N2324);
nor NOR4 (N2755, N2751, N2210, N1434, N1262);
or OR4 (N2756, N2749, N1046, N791, N2401);
or OR4 (N2757, N2752, N2284, N2048, N2506);
not NOT1 (N2758, N2756);
buf BUF1 (N2759, N2746);
nor NOR4 (N2760, N2735, N1929, N547, N1197);
nand NAND2 (N2761, N2742, N1209);
buf BUF1 (N2762, N2757);
buf BUF1 (N2763, N2762);
buf BUF1 (N2764, N2755);
not NOT1 (N2765, N2712);
and AND3 (N2766, N2759, N124, N2349);
not NOT1 (N2767, N2753);
buf BUF1 (N2768, N2767);
or OR2 (N2769, N2760, N2471);
and AND2 (N2770, N2764, N1475);
and AND4 (N2771, N2770, N674, N948, N1496);
and AND4 (N2772, N2758, N1290, N2699, N1153);
xor XOR2 (N2773, N2763, N1799);
not NOT1 (N2774, N2733);
buf BUF1 (N2775, N2765);
not NOT1 (N2776, N2766);
buf BUF1 (N2777, N2769);
nor NOR3 (N2778, N2761, N2102, N1330);
xor XOR2 (N2779, N2754, N311);
buf BUF1 (N2780, N2771);
nand NAND4 (N2781, N2778, N639, N1443, N960);
or OR4 (N2782, N2774, N1618, N1662, N367);
not NOT1 (N2783, N2775);
xor XOR2 (N2784, N2777, N754);
and AND3 (N2785, N2783, N981, N485);
nand NAND3 (N2786, N2768, N1832, N1241);
or OR3 (N2787, N2786, N155, N596);
or OR3 (N2788, N2785, N1981, N1249);
not NOT1 (N2789, N2781);
buf BUF1 (N2790, N2772);
xor XOR2 (N2791, N2776, N2702);
buf BUF1 (N2792, N2790);
and AND4 (N2793, N2787, N1083, N566, N1830);
or OR4 (N2794, N2773, N2671, N2447, N1234);
xor XOR2 (N2795, N2780, N2483);
and AND2 (N2796, N2792, N1358);
xor XOR2 (N2797, N2793, N170);
xor XOR2 (N2798, N2796, N2481);
not NOT1 (N2799, N2797);
nand NAND4 (N2800, N2795, N546, N2346, N429);
nand NAND4 (N2801, N2789, N1672, N881, N2575);
nand NAND2 (N2802, N2799, N137);
and AND4 (N2803, N2782, N609, N15, N2271);
nand NAND2 (N2804, N2800, N378);
not NOT1 (N2805, N2788);
not NOT1 (N2806, N2802);
xor XOR2 (N2807, N2798, N1021);
or OR2 (N2808, N2801, N1898);
buf BUF1 (N2809, N2804);
buf BUF1 (N2810, N2794);
buf BUF1 (N2811, N2808);
and AND2 (N2812, N2805, N2647);
and AND4 (N2813, N2779, N1875, N2084, N2501);
and AND3 (N2814, N2807, N1134, N27);
and AND4 (N2815, N2811, N2579, N1326, N888);
buf BUF1 (N2816, N2810);
and AND4 (N2817, N2814, N1918, N1318, N883);
or OR3 (N2818, N2813, N1016, N1235);
not NOT1 (N2819, N2816);
xor XOR2 (N2820, N2815, N645);
buf BUF1 (N2821, N2784);
and AND4 (N2822, N2820, N1098, N2061, N1611);
buf BUF1 (N2823, N2812);
not NOT1 (N2824, N2818);
xor XOR2 (N2825, N2803, N552);
buf BUF1 (N2826, N2791);
or OR3 (N2827, N2809, N2421, N2125);
buf BUF1 (N2828, N2821);
or OR2 (N2829, N2827, N746);
or OR4 (N2830, N2825, N1298, N1318, N34);
buf BUF1 (N2831, N2822);
nand NAND4 (N2832, N2817, N2080, N1957, N476);
nand NAND2 (N2833, N2831, N1323);
not NOT1 (N2834, N2828);
or OR2 (N2835, N2834, N1914);
xor XOR2 (N2836, N2806, N887);
nand NAND4 (N2837, N2832, N1060, N2792, N2484);
and AND4 (N2838, N2829, N2600, N1155, N683);
buf BUF1 (N2839, N2833);
xor XOR2 (N2840, N2826, N1089);
not NOT1 (N2841, N2838);
xor XOR2 (N2842, N2824, N1518);
nor NOR3 (N2843, N2830, N2564, N434);
or OR4 (N2844, N2823, N1008, N2731, N667);
and AND3 (N2845, N2842, N1480, N1159);
nand NAND4 (N2846, N2845, N1572, N654, N593);
nand NAND3 (N2847, N2840, N395, N2204);
and AND2 (N2848, N2835, N399);
xor XOR2 (N2849, N2837, N51);
nor NOR3 (N2850, N2841, N843, N897);
nand NAND3 (N2851, N2849, N2211, N76);
not NOT1 (N2852, N2819);
or OR4 (N2853, N2846, N2477, N2504, N194);
xor XOR2 (N2854, N2853, N434);
buf BUF1 (N2855, N2836);
not NOT1 (N2856, N2854);
and AND4 (N2857, N2843, N114, N1748, N542);
and AND2 (N2858, N2851, N23);
nand NAND4 (N2859, N2858, N1317, N1471, N2042);
and AND4 (N2860, N2855, N1142, N1213, N2031);
xor XOR2 (N2861, N2860, N2310);
buf BUF1 (N2862, N2839);
nand NAND2 (N2863, N2848, N805);
xor XOR2 (N2864, N2859, N1178);
xor XOR2 (N2865, N2857, N2114);
not NOT1 (N2866, N2847);
nand NAND4 (N2867, N2861, N2116, N823, N1816);
nand NAND2 (N2868, N2866, N2659);
not NOT1 (N2869, N2852);
nor NOR2 (N2870, N2869, N1784);
nor NOR3 (N2871, N2870, N1737, N1875);
buf BUF1 (N2872, N2868);
xor XOR2 (N2873, N2867, N260);
nor NOR2 (N2874, N2862, N1427);
buf BUF1 (N2875, N2872);
xor XOR2 (N2876, N2875, N1256);
not NOT1 (N2877, N2864);
not NOT1 (N2878, N2856);
nand NAND4 (N2879, N2878, N1043, N2146, N2155);
nand NAND2 (N2880, N2876, N2212);
nand NAND2 (N2881, N2865, N248);
xor XOR2 (N2882, N2877, N26);
xor XOR2 (N2883, N2871, N1933);
nor NOR2 (N2884, N2882, N1384);
not NOT1 (N2885, N2879);
nor NOR3 (N2886, N2885, N2783, N2306);
nand NAND4 (N2887, N2863, N1279, N286, N1059);
or OR3 (N2888, N2880, N173, N1073);
xor XOR2 (N2889, N2884, N422);
or OR2 (N2890, N2844, N149);
or OR2 (N2891, N2890, N2487);
not NOT1 (N2892, N2891);
and AND4 (N2893, N2888, N971, N2121, N14);
xor XOR2 (N2894, N2893, N2731);
nand NAND4 (N2895, N2887, N1376, N2083, N1028);
buf BUF1 (N2896, N2873);
or OR4 (N2897, N2894, N1778, N1726, N1777);
or OR4 (N2898, N2896, N1773, N1073, N2815);
buf BUF1 (N2899, N2850);
and AND2 (N2900, N2892, N865);
nand NAND2 (N2901, N2874, N826);
or OR4 (N2902, N2881, N2367, N839, N1626);
or OR4 (N2903, N2902, N2840, N1995, N1245);
and AND3 (N2904, N2895, N260, N560);
or OR3 (N2905, N2901, N1322, N2615);
nand NAND3 (N2906, N2883, N238, N641);
and AND4 (N2907, N2903, N476, N2431, N2603);
not NOT1 (N2908, N2904);
nand NAND2 (N2909, N2908, N1529);
xor XOR2 (N2910, N2886, N856);
not NOT1 (N2911, N2907);
and AND4 (N2912, N2906, N2446, N1137, N522);
nor NOR3 (N2913, N2905, N2853, N1339);
nor NOR2 (N2914, N2913, N101);
nor NOR2 (N2915, N2897, N1270);
nor NOR2 (N2916, N2911, N2237);
and AND2 (N2917, N2889, N1734);
not NOT1 (N2918, N2910);
or OR2 (N2919, N2900, N2265);
not NOT1 (N2920, N2909);
xor XOR2 (N2921, N2914, N275);
xor XOR2 (N2922, N2917, N1942);
nor NOR2 (N2923, N2919, N1518);
xor XOR2 (N2924, N2918, N2863);
nand NAND3 (N2925, N2921, N1025, N1858);
nand NAND4 (N2926, N2925, N2845, N2864, N1387);
buf BUF1 (N2927, N2899);
nor NOR4 (N2928, N2920, N2347, N1554, N271);
xor XOR2 (N2929, N2926, N892);
nor NOR3 (N2930, N2927, N1731, N556);
nor NOR2 (N2931, N2923, N1161);
xor XOR2 (N2932, N2915, N2583);
not NOT1 (N2933, N2912);
and AND3 (N2934, N2898, N1013, N113);
nand NAND3 (N2935, N2929, N636, N1131);
buf BUF1 (N2936, N2933);
xor XOR2 (N2937, N2924, N1459);
xor XOR2 (N2938, N2936, N33);
xor XOR2 (N2939, N2935, N157);
or OR3 (N2940, N2938, N1455, N1637);
xor XOR2 (N2941, N2930, N545);
nor NOR3 (N2942, N2931, N797, N145);
nor NOR3 (N2943, N2937, N1415, N2366);
not NOT1 (N2944, N2932);
nand NAND2 (N2945, N2944, N2284);
and AND4 (N2946, N2934, N1342, N1098, N1008);
or OR4 (N2947, N2943, N1719, N725, N2382);
buf BUF1 (N2948, N2945);
nor NOR3 (N2949, N2922, N1794, N271);
xor XOR2 (N2950, N2916, N2613);
nand NAND2 (N2951, N2939, N2407);
and AND4 (N2952, N2950, N483, N2496, N1128);
xor XOR2 (N2953, N2951, N2041);
nor NOR4 (N2954, N2953, N1192, N1372, N916);
nor NOR2 (N2955, N2946, N2327);
nor NOR3 (N2956, N2955, N1887, N261);
or OR2 (N2957, N2954, N1492);
and AND3 (N2958, N2940, N2305, N2104);
buf BUF1 (N2959, N2956);
xor XOR2 (N2960, N2947, N2900);
not NOT1 (N2961, N2959);
nand NAND3 (N2962, N2942, N938, N1474);
nor NOR4 (N2963, N2960, N232, N926, N2937);
and AND4 (N2964, N2952, N2322, N1890, N1743);
or OR2 (N2965, N2949, N2065);
nor NOR4 (N2966, N2962, N2233, N2570, N2047);
nand NAND4 (N2967, N2957, N837, N1842, N1248);
nor NOR2 (N2968, N2928, N375);
nor NOR4 (N2969, N2958, N8, N2327, N430);
nor NOR4 (N2970, N2965, N122, N2068, N158);
xor XOR2 (N2971, N2970, N1396);
not NOT1 (N2972, N2971);
nor NOR4 (N2973, N2941, N603, N2900, N268);
nor NOR2 (N2974, N2963, N2895);
nand NAND4 (N2975, N2964, N141, N1755, N2962);
nand NAND4 (N2976, N2966, N2341, N1439, N868);
buf BUF1 (N2977, N2967);
nand NAND3 (N2978, N2948, N538, N800);
buf BUF1 (N2979, N2974);
not NOT1 (N2980, N2975);
nor NOR2 (N2981, N2980, N1138);
nor NOR3 (N2982, N2961, N156, N2188);
buf BUF1 (N2983, N2973);
or OR4 (N2984, N2968, N12, N314, N330);
nand NAND3 (N2985, N2983, N331, N2091);
and AND3 (N2986, N2984, N2058, N758);
nor NOR2 (N2987, N2976, N1639);
and AND3 (N2988, N2969, N2129, N2237);
not NOT1 (N2989, N2987);
buf BUF1 (N2990, N2972);
xor XOR2 (N2991, N2981, N1498);
not NOT1 (N2992, N2989);
and AND3 (N2993, N2990, N1707, N1229);
xor XOR2 (N2994, N2992, N2675);
or OR2 (N2995, N2985, N429);
buf BUF1 (N2996, N2977);
or OR2 (N2997, N2996, N2695);
buf BUF1 (N2998, N2991);
xor XOR2 (N2999, N2978, N1277);
not NOT1 (N3000, N2994);
and AND3 (N3001, N2979, N2547, N2155);
xor XOR2 (N3002, N3000, N1264);
nor NOR4 (N3003, N3001, N1630, N621, N715);
xor XOR2 (N3004, N2999, N359);
buf BUF1 (N3005, N2998);
xor XOR2 (N3006, N3003, N681);
buf BUF1 (N3007, N3006);
or OR3 (N3008, N3002, N231, N1902);
nand NAND2 (N3009, N3004, N2449);
nand NAND4 (N3010, N2997, N1500, N153, N2610);
not NOT1 (N3011, N3009);
nand NAND2 (N3012, N2986, N2032);
endmodule