// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N279,N317,N314,N309,N316,N318,N306,N298,N310,N319;

not NOT1 (N20, N2);
buf BUF1 (N21, N6);
not NOT1 (N22, N12);
nand NAND2 (N23, N11, N16);
not NOT1 (N24, N18);
or OR3 (N25, N16, N16, N15);
nor NOR3 (N26, N10, N18, N15);
buf BUF1 (N27, N15);
and AND2 (N28, N7, N25);
nor NOR3 (N29, N14, N16, N10);
not NOT1 (N30, N19);
and AND4 (N31, N23, N18, N12, N26);
or OR2 (N32, N8, N8);
nand NAND4 (N33, N30, N10, N25, N6);
nor NOR3 (N34, N31, N25, N1);
nand NAND2 (N35, N28, N10);
nand NAND3 (N36, N29, N10, N18);
or OR4 (N37, N22, N32, N22, N29);
or OR4 (N38, N34, N20, N36, N29);
not NOT1 (N39, N9);
or OR4 (N40, N16, N17, N21, N4);
buf BUF1 (N41, N24);
not NOT1 (N42, N39);
not NOT1 (N43, N39);
nor NOR4 (N44, N16, N9, N38, N35);
buf BUF1 (N45, N44);
nor NOR2 (N46, N7, N21);
and AND4 (N47, N20, N40, N39, N27);
buf BUF1 (N48, N24);
and AND2 (N49, N10, N43);
xor XOR2 (N50, N36, N14);
not NOT1 (N51, N45);
nand NAND3 (N52, N41, N45, N25);
xor XOR2 (N53, N47, N27);
nor NOR4 (N54, N49, N6, N49, N53);
and AND2 (N55, N42, N33);
xor XOR2 (N56, N2, N24);
not NOT1 (N57, N26);
buf BUF1 (N58, N56);
nor NOR4 (N59, N46, N42, N12, N55);
and AND3 (N60, N54, N29, N27);
not NOT1 (N61, N41);
not NOT1 (N62, N37);
and AND2 (N63, N58, N29);
not NOT1 (N64, N52);
xor XOR2 (N65, N63, N60);
or OR4 (N66, N16, N34, N19, N34);
or OR4 (N67, N65, N59, N49, N6);
xor XOR2 (N68, N22, N58);
nor NOR2 (N69, N68, N56);
or OR4 (N70, N67, N7, N8, N65);
buf BUF1 (N71, N50);
or OR3 (N72, N64, N2, N38);
buf BUF1 (N73, N51);
buf BUF1 (N74, N73);
nor NOR4 (N75, N71, N57, N74, N22);
nor NOR3 (N76, N3, N53, N56);
not NOT1 (N77, N37);
nor NOR3 (N78, N77, N9, N17);
nand NAND2 (N79, N48, N13);
nor NOR4 (N80, N76, N58, N79, N21);
buf BUF1 (N81, N25);
and AND4 (N82, N81, N72, N41, N72);
nor NOR4 (N83, N39, N56, N79, N31);
nand NAND4 (N84, N66, N53, N1, N7);
nand NAND4 (N85, N80, N71, N47, N32);
buf BUF1 (N86, N69);
nand NAND4 (N87, N62, N2, N28, N84);
and AND4 (N88, N62, N40, N21, N58);
nand NAND2 (N89, N83, N2);
not NOT1 (N90, N70);
nand NAND2 (N91, N88, N69);
nor NOR4 (N92, N75, N28, N51, N37);
nor NOR4 (N93, N89, N14, N18, N20);
not NOT1 (N94, N87);
buf BUF1 (N95, N78);
not NOT1 (N96, N61);
nor NOR3 (N97, N90, N17, N45);
and AND3 (N98, N92, N93, N12);
xor XOR2 (N99, N70, N48);
nand NAND4 (N100, N95, N90, N79, N13);
or OR3 (N101, N98, N30, N83);
xor XOR2 (N102, N86, N57);
and AND2 (N103, N94, N35);
nand NAND3 (N104, N103, N72, N28);
not NOT1 (N105, N85);
not NOT1 (N106, N96);
nand NAND3 (N107, N91, N54, N51);
xor XOR2 (N108, N105, N8);
not NOT1 (N109, N104);
xor XOR2 (N110, N108, N66);
nor NOR4 (N111, N82, N54, N47, N56);
nand NAND3 (N112, N110, N97, N76);
nand NAND3 (N113, N97, N12, N30);
and AND2 (N114, N102, N109);
and AND3 (N115, N26, N99, N106);
and AND2 (N116, N9, N55);
xor XOR2 (N117, N18, N20);
or OR2 (N118, N113, N66);
nor NOR4 (N119, N100, N51, N98, N103);
xor XOR2 (N120, N116, N80);
buf BUF1 (N121, N120);
and AND4 (N122, N101, N78, N53, N11);
and AND4 (N123, N121, N22, N64, N19);
xor XOR2 (N124, N119, N91);
or OR2 (N125, N123, N44);
buf BUF1 (N126, N112);
nor NOR4 (N127, N122, N33, N43, N122);
not NOT1 (N128, N111);
xor XOR2 (N129, N107, N16);
not NOT1 (N130, N114);
nor NOR3 (N131, N125, N118, N65);
or OR2 (N132, N105, N6);
or OR4 (N133, N132, N53, N27, N39);
and AND4 (N134, N128, N98, N14, N28);
not NOT1 (N135, N126);
nand NAND3 (N136, N134, N80, N94);
or OR3 (N137, N115, N115, N3);
and AND3 (N138, N124, N34, N96);
buf BUF1 (N139, N136);
xor XOR2 (N140, N139, N98);
not NOT1 (N141, N138);
nand NAND3 (N142, N133, N20, N125);
not NOT1 (N143, N129);
and AND3 (N144, N130, N27, N17);
xor XOR2 (N145, N142, N72);
not NOT1 (N146, N127);
xor XOR2 (N147, N144, N7);
buf BUF1 (N148, N147);
buf BUF1 (N149, N137);
xor XOR2 (N150, N140, N117);
or OR4 (N151, N139, N40, N13, N113);
buf BUF1 (N152, N150);
nor NOR2 (N153, N151, N35);
or OR2 (N154, N131, N95);
nand NAND3 (N155, N154, N68, N14);
buf BUF1 (N156, N155);
or OR4 (N157, N146, N143, N145, N25);
or OR4 (N158, N91, N155, N143, N53);
and AND4 (N159, N124, N56, N152, N42);
buf BUF1 (N160, N8);
xor XOR2 (N161, N135, N83);
and AND4 (N162, N156, N59, N15, N139);
xor XOR2 (N163, N160, N125);
nor NOR2 (N164, N159, N37);
nand NAND4 (N165, N148, N37, N45, N144);
not NOT1 (N166, N158);
nand NAND2 (N167, N141, N158);
nor NOR2 (N168, N163, N67);
and AND2 (N169, N168, N37);
not NOT1 (N170, N161);
buf BUF1 (N171, N167);
or OR2 (N172, N165, N102);
not NOT1 (N173, N169);
nor NOR2 (N174, N166, N107);
nand NAND4 (N175, N174, N110, N53, N17);
buf BUF1 (N176, N157);
nor NOR2 (N177, N170, N120);
not NOT1 (N178, N153);
nand NAND2 (N179, N172, N87);
nand NAND4 (N180, N162, N6, N10, N175);
nand NAND3 (N181, N96, N130, N89);
or OR3 (N182, N179, N21, N55);
nand NAND2 (N183, N149, N122);
not NOT1 (N184, N173);
or OR2 (N185, N178, N138);
nor NOR4 (N186, N185, N21, N21, N112);
not NOT1 (N187, N184);
or OR4 (N188, N182, N142, N180, N138);
xor XOR2 (N189, N50, N157);
and AND3 (N190, N177, N109, N70);
nand NAND4 (N191, N181, N43, N149, N42);
not NOT1 (N192, N190);
nand NAND2 (N193, N186, N11);
nor NOR3 (N194, N171, N7, N132);
not NOT1 (N195, N194);
buf BUF1 (N196, N189);
or OR4 (N197, N188, N102, N186, N152);
nor NOR3 (N198, N164, N23, N197);
and AND4 (N199, N190, N187, N62, N128);
buf BUF1 (N200, N153);
or OR4 (N201, N195, N65, N87, N50);
nand NAND3 (N202, N199, N124, N192);
not NOT1 (N203, N14);
not NOT1 (N204, N198);
not NOT1 (N205, N183);
not NOT1 (N206, N203);
or OR2 (N207, N196, N100);
and AND4 (N208, N204, N119, N133, N207);
or OR2 (N209, N132, N187);
buf BUF1 (N210, N209);
and AND2 (N211, N176, N181);
xor XOR2 (N212, N200, N50);
nand NAND3 (N213, N201, N105, N203);
nand NAND2 (N214, N208, N44);
xor XOR2 (N215, N211, N25);
or OR3 (N216, N214, N53, N38);
xor XOR2 (N217, N210, N74);
buf BUF1 (N218, N212);
nand NAND3 (N219, N218, N166, N14);
nor NOR3 (N220, N213, N85, N138);
not NOT1 (N221, N220);
nor NOR3 (N222, N215, N51, N14);
or OR4 (N223, N205, N177, N189, N210);
and AND3 (N224, N221, N182, N125);
xor XOR2 (N225, N224, N10);
and AND3 (N226, N206, N205, N87);
not NOT1 (N227, N217);
nor NOR3 (N228, N191, N165, N4);
nand NAND4 (N229, N216, N39, N7, N222);
buf BUF1 (N230, N71);
nand NAND2 (N231, N229, N176);
not NOT1 (N232, N219);
xor XOR2 (N233, N225, N12);
or OR3 (N234, N193, N216, N17);
or OR4 (N235, N232, N76, N28, N143);
and AND2 (N236, N226, N211);
buf BUF1 (N237, N228);
and AND3 (N238, N230, N80, N80);
not NOT1 (N239, N238);
nand NAND2 (N240, N231, N205);
nand NAND3 (N241, N227, N109, N167);
buf BUF1 (N242, N202);
and AND4 (N243, N233, N61, N17, N153);
nand NAND4 (N244, N234, N141, N106, N126);
and AND3 (N245, N240, N195, N65);
xor XOR2 (N246, N223, N210);
nand NAND3 (N247, N243, N153, N39);
buf BUF1 (N248, N247);
nor NOR4 (N249, N239, N88, N146, N45);
nor NOR2 (N250, N249, N157);
buf BUF1 (N251, N241);
xor XOR2 (N252, N235, N119);
xor XOR2 (N253, N252, N153);
and AND4 (N254, N250, N155, N170, N200);
xor XOR2 (N255, N251, N203);
or OR3 (N256, N237, N197, N47);
nor NOR2 (N257, N244, N231);
xor XOR2 (N258, N245, N82);
nor NOR3 (N259, N255, N205, N103);
not NOT1 (N260, N253);
or OR2 (N261, N242, N65);
nor NOR4 (N262, N257, N193, N143, N196);
xor XOR2 (N263, N246, N119);
xor XOR2 (N264, N248, N232);
nor NOR3 (N265, N263, N179, N5);
and AND2 (N266, N258, N261);
not NOT1 (N267, N202);
nor NOR3 (N268, N262, N56, N225);
nor NOR3 (N269, N268, N173, N188);
not NOT1 (N270, N254);
and AND4 (N271, N267, N229, N72, N69);
and AND3 (N272, N260, N266, N220);
and AND2 (N273, N225, N207);
nor NOR2 (N274, N273, N68);
nor NOR3 (N275, N270, N55, N36);
xor XOR2 (N276, N274, N96);
xor XOR2 (N277, N265, N60);
and AND2 (N278, N271, N57);
xor XOR2 (N279, N278, N262);
buf BUF1 (N280, N276);
and AND3 (N281, N264, N60, N120);
or OR4 (N282, N275, N188, N12, N238);
xor XOR2 (N283, N269, N131);
nor NOR2 (N284, N281, N225);
and AND4 (N285, N256, N123, N75, N79);
not NOT1 (N286, N280);
buf BUF1 (N287, N285);
xor XOR2 (N288, N272, N107);
xor XOR2 (N289, N236, N211);
xor XOR2 (N290, N277, N205);
and AND3 (N291, N289, N21, N290);
buf BUF1 (N292, N29);
nor NOR3 (N293, N283, N269, N189);
nor NOR3 (N294, N288, N189, N140);
nand NAND2 (N295, N294, N20);
nor NOR4 (N296, N286, N15, N181, N133);
nand NAND4 (N297, N284, N44, N9, N162);
nand NAND4 (N298, N292, N76, N160, N34);
buf BUF1 (N299, N287);
or OR3 (N300, N259, N209, N112);
buf BUF1 (N301, N291);
nand NAND4 (N302, N295, N223, N106, N267);
buf BUF1 (N303, N296);
and AND3 (N304, N282, N239, N177);
and AND3 (N305, N299, N187, N58);
xor XOR2 (N306, N300, N302);
not NOT1 (N307, N2);
or OR2 (N308, N297, N270);
not NOT1 (N309, N307);
buf BUF1 (N310, N304);
nand NAND4 (N311, N303, N305, N145, N148);
xor XOR2 (N312, N105, N163);
not NOT1 (N313, N293);
buf BUF1 (N314, N312);
nand NAND3 (N315, N308, N162, N295);
not NOT1 (N316, N315);
nand NAND2 (N317, N301, N10);
or OR4 (N318, N311, N19, N182, N109);
buf BUF1 (N319, N313);
endmodule