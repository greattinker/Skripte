// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N3517,N3515,N3520,N3519,N3518,N3498,N3513,N3511,N3509,N3521;

buf BUF1 (N22, N9);
and AND3 (N23, N16, N22, N4);
not NOT1 (N24, N5);
or OR4 (N25, N19, N16, N12, N17);
not NOT1 (N26, N8);
nand NAND4 (N27, N19, N19, N9, N20);
buf BUF1 (N28, N11);
xor XOR2 (N29, N20, N18);
nor NOR4 (N30, N26, N8, N14, N22);
xor XOR2 (N31, N26, N16);
not NOT1 (N32, N20);
nor NOR4 (N33, N28, N13, N4, N8);
or OR4 (N34, N31, N8, N17, N16);
xor XOR2 (N35, N19, N30);
buf BUF1 (N36, N23);
buf BUF1 (N37, N29);
not NOT1 (N38, N1);
or OR4 (N39, N37, N33, N13, N26);
nor NOR4 (N40, N11, N28, N22, N8);
nand NAND3 (N41, N25, N16, N15);
buf BUF1 (N42, N41);
or OR2 (N43, N40, N19);
xor XOR2 (N44, N38, N19);
or OR4 (N45, N36, N14, N20, N44);
not NOT1 (N46, N21);
or OR3 (N47, N42, N37, N13);
buf BUF1 (N48, N27);
xor XOR2 (N49, N43, N47);
or OR3 (N50, N6, N24, N26);
nor NOR2 (N51, N43, N30);
or OR3 (N52, N45, N30, N9);
xor XOR2 (N53, N46, N43);
xor XOR2 (N54, N34, N12);
or OR2 (N55, N50, N30);
or OR4 (N56, N49, N45, N46, N32);
buf BUF1 (N57, N55);
buf BUF1 (N58, N10);
and AND3 (N59, N53, N12, N31);
nor NOR4 (N60, N48, N57, N35, N2);
nor NOR3 (N61, N50, N47, N48);
or OR4 (N62, N55, N4, N22, N28);
xor XOR2 (N63, N56, N58);
not NOT1 (N64, N42);
or OR2 (N65, N61, N25);
nand NAND4 (N66, N54, N44, N19, N13);
and AND4 (N67, N66, N36, N62, N16);
and AND4 (N68, N48, N34, N21, N57);
nor NOR2 (N69, N63, N46);
and AND2 (N70, N65, N56);
nor NOR4 (N71, N52, N45, N64, N57);
and AND4 (N72, N65, N69, N35, N71);
nand NAND3 (N73, N24, N58, N64);
and AND4 (N74, N55, N24, N31, N3);
xor XOR2 (N75, N39, N4);
buf BUF1 (N76, N73);
and AND2 (N77, N60, N13);
and AND3 (N78, N70, N14, N26);
not NOT1 (N79, N51);
nor NOR4 (N80, N74, N60, N57, N18);
or OR4 (N81, N79, N40, N60, N13);
nand NAND2 (N82, N68, N61);
nand NAND4 (N83, N77, N14, N50, N33);
nand NAND3 (N84, N72, N57, N19);
buf BUF1 (N85, N82);
not NOT1 (N86, N81);
xor XOR2 (N87, N86, N52);
xor XOR2 (N88, N84, N44);
buf BUF1 (N89, N76);
or OR4 (N90, N67, N70, N79, N70);
nor NOR3 (N91, N90, N1, N28);
buf BUF1 (N92, N75);
or OR3 (N93, N85, N35, N77);
buf BUF1 (N94, N83);
nand NAND4 (N95, N87, N94, N72, N79);
or OR2 (N96, N25, N63);
xor XOR2 (N97, N78, N87);
and AND2 (N98, N97, N47);
and AND3 (N99, N93, N51, N83);
buf BUF1 (N100, N89);
nand NAND4 (N101, N98, N82, N15, N79);
buf BUF1 (N102, N92);
and AND3 (N103, N59, N22, N89);
xor XOR2 (N104, N103, N96);
or OR3 (N105, N79, N44, N51);
not NOT1 (N106, N91);
not NOT1 (N107, N102);
nor NOR3 (N108, N100, N78, N69);
nand NAND2 (N109, N104, N71);
not NOT1 (N110, N99);
nand NAND2 (N111, N109, N49);
and AND3 (N112, N95, N13, N105);
nor NOR4 (N113, N54, N13, N45, N61);
buf BUF1 (N114, N101);
and AND3 (N115, N80, N71, N103);
nor NOR2 (N116, N113, N111);
xor XOR2 (N117, N10, N91);
or OR4 (N118, N115, N112, N43, N93);
xor XOR2 (N119, N24, N73);
nor NOR4 (N120, N117, N87, N79, N67);
nand NAND4 (N121, N110, N92, N57, N4);
nor NOR4 (N122, N88, N19, N58, N49);
not NOT1 (N123, N106);
not NOT1 (N124, N120);
nor NOR4 (N125, N119, N72, N40, N36);
not NOT1 (N126, N108);
and AND3 (N127, N122, N16, N80);
not NOT1 (N128, N126);
nor NOR2 (N129, N116, N128);
xor XOR2 (N130, N1, N72);
buf BUF1 (N131, N107);
or OR2 (N132, N125, N85);
buf BUF1 (N133, N127);
xor XOR2 (N134, N121, N102);
buf BUF1 (N135, N123);
nor NOR4 (N136, N124, N64, N106, N1);
and AND4 (N137, N134, N129, N124, N89);
or OR4 (N138, N13, N94, N67, N118);
or OR4 (N139, N96, N21, N70, N103);
nor NOR3 (N140, N131, N36, N29);
nor NOR3 (N141, N137, N139, N37);
and AND4 (N142, N124, N123, N64, N8);
not NOT1 (N143, N140);
xor XOR2 (N144, N132, N135);
not NOT1 (N145, N61);
xor XOR2 (N146, N142, N72);
and AND4 (N147, N114, N28, N122, N81);
or OR2 (N148, N133, N46);
xor XOR2 (N149, N147, N85);
and AND3 (N150, N138, N81, N60);
xor XOR2 (N151, N150, N98);
or OR4 (N152, N146, N86, N18, N80);
buf BUF1 (N153, N151);
nand NAND2 (N154, N145, N29);
buf BUF1 (N155, N148);
and AND3 (N156, N143, N6, N21);
not NOT1 (N157, N141);
nand NAND3 (N158, N149, N149, N26);
nor NOR3 (N159, N156, N100, N131);
nand NAND4 (N160, N159, N156, N66, N147);
not NOT1 (N161, N157);
not NOT1 (N162, N158);
xor XOR2 (N163, N144, N34);
nor NOR2 (N164, N162, N145);
not NOT1 (N165, N154);
nor NOR3 (N166, N163, N77, N65);
and AND3 (N167, N130, N129, N114);
nand NAND4 (N168, N153, N73, N157, N142);
and AND4 (N169, N168, N30, N126, N33);
buf BUF1 (N170, N155);
nor NOR3 (N171, N152, N103, N110);
not NOT1 (N172, N160);
or OR3 (N173, N136, N137, N4);
nor NOR2 (N174, N164, N6);
and AND4 (N175, N173, N174, N19, N33);
nor NOR2 (N176, N25, N90);
nor NOR3 (N177, N170, N7, N137);
or OR4 (N178, N171, N155, N38, N124);
not NOT1 (N179, N161);
and AND4 (N180, N165, N169, N93, N166);
xor XOR2 (N181, N129, N28);
or OR4 (N182, N170, N82, N161, N165);
and AND3 (N183, N177, N91, N5);
and AND3 (N184, N183, N72, N72);
nand NAND2 (N185, N182, N155);
buf BUF1 (N186, N167);
nand NAND4 (N187, N176, N133, N98, N122);
and AND3 (N188, N172, N18, N184);
nor NOR2 (N189, N97, N5);
nor NOR4 (N190, N188, N158, N48, N74);
xor XOR2 (N191, N179, N172);
not NOT1 (N192, N181);
nor NOR4 (N193, N192, N118, N75, N30);
nand NAND2 (N194, N175, N176);
nor NOR4 (N195, N180, N29, N150, N12);
and AND4 (N196, N185, N33, N25, N194);
and AND3 (N197, N85, N107, N96);
not NOT1 (N198, N187);
buf BUF1 (N199, N198);
not NOT1 (N200, N178);
or OR3 (N201, N200, N97, N132);
nor NOR3 (N202, N196, N170, N1);
and AND4 (N203, N193, N107, N187, N25);
xor XOR2 (N204, N203, N135);
xor XOR2 (N205, N195, N104);
nand NAND4 (N206, N201, N156, N169, N113);
xor XOR2 (N207, N190, N201);
nand NAND4 (N208, N202, N187, N43, N106);
or OR3 (N209, N206, N120, N171);
and AND3 (N210, N186, N59, N189);
not NOT1 (N211, N82);
nor NOR2 (N212, N207, N109);
nand NAND3 (N213, N205, N59, N63);
not NOT1 (N214, N210);
nor NOR3 (N215, N191, N29, N17);
buf BUF1 (N216, N204);
buf BUF1 (N217, N199);
not NOT1 (N218, N214);
buf BUF1 (N219, N216);
or OR2 (N220, N219, N77);
not NOT1 (N221, N212);
or OR2 (N222, N221, N111);
nand NAND4 (N223, N220, N141, N61, N70);
or OR2 (N224, N213, N151);
not NOT1 (N225, N222);
buf BUF1 (N226, N215);
and AND3 (N227, N218, N56, N179);
buf BUF1 (N228, N227);
nor NOR2 (N229, N209, N71);
nor NOR4 (N230, N225, N142, N35, N2);
buf BUF1 (N231, N208);
xor XOR2 (N232, N230, N4);
nor NOR2 (N233, N228, N33);
nand NAND2 (N234, N232, N144);
buf BUF1 (N235, N226);
or OR3 (N236, N229, N20, N113);
nand NAND2 (N237, N233, N117);
and AND4 (N238, N235, N99, N61, N98);
buf BUF1 (N239, N234);
xor XOR2 (N240, N211, N73);
xor XOR2 (N241, N197, N39);
buf BUF1 (N242, N238);
not NOT1 (N243, N217);
nor NOR3 (N244, N223, N167, N127);
not NOT1 (N245, N243);
buf BUF1 (N246, N236);
or OR4 (N247, N246, N123, N81, N193);
nor NOR2 (N248, N247, N214);
nand NAND3 (N249, N224, N31, N46);
xor XOR2 (N250, N248, N222);
buf BUF1 (N251, N242);
nor NOR3 (N252, N241, N18, N49);
not NOT1 (N253, N239);
buf BUF1 (N254, N237);
and AND4 (N255, N253, N57, N80, N137);
and AND3 (N256, N249, N114, N48);
buf BUF1 (N257, N240);
and AND4 (N258, N251, N187, N129, N31);
buf BUF1 (N259, N256);
buf BUF1 (N260, N259);
buf BUF1 (N261, N255);
or OR3 (N262, N258, N116, N5);
nor NOR4 (N263, N254, N230, N37, N213);
and AND4 (N264, N261, N226, N159, N99);
or OR2 (N265, N262, N192);
not NOT1 (N266, N265);
buf BUF1 (N267, N252);
or OR2 (N268, N257, N24);
nand NAND3 (N269, N263, N87, N243);
not NOT1 (N270, N267);
or OR3 (N271, N244, N231, N136);
nor NOR2 (N272, N249, N248);
or OR3 (N273, N272, N191, N129);
xor XOR2 (N274, N270, N215);
buf BUF1 (N275, N260);
nand NAND3 (N276, N250, N169, N10);
buf BUF1 (N277, N269);
and AND4 (N278, N268, N83, N211, N179);
and AND3 (N279, N273, N8, N258);
or OR3 (N280, N264, N81, N62);
buf BUF1 (N281, N279);
buf BUF1 (N282, N278);
xor XOR2 (N283, N275, N23);
not NOT1 (N284, N280);
nor NOR2 (N285, N276, N140);
or OR2 (N286, N266, N45);
and AND4 (N287, N274, N284, N230, N3);
xor XOR2 (N288, N134, N255);
nor NOR2 (N289, N286, N100);
xor XOR2 (N290, N245, N14);
xor XOR2 (N291, N290, N243);
not NOT1 (N292, N288);
or OR3 (N293, N289, N51, N164);
buf BUF1 (N294, N285);
or OR2 (N295, N291, N241);
nor NOR4 (N296, N277, N98, N20, N150);
xor XOR2 (N297, N294, N282);
nor NOR2 (N298, N221, N65);
xor XOR2 (N299, N292, N220);
not NOT1 (N300, N271);
nand NAND4 (N301, N287, N298, N148, N228);
or OR3 (N302, N83, N15, N243);
nand NAND3 (N303, N293, N143, N74);
nand NAND2 (N304, N302, N187);
not NOT1 (N305, N296);
buf BUF1 (N306, N304);
and AND4 (N307, N297, N178, N211, N235);
or OR4 (N308, N303, N50, N250, N175);
nor NOR4 (N309, N299, N240, N187, N49);
and AND4 (N310, N308, N79, N58, N51);
buf BUF1 (N311, N310);
xor XOR2 (N312, N300, N280);
buf BUF1 (N313, N307);
buf BUF1 (N314, N283);
xor XOR2 (N315, N281, N11);
or OR4 (N316, N315, N200, N268, N49);
not NOT1 (N317, N311);
and AND2 (N318, N314, N294);
nor NOR3 (N319, N301, N276, N195);
buf BUF1 (N320, N316);
or OR3 (N321, N312, N174, N199);
not NOT1 (N322, N295);
not NOT1 (N323, N319);
and AND4 (N324, N305, N177, N268, N132);
and AND2 (N325, N318, N86);
xor XOR2 (N326, N323, N266);
or OR4 (N327, N320, N196, N302, N268);
buf BUF1 (N328, N309);
or OR4 (N329, N313, N97, N272, N256);
nand NAND4 (N330, N317, N155, N303, N273);
not NOT1 (N331, N322);
not NOT1 (N332, N324);
buf BUF1 (N333, N321);
nand NAND3 (N334, N328, N269, N45);
xor XOR2 (N335, N334, N141);
or OR2 (N336, N332, N107);
buf BUF1 (N337, N333);
nand NAND3 (N338, N329, N318, N262);
and AND2 (N339, N338, N245);
xor XOR2 (N340, N337, N304);
buf BUF1 (N341, N331);
nand NAND3 (N342, N330, N306, N149);
nor NOR3 (N343, N176, N266, N291);
not NOT1 (N344, N326);
nor NOR4 (N345, N335, N310, N37, N220);
and AND2 (N346, N343, N331);
or OR4 (N347, N346, N41, N188, N138);
buf BUF1 (N348, N347);
or OR2 (N349, N344, N333);
xor XOR2 (N350, N325, N220);
nand NAND3 (N351, N348, N36, N21);
or OR2 (N352, N340, N80);
buf BUF1 (N353, N339);
nand NAND3 (N354, N352, N105, N28);
xor XOR2 (N355, N341, N299);
not NOT1 (N356, N349);
not NOT1 (N357, N355);
and AND2 (N358, N353, N279);
xor XOR2 (N359, N350, N144);
or OR2 (N360, N356, N269);
nand NAND3 (N361, N351, N11, N209);
nand NAND2 (N362, N354, N83);
nor NOR4 (N363, N327, N145, N50, N251);
nand NAND3 (N364, N360, N161, N316);
buf BUF1 (N365, N361);
not NOT1 (N366, N336);
xor XOR2 (N367, N366, N260);
nor NOR3 (N368, N365, N316, N323);
and AND2 (N369, N368, N189);
not NOT1 (N370, N357);
not NOT1 (N371, N345);
nor NOR2 (N372, N362, N350);
nand NAND3 (N373, N372, N115, N342);
or OR2 (N374, N321, N231);
xor XOR2 (N375, N371, N93);
or OR4 (N376, N367, N113, N357, N137);
nand NAND4 (N377, N369, N5, N175, N77);
or OR3 (N378, N370, N55, N140);
and AND3 (N379, N377, N28, N87);
nor NOR2 (N380, N359, N71);
nor NOR3 (N381, N376, N202, N208);
not NOT1 (N382, N363);
buf BUF1 (N383, N375);
nand NAND4 (N384, N373, N46, N261, N176);
and AND4 (N385, N383, N168, N243, N139);
xor XOR2 (N386, N380, N87);
not NOT1 (N387, N385);
and AND3 (N388, N378, N205, N206);
nand NAND4 (N389, N381, N20, N119, N57);
nand NAND2 (N390, N382, N154);
not NOT1 (N391, N386);
nor NOR2 (N392, N379, N72);
not NOT1 (N393, N384);
or OR4 (N394, N389, N127, N125, N171);
and AND2 (N395, N390, N193);
and AND2 (N396, N387, N16);
buf BUF1 (N397, N393);
and AND4 (N398, N358, N321, N324, N373);
and AND3 (N399, N392, N96, N40);
nand NAND2 (N400, N364, N169);
nand NAND4 (N401, N397, N218, N362, N28);
nor NOR3 (N402, N394, N368, N183);
not NOT1 (N403, N402);
or OR2 (N404, N399, N286);
and AND4 (N405, N403, N12, N218, N225);
nand NAND3 (N406, N398, N401, N164);
xor XOR2 (N407, N51, N41);
nand NAND2 (N408, N407, N139);
nand NAND4 (N409, N388, N286, N392, N86);
nand NAND4 (N410, N404, N326, N94, N202);
not NOT1 (N411, N391);
xor XOR2 (N412, N405, N145);
nor NOR4 (N413, N411, N190, N227, N262);
xor XOR2 (N414, N395, N199);
buf BUF1 (N415, N396);
buf BUF1 (N416, N406);
or OR2 (N417, N412, N3);
nand NAND4 (N418, N409, N70, N360, N110);
xor XOR2 (N419, N408, N390);
xor XOR2 (N420, N415, N415);
nor NOR4 (N421, N374, N194, N111, N175);
not NOT1 (N422, N420);
or OR4 (N423, N416, N382, N264, N285);
xor XOR2 (N424, N423, N88);
not NOT1 (N425, N418);
or OR3 (N426, N413, N33, N86);
and AND3 (N427, N425, N414, N256);
nor NOR4 (N428, N182, N175, N317, N166);
nand NAND3 (N429, N427, N48, N277);
not NOT1 (N430, N424);
or OR4 (N431, N400, N270, N298, N238);
nand NAND2 (N432, N419, N266);
not NOT1 (N433, N432);
nand NAND3 (N434, N410, N249, N424);
not NOT1 (N435, N417);
buf BUF1 (N436, N428);
and AND4 (N437, N426, N368, N118, N293);
xor XOR2 (N438, N436, N6);
nand NAND4 (N439, N429, N77, N118, N76);
nand NAND4 (N440, N433, N409, N205, N75);
xor XOR2 (N441, N421, N234);
nand NAND3 (N442, N440, N406, N211);
xor XOR2 (N443, N435, N7);
not NOT1 (N444, N438);
and AND4 (N445, N437, N352, N429, N164);
nor NOR3 (N446, N443, N264, N33);
not NOT1 (N447, N444);
nand NAND3 (N448, N434, N7, N117);
or OR2 (N449, N445, N317);
buf BUF1 (N450, N447);
and AND2 (N451, N446, N210);
not NOT1 (N452, N450);
not NOT1 (N453, N430);
xor XOR2 (N454, N451, N345);
nor NOR3 (N455, N422, N117, N103);
nand NAND4 (N456, N454, N170, N353, N92);
xor XOR2 (N457, N439, N220);
and AND4 (N458, N441, N284, N257, N121);
xor XOR2 (N459, N431, N198);
nand NAND3 (N460, N456, N107, N58);
xor XOR2 (N461, N455, N446);
not NOT1 (N462, N453);
nand NAND2 (N463, N449, N39);
nor NOR3 (N464, N463, N183, N224);
buf BUF1 (N465, N448);
or OR3 (N466, N465, N343, N66);
buf BUF1 (N467, N442);
or OR2 (N468, N452, N433);
not NOT1 (N469, N462);
xor XOR2 (N470, N464, N267);
and AND4 (N471, N469, N4, N416, N126);
buf BUF1 (N472, N458);
xor XOR2 (N473, N470, N407);
buf BUF1 (N474, N473);
or OR2 (N475, N474, N313);
not NOT1 (N476, N457);
buf BUF1 (N477, N460);
nor NOR3 (N478, N475, N114, N278);
nand NAND4 (N479, N472, N243, N406, N95);
buf BUF1 (N480, N471);
and AND3 (N481, N461, N271, N389);
or OR3 (N482, N481, N2, N153);
or OR4 (N483, N477, N287, N414, N328);
nor NOR2 (N484, N482, N467);
buf BUF1 (N485, N411);
not NOT1 (N486, N466);
not NOT1 (N487, N478);
or OR2 (N488, N459, N30);
xor XOR2 (N489, N484, N52);
and AND3 (N490, N488, N221, N92);
nand NAND4 (N491, N489, N72, N316, N436);
nand NAND4 (N492, N486, N304, N115, N374);
or OR4 (N493, N487, N14, N148, N275);
xor XOR2 (N494, N468, N290);
and AND4 (N495, N492, N327, N261, N241);
buf BUF1 (N496, N485);
not NOT1 (N497, N490);
xor XOR2 (N498, N494, N224);
buf BUF1 (N499, N493);
nor NOR2 (N500, N495, N162);
nand NAND3 (N501, N479, N177, N165);
nor NOR2 (N502, N491, N296);
xor XOR2 (N503, N502, N37);
or OR3 (N504, N499, N112, N443);
buf BUF1 (N505, N500);
or OR4 (N506, N505, N20, N129, N502);
buf BUF1 (N507, N504);
nand NAND4 (N508, N498, N316, N309, N268);
nor NOR3 (N509, N496, N46, N429);
buf BUF1 (N510, N480);
nand NAND2 (N511, N501, N137);
nor NOR4 (N512, N507, N476, N112, N308);
and AND4 (N513, N158, N167, N198, N26);
not NOT1 (N514, N509);
buf BUF1 (N515, N512);
buf BUF1 (N516, N483);
nor NOR3 (N517, N511, N516, N279);
buf BUF1 (N518, N185);
not NOT1 (N519, N518);
and AND2 (N520, N506, N177);
and AND2 (N521, N520, N102);
nand NAND2 (N522, N515, N285);
not NOT1 (N523, N522);
buf BUF1 (N524, N517);
not NOT1 (N525, N514);
or OR2 (N526, N524, N310);
nand NAND2 (N527, N508, N520);
nor NOR2 (N528, N526, N333);
xor XOR2 (N529, N528, N126);
nor NOR3 (N530, N529, N462, N339);
or OR3 (N531, N521, N264, N331);
xor XOR2 (N532, N530, N140);
or OR4 (N533, N527, N449, N425, N508);
or OR2 (N534, N519, N258);
nand NAND3 (N535, N523, N393, N175);
nand NAND2 (N536, N513, N400);
buf BUF1 (N537, N497);
or OR2 (N538, N503, N408);
or OR3 (N539, N531, N463, N238);
or OR3 (N540, N536, N425, N530);
or OR2 (N541, N525, N485);
nand NAND2 (N542, N534, N499);
nor NOR4 (N543, N540, N147, N300, N15);
and AND3 (N544, N541, N404, N532);
xor XOR2 (N545, N299, N451);
xor XOR2 (N546, N535, N219);
buf BUF1 (N547, N545);
not NOT1 (N548, N543);
or OR4 (N549, N537, N475, N8, N303);
buf BUF1 (N550, N539);
and AND3 (N551, N548, N406, N161);
nor NOR2 (N552, N542, N323);
buf BUF1 (N553, N552);
nand NAND2 (N554, N551, N65);
or OR3 (N555, N550, N306, N10);
not NOT1 (N556, N533);
nor NOR3 (N557, N556, N548, N118);
or OR4 (N558, N544, N207, N423, N294);
buf BUF1 (N559, N538);
or OR4 (N560, N510, N386, N403, N99);
nor NOR2 (N561, N553, N87);
not NOT1 (N562, N547);
nand NAND2 (N563, N562, N64);
or OR2 (N564, N559, N326);
xor XOR2 (N565, N560, N563);
buf BUF1 (N566, N212);
xor XOR2 (N567, N566, N279);
not NOT1 (N568, N555);
or OR3 (N569, N546, N568, N47);
nor NOR3 (N570, N462, N277, N259);
xor XOR2 (N571, N558, N429);
nor NOR2 (N572, N565, N7);
nor NOR2 (N573, N572, N381);
buf BUF1 (N574, N573);
buf BUF1 (N575, N561);
not NOT1 (N576, N549);
xor XOR2 (N577, N569, N137);
xor XOR2 (N578, N574, N4);
and AND3 (N579, N577, N496, N63);
or OR3 (N580, N576, N21, N506);
not NOT1 (N581, N579);
nand NAND3 (N582, N567, N165, N294);
and AND4 (N583, N557, N440, N241, N350);
or OR3 (N584, N570, N130, N441);
xor XOR2 (N585, N583, N316);
or OR2 (N586, N581, N402);
nand NAND3 (N587, N586, N555, N127);
buf BUF1 (N588, N587);
xor XOR2 (N589, N584, N233);
xor XOR2 (N590, N554, N583);
and AND4 (N591, N564, N54, N230, N221);
and AND3 (N592, N575, N98, N156);
not NOT1 (N593, N571);
buf BUF1 (N594, N580);
buf BUF1 (N595, N593);
not NOT1 (N596, N590);
nand NAND3 (N597, N595, N34, N61);
buf BUF1 (N598, N592);
xor XOR2 (N599, N596, N392);
nor NOR4 (N600, N598, N408, N539, N161);
nor NOR4 (N601, N582, N525, N574, N78);
or OR4 (N602, N585, N32, N591, N335);
or OR4 (N603, N304, N310, N432, N298);
and AND2 (N604, N578, N133);
nand NAND3 (N605, N588, N402, N132);
or OR4 (N606, N603, N234, N245, N557);
nand NAND4 (N607, N594, N166, N218, N543);
and AND4 (N608, N589, N460, N599, N114);
buf BUF1 (N609, N29);
nor NOR2 (N610, N607, N300);
nand NAND3 (N611, N610, N61, N508);
nand NAND2 (N612, N608, N101);
or OR2 (N613, N605, N202);
xor XOR2 (N614, N602, N241);
xor XOR2 (N615, N600, N539);
buf BUF1 (N616, N606);
nand NAND3 (N617, N604, N336, N601);
not NOT1 (N618, N355);
buf BUF1 (N619, N618);
nand NAND3 (N620, N613, N199, N351);
xor XOR2 (N621, N620, N518);
buf BUF1 (N622, N612);
or OR4 (N623, N615, N19, N152, N290);
or OR4 (N624, N609, N153, N255, N282);
buf BUF1 (N625, N611);
nand NAND4 (N626, N597, N368, N492, N543);
xor XOR2 (N627, N622, N312);
not NOT1 (N628, N616);
and AND3 (N629, N621, N325, N622);
not NOT1 (N630, N623);
and AND4 (N631, N626, N443, N287, N493);
or OR3 (N632, N628, N305, N600);
or OR3 (N633, N631, N327, N351);
nand NAND2 (N634, N627, N241);
nor NOR4 (N635, N633, N154, N585, N614);
buf BUF1 (N636, N76);
buf BUF1 (N637, N624);
not NOT1 (N638, N632);
buf BUF1 (N639, N619);
and AND3 (N640, N639, N213, N386);
not NOT1 (N641, N625);
xor XOR2 (N642, N638, N82);
not NOT1 (N643, N641);
not NOT1 (N644, N640);
nand NAND2 (N645, N617, N557);
nor NOR2 (N646, N635, N489);
not NOT1 (N647, N645);
buf BUF1 (N648, N646);
nand NAND2 (N649, N642, N50);
or OR3 (N650, N648, N266, N633);
nor NOR4 (N651, N634, N430, N67, N292);
and AND3 (N652, N644, N175, N21);
nand NAND4 (N653, N649, N470, N82, N100);
nand NAND3 (N654, N629, N26, N544);
or OR4 (N655, N643, N492, N151, N605);
and AND4 (N656, N647, N13, N478, N327);
or OR4 (N657, N656, N580, N436, N242);
nor NOR4 (N658, N650, N415, N329, N297);
or OR4 (N659, N636, N19, N247, N176);
nand NAND3 (N660, N637, N395, N319);
and AND3 (N661, N652, N58, N619);
not NOT1 (N662, N630);
xor XOR2 (N663, N658, N469);
or OR3 (N664, N657, N181, N72);
nor NOR2 (N665, N661, N50);
not NOT1 (N666, N653);
not NOT1 (N667, N666);
buf BUF1 (N668, N654);
not NOT1 (N669, N662);
and AND4 (N670, N665, N202, N402, N545);
nand NAND3 (N671, N651, N603, N458);
not NOT1 (N672, N663);
xor XOR2 (N673, N659, N282);
xor XOR2 (N674, N672, N26);
not NOT1 (N675, N660);
xor XOR2 (N676, N670, N349);
nor NOR3 (N677, N664, N561, N85);
not NOT1 (N678, N673);
nor NOR2 (N679, N669, N516);
nand NAND2 (N680, N678, N604);
nand NAND4 (N681, N655, N630, N656, N629);
or OR2 (N682, N675, N66);
nand NAND2 (N683, N682, N178);
and AND3 (N684, N668, N491, N627);
and AND3 (N685, N671, N43, N632);
nand NAND3 (N686, N679, N159, N451);
or OR3 (N687, N686, N637, N107);
buf BUF1 (N688, N674);
nand NAND2 (N689, N680, N596);
not NOT1 (N690, N677);
buf BUF1 (N691, N685);
nor NOR3 (N692, N667, N42, N309);
buf BUF1 (N693, N690);
buf BUF1 (N694, N692);
and AND2 (N695, N689, N380);
nor NOR2 (N696, N691, N177);
nand NAND3 (N697, N694, N613, N31);
xor XOR2 (N698, N681, N563);
buf BUF1 (N699, N695);
nand NAND3 (N700, N697, N449, N554);
buf BUF1 (N701, N699);
not NOT1 (N702, N684);
nor NOR2 (N703, N701, N201);
nand NAND2 (N704, N687, N97);
or OR4 (N705, N696, N236, N326, N44);
xor XOR2 (N706, N688, N506);
buf BUF1 (N707, N706);
nor NOR3 (N708, N702, N406, N420);
and AND3 (N709, N703, N282, N622);
nor NOR4 (N710, N707, N641, N323, N368);
and AND2 (N711, N683, N692);
and AND3 (N712, N705, N143, N216);
buf BUF1 (N713, N693);
xor XOR2 (N714, N709, N346);
buf BUF1 (N715, N710);
not NOT1 (N716, N708);
buf BUF1 (N717, N713);
nor NOR3 (N718, N704, N677, N571);
xor XOR2 (N719, N716, N379);
and AND4 (N720, N711, N492, N124, N431);
and AND4 (N721, N714, N92, N215, N389);
nor NOR3 (N722, N718, N105, N534);
nand NAND2 (N723, N700, N137);
nand NAND3 (N724, N721, N272, N382);
not NOT1 (N725, N720);
xor XOR2 (N726, N712, N387);
not NOT1 (N727, N722);
not NOT1 (N728, N717);
not NOT1 (N729, N676);
nand NAND4 (N730, N715, N310, N397, N127);
and AND3 (N731, N728, N296, N232);
not NOT1 (N732, N729);
and AND3 (N733, N732, N609, N491);
or OR3 (N734, N731, N437, N423);
and AND2 (N735, N698, N217);
xor XOR2 (N736, N724, N476);
nor NOR4 (N737, N730, N390, N404, N109);
nor NOR3 (N738, N723, N177, N662);
or OR2 (N739, N719, N64);
xor XOR2 (N740, N738, N730);
nand NAND4 (N741, N735, N477, N656, N196);
or OR4 (N742, N727, N626, N203, N295);
or OR4 (N743, N734, N249, N161, N393);
not NOT1 (N744, N743);
and AND2 (N745, N739, N702);
not NOT1 (N746, N741);
nor NOR2 (N747, N744, N610);
xor XOR2 (N748, N737, N557);
nand NAND2 (N749, N740, N141);
not NOT1 (N750, N726);
or OR4 (N751, N745, N353, N44, N443);
nand NAND4 (N752, N725, N203, N333, N685);
buf BUF1 (N753, N747);
nand NAND3 (N754, N752, N221, N289);
not NOT1 (N755, N749);
nand NAND2 (N756, N748, N665);
and AND4 (N757, N750, N486, N156, N547);
nor NOR4 (N758, N746, N125, N674, N361);
nand NAND3 (N759, N742, N76, N301);
or OR2 (N760, N758, N751);
nand NAND2 (N761, N227, N618);
nand NAND3 (N762, N736, N363, N718);
nor NOR2 (N763, N757, N296);
not NOT1 (N764, N760);
buf BUF1 (N765, N754);
nor NOR3 (N766, N764, N252, N473);
or OR2 (N767, N762, N302);
nand NAND4 (N768, N756, N415, N292, N245);
nor NOR4 (N769, N755, N74, N346, N203);
and AND4 (N770, N761, N622, N441, N725);
nand NAND3 (N771, N763, N633, N59);
not NOT1 (N772, N753);
buf BUF1 (N773, N772);
and AND3 (N774, N733, N726, N468);
buf BUF1 (N775, N770);
or OR4 (N776, N767, N567, N271, N573);
buf BUF1 (N777, N775);
or OR3 (N778, N773, N298, N500);
xor XOR2 (N779, N768, N285);
nand NAND2 (N780, N774, N90);
not NOT1 (N781, N759);
or OR4 (N782, N765, N338, N176, N88);
and AND4 (N783, N777, N325, N623, N467);
nor NOR4 (N784, N778, N125, N41, N685);
and AND3 (N785, N776, N661, N688);
nor NOR4 (N786, N783, N22, N785, N94);
or OR2 (N787, N786, N343);
and AND2 (N788, N249, N700);
or OR3 (N789, N782, N610, N722);
or OR2 (N790, N780, N402);
and AND2 (N791, N787, N441);
nand NAND4 (N792, N789, N282, N214, N774);
or OR3 (N793, N788, N2, N262);
or OR2 (N794, N792, N728);
nor NOR4 (N795, N766, N603, N343, N689);
nand NAND2 (N796, N771, N722);
xor XOR2 (N797, N779, N199);
and AND2 (N798, N769, N167);
buf BUF1 (N799, N794);
buf BUF1 (N800, N797);
nand NAND3 (N801, N784, N596, N689);
buf BUF1 (N802, N791);
buf BUF1 (N803, N793);
nor NOR4 (N804, N803, N487, N468, N29);
not NOT1 (N805, N799);
xor XOR2 (N806, N790, N93);
or OR2 (N807, N802, N456);
nand NAND3 (N808, N796, N1, N625);
not NOT1 (N809, N804);
not NOT1 (N810, N800);
nand NAND3 (N811, N809, N135, N436);
or OR4 (N812, N810, N726, N421, N749);
nor NOR4 (N813, N795, N259, N352, N25);
nor NOR2 (N814, N808, N285);
buf BUF1 (N815, N798);
and AND4 (N816, N814, N391, N203, N586);
buf BUF1 (N817, N805);
not NOT1 (N818, N815);
nor NOR4 (N819, N811, N550, N599, N406);
not NOT1 (N820, N817);
xor XOR2 (N821, N819, N289);
buf BUF1 (N822, N818);
nand NAND4 (N823, N822, N732, N502, N795);
buf BUF1 (N824, N821);
buf BUF1 (N825, N816);
nand NAND4 (N826, N806, N434, N162, N708);
or OR2 (N827, N781, N291);
buf BUF1 (N828, N826);
nor NOR2 (N829, N824, N641);
nor NOR4 (N830, N801, N369, N67, N121);
not NOT1 (N831, N813);
not NOT1 (N832, N812);
not NOT1 (N833, N829);
xor XOR2 (N834, N832, N491);
not NOT1 (N835, N823);
or OR2 (N836, N835, N265);
and AND4 (N837, N825, N596, N83, N362);
and AND4 (N838, N837, N338, N583, N196);
nand NAND3 (N839, N838, N227, N243);
xor XOR2 (N840, N839, N443);
or OR2 (N841, N828, N416);
nand NAND2 (N842, N831, N430);
nand NAND2 (N843, N841, N796);
xor XOR2 (N844, N833, N95);
buf BUF1 (N845, N842);
nor NOR3 (N846, N827, N359, N782);
buf BUF1 (N847, N834);
buf BUF1 (N848, N830);
not NOT1 (N849, N845);
nor NOR4 (N850, N840, N530, N522, N827);
nor NOR4 (N851, N850, N806, N770, N371);
nand NAND3 (N852, N836, N707, N685);
and AND4 (N853, N849, N622, N384, N45);
not NOT1 (N854, N853);
not NOT1 (N855, N851);
buf BUF1 (N856, N846);
buf BUF1 (N857, N807);
nand NAND3 (N858, N854, N716, N328);
or OR2 (N859, N843, N179);
or OR3 (N860, N855, N716, N332);
xor XOR2 (N861, N848, N219);
and AND4 (N862, N860, N386, N184, N487);
and AND2 (N863, N861, N742);
not NOT1 (N864, N820);
nand NAND3 (N865, N847, N481, N690);
and AND4 (N866, N864, N670, N778, N2);
nor NOR3 (N867, N865, N849, N334);
nor NOR2 (N868, N857, N296);
not NOT1 (N869, N863);
not NOT1 (N870, N859);
buf BUF1 (N871, N852);
buf BUF1 (N872, N870);
and AND3 (N873, N872, N77, N633);
nor NOR2 (N874, N866, N568);
buf BUF1 (N875, N871);
xor XOR2 (N876, N844, N84);
or OR2 (N877, N874, N195);
not NOT1 (N878, N862);
not NOT1 (N879, N873);
and AND3 (N880, N877, N553, N301);
nand NAND4 (N881, N878, N480, N798, N249);
or OR3 (N882, N869, N871, N527);
nand NAND3 (N883, N876, N530, N11);
and AND3 (N884, N881, N792, N557);
or OR3 (N885, N875, N264, N126);
not NOT1 (N886, N867);
buf BUF1 (N887, N856);
and AND3 (N888, N884, N173, N221);
or OR4 (N889, N882, N197, N501, N152);
xor XOR2 (N890, N885, N885);
or OR3 (N891, N886, N439, N484);
or OR3 (N892, N891, N152, N644);
and AND3 (N893, N888, N30, N765);
and AND4 (N894, N889, N704, N585, N754);
xor XOR2 (N895, N890, N414);
nor NOR2 (N896, N880, N54);
nand NAND4 (N897, N894, N508, N667, N543);
nor NOR4 (N898, N895, N822, N380, N334);
nand NAND3 (N899, N892, N149, N654);
xor XOR2 (N900, N883, N117);
not NOT1 (N901, N899);
nand NAND2 (N902, N893, N870);
nand NAND2 (N903, N897, N552);
and AND3 (N904, N903, N503, N666);
and AND2 (N905, N879, N192);
nand NAND2 (N906, N904, N263);
nor NOR3 (N907, N902, N166, N132);
nand NAND2 (N908, N901, N822);
nor NOR4 (N909, N898, N858, N734, N907);
or OR4 (N910, N381, N245, N850, N772);
nor NOR4 (N911, N780, N895, N401, N633);
not NOT1 (N912, N906);
nand NAND3 (N913, N909, N228, N682);
and AND2 (N914, N913, N756);
buf BUF1 (N915, N912);
or OR4 (N916, N908, N255, N605, N832);
xor XOR2 (N917, N905, N42);
not NOT1 (N918, N911);
or OR2 (N919, N918, N518);
xor XOR2 (N920, N915, N899);
and AND3 (N921, N900, N606, N658);
and AND2 (N922, N868, N902);
nand NAND2 (N923, N922, N633);
xor XOR2 (N924, N923, N633);
nand NAND2 (N925, N919, N478);
or OR3 (N926, N916, N394, N555);
not NOT1 (N927, N921);
nand NAND3 (N928, N927, N391, N96);
or OR2 (N929, N924, N318);
xor XOR2 (N930, N929, N736);
and AND4 (N931, N910, N582, N267, N887);
nand NAND3 (N932, N825, N590, N721);
xor XOR2 (N933, N931, N97);
buf BUF1 (N934, N914);
xor XOR2 (N935, N933, N357);
buf BUF1 (N936, N932);
and AND3 (N937, N925, N308, N224);
or OR4 (N938, N937, N548, N646, N764);
and AND2 (N939, N938, N261);
buf BUF1 (N940, N928);
or OR3 (N941, N940, N754, N894);
or OR4 (N942, N926, N16, N438, N896);
nand NAND3 (N943, N131, N750, N424);
nand NAND4 (N944, N920, N55, N131, N893);
and AND4 (N945, N943, N858, N681, N287);
buf BUF1 (N946, N942);
and AND2 (N947, N936, N57);
or OR2 (N948, N947, N608);
buf BUF1 (N949, N945);
not NOT1 (N950, N946);
nor NOR4 (N951, N948, N560, N521, N63);
not NOT1 (N952, N917);
or OR4 (N953, N934, N60, N789, N367);
not NOT1 (N954, N950);
nand NAND2 (N955, N951, N812);
nor NOR3 (N956, N952, N229, N623);
or OR2 (N957, N956, N281);
not NOT1 (N958, N935);
xor XOR2 (N959, N953, N258);
not NOT1 (N960, N958);
nand NAND3 (N961, N930, N830, N116);
not NOT1 (N962, N955);
buf BUF1 (N963, N960);
not NOT1 (N964, N939);
and AND2 (N965, N961, N776);
not NOT1 (N966, N965);
not NOT1 (N967, N941);
buf BUF1 (N968, N967);
nand NAND2 (N969, N957, N705);
buf BUF1 (N970, N954);
not NOT1 (N971, N962);
or OR4 (N972, N969, N352, N415, N880);
nand NAND3 (N973, N944, N34, N478);
xor XOR2 (N974, N964, N666);
or OR3 (N975, N974, N899, N63);
buf BUF1 (N976, N975);
not NOT1 (N977, N972);
nand NAND2 (N978, N968, N226);
nand NAND4 (N979, N978, N38, N808, N822);
xor XOR2 (N980, N963, N673);
buf BUF1 (N981, N980);
nand NAND2 (N982, N959, N320);
nor NOR2 (N983, N971, N469);
nor NOR4 (N984, N949, N978, N800, N613);
nor NOR4 (N985, N976, N762, N129, N670);
and AND4 (N986, N984, N222, N347, N523);
and AND3 (N987, N986, N20, N623);
or OR4 (N988, N977, N131, N937, N789);
nand NAND4 (N989, N982, N645, N200, N251);
or OR4 (N990, N966, N788, N237, N385);
or OR4 (N991, N983, N772, N956, N132);
xor XOR2 (N992, N979, N783);
or OR2 (N993, N991, N531);
xor XOR2 (N994, N970, N737);
nand NAND4 (N995, N973, N433, N346, N827);
nand NAND2 (N996, N987, N727);
buf BUF1 (N997, N981);
buf BUF1 (N998, N989);
and AND4 (N999, N995, N774, N336, N493);
or OR4 (N1000, N997, N572, N90, N105);
or OR3 (N1001, N994, N280, N394);
nor NOR4 (N1002, N998, N729, N711, N634);
buf BUF1 (N1003, N1000);
or OR2 (N1004, N990, N811);
nand NAND2 (N1005, N985, N829);
and AND4 (N1006, N988, N161, N544, N499);
xor XOR2 (N1007, N1006, N532);
and AND2 (N1008, N993, N526);
xor XOR2 (N1009, N1001, N307);
nand NAND3 (N1010, N1002, N136, N203);
nand NAND3 (N1011, N992, N424, N437);
and AND4 (N1012, N1008, N640, N78, N718);
not NOT1 (N1013, N1003);
xor XOR2 (N1014, N999, N945);
not NOT1 (N1015, N1012);
xor XOR2 (N1016, N1015, N771);
buf BUF1 (N1017, N1005);
not NOT1 (N1018, N1017);
nand NAND3 (N1019, N1004, N787, N556);
nor NOR4 (N1020, N996, N793, N325, N216);
or OR2 (N1021, N1019, N995);
xor XOR2 (N1022, N1016, N150);
xor XOR2 (N1023, N1009, N144);
xor XOR2 (N1024, N1020, N452);
and AND2 (N1025, N1023, N674);
or OR2 (N1026, N1007, N262);
or OR3 (N1027, N1014, N912, N883);
not NOT1 (N1028, N1022);
nand NAND2 (N1029, N1010, N53);
buf BUF1 (N1030, N1018);
not NOT1 (N1031, N1011);
nor NOR2 (N1032, N1030, N212);
xor XOR2 (N1033, N1024, N65);
not NOT1 (N1034, N1032);
not NOT1 (N1035, N1026);
or OR4 (N1036, N1021, N507, N361, N835);
nand NAND3 (N1037, N1036, N501, N321);
and AND3 (N1038, N1025, N1034, N557);
nor NOR4 (N1039, N416, N483, N250, N983);
nor NOR2 (N1040, N1028, N127);
nor NOR3 (N1041, N1038, N870, N551);
nor NOR4 (N1042, N1041, N821, N68, N292);
and AND2 (N1043, N1039, N311);
nand NAND2 (N1044, N1037, N343);
xor XOR2 (N1045, N1031, N930);
xor XOR2 (N1046, N1033, N574);
or OR3 (N1047, N1029, N670, N250);
nor NOR3 (N1048, N1035, N1043, N342);
or OR3 (N1049, N798, N147, N415);
nor NOR4 (N1050, N1013, N155, N724, N934);
and AND2 (N1051, N1027, N883);
not NOT1 (N1052, N1044);
and AND4 (N1053, N1049, N908, N178, N49);
and AND4 (N1054, N1052, N865, N726, N588);
xor XOR2 (N1055, N1048, N490);
buf BUF1 (N1056, N1042);
or OR2 (N1057, N1040, N270);
or OR2 (N1058, N1046, N462);
xor XOR2 (N1059, N1055, N166);
nor NOR4 (N1060, N1054, N480, N40, N692);
xor XOR2 (N1061, N1056, N954);
or OR3 (N1062, N1057, N34, N532);
or OR3 (N1063, N1058, N609, N502);
not NOT1 (N1064, N1063);
and AND4 (N1065, N1060, N711, N45, N95);
nand NAND2 (N1066, N1050, N301);
nand NAND4 (N1067, N1065, N938, N619, N640);
buf BUF1 (N1068, N1062);
not NOT1 (N1069, N1061);
and AND2 (N1070, N1069, N949);
nand NAND2 (N1071, N1047, N434);
or OR2 (N1072, N1071, N942);
not NOT1 (N1073, N1068);
and AND4 (N1074, N1067, N578, N519, N106);
or OR3 (N1075, N1073, N194, N609);
and AND2 (N1076, N1070, N24);
xor XOR2 (N1077, N1072, N944);
and AND2 (N1078, N1077, N923);
and AND3 (N1079, N1066, N745, N824);
not NOT1 (N1080, N1064);
not NOT1 (N1081, N1053);
nor NOR2 (N1082, N1074, N610);
or OR3 (N1083, N1076, N485, N172);
xor XOR2 (N1084, N1051, N566);
buf BUF1 (N1085, N1082);
or OR3 (N1086, N1075, N198, N122);
nor NOR3 (N1087, N1081, N555, N24);
nand NAND4 (N1088, N1080, N231, N769, N878);
nor NOR2 (N1089, N1059, N346);
nand NAND3 (N1090, N1045, N1086, N1039);
xor XOR2 (N1091, N1070, N220);
nand NAND2 (N1092, N1090, N858);
buf BUF1 (N1093, N1085);
and AND2 (N1094, N1092, N179);
nand NAND4 (N1095, N1079, N888, N28, N312);
nand NAND4 (N1096, N1089, N362, N762, N661);
not NOT1 (N1097, N1093);
xor XOR2 (N1098, N1095, N265);
xor XOR2 (N1099, N1078, N185);
buf BUF1 (N1100, N1084);
and AND3 (N1101, N1099, N351, N84);
nor NOR2 (N1102, N1098, N705);
or OR4 (N1103, N1091, N113, N279, N566);
nor NOR3 (N1104, N1102, N631, N529);
or OR3 (N1105, N1097, N424, N825);
not NOT1 (N1106, N1105);
nor NOR4 (N1107, N1087, N555, N304, N742);
not NOT1 (N1108, N1094);
buf BUF1 (N1109, N1101);
nand NAND3 (N1110, N1083, N727, N628);
nor NOR4 (N1111, N1096, N968, N594, N281);
and AND3 (N1112, N1109, N249, N344);
and AND4 (N1113, N1107, N455, N870, N220);
and AND2 (N1114, N1100, N1051);
and AND3 (N1115, N1114, N259, N3);
xor XOR2 (N1116, N1113, N426);
and AND4 (N1117, N1103, N114, N805, N128);
not NOT1 (N1118, N1115);
buf BUF1 (N1119, N1112);
not NOT1 (N1120, N1110);
buf BUF1 (N1121, N1116);
not NOT1 (N1122, N1119);
buf BUF1 (N1123, N1118);
nor NOR2 (N1124, N1108, N245);
not NOT1 (N1125, N1120);
buf BUF1 (N1126, N1121);
or OR3 (N1127, N1117, N802, N200);
or OR2 (N1128, N1111, N394);
nor NOR2 (N1129, N1127, N570);
and AND3 (N1130, N1122, N508, N916);
buf BUF1 (N1131, N1130);
nand NAND2 (N1132, N1124, N830);
or OR4 (N1133, N1104, N16, N567, N62);
xor XOR2 (N1134, N1125, N412);
xor XOR2 (N1135, N1131, N1);
buf BUF1 (N1136, N1123);
buf BUF1 (N1137, N1132);
nand NAND2 (N1138, N1133, N216);
nand NAND4 (N1139, N1128, N1114, N601, N560);
xor XOR2 (N1140, N1139, N576);
and AND2 (N1141, N1140, N207);
and AND2 (N1142, N1135, N713);
not NOT1 (N1143, N1088);
buf BUF1 (N1144, N1141);
or OR2 (N1145, N1126, N588);
xor XOR2 (N1146, N1134, N862);
or OR2 (N1147, N1137, N335);
not NOT1 (N1148, N1147);
nand NAND4 (N1149, N1145, N858, N1077, N688);
nor NOR2 (N1150, N1142, N497);
or OR3 (N1151, N1136, N294, N275);
or OR2 (N1152, N1144, N10);
or OR4 (N1153, N1149, N151, N401, N557);
xor XOR2 (N1154, N1153, N504);
xor XOR2 (N1155, N1129, N1142);
xor XOR2 (N1156, N1146, N407);
not NOT1 (N1157, N1106);
buf BUF1 (N1158, N1151);
or OR2 (N1159, N1152, N442);
xor XOR2 (N1160, N1155, N264);
buf BUF1 (N1161, N1157);
nor NOR4 (N1162, N1154, N455, N811, N721);
nor NOR4 (N1163, N1162, N830, N799, N328);
xor XOR2 (N1164, N1156, N514);
buf BUF1 (N1165, N1150);
and AND4 (N1166, N1163, N381, N196, N1078);
and AND4 (N1167, N1166, N410, N64, N342);
not NOT1 (N1168, N1159);
nand NAND3 (N1169, N1158, N848, N955);
and AND2 (N1170, N1164, N1034);
xor XOR2 (N1171, N1143, N826);
not NOT1 (N1172, N1169);
or OR3 (N1173, N1168, N835, N699);
xor XOR2 (N1174, N1167, N1100);
or OR4 (N1175, N1171, N965, N861, N423);
not NOT1 (N1176, N1148);
nor NOR2 (N1177, N1160, N438);
nor NOR3 (N1178, N1138, N588, N850);
buf BUF1 (N1179, N1161);
nor NOR3 (N1180, N1174, N395, N573);
buf BUF1 (N1181, N1179);
xor XOR2 (N1182, N1170, N285);
and AND3 (N1183, N1177, N626, N50);
nand NAND3 (N1184, N1173, N611, N835);
buf BUF1 (N1185, N1180);
or OR3 (N1186, N1165, N1167, N445);
nand NAND2 (N1187, N1181, N645);
nor NOR4 (N1188, N1185, N806, N468, N323);
not NOT1 (N1189, N1176);
nor NOR3 (N1190, N1184, N269, N1139);
xor XOR2 (N1191, N1178, N1154);
buf BUF1 (N1192, N1182);
not NOT1 (N1193, N1190);
and AND4 (N1194, N1193, N598, N781, N684);
nor NOR4 (N1195, N1187, N195, N1177, N325);
nor NOR4 (N1196, N1183, N1041, N412, N436);
nor NOR2 (N1197, N1191, N919);
nand NAND2 (N1198, N1188, N584);
or OR3 (N1199, N1194, N289, N136);
nand NAND4 (N1200, N1186, N725, N521, N823);
nand NAND4 (N1201, N1200, N693, N95, N660);
nor NOR4 (N1202, N1172, N316, N165, N131);
nor NOR3 (N1203, N1202, N1190, N1101);
and AND3 (N1204, N1203, N327, N482);
nand NAND4 (N1205, N1192, N1149, N77, N88);
or OR3 (N1206, N1201, N804, N522);
or OR3 (N1207, N1196, N796, N287);
buf BUF1 (N1208, N1189);
and AND3 (N1209, N1195, N382, N1032);
nor NOR3 (N1210, N1197, N490, N232);
not NOT1 (N1211, N1207);
not NOT1 (N1212, N1210);
and AND3 (N1213, N1209, N22, N441);
or OR3 (N1214, N1204, N734, N72);
or OR2 (N1215, N1205, N954);
nor NOR3 (N1216, N1199, N617, N505);
not NOT1 (N1217, N1216);
and AND3 (N1218, N1217, N1212, N844);
xor XOR2 (N1219, N1038, N766);
nor NOR4 (N1220, N1208, N357, N654, N246);
and AND2 (N1221, N1211, N638);
nand NAND2 (N1222, N1206, N781);
or OR4 (N1223, N1198, N340, N671, N919);
buf BUF1 (N1224, N1218);
and AND2 (N1225, N1175, N1224);
and AND3 (N1226, N601, N556, N326);
or OR4 (N1227, N1220, N716, N75, N785);
nand NAND3 (N1228, N1225, N494, N106);
nand NAND3 (N1229, N1221, N1136, N1041);
nand NAND2 (N1230, N1228, N217);
nor NOR2 (N1231, N1227, N912);
nand NAND3 (N1232, N1222, N572, N202);
xor XOR2 (N1233, N1232, N441);
nand NAND3 (N1234, N1226, N170, N406);
or OR2 (N1235, N1234, N410);
xor XOR2 (N1236, N1213, N1118);
and AND4 (N1237, N1215, N630, N1199, N989);
and AND3 (N1238, N1214, N865, N196);
buf BUF1 (N1239, N1235);
nor NOR4 (N1240, N1230, N615, N643, N917);
nor NOR4 (N1241, N1238, N69, N84, N1182);
nor NOR3 (N1242, N1231, N710, N919);
nand NAND4 (N1243, N1219, N918, N293, N522);
and AND3 (N1244, N1241, N71, N3);
and AND3 (N1245, N1243, N15, N1227);
nand NAND2 (N1246, N1245, N1139);
and AND2 (N1247, N1246, N583);
nand NAND4 (N1248, N1242, N663, N515, N1222);
nor NOR2 (N1249, N1236, N1136);
not NOT1 (N1250, N1248);
and AND3 (N1251, N1239, N949, N687);
nand NAND3 (N1252, N1233, N941, N989);
buf BUF1 (N1253, N1250);
nand NAND3 (N1254, N1244, N1050, N692);
nor NOR2 (N1255, N1249, N838);
nor NOR3 (N1256, N1247, N1158, N1158);
nand NAND4 (N1257, N1256, N1223, N209, N408);
nor NOR2 (N1258, N1123, N1026);
nand NAND3 (N1259, N1251, N103, N388);
xor XOR2 (N1260, N1259, N868);
nor NOR3 (N1261, N1229, N754, N1011);
or OR3 (N1262, N1261, N458, N53);
or OR2 (N1263, N1260, N528);
not NOT1 (N1264, N1237);
and AND2 (N1265, N1255, N900);
xor XOR2 (N1266, N1258, N1158);
and AND4 (N1267, N1266, N990, N640, N1223);
xor XOR2 (N1268, N1252, N1123);
xor XOR2 (N1269, N1263, N756);
buf BUF1 (N1270, N1253);
and AND2 (N1271, N1262, N791);
and AND4 (N1272, N1268, N536, N894, N862);
or OR3 (N1273, N1271, N383, N1147);
nand NAND4 (N1274, N1264, N895, N725, N286);
nor NOR4 (N1275, N1240, N568, N1022, N341);
and AND2 (N1276, N1267, N289);
xor XOR2 (N1277, N1265, N988);
not NOT1 (N1278, N1277);
buf BUF1 (N1279, N1257);
buf BUF1 (N1280, N1276);
nor NOR4 (N1281, N1275, N1055, N277, N939);
not NOT1 (N1282, N1281);
or OR3 (N1283, N1270, N388, N630);
or OR2 (N1284, N1282, N914);
or OR4 (N1285, N1269, N241, N902, N182);
xor XOR2 (N1286, N1278, N792);
or OR4 (N1287, N1284, N1199, N1119, N701);
nand NAND2 (N1288, N1285, N677);
and AND2 (N1289, N1287, N324);
nor NOR4 (N1290, N1288, N264, N341, N459);
nor NOR2 (N1291, N1273, N136);
buf BUF1 (N1292, N1280);
xor XOR2 (N1293, N1292, N794);
xor XOR2 (N1294, N1291, N596);
nand NAND4 (N1295, N1286, N977, N625, N167);
nand NAND3 (N1296, N1283, N461, N1279);
not NOT1 (N1297, N1229);
not NOT1 (N1298, N1296);
xor XOR2 (N1299, N1272, N1142);
not NOT1 (N1300, N1274);
and AND2 (N1301, N1297, N1039);
or OR3 (N1302, N1293, N525, N878);
buf BUF1 (N1303, N1254);
or OR4 (N1304, N1301, N1167, N585, N596);
or OR2 (N1305, N1303, N473);
buf BUF1 (N1306, N1298);
and AND2 (N1307, N1295, N1249);
and AND4 (N1308, N1294, N1295, N1049, N499);
nand NAND2 (N1309, N1304, N439);
xor XOR2 (N1310, N1290, N776);
or OR4 (N1311, N1302, N719, N818, N49);
buf BUF1 (N1312, N1309);
nand NAND3 (N1313, N1299, N1070, N23);
nand NAND4 (N1314, N1289, N474, N981, N520);
nand NAND2 (N1315, N1312, N967);
nand NAND4 (N1316, N1307, N167, N1144, N1216);
nor NOR2 (N1317, N1314, N1200);
not NOT1 (N1318, N1311);
not NOT1 (N1319, N1305);
or OR4 (N1320, N1313, N591, N120, N203);
buf BUF1 (N1321, N1319);
xor XOR2 (N1322, N1321, N838);
nand NAND2 (N1323, N1318, N305);
buf BUF1 (N1324, N1308);
nand NAND3 (N1325, N1324, N1220, N782);
nand NAND2 (N1326, N1322, N643);
buf BUF1 (N1327, N1316);
nor NOR4 (N1328, N1323, N723, N1211, N1183);
not NOT1 (N1329, N1326);
not NOT1 (N1330, N1317);
not NOT1 (N1331, N1329);
and AND2 (N1332, N1325, N681);
nand NAND3 (N1333, N1328, N498, N1268);
nand NAND3 (N1334, N1306, N811, N940);
nor NOR2 (N1335, N1320, N1318);
buf BUF1 (N1336, N1327);
or OR4 (N1337, N1315, N816, N397, N1150);
nand NAND2 (N1338, N1335, N793);
xor XOR2 (N1339, N1300, N658);
nand NAND2 (N1340, N1334, N725);
buf BUF1 (N1341, N1336);
nand NAND2 (N1342, N1330, N613);
xor XOR2 (N1343, N1341, N870);
buf BUF1 (N1344, N1338);
nand NAND3 (N1345, N1342, N468, N77);
xor XOR2 (N1346, N1337, N201);
or OR4 (N1347, N1331, N376, N734, N1251);
nor NOR4 (N1348, N1347, N658, N331, N874);
and AND2 (N1349, N1333, N1140);
buf BUF1 (N1350, N1349);
not NOT1 (N1351, N1340);
nand NAND3 (N1352, N1339, N29, N664);
xor XOR2 (N1353, N1345, N488);
not NOT1 (N1354, N1352);
nor NOR4 (N1355, N1351, N1175, N63, N1079);
nand NAND3 (N1356, N1343, N863, N1221);
xor XOR2 (N1357, N1348, N438);
and AND4 (N1358, N1344, N869, N145, N1304);
nor NOR3 (N1359, N1357, N789, N710);
xor XOR2 (N1360, N1355, N908);
nor NOR3 (N1361, N1332, N1190, N1340);
nor NOR4 (N1362, N1350, N286, N672, N517);
nand NAND4 (N1363, N1362, N144, N60, N1132);
nor NOR2 (N1364, N1363, N840);
buf BUF1 (N1365, N1353);
nand NAND2 (N1366, N1365, N100);
not NOT1 (N1367, N1358);
not NOT1 (N1368, N1364);
nor NOR4 (N1369, N1366, N195, N308, N978);
xor XOR2 (N1370, N1361, N1071);
not NOT1 (N1371, N1369);
not NOT1 (N1372, N1368);
buf BUF1 (N1373, N1354);
or OR2 (N1374, N1371, N1274);
and AND3 (N1375, N1367, N937, N1043);
buf BUF1 (N1376, N1359);
and AND3 (N1377, N1372, N389, N736);
buf BUF1 (N1378, N1376);
buf BUF1 (N1379, N1373);
xor XOR2 (N1380, N1374, N788);
nor NOR3 (N1381, N1378, N1245, N1193);
xor XOR2 (N1382, N1356, N706);
and AND2 (N1383, N1377, N560);
buf BUF1 (N1384, N1380);
nand NAND2 (N1385, N1381, N1352);
or OR2 (N1386, N1346, N440);
nor NOR2 (N1387, N1375, N244);
and AND2 (N1388, N1310, N23);
nor NOR2 (N1389, N1370, N1381);
or OR4 (N1390, N1382, N440, N521, N356);
nand NAND3 (N1391, N1379, N380, N284);
not NOT1 (N1392, N1360);
or OR4 (N1393, N1387, N694, N940, N199);
nand NAND4 (N1394, N1385, N659, N517, N515);
nor NOR4 (N1395, N1391, N741, N134, N1058);
not NOT1 (N1396, N1389);
nand NAND2 (N1397, N1394, N1319);
nor NOR3 (N1398, N1392, N1189, N420);
nor NOR2 (N1399, N1397, N494);
not NOT1 (N1400, N1390);
xor XOR2 (N1401, N1386, N588);
nand NAND2 (N1402, N1396, N761);
or OR3 (N1403, N1384, N447, N120);
xor XOR2 (N1404, N1395, N118);
nor NOR2 (N1405, N1383, N667);
and AND3 (N1406, N1398, N66, N146);
xor XOR2 (N1407, N1406, N761);
xor XOR2 (N1408, N1399, N1014);
and AND4 (N1409, N1401, N232, N1100, N292);
buf BUF1 (N1410, N1408);
xor XOR2 (N1411, N1405, N1343);
xor XOR2 (N1412, N1411, N679);
nor NOR3 (N1413, N1410, N293, N1408);
not NOT1 (N1414, N1409);
xor XOR2 (N1415, N1413, N289);
nand NAND2 (N1416, N1402, N151);
xor XOR2 (N1417, N1404, N1247);
nor NOR3 (N1418, N1403, N72, N1301);
buf BUF1 (N1419, N1416);
buf BUF1 (N1420, N1419);
not NOT1 (N1421, N1412);
buf BUF1 (N1422, N1415);
and AND3 (N1423, N1422, N801, N836);
nand NAND4 (N1424, N1400, N1053, N140, N399);
xor XOR2 (N1425, N1418, N787);
or OR3 (N1426, N1421, N762, N893);
nand NAND4 (N1427, N1424, N38, N1203, N421);
nand NAND3 (N1428, N1414, N1055, N24);
and AND4 (N1429, N1427, N275, N856, N276);
nor NOR2 (N1430, N1417, N27);
not NOT1 (N1431, N1430);
or OR3 (N1432, N1388, N568, N38);
xor XOR2 (N1433, N1393, N156);
nor NOR4 (N1434, N1426, N42, N446, N1355);
and AND3 (N1435, N1432, N1419, N1141);
not NOT1 (N1436, N1428);
xor XOR2 (N1437, N1429, N826);
nand NAND2 (N1438, N1423, N139);
nor NOR2 (N1439, N1433, N1297);
buf BUF1 (N1440, N1425);
not NOT1 (N1441, N1436);
or OR2 (N1442, N1431, N212);
or OR4 (N1443, N1434, N547, N828, N728);
buf BUF1 (N1444, N1441);
or OR2 (N1445, N1443, N449);
xor XOR2 (N1446, N1442, N1128);
xor XOR2 (N1447, N1437, N160);
nand NAND2 (N1448, N1447, N1113);
nand NAND2 (N1449, N1439, N395);
and AND2 (N1450, N1435, N503);
buf BUF1 (N1451, N1446);
not NOT1 (N1452, N1407);
nand NAND3 (N1453, N1448, N830, N328);
or OR2 (N1454, N1451, N663);
or OR4 (N1455, N1454, N297, N236, N1287);
nand NAND3 (N1456, N1438, N687, N823);
and AND4 (N1457, N1453, N1300, N556, N508);
xor XOR2 (N1458, N1452, N886);
or OR2 (N1459, N1440, N1207);
and AND2 (N1460, N1450, N1315);
nor NOR2 (N1461, N1458, N838);
not NOT1 (N1462, N1457);
nand NAND4 (N1463, N1420, N1290, N1436, N197);
nand NAND4 (N1464, N1460, N23, N916, N332);
nor NOR3 (N1465, N1463, N1338, N60);
not NOT1 (N1466, N1459);
nand NAND4 (N1467, N1462, N1170, N466, N573);
or OR2 (N1468, N1464, N826);
nand NAND2 (N1469, N1465, N800);
and AND4 (N1470, N1455, N1405, N1452, N119);
and AND4 (N1471, N1470, N466, N755, N866);
and AND3 (N1472, N1471, N705, N1421);
and AND3 (N1473, N1467, N394, N702);
xor XOR2 (N1474, N1456, N373);
not NOT1 (N1475, N1445);
xor XOR2 (N1476, N1468, N264);
xor XOR2 (N1477, N1472, N1324);
or OR3 (N1478, N1466, N1273, N859);
nor NOR4 (N1479, N1478, N1295, N710, N1315);
buf BUF1 (N1480, N1477);
nand NAND2 (N1481, N1473, N838);
buf BUF1 (N1482, N1476);
not NOT1 (N1483, N1461);
nand NAND4 (N1484, N1481, N540, N971, N634);
nand NAND2 (N1485, N1469, N968);
nand NAND3 (N1486, N1482, N586, N1233);
buf BUF1 (N1487, N1479);
and AND2 (N1488, N1475, N210);
or OR3 (N1489, N1486, N1088, N399);
and AND3 (N1490, N1449, N1047, N211);
not NOT1 (N1491, N1483);
or OR2 (N1492, N1487, N74);
nor NOR3 (N1493, N1484, N1124, N1327);
xor XOR2 (N1494, N1474, N978);
buf BUF1 (N1495, N1490);
xor XOR2 (N1496, N1488, N1091);
and AND4 (N1497, N1491, N1295, N268, N536);
not NOT1 (N1498, N1493);
xor XOR2 (N1499, N1497, N1083);
nand NAND2 (N1500, N1489, N589);
nor NOR4 (N1501, N1444, N837, N9, N682);
or OR3 (N1502, N1485, N627, N878);
nand NAND3 (N1503, N1496, N413, N1307);
nand NAND2 (N1504, N1494, N830);
nand NAND4 (N1505, N1501, N182, N353, N1137);
or OR2 (N1506, N1492, N401);
nand NAND2 (N1507, N1500, N1468);
xor XOR2 (N1508, N1495, N147);
nor NOR4 (N1509, N1508, N604, N875, N1237);
or OR3 (N1510, N1499, N389, N814);
not NOT1 (N1511, N1502);
nand NAND2 (N1512, N1504, N941);
xor XOR2 (N1513, N1505, N1348);
nor NOR3 (N1514, N1503, N861, N1388);
nand NAND2 (N1515, N1514, N410);
nor NOR3 (N1516, N1506, N859, N141);
buf BUF1 (N1517, N1512);
or OR3 (N1518, N1509, N856, N1142);
xor XOR2 (N1519, N1518, N1090);
nand NAND4 (N1520, N1519, N805, N1288, N1272);
or OR2 (N1521, N1515, N177);
nor NOR2 (N1522, N1480, N219);
and AND2 (N1523, N1522, N1434);
nand NAND3 (N1524, N1507, N1511, N1225);
nand NAND3 (N1525, N767, N868, N1190);
nor NOR3 (N1526, N1525, N215, N929);
nand NAND4 (N1527, N1523, N1100, N457, N1101);
and AND3 (N1528, N1524, N39, N263);
not NOT1 (N1529, N1521);
xor XOR2 (N1530, N1498, N1490);
or OR4 (N1531, N1513, N876, N1087, N1278);
and AND4 (N1532, N1530, N712, N386, N523);
xor XOR2 (N1533, N1510, N114);
or OR3 (N1534, N1531, N1226, N1402);
xor XOR2 (N1535, N1534, N125);
nand NAND2 (N1536, N1516, N97);
and AND4 (N1537, N1533, N360, N534, N985);
or OR2 (N1538, N1535, N285);
xor XOR2 (N1539, N1520, N959);
buf BUF1 (N1540, N1532);
not NOT1 (N1541, N1528);
or OR3 (N1542, N1537, N854, N854);
not NOT1 (N1543, N1526);
or OR4 (N1544, N1527, N982, N147, N851);
buf BUF1 (N1545, N1543);
xor XOR2 (N1546, N1544, N1518);
not NOT1 (N1547, N1517);
not NOT1 (N1548, N1539);
buf BUF1 (N1549, N1542);
xor XOR2 (N1550, N1549, N426);
buf BUF1 (N1551, N1550);
buf BUF1 (N1552, N1540);
not NOT1 (N1553, N1547);
or OR4 (N1554, N1551, N558, N48, N463);
buf BUF1 (N1555, N1536);
or OR3 (N1556, N1552, N596, N1395);
buf BUF1 (N1557, N1554);
and AND2 (N1558, N1556, N1112);
nand NAND2 (N1559, N1555, N126);
and AND4 (N1560, N1557, N1512, N856, N263);
xor XOR2 (N1561, N1548, N284);
xor XOR2 (N1562, N1553, N637);
not NOT1 (N1563, N1545);
or OR4 (N1564, N1558, N448, N1176, N1293);
not NOT1 (N1565, N1546);
nand NAND2 (N1566, N1564, N677);
xor XOR2 (N1567, N1560, N1001);
buf BUF1 (N1568, N1541);
nor NOR4 (N1569, N1561, N1264, N485, N1551);
and AND4 (N1570, N1538, N1450, N1386, N469);
nand NAND3 (N1571, N1562, N185, N923);
nor NOR4 (N1572, N1567, N1116, N782, N1567);
buf BUF1 (N1573, N1563);
nand NAND3 (N1574, N1569, N380, N514);
nor NOR4 (N1575, N1573, N17, N1499, N1014);
or OR2 (N1576, N1529, N976);
xor XOR2 (N1577, N1570, N742);
xor XOR2 (N1578, N1559, N1092);
or OR2 (N1579, N1566, N979);
nor NOR4 (N1580, N1565, N779, N1186, N174);
buf BUF1 (N1581, N1578);
xor XOR2 (N1582, N1574, N554);
buf BUF1 (N1583, N1581);
xor XOR2 (N1584, N1575, N1064);
buf BUF1 (N1585, N1571);
not NOT1 (N1586, N1580);
xor XOR2 (N1587, N1577, N794);
and AND4 (N1588, N1585, N1545, N1424, N577);
xor XOR2 (N1589, N1584, N372);
nor NOR3 (N1590, N1568, N928, N197);
or OR2 (N1591, N1583, N221);
nor NOR2 (N1592, N1591, N1245);
nand NAND2 (N1593, N1592, N1264);
nand NAND4 (N1594, N1576, N805, N551, N279);
xor XOR2 (N1595, N1594, N446);
or OR3 (N1596, N1572, N301, N466);
xor XOR2 (N1597, N1587, N445);
nand NAND3 (N1598, N1595, N978, N1413);
or OR3 (N1599, N1597, N662, N1370);
not NOT1 (N1600, N1588);
not NOT1 (N1601, N1598);
or OR3 (N1602, N1590, N921, N437);
and AND3 (N1603, N1602, N1401, N1242);
and AND3 (N1604, N1586, N121, N336);
xor XOR2 (N1605, N1589, N1560);
not NOT1 (N1606, N1582);
buf BUF1 (N1607, N1605);
nand NAND4 (N1608, N1593, N1571, N389, N520);
and AND3 (N1609, N1601, N583, N1537);
nand NAND4 (N1610, N1596, N862, N1321, N531);
not NOT1 (N1611, N1604);
buf BUF1 (N1612, N1600);
and AND3 (N1613, N1603, N1565, N954);
nor NOR2 (N1614, N1609, N748);
buf BUF1 (N1615, N1579);
or OR4 (N1616, N1608, N480, N138, N1458);
nand NAND3 (N1617, N1606, N1413, N573);
nand NAND3 (N1618, N1616, N1141, N469);
nor NOR2 (N1619, N1617, N75);
buf BUF1 (N1620, N1611);
or OR2 (N1621, N1618, N545);
buf BUF1 (N1622, N1614);
nor NOR4 (N1623, N1610, N672, N176, N29);
and AND2 (N1624, N1621, N592);
and AND4 (N1625, N1615, N1143, N918, N1144);
and AND2 (N1626, N1607, N113);
nor NOR4 (N1627, N1612, N1228, N17, N1555);
nand NAND4 (N1628, N1613, N835, N159, N708);
or OR4 (N1629, N1623, N1299, N349, N864);
xor XOR2 (N1630, N1599, N1543);
xor XOR2 (N1631, N1620, N211);
nor NOR4 (N1632, N1624, N248, N387, N280);
and AND3 (N1633, N1632, N568, N1488);
and AND2 (N1634, N1622, N426);
buf BUF1 (N1635, N1619);
or OR4 (N1636, N1627, N541, N330, N905);
not NOT1 (N1637, N1633);
buf BUF1 (N1638, N1635);
nor NOR2 (N1639, N1634, N905);
nor NOR3 (N1640, N1639, N332, N1531);
or OR4 (N1641, N1636, N324, N478, N73);
nor NOR2 (N1642, N1640, N1026);
xor XOR2 (N1643, N1630, N1530);
or OR2 (N1644, N1631, N36);
nand NAND4 (N1645, N1641, N1605, N1384, N158);
and AND4 (N1646, N1638, N1170, N567, N1070);
and AND3 (N1647, N1642, N546, N954);
not NOT1 (N1648, N1645);
buf BUF1 (N1649, N1637);
xor XOR2 (N1650, N1648, N997);
xor XOR2 (N1651, N1625, N1487);
or OR3 (N1652, N1628, N1421, N1150);
and AND4 (N1653, N1644, N700, N578, N697);
nand NAND4 (N1654, N1651, N642, N961, N160);
nor NOR3 (N1655, N1650, N745, N324);
xor XOR2 (N1656, N1629, N1591);
nand NAND2 (N1657, N1652, N1415);
and AND2 (N1658, N1654, N1629);
nand NAND4 (N1659, N1653, N873, N624, N371);
and AND2 (N1660, N1626, N486);
xor XOR2 (N1661, N1656, N1226);
xor XOR2 (N1662, N1655, N286);
not NOT1 (N1663, N1661);
not NOT1 (N1664, N1649);
xor XOR2 (N1665, N1660, N1037);
nor NOR2 (N1666, N1659, N1186);
buf BUF1 (N1667, N1666);
not NOT1 (N1668, N1665);
xor XOR2 (N1669, N1647, N663);
not NOT1 (N1670, N1658);
xor XOR2 (N1671, N1664, N721);
and AND4 (N1672, N1662, N1108, N1556, N1635);
xor XOR2 (N1673, N1657, N46);
nor NOR4 (N1674, N1670, N819, N550, N929);
xor XOR2 (N1675, N1667, N1420);
or OR2 (N1676, N1675, N1347);
buf BUF1 (N1677, N1673);
nor NOR2 (N1678, N1674, N815);
xor XOR2 (N1679, N1671, N1541);
buf BUF1 (N1680, N1677);
and AND4 (N1681, N1643, N724, N166, N108);
nand NAND4 (N1682, N1669, N539, N47, N1062);
nor NOR2 (N1683, N1672, N846);
buf BUF1 (N1684, N1668);
and AND3 (N1685, N1678, N6, N529);
xor XOR2 (N1686, N1646, N1126);
xor XOR2 (N1687, N1676, N549);
nand NAND2 (N1688, N1687, N234);
and AND4 (N1689, N1684, N532, N86, N1529);
nand NAND3 (N1690, N1686, N1081, N1402);
nor NOR4 (N1691, N1689, N1071, N616, N884);
nor NOR4 (N1692, N1681, N1486, N846, N917);
not NOT1 (N1693, N1691);
or OR2 (N1694, N1685, N344);
xor XOR2 (N1695, N1663, N699);
and AND4 (N1696, N1690, N1425, N577, N464);
or OR3 (N1697, N1683, N1149, N552);
or OR4 (N1698, N1694, N963, N1589, N1508);
and AND3 (N1699, N1695, N1487, N788);
nand NAND3 (N1700, N1696, N1109, N1366);
not NOT1 (N1701, N1682);
not NOT1 (N1702, N1679);
nor NOR2 (N1703, N1699, N334);
and AND3 (N1704, N1701, N789, N1207);
not NOT1 (N1705, N1692);
or OR2 (N1706, N1698, N43);
not NOT1 (N1707, N1703);
nand NAND2 (N1708, N1704, N236);
nor NOR4 (N1709, N1708, N1158, N519, N28);
xor XOR2 (N1710, N1700, N1604);
nor NOR2 (N1711, N1706, N1495);
nand NAND2 (N1712, N1711, N281);
nand NAND4 (N1713, N1697, N1705, N1228, N336);
and AND4 (N1714, N1158, N1213, N1704, N1193);
xor XOR2 (N1715, N1710, N1673);
nor NOR2 (N1716, N1702, N239);
nor NOR2 (N1717, N1713, N502);
and AND2 (N1718, N1680, N1268);
not NOT1 (N1719, N1718);
nor NOR4 (N1720, N1714, N1478, N1165, N1058);
or OR4 (N1721, N1715, N576, N988, N946);
nor NOR3 (N1722, N1693, N357, N1038);
not NOT1 (N1723, N1716);
nor NOR2 (N1724, N1722, N282);
nand NAND2 (N1725, N1707, N555);
xor XOR2 (N1726, N1723, N280);
and AND3 (N1727, N1726, N1036, N1527);
buf BUF1 (N1728, N1727);
or OR4 (N1729, N1720, N920, N1242, N1430);
not NOT1 (N1730, N1709);
xor XOR2 (N1731, N1719, N276);
nor NOR2 (N1732, N1729, N542);
and AND4 (N1733, N1731, N1700, N1186, N1679);
xor XOR2 (N1734, N1721, N1227);
and AND3 (N1735, N1730, N875, N1455);
or OR3 (N1736, N1725, N533, N573);
not NOT1 (N1737, N1728);
and AND4 (N1738, N1737, N209, N384, N294);
nor NOR4 (N1739, N1717, N975, N235, N268);
and AND3 (N1740, N1732, N806, N638);
xor XOR2 (N1741, N1738, N1546);
or OR4 (N1742, N1724, N975, N1706, N530);
and AND2 (N1743, N1733, N252);
nand NAND4 (N1744, N1743, N376, N28, N989);
and AND3 (N1745, N1744, N11, N1472);
nor NOR2 (N1746, N1688, N820);
or OR3 (N1747, N1742, N864, N1433);
nand NAND2 (N1748, N1745, N1495);
nand NAND3 (N1749, N1747, N773, N1043);
nor NOR4 (N1750, N1741, N1570, N624, N944);
xor XOR2 (N1751, N1740, N322);
and AND4 (N1752, N1735, N1368, N846, N1170);
xor XOR2 (N1753, N1748, N876);
or OR4 (N1754, N1749, N563, N1701, N1558);
nor NOR4 (N1755, N1752, N1394, N182, N800);
not NOT1 (N1756, N1739);
and AND4 (N1757, N1712, N1741, N1230, N187);
nand NAND3 (N1758, N1734, N1726, N602);
nor NOR2 (N1759, N1750, N1539);
or OR2 (N1760, N1758, N132);
nand NAND4 (N1761, N1755, N722, N243, N204);
or OR4 (N1762, N1753, N1495, N489, N878);
nor NOR4 (N1763, N1760, N475, N1699, N1123);
buf BUF1 (N1764, N1762);
not NOT1 (N1765, N1761);
not NOT1 (N1766, N1764);
buf BUF1 (N1767, N1736);
xor XOR2 (N1768, N1765, N129);
nand NAND2 (N1769, N1751, N1176);
nand NAND2 (N1770, N1759, N782);
or OR2 (N1771, N1754, N175);
and AND4 (N1772, N1757, N1459, N208, N1521);
buf BUF1 (N1773, N1771);
nand NAND2 (N1774, N1767, N1581);
or OR2 (N1775, N1769, N1547);
and AND3 (N1776, N1763, N1552, N64);
not NOT1 (N1777, N1770);
xor XOR2 (N1778, N1776, N1423);
not NOT1 (N1779, N1775);
and AND4 (N1780, N1772, N85, N308, N1517);
buf BUF1 (N1781, N1778);
and AND2 (N1782, N1780, N308);
and AND2 (N1783, N1746, N1132);
nand NAND2 (N1784, N1779, N712);
nand NAND2 (N1785, N1784, N582);
not NOT1 (N1786, N1768);
or OR4 (N1787, N1783, N1118, N722, N1387);
buf BUF1 (N1788, N1766);
buf BUF1 (N1789, N1756);
nand NAND4 (N1790, N1787, N861, N401, N1277);
buf BUF1 (N1791, N1777);
or OR2 (N1792, N1791, N51);
or OR3 (N1793, N1782, N1628, N203);
not NOT1 (N1794, N1781);
nor NOR4 (N1795, N1788, N1290, N320, N1455);
nand NAND4 (N1796, N1793, N1721, N873, N1788);
buf BUF1 (N1797, N1790);
nor NOR3 (N1798, N1794, N463, N1611);
xor XOR2 (N1799, N1789, N45);
nor NOR4 (N1800, N1798, N364, N472, N1598);
xor XOR2 (N1801, N1795, N961);
buf BUF1 (N1802, N1801);
and AND3 (N1803, N1796, N1802, N738);
and AND3 (N1804, N1267, N344, N186);
buf BUF1 (N1805, N1785);
and AND2 (N1806, N1786, N1484);
or OR3 (N1807, N1792, N1790, N162);
not NOT1 (N1808, N1807);
and AND2 (N1809, N1804, N1579);
nand NAND4 (N1810, N1799, N233, N212, N698);
or OR2 (N1811, N1810, N161);
not NOT1 (N1812, N1797);
nand NAND4 (N1813, N1805, N939, N581, N493);
nor NOR2 (N1814, N1803, N1484);
xor XOR2 (N1815, N1774, N733);
nor NOR2 (N1816, N1813, N282);
or OR4 (N1817, N1814, N612, N1245, N707);
buf BUF1 (N1818, N1773);
not NOT1 (N1819, N1812);
not NOT1 (N1820, N1819);
nor NOR3 (N1821, N1818, N1664, N254);
or OR2 (N1822, N1821, N911);
nor NOR3 (N1823, N1808, N1417, N105);
or OR2 (N1824, N1806, N1687);
xor XOR2 (N1825, N1800, N1032);
or OR4 (N1826, N1824, N1553, N329, N1121);
nor NOR2 (N1827, N1820, N1236);
nor NOR4 (N1828, N1809, N868, N1583, N1672);
nand NAND4 (N1829, N1823, N1770, N1075, N1206);
buf BUF1 (N1830, N1811);
nand NAND2 (N1831, N1822, N139);
and AND3 (N1832, N1827, N1062, N546);
xor XOR2 (N1833, N1815, N838);
buf BUF1 (N1834, N1833);
nand NAND2 (N1835, N1825, N954);
not NOT1 (N1836, N1817);
not NOT1 (N1837, N1832);
and AND4 (N1838, N1831, N238, N530, N1088);
nand NAND4 (N1839, N1837, N1632, N124, N528);
nand NAND4 (N1840, N1828, N534, N1340, N1515);
nor NOR4 (N1841, N1816, N144, N310, N846);
xor XOR2 (N1842, N1834, N678);
or OR3 (N1843, N1842, N182, N266);
and AND2 (N1844, N1826, N1716);
nand NAND4 (N1845, N1844, N922, N208, N906);
nand NAND2 (N1846, N1839, N1239);
xor XOR2 (N1847, N1838, N972);
nor NOR2 (N1848, N1836, N1779);
nand NAND4 (N1849, N1845, N458, N606, N177);
nor NOR3 (N1850, N1840, N437, N179);
nand NAND2 (N1851, N1843, N1256);
xor XOR2 (N1852, N1849, N1826);
xor XOR2 (N1853, N1848, N1680);
or OR3 (N1854, N1850, N1633, N765);
nor NOR4 (N1855, N1851, N1090, N947, N850);
not NOT1 (N1856, N1841);
and AND3 (N1857, N1853, N1212, N487);
and AND4 (N1858, N1855, N1289, N959, N1505);
nand NAND4 (N1859, N1854, N440, N205, N1782);
buf BUF1 (N1860, N1830);
not NOT1 (N1861, N1857);
or OR4 (N1862, N1847, N867, N997, N1737);
xor XOR2 (N1863, N1862, N502);
nor NOR2 (N1864, N1829, N1733);
nand NAND3 (N1865, N1835, N1774, N1440);
nor NOR3 (N1866, N1861, N1437, N356);
nand NAND3 (N1867, N1859, N1210, N824);
not NOT1 (N1868, N1867);
and AND2 (N1869, N1852, N580);
or OR4 (N1870, N1858, N1820, N1173, N334);
or OR4 (N1871, N1870, N274, N1092, N411);
or OR3 (N1872, N1864, N216, N460);
buf BUF1 (N1873, N1846);
xor XOR2 (N1874, N1866, N142);
nor NOR3 (N1875, N1865, N1044, N838);
xor XOR2 (N1876, N1872, N812);
xor XOR2 (N1877, N1871, N134);
not NOT1 (N1878, N1876);
not NOT1 (N1879, N1863);
or OR3 (N1880, N1877, N737, N743);
not NOT1 (N1881, N1868);
and AND2 (N1882, N1879, N152);
nor NOR2 (N1883, N1880, N54);
xor XOR2 (N1884, N1874, N650);
nor NOR3 (N1885, N1882, N158, N1696);
xor XOR2 (N1886, N1856, N358);
not NOT1 (N1887, N1886);
not NOT1 (N1888, N1869);
nor NOR4 (N1889, N1860, N1142, N378, N1505);
and AND2 (N1890, N1888, N509);
nand NAND2 (N1891, N1883, N363);
xor XOR2 (N1892, N1891, N659);
and AND2 (N1893, N1875, N564);
nor NOR2 (N1894, N1878, N779);
buf BUF1 (N1895, N1873);
buf BUF1 (N1896, N1892);
nand NAND3 (N1897, N1890, N1150, N433);
buf BUF1 (N1898, N1895);
and AND2 (N1899, N1893, N1345);
or OR3 (N1900, N1889, N554, N1786);
buf BUF1 (N1901, N1881);
buf BUF1 (N1902, N1898);
xor XOR2 (N1903, N1901, N680);
not NOT1 (N1904, N1897);
nand NAND4 (N1905, N1904, N146, N1880, N1024);
xor XOR2 (N1906, N1896, N1383);
and AND3 (N1907, N1884, N922, N64);
buf BUF1 (N1908, N1900);
or OR3 (N1909, N1905, N1021, N1710);
nor NOR2 (N1910, N1907, N444);
not NOT1 (N1911, N1908);
buf BUF1 (N1912, N1906);
xor XOR2 (N1913, N1909, N975);
or OR2 (N1914, N1885, N890);
nor NOR4 (N1915, N1902, N631, N1298, N852);
nor NOR2 (N1916, N1911, N137);
nor NOR4 (N1917, N1912, N964, N1082, N1712);
and AND4 (N1918, N1903, N1551, N1172, N661);
nor NOR4 (N1919, N1915, N601, N155, N1322);
nor NOR3 (N1920, N1917, N647, N1026);
xor XOR2 (N1921, N1887, N492);
nand NAND4 (N1922, N1921, N276, N714, N1334);
not NOT1 (N1923, N1894);
or OR2 (N1924, N1918, N1572);
and AND3 (N1925, N1914, N1744, N420);
buf BUF1 (N1926, N1919);
nor NOR4 (N1927, N1910, N798, N236, N645);
buf BUF1 (N1928, N1927);
xor XOR2 (N1929, N1922, N942);
and AND2 (N1930, N1924, N1454);
or OR2 (N1931, N1929, N842);
nor NOR3 (N1932, N1923, N781, N211);
not NOT1 (N1933, N1931);
and AND3 (N1934, N1925, N370, N1145);
not NOT1 (N1935, N1930);
or OR4 (N1936, N1916, N1637, N507, N1187);
xor XOR2 (N1937, N1928, N773);
xor XOR2 (N1938, N1899, N1655);
nand NAND4 (N1939, N1932, N674, N1326, N1928);
nor NOR4 (N1940, N1920, N403, N606, N811);
xor XOR2 (N1941, N1936, N854);
or OR4 (N1942, N1941, N574, N1350, N455);
buf BUF1 (N1943, N1938);
nand NAND2 (N1944, N1935, N58);
not NOT1 (N1945, N1913);
and AND3 (N1946, N1934, N755, N736);
not NOT1 (N1947, N1937);
or OR2 (N1948, N1946, N1410);
nor NOR2 (N1949, N1948, N1942);
buf BUF1 (N1950, N1564);
and AND4 (N1951, N1949, N222, N515, N1567);
nor NOR2 (N1952, N1939, N315);
nor NOR2 (N1953, N1943, N803);
and AND4 (N1954, N1933, N1076, N1370, N935);
and AND4 (N1955, N1926, N663, N125, N80);
and AND4 (N1956, N1954, N693, N778, N1058);
nor NOR3 (N1957, N1945, N1128, N396);
or OR4 (N1958, N1950, N399, N250, N1848);
and AND4 (N1959, N1940, N1525, N1425, N260);
or OR4 (N1960, N1959, N186, N1705, N1907);
nand NAND2 (N1961, N1957, N1838);
xor XOR2 (N1962, N1961, N1648);
or OR3 (N1963, N1958, N1790, N1166);
or OR4 (N1964, N1955, N727, N881, N1379);
not NOT1 (N1965, N1952);
and AND4 (N1966, N1965, N645, N957, N1836);
nand NAND4 (N1967, N1966, N600, N239, N80);
and AND3 (N1968, N1951, N184, N59);
or OR2 (N1969, N1944, N798);
xor XOR2 (N1970, N1953, N242);
or OR3 (N1971, N1967, N1623, N1940);
xor XOR2 (N1972, N1971, N1815);
buf BUF1 (N1973, N1963);
or OR2 (N1974, N1970, N682);
nor NOR2 (N1975, N1956, N87);
not NOT1 (N1976, N1960);
nor NOR2 (N1977, N1975, N1493);
not NOT1 (N1978, N1973);
xor XOR2 (N1979, N1972, N702);
not NOT1 (N1980, N1962);
or OR3 (N1981, N1947, N49, N261);
nand NAND3 (N1982, N1976, N1778, N1884);
buf BUF1 (N1983, N1981);
xor XOR2 (N1984, N1968, N1756);
nand NAND3 (N1985, N1980, N1133, N189);
nor NOR2 (N1986, N1978, N1857);
xor XOR2 (N1987, N1984, N1773);
xor XOR2 (N1988, N1985, N209);
nor NOR4 (N1989, N1982, N1376, N1209, N1971);
or OR2 (N1990, N1987, N979);
nor NOR4 (N1991, N1977, N508, N1532, N1863);
or OR3 (N1992, N1969, N1214, N1975);
or OR2 (N1993, N1992, N830);
nand NAND4 (N1994, N1986, N245, N1817, N1245);
not NOT1 (N1995, N1974);
and AND2 (N1996, N1983, N1292);
nand NAND3 (N1997, N1988, N1037, N873);
or OR3 (N1998, N1979, N261, N1220);
nand NAND3 (N1999, N1997, N992, N233);
and AND4 (N2000, N1995, N298, N1299, N1780);
buf BUF1 (N2001, N1994);
and AND4 (N2002, N1990, N1949, N45, N471);
nor NOR4 (N2003, N2002, N427, N323, N1464);
buf BUF1 (N2004, N1964);
nor NOR2 (N2005, N2001, N1457);
or OR4 (N2006, N1993, N197, N1546, N170);
xor XOR2 (N2007, N2000, N1668);
or OR3 (N2008, N1998, N385, N1587);
nand NAND2 (N2009, N2005, N589);
nor NOR3 (N2010, N1996, N662, N1056);
buf BUF1 (N2011, N2007);
and AND4 (N2012, N2006, N1720, N1315, N129);
not NOT1 (N2013, N2003);
nor NOR2 (N2014, N2008, N723);
buf BUF1 (N2015, N2010);
xor XOR2 (N2016, N2014, N1794);
and AND4 (N2017, N2012, N1321, N870, N1945);
nand NAND2 (N2018, N2017, N463);
xor XOR2 (N2019, N1999, N678);
and AND2 (N2020, N2013, N1060);
nor NOR3 (N2021, N2020, N34, N1311);
and AND4 (N2022, N2021, N849, N512, N1315);
nor NOR4 (N2023, N2004, N1126, N1481, N1661);
xor XOR2 (N2024, N2016, N58);
not NOT1 (N2025, N2011);
nand NAND3 (N2026, N1991, N642, N1773);
nand NAND4 (N2027, N2026, N1847, N1496, N1975);
nand NAND4 (N2028, N2024, N1590, N990, N306);
buf BUF1 (N2029, N2022);
or OR2 (N2030, N2009, N760);
or OR2 (N2031, N2029, N2028);
not NOT1 (N2032, N596);
nor NOR4 (N2033, N2027, N454, N1639, N988);
nand NAND3 (N2034, N2015, N1168, N1725);
buf BUF1 (N2035, N2034);
not NOT1 (N2036, N2032);
nor NOR2 (N2037, N1989, N1290);
and AND4 (N2038, N2025, N1468, N1970, N864);
and AND4 (N2039, N2030, N828, N329, N443);
not NOT1 (N2040, N2018);
xor XOR2 (N2041, N2031, N1375);
nor NOR4 (N2042, N2035, N792, N1984, N1942);
not NOT1 (N2043, N2039);
xor XOR2 (N2044, N2033, N102);
nand NAND3 (N2045, N2023, N698, N1736);
xor XOR2 (N2046, N2045, N1403);
nand NAND4 (N2047, N2038, N1117, N1891, N746);
nand NAND3 (N2048, N2036, N1844, N994);
nor NOR3 (N2049, N2048, N727, N1207);
or OR3 (N2050, N2042, N469, N199);
nor NOR4 (N2051, N2037, N1854, N422, N1515);
not NOT1 (N2052, N2051);
nor NOR2 (N2053, N2047, N1501);
buf BUF1 (N2054, N2052);
or OR4 (N2055, N2050, N109, N321, N916);
not NOT1 (N2056, N2046);
and AND3 (N2057, N2049, N462, N356);
or OR2 (N2058, N2044, N676);
nand NAND2 (N2059, N2043, N1302);
and AND4 (N2060, N2055, N1370, N91, N1177);
buf BUF1 (N2061, N2058);
or OR4 (N2062, N2053, N739, N469, N1227);
nand NAND2 (N2063, N2056, N1629);
and AND2 (N2064, N2061, N243);
or OR3 (N2065, N2054, N1107, N1005);
and AND3 (N2066, N2060, N457, N893);
nor NOR3 (N2067, N2041, N1072, N88);
or OR2 (N2068, N2057, N1423);
nor NOR2 (N2069, N2019, N676);
xor XOR2 (N2070, N2064, N1214);
or OR3 (N2071, N2066, N1444, N1657);
nor NOR2 (N2072, N2062, N837);
buf BUF1 (N2073, N2068);
not NOT1 (N2074, N2072);
buf BUF1 (N2075, N2069);
not NOT1 (N2076, N2073);
not NOT1 (N2077, N2059);
or OR4 (N2078, N2067, N1280, N592, N804);
and AND4 (N2079, N2078, N563, N1936, N93);
xor XOR2 (N2080, N2070, N229);
or OR4 (N2081, N2076, N1863, N363, N268);
xor XOR2 (N2082, N2080, N468);
nor NOR2 (N2083, N2040, N608);
and AND2 (N2084, N2082, N773);
and AND4 (N2085, N2065, N692, N786, N1881);
and AND3 (N2086, N2083, N633, N774);
and AND3 (N2087, N2081, N1958, N781);
not NOT1 (N2088, N2079);
buf BUF1 (N2089, N2086);
or OR2 (N2090, N2074, N1805);
buf BUF1 (N2091, N2063);
and AND2 (N2092, N2084, N260);
xor XOR2 (N2093, N2075, N637);
xor XOR2 (N2094, N2091, N1730);
buf BUF1 (N2095, N2085);
xor XOR2 (N2096, N2093, N528);
and AND2 (N2097, N2092, N1051);
nand NAND3 (N2098, N2094, N1835, N552);
nor NOR2 (N2099, N2089, N1170);
nand NAND4 (N2100, N2098, N578, N1780, N1120);
or OR3 (N2101, N2097, N450, N234);
buf BUF1 (N2102, N2090);
or OR2 (N2103, N2087, N770);
not NOT1 (N2104, N2096);
or OR3 (N2105, N2104, N120, N1237);
xor XOR2 (N2106, N2103, N1866);
buf BUF1 (N2107, N2101);
or OR4 (N2108, N2102, N614, N1972, N844);
or OR4 (N2109, N2071, N2035, N1313, N1684);
or OR2 (N2110, N2088, N1797);
xor XOR2 (N2111, N2106, N1706);
and AND4 (N2112, N2110, N393, N1659, N1190);
nand NAND4 (N2113, N2095, N1018, N2058, N1949);
or OR2 (N2114, N2109, N1155);
not NOT1 (N2115, N2112);
nand NAND2 (N2116, N2111, N356);
or OR4 (N2117, N2115, N650, N734, N1406);
xor XOR2 (N2118, N2114, N555);
buf BUF1 (N2119, N2116);
and AND4 (N2120, N2108, N189, N2056, N1593);
nand NAND2 (N2121, N2077, N780);
and AND3 (N2122, N2105, N1108, N581);
xor XOR2 (N2123, N2121, N1247);
or OR2 (N2124, N2099, N116);
not NOT1 (N2125, N2123);
or OR2 (N2126, N2124, N1494);
nand NAND3 (N2127, N2119, N785, N958);
or OR4 (N2128, N2117, N774, N608, N1860);
not NOT1 (N2129, N2125);
and AND2 (N2130, N2128, N1942);
not NOT1 (N2131, N2100);
and AND2 (N2132, N2107, N661);
buf BUF1 (N2133, N2129);
xor XOR2 (N2134, N2130, N1851);
nor NOR4 (N2135, N2122, N919, N1909, N424);
not NOT1 (N2136, N2127);
not NOT1 (N2137, N2135);
nand NAND4 (N2138, N2126, N1219, N2006, N2005);
nor NOR4 (N2139, N2138, N1854, N314, N1432);
xor XOR2 (N2140, N2118, N1127);
or OR2 (N2141, N2139, N1686);
buf BUF1 (N2142, N2137);
nor NOR2 (N2143, N2132, N282);
xor XOR2 (N2144, N2142, N1551);
or OR4 (N2145, N2131, N231, N2118, N5);
nand NAND3 (N2146, N2140, N743, N1926);
and AND2 (N2147, N2134, N2129);
buf BUF1 (N2148, N2120);
nor NOR3 (N2149, N2147, N1438, N1680);
or OR3 (N2150, N2144, N426, N275);
not NOT1 (N2151, N2146);
or OR3 (N2152, N2113, N794, N2009);
buf BUF1 (N2153, N2136);
xor XOR2 (N2154, N2150, N1178);
not NOT1 (N2155, N2141);
not NOT1 (N2156, N2155);
nand NAND2 (N2157, N2148, N1040);
nor NOR2 (N2158, N2154, N1553);
xor XOR2 (N2159, N2133, N171);
nor NOR3 (N2160, N2158, N1684, N50);
nand NAND2 (N2161, N2151, N1013);
nor NOR3 (N2162, N2161, N1826, N1903);
nand NAND2 (N2163, N2153, N258);
nand NAND3 (N2164, N2160, N1212, N742);
and AND4 (N2165, N2163, N2132, N673, N2146);
and AND3 (N2166, N2164, N1397, N848);
buf BUF1 (N2167, N2156);
not NOT1 (N2168, N2165);
or OR2 (N2169, N2157, N931);
xor XOR2 (N2170, N2149, N1856);
xor XOR2 (N2171, N2166, N324);
or OR2 (N2172, N2145, N1974);
or OR3 (N2173, N2167, N256, N437);
xor XOR2 (N2174, N2143, N863);
nor NOR4 (N2175, N2159, N1826, N1153, N782);
and AND2 (N2176, N2174, N1747);
or OR4 (N2177, N2162, N299, N1344, N1837);
nand NAND2 (N2178, N2173, N315);
or OR3 (N2179, N2152, N1949, N494);
or OR3 (N2180, N2170, N215, N868);
or OR2 (N2181, N2168, N1270);
and AND3 (N2182, N2175, N809, N1061);
nand NAND4 (N2183, N2176, N1914, N301, N1476);
nand NAND4 (N2184, N2180, N1671, N609, N704);
nor NOR2 (N2185, N2172, N2170);
not NOT1 (N2186, N2169);
nor NOR4 (N2187, N2171, N1062, N1522, N1908);
or OR4 (N2188, N2183, N2019, N1725, N1483);
and AND4 (N2189, N2179, N1263, N651, N832);
not NOT1 (N2190, N2182);
or OR2 (N2191, N2186, N55);
buf BUF1 (N2192, N2178);
or OR4 (N2193, N2188, N11, N1060, N706);
nand NAND2 (N2194, N2181, N955);
not NOT1 (N2195, N2185);
or OR4 (N2196, N2195, N616, N469, N81);
and AND2 (N2197, N2189, N1224);
xor XOR2 (N2198, N2192, N1361);
or OR2 (N2199, N2177, N242);
not NOT1 (N2200, N2193);
and AND2 (N2201, N2184, N1010);
not NOT1 (N2202, N2201);
nand NAND3 (N2203, N2199, N173, N943);
xor XOR2 (N2204, N2203, N1947);
xor XOR2 (N2205, N2202, N118);
buf BUF1 (N2206, N2200);
buf BUF1 (N2207, N2204);
nand NAND2 (N2208, N2205, N679);
xor XOR2 (N2209, N2208, N1207);
xor XOR2 (N2210, N2196, N157);
not NOT1 (N2211, N2194);
nand NAND2 (N2212, N2187, N720);
not NOT1 (N2213, N2212);
or OR4 (N2214, N2211, N1258, N892, N1345);
and AND2 (N2215, N2191, N2109);
xor XOR2 (N2216, N2198, N11);
or OR4 (N2217, N2215, N1968, N651, N1355);
and AND3 (N2218, N2216, N218, N1647);
nor NOR3 (N2219, N2210, N692, N96);
nand NAND3 (N2220, N2214, N1033, N341);
or OR3 (N2221, N2190, N1854, N1687);
buf BUF1 (N2222, N2218);
xor XOR2 (N2223, N2209, N200);
and AND4 (N2224, N2222, N2118, N1461, N1043);
and AND4 (N2225, N2220, N1169, N1324, N130);
nor NOR2 (N2226, N2213, N601);
nor NOR4 (N2227, N2224, N1234, N1906, N546);
nor NOR4 (N2228, N2223, N2204, N457, N2060);
nand NAND3 (N2229, N2228, N2227, N344);
xor XOR2 (N2230, N285, N345);
not NOT1 (N2231, N2221);
and AND3 (N2232, N2230, N1396, N1736);
nor NOR3 (N2233, N2219, N1809, N1654);
buf BUF1 (N2234, N2229);
nor NOR4 (N2235, N2225, N1704, N739, N270);
nand NAND3 (N2236, N2207, N2151, N192);
or OR4 (N2237, N2197, N2165, N1840, N840);
not NOT1 (N2238, N2234);
and AND4 (N2239, N2217, N101, N1059, N1723);
or OR4 (N2240, N2235, N428, N2212, N1721);
or OR3 (N2241, N2232, N387, N1002);
nor NOR2 (N2242, N2238, N390);
not NOT1 (N2243, N2242);
not NOT1 (N2244, N2236);
or OR4 (N2245, N2243, N1523, N129, N452);
not NOT1 (N2246, N2241);
not NOT1 (N2247, N2244);
nor NOR2 (N2248, N2247, N551);
or OR2 (N2249, N2240, N904);
not NOT1 (N2250, N2226);
or OR3 (N2251, N2250, N1083, N7);
and AND3 (N2252, N2248, N2232, N789);
not NOT1 (N2253, N2206);
and AND3 (N2254, N2251, N2137, N1798);
xor XOR2 (N2255, N2239, N1850);
or OR4 (N2256, N2231, N377, N2206, N1923);
buf BUF1 (N2257, N2252);
and AND4 (N2258, N2257, N1724, N1913, N1517);
and AND2 (N2259, N2246, N2229);
buf BUF1 (N2260, N2255);
or OR4 (N2261, N2237, N1777, N2060, N2186);
nor NOR3 (N2262, N2261, N1979, N1330);
nand NAND2 (N2263, N2256, N704);
and AND4 (N2264, N2249, N20, N105, N1012);
nand NAND3 (N2265, N2258, N1353, N59);
and AND2 (N2266, N2253, N894);
and AND2 (N2267, N2262, N296);
nor NOR4 (N2268, N2260, N1748, N2065, N1350);
buf BUF1 (N2269, N2267);
nor NOR4 (N2270, N2266, N502, N1341, N1723);
xor XOR2 (N2271, N2265, N1368);
and AND2 (N2272, N2268, N88);
not NOT1 (N2273, N2259);
xor XOR2 (N2274, N2272, N2079);
nor NOR3 (N2275, N2269, N1592, N209);
nor NOR4 (N2276, N2271, N1536, N402, N1548);
nor NOR4 (N2277, N2276, N81, N40, N1725);
xor XOR2 (N2278, N2264, N689);
buf BUF1 (N2279, N2263);
and AND2 (N2280, N2233, N1924);
buf BUF1 (N2281, N2273);
nor NOR4 (N2282, N2254, N729, N650, N1521);
nand NAND3 (N2283, N2274, N18, N1437);
or OR3 (N2284, N2270, N1917, N1548);
nand NAND2 (N2285, N2281, N1042);
or OR2 (N2286, N2283, N587);
or OR3 (N2287, N2286, N1616, N509);
nand NAND2 (N2288, N2245, N1457);
not NOT1 (N2289, N2287);
xor XOR2 (N2290, N2284, N820);
nor NOR4 (N2291, N2288, N1214, N164, N666);
not NOT1 (N2292, N2280);
buf BUF1 (N2293, N2277);
nor NOR3 (N2294, N2285, N2157, N1920);
buf BUF1 (N2295, N2282);
and AND2 (N2296, N2292, N808);
nand NAND2 (N2297, N2293, N678);
nor NOR2 (N2298, N2278, N1301);
nand NAND2 (N2299, N2291, N721);
nor NOR2 (N2300, N2294, N1363);
nor NOR3 (N2301, N2275, N1650, N851);
or OR3 (N2302, N2279, N1562, N1019);
not NOT1 (N2303, N2301);
nand NAND2 (N2304, N2300, N1054);
or OR2 (N2305, N2299, N631);
buf BUF1 (N2306, N2295);
and AND3 (N2307, N2306, N19, N369);
and AND2 (N2308, N2296, N298);
nand NAND3 (N2309, N2308, N784, N2042);
nand NAND4 (N2310, N2309, N1794, N680, N1637);
xor XOR2 (N2311, N2297, N1902);
nand NAND3 (N2312, N2303, N2244, N1472);
not NOT1 (N2313, N2289);
nor NOR3 (N2314, N2305, N1771, N781);
or OR3 (N2315, N2290, N2001, N674);
and AND2 (N2316, N2311, N863);
not NOT1 (N2317, N2315);
or OR2 (N2318, N2302, N821);
or OR4 (N2319, N2314, N898, N973, N483);
and AND3 (N2320, N2319, N1277, N1847);
or OR3 (N2321, N2317, N190, N1111);
and AND3 (N2322, N2318, N449, N713);
nor NOR4 (N2323, N2298, N1445, N1732, N2246);
nand NAND2 (N2324, N2321, N1046);
nor NOR4 (N2325, N2307, N1934, N573, N1198);
nor NOR3 (N2326, N2312, N215, N1723);
nand NAND2 (N2327, N2316, N607);
nand NAND4 (N2328, N2322, N226, N432, N2009);
not NOT1 (N2329, N2325);
and AND2 (N2330, N2326, N1064);
nand NAND4 (N2331, N2310, N1808, N1726, N39);
nand NAND2 (N2332, N2324, N1003);
xor XOR2 (N2333, N2329, N354);
or OR4 (N2334, N2323, N2135, N648, N1606);
and AND4 (N2335, N2320, N763, N639, N568);
or OR3 (N2336, N2304, N1615, N190);
xor XOR2 (N2337, N2327, N705);
xor XOR2 (N2338, N2336, N1654);
xor XOR2 (N2339, N2338, N1199);
nor NOR3 (N2340, N2337, N129, N234);
and AND3 (N2341, N2335, N1385, N2088);
and AND2 (N2342, N2334, N261);
nor NOR2 (N2343, N2342, N1711);
nor NOR2 (N2344, N2333, N631);
or OR2 (N2345, N2330, N821);
not NOT1 (N2346, N2341);
not NOT1 (N2347, N2331);
xor XOR2 (N2348, N2346, N1799);
xor XOR2 (N2349, N2313, N708);
not NOT1 (N2350, N2349);
nand NAND4 (N2351, N2340, N1045, N1897, N2083);
nand NAND3 (N2352, N2339, N707, N1801);
nand NAND2 (N2353, N2352, N2349);
nand NAND3 (N2354, N2345, N2353, N15);
xor XOR2 (N2355, N626, N1782);
not NOT1 (N2356, N2332);
and AND4 (N2357, N2356, N686, N1270, N1960);
nand NAND4 (N2358, N2344, N139, N606, N1335);
nand NAND3 (N2359, N2357, N1951, N2238);
nor NOR4 (N2360, N2347, N2197, N878, N1812);
or OR3 (N2361, N2355, N150, N964);
buf BUF1 (N2362, N2360);
buf BUF1 (N2363, N2354);
buf BUF1 (N2364, N2343);
nand NAND3 (N2365, N2348, N1903, N1501);
not NOT1 (N2366, N2364);
nand NAND4 (N2367, N2351, N1101, N1167, N722);
buf BUF1 (N2368, N2358);
or OR2 (N2369, N2362, N1711);
nor NOR2 (N2370, N2366, N1882);
not NOT1 (N2371, N2363);
xor XOR2 (N2372, N2350, N962);
and AND3 (N2373, N2367, N2211, N906);
buf BUF1 (N2374, N2359);
buf BUF1 (N2375, N2365);
not NOT1 (N2376, N2368);
nor NOR2 (N2377, N2369, N531);
nand NAND3 (N2378, N2374, N162, N1368);
and AND2 (N2379, N2376, N2157);
nand NAND4 (N2380, N2372, N1539, N223, N1909);
nor NOR4 (N2381, N2380, N2055, N2347, N319);
or OR2 (N2382, N2373, N1410);
or OR3 (N2383, N2371, N911, N863);
not NOT1 (N2384, N2378);
nor NOR3 (N2385, N2382, N2165, N2320);
nor NOR4 (N2386, N2379, N163, N1, N2381);
xor XOR2 (N2387, N216, N572);
buf BUF1 (N2388, N2385);
nand NAND3 (N2389, N2386, N1980, N1956);
buf BUF1 (N2390, N2388);
or OR2 (N2391, N2390, N695);
xor XOR2 (N2392, N2389, N1914);
nand NAND4 (N2393, N2387, N1854, N1043, N1591);
and AND2 (N2394, N2370, N1065);
not NOT1 (N2395, N2392);
xor XOR2 (N2396, N2383, N2209);
not NOT1 (N2397, N2396);
nor NOR2 (N2398, N2393, N1183);
buf BUF1 (N2399, N2361);
or OR4 (N2400, N2399, N1141, N2062, N988);
buf BUF1 (N2401, N2384);
xor XOR2 (N2402, N2391, N1154);
nor NOR4 (N2403, N2402, N1676, N794, N917);
and AND4 (N2404, N2395, N568, N1613, N2163);
buf BUF1 (N2405, N2401);
and AND3 (N2406, N2400, N60, N148);
not NOT1 (N2407, N2375);
not NOT1 (N2408, N2405);
nor NOR2 (N2409, N2377, N1220);
buf BUF1 (N2410, N2406);
not NOT1 (N2411, N2409);
nand NAND2 (N2412, N2408, N302);
or OR4 (N2413, N2397, N1531, N355, N1374);
and AND3 (N2414, N2328, N1707, N2100);
nor NOR2 (N2415, N2403, N1346);
nor NOR3 (N2416, N2413, N1769, N2373);
buf BUF1 (N2417, N2412);
and AND4 (N2418, N2394, N1709, N1082, N850);
and AND2 (N2419, N2404, N841);
buf BUF1 (N2420, N2415);
nor NOR3 (N2421, N2419, N1927, N115);
or OR3 (N2422, N2398, N1210, N1691);
nand NAND2 (N2423, N2417, N648);
nor NOR2 (N2424, N2422, N302);
xor XOR2 (N2425, N2423, N1309);
nand NAND4 (N2426, N2407, N431, N290, N240);
buf BUF1 (N2427, N2410);
not NOT1 (N2428, N2427);
buf BUF1 (N2429, N2418);
buf BUF1 (N2430, N2424);
and AND4 (N2431, N2416, N2258, N2367, N701);
buf BUF1 (N2432, N2428);
and AND4 (N2433, N2430, N403, N2172, N2363);
nand NAND2 (N2434, N2431, N1209);
and AND2 (N2435, N2420, N379);
and AND4 (N2436, N2421, N591, N241, N495);
xor XOR2 (N2437, N2429, N1839);
and AND4 (N2438, N2414, N347, N1078, N269);
and AND4 (N2439, N2426, N577, N2166, N289);
xor XOR2 (N2440, N2435, N861);
or OR2 (N2441, N2425, N1155);
buf BUF1 (N2442, N2441);
nand NAND4 (N2443, N2437, N1834, N271, N530);
and AND3 (N2444, N2442, N687, N210);
or OR2 (N2445, N2432, N1249);
nor NOR2 (N2446, N2411, N1135);
xor XOR2 (N2447, N2440, N1987);
not NOT1 (N2448, N2436);
buf BUF1 (N2449, N2448);
or OR3 (N2450, N2449, N656, N851);
not NOT1 (N2451, N2439);
buf BUF1 (N2452, N2445);
buf BUF1 (N2453, N2434);
nor NOR3 (N2454, N2452, N107, N1218);
xor XOR2 (N2455, N2433, N2033);
buf BUF1 (N2456, N2446);
nand NAND4 (N2457, N2451, N1714, N740, N1533);
nor NOR3 (N2458, N2443, N2354, N852);
not NOT1 (N2459, N2447);
and AND4 (N2460, N2458, N1996, N280, N1250);
xor XOR2 (N2461, N2453, N2251);
or OR3 (N2462, N2444, N391, N1858);
nand NAND3 (N2463, N2455, N1680, N1718);
not NOT1 (N2464, N2438);
xor XOR2 (N2465, N2450, N717);
buf BUF1 (N2466, N2459);
and AND3 (N2467, N2462, N1992, N1284);
nor NOR4 (N2468, N2463, N1113, N1114, N1823);
or OR4 (N2469, N2461, N2248, N863, N973);
nor NOR3 (N2470, N2454, N651, N917);
xor XOR2 (N2471, N2457, N1132);
nor NOR4 (N2472, N2456, N1896, N1687, N1303);
nand NAND2 (N2473, N2460, N358);
not NOT1 (N2474, N2465);
buf BUF1 (N2475, N2472);
buf BUF1 (N2476, N2466);
xor XOR2 (N2477, N2470, N2425);
and AND3 (N2478, N2471, N2305, N1340);
or OR4 (N2479, N2468, N345, N861, N1460);
not NOT1 (N2480, N2479);
nor NOR4 (N2481, N2474, N267, N2212, N145);
and AND2 (N2482, N2475, N1096);
nand NAND2 (N2483, N2482, N629);
and AND4 (N2484, N2480, N2255, N321, N1691);
xor XOR2 (N2485, N2473, N1064);
or OR4 (N2486, N2478, N325, N1056, N993);
and AND2 (N2487, N2485, N2376);
or OR2 (N2488, N2481, N2383);
and AND4 (N2489, N2464, N344, N723, N551);
buf BUF1 (N2490, N2477);
not NOT1 (N2491, N2488);
xor XOR2 (N2492, N2491, N1413);
nor NOR4 (N2493, N2483, N1365, N680, N1571);
not NOT1 (N2494, N2486);
nand NAND3 (N2495, N2489, N1189, N1462);
not NOT1 (N2496, N2490);
not NOT1 (N2497, N2494);
nand NAND3 (N2498, N2467, N1861, N1512);
and AND3 (N2499, N2496, N2320, N70);
buf BUF1 (N2500, N2487);
not NOT1 (N2501, N2498);
nand NAND2 (N2502, N2476, N1648);
xor XOR2 (N2503, N2493, N496);
not NOT1 (N2504, N2497);
nor NOR4 (N2505, N2495, N2458, N2128, N1189);
nor NOR4 (N2506, N2500, N912, N972, N375);
buf BUF1 (N2507, N2499);
buf BUF1 (N2508, N2501);
not NOT1 (N2509, N2506);
not NOT1 (N2510, N2505);
not NOT1 (N2511, N2509);
nor NOR4 (N2512, N2492, N271, N584, N637);
not NOT1 (N2513, N2512);
and AND4 (N2514, N2502, N271, N337, N291);
buf BUF1 (N2515, N2469);
nor NOR4 (N2516, N2508, N1779, N1716, N2207);
nor NOR2 (N2517, N2510, N789);
nor NOR3 (N2518, N2514, N1392, N1445);
or OR2 (N2519, N2504, N2147);
nor NOR2 (N2520, N2513, N1169);
nor NOR4 (N2521, N2503, N1579, N516, N1806);
buf BUF1 (N2522, N2519);
nand NAND4 (N2523, N2516, N2027, N44, N1868);
buf BUF1 (N2524, N2522);
buf BUF1 (N2525, N2523);
xor XOR2 (N2526, N2518, N1707);
buf BUF1 (N2527, N2507);
nand NAND2 (N2528, N2525, N2174);
xor XOR2 (N2529, N2524, N2335);
or OR4 (N2530, N2484, N789, N1355, N300);
buf BUF1 (N2531, N2520);
not NOT1 (N2532, N2530);
nand NAND2 (N2533, N2529, N91);
or OR3 (N2534, N2533, N745, N61);
not NOT1 (N2535, N2527);
buf BUF1 (N2536, N2521);
or OR2 (N2537, N2535, N1387);
nand NAND3 (N2538, N2537, N1978, N356);
or OR2 (N2539, N2534, N2182);
buf BUF1 (N2540, N2538);
nor NOR4 (N2541, N2511, N2240, N196, N2392);
and AND2 (N2542, N2515, N2367);
not NOT1 (N2543, N2539);
buf BUF1 (N2544, N2531);
and AND4 (N2545, N2543, N1661, N26, N327);
buf BUF1 (N2546, N2544);
buf BUF1 (N2547, N2528);
buf BUF1 (N2548, N2545);
nand NAND3 (N2549, N2548, N539, N2315);
nor NOR3 (N2550, N2542, N153, N571);
xor XOR2 (N2551, N2536, N2152);
nand NAND3 (N2552, N2526, N1207, N2265);
nand NAND3 (N2553, N2532, N326, N929);
and AND4 (N2554, N2552, N500, N264, N2066);
or OR4 (N2555, N2554, N1890, N2346, N77);
nor NOR2 (N2556, N2517, N2022);
and AND2 (N2557, N2541, N970);
or OR2 (N2558, N2553, N2419);
or OR3 (N2559, N2555, N509, N1394);
nand NAND4 (N2560, N2540, N2349, N286, N1542);
or OR3 (N2561, N2560, N1792, N796);
xor XOR2 (N2562, N2550, N515);
buf BUF1 (N2563, N2559);
xor XOR2 (N2564, N2549, N1472);
and AND4 (N2565, N2561, N1673, N2308, N2478);
buf BUF1 (N2566, N2562);
buf BUF1 (N2567, N2564);
and AND2 (N2568, N2566, N2031);
xor XOR2 (N2569, N2551, N7);
nand NAND2 (N2570, N2558, N2271);
not NOT1 (N2571, N2570);
nand NAND2 (N2572, N2547, N775);
and AND2 (N2573, N2567, N273);
nand NAND3 (N2574, N2572, N2041, N650);
xor XOR2 (N2575, N2574, N31);
xor XOR2 (N2576, N2575, N269);
not NOT1 (N2577, N2557);
nand NAND2 (N2578, N2577, N1611);
nor NOR3 (N2579, N2568, N2030, N631);
and AND2 (N2580, N2546, N1697);
nor NOR2 (N2581, N2563, N2298);
nand NAND2 (N2582, N2580, N1317);
and AND2 (N2583, N2582, N1080);
nand NAND4 (N2584, N2571, N2044, N1312, N2156);
nor NOR2 (N2585, N2578, N1513);
and AND2 (N2586, N2583, N1632);
or OR2 (N2587, N2585, N33);
not NOT1 (N2588, N2584);
buf BUF1 (N2589, N2569);
nor NOR3 (N2590, N2589, N2426, N262);
nor NOR2 (N2591, N2588, N497);
buf BUF1 (N2592, N2590);
buf BUF1 (N2593, N2586);
and AND2 (N2594, N2592, N200);
and AND2 (N2595, N2587, N1203);
xor XOR2 (N2596, N2579, N621);
xor XOR2 (N2597, N2565, N747);
not NOT1 (N2598, N2597);
or OR3 (N2599, N2593, N1171, N1346);
nor NOR4 (N2600, N2598, N1990, N1903, N353);
not NOT1 (N2601, N2581);
nor NOR4 (N2602, N2601, N413, N1364, N2049);
nand NAND4 (N2603, N2600, N1469, N835, N4);
and AND2 (N2604, N2603, N1355);
or OR2 (N2605, N2594, N142);
nand NAND4 (N2606, N2595, N2307, N1060, N562);
buf BUF1 (N2607, N2599);
nand NAND2 (N2608, N2607, N2424);
not NOT1 (N2609, N2556);
and AND2 (N2610, N2608, N1339);
nor NOR2 (N2611, N2605, N2505);
and AND2 (N2612, N2611, N128);
nor NOR2 (N2613, N2610, N876);
nor NOR4 (N2614, N2573, N919, N358, N2101);
buf BUF1 (N2615, N2612);
not NOT1 (N2616, N2576);
buf BUF1 (N2617, N2604);
xor XOR2 (N2618, N2591, N2118);
xor XOR2 (N2619, N2602, N747);
not NOT1 (N2620, N2614);
xor XOR2 (N2621, N2613, N516);
and AND4 (N2622, N2616, N1420, N1316, N2001);
nand NAND3 (N2623, N2618, N1350, N1227);
and AND4 (N2624, N2617, N411, N908, N1038);
nand NAND4 (N2625, N2615, N1147, N1416, N1701);
nor NOR2 (N2626, N2625, N589);
xor XOR2 (N2627, N2626, N2070);
or OR3 (N2628, N2619, N828, N2125);
buf BUF1 (N2629, N2624);
not NOT1 (N2630, N2629);
not NOT1 (N2631, N2628);
not NOT1 (N2632, N2630);
nand NAND3 (N2633, N2627, N83, N1643);
nand NAND4 (N2634, N2632, N1602, N2547, N1092);
and AND3 (N2635, N2622, N1539, N1440);
nand NAND3 (N2636, N2621, N40, N2296);
nor NOR3 (N2637, N2633, N2574, N2218);
nand NAND3 (N2638, N2596, N1050, N2409);
nor NOR4 (N2639, N2636, N1598, N1763, N862);
nand NAND3 (N2640, N2638, N638, N454);
or OR2 (N2641, N2640, N1932);
not NOT1 (N2642, N2631);
or OR4 (N2643, N2639, N653, N884, N92);
not NOT1 (N2644, N2641);
and AND2 (N2645, N2623, N1654);
nor NOR2 (N2646, N2643, N2011);
nor NOR4 (N2647, N2609, N124, N1131, N2553);
nor NOR4 (N2648, N2647, N635, N137, N1438);
not NOT1 (N2649, N2606);
nand NAND3 (N2650, N2637, N2057, N1852);
nand NAND3 (N2651, N2635, N1344, N2511);
or OR3 (N2652, N2649, N893, N745);
buf BUF1 (N2653, N2620);
nand NAND3 (N2654, N2651, N2472, N231);
and AND2 (N2655, N2653, N804);
or OR3 (N2656, N2650, N2616, N186);
nand NAND3 (N2657, N2656, N437, N2411);
xor XOR2 (N2658, N2655, N112);
nand NAND3 (N2659, N2645, N1096, N2478);
not NOT1 (N2660, N2646);
nand NAND3 (N2661, N2652, N960, N1873);
xor XOR2 (N2662, N2642, N271);
buf BUF1 (N2663, N2662);
buf BUF1 (N2664, N2648);
and AND3 (N2665, N2634, N707, N1134);
xor XOR2 (N2666, N2659, N987);
or OR3 (N2667, N2665, N1706, N2389);
xor XOR2 (N2668, N2654, N696);
xor XOR2 (N2669, N2668, N376);
or OR2 (N2670, N2667, N1769);
buf BUF1 (N2671, N2660);
nand NAND3 (N2672, N2666, N1258, N881);
not NOT1 (N2673, N2657);
not NOT1 (N2674, N2663);
or OR2 (N2675, N2644, N1916);
and AND3 (N2676, N2664, N1495, N366);
xor XOR2 (N2677, N2658, N1824);
not NOT1 (N2678, N2669);
and AND2 (N2679, N2678, N1294);
not NOT1 (N2680, N2672);
nor NOR2 (N2681, N2673, N663);
or OR2 (N2682, N2676, N43);
not NOT1 (N2683, N2679);
and AND4 (N2684, N2677, N1717, N1776, N1012);
not NOT1 (N2685, N2682);
not NOT1 (N2686, N2681);
nor NOR4 (N2687, N2683, N1163, N1832, N2650);
nand NAND3 (N2688, N2670, N837, N710);
not NOT1 (N2689, N2687);
xor XOR2 (N2690, N2674, N2469);
not NOT1 (N2691, N2661);
or OR3 (N2692, N2685, N719, N453);
and AND4 (N2693, N2671, N2306, N166, N737);
not NOT1 (N2694, N2686);
and AND3 (N2695, N2689, N1781, N1187);
not NOT1 (N2696, N2684);
buf BUF1 (N2697, N2688);
buf BUF1 (N2698, N2694);
buf BUF1 (N2699, N2697);
xor XOR2 (N2700, N2695, N2148);
nor NOR3 (N2701, N2698, N1233, N353);
nor NOR3 (N2702, N2699, N164, N574);
not NOT1 (N2703, N2692);
not NOT1 (N2704, N2690);
nor NOR2 (N2705, N2696, N995);
xor XOR2 (N2706, N2693, N2577);
or OR2 (N2707, N2704, N329);
nand NAND3 (N2708, N2675, N1414, N2450);
nor NOR4 (N2709, N2703, N1974, N763, N215);
xor XOR2 (N2710, N2706, N2357);
xor XOR2 (N2711, N2705, N885);
nor NOR3 (N2712, N2707, N365, N710);
nand NAND2 (N2713, N2701, N137);
xor XOR2 (N2714, N2710, N1588);
buf BUF1 (N2715, N2709);
buf BUF1 (N2716, N2713);
nand NAND2 (N2717, N2702, N2627);
or OR3 (N2718, N2711, N1755, N896);
or OR2 (N2719, N2716, N1345);
or OR2 (N2720, N2718, N2579);
and AND3 (N2721, N2700, N214, N888);
and AND3 (N2722, N2717, N2247, N1177);
nor NOR2 (N2723, N2714, N2627);
or OR4 (N2724, N2680, N1442, N2247, N1132);
nor NOR2 (N2725, N2715, N2314);
nor NOR4 (N2726, N2708, N735, N2263, N2244);
or OR4 (N2727, N2723, N1739, N2710, N2268);
nand NAND2 (N2728, N2719, N1603);
not NOT1 (N2729, N2724);
nand NAND4 (N2730, N2729, N141, N122, N2253);
nand NAND2 (N2731, N2725, N2426);
buf BUF1 (N2732, N2728);
and AND3 (N2733, N2720, N1779, N986);
xor XOR2 (N2734, N2712, N2710);
and AND3 (N2735, N2731, N1792, N92);
xor XOR2 (N2736, N2730, N16);
nand NAND2 (N2737, N2733, N2487);
and AND3 (N2738, N2726, N99, N1107);
xor XOR2 (N2739, N2734, N1590);
buf BUF1 (N2740, N2722);
xor XOR2 (N2741, N2740, N1486);
nor NOR4 (N2742, N2721, N1265, N233, N692);
xor XOR2 (N2743, N2691, N214);
or OR4 (N2744, N2738, N138, N2709, N2596);
nor NOR3 (N2745, N2737, N1876, N2410);
xor XOR2 (N2746, N2741, N2369);
nor NOR4 (N2747, N2735, N217, N2645, N1268);
buf BUF1 (N2748, N2736);
nand NAND3 (N2749, N2742, N229, N2200);
buf BUF1 (N2750, N2747);
nand NAND3 (N2751, N2749, N2070, N2189);
nand NAND3 (N2752, N2743, N2435, N325);
xor XOR2 (N2753, N2744, N1915);
nor NOR4 (N2754, N2753, N1182, N2036, N769);
xor XOR2 (N2755, N2739, N1742);
nor NOR4 (N2756, N2746, N340, N868, N1385);
buf BUF1 (N2757, N2745);
nand NAND2 (N2758, N2756, N1206);
or OR2 (N2759, N2751, N2706);
and AND3 (N2760, N2748, N2582, N1538);
or OR3 (N2761, N2760, N2640, N919);
and AND4 (N2762, N2727, N1175, N595, N1833);
nor NOR3 (N2763, N2752, N2008, N2256);
or OR4 (N2764, N2755, N1446, N596, N1054);
buf BUF1 (N2765, N2761);
nor NOR4 (N2766, N2765, N1857, N2067, N2032);
nand NAND4 (N2767, N2750, N2072, N1638, N2399);
nor NOR4 (N2768, N2754, N1047, N724, N243);
not NOT1 (N2769, N2759);
nand NAND2 (N2770, N2768, N1430);
and AND3 (N2771, N2732, N1640, N1566);
xor XOR2 (N2772, N2762, N1759);
nand NAND4 (N2773, N2758, N963, N1813, N380);
buf BUF1 (N2774, N2769);
or OR2 (N2775, N2767, N1319);
or OR4 (N2776, N2773, N209, N1389, N461);
buf BUF1 (N2777, N2764);
or OR3 (N2778, N2766, N2595, N226);
xor XOR2 (N2779, N2777, N1409);
and AND2 (N2780, N2771, N1558);
xor XOR2 (N2781, N2763, N2205);
not NOT1 (N2782, N2775);
and AND3 (N2783, N2757, N1745, N1670);
and AND3 (N2784, N2770, N139, N1859);
not NOT1 (N2785, N2774);
nand NAND2 (N2786, N2785, N1682);
nor NOR3 (N2787, N2786, N2405, N773);
not NOT1 (N2788, N2779);
nand NAND4 (N2789, N2787, N2147, N1534, N771);
or OR4 (N2790, N2772, N1279, N927, N119);
and AND4 (N2791, N2783, N82, N961, N324);
and AND3 (N2792, N2784, N1156, N645);
nand NAND4 (N2793, N2791, N2086, N2529, N1128);
or OR3 (N2794, N2776, N634, N1297);
nand NAND2 (N2795, N2788, N1425);
nor NOR3 (N2796, N2792, N2655, N511);
not NOT1 (N2797, N2781);
nand NAND4 (N2798, N2780, N696, N2491, N863);
nand NAND2 (N2799, N2798, N2694);
nor NOR2 (N2800, N2790, N295);
buf BUF1 (N2801, N2797);
or OR4 (N2802, N2796, N400, N416, N1587);
xor XOR2 (N2803, N2794, N398);
nor NOR3 (N2804, N2799, N1413, N1562);
nand NAND4 (N2805, N2803, N2161, N1733, N203);
xor XOR2 (N2806, N2778, N2556);
buf BUF1 (N2807, N2801);
or OR4 (N2808, N2802, N11, N2021, N1327);
or OR2 (N2809, N2795, N257);
nor NOR4 (N2810, N2806, N2712, N2670, N92);
nor NOR2 (N2811, N2793, N976);
and AND4 (N2812, N2811, N880, N2389, N1424);
nor NOR2 (N2813, N2782, N1909);
and AND3 (N2814, N2789, N2754, N775);
nor NOR3 (N2815, N2810, N2398, N485);
xor XOR2 (N2816, N2805, N1900);
buf BUF1 (N2817, N2804);
nand NAND3 (N2818, N2808, N606, N2149);
nor NOR2 (N2819, N2815, N208);
xor XOR2 (N2820, N2809, N2552);
or OR4 (N2821, N2819, N686, N1604, N870);
nand NAND3 (N2822, N2821, N2150, N1101);
and AND3 (N2823, N2814, N2303, N1973);
xor XOR2 (N2824, N2813, N1163);
xor XOR2 (N2825, N2807, N1322);
nor NOR4 (N2826, N2823, N66, N798, N172);
nor NOR4 (N2827, N2816, N802, N2078, N357);
buf BUF1 (N2828, N2817);
xor XOR2 (N2829, N2825, N336);
not NOT1 (N2830, N2820);
buf BUF1 (N2831, N2824);
buf BUF1 (N2832, N2826);
not NOT1 (N2833, N2828);
nand NAND4 (N2834, N2818, N1552, N1333, N1562);
nand NAND3 (N2835, N2834, N1800, N1262);
nand NAND4 (N2836, N2831, N1040, N1894, N1458);
buf BUF1 (N2837, N2829);
or OR4 (N2838, N2837, N1070, N345, N990);
not NOT1 (N2839, N2830);
nor NOR4 (N2840, N2839, N440, N2390, N2114);
not NOT1 (N2841, N2836);
or OR3 (N2842, N2840, N2125, N1171);
buf BUF1 (N2843, N2832);
and AND4 (N2844, N2827, N2044, N369, N214);
nand NAND2 (N2845, N2843, N2740);
or OR3 (N2846, N2833, N1380, N2476);
and AND4 (N2847, N2845, N2402, N2630, N1798);
and AND4 (N2848, N2842, N1803, N855, N376);
and AND3 (N2849, N2812, N171, N1517);
buf BUF1 (N2850, N2849);
nand NAND2 (N2851, N2838, N789);
not NOT1 (N2852, N2846);
not NOT1 (N2853, N2850);
and AND3 (N2854, N2853, N368, N702);
nor NOR2 (N2855, N2851, N189);
not NOT1 (N2856, N2854);
not NOT1 (N2857, N2844);
nor NOR2 (N2858, N2835, N199);
and AND2 (N2859, N2800, N759);
and AND2 (N2860, N2857, N1479);
buf BUF1 (N2861, N2856);
nand NAND4 (N2862, N2847, N318, N1285, N773);
nor NOR4 (N2863, N2860, N1216, N222, N1392);
buf BUF1 (N2864, N2862);
buf BUF1 (N2865, N2861);
nand NAND4 (N2866, N2822, N1010, N1158, N2416);
xor XOR2 (N2867, N2866, N582);
nor NOR3 (N2868, N2848, N2075, N302);
or OR2 (N2869, N2841, N2623);
buf BUF1 (N2870, N2859);
nand NAND4 (N2871, N2869, N1383, N651, N938);
and AND2 (N2872, N2870, N1091);
or OR2 (N2873, N2855, N1764);
xor XOR2 (N2874, N2858, N1611);
or OR2 (N2875, N2868, N1754);
not NOT1 (N2876, N2863);
and AND4 (N2877, N2864, N920, N802, N2402);
xor XOR2 (N2878, N2865, N826);
nor NOR3 (N2879, N2877, N1, N755);
buf BUF1 (N2880, N2852);
or OR4 (N2881, N2879, N438, N1259, N1576);
nand NAND2 (N2882, N2878, N2863);
and AND2 (N2883, N2867, N2334);
buf BUF1 (N2884, N2881);
xor XOR2 (N2885, N2883, N1518);
or OR3 (N2886, N2873, N2851, N2449);
nand NAND2 (N2887, N2874, N723);
xor XOR2 (N2888, N2876, N208);
nor NOR4 (N2889, N2887, N812, N692, N2158);
and AND3 (N2890, N2871, N2466, N602);
or OR2 (N2891, N2875, N1477);
or OR2 (N2892, N2882, N2386);
xor XOR2 (N2893, N2888, N2229);
or OR2 (N2894, N2884, N1495);
not NOT1 (N2895, N2893);
nor NOR4 (N2896, N2894, N873, N1398, N1728);
xor XOR2 (N2897, N2891, N566);
xor XOR2 (N2898, N2895, N2150);
or OR4 (N2899, N2872, N1061, N2619, N2651);
nor NOR3 (N2900, N2890, N2377, N1397);
or OR3 (N2901, N2897, N1151, N2775);
xor XOR2 (N2902, N2900, N840);
or OR2 (N2903, N2880, N1837);
nand NAND4 (N2904, N2902, N2292, N1098, N1586);
nand NAND2 (N2905, N2903, N978);
and AND4 (N2906, N2892, N665, N2072, N376);
nor NOR3 (N2907, N2886, N1220, N1035);
not NOT1 (N2908, N2906);
nand NAND3 (N2909, N2898, N1698, N2382);
nand NAND4 (N2910, N2896, N1650, N2883, N2516);
or OR4 (N2911, N2905, N148, N129, N307);
buf BUF1 (N2912, N2899);
or OR2 (N2913, N2901, N93);
not NOT1 (N2914, N2910);
xor XOR2 (N2915, N2914, N1537);
not NOT1 (N2916, N2885);
nor NOR2 (N2917, N2912, N1151);
nor NOR4 (N2918, N2904, N1044, N2796, N933);
or OR4 (N2919, N2917, N2155, N1343, N184);
buf BUF1 (N2920, N2919);
or OR3 (N2921, N2915, N2026, N188);
nor NOR4 (N2922, N2913, N1144, N1405, N487);
nor NOR2 (N2923, N2911, N94);
nand NAND4 (N2924, N2909, N1907, N734, N449);
or OR4 (N2925, N2922, N2583, N2132, N2346);
and AND2 (N2926, N2923, N327);
and AND2 (N2927, N2926, N441);
or OR4 (N2928, N2925, N1907, N911, N155);
and AND4 (N2929, N2907, N498, N1463, N1239);
nand NAND2 (N2930, N2928, N19);
buf BUF1 (N2931, N2930);
xor XOR2 (N2932, N2924, N855);
nor NOR4 (N2933, N2908, N315, N733, N107);
not NOT1 (N2934, N2921);
buf BUF1 (N2935, N2934);
or OR2 (N2936, N2931, N877);
xor XOR2 (N2937, N2936, N286);
or OR3 (N2938, N2889, N1218, N2755);
or OR4 (N2939, N2938, N1337, N928, N1563);
or OR4 (N2940, N2933, N2508, N2802, N1555);
xor XOR2 (N2941, N2927, N1400);
nand NAND3 (N2942, N2932, N872, N1707);
xor XOR2 (N2943, N2937, N2485);
and AND3 (N2944, N2920, N1364, N1658);
not NOT1 (N2945, N2941);
and AND2 (N2946, N2929, N716);
xor XOR2 (N2947, N2943, N454);
xor XOR2 (N2948, N2918, N1825);
nand NAND3 (N2949, N2944, N2789, N689);
xor XOR2 (N2950, N2916, N2592);
buf BUF1 (N2951, N2939);
nand NAND4 (N2952, N2945, N1724, N1606, N1378);
or OR2 (N2953, N2946, N1992);
nor NOR4 (N2954, N2953, N2478, N102, N470);
buf BUF1 (N2955, N2942);
xor XOR2 (N2956, N2951, N943);
nand NAND4 (N2957, N2940, N2128, N228, N978);
or OR3 (N2958, N2955, N920, N2740);
nand NAND2 (N2959, N2956, N2689);
and AND3 (N2960, N2948, N1904, N1499);
nor NOR2 (N2961, N2935, N940);
or OR3 (N2962, N2958, N1490, N802);
not NOT1 (N2963, N2962);
nand NAND4 (N2964, N2960, N2517, N55, N2452);
nor NOR3 (N2965, N2964, N2413, N579);
nor NOR4 (N2966, N2952, N2079, N2725, N1167);
nor NOR2 (N2967, N2965, N2628);
xor XOR2 (N2968, N2963, N1924);
nand NAND3 (N2969, N2968, N2952, N8);
not NOT1 (N2970, N2950);
nor NOR4 (N2971, N2949, N1594, N2830, N1684);
nand NAND3 (N2972, N2959, N1089, N847);
and AND2 (N2973, N2971, N382);
xor XOR2 (N2974, N2954, N443);
nor NOR2 (N2975, N2969, N1903);
not NOT1 (N2976, N2957);
buf BUF1 (N2977, N2972);
and AND2 (N2978, N2947, N2071);
xor XOR2 (N2979, N2967, N2669);
nand NAND2 (N2980, N2966, N1252);
xor XOR2 (N2981, N2978, N2963);
nand NAND2 (N2982, N2974, N209);
buf BUF1 (N2983, N2961);
and AND2 (N2984, N2983, N619);
and AND3 (N2985, N2975, N2693, N341);
nand NAND3 (N2986, N2984, N146, N50);
buf BUF1 (N2987, N2986);
xor XOR2 (N2988, N2980, N2557);
nand NAND3 (N2989, N2982, N2306, N1774);
and AND3 (N2990, N2979, N1850, N1991);
and AND3 (N2991, N2987, N1732, N2918);
buf BUF1 (N2992, N2981);
nand NAND4 (N2993, N2970, N1879, N292, N2052);
nor NOR2 (N2994, N2991, N8);
not NOT1 (N2995, N2990);
nand NAND4 (N2996, N2992, N2896, N1537, N1048);
nand NAND4 (N2997, N2988, N1731, N1965, N2509);
xor XOR2 (N2998, N2973, N2329);
and AND2 (N2999, N2998, N1640);
or OR4 (N3000, N2997, N727, N890, N1304);
nand NAND4 (N3001, N3000, N2428, N466, N2527);
nand NAND2 (N3002, N2985, N2596);
and AND2 (N3003, N2994, N1215);
or OR3 (N3004, N2976, N2603, N159);
not NOT1 (N3005, N2999);
nor NOR3 (N3006, N3005, N423, N1106);
and AND2 (N3007, N3002, N1329);
or OR3 (N3008, N3003, N2875, N1747);
not NOT1 (N3009, N3007);
xor XOR2 (N3010, N2996, N1867);
buf BUF1 (N3011, N3009);
or OR4 (N3012, N2989, N2676, N2764, N2417);
xor XOR2 (N3013, N3012, N986);
not NOT1 (N3014, N3006);
and AND3 (N3015, N2995, N2919, N749);
xor XOR2 (N3016, N3013, N2856);
and AND2 (N3017, N3004, N611);
buf BUF1 (N3018, N3015);
and AND4 (N3019, N2993, N2321, N2608, N1668);
not NOT1 (N3020, N3010);
buf BUF1 (N3021, N3008);
nand NAND2 (N3022, N3019, N660);
not NOT1 (N3023, N3020);
nand NAND4 (N3024, N3018, N2534, N1176, N1855);
nand NAND4 (N3025, N3011, N324, N48, N1488);
nor NOR4 (N3026, N3022, N1587, N2999, N838);
not NOT1 (N3027, N3016);
buf BUF1 (N3028, N3023);
nand NAND3 (N3029, N3028, N1299, N924);
or OR2 (N3030, N3027, N1744);
nor NOR4 (N3031, N3017, N2940, N116, N784);
nor NOR4 (N3032, N3001, N1064, N2630, N2457);
nor NOR3 (N3033, N2977, N1745, N2686);
not NOT1 (N3034, N3025);
buf BUF1 (N3035, N3032);
not NOT1 (N3036, N3033);
and AND3 (N3037, N3029, N2490, N2052);
xor XOR2 (N3038, N3035, N838);
not NOT1 (N3039, N3034);
and AND4 (N3040, N3038, N480, N241, N196);
xor XOR2 (N3041, N3024, N713);
not NOT1 (N3042, N3021);
not NOT1 (N3043, N3031);
xor XOR2 (N3044, N3014, N1366);
not NOT1 (N3045, N3043);
not NOT1 (N3046, N3042);
not NOT1 (N3047, N3037);
xor XOR2 (N3048, N3039, N1786);
nand NAND2 (N3049, N3030, N975);
nor NOR3 (N3050, N3046, N570, N506);
or OR3 (N3051, N3048, N2727, N1338);
and AND3 (N3052, N3036, N2299, N1612);
or OR4 (N3053, N3040, N2307, N2683, N2710);
nor NOR4 (N3054, N3050, N733, N1582, N1077);
buf BUF1 (N3055, N3054);
nand NAND4 (N3056, N3041, N649, N1929, N399);
not NOT1 (N3057, N3044);
nand NAND4 (N3058, N3053, N2592, N704, N339);
nand NAND2 (N3059, N3045, N1126);
nor NOR3 (N3060, N3051, N2381, N972);
and AND2 (N3061, N3047, N453);
nand NAND4 (N3062, N3058, N1612, N2868, N2950);
nor NOR2 (N3063, N3052, N1625);
buf BUF1 (N3064, N3059);
or OR3 (N3065, N3057, N1458, N2628);
not NOT1 (N3066, N3064);
xor XOR2 (N3067, N3060, N2185);
and AND2 (N3068, N3062, N1099);
or OR3 (N3069, N3067, N225, N2074);
or OR3 (N3070, N3065, N2193, N739);
xor XOR2 (N3071, N3049, N2489);
nand NAND3 (N3072, N3066, N123, N474);
nand NAND3 (N3073, N3063, N2424, N1268);
and AND2 (N3074, N3061, N2581);
and AND3 (N3075, N3070, N2616, N495);
and AND3 (N3076, N3075, N2492, N3050);
and AND3 (N3077, N3074, N239, N1706);
nor NOR3 (N3078, N3073, N2905, N1620);
nand NAND2 (N3079, N3078, N2129);
nor NOR3 (N3080, N3072, N129, N2599);
buf BUF1 (N3081, N3026);
or OR4 (N3082, N3069, N1262, N683, N1986);
and AND4 (N3083, N3056, N117, N2308, N3053);
xor XOR2 (N3084, N3068, N2617);
and AND2 (N3085, N3084, N2065);
and AND3 (N3086, N3082, N2593, N789);
and AND4 (N3087, N3055, N2874, N1448, N2379);
or OR4 (N3088, N3076, N2761, N3084, N1632);
xor XOR2 (N3089, N3077, N1472);
nor NOR3 (N3090, N3087, N1659, N276);
or OR4 (N3091, N3088, N2797, N602, N335);
or OR3 (N3092, N3090, N870, N282);
or OR2 (N3093, N3080, N1690);
or OR2 (N3094, N3089, N2598);
or OR3 (N3095, N3091, N1357, N867);
or OR3 (N3096, N3085, N2646, N2717);
xor XOR2 (N3097, N3083, N2927);
and AND2 (N3098, N3095, N1853);
nor NOR4 (N3099, N3098, N1765, N1301, N783);
buf BUF1 (N3100, N3092);
not NOT1 (N3101, N3079);
buf BUF1 (N3102, N3100);
and AND4 (N3103, N3093, N1787, N815, N2249);
nand NAND3 (N3104, N3102, N1295, N2478);
nor NOR3 (N3105, N3101, N303, N2031);
or OR2 (N3106, N3099, N1965);
not NOT1 (N3107, N3104);
and AND3 (N3108, N3097, N105, N261);
nand NAND3 (N3109, N3094, N845, N1552);
buf BUF1 (N3110, N3103);
and AND2 (N3111, N3105, N1050);
buf BUF1 (N3112, N3081);
nand NAND3 (N3113, N3086, N86, N236);
nor NOR4 (N3114, N3096, N1454, N1379, N725);
or OR2 (N3115, N3114, N2527);
nor NOR3 (N3116, N3110, N2968, N1552);
not NOT1 (N3117, N3111);
and AND2 (N3118, N3106, N2949);
nand NAND2 (N3119, N3117, N2232);
and AND2 (N3120, N3119, N954);
or OR3 (N3121, N3108, N1039, N2854);
xor XOR2 (N3122, N3116, N1630);
and AND4 (N3123, N3109, N1373, N32, N684);
and AND4 (N3124, N3113, N2901, N271, N328);
not NOT1 (N3125, N3121);
buf BUF1 (N3126, N3125);
nor NOR3 (N3127, N3122, N1818, N1092);
nand NAND3 (N3128, N3115, N2720, N463);
and AND4 (N3129, N3124, N1536, N1016, N1226);
and AND2 (N3130, N3128, N202);
xor XOR2 (N3131, N3118, N2535);
not NOT1 (N3132, N3126);
or OR2 (N3133, N3132, N1029);
and AND2 (N3134, N3112, N1976);
and AND4 (N3135, N3071, N570, N2177, N2985);
or OR3 (N3136, N3129, N1929, N2592);
and AND4 (N3137, N3120, N1071, N1034, N2425);
nor NOR3 (N3138, N3135, N2884, N2147);
xor XOR2 (N3139, N3107, N2056);
buf BUF1 (N3140, N3133);
buf BUF1 (N3141, N3134);
buf BUF1 (N3142, N3138);
nor NOR3 (N3143, N3130, N1452, N539);
and AND4 (N3144, N3131, N107, N167, N2641);
nor NOR3 (N3145, N3127, N1684, N2748);
or OR3 (N3146, N3136, N21, N2300);
not NOT1 (N3147, N3137);
nor NOR4 (N3148, N3123, N887, N1798, N921);
xor XOR2 (N3149, N3139, N843);
and AND3 (N3150, N3140, N276, N1825);
xor XOR2 (N3151, N3148, N584);
not NOT1 (N3152, N3149);
nor NOR3 (N3153, N3143, N1895, N2642);
nand NAND3 (N3154, N3150, N2197, N474);
not NOT1 (N3155, N3151);
and AND3 (N3156, N3146, N2177, N2648);
buf BUF1 (N3157, N3144);
not NOT1 (N3158, N3152);
or OR3 (N3159, N3156, N1920, N826);
xor XOR2 (N3160, N3147, N1994);
nor NOR2 (N3161, N3157, N1829);
xor XOR2 (N3162, N3158, N1036);
nand NAND2 (N3163, N3153, N2310);
or OR4 (N3164, N3162, N2396, N3017, N2503);
nand NAND4 (N3165, N3145, N2963, N3103, N2295);
and AND4 (N3166, N3165, N406, N2042, N636);
not NOT1 (N3167, N3164);
or OR3 (N3168, N3163, N845, N1143);
nor NOR4 (N3169, N3168, N231, N3006, N2113);
nand NAND3 (N3170, N3142, N1198, N737);
or OR3 (N3171, N3141, N1781, N2195);
xor XOR2 (N3172, N3159, N1632);
xor XOR2 (N3173, N3170, N2954);
xor XOR2 (N3174, N3155, N2288);
or OR3 (N3175, N3166, N2193, N604);
or OR3 (N3176, N3175, N2404, N769);
or OR3 (N3177, N3174, N2761, N1522);
or OR4 (N3178, N3161, N2710, N351, N1834);
buf BUF1 (N3179, N3176);
nor NOR2 (N3180, N3160, N2550);
not NOT1 (N3181, N3167);
buf BUF1 (N3182, N3154);
or OR4 (N3183, N3177, N1739, N1994, N338);
not NOT1 (N3184, N3172);
nand NAND3 (N3185, N3178, N586, N1715);
nand NAND4 (N3186, N3180, N281, N2240, N185);
or OR3 (N3187, N3171, N1295, N2800);
buf BUF1 (N3188, N3187);
xor XOR2 (N3189, N3186, N2861);
or OR4 (N3190, N3179, N1869, N2462, N982);
xor XOR2 (N3191, N3185, N2367);
not NOT1 (N3192, N3182);
nor NOR3 (N3193, N3189, N188, N848);
buf BUF1 (N3194, N3191);
not NOT1 (N3195, N3194);
nand NAND4 (N3196, N3193, N791, N531, N2836);
or OR2 (N3197, N3192, N1962);
buf BUF1 (N3198, N3183);
or OR3 (N3199, N3169, N422, N2926);
and AND4 (N3200, N3195, N1909, N2067, N2060);
xor XOR2 (N3201, N3197, N2662);
nand NAND3 (N3202, N3201, N3087, N110);
or OR4 (N3203, N3196, N1608, N2792, N1504);
or OR2 (N3204, N3203, N930);
or OR3 (N3205, N3173, N1319, N1955);
buf BUF1 (N3206, N3205);
and AND2 (N3207, N3188, N2463);
or OR3 (N3208, N3190, N1215, N2404);
xor XOR2 (N3209, N3199, N1814);
buf BUF1 (N3210, N3204);
nor NOR4 (N3211, N3202, N2979, N999, N884);
or OR3 (N3212, N3181, N2230, N3170);
buf BUF1 (N3213, N3212);
and AND3 (N3214, N3184, N1682, N2370);
xor XOR2 (N3215, N3207, N213);
not NOT1 (N3216, N3211);
nand NAND3 (N3217, N3214, N1728, N2507);
xor XOR2 (N3218, N3215, N2719);
buf BUF1 (N3219, N3206);
nand NAND3 (N3220, N3218, N347, N971);
nand NAND3 (N3221, N3219, N2826, N137);
buf BUF1 (N3222, N3209);
not NOT1 (N3223, N3200);
not NOT1 (N3224, N3220);
nor NOR4 (N3225, N3208, N2929, N147, N1589);
nor NOR3 (N3226, N3210, N991, N3225);
nor NOR4 (N3227, N2066, N2790, N1254, N293);
xor XOR2 (N3228, N3227, N1586);
buf BUF1 (N3229, N3217);
nor NOR4 (N3230, N3229, N102, N1542, N1236);
not NOT1 (N3231, N3230);
not NOT1 (N3232, N3222);
not NOT1 (N3233, N3216);
not NOT1 (N3234, N3221);
xor XOR2 (N3235, N3231, N573);
nand NAND4 (N3236, N3232, N30, N2415, N1080);
and AND2 (N3237, N3233, N2482);
and AND4 (N3238, N3224, N2768, N2628, N782);
nand NAND4 (N3239, N3238, N2866, N1476, N1348);
or OR3 (N3240, N3237, N127, N677);
not NOT1 (N3241, N3239);
not NOT1 (N3242, N3228);
nor NOR4 (N3243, N3223, N49, N2906, N1921);
nor NOR3 (N3244, N3234, N1195, N1324);
nor NOR4 (N3245, N3244, N1327, N1545, N728);
nor NOR4 (N3246, N3240, N2115, N1402, N1224);
nor NOR4 (N3247, N3241, N2407, N2351, N1401);
not NOT1 (N3248, N3236);
xor XOR2 (N3249, N3247, N2730);
nand NAND2 (N3250, N3242, N2063);
nor NOR4 (N3251, N3198, N2508, N3213, N932);
or OR2 (N3252, N1159, N2884);
nand NAND2 (N3253, N3250, N2861);
nand NAND3 (N3254, N3246, N1436, N136);
nand NAND3 (N3255, N3253, N2039, N2081);
and AND4 (N3256, N3226, N2043, N844, N2959);
not NOT1 (N3257, N3255);
xor XOR2 (N3258, N3249, N2715);
xor XOR2 (N3259, N3254, N1671);
and AND2 (N3260, N3248, N2066);
nor NOR4 (N3261, N3235, N840, N3157, N314);
buf BUF1 (N3262, N3251);
xor XOR2 (N3263, N3262, N611);
xor XOR2 (N3264, N3259, N1325);
nand NAND3 (N3265, N3252, N39, N1226);
not NOT1 (N3266, N3243);
nor NOR3 (N3267, N3245, N693, N1673);
nand NAND3 (N3268, N3267, N2353, N54);
and AND3 (N3269, N3266, N544, N26);
xor XOR2 (N3270, N3256, N1086);
nand NAND4 (N3271, N3258, N2161, N217, N1656);
or OR2 (N3272, N3265, N1513);
buf BUF1 (N3273, N3263);
xor XOR2 (N3274, N3257, N1106);
and AND3 (N3275, N3270, N1238, N2033);
or OR3 (N3276, N3269, N965, N287);
and AND2 (N3277, N3268, N2526);
or OR2 (N3278, N3275, N2824);
xor XOR2 (N3279, N3271, N322);
nor NOR3 (N3280, N3277, N2833, N2012);
buf BUF1 (N3281, N3280);
nand NAND3 (N3282, N3273, N2253, N1969);
not NOT1 (N3283, N3260);
buf BUF1 (N3284, N3283);
buf BUF1 (N3285, N3284);
and AND4 (N3286, N3272, N3170, N1571, N2673);
xor XOR2 (N3287, N3279, N2029);
nand NAND2 (N3288, N3281, N2746);
not NOT1 (N3289, N3264);
nand NAND2 (N3290, N3285, N2913);
xor XOR2 (N3291, N3286, N267);
and AND2 (N3292, N3290, N486);
or OR2 (N3293, N3278, N2566);
nor NOR4 (N3294, N3276, N2760, N849, N2218);
xor XOR2 (N3295, N3293, N1639);
nand NAND3 (N3296, N3291, N1110, N2349);
buf BUF1 (N3297, N3294);
nor NOR3 (N3298, N3295, N1201, N1471);
xor XOR2 (N3299, N3274, N1963);
buf BUF1 (N3300, N3287);
or OR3 (N3301, N3288, N660, N2679);
and AND4 (N3302, N3282, N3169, N2361, N1507);
nor NOR3 (N3303, N3301, N583, N413);
nand NAND3 (N3304, N3300, N3206, N554);
xor XOR2 (N3305, N3299, N2390);
nand NAND3 (N3306, N3292, N3293, N3129);
and AND3 (N3307, N3305, N442, N2900);
nand NAND2 (N3308, N3298, N486);
nand NAND2 (N3309, N3297, N752);
not NOT1 (N3310, N3307);
not NOT1 (N3311, N3302);
buf BUF1 (N3312, N3289);
xor XOR2 (N3313, N3303, N2953);
nor NOR4 (N3314, N3304, N2476, N1659, N601);
not NOT1 (N3315, N3309);
nor NOR3 (N3316, N3315, N542, N2528);
nand NAND3 (N3317, N3313, N1949, N2318);
and AND4 (N3318, N3261, N762, N14, N1922);
not NOT1 (N3319, N3296);
and AND4 (N3320, N3316, N876, N539, N2705);
nor NOR4 (N3321, N3312, N517, N2629, N529);
and AND4 (N3322, N3320, N2590, N144, N2907);
xor XOR2 (N3323, N3311, N2927);
and AND3 (N3324, N3308, N1017, N3181);
xor XOR2 (N3325, N3306, N1392);
nor NOR2 (N3326, N3321, N2662);
or OR2 (N3327, N3318, N238);
nor NOR4 (N3328, N3325, N1480, N1241, N2238);
xor XOR2 (N3329, N3326, N2397);
or OR4 (N3330, N3314, N111, N814, N58);
nand NAND3 (N3331, N3322, N1491, N1986);
buf BUF1 (N3332, N3324);
or OR2 (N3333, N3317, N2228);
and AND4 (N3334, N3323, N2143, N3076, N1138);
or OR4 (N3335, N3329, N520, N469, N260);
nand NAND4 (N3336, N3310, N1491, N328, N1287);
and AND3 (N3337, N3332, N1767, N902);
xor XOR2 (N3338, N3333, N653);
buf BUF1 (N3339, N3331);
buf BUF1 (N3340, N3330);
buf BUF1 (N3341, N3334);
buf BUF1 (N3342, N3335);
and AND2 (N3343, N3341, N1538);
not NOT1 (N3344, N3336);
and AND3 (N3345, N3319, N2006, N2428);
or OR2 (N3346, N3327, N546);
and AND4 (N3347, N3344, N3251, N1892, N2335);
nor NOR4 (N3348, N3328, N1087, N1705, N942);
xor XOR2 (N3349, N3348, N2246);
not NOT1 (N3350, N3342);
and AND2 (N3351, N3337, N2821);
and AND3 (N3352, N3351, N1836, N1348);
not NOT1 (N3353, N3343);
buf BUF1 (N3354, N3349);
or OR3 (N3355, N3347, N677, N446);
xor XOR2 (N3356, N3353, N1858);
or OR4 (N3357, N3345, N1351, N2068, N507);
nor NOR2 (N3358, N3338, N1534);
xor XOR2 (N3359, N3358, N3098);
or OR3 (N3360, N3340, N1718, N1484);
nor NOR2 (N3361, N3360, N654);
nor NOR2 (N3362, N3361, N2519);
or OR2 (N3363, N3356, N194);
or OR3 (N3364, N3355, N3144, N2476);
or OR4 (N3365, N3350, N128, N1226, N2165);
nand NAND2 (N3366, N3352, N1025);
nand NAND2 (N3367, N3366, N546);
xor XOR2 (N3368, N3365, N3107);
buf BUF1 (N3369, N3346);
nor NOR4 (N3370, N3362, N2529, N475, N553);
and AND4 (N3371, N3363, N86, N2338, N974);
xor XOR2 (N3372, N3357, N1423);
xor XOR2 (N3373, N3368, N216);
and AND2 (N3374, N3367, N2061);
or OR4 (N3375, N3364, N3292, N3176, N2431);
nand NAND3 (N3376, N3359, N2803, N1564);
and AND3 (N3377, N3376, N363, N1173);
xor XOR2 (N3378, N3372, N414);
not NOT1 (N3379, N3377);
and AND2 (N3380, N3379, N239);
not NOT1 (N3381, N3369);
nand NAND3 (N3382, N3371, N464, N2897);
or OR3 (N3383, N3373, N1075, N2077);
nor NOR4 (N3384, N3383, N3141, N1391, N1280);
or OR2 (N3385, N3354, N2075);
xor XOR2 (N3386, N3382, N3296);
and AND4 (N3387, N3370, N2824, N1439, N2843);
not NOT1 (N3388, N3381);
and AND3 (N3389, N3387, N2878, N229);
buf BUF1 (N3390, N3385);
and AND3 (N3391, N3339, N648, N1044);
nand NAND4 (N3392, N3389, N1204, N842, N1262);
nor NOR3 (N3393, N3374, N1343, N1316);
xor XOR2 (N3394, N3392, N1353);
buf BUF1 (N3395, N3384);
not NOT1 (N3396, N3394);
nor NOR3 (N3397, N3393, N2316, N1854);
and AND3 (N3398, N3380, N3147, N1436);
nand NAND3 (N3399, N3398, N2905, N2504);
not NOT1 (N3400, N3397);
nand NAND3 (N3401, N3375, N2529, N3390);
nand NAND3 (N3402, N3218, N1404, N1110);
not NOT1 (N3403, N3402);
not NOT1 (N3404, N3388);
or OR4 (N3405, N3391, N2844, N758, N3347);
and AND4 (N3406, N3403, N758, N837, N2879);
nor NOR2 (N3407, N3401, N215);
buf BUF1 (N3408, N3399);
buf BUF1 (N3409, N3408);
nand NAND2 (N3410, N3378, N189);
nand NAND4 (N3411, N3405, N555, N1872, N3235);
nor NOR2 (N3412, N3407, N810);
nor NOR2 (N3413, N3412, N1084);
or OR3 (N3414, N3411, N1415, N440);
nand NAND2 (N3415, N3413, N2769);
and AND2 (N3416, N3409, N772);
and AND2 (N3417, N3400, N1961);
buf BUF1 (N3418, N3410);
nand NAND4 (N3419, N3414, N3312, N2960, N1367);
nand NAND4 (N3420, N3404, N3295, N1495, N2832);
and AND3 (N3421, N3417, N1660, N3303);
not NOT1 (N3422, N3420);
nor NOR3 (N3423, N3421, N169, N2826);
nand NAND2 (N3424, N3395, N145);
nor NOR3 (N3425, N3419, N2919, N986);
nand NAND2 (N3426, N3424, N571);
buf BUF1 (N3427, N3425);
nor NOR2 (N3428, N3427, N2437);
nand NAND3 (N3429, N3406, N2908, N2200);
not NOT1 (N3430, N3416);
and AND3 (N3431, N3418, N1063, N2813);
nand NAND3 (N3432, N3396, N2917, N1645);
and AND3 (N3433, N3422, N1093, N979);
nand NAND2 (N3434, N3433, N2199);
or OR4 (N3435, N3434, N1043, N3364, N2081);
or OR4 (N3436, N3415, N1185, N1501, N2197);
xor XOR2 (N3437, N3430, N2570);
xor XOR2 (N3438, N3437, N299);
nor NOR4 (N3439, N3431, N1653, N1027, N1444);
nor NOR4 (N3440, N3438, N2858, N2383, N1626);
buf BUF1 (N3441, N3440);
or OR2 (N3442, N3426, N2068);
nor NOR4 (N3443, N3439, N2349, N3436, N2425);
or OR2 (N3444, N1996, N525);
and AND2 (N3445, N3428, N551);
and AND3 (N3446, N3442, N3171, N2256);
xor XOR2 (N3447, N3432, N3197);
xor XOR2 (N3448, N3441, N2753);
buf BUF1 (N3449, N3423);
and AND3 (N3450, N3386, N1830, N447);
nor NOR3 (N3451, N3444, N735, N1881);
not NOT1 (N3452, N3448);
nor NOR3 (N3453, N3435, N43, N209);
buf BUF1 (N3454, N3449);
nor NOR2 (N3455, N3447, N1064);
or OR2 (N3456, N3454, N71);
nand NAND3 (N3457, N3456, N2268, N2040);
nand NAND2 (N3458, N3429, N2522);
nor NOR3 (N3459, N3443, N2926, N131);
not NOT1 (N3460, N3450);
nand NAND4 (N3461, N3460, N491, N1973, N450);
buf BUF1 (N3462, N3457);
not NOT1 (N3463, N3462);
buf BUF1 (N3464, N3455);
and AND4 (N3465, N3452, N1338, N1051, N1570);
and AND3 (N3466, N3463, N2989, N1688);
nand NAND4 (N3467, N3445, N2578, N2459, N1102);
buf BUF1 (N3468, N3459);
nand NAND2 (N3469, N3446, N3199);
or OR3 (N3470, N3468, N2472, N2682);
not NOT1 (N3471, N3461);
nand NAND3 (N3472, N3465, N2278, N1594);
and AND3 (N3473, N3467, N1621, N1106);
nand NAND3 (N3474, N3473, N2354, N470);
or OR3 (N3475, N3464, N2318, N1733);
not NOT1 (N3476, N3474);
nor NOR3 (N3477, N3476, N950, N404);
buf BUF1 (N3478, N3477);
not NOT1 (N3479, N3458);
not NOT1 (N3480, N3475);
not NOT1 (N3481, N3480);
nand NAND3 (N3482, N3469, N2512, N1165);
nand NAND4 (N3483, N3466, N876, N1370, N57);
buf BUF1 (N3484, N3479);
not NOT1 (N3485, N3482);
or OR2 (N3486, N3485, N689);
and AND3 (N3487, N3478, N2229, N2243);
and AND4 (N3488, N3453, N2668, N3324, N1064);
or OR3 (N3489, N3487, N3134, N2564);
xor XOR2 (N3490, N3484, N1031);
buf BUF1 (N3491, N3486);
buf BUF1 (N3492, N3490);
and AND3 (N3493, N3471, N509, N961);
buf BUF1 (N3494, N3488);
not NOT1 (N3495, N3492);
and AND3 (N3496, N3491, N1058, N2576);
or OR3 (N3497, N3489, N2087, N2825);
nand NAND4 (N3498, N3493, N2621, N2001, N906);
xor XOR2 (N3499, N3472, N2123);
xor XOR2 (N3500, N3481, N2457);
or OR4 (N3501, N3470, N3022, N685, N2469);
nor NOR2 (N3502, N3483, N3154);
xor XOR2 (N3503, N3502, N1128);
not NOT1 (N3504, N3496);
and AND2 (N3505, N3495, N2374);
and AND4 (N3506, N3494, N1137, N1071, N3420);
buf BUF1 (N3507, N3499);
nand NAND3 (N3508, N3504, N119, N699);
and AND2 (N3509, N3506, N791);
buf BUF1 (N3510, N3503);
or OR3 (N3511, N3507, N2462, N2508);
nor NOR3 (N3512, N3508, N2528, N1908);
or OR2 (N3513, N3501, N732);
xor XOR2 (N3514, N3510, N3080);
and AND2 (N3515, N3451, N2338);
nand NAND3 (N3516, N3505, N472, N3138);
nor NOR3 (N3517, N3497, N3024, N2049);
buf BUF1 (N3518, N3512);
nor NOR3 (N3519, N3516, N3244, N1461);
nand NAND2 (N3520, N3500, N1790);
nor NOR3 (N3521, N3514, N2541, N2193);
endmodule