// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N4007,N4010,N4012,N4011,N4005,N4009,N4015,N4006,N4008,N4016;

nand NAND4 (N17, N15, N13, N3, N6);
not NOT1 (N18, N15);
nand NAND2 (N19, N3, N1);
buf BUF1 (N20, N18);
nand NAND4 (N21, N20, N13, N16, N1);
buf BUF1 (N22, N4);
nand NAND4 (N23, N4, N18, N18, N2);
nor NOR3 (N24, N5, N1, N22);
nand NAND2 (N25, N14, N11);
buf BUF1 (N26, N1);
buf BUF1 (N27, N1);
nor NOR3 (N28, N14, N1, N25);
nor NOR3 (N29, N3, N22, N4);
or OR3 (N30, N21, N25, N10);
or OR3 (N31, N2, N20, N14);
not NOT1 (N32, N26);
or OR2 (N33, N23, N30);
nand NAND2 (N34, N29, N22);
not NOT1 (N35, N13);
or OR2 (N36, N27, N7);
xor XOR2 (N37, N32, N8);
buf BUF1 (N38, N24);
and AND4 (N39, N34, N33, N20, N26);
buf BUF1 (N40, N17);
not NOT1 (N41, N33);
nand NAND2 (N42, N19, N30);
xor XOR2 (N43, N41, N1);
nor NOR2 (N44, N31, N5);
xor XOR2 (N45, N39, N21);
buf BUF1 (N46, N36);
xor XOR2 (N47, N40, N28);
or OR2 (N48, N26, N28);
buf BUF1 (N49, N45);
nor NOR2 (N50, N37, N20);
or OR2 (N51, N49, N44);
nor NOR2 (N52, N11, N12);
nor NOR3 (N53, N47, N45, N17);
xor XOR2 (N54, N52, N48);
or OR4 (N55, N23, N22, N6, N1);
not NOT1 (N56, N51);
and AND2 (N57, N50, N55);
xor XOR2 (N58, N25, N42);
buf BUF1 (N59, N40);
and AND4 (N60, N58, N37, N6, N4);
nand NAND4 (N61, N53, N17, N29, N13);
and AND4 (N62, N46, N39, N31, N44);
xor XOR2 (N63, N54, N14);
xor XOR2 (N64, N43, N35);
xor XOR2 (N65, N1, N26);
xor XOR2 (N66, N62, N56);
and AND2 (N67, N28, N11);
nand NAND2 (N68, N57, N34);
buf BUF1 (N69, N67);
not NOT1 (N70, N38);
xor XOR2 (N71, N64, N43);
nand NAND4 (N72, N68, N56, N28, N30);
or OR2 (N73, N72, N62);
nand NAND4 (N74, N71, N68, N19, N44);
xor XOR2 (N75, N60, N41);
nand NAND4 (N76, N61, N14, N24, N25);
nor NOR4 (N77, N66, N75, N2, N63);
buf BUF1 (N78, N7);
or OR3 (N79, N42, N68, N75);
xor XOR2 (N80, N76, N72);
or OR2 (N81, N80, N31);
nand NAND2 (N82, N81, N68);
nand NAND3 (N83, N65, N9, N22);
and AND3 (N84, N73, N71, N12);
or OR4 (N85, N82, N28, N9, N20);
not NOT1 (N86, N78);
or OR3 (N87, N86, N35, N17);
nor NOR4 (N88, N70, N51, N61, N36);
nand NAND4 (N89, N84, N41, N26, N21);
xor XOR2 (N90, N59, N15);
xor XOR2 (N91, N74, N13);
not NOT1 (N92, N85);
nor NOR2 (N93, N91, N24);
buf BUF1 (N94, N89);
and AND2 (N95, N88, N13);
xor XOR2 (N96, N79, N35);
or OR4 (N97, N90, N32, N27, N44);
nor NOR2 (N98, N96, N70);
nand NAND2 (N99, N93, N94);
nor NOR3 (N100, N70, N10, N99);
nor NOR3 (N101, N84, N61, N32);
and AND2 (N102, N87, N73);
xor XOR2 (N103, N102, N11);
nor NOR2 (N104, N77, N92);
buf BUF1 (N105, N68);
xor XOR2 (N106, N83, N48);
buf BUF1 (N107, N105);
buf BUF1 (N108, N69);
and AND4 (N109, N100, N54, N27, N8);
buf BUF1 (N110, N103);
nor NOR2 (N111, N101, N99);
nand NAND3 (N112, N97, N82, N7);
nand NAND4 (N113, N109, N57, N28, N2);
buf BUF1 (N114, N98);
xor XOR2 (N115, N111, N3);
not NOT1 (N116, N108);
and AND4 (N117, N107, N46, N29, N43);
xor XOR2 (N118, N95, N24);
not NOT1 (N119, N113);
nor NOR2 (N120, N115, N102);
or OR4 (N121, N117, N62, N120, N73);
xor XOR2 (N122, N3, N109);
nand NAND2 (N123, N110, N71);
xor XOR2 (N124, N114, N122);
nor NOR4 (N125, N49, N34, N66, N31);
buf BUF1 (N126, N104);
buf BUF1 (N127, N125);
nand NAND2 (N128, N112, N40);
and AND4 (N129, N121, N107, N6, N11);
not NOT1 (N130, N126);
xor XOR2 (N131, N127, N53);
nand NAND3 (N132, N106, N115, N16);
xor XOR2 (N133, N128, N44);
and AND3 (N134, N119, N118, N27);
not NOT1 (N135, N52);
and AND3 (N136, N124, N17, N4);
and AND2 (N137, N129, N125);
or OR4 (N138, N136, N119, N75, N8);
and AND2 (N139, N134, N132);
and AND4 (N140, N117, N85, N48, N40);
nor NOR2 (N141, N137, N137);
and AND4 (N142, N138, N67, N41, N91);
or OR4 (N143, N131, N7, N15, N70);
nor NOR3 (N144, N140, N81, N91);
not NOT1 (N145, N130);
buf BUF1 (N146, N135);
or OR2 (N147, N116, N123);
buf BUF1 (N148, N125);
nand NAND3 (N149, N139, N103, N107);
and AND3 (N150, N133, N29, N17);
nor NOR2 (N151, N146, N21);
xor XOR2 (N152, N150, N133);
nand NAND3 (N153, N144, N1, N23);
buf BUF1 (N154, N148);
not NOT1 (N155, N143);
and AND3 (N156, N154, N28, N40);
not NOT1 (N157, N156);
nor NOR3 (N158, N157, N111, N56);
and AND2 (N159, N147, N124);
buf BUF1 (N160, N155);
nand NAND3 (N161, N152, N95, N69);
buf BUF1 (N162, N158);
nand NAND4 (N163, N145, N33, N67, N121);
buf BUF1 (N164, N159);
not NOT1 (N165, N141);
xor XOR2 (N166, N164, N47);
not NOT1 (N167, N149);
or OR2 (N168, N167, N92);
or OR2 (N169, N166, N46);
or OR3 (N170, N160, N141, N27);
or OR2 (N171, N153, N147);
xor XOR2 (N172, N170, N98);
buf BUF1 (N173, N172);
nand NAND2 (N174, N162, N29);
not NOT1 (N175, N173);
buf BUF1 (N176, N165);
nor NOR2 (N177, N169, N143);
or OR4 (N178, N171, N140, N16, N162);
nor NOR4 (N179, N174, N4, N165, N34);
not NOT1 (N180, N178);
not NOT1 (N181, N177);
nor NOR4 (N182, N180, N176, N49, N124);
and AND4 (N183, N36, N4, N78, N27);
and AND4 (N184, N168, N177, N100, N19);
xor XOR2 (N185, N161, N56);
and AND4 (N186, N185, N23, N97, N155);
not NOT1 (N187, N179);
nor NOR3 (N188, N184, N79, N57);
nand NAND4 (N189, N182, N12, N8, N94);
or OR2 (N190, N189, N126);
or OR4 (N191, N181, N55, N87, N167);
or OR3 (N192, N175, N128, N8);
not NOT1 (N193, N188);
not NOT1 (N194, N183);
nand NAND4 (N195, N194, N181, N75, N138);
xor XOR2 (N196, N186, N100);
and AND3 (N197, N142, N95, N43);
nand NAND4 (N198, N195, N56, N132, N185);
and AND3 (N199, N190, N95, N64);
not NOT1 (N200, N187);
xor XOR2 (N201, N191, N100);
nand NAND3 (N202, N163, N116, N145);
and AND3 (N203, N198, N200, N76);
and AND2 (N204, N22, N77);
or OR2 (N205, N201, N150);
buf BUF1 (N206, N205);
xor XOR2 (N207, N193, N85);
buf BUF1 (N208, N151);
or OR3 (N209, N203, N145, N101);
xor XOR2 (N210, N209, N117);
nand NAND2 (N211, N207, N52);
xor XOR2 (N212, N197, N182);
and AND2 (N213, N210, N89);
buf BUF1 (N214, N212);
nor NOR4 (N215, N196, N5, N126, N49);
buf BUF1 (N216, N202);
and AND3 (N217, N204, N78, N176);
not NOT1 (N218, N211);
xor XOR2 (N219, N192, N7);
nor NOR2 (N220, N208, N169);
or OR2 (N221, N218, N33);
nor NOR4 (N222, N206, N190, N221, N203);
buf BUF1 (N223, N148);
nand NAND3 (N224, N219, N165, N69);
not NOT1 (N225, N214);
nand NAND3 (N226, N223, N153, N97);
not NOT1 (N227, N217);
nand NAND3 (N228, N215, N145, N73);
nand NAND2 (N229, N222, N69);
nand NAND4 (N230, N228, N84, N63, N18);
not NOT1 (N231, N199);
and AND4 (N232, N226, N10, N150, N166);
xor XOR2 (N233, N220, N218);
buf BUF1 (N234, N231);
or OR3 (N235, N225, N72, N210);
nor NOR2 (N236, N235, N221);
nor NOR2 (N237, N213, N172);
or OR3 (N238, N234, N229, N218);
or OR4 (N239, N30, N51, N135, N130);
xor XOR2 (N240, N232, N4);
buf BUF1 (N241, N230);
or OR3 (N242, N236, N163, N125);
nand NAND3 (N243, N216, N199, N193);
not NOT1 (N244, N238);
xor XOR2 (N245, N233, N45);
nor NOR4 (N246, N244, N57, N184, N232);
not NOT1 (N247, N224);
not NOT1 (N248, N239);
nor NOR4 (N249, N242, N135, N132, N182);
buf BUF1 (N250, N247);
nand NAND3 (N251, N248, N187, N200);
not NOT1 (N252, N249);
and AND3 (N253, N245, N222, N215);
xor XOR2 (N254, N227, N231);
not NOT1 (N255, N246);
buf BUF1 (N256, N255);
xor XOR2 (N257, N240, N102);
and AND4 (N258, N237, N250, N98, N54);
or OR2 (N259, N168, N244);
buf BUF1 (N260, N254);
nand NAND2 (N261, N252, N166);
and AND3 (N262, N241, N180, N131);
or OR2 (N263, N259, N20);
buf BUF1 (N264, N262);
xor XOR2 (N265, N257, N238);
or OR2 (N266, N256, N55);
nor NOR3 (N267, N265, N192, N243);
nor NOR3 (N268, N219, N176, N177);
and AND3 (N269, N268, N47, N33);
xor XOR2 (N270, N253, N239);
or OR3 (N271, N269, N176, N198);
not NOT1 (N272, N266);
xor XOR2 (N273, N263, N10);
or OR3 (N274, N258, N33, N205);
or OR4 (N275, N270, N27, N87, N44);
xor XOR2 (N276, N260, N197);
not NOT1 (N277, N251);
xor XOR2 (N278, N264, N269);
or OR4 (N279, N272, N182, N195, N98);
and AND4 (N280, N277, N117, N42, N133);
buf BUF1 (N281, N278);
not NOT1 (N282, N276);
not NOT1 (N283, N274);
nor NOR2 (N284, N279, N282);
xor XOR2 (N285, N187, N149);
buf BUF1 (N286, N271);
nand NAND3 (N287, N281, N52, N59);
and AND4 (N288, N284, N21, N14, N95);
buf BUF1 (N289, N285);
nor NOR2 (N290, N280, N139);
xor XOR2 (N291, N261, N168);
buf BUF1 (N292, N286);
not NOT1 (N293, N288);
nand NAND2 (N294, N289, N56);
nor NOR2 (N295, N291, N44);
nand NAND2 (N296, N290, N159);
nand NAND2 (N297, N293, N249);
and AND2 (N298, N287, N27);
not NOT1 (N299, N297);
nand NAND3 (N300, N299, N23, N221);
nor NOR2 (N301, N296, N70);
not NOT1 (N302, N295);
buf BUF1 (N303, N294);
xor XOR2 (N304, N267, N113);
buf BUF1 (N305, N298);
buf BUF1 (N306, N303);
not NOT1 (N307, N302);
and AND4 (N308, N301, N270, N17, N91);
xor XOR2 (N309, N292, N110);
nor NOR3 (N310, N273, N36, N200);
nand NAND3 (N311, N305, N185, N147);
and AND4 (N312, N309, N7, N230, N143);
nor NOR2 (N313, N306, N148);
nand NAND3 (N314, N310, N193, N303);
and AND4 (N315, N311, N53, N155, N260);
not NOT1 (N316, N300);
buf BUF1 (N317, N308);
xor XOR2 (N318, N316, N81);
not NOT1 (N319, N283);
or OR2 (N320, N312, N122);
or OR3 (N321, N315, N59, N300);
buf BUF1 (N322, N321);
or OR3 (N323, N314, N209, N174);
not NOT1 (N324, N320);
not NOT1 (N325, N324);
or OR3 (N326, N325, N205, N294);
and AND2 (N327, N323, N56);
not NOT1 (N328, N313);
not NOT1 (N329, N327);
xor XOR2 (N330, N322, N183);
nand NAND4 (N331, N329, N110, N29, N57);
buf BUF1 (N332, N318);
nand NAND4 (N333, N304, N36, N116, N246);
and AND4 (N334, N326, N186, N98, N90);
nand NAND4 (N335, N328, N93, N79, N27);
and AND2 (N336, N333, N202);
or OR2 (N337, N335, N266);
and AND4 (N338, N336, N313, N121, N209);
nand NAND4 (N339, N331, N50, N157, N66);
not NOT1 (N340, N334);
not NOT1 (N341, N275);
nor NOR2 (N342, N341, N334);
not NOT1 (N343, N307);
or OR2 (N344, N342, N146);
buf BUF1 (N345, N317);
nor NOR2 (N346, N343, N173);
nand NAND3 (N347, N340, N147, N34);
not NOT1 (N348, N345);
or OR2 (N349, N344, N261);
and AND4 (N350, N319, N229, N266, N144);
xor XOR2 (N351, N350, N105);
buf BUF1 (N352, N349);
buf BUF1 (N353, N351);
buf BUF1 (N354, N339);
or OR2 (N355, N352, N242);
nor NOR4 (N356, N353, N169, N5, N29);
or OR4 (N357, N330, N118, N261, N154);
or OR3 (N358, N356, N263, N324);
nor NOR4 (N359, N348, N203, N339, N228);
nand NAND3 (N360, N354, N241, N175);
and AND3 (N361, N359, N302, N49);
and AND2 (N362, N360, N247);
not NOT1 (N363, N358);
xor XOR2 (N364, N363, N16);
and AND2 (N365, N364, N270);
buf BUF1 (N366, N361);
nand NAND2 (N367, N337, N144);
and AND3 (N368, N346, N4, N180);
or OR3 (N369, N338, N30, N242);
and AND3 (N370, N365, N195, N62);
or OR2 (N371, N367, N237);
or OR3 (N372, N371, N58, N218);
xor XOR2 (N373, N370, N132);
buf BUF1 (N374, N372);
or OR2 (N375, N368, N137);
or OR4 (N376, N362, N286, N363, N283);
buf BUF1 (N377, N376);
or OR2 (N378, N332, N108);
nand NAND2 (N379, N373, N246);
and AND2 (N380, N369, N292);
buf BUF1 (N381, N378);
nor NOR2 (N382, N380, N23);
not NOT1 (N383, N355);
xor XOR2 (N384, N382, N138);
and AND4 (N385, N377, N58, N206, N60);
xor XOR2 (N386, N366, N101);
buf BUF1 (N387, N379);
buf BUF1 (N388, N381);
nand NAND4 (N389, N375, N113, N325, N111);
and AND4 (N390, N387, N155, N69, N341);
buf BUF1 (N391, N385);
or OR4 (N392, N386, N197, N156, N151);
and AND3 (N393, N347, N304, N240);
buf BUF1 (N394, N392);
or OR2 (N395, N374, N234);
not NOT1 (N396, N384);
xor XOR2 (N397, N394, N163);
and AND3 (N398, N395, N202, N186);
and AND4 (N399, N391, N46, N50, N134);
nand NAND4 (N400, N396, N346, N16, N312);
not NOT1 (N401, N388);
not NOT1 (N402, N400);
xor XOR2 (N403, N401, N383);
nand NAND4 (N404, N71, N330, N325, N86);
not NOT1 (N405, N357);
or OR3 (N406, N403, N9, N215);
nor NOR4 (N407, N399, N178, N112, N146);
or OR3 (N408, N397, N177, N284);
or OR4 (N409, N406, N371, N47, N125);
nand NAND4 (N410, N408, N226, N250, N382);
nand NAND3 (N411, N390, N24, N52);
and AND2 (N412, N410, N186);
xor XOR2 (N413, N411, N255);
not NOT1 (N414, N398);
and AND2 (N415, N393, N105);
buf BUF1 (N416, N409);
nor NOR4 (N417, N407, N150, N6, N403);
xor XOR2 (N418, N415, N360);
xor XOR2 (N419, N413, N59);
nor NOR4 (N420, N416, N360, N234, N303);
nor NOR4 (N421, N389, N112, N277, N173);
or OR4 (N422, N420, N261, N312, N39);
nand NAND4 (N423, N404, N289, N209, N119);
or OR2 (N424, N414, N402);
buf BUF1 (N425, N208);
nor NOR4 (N426, N417, N270, N416, N110);
nor NOR2 (N427, N422, N415);
nor NOR4 (N428, N424, N344, N224, N269);
nor NOR3 (N429, N418, N137, N205);
not NOT1 (N430, N425);
and AND3 (N431, N427, N264, N387);
or OR4 (N432, N430, N5, N173, N125);
buf BUF1 (N433, N421);
not NOT1 (N434, N405);
nor NOR2 (N435, N426, N110);
and AND4 (N436, N419, N73, N149, N269);
nand NAND4 (N437, N431, N35, N116, N269);
xor XOR2 (N438, N436, N437);
not NOT1 (N439, N247);
nor NOR3 (N440, N432, N206, N345);
not NOT1 (N441, N438);
xor XOR2 (N442, N441, N138);
buf BUF1 (N443, N442);
and AND4 (N444, N429, N375, N419, N363);
and AND2 (N445, N412, N248);
and AND2 (N446, N443, N35);
not NOT1 (N447, N446);
xor XOR2 (N448, N434, N210);
not NOT1 (N449, N440);
not NOT1 (N450, N444);
buf BUF1 (N451, N450);
xor XOR2 (N452, N447, N37);
and AND2 (N453, N451, N340);
not NOT1 (N454, N428);
xor XOR2 (N455, N439, N108);
nor NOR2 (N456, N433, N299);
nor NOR4 (N457, N454, N138, N195, N390);
or OR2 (N458, N449, N388);
nor NOR2 (N459, N453, N79);
or OR2 (N460, N458, N387);
and AND3 (N461, N452, N409, N99);
or OR4 (N462, N448, N333, N58, N53);
and AND3 (N463, N461, N309, N368);
nand NAND2 (N464, N457, N112);
nand NAND2 (N465, N460, N335);
xor XOR2 (N466, N459, N9);
and AND3 (N467, N455, N147, N159);
and AND3 (N468, N462, N246, N236);
nand NAND3 (N469, N464, N454, N233);
nor NOR4 (N470, N463, N98, N426, N423);
xor XOR2 (N471, N382, N199);
xor XOR2 (N472, N445, N78);
not NOT1 (N473, N470);
or OR4 (N474, N435, N366, N448, N94);
not NOT1 (N475, N474);
xor XOR2 (N476, N456, N196);
buf BUF1 (N477, N472);
or OR2 (N478, N469, N236);
nand NAND3 (N479, N477, N380, N142);
and AND3 (N480, N468, N275, N290);
buf BUF1 (N481, N478);
nand NAND2 (N482, N465, N47);
or OR3 (N483, N480, N260, N236);
or OR3 (N484, N475, N274, N39);
buf BUF1 (N485, N467);
buf BUF1 (N486, N473);
xor XOR2 (N487, N479, N136);
not NOT1 (N488, N481);
and AND2 (N489, N483, N132);
xor XOR2 (N490, N485, N197);
nand NAND2 (N491, N476, N172);
nor NOR2 (N492, N486, N107);
not NOT1 (N493, N492);
not NOT1 (N494, N466);
xor XOR2 (N495, N491, N67);
nand NAND4 (N496, N487, N317, N410, N340);
nand NAND4 (N497, N494, N269, N486, N299);
nor NOR2 (N498, N497, N239);
not NOT1 (N499, N484);
nand NAND2 (N500, N482, N287);
not NOT1 (N501, N496);
buf BUF1 (N502, N500);
not NOT1 (N503, N493);
nor NOR2 (N504, N501, N181);
nor NOR2 (N505, N499, N208);
nor NOR2 (N506, N504, N152);
xor XOR2 (N507, N506, N315);
nand NAND2 (N508, N488, N55);
nand NAND4 (N509, N508, N424, N139, N410);
or OR2 (N510, N490, N342);
or OR2 (N511, N510, N57);
nand NAND4 (N512, N495, N175, N162, N323);
or OR2 (N513, N498, N128);
or OR2 (N514, N503, N32);
buf BUF1 (N515, N489);
xor XOR2 (N516, N511, N439);
or OR3 (N517, N515, N272, N239);
nor NOR3 (N518, N516, N285, N291);
xor XOR2 (N519, N513, N331);
or OR4 (N520, N502, N124, N394, N501);
buf BUF1 (N521, N520);
or OR2 (N522, N509, N213);
and AND2 (N523, N505, N168);
nor NOR4 (N524, N522, N355, N511, N70);
nand NAND2 (N525, N521, N79);
and AND4 (N526, N471, N213, N405, N102);
buf BUF1 (N527, N517);
nand NAND3 (N528, N525, N456, N213);
and AND3 (N529, N526, N50, N266);
xor XOR2 (N530, N512, N172);
xor XOR2 (N531, N524, N115);
nand NAND2 (N532, N507, N197);
nand NAND4 (N533, N527, N308, N131, N135);
or OR4 (N534, N518, N95, N274, N3);
buf BUF1 (N535, N523);
nand NAND3 (N536, N514, N22, N247);
not NOT1 (N537, N532);
xor XOR2 (N538, N535, N362);
xor XOR2 (N539, N534, N439);
or OR4 (N540, N528, N419, N223, N164);
buf BUF1 (N541, N529);
nor NOR2 (N542, N541, N161);
not NOT1 (N543, N533);
not NOT1 (N544, N539);
not NOT1 (N545, N538);
xor XOR2 (N546, N545, N515);
nor NOR2 (N547, N540, N454);
xor XOR2 (N548, N531, N184);
and AND2 (N549, N548, N340);
xor XOR2 (N550, N544, N123);
xor XOR2 (N551, N543, N41);
buf BUF1 (N552, N550);
nand NAND3 (N553, N546, N295, N309);
not NOT1 (N554, N537);
nand NAND4 (N555, N519, N490, N177, N388);
and AND2 (N556, N555, N127);
nand NAND3 (N557, N542, N227, N210);
and AND4 (N558, N547, N142, N550, N98);
buf BUF1 (N559, N530);
nand NAND4 (N560, N536, N507, N49, N169);
nor NOR2 (N561, N551, N308);
nor NOR3 (N562, N558, N433, N127);
not NOT1 (N563, N562);
not NOT1 (N564, N557);
or OR2 (N565, N560, N342);
not NOT1 (N566, N554);
or OR3 (N567, N553, N207, N386);
nand NAND4 (N568, N566, N457, N255, N189);
not NOT1 (N569, N563);
nor NOR3 (N570, N569, N439, N531);
or OR4 (N571, N568, N73, N507, N209);
and AND3 (N572, N552, N198, N250);
nand NAND3 (N573, N565, N436, N453);
not NOT1 (N574, N572);
and AND3 (N575, N574, N496, N237);
not NOT1 (N576, N564);
nor NOR2 (N577, N576, N227);
not NOT1 (N578, N559);
nor NOR2 (N579, N570, N138);
not NOT1 (N580, N578);
buf BUF1 (N581, N549);
not NOT1 (N582, N579);
nor NOR3 (N583, N580, N378, N293);
and AND3 (N584, N561, N30, N466);
xor XOR2 (N585, N571, N313);
nor NOR3 (N586, N575, N218, N492);
or OR3 (N587, N586, N188, N547);
nor NOR2 (N588, N577, N60);
or OR3 (N589, N585, N157, N156);
buf BUF1 (N590, N567);
not NOT1 (N591, N584);
not NOT1 (N592, N589);
xor XOR2 (N593, N590, N248);
nor NOR4 (N594, N588, N576, N449, N123);
and AND2 (N595, N556, N403);
xor XOR2 (N596, N593, N43);
buf BUF1 (N597, N581);
nand NAND2 (N598, N587, N64);
not NOT1 (N599, N592);
or OR4 (N600, N597, N20, N422, N400);
xor XOR2 (N601, N596, N409);
buf BUF1 (N602, N601);
or OR4 (N603, N602, N117, N390, N166);
nor NOR4 (N604, N599, N597, N199, N558);
nor NOR4 (N605, N604, N588, N176, N186);
and AND3 (N606, N582, N461, N127);
nand NAND4 (N607, N594, N449, N557, N535);
or OR2 (N608, N598, N573);
and AND4 (N609, N549, N542, N584, N530);
nand NAND3 (N610, N595, N409, N73);
nand NAND2 (N611, N609, N593);
not NOT1 (N612, N608);
xor XOR2 (N613, N600, N369);
not NOT1 (N614, N591);
nand NAND4 (N615, N603, N460, N175, N42);
nor NOR2 (N616, N614, N290);
and AND2 (N617, N605, N387);
nor NOR2 (N618, N616, N160);
not NOT1 (N619, N606);
xor XOR2 (N620, N611, N230);
xor XOR2 (N621, N613, N486);
nand NAND2 (N622, N617, N68);
nor NOR4 (N623, N607, N237, N35, N37);
not NOT1 (N624, N622);
and AND4 (N625, N619, N391, N341, N205);
nand NAND3 (N626, N620, N390, N15);
not NOT1 (N627, N625);
not NOT1 (N628, N623);
and AND3 (N629, N610, N445, N73);
not NOT1 (N630, N615);
or OR4 (N631, N629, N44, N552, N240);
nand NAND2 (N632, N628, N502);
or OR3 (N633, N631, N4, N245);
and AND4 (N634, N627, N560, N597, N235);
buf BUF1 (N635, N630);
buf BUF1 (N636, N632);
not NOT1 (N637, N621);
nand NAND2 (N638, N583, N358);
xor XOR2 (N639, N633, N583);
or OR3 (N640, N624, N228, N351);
xor XOR2 (N641, N634, N635);
xor XOR2 (N642, N89, N281);
and AND3 (N643, N641, N203, N26);
buf BUF1 (N644, N618);
buf BUF1 (N645, N637);
buf BUF1 (N646, N639);
and AND2 (N647, N643, N512);
or OR3 (N648, N646, N310, N640);
nand NAND3 (N649, N288, N77, N542);
nor NOR4 (N650, N636, N140, N171, N72);
nand NAND4 (N651, N650, N428, N326, N644);
buf BUF1 (N652, N529);
or OR3 (N653, N612, N297, N302);
xor XOR2 (N654, N653, N571);
nand NAND4 (N655, N626, N33, N19, N543);
nand NAND2 (N656, N642, N594);
not NOT1 (N657, N655);
nand NAND2 (N658, N652, N380);
buf BUF1 (N659, N657);
not NOT1 (N660, N638);
xor XOR2 (N661, N654, N59);
xor XOR2 (N662, N648, N367);
and AND2 (N663, N661, N144);
nor NOR2 (N664, N662, N457);
or OR3 (N665, N649, N449, N589);
and AND4 (N666, N659, N28, N459, N32);
not NOT1 (N667, N651);
nor NOR2 (N668, N663, N321);
and AND2 (N669, N666, N108);
or OR3 (N670, N660, N142, N129);
and AND2 (N671, N669, N76);
not NOT1 (N672, N664);
nor NOR4 (N673, N670, N637, N360, N597);
nor NOR4 (N674, N645, N640, N169, N8);
nand NAND2 (N675, N668, N31);
and AND4 (N676, N665, N594, N357, N285);
nor NOR2 (N677, N673, N2);
or OR2 (N678, N656, N228);
nand NAND3 (N679, N672, N286, N147);
not NOT1 (N680, N667);
nor NOR4 (N681, N678, N527, N251, N326);
nor NOR2 (N682, N681, N407);
or OR2 (N683, N679, N628);
nor NOR4 (N684, N647, N575, N12, N17);
nor NOR4 (N685, N677, N364, N136, N438);
not NOT1 (N686, N676);
nand NAND2 (N687, N683, N15);
nand NAND4 (N688, N680, N462, N627, N403);
nor NOR2 (N689, N658, N327);
buf BUF1 (N690, N686);
and AND4 (N691, N690, N413, N682, N364);
and AND2 (N692, N684, N52);
buf BUF1 (N693, N437);
not NOT1 (N694, N693);
xor XOR2 (N695, N692, N669);
not NOT1 (N696, N675);
nand NAND4 (N697, N689, N655, N411, N519);
not NOT1 (N698, N694);
or OR4 (N699, N685, N607, N24, N214);
buf BUF1 (N700, N696);
buf BUF1 (N701, N688);
and AND2 (N702, N700, N244);
xor XOR2 (N703, N701, N77);
xor XOR2 (N704, N703, N456);
nand NAND4 (N705, N699, N541, N238, N35);
xor XOR2 (N706, N691, N493);
or OR3 (N707, N695, N538, N98);
or OR3 (N708, N706, N345, N577);
not NOT1 (N709, N704);
nor NOR3 (N710, N671, N277, N627);
nor NOR3 (N711, N707, N238, N443);
and AND3 (N712, N687, N683, N491);
buf BUF1 (N713, N712);
not NOT1 (N714, N708);
xor XOR2 (N715, N710, N673);
not NOT1 (N716, N715);
not NOT1 (N717, N698);
nor NOR4 (N718, N717, N405, N495, N385);
not NOT1 (N719, N702);
and AND3 (N720, N713, N176, N596);
or OR3 (N721, N714, N578, N589);
nand NAND4 (N722, N697, N400, N348, N277);
buf BUF1 (N723, N711);
or OR3 (N724, N716, N152, N86);
nor NOR3 (N725, N722, N390, N58);
buf BUF1 (N726, N709);
nand NAND2 (N727, N674, N437);
nand NAND4 (N728, N720, N62, N129, N348);
or OR2 (N729, N725, N297);
not NOT1 (N730, N728);
nor NOR3 (N731, N729, N234, N265);
and AND4 (N732, N730, N54, N507, N523);
buf BUF1 (N733, N705);
nor NOR3 (N734, N723, N243, N337);
not NOT1 (N735, N733);
and AND4 (N736, N726, N298, N585, N200);
and AND2 (N737, N721, N190);
nor NOR2 (N738, N734, N324);
xor XOR2 (N739, N731, N495);
nand NAND4 (N740, N738, N700, N654, N349);
nor NOR4 (N741, N727, N427, N37, N508);
or OR2 (N742, N732, N479);
xor XOR2 (N743, N741, N128);
nor NOR4 (N744, N739, N49, N441, N452);
nor NOR2 (N745, N724, N426);
nor NOR2 (N746, N744, N130);
nand NAND4 (N747, N743, N57, N549, N544);
nor NOR2 (N748, N742, N740);
not NOT1 (N749, N36);
nor NOR4 (N750, N745, N318, N657, N116);
nor NOR3 (N751, N719, N683, N676);
xor XOR2 (N752, N747, N9);
or OR4 (N753, N736, N262, N685, N21);
xor XOR2 (N754, N752, N54);
not NOT1 (N755, N735);
xor XOR2 (N756, N718, N42);
not NOT1 (N757, N756);
nor NOR4 (N758, N753, N403, N85, N491);
and AND4 (N759, N750, N556, N3, N12);
not NOT1 (N760, N758);
xor XOR2 (N761, N759, N538);
xor XOR2 (N762, N757, N200);
and AND4 (N763, N761, N556, N419, N672);
buf BUF1 (N764, N748);
xor XOR2 (N765, N746, N520);
not NOT1 (N766, N764);
or OR2 (N767, N766, N555);
buf BUF1 (N768, N765);
nand NAND2 (N769, N768, N380);
not NOT1 (N770, N769);
and AND3 (N771, N751, N535, N61);
nand NAND3 (N772, N762, N269, N265);
not NOT1 (N773, N760);
nor NOR2 (N774, N767, N212);
or OR3 (N775, N771, N150, N621);
nor NOR4 (N776, N772, N644, N393, N658);
not NOT1 (N777, N775);
xor XOR2 (N778, N763, N280);
and AND3 (N779, N776, N726, N278);
not NOT1 (N780, N755);
and AND2 (N781, N754, N24);
and AND3 (N782, N770, N460, N117);
and AND3 (N783, N778, N627, N220);
buf BUF1 (N784, N777);
nor NOR2 (N785, N782, N183);
xor XOR2 (N786, N779, N206);
buf BUF1 (N787, N737);
buf BUF1 (N788, N783);
and AND3 (N789, N787, N786, N83);
nor NOR4 (N790, N561, N142, N115, N277);
xor XOR2 (N791, N773, N759);
xor XOR2 (N792, N790, N511);
not NOT1 (N793, N785);
nand NAND4 (N794, N789, N643, N709, N129);
nor NOR3 (N795, N784, N172, N263);
xor XOR2 (N796, N774, N627);
nor NOR4 (N797, N795, N646, N429, N480);
buf BUF1 (N798, N781);
nor NOR3 (N799, N797, N442, N55);
or OR4 (N800, N749, N264, N444, N621);
nand NAND2 (N801, N788, N143);
or OR4 (N802, N799, N294, N768, N722);
not NOT1 (N803, N794);
buf BUF1 (N804, N798);
xor XOR2 (N805, N791, N60);
nor NOR4 (N806, N792, N374, N753, N556);
not NOT1 (N807, N801);
or OR3 (N808, N804, N753, N529);
or OR4 (N809, N803, N260, N788, N45);
not NOT1 (N810, N805);
or OR2 (N811, N810, N808);
or OR2 (N812, N48, N556);
and AND2 (N813, N806, N277);
or OR3 (N814, N796, N446, N590);
or OR2 (N815, N802, N189);
buf BUF1 (N816, N815);
and AND2 (N817, N811, N34);
and AND4 (N818, N813, N614, N785, N758);
xor XOR2 (N819, N814, N278);
buf BUF1 (N820, N812);
or OR3 (N821, N818, N173, N349);
xor XOR2 (N822, N817, N669);
nor NOR2 (N823, N793, N623);
xor XOR2 (N824, N823, N261);
or OR2 (N825, N822, N310);
and AND2 (N826, N780, N426);
and AND2 (N827, N816, N44);
not NOT1 (N828, N826);
and AND3 (N829, N820, N307, N18);
nand NAND2 (N830, N821, N616);
not NOT1 (N831, N807);
and AND2 (N832, N828, N745);
not NOT1 (N833, N825);
xor XOR2 (N834, N829, N289);
buf BUF1 (N835, N819);
xor XOR2 (N836, N830, N441);
nand NAND2 (N837, N834, N221);
xor XOR2 (N838, N835, N373);
and AND3 (N839, N832, N787, N711);
or OR2 (N840, N824, N300);
or OR3 (N841, N837, N639, N272);
nor NOR4 (N842, N800, N80, N747, N550);
buf BUF1 (N843, N841);
not NOT1 (N844, N840);
not NOT1 (N845, N839);
or OR3 (N846, N842, N196, N80);
nor NOR3 (N847, N838, N811, N676);
xor XOR2 (N848, N845, N542);
and AND3 (N849, N846, N399, N453);
buf BUF1 (N850, N848);
not NOT1 (N851, N827);
xor XOR2 (N852, N850, N805);
xor XOR2 (N853, N847, N25);
nand NAND3 (N854, N833, N653, N436);
or OR3 (N855, N851, N138, N740);
nand NAND4 (N856, N852, N445, N26, N62);
or OR4 (N857, N854, N110, N564, N312);
or OR4 (N858, N853, N724, N5, N208);
nand NAND4 (N859, N856, N454, N418, N810);
nor NOR2 (N860, N858, N671);
nand NAND3 (N861, N849, N60, N738);
and AND4 (N862, N844, N68, N290, N578);
or OR4 (N863, N836, N774, N179, N608);
and AND3 (N864, N860, N671, N125);
and AND4 (N865, N831, N352, N391, N453);
and AND2 (N866, N857, N670);
xor XOR2 (N867, N843, N686);
not NOT1 (N868, N864);
buf BUF1 (N869, N859);
and AND4 (N870, N862, N772, N107, N360);
and AND2 (N871, N867, N763);
xor XOR2 (N872, N871, N33);
buf BUF1 (N873, N863);
nand NAND4 (N874, N855, N765, N243, N342);
nor NOR2 (N875, N870, N22);
and AND3 (N876, N868, N342, N531);
not NOT1 (N877, N872);
xor XOR2 (N878, N809, N8);
buf BUF1 (N879, N876);
xor XOR2 (N880, N875, N209);
or OR4 (N881, N878, N172, N832, N510);
buf BUF1 (N882, N881);
nor NOR4 (N883, N877, N831, N590, N466);
xor XOR2 (N884, N879, N388);
nor NOR2 (N885, N873, N632);
xor XOR2 (N886, N884, N129);
or OR2 (N887, N861, N370);
xor XOR2 (N888, N883, N771);
nand NAND2 (N889, N866, N111);
not NOT1 (N890, N885);
not NOT1 (N891, N890);
or OR2 (N892, N874, N187);
nand NAND2 (N893, N892, N301);
xor XOR2 (N894, N888, N66);
and AND3 (N895, N886, N153, N576);
nand NAND3 (N896, N895, N575, N312);
nand NAND2 (N897, N887, N659);
buf BUF1 (N898, N893);
nor NOR4 (N899, N891, N299, N406, N526);
buf BUF1 (N900, N897);
xor XOR2 (N901, N889, N756);
nand NAND3 (N902, N900, N731, N710);
and AND4 (N903, N894, N586, N277, N856);
or OR2 (N904, N899, N665);
and AND3 (N905, N896, N854, N855);
or OR2 (N906, N905, N788);
nor NOR2 (N907, N906, N188);
and AND2 (N908, N903, N34);
buf BUF1 (N909, N865);
xor XOR2 (N910, N902, N213);
xor XOR2 (N911, N880, N499);
not NOT1 (N912, N910);
nand NAND2 (N913, N869, N534);
nor NOR4 (N914, N901, N567, N374, N347);
buf BUF1 (N915, N904);
and AND2 (N916, N907, N552);
not NOT1 (N917, N913);
not NOT1 (N918, N908);
or OR2 (N919, N909, N62);
buf BUF1 (N920, N914);
nand NAND3 (N921, N920, N415, N301);
and AND3 (N922, N918, N906, N123);
and AND3 (N923, N912, N327, N461);
buf BUF1 (N924, N882);
nand NAND4 (N925, N917, N265, N548, N320);
buf BUF1 (N926, N923);
nand NAND2 (N927, N911, N404);
and AND3 (N928, N916, N556, N104);
xor XOR2 (N929, N898, N214);
xor XOR2 (N930, N927, N420);
nand NAND3 (N931, N929, N373, N630);
xor XOR2 (N932, N926, N418);
xor XOR2 (N933, N922, N432);
and AND2 (N934, N930, N199);
nand NAND2 (N935, N924, N98);
nor NOR2 (N936, N919, N612);
buf BUF1 (N937, N928);
not NOT1 (N938, N925);
buf BUF1 (N939, N937);
nand NAND4 (N940, N931, N100, N642, N109);
xor XOR2 (N941, N932, N321);
nor NOR4 (N942, N915, N67, N917, N741);
or OR2 (N943, N921, N430);
not NOT1 (N944, N941);
buf BUF1 (N945, N944);
buf BUF1 (N946, N945);
nor NOR4 (N947, N938, N662, N444, N709);
buf BUF1 (N948, N934);
xor XOR2 (N949, N936, N594);
buf BUF1 (N950, N935);
nor NOR2 (N951, N948, N641);
and AND4 (N952, N946, N469, N421, N88);
nor NOR2 (N953, N950, N446);
nand NAND3 (N954, N953, N385, N137);
nand NAND4 (N955, N939, N674, N67, N626);
nor NOR4 (N956, N943, N304, N923, N886);
or OR4 (N957, N949, N75, N178, N629);
nand NAND2 (N958, N933, N445);
xor XOR2 (N959, N955, N382);
nand NAND2 (N960, N951, N325);
or OR3 (N961, N958, N248, N813);
buf BUF1 (N962, N947);
nor NOR4 (N963, N960, N181, N396, N483);
xor XOR2 (N964, N961, N233);
and AND4 (N965, N954, N144, N500, N387);
not NOT1 (N966, N942);
or OR4 (N967, N965, N330, N537, N156);
buf BUF1 (N968, N964);
or OR2 (N969, N963, N471);
not NOT1 (N970, N940);
nand NAND2 (N971, N957, N481);
or OR3 (N972, N959, N849, N760);
nor NOR3 (N973, N956, N751, N876);
nand NAND2 (N974, N962, N768);
xor XOR2 (N975, N970, N308);
not NOT1 (N976, N967);
nand NAND2 (N977, N971, N577);
nand NAND4 (N978, N974, N129, N25, N834);
and AND4 (N979, N978, N23, N373, N553);
xor XOR2 (N980, N966, N865);
nand NAND2 (N981, N969, N337);
nand NAND2 (N982, N981, N67);
not NOT1 (N983, N972);
nor NOR4 (N984, N977, N470, N552, N595);
xor XOR2 (N985, N984, N771);
nor NOR4 (N986, N973, N867, N312, N153);
nand NAND3 (N987, N983, N845, N273);
buf BUF1 (N988, N986);
not NOT1 (N989, N979);
not NOT1 (N990, N976);
not NOT1 (N991, N952);
or OR4 (N992, N982, N752, N952, N78);
nand NAND4 (N993, N989, N527, N879, N366);
and AND4 (N994, N987, N103, N543, N378);
not NOT1 (N995, N980);
xor XOR2 (N996, N968, N992);
or OR3 (N997, N127, N281, N138);
or OR2 (N998, N996, N897);
xor XOR2 (N999, N993, N700);
not NOT1 (N1000, N997);
or OR2 (N1001, N994, N865);
nand NAND4 (N1002, N995, N312, N794, N154);
not NOT1 (N1003, N975);
or OR4 (N1004, N985, N993, N147, N720);
not NOT1 (N1005, N998);
buf BUF1 (N1006, N1004);
not NOT1 (N1007, N1005);
buf BUF1 (N1008, N1007);
buf BUF1 (N1009, N1003);
buf BUF1 (N1010, N1008);
buf BUF1 (N1011, N999);
nand NAND4 (N1012, N1002, N111, N527, N593);
buf BUF1 (N1013, N990);
nor NOR4 (N1014, N1001, N47, N319, N461);
nand NAND3 (N1015, N1000, N534, N572);
and AND4 (N1016, N991, N67, N518, N922);
nor NOR4 (N1017, N1012, N344, N349, N134);
nor NOR2 (N1018, N1013, N408);
or OR4 (N1019, N1010, N346, N688, N386);
xor XOR2 (N1020, N988, N458);
and AND4 (N1021, N1017, N361, N158, N614);
not NOT1 (N1022, N1006);
xor XOR2 (N1023, N1011, N1019);
and AND2 (N1024, N799, N242);
xor XOR2 (N1025, N1021, N1005);
and AND3 (N1026, N1014, N839, N67);
nor NOR2 (N1027, N1023, N141);
or OR4 (N1028, N1020, N947, N1019, N238);
xor XOR2 (N1029, N1028, N290);
nor NOR4 (N1030, N1026, N174, N619, N823);
nor NOR4 (N1031, N1016, N779, N407, N691);
and AND2 (N1032, N1025, N358);
not NOT1 (N1033, N1032);
or OR3 (N1034, N1018, N66, N612);
not NOT1 (N1035, N1034);
buf BUF1 (N1036, N1030);
or OR3 (N1037, N1036, N719, N432);
nor NOR3 (N1038, N1035, N519, N412);
or OR2 (N1039, N1024, N682);
xor XOR2 (N1040, N1029, N751);
nand NAND4 (N1041, N1039, N104, N792, N167);
nor NOR2 (N1042, N1037, N315);
xor XOR2 (N1043, N1027, N493);
not NOT1 (N1044, N1043);
or OR3 (N1045, N1038, N76, N761);
xor XOR2 (N1046, N1045, N606);
or OR3 (N1047, N1022, N693, N721);
nand NAND2 (N1048, N1047, N161);
not NOT1 (N1049, N1040);
or OR4 (N1050, N1009, N980, N584, N895);
nor NOR2 (N1051, N1015, N595);
nand NAND4 (N1052, N1046, N177, N793, N842);
buf BUF1 (N1053, N1033);
buf BUF1 (N1054, N1052);
not NOT1 (N1055, N1042);
nor NOR2 (N1056, N1055, N203);
buf BUF1 (N1057, N1041);
xor XOR2 (N1058, N1051, N486);
or OR3 (N1059, N1056, N386, N801);
nand NAND3 (N1060, N1059, N1029, N775);
or OR4 (N1061, N1044, N473, N287, N203);
or OR2 (N1062, N1054, N730);
nand NAND4 (N1063, N1057, N268, N554, N920);
xor XOR2 (N1064, N1049, N311);
nand NAND3 (N1065, N1063, N801, N219);
xor XOR2 (N1066, N1061, N278);
buf BUF1 (N1067, N1048);
or OR4 (N1068, N1062, N572, N135, N679);
nor NOR3 (N1069, N1058, N46, N610);
or OR3 (N1070, N1066, N961, N191);
xor XOR2 (N1071, N1050, N877);
not NOT1 (N1072, N1071);
buf BUF1 (N1073, N1070);
and AND3 (N1074, N1073, N95, N398);
buf BUF1 (N1075, N1064);
nand NAND2 (N1076, N1053, N180);
buf BUF1 (N1077, N1074);
not NOT1 (N1078, N1075);
nor NOR3 (N1079, N1067, N798, N619);
nor NOR2 (N1080, N1078, N943);
or OR2 (N1081, N1077, N449);
buf BUF1 (N1082, N1076);
not NOT1 (N1083, N1069);
xor XOR2 (N1084, N1060, N827);
xor XOR2 (N1085, N1080, N752);
not NOT1 (N1086, N1079);
and AND3 (N1087, N1083, N425, N958);
nand NAND4 (N1088, N1086, N881, N52, N673);
nand NAND2 (N1089, N1088, N925);
not NOT1 (N1090, N1082);
buf BUF1 (N1091, N1090);
nor NOR2 (N1092, N1081, N1);
not NOT1 (N1093, N1031);
and AND2 (N1094, N1093, N622);
not NOT1 (N1095, N1085);
and AND2 (N1096, N1072, N1070);
nor NOR3 (N1097, N1091, N434, N465);
nand NAND2 (N1098, N1095, N310);
nor NOR2 (N1099, N1092, N1039);
nor NOR4 (N1100, N1065, N97, N667, N979);
nor NOR4 (N1101, N1084, N929, N650, N782);
not NOT1 (N1102, N1096);
nand NAND4 (N1103, N1100, N52, N929, N72);
nand NAND2 (N1104, N1103, N911);
nor NOR4 (N1105, N1097, N8, N1052, N1085);
buf BUF1 (N1106, N1089);
nor NOR3 (N1107, N1101, N421, N518);
and AND3 (N1108, N1068, N292, N1004);
buf BUF1 (N1109, N1098);
xor XOR2 (N1110, N1105, N98);
nand NAND4 (N1111, N1106, N795, N494, N453);
and AND4 (N1112, N1102, N796, N512, N35);
xor XOR2 (N1113, N1104, N451);
nand NAND4 (N1114, N1107, N414, N870, N1112);
nand NAND4 (N1115, N67, N869, N1006, N799);
and AND4 (N1116, N1094, N461, N633, N989);
nor NOR3 (N1117, N1109, N387, N368);
nor NOR4 (N1118, N1087, N283, N24, N133);
nand NAND2 (N1119, N1116, N735);
nor NOR4 (N1120, N1117, N925, N177, N455);
nand NAND3 (N1121, N1115, N349, N363);
nor NOR3 (N1122, N1120, N883, N534);
or OR3 (N1123, N1113, N965, N1058);
or OR2 (N1124, N1118, N90);
and AND3 (N1125, N1121, N1068, N705);
and AND2 (N1126, N1110, N572);
not NOT1 (N1127, N1099);
xor XOR2 (N1128, N1124, N203);
xor XOR2 (N1129, N1128, N89);
buf BUF1 (N1130, N1129);
xor XOR2 (N1131, N1122, N639);
nand NAND4 (N1132, N1127, N858, N246, N1114);
and AND2 (N1133, N36, N90);
and AND2 (N1134, N1119, N255);
buf BUF1 (N1135, N1126);
nand NAND2 (N1136, N1125, N75);
and AND4 (N1137, N1130, N1056, N414, N725);
not NOT1 (N1138, N1134);
or OR4 (N1139, N1108, N957, N274, N60);
not NOT1 (N1140, N1135);
nand NAND2 (N1141, N1138, N547);
nor NOR2 (N1142, N1136, N325);
and AND2 (N1143, N1139, N265);
nor NOR2 (N1144, N1142, N690);
and AND3 (N1145, N1137, N626, N864);
nand NAND2 (N1146, N1123, N1080);
or OR2 (N1147, N1145, N1137);
buf BUF1 (N1148, N1147);
buf BUF1 (N1149, N1111);
buf BUF1 (N1150, N1146);
or OR2 (N1151, N1144, N770);
or OR2 (N1152, N1151, N906);
xor XOR2 (N1153, N1132, N1002);
xor XOR2 (N1154, N1153, N290);
and AND3 (N1155, N1148, N805, N891);
nor NOR3 (N1156, N1149, N573, N266);
nand NAND2 (N1157, N1150, N1073);
not NOT1 (N1158, N1155);
and AND3 (N1159, N1143, N6, N1105);
or OR2 (N1160, N1156, N937);
not NOT1 (N1161, N1140);
xor XOR2 (N1162, N1157, N760);
or OR2 (N1163, N1141, N1042);
nor NOR2 (N1164, N1159, N840);
and AND3 (N1165, N1160, N174, N116);
buf BUF1 (N1166, N1131);
nor NOR4 (N1167, N1164, N324, N289, N720);
or OR3 (N1168, N1152, N744, N241);
or OR3 (N1169, N1166, N905, N665);
xor XOR2 (N1170, N1169, N72);
or OR3 (N1171, N1162, N294, N103);
not NOT1 (N1172, N1163);
xor XOR2 (N1173, N1167, N463);
xor XOR2 (N1174, N1165, N826);
or OR2 (N1175, N1171, N888);
buf BUF1 (N1176, N1174);
nand NAND2 (N1177, N1133, N507);
not NOT1 (N1178, N1177);
or OR2 (N1179, N1176, N435);
nand NAND3 (N1180, N1161, N1096, N901);
or OR3 (N1181, N1179, N2, N45);
buf BUF1 (N1182, N1178);
buf BUF1 (N1183, N1182);
not NOT1 (N1184, N1158);
nor NOR4 (N1185, N1183, N131, N274, N1076);
and AND4 (N1186, N1168, N754, N362, N1029);
buf BUF1 (N1187, N1154);
and AND3 (N1188, N1185, N1079, N884);
xor XOR2 (N1189, N1170, N97);
nand NAND2 (N1190, N1184, N517);
and AND2 (N1191, N1173, N837);
nand NAND4 (N1192, N1191, N473, N294, N860);
and AND2 (N1193, N1181, N1172);
not NOT1 (N1194, N406);
or OR4 (N1195, N1186, N16, N467, N787);
nor NOR4 (N1196, N1193, N1116, N404, N1046);
buf BUF1 (N1197, N1187);
buf BUF1 (N1198, N1195);
nor NOR4 (N1199, N1194, N240, N183, N786);
or OR2 (N1200, N1197, N1081);
xor XOR2 (N1201, N1189, N164);
xor XOR2 (N1202, N1201, N290);
and AND4 (N1203, N1192, N658, N618, N859);
nand NAND3 (N1204, N1196, N792, N803);
buf BUF1 (N1205, N1199);
buf BUF1 (N1206, N1200);
or OR2 (N1207, N1175, N958);
not NOT1 (N1208, N1198);
not NOT1 (N1209, N1202);
nand NAND4 (N1210, N1203, N188, N1146, N496);
nand NAND2 (N1211, N1208, N280);
or OR4 (N1212, N1190, N1057, N189, N1017);
nor NOR4 (N1213, N1212, N1049, N807, N653);
nor NOR3 (N1214, N1209, N797, N259);
not NOT1 (N1215, N1180);
or OR3 (N1216, N1206, N1023, N1110);
or OR3 (N1217, N1207, N984, N419);
xor XOR2 (N1218, N1215, N109);
or OR2 (N1219, N1214, N363);
nand NAND2 (N1220, N1219, N1115);
nand NAND4 (N1221, N1218, N774, N1019, N488);
or OR4 (N1222, N1205, N1147, N929, N62);
nand NAND4 (N1223, N1188, N229, N640, N214);
not NOT1 (N1224, N1211);
nand NAND2 (N1225, N1223, N816);
nand NAND2 (N1226, N1222, N959);
xor XOR2 (N1227, N1226, N1045);
nand NAND3 (N1228, N1224, N1060, N541);
xor XOR2 (N1229, N1210, N836);
buf BUF1 (N1230, N1227);
or OR2 (N1231, N1217, N429);
or OR4 (N1232, N1220, N13, N557, N1010);
nor NOR2 (N1233, N1216, N585);
and AND2 (N1234, N1229, N968);
buf BUF1 (N1235, N1204);
and AND2 (N1236, N1228, N685);
xor XOR2 (N1237, N1231, N789);
xor XOR2 (N1238, N1236, N738);
nand NAND4 (N1239, N1230, N100, N138, N1021);
nand NAND3 (N1240, N1234, N557, N413);
buf BUF1 (N1241, N1240);
or OR4 (N1242, N1221, N989, N1216, N345);
not NOT1 (N1243, N1213);
or OR4 (N1244, N1241, N916, N648, N347);
xor XOR2 (N1245, N1242, N991);
xor XOR2 (N1246, N1238, N482);
nor NOR3 (N1247, N1233, N559, N1211);
and AND2 (N1248, N1237, N600);
buf BUF1 (N1249, N1244);
xor XOR2 (N1250, N1239, N1124);
not NOT1 (N1251, N1235);
or OR2 (N1252, N1250, N1192);
xor XOR2 (N1253, N1245, N950);
not NOT1 (N1254, N1225);
buf BUF1 (N1255, N1251);
nand NAND4 (N1256, N1248, N951, N994, N279);
nor NOR4 (N1257, N1243, N143, N1058, N1010);
xor XOR2 (N1258, N1232, N530);
not NOT1 (N1259, N1256);
buf BUF1 (N1260, N1249);
or OR2 (N1261, N1258, N1139);
and AND3 (N1262, N1247, N783, N286);
and AND2 (N1263, N1260, N1217);
xor XOR2 (N1264, N1246, N26);
not NOT1 (N1265, N1255);
not NOT1 (N1266, N1252);
not NOT1 (N1267, N1254);
and AND2 (N1268, N1265, N245);
not NOT1 (N1269, N1262);
nor NOR2 (N1270, N1259, N239);
buf BUF1 (N1271, N1267);
nor NOR3 (N1272, N1264, N1014, N426);
not NOT1 (N1273, N1261);
xor XOR2 (N1274, N1270, N516);
nor NOR4 (N1275, N1268, N650, N1075, N488);
and AND4 (N1276, N1272, N1203, N1250, N457);
not NOT1 (N1277, N1253);
not NOT1 (N1278, N1273);
and AND4 (N1279, N1266, N403, N61, N622);
xor XOR2 (N1280, N1276, N1137);
not NOT1 (N1281, N1271);
buf BUF1 (N1282, N1278);
xor XOR2 (N1283, N1274, N1242);
or OR2 (N1284, N1269, N497);
and AND2 (N1285, N1284, N810);
nand NAND3 (N1286, N1282, N1197, N116);
xor XOR2 (N1287, N1279, N1232);
not NOT1 (N1288, N1285);
buf BUF1 (N1289, N1286);
buf BUF1 (N1290, N1281);
not NOT1 (N1291, N1257);
nand NAND2 (N1292, N1290, N398);
nor NOR2 (N1293, N1280, N476);
or OR3 (N1294, N1291, N429, N265);
xor XOR2 (N1295, N1292, N875);
nor NOR2 (N1296, N1283, N716);
nor NOR2 (N1297, N1287, N970);
or OR4 (N1298, N1293, N1287, N846, N443);
buf BUF1 (N1299, N1277);
not NOT1 (N1300, N1298);
nor NOR4 (N1301, N1300, N1150, N799, N56);
not NOT1 (N1302, N1263);
nand NAND3 (N1303, N1288, N171, N49);
xor XOR2 (N1304, N1289, N1114);
buf BUF1 (N1305, N1275);
not NOT1 (N1306, N1295);
and AND3 (N1307, N1302, N1035, N586);
buf BUF1 (N1308, N1305);
xor XOR2 (N1309, N1308, N211);
xor XOR2 (N1310, N1294, N639);
xor XOR2 (N1311, N1304, N1007);
buf BUF1 (N1312, N1296);
xor XOR2 (N1313, N1310, N193);
nor NOR2 (N1314, N1313, N1003);
and AND2 (N1315, N1299, N431);
and AND4 (N1316, N1309, N1036, N1167, N1249);
or OR2 (N1317, N1311, N439);
nand NAND4 (N1318, N1301, N407, N1129, N928);
nand NAND4 (N1319, N1318, N164, N355, N1011);
buf BUF1 (N1320, N1316);
not NOT1 (N1321, N1315);
not NOT1 (N1322, N1312);
or OR2 (N1323, N1307, N1002);
nand NAND4 (N1324, N1314, N123, N23, N1144);
nand NAND3 (N1325, N1319, N362, N1187);
xor XOR2 (N1326, N1323, N238);
nand NAND3 (N1327, N1320, N170, N1140);
or OR2 (N1328, N1325, N105);
xor XOR2 (N1329, N1303, N740);
buf BUF1 (N1330, N1297);
nand NAND2 (N1331, N1329, N1078);
xor XOR2 (N1332, N1322, N91);
or OR2 (N1333, N1332, N1134);
buf BUF1 (N1334, N1328);
or OR3 (N1335, N1330, N825, N547);
nand NAND3 (N1336, N1321, N1116, N121);
nand NAND4 (N1337, N1331, N522, N956, N1185);
and AND3 (N1338, N1306, N710, N628);
buf BUF1 (N1339, N1333);
buf BUF1 (N1340, N1335);
or OR2 (N1341, N1327, N714);
not NOT1 (N1342, N1341);
and AND4 (N1343, N1342, N1268, N1263, N307);
xor XOR2 (N1344, N1336, N132);
nor NOR4 (N1345, N1338, N1307, N383, N943);
nor NOR2 (N1346, N1317, N294);
not NOT1 (N1347, N1339);
and AND4 (N1348, N1337, N818, N1259, N404);
buf BUF1 (N1349, N1346);
not NOT1 (N1350, N1347);
buf BUF1 (N1351, N1345);
and AND4 (N1352, N1334, N961, N1091, N554);
nor NOR4 (N1353, N1326, N1334, N1189, N608);
and AND4 (N1354, N1340, N747, N1086, N1163);
nand NAND4 (N1355, N1352, N964, N1225, N1284);
or OR3 (N1356, N1354, N74, N1059);
buf BUF1 (N1357, N1350);
nor NOR3 (N1358, N1357, N992, N184);
xor XOR2 (N1359, N1353, N743);
not NOT1 (N1360, N1359);
or OR2 (N1361, N1343, N640);
buf BUF1 (N1362, N1356);
xor XOR2 (N1363, N1361, N324);
and AND3 (N1364, N1358, N1140, N231);
and AND3 (N1365, N1324, N200, N767);
not NOT1 (N1366, N1349);
not NOT1 (N1367, N1360);
buf BUF1 (N1368, N1363);
and AND4 (N1369, N1355, N441, N1002, N1341);
not NOT1 (N1370, N1344);
nor NOR2 (N1371, N1369, N593);
and AND2 (N1372, N1370, N1312);
xor XOR2 (N1373, N1368, N788);
not NOT1 (N1374, N1365);
not NOT1 (N1375, N1374);
xor XOR2 (N1376, N1366, N149);
nor NOR4 (N1377, N1348, N966, N327, N738);
xor XOR2 (N1378, N1367, N1274);
and AND2 (N1379, N1377, N871);
nor NOR3 (N1380, N1364, N94, N1342);
nand NAND3 (N1381, N1373, N31, N1323);
nand NAND2 (N1382, N1371, N953);
nand NAND4 (N1383, N1375, N824, N889, N1073);
nand NAND2 (N1384, N1372, N138);
xor XOR2 (N1385, N1381, N936);
not NOT1 (N1386, N1383);
or OR2 (N1387, N1362, N1145);
nor NOR3 (N1388, N1386, N705, N243);
xor XOR2 (N1389, N1388, N659);
buf BUF1 (N1390, N1389);
nor NOR3 (N1391, N1382, N364, N1003);
xor XOR2 (N1392, N1379, N236);
not NOT1 (N1393, N1380);
nor NOR3 (N1394, N1376, N365, N779);
nor NOR3 (N1395, N1391, N655, N693);
buf BUF1 (N1396, N1395);
buf BUF1 (N1397, N1378);
buf BUF1 (N1398, N1397);
not NOT1 (N1399, N1387);
not NOT1 (N1400, N1351);
buf BUF1 (N1401, N1400);
and AND3 (N1402, N1396, N210, N11);
and AND3 (N1403, N1402, N696, N337);
nor NOR4 (N1404, N1398, N380, N658, N551);
not NOT1 (N1405, N1385);
xor XOR2 (N1406, N1401, N1148);
not NOT1 (N1407, N1405);
nand NAND2 (N1408, N1392, N826);
buf BUF1 (N1409, N1384);
xor XOR2 (N1410, N1399, N359);
and AND3 (N1411, N1403, N1232, N1005);
not NOT1 (N1412, N1406);
xor XOR2 (N1413, N1411, N904);
nand NAND2 (N1414, N1393, N1171);
buf BUF1 (N1415, N1413);
nand NAND3 (N1416, N1394, N57, N355);
and AND3 (N1417, N1414, N1359, N830);
buf BUF1 (N1418, N1416);
buf BUF1 (N1419, N1404);
buf BUF1 (N1420, N1417);
or OR4 (N1421, N1412, N412, N1086, N653);
nor NOR3 (N1422, N1419, N1195, N324);
nand NAND2 (N1423, N1409, N302);
and AND3 (N1424, N1422, N1112, N1157);
nand NAND2 (N1425, N1410, N721);
buf BUF1 (N1426, N1415);
xor XOR2 (N1427, N1423, N1185);
or OR2 (N1428, N1418, N1411);
nor NOR2 (N1429, N1427, N1124);
or OR4 (N1430, N1429, N791, N94, N508);
not NOT1 (N1431, N1428);
buf BUF1 (N1432, N1421);
and AND2 (N1433, N1424, N1227);
nor NOR4 (N1434, N1432, N1237, N478, N127);
not NOT1 (N1435, N1426);
buf BUF1 (N1436, N1390);
or OR2 (N1437, N1408, N422);
buf BUF1 (N1438, N1407);
xor XOR2 (N1439, N1435, N408);
xor XOR2 (N1440, N1433, N673);
or OR3 (N1441, N1439, N1003, N229);
xor XOR2 (N1442, N1425, N843);
xor XOR2 (N1443, N1436, N1063);
nor NOR4 (N1444, N1442, N948, N461, N625);
not NOT1 (N1445, N1437);
nor NOR2 (N1446, N1431, N1347);
and AND2 (N1447, N1443, N1168);
or OR3 (N1448, N1420, N196, N915);
nand NAND2 (N1449, N1434, N478);
not NOT1 (N1450, N1441);
xor XOR2 (N1451, N1440, N282);
not NOT1 (N1452, N1430);
nor NOR3 (N1453, N1444, N1433, N501);
and AND4 (N1454, N1438, N16, N985, N655);
not NOT1 (N1455, N1448);
xor XOR2 (N1456, N1446, N959);
or OR2 (N1457, N1455, N1234);
and AND3 (N1458, N1450, N1043, N1118);
or OR4 (N1459, N1457, N817, N1362, N900);
xor XOR2 (N1460, N1454, N1449);
not NOT1 (N1461, N909);
buf BUF1 (N1462, N1459);
and AND3 (N1463, N1445, N115, N267);
and AND4 (N1464, N1452, N668, N482, N1017);
and AND3 (N1465, N1453, N1193, N1155);
buf BUF1 (N1466, N1456);
not NOT1 (N1467, N1460);
nand NAND4 (N1468, N1451, N205, N1352, N819);
nand NAND2 (N1469, N1467, N924);
nand NAND4 (N1470, N1447, N631, N1081, N1301);
nand NAND4 (N1471, N1468, N748, N1374, N83);
and AND3 (N1472, N1465, N734, N1315);
buf BUF1 (N1473, N1461);
not NOT1 (N1474, N1469);
or OR3 (N1475, N1466, N1118, N1033);
not NOT1 (N1476, N1475);
not NOT1 (N1477, N1470);
buf BUF1 (N1478, N1473);
buf BUF1 (N1479, N1463);
nor NOR2 (N1480, N1478, N20);
buf BUF1 (N1481, N1477);
buf BUF1 (N1482, N1480);
nor NOR2 (N1483, N1462, N685);
not NOT1 (N1484, N1464);
and AND4 (N1485, N1472, N1238, N116, N407);
not NOT1 (N1486, N1481);
and AND3 (N1487, N1484, N569, N120);
not NOT1 (N1488, N1458);
and AND2 (N1489, N1471, N88);
nor NOR4 (N1490, N1476, N1220, N1234, N1263);
xor XOR2 (N1491, N1486, N1144);
xor XOR2 (N1492, N1482, N485);
or OR4 (N1493, N1487, N80, N896, N1005);
not NOT1 (N1494, N1492);
xor XOR2 (N1495, N1485, N1040);
buf BUF1 (N1496, N1493);
buf BUF1 (N1497, N1494);
xor XOR2 (N1498, N1497, N613);
or OR4 (N1499, N1498, N833, N329, N442);
not NOT1 (N1500, N1490);
nor NOR3 (N1501, N1496, N962, N1378);
not NOT1 (N1502, N1479);
not NOT1 (N1503, N1495);
not NOT1 (N1504, N1502);
buf BUF1 (N1505, N1483);
not NOT1 (N1506, N1500);
nor NOR4 (N1507, N1488, N1343, N1406, N631);
nor NOR4 (N1508, N1474, N338, N1481, N1311);
nor NOR3 (N1509, N1501, N913, N646);
nor NOR3 (N1510, N1506, N1349, N894);
nand NAND3 (N1511, N1499, N1331, N756);
xor XOR2 (N1512, N1491, N1356);
xor XOR2 (N1513, N1505, N344);
buf BUF1 (N1514, N1512);
xor XOR2 (N1515, N1513, N905);
buf BUF1 (N1516, N1489);
and AND3 (N1517, N1508, N1366, N886);
xor XOR2 (N1518, N1503, N121);
or OR4 (N1519, N1510, N624, N27, N778);
nand NAND4 (N1520, N1518, N683, N831, N218);
buf BUF1 (N1521, N1504);
nor NOR4 (N1522, N1507, N1409, N574, N55);
nor NOR3 (N1523, N1509, N30, N784);
not NOT1 (N1524, N1522);
buf BUF1 (N1525, N1515);
not NOT1 (N1526, N1514);
not NOT1 (N1527, N1525);
buf BUF1 (N1528, N1516);
buf BUF1 (N1529, N1528);
and AND4 (N1530, N1517, N1424, N1004, N714);
nand NAND3 (N1531, N1523, N1297, N645);
nand NAND2 (N1532, N1529, N875);
not NOT1 (N1533, N1521);
and AND4 (N1534, N1511, N1304, N1480, N1365);
buf BUF1 (N1535, N1526);
nor NOR3 (N1536, N1527, N655, N868);
nand NAND4 (N1537, N1519, N719, N662, N373);
nor NOR2 (N1538, N1531, N642);
buf BUF1 (N1539, N1524);
not NOT1 (N1540, N1538);
nor NOR4 (N1541, N1530, N876, N1451, N1462);
and AND4 (N1542, N1535, N1041, N1412, N869);
not NOT1 (N1543, N1536);
xor XOR2 (N1544, N1532, N447);
xor XOR2 (N1545, N1540, N580);
or OR4 (N1546, N1533, N1242, N227, N338);
not NOT1 (N1547, N1537);
xor XOR2 (N1548, N1520, N402);
buf BUF1 (N1549, N1545);
buf BUF1 (N1550, N1548);
nor NOR4 (N1551, N1546, N912, N95, N1001);
or OR2 (N1552, N1547, N691);
nand NAND2 (N1553, N1543, N1295);
and AND3 (N1554, N1539, N835, N81);
buf BUF1 (N1555, N1541);
or OR4 (N1556, N1555, N103, N552, N942);
buf BUF1 (N1557, N1534);
nand NAND4 (N1558, N1549, N1337, N642, N1278);
not NOT1 (N1559, N1551);
nor NOR4 (N1560, N1556, N383, N245, N1115);
nand NAND3 (N1561, N1557, N948, N807);
nand NAND4 (N1562, N1554, N81, N733, N1142);
or OR4 (N1563, N1544, N109, N612, N1441);
xor XOR2 (N1564, N1559, N1414);
or OR4 (N1565, N1542, N1031, N1549, N1540);
xor XOR2 (N1566, N1552, N111);
xor XOR2 (N1567, N1558, N1249);
and AND2 (N1568, N1564, N919);
and AND3 (N1569, N1567, N1191, N524);
not NOT1 (N1570, N1553);
buf BUF1 (N1571, N1562);
and AND4 (N1572, N1568, N64, N1480, N981);
buf BUF1 (N1573, N1569);
nand NAND3 (N1574, N1563, N305, N966);
nor NOR2 (N1575, N1574, N1002);
xor XOR2 (N1576, N1560, N1110);
buf BUF1 (N1577, N1566);
or OR4 (N1578, N1565, N357, N1533, N393);
and AND4 (N1579, N1550, N1036, N693, N365);
xor XOR2 (N1580, N1575, N583);
and AND3 (N1581, N1571, N1143, N199);
buf BUF1 (N1582, N1572);
and AND4 (N1583, N1576, N686, N735, N407);
and AND2 (N1584, N1579, N168);
buf BUF1 (N1585, N1577);
xor XOR2 (N1586, N1580, N333);
not NOT1 (N1587, N1578);
xor XOR2 (N1588, N1587, N876);
and AND3 (N1589, N1586, N1047, N1338);
buf BUF1 (N1590, N1570);
nor NOR2 (N1591, N1585, N1494);
nor NOR2 (N1592, N1583, N1218);
and AND3 (N1593, N1592, N1447, N183);
buf BUF1 (N1594, N1573);
or OR2 (N1595, N1561, N122);
buf BUF1 (N1596, N1584);
nor NOR2 (N1597, N1594, N52);
xor XOR2 (N1598, N1588, N413);
buf BUF1 (N1599, N1598);
xor XOR2 (N1600, N1591, N1516);
and AND4 (N1601, N1593, N587, N51, N1421);
nand NAND2 (N1602, N1597, N1532);
and AND2 (N1603, N1601, N789);
nand NAND3 (N1604, N1596, N294, N119);
nor NOR3 (N1605, N1600, N1600, N978);
buf BUF1 (N1606, N1602);
and AND2 (N1607, N1590, N1243);
or OR4 (N1608, N1599, N777, N719, N120);
nor NOR4 (N1609, N1605, N472, N41, N537);
nand NAND2 (N1610, N1603, N1192);
not NOT1 (N1611, N1595);
nand NAND3 (N1612, N1611, N923, N736);
nor NOR2 (N1613, N1612, N229);
nand NAND3 (N1614, N1582, N297, N112);
not NOT1 (N1615, N1609);
nor NOR3 (N1616, N1589, N607, N960);
or OR4 (N1617, N1616, N711, N969, N101);
not NOT1 (N1618, N1607);
and AND3 (N1619, N1604, N905, N382);
nor NOR2 (N1620, N1614, N1110);
nor NOR2 (N1621, N1613, N1260);
not NOT1 (N1622, N1615);
xor XOR2 (N1623, N1617, N634);
nor NOR3 (N1624, N1581, N983, N1017);
nor NOR2 (N1625, N1610, N1196);
not NOT1 (N1626, N1606);
nand NAND4 (N1627, N1622, N805, N543, N297);
xor XOR2 (N1628, N1619, N541);
or OR4 (N1629, N1618, N1431, N584, N551);
not NOT1 (N1630, N1625);
and AND3 (N1631, N1626, N964, N782);
or OR2 (N1632, N1630, N302);
nor NOR3 (N1633, N1631, N729, N1215);
buf BUF1 (N1634, N1633);
and AND4 (N1635, N1634, N419, N1470, N436);
nand NAND3 (N1636, N1608, N133, N1141);
xor XOR2 (N1637, N1629, N314);
xor XOR2 (N1638, N1632, N1392);
nor NOR3 (N1639, N1621, N1479, N507);
buf BUF1 (N1640, N1628);
nand NAND4 (N1641, N1627, N1266, N515, N264);
xor XOR2 (N1642, N1620, N1435);
or OR2 (N1643, N1635, N22);
nor NOR4 (N1644, N1640, N144, N1140, N894);
not NOT1 (N1645, N1642);
nor NOR3 (N1646, N1623, N652, N767);
buf BUF1 (N1647, N1639);
xor XOR2 (N1648, N1645, N1035);
nand NAND2 (N1649, N1624, N737);
nor NOR2 (N1650, N1644, N642);
or OR3 (N1651, N1643, N984, N422);
nor NOR4 (N1652, N1638, N264, N831, N1519);
buf BUF1 (N1653, N1637);
and AND3 (N1654, N1653, N1426, N116);
or OR3 (N1655, N1641, N309, N938);
nand NAND3 (N1656, N1652, N1322, N512);
and AND3 (N1657, N1648, N1162, N1125);
and AND2 (N1658, N1650, N1173);
xor XOR2 (N1659, N1649, N1007);
or OR3 (N1660, N1657, N423, N182);
buf BUF1 (N1661, N1654);
nor NOR3 (N1662, N1646, N834, N1128);
or OR2 (N1663, N1636, N1309);
and AND4 (N1664, N1651, N367, N532, N1388);
nor NOR2 (N1665, N1662, N738);
and AND4 (N1666, N1664, N1576, N121, N1147);
and AND3 (N1667, N1663, N265, N1645);
nand NAND2 (N1668, N1661, N794);
nor NOR2 (N1669, N1668, N475);
or OR3 (N1670, N1647, N1296, N59);
or OR3 (N1671, N1655, N958, N11);
xor XOR2 (N1672, N1665, N1325);
not NOT1 (N1673, N1671);
or OR3 (N1674, N1659, N209, N174);
nand NAND2 (N1675, N1672, N929);
and AND4 (N1676, N1658, N933, N709, N1167);
nand NAND3 (N1677, N1666, N404, N644);
nand NAND2 (N1678, N1676, N785);
nor NOR3 (N1679, N1677, N20, N411);
and AND3 (N1680, N1674, N1343, N1491);
xor XOR2 (N1681, N1656, N564);
nand NAND2 (N1682, N1660, N828);
or OR2 (N1683, N1670, N1639);
buf BUF1 (N1684, N1680);
buf BUF1 (N1685, N1683);
or OR2 (N1686, N1669, N1328);
or OR3 (N1687, N1667, N1517, N1272);
buf BUF1 (N1688, N1682);
nand NAND3 (N1689, N1678, N1181, N659);
not NOT1 (N1690, N1673);
xor XOR2 (N1691, N1684, N1254);
xor XOR2 (N1692, N1681, N1406);
nand NAND4 (N1693, N1679, N994, N814, N47);
nand NAND3 (N1694, N1688, N82, N77);
buf BUF1 (N1695, N1694);
or OR4 (N1696, N1686, N1443, N642, N1504);
nor NOR2 (N1697, N1689, N732);
xor XOR2 (N1698, N1675, N1635);
xor XOR2 (N1699, N1687, N1072);
and AND3 (N1700, N1696, N1175, N265);
and AND4 (N1701, N1693, N1101, N1455, N1463);
and AND4 (N1702, N1690, N136, N410, N1329);
and AND2 (N1703, N1701, N358);
not NOT1 (N1704, N1698);
or OR2 (N1705, N1695, N913);
nor NOR3 (N1706, N1705, N1218, N1491);
or OR4 (N1707, N1700, N1330, N606, N1258);
or OR4 (N1708, N1707, N319, N199, N647);
or OR3 (N1709, N1702, N959, N182);
nand NAND2 (N1710, N1706, N1121);
nor NOR3 (N1711, N1685, N326, N1675);
and AND3 (N1712, N1710, N1607, N1199);
nand NAND4 (N1713, N1704, N1637, N1444, N1215);
and AND3 (N1714, N1713, N307, N391);
buf BUF1 (N1715, N1711);
not NOT1 (N1716, N1703);
xor XOR2 (N1717, N1699, N485);
nor NOR3 (N1718, N1697, N144, N1700);
or OR3 (N1719, N1714, N1194, N1625);
nand NAND4 (N1720, N1715, N1471, N1713, N1624);
or OR4 (N1721, N1718, N617, N1621, N402);
and AND4 (N1722, N1692, N658, N1404, N127);
buf BUF1 (N1723, N1720);
or OR4 (N1724, N1712, N662, N542, N1704);
xor XOR2 (N1725, N1716, N1693);
xor XOR2 (N1726, N1722, N1461);
or OR4 (N1727, N1708, N136, N587, N1659);
or OR2 (N1728, N1724, N72);
and AND4 (N1729, N1717, N1105, N78, N966);
or OR2 (N1730, N1727, N444);
not NOT1 (N1731, N1691);
buf BUF1 (N1732, N1728);
buf BUF1 (N1733, N1709);
not NOT1 (N1734, N1726);
buf BUF1 (N1735, N1725);
and AND3 (N1736, N1719, N1255, N608);
or OR3 (N1737, N1721, N119, N1455);
buf BUF1 (N1738, N1734);
not NOT1 (N1739, N1732);
buf BUF1 (N1740, N1733);
not NOT1 (N1741, N1730);
or OR2 (N1742, N1736, N455);
and AND4 (N1743, N1723, N591, N776, N1256);
or OR4 (N1744, N1729, N505, N218, N122);
nand NAND3 (N1745, N1737, N1202, N81);
and AND4 (N1746, N1741, N354, N642, N1189);
buf BUF1 (N1747, N1745);
xor XOR2 (N1748, N1746, N372);
not NOT1 (N1749, N1738);
not NOT1 (N1750, N1731);
buf BUF1 (N1751, N1748);
nor NOR2 (N1752, N1750, N480);
and AND4 (N1753, N1743, N356, N55, N1563);
and AND4 (N1754, N1735, N1724, N1036, N1587);
nand NAND4 (N1755, N1751, N545, N1710, N239);
buf BUF1 (N1756, N1752);
or OR3 (N1757, N1742, N1542, N964);
not NOT1 (N1758, N1740);
and AND3 (N1759, N1756, N1405, N370);
or OR4 (N1760, N1759, N75, N922, N1027);
xor XOR2 (N1761, N1754, N1191);
or OR4 (N1762, N1755, N476, N447, N891);
not NOT1 (N1763, N1757);
or OR3 (N1764, N1763, N1081, N885);
nand NAND3 (N1765, N1758, N1382, N986);
nand NAND2 (N1766, N1761, N227);
not NOT1 (N1767, N1764);
nor NOR2 (N1768, N1749, N1497);
buf BUF1 (N1769, N1744);
nand NAND4 (N1770, N1769, N781, N570, N1651);
nor NOR4 (N1771, N1770, N769, N1682, N1564);
xor XOR2 (N1772, N1739, N175);
nand NAND4 (N1773, N1765, N1508, N261, N1770);
or OR3 (N1774, N1766, N1092, N355);
buf BUF1 (N1775, N1747);
nand NAND4 (N1776, N1773, N528, N170, N1031);
buf BUF1 (N1777, N1760);
nor NOR3 (N1778, N1753, N1562, N1487);
buf BUF1 (N1779, N1777);
nand NAND3 (N1780, N1779, N15, N909);
nor NOR4 (N1781, N1767, N1066, N658, N1470);
xor XOR2 (N1782, N1771, N250);
and AND3 (N1783, N1776, N1772, N243);
and AND3 (N1784, N903, N1392, N549);
and AND2 (N1785, N1780, N1238);
nand NAND2 (N1786, N1778, N82);
and AND4 (N1787, N1762, N1307, N307, N810);
nor NOR2 (N1788, N1787, N849);
buf BUF1 (N1789, N1768);
nor NOR2 (N1790, N1788, N374);
buf BUF1 (N1791, N1782);
nand NAND3 (N1792, N1781, N421, N23);
or OR4 (N1793, N1774, N254, N527, N527);
nor NOR2 (N1794, N1783, N1339);
nor NOR4 (N1795, N1791, N1449, N1352, N1612);
or OR2 (N1796, N1789, N950);
and AND4 (N1797, N1796, N153, N217, N566);
not NOT1 (N1798, N1795);
buf BUF1 (N1799, N1785);
nand NAND3 (N1800, N1784, N843, N554);
xor XOR2 (N1801, N1797, N155);
and AND2 (N1802, N1800, N194);
nor NOR2 (N1803, N1790, N457);
not NOT1 (N1804, N1803);
buf BUF1 (N1805, N1793);
xor XOR2 (N1806, N1802, N353);
nand NAND4 (N1807, N1794, N120, N1246, N1590);
nor NOR2 (N1808, N1804, N1043);
not NOT1 (N1809, N1805);
nand NAND2 (N1810, N1792, N1211);
or OR3 (N1811, N1806, N1606, N1626);
nand NAND3 (N1812, N1811, N207, N1108);
or OR3 (N1813, N1786, N1463, N833);
xor XOR2 (N1814, N1775, N1011);
xor XOR2 (N1815, N1798, N1711);
nand NAND4 (N1816, N1812, N237, N778, N238);
nor NOR3 (N1817, N1810, N1725, N418);
nand NAND3 (N1818, N1809, N7, N417);
or OR3 (N1819, N1816, N889, N637);
xor XOR2 (N1820, N1808, N1730);
not NOT1 (N1821, N1815);
nand NAND3 (N1822, N1821, N161, N1461);
and AND3 (N1823, N1814, N922, N970);
xor XOR2 (N1824, N1823, N478);
xor XOR2 (N1825, N1820, N622);
nor NOR2 (N1826, N1817, N1159);
buf BUF1 (N1827, N1824);
and AND2 (N1828, N1826, N114);
or OR3 (N1829, N1799, N798, N888);
not NOT1 (N1830, N1801);
or OR4 (N1831, N1819, N306, N1726, N655);
buf BUF1 (N1832, N1825);
xor XOR2 (N1833, N1830, N970);
xor XOR2 (N1834, N1833, N1206);
and AND3 (N1835, N1827, N1168, N1454);
nor NOR4 (N1836, N1828, N1492, N1178, N1557);
xor XOR2 (N1837, N1832, N1357);
buf BUF1 (N1838, N1807);
or OR2 (N1839, N1831, N1070);
nand NAND2 (N1840, N1829, N1376);
or OR3 (N1841, N1836, N936, N1659);
nor NOR4 (N1842, N1840, N1012, N809, N1443);
nand NAND3 (N1843, N1813, N369, N1043);
buf BUF1 (N1844, N1839);
or OR3 (N1845, N1838, N944, N591);
nand NAND2 (N1846, N1845, N1442);
buf BUF1 (N1847, N1843);
or OR3 (N1848, N1841, N150, N922);
or OR3 (N1849, N1848, N1235, N947);
xor XOR2 (N1850, N1849, N366);
xor XOR2 (N1851, N1850, N1127);
xor XOR2 (N1852, N1844, N717);
buf BUF1 (N1853, N1851);
xor XOR2 (N1854, N1842, N586);
nand NAND2 (N1855, N1853, N434);
buf BUF1 (N1856, N1847);
not NOT1 (N1857, N1818);
nor NOR4 (N1858, N1822, N1045, N204, N1492);
xor XOR2 (N1859, N1846, N290);
xor XOR2 (N1860, N1859, N1272);
buf BUF1 (N1861, N1852);
and AND4 (N1862, N1837, N159, N1369, N786);
or OR4 (N1863, N1861, N857, N163, N204);
nor NOR2 (N1864, N1834, N359);
not NOT1 (N1865, N1856);
not NOT1 (N1866, N1865);
buf BUF1 (N1867, N1854);
xor XOR2 (N1868, N1864, N494);
or OR3 (N1869, N1835, N1707, N1534);
nor NOR2 (N1870, N1857, N670);
nor NOR3 (N1871, N1862, N1496, N535);
buf BUF1 (N1872, N1863);
buf BUF1 (N1873, N1855);
nor NOR4 (N1874, N1867, N1062, N1163, N524);
not NOT1 (N1875, N1866);
and AND3 (N1876, N1872, N607, N946);
not NOT1 (N1877, N1871);
and AND2 (N1878, N1868, N386);
xor XOR2 (N1879, N1869, N1812);
and AND2 (N1880, N1870, N1430);
nor NOR3 (N1881, N1875, N1024, N1754);
or OR4 (N1882, N1879, N329, N1549, N950);
nand NAND2 (N1883, N1880, N230);
buf BUF1 (N1884, N1878);
or OR3 (N1885, N1860, N209, N844);
nand NAND2 (N1886, N1858, N1122);
nand NAND4 (N1887, N1876, N736, N845, N91);
not NOT1 (N1888, N1884);
not NOT1 (N1889, N1882);
xor XOR2 (N1890, N1887, N801);
and AND2 (N1891, N1890, N1626);
nand NAND2 (N1892, N1886, N156);
xor XOR2 (N1893, N1892, N1137);
and AND2 (N1894, N1888, N25);
xor XOR2 (N1895, N1889, N1256);
nor NOR2 (N1896, N1895, N931);
nor NOR3 (N1897, N1873, N47, N1185);
and AND3 (N1898, N1894, N1563, N32);
not NOT1 (N1899, N1896);
nor NOR3 (N1900, N1877, N970, N1451);
xor XOR2 (N1901, N1893, N209);
nand NAND3 (N1902, N1874, N1769, N1828);
and AND2 (N1903, N1883, N669);
nor NOR2 (N1904, N1885, N760);
or OR4 (N1905, N1897, N910, N286, N1185);
xor XOR2 (N1906, N1891, N58);
xor XOR2 (N1907, N1881, N1416);
buf BUF1 (N1908, N1901);
xor XOR2 (N1909, N1907, N343);
xor XOR2 (N1910, N1908, N306);
not NOT1 (N1911, N1904);
and AND4 (N1912, N1902, N1558, N204, N713);
or OR4 (N1913, N1905, N219, N763, N538);
nor NOR3 (N1914, N1909, N1823, N254);
and AND3 (N1915, N1900, N1126, N250);
not NOT1 (N1916, N1906);
or OR4 (N1917, N1911, N248, N802, N625);
nor NOR3 (N1918, N1917, N121, N922);
and AND3 (N1919, N1910, N1377, N892);
and AND2 (N1920, N1918, N1608);
not NOT1 (N1921, N1916);
xor XOR2 (N1922, N1920, N1185);
and AND2 (N1923, N1898, N517);
not NOT1 (N1924, N1899);
nand NAND2 (N1925, N1913, N675);
nand NAND4 (N1926, N1924, N695, N93, N1700);
nand NAND4 (N1927, N1912, N575, N280, N331);
and AND3 (N1928, N1926, N1260, N1467);
or OR2 (N1929, N1903, N864);
or OR2 (N1930, N1928, N1613);
buf BUF1 (N1931, N1923);
xor XOR2 (N1932, N1914, N1531);
or OR2 (N1933, N1930, N1226);
or OR2 (N1934, N1929, N1639);
and AND2 (N1935, N1931, N1157);
xor XOR2 (N1936, N1933, N1340);
and AND3 (N1937, N1922, N532, N10);
nor NOR2 (N1938, N1925, N419);
or OR2 (N1939, N1935, N818);
not NOT1 (N1940, N1932);
nor NOR3 (N1941, N1921, N1865, N894);
not NOT1 (N1942, N1940);
nor NOR4 (N1943, N1938, N824, N221, N285);
or OR2 (N1944, N1939, N1194);
not NOT1 (N1945, N1944);
or OR2 (N1946, N1936, N224);
xor XOR2 (N1947, N1945, N424);
xor XOR2 (N1948, N1919, N1723);
xor XOR2 (N1949, N1948, N577);
nor NOR3 (N1950, N1947, N618, N1070);
or OR4 (N1951, N1937, N1564, N927, N355);
nand NAND4 (N1952, N1949, N1570, N1376, N447);
nor NOR4 (N1953, N1934, N1794, N1744, N792);
xor XOR2 (N1954, N1951, N409);
and AND2 (N1955, N1954, N459);
nand NAND3 (N1956, N1953, N1008, N875);
not NOT1 (N1957, N1927);
buf BUF1 (N1958, N1950);
or OR4 (N1959, N1946, N1130, N1655, N30);
or OR4 (N1960, N1955, N703, N1026, N1453);
nor NOR4 (N1961, N1943, N4, N721, N1342);
nor NOR4 (N1962, N1959, N853, N143, N333);
and AND2 (N1963, N1960, N1405);
or OR3 (N1964, N1961, N556, N674);
and AND4 (N1965, N1941, N105, N301, N360);
not NOT1 (N1966, N1963);
xor XOR2 (N1967, N1915, N1339);
not NOT1 (N1968, N1958);
buf BUF1 (N1969, N1962);
xor XOR2 (N1970, N1952, N1241);
and AND2 (N1971, N1967, N428);
nand NAND4 (N1972, N1971, N522, N841, N1909);
nand NAND4 (N1973, N1969, N683, N957, N1601);
and AND2 (N1974, N1966, N1137);
buf BUF1 (N1975, N1957);
nand NAND4 (N1976, N1972, N1540, N612, N1349);
or OR2 (N1977, N1975, N1591);
xor XOR2 (N1978, N1942, N1463);
and AND4 (N1979, N1973, N224, N671, N1437);
or OR3 (N1980, N1976, N1838, N1787);
not NOT1 (N1981, N1965);
nand NAND4 (N1982, N1981, N1734, N973, N54);
buf BUF1 (N1983, N1982);
or OR4 (N1984, N1978, N602, N1362, N1282);
and AND4 (N1985, N1983, N266, N1453, N503);
and AND4 (N1986, N1979, N78, N604, N295);
and AND3 (N1987, N1984, N1531, N394);
xor XOR2 (N1988, N1986, N686);
buf BUF1 (N1989, N1974);
nor NOR2 (N1990, N1980, N409);
or OR4 (N1991, N1956, N617, N616, N1232);
nor NOR4 (N1992, N1988, N1757, N1681, N1500);
or OR2 (N1993, N1964, N1003);
nand NAND4 (N1994, N1989, N1525, N1703, N306);
not NOT1 (N1995, N1990);
or OR4 (N1996, N1991, N868, N923, N761);
nand NAND4 (N1997, N1987, N383, N521, N849);
or OR2 (N1998, N1968, N946);
or OR3 (N1999, N1998, N1841, N1181);
xor XOR2 (N2000, N1996, N139);
and AND2 (N2001, N1970, N676);
buf BUF1 (N2002, N1992);
nand NAND3 (N2003, N1999, N1203, N374);
not NOT1 (N2004, N2001);
buf BUF1 (N2005, N1993);
or OR4 (N2006, N2002, N1816, N874, N301);
or OR2 (N2007, N2000, N1067);
not NOT1 (N2008, N2004);
and AND4 (N2009, N1994, N918, N314, N1596);
or OR4 (N2010, N2003, N1374, N1963, N1795);
xor XOR2 (N2011, N2007, N1043);
and AND3 (N2012, N1977, N944, N847);
nand NAND3 (N2013, N2012, N1523, N873);
not NOT1 (N2014, N2013);
xor XOR2 (N2015, N1997, N1519);
and AND4 (N2016, N2011, N327, N166, N883);
buf BUF1 (N2017, N1985);
or OR3 (N2018, N2010, N1102, N876);
buf BUF1 (N2019, N2005);
nand NAND3 (N2020, N1995, N1605, N1671);
not NOT1 (N2021, N2009);
nand NAND4 (N2022, N2016, N1796, N1448, N1117);
or OR2 (N2023, N2018, N1621);
nand NAND2 (N2024, N2015, N1143);
xor XOR2 (N2025, N2008, N551);
and AND2 (N2026, N2024, N104);
or OR3 (N2027, N2019, N1406, N282);
nand NAND4 (N2028, N2022, N1146, N1518, N1949);
buf BUF1 (N2029, N2026);
xor XOR2 (N2030, N2023, N1704);
and AND4 (N2031, N2029, N1851, N1032, N1374);
nand NAND4 (N2032, N2027, N1797, N1985, N671);
or OR2 (N2033, N2020, N136);
nand NAND4 (N2034, N2032, N222, N566, N1900);
buf BUF1 (N2035, N2028);
and AND3 (N2036, N2025, N1585, N591);
buf BUF1 (N2037, N2036);
xor XOR2 (N2038, N2030, N1798);
or OR4 (N2039, N2021, N119, N1367, N985);
not NOT1 (N2040, N2031);
and AND4 (N2041, N2033, N712, N994, N1585);
nand NAND4 (N2042, N2040, N1560, N1991, N1779);
not NOT1 (N2043, N2042);
not NOT1 (N2044, N2006);
nand NAND2 (N2045, N2037, N239);
buf BUF1 (N2046, N2044);
buf BUF1 (N2047, N2034);
nor NOR3 (N2048, N2035, N75, N756);
nor NOR3 (N2049, N2039, N531, N912);
not NOT1 (N2050, N2045);
nand NAND4 (N2051, N2017, N2018, N1186, N1076);
buf BUF1 (N2052, N2046);
not NOT1 (N2053, N2014);
or OR2 (N2054, N2050, N4);
or OR2 (N2055, N2047, N1516);
nor NOR2 (N2056, N2049, N310);
or OR2 (N2057, N2051, N254);
nor NOR4 (N2058, N2043, N1821, N1729, N566);
not NOT1 (N2059, N2056);
nand NAND2 (N2060, N2054, N1943);
or OR4 (N2061, N2052, N503, N1627, N1151);
buf BUF1 (N2062, N2058);
nand NAND3 (N2063, N2057, N160, N1426);
not NOT1 (N2064, N2061);
or OR3 (N2065, N2041, N1069, N25);
and AND4 (N2066, N2065, N1810, N647, N1729);
or OR4 (N2067, N2053, N1961, N193, N358);
or OR4 (N2068, N2064, N933, N551, N471);
nor NOR4 (N2069, N2055, N1182, N234, N145);
nand NAND3 (N2070, N2048, N916, N1152);
not NOT1 (N2071, N2060);
nand NAND3 (N2072, N2062, N2003, N723);
not NOT1 (N2073, N2069);
not NOT1 (N2074, N2070);
nand NAND4 (N2075, N2063, N373, N1936, N415);
buf BUF1 (N2076, N2072);
not NOT1 (N2077, N2059);
or OR3 (N2078, N2067, N553, N420);
or OR2 (N2079, N2071, N105);
xor XOR2 (N2080, N2079, N260);
nor NOR3 (N2081, N2038, N1083, N167);
nor NOR2 (N2082, N2073, N1878);
nand NAND3 (N2083, N2076, N863, N1864);
nand NAND2 (N2084, N2074, N365);
nor NOR4 (N2085, N2083, N262, N407, N189);
or OR4 (N2086, N2081, N1245, N1391, N1453);
xor XOR2 (N2087, N2084, N1371);
xor XOR2 (N2088, N2077, N1289);
xor XOR2 (N2089, N2082, N1449);
nor NOR4 (N2090, N2075, N391, N1990, N1460);
xor XOR2 (N2091, N2078, N2031);
xor XOR2 (N2092, N2089, N1218);
xor XOR2 (N2093, N2086, N1276);
and AND3 (N2094, N2091, N1043, N1805);
not NOT1 (N2095, N2092);
not NOT1 (N2096, N2088);
and AND3 (N2097, N2096, N384, N1792);
nor NOR4 (N2098, N2087, N1319, N1453, N253);
nand NAND4 (N2099, N2093, N355, N998, N1112);
or OR4 (N2100, N2098, N641, N736, N1433);
not NOT1 (N2101, N2100);
nand NAND4 (N2102, N2099, N547, N354, N264);
buf BUF1 (N2103, N2066);
buf BUF1 (N2104, N2103);
buf BUF1 (N2105, N2097);
and AND3 (N2106, N2080, N1819, N1265);
buf BUF1 (N2107, N2105);
nand NAND4 (N2108, N2085, N1667, N1426, N165);
not NOT1 (N2109, N2094);
xor XOR2 (N2110, N2102, N238);
nor NOR2 (N2111, N2110, N335);
buf BUF1 (N2112, N2104);
nor NOR4 (N2113, N2112, N1501, N516, N991);
not NOT1 (N2114, N2095);
nor NOR2 (N2115, N2114, N458);
nor NOR4 (N2116, N2109, N1230, N1288, N1145);
buf BUF1 (N2117, N2115);
buf BUF1 (N2118, N2068);
or OR4 (N2119, N2090, N1010, N312, N184);
or OR2 (N2120, N2101, N1554);
or OR4 (N2121, N2111, N797, N1723, N1751);
and AND2 (N2122, N2113, N1512);
buf BUF1 (N2123, N2106);
or OR2 (N2124, N2123, N977);
xor XOR2 (N2125, N2116, N985);
and AND4 (N2126, N2119, N575, N970, N1135);
nor NOR4 (N2127, N2124, N1929, N1831, N1916);
nor NOR3 (N2128, N2117, N1523, N1729);
xor XOR2 (N2129, N2120, N1521);
nand NAND3 (N2130, N2129, N161, N2113);
buf BUF1 (N2131, N2130);
nor NOR2 (N2132, N2118, N1038);
and AND4 (N2133, N2126, N563, N1253, N365);
xor XOR2 (N2134, N2128, N820);
xor XOR2 (N2135, N2108, N1790);
xor XOR2 (N2136, N2125, N635);
nor NOR4 (N2137, N2135, N687, N2111, N544);
nand NAND2 (N2138, N2121, N1146);
or OR4 (N2139, N2107, N266, N1008, N620);
and AND3 (N2140, N2122, N1134, N1351);
not NOT1 (N2141, N2139);
nand NAND2 (N2142, N2140, N1194);
nor NOR4 (N2143, N2131, N214, N1643, N225);
xor XOR2 (N2144, N2137, N569);
or OR2 (N2145, N2143, N390);
xor XOR2 (N2146, N2127, N1097);
buf BUF1 (N2147, N2133);
not NOT1 (N2148, N2145);
or OR2 (N2149, N2132, N1155);
or OR3 (N2150, N2134, N1075, N754);
not NOT1 (N2151, N2146);
nor NOR4 (N2152, N2138, N921, N2125, N1492);
buf BUF1 (N2153, N2147);
buf BUF1 (N2154, N2153);
or OR2 (N2155, N2151, N1859);
and AND4 (N2156, N2150, N538, N1885, N464);
not NOT1 (N2157, N2136);
not NOT1 (N2158, N2148);
not NOT1 (N2159, N2156);
buf BUF1 (N2160, N2157);
nand NAND4 (N2161, N2159, N1875, N772, N1733);
nand NAND3 (N2162, N2142, N1334, N1191);
and AND4 (N2163, N2144, N967, N1907, N1768);
xor XOR2 (N2164, N2149, N781);
xor XOR2 (N2165, N2160, N1781);
buf BUF1 (N2166, N2161);
and AND2 (N2167, N2164, N1548);
xor XOR2 (N2168, N2165, N688);
buf BUF1 (N2169, N2167);
nand NAND4 (N2170, N2169, N1671, N712, N1746);
nor NOR2 (N2171, N2170, N1528);
and AND4 (N2172, N2154, N1753, N1773, N1118);
buf BUF1 (N2173, N2141);
buf BUF1 (N2174, N2158);
xor XOR2 (N2175, N2155, N71);
xor XOR2 (N2176, N2162, N370);
and AND4 (N2177, N2168, N424, N690, N1910);
nand NAND4 (N2178, N2173, N600, N1534, N869);
xor XOR2 (N2179, N2176, N1980);
or OR4 (N2180, N2179, N287, N632, N73);
and AND2 (N2181, N2178, N55);
nand NAND4 (N2182, N2172, N1534, N914, N1513);
nand NAND4 (N2183, N2177, N690, N1811, N1252);
and AND2 (N2184, N2171, N1034);
buf BUF1 (N2185, N2180);
or OR3 (N2186, N2174, N1723, N1977);
not NOT1 (N2187, N2186);
nand NAND3 (N2188, N2184, N1859, N764);
nand NAND4 (N2189, N2166, N53, N1014, N1254);
and AND2 (N2190, N2175, N1762);
xor XOR2 (N2191, N2181, N1574);
xor XOR2 (N2192, N2188, N1019);
buf BUF1 (N2193, N2163);
nand NAND3 (N2194, N2192, N1502, N343);
and AND4 (N2195, N2191, N1685, N1621, N1163);
or OR3 (N2196, N2194, N737, N1406);
or OR4 (N2197, N2187, N835, N491, N342);
buf BUF1 (N2198, N2183);
nor NOR3 (N2199, N2182, N2014, N1898);
and AND2 (N2200, N2197, N1216);
not NOT1 (N2201, N2195);
or OR4 (N2202, N2189, N926, N1828, N1400);
not NOT1 (N2203, N2202);
not NOT1 (N2204, N2198);
and AND4 (N2205, N2193, N55, N1278, N412);
nor NOR4 (N2206, N2200, N1034, N88, N110);
or OR3 (N2207, N2196, N1116, N1835);
xor XOR2 (N2208, N2152, N1798);
and AND3 (N2209, N2206, N1231, N1100);
buf BUF1 (N2210, N2199);
xor XOR2 (N2211, N2205, N2044);
nor NOR3 (N2212, N2190, N1426, N1738);
or OR3 (N2213, N2204, N1062, N582);
not NOT1 (N2214, N2208);
buf BUF1 (N2215, N2210);
and AND3 (N2216, N2215, N245, N334);
or OR4 (N2217, N2216, N744, N1590, N837);
or OR4 (N2218, N2214, N720, N1555, N1760);
nand NAND4 (N2219, N2201, N168, N574, N1693);
xor XOR2 (N2220, N2203, N828);
or OR4 (N2221, N2219, N8, N171, N1634);
nand NAND2 (N2222, N2217, N1112);
xor XOR2 (N2223, N2209, N1417);
nor NOR2 (N2224, N2185, N1954);
nor NOR3 (N2225, N2224, N720, N1166);
nand NAND3 (N2226, N2213, N1262, N2098);
or OR2 (N2227, N2225, N1459);
not NOT1 (N2228, N2223);
nand NAND4 (N2229, N2222, N1542, N1117, N1055);
buf BUF1 (N2230, N2220);
xor XOR2 (N2231, N2218, N1781);
and AND2 (N2232, N2227, N229);
nand NAND3 (N2233, N2211, N1079, N1019);
nand NAND3 (N2234, N2230, N1834, N475);
buf BUF1 (N2235, N2221);
and AND3 (N2236, N2232, N764, N1943);
not NOT1 (N2237, N2236);
nand NAND4 (N2238, N2234, N1513, N858, N1352);
nand NAND3 (N2239, N2235, N289, N1006);
not NOT1 (N2240, N2207);
not NOT1 (N2241, N2228);
and AND3 (N2242, N2229, N917, N1079);
buf BUF1 (N2243, N2240);
or OR2 (N2244, N2239, N1128);
nor NOR3 (N2245, N2243, N1001, N2216);
and AND2 (N2246, N2231, N1155);
nor NOR3 (N2247, N2245, N1123, N1867);
or OR2 (N2248, N2246, N1198);
not NOT1 (N2249, N2241);
not NOT1 (N2250, N2248);
or OR2 (N2251, N2237, N1417);
nand NAND3 (N2252, N2226, N1842, N1973);
and AND2 (N2253, N2251, N1664);
buf BUF1 (N2254, N2252);
or OR3 (N2255, N2238, N2194, N1494);
xor XOR2 (N2256, N2250, N246);
or OR3 (N2257, N2256, N1744, N1290);
nor NOR4 (N2258, N2244, N897, N312, N323);
and AND4 (N2259, N2247, N1889, N550, N120);
nor NOR4 (N2260, N2249, N1611, N1447, N1671);
buf BUF1 (N2261, N2257);
nand NAND2 (N2262, N2242, N114);
or OR2 (N2263, N2260, N1863);
xor XOR2 (N2264, N2261, N230);
xor XOR2 (N2265, N2259, N1277);
or OR2 (N2266, N2254, N1197);
not NOT1 (N2267, N2233);
nor NOR4 (N2268, N2255, N2133, N1951, N2166);
nor NOR2 (N2269, N2258, N1146);
xor XOR2 (N2270, N2263, N969);
nor NOR2 (N2271, N2262, N612);
not NOT1 (N2272, N2270);
xor XOR2 (N2273, N2271, N753);
nor NOR3 (N2274, N2212, N1419, N773);
not NOT1 (N2275, N2253);
and AND3 (N2276, N2266, N363, N672);
buf BUF1 (N2277, N2267);
or OR4 (N2278, N2275, N423, N487, N2221);
nand NAND3 (N2279, N2276, N1921, N395);
nand NAND2 (N2280, N2265, N1648);
xor XOR2 (N2281, N2277, N2127);
or OR2 (N2282, N2280, N1785);
buf BUF1 (N2283, N2279);
not NOT1 (N2284, N2272);
and AND4 (N2285, N2281, N615, N757, N1176);
nor NOR4 (N2286, N2278, N876, N2253, N818);
and AND4 (N2287, N2273, N1649, N1781, N136);
nor NOR4 (N2288, N2285, N2268, N2179, N195);
and AND3 (N2289, N1074, N226, N1066);
not NOT1 (N2290, N2283);
xor XOR2 (N2291, N2264, N2220);
nor NOR4 (N2292, N2286, N817, N1725, N312);
or OR4 (N2293, N2289, N1443, N940, N717);
not NOT1 (N2294, N2284);
nand NAND3 (N2295, N2287, N1074, N1454);
buf BUF1 (N2296, N2269);
and AND4 (N2297, N2294, N1948, N981, N1437);
not NOT1 (N2298, N2292);
not NOT1 (N2299, N2293);
nand NAND2 (N2300, N2299, N1643);
nor NOR4 (N2301, N2296, N1487, N1626, N1129);
or OR2 (N2302, N2288, N1778);
and AND3 (N2303, N2274, N215, N2045);
buf BUF1 (N2304, N2295);
or OR4 (N2305, N2290, N285, N896, N1512);
xor XOR2 (N2306, N2297, N1611);
not NOT1 (N2307, N2303);
or OR2 (N2308, N2302, N471);
nand NAND4 (N2309, N2306, N2169, N1019, N2088);
nor NOR2 (N2310, N2282, N394);
not NOT1 (N2311, N2304);
nand NAND3 (N2312, N2308, N1215, N1460);
buf BUF1 (N2313, N2291);
nand NAND2 (N2314, N2307, N1209);
nor NOR3 (N2315, N2314, N1769, N1656);
xor XOR2 (N2316, N2313, N618);
nor NOR3 (N2317, N2300, N2144, N1981);
or OR3 (N2318, N2317, N70, N1260);
nor NOR2 (N2319, N2318, N950);
not NOT1 (N2320, N2301);
xor XOR2 (N2321, N2315, N1747);
and AND3 (N2322, N2320, N1962, N2081);
not NOT1 (N2323, N2310);
not NOT1 (N2324, N2316);
and AND4 (N2325, N2324, N1993, N1169, N953);
nand NAND2 (N2326, N2321, N1598);
or OR3 (N2327, N2325, N271, N1105);
and AND3 (N2328, N2319, N359, N1040);
and AND4 (N2329, N2305, N1418, N395, N2201);
xor XOR2 (N2330, N2322, N1927);
xor XOR2 (N2331, N2328, N1602);
or OR2 (N2332, N2326, N1963);
and AND4 (N2333, N2312, N1672, N1680, N1496);
nand NAND3 (N2334, N2311, N2292, N258);
nor NOR3 (N2335, N2327, N649, N691);
nor NOR4 (N2336, N2309, N2103, N2077, N867);
or OR4 (N2337, N2335, N1173, N757, N1369);
buf BUF1 (N2338, N2329);
xor XOR2 (N2339, N2337, N1974);
buf BUF1 (N2340, N2331);
nor NOR3 (N2341, N2339, N331, N2242);
or OR3 (N2342, N2323, N77, N30);
xor XOR2 (N2343, N2332, N2088);
buf BUF1 (N2344, N2342);
or OR3 (N2345, N2298, N2146, N1635);
xor XOR2 (N2346, N2343, N1401);
buf BUF1 (N2347, N2340);
buf BUF1 (N2348, N2336);
xor XOR2 (N2349, N2348, N948);
and AND2 (N2350, N2338, N1586);
not NOT1 (N2351, N2350);
not NOT1 (N2352, N2341);
nand NAND3 (N2353, N2330, N668, N2105);
nand NAND4 (N2354, N2334, N1784, N717, N2308);
xor XOR2 (N2355, N2353, N1451);
buf BUF1 (N2356, N2346);
nor NOR3 (N2357, N2333, N828, N973);
or OR2 (N2358, N2352, N1106);
nand NAND4 (N2359, N2349, N91, N472, N1711);
and AND2 (N2360, N2358, N483);
and AND2 (N2361, N2347, N825);
buf BUF1 (N2362, N2345);
buf BUF1 (N2363, N2356);
or OR4 (N2364, N2344, N1151, N324, N2153);
or OR3 (N2365, N2361, N2268, N1127);
nor NOR4 (N2366, N2355, N1444, N953, N389);
buf BUF1 (N2367, N2351);
xor XOR2 (N2368, N2360, N1529);
not NOT1 (N2369, N2357);
nor NOR2 (N2370, N2369, N363);
nand NAND2 (N2371, N2370, N2335);
not NOT1 (N2372, N2366);
nand NAND4 (N2373, N2368, N771, N1706, N730);
not NOT1 (N2374, N2359);
xor XOR2 (N2375, N2373, N130);
or OR4 (N2376, N2362, N609, N1119, N832);
or OR4 (N2377, N2367, N1185, N582, N678);
or OR4 (N2378, N2375, N1816, N1472, N1051);
or OR2 (N2379, N2364, N1003);
xor XOR2 (N2380, N2378, N48);
or OR2 (N2381, N2376, N1849);
xor XOR2 (N2382, N2354, N976);
not NOT1 (N2383, N2365);
and AND3 (N2384, N2381, N1116, N1251);
buf BUF1 (N2385, N2383);
buf BUF1 (N2386, N2377);
or OR4 (N2387, N2384, N716, N713, N1107);
not NOT1 (N2388, N2379);
or OR4 (N2389, N2372, N391, N80, N362);
and AND4 (N2390, N2382, N1580, N1839, N1831);
nor NOR4 (N2391, N2390, N2186, N1557, N744);
xor XOR2 (N2392, N2386, N2245);
and AND4 (N2393, N2385, N1603, N1000, N967);
or OR3 (N2394, N2363, N760, N2253);
nor NOR4 (N2395, N2388, N537, N1237, N1063);
nor NOR4 (N2396, N2374, N622, N1350, N2306);
buf BUF1 (N2397, N2392);
xor XOR2 (N2398, N2395, N1055);
and AND2 (N2399, N2397, N490);
and AND2 (N2400, N2389, N1157);
nand NAND2 (N2401, N2391, N132);
and AND3 (N2402, N2396, N2099, N802);
nor NOR3 (N2403, N2387, N1395, N1621);
not NOT1 (N2404, N2399);
and AND2 (N2405, N2394, N2092);
nand NAND4 (N2406, N2403, N979, N1351, N196);
not NOT1 (N2407, N2401);
nor NOR4 (N2408, N2380, N2211, N1846, N1679);
or OR4 (N2409, N2402, N994, N681, N2051);
and AND3 (N2410, N2409, N1602, N2356);
and AND4 (N2411, N2410, N42, N694, N960);
buf BUF1 (N2412, N2405);
buf BUF1 (N2413, N2400);
not NOT1 (N2414, N2413);
and AND2 (N2415, N2407, N175);
buf BUF1 (N2416, N2411);
nor NOR2 (N2417, N2393, N1680);
or OR4 (N2418, N2371, N1852, N1269, N631);
buf BUF1 (N2419, N2414);
nand NAND3 (N2420, N2415, N2240, N1797);
xor XOR2 (N2421, N2412, N2018);
nand NAND4 (N2422, N2416, N1959, N1626, N487);
xor XOR2 (N2423, N2404, N1584);
xor XOR2 (N2424, N2406, N900);
nand NAND3 (N2425, N2422, N538, N491);
buf BUF1 (N2426, N2420);
or OR3 (N2427, N2417, N885, N2394);
and AND3 (N2428, N2426, N1691, N2290);
xor XOR2 (N2429, N2398, N1062);
not NOT1 (N2430, N2418);
nand NAND4 (N2431, N2408, N1095, N60, N2252);
buf BUF1 (N2432, N2431);
or OR3 (N2433, N2430, N1726, N1334);
xor XOR2 (N2434, N2425, N1823);
xor XOR2 (N2435, N2427, N2049);
nand NAND3 (N2436, N2434, N1421, N1834);
nand NAND3 (N2437, N2423, N1351, N2080);
xor XOR2 (N2438, N2432, N2296);
nor NOR2 (N2439, N2433, N2050);
not NOT1 (N2440, N2428);
buf BUF1 (N2441, N2436);
nor NOR2 (N2442, N2424, N1048);
xor XOR2 (N2443, N2429, N217);
and AND2 (N2444, N2442, N1664);
xor XOR2 (N2445, N2437, N1047);
nor NOR3 (N2446, N2440, N1387, N1999);
not NOT1 (N2447, N2438);
or OR4 (N2448, N2419, N596, N1462, N1259);
nor NOR2 (N2449, N2435, N2300);
nand NAND2 (N2450, N2448, N682);
xor XOR2 (N2451, N2439, N1747);
nand NAND2 (N2452, N2421, N950);
not NOT1 (N2453, N2451);
nand NAND4 (N2454, N2441, N1043, N718, N766);
nand NAND4 (N2455, N2444, N502, N246, N1863);
nor NOR3 (N2456, N2452, N1411, N2012);
not NOT1 (N2457, N2456);
nor NOR3 (N2458, N2449, N1114, N350);
buf BUF1 (N2459, N2450);
nand NAND3 (N2460, N2443, N1615, N1437);
nand NAND2 (N2461, N2460, N27);
or OR4 (N2462, N2446, N1666, N886, N808);
and AND3 (N2463, N2445, N1319, N1907);
nand NAND3 (N2464, N2455, N245, N177);
or OR2 (N2465, N2458, N650);
nor NOR2 (N2466, N2463, N1920);
nor NOR4 (N2467, N2461, N1896, N2461, N1015);
and AND3 (N2468, N2454, N548, N1841);
and AND4 (N2469, N2453, N430, N789, N675);
xor XOR2 (N2470, N2467, N868);
buf BUF1 (N2471, N2470);
xor XOR2 (N2472, N2447, N767);
xor XOR2 (N2473, N2459, N1834);
nand NAND3 (N2474, N2457, N1584, N1721);
nand NAND3 (N2475, N2468, N2465, N1761);
buf BUF1 (N2476, N1901);
or OR4 (N2477, N2469, N510, N1332, N1819);
xor XOR2 (N2478, N2472, N707);
not NOT1 (N2479, N2474);
nand NAND4 (N2480, N2478, N1121, N2015, N336);
nand NAND2 (N2481, N2464, N1502);
or OR2 (N2482, N2479, N238);
xor XOR2 (N2483, N2473, N2315);
and AND2 (N2484, N2462, N2160);
xor XOR2 (N2485, N2484, N1109);
and AND3 (N2486, N2480, N1997, N2106);
not NOT1 (N2487, N2485);
not NOT1 (N2488, N2487);
not NOT1 (N2489, N2471);
xor XOR2 (N2490, N2481, N171);
xor XOR2 (N2491, N2482, N802);
and AND3 (N2492, N2476, N2463, N1574);
nor NOR4 (N2493, N2475, N988, N1469, N1527);
nand NAND2 (N2494, N2488, N2150);
buf BUF1 (N2495, N2483);
buf BUF1 (N2496, N2492);
xor XOR2 (N2497, N2493, N1766);
and AND2 (N2498, N2496, N2229);
not NOT1 (N2499, N2489);
not NOT1 (N2500, N2491);
not NOT1 (N2501, N2500);
xor XOR2 (N2502, N2486, N107);
xor XOR2 (N2503, N2490, N96);
buf BUF1 (N2504, N2466);
nor NOR4 (N2505, N2477, N1664, N1062, N1470);
xor XOR2 (N2506, N2497, N1040);
and AND4 (N2507, N2504, N185, N222, N1749);
nand NAND4 (N2508, N2494, N998, N1589, N1517);
xor XOR2 (N2509, N2501, N708);
buf BUF1 (N2510, N2502);
or OR2 (N2511, N2495, N2439);
and AND2 (N2512, N2509, N1242);
nor NOR3 (N2513, N2510, N1970, N2187);
nor NOR4 (N2514, N2503, N446, N1845, N1021);
xor XOR2 (N2515, N2506, N1647);
not NOT1 (N2516, N2498);
or OR4 (N2517, N2508, N2223, N1936, N975);
buf BUF1 (N2518, N2516);
buf BUF1 (N2519, N2514);
xor XOR2 (N2520, N2515, N130);
not NOT1 (N2521, N2520);
not NOT1 (N2522, N2505);
xor XOR2 (N2523, N2511, N1504);
and AND3 (N2524, N2521, N633, N2187);
and AND4 (N2525, N2512, N313, N363, N546);
nand NAND3 (N2526, N2518, N2057, N1533);
not NOT1 (N2527, N2517);
not NOT1 (N2528, N2513);
nor NOR2 (N2529, N2499, N1368);
nor NOR2 (N2530, N2526, N1625);
buf BUF1 (N2531, N2530);
xor XOR2 (N2532, N2507, N54);
not NOT1 (N2533, N2522);
nor NOR3 (N2534, N2524, N1665, N2405);
nand NAND3 (N2535, N2528, N1812, N1451);
not NOT1 (N2536, N2523);
nor NOR4 (N2537, N2519, N512, N232, N112);
nor NOR2 (N2538, N2529, N208);
nor NOR4 (N2539, N2537, N630, N1695, N1522);
and AND4 (N2540, N2539, N292, N1085, N18);
nand NAND3 (N2541, N2536, N2082, N1661);
not NOT1 (N2542, N2533);
nor NOR2 (N2543, N2525, N1910);
nor NOR4 (N2544, N2543, N2269, N2452, N496);
not NOT1 (N2545, N2535);
nor NOR4 (N2546, N2534, N530, N745, N238);
or OR4 (N2547, N2544, N84, N2070, N1639);
or OR2 (N2548, N2532, N2326);
nor NOR4 (N2549, N2542, N822, N1478, N305);
xor XOR2 (N2550, N2548, N38);
and AND2 (N2551, N2541, N216);
nor NOR3 (N2552, N2550, N1647, N2157);
and AND3 (N2553, N2549, N1287, N1126);
not NOT1 (N2554, N2552);
nand NAND2 (N2555, N2545, N2265);
buf BUF1 (N2556, N2538);
not NOT1 (N2557, N2546);
not NOT1 (N2558, N2557);
buf BUF1 (N2559, N2551);
nand NAND2 (N2560, N2553, N430);
and AND3 (N2561, N2558, N435, N929);
nand NAND3 (N2562, N2554, N501, N1463);
or OR3 (N2563, N2562, N2558, N1016);
buf BUF1 (N2564, N2563);
nor NOR2 (N2565, N2559, N150);
nand NAND4 (N2566, N2564, N1950, N2100, N2081);
nand NAND4 (N2567, N2547, N1102, N453, N1265);
buf BUF1 (N2568, N2560);
or OR3 (N2569, N2568, N1481, N841);
or OR3 (N2570, N2567, N710, N693);
or OR4 (N2571, N2555, N682, N659, N2325);
buf BUF1 (N2572, N2570);
nand NAND2 (N2573, N2527, N370);
not NOT1 (N2574, N2569);
buf BUF1 (N2575, N2573);
nand NAND4 (N2576, N2565, N428, N2313, N153);
or OR4 (N2577, N2572, N720, N1962, N151);
nand NAND3 (N2578, N2571, N2327, N2061);
nor NOR2 (N2579, N2575, N210);
buf BUF1 (N2580, N2556);
and AND2 (N2581, N2531, N565);
nor NOR4 (N2582, N2577, N1141, N1920, N73);
or OR3 (N2583, N2582, N1241, N838);
buf BUF1 (N2584, N2583);
or OR2 (N2585, N2574, N1034);
or OR4 (N2586, N2580, N1935, N1291, N1587);
or OR3 (N2587, N2586, N1439, N726);
nand NAND2 (N2588, N2587, N221);
not NOT1 (N2589, N2581);
xor XOR2 (N2590, N2561, N2429);
and AND4 (N2591, N2585, N2575, N877, N718);
buf BUF1 (N2592, N2589);
xor XOR2 (N2593, N2588, N2144);
nand NAND4 (N2594, N2579, N1539, N1461, N2437);
xor XOR2 (N2595, N2578, N112);
and AND3 (N2596, N2594, N1745, N1678);
xor XOR2 (N2597, N2576, N220);
buf BUF1 (N2598, N2596);
and AND4 (N2599, N2591, N1063, N146, N1804);
buf BUF1 (N2600, N2590);
nor NOR2 (N2601, N2595, N2443);
and AND2 (N2602, N2592, N1899);
and AND2 (N2603, N2598, N274);
nand NAND4 (N2604, N2584, N1298, N1761, N1330);
or OR2 (N2605, N2540, N1660);
xor XOR2 (N2606, N2603, N1349);
nand NAND2 (N2607, N2597, N452);
and AND2 (N2608, N2605, N402);
nor NOR3 (N2609, N2602, N2320, N2200);
nand NAND3 (N2610, N2600, N232, N699);
nand NAND4 (N2611, N2609, N1314, N1437, N703);
xor XOR2 (N2612, N2610, N721);
and AND2 (N2613, N2599, N417);
not NOT1 (N2614, N2606);
buf BUF1 (N2615, N2601);
nor NOR3 (N2616, N2604, N2438, N1765);
xor XOR2 (N2617, N2613, N2364);
buf BUF1 (N2618, N2612);
buf BUF1 (N2619, N2617);
buf BUF1 (N2620, N2566);
nand NAND2 (N2621, N2619, N1966);
and AND4 (N2622, N2593, N2437, N2439, N1893);
and AND3 (N2623, N2611, N1043, N2337);
nor NOR4 (N2624, N2621, N1707, N1872, N1620);
nor NOR4 (N2625, N2624, N341, N602, N1601);
nor NOR4 (N2626, N2618, N1333, N1961, N1411);
nor NOR4 (N2627, N2620, N1597, N1829, N578);
xor XOR2 (N2628, N2626, N1049);
and AND2 (N2629, N2607, N208);
xor XOR2 (N2630, N2616, N1021);
xor XOR2 (N2631, N2615, N875);
not NOT1 (N2632, N2608);
or OR2 (N2633, N2630, N1552);
and AND4 (N2634, N2631, N1361, N762, N2090);
xor XOR2 (N2635, N2634, N1339);
nand NAND2 (N2636, N2628, N16);
xor XOR2 (N2637, N2614, N2245);
buf BUF1 (N2638, N2629);
nor NOR2 (N2639, N2622, N2215);
nor NOR3 (N2640, N2627, N2226, N1462);
xor XOR2 (N2641, N2640, N1745);
nor NOR3 (N2642, N2636, N876, N497);
nor NOR4 (N2643, N2639, N2202, N561, N205);
nor NOR2 (N2644, N2637, N39);
or OR3 (N2645, N2638, N1380, N2395);
xor XOR2 (N2646, N2625, N2105);
xor XOR2 (N2647, N2646, N1333);
or OR2 (N2648, N2623, N715);
or OR3 (N2649, N2645, N2175, N1435);
or OR3 (N2650, N2641, N749, N523);
not NOT1 (N2651, N2650);
or OR3 (N2652, N2642, N470, N990);
not NOT1 (N2653, N2648);
nand NAND3 (N2654, N2632, N409, N407);
buf BUF1 (N2655, N2643);
nor NOR4 (N2656, N2652, N212, N1751, N1801);
and AND2 (N2657, N2656, N2120);
nor NOR3 (N2658, N2651, N1343, N989);
buf BUF1 (N2659, N2644);
and AND2 (N2660, N2658, N385);
nor NOR4 (N2661, N2653, N2339, N439, N2626);
nor NOR2 (N2662, N2660, N620);
nand NAND3 (N2663, N2633, N264, N660);
not NOT1 (N2664, N2659);
or OR3 (N2665, N2635, N1889, N732);
buf BUF1 (N2666, N2657);
nand NAND3 (N2667, N2665, N264, N434);
buf BUF1 (N2668, N2655);
or OR3 (N2669, N2654, N1945, N735);
and AND2 (N2670, N2647, N633);
buf BUF1 (N2671, N2669);
nand NAND2 (N2672, N2667, N311);
xor XOR2 (N2673, N2670, N2420);
nand NAND2 (N2674, N2666, N2294);
not NOT1 (N2675, N2671);
buf BUF1 (N2676, N2668);
xor XOR2 (N2677, N2675, N731);
xor XOR2 (N2678, N2673, N1241);
nand NAND3 (N2679, N2662, N2192, N2281);
xor XOR2 (N2680, N2663, N784);
not NOT1 (N2681, N2680);
nor NOR3 (N2682, N2677, N506, N531);
or OR2 (N2683, N2682, N2107);
buf BUF1 (N2684, N2678);
or OR3 (N2685, N2684, N827, N1975);
or OR3 (N2686, N2664, N992, N121);
nand NAND3 (N2687, N2679, N998, N1919);
nor NOR3 (N2688, N2649, N2456, N628);
xor XOR2 (N2689, N2688, N2273);
or OR2 (N2690, N2676, N808);
nor NOR4 (N2691, N2681, N1519, N896, N1383);
not NOT1 (N2692, N2672);
and AND2 (N2693, N2685, N1160);
xor XOR2 (N2694, N2693, N2372);
xor XOR2 (N2695, N2687, N758);
buf BUF1 (N2696, N2686);
not NOT1 (N2697, N2690);
not NOT1 (N2698, N2661);
nor NOR3 (N2699, N2697, N659, N2035);
nand NAND4 (N2700, N2698, N2246, N724, N624);
nand NAND2 (N2701, N2696, N1784);
xor XOR2 (N2702, N2701, N2083);
buf BUF1 (N2703, N2699);
or OR4 (N2704, N2692, N1645, N2525, N2257);
not NOT1 (N2705, N2700);
nand NAND3 (N2706, N2691, N1520, N738);
and AND3 (N2707, N2695, N1300, N2069);
or OR3 (N2708, N2702, N1789, N2454);
buf BUF1 (N2709, N2704);
or OR2 (N2710, N2689, N255);
or OR4 (N2711, N2674, N1395, N1797, N367);
nand NAND3 (N2712, N2703, N2401, N976);
buf BUF1 (N2713, N2710);
and AND2 (N2714, N2709, N590);
or OR3 (N2715, N2711, N2353, N249);
or OR4 (N2716, N2715, N895, N1852, N153);
and AND3 (N2717, N2705, N104, N2032);
nand NAND4 (N2718, N2683, N1060, N223, N2315);
buf BUF1 (N2719, N2706);
xor XOR2 (N2720, N2719, N1211);
buf BUF1 (N2721, N2714);
buf BUF1 (N2722, N2721);
nor NOR4 (N2723, N2718, N954, N2689, N1399);
and AND2 (N2724, N2713, N484);
nor NOR4 (N2725, N2724, N237, N1207, N1920);
and AND4 (N2726, N2707, N1782, N468, N1797);
or OR2 (N2727, N2726, N439);
buf BUF1 (N2728, N2720);
or OR3 (N2729, N2708, N1154, N2113);
buf BUF1 (N2730, N2717);
and AND3 (N2731, N2722, N53, N2584);
and AND3 (N2732, N2712, N1558, N2395);
or OR4 (N2733, N2730, N240, N2585, N2408);
not NOT1 (N2734, N2725);
nor NOR3 (N2735, N2723, N188, N1288);
not NOT1 (N2736, N2734);
not NOT1 (N2737, N2736);
or OR4 (N2738, N2732, N109, N742, N1302);
nand NAND2 (N2739, N2731, N2232);
and AND4 (N2740, N2694, N473, N2441, N505);
xor XOR2 (N2741, N2716, N2321);
nand NAND3 (N2742, N2729, N438, N1365);
nand NAND2 (N2743, N2727, N1061);
nor NOR4 (N2744, N2739, N262, N1177, N45);
xor XOR2 (N2745, N2728, N729);
not NOT1 (N2746, N2742);
nor NOR2 (N2747, N2733, N1805);
xor XOR2 (N2748, N2744, N1495);
xor XOR2 (N2749, N2740, N594);
xor XOR2 (N2750, N2735, N1423);
and AND2 (N2751, N2749, N1942);
buf BUF1 (N2752, N2743);
xor XOR2 (N2753, N2747, N1224);
xor XOR2 (N2754, N2746, N2454);
nor NOR4 (N2755, N2741, N935, N2088, N2509);
nand NAND4 (N2756, N2755, N1256, N1628, N2247);
and AND4 (N2757, N2751, N826, N2204, N136);
xor XOR2 (N2758, N2748, N988);
xor XOR2 (N2759, N2754, N198);
nor NOR3 (N2760, N2759, N403, N1954);
nand NAND2 (N2761, N2756, N1523);
nor NOR4 (N2762, N2750, N130, N2745, N1492);
buf BUF1 (N2763, N2583);
buf BUF1 (N2764, N2737);
and AND4 (N2765, N2757, N912, N1690, N765);
or OR2 (N2766, N2762, N1518);
nand NAND2 (N2767, N2758, N2494);
or OR4 (N2768, N2767, N1783, N2712, N2264);
and AND4 (N2769, N2761, N1786, N1548, N2404);
nor NOR2 (N2770, N2765, N996);
not NOT1 (N2771, N2738);
not NOT1 (N2772, N2760);
nand NAND3 (N2773, N2769, N1301, N2021);
nand NAND4 (N2774, N2771, N2536, N475, N1943);
buf BUF1 (N2775, N2766);
nand NAND3 (N2776, N2773, N912, N186);
buf BUF1 (N2777, N2764);
or OR4 (N2778, N2774, N2138, N1751, N296);
buf BUF1 (N2779, N2768);
nand NAND2 (N2780, N2776, N2629);
nor NOR2 (N2781, N2763, N1143);
xor XOR2 (N2782, N2775, N1191);
or OR2 (N2783, N2781, N2728);
buf BUF1 (N2784, N2777);
or OR3 (N2785, N2770, N836, N1656);
buf BUF1 (N2786, N2772);
and AND2 (N2787, N2783, N311);
buf BUF1 (N2788, N2786);
or OR3 (N2789, N2753, N1200, N1468);
buf BUF1 (N2790, N2785);
xor XOR2 (N2791, N2778, N2722);
and AND3 (N2792, N2788, N656, N2191);
nor NOR3 (N2793, N2779, N2119, N68);
buf BUF1 (N2794, N2752);
and AND3 (N2795, N2793, N1845, N6);
and AND4 (N2796, N2784, N26, N1070, N2701);
and AND2 (N2797, N2795, N2145);
and AND4 (N2798, N2782, N1898, N1719, N1446);
buf BUF1 (N2799, N2796);
nor NOR4 (N2800, N2789, N1680, N1340, N1789);
not NOT1 (N2801, N2790);
and AND3 (N2802, N2780, N1367, N2704);
nand NAND3 (N2803, N2794, N39, N2094);
xor XOR2 (N2804, N2802, N2735);
buf BUF1 (N2805, N2801);
or OR4 (N2806, N2805, N602, N2488, N806);
and AND4 (N2807, N2797, N1384, N2579, N1267);
or OR4 (N2808, N2791, N2451, N1823, N866);
xor XOR2 (N2809, N2800, N356);
or OR4 (N2810, N2806, N796, N1289, N718);
nand NAND4 (N2811, N2810, N1351, N2466, N1368);
and AND4 (N2812, N2804, N102, N1687, N2018);
not NOT1 (N2813, N2792);
not NOT1 (N2814, N2811);
nor NOR3 (N2815, N2809, N625, N2685);
xor XOR2 (N2816, N2815, N362);
and AND2 (N2817, N2812, N279);
not NOT1 (N2818, N2816);
and AND4 (N2819, N2787, N357, N188, N2297);
nor NOR2 (N2820, N2813, N1587);
not NOT1 (N2821, N2814);
and AND3 (N2822, N2808, N2073, N1441);
nand NAND2 (N2823, N2798, N1311);
xor XOR2 (N2824, N2820, N2);
nor NOR3 (N2825, N2823, N825, N569);
and AND3 (N2826, N2803, N1596, N10);
or OR3 (N2827, N2821, N2574, N742);
not NOT1 (N2828, N2825);
or OR4 (N2829, N2824, N1943, N2442, N33);
xor XOR2 (N2830, N2822, N2218);
nand NAND3 (N2831, N2830, N1682, N1925);
nand NAND2 (N2832, N2817, N2511);
not NOT1 (N2833, N2818);
nand NAND4 (N2834, N2807, N1587, N2018, N1344);
and AND2 (N2835, N2829, N2407);
not NOT1 (N2836, N2826);
xor XOR2 (N2837, N2819, N1043);
nor NOR2 (N2838, N2799, N1269);
nor NOR2 (N2839, N2832, N2309);
xor XOR2 (N2840, N2835, N1513);
or OR3 (N2841, N2827, N2167, N2318);
nand NAND2 (N2842, N2839, N2825);
xor XOR2 (N2843, N2834, N820);
xor XOR2 (N2844, N2840, N1034);
and AND2 (N2845, N2841, N174);
nand NAND4 (N2846, N2843, N1493, N549, N2587);
nand NAND3 (N2847, N2846, N1924, N2164);
not NOT1 (N2848, N2831);
xor XOR2 (N2849, N2845, N1993);
not NOT1 (N2850, N2833);
nand NAND2 (N2851, N2836, N937);
not NOT1 (N2852, N2847);
buf BUF1 (N2853, N2851);
xor XOR2 (N2854, N2837, N2226);
xor XOR2 (N2855, N2852, N1179);
and AND3 (N2856, N2844, N107, N1513);
nand NAND2 (N2857, N2848, N1120);
nand NAND2 (N2858, N2842, N2158);
and AND3 (N2859, N2850, N2399, N1841);
or OR3 (N2860, N2858, N1180, N1474);
nor NOR2 (N2861, N2828, N1963);
nor NOR2 (N2862, N2855, N1880);
nor NOR2 (N2863, N2856, N2162);
nor NOR3 (N2864, N2853, N1671, N684);
xor XOR2 (N2865, N2860, N2023);
xor XOR2 (N2866, N2864, N2195);
nor NOR2 (N2867, N2863, N837);
nand NAND3 (N2868, N2867, N1237, N435);
and AND3 (N2869, N2849, N2602, N984);
nor NOR2 (N2870, N2862, N1645);
nand NAND2 (N2871, N2854, N2005);
nand NAND2 (N2872, N2857, N720);
buf BUF1 (N2873, N2868);
nor NOR4 (N2874, N2838, N1506, N1491, N2872);
nor NOR2 (N2875, N359, N1498);
buf BUF1 (N2876, N2875);
nand NAND4 (N2877, N2873, N737, N1958, N1646);
buf BUF1 (N2878, N2866);
nor NOR3 (N2879, N2878, N443, N914);
nand NAND4 (N2880, N2879, N232, N2749, N2644);
or OR2 (N2881, N2880, N1014);
nor NOR3 (N2882, N2869, N38, N1375);
xor XOR2 (N2883, N2874, N2236);
and AND2 (N2884, N2877, N482);
or OR4 (N2885, N2870, N1417, N296, N794);
buf BUF1 (N2886, N2865);
not NOT1 (N2887, N2882);
or OR3 (N2888, N2884, N786, N2754);
nand NAND3 (N2889, N2886, N2790, N1005);
buf BUF1 (N2890, N2871);
nand NAND3 (N2891, N2876, N700, N1713);
xor XOR2 (N2892, N2889, N2336);
nor NOR4 (N2893, N2881, N2005, N790, N1171);
nand NAND4 (N2894, N2892, N1027, N455, N74);
nor NOR4 (N2895, N2861, N2445, N208, N931);
buf BUF1 (N2896, N2893);
and AND2 (N2897, N2883, N1839);
xor XOR2 (N2898, N2895, N820);
buf BUF1 (N2899, N2887);
nand NAND2 (N2900, N2898, N1582);
and AND4 (N2901, N2891, N1399, N1861, N2133);
not NOT1 (N2902, N2899);
xor XOR2 (N2903, N2900, N1786);
nor NOR2 (N2904, N2890, N2773);
xor XOR2 (N2905, N2888, N1216);
or OR3 (N2906, N2903, N1662, N594);
and AND3 (N2907, N2901, N1596, N2589);
nor NOR4 (N2908, N2902, N1532, N2026, N2394);
not NOT1 (N2909, N2894);
nor NOR4 (N2910, N2885, N2230, N1285, N2343);
not NOT1 (N2911, N2908);
or OR3 (N2912, N2905, N1931, N1557);
and AND3 (N2913, N2910, N1433, N1545);
buf BUF1 (N2914, N2897);
nand NAND3 (N2915, N2914, N2586, N2597);
or OR2 (N2916, N2896, N653);
buf BUF1 (N2917, N2911);
not NOT1 (N2918, N2859);
buf BUF1 (N2919, N2916);
not NOT1 (N2920, N2907);
and AND3 (N2921, N2919, N2652, N1669);
nor NOR4 (N2922, N2906, N432, N2704, N1080);
or OR3 (N2923, N2904, N337, N1273);
or OR3 (N2924, N2921, N1827, N2540);
nand NAND4 (N2925, N2913, N1071, N2410, N802);
xor XOR2 (N2926, N2923, N2552);
nor NOR3 (N2927, N2915, N1408, N2326);
buf BUF1 (N2928, N2918);
nor NOR2 (N2929, N2912, N1906);
xor XOR2 (N2930, N2924, N1242);
xor XOR2 (N2931, N2927, N1560);
or OR4 (N2932, N2931, N2092, N1695, N1627);
nor NOR2 (N2933, N2929, N1550);
nor NOR2 (N2934, N2930, N123);
xor XOR2 (N2935, N2928, N256);
nor NOR2 (N2936, N2920, N380);
xor XOR2 (N2937, N2909, N256);
nor NOR4 (N2938, N2932, N91, N197, N1576);
buf BUF1 (N2939, N2937);
nand NAND3 (N2940, N2936, N1404, N1298);
xor XOR2 (N2941, N2940, N2579);
buf BUF1 (N2942, N2939);
nor NOR3 (N2943, N2942, N1054, N9);
or OR3 (N2944, N2941, N2721, N1877);
buf BUF1 (N2945, N2938);
xor XOR2 (N2946, N2933, N469);
nand NAND2 (N2947, N2922, N127);
nand NAND4 (N2948, N2943, N1377, N561, N863);
nand NAND3 (N2949, N2946, N631, N715);
nand NAND3 (N2950, N2944, N80, N1074);
nand NAND3 (N2951, N2948, N1953, N702);
or OR2 (N2952, N2950, N76);
not NOT1 (N2953, N2952);
nor NOR3 (N2954, N2934, N1730, N850);
xor XOR2 (N2955, N2954, N627);
xor XOR2 (N2956, N2935, N2176);
nor NOR2 (N2957, N2955, N69);
xor XOR2 (N2958, N2953, N1253);
buf BUF1 (N2959, N2956);
and AND4 (N2960, N2949, N729, N889, N2701);
nor NOR4 (N2961, N2926, N495, N2179, N1562);
buf BUF1 (N2962, N2957);
nand NAND2 (N2963, N2958, N597);
nand NAND3 (N2964, N2947, N2174, N2872);
xor XOR2 (N2965, N2959, N1838);
xor XOR2 (N2966, N2945, N1210);
xor XOR2 (N2967, N2963, N1);
or OR2 (N2968, N2967, N2793);
nand NAND2 (N2969, N2925, N170);
not NOT1 (N2970, N2965);
not NOT1 (N2971, N2969);
or OR4 (N2972, N2970, N2161, N2970, N2285);
xor XOR2 (N2973, N2968, N836);
not NOT1 (N2974, N2917);
and AND2 (N2975, N2974, N2447);
buf BUF1 (N2976, N2975);
or OR4 (N2977, N2962, N2138, N790, N2089);
and AND4 (N2978, N2964, N226, N2594, N1300);
xor XOR2 (N2979, N2960, N447);
xor XOR2 (N2980, N2978, N1043);
not NOT1 (N2981, N2961);
not NOT1 (N2982, N2966);
nor NOR3 (N2983, N2973, N2286, N2038);
and AND4 (N2984, N2977, N2077, N514, N2886);
not NOT1 (N2985, N2984);
buf BUF1 (N2986, N2972);
xor XOR2 (N2987, N2979, N850);
not NOT1 (N2988, N2951);
buf BUF1 (N2989, N2988);
nand NAND4 (N2990, N2983, N2130, N1668, N2981);
not NOT1 (N2991, N1646);
and AND3 (N2992, N2986, N2749, N1638);
not NOT1 (N2993, N2982);
not NOT1 (N2994, N2991);
nand NAND4 (N2995, N2976, N2154, N137, N1739);
or OR4 (N2996, N2992, N2263, N2693, N1126);
and AND2 (N2997, N2996, N2076);
buf BUF1 (N2998, N2994);
nand NAND3 (N2999, N2987, N735, N1150);
or OR2 (N3000, N2980, N770);
nand NAND3 (N3001, N2998, N1280, N354);
buf BUF1 (N3002, N3001);
buf BUF1 (N3003, N2999);
nand NAND2 (N3004, N3002, N1507);
and AND4 (N3005, N2971, N870, N2586, N468);
and AND4 (N3006, N2997, N2342, N2250, N621);
xor XOR2 (N3007, N2990, N601);
and AND2 (N3008, N2995, N1470);
nor NOR4 (N3009, N3003, N1984, N2058, N2966);
nand NAND3 (N3010, N2985, N776, N2178);
not NOT1 (N3011, N3007);
not NOT1 (N3012, N3009);
nor NOR2 (N3013, N3006, N2573);
xor XOR2 (N3014, N3008, N2370);
or OR3 (N3015, N3004, N1666, N1159);
buf BUF1 (N3016, N3015);
xor XOR2 (N3017, N3012, N2415);
not NOT1 (N3018, N3000);
and AND2 (N3019, N3010, N109);
not NOT1 (N3020, N3016);
and AND3 (N3021, N2993, N1705, N2652);
or OR2 (N3022, N3017, N879);
xor XOR2 (N3023, N3011, N412);
not NOT1 (N3024, N3021);
buf BUF1 (N3025, N3018);
nor NOR3 (N3026, N3025, N2988, N1586);
nand NAND3 (N3027, N3013, N1296, N2271);
nor NOR2 (N3028, N3005, N1645);
or OR4 (N3029, N3014, N103, N79, N1918);
nand NAND2 (N3030, N3023, N811);
nor NOR2 (N3031, N3029, N1947);
not NOT1 (N3032, N3024);
nor NOR2 (N3033, N3019, N327);
buf BUF1 (N3034, N3020);
buf BUF1 (N3035, N3031);
buf BUF1 (N3036, N3027);
nand NAND2 (N3037, N3035, N1702);
nand NAND2 (N3038, N3036, N2245);
not NOT1 (N3039, N3033);
or OR2 (N3040, N2989, N887);
nor NOR3 (N3041, N3037, N1953, N113);
xor XOR2 (N3042, N3032, N1852);
buf BUF1 (N3043, N3030);
nand NAND2 (N3044, N3039, N936);
nor NOR3 (N3045, N3042, N69, N853);
nor NOR3 (N3046, N3026, N496, N2987);
or OR3 (N3047, N3034, N2901, N1993);
xor XOR2 (N3048, N3028, N397);
nor NOR4 (N3049, N3040, N421, N2056, N1440);
and AND4 (N3050, N3045, N1288, N2258, N2919);
nor NOR4 (N3051, N3041, N2997, N2212, N2087);
or OR2 (N3052, N3049, N2048);
and AND2 (N3053, N3022, N1214);
nand NAND4 (N3054, N3038, N2243, N2074, N459);
not NOT1 (N3055, N3053);
or OR4 (N3056, N3048, N2058, N2614, N2021);
not NOT1 (N3057, N3056);
nor NOR2 (N3058, N3050, N1724);
not NOT1 (N3059, N3057);
and AND3 (N3060, N3055, N2262, N2647);
buf BUF1 (N3061, N3046);
not NOT1 (N3062, N3051);
nor NOR4 (N3063, N3047, N2966, N355, N2697);
xor XOR2 (N3064, N3059, N1721);
and AND4 (N3065, N3058, N3036, N954, N1069);
or OR4 (N3066, N3063, N119, N2360, N1943);
or OR2 (N3067, N3066, N2430);
and AND3 (N3068, N3060, N346, N2822);
nand NAND2 (N3069, N3054, N582);
xor XOR2 (N3070, N3064, N722);
buf BUF1 (N3071, N3070);
buf BUF1 (N3072, N3044);
nor NOR3 (N3073, N3072, N2926, N666);
xor XOR2 (N3074, N3067, N1413);
nand NAND4 (N3075, N3069, N2373, N252, N1517);
nor NOR2 (N3076, N3061, N2340);
xor XOR2 (N3077, N3075, N2921);
buf BUF1 (N3078, N3073);
nor NOR4 (N3079, N3077, N594, N1530, N1488);
and AND3 (N3080, N3071, N109, N630);
nand NAND3 (N3081, N3079, N1902, N1563);
not NOT1 (N3082, N3081);
not NOT1 (N3083, N3043);
nor NOR4 (N3084, N3062, N862, N2824, N2886);
not NOT1 (N3085, N3068);
nor NOR2 (N3086, N3065, N1506);
or OR2 (N3087, N3082, N1852);
xor XOR2 (N3088, N3074, N856);
not NOT1 (N3089, N3076);
nand NAND3 (N3090, N3085, N2457, N873);
buf BUF1 (N3091, N3089);
not NOT1 (N3092, N3088);
nor NOR3 (N3093, N3084, N2599, N828);
nand NAND3 (N3094, N3090, N2875, N2907);
not NOT1 (N3095, N3080);
xor XOR2 (N3096, N3087, N415);
or OR4 (N3097, N3086, N1684, N2719, N1216);
nor NOR2 (N3098, N3092, N565);
xor XOR2 (N3099, N3083, N1480);
and AND3 (N3100, N3052, N1637, N2492);
nand NAND3 (N3101, N3093, N1351, N2833);
and AND3 (N3102, N3096, N1907, N2357);
buf BUF1 (N3103, N3094);
xor XOR2 (N3104, N3102, N1236);
and AND3 (N3105, N3095, N1004, N1748);
xor XOR2 (N3106, N3098, N773);
not NOT1 (N3107, N3091);
nand NAND3 (N3108, N3100, N1657, N1311);
nand NAND2 (N3109, N3097, N1722);
not NOT1 (N3110, N3108);
or OR4 (N3111, N3101, N684, N816, N3073);
and AND4 (N3112, N3110, N832, N1401, N1909);
or OR2 (N3113, N3111, N1423);
nor NOR2 (N3114, N3078, N1434);
nor NOR4 (N3115, N3107, N2703, N616, N1454);
buf BUF1 (N3116, N3115);
or OR2 (N3117, N3116, N2205);
nor NOR3 (N3118, N3105, N1702, N2898);
nor NOR2 (N3119, N3112, N1662);
or OR3 (N3120, N3119, N2824, N904);
or OR3 (N3121, N3109, N2732, N2892);
and AND3 (N3122, N3117, N3029, N2434);
xor XOR2 (N3123, N3114, N1866);
and AND3 (N3124, N3122, N1251, N2680);
xor XOR2 (N3125, N3124, N200);
or OR3 (N3126, N3125, N1961, N858);
not NOT1 (N3127, N3126);
or OR3 (N3128, N3123, N2387, N1277);
and AND2 (N3129, N3103, N1491);
or OR4 (N3130, N3127, N575, N653, N1839);
and AND2 (N3131, N3129, N1526);
and AND3 (N3132, N3121, N1492, N2192);
nor NOR4 (N3133, N3113, N2953, N2800, N1978);
buf BUF1 (N3134, N3131);
or OR3 (N3135, N3120, N2009, N1662);
or OR2 (N3136, N3099, N2149);
not NOT1 (N3137, N3118);
not NOT1 (N3138, N3134);
not NOT1 (N3139, N3136);
xor XOR2 (N3140, N3133, N1881);
xor XOR2 (N3141, N3132, N1062);
nor NOR4 (N3142, N3104, N1434, N1526, N1919);
not NOT1 (N3143, N3130);
nand NAND2 (N3144, N3128, N3088);
buf BUF1 (N3145, N3140);
not NOT1 (N3146, N3138);
and AND4 (N3147, N3135, N2170, N296, N1416);
nor NOR3 (N3148, N3142, N2535, N1571);
and AND2 (N3149, N3143, N2393);
buf BUF1 (N3150, N3141);
nand NAND2 (N3151, N3150, N835);
and AND4 (N3152, N3151, N1770, N2247, N2751);
nor NOR2 (N3153, N3149, N2910);
nand NAND3 (N3154, N3144, N2255, N1924);
xor XOR2 (N3155, N3152, N2146);
or OR2 (N3156, N3106, N620);
and AND2 (N3157, N3145, N1122);
nand NAND4 (N3158, N3153, N324, N3130, N1836);
not NOT1 (N3159, N3157);
buf BUF1 (N3160, N3137);
buf BUF1 (N3161, N3146);
xor XOR2 (N3162, N3139, N1421);
nand NAND4 (N3163, N3155, N525, N1065, N429);
not NOT1 (N3164, N3163);
xor XOR2 (N3165, N3161, N757);
and AND2 (N3166, N3165, N1739);
or OR2 (N3167, N3162, N1586);
and AND2 (N3168, N3156, N2251);
not NOT1 (N3169, N3148);
nor NOR3 (N3170, N3166, N807, N1470);
and AND3 (N3171, N3147, N1300, N2924);
nor NOR4 (N3172, N3160, N2468, N2216, N1153);
nand NAND3 (N3173, N3154, N909, N2085);
buf BUF1 (N3174, N3169);
or OR2 (N3175, N3171, N207);
xor XOR2 (N3176, N3159, N2764);
buf BUF1 (N3177, N3175);
and AND4 (N3178, N3172, N1505, N654, N971);
and AND4 (N3179, N3168, N341, N357, N696);
not NOT1 (N3180, N3177);
xor XOR2 (N3181, N3176, N1780);
xor XOR2 (N3182, N3167, N2500);
or OR2 (N3183, N3180, N266);
not NOT1 (N3184, N3179);
nor NOR3 (N3185, N3164, N2595, N2204);
nand NAND3 (N3186, N3185, N2262, N370);
not NOT1 (N3187, N3182);
or OR2 (N3188, N3184, N297);
buf BUF1 (N3189, N3186);
nor NOR4 (N3190, N3178, N2757, N83, N2083);
not NOT1 (N3191, N3187);
buf BUF1 (N3192, N3183);
or OR3 (N3193, N3174, N2725, N554);
buf BUF1 (N3194, N3189);
buf BUF1 (N3195, N3181);
or OR4 (N3196, N3170, N2975, N3077, N1373);
and AND3 (N3197, N3193, N1592, N2996);
nand NAND4 (N3198, N3197, N552, N281, N2228);
and AND4 (N3199, N3196, N1225, N1564, N933);
and AND3 (N3200, N3190, N2362, N790);
nor NOR2 (N3201, N3158, N1348);
or OR4 (N3202, N3191, N1776, N2987, N2046);
and AND3 (N3203, N3195, N1831, N1303);
and AND3 (N3204, N3192, N1598, N2166);
buf BUF1 (N3205, N3203);
not NOT1 (N3206, N3199);
buf BUF1 (N3207, N3201);
nand NAND4 (N3208, N3173, N2168, N1196, N1149);
nand NAND3 (N3209, N3200, N1029, N531);
nand NAND3 (N3210, N3207, N2260, N3132);
nand NAND3 (N3211, N3202, N309, N217);
nor NOR2 (N3212, N3208, N2192);
nor NOR3 (N3213, N3205, N1895, N2930);
not NOT1 (N3214, N3209);
buf BUF1 (N3215, N3213);
and AND2 (N3216, N3204, N786);
nor NOR4 (N3217, N3214, N2985, N2504, N983);
nor NOR4 (N3218, N3211, N1506, N3189, N1819);
xor XOR2 (N3219, N3210, N1726);
not NOT1 (N3220, N3212);
buf BUF1 (N3221, N3198);
not NOT1 (N3222, N3188);
buf BUF1 (N3223, N3222);
xor XOR2 (N3224, N3216, N1841);
buf BUF1 (N3225, N3217);
buf BUF1 (N3226, N3223);
and AND2 (N3227, N3218, N1501);
and AND4 (N3228, N3224, N967, N1535, N2023);
nand NAND4 (N3229, N3225, N1812, N398, N2808);
and AND4 (N3230, N3227, N2718, N1947, N788);
and AND3 (N3231, N3219, N648, N955);
and AND3 (N3232, N3221, N703, N2673);
or OR4 (N3233, N3228, N85, N192, N1925);
nand NAND2 (N3234, N3230, N1951);
nand NAND3 (N3235, N3215, N1841, N1899);
nor NOR4 (N3236, N3220, N2859, N416, N567);
and AND4 (N3237, N3235, N1654, N386, N1707);
and AND3 (N3238, N3234, N2880, N308);
buf BUF1 (N3239, N3237);
nor NOR4 (N3240, N3233, N2565, N1369, N819);
and AND3 (N3241, N3229, N293, N2365);
xor XOR2 (N3242, N3226, N2381);
nand NAND3 (N3243, N3241, N1519, N1659);
nor NOR2 (N3244, N3206, N3111);
not NOT1 (N3245, N3242);
nor NOR3 (N3246, N3244, N3077, N3062);
nor NOR3 (N3247, N3246, N2017, N2100);
xor XOR2 (N3248, N3243, N553);
and AND2 (N3249, N3238, N2434);
nor NOR2 (N3250, N3249, N1489);
xor XOR2 (N3251, N3239, N727);
nand NAND4 (N3252, N3250, N1983, N1538, N2496);
nor NOR3 (N3253, N3236, N806, N2217);
not NOT1 (N3254, N3194);
or OR4 (N3255, N3231, N2447, N3137, N799);
and AND2 (N3256, N3240, N43);
and AND2 (N3257, N3251, N728);
not NOT1 (N3258, N3254);
nor NOR2 (N3259, N3232, N1274);
xor XOR2 (N3260, N3247, N166);
nand NAND2 (N3261, N3256, N766);
and AND4 (N3262, N3259, N1061, N619, N2242);
nor NOR2 (N3263, N3258, N1536);
or OR3 (N3264, N3263, N1177, N920);
or OR2 (N3265, N3262, N67);
and AND2 (N3266, N3252, N1338);
nor NOR4 (N3267, N3260, N873, N1649, N2734);
buf BUF1 (N3268, N3261);
not NOT1 (N3269, N3266);
nand NAND4 (N3270, N3253, N2548, N3237, N974);
nand NAND4 (N3271, N3269, N114, N1596, N1462);
not NOT1 (N3272, N3267);
nand NAND3 (N3273, N3271, N2783, N1840);
or OR2 (N3274, N3248, N2354);
and AND2 (N3275, N3264, N2619);
nand NAND4 (N3276, N3270, N1511, N3075, N2311);
buf BUF1 (N3277, N3255);
and AND3 (N3278, N3277, N474, N502);
nor NOR3 (N3279, N3265, N1233, N2421);
buf BUF1 (N3280, N3268);
nand NAND2 (N3281, N3275, N3231);
or OR4 (N3282, N3257, N2108, N3232, N2606);
nand NAND2 (N3283, N3274, N2674);
nand NAND4 (N3284, N3282, N3114, N1863, N1098);
not NOT1 (N3285, N3278);
buf BUF1 (N3286, N3281);
or OR4 (N3287, N3283, N2242, N716, N1987);
not NOT1 (N3288, N3286);
not NOT1 (N3289, N3280);
not NOT1 (N3290, N3284);
xor XOR2 (N3291, N3276, N3257);
buf BUF1 (N3292, N3279);
and AND2 (N3293, N3288, N1571);
nand NAND4 (N3294, N3292, N936, N1511, N337);
nor NOR4 (N3295, N3290, N2512, N2948, N1736);
xor XOR2 (N3296, N3287, N1893);
nor NOR3 (N3297, N3245, N1222, N2118);
not NOT1 (N3298, N3285);
nor NOR3 (N3299, N3272, N1855, N1013);
nand NAND4 (N3300, N3293, N75, N2987, N551);
buf BUF1 (N3301, N3297);
and AND3 (N3302, N3298, N3193, N2042);
nand NAND4 (N3303, N3273, N2785, N2190, N1304);
not NOT1 (N3304, N3303);
nor NOR4 (N3305, N3299, N1004, N2885, N2876);
or OR2 (N3306, N3300, N3001);
not NOT1 (N3307, N3306);
xor XOR2 (N3308, N3305, N3159);
xor XOR2 (N3309, N3301, N1803);
nand NAND3 (N3310, N3294, N769, N2945);
nand NAND4 (N3311, N3308, N897, N520, N1074);
nor NOR3 (N3312, N3296, N1520, N286);
nor NOR2 (N3313, N3309, N378);
not NOT1 (N3314, N3311);
buf BUF1 (N3315, N3313);
xor XOR2 (N3316, N3304, N3005);
nand NAND4 (N3317, N3310, N1722, N3023, N3146);
buf BUF1 (N3318, N3307);
nand NAND3 (N3319, N3289, N2322, N780);
xor XOR2 (N3320, N3295, N46);
and AND4 (N3321, N3314, N1301, N3268, N1609);
nand NAND4 (N3322, N3318, N2486, N884, N2393);
nor NOR4 (N3323, N3291, N420, N452, N1415);
nor NOR2 (N3324, N3316, N2653);
buf BUF1 (N3325, N3321);
buf BUF1 (N3326, N3319);
xor XOR2 (N3327, N3302, N43);
nor NOR4 (N3328, N3320, N2508, N277, N2393);
buf BUF1 (N3329, N3325);
and AND4 (N3330, N3322, N1553, N1885, N1975);
nand NAND2 (N3331, N3329, N190);
nor NOR3 (N3332, N3328, N2368, N2301);
nor NOR3 (N3333, N3330, N1021, N1276);
xor XOR2 (N3334, N3323, N364);
xor XOR2 (N3335, N3317, N2921);
nand NAND2 (N3336, N3332, N1001);
nand NAND4 (N3337, N3335, N28, N1490, N2900);
or OR2 (N3338, N3331, N959);
and AND4 (N3339, N3337, N472, N1525, N3054);
or OR3 (N3340, N3334, N75, N2702);
nor NOR4 (N3341, N3315, N1456, N2970, N539);
buf BUF1 (N3342, N3326);
and AND2 (N3343, N3340, N683);
or OR3 (N3344, N3339, N613, N136);
nand NAND2 (N3345, N3312, N3291);
or OR3 (N3346, N3345, N3195, N905);
not NOT1 (N3347, N3346);
nor NOR2 (N3348, N3344, N1028);
nor NOR4 (N3349, N3327, N843, N3150, N1648);
or OR2 (N3350, N3333, N1891);
nand NAND4 (N3351, N3343, N278, N1204, N3017);
buf BUF1 (N3352, N3336);
nand NAND2 (N3353, N3338, N3186);
buf BUF1 (N3354, N3348);
not NOT1 (N3355, N3350);
xor XOR2 (N3356, N3351, N2670);
and AND4 (N3357, N3347, N1517, N2399, N1509);
nor NOR4 (N3358, N3349, N389, N2252, N2680);
and AND4 (N3359, N3352, N2352, N2555, N922);
xor XOR2 (N3360, N3357, N1690);
and AND4 (N3361, N3324, N976, N965, N2134);
or OR2 (N3362, N3356, N1677);
or OR2 (N3363, N3342, N3287);
xor XOR2 (N3364, N3354, N717);
or OR2 (N3365, N3364, N1977);
buf BUF1 (N3366, N3355);
nor NOR2 (N3367, N3361, N1526);
xor XOR2 (N3368, N3353, N2191);
buf BUF1 (N3369, N3341);
not NOT1 (N3370, N3368);
not NOT1 (N3371, N3369);
not NOT1 (N3372, N3371);
nor NOR3 (N3373, N3359, N1520, N1203);
buf BUF1 (N3374, N3366);
nor NOR3 (N3375, N3372, N291, N3304);
and AND4 (N3376, N3374, N829, N3094, N465);
xor XOR2 (N3377, N3362, N2328);
xor XOR2 (N3378, N3363, N465);
xor XOR2 (N3379, N3360, N501);
buf BUF1 (N3380, N3376);
or OR4 (N3381, N3380, N1524, N1962, N23);
nand NAND2 (N3382, N3378, N851);
not NOT1 (N3383, N3377);
and AND4 (N3384, N3383, N1411, N3157, N1911);
or OR2 (N3385, N3370, N1422);
not NOT1 (N3386, N3384);
xor XOR2 (N3387, N3375, N1757);
xor XOR2 (N3388, N3365, N1941);
nand NAND2 (N3389, N3373, N2916);
not NOT1 (N3390, N3386);
or OR4 (N3391, N3382, N644, N2274, N880);
not NOT1 (N3392, N3358);
and AND4 (N3393, N3367, N3327, N1797, N1536);
not NOT1 (N3394, N3388);
nand NAND4 (N3395, N3385, N2816, N3324, N1228);
xor XOR2 (N3396, N3387, N1726);
nor NOR2 (N3397, N3379, N3225);
nor NOR4 (N3398, N3392, N3336, N1312, N2154);
not NOT1 (N3399, N3398);
nand NAND4 (N3400, N3397, N521, N1469, N2839);
nand NAND3 (N3401, N3389, N496, N1801);
buf BUF1 (N3402, N3391);
not NOT1 (N3403, N3399);
nor NOR3 (N3404, N3390, N3173, N353);
xor XOR2 (N3405, N3393, N2927);
nand NAND2 (N3406, N3402, N1656);
nand NAND3 (N3407, N3395, N2526, N2086);
or OR3 (N3408, N3403, N1892, N2924);
xor XOR2 (N3409, N3401, N1284);
nor NOR2 (N3410, N3396, N260);
xor XOR2 (N3411, N3407, N2848);
nor NOR2 (N3412, N3410, N26);
and AND3 (N3413, N3411, N541, N2406);
not NOT1 (N3414, N3405);
or OR4 (N3415, N3381, N1158, N1914, N902);
or OR2 (N3416, N3415, N230);
buf BUF1 (N3417, N3406);
nor NOR4 (N3418, N3414, N397, N2486, N1269);
buf BUF1 (N3419, N3412);
not NOT1 (N3420, N3413);
not NOT1 (N3421, N3420);
buf BUF1 (N3422, N3409);
and AND3 (N3423, N3394, N2983, N3055);
buf BUF1 (N3424, N3400);
nor NOR3 (N3425, N3418, N1429, N173);
nor NOR2 (N3426, N3422, N3104);
nor NOR2 (N3427, N3425, N1431);
buf BUF1 (N3428, N3419);
nor NOR3 (N3429, N3426, N3334, N3389);
or OR2 (N3430, N3416, N2642);
buf BUF1 (N3431, N3408);
not NOT1 (N3432, N3427);
and AND4 (N3433, N3430, N3015, N2912, N2651);
xor XOR2 (N3434, N3424, N453);
and AND3 (N3435, N3431, N955, N343);
not NOT1 (N3436, N3428);
and AND4 (N3437, N3432, N980, N2128, N1164);
and AND4 (N3438, N3435, N955, N2280, N1738);
buf BUF1 (N3439, N3423);
not NOT1 (N3440, N3438);
nor NOR3 (N3441, N3433, N926, N3229);
and AND2 (N3442, N3434, N2138);
nand NAND4 (N3443, N3436, N384, N340, N1557);
or OR2 (N3444, N3441, N3207);
nand NAND3 (N3445, N3404, N3120, N2216);
or OR2 (N3446, N3437, N1570);
nor NOR4 (N3447, N3439, N2910, N1638, N3263);
xor XOR2 (N3448, N3429, N1109);
not NOT1 (N3449, N3442);
or OR4 (N3450, N3443, N1394, N1494, N997);
and AND2 (N3451, N3440, N687);
buf BUF1 (N3452, N3421);
not NOT1 (N3453, N3449);
and AND2 (N3454, N3452, N1616);
nor NOR4 (N3455, N3447, N2337, N2069, N1346);
not NOT1 (N3456, N3417);
and AND3 (N3457, N3444, N1542, N472);
not NOT1 (N3458, N3456);
xor XOR2 (N3459, N3446, N2378);
nand NAND2 (N3460, N3454, N1526);
and AND2 (N3461, N3450, N3071);
not NOT1 (N3462, N3460);
nor NOR3 (N3463, N3445, N2162, N2677);
or OR4 (N3464, N3451, N688, N1058, N1821);
or OR3 (N3465, N3457, N888, N1154);
not NOT1 (N3466, N3453);
xor XOR2 (N3467, N3455, N1341);
xor XOR2 (N3468, N3448, N1244);
buf BUF1 (N3469, N3467);
and AND3 (N3470, N3468, N3330, N2423);
or OR3 (N3471, N3463, N2721, N565);
nor NOR2 (N3472, N3466, N181);
and AND3 (N3473, N3464, N2063, N1321);
nand NAND4 (N3474, N3465, N54, N170, N3043);
nand NAND3 (N3475, N3471, N3451, N2216);
buf BUF1 (N3476, N3475);
not NOT1 (N3477, N3459);
or OR2 (N3478, N3472, N158);
buf BUF1 (N3479, N3461);
nor NOR4 (N3480, N3462, N31, N97, N1798);
buf BUF1 (N3481, N3480);
buf BUF1 (N3482, N3474);
nand NAND2 (N3483, N3477, N2183);
not NOT1 (N3484, N3473);
xor XOR2 (N3485, N3484, N3);
not NOT1 (N3486, N3483);
and AND3 (N3487, N3486, N2714, N3026);
buf BUF1 (N3488, N3476);
nor NOR2 (N3489, N3487, N3207);
and AND4 (N3490, N3478, N3157, N541, N2700);
and AND2 (N3491, N3482, N2767);
or OR2 (N3492, N3489, N2396);
not NOT1 (N3493, N3479);
and AND4 (N3494, N3493, N1556, N1669, N156);
and AND4 (N3495, N3470, N2459, N2292, N730);
nand NAND3 (N3496, N3458, N916, N1805);
and AND2 (N3497, N3490, N1819);
or OR4 (N3498, N3496, N2572, N3250, N2336);
buf BUF1 (N3499, N3494);
buf BUF1 (N3500, N3498);
buf BUF1 (N3501, N3481);
nand NAND2 (N3502, N3488, N677);
buf BUF1 (N3503, N3469);
xor XOR2 (N3504, N3500, N508);
or OR3 (N3505, N3492, N1877, N3020);
nand NAND3 (N3506, N3499, N3203, N1929);
nand NAND3 (N3507, N3491, N819, N3344);
nand NAND4 (N3508, N3502, N2605, N3010, N3436);
buf BUF1 (N3509, N3508);
or OR4 (N3510, N3504, N2143, N1635, N719);
nand NAND3 (N3511, N3510, N1458, N2838);
nand NAND2 (N3512, N3505, N2090);
xor XOR2 (N3513, N3485, N1996);
nor NOR3 (N3514, N3503, N2876, N3388);
buf BUF1 (N3515, N3497);
or OR4 (N3516, N3509, N2685, N2335, N2843);
buf BUF1 (N3517, N3506);
nand NAND4 (N3518, N3517, N2075, N2207, N1942);
xor XOR2 (N3519, N3495, N2388);
and AND2 (N3520, N3507, N3047);
buf BUF1 (N3521, N3516);
and AND3 (N3522, N3515, N1641, N3214);
nor NOR2 (N3523, N3522, N887);
nor NOR4 (N3524, N3512, N97, N2289, N402);
and AND2 (N3525, N3518, N1882);
nor NOR3 (N3526, N3519, N2231, N811);
buf BUF1 (N3527, N3513);
not NOT1 (N3528, N3524);
nor NOR4 (N3529, N3525, N3023, N754, N1201);
and AND3 (N3530, N3521, N2234, N910);
and AND2 (N3531, N3530, N108);
nor NOR2 (N3532, N3527, N2998);
and AND3 (N3533, N3501, N1030, N588);
xor XOR2 (N3534, N3526, N185);
and AND3 (N3535, N3523, N410, N2525);
buf BUF1 (N3536, N3532);
not NOT1 (N3537, N3514);
nor NOR4 (N3538, N3528, N2201, N1980, N1262);
buf BUF1 (N3539, N3537);
and AND3 (N3540, N3539, N1479, N497);
xor XOR2 (N3541, N3535, N459);
nand NAND4 (N3542, N3511, N2152, N3160, N2283);
nand NAND3 (N3543, N3520, N2090, N2376);
not NOT1 (N3544, N3541);
or OR3 (N3545, N3542, N3464, N1917);
nor NOR3 (N3546, N3540, N1736, N2658);
buf BUF1 (N3547, N3546);
nor NOR4 (N3548, N3531, N141, N1063, N1763);
nand NAND3 (N3549, N3545, N1523, N1044);
buf BUF1 (N3550, N3543);
not NOT1 (N3551, N3550);
nor NOR3 (N3552, N3536, N247, N240);
not NOT1 (N3553, N3534);
nand NAND4 (N3554, N3548, N1162, N1677, N812);
nand NAND3 (N3555, N3538, N335, N458);
xor XOR2 (N3556, N3552, N2156);
xor XOR2 (N3557, N3544, N2711);
not NOT1 (N3558, N3555);
xor XOR2 (N3559, N3529, N2419);
nand NAND3 (N3560, N3553, N3181, N2758);
xor XOR2 (N3561, N3549, N1820);
nand NAND4 (N3562, N3547, N1741, N3089, N2786);
not NOT1 (N3563, N3557);
nand NAND2 (N3564, N3556, N1066);
xor XOR2 (N3565, N3560, N928);
xor XOR2 (N3566, N3551, N1838);
and AND2 (N3567, N3561, N2433);
and AND3 (N3568, N3564, N3534, N3380);
nand NAND4 (N3569, N3558, N3133, N2245, N1651);
not NOT1 (N3570, N3563);
nand NAND4 (N3571, N3554, N233, N992, N3105);
not NOT1 (N3572, N3570);
or OR3 (N3573, N3572, N3330, N1997);
and AND4 (N3574, N3565, N570, N1960, N2349);
or OR4 (N3575, N3568, N1775, N1928, N1909);
not NOT1 (N3576, N3562);
xor XOR2 (N3577, N3567, N3412);
buf BUF1 (N3578, N3569);
and AND2 (N3579, N3576, N3403);
and AND3 (N3580, N3573, N755, N1238);
and AND2 (N3581, N3566, N2273);
not NOT1 (N3582, N3559);
nor NOR2 (N3583, N3581, N2766);
xor XOR2 (N3584, N3577, N2723);
buf BUF1 (N3585, N3578);
nor NOR3 (N3586, N3584, N1475, N1020);
buf BUF1 (N3587, N3585);
not NOT1 (N3588, N3533);
xor XOR2 (N3589, N3583, N3283);
and AND4 (N3590, N3574, N1444, N1359, N2423);
and AND2 (N3591, N3586, N1061);
or OR3 (N3592, N3580, N3352, N3547);
buf BUF1 (N3593, N3592);
buf BUF1 (N3594, N3591);
or OR4 (N3595, N3593, N803, N723, N2800);
buf BUF1 (N3596, N3587);
or OR4 (N3597, N3582, N2652, N75, N3576);
not NOT1 (N3598, N3596);
or OR4 (N3599, N3579, N2978, N2141, N2115);
nand NAND2 (N3600, N3571, N3522);
nand NAND3 (N3601, N3575, N130, N1833);
not NOT1 (N3602, N3601);
and AND2 (N3603, N3597, N107);
or OR3 (N3604, N3595, N1502, N3350);
or OR4 (N3605, N3600, N3271, N1294, N3358);
and AND4 (N3606, N3602, N677, N935, N276);
nor NOR2 (N3607, N3594, N713);
xor XOR2 (N3608, N3588, N1929);
and AND4 (N3609, N3605, N355, N1270, N350);
nand NAND4 (N3610, N3609, N574, N2448, N1056);
and AND3 (N3611, N3608, N1684, N1221);
and AND2 (N3612, N3598, N3538);
or OR3 (N3613, N3604, N404, N1684);
buf BUF1 (N3614, N3610);
and AND4 (N3615, N3607, N3206, N1850, N1368);
xor XOR2 (N3616, N3603, N2469);
xor XOR2 (N3617, N3614, N2636);
or OR4 (N3618, N3589, N1428, N1112, N3601);
nor NOR4 (N3619, N3618, N441, N1162, N2590);
buf BUF1 (N3620, N3615);
buf BUF1 (N3621, N3606);
xor XOR2 (N3622, N3621, N3377);
nor NOR3 (N3623, N3620, N131, N3126);
nor NOR3 (N3624, N3613, N2725, N3013);
not NOT1 (N3625, N3622);
and AND2 (N3626, N3623, N1354);
xor XOR2 (N3627, N3611, N1642);
not NOT1 (N3628, N3619);
and AND4 (N3629, N3599, N2636, N1419, N1234);
or OR2 (N3630, N3627, N1062);
nor NOR3 (N3631, N3612, N122, N1051);
nand NAND3 (N3632, N3630, N3569, N2568);
nor NOR3 (N3633, N3628, N57, N1827);
nor NOR3 (N3634, N3633, N1439, N1228);
nand NAND4 (N3635, N3616, N1311, N880, N851);
buf BUF1 (N3636, N3590);
or OR2 (N3637, N3631, N2123);
and AND2 (N3638, N3637, N3062);
buf BUF1 (N3639, N3617);
not NOT1 (N3640, N3625);
not NOT1 (N3641, N3636);
nand NAND2 (N3642, N3629, N567);
buf BUF1 (N3643, N3642);
buf BUF1 (N3644, N3638);
not NOT1 (N3645, N3635);
nor NOR4 (N3646, N3639, N2937, N1795, N1408);
not NOT1 (N3647, N3646);
and AND2 (N3648, N3643, N2416);
not NOT1 (N3649, N3648);
xor XOR2 (N3650, N3634, N1202);
or OR3 (N3651, N3640, N2383, N223);
nor NOR2 (N3652, N3644, N3499);
buf BUF1 (N3653, N3632);
buf BUF1 (N3654, N3626);
nand NAND2 (N3655, N3641, N3609);
not NOT1 (N3656, N3655);
xor XOR2 (N3657, N3647, N1697);
and AND4 (N3658, N3645, N3122, N3411, N2664);
nand NAND3 (N3659, N3656, N2177, N1291);
and AND4 (N3660, N3653, N114, N796, N2785);
or OR3 (N3661, N3651, N937, N326);
not NOT1 (N3662, N3652);
not NOT1 (N3663, N3662);
nor NOR3 (N3664, N3658, N2260, N962);
or OR3 (N3665, N3664, N3365, N2452);
and AND3 (N3666, N3654, N2894, N1535);
xor XOR2 (N3667, N3649, N1110);
nand NAND4 (N3668, N3660, N2342, N3077, N2989);
nand NAND3 (N3669, N3661, N3087, N2039);
nand NAND2 (N3670, N3667, N470);
nand NAND3 (N3671, N3669, N2187, N1902);
or OR2 (N3672, N3659, N995);
buf BUF1 (N3673, N3665);
or OR2 (N3674, N3672, N3095);
nor NOR4 (N3675, N3671, N670, N3122, N3566);
buf BUF1 (N3676, N3668);
and AND2 (N3677, N3673, N3200);
and AND3 (N3678, N3657, N642, N2292);
not NOT1 (N3679, N3677);
and AND3 (N3680, N3675, N280, N2693);
nand NAND2 (N3681, N3670, N2700);
and AND3 (N3682, N3679, N223, N70);
not NOT1 (N3683, N3678);
buf BUF1 (N3684, N3650);
xor XOR2 (N3685, N3666, N172);
xor XOR2 (N3686, N3682, N2277);
buf BUF1 (N3687, N3681);
and AND3 (N3688, N3683, N167, N690);
or OR4 (N3689, N3687, N2476, N2055, N464);
and AND3 (N3690, N3676, N1705, N1150);
xor XOR2 (N3691, N3686, N2511);
nor NOR4 (N3692, N3685, N2888, N1995, N54);
nor NOR4 (N3693, N3691, N2076, N1265, N1340);
or OR2 (N3694, N3689, N1944);
or OR3 (N3695, N3688, N236, N553);
not NOT1 (N3696, N3674);
nand NAND2 (N3697, N3696, N2470);
or OR4 (N3698, N3693, N3522, N551, N1222);
nand NAND2 (N3699, N3694, N1092);
buf BUF1 (N3700, N3692);
not NOT1 (N3701, N3698);
buf BUF1 (N3702, N3700);
or OR3 (N3703, N3624, N3581, N476);
nand NAND3 (N3704, N3701, N1336, N248);
buf BUF1 (N3705, N3702);
buf BUF1 (N3706, N3697);
buf BUF1 (N3707, N3695);
or OR3 (N3708, N3684, N1214, N3164);
nor NOR2 (N3709, N3708, N2007);
nand NAND2 (N3710, N3663, N2954);
buf BUF1 (N3711, N3704);
nand NAND3 (N3712, N3705, N1541, N2273);
buf BUF1 (N3713, N3690);
not NOT1 (N3714, N3711);
and AND3 (N3715, N3680, N927, N2926);
nor NOR4 (N3716, N3715, N1636, N3613, N714);
or OR2 (N3717, N3699, N618);
nand NAND3 (N3718, N3713, N2925, N1213);
or OR4 (N3719, N3706, N50, N258, N3470);
nand NAND3 (N3720, N3712, N138, N1176);
nor NOR4 (N3721, N3718, N1610, N548, N2462);
or OR3 (N3722, N3716, N845, N932);
nor NOR2 (N3723, N3721, N806);
xor XOR2 (N3724, N3703, N2232);
and AND2 (N3725, N3707, N1202);
nor NOR2 (N3726, N3720, N2747);
nand NAND3 (N3727, N3717, N1174, N792);
xor XOR2 (N3728, N3709, N2064);
buf BUF1 (N3729, N3722);
nand NAND2 (N3730, N3719, N893);
buf BUF1 (N3731, N3730);
nor NOR4 (N3732, N3726, N649, N1208, N551);
nand NAND3 (N3733, N3727, N2646, N1056);
xor XOR2 (N3734, N3723, N2519);
not NOT1 (N3735, N3714);
nor NOR2 (N3736, N3733, N1855);
buf BUF1 (N3737, N3724);
nand NAND3 (N3738, N3736, N2378, N2474);
buf BUF1 (N3739, N3728);
buf BUF1 (N3740, N3710);
not NOT1 (N3741, N3734);
or OR3 (N3742, N3737, N818, N2110);
and AND3 (N3743, N3732, N1848, N1861);
nor NOR4 (N3744, N3731, N1373, N521, N3297);
not NOT1 (N3745, N3725);
nor NOR3 (N3746, N3740, N1509, N3501);
or OR2 (N3747, N3746, N1996);
nand NAND4 (N3748, N3745, N929, N2918, N3010);
not NOT1 (N3749, N3744);
buf BUF1 (N3750, N3742);
nand NAND2 (N3751, N3747, N585);
nand NAND4 (N3752, N3739, N1111, N2678, N1520);
nor NOR3 (N3753, N3748, N2922, N946);
nor NOR3 (N3754, N3752, N836, N2549);
not NOT1 (N3755, N3729);
not NOT1 (N3756, N3755);
nor NOR3 (N3757, N3735, N2406, N2910);
xor XOR2 (N3758, N3756, N317);
not NOT1 (N3759, N3753);
buf BUF1 (N3760, N3759);
not NOT1 (N3761, N3751);
nand NAND4 (N3762, N3741, N875, N504, N3236);
and AND2 (N3763, N3762, N2313);
not NOT1 (N3764, N3760);
and AND3 (N3765, N3764, N810, N1980);
xor XOR2 (N3766, N3749, N1682);
and AND4 (N3767, N3761, N1601, N1132, N3523);
not NOT1 (N3768, N3754);
nor NOR4 (N3769, N3743, N2617, N2536, N3322);
nor NOR2 (N3770, N3765, N1196);
nand NAND2 (N3771, N3763, N1483);
not NOT1 (N3772, N3757);
buf BUF1 (N3773, N3772);
xor XOR2 (N3774, N3768, N150);
not NOT1 (N3775, N3771);
xor XOR2 (N3776, N3775, N2018);
or OR3 (N3777, N3774, N2619, N3590);
buf BUF1 (N3778, N3758);
not NOT1 (N3779, N3738);
not NOT1 (N3780, N3769);
nor NOR4 (N3781, N3767, N2365, N2333, N455);
xor XOR2 (N3782, N3766, N1327);
or OR3 (N3783, N3778, N3045, N2050);
nor NOR3 (N3784, N3779, N1260, N254);
not NOT1 (N3785, N3782);
nand NAND2 (N3786, N3776, N30);
xor XOR2 (N3787, N3781, N508);
or OR3 (N3788, N3786, N1205, N2554);
nor NOR3 (N3789, N3780, N2525, N3624);
not NOT1 (N3790, N3788);
nand NAND4 (N3791, N3773, N1919, N57, N1321);
buf BUF1 (N3792, N3777);
xor XOR2 (N3793, N3785, N1943);
nand NAND3 (N3794, N3793, N3577, N3099);
nand NAND4 (N3795, N3770, N2481, N3080, N852);
and AND4 (N3796, N3791, N2880, N3587, N3065);
nor NOR2 (N3797, N3750, N1158);
or OR3 (N3798, N3795, N1460, N2535);
nor NOR2 (N3799, N3797, N701);
nor NOR4 (N3800, N3790, N1179, N3289, N2264);
nor NOR3 (N3801, N3800, N1046, N1529);
not NOT1 (N3802, N3789);
buf BUF1 (N3803, N3796);
nand NAND2 (N3804, N3802, N2449);
xor XOR2 (N3805, N3794, N1035);
buf BUF1 (N3806, N3799);
or OR3 (N3807, N3787, N1907, N1974);
xor XOR2 (N3808, N3783, N30);
not NOT1 (N3809, N3784);
nand NAND2 (N3810, N3798, N1036);
or OR2 (N3811, N3808, N640);
or OR3 (N3812, N3792, N1753, N1571);
not NOT1 (N3813, N3804);
nor NOR2 (N3814, N3811, N2892);
nor NOR2 (N3815, N3812, N2868);
or OR3 (N3816, N3807, N851, N916);
buf BUF1 (N3817, N3810);
nand NAND4 (N3818, N3803, N861, N3787, N1203);
and AND3 (N3819, N3806, N3212, N2143);
or OR3 (N3820, N3814, N3495, N1011);
buf BUF1 (N3821, N3819);
and AND2 (N3822, N3815, N1794);
not NOT1 (N3823, N3809);
buf BUF1 (N3824, N3818);
buf BUF1 (N3825, N3824);
or OR2 (N3826, N3813, N2641);
or OR2 (N3827, N3801, N2862);
nor NOR2 (N3828, N3822, N1299);
buf BUF1 (N3829, N3823);
and AND3 (N3830, N3816, N3039, N1873);
not NOT1 (N3831, N3817);
buf BUF1 (N3832, N3826);
xor XOR2 (N3833, N3832, N2820);
buf BUF1 (N3834, N3805);
nand NAND3 (N3835, N3833, N1517, N503);
xor XOR2 (N3836, N3827, N1710);
nand NAND3 (N3837, N3835, N366, N3786);
and AND4 (N3838, N3829, N130, N2532, N3460);
and AND4 (N3839, N3825, N192, N404, N2274);
nor NOR3 (N3840, N3834, N2973, N54);
nand NAND3 (N3841, N3840, N1566, N1467);
nand NAND4 (N3842, N3837, N2794, N2935, N2012);
or OR2 (N3843, N3830, N2481);
nand NAND3 (N3844, N3841, N2091, N1438);
and AND3 (N3845, N3836, N31, N2642);
nand NAND2 (N3846, N3831, N2939);
xor XOR2 (N3847, N3846, N1705);
not NOT1 (N3848, N3842);
xor XOR2 (N3849, N3820, N3014);
nand NAND2 (N3850, N3849, N3499);
not NOT1 (N3851, N3839);
nand NAND3 (N3852, N3838, N2681, N13);
and AND4 (N3853, N3828, N1144, N1723, N1193);
or OR4 (N3854, N3851, N2139, N946, N3816);
xor XOR2 (N3855, N3852, N3631);
not NOT1 (N3856, N3848);
nor NOR3 (N3857, N3847, N3755, N611);
not NOT1 (N3858, N3844);
not NOT1 (N3859, N3821);
not NOT1 (N3860, N3853);
not NOT1 (N3861, N3860);
nor NOR4 (N3862, N3856, N1028, N3290, N2007);
and AND2 (N3863, N3859, N3196);
buf BUF1 (N3864, N3862);
xor XOR2 (N3865, N3861, N1626);
nand NAND4 (N3866, N3855, N2594, N1406, N1269);
xor XOR2 (N3867, N3865, N24);
xor XOR2 (N3868, N3845, N3734);
xor XOR2 (N3869, N3863, N225);
or OR4 (N3870, N3857, N1225, N1190, N1182);
or OR2 (N3871, N3870, N3246);
not NOT1 (N3872, N3866);
and AND2 (N3873, N3871, N3131);
and AND2 (N3874, N3867, N2054);
xor XOR2 (N3875, N3874, N2039);
nand NAND4 (N3876, N3872, N853, N1130, N114);
or OR4 (N3877, N3873, N3686, N3759, N2489);
nor NOR3 (N3878, N3843, N2382, N3461);
nor NOR4 (N3879, N3850, N592, N3373, N2456);
not NOT1 (N3880, N3875);
and AND2 (N3881, N3879, N2649);
nor NOR3 (N3882, N3878, N2221, N2776);
not NOT1 (N3883, N3854);
nand NAND2 (N3884, N3868, N1171);
and AND3 (N3885, N3883, N3548, N1218);
xor XOR2 (N3886, N3858, N1106);
and AND3 (N3887, N3869, N2780, N641);
not NOT1 (N3888, N3884);
nor NOR2 (N3889, N3876, N2117);
or OR2 (N3890, N3886, N1182);
not NOT1 (N3891, N3889);
nand NAND2 (N3892, N3864, N3435);
xor XOR2 (N3893, N3877, N927);
xor XOR2 (N3894, N3887, N281);
nand NAND4 (N3895, N3893, N2176, N3014, N612);
not NOT1 (N3896, N3882);
and AND4 (N3897, N3895, N3013, N1298, N1900);
buf BUF1 (N3898, N3892);
and AND4 (N3899, N3888, N1258, N338, N731);
nand NAND3 (N3900, N3890, N2587, N3306);
nand NAND3 (N3901, N3881, N137, N3724);
nor NOR2 (N3902, N3891, N3392);
buf BUF1 (N3903, N3897);
or OR2 (N3904, N3903, N769);
and AND2 (N3905, N3900, N1826);
nor NOR2 (N3906, N3905, N3852);
nor NOR3 (N3907, N3906, N3399, N725);
nor NOR4 (N3908, N3902, N1148, N726, N3090);
buf BUF1 (N3909, N3904);
nand NAND3 (N3910, N3901, N1015, N1370);
nand NAND3 (N3911, N3908, N1469, N100);
nor NOR2 (N3912, N3880, N3524);
nand NAND4 (N3913, N3907, N1450, N2480, N1424);
buf BUF1 (N3914, N3913);
or OR4 (N3915, N3911, N2611, N159, N1122);
nand NAND4 (N3916, N3885, N1644, N3753, N291);
and AND2 (N3917, N3899, N1235);
buf BUF1 (N3918, N3917);
nor NOR4 (N3919, N3909, N2850, N1412, N3688);
buf BUF1 (N3920, N3915);
or OR2 (N3921, N3918, N2848);
or OR3 (N3922, N3896, N863, N633);
nand NAND3 (N3923, N3912, N176, N3391);
nor NOR2 (N3924, N3921, N14);
or OR2 (N3925, N3924, N1827);
or OR2 (N3926, N3920, N110);
or OR3 (N3927, N3898, N2297, N2693);
buf BUF1 (N3928, N3925);
nor NOR3 (N3929, N3894, N1707, N3404);
nand NAND2 (N3930, N3927, N85);
not NOT1 (N3931, N3929);
and AND2 (N3932, N3919, N3031);
nor NOR4 (N3933, N3916, N2533, N793, N2837);
nor NOR3 (N3934, N3930, N2456, N995);
nor NOR2 (N3935, N3910, N2249);
nor NOR2 (N3936, N3935, N1860);
buf BUF1 (N3937, N3934);
buf BUF1 (N3938, N3922);
not NOT1 (N3939, N3923);
or OR3 (N3940, N3939, N2136, N1657);
nor NOR2 (N3941, N3940, N1334);
buf BUF1 (N3942, N3937);
or OR4 (N3943, N3941, N3852, N1586, N2906);
nand NAND3 (N3944, N3914, N251, N3487);
buf BUF1 (N3945, N3933);
buf BUF1 (N3946, N3936);
not NOT1 (N3947, N3932);
or OR2 (N3948, N3926, N198);
not NOT1 (N3949, N3945);
xor XOR2 (N3950, N3946, N2314);
and AND3 (N3951, N3942, N1391, N664);
and AND3 (N3952, N3931, N1355, N1952);
buf BUF1 (N3953, N3949);
buf BUF1 (N3954, N3950);
not NOT1 (N3955, N3953);
nor NOR2 (N3956, N3952, N1991);
not NOT1 (N3957, N3943);
xor XOR2 (N3958, N3954, N3154);
and AND4 (N3959, N3947, N1032, N1889, N3487);
or OR3 (N3960, N3958, N1265, N3401);
xor XOR2 (N3961, N3948, N1464);
nor NOR2 (N3962, N3957, N3259);
and AND3 (N3963, N3938, N3804, N2101);
nor NOR4 (N3964, N3951, N861, N742, N2187);
nor NOR3 (N3965, N3955, N2309, N3234);
not NOT1 (N3966, N3961);
xor XOR2 (N3967, N3956, N263);
xor XOR2 (N3968, N3960, N410);
buf BUF1 (N3969, N3964);
nand NAND4 (N3970, N3967, N3293, N185, N1663);
xor XOR2 (N3971, N3944, N3498);
or OR4 (N3972, N3969, N3782, N1040, N1862);
xor XOR2 (N3973, N3972, N1291);
nor NOR4 (N3974, N3965, N2304, N3343, N3143);
or OR4 (N3975, N3971, N804, N2564, N1605);
not NOT1 (N3976, N3975);
or OR4 (N3977, N3928, N12, N2050, N2354);
and AND4 (N3978, N3977, N2659, N340, N577);
or OR3 (N3979, N3959, N1251, N2533);
buf BUF1 (N3980, N3963);
xor XOR2 (N3981, N3962, N3801);
or OR4 (N3982, N3966, N789, N1418, N1351);
or OR3 (N3983, N3970, N3292, N3909);
nand NAND3 (N3984, N3979, N1242, N1566);
or OR4 (N3985, N3976, N769, N1124, N3412);
buf BUF1 (N3986, N3980);
nor NOR4 (N3987, N3978, N916, N936, N2516);
nand NAND3 (N3988, N3984, N3438, N809);
and AND3 (N3989, N3985, N2921, N2205);
or OR2 (N3990, N3983, N2169);
or OR3 (N3991, N3982, N2001, N2328);
nand NAND4 (N3992, N3988, N1504, N126, N1080);
nor NOR4 (N3993, N3987, N2676, N2915, N3745);
and AND3 (N3994, N3991, N752, N3844);
and AND2 (N3995, N3974, N83);
or OR3 (N3996, N3990, N325, N226);
nor NOR4 (N3997, N3968, N415, N2628, N1975);
not NOT1 (N3998, N3992);
buf BUF1 (N3999, N3997);
not NOT1 (N4000, N3996);
not NOT1 (N4001, N3986);
xor XOR2 (N4002, N3973, N2899);
buf BUF1 (N4003, N3995);
or OR2 (N4004, N3994, N3591);
buf BUF1 (N4005, N4001);
or OR4 (N4006, N4000, N315, N3967, N1225);
nand NAND2 (N4007, N3989, N2193);
nand NAND3 (N4008, N4004, N3329, N2718);
or OR4 (N4009, N4003, N3968, N2800, N2);
nand NAND4 (N4010, N3993, N2102, N2337, N872);
or OR2 (N4011, N3998, N3432);
and AND3 (N4012, N3981, N1990, N3524);
nor NOR2 (N4013, N3999, N2017);
nand NAND4 (N4014, N4013, N2726, N3496, N538);
buf BUF1 (N4015, N4014);
and AND3 (N4016, N4002, N1881, N536);
endmodule