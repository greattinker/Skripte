// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N16001,N16003,N16008,N16009,N15993,N16010,N15999,N15958,N16002,N16011;

buf BUF1 (N12, N1);
nor NOR4 (N13, N10, N4, N9, N12);
and AND4 (N14, N13, N13, N7, N6);
nand NAND2 (N15, N14, N14);
and AND3 (N16, N10, N4, N13);
nand NAND3 (N17, N12, N12, N12);
and AND4 (N18, N9, N14, N6, N1);
buf BUF1 (N19, N9);
or OR2 (N20, N9, N7);
and AND2 (N21, N7, N17);
or OR3 (N22, N20, N21, N8);
not NOT1 (N23, N3);
or OR4 (N24, N19, N10, N7, N3);
buf BUF1 (N25, N1);
or OR4 (N26, N21, N13, N3, N13);
buf BUF1 (N27, N16);
xor XOR2 (N28, N9, N14);
xor XOR2 (N29, N19, N8);
nand NAND3 (N30, N28, N7, N14);
nand NAND4 (N31, N18, N20, N16, N26);
buf BUF1 (N32, N21);
and AND2 (N33, N24, N32);
or OR3 (N34, N23, N26, N21);
or OR2 (N35, N16, N1);
xor XOR2 (N36, N22, N20);
not NOT1 (N37, N31);
nor NOR2 (N38, N34, N22);
nor NOR2 (N39, N29, N26);
xor XOR2 (N40, N30, N24);
and AND2 (N41, N36, N18);
nor NOR4 (N42, N15, N1, N13, N31);
not NOT1 (N43, N38);
and AND3 (N44, N25, N2, N33);
xor XOR2 (N45, N13, N26);
and AND3 (N46, N37, N27, N22);
or OR3 (N47, N24, N15, N4);
buf BUF1 (N48, N46);
nor NOR2 (N49, N41, N22);
nor NOR2 (N50, N49, N30);
and AND3 (N51, N50, N30, N27);
or OR4 (N52, N39, N34, N7, N38);
buf BUF1 (N53, N42);
nor NOR2 (N54, N51, N38);
nor NOR3 (N55, N52, N16, N42);
xor XOR2 (N56, N47, N21);
nor NOR2 (N57, N35, N38);
not NOT1 (N58, N45);
nor NOR2 (N59, N53, N16);
buf BUF1 (N60, N40);
or OR2 (N61, N57, N26);
or OR4 (N62, N58, N32, N3, N24);
not NOT1 (N63, N61);
nand NAND3 (N64, N63, N35, N3);
and AND4 (N65, N64, N53, N27, N23);
nand NAND3 (N66, N55, N2, N30);
and AND3 (N67, N66, N41, N48);
nand NAND2 (N68, N27, N67);
xor XOR2 (N69, N11, N57);
buf BUF1 (N70, N68);
and AND2 (N71, N43, N70);
nor NOR4 (N72, N50, N39, N32, N4);
nor NOR2 (N73, N44, N20);
or OR2 (N74, N56, N3);
buf BUF1 (N75, N72);
or OR3 (N76, N62, N37, N9);
and AND2 (N77, N74, N45);
not NOT1 (N78, N76);
nor NOR3 (N79, N60, N32, N42);
not NOT1 (N80, N54);
xor XOR2 (N81, N59, N15);
nor NOR2 (N82, N81, N41);
or OR3 (N83, N69, N6, N52);
and AND2 (N84, N65, N83);
xor XOR2 (N85, N19, N36);
or OR3 (N86, N71, N51, N29);
xor XOR2 (N87, N80, N50);
buf BUF1 (N88, N77);
or OR2 (N89, N85, N83);
nor NOR2 (N90, N84, N85);
xor XOR2 (N91, N73, N60);
or OR4 (N92, N91, N45, N44, N52);
xor XOR2 (N93, N88, N55);
nor NOR2 (N94, N92, N63);
buf BUF1 (N95, N87);
nand NAND2 (N96, N86, N32);
nand NAND3 (N97, N75, N11, N15);
or OR2 (N98, N95, N95);
nor NOR2 (N99, N94, N52);
nand NAND3 (N100, N78, N30, N26);
xor XOR2 (N101, N99, N82);
or OR4 (N102, N55, N39, N78, N73);
not NOT1 (N103, N89);
nand NAND4 (N104, N97, N15, N34, N98);
or OR4 (N105, N44, N95, N96, N1);
nor NOR4 (N106, N29, N62, N12, N82);
buf BUF1 (N107, N102);
xor XOR2 (N108, N90, N6);
nand NAND2 (N109, N101, N59);
or OR4 (N110, N106, N13, N93, N96);
and AND4 (N111, N73, N5, N104, N1);
not NOT1 (N112, N70);
nor NOR4 (N113, N110, N77, N13, N104);
xor XOR2 (N114, N103, N12);
and AND4 (N115, N114, N92, N52, N9);
or OR4 (N116, N109, N68, N32, N13);
nor NOR4 (N117, N107, N57, N4, N71);
nor NOR4 (N118, N115, N117, N44, N95);
not NOT1 (N119, N113);
or OR4 (N120, N25, N34, N69, N48);
buf BUF1 (N121, N120);
xor XOR2 (N122, N108, N90);
xor XOR2 (N123, N100, N86);
nor NOR2 (N124, N116, N33);
and AND3 (N125, N79, N113, N7);
nor NOR3 (N126, N119, N83, N74);
nand NAND3 (N127, N125, N12, N122);
or OR3 (N128, N14, N7, N120);
xor XOR2 (N129, N111, N41);
and AND4 (N130, N118, N119, N15, N100);
and AND3 (N131, N128, N52, N59);
xor XOR2 (N132, N129, N128);
and AND2 (N133, N130, N56);
nand NAND4 (N134, N132, N73, N66, N99);
nand NAND4 (N135, N133, N92, N127, N38);
nor NOR4 (N136, N40, N37, N105, N110);
buf BUF1 (N137, N122);
nor NOR3 (N138, N136, N54, N91);
or OR3 (N139, N121, N107, N1);
and AND2 (N140, N123, N122);
nand NAND2 (N141, N138, N86);
or OR4 (N142, N137, N24, N8, N105);
buf BUF1 (N143, N139);
xor XOR2 (N144, N142, N14);
nor NOR2 (N145, N140, N110);
and AND3 (N146, N134, N21, N22);
and AND3 (N147, N135, N74, N45);
xor XOR2 (N148, N141, N10);
and AND3 (N149, N145, N71, N15);
nor NOR2 (N150, N149, N149);
xor XOR2 (N151, N148, N132);
not NOT1 (N152, N126);
buf BUF1 (N153, N112);
and AND4 (N154, N146, N122, N132, N81);
and AND4 (N155, N147, N136, N151, N56);
not NOT1 (N156, N126);
and AND2 (N157, N150, N30);
xor XOR2 (N158, N143, N27);
nand NAND4 (N159, N144, N91, N4, N125);
not NOT1 (N160, N155);
buf BUF1 (N161, N154);
and AND2 (N162, N160, N134);
and AND3 (N163, N159, N52, N23);
and AND2 (N164, N161, N61);
buf BUF1 (N165, N157);
or OR2 (N166, N162, N146);
nand NAND4 (N167, N165, N95, N54, N35);
nand NAND2 (N168, N124, N13);
or OR3 (N169, N164, N50, N118);
nor NOR4 (N170, N152, N90, N121, N97);
nor NOR4 (N171, N163, N23, N114, N108);
buf BUF1 (N172, N166);
buf BUF1 (N173, N158);
nor NOR3 (N174, N153, N172, N63);
nor NOR2 (N175, N99, N49);
and AND4 (N176, N170, N47, N64, N77);
or OR3 (N177, N176, N145, N127);
not NOT1 (N178, N173);
not NOT1 (N179, N177);
nand NAND2 (N180, N168, N114);
nand NAND4 (N181, N180, N25, N66, N115);
or OR3 (N182, N181, N63, N179);
or OR4 (N183, N5, N99, N158, N179);
or OR4 (N184, N156, N20, N95, N183);
nor NOR4 (N185, N41, N111, N34, N164);
nand NAND2 (N186, N182, N112);
not NOT1 (N187, N169);
not NOT1 (N188, N187);
xor XOR2 (N189, N174, N133);
or OR3 (N190, N131, N147, N93);
nand NAND2 (N191, N186, N159);
xor XOR2 (N192, N185, N1);
or OR2 (N193, N171, N168);
nor NOR3 (N194, N190, N124, N151);
xor XOR2 (N195, N189, N189);
and AND3 (N196, N188, N169, N43);
buf BUF1 (N197, N192);
or OR3 (N198, N167, N169, N118);
not NOT1 (N199, N198);
nand NAND2 (N200, N199, N195);
xor XOR2 (N201, N165, N93);
nor NOR2 (N202, N175, N122);
nand NAND2 (N203, N194, N36);
buf BUF1 (N204, N196);
and AND3 (N205, N201, N8, N167);
nor NOR4 (N206, N178, N175, N23, N94);
nor NOR2 (N207, N193, N164);
or OR4 (N208, N203, N27, N27, N123);
buf BUF1 (N209, N206);
not NOT1 (N210, N205);
not NOT1 (N211, N197);
and AND2 (N212, N207, N27);
or OR3 (N213, N202, N82, N58);
and AND2 (N214, N211, N104);
and AND3 (N215, N209, N67, N142);
or OR2 (N216, N204, N158);
not NOT1 (N217, N184);
nor NOR4 (N218, N215, N202, N83, N108);
nor NOR2 (N219, N214, N127);
not NOT1 (N220, N218);
buf BUF1 (N221, N210);
nand NAND4 (N222, N216, N47, N102, N47);
buf BUF1 (N223, N221);
buf BUF1 (N224, N219);
nand NAND2 (N225, N208, N35);
not NOT1 (N226, N217);
nor NOR2 (N227, N213, N64);
nor NOR2 (N228, N191, N116);
xor XOR2 (N229, N225, N185);
buf BUF1 (N230, N212);
nor NOR3 (N231, N230, N140, N59);
buf BUF1 (N232, N228);
or OR4 (N233, N224, N24, N3, N45);
xor XOR2 (N234, N231, N61);
nor NOR2 (N235, N232, N170);
not NOT1 (N236, N227);
buf BUF1 (N237, N222);
xor XOR2 (N238, N226, N77);
not NOT1 (N239, N220);
not NOT1 (N240, N223);
xor XOR2 (N241, N239, N29);
or OR4 (N242, N237, N156, N13, N176);
xor XOR2 (N243, N240, N210);
nand NAND4 (N244, N234, N21, N40, N215);
buf BUF1 (N245, N235);
nor NOR4 (N246, N236, N6, N88, N24);
not NOT1 (N247, N244);
nor NOR4 (N248, N243, N98, N230, N75);
and AND4 (N249, N248, N161, N90, N20);
and AND4 (N250, N245, N95, N219, N154);
or OR2 (N251, N241, N191);
nor NOR2 (N252, N242, N206);
and AND3 (N253, N250, N115, N25);
and AND2 (N254, N253, N85);
or OR4 (N255, N254, N227, N185, N71);
buf BUF1 (N256, N229);
and AND2 (N257, N233, N169);
nand NAND2 (N258, N247, N22);
nand NAND2 (N259, N257, N98);
xor XOR2 (N260, N258, N77);
nor NOR4 (N261, N246, N142, N150, N87);
or OR4 (N262, N249, N69, N233, N92);
and AND4 (N263, N262, N146, N254, N219);
nor NOR4 (N264, N255, N31, N65, N70);
xor XOR2 (N265, N261, N42);
buf BUF1 (N266, N264);
nor NOR3 (N267, N238, N250, N49);
buf BUF1 (N268, N251);
nand NAND4 (N269, N259, N206, N80, N202);
and AND3 (N270, N265, N137, N33);
and AND4 (N271, N267, N48, N40, N247);
nand NAND4 (N272, N252, N228, N6, N132);
not NOT1 (N273, N256);
or OR2 (N274, N273, N51);
nand NAND2 (N275, N266, N148);
or OR2 (N276, N200, N151);
and AND3 (N277, N260, N174, N253);
nand NAND3 (N278, N263, N61, N102);
not NOT1 (N279, N276);
nand NAND3 (N280, N272, N6, N124);
nand NAND4 (N281, N278, N121, N14, N190);
or OR4 (N282, N268, N76, N90, N149);
not NOT1 (N283, N279);
nand NAND3 (N284, N280, N187, N55);
and AND4 (N285, N269, N63, N261, N165);
not NOT1 (N286, N275);
xor XOR2 (N287, N274, N19);
nand NAND4 (N288, N283, N5, N146, N20);
xor XOR2 (N289, N277, N153);
nand NAND2 (N290, N287, N5);
xor XOR2 (N291, N289, N44);
or OR3 (N292, N271, N192, N72);
not NOT1 (N293, N282);
nand NAND3 (N294, N286, N233, N119);
xor XOR2 (N295, N290, N258);
nor NOR3 (N296, N285, N209, N101);
buf BUF1 (N297, N281);
nor NOR2 (N298, N284, N36);
and AND4 (N299, N298, N232, N225, N110);
nor NOR3 (N300, N291, N206, N270);
nand NAND3 (N301, N280, N3, N14);
xor XOR2 (N302, N293, N300);
buf BUF1 (N303, N241);
xor XOR2 (N304, N299, N300);
or OR4 (N305, N288, N55, N166, N106);
or OR3 (N306, N294, N267, N188);
nor NOR3 (N307, N303, N90, N63);
or OR3 (N308, N295, N60, N46);
nor NOR3 (N309, N302, N211, N201);
not NOT1 (N310, N305);
not NOT1 (N311, N297);
or OR4 (N312, N309, N89, N41, N37);
not NOT1 (N313, N304);
or OR4 (N314, N308, N28, N173, N276);
or OR2 (N315, N296, N64);
buf BUF1 (N316, N301);
not NOT1 (N317, N310);
and AND4 (N318, N311, N317, N83, N299);
and AND4 (N319, N311, N279, N65, N253);
nand NAND2 (N320, N313, N6);
buf BUF1 (N321, N307);
buf BUF1 (N322, N315);
xor XOR2 (N323, N312, N20);
or OR3 (N324, N321, N161, N304);
and AND2 (N325, N306, N60);
xor XOR2 (N326, N324, N319);
and AND2 (N327, N239, N219);
and AND4 (N328, N316, N71, N192, N282);
buf BUF1 (N329, N326);
nand NAND3 (N330, N292, N83, N36);
or OR3 (N331, N318, N163, N316);
xor XOR2 (N332, N314, N134);
and AND3 (N333, N329, N156, N47);
buf BUF1 (N334, N325);
and AND4 (N335, N331, N23, N114, N209);
or OR4 (N336, N332, N124, N151, N312);
nand NAND2 (N337, N334, N144);
xor XOR2 (N338, N320, N291);
xor XOR2 (N339, N336, N199);
and AND4 (N340, N333, N142, N26, N110);
nand NAND3 (N341, N335, N264, N22);
nand NAND4 (N342, N338, N145, N175, N128);
not NOT1 (N343, N337);
buf BUF1 (N344, N330);
or OR2 (N345, N340, N215);
not NOT1 (N346, N339);
nor NOR4 (N347, N328, N155, N227, N183);
or OR4 (N348, N342, N126, N25, N217);
or OR3 (N349, N347, N179, N237);
nor NOR3 (N350, N323, N154, N248);
not NOT1 (N351, N348);
or OR2 (N352, N343, N123);
not NOT1 (N353, N345);
nor NOR3 (N354, N353, N47, N224);
not NOT1 (N355, N344);
buf BUF1 (N356, N350);
nand NAND2 (N357, N355, N2);
buf BUF1 (N358, N357);
or OR3 (N359, N327, N252, N82);
nand NAND2 (N360, N356, N313);
xor XOR2 (N361, N359, N102);
or OR4 (N362, N354, N92, N287, N299);
or OR2 (N363, N352, N77);
and AND2 (N364, N358, N92);
or OR4 (N365, N364, N199, N7, N66);
nand NAND4 (N366, N346, N303, N275, N356);
not NOT1 (N367, N349);
nor NOR4 (N368, N341, N133, N78, N15);
xor XOR2 (N369, N367, N163);
buf BUF1 (N370, N363);
buf BUF1 (N371, N370);
not NOT1 (N372, N369);
buf BUF1 (N373, N372);
xor XOR2 (N374, N362, N18);
nor NOR4 (N375, N360, N201, N333, N320);
not NOT1 (N376, N366);
buf BUF1 (N377, N351);
buf BUF1 (N378, N373);
buf BUF1 (N379, N375);
xor XOR2 (N380, N376, N134);
buf BUF1 (N381, N379);
not NOT1 (N382, N377);
nand NAND3 (N383, N381, N162, N131);
not NOT1 (N384, N383);
nand NAND4 (N385, N365, N348, N328, N262);
not NOT1 (N386, N368);
or OR2 (N387, N385, N298);
buf BUF1 (N388, N380);
nor NOR2 (N389, N371, N235);
nor NOR4 (N390, N361, N68, N271, N136);
not NOT1 (N391, N384);
buf BUF1 (N392, N374);
xor XOR2 (N393, N386, N374);
nand NAND2 (N394, N390, N90);
or OR3 (N395, N393, N317, N354);
not NOT1 (N396, N378);
not NOT1 (N397, N382);
buf BUF1 (N398, N392);
or OR2 (N399, N396, N41);
or OR4 (N400, N388, N368, N218, N315);
not NOT1 (N401, N322);
buf BUF1 (N402, N395);
not NOT1 (N403, N394);
nor NOR3 (N404, N400, N180, N231);
xor XOR2 (N405, N391, N37);
xor XOR2 (N406, N401, N109);
buf BUF1 (N407, N405);
not NOT1 (N408, N398);
not NOT1 (N409, N397);
xor XOR2 (N410, N404, N126);
not NOT1 (N411, N399);
not NOT1 (N412, N402);
nor NOR3 (N413, N407, N189, N87);
and AND3 (N414, N387, N69, N354);
or OR3 (N415, N409, N137, N395);
or OR4 (N416, N406, N371, N88, N291);
or OR2 (N417, N416, N137);
and AND4 (N418, N410, N347, N2, N291);
or OR4 (N419, N411, N285, N13, N294);
not NOT1 (N420, N419);
nor NOR4 (N421, N412, N27, N147, N330);
nor NOR4 (N422, N415, N295, N344, N349);
xor XOR2 (N423, N421, N222);
nor NOR2 (N424, N418, N336);
buf BUF1 (N425, N413);
or OR4 (N426, N424, N417, N368, N298);
or OR3 (N427, N148, N267, N400);
buf BUF1 (N428, N414);
nand NAND2 (N429, N423, N13);
not NOT1 (N430, N408);
and AND4 (N431, N427, N402, N253, N134);
and AND3 (N432, N430, N324, N149);
nand NAND2 (N433, N403, N419);
not NOT1 (N434, N425);
buf BUF1 (N435, N429);
nand NAND3 (N436, N431, N354, N296);
not NOT1 (N437, N433);
nor NOR2 (N438, N436, N386);
buf BUF1 (N439, N426);
xor XOR2 (N440, N435, N92);
xor XOR2 (N441, N434, N199);
or OR3 (N442, N389, N109, N49);
nand NAND4 (N443, N428, N419, N70, N226);
and AND4 (N444, N437, N210, N84, N125);
xor XOR2 (N445, N420, N311);
nand NAND4 (N446, N443, N284, N246, N335);
nor NOR3 (N447, N422, N440, N194);
nand NAND2 (N448, N401, N199);
and AND2 (N449, N432, N132);
buf BUF1 (N450, N448);
nor NOR2 (N451, N444, N102);
nor NOR2 (N452, N445, N4);
buf BUF1 (N453, N446);
nand NAND3 (N454, N441, N128, N42);
not NOT1 (N455, N449);
xor XOR2 (N456, N439, N97);
nor NOR3 (N457, N456, N351, N220);
nor NOR2 (N458, N454, N454);
or OR2 (N459, N453, N368);
nor NOR2 (N460, N455, N282);
xor XOR2 (N461, N458, N153);
xor XOR2 (N462, N438, N244);
or OR2 (N463, N447, N447);
not NOT1 (N464, N462);
buf BUF1 (N465, N452);
xor XOR2 (N466, N451, N171);
nor NOR3 (N467, N460, N192, N461);
buf BUF1 (N468, N125);
buf BUF1 (N469, N465);
nand NAND3 (N470, N469, N181, N86);
nor NOR2 (N471, N466, N264);
buf BUF1 (N472, N463);
nor NOR2 (N473, N467, N33);
or OR3 (N474, N468, N246, N104);
xor XOR2 (N475, N473, N287);
not NOT1 (N476, N457);
not NOT1 (N477, N472);
or OR2 (N478, N476, N281);
and AND3 (N479, N459, N407, N178);
nand NAND2 (N480, N477, N124);
and AND4 (N481, N474, N29, N389, N82);
xor XOR2 (N482, N470, N302);
and AND2 (N483, N478, N266);
not NOT1 (N484, N475);
buf BUF1 (N485, N442);
nand NAND2 (N486, N479, N296);
nand NAND3 (N487, N464, N402, N346);
nor NOR2 (N488, N485, N445);
and AND4 (N489, N480, N370, N291, N181);
buf BUF1 (N490, N483);
and AND4 (N491, N486, N148, N327, N434);
or OR2 (N492, N491, N388);
nand NAND2 (N493, N471, N374);
nand NAND2 (N494, N481, N44);
nand NAND3 (N495, N487, N473, N172);
not NOT1 (N496, N489);
buf BUF1 (N497, N493);
xor XOR2 (N498, N490, N211);
or OR2 (N499, N488, N281);
or OR2 (N500, N482, N200);
buf BUF1 (N501, N484);
buf BUF1 (N502, N496);
xor XOR2 (N503, N501, N81);
buf BUF1 (N504, N492);
nor NOR4 (N505, N502, N267, N425, N305);
nor NOR3 (N506, N494, N281, N442);
and AND3 (N507, N499, N226, N501);
xor XOR2 (N508, N503, N386);
not NOT1 (N509, N497);
buf BUF1 (N510, N495);
buf BUF1 (N511, N506);
not NOT1 (N512, N500);
buf BUF1 (N513, N504);
xor XOR2 (N514, N512, N440);
nand NAND3 (N515, N510, N476, N328);
nand NAND3 (N516, N505, N227, N327);
and AND2 (N517, N514, N107);
xor XOR2 (N518, N508, N3);
not NOT1 (N519, N498);
buf BUF1 (N520, N518);
nand NAND2 (N521, N509, N187);
xor XOR2 (N522, N517, N186);
buf BUF1 (N523, N520);
or OR4 (N524, N450, N78, N321, N263);
not NOT1 (N525, N515);
and AND4 (N526, N507, N390, N127, N497);
and AND3 (N527, N519, N171, N106);
or OR4 (N528, N522, N8, N167, N3);
not NOT1 (N529, N511);
and AND4 (N530, N513, N443, N183, N16);
buf BUF1 (N531, N525);
or OR4 (N532, N529, N278, N394, N215);
buf BUF1 (N533, N523);
nand NAND2 (N534, N516, N38);
xor XOR2 (N535, N530, N171);
and AND4 (N536, N532, N438, N381, N43);
xor XOR2 (N537, N534, N5);
buf BUF1 (N538, N526);
nand NAND4 (N539, N533, N239, N455, N104);
xor XOR2 (N540, N528, N178);
nand NAND2 (N541, N540, N266);
and AND3 (N542, N541, N287, N425);
nand NAND3 (N543, N524, N217, N272);
or OR2 (N544, N537, N389);
or OR3 (N545, N531, N453, N324);
nor NOR3 (N546, N542, N539, N543);
nand NAND2 (N547, N315, N60);
or OR3 (N548, N85, N290, N142);
xor XOR2 (N549, N527, N175);
nor NOR4 (N550, N547, N344, N318, N29);
xor XOR2 (N551, N535, N144);
or OR2 (N552, N549, N434);
nor NOR2 (N553, N546, N540);
buf BUF1 (N554, N548);
xor XOR2 (N555, N554, N75);
or OR4 (N556, N555, N53, N404, N223);
not NOT1 (N557, N551);
xor XOR2 (N558, N552, N210);
xor XOR2 (N559, N553, N297);
xor XOR2 (N560, N544, N148);
xor XOR2 (N561, N550, N368);
or OR2 (N562, N560, N8);
or OR2 (N563, N538, N395);
or OR2 (N564, N561, N436);
xor XOR2 (N565, N562, N96);
or OR4 (N566, N556, N250, N316, N549);
xor XOR2 (N567, N559, N41);
or OR4 (N568, N563, N516, N153, N74);
and AND3 (N569, N557, N73, N464);
and AND3 (N570, N565, N130, N390);
nand NAND3 (N571, N545, N291, N291);
and AND3 (N572, N568, N333, N185);
nand NAND4 (N573, N536, N23, N323, N109);
and AND2 (N574, N569, N327);
xor XOR2 (N575, N558, N372);
or OR2 (N576, N521, N480);
buf BUF1 (N577, N575);
and AND3 (N578, N564, N124, N102);
xor XOR2 (N579, N570, N574);
xor XOR2 (N580, N502, N441);
xor XOR2 (N581, N572, N363);
nor NOR3 (N582, N579, N283, N126);
buf BUF1 (N583, N567);
xor XOR2 (N584, N573, N395);
xor XOR2 (N585, N571, N223);
nor NOR2 (N586, N581, N227);
or OR2 (N587, N582, N291);
or OR2 (N588, N576, N247);
nor NOR2 (N589, N587, N275);
nor NOR2 (N590, N585, N412);
nand NAND2 (N591, N566, N271);
xor XOR2 (N592, N590, N429);
xor XOR2 (N593, N592, N503);
nor NOR4 (N594, N580, N425, N32, N298);
or OR4 (N595, N583, N342, N525, N149);
buf BUF1 (N596, N586);
nor NOR2 (N597, N589, N11);
or OR4 (N598, N594, N472, N175, N292);
and AND4 (N599, N588, N344, N545, N552);
or OR3 (N600, N597, N460, N238);
nor NOR2 (N601, N584, N460);
xor XOR2 (N602, N578, N530);
nand NAND2 (N603, N596, N366);
not NOT1 (N604, N603);
not NOT1 (N605, N577);
xor XOR2 (N606, N601, N490);
xor XOR2 (N607, N602, N441);
not NOT1 (N608, N606);
not NOT1 (N609, N599);
and AND3 (N610, N608, N436, N140);
not NOT1 (N611, N605);
not NOT1 (N612, N593);
xor XOR2 (N613, N604, N431);
buf BUF1 (N614, N612);
and AND4 (N615, N607, N32, N142, N339);
nor NOR3 (N616, N613, N390, N104);
xor XOR2 (N617, N615, N223);
not NOT1 (N618, N591);
buf BUF1 (N619, N609);
nand NAND3 (N620, N610, N340, N587);
nor NOR2 (N621, N598, N366);
nand NAND3 (N622, N619, N106, N498);
nor NOR4 (N623, N622, N596, N428, N169);
nand NAND3 (N624, N623, N384, N372);
or OR4 (N625, N595, N295, N483, N173);
not NOT1 (N626, N624);
and AND3 (N627, N626, N101, N202);
xor XOR2 (N628, N611, N89);
buf BUF1 (N629, N600);
nand NAND4 (N630, N620, N168, N34, N300);
xor XOR2 (N631, N616, N595);
nand NAND2 (N632, N631, N485);
not NOT1 (N633, N614);
nand NAND2 (N634, N618, N630);
not NOT1 (N635, N407);
and AND2 (N636, N634, N325);
not NOT1 (N637, N617);
not NOT1 (N638, N628);
xor XOR2 (N639, N632, N344);
nor NOR4 (N640, N629, N18, N518, N34);
and AND4 (N641, N621, N485, N486, N633);
and AND3 (N642, N418, N463, N70);
not NOT1 (N643, N636);
or OR4 (N644, N642, N379, N216, N43);
nor NOR4 (N645, N627, N185, N296, N480);
nand NAND3 (N646, N639, N437, N423);
xor XOR2 (N647, N625, N608);
not NOT1 (N648, N646);
and AND3 (N649, N641, N21, N548);
buf BUF1 (N650, N637);
xor XOR2 (N651, N640, N632);
nand NAND4 (N652, N643, N547, N250, N614);
or OR2 (N653, N652, N210);
or OR4 (N654, N638, N491, N594, N37);
not NOT1 (N655, N649);
not NOT1 (N656, N651);
and AND4 (N657, N648, N88, N622, N81);
nand NAND4 (N658, N655, N594, N305, N480);
nor NOR2 (N659, N658, N560);
buf BUF1 (N660, N650);
nor NOR2 (N661, N654, N633);
and AND3 (N662, N653, N112, N27);
nand NAND3 (N663, N644, N450, N188);
nand NAND2 (N664, N656, N179);
and AND4 (N665, N664, N124, N468, N657);
xor XOR2 (N666, N89, N35);
xor XOR2 (N667, N665, N158);
xor XOR2 (N668, N666, N92);
buf BUF1 (N669, N645);
not NOT1 (N670, N659);
not NOT1 (N671, N635);
xor XOR2 (N672, N667, N623);
and AND4 (N673, N663, N589, N25, N459);
xor XOR2 (N674, N670, N598);
not NOT1 (N675, N661);
or OR4 (N676, N675, N535, N1, N73);
nand NAND4 (N677, N674, N609, N346, N229);
buf BUF1 (N678, N660);
or OR2 (N679, N647, N519);
or OR3 (N680, N676, N352, N321);
xor XOR2 (N681, N672, N41);
not NOT1 (N682, N671);
buf BUF1 (N683, N680);
nor NOR4 (N684, N681, N407, N406, N546);
not NOT1 (N685, N678);
buf BUF1 (N686, N685);
or OR4 (N687, N668, N237, N353, N576);
xor XOR2 (N688, N686, N35);
not NOT1 (N689, N682);
not NOT1 (N690, N673);
or OR4 (N691, N688, N234, N680, N562);
buf BUF1 (N692, N683);
xor XOR2 (N693, N662, N37);
not NOT1 (N694, N684);
nor NOR2 (N695, N689, N639);
not NOT1 (N696, N679);
xor XOR2 (N697, N691, N413);
nand NAND3 (N698, N695, N259, N292);
buf BUF1 (N699, N696);
buf BUF1 (N700, N698);
nand NAND4 (N701, N700, N243, N507, N109);
nand NAND2 (N702, N677, N329);
nor NOR4 (N703, N701, N450, N144, N111);
xor XOR2 (N704, N697, N577);
xor XOR2 (N705, N687, N703);
nand NAND2 (N706, N205, N648);
nor NOR2 (N707, N704, N105);
nand NAND3 (N708, N669, N696, N332);
and AND4 (N709, N707, N544, N481, N611);
buf BUF1 (N710, N705);
nand NAND2 (N711, N709, N127);
nand NAND2 (N712, N699, N295);
xor XOR2 (N713, N708, N164);
and AND2 (N714, N702, N444);
xor XOR2 (N715, N712, N307);
nor NOR4 (N716, N690, N158, N659, N326);
nor NOR4 (N717, N694, N538, N443, N239);
not NOT1 (N718, N693);
not NOT1 (N719, N706);
nand NAND2 (N720, N715, N21);
nand NAND3 (N721, N711, N561, N372);
buf BUF1 (N722, N719);
not NOT1 (N723, N710);
or OR2 (N724, N723, N528);
nand NAND3 (N725, N721, N95, N164);
nand NAND4 (N726, N724, N628, N205, N298);
nand NAND3 (N727, N692, N322, N52);
and AND4 (N728, N714, N365, N572, N435);
and AND2 (N729, N718, N582);
or OR3 (N730, N728, N542, N487);
nand NAND3 (N731, N713, N336, N152);
and AND2 (N732, N725, N224);
not NOT1 (N733, N716);
buf BUF1 (N734, N722);
nor NOR3 (N735, N734, N569, N166);
nand NAND4 (N736, N733, N349, N659, N523);
and AND4 (N737, N736, N383, N233, N481);
not NOT1 (N738, N732);
buf BUF1 (N739, N729);
nor NOR4 (N740, N720, N558, N549, N173);
nand NAND3 (N741, N727, N182, N398);
not NOT1 (N742, N731);
nor NOR3 (N743, N742, N533, N269);
buf BUF1 (N744, N737);
buf BUF1 (N745, N744);
not NOT1 (N746, N730);
and AND2 (N747, N739, N573);
xor XOR2 (N748, N740, N508);
buf BUF1 (N749, N738);
nor NOR4 (N750, N741, N581, N413, N219);
nor NOR3 (N751, N750, N411, N422);
not NOT1 (N752, N746);
and AND2 (N753, N735, N484);
or OR4 (N754, N745, N172, N210, N276);
nand NAND4 (N755, N717, N598, N493, N689);
not NOT1 (N756, N753);
or OR3 (N757, N743, N443, N11);
nand NAND3 (N758, N749, N107, N38);
buf BUF1 (N759, N748);
not NOT1 (N760, N754);
and AND4 (N761, N760, N461, N419, N647);
nand NAND2 (N762, N758, N155);
nand NAND3 (N763, N762, N399, N557);
and AND4 (N764, N757, N176, N567, N318);
nand NAND4 (N765, N763, N42, N485, N358);
not NOT1 (N766, N764);
and AND3 (N767, N726, N720, N166);
not NOT1 (N768, N755);
xor XOR2 (N769, N756, N710);
or OR4 (N770, N765, N537, N27, N179);
buf BUF1 (N771, N770);
or OR2 (N772, N752, N45);
or OR3 (N773, N769, N192, N347);
xor XOR2 (N774, N768, N441);
xor XOR2 (N775, N751, N61);
and AND2 (N776, N759, N569);
or OR4 (N777, N761, N380, N210, N598);
and AND2 (N778, N747, N545);
buf BUF1 (N779, N766);
xor XOR2 (N780, N777, N383);
and AND3 (N781, N772, N687, N264);
buf BUF1 (N782, N776);
xor XOR2 (N783, N774, N440);
or OR2 (N784, N767, N71);
and AND4 (N785, N783, N166, N275, N690);
and AND4 (N786, N782, N752, N394, N612);
and AND3 (N787, N780, N731, N459);
and AND3 (N788, N771, N298, N475);
nor NOR3 (N789, N784, N607, N713);
or OR3 (N790, N779, N84, N738);
buf BUF1 (N791, N775);
and AND2 (N792, N785, N465);
buf BUF1 (N793, N790);
nor NOR2 (N794, N789, N383);
nand NAND4 (N795, N786, N399, N451, N567);
nand NAND4 (N796, N792, N261, N245, N38);
nand NAND2 (N797, N787, N765);
xor XOR2 (N798, N796, N202);
or OR3 (N799, N797, N543, N625);
xor XOR2 (N800, N791, N251);
nand NAND3 (N801, N788, N789, N187);
xor XOR2 (N802, N801, N431);
and AND3 (N803, N781, N560, N702);
or OR2 (N804, N795, N448);
not NOT1 (N805, N804);
or OR4 (N806, N794, N756, N342, N219);
nor NOR4 (N807, N805, N57, N379, N357);
buf BUF1 (N808, N778);
not NOT1 (N809, N793);
nand NAND2 (N810, N799, N256);
nand NAND2 (N811, N808, N584);
or OR4 (N812, N810, N499, N572, N333);
nor NOR3 (N813, N811, N449, N740);
not NOT1 (N814, N800);
xor XOR2 (N815, N809, N97);
xor XOR2 (N816, N814, N805);
nor NOR3 (N817, N798, N800, N518);
buf BUF1 (N818, N817);
buf BUF1 (N819, N816);
buf BUF1 (N820, N803);
or OR2 (N821, N815, N814);
buf BUF1 (N822, N773);
buf BUF1 (N823, N818);
nand NAND2 (N824, N813, N401);
xor XOR2 (N825, N820, N384);
nor NOR3 (N826, N812, N302, N225);
and AND2 (N827, N806, N307);
or OR2 (N828, N826, N585);
nor NOR3 (N829, N822, N676, N237);
not NOT1 (N830, N821);
nor NOR2 (N831, N828, N101);
buf BUF1 (N832, N827);
buf BUF1 (N833, N830);
nand NAND3 (N834, N832, N140, N374);
nand NAND4 (N835, N807, N807, N663, N727);
xor XOR2 (N836, N834, N355);
buf BUF1 (N837, N831);
buf BUF1 (N838, N829);
nand NAND3 (N839, N836, N690, N124);
nor NOR2 (N840, N838, N398);
buf BUF1 (N841, N837);
nand NAND4 (N842, N823, N124, N247, N292);
nand NAND2 (N843, N833, N728);
not NOT1 (N844, N824);
not NOT1 (N845, N839);
nor NOR4 (N846, N841, N90, N603, N235);
buf BUF1 (N847, N802);
xor XOR2 (N848, N844, N770);
xor XOR2 (N849, N845, N595);
or OR3 (N850, N847, N16, N296);
not NOT1 (N851, N843);
or OR2 (N852, N840, N767);
nor NOR4 (N853, N852, N706, N75, N382);
nand NAND3 (N854, N849, N735, N147);
xor XOR2 (N855, N825, N697);
not NOT1 (N856, N848);
and AND3 (N857, N846, N164, N239);
and AND4 (N858, N842, N411, N781, N674);
not NOT1 (N859, N856);
buf BUF1 (N860, N850);
buf BUF1 (N861, N859);
or OR2 (N862, N858, N153);
xor XOR2 (N863, N861, N130);
and AND2 (N864, N854, N78);
or OR3 (N865, N835, N359, N713);
xor XOR2 (N866, N863, N402);
or OR4 (N867, N853, N269, N689, N323);
and AND2 (N868, N866, N334);
nand NAND3 (N869, N865, N356, N129);
xor XOR2 (N870, N864, N273);
and AND4 (N871, N857, N732, N98, N49);
nand NAND4 (N872, N871, N52, N815, N813);
nand NAND3 (N873, N869, N279, N713);
nor NOR2 (N874, N872, N781);
and AND2 (N875, N870, N612);
buf BUF1 (N876, N819);
xor XOR2 (N877, N875, N513);
buf BUF1 (N878, N877);
nand NAND4 (N879, N855, N732, N461, N75);
nand NAND2 (N880, N868, N716);
buf BUF1 (N881, N851);
buf BUF1 (N882, N867);
nor NOR3 (N883, N878, N748, N854);
nor NOR2 (N884, N881, N752);
xor XOR2 (N885, N874, N102);
xor XOR2 (N886, N880, N222);
not NOT1 (N887, N886);
nor NOR2 (N888, N879, N264);
not NOT1 (N889, N876);
xor XOR2 (N890, N883, N555);
nor NOR2 (N891, N887, N689);
nand NAND4 (N892, N884, N607, N864, N140);
or OR4 (N893, N892, N516, N290, N665);
nor NOR3 (N894, N873, N870, N285);
and AND3 (N895, N862, N538, N347);
nor NOR3 (N896, N893, N681, N786);
xor XOR2 (N897, N889, N320);
nor NOR4 (N898, N896, N638, N320, N569);
buf BUF1 (N899, N860);
nor NOR4 (N900, N890, N897, N195, N135);
and AND4 (N901, N120, N130, N480, N776);
xor XOR2 (N902, N882, N654);
or OR2 (N903, N885, N529);
nand NAND3 (N904, N901, N745, N447);
buf BUF1 (N905, N904);
or OR4 (N906, N895, N17, N449, N57);
nand NAND4 (N907, N900, N352, N287, N591);
buf BUF1 (N908, N906);
nand NAND3 (N909, N888, N621, N120);
and AND2 (N910, N907, N571);
buf BUF1 (N911, N891);
or OR2 (N912, N894, N414);
xor XOR2 (N913, N911, N676);
xor XOR2 (N914, N905, N210);
nand NAND4 (N915, N910, N446, N298, N810);
xor XOR2 (N916, N899, N212);
or OR2 (N917, N914, N410);
buf BUF1 (N918, N903);
xor XOR2 (N919, N908, N66);
nand NAND2 (N920, N912, N172);
or OR3 (N921, N913, N340, N765);
xor XOR2 (N922, N920, N476);
nor NOR4 (N923, N922, N734, N516, N599);
xor XOR2 (N924, N921, N647);
xor XOR2 (N925, N915, N240);
not NOT1 (N926, N923);
or OR4 (N927, N902, N841, N322, N866);
buf BUF1 (N928, N924);
and AND3 (N929, N909, N512, N534);
nand NAND4 (N930, N919, N237, N479, N893);
or OR4 (N931, N926, N599, N636, N638);
or OR2 (N932, N917, N883);
xor XOR2 (N933, N918, N585);
nor NOR4 (N934, N933, N815, N367, N417);
buf BUF1 (N935, N930);
xor XOR2 (N936, N898, N49);
or OR2 (N937, N934, N724);
or OR4 (N938, N935, N305, N90, N132);
nor NOR2 (N939, N932, N265);
buf BUF1 (N940, N931);
xor XOR2 (N941, N936, N103);
xor XOR2 (N942, N927, N86);
nor NOR3 (N943, N942, N937, N581);
not NOT1 (N944, N154);
buf BUF1 (N945, N941);
not NOT1 (N946, N925);
nand NAND4 (N947, N943, N895, N182, N209);
nand NAND4 (N948, N946, N720, N364, N378);
nor NOR2 (N949, N928, N383);
and AND4 (N950, N947, N703, N687, N119);
nand NAND2 (N951, N950, N394);
xor XOR2 (N952, N944, N99);
nor NOR4 (N953, N948, N708, N914, N566);
and AND3 (N954, N953, N642, N400);
nor NOR3 (N955, N916, N395, N640);
nor NOR4 (N956, N938, N901, N856, N249);
buf BUF1 (N957, N955);
nand NAND2 (N958, N940, N289);
xor XOR2 (N959, N939, N803);
nand NAND4 (N960, N952, N170, N902, N337);
and AND2 (N961, N956, N655);
nand NAND2 (N962, N951, N901);
or OR2 (N963, N945, N365);
xor XOR2 (N964, N963, N820);
nor NOR4 (N965, N962, N769, N532, N199);
or OR2 (N966, N959, N386);
xor XOR2 (N967, N957, N534);
nor NOR2 (N968, N949, N94);
xor XOR2 (N969, N965, N108);
xor XOR2 (N970, N954, N73);
xor XOR2 (N971, N969, N33);
not NOT1 (N972, N964);
not NOT1 (N973, N961);
xor XOR2 (N974, N929, N691);
nor NOR3 (N975, N971, N556, N940);
nand NAND3 (N976, N970, N144, N86);
not NOT1 (N977, N960);
nand NAND3 (N978, N976, N761, N708);
not NOT1 (N979, N966);
xor XOR2 (N980, N974, N796);
or OR4 (N981, N972, N789, N537, N159);
and AND2 (N982, N968, N54);
nand NAND2 (N983, N977, N470);
xor XOR2 (N984, N979, N719);
or OR3 (N985, N983, N789, N508);
nand NAND4 (N986, N975, N579, N960, N690);
buf BUF1 (N987, N986);
and AND2 (N988, N978, N975);
or OR2 (N989, N984, N837);
not NOT1 (N990, N981);
not NOT1 (N991, N988);
buf BUF1 (N992, N989);
nor NOR2 (N993, N980, N487);
or OR4 (N994, N973, N182, N914, N375);
nand NAND4 (N995, N958, N192, N777, N409);
nor NOR4 (N996, N994, N82, N314, N760);
xor XOR2 (N997, N993, N606);
not NOT1 (N998, N992);
xor XOR2 (N999, N990, N207);
nor NOR2 (N1000, N998, N266);
and AND3 (N1001, N967, N987, N219);
and AND2 (N1002, N58, N207);
or OR2 (N1003, N985, N20);
xor XOR2 (N1004, N1002, N728);
not NOT1 (N1005, N1003);
nand NAND3 (N1006, N1004, N531, N431);
or OR4 (N1007, N995, N160, N537, N818);
nor NOR2 (N1008, N991, N81);
and AND3 (N1009, N1008, N752, N240);
buf BUF1 (N1010, N1005);
not NOT1 (N1011, N997);
buf BUF1 (N1012, N1009);
and AND4 (N1013, N996, N885, N96, N111);
buf BUF1 (N1014, N1013);
not NOT1 (N1015, N1007);
nand NAND4 (N1016, N1000, N208, N998, N587);
or OR2 (N1017, N999, N190);
and AND4 (N1018, N1006, N21, N207, N87);
not NOT1 (N1019, N1018);
and AND4 (N1020, N1015, N38, N599, N408);
xor XOR2 (N1021, N1020, N197);
nand NAND4 (N1022, N1010, N425, N340, N255);
and AND2 (N1023, N1016, N298);
not NOT1 (N1024, N1019);
buf BUF1 (N1025, N1024);
nand NAND4 (N1026, N1022, N662, N666, N986);
buf BUF1 (N1027, N1012);
or OR4 (N1028, N1017, N132, N313, N106);
and AND3 (N1029, N1021, N186, N136);
or OR2 (N1030, N1028, N641);
xor XOR2 (N1031, N1027, N433);
and AND3 (N1032, N1014, N465, N214);
nand NAND2 (N1033, N1032, N811);
nor NOR4 (N1034, N1001, N722, N802, N117);
not NOT1 (N1035, N1026);
nand NAND2 (N1036, N1035, N543);
or OR2 (N1037, N1029, N920);
xor XOR2 (N1038, N1025, N851);
nand NAND2 (N1039, N1038, N349);
buf BUF1 (N1040, N1033);
xor XOR2 (N1041, N1031, N889);
not NOT1 (N1042, N1041);
xor XOR2 (N1043, N1040, N942);
xor XOR2 (N1044, N982, N970);
buf BUF1 (N1045, N1011);
nand NAND4 (N1046, N1042, N135, N913, N68);
buf BUF1 (N1047, N1036);
xor XOR2 (N1048, N1030, N1009);
and AND2 (N1049, N1045, N569);
buf BUF1 (N1050, N1043);
or OR4 (N1051, N1023, N168, N219, N150);
buf BUF1 (N1052, N1048);
nor NOR4 (N1053, N1050, N485, N171, N638);
or OR4 (N1054, N1046, N953, N26, N1028);
nand NAND2 (N1055, N1049, N663);
and AND2 (N1056, N1051, N634);
not NOT1 (N1057, N1034);
nor NOR2 (N1058, N1039, N906);
not NOT1 (N1059, N1037);
or OR2 (N1060, N1055, N307);
nor NOR2 (N1061, N1059, N707);
xor XOR2 (N1062, N1056, N1042);
nand NAND2 (N1063, N1047, N973);
not NOT1 (N1064, N1052);
buf BUF1 (N1065, N1060);
xor XOR2 (N1066, N1044, N972);
and AND3 (N1067, N1058, N655, N900);
or OR2 (N1068, N1065, N865);
buf BUF1 (N1069, N1062);
nand NAND4 (N1070, N1063, N1044, N209, N239);
and AND4 (N1071, N1070, N30, N52, N30);
xor XOR2 (N1072, N1054, N535);
nand NAND4 (N1073, N1069, N664, N906, N525);
and AND2 (N1074, N1071, N202);
xor XOR2 (N1075, N1053, N510);
or OR2 (N1076, N1064, N202);
buf BUF1 (N1077, N1074);
not NOT1 (N1078, N1072);
buf BUF1 (N1079, N1068);
not NOT1 (N1080, N1075);
buf BUF1 (N1081, N1076);
and AND3 (N1082, N1079, N473, N1077);
not NOT1 (N1083, N565);
buf BUF1 (N1084, N1073);
xor XOR2 (N1085, N1061, N885);
or OR2 (N1086, N1083, N57);
xor XOR2 (N1087, N1067, N934);
nor NOR4 (N1088, N1057, N412, N1048, N435);
xor XOR2 (N1089, N1088, N474);
nor NOR2 (N1090, N1084, N515);
buf BUF1 (N1091, N1078);
not NOT1 (N1092, N1089);
xor XOR2 (N1093, N1092, N475);
not NOT1 (N1094, N1091);
not NOT1 (N1095, N1087);
nor NOR3 (N1096, N1086, N608, N649);
and AND3 (N1097, N1081, N781, N626);
nand NAND2 (N1098, N1093, N222);
nand NAND3 (N1099, N1080, N591, N206);
buf BUF1 (N1100, N1098);
and AND4 (N1101, N1097, N472, N744, N269);
xor XOR2 (N1102, N1096, N630);
and AND3 (N1103, N1085, N473, N362);
nand NAND4 (N1104, N1066, N1004, N687, N1060);
xor XOR2 (N1105, N1100, N923);
nor NOR2 (N1106, N1105, N782);
buf BUF1 (N1107, N1102);
or OR3 (N1108, N1104, N756, N260);
nor NOR2 (N1109, N1103, N783);
xor XOR2 (N1110, N1090, N602);
nand NAND2 (N1111, N1082, N620);
and AND3 (N1112, N1108, N390, N773);
nand NAND4 (N1113, N1110, N327, N579, N661);
xor XOR2 (N1114, N1094, N977);
and AND2 (N1115, N1112, N361);
not NOT1 (N1116, N1107);
and AND4 (N1117, N1114, N821, N1061, N314);
nand NAND3 (N1118, N1113, N494, N53);
nor NOR4 (N1119, N1117, N1033, N506, N176);
nand NAND4 (N1120, N1119, N40, N351, N628);
buf BUF1 (N1121, N1111);
not NOT1 (N1122, N1115);
not NOT1 (N1123, N1121);
or OR3 (N1124, N1101, N588, N649);
nor NOR3 (N1125, N1120, N48, N101);
and AND3 (N1126, N1116, N944, N634);
buf BUF1 (N1127, N1123);
xor XOR2 (N1128, N1106, N399);
nand NAND3 (N1129, N1124, N607, N885);
nand NAND4 (N1130, N1122, N255, N630, N693);
xor XOR2 (N1131, N1130, N1123);
buf BUF1 (N1132, N1128);
xor XOR2 (N1133, N1099, N335);
and AND3 (N1134, N1109, N564, N73);
nor NOR4 (N1135, N1129, N424, N771, N878);
not NOT1 (N1136, N1125);
nand NAND4 (N1137, N1134, N271, N439, N206);
not NOT1 (N1138, N1131);
not NOT1 (N1139, N1136);
nand NAND4 (N1140, N1127, N522, N760, N1008);
nor NOR3 (N1141, N1139, N433, N323);
nand NAND4 (N1142, N1141, N560, N825, N984);
xor XOR2 (N1143, N1118, N549);
nand NAND3 (N1144, N1138, N99, N982);
nand NAND3 (N1145, N1133, N1006, N208);
buf BUF1 (N1146, N1140);
nor NOR2 (N1147, N1137, N87);
not NOT1 (N1148, N1126);
or OR4 (N1149, N1145, N875, N931, N528);
buf BUF1 (N1150, N1148);
or OR2 (N1151, N1095, N5);
nor NOR4 (N1152, N1135, N882, N327, N214);
or OR2 (N1153, N1149, N1061);
nand NAND3 (N1154, N1150, N1144, N782);
or OR2 (N1155, N638, N816);
or OR3 (N1156, N1146, N930, N755);
nor NOR4 (N1157, N1151, N298, N599, N1111);
nor NOR2 (N1158, N1152, N59);
buf BUF1 (N1159, N1143);
not NOT1 (N1160, N1153);
not NOT1 (N1161, N1147);
buf BUF1 (N1162, N1157);
nor NOR3 (N1163, N1158, N805, N693);
xor XOR2 (N1164, N1161, N691);
nor NOR3 (N1165, N1159, N928, N136);
nand NAND2 (N1166, N1156, N688);
xor XOR2 (N1167, N1166, N61);
or OR3 (N1168, N1132, N127, N1123);
xor XOR2 (N1169, N1167, N604);
not NOT1 (N1170, N1163);
nor NOR2 (N1171, N1165, N697);
xor XOR2 (N1172, N1155, N339);
nor NOR2 (N1173, N1170, N782);
not NOT1 (N1174, N1154);
nor NOR3 (N1175, N1142, N794, N583);
buf BUF1 (N1176, N1175);
or OR3 (N1177, N1173, N214, N193);
not NOT1 (N1178, N1172);
buf BUF1 (N1179, N1171);
and AND4 (N1180, N1179, N871, N67, N179);
nand NAND4 (N1181, N1178, N151, N983, N41);
xor XOR2 (N1182, N1176, N403);
and AND3 (N1183, N1160, N1038, N698);
nor NOR3 (N1184, N1183, N1076, N423);
xor XOR2 (N1185, N1169, N604);
nor NOR3 (N1186, N1164, N342, N1078);
nor NOR2 (N1187, N1180, N841);
and AND4 (N1188, N1181, N932, N962, N820);
nand NAND3 (N1189, N1186, N1082, N641);
or OR3 (N1190, N1177, N660, N1123);
and AND2 (N1191, N1174, N639);
not NOT1 (N1192, N1185);
not NOT1 (N1193, N1191);
nor NOR2 (N1194, N1182, N537);
xor XOR2 (N1195, N1189, N770);
nor NOR3 (N1196, N1193, N403, N986);
not NOT1 (N1197, N1195);
xor XOR2 (N1198, N1196, N933);
not NOT1 (N1199, N1198);
buf BUF1 (N1200, N1188);
nor NOR3 (N1201, N1197, N372, N913);
and AND4 (N1202, N1162, N745, N579, N569);
xor XOR2 (N1203, N1199, N1070);
or OR4 (N1204, N1192, N512, N1139, N820);
or OR2 (N1205, N1203, N2);
xor XOR2 (N1206, N1168, N827);
xor XOR2 (N1207, N1204, N1027);
buf BUF1 (N1208, N1184);
or OR3 (N1209, N1202, N1170, N1005);
not NOT1 (N1210, N1209);
xor XOR2 (N1211, N1207, N885);
not NOT1 (N1212, N1200);
nor NOR4 (N1213, N1187, N804, N975, N71);
buf BUF1 (N1214, N1212);
nand NAND3 (N1215, N1190, N197, N1190);
and AND2 (N1216, N1194, N509);
nor NOR3 (N1217, N1216, N46, N874);
xor XOR2 (N1218, N1215, N264);
buf BUF1 (N1219, N1214);
or OR3 (N1220, N1219, N305, N989);
xor XOR2 (N1221, N1211, N304);
nor NOR4 (N1222, N1208, N635, N511, N447);
buf BUF1 (N1223, N1206);
or OR4 (N1224, N1205, N936, N559, N484);
nor NOR3 (N1225, N1224, N932, N4);
nand NAND3 (N1226, N1217, N624, N859);
nand NAND2 (N1227, N1226, N128);
and AND3 (N1228, N1223, N727, N255);
xor XOR2 (N1229, N1225, N634);
and AND3 (N1230, N1201, N1131, N721);
not NOT1 (N1231, N1229);
not NOT1 (N1232, N1231);
nand NAND3 (N1233, N1213, N1075, N721);
buf BUF1 (N1234, N1227);
not NOT1 (N1235, N1220);
buf BUF1 (N1236, N1230);
xor XOR2 (N1237, N1210, N957);
nand NAND3 (N1238, N1232, N1007, N334);
nor NOR3 (N1239, N1228, N181, N652);
xor XOR2 (N1240, N1235, N359);
or OR3 (N1241, N1239, N910, N1149);
nand NAND3 (N1242, N1221, N670, N1172);
and AND3 (N1243, N1241, N921, N147);
or OR4 (N1244, N1238, N786, N124, N303);
and AND2 (N1245, N1243, N195);
or OR3 (N1246, N1240, N1103, N723);
nand NAND2 (N1247, N1234, N328);
buf BUF1 (N1248, N1246);
and AND4 (N1249, N1237, N8, N1019, N983);
nand NAND3 (N1250, N1233, N10, N801);
nand NAND4 (N1251, N1250, N905, N878, N539);
nand NAND4 (N1252, N1236, N970, N434, N888);
nand NAND3 (N1253, N1222, N482, N638);
and AND4 (N1254, N1242, N588, N842, N570);
not NOT1 (N1255, N1252);
xor XOR2 (N1256, N1253, N1106);
and AND2 (N1257, N1218, N1073);
or OR4 (N1258, N1249, N654, N1045, N1014);
nor NOR3 (N1259, N1248, N711, N1013);
xor XOR2 (N1260, N1258, N1179);
nor NOR2 (N1261, N1245, N1177);
nand NAND4 (N1262, N1256, N372, N199, N889);
xor XOR2 (N1263, N1251, N786);
nand NAND4 (N1264, N1255, N233, N804, N1105);
and AND2 (N1265, N1262, N813);
buf BUF1 (N1266, N1259);
xor XOR2 (N1267, N1263, N474);
not NOT1 (N1268, N1267);
nor NOR4 (N1269, N1247, N727, N178, N673);
xor XOR2 (N1270, N1266, N701);
buf BUF1 (N1271, N1264);
and AND2 (N1272, N1257, N682);
xor XOR2 (N1273, N1244, N780);
nor NOR3 (N1274, N1268, N74, N546);
nand NAND4 (N1275, N1270, N656, N527, N1187);
buf BUF1 (N1276, N1274);
and AND4 (N1277, N1261, N800, N1174, N1017);
buf BUF1 (N1278, N1273);
nand NAND2 (N1279, N1275, N763);
not NOT1 (N1280, N1278);
and AND2 (N1281, N1276, N1018);
buf BUF1 (N1282, N1271);
nand NAND4 (N1283, N1254, N1236, N607, N37);
nand NAND3 (N1284, N1281, N974, N639);
and AND2 (N1285, N1260, N838);
and AND4 (N1286, N1282, N845, N463, N1162);
nand NAND2 (N1287, N1284, N1153);
buf BUF1 (N1288, N1279);
buf BUF1 (N1289, N1285);
and AND4 (N1290, N1289, N338, N777, N1095);
not NOT1 (N1291, N1287);
buf BUF1 (N1292, N1291);
xor XOR2 (N1293, N1280, N394);
nand NAND2 (N1294, N1265, N479);
nor NOR4 (N1295, N1288, N502, N598, N667);
or OR3 (N1296, N1293, N843, N173);
nor NOR3 (N1297, N1290, N455, N695);
and AND3 (N1298, N1277, N224, N1003);
nand NAND2 (N1299, N1286, N430);
buf BUF1 (N1300, N1269);
nor NOR3 (N1301, N1294, N209, N140);
xor XOR2 (N1302, N1301, N346);
not NOT1 (N1303, N1300);
and AND2 (N1304, N1302, N474);
and AND2 (N1305, N1292, N656);
nand NAND4 (N1306, N1304, N617, N1083, N518);
nor NOR3 (N1307, N1299, N279, N440);
nor NOR4 (N1308, N1303, N131, N417, N1224);
buf BUF1 (N1309, N1296);
or OR2 (N1310, N1309, N674);
and AND4 (N1311, N1305, N687, N1213, N394);
nor NOR2 (N1312, N1297, N561);
and AND4 (N1313, N1306, N624, N948, N895);
not NOT1 (N1314, N1283);
nand NAND3 (N1315, N1311, N153, N707);
and AND3 (N1316, N1313, N530, N487);
and AND2 (N1317, N1315, N551);
nor NOR4 (N1318, N1308, N1275, N1103, N1247);
nor NOR2 (N1319, N1318, N916);
nand NAND4 (N1320, N1314, N1268, N407, N1248);
nor NOR3 (N1321, N1307, N260, N544);
or OR3 (N1322, N1272, N1309, N3);
buf BUF1 (N1323, N1317);
buf BUF1 (N1324, N1322);
nand NAND3 (N1325, N1295, N653, N927);
or OR4 (N1326, N1310, N650, N612, N692);
or OR4 (N1327, N1325, N298, N795, N1122);
nand NAND3 (N1328, N1324, N879, N509);
nor NOR3 (N1329, N1320, N105, N1100);
nand NAND2 (N1330, N1316, N583);
or OR4 (N1331, N1323, N563, N605, N1134);
and AND2 (N1332, N1298, N50);
and AND2 (N1333, N1328, N1278);
nor NOR4 (N1334, N1321, N153, N10, N962);
not NOT1 (N1335, N1332);
nand NAND4 (N1336, N1312, N292, N970, N1059);
not NOT1 (N1337, N1335);
and AND3 (N1338, N1326, N153, N1281);
buf BUF1 (N1339, N1334);
xor XOR2 (N1340, N1337, N377);
nand NAND3 (N1341, N1327, N1311, N487);
buf BUF1 (N1342, N1329);
nand NAND2 (N1343, N1342, N1064);
nor NOR2 (N1344, N1333, N1187);
xor XOR2 (N1345, N1340, N1038);
xor XOR2 (N1346, N1341, N191);
and AND3 (N1347, N1338, N140, N1340);
and AND2 (N1348, N1331, N1107);
or OR2 (N1349, N1348, N556);
nand NAND2 (N1350, N1344, N1031);
xor XOR2 (N1351, N1349, N1166);
nor NOR4 (N1352, N1319, N406, N529, N319);
nor NOR2 (N1353, N1336, N733);
nand NAND4 (N1354, N1346, N1165, N562, N771);
not NOT1 (N1355, N1330);
xor XOR2 (N1356, N1351, N793);
nor NOR2 (N1357, N1352, N157);
nand NAND3 (N1358, N1357, N1297, N342);
and AND2 (N1359, N1354, N593);
not NOT1 (N1360, N1353);
buf BUF1 (N1361, N1359);
nor NOR2 (N1362, N1358, N1298);
not NOT1 (N1363, N1360);
not NOT1 (N1364, N1355);
nor NOR4 (N1365, N1364, N457, N299, N1127);
and AND3 (N1366, N1350, N409, N1354);
and AND3 (N1367, N1339, N762, N1256);
nand NAND3 (N1368, N1343, N992, N784);
nor NOR2 (N1369, N1356, N38);
xor XOR2 (N1370, N1345, N130);
nor NOR4 (N1371, N1347, N373, N422, N379);
not NOT1 (N1372, N1367);
xor XOR2 (N1373, N1371, N1123);
and AND4 (N1374, N1365, N935, N1186, N18);
buf BUF1 (N1375, N1368);
nor NOR4 (N1376, N1375, N571, N652, N1127);
nor NOR4 (N1377, N1369, N602, N1337, N795);
buf BUF1 (N1378, N1372);
nand NAND3 (N1379, N1363, N80, N139);
xor XOR2 (N1380, N1373, N678);
or OR3 (N1381, N1370, N800, N242);
and AND3 (N1382, N1362, N427, N687);
buf BUF1 (N1383, N1366);
xor XOR2 (N1384, N1383, N820);
and AND2 (N1385, N1377, N205);
and AND4 (N1386, N1379, N616, N1184, N756);
not NOT1 (N1387, N1384);
not NOT1 (N1388, N1361);
not NOT1 (N1389, N1385);
not NOT1 (N1390, N1374);
or OR2 (N1391, N1376, N1374);
nor NOR2 (N1392, N1386, N880);
nor NOR2 (N1393, N1382, N380);
not NOT1 (N1394, N1389);
nor NOR2 (N1395, N1388, N1249);
nor NOR3 (N1396, N1391, N598, N1288);
buf BUF1 (N1397, N1393);
and AND4 (N1398, N1380, N715, N1324, N57);
not NOT1 (N1399, N1397);
not NOT1 (N1400, N1399);
or OR2 (N1401, N1400, N150);
not NOT1 (N1402, N1396);
or OR3 (N1403, N1390, N98, N1033);
nand NAND2 (N1404, N1381, N11);
nor NOR4 (N1405, N1392, N570, N564, N602);
nand NAND2 (N1406, N1395, N414);
nor NOR2 (N1407, N1403, N779);
or OR4 (N1408, N1401, N138, N15, N163);
buf BUF1 (N1409, N1378);
xor XOR2 (N1410, N1398, N68);
buf BUF1 (N1411, N1409);
xor XOR2 (N1412, N1387, N342);
buf BUF1 (N1413, N1412);
not NOT1 (N1414, N1402);
or OR2 (N1415, N1410, N1245);
or OR3 (N1416, N1394, N376, N1392);
nor NOR3 (N1417, N1416, N1212, N264);
nor NOR2 (N1418, N1405, N441);
not NOT1 (N1419, N1406);
buf BUF1 (N1420, N1411);
nor NOR2 (N1421, N1420, N1034);
or OR3 (N1422, N1414, N476, N1076);
or OR2 (N1423, N1422, N34);
buf BUF1 (N1424, N1421);
nor NOR4 (N1425, N1417, N128, N54, N1243);
nand NAND2 (N1426, N1418, N412);
buf BUF1 (N1427, N1404);
nor NOR4 (N1428, N1415, N453, N693, N248);
and AND2 (N1429, N1419, N549);
nor NOR3 (N1430, N1413, N1344, N932);
or OR2 (N1431, N1425, N839);
or OR3 (N1432, N1428, N1038, N35);
and AND4 (N1433, N1427, N1139, N1305, N1150);
and AND4 (N1434, N1432, N259, N560, N895);
and AND2 (N1435, N1431, N1331);
not NOT1 (N1436, N1408);
xor XOR2 (N1437, N1426, N956);
and AND3 (N1438, N1433, N1307, N138);
buf BUF1 (N1439, N1438);
nand NAND4 (N1440, N1429, N216, N905, N988);
and AND3 (N1441, N1434, N1272, N117);
xor XOR2 (N1442, N1437, N500);
nor NOR4 (N1443, N1407, N856, N1182, N739);
xor XOR2 (N1444, N1442, N1014);
buf BUF1 (N1445, N1444);
or OR3 (N1446, N1441, N61, N489);
or OR2 (N1447, N1436, N1364);
nand NAND2 (N1448, N1443, N1406);
nand NAND3 (N1449, N1445, N335, N617);
buf BUF1 (N1450, N1430);
nor NOR3 (N1451, N1424, N771, N282);
not NOT1 (N1452, N1450);
not NOT1 (N1453, N1446);
and AND3 (N1454, N1449, N946, N235);
xor XOR2 (N1455, N1440, N913);
or OR4 (N1456, N1451, N616, N1399, N659);
nand NAND2 (N1457, N1454, N639);
or OR2 (N1458, N1456, N1042);
nand NAND2 (N1459, N1455, N675);
or OR2 (N1460, N1448, N1378);
buf BUF1 (N1461, N1460);
not NOT1 (N1462, N1447);
buf BUF1 (N1463, N1462);
nor NOR3 (N1464, N1457, N440, N229);
or OR2 (N1465, N1453, N176);
and AND2 (N1466, N1465, N679);
nor NOR2 (N1467, N1463, N842);
buf BUF1 (N1468, N1466);
and AND2 (N1469, N1452, N1158);
and AND3 (N1470, N1459, N171, N1425);
and AND3 (N1471, N1423, N646, N1132);
nor NOR2 (N1472, N1470, N781);
or OR2 (N1473, N1439, N223);
nor NOR2 (N1474, N1458, N620);
or OR3 (N1475, N1473, N1004, N120);
xor XOR2 (N1476, N1464, N1085);
buf BUF1 (N1477, N1469);
or OR4 (N1478, N1461, N504, N1203, N1024);
nor NOR3 (N1479, N1475, N105, N517);
xor XOR2 (N1480, N1477, N187);
buf BUF1 (N1481, N1435);
xor XOR2 (N1482, N1472, N1124);
and AND2 (N1483, N1482, N253);
xor XOR2 (N1484, N1467, N877);
buf BUF1 (N1485, N1483);
nor NOR4 (N1486, N1476, N996, N2, N1356);
not NOT1 (N1487, N1486);
xor XOR2 (N1488, N1471, N370);
nand NAND3 (N1489, N1468, N844, N1107);
buf BUF1 (N1490, N1481);
or OR3 (N1491, N1488, N1155, N398);
or OR2 (N1492, N1489, N1234);
nand NAND4 (N1493, N1491, N74, N164, N291);
nand NAND3 (N1494, N1485, N69, N84);
not NOT1 (N1495, N1474);
xor XOR2 (N1496, N1478, N582);
buf BUF1 (N1497, N1484);
nand NAND2 (N1498, N1487, N642);
and AND2 (N1499, N1490, N629);
not NOT1 (N1500, N1499);
or OR3 (N1501, N1493, N558, N117);
nand NAND2 (N1502, N1480, N108);
and AND4 (N1503, N1497, N157, N1488, N1006);
not NOT1 (N1504, N1498);
or OR2 (N1505, N1502, N1203);
not NOT1 (N1506, N1501);
nand NAND2 (N1507, N1495, N769);
nor NOR3 (N1508, N1503, N1249, N1202);
xor XOR2 (N1509, N1494, N1353);
or OR2 (N1510, N1496, N915);
and AND3 (N1511, N1506, N510, N568);
buf BUF1 (N1512, N1507);
and AND2 (N1513, N1512, N934);
or OR4 (N1514, N1511, N322, N209, N80);
and AND2 (N1515, N1500, N103);
nand NAND2 (N1516, N1492, N200);
and AND3 (N1517, N1479, N637, N1075);
not NOT1 (N1518, N1514);
and AND3 (N1519, N1513, N611, N44);
nor NOR2 (N1520, N1510, N499);
not NOT1 (N1521, N1505);
buf BUF1 (N1522, N1517);
nor NOR4 (N1523, N1508, N794, N975, N930);
not NOT1 (N1524, N1509);
buf BUF1 (N1525, N1522);
nand NAND4 (N1526, N1523, N1283, N380, N1169);
buf BUF1 (N1527, N1518);
nor NOR3 (N1528, N1520, N863, N1046);
or OR2 (N1529, N1528, N465);
buf BUF1 (N1530, N1504);
nor NOR2 (N1531, N1529, N102);
xor XOR2 (N1532, N1524, N283);
or OR2 (N1533, N1515, N901);
not NOT1 (N1534, N1519);
buf BUF1 (N1535, N1516);
buf BUF1 (N1536, N1526);
buf BUF1 (N1537, N1521);
or OR4 (N1538, N1525, N32, N424, N905);
buf BUF1 (N1539, N1531);
or OR3 (N1540, N1535, N1227, N674);
xor XOR2 (N1541, N1532, N1046);
or OR4 (N1542, N1538, N583, N1461, N1168);
not NOT1 (N1543, N1542);
nand NAND4 (N1544, N1543, N958, N1261, N130);
not NOT1 (N1545, N1533);
and AND2 (N1546, N1534, N613);
xor XOR2 (N1547, N1541, N102);
and AND3 (N1548, N1536, N1232, N219);
nand NAND4 (N1549, N1548, N575, N662, N1024);
xor XOR2 (N1550, N1544, N157);
or OR4 (N1551, N1546, N705, N450, N1200);
not NOT1 (N1552, N1527);
and AND2 (N1553, N1549, N946);
buf BUF1 (N1554, N1545);
nor NOR2 (N1555, N1530, N523);
buf BUF1 (N1556, N1550);
and AND2 (N1557, N1540, N449);
buf BUF1 (N1558, N1552);
buf BUF1 (N1559, N1554);
xor XOR2 (N1560, N1558, N30);
not NOT1 (N1561, N1557);
not NOT1 (N1562, N1560);
buf BUF1 (N1563, N1555);
or OR3 (N1564, N1563, N245, N1050);
buf BUF1 (N1565, N1537);
and AND3 (N1566, N1553, N1494, N1268);
not NOT1 (N1567, N1561);
xor XOR2 (N1568, N1565, N1278);
nor NOR2 (N1569, N1559, N1235);
or OR3 (N1570, N1569, N44, N93);
not NOT1 (N1571, N1556);
not NOT1 (N1572, N1547);
buf BUF1 (N1573, N1562);
not NOT1 (N1574, N1551);
and AND3 (N1575, N1564, N333, N631);
nor NOR2 (N1576, N1574, N388);
nand NAND3 (N1577, N1571, N864, N93);
nand NAND2 (N1578, N1570, N1274);
nor NOR3 (N1579, N1567, N83, N779);
nand NAND4 (N1580, N1577, N363, N1263, N1546);
xor XOR2 (N1581, N1575, N283);
buf BUF1 (N1582, N1572);
nor NOR3 (N1583, N1539, N309, N1156);
and AND3 (N1584, N1573, N190, N356);
buf BUF1 (N1585, N1579);
not NOT1 (N1586, N1578);
and AND4 (N1587, N1582, N1363, N1176, N1491);
xor XOR2 (N1588, N1576, N1451);
nor NOR3 (N1589, N1583, N542, N965);
or OR4 (N1590, N1566, N254, N414, N1015);
and AND3 (N1591, N1586, N1544, N343);
nand NAND3 (N1592, N1585, N618, N464);
or OR3 (N1593, N1592, N1512, N1403);
and AND2 (N1594, N1591, N815);
not NOT1 (N1595, N1584);
buf BUF1 (N1596, N1593);
buf BUF1 (N1597, N1595);
nand NAND2 (N1598, N1588, N1431);
or OR3 (N1599, N1589, N1444, N387);
xor XOR2 (N1600, N1581, N90);
nand NAND3 (N1601, N1600, N1039, N1089);
buf BUF1 (N1602, N1594);
or OR3 (N1603, N1587, N960, N572);
buf BUF1 (N1604, N1602);
nand NAND4 (N1605, N1598, N1154, N1020, N24);
nand NAND2 (N1606, N1599, N1376);
xor XOR2 (N1607, N1597, N607);
buf BUF1 (N1608, N1590);
and AND2 (N1609, N1604, N70);
xor XOR2 (N1610, N1606, N765);
xor XOR2 (N1611, N1609, N587);
or OR2 (N1612, N1596, N1439);
or OR3 (N1613, N1611, N1317, N491);
nor NOR3 (N1614, N1608, N276, N1429);
buf BUF1 (N1615, N1603);
and AND2 (N1616, N1614, N1268);
nand NAND4 (N1617, N1613, N142, N1372, N700);
buf BUF1 (N1618, N1568);
and AND4 (N1619, N1605, N1162, N202, N629);
xor XOR2 (N1620, N1610, N560);
or OR3 (N1621, N1607, N557, N1601);
buf BUF1 (N1622, N85);
nand NAND4 (N1623, N1616, N1228, N51, N1321);
xor XOR2 (N1624, N1617, N330);
and AND3 (N1625, N1580, N549, N1127);
nand NAND2 (N1626, N1618, N1029);
xor XOR2 (N1627, N1620, N264);
or OR4 (N1628, N1615, N1136, N1530, N1617);
or OR2 (N1629, N1619, N1583);
or OR2 (N1630, N1628, N327);
and AND3 (N1631, N1622, N1630, N1166);
and AND2 (N1632, N1469, N179);
and AND2 (N1633, N1629, N1261);
not NOT1 (N1634, N1625);
buf BUF1 (N1635, N1633);
or OR3 (N1636, N1621, N1457, N261);
or OR3 (N1637, N1631, N839, N983);
nor NOR2 (N1638, N1634, N206);
xor XOR2 (N1639, N1624, N1360);
buf BUF1 (N1640, N1632);
nand NAND4 (N1641, N1636, N507, N732, N1062);
and AND4 (N1642, N1612, N16, N42, N1055);
or OR2 (N1643, N1639, N1271);
nor NOR4 (N1644, N1635, N963, N1212, N539);
buf BUF1 (N1645, N1638);
xor XOR2 (N1646, N1640, N509);
xor XOR2 (N1647, N1623, N1609);
or OR3 (N1648, N1642, N428, N996);
and AND4 (N1649, N1645, N409, N1095, N1512);
not NOT1 (N1650, N1626);
not NOT1 (N1651, N1643);
not NOT1 (N1652, N1627);
xor XOR2 (N1653, N1649, N1246);
not NOT1 (N1654, N1647);
and AND4 (N1655, N1654, N740, N1263, N170);
not NOT1 (N1656, N1644);
and AND2 (N1657, N1648, N457);
not NOT1 (N1658, N1655);
buf BUF1 (N1659, N1653);
and AND2 (N1660, N1641, N1024);
not NOT1 (N1661, N1660);
nand NAND4 (N1662, N1651, N246, N694, N1634);
nor NOR4 (N1663, N1659, N473, N1615, N1308);
nor NOR2 (N1664, N1650, N620);
nand NAND2 (N1665, N1664, N1231);
xor XOR2 (N1666, N1656, N170);
buf BUF1 (N1667, N1662);
nand NAND4 (N1668, N1646, N169, N887, N811);
buf BUF1 (N1669, N1666);
not NOT1 (N1670, N1665);
and AND3 (N1671, N1668, N1385, N373);
or OR4 (N1672, N1670, N1661, N1034, N392);
and AND4 (N1673, N116, N1295, N335, N554);
not NOT1 (N1674, N1658);
and AND3 (N1675, N1672, N1372, N890);
nor NOR2 (N1676, N1637, N146);
and AND2 (N1677, N1675, N1543);
and AND4 (N1678, N1657, N1479, N1482, N1434);
and AND3 (N1679, N1671, N1644, N1095);
buf BUF1 (N1680, N1667);
not NOT1 (N1681, N1676);
not NOT1 (N1682, N1669);
nand NAND4 (N1683, N1682, N188, N449, N877);
nand NAND2 (N1684, N1663, N934);
buf BUF1 (N1685, N1678);
buf BUF1 (N1686, N1673);
buf BUF1 (N1687, N1652);
nor NOR4 (N1688, N1679, N248, N282, N512);
not NOT1 (N1689, N1680);
nand NAND4 (N1690, N1685, N121, N607, N1305);
or OR3 (N1691, N1687, N664, N47);
not NOT1 (N1692, N1686);
buf BUF1 (N1693, N1677);
nand NAND3 (N1694, N1681, N697, N881);
not NOT1 (N1695, N1684);
not NOT1 (N1696, N1695);
xor XOR2 (N1697, N1674, N1009);
not NOT1 (N1698, N1689);
and AND4 (N1699, N1696, N119, N502, N1656);
buf BUF1 (N1700, N1698);
nor NOR4 (N1701, N1683, N1640, N18, N1033);
or OR3 (N1702, N1690, N852, N350);
not NOT1 (N1703, N1694);
buf BUF1 (N1704, N1702);
buf BUF1 (N1705, N1697);
buf BUF1 (N1706, N1701);
buf BUF1 (N1707, N1699);
or OR4 (N1708, N1706, N271, N910, N1500);
buf BUF1 (N1709, N1692);
nor NOR2 (N1710, N1707, N1149);
buf BUF1 (N1711, N1693);
nor NOR2 (N1712, N1691, N146);
or OR4 (N1713, N1710, N1566, N859, N311);
and AND4 (N1714, N1705, N87, N1344, N1624);
or OR4 (N1715, N1688, N1381, N820, N1376);
not NOT1 (N1716, N1703);
or OR2 (N1717, N1716, N176);
xor XOR2 (N1718, N1711, N1193);
and AND4 (N1719, N1714, N117, N1007, N725);
nand NAND4 (N1720, N1700, N1041, N624, N1286);
or OR4 (N1721, N1719, N440, N884, N369);
nor NOR4 (N1722, N1708, N632, N365, N1066);
nor NOR2 (N1723, N1722, N230);
nor NOR2 (N1724, N1717, N1606);
or OR2 (N1725, N1718, N884);
xor XOR2 (N1726, N1712, N66);
nand NAND4 (N1727, N1715, N1186, N893, N1511);
buf BUF1 (N1728, N1709);
xor XOR2 (N1729, N1725, N929);
buf BUF1 (N1730, N1713);
not NOT1 (N1731, N1726);
buf BUF1 (N1732, N1720);
nor NOR4 (N1733, N1728, N196, N1427, N695);
not NOT1 (N1734, N1723);
nand NAND3 (N1735, N1727, N26, N1154);
buf BUF1 (N1736, N1730);
and AND3 (N1737, N1704, N1246, N1699);
or OR3 (N1738, N1737, N578, N1169);
xor XOR2 (N1739, N1731, N1256);
buf BUF1 (N1740, N1739);
xor XOR2 (N1741, N1736, N1151);
or OR2 (N1742, N1740, N604);
buf BUF1 (N1743, N1741);
not NOT1 (N1744, N1732);
nor NOR3 (N1745, N1734, N899, N609);
and AND4 (N1746, N1721, N1208, N373, N1081);
xor XOR2 (N1747, N1738, N711);
buf BUF1 (N1748, N1735);
nand NAND2 (N1749, N1745, N1554);
xor XOR2 (N1750, N1747, N1094);
or OR2 (N1751, N1750, N1694);
nand NAND3 (N1752, N1746, N1580, N906);
xor XOR2 (N1753, N1748, N1545);
xor XOR2 (N1754, N1752, N1320);
or OR3 (N1755, N1749, N962, N1309);
nor NOR4 (N1756, N1744, N903, N1694, N33);
nand NAND3 (N1757, N1724, N956, N113);
or OR2 (N1758, N1753, N1638);
and AND4 (N1759, N1742, N991, N900, N268);
not NOT1 (N1760, N1751);
nor NOR4 (N1761, N1760, N1085, N761, N852);
or OR2 (N1762, N1729, N1667);
xor XOR2 (N1763, N1758, N618);
nand NAND4 (N1764, N1754, N1536, N786, N718);
nor NOR4 (N1765, N1762, N623, N922, N1367);
nand NAND2 (N1766, N1759, N1357);
buf BUF1 (N1767, N1755);
or OR4 (N1768, N1766, N1043, N210, N580);
xor XOR2 (N1769, N1765, N1093);
not NOT1 (N1770, N1733);
or OR4 (N1771, N1769, N1341, N1107, N181);
and AND4 (N1772, N1761, N1529, N614, N1096);
nand NAND2 (N1773, N1764, N117);
nand NAND2 (N1774, N1756, N995);
and AND2 (N1775, N1770, N336);
or OR4 (N1776, N1763, N1144, N1195, N840);
and AND3 (N1777, N1775, N1717, N1135);
nor NOR4 (N1778, N1743, N678, N90, N284);
xor XOR2 (N1779, N1768, N82);
nor NOR4 (N1780, N1773, N24, N308, N1052);
or OR2 (N1781, N1776, N790);
nor NOR2 (N1782, N1779, N1001);
xor XOR2 (N1783, N1777, N1566);
buf BUF1 (N1784, N1772);
nand NAND3 (N1785, N1774, N1544, N7);
or OR3 (N1786, N1782, N668, N1096);
nor NOR4 (N1787, N1781, N1486, N1415, N1557);
nand NAND3 (N1788, N1785, N1727, N1357);
nand NAND3 (N1789, N1787, N581, N1367);
nand NAND2 (N1790, N1788, N961);
buf BUF1 (N1791, N1780);
not NOT1 (N1792, N1778);
xor XOR2 (N1793, N1771, N20);
nor NOR2 (N1794, N1793, N1002);
xor XOR2 (N1795, N1784, N996);
or OR4 (N1796, N1794, N1617, N1700, N1585);
and AND2 (N1797, N1767, N1316);
not NOT1 (N1798, N1797);
xor XOR2 (N1799, N1757, N1169);
xor XOR2 (N1800, N1791, N1066);
xor XOR2 (N1801, N1792, N282);
xor XOR2 (N1802, N1800, N1355);
buf BUF1 (N1803, N1786);
or OR2 (N1804, N1799, N1442);
not NOT1 (N1805, N1804);
or OR3 (N1806, N1789, N471, N1783);
and AND2 (N1807, N986, N1690);
nand NAND3 (N1808, N1807, N970, N904);
nor NOR3 (N1809, N1808, N341, N1754);
nor NOR3 (N1810, N1802, N726, N686);
buf BUF1 (N1811, N1809);
nand NAND4 (N1812, N1805, N152, N357, N89);
nor NOR2 (N1813, N1798, N326);
and AND3 (N1814, N1803, N235, N865);
not NOT1 (N1815, N1790);
and AND2 (N1816, N1801, N1244);
nand NAND4 (N1817, N1795, N1036, N1128, N1586);
not NOT1 (N1818, N1810);
nand NAND3 (N1819, N1818, N100, N6);
xor XOR2 (N1820, N1811, N584);
xor XOR2 (N1821, N1817, N1246);
or OR4 (N1822, N1820, N179, N1566, N1661);
nand NAND3 (N1823, N1816, N328, N537);
and AND3 (N1824, N1822, N671, N588);
xor XOR2 (N1825, N1819, N525);
nand NAND3 (N1826, N1825, N1591, N1635);
and AND2 (N1827, N1813, N1210);
nand NAND2 (N1828, N1823, N1789);
or OR3 (N1829, N1826, N1408, N806);
and AND4 (N1830, N1827, N1140, N542, N1013);
buf BUF1 (N1831, N1830);
nor NOR3 (N1832, N1829, N526, N1274);
buf BUF1 (N1833, N1821);
and AND2 (N1834, N1824, N973);
not NOT1 (N1835, N1832);
nand NAND4 (N1836, N1812, N1025, N1192, N1203);
nor NOR2 (N1837, N1831, N129);
not NOT1 (N1838, N1835);
xor XOR2 (N1839, N1815, N1715);
nand NAND2 (N1840, N1837, N231);
and AND4 (N1841, N1840, N158, N805, N413);
xor XOR2 (N1842, N1834, N1165);
buf BUF1 (N1843, N1836);
or OR2 (N1844, N1814, N1604);
xor XOR2 (N1845, N1796, N1285);
or OR3 (N1846, N1806, N1294, N1762);
buf BUF1 (N1847, N1846);
nand NAND2 (N1848, N1842, N1178);
or OR2 (N1849, N1843, N1757);
nand NAND3 (N1850, N1833, N72, N776);
or OR3 (N1851, N1839, N962, N1565);
or OR2 (N1852, N1848, N1694);
and AND3 (N1853, N1844, N256, N829);
nand NAND3 (N1854, N1845, N560, N1483);
and AND4 (N1855, N1849, N727, N724, N1764);
and AND2 (N1856, N1841, N1412);
and AND4 (N1857, N1853, N211, N819, N1712);
and AND3 (N1858, N1855, N826, N1668);
xor XOR2 (N1859, N1856, N106);
nand NAND3 (N1860, N1854, N552, N1393);
not NOT1 (N1861, N1828);
and AND3 (N1862, N1859, N1418, N1321);
nand NAND4 (N1863, N1852, N1000, N1559, N1773);
and AND2 (N1864, N1863, N130);
nor NOR3 (N1865, N1861, N1516, N74);
and AND2 (N1866, N1864, N1788);
not NOT1 (N1867, N1858);
and AND2 (N1868, N1866, N1296);
xor XOR2 (N1869, N1838, N907);
buf BUF1 (N1870, N1862);
and AND4 (N1871, N1847, N334, N541, N846);
nor NOR4 (N1872, N1860, N1230, N851, N1015);
and AND4 (N1873, N1867, N1326, N575, N383);
and AND2 (N1874, N1871, N1848);
not NOT1 (N1875, N1851);
nand NAND2 (N1876, N1850, N750);
and AND4 (N1877, N1870, N402, N1633, N1545);
nand NAND2 (N1878, N1873, N1054);
or OR2 (N1879, N1877, N838);
xor XOR2 (N1880, N1876, N747);
not NOT1 (N1881, N1878);
buf BUF1 (N1882, N1872);
and AND4 (N1883, N1857, N1337, N954, N661);
xor XOR2 (N1884, N1875, N1590);
not NOT1 (N1885, N1881);
nand NAND4 (N1886, N1880, N1050, N1460, N123);
nand NAND3 (N1887, N1874, N16, N1451);
and AND4 (N1888, N1886, N1358, N1785, N788);
and AND4 (N1889, N1882, N284, N135, N1607);
not NOT1 (N1890, N1879);
nand NAND3 (N1891, N1884, N800, N1589);
nor NOR3 (N1892, N1865, N1519, N13);
or OR4 (N1893, N1883, N853, N1375, N1458);
not NOT1 (N1894, N1889);
buf BUF1 (N1895, N1888);
and AND4 (N1896, N1869, N1134, N1765, N1858);
and AND2 (N1897, N1868, N612);
buf BUF1 (N1898, N1890);
nand NAND3 (N1899, N1897, N1868, N595);
buf BUF1 (N1900, N1887);
and AND3 (N1901, N1898, N1206, N796);
nor NOR3 (N1902, N1893, N417, N1579);
buf BUF1 (N1903, N1891);
xor XOR2 (N1904, N1903, N610);
or OR3 (N1905, N1904, N1730, N781);
buf BUF1 (N1906, N1894);
not NOT1 (N1907, N1902);
nor NOR2 (N1908, N1901, N1194);
nand NAND4 (N1909, N1885, N827, N1409, N420);
buf BUF1 (N1910, N1900);
xor XOR2 (N1911, N1910, N303);
or OR2 (N1912, N1908, N1178);
or OR4 (N1913, N1906, N1085, N837, N1836);
buf BUF1 (N1914, N1895);
not NOT1 (N1915, N1907);
or OR4 (N1916, N1892, N520, N1587, N1844);
xor XOR2 (N1917, N1905, N310);
not NOT1 (N1918, N1911);
and AND4 (N1919, N1916, N1269, N1446, N884);
buf BUF1 (N1920, N1914);
nor NOR4 (N1921, N1920, N313, N133, N1704);
and AND2 (N1922, N1909, N530);
nor NOR4 (N1923, N1922, N1794, N1138, N722);
or OR2 (N1924, N1915, N1382);
and AND3 (N1925, N1921, N990, N1488);
nand NAND4 (N1926, N1919, N1019, N930, N931);
buf BUF1 (N1927, N1913);
or OR4 (N1928, N1912, N1915, N1291, N1869);
or OR2 (N1929, N1927, N1816);
nand NAND4 (N1930, N1924, N1291, N660, N258);
nand NAND2 (N1931, N1899, N1296);
not NOT1 (N1932, N1917);
or OR3 (N1933, N1932, N938, N986);
or OR2 (N1934, N1925, N574);
buf BUF1 (N1935, N1926);
xor XOR2 (N1936, N1896, N226);
and AND4 (N1937, N1923, N1449, N823, N1780);
buf BUF1 (N1938, N1934);
nand NAND2 (N1939, N1918, N1190);
or OR2 (N1940, N1938, N460);
and AND2 (N1941, N1940, N883);
not NOT1 (N1942, N1931);
or OR3 (N1943, N1939, N209, N523);
or OR2 (N1944, N1941, N516);
not NOT1 (N1945, N1930);
nand NAND2 (N1946, N1945, N773);
and AND4 (N1947, N1935, N317, N849, N225);
not NOT1 (N1948, N1944);
buf BUF1 (N1949, N1933);
nand NAND3 (N1950, N1947, N353, N1613);
not NOT1 (N1951, N1937);
and AND2 (N1952, N1942, N306);
and AND4 (N1953, N1950, N817, N438, N1242);
buf BUF1 (N1954, N1943);
not NOT1 (N1955, N1952);
and AND2 (N1956, N1949, N829);
nand NAND2 (N1957, N1948, N763);
nand NAND3 (N1958, N1956, N1836, N901);
or OR3 (N1959, N1936, N304, N1173);
not NOT1 (N1960, N1929);
nand NAND3 (N1961, N1957, N1052, N29);
nor NOR4 (N1962, N1959, N306, N1011, N184);
nor NOR3 (N1963, N1951, N1249, N1429);
xor XOR2 (N1964, N1962, N1954);
or OR3 (N1965, N981, N666, N844);
or OR3 (N1966, N1960, N775, N1846);
not NOT1 (N1967, N1965);
buf BUF1 (N1968, N1946);
xor XOR2 (N1969, N1966, N1281);
buf BUF1 (N1970, N1969);
nor NOR3 (N1971, N1967, N1757, N177);
and AND2 (N1972, N1961, N386);
or OR3 (N1973, N1963, N1152, N804);
nor NOR3 (N1974, N1972, N1765, N799);
and AND3 (N1975, N1973, N850, N1836);
not NOT1 (N1976, N1968);
nand NAND2 (N1977, N1971, N1787);
not NOT1 (N1978, N1928);
nor NOR3 (N1979, N1975, N239, N1685);
nor NOR2 (N1980, N1979, N1329);
not NOT1 (N1981, N1953);
and AND2 (N1982, N1980, N1684);
or OR4 (N1983, N1976, N1738, N1710, N918);
buf BUF1 (N1984, N1978);
nand NAND4 (N1985, N1964, N225, N678, N1083);
not NOT1 (N1986, N1958);
or OR2 (N1987, N1986, N440);
not NOT1 (N1988, N1974);
buf BUF1 (N1989, N1981);
nand NAND3 (N1990, N1970, N216, N987);
or OR2 (N1991, N1988, N360);
xor XOR2 (N1992, N1989, N925);
or OR2 (N1993, N1984, N1178);
or OR2 (N1994, N1982, N1625);
xor XOR2 (N1995, N1992, N1011);
and AND2 (N1996, N1990, N1010);
or OR2 (N1997, N1955, N317);
nand NAND3 (N1998, N1985, N803, N1010);
or OR4 (N1999, N1993, N1254, N533, N1435);
nand NAND4 (N2000, N1991, N1766, N1485, N803);
xor XOR2 (N2001, N1996, N973);
xor XOR2 (N2002, N1977, N1709);
not NOT1 (N2003, N1987);
or OR2 (N2004, N1999, N856);
not NOT1 (N2005, N2002);
nand NAND3 (N2006, N2005, N1003, N115);
or OR3 (N2007, N1983, N223, N552);
nor NOR2 (N2008, N2006, N1436);
or OR4 (N2009, N2008, N1460, N51, N1155);
xor XOR2 (N2010, N2009, N713);
xor XOR2 (N2011, N1997, N616);
nor NOR3 (N2012, N2010, N1254, N75);
or OR4 (N2013, N1998, N449, N1759, N1223);
nand NAND2 (N2014, N2001, N1030);
not NOT1 (N2015, N2011);
buf BUF1 (N2016, N2004);
nor NOR4 (N2017, N2014, N1779, N697, N308);
nor NOR2 (N2018, N2015, N738);
xor XOR2 (N2019, N2007, N1365);
nand NAND4 (N2020, N2018, N642, N1803, N1835);
nor NOR2 (N2021, N2013, N1312);
xor XOR2 (N2022, N2020, N1503);
and AND2 (N2023, N2000, N1040);
nor NOR2 (N2024, N2022, N555);
or OR2 (N2025, N2021, N1732);
nor NOR3 (N2026, N2003, N788, N918);
buf BUF1 (N2027, N1994);
nand NAND4 (N2028, N2017, N1547, N1570, N524);
not NOT1 (N2029, N2023);
nand NAND4 (N2030, N2012, N1642, N1751, N140);
xor XOR2 (N2031, N2025, N1537);
buf BUF1 (N2032, N2016);
not NOT1 (N2033, N2027);
nor NOR2 (N2034, N2026, N381);
xor XOR2 (N2035, N2028, N819);
buf BUF1 (N2036, N2030);
not NOT1 (N2037, N1995);
xor XOR2 (N2038, N2035, N952);
xor XOR2 (N2039, N2033, N1565);
or OR2 (N2040, N2031, N1257);
xor XOR2 (N2041, N2032, N69);
or OR2 (N2042, N2029, N641);
buf BUF1 (N2043, N2024);
xor XOR2 (N2044, N2042, N1536);
nand NAND2 (N2045, N2044, N1619);
or OR3 (N2046, N2041, N339, N1782);
nor NOR3 (N2047, N2040, N1956, N807);
nor NOR2 (N2048, N2038, N1594);
xor XOR2 (N2049, N2046, N1183);
xor XOR2 (N2050, N2048, N95);
nand NAND3 (N2051, N2050, N1906, N159);
and AND2 (N2052, N2051, N951);
nor NOR2 (N2053, N2045, N737);
nand NAND3 (N2054, N2043, N791, N703);
xor XOR2 (N2055, N2019, N553);
or OR4 (N2056, N2049, N1284, N1350, N394);
nor NOR4 (N2057, N2034, N1052, N612, N1852);
nor NOR4 (N2058, N2047, N2045, N1582, N690);
not NOT1 (N2059, N2036);
and AND2 (N2060, N2055, N574);
xor XOR2 (N2061, N2053, N212);
nor NOR2 (N2062, N2037, N1277);
xor XOR2 (N2063, N2061, N641);
buf BUF1 (N2064, N2062);
not NOT1 (N2065, N2060);
nor NOR2 (N2066, N2064, N1116);
nand NAND4 (N2067, N2059, N1900, N616, N958);
or OR3 (N2068, N2065, N1157, N1582);
buf BUF1 (N2069, N2067);
nand NAND4 (N2070, N2057, N1995, N1599, N1068);
xor XOR2 (N2071, N2052, N1120);
or OR3 (N2072, N2056, N888, N2052);
buf BUF1 (N2073, N2066);
and AND3 (N2074, N2071, N544, N2023);
nand NAND3 (N2075, N2070, N926, N1653);
nand NAND3 (N2076, N2063, N1446, N1750);
xor XOR2 (N2077, N2074, N1824);
and AND3 (N2078, N2039, N1671, N1790);
and AND3 (N2079, N2075, N1261, N851);
nand NAND4 (N2080, N2072, N77, N955, N1791);
not NOT1 (N2081, N2076);
and AND2 (N2082, N2058, N1894);
xor XOR2 (N2083, N2068, N1380);
xor XOR2 (N2084, N2073, N848);
nand NAND2 (N2085, N2084, N1323);
buf BUF1 (N2086, N2069);
nor NOR4 (N2087, N2078, N1566, N1015, N1782);
and AND3 (N2088, N2082, N1194, N866);
or OR2 (N2089, N2079, N757);
nand NAND2 (N2090, N2077, N2084);
buf BUF1 (N2091, N2088);
xor XOR2 (N2092, N2081, N55);
or OR3 (N2093, N2054, N161, N242);
not NOT1 (N2094, N2086);
xor XOR2 (N2095, N2093, N1743);
buf BUF1 (N2096, N2087);
buf BUF1 (N2097, N2095);
buf BUF1 (N2098, N2080);
nand NAND2 (N2099, N2091, N2068);
not NOT1 (N2100, N2098);
xor XOR2 (N2101, N2099, N1585);
nor NOR3 (N2102, N2097, N299, N977);
nor NOR2 (N2103, N2102, N170);
not NOT1 (N2104, N2096);
not NOT1 (N2105, N2104);
nor NOR2 (N2106, N2083, N1766);
nand NAND2 (N2107, N2092, N1574);
nand NAND3 (N2108, N2103, N820, N228);
or OR3 (N2109, N2100, N655, N1839);
xor XOR2 (N2110, N2094, N462);
and AND3 (N2111, N2107, N1839, N1603);
nor NOR3 (N2112, N2108, N769, N800);
or OR3 (N2113, N2090, N1131, N1943);
or OR2 (N2114, N2089, N210);
nand NAND4 (N2115, N2111, N1075, N1467, N1671);
and AND4 (N2116, N2115, N152, N1635, N1291);
and AND4 (N2117, N2116, N809, N1865, N1229);
nand NAND4 (N2118, N2110, N384, N959, N351);
not NOT1 (N2119, N2117);
buf BUF1 (N2120, N2114);
nand NAND2 (N2121, N2105, N1466);
nand NAND2 (N2122, N2119, N1251);
or OR2 (N2123, N2106, N550);
nand NAND3 (N2124, N2101, N1605, N1726);
and AND3 (N2125, N2124, N1196, N102);
xor XOR2 (N2126, N2118, N1914);
nand NAND2 (N2127, N2113, N700);
nor NOR3 (N2128, N2123, N2106, N736);
not NOT1 (N2129, N2109);
xor XOR2 (N2130, N2112, N1468);
xor XOR2 (N2131, N2129, N706);
and AND3 (N2132, N2128, N129, N615);
or OR2 (N2133, N2127, N69);
buf BUF1 (N2134, N2126);
and AND4 (N2135, N2120, N541, N1323, N1876);
not NOT1 (N2136, N2132);
or OR4 (N2137, N2125, N682, N1209, N1868);
nand NAND4 (N2138, N2134, N1520, N980, N150);
and AND4 (N2139, N2130, N1960, N1823, N579);
not NOT1 (N2140, N2138);
buf BUF1 (N2141, N2122);
xor XOR2 (N2142, N2121, N1132);
nor NOR3 (N2143, N2137, N810, N1177);
and AND3 (N2144, N2143, N1743, N75);
xor XOR2 (N2145, N2140, N402);
buf BUF1 (N2146, N2145);
nand NAND4 (N2147, N2144, N401, N780, N796);
and AND2 (N2148, N2085, N1904);
and AND4 (N2149, N2142, N1465, N154, N329);
or OR4 (N2150, N2147, N1761, N1490, N436);
and AND3 (N2151, N2135, N1334, N595);
nand NAND2 (N2152, N2139, N226);
buf BUF1 (N2153, N2149);
buf BUF1 (N2154, N2141);
and AND3 (N2155, N2151, N278, N1294);
not NOT1 (N2156, N2152);
or OR3 (N2157, N2131, N1967, N268);
not NOT1 (N2158, N2136);
nor NOR4 (N2159, N2146, N1, N653, N2017);
not NOT1 (N2160, N2150);
and AND3 (N2161, N2153, N346, N901);
or OR3 (N2162, N2157, N1448, N1513);
nor NOR3 (N2163, N2160, N961, N170);
xor XOR2 (N2164, N2158, N170);
nor NOR3 (N2165, N2154, N1526, N491);
buf BUF1 (N2166, N2133);
not NOT1 (N2167, N2148);
or OR2 (N2168, N2159, N1267);
buf BUF1 (N2169, N2155);
nor NOR3 (N2170, N2164, N2035, N53);
and AND3 (N2171, N2167, N1996, N1195);
and AND2 (N2172, N2169, N141);
buf BUF1 (N2173, N2165);
buf BUF1 (N2174, N2173);
or OR2 (N2175, N2172, N1881);
nor NOR2 (N2176, N2174, N1361);
or OR3 (N2177, N2176, N855, N475);
not NOT1 (N2178, N2163);
not NOT1 (N2179, N2162);
not NOT1 (N2180, N2156);
nor NOR2 (N2181, N2178, N1313);
and AND2 (N2182, N2179, N330);
buf BUF1 (N2183, N2182);
or OR3 (N2184, N2175, N1601, N176);
nand NAND4 (N2185, N2170, N151, N1854, N1408);
buf BUF1 (N2186, N2180);
not NOT1 (N2187, N2171);
and AND3 (N2188, N2185, N1954, N438);
nor NOR2 (N2189, N2186, N886);
xor XOR2 (N2190, N2177, N961);
nor NOR3 (N2191, N2183, N2189, N2132);
and AND2 (N2192, N865, N578);
and AND4 (N2193, N2166, N229, N2044, N479);
nor NOR2 (N2194, N2190, N1552);
buf BUF1 (N2195, N2187);
nor NOR4 (N2196, N2188, N1333, N1289, N1484);
or OR4 (N2197, N2196, N576, N657, N1368);
and AND2 (N2198, N2168, N875);
nand NAND3 (N2199, N2161, N2164, N1466);
or OR2 (N2200, N2195, N2130);
xor XOR2 (N2201, N2199, N497);
xor XOR2 (N2202, N2192, N1524);
not NOT1 (N2203, N2198);
buf BUF1 (N2204, N2184);
not NOT1 (N2205, N2191);
nor NOR2 (N2206, N2181, N837);
xor XOR2 (N2207, N2206, N2060);
nand NAND3 (N2208, N2194, N2192, N850);
or OR3 (N2209, N2204, N2178, N144);
xor XOR2 (N2210, N2207, N706);
nor NOR2 (N2211, N2209, N1563);
nor NOR2 (N2212, N2197, N2157);
nand NAND4 (N2213, N2208, N676, N992, N589);
or OR3 (N2214, N2205, N749, N1097);
not NOT1 (N2215, N2213);
or OR2 (N2216, N2212, N1);
not NOT1 (N2217, N2214);
nor NOR2 (N2218, N2215, N1885);
nor NOR4 (N2219, N2217, N2, N1818, N725);
nor NOR4 (N2220, N2201, N188, N1309, N302);
not NOT1 (N2221, N2203);
or OR4 (N2222, N2218, N83, N721, N1510);
or OR2 (N2223, N2220, N207);
not NOT1 (N2224, N2221);
nand NAND4 (N2225, N2216, N92, N538, N1632);
or OR2 (N2226, N2222, N565);
nand NAND2 (N2227, N2200, N2155);
and AND2 (N2228, N2211, N1453);
nand NAND4 (N2229, N2227, N1909, N1086, N1969);
and AND2 (N2230, N2228, N300);
or OR4 (N2231, N2224, N1115, N1249, N1899);
or OR2 (N2232, N2219, N964);
xor XOR2 (N2233, N2232, N1476);
buf BUF1 (N2234, N2202);
and AND3 (N2235, N2229, N442, N949);
buf BUF1 (N2236, N2210);
and AND2 (N2237, N2230, N2176);
xor XOR2 (N2238, N2237, N2154);
not NOT1 (N2239, N2193);
buf BUF1 (N2240, N2226);
not NOT1 (N2241, N2235);
or OR3 (N2242, N2234, N642, N1273);
and AND3 (N2243, N2241, N1129, N1255);
not NOT1 (N2244, N2233);
nand NAND2 (N2245, N2239, N1593);
buf BUF1 (N2246, N2244);
not NOT1 (N2247, N2223);
and AND4 (N2248, N2246, N2076, N1643, N324);
or OR4 (N2249, N2242, N1926, N452, N198);
or OR4 (N2250, N2225, N1252, N735, N885);
xor XOR2 (N2251, N2240, N431);
xor XOR2 (N2252, N2250, N186);
nand NAND3 (N2253, N2249, N395, N1355);
nand NAND3 (N2254, N2236, N400, N2130);
nand NAND4 (N2255, N2245, N1751, N660, N1199);
or OR4 (N2256, N2247, N1541, N2052, N1557);
and AND3 (N2257, N2253, N1647, N1148);
buf BUF1 (N2258, N2252);
and AND3 (N2259, N2248, N1733, N1985);
or OR3 (N2260, N2256, N1724, N125);
not NOT1 (N2261, N2243);
nor NOR3 (N2262, N2238, N850, N2009);
or OR3 (N2263, N2260, N174, N1754);
not NOT1 (N2264, N2259);
and AND4 (N2265, N2251, N568, N747, N762);
nor NOR4 (N2266, N2254, N952, N2189, N833);
nor NOR3 (N2267, N2231, N758, N1776);
buf BUF1 (N2268, N2255);
and AND4 (N2269, N2266, N760, N776, N1202);
xor XOR2 (N2270, N2265, N1692);
nor NOR4 (N2271, N2263, N1454, N483, N284);
and AND4 (N2272, N2270, N1277, N250, N791);
not NOT1 (N2273, N2261);
and AND2 (N2274, N2268, N2065);
and AND4 (N2275, N2262, N1867, N1557, N759);
nor NOR3 (N2276, N2264, N1456, N857);
or OR3 (N2277, N2257, N1583, N890);
buf BUF1 (N2278, N2271);
or OR4 (N2279, N2272, N663, N2236, N2039);
nor NOR3 (N2280, N2278, N131, N520);
nor NOR4 (N2281, N2277, N1591, N711, N2255);
and AND4 (N2282, N2281, N345, N1491, N1313);
not NOT1 (N2283, N2279);
buf BUF1 (N2284, N2282);
and AND4 (N2285, N2275, N221, N956, N585);
xor XOR2 (N2286, N2273, N2179);
nor NOR2 (N2287, N2269, N407);
not NOT1 (N2288, N2283);
nor NOR2 (N2289, N2284, N670);
nand NAND3 (N2290, N2288, N640, N630);
buf BUF1 (N2291, N2287);
nand NAND3 (N2292, N2291, N743, N1722);
not NOT1 (N2293, N2267);
or OR3 (N2294, N2292, N2095, N1087);
xor XOR2 (N2295, N2293, N147);
not NOT1 (N2296, N2294);
buf BUF1 (N2297, N2280);
or OR4 (N2298, N2297, N656, N1449, N1416);
or OR2 (N2299, N2289, N252);
xor XOR2 (N2300, N2274, N2208);
nor NOR3 (N2301, N2300, N1677, N680);
or OR2 (N2302, N2301, N2203);
nor NOR3 (N2303, N2298, N996, N585);
buf BUF1 (N2304, N2295);
xor XOR2 (N2305, N2276, N17);
nand NAND4 (N2306, N2303, N773, N1602, N2160);
buf BUF1 (N2307, N2290);
buf BUF1 (N2308, N2286);
nand NAND4 (N2309, N2299, N1052, N1688, N2001);
nor NOR3 (N2310, N2258, N302, N1428);
xor XOR2 (N2311, N2308, N1783);
buf BUF1 (N2312, N2309);
and AND4 (N2313, N2304, N645, N1383, N563);
not NOT1 (N2314, N2307);
nor NOR4 (N2315, N2313, N1570, N141, N1493);
and AND2 (N2316, N2305, N1158);
buf BUF1 (N2317, N2302);
xor XOR2 (N2318, N2296, N1389);
nor NOR3 (N2319, N2318, N1359, N2126);
nand NAND2 (N2320, N2317, N1763);
or OR2 (N2321, N2285, N1993);
nand NAND4 (N2322, N2306, N1393, N193, N497);
and AND3 (N2323, N2315, N852, N2206);
xor XOR2 (N2324, N2314, N1705);
and AND4 (N2325, N2324, N445, N99, N705);
or OR2 (N2326, N2319, N2132);
or OR4 (N2327, N2320, N1997, N934, N329);
nand NAND3 (N2328, N2325, N1827, N828);
buf BUF1 (N2329, N2312);
xor XOR2 (N2330, N2327, N339);
or OR4 (N2331, N2329, N651, N745, N673);
and AND3 (N2332, N2321, N257, N192);
or OR4 (N2333, N2328, N40, N1457, N808);
and AND2 (N2334, N2326, N1835);
and AND3 (N2335, N2316, N646, N2321);
not NOT1 (N2336, N2330);
xor XOR2 (N2337, N2334, N201);
xor XOR2 (N2338, N2336, N1676);
or OR4 (N2339, N2323, N966, N767, N259);
not NOT1 (N2340, N2311);
nand NAND2 (N2341, N2331, N417);
nor NOR3 (N2342, N2337, N491, N2077);
and AND3 (N2343, N2333, N1706, N645);
not NOT1 (N2344, N2332);
buf BUF1 (N2345, N2341);
and AND4 (N2346, N2344, N1293, N1973, N2110);
nand NAND2 (N2347, N2343, N2332);
and AND3 (N2348, N2339, N1123, N816);
and AND2 (N2349, N2338, N910);
and AND2 (N2350, N2340, N1419);
nor NOR4 (N2351, N2346, N419, N16, N1087);
buf BUF1 (N2352, N2348);
or OR2 (N2353, N2347, N9);
nand NAND2 (N2354, N2342, N249);
buf BUF1 (N2355, N2354);
nor NOR3 (N2356, N2349, N37, N740);
nand NAND3 (N2357, N2355, N1967, N170);
buf BUF1 (N2358, N2353);
buf BUF1 (N2359, N2322);
xor XOR2 (N2360, N2352, N231);
xor XOR2 (N2361, N2360, N1179);
nor NOR4 (N2362, N2335, N1489, N1264, N572);
xor XOR2 (N2363, N2361, N1829);
nand NAND2 (N2364, N2345, N2196);
xor XOR2 (N2365, N2362, N1017);
not NOT1 (N2366, N2363);
not NOT1 (N2367, N2357);
nand NAND3 (N2368, N2350, N1093, N1993);
nand NAND2 (N2369, N2365, N1890);
xor XOR2 (N2370, N2351, N1314);
or OR3 (N2371, N2366, N1004, N1838);
nand NAND4 (N2372, N2359, N349, N1231, N1074);
xor XOR2 (N2373, N2356, N61);
buf BUF1 (N2374, N2310);
xor XOR2 (N2375, N2373, N1405);
xor XOR2 (N2376, N2358, N2155);
xor XOR2 (N2377, N2367, N79);
and AND4 (N2378, N2372, N1585, N1727, N1992);
or OR4 (N2379, N2374, N1018, N2229, N2134);
buf BUF1 (N2380, N2369);
nand NAND3 (N2381, N2380, N454, N703);
nor NOR3 (N2382, N2381, N771, N2229);
buf BUF1 (N2383, N2378);
not NOT1 (N2384, N2364);
xor XOR2 (N2385, N2384, N1971);
not NOT1 (N2386, N2375);
and AND2 (N2387, N2368, N2218);
buf BUF1 (N2388, N2387);
nor NOR2 (N2389, N2379, N120);
not NOT1 (N2390, N2377);
not NOT1 (N2391, N2371);
and AND3 (N2392, N2383, N448, N2186);
xor XOR2 (N2393, N2385, N197);
nor NOR4 (N2394, N2382, N1537, N2100, N1426);
buf BUF1 (N2395, N2376);
buf BUF1 (N2396, N2388);
and AND2 (N2397, N2391, N2039);
and AND2 (N2398, N2393, N172);
not NOT1 (N2399, N2396);
nand NAND4 (N2400, N2397, N2330, N2105, N274);
nand NAND2 (N2401, N2394, N899);
nand NAND3 (N2402, N2398, N341, N631);
xor XOR2 (N2403, N2386, N1613);
and AND4 (N2404, N2400, N1648, N271, N1964);
xor XOR2 (N2405, N2390, N1279);
nand NAND3 (N2406, N2389, N1779, N1594);
buf BUF1 (N2407, N2392);
buf BUF1 (N2408, N2401);
or OR2 (N2409, N2405, N684);
and AND3 (N2410, N2409, N2354, N2150);
not NOT1 (N2411, N2408);
and AND4 (N2412, N2370, N1348, N1359, N1645);
xor XOR2 (N2413, N2395, N314);
or OR2 (N2414, N2412, N840);
buf BUF1 (N2415, N2413);
nand NAND3 (N2416, N2399, N1395, N1186);
and AND4 (N2417, N2407, N1938, N859, N630);
not NOT1 (N2418, N2417);
and AND3 (N2419, N2410, N1665, N2174);
and AND3 (N2420, N2404, N2026, N714);
or OR3 (N2421, N2418, N242, N636);
nor NOR3 (N2422, N2411, N778, N335);
not NOT1 (N2423, N2402);
or OR4 (N2424, N2416, N79, N2239, N505);
xor XOR2 (N2425, N2406, N1628);
or OR3 (N2426, N2423, N887, N22);
buf BUF1 (N2427, N2419);
and AND3 (N2428, N2426, N2178, N1005);
or OR2 (N2429, N2424, N862);
nand NAND4 (N2430, N2403, N1564, N798, N1723);
and AND4 (N2431, N2415, N1694, N1343, N2111);
and AND2 (N2432, N2425, N2369);
nand NAND4 (N2433, N2420, N470, N1025, N1211);
and AND3 (N2434, N2414, N567, N1855);
xor XOR2 (N2435, N2421, N1618);
nand NAND2 (N2436, N2429, N1385);
nor NOR2 (N2437, N2431, N2246);
xor XOR2 (N2438, N2430, N2135);
nand NAND2 (N2439, N2427, N1014);
or OR2 (N2440, N2436, N1400);
xor XOR2 (N2441, N2428, N1097);
nor NOR3 (N2442, N2434, N476, N588);
nor NOR3 (N2443, N2438, N2180, N2362);
not NOT1 (N2444, N2433);
and AND2 (N2445, N2444, N1241);
and AND2 (N2446, N2443, N124);
nor NOR2 (N2447, N2437, N578);
nand NAND2 (N2448, N2441, N1954);
nor NOR2 (N2449, N2446, N1955);
nand NAND4 (N2450, N2449, N1274, N1582, N2445);
xor XOR2 (N2451, N1489, N430);
and AND2 (N2452, N2432, N394);
buf BUF1 (N2453, N2435);
or OR3 (N2454, N2452, N1289, N615);
nor NOR3 (N2455, N2453, N1397, N2430);
not NOT1 (N2456, N2422);
or OR2 (N2457, N2448, N1665);
and AND2 (N2458, N2442, N56);
xor XOR2 (N2459, N2458, N255);
buf BUF1 (N2460, N2440);
and AND4 (N2461, N2439, N203, N1029, N1526);
nor NOR4 (N2462, N2451, N1594, N826, N611);
not NOT1 (N2463, N2461);
buf BUF1 (N2464, N2447);
or OR2 (N2465, N2455, N533);
nor NOR2 (N2466, N2459, N2185);
nand NAND4 (N2467, N2465, N582, N1045, N425);
xor XOR2 (N2468, N2456, N1894);
or OR4 (N2469, N2466, N1482, N722, N351);
nor NOR2 (N2470, N2457, N1684);
and AND4 (N2471, N2463, N561, N369, N538);
nand NAND4 (N2472, N2464, N2205, N796, N737);
xor XOR2 (N2473, N2467, N1865);
buf BUF1 (N2474, N2473);
nand NAND2 (N2475, N2462, N1906);
buf BUF1 (N2476, N2454);
or OR3 (N2477, N2470, N2121, N329);
not NOT1 (N2478, N2471);
nor NOR2 (N2479, N2460, N1045);
buf BUF1 (N2480, N2479);
nand NAND2 (N2481, N2468, N142);
nand NAND4 (N2482, N2472, N2435, N1376, N1661);
and AND2 (N2483, N2481, N1005);
nand NAND4 (N2484, N2480, N325, N1236, N2271);
nor NOR2 (N2485, N2475, N1914);
or OR2 (N2486, N2474, N861);
and AND2 (N2487, N2478, N2019);
nand NAND4 (N2488, N2469, N2015, N1144, N182);
nand NAND2 (N2489, N2482, N1938);
buf BUF1 (N2490, N2487);
nand NAND3 (N2491, N2489, N2295, N2139);
not NOT1 (N2492, N2485);
or OR2 (N2493, N2450, N795);
or OR3 (N2494, N2477, N1612, N1671);
xor XOR2 (N2495, N2491, N2241);
not NOT1 (N2496, N2494);
buf BUF1 (N2497, N2484);
not NOT1 (N2498, N2483);
or OR3 (N2499, N2476, N569, N830);
buf BUF1 (N2500, N2490);
and AND4 (N2501, N2488, N171, N1369, N2062);
or OR3 (N2502, N2492, N1897, N290);
or OR3 (N2503, N2501, N2464, N1815);
or OR4 (N2504, N2499, N559, N1369, N1813);
xor XOR2 (N2505, N2504, N650);
or OR4 (N2506, N2495, N1947, N1633, N2418);
buf BUF1 (N2507, N2503);
buf BUF1 (N2508, N2493);
or OR4 (N2509, N2506, N812, N1739, N2498);
xor XOR2 (N2510, N2386, N1657);
nand NAND4 (N2511, N2496, N2031, N1551, N143);
buf BUF1 (N2512, N2509);
nor NOR3 (N2513, N2512, N779, N1817);
buf BUF1 (N2514, N2513);
or OR2 (N2515, N2502, N2094);
nand NAND3 (N2516, N2514, N1912, N288);
not NOT1 (N2517, N2510);
and AND2 (N2518, N2516, N949);
or OR3 (N2519, N2515, N1571, N1426);
nand NAND3 (N2520, N2505, N1593, N2373);
xor XOR2 (N2521, N2518, N2436);
not NOT1 (N2522, N2521);
and AND3 (N2523, N2520, N1108, N2353);
xor XOR2 (N2524, N2486, N232);
buf BUF1 (N2525, N2517);
not NOT1 (N2526, N2500);
or OR3 (N2527, N2523, N2062, N1032);
or OR2 (N2528, N2527, N1394);
nor NOR2 (N2529, N2507, N2126);
nand NAND3 (N2530, N2511, N718, N2448);
nand NAND2 (N2531, N2497, N1164);
xor XOR2 (N2532, N2524, N2491);
and AND4 (N2533, N2528, N763, N142, N1249);
nand NAND4 (N2534, N2522, N1477, N1699, N2383);
nor NOR2 (N2535, N2532, N1389);
xor XOR2 (N2536, N2533, N443);
xor XOR2 (N2537, N2508, N1422);
nand NAND2 (N2538, N2535, N2407);
not NOT1 (N2539, N2538);
or OR2 (N2540, N2534, N2223);
not NOT1 (N2541, N2525);
nor NOR4 (N2542, N2529, N2395, N2258, N608);
nor NOR2 (N2543, N2530, N273);
or OR2 (N2544, N2519, N846);
nor NOR3 (N2545, N2540, N560, N1224);
or OR2 (N2546, N2536, N667);
nor NOR2 (N2547, N2526, N2107);
buf BUF1 (N2548, N2545);
nand NAND4 (N2549, N2531, N1081, N2285, N54);
nand NAND3 (N2550, N2548, N1972, N511);
buf BUF1 (N2551, N2542);
or OR4 (N2552, N2551, N217, N1392, N937);
and AND4 (N2553, N2550, N2143, N2052, N341);
nor NOR2 (N2554, N2543, N2199);
or OR2 (N2555, N2549, N798);
nor NOR2 (N2556, N2539, N1655);
nor NOR2 (N2557, N2544, N1308);
nand NAND3 (N2558, N2554, N1876, N1386);
and AND2 (N2559, N2557, N2293);
buf BUF1 (N2560, N2556);
not NOT1 (N2561, N2552);
and AND4 (N2562, N2546, N1814, N301, N1486);
and AND4 (N2563, N2555, N1077, N2160, N811);
nor NOR2 (N2564, N2541, N610);
not NOT1 (N2565, N2564);
xor XOR2 (N2566, N2565, N1233);
or OR4 (N2567, N2560, N2415, N2029, N612);
nor NOR4 (N2568, N2547, N1153, N186, N1618);
xor XOR2 (N2569, N2567, N1352);
buf BUF1 (N2570, N2562);
and AND4 (N2571, N2553, N762, N2011, N141);
not NOT1 (N2572, N2558);
not NOT1 (N2573, N2572);
buf BUF1 (N2574, N2570);
or OR3 (N2575, N2559, N1703, N2430);
nand NAND3 (N2576, N2571, N39, N1177);
xor XOR2 (N2577, N2573, N153);
or OR2 (N2578, N2563, N880);
xor XOR2 (N2579, N2578, N515);
and AND2 (N2580, N2574, N972);
not NOT1 (N2581, N2577);
not NOT1 (N2582, N2537);
nand NAND2 (N2583, N2575, N1566);
not NOT1 (N2584, N2576);
nand NAND2 (N2585, N2580, N1509);
or OR2 (N2586, N2585, N539);
xor XOR2 (N2587, N2569, N534);
xor XOR2 (N2588, N2561, N568);
xor XOR2 (N2589, N2581, N2500);
and AND2 (N2590, N2586, N1640);
not NOT1 (N2591, N2584);
and AND4 (N2592, N2588, N1068, N1492, N1107);
and AND3 (N2593, N2583, N613, N382);
not NOT1 (N2594, N2590);
xor XOR2 (N2595, N2568, N2465);
and AND2 (N2596, N2589, N1307);
or OR2 (N2597, N2587, N2259);
or OR4 (N2598, N2597, N1359, N157, N2427);
nor NOR3 (N2599, N2582, N120, N2380);
xor XOR2 (N2600, N2579, N635);
nand NAND3 (N2601, N2593, N1951, N1876);
nand NAND3 (N2602, N2601, N1477, N1278);
and AND2 (N2603, N2598, N1783);
and AND2 (N2604, N2600, N435);
or OR2 (N2605, N2604, N1511);
xor XOR2 (N2606, N2592, N771);
or OR2 (N2607, N2603, N969);
xor XOR2 (N2608, N2594, N1908);
not NOT1 (N2609, N2606);
buf BUF1 (N2610, N2596);
buf BUF1 (N2611, N2607);
buf BUF1 (N2612, N2595);
xor XOR2 (N2613, N2612, N1784);
nand NAND4 (N2614, N2611, N1581, N2121, N1609);
buf BUF1 (N2615, N2602);
nand NAND4 (N2616, N2610, N956, N1358, N49);
nand NAND2 (N2617, N2591, N2103);
nor NOR2 (N2618, N2617, N527);
xor XOR2 (N2619, N2618, N698);
or OR3 (N2620, N2609, N1527, N1573);
not NOT1 (N2621, N2619);
or OR2 (N2622, N2608, N524);
and AND2 (N2623, N2566, N2513);
xor XOR2 (N2624, N2621, N1065);
xor XOR2 (N2625, N2599, N290);
nor NOR4 (N2626, N2616, N206, N911, N863);
or OR4 (N2627, N2622, N1117, N279, N2611);
or OR2 (N2628, N2624, N1036);
buf BUF1 (N2629, N2613);
nor NOR4 (N2630, N2623, N2500, N2249, N2207);
nor NOR3 (N2631, N2605, N2255, N6);
xor XOR2 (N2632, N2627, N1110);
nand NAND2 (N2633, N2629, N262);
buf BUF1 (N2634, N2625);
and AND2 (N2635, N2626, N637);
xor XOR2 (N2636, N2615, N2430);
nor NOR4 (N2637, N2635, N1328, N693, N1237);
and AND4 (N2638, N2634, N2277, N350, N1024);
buf BUF1 (N2639, N2637);
not NOT1 (N2640, N2636);
and AND4 (N2641, N2620, N1832, N1828, N1696);
nor NOR2 (N2642, N2631, N1882);
not NOT1 (N2643, N2642);
buf BUF1 (N2644, N2643);
nor NOR4 (N2645, N2638, N2449, N1041, N1572);
or OR3 (N2646, N2639, N1299, N214);
not NOT1 (N2647, N2630);
not NOT1 (N2648, N2633);
xor XOR2 (N2649, N2614, N788);
nand NAND2 (N2650, N2640, N2179);
not NOT1 (N2651, N2641);
buf BUF1 (N2652, N2650);
and AND4 (N2653, N2649, N2336, N2129, N1541);
and AND4 (N2654, N2644, N1693, N2141, N2338);
buf BUF1 (N2655, N2651);
nand NAND4 (N2656, N2628, N216, N2181, N2393);
buf BUF1 (N2657, N2646);
or OR3 (N2658, N2648, N433, N759);
nor NOR3 (N2659, N2656, N2536, N2338);
and AND4 (N2660, N2632, N2060, N2487, N1918);
not NOT1 (N2661, N2655);
not NOT1 (N2662, N2652);
and AND2 (N2663, N2657, N2014);
nor NOR2 (N2664, N2645, N2334);
and AND3 (N2665, N2660, N1129, N53);
nor NOR4 (N2666, N2653, N669, N5, N509);
and AND4 (N2667, N2666, N1255, N2226, N2634);
or OR2 (N2668, N2659, N454);
and AND3 (N2669, N2664, N1322, N587);
buf BUF1 (N2670, N2669);
xor XOR2 (N2671, N2661, N1289);
not NOT1 (N2672, N2670);
and AND4 (N2673, N2662, N1698, N542, N1876);
buf BUF1 (N2674, N2647);
not NOT1 (N2675, N2674);
buf BUF1 (N2676, N2672);
not NOT1 (N2677, N2673);
buf BUF1 (N2678, N2668);
and AND2 (N2679, N2676, N1731);
nand NAND3 (N2680, N2679, N558, N517);
and AND4 (N2681, N2680, N62, N588, N177);
xor XOR2 (N2682, N2678, N77);
nor NOR3 (N2683, N2677, N527, N1929);
or OR2 (N2684, N2663, N1770);
not NOT1 (N2685, N2682);
nor NOR4 (N2686, N2671, N2548, N1311, N2587);
nand NAND2 (N2687, N2684, N1545);
xor XOR2 (N2688, N2667, N1710);
xor XOR2 (N2689, N2685, N1265);
xor XOR2 (N2690, N2689, N2133);
nand NAND3 (N2691, N2687, N493, N1556);
nor NOR3 (N2692, N2665, N2239, N2116);
nor NOR2 (N2693, N2692, N2003);
xor XOR2 (N2694, N2683, N1655);
nand NAND4 (N2695, N2688, N523, N1918, N208);
and AND2 (N2696, N2686, N2017);
not NOT1 (N2697, N2690);
not NOT1 (N2698, N2691);
buf BUF1 (N2699, N2675);
and AND3 (N2700, N2693, N1401, N2616);
nor NOR3 (N2701, N2654, N1066, N1256);
nor NOR4 (N2702, N2681, N149, N1789, N1077);
and AND4 (N2703, N2697, N1827, N1247, N613);
xor XOR2 (N2704, N2658, N1399);
and AND2 (N2705, N2698, N933);
not NOT1 (N2706, N2704);
nor NOR2 (N2707, N2699, N931);
nand NAND2 (N2708, N2702, N415);
nor NOR3 (N2709, N2694, N1999, N1139);
and AND2 (N2710, N2709, N1824);
not NOT1 (N2711, N2700);
buf BUF1 (N2712, N2701);
xor XOR2 (N2713, N2711, N1387);
or OR4 (N2714, N2705, N1447, N813, N1975);
buf BUF1 (N2715, N2713);
nor NOR3 (N2716, N2715, N304, N200);
nor NOR4 (N2717, N2712, N1218, N1758, N1244);
buf BUF1 (N2718, N2708);
xor XOR2 (N2719, N2710, N564);
or OR2 (N2720, N2719, N928);
nor NOR3 (N2721, N2720, N672, N1255);
nand NAND3 (N2722, N2696, N1347, N1987);
nand NAND3 (N2723, N2707, N1923, N2550);
nand NAND4 (N2724, N2716, N379, N2628, N1749);
nor NOR3 (N2725, N2695, N1274, N1778);
not NOT1 (N2726, N2714);
buf BUF1 (N2727, N2721);
and AND2 (N2728, N2725, N2498);
nor NOR3 (N2729, N2703, N2266, N491);
nand NAND3 (N2730, N2717, N1096, N965);
not NOT1 (N2731, N2728);
not NOT1 (N2732, N2727);
nand NAND4 (N2733, N2726, N85, N329, N2276);
buf BUF1 (N2734, N2723);
nor NOR3 (N2735, N2722, N2265, N1631);
or OR4 (N2736, N2724, N1638, N1745, N1185);
and AND2 (N2737, N2706, N1421);
and AND2 (N2738, N2735, N384);
xor XOR2 (N2739, N2734, N256);
and AND4 (N2740, N2733, N2053, N390, N2281);
or OR4 (N2741, N2730, N911, N1887, N1091);
buf BUF1 (N2742, N2739);
buf BUF1 (N2743, N2718);
or OR2 (N2744, N2736, N627);
nor NOR3 (N2745, N2731, N313, N1534);
or OR2 (N2746, N2738, N14);
not NOT1 (N2747, N2742);
and AND3 (N2748, N2740, N1930, N2141);
nand NAND3 (N2749, N2737, N1108, N2154);
nor NOR3 (N2750, N2747, N511, N71);
nand NAND3 (N2751, N2741, N1196, N2135);
nand NAND2 (N2752, N2750, N1187);
nor NOR2 (N2753, N2746, N1330);
and AND4 (N2754, N2745, N110, N2540, N492);
nor NOR4 (N2755, N2732, N1407, N2438, N1339);
not NOT1 (N2756, N2743);
buf BUF1 (N2757, N2729);
nor NOR4 (N2758, N2748, N272, N254, N2050);
xor XOR2 (N2759, N2758, N380);
nor NOR2 (N2760, N2757, N340);
nor NOR2 (N2761, N2759, N79);
and AND2 (N2762, N2751, N196);
xor XOR2 (N2763, N2762, N632);
and AND3 (N2764, N2756, N982, N1105);
or OR4 (N2765, N2754, N915, N222, N1919);
or OR2 (N2766, N2763, N848);
not NOT1 (N2767, N2749);
xor XOR2 (N2768, N2766, N2013);
not NOT1 (N2769, N2768);
not NOT1 (N2770, N2744);
and AND3 (N2771, N2753, N224, N1941);
not NOT1 (N2772, N2767);
nand NAND2 (N2773, N2761, N1521);
nor NOR2 (N2774, N2755, N685);
nor NOR3 (N2775, N2765, N108, N2095);
nand NAND2 (N2776, N2764, N611);
xor XOR2 (N2777, N2774, N1575);
xor XOR2 (N2778, N2775, N1599);
nand NAND2 (N2779, N2752, N1819);
nand NAND3 (N2780, N2769, N297, N2227);
buf BUF1 (N2781, N2770);
and AND2 (N2782, N2760, N2347);
not NOT1 (N2783, N2776);
or OR4 (N2784, N2777, N1690, N2323, N1095);
xor XOR2 (N2785, N2781, N2349);
nand NAND2 (N2786, N2773, N39);
not NOT1 (N2787, N2772);
and AND3 (N2788, N2778, N1294, N1596);
xor XOR2 (N2789, N2785, N2069);
nand NAND3 (N2790, N2779, N2747, N2076);
buf BUF1 (N2791, N2786);
and AND3 (N2792, N2791, N1212, N583);
or OR4 (N2793, N2771, N1011, N2210, N181);
xor XOR2 (N2794, N2792, N960);
xor XOR2 (N2795, N2793, N1569);
nor NOR3 (N2796, N2789, N1986, N1186);
or OR2 (N2797, N2795, N1175);
nor NOR4 (N2798, N2796, N1869, N1094, N1401);
and AND3 (N2799, N2797, N1426, N759);
nand NAND3 (N2800, N2780, N2019, N769);
nand NAND4 (N2801, N2800, N2389, N2620, N268);
buf BUF1 (N2802, N2787);
or OR2 (N2803, N2788, N442);
xor XOR2 (N2804, N2802, N1859);
not NOT1 (N2805, N2794);
buf BUF1 (N2806, N2798);
and AND4 (N2807, N2803, N1463, N1537, N992);
xor XOR2 (N2808, N2782, N1199);
nor NOR2 (N2809, N2801, N1243);
or OR4 (N2810, N2790, N1978, N1890, N2053);
and AND4 (N2811, N2805, N2437, N98, N2495);
and AND3 (N2812, N2806, N2487, N2145);
or OR2 (N2813, N2799, N977);
not NOT1 (N2814, N2804);
buf BUF1 (N2815, N2810);
buf BUF1 (N2816, N2783);
xor XOR2 (N2817, N2812, N652);
or OR2 (N2818, N2817, N1652);
or OR3 (N2819, N2815, N637, N1065);
nand NAND3 (N2820, N2784, N664, N466);
nand NAND2 (N2821, N2819, N2617);
or OR3 (N2822, N2818, N759, N2385);
and AND3 (N2823, N2821, N816, N1228);
not NOT1 (N2824, N2809);
nand NAND3 (N2825, N2808, N1185, N642);
buf BUF1 (N2826, N2807);
and AND2 (N2827, N2820, N614);
buf BUF1 (N2828, N2827);
not NOT1 (N2829, N2811);
nor NOR4 (N2830, N2824, N2424, N1424, N1680);
buf BUF1 (N2831, N2829);
xor XOR2 (N2832, N2831, N732);
and AND3 (N2833, N2830, N478, N92);
not NOT1 (N2834, N2822);
xor XOR2 (N2835, N2828, N1420);
and AND3 (N2836, N2816, N2565, N2298);
not NOT1 (N2837, N2832);
not NOT1 (N2838, N2826);
nor NOR4 (N2839, N2838, N1095, N660, N544);
xor XOR2 (N2840, N2839, N1227);
or OR2 (N2841, N2833, N2485);
not NOT1 (N2842, N2837);
nor NOR3 (N2843, N2836, N1126, N2783);
nor NOR4 (N2844, N2843, N1623, N2715, N2360);
nand NAND4 (N2845, N2813, N2519, N553, N2358);
nor NOR2 (N2846, N2825, N1160);
xor XOR2 (N2847, N2844, N1183);
and AND3 (N2848, N2834, N2579, N1538);
nor NOR2 (N2849, N2814, N310);
not NOT1 (N2850, N2823);
not NOT1 (N2851, N2845);
xor XOR2 (N2852, N2841, N2296);
nor NOR2 (N2853, N2847, N2677);
and AND3 (N2854, N2840, N158, N489);
nor NOR3 (N2855, N2853, N405, N2209);
nor NOR4 (N2856, N2851, N1722, N2853, N2289);
buf BUF1 (N2857, N2856);
buf BUF1 (N2858, N2852);
not NOT1 (N2859, N2849);
nand NAND4 (N2860, N2859, N1321, N2681, N1688);
nor NOR4 (N2861, N2850, N2320, N2833, N57);
nand NAND2 (N2862, N2846, N1840);
xor XOR2 (N2863, N2855, N1911);
buf BUF1 (N2864, N2858);
and AND2 (N2865, N2862, N1301);
or OR3 (N2866, N2864, N1556, N1417);
nand NAND3 (N2867, N2857, N2250, N22);
xor XOR2 (N2868, N2863, N2611);
and AND3 (N2869, N2866, N1951, N686);
buf BUF1 (N2870, N2835);
xor XOR2 (N2871, N2868, N2352);
xor XOR2 (N2872, N2854, N1749);
nor NOR2 (N2873, N2865, N2600);
nor NOR2 (N2874, N2861, N517);
and AND3 (N2875, N2872, N605, N573);
buf BUF1 (N2876, N2867);
or OR2 (N2877, N2875, N906);
nand NAND3 (N2878, N2870, N615, N735);
buf BUF1 (N2879, N2877);
nor NOR4 (N2880, N2842, N2876, N381, N1751);
buf BUF1 (N2881, N469);
nand NAND3 (N2882, N2880, N804, N1054);
xor XOR2 (N2883, N2871, N321);
xor XOR2 (N2884, N2881, N2547);
or OR2 (N2885, N2873, N16);
nor NOR2 (N2886, N2878, N1677);
buf BUF1 (N2887, N2886);
xor XOR2 (N2888, N2848, N2252);
nor NOR4 (N2889, N2860, N216, N2223, N1568);
nor NOR2 (N2890, N2887, N1308);
buf BUF1 (N2891, N2884);
xor XOR2 (N2892, N2888, N1256);
or OR4 (N2893, N2891, N1929, N1506, N817);
nand NAND2 (N2894, N2879, N1159);
and AND3 (N2895, N2893, N2832, N2213);
buf BUF1 (N2896, N2895);
and AND4 (N2897, N2882, N72, N693, N258);
buf BUF1 (N2898, N2894);
or OR3 (N2899, N2898, N2602, N2811);
nor NOR2 (N2900, N2889, N2172);
nand NAND3 (N2901, N2899, N2102, N1175);
nand NAND4 (N2902, N2885, N1280, N1522, N156);
or OR4 (N2903, N2896, N309, N1194, N2329);
nand NAND4 (N2904, N2874, N2027, N1639, N2403);
nand NAND4 (N2905, N2883, N989, N179, N797);
buf BUF1 (N2906, N2902);
buf BUF1 (N2907, N2900);
and AND3 (N2908, N2892, N189, N827);
nor NOR3 (N2909, N2904, N1657, N577);
buf BUF1 (N2910, N2890);
xor XOR2 (N2911, N2908, N2375);
nand NAND2 (N2912, N2909, N1453);
buf BUF1 (N2913, N2905);
nand NAND2 (N2914, N2911, N2729);
buf BUF1 (N2915, N2906);
xor XOR2 (N2916, N2910, N32);
or OR2 (N2917, N2907, N1750);
nor NOR3 (N2918, N2916, N1873, N16);
nor NOR3 (N2919, N2915, N2145, N2492);
and AND4 (N2920, N2917, N1716, N1830, N941);
xor XOR2 (N2921, N2901, N1533);
and AND4 (N2922, N2920, N2205, N1441, N2552);
or OR3 (N2923, N2918, N1472, N1310);
or OR4 (N2924, N2919, N1279, N1884, N918);
nor NOR3 (N2925, N2922, N2833, N1083);
nor NOR4 (N2926, N2925, N2530, N2106, N2);
xor XOR2 (N2927, N2913, N559);
and AND2 (N2928, N2897, N1981);
xor XOR2 (N2929, N2923, N761);
nand NAND4 (N2930, N2914, N478, N1865, N460);
xor XOR2 (N2931, N2929, N2510);
buf BUF1 (N2932, N2924);
xor XOR2 (N2933, N2931, N1861);
buf BUF1 (N2934, N2921);
or OR3 (N2935, N2927, N349, N991);
not NOT1 (N2936, N2934);
and AND3 (N2937, N2869, N1483, N240);
or OR3 (N2938, N2926, N382, N2591);
xor XOR2 (N2939, N2933, N94);
xor XOR2 (N2940, N2939, N2475);
xor XOR2 (N2941, N2930, N695);
and AND3 (N2942, N2903, N2934, N391);
xor XOR2 (N2943, N2932, N890);
not NOT1 (N2944, N2941);
nor NOR2 (N2945, N2943, N1704);
and AND2 (N2946, N2936, N1278);
nand NAND3 (N2947, N2938, N161, N1475);
nand NAND2 (N2948, N2942, N157);
nor NOR4 (N2949, N2947, N2632, N1720, N937);
buf BUF1 (N2950, N2945);
xor XOR2 (N2951, N2935, N252);
or OR3 (N2952, N2940, N2530, N2093);
and AND3 (N2953, N2949, N1370, N673);
xor XOR2 (N2954, N2928, N2648);
xor XOR2 (N2955, N2954, N614);
not NOT1 (N2956, N2951);
nand NAND2 (N2957, N2950, N1547);
xor XOR2 (N2958, N2948, N1134);
or OR3 (N2959, N2946, N669, N1612);
nand NAND3 (N2960, N2953, N1280, N68);
not NOT1 (N2961, N2955);
or OR4 (N2962, N2956, N252, N102, N1640);
nand NAND2 (N2963, N2961, N2572);
or OR2 (N2964, N2952, N2437);
not NOT1 (N2965, N2960);
not NOT1 (N2966, N2944);
xor XOR2 (N2967, N2937, N1570);
xor XOR2 (N2968, N2959, N1834);
xor XOR2 (N2969, N2912, N1787);
nand NAND2 (N2970, N2966, N2081);
nand NAND2 (N2971, N2970, N2123);
buf BUF1 (N2972, N2964);
xor XOR2 (N2973, N2971, N332);
xor XOR2 (N2974, N2969, N577);
not NOT1 (N2975, N2963);
xor XOR2 (N2976, N2975, N2674);
or OR3 (N2977, N2967, N300, N729);
and AND2 (N2978, N2957, N2294);
nor NOR4 (N2979, N2977, N896, N1309, N1185);
xor XOR2 (N2980, N2968, N1666);
and AND2 (N2981, N2980, N2535);
nand NAND3 (N2982, N2962, N1725, N410);
or OR4 (N2983, N2974, N1539, N2931, N2044);
and AND3 (N2984, N2973, N440, N212);
or OR2 (N2985, N2982, N2926);
xor XOR2 (N2986, N2979, N754);
nor NOR3 (N2987, N2981, N1441, N2756);
or OR4 (N2988, N2965, N1574, N13, N522);
buf BUF1 (N2989, N2984);
buf BUF1 (N2990, N2988);
not NOT1 (N2991, N2978);
nor NOR4 (N2992, N2972, N2595, N1603, N2447);
and AND3 (N2993, N2992, N2937, N1682);
and AND2 (N2994, N2985, N2052);
and AND3 (N2995, N2987, N1258, N2195);
not NOT1 (N2996, N2986);
nand NAND3 (N2997, N2995, N433, N2175);
xor XOR2 (N2998, N2991, N1371);
buf BUF1 (N2999, N2997);
nor NOR2 (N3000, N2996, N2589);
nand NAND4 (N3001, N3000, N1004, N616, N850);
and AND4 (N3002, N2998, N1131, N1486, N966);
nor NOR3 (N3003, N2993, N295, N633);
xor XOR2 (N3004, N2990, N2002);
nand NAND4 (N3005, N3004, N1021, N305, N640);
nor NOR3 (N3006, N2976, N2950, N829);
nand NAND3 (N3007, N2999, N1773, N715);
nand NAND2 (N3008, N2983, N13);
nor NOR4 (N3009, N3007, N556, N2666, N747);
not NOT1 (N3010, N2989);
not NOT1 (N3011, N3010);
and AND2 (N3012, N3001, N2314);
not NOT1 (N3013, N3003);
not NOT1 (N3014, N2958);
buf BUF1 (N3015, N3014);
and AND3 (N3016, N3013, N2789, N2825);
nand NAND3 (N3017, N3005, N2005, N1646);
not NOT1 (N3018, N3009);
nand NAND3 (N3019, N3017, N2372, N1503);
buf BUF1 (N3020, N3008);
nand NAND3 (N3021, N2994, N1274, N487);
nand NAND3 (N3022, N3018, N2958, N3008);
xor XOR2 (N3023, N3015, N2143);
and AND2 (N3024, N3002, N2503);
not NOT1 (N3025, N3019);
and AND2 (N3026, N3024, N220);
xor XOR2 (N3027, N3025, N2797);
nor NOR3 (N3028, N3012, N2748, N901);
nor NOR4 (N3029, N3026, N356, N1381, N823);
xor XOR2 (N3030, N3028, N645);
or OR4 (N3031, N3021, N2741, N1926, N2766);
buf BUF1 (N3032, N3023);
nor NOR4 (N3033, N3029, N1222, N577, N1305);
not NOT1 (N3034, N3006);
nand NAND3 (N3035, N3016, N2753, N1286);
not NOT1 (N3036, N3033);
buf BUF1 (N3037, N3032);
nand NAND3 (N3038, N3037, N2826, N2941);
buf BUF1 (N3039, N3011);
buf BUF1 (N3040, N3039);
or OR2 (N3041, N3040, N984);
xor XOR2 (N3042, N3027, N2233);
or OR4 (N3043, N3041, N3032, N1699, N2939);
buf BUF1 (N3044, N3020);
nor NOR3 (N3045, N3043, N1421, N2090);
and AND4 (N3046, N3031, N1733, N1009, N2801);
buf BUF1 (N3047, N3046);
and AND4 (N3048, N3044, N2089, N1477, N1468);
xor XOR2 (N3049, N3042, N886);
nor NOR4 (N3050, N3035, N107, N476, N817);
nor NOR4 (N3051, N3045, N1278, N1197, N1681);
nand NAND2 (N3052, N3034, N27);
not NOT1 (N3053, N3022);
xor XOR2 (N3054, N3038, N3014);
or OR2 (N3055, N3030, N2400);
or OR3 (N3056, N3054, N156, N2174);
xor XOR2 (N3057, N3053, N638);
not NOT1 (N3058, N3050);
xor XOR2 (N3059, N3047, N2455);
buf BUF1 (N3060, N3056);
or OR2 (N3061, N3055, N404);
not NOT1 (N3062, N3036);
nand NAND4 (N3063, N3062, N2598, N1684, N702);
or OR4 (N3064, N3058, N1423, N1753, N958);
and AND4 (N3065, N3057, N2003, N1918, N1735);
nor NOR2 (N3066, N3063, N2962);
and AND2 (N3067, N3061, N1773);
buf BUF1 (N3068, N3060);
nand NAND3 (N3069, N3065, N2599, N1620);
xor XOR2 (N3070, N3059, N2142);
nor NOR2 (N3071, N3051, N1947);
buf BUF1 (N3072, N3067);
buf BUF1 (N3073, N3071);
or OR4 (N3074, N3064, N1306, N472, N2325);
nor NOR4 (N3075, N3052, N1012, N1508, N2985);
nor NOR4 (N3076, N3073, N2755, N952, N573);
not NOT1 (N3077, N3074);
nand NAND4 (N3078, N3077, N467, N2520, N1496);
or OR2 (N3079, N3072, N882);
buf BUF1 (N3080, N3075);
or OR4 (N3081, N3049, N597, N2193, N1067);
nand NAND2 (N3082, N3081, N234);
xor XOR2 (N3083, N3080, N803);
nor NOR4 (N3084, N3066, N1736, N533, N1221);
xor XOR2 (N3085, N3070, N583);
xor XOR2 (N3086, N3048, N544);
xor XOR2 (N3087, N3085, N2230);
xor XOR2 (N3088, N3078, N696);
nor NOR4 (N3089, N3068, N79, N2850, N2259);
nand NAND2 (N3090, N3089, N2607);
xor XOR2 (N3091, N3076, N2695);
or OR3 (N3092, N3069, N2628, N1962);
or OR2 (N3093, N3088, N1982);
buf BUF1 (N3094, N3082);
and AND2 (N3095, N3090, N2965);
buf BUF1 (N3096, N3086);
xor XOR2 (N3097, N3087, N2279);
buf BUF1 (N3098, N3096);
xor XOR2 (N3099, N3091, N1551);
nor NOR3 (N3100, N3084, N1923, N1804);
nor NOR3 (N3101, N3095, N1258, N2219);
nand NAND2 (N3102, N3079, N1133);
buf BUF1 (N3103, N3100);
nor NOR4 (N3104, N3099, N2422, N2562, N2770);
buf BUF1 (N3105, N3101);
and AND3 (N3106, N3098, N515, N102);
nand NAND2 (N3107, N3092, N1189);
not NOT1 (N3108, N3106);
and AND2 (N3109, N3102, N2541);
nand NAND2 (N3110, N3093, N1738);
and AND3 (N3111, N3097, N1278, N2249);
buf BUF1 (N3112, N3083);
xor XOR2 (N3113, N3112, N242);
nand NAND4 (N3114, N3105, N2574, N498, N568);
and AND4 (N3115, N3094, N3025, N552, N107);
or OR2 (N3116, N3114, N61);
not NOT1 (N3117, N3111);
nor NOR2 (N3118, N3107, N1667);
buf BUF1 (N3119, N3117);
not NOT1 (N3120, N3115);
xor XOR2 (N3121, N3120, N2744);
buf BUF1 (N3122, N3109);
nand NAND2 (N3123, N3119, N958);
buf BUF1 (N3124, N3118);
or OR4 (N3125, N3116, N2733, N1554, N3038);
buf BUF1 (N3126, N3113);
nor NOR2 (N3127, N3123, N2907);
nand NAND2 (N3128, N3104, N1946);
xor XOR2 (N3129, N3128, N817);
not NOT1 (N3130, N3129);
or OR2 (N3131, N3125, N2575);
xor XOR2 (N3132, N3103, N738);
nand NAND4 (N3133, N3121, N2984, N475, N2348);
or OR3 (N3134, N3110, N998, N2983);
and AND3 (N3135, N3124, N464, N1794);
buf BUF1 (N3136, N3130);
or OR2 (N3137, N3133, N1618);
not NOT1 (N3138, N3108);
or OR4 (N3139, N3138, N2238, N585, N860);
nand NAND4 (N3140, N3126, N1211, N3032, N1217);
xor XOR2 (N3141, N3132, N2773);
or OR4 (N3142, N3131, N2872, N1393, N1454);
nor NOR3 (N3143, N3134, N1896, N204);
buf BUF1 (N3144, N3136);
nand NAND3 (N3145, N3127, N2767, N1644);
and AND4 (N3146, N3139, N488, N397, N1759);
and AND2 (N3147, N3145, N2732);
nor NOR4 (N3148, N3143, N1653, N1590, N2571);
xor XOR2 (N3149, N3141, N3079);
nand NAND4 (N3150, N3140, N2690, N1289, N1932);
and AND3 (N3151, N3149, N247, N2166);
or OR2 (N3152, N3137, N689);
nand NAND4 (N3153, N3150, N2684, N2525, N1768);
buf BUF1 (N3154, N3147);
xor XOR2 (N3155, N3122, N787);
and AND3 (N3156, N3135, N542, N911);
and AND2 (N3157, N3156, N1474);
or OR4 (N3158, N3153, N1371, N1624, N2026);
or OR3 (N3159, N3155, N2585, N1984);
nor NOR3 (N3160, N3159, N1729, N2373);
or OR3 (N3161, N3154, N2702, N1630);
nand NAND2 (N3162, N3144, N2132);
xor XOR2 (N3163, N3157, N98);
xor XOR2 (N3164, N3161, N1999);
and AND3 (N3165, N3142, N2710, N897);
or OR4 (N3166, N3162, N1915, N1735, N2533);
not NOT1 (N3167, N3166);
or OR3 (N3168, N3164, N2886, N1050);
nand NAND2 (N3169, N3151, N1817);
xor XOR2 (N3170, N3169, N2046);
and AND2 (N3171, N3167, N2880);
not NOT1 (N3172, N3146);
and AND3 (N3173, N3172, N2970, N1168);
xor XOR2 (N3174, N3148, N127);
or OR2 (N3175, N3168, N1616);
buf BUF1 (N3176, N3160);
or OR4 (N3177, N3171, N967, N663, N2848);
or OR3 (N3178, N3152, N633, N2989);
or OR3 (N3179, N3177, N2144, N577);
or OR3 (N3180, N3174, N2926, N1576);
not NOT1 (N3181, N3165);
and AND2 (N3182, N3170, N648);
buf BUF1 (N3183, N3173);
nand NAND3 (N3184, N3181, N2495, N820);
nor NOR2 (N3185, N3178, N2767);
not NOT1 (N3186, N3184);
or OR2 (N3187, N3175, N2094);
buf BUF1 (N3188, N3179);
nor NOR4 (N3189, N3176, N1748, N2667, N2995);
or OR2 (N3190, N3186, N247);
and AND3 (N3191, N3180, N2582, N2385);
nand NAND4 (N3192, N3188, N30, N637, N1199);
and AND2 (N3193, N3187, N1785);
nor NOR3 (N3194, N3183, N1026, N355);
nand NAND4 (N3195, N3194, N159, N2125, N654);
buf BUF1 (N3196, N3158);
buf BUF1 (N3197, N3182);
not NOT1 (N3198, N3190);
nor NOR4 (N3199, N3163, N3165, N1424, N1447);
not NOT1 (N3200, N3199);
nand NAND4 (N3201, N3193, N249, N2471, N2554);
and AND3 (N3202, N3200, N762, N2269);
nor NOR4 (N3203, N3197, N595, N1347, N2827);
not NOT1 (N3204, N3195);
or OR2 (N3205, N3189, N2486);
buf BUF1 (N3206, N3198);
nand NAND3 (N3207, N3191, N824, N2049);
nand NAND3 (N3208, N3196, N2683, N2804);
buf BUF1 (N3209, N3192);
nand NAND2 (N3210, N3205, N2040);
buf BUF1 (N3211, N3201);
not NOT1 (N3212, N3210);
not NOT1 (N3213, N3185);
not NOT1 (N3214, N3208);
not NOT1 (N3215, N3207);
xor XOR2 (N3216, N3212, N1085);
nand NAND4 (N3217, N3213, N2663, N63, N2680);
nand NAND4 (N3218, N3215, N47, N454, N632);
xor XOR2 (N3219, N3206, N2871);
nor NOR2 (N3220, N3209, N483);
buf BUF1 (N3221, N3220);
xor XOR2 (N3222, N3204, N2760);
and AND2 (N3223, N3202, N1644);
nor NOR3 (N3224, N3219, N166, N2001);
not NOT1 (N3225, N3224);
buf BUF1 (N3226, N3216);
and AND2 (N3227, N3221, N1955);
nand NAND3 (N3228, N3222, N2185, N3025);
nor NOR4 (N3229, N3211, N1753, N2713, N1313);
not NOT1 (N3230, N3203);
and AND4 (N3231, N3225, N1877, N1155, N3203);
or OR3 (N3232, N3217, N2290, N2954);
or OR3 (N3233, N3230, N1419, N839);
nor NOR3 (N3234, N3226, N2856, N1900);
buf BUF1 (N3235, N3218);
buf BUF1 (N3236, N3235);
buf BUF1 (N3237, N3234);
xor XOR2 (N3238, N3229, N606);
xor XOR2 (N3239, N3237, N2142);
buf BUF1 (N3240, N3233);
and AND3 (N3241, N3231, N2981, N1354);
xor XOR2 (N3242, N3236, N3063);
nor NOR3 (N3243, N3238, N2334, N98);
not NOT1 (N3244, N3227);
not NOT1 (N3245, N3242);
xor XOR2 (N3246, N3214, N1974);
nor NOR4 (N3247, N3239, N3149, N2580, N1250);
buf BUF1 (N3248, N3246);
buf BUF1 (N3249, N3247);
and AND2 (N3250, N3249, N196);
or OR2 (N3251, N3245, N1931);
not NOT1 (N3252, N3248);
and AND4 (N3253, N3241, N2991, N2660, N2042);
xor XOR2 (N3254, N3250, N2034);
not NOT1 (N3255, N3232);
not NOT1 (N3256, N3240);
xor XOR2 (N3257, N3243, N3196);
not NOT1 (N3258, N3254);
not NOT1 (N3259, N3223);
buf BUF1 (N3260, N3252);
buf BUF1 (N3261, N3259);
and AND2 (N3262, N3256, N1066);
or OR4 (N3263, N3260, N1690, N1100, N1031);
or OR2 (N3264, N3244, N2036);
buf BUF1 (N3265, N3253);
nor NOR3 (N3266, N3261, N1168, N952);
and AND3 (N3267, N3265, N568, N1712);
or OR2 (N3268, N3267, N2509);
buf BUF1 (N3269, N3262);
nand NAND2 (N3270, N3255, N2141);
buf BUF1 (N3271, N3263);
nand NAND3 (N3272, N3270, N2030, N2284);
or OR4 (N3273, N3272, N324, N182, N722);
xor XOR2 (N3274, N3266, N1093);
nand NAND3 (N3275, N3228, N88, N1649);
nor NOR2 (N3276, N3251, N1509);
buf BUF1 (N3277, N3273);
nand NAND2 (N3278, N3276, N2402);
buf BUF1 (N3279, N3275);
or OR2 (N3280, N3277, N1631);
buf BUF1 (N3281, N3280);
and AND4 (N3282, N3274, N426, N1769, N1074);
nor NOR3 (N3283, N3281, N692, N1500);
xor XOR2 (N3284, N3258, N2561);
xor XOR2 (N3285, N3283, N3072);
and AND4 (N3286, N3284, N2152, N2257, N694);
and AND3 (N3287, N3269, N509, N2932);
not NOT1 (N3288, N3271);
nor NOR4 (N3289, N3268, N775, N775, N2165);
or OR3 (N3290, N3282, N3077, N827);
not NOT1 (N3291, N3290);
not NOT1 (N3292, N3287);
xor XOR2 (N3293, N3289, N465);
nor NOR4 (N3294, N3286, N3048, N47, N2550);
nor NOR3 (N3295, N3294, N845, N710);
nand NAND3 (N3296, N3257, N579, N3226);
xor XOR2 (N3297, N3292, N2533);
not NOT1 (N3298, N3297);
buf BUF1 (N3299, N3295);
and AND4 (N3300, N3296, N1388, N418, N2221);
nor NOR2 (N3301, N3288, N241);
xor XOR2 (N3302, N3300, N2962);
and AND2 (N3303, N3299, N1794);
nor NOR2 (N3304, N3293, N1993);
xor XOR2 (N3305, N3301, N2227);
or OR3 (N3306, N3264, N3284, N2521);
not NOT1 (N3307, N3305);
buf BUF1 (N3308, N3279);
nand NAND4 (N3309, N3308, N774, N716, N2831);
and AND3 (N3310, N3307, N1770, N3032);
buf BUF1 (N3311, N3309);
nor NOR4 (N3312, N3303, N409, N47, N877);
or OR4 (N3313, N3312, N1013, N829, N2325);
or OR2 (N3314, N3291, N144);
xor XOR2 (N3315, N3278, N1770);
xor XOR2 (N3316, N3311, N886);
or OR3 (N3317, N3313, N2227, N492);
buf BUF1 (N3318, N3306);
and AND3 (N3319, N3310, N291, N2754);
nand NAND4 (N3320, N3298, N996, N2549, N2049);
or OR4 (N3321, N3315, N2187, N2478, N1398);
or OR4 (N3322, N3320, N2957, N2668, N2083);
nor NOR3 (N3323, N3304, N993, N673);
or OR4 (N3324, N3317, N1652, N2849, N3014);
xor XOR2 (N3325, N3314, N3180);
and AND2 (N3326, N3285, N899);
nor NOR2 (N3327, N3321, N2080);
and AND3 (N3328, N3324, N3059, N973);
not NOT1 (N3329, N3325);
and AND3 (N3330, N3322, N560, N3208);
and AND3 (N3331, N3319, N1412, N795);
nand NAND4 (N3332, N3326, N705, N2991, N1510);
not NOT1 (N3333, N3332);
or OR2 (N3334, N3323, N3331);
nand NAND2 (N3335, N1239, N778);
or OR4 (N3336, N3328, N2420, N472, N104);
nor NOR4 (N3337, N3333, N2603, N2139, N1921);
not NOT1 (N3338, N3335);
buf BUF1 (N3339, N3316);
and AND4 (N3340, N3302, N912, N715, N918);
or OR3 (N3341, N3318, N108, N2991);
not NOT1 (N3342, N3330);
xor XOR2 (N3343, N3342, N2761);
nand NAND4 (N3344, N3329, N831, N1233, N2665);
or OR2 (N3345, N3334, N2144);
buf BUF1 (N3346, N3345);
buf BUF1 (N3347, N3343);
xor XOR2 (N3348, N3339, N2775);
buf BUF1 (N3349, N3338);
xor XOR2 (N3350, N3336, N2200);
xor XOR2 (N3351, N3344, N3134);
not NOT1 (N3352, N3327);
not NOT1 (N3353, N3340);
not NOT1 (N3354, N3348);
and AND4 (N3355, N3354, N1748, N308, N3331);
xor XOR2 (N3356, N3346, N1894);
nand NAND3 (N3357, N3349, N3150, N2072);
xor XOR2 (N3358, N3347, N1836);
nor NOR3 (N3359, N3352, N530, N2030);
and AND3 (N3360, N3337, N824, N1288);
buf BUF1 (N3361, N3341);
buf BUF1 (N3362, N3350);
xor XOR2 (N3363, N3355, N1969);
buf BUF1 (N3364, N3353);
nor NOR3 (N3365, N3363, N2492, N2972);
not NOT1 (N3366, N3360);
xor XOR2 (N3367, N3359, N2963);
and AND3 (N3368, N3366, N1615, N2230);
or OR2 (N3369, N3357, N2457);
nand NAND4 (N3370, N3362, N2413, N2690, N2893);
or OR3 (N3371, N3365, N1435, N1623);
nor NOR4 (N3372, N3358, N1336, N3000, N522);
not NOT1 (N3373, N3356);
and AND3 (N3374, N3369, N2309, N434);
xor XOR2 (N3375, N3370, N448);
xor XOR2 (N3376, N3364, N89);
or OR4 (N3377, N3371, N464, N666, N451);
buf BUF1 (N3378, N3361);
nor NOR4 (N3379, N3375, N2050, N443, N433);
not NOT1 (N3380, N3368);
not NOT1 (N3381, N3374);
xor XOR2 (N3382, N3381, N2533);
buf BUF1 (N3383, N3378);
nand NAND4 (N3384, N3367, N2782, N2510, N1314);
nor NOR4 (N3385, N3382, N592, N1776, N1278);
not NOT1 (N3386, N3372);
or OR4 (N3387, N3373, N1388, N822, N2892);
or OR4 (N3388, N3377, N2755, N2245, N415);
and AND4 (N3389, N3379, N1928, N557, N1858);
and AND2 (N3390, N3384, N755);
xor XOR2 (N3391, N3376, N3231);
not NOT1 (N3392, N3389);
nand NAND3 (N3393, N3386, N39, N1079);
not NOT1 (N3394, N3383);
and AND3 (N3395, N3393, N2912, N3375);
nor NOR4 (N3396, N3388, N2363, N635, N1555);
and AND2 (N3397, N3391, N427);
or OR3 (N3398, N3390, N1196, N395);
nand NAND3 (N3399, N3387, N1726, N1450);
nand NAND4 (N3400, N3351, N2936, N240, N2214);
nor NOR3 (N3401, N3398, N83, N1089);
not NOT1 (N3402, N3395);
xor XOR2 (N3403, N3397, N1074);
xor XOR2 (N3404, N3396, N196);
not NOT1 (N3405, N3380);
and AND3 (N3406, N3385, N1714, N2592);
not NOT1 (N3407, N3405);
buf BUF1 (N3408, N3399);
nand NAND2 (N3409, N3407, N1667);
nand NAND4 (N3410, N3401, N1181, N1172, N1443);
nor NOR4 (N3411, N3408, N1981, N1240, N2330);
buf BUF1 (N3412, N3411);
nand NAND2 (N3413, N3394, N348);
and AND3 (N3414, N3406, N1363, N1670);
nand NAND2 (N3415, N3409, N3073);
not NOT1 (N3416, N3404);
nand NAND4 (N3417, N3412, N2497, N1174, N3208);
xor XOR2 (N3418, N3400, N217);
nand NAND4 (N3419, N3415, N3050, N2512, N2157);
buf BUF1 (N3420, N3410);
not NOT1 (N3421, N3413);
and AND2 (N3422, N3414, N2472);
not NOT1 (N3423, N3403);
xor XOR2 (N3424, N3402, N3232);
or OR3 (N3425, N3417, N43, N1384);
and AND2 (N3426, N3421, N160);
buf BUF1 (N3427, N3425);
or OR3 (N3428, N3424, N2273, N2977);
not NOT1 (N3429, N3418);
and AND4 (N3430, N3392, N868, N2619, N1184);
buf BUF1 (N3431, N3416);
nor NOR4 (N3432, N3426, N151, N2359, N808);
xor XOR2 (N3433, N3430, N2232);
and AND4 (N3434, N3429, N1595, N852, N1465);
or OR4 (N3435, N3433, N1035, N560, N1414);
or OR3 (N3436, N3428, N2033, N1348);
not NOT1 (N3437, N3422);
or OR2 (N3438, N3431, N2236);
and AND3 (N3439, N3434, N990, N1906);
and AND3 (N3440, N3435, N1442, N836);
buf BUF1 (N3441, N3420);
or OR4 (N3442, N3440, N422, N560, N2122);
buf BUF1 (N3443, N3432);
xor XOR2 (N3444, N3442, N1147);
not NOT1 (N3445, N3439);
not NOT1 (N3446, N3445);
nand NAND2 (N3447, N3444, N1297);
and AND2 (N3448, N3441, N2987);
nor NOR4 (N3449, N3447, N1947, N732, N2855);
not NOT1 (N3450, N3438);
and AND3 (N3451, N3443, N2635, N1949);
not NOT1 (N3452, N3448);
and AND3 (N3453, N3451, N2525, N1849);
xor XOR2 (N3454, N3419, N1701);
or OR2 (N3455, N3436, N1994);
not NOT1 (N3456, N3446);
or OR3 (N3457, N3437, N1562, N837);
buf BUF1 (N3458, N3453);
nor NOR3 (N3459, N3454, N1033, N1276);
nor NOR2 (N3460, N3452, N767);
buf BUF1 (N3461, N3456);
not NOT1 (N3462, N3459);
and AND3 (N3463, N3450, N2934, N2641);
nand NAND2 (N3464, N3461, N3046);
not NOT1 (N3465, N3460);
and AND2 (N3466, N3465, N3370);
nand NAND4 (N3467, N3463, N532, N1976, N1429);
or OR4 (N3468, N3464, N19, N2430, N1299);
not NOT1 (N3469, N3458);
xor XOR2 (N3470, N3423, N2358);
and AND4 (N3471, N3449, N1969, N743, N644);
not NOT1 (N3472, N3471);
nand NAND2 (N3473, N3467, N2091);
not NOT1 (N3474, N3427);
nor NOR2 (N3475, N3462, N3167);
or OR2 (N3476, N3475, N2869);
not NOT1 (N3477, N3469);
xor XOR2 (N3478, N3466, N2441);
nor NOR4 (N3479, N3474, N1780, N1456, N1001);
or OR3 (N3480, N3468, N707, N246);
nor NOR3 (N3481, N3473, N1881, N2392);
and AND4 (N3482, N3472, N3042, N3271, N57);
nor NOR2 (N3483, N3480, N1382);
not NOT1 (N3484, N3482);
nor NOR2 (N3485, N3477, N3458);
nor NOR4 (N3486, N3457, N553, N1951, N3249);
nand NAND2 (N3487, N3478, N1151);
and AND4 (N3488, N3470, N2056, N1172, N2540);
nand NAND3 (N3489, N3484, N1611, N3156);
not NOT1 (N3490, N3476);
nand NAND3 (N3491, N3481, N616, N228);
xor XOR2 (N3492, N3488, N2207);
nand NAND2 (N3493, N3485, N198);
buf BUF1 (N3494, N3487);
buf BUF1 (N3495, N3486);
not NOT1 (N3496, N3492);
nor NOR4 (N3497, N3493, N1635, N3375, N800);
or OR4 (N3498, N3490, N3346, N643, N2977);
not NOT1 (N3499, N3491);
and AND4 (N3500, N3479, N1588, N1801, N2481);
not NOT1 (N3501, N3489);
and AND2 (N3502, N3501, N3015);
and AND4 (N3503, N3500, N1858, N380, N1513);
not NOT1 (N3504, N3455);
nand NAND3 (N3505, N3495, N443, N1524);
not NOT1 (N3506, N3499);
nor NOR2 (N3507, N3502, N925);
or OR2 (N3508, N3483, N1720);
buf BUF1 (N3509, N3505);
nor NOR3 (N3510, N3497, N3429, N2079);
or OR3 (N3511, N3498, N334, N3375);
xor XOR2 (N3512, N3510, N3211);
nand NAND2 (N3513, N3494, N2640);
and AND3 (N3514, N3503, N1648, N202);
nand NAND3 (N3515, N3496, N113, N2622);
buf BUF1 (N3516, N3506);
and AND3 (N3517, N3514, N3136, N3111);
nor NOR4 (N3518, N3507, N1478, N2868, N2846);
or OR3 (N3519, N3515, N503, N1950);
nor NOR4 (N3520, N3517, N1781, N555, N1561);
and AND4 (N3521, N3509, N3188, N664, N890);
or OR2 (N3522, N3513, N2854);
nor NOR2 (N3523, N3518, N102);
and AND3 (N3524, N3516, N2762, N832);
and AND2 (N3525, N3511, N120);
not NOT1 (N3526, N3508);
nor NOR3 (N3527, N3523, N1521, N3311);
nor NOR2 (N3528, N3520, N522);
nand NAND4 (N3529, N3522, N330, N909, N2975);
and AND4 (N3530, N3519, N3526, N1258, N2260);
or OR2 (N3531, N740, N373);
buf BUF1 (N3532, N3504);
xor XOR2 (N3533, N3524, N3318);
nor NOR2 (N3534, N3528, N432);
buf BUF1 (N3535, N3533);
or OR3 (N3536, N3512, N618, N2668);
or OR3 (N3537, N3531, N397, N911);
and AND2 (N3538, N3535, N212);
nor NOR2 (N3539, N3538, N252);
not NOT1 (N3540, N3527);
or OR2 (N3541, N3534, N1352);
nor NOR2 (N3542, N3532, N971);
xor XOR2 (N3543, N3525, N1395);
xor XOR2 (N3544, N3540, N1729);
and AND3 (N3545, N3542, N1224, N1966);
xor XOR2 (N3546, N3543, N615);
or OR4 (N3547, N3539, N2000, N1072, N547);
and AND4 (N3548, N3529, N53, N1874, N2580);
nand NAND3 (N3549, N3530, N1136, N2808);
buf BUF1 (N3550, N3541);
xor XOR2 (N3551, N3550, N1192);
nor NOR2 (N3552, N3549, N1649);
nor NOR2 (N3553, N3551, N240);
nor NOR4 (N3554, N3537, N707, N3186, N2679);
or OR4 (N3555, N3536, N1514, N47, N2160);
and AND4 (N3556, N3548, N1721, N877, N3211);
buf BUF1 (N3557, N3553);
and AND3 (N3558, N3555, N2133, N301);
and AND2 (N3559, N3544, N2174);
xor XOR2 (N3560, N3559, N1230);
and AND3 (N3561, N3545, N3442, N829);
nand NAND2 (N3562, N3521, N3302);
xor XOR2 (N3563, N3552, N544);
xor XOR2 (N3564, N3560, N519);
buf BUF1 (N3565, N3564);
buf BUF1 (N3566, N3565);
nand NAND3 (N3567, N3557, N2740, N3054);
not NOT1 (N3568, N3566);
not NOT1 (N3569, N3568);
nor NOR3 (N3570, N3569, N3235, N1494);
and AND2 (N3571, N3567, N54);
not NOT1 (N3572, N3561);
and AND3 (N3573, N3558, N1319, N2722);
or OR3 (N3574, N3570, N2050, N866);
buf BUF1 (N3575, N3554);
or OR4 (N3576, N3575, N3405, N954, N2087);
or OR2 (N3577, N3571, N3077);
buf BUF1 (N3578, N3563);
xor XOR2 (N3579, N3572, N1630);
or OR2 (N3580, N3576, N1902);
buf BUF1 (N3581, N3577);
not NOT1 (N3582, N3580);
not NOT1 (N3583, N3578);
nand NAND3 (N3584, N3573, N3181, N2206);
xor XOR2 (N3585, N3574, N1657);
xor XOR2 (N3586, N3583, N876);
not NOT1 (N3587, N3586);
buf BUF1 (N3588, N3585);
not NOT1 (N3589, N3562);
nand NAND4 (N3590, N3582, N499, N1576, N1505);
nand NAND4 (N3591, N3546, N2316, N2621, N2486);
and AND2 (N3592, N3588, N552);
or OR2 (N3593, N3584, N2649);
or OR4 (N3594, N3589, N1480, N3212, N3128);
or OR3 (N3595, N3581, N2004, N1826);
xor XOR2 (N3596, N3594, N977);
buf BUF1 (N3597, N3587);
or OR4 (N3598, N3556, N2718, N387, N255);
nor NOR4 (N3599, N3590, N2074, N1933, N3381);
not NOT1 (N3600, N3591);
nand NAND2 (N3601, N3547, N3584);
xor XOR2 (N3602, N3593, N3201);
xor XOR2 (N3603, N3595, N827);
buf BUF1 (N3604, N3600);
xor XOR2 (N3605, N3604, N3018);
nand NAND2 (N3606, N3599, N444);
and AND3 (N3607, N3597, N3589, N631);
xor XOR2 (N3608, N3592, N3452);
nand NAND4 (N3609, N3602, N3, N1942, N1112);
buf BUF1 (N3610, N3609);
buf BUF1 (N3611, N3605);
or OR2 (N3612, N3611, N2263);
not NOT1 (N3613, N3579);
buf BUF1 (N3614, N3601);
nor NOR2 (N3615, N3596, N2962);
xor XOR2 (N3616, N3615, N1803);
xor XOR2 (N3617, N3607, N1056);
nor NOR3 (N3618, N3608, N2439, N671);
not NOT1 (N3619, N3616);
xor XOR2 (N3620, N3598, N929);
or OR2 (N3621, N3619, N278);
nor NOR4 (N3622, N3603, N2913, N2103, N1247);
or OR2 (N3623, N3612, N1936);
or OR3 (N3624, N3613, N2686, N150);
or OR2 (N3625, N3606, N3361);
nand NAND4 (N3626, N3614, N2080, N3069, N2804);
nor NOR3 (N3627, N3620, N1721, N71);
buf BUF1 (N3628, N3627);
nand NAND4 (N3629, N3625, N439, N461, N1522);
nand NAND2 (N3630, N3623, N3154);
and AND3 (N3631, N3618, N1511, N1120);
xor XOR2 (N3632, N3624, N2471);
nand NAND2 (N3633, N3632, N1365);
and AND2 (N3634, N3622, N3312);
xor XOR2 (N3635, N3629, N2641);
nor NOR4 (N3636, N3626, N1276, N1261, N541);
or OR2 (N3637, N3631, N2852);
buf BUF1 (N3638, N3633);
nor NOR4 (N3639, N3610, N2969, N212, N1884);
buf BUF1 (N3640, N3637);
or OR3 (N3641, N3639, N1532, N1617);
not NOT1 (N3642, N3636);
buf BUF1 (N3643, N3634);
nor NOR3 (N3644, N3630, N675, N1057);
and AND2 (N3645, N3628, N866);
and AND2 (N3646, N3617, N383);
xor XOR2 (N3647, N3642, N2159);
and AND3 (N3648, N3635, N606, N2904);
nor NOR2 (N3649, N3640, N3357);
nand NAND2 (N3650, N3645, N3200);
and AND2 (N3651, N3650, N210);
nor NOR4 (N3652, N3638, N651, N2308, N3427);
and AND4 (N3653, N3621, N2654, N2914, N1835);
or OR3 (N3654, N3652, N1910, N3248);
nand NAND3 (N3655, N3643, N1029, N1382);
xor XOR2 (N3656, N3651, N3493);
nor NOR4 (N3657, N3654, N3175, N3116, N322);
nand NAND4 (N3658, N3653, N751, N7, N227);
nand NAND2 (N3659, N3646, N2014);
nand NAND3 (N3660, N3644, N1163, N158);
or OR3 (N3661, N3660, N1648, N3320);
nand NAND2 (N3662, N3648, N11);
nand NAND4 (N3663, N3658, N1953, N1256, N1369);
not NOT1 (N3664, N3641);
not NOT1 (N3665, N3655);
and AND4 (N3666, N3647, N1084, N2132, N1617);
or OR3 (N3667, N3661, N2350, N3347);
xor XOR2 (N3668, N3662, N2760);
nand NAND4 (N3669, N3649, N3274, N1490, N1537);
or OR4 (N3670, N3665, N1777, N2972, N1436);
nor NOR2 (N3671, N3666, N947);
xor XOR2 (N3672, N3657, N3622);
xor XOR2 (N3673, N3668, N2644);
or OR4 (N3674, N3656, N2694, N1547, N2412);
not NOT1 (N3675, N3663);
nand NAND2 (N3676, N3673, N2206);
buf BUF1 (N3677, N3672);
not NOT1 (N3678, N3670);
buf BUF1 (N3679, N3671);
nor NOR3 (N3680, N3667, N1148, N480);
and AND4 (N3681, N3674, N154, N3021, N3645);
not NOT1 (N3682, N3678);
nand NAND3 (N3683, N3679, N1216, N803);
xor XOR2 (N3684, N3659, N446);
buf BUF1 (N3685, N3677);
nand NAND2 (N3686, N3681, N1657);
xor XOR2 (N3687, N3680, N3154);
nor NOR4 (N3688, N3664, N3145, N2773, N3167);
nor NOR4 (N3689, N3675, N2139, N3632, N788);
not NOT1 (N3690, N3686);
buf BUF1 (N3691, N3683);
not NOT1 (N3692, N3684);
nor NOR4 (N3693, N3688, N3555, N1868, N2645);
xor XOR2 (N3694, N3682, N666);
and AND2 (N3695, N3676, N2278);
buf BUF1 (N3696, N3669);
and AND4 (N3697, N3690, N297, N2559, N723);
nand NAND3 (N3698, N3697, N2823, N1971);
buf BUF1 (N3699, N3687);
not NOT1 (N3700, N3685);
xor XOR2 (N3701, N3693, N1265);
xor XOR2 (N3702, N3700, N1941);
xor XOR2 (N3703, N3702, N2810);
or OR3 (N3704, N3698, N1187, N1257);
and AND3 (N3705, N3689, N3169, N705);
and AND4 (N3706, N3692, N1385, N3625, N3288);
not NOT1 (N3707, N3696);
nand NAND4 (N3708, N3704, N1796, N1638, N3220);
not NOT1 (N3709, N3706);
nor NOR4 (N3710, N3694, N692, N3614, N60);
or OR3 (N3711, N3703, N1912, N3130);
or OR2 (N3712, N3709, N1992);
or OR4 (N3713, N3711, N2754, N3337, N3559);
and AND3 (N3714, N3707, N1990, N267);
not NOT1 (N3715, N3699);
or OR3 (N3716, N3691, N45, N586);
buf BUF1 (N3717, N3705);
or OR4 (N3718, N3715, N1064, N423, N1488);
nor NOR3 (N3719, N3712, N1589, N1152);
xor XOR2 (N3720, N3716, N442);
nor NOR2 (N3721, N3710, N2533);
or OR3 (N3722, N3720, N2282, N61);
and AND3 (N3723, N3721, N1124, N541);
not NOT1 (N3724, N3695);
buf BUF1 (N3725, N3719);
buf BUF1 (N3726, N3701);
not NOT1 (N3727, N3726);
or OR4 (N3728, N3727, N2213, N206, N975);
nor NOR2 (N3729, N3722, N3713);
or OR3 (N3730, N1176, N3218, N973);
not NOT1 (N3731, N3729);
and AND4 (N3732, N3730, N1365, N2042, N944);
nor NOR3 (N3733, N3725, N3256, N3405);
xor XOR2 (N3734, N3728, N3510);
xor XOR2 (N3735, N3731, N683);
nand NAND4 (N3736, N3735, N3274, N1265, N3494);
and AND2 (N3737, N3734, N1112);
and AND2 (N3738, N3733, N691);
nand NAND2 (N3739, N3732, N3188);
buf BUF1 (N3740, N3736);
or OR3 (N3741, N3724, N965, N1553);
buf BUF1 (N3742, N3714);
xor XOR2 (N3743, N3738, N1256);
buf BUF1 (N3744, N3723);
nor NOR4 (N3745, N3741, N3621, N3362, N1869);
and AND3 (N3746, N3744, N2285, N908);
xor XOR2 (N3747, N3708, N1906);
nand NAND2 (N3748, N3747, N308);
and AND2 (N3749, N3737, N1386);
or OR2 (N3750, N3743, N1503);
not NOT1 (N3751, N3746);
not NOT1 (N3752, N3718);
not NOT1 (N3753, N3739);
nand NAND2 (N3754, N3740, N3712);
not NOT1 (N3755, N3717);
and AND4 (N3756, N3755, N1122, N3081, N2085);
xor XOR2 (N3757, N3745, N3522);
not NOT1 (N3758, N3751);
and AND4 (N3759, N3750, N3300, N1403, N874);
xor XOR2 (N3760, N3757, N1623);
xor XOR2 (N3761, N3753, N938);
nor NOR3 (N3762, N3749, N2422, N2110);
buf BUF1 (N3763, N3758);
buf BUF1 (N3764, N3760);
not NOT1 (N3765, N3756);
not NOT1 (N3766, N3754);
xor XOR2 (N3767, N3762, N2676);
or OR2 (N3768, N3763, N1190);
and AND2 (N3769, N3765, N3180);
or OR3 (N3770, N3742, N142, N2902);
and AND4 (N3771, N3766, N1225, N1973, N3113);
and AND2 (N3772, N3759, N3716);
xor XOR2 (N3773, N3752, N925);
nor NOR3 (N3774, N3771, N3050, N173);
and AND4 (N3775, N3770, N747, N1596, N1758);
or OR4 (N3776, N3768, N3285, N3696, N3477);
not NOT1 (N3777, N3764);
and AND3 (N3778, N3775, N1303, N1816);
and AND2 (N3779, N3773, N1751);
nand NAND4 (N3780, N3777, N952, N3353, N1957);
xor XOR2 (N3781, N3780, N3096);
nor NOR3 (N3782, N3772, N2499, N177);
nor NOR4 (N3783, N3781, N2036, N115, N2675);
not NOT1 (N3784, N3783);
and AND2 (N3785, N3767, N446);
nand NAND2 (N3786, N3761, N127);
nor NOR2 (N3787, N3785, N308);
nand NAND4 (N3788, N3779, N3025, N2899, N1196);
nand NAND3 (N3789, N3776, N2698, N2810);
buf BUF1 (N3790, N3787);
nor NOR2 (N3791, N3786, N2688);
nor NOR4 (N3792, N3788, N1661, N2954, N3669);
xor XOR2 (N3793, N3778, N2873);
or OR4 (N3794, N3774, N3574, N2763, N2563);
nand NAND4 (N3795, N3782, N909, N3328, N2507);
nand NAND3 (N3796, N3748, N169, N2416);
not NOT1 (N3797, N3789);
xor XOR2 (N3798, N3794, N302);
xor XOR2 (N3799, N3769, N3796);
or OR3 (N3800, N1399, N2533, N3468);
nor NOR2 (N3801, N3798, N5);
nand NAND2 (N3802, N3792, N3566);
or OR3 (N3803, N3791, N2323, N938);
xor XOR2 (N3804, N3800, N2028);
nor NOR4 (N3805, N3797, N899, N2013, N1963);
xor XOR2 (N3806, N3799, N2858);
nand NAND3 (N3807, N3803, N2130, N1224);
buf BUF1 (N3808, N3807);
not NOT1 (N3809, N3784);
nor NOR2 (N3810, N3802, N2808);
and AND3 (N3811, N3804, N39, N1040);
buf BUF1 (N3812, N3806);
not NOT1 (N3813, N3795);
buf BUF1 (N3814, N3810);
nor NOR4 (N3815, N3793, N3781, N3585, N1643);
buf BUF1 (N3816, N3801);
not NOT1 (N3817, N3812);
nor NOR2 (N3818, N3817, N414);
buf BUF1 (N3819, N3814);
and AND2 (N3820, N3805, N2823);
nand NAND2 (N3821, N3790, N3538);
nor NOR4 (N3822, N3820, N3190, N2299, N1445);
nand NAND4 (N3823, N3819, N1043, N1615, N1931);
xor XOR2 (N3824, N3816, N679);
or OR4 (N3825, N3811, N3327, N2008, N264);
or OR4 (N3826, N3808, N1946, N2740, N2246);
and AND3 (N3827, N3823, N262, N3043);
and AND3 (N3828, N3824, N1588, N1166);
nand NAND3 (N3829, N3825, N3052, N2970);
not NOT1 (N3830, N3827);
or OR4 (N3831, N3809, N343, N892, N1070);
buf BUF1 (N3832, N3818);
nor NOR2 (N3833, N3813, N3294);
buf BUF1 (N3834, N3833);
buf BUF1 (N3835, N3822);
nor NOR3 (N3836, N3831, N211, N2021);
nand NAND4 (N3837, N3830, N1990, N1606, N390);
nor NOR2 (N3838, N3832, N1865);
buf BUF1 (N3839, N3837);
xor XOR2 (N3840, N3839, N3074);
and AND4 (N3841, N3835, N2439, N2660, N2786);
not NOT1 (N3842, N3829);
and AND2 (N3843, N3842, N78);
buf BUF1 (N3844, N3834);
xor XOR2 (N3845, N3828, N1188);
and AND3 (N3846, N3821, N1214, N3747);
and AND2 (N3847, N3844, N3353);
not NOT1 (N3848, N3838);
buf BUF1 (N3849, N3841);
nand NAND3 (N3850, N3826, N595, N1201);
xor XOR2 (N3851, N3850, N3418);
nand NAND4 (N3852, N3845, N2925, N1453, N1367);
or OR2 (N3853, N3846, N2891);
nor NOR2 (N3854, N3849, N2271);
nor NOR2 (N3855, N3847, N380);
xor XOR2 (N3856, N3854, N2020);
xor XOR2 (N3857, N3843, N912);
or OR3 (N3858, N3851, N1517, N3232);
buf BUF1 (N3859, N3857);
and AND4 (N3860, N3853, N226, N2423, N163);
and AND2 (N3861, N3855, N2860);
or OR2 (N3862, N3861, N1346);
nor NOR3 (N3863, N3862, N3128, N1761);
nor NOR4 (N3864, N3848, N1269, N157, N2815);
not NOT1 (N3865, N3863);
nor NOR3 (N3866, N3840, N3129, N1009);
xor XOR2 (N3867, N3860, N933);
or OR3 (N3868, N3858, N25, N3654);
xor XOR2 (N3869, N3867, N2386);
buf BUF1 (N3870, N3836);
buf BUF1 (N3871, N3865);
not NOT1 (N3872, N3856);
not NOT1 (N3873, N3870);
nand NAND3 (N3874, N3859, N2869, N3583);
nor NOR3 (N3875, N3871, N3176, N2996);
nor NOR2 (N3876, N3872, N414);
nand NAND2 (N3877, N3868, N1592);
not NOT1 (N3878, N3875);
not NOT1 (N3879, N3873);
buf BUF1 (N3880, N3864);
nand NAND3 (N3881, N3879, N2668, N3678);
buf BUF1 (N3882, N3866);
xor XOR2 (N3883, N3869, N398);
not NOT1 (N3884, N3877);
and AND2 (N3885, N3884, N1152);
nor NOR4 (N3886, N3878, N1219, N1831, N2252);
not NOT1 (N3887, N3874);
xor XOR2 (N3888, N3881, N557);
nor NOR3 (N3889, N3883, N1528, N729);
xor XOR2 (N3890, N3880, N464);
not NOT1 (N3891, N3885);
nor NOR3 (N3892, N3876, N2069, N1104);
or OR2 (N3893, N3886, N473);
nor NOR4 (N3894, N3890, N2355, N3031, N164);
buf BUF1 (N3895, N3892);
not NOT1 (N3896, N3893);
not NOT1 (N3897, N3889);
not NOT1 (N3898, N3897);
not NOT1 (N3899, N3898);
not NOT1 (N3900, N3852);
and AND2 (N3901, N3891, N49);
and AND3 (N3902, N3901, N1363, N2445);
xor XOR2 (N3903, N3900, N3610);
nor NOR3 (N3904, N3899, N2396, N1020);
or OR4 (N3905, N3894, N1203, N85, N1967);
and AND4 (N3906, N3896, N2005, N1720, N2686);
buf BUF1 (N3907, N3905);
xor XOR2 (N3908, N3887, N823);
xor XOR2 (N3909, N3815, N2003);
nand NAND4 (N3910, N3895, N3830, N1730, N1597);
xor XOR2 (N3911, N3902, N3491);
xor XOR2 (N3912, N3903, N1043);
nor NOR2 (N3913, N3912, N2012);
and AND4 (N3914, N3907, N1084, N2670, N3700);
and AND2 (N3915, N3910, N1141);
or OR2 (N3916, N3914, N3506);
nand NAND2 (N3917, N3888, N3444);
nor NOR2 (N3918, N3882, N3898);
nand NAND4 (N3919, N3908, N1690, N310, N3425);
not NOT1 (N3920, N3917);
nor NOR4 (N3921, N3904, N2850, N2195, N2261);
or OR3 (N3922, N3920, N3279, N1953);
xor XOR2 (N3923, N3909, N1057);
and AND2 (N3924, N3916, N2051);
not NOT1 (N3925, N3906);
nand NAND3 (N3926, N3915, N1570, N875);
or OR4 (N3927, N3924, N807, N3005, N3482);
xor XOR2 (N3928, N3919, N2496);
nand NAND2 (N3929, N3918, N3435);
buf BUF1 (N3930, N3927);
or OR3 (N3931, N3921, N2119, N2181);
xor XOR2 (N3932, N3926, N999);
and AND4 (N3933, N3925, N1366, N1328, N3383);
and AND3 (N3934, N3913, N1048, N2806);
not NOT1 (N3935, N3929);
buf BUF1 (N3936, N3933);
not NOT1 (N3937, N3934);
and AND2 (N3938, N3930, N2932);
nand NAND4 (N3939, N3937, N2390, N431, N2534);
nor NOR4 (N3940, N3931, N3241, N1321, N2015);
xor XOR2 (N3941, N3932, N3151);
not NOT1 (N3942, N3935);
not NOT1 (N3943, N3922);
and AND4 (N3944, N3943, N1099, N3465, N1694);
or OR3 (N3945, N3940, N3465, N43);
or OR4 (N3946, N3923, N3801, N2449, N1605);
buf BUF1 (N3947, N3945);
and AND3 (N3948, N3911, N2470, N3298);
and AND4 (N3949, N3939, N3251, N2732, N170);
xor XOR2 (N3950, N3938, N954);
nor NOR2 (N3951, N3928, N2092);
nor NOR2 (N3952, N3950, N3337);
not NOT1 (N3953, N3936);
and AND4 (N3954, N3949, N3541, N2655, N2506);
nor NOR4 (N3955, N3953, N971, N3533, N1977);
or OR4 (N3956, N3941, N2147, N2041, N2969);
and AND4 (N3957, N3955, N1288, N3374, N3771);
xor XOR2 (N3958, N3956, N3544);
nor NOR2 (N3959, N3958, N2469);
nor NOR4 (N3960, N3957, N1449, N132, N3593);
nand NAND4 (N3961, N3946, N1536, N816, N1330);
nor NOR3 (N3962, N3952, N3162, N603);
buf BUF1 (N3963, N3944);
and AND3 (N3964, N3951, N1923, N1563);
buf BUF1 (N3965, N3964);
buf BUF1 (N3966, N3959);
not NOT1 (N3967, N3954);
or OR4 (N3968, N3961, N2283, N1582, N3538);
buf BUF1 (N3969, N3947);
and AND2 (N3970, N3963, N2623);
nand NAND4 (N3971, N3966, N249, N3934, N1936);
not NOT1 (N3972, N3968);
or OR2 (N3973, N3948, N2695);
and AND4 (N3974, N3965, N1531, N3689, N663);
nor NOR3 (N3975, N3942, N2201, N1615);
nor NOR2 (N3976, N3971, N3347);
buf BUF1 (N3977, N3972);
and AND4 (N3978, N3967, N2099, N1584, N873);
nand NAND2 (N3979, N3978, N2348);
or OR2 (N3980, N3974, N3284);
or OR4 (N3981, N3979, N336, N3898, N1738);
nor NOR4 (N3982, N3973, N802, N3951, N2403);
buf BUF1 (N3983, N3975);
xor XOR2 (N3984, N3960, N138);
and AND3 (N3985, N3970, N3725, N2594);
nand NAND4 (N3986, N3982, N2669, N2232, N2001);
nor NOR4 (N3987, N3962, N2177, N3243, N703);
nor NOR4 (N3988, N3980, N3716, N886, N3401);
and AND4 (N3989, N3988, N1109, N1852, N3883);
nor NOR4 (N3990, N3981, N1131, N938, N2966);
nor NOR3 (N3991, N3985, N1209, N2457);
nor NOR4 (N3992, N3983, N2559, N262, N1215);
and AND4 (N3993, N3976, N127, N3191, N884);
nand NAND2 (N3994, N3993, N1826);
buf BUF1 (N3995, N3992);
xor XOR2 (N3996, N3986, N3139);
not NOT1 (N3997, N3995);
or OR4 (N3998, N3989, N2521, N3370, N906);
or OR2 (N3999, N3984, N1872);
buf BUF1 (N4000, N3994);
not NOT1 (N4001, N3997);
not NOT1 (N4002, N4000);
not NOT1 (N4003, N3977);
xor XOR2 (N4004, N4001, N1141);
or OR2 (N4005, N4002, N571);
buf BUF1 (N4006, N3999);
xor XOR2 (N4007, N3996, N1896);
nand NAND3 (N4008, N3969, N3746, N3189);
nand NAND3 (N4009, N4004, N2700, N1787);
nand NAND3 (N4010, N4009, N2220, N3705);
nor NOR3 (N4011, N4003, N2041, N274);
and AND2 (N4012, N3990, N3217);
not NOT1 (N4013, N4008);
xor XOR2 (N4014, N4007, N2936);
not NOT1 (N4015, N3991);
nor NOR3 (N4016, N4013, N1200, N3088);
nor NOR3 (N4017, N4006, N1421, N1077);
not NOT1 (N4018, N3998);
nand NAND3 (N4019, N4016, N1331, N2008);
and AND4 (N4020, N4014, N407, N3493, N1792);
nand NAND3 (N4021, N4019, N1808, N1457);
nor NOR4 (N4022, N4011, N56, N1100, N2851);
not NOT1 (N4023, N4018);
buf BUF1 (N4024, N4010);
and AND4 (N4025, N4015, N3497, N2564, N244);
or OR3 (N4026, N4020, N2415, N488);
or OR2 (N4027, N4026, N3280);
buf BUF1 (N4028, N4022);
or OR3 (N4029, N4027, N2863, N892);
nor NOR3 (N4030, N4024, N3140, N3454);
and AND2 (N4031, N4012, N746);
or OR3 (N4032, N4031, N580, N149);
nor NOR3 (N4033, N4030, N3837, N122);
nand NAND3 (N4034, N4033, N3811, N117);
not NOT1 (N4035, N4005);
nand NAND2 (N4036, N4025, N3731);
xor XOR2 (N4037, N4028, N984);
or OR2 (N4038, N4017, N2281);
xor XOR2 (N4039, N4032, N1451);
not NOT1 (N4040, N4021);
and AND2 (N4041, N4036, N205);
and AND4 (N4042, N4035, N3803, N3744, N828);
xor XOR2 (N4043, N4039, N3666);
xor XOR2 (N4044, N4040, N3467);
buf BUF1 (N4045, N3987);
nand NAND2 (N4046, N4042, N1819);
or OR3 (N4047, N4046, N2459, N3966);
or OR3 (N4048, N4037, N2844, N2902);
buf BUF1 (N4049, N4038);
nor NOR4 (N4050, N4047, N1388, N2142, N3040);
xor XOR2 (N4051, N4044, N147);
or OR3 (N4052, N4029, N1244, N1969);
or OR4 (N4053, N4052, N3573, N1827, N3968);
xor XOR2 (N4054, N4048, N2668);
xor XOR2 (N4055, N4053, N1568);
and AND3 (N4056, N4041, N1342, N364);
xor XOR2 (N4057, N4050, N1003);
nand NAND4 (N4058, N4043, N3983, N1928, N3662);
and AND4 (N4059, N4056, N2398, N3530, N2903);
and AND2 (N4060, N4058, N3464);
buf BUF1 (N4061, N4055);
xor XOR2 (N4062, N4045, N1965);
and AND2 (N4063, N4057, N2168);
xor XOR2 (N4064, N4051, N3790);
nor NOR3 (N4065, N4063, N703, N2518);
not NOT1 (N4066, N4065);
nand NAND4 (N4067, N4064, N2291, N3490, N3846);
and AND2 (N4068, N4034, N3424);
and AND2 (N4069, N4066, N2689);
and AND3 (N4070, N4061, N2363, N341);
and AND4 (N4071, N4070, N2014, N601, N2652);
buf BUF1 (N4072, N4062);
and AND3 (N4073, N4049, N2890, N1949);
xor XOR2 (N4074, N4060, N2448);
buf BUF1 (N4075, N4068);
or OR3 (N4076, N4074, N2735, N3469);
not NOT1 (N4077, N4059);
or OR4 (N4078, N4054, N1246, N623, N3365);
nand NAND4 (N4079, N4071, N3059, N3260, N1523);
xor XOR2 (N4080, N4073, N814);
buf BUF1 (N4081, N4075);
not NOT1 (N4082, N4076);
not NOT1 (N4083, N4082);
or OR3 (N4084, N4080, N593, N3484);
xor XOR2 (N4085, N4084, N2093);
or OR4 (N4086, N4023, N3354, N3198, N3574);
and AND2 (N4087, N4085, N1329);
nor NOR4 (N4088, N4067, N343, N3551, N2224);
nand NAND3 (N4089, N4078, N3901, N2631);
or OR4 (N4090, N4079, N2528, N3342, N1682);
or OR2 (N4091, N4072, N2013);
xor XOR2 (N4092, N4089, N1433);
not NOT1 (N4093, N4086);
nand NAND3 (N4094, N4083, N2960, N3202);
xor XOR2 (N4095, N4081, N2273);
nand NAND3 (N4096, N4088, N1739, N2738);
nor NOR2 (N4097, N4091, N227);
not NOT1 (N4098, N4087);
not NOT1 (N4099, N4094);
not NOT1 (N4100, N4099);
xor XOR2 (N4101, N4090, N821);
and AND4 (N4102, N4097, N1280, N2440, N319);
or OR2 (N4103, N4100, N3588);
xor XOR2 (N4104, N4101, N3927);
not NOT1 (N4105, N4102);
xor XOR2 (N4106, N4105, N3745);
nand NAND2 (N4107, N4095, N3023);
nor NOR2 (N4108, N4069, N3680);
xor XOR2 (N4109, N4077, N735);
nor NOR4 (N4110, N4104, N2409, N250, N1958);
nand NAND3 (N4111, N4092, N2347, N4087);
buf BUF1 (N4112, N4093);
or OR2 (N4113, N4107, N3848);
nand NAND3 (N4114, N4108, N448, N483);
or OR3 (N4115, N4098, N2898, N530);
nand NAND3 (N4116, N4113, N808, N2928);
xor XOR2 (N4117, N4111, N3816);
buf BUF1 (N4118, N4112);
buf BUF1 (N4119, N4116);
nor NOR2 (N4120, N4114, N768);
not NOT1 (N4121, N4119);
and AND2 (N4122, N4103, N1456);
and AND2 (N4123, N4110, N3260);
and AND3 (N4124, N4121, N564, N1592);
not NOT1 (N4125, N4124);
or OR4 (N4126, N4117, N2028, N1845, N3767);
or OR3 (N4127, N4109, N3823, N3004);
or OR3 (N4128, N4115, N1405, N1642);
not NOT1 (N4129, N4123);
nand NAND2 (N4130, N4118, N140);
nor NOR3 (N4131, N4128, N3130, N2026);
or OR2 (N4132, N4096, N2360);
nor NOR2 (N4133, N4126, N3192);
nor NOR3 (N4134, N4120, N2290, N336);
buf BUF1 (N4135, N4122);
or OR2 (N4136, N4106, N1839);
or OR4 (N4137, N4135, N983, N3222, N3075);
not NOT1 (N4138, N4129);
xor XOR2 (N4139, N4133, N830);
xor XOR2 (N4140, N4138, N3364);
and AND2 (N4141, N4125, N3292);
not NOT1 (N4142, N4132);
buf BUF1 (N4143, N4134);
and AND3 (N4144, N4139, N3468, N3000);
nor NOR4 (N4145, N4144, N4082, N2576, N963);
nor NOR4 (N4146, N4136, N1858, N4101, N1502);
xor XOR2 (N4147, N4146, N2195);
buf BUF1 (N4148, N4147);
or OR2 (N4149, N4142, N743);
nor NOR4 (N4150, N4127, N3070, N4005, N3720);
nor NOR2 (N4151, N4141, N2558);
nor NOR4 (N4152, N4148, N3758, N305, N2778);
and AND3 (N4153, N4130, N2186, N260);
or OR4 (N4154, N4143, N3813, N2424, N3161);
buf BUF1 (N4155, N4153);
xor XOR2 (N4156, N4152, N2155);
not NOT1 (N4157, N4151);
and AND4 (N4158, N4157, N3865, N3761, N879);
xor XOR2 (N4159, N4137, N2890);
nand NAND3 (N4160, N4140, N687, N2819);
xor XOR2 (N4161, N4155, N2354);
or OR3 (N4162, N4160, N612, N3415);
nor NOR4 (N4163, N4149, N565, N3563, N3826);
or OR4 (N4164, N4150, N3957, N3783, N3971);
nand NAND2 (N4165, N4156, N2596);
nor NOR2 (N4166, N4164, N124);
nor NOR4 (N4167, N4161, N555, N3323, N3735);
xor XOR2 (N4168, N4145, N2276);
not NOT1 (N4169, N4167);
nor NOR3 (N4170, N4159, N2637, N2504);
not NOT1 (N4171, N4163);
xor XOR2 (N4172, N4166, N3882);
or OR4 (N4173, N4169, N3709, N3716, N774);
and AND4 (N4174, N4170, N1364, N2116, N1140);
not NOT1 (N4175, N4165);
or OR2 (N4176, N4168, N3787);
nand NAND2 (N4177, N4174, N2372);
not NOT1 (N4178, N4162);
or OR2 (N4179, N4176, N4005);
xor XOR2 (N4180, N4154, N1622);
nand NAND2 (N4181, N4177, N2505);
or OR4 (N4182, N4173, N4015, N2636, N3552);
nand NAND4 (N4183, N4180, N252, N311, N3347);
not NOT1 (N4184, N4181);
nor NOR2 (N4185, N4183, N2530);
nand NAND4 (N4186, N4185, N1823, N2301, N748);
nand NAND2 (N4187, N4179, N3752);
buf BUF1 (N4188, N4171);
buf BUF1 (N4189, N4186);
xor XOR2 (N4190, N4187, N3268);
not NOT1 (N4191, N4172);
and AND4 (N4192, N4175, N1676, N1226, N2371);
and AND2 (N4193, N4158, N3198);
xor XOR2 (N4194, N4188, N3918);
buf BUF1 (N4195, N4194);
not NOT1 (N4196, N4195);
and AND4 (N4197, N4184, N221, N662, N3357);
and AND2 (N4198, N4193, N2204);
buf BUF1 (N4199, N4131);
nand NAND4 (N4200, N4196, N1710, N3843, N714);
buf BUF1 (N4201, N4198);
xor XOR2 (N4202, N4182, N626);
buf BUF1 (N4203, N4191);
xor XOR2 (N4204, N4197, N1167);
nor NOR4 (N4205, N4192, N4003, N1309, N997);
not NOT1 (N4206, N4189);
nand NAND2 (N4207, N4199, N3183);
nor NOR4 (N4208, N4203, N1998, N2705, N1440);
nand NAND4 (N4209, N4200, N1810, N243, N3222);
or OR4 (N4210, N4190, N707, N335, N3752);
nand NAND2 (N4211, N4202, N511);
xor XOR2 (N4212, N4201, N3073);
nand NAND4 (N4213, N4211, N324, N1838, N1436);
buf BUF1 (N4214, N4206);
nand NAND4 (N4215, N4214, N3551, N2238, N688);
or OR3 (N4216, N4212, N1728, N529);
and AND3 (N4217, N4178, N1436, N3439);
nand NAND2 (N4218, N4215, N2287);
nand NAND3 (N4219, N4217, N1801, N3829);
nand NAND3 (N4220, N4207, N1900, N717);
nor NOR4 (N4221, N4213, N4065, N2454, N3535);
and AND3 (N4222, N4204, N170, N147);
xor XOR2 (N4223, N4210, N220);
or OR4 (N4224, N4218, N3636, N1549, N4069);
nand NAND2 (N4225, N4222, N2582);
nor NOR2 (N4226, N4221, N4189);
and AND3 (N4227, N4205, N2990, N596);
nand NAND3 (N4228, N4216, N314, N3808);
nand NAND2 (N4229, N4224, N2297);
buf BUF1 (N4230, N4223);
nor NOR3 (N4231, N4227, N3563, N2087);
or OR3 (N4232, N4208, N4017, N667);
nand NAND3 (N4233, N4225, N1461, N3352);
buf BUF1 (N4234, N4229);
or OR4 (N4235, N4220, N1718, N2299, N2475);
and AND4 (N4236, N4209, N4045, N1311, N136);
or OR3 (N4237, N4234, N996, N2655);
nand NAND3 (N4238, N4226, N3701, N1808);
buf BUF1 (N4239, N4235);
buf BUF1 (N4240, N4237);
not NOT1 (N4241, N4238);
not NOT1 (N4242, N4239);
or OR3 (N4243, N4236, N1162, N3916);
xor XOR2 (N4244, N4233, N3163);
and AND3 (N4245, N4243, N2706, N3809);
xor XOR2 (N4246, N4232, N979);
not NOT1 (N4247, N4230);
buf BUF1 (N4248, N4241);
nand NAND3 (N4249, N4248, N2644, N2416);
or OR4 (N4250, N4249, N3451, N2844, N3438);
and AND4 (N4251, N4247, N913, N3434, N1268);
and AND3 (N4252, N4246, N2468, N2601);
and AND4 (N4253, N4250, N1628, N438, N4198);
nor NOR2 (N4254, N4228, N3747);
and AND4 (N4255, N4254, N73, N1137, N1507);
buf BUF1 (N4256, N4252);
buf BUF1 (N4257, N4244);
or OR3 (N4258, N4240, N2579, N2126);
nand NAND4 (N4259, N4219, N1369, N2194, N3726);
or OR2 (N4260, N4259, N1406);
and AND2 (N4261, N4258, N2670);
buf BUF1 (N4262, N4256);
nor NOR2 (N4263, N4231, N1615);
xor XOR2 (N4264, N4255, N1602);
nor NOR4 (N4265, N4264, N3497, N907, N3174);
nor NOR3 (N4266, N4253, N2513, N73);
buf BUF1 (N4267, N4251);
buf BUF1 (N4268, N4245);
nand NAND3 (N4269, N4263, N2162, N3572);
or OR3 (N4270, N4266, N379, N1622);
or OR4 (N4271, N4268, N3823, N2117, N1534);
nand NAND4 (N4272, N4271, N2072, N2046, N3706);
nand NAND3 (N4273, N4265, N3992, N3787);
and AND4 (N4274, N4273, N4194, N3759, N4048);
nor NOR2 (N4275, N4269, N2199);
nor NOR3 (N4276, N4272, N103, N2252);
nor NOR3 (N4277, N4262, N3585, N4040);
buf BUF1 (N4278, N4274);
not NOT1 (N4279, N4260);
and AND3 (N4280, N4242, N2955, N2365);
not NOT1 (N4281, N4278);
not NOT1 (N4282, N4276);
nand NAND3 (N4283, N4277, N827, N4110);
or OR4 (N4284, N4261, N3673, N2321, N2911);
or OR2 (N4285, N4283, N3959);
xor XOR2 (N4286, N4270, N2799);
buf BUF1 (N4287, N4286);
or OR2 (N4288, N4275, N2454);
nor NOR2 (N4289, N4282, N2219);
not NOT1 (N4290, N4284);
nor NOR3 (N4291, N4290, N2576, N467);
nand NAND4 (N4292, N4289, N1422, N2829, N793);
xor XOR2 (N4293, N4285, N2339);
not NOT1 (N4294, N4291);
or OR4 (N4295, N4292, N2021, N1870, N1328);
nand NAND3 (N4296, N4295, N1435, N3304);
buf BUF1 (N4297, N4279);
buf BUF1 (N4298, N4294);
nand NAND2 (N4299, N4288, N602);
buf BUF1 (N4300, N4281);
nand NAND2 (N4301, N4299, N189);
not NOT1 (N4302, N4257);
buf BUF1 (N4303, N4296);
or OR4 (N4304, N4267, N4252, N580, N849);
nand NAND3 (N4305, N4293, N3917, N2785);
or OR4 (N4306, N4301, N2492, N2003, N357);
xor XOR2 (N4307, N4298, N3872);
and AND3 (N4308, N4302, N1682, N4010);
not NOT1 (N4309, N4280);
nor NOR4 (N4310, N4303, N4246, N4148, N3234);
and AND2 (N4311, N4305, N1839);
and AND3 (N4312, N4287, N759, N2078);
nand NAND2 (N4313, N4309, N4048);
or OR4 (N4314, N4297, N3523, N2316, N1977);
nand NAND2 (N4315, N4307, N363);
nor NOR3 (N4316, N4306, N623, N804);
not NOT1 (N4317, N4304);
nor NOR2 (N4318, N4316, N128);
buf BUF1 (N4319, N4315);
nand NAND3 (N4320, N4319, N4191, N124);
xor XOR2 (N4321, N4317, N380);
and AND3 (N4322, N4314, N2383, N602);
xor XOR2 (N4323, N4310, N2915);
not NOT1 (N4324, N4312);
xor XOR2 (N4325, N4323, N3256);
nor NOR4 (N4326, N4300, N1198, N2069, N983);
or OR3 (N4327, N4320, N2930, N947);
or OR2 (N4328, N4326, N1536);
or OR3 (N4329, N4311, N807, N3740);
not NOT1 (N4330, N4313);
or OR3 (N4331, N4308, N2647, N1022);
nand NAND2 (N4332, N4329, N2029);
xor XOR2 (N4333, N4327, N3548);
and AND3 (N4334, N4318, N499, N2586);
not NOT1 (N4335, N4328);
nand NAND4 (N4336, N4325, N604, N3174, N2770);
nand NAND3 (N4337, N4333, N2651, N1911);
or OR2 (N4338, N4332, N413);
not NOT1 (N4339, N4337);
or OR2 (N4340, N4339, N1151);
xor XOR2 (N4341, N4331, N3438);
nand NAND3 (N4342, N4334, N1343, N450);
or OR4 (N4343, N4335, N3366, N3586, N4251);
nand NAND3 (N4344, N4341, N2467, N3522);
not NOT1 (N4345, N4321);
and AND4 (N4346, N4330, N3847, N3618, N276);
buf BUF1 (N4347, N4343);
or OR3 (N4348, N4324, N197, N546);
and AND3 (N4349, N4336, N4227, N1357);
not NOT1 (N4350, N4338);
buf BUF1 (N4351, N4349);
xor XOR2 (N4352, N4346, N802);
xor XOR2 (N4353, N4342, N3313);
nand NAND4 (N4354, N4344, N1252, N1598, N488);
xor XOR2 (N4355, N4348, N3401);
xor XOR2 (N4356, N4347, N2032);
buf BUF1 (N4357, N4353);
buf BUF1 (N4358, N4350);
or OR3 (N4359, N4352, N416, N2843);
xor XOR2 (N4360, N4355, N3262);
nand NAND4 (N4361, N4356, N2172, N2095, N2055);
not NOT1 (N4362, N4358);
nor NOR3 (N4363, N4351, N1627, N1117);
nand NAND2 (N4364, N4359, N3294);
nand NAND2 (N4365, N4363, N823);
and AND2 (N4366, N4354, N967);
nand NAND4 (N4367, N4340, N2320, N3639, N3420);
xor XOR2 (N4368, N4364, N677);
or OR2 (N4369, N4365, N358);
buf BUF1 (N4370, N4367);
not NOT1 (N4371, N4370);
xor XOR2 (N4372, N4345, N724);
and AND4 (N4373, N4368, N714, N3080, N2931);
and AND3 (N4374, N4369, N2874, N642);
xor XOR2 (N4375, N4371, N580);
nand NAND3 (N4376, N4322, N3019, N2346);
and AND4 (N4377, N4360, N3637, N2287, N1037);
xor XOR2 (N4378, N4374, N2878);
xor XOR2 (N4379, N4362, N14);
nand NAND3 (N4380, N4375, N1811, N3868);
nor NOR4 (N4381, N4378, N3806, N2306, N518);
or OR3 (N4382, N4366, N3731, N4301);
nand NAND4 (N4383, N4372, N4265, N2937, N1811);
xor XOR2 (N4384, N4376, N346);
nand NAND2 (N4385, N4383, N1849);
and AND4 (N4386, N4384, N49, N2106, N3734);
nor NOR3 (N4387, N4380, N3158, N3978);
or OR2 (N4388, N4361, N1123);
nand NAND3 (N4389, N4377, N1916, N4111);
not NOT1 (N4390, N4381);
or OR4 (N4391, N4386, N2631, N2429, N3166);
not NOT1 (N4392, N4387);
buf BUF1 (N4393, N4357);
nand NAND4 (N4394, N4392, N3344, N2832, N3786);
and AND4 (N4395, N4389, N2240, N3965, N517);
not NOT1 (N4396, N4394);
and AND3 (N4397, N4395, N1753, N1064);
nand NAND4 (N4398, N4397, N2249, N3967, N3722);
not NOT1 (N4399, N4391);
xor XOR2 (N4400, N4390, N924);
and AND2 (N4401, N4400, N1721);
nand NAND3 (N4402, N4388, N3045, N4214);
xor XOR2 (N4403, N4379, N1103);
or OR4 (N4404, N4398, N4345, N3597, N723);
and AND2 (N4405, N4399, N2414);
buf BUF1 (N4406, N4396);
or OR3 (N4407, N4405, N109, N2824);
buf BUF1 (N4408, N4373);
xor XOR2 (N4409, N4408, N3840);
xor XOR2 (N4410, N4404, N1052);
nand NAND4 (N4411, N4410, N1378, N3626, N2214);
buf BUF1 (N4412, N4407);
and AND4 (N4413, N4409, N2941, N2759, N3944);
xor XOR2 (N4414, N4393, N1355);
buf BUF1 (N4415, N4413);
not NOT1 (N4416, N4411);
not NOT1 (N4417, N4401);
buf BUF1 (N4418, N4416);
nor NOR3 (N4419, N4382, N1938, N740);
buf BUF1 (N4420, N4415);
nand NAND4 (N4421, N4406, N2888, N2944, N543);
not NOT1 (N4422, N4403);
and AND2 (N4423, N4385, N56);
buf BUF1 (N4424, N4418);
not NOT1 (N4425, N4420);
nor NOR2 (N4426, N4424, N2225);
buf BUF1 (N4427, N4417);
not NOT1 (N4428, N4419);
not NOT1 (N4429, N4412);
not NOT1 (N4430, N4414);
and AND3 (N4431, N4426, N2279, N3827);
nor NOR4 (N4432, N4402, N1365, N2597, N3850);
nand NAND2 (N4433, N4425, N3846);
and AND3 (N4434, N4429, N2379, N3865);
nand NAND4 (N4435, N4421, N181, N703, N3317);
xor XOR2 (N4436, N4431, N1180);
and AND2 (N4437, N4434, N1842);
nor NOR4 (N4438, N4436, N1700, N1042, N2612);
buf BUF1 (N4439, N4423);
or OR3 (N4440, N4435, N2848, N4114);
and AND2 (N4441, N4430, N3350);
and AND2 (N4442, N4441, N1778);
nor NOR4 (N4443, N4440, N861, N2795, N374);
not NOT1 (N4444, N4439);
nand NAND2 (N4445, N4433, N3635);
nand NAND3 (N4446, N4438, N2049, N4064);
and AND3 (N4447, N4428, N3260, N4373);
nand NAND4 (N4448, N4432, N2052, N3555, N2345);
buf BUF1 (N4449, N4422);
nand NAND3 (N4450, N4444, N3490, N2509);
nand NAND2 (N4451, N4437, N1119);
buf BUF1 (N4452, N4449);
buf BUF1 (N4453, N4443);
buf BUF1 (N4454, N4446);
nand NAND2 (N4455, N4454, N2308);
not NOT1 (N4456, N4453);
or OR4 (N4457, N4448, N719, N4276, N1984);
and AND4 (N4458, N4427, N3834, N3699, N288);
and AND2 (N4459, N4450, N4115);
and AND3 (N4460, N4451, N1641, N840);
not NOT1 (N4461, N4460);
nor NOR2 (N4462, N4456, N4062);
and AND3 (N4463, N4459, N3607, N4029);
and AND4 (N4464, N4442, N2341, N3276, N3206);
not NOT1 (N4465, N4447);
nand NAND2 (N4466, N4457, N2671);
nand NAND4 (N4467, N4464, N757, N69, N2176);
not NOT1 (N4468, N4465);
and AND2 (N4469, N4468, N2488);
nand NAND3 (N4470, N4445, N2669, N84);
nor NOR4 (N4471, N4455, N2234, N1421, N4096);
and AND3 (N4472, N4458, N3057, N3696);
buf BUF1 (N4473, N4461);
nor NOR4 (N4474, N4452, N812, N2607, N189);
buf BUF1 (N4475, N4470);
and AND3 (N4476, N4474, N2805, N2755);
nor NOR4 (N4477, N4476, N4431, N2676, N1710);
not NOT1 (N4478, N4466);
and AND4 (N4479, N4478, N276, N80, N1572);
xor XOR2 (N4480, N4473, N1635);
not NOT1 (N4481, N4462);
nand NAND4 (N4482, N4480, N1414, N2319, N3481);
nor NOR4 (N4483, N4482, N2951, N1051, N57);
or OR4 (N4484, N4475, N3382, N3771, N1175);
nor NOR3 (N4485, N4469, N3472, N698);
or OR4 (N4486, N4471, N1660, N1199, N4431);
nand NAND3 (N4487, N4479, N549, N4294);
xor XOR2 (N4488, N4467, N861);
and AND4 (N4489, N4472, N77, N1049, N3657);
nor NOR3 (N4490, N4486, N1480, N2971);
or OR3 (N4491, N4481, N315, N1391);
buf BUF1 (N4492, N4483);
and AND2 (N4493, N4488, N35);
buf BUF1 (N4494, N4489);
nand NAND3 (N4495, N4487, N213, N4057);
xor XOR2 (N4496, N4491, N3698);
nand NAND3 (N4497, N4495, N4256, N1074);
nor NOR2 (N4498, N4493, N37);
and AND2 (N4499, N4484, N2153);
nor NOR4 (N4500, N4490, N1712, N1700, N2196);
nor NOR3 (N4501, N4494, N3652, N2940);
not NOT1 (N4502, N4500);
or OR4 (N4503, N4492, N896, N188, N4451);
nand NAND4 (N4504, N4503, N3927, N2519, N3930);
buf BUF1 (N4505, N4501);
not NOT1 (N4506, N4504);
not NOT1 (N4507, N4496);
and AND2 (N4508, N4505, N1332);
not NOT1 (N4509, N4485);
or OR4 (N4510, N4508, N4364, N3724, N424);
not NOT1 (N4511, N4507);
nand NAND3 (N4512, N4499, N138, N1272);
or OR2 (N4513, N4509, N2896);
buf BUF1 (N4514, N4498);
or OR2 (N4515, N4512, N1262);
and AND4 (N4516, N4506, N4314, N1854, N1196);
nor NOR4 (N4517, N4477, N3694, N3484, N3861);
nor NOR2 (N4518, N4517, N18);
or OR4 (N4519, N4516, N2172, N1668, N971);
xor XOR2 (N4520, N4515, N2297);
not NOT1 (N4521, N4511);
xor XOR2 (N4522, N4514, N2699);
buf BUF1 (N4523, N4510);
or OR2 (N4524, N4522, N448);
nor NOR2 (N4525, N4502, N1862);
xor XOR2 (N4526, N4497, N2275);
not NOT1 (N4527, N4518);
xor XOR2 (N4528, N4525, N1817);
and AND2 (N4529, N4520, N1173);
xor XOR2 (N4530, N4523, N1909);
not NOT1 (N4531, N4513);
or OR3 (N4532, N4529, N1402, N4406);
not NOT1 (N4533, N4463);
or OR3 (N4534, N4530, N3657, N2875);
or OR4 (N4535, N4527, N1697, N2254, N3533);
not NOT1 (N4536, N4519);
or OR2 (N4537, N4532, N1391);
not NOT1 (N4538, N4528);
and AND2 (N4539, N4521, N1591);
nor NOR3 (N4540, N4537, N1542, N1295);
or OR4 (N4541, N4539, N1028, N1229, N980);
or OR2 (N4542, N4526, N3116);
not NOT1 (N4543, N4538);
buf BUF1 (N4544, N4540);
not NOT1 (N4545, N4524);
not NOT1 (N4546, N4543);
nor NOR4 (N4547, N4544, N4214, N3606, N2249);
and AND3 (N4548, N4546, N197, N2025);
and AND3 (N4549, N4534, N4078, N4181);
not NOT1 (N4550, N4548);
and AND3 (N4551, N4533, N720, N387);
not NOT1 (N4552, N4535);
nand NAND2 (N4553, N4547, N101);
and AND3 (N4554, N4541, N3134, N655);
nand NAND4 (N4555, N4553, N618, N1803, N1923);
and AND3 (N4556, N4555, N3254, N795);
nand NAND3 (N4557, N4556, N4266, N352);
not NOT1 (N4558, N4536);
nor NOR2 (N4559, N4550, N1931);
not NOT1 (N4560, N4549);
nor NOR2 (N4561, N4554, N4421);
xor XOR2 (N4562, N4561, N4466);
not NOT1 (N4563, N4552);
or OR2 (N4564, N4563, N490);
buf BUF1 (N4565, N4564);
xor XOR2 (N4566, N4562, N1493);
nor NOR3 (N4567, N4542, N2118, N1738);
xor XOR2 (N4568, N4545, N3257);
nand NAND3 (N4569, N4559, N3224, N3176);
and AND4 (N4570, N4558, N1944, N53, N2338);
buf BUF1 (N4571, N4566);
not NOT1 (N4572, N4551);
xor XOR2 (N4573, N4531, N2179);
not NOT1 (N4574, N4557);
nand NAND2 (N4575, N4568, N4100);
nor NOR2 (N4576, N4567, N2689);
not NOT1 (N4577, N4569);
or OR4 (N4578, N4560, N1330, N1865, N2386);
nand NAND2 (N4579, N4574, N1050);
buf BUF1 (N4580, N4577);
nand NAND3 (N4581, N4571, N3790, N2324);
nor NOR2 (N4582, N4578, N1531);
and AND3 (N4583, N4582, N893, N2750);
buf BUF1 (N4584, N4575);
nand NAND4 (N4585, N4570, N3881, N1496, N2383);
and AND4 (N4586, N4579, N178, N329, N743);
nor NOR2 (N4587, N4572, N257);
nand NAND3 (N4588, N4573, N1737, N1747);
nor NOR4 (N4589, N4588, N951, N4138, N2812);
not NOT1 (N4590, N4581);
not NOT1 (N4591, N4584);
or OR4 (N4592, N4590, N1542, N3596, N112);
not NOT1 (N4593, N4585);
or OR2 (N4594, N4576, N2937);
and AND3 (N4595, N4565, N1762, N700);
xor XOR2 (N4596, N4587, N2985);
xor XOR2 (N4597, N4586, N2038);
and AND3 (N4598, N4595, N2435, N2885);
nor NOR2 (N4599, N4593, N2513);
xor XOR2 (N4600, N4599, N3523);
xor XOR2 (N4601, N4589, N4333);
buf BUF1 (N4602, N4592);
nor NOR4 (N4603, N4596, N2392, N4011, N1385);
not NOT1 (N4604, N4602);
buf BUF1 (N4605, N4604);
and AND3 (N4606, N4583, N4093, N2073);
nor NOR2 (N4607, N4591, N2516);
nor NOR4 (N4608, N4603, N1830, N2774, N4461);
xor XOR2 (N4609, N4608, N462);
or OR4 (N4610, N4597, N1317, N2913, N1564);
not NOT1 (N4611, N4598);
buf BUF1 (N4612, N4601);
or OR4 (N4613, N4580, N824, N2268, N2124);
xor XOR2 (N4614, N4611, N188);
and AND3 (N4615, N4613, N3842, N3386);
and AND4 (N4616, N4600, N4180, N3546, N3386);
and AND2 (N4617, N4609, N3446);
nand NAND2 (N4618, N4615, N3289);
not NOT1 (N4619, N4618);
nand NAND3 (N4620, N4606, N4580, N3737);
xor XOR2 (N4621, N4616, N333);
and AND2 (N4622, N4610, N1183);
xor XOR2 (N4623, N4594, N2438);
or OR2 (N4624, N4622, N2162);
or OR3 (N4625, N4607, N2526, N3188);
nor NOR4 (N4626, N4612, N1264, N2234, N2827);
not NOT1 (N4627, N4605);
not NOT1 (N4628, N4619);
xor XOR2 (N4629, N4624, N1202);
not NOT1 (N4630, N4620);
nand NAND4 (N4631, N4629, N1575, N1546, N2019);
not NOT1 (N4632, N4617);
buf BUF1 (N4633, N4614);
nor NOR4 (N4634, N4631, N2484, N3416, N2933);
or OR4 (N4635, N4632, N2824, N2026, N1153);
or OR2 (N4636, N4634, N1518);
or OR3 (N4637, N4627, N4447, N9);
nor NOR4 (N4638, N4625, N2426, N4053, N2541);
nor NOR4 (N4639, N4638, N1281, N4171, N979);
nor NOR4 (N4640, N4636, N1671, N1783, N2052);
or OR4 (N4641, N4637, N636, N1027, N2859);
not NOT1 (N4642, N4623);
buf BUF1 (N4643, N4621);
or OR2 (N4644, N4641, N1922);
and AND2 (N4645, N4644, N340);
xor XOR2 (N4646, N4642, N2661);
nor NOR2 (N4647, N4633, N1305);
or OR3 (N4648, N4630, N577, N1686);
or OR4 (N4649, N4647, N3657, N3491, N3557);
xor XOR2 (N4650, N4646, N2446);
and AND4 (N4651, N4640, N4115, N3161, N1380);
nor NOR2 (N4652, N4651, N3775);
nor NOR2 (N4653, N4639, N667);
buf BUF1 (N4654, N4628);
xor XOR2 (N4655, N4648, N590);
nor NOR4 (N4656, N4626, N4560, N1456, N1684);
or OR4 (N4657, N4652, N2963, N2441, N2789);
buf BUF1 (N4658, N4655);
or OR3 (N4659, N4656, N2696, N2404);
or OR4 (N4660, N4649, N2856, N1391, N1648);
or OR4 (N4661, N4659, N1615, N2255, N772);
nand NAND4 (N4662, N4660, N2934, N1016, N1842);
not NOT1 (N4663, N4635);
not NOT1 (N4664, N4663);
and AND3 (N4665, N4650, N3905, N869);
xor XOR2 (N4666, N4657, N1841);
and AND3 (N4667, N4645, N3806, N1216);
nor NOR4 (N4668, N4653, N3218, N3190, N1605);
not NOT1 (N4669, N4667);
buf BUF1 (N4670, N4661);
not NOT1 (N4671, N4662);
or OR4 (N4672, N4658, N978, N1130, N3419);
buf BUF1 (N4673, N4668);
nor NOR3 (N4674, N4643, N1346, N472);
or OR4 (N4675, N4664, N2891, N216, N3719);
or OR3 (N4676, N4672, N4015, N1314);
nor NOR2 (N4677, N4671, N1403);
or OR2 (N4678, N4677, N777);
or OR3 (N4679, N4675, N449, N4668);
xor XOR2 (N4680, N4670, N1283);
xor XOR2 (N4681, N4665, N4213);
nand NAND4 (N4682, N4681, N2252, N4595, N923);
xor XOR2 (N4683, N4682, N4356);
and AND2 (N4684, N4680, N2996);
nand NAND3 (N4685, N4678, N723, N1924);
xor XOR2 (N4686, N4679, N3668);
not NOT1 (N4687, N4676);
or OR3 (N4688, N4683, N3099, N4307);
xor XOR2 (N4689, N4684, N3583);
xor XOR2 (N4690, N4688, N4637);
buf BUF1 (N4691, N4654);
or OR4 (N4692, N4691, N308, N1470, N2026);
nand NAND3 (N4693, N4690, N3617, N2821);
nand NAND2 (N4694, N4693, N296);
and AND2 (N4695, N4687, N1784);
buf BUF1 (N4696, N4694);
nand NAND4 (N4697, N4689, N1319, N2002, N4520);
not NOT1 (N4698, N4673);
xor XOR2 (N4699, N4686, N1864);
or OR3 (N4700, N4674, N752, N1879);
buf BUF1 (N4701, N4698);
and AND2 (N4702, N4666, N2566);
and AND2 (N4703, N4702, N3694);
not NOT1 (N4704, N4685);
buf BUF1 (N4705, N4700);
nor NOR3 (N4706, N4705, N324, N2306);
not NOT1 (N4707, N4669);
or OR2 (N4708, N4696, N28);
nor NOR2 (N4709, N4699, N1298);
and AND2 (N4710, N4701, N4185);
buf BUF1 (N4711, N4692);
buf BUF1 (N4712, N4707);
not NOT1 (N4713, N4695);
not NOT1 (N4714, N4710);
and AND2 (N4715, N4697, N1564);
not NOT1 (N4716, N4713);
buf BUF1 (N4717, N4708);
or OR2 (N4718, N4714, N3763);
xor XOR2 (N4719, N4703, N2174);
not NOT1 (N4720, N4711);
not NOT1 (N4721, N4717);
nand NAND2 (N4722, N4706, N1819);
and AND4 (N4723, N4721, N1224, N2313, N4618);
nand NAND4 (N4724, N4718, N3157, N1538, N2441);
nor NOR2 (N4725, N4709, N1167);
xor XOR2 (N4726, N4722, N1787);
nor NOR2 (N4727, N4725, N4044);
and AND4 (N4728, N4727, N4376, N2004, N2197);
nand NAND3 (N4729, N4723, N2300, N4336);
buf BUF1 (N4730, N4724);
nand NAND2 (N4731, N4704, N4227);
or OR3 (N4732, N4731, N2564, N539);
nand NAND3 (N4733, N4715, N3845, N3803);
xor XOR2 (N4734, N4732, N1742);
xor XOR2 (N4735, N4716, N4713);
and AND3 (N4736, N4726, N3150, N4039);
and AND4 (N4737, N4728, N4678, N2916, N4230);
buf BUF1 (N4738, N4735);
or OR4 (N4739, N4736, N495, N4009, N1906);
or OR4 (N4740, N4719, N3582, N4246, N1154);
buf BUF1 (N4741, N4720);
or OR2 (N4742, N4733, N2229);
and AND4 (N4743, N4740, N3028, N491, N1691);
nor NOR3 (N4744, N4712, N582, N1871);
buf BUF1 (N4745, N4730);
or OR3 (N4746, N4744, N841, N1987);
or OR2 (N4747, N4734, N12);
xor XOR2 (N4748, N4738, N928);
not NOT1 (N4749, N4742);
and AND3 (N4750, N4737, N2387, N168);
and AND2 (N4751, N4749, N2679);
not NOT1 (N4752, N4747);
and AND4 (N4753, N4745, N4450, N1114, N65);
xor XOR2 (N4754, N4752, N4139);
not NOT1 (N4755, N4743);
nor NOR2 (N4756, N4753, N681);
not NOT1 (N4757, N4741);
and AND2 (N4758, N4750, N3609);
nor NOR2 (N4759, N4754, N723);
not NOT1 (N4760, N4755);
not NOT1 (N4761, N4757);
or OR3 (N4762, N4748, N4001, N4093);
nor NOR3 (N4763, N4759, N355, N1266);
buf BUF1 (N4764, N4746);
or OR3 (N4765, N4763, N2489, N3862);
nor NOR3 (N4766, N4760, N2664, N2871);
nand NAND4 (N4767, N4729, N2809, N338, N3844);
and AND2 (N4768, N4767, N4309);
nand NAND2 (N4769, N4751, N4636);
or OR2 (N4770, N4764, N421);
nand NAND4 (N4771, N4756, N407, N2168, N621);
nor NOR3 (N4772, N4761, N4232, N4016);
not NOT1 (N4773, N4769);
buf BUF1 (N4774, N4758);
not NOT1 (N4775, N4770);
nand NAND4 (N4776, N4775, N2707, N2495, N2268);
and AND4 (N4777, N4765, N3104, N3064, N4598);
or OR3 (N4778, N4766, N748, N1760);
nand NAND3 (N4779, N4768, N1665, N1358);
buf BUF1 (N4780, N4778);
xor XOR2 (N4781, N4773, N1685);
buf BUF1 (N4782, N4774);
xor XOR2 (N4783, N4780, N2340);
buf BUF1 (N4784, N4772);
and AND2 (N4785, N4779, N3421);
buf BUF1 (N4786, N4783);
not NOT1 (N4787, N4739);
xor XOR2 (N4788, N4787, N1142);
nor NOR3 (N4789, N4782, N583, N3747);
nand NAND4 (N4790, N4776, N3176, N1001, N4715);
nand NAND3 (N4791, N4771, N29, N2609);
buf BUF1 (N4792, N4788);
nand NAND2 (N4793, N4791, N3231);
and AND4 (N4794, N4792, N3559, N139, N1083);
not NOT1 (N4795, N4762);
nand NAND2 (N4796, N4789, N948);
or OR4 (N4797, N4784, N3837, N2999, N797);
or OR4 (N4798, N4781, N3207, N2188, N1013);
and AND3 (N4799, N4790, N3884, N3018);
xor XOR2 (N4800, N4793, N950);
or OR2 (N4801, N4786, N3388);
not NOT1 (N4802, N4799);
nor NOR2 (N4803, N4795, N114);
not NOT1 (N4804, N4803);
nand NAND2 (N4805, N4802, N3125);
not NOT1 (N4806, N4785);
buf BUF1 (N4807, N4805);
and AND3 (N4808, N4797, N3414, N2119);
nand NAND4 (N4809, N4804, N2269, N1073, N4188);
and AND4 (N4810, N4796, N442, N1594, N35);
not NOT1 (N4811, N4798);
or OR3 (N4812, N4811, N2724, N4198);
xor XOR2 (N4813, N4812, N3943);
and AND4 (N4814, N4813, N599, N615, N1888);
not NOT1 (N4815, N4794);
or OR4 (N4816, N4806, N987, N4473, N2188);
or OR4 (N4817, N4801, N4385, N2616, N2927);
and AND3 (N4818, N4800, N2536, N4630);
xor XOR2 (N4819, N4814, N3433);
or OR3 (N4820, N4807, N1249, N140);
nor NOR4 (N4821, N4810, N738, N4201, N3465);
buf BUF1 (N4822, N4815);
not NOT1 (N4823, N4818);
nor NOR2 (N4824, N4819, N2269);
nand NAND2 (N4825, N4817, N506);
xor XOR2 (N4826, N4808, N2435);
and AND2 (N4827, N4816, N2164);
buf BUF1 (N4828, N4809);
or OR2 (N4829, N4823, N1652);
not NOT1 (N4830, N4829);
buf BUF1 (N4831, N4830);
nor NOR4 (N4832, N4828, N2221, N1845, N4377);
nand NAND4 (N4833, N4826, N3091, N2001, N2314);
not NOT1 (N4834, N4832);
xor XOR2 (N4835, N4822, N3726);
or OR3 (N4836, N4835, N607, N2383);
xor XOR2 (N4837, N4833, N103);
buf BUF1 (N4838, N4837);
nand NAND2 (N4839, N4827, N3548);
and AND4 (N4840, N4820, N1626, N2874, N72);
nand NAND3 (N4841, N4838, N1368, N4027);
and AND4 (N4842, N4831, N2082, N1818, N4700);
and AND3 (N4843, N4824, N3924, N1920);
nand NAND4 (N4844, N4839, N493, N2095, N3693);
nand NAND2 (N4845, N4843, N2274);
xor XOR2 (N4846, N4825, N528);
or OR4 (N4847, N4834, N3738, N1141, N958);
nor NOR2 (N4848, N4836, N1224);
nor NOR3 (N4849, N4845, N1620, N3753);
or OR4 (N4850, N4842, N366, N931, N534);
buf BUF1 (N4851, N4777);
buf BUF1 (N4852, N4847);
xor XOR2 (N4853, N4841, N3600);
buf BUF1 (N4854, N4846);
buf BUF1 (N4855, N4848);
nand NAND2 (N4856, N4821, N256);
xor XOR2 (N4857, N4853, N3250);
nand NAND3 (N4858, N4844, N4086, N65);
buf BUF1 (N4859, N4852);
nor NOR4 (N4860, N4851, N3928, N1168, N3388);
buf BUF1 (N4861, N4860);
and AND3 (N4862, N4854, N1713, N571);
nor NOR4 (N4863, N4849, N2158, N4755, N4515);
not NOT1 (N4864, N4858);
and AND4 (N4865, N4855, N3190, N2310, N3988);
nand NAND2 (N4866, N4856, N4863);
or OR4 (N4867, N4501, N2330, N4115, N1935);
buf BUF1 (N4868, N4861);
nor NOR2 (N4869, N4840, N142);
xor XOR2 (N4870, N4869, N4713);
not NOT1 (N4871, N4857);
nand NAND4 (N4872, N4864, N3840, N774, N815);
or OR4 (N4873, N4868, N592, N3683, N4149);
xor XOR2 (N4874, N4862, N4279);
nand NAND4 (N4875, N4865, N2687, N291, N3179);
not NOT1 (N4876, N4872);
nand NAND2 (N4877, N4871, N1153);
nor NOR4 (N4878, N4850, N3988, N2824, N1610);
buf BUF1 (N4879, N4873);
xor XOR2 (N4880, N4867, N1954);
and AND3 (N4881, N4876, N2247, N470);
not NOT1 (N4882, N4874);
not NOT1 (N4883, N4882);
or OR2 (N4884, N4870, N2679);
and AND3 (N4885, N4866, N1439, N201);
buf BUF1 (N4886, N4875);
nor NOR2 (N4887, N4883, N3011);
buf BUF1 (N4888, N4880);
nor NOR2 (N4889, N4885, N4825);
or OR2 (N4890, N4877, N1254);
not NOT1 (N4891, N4889);
or OR3 (N4892, N4886, N721, N3898);
nand NAND4 (N4893, N4881, N928, N2337, N1783);
buf BUF1 (N4894, N4879);
buf BUF1 (N4895, N4884);
nor NOR2 (N4896, N4894, N4486);
and AND3 (N4897, N4888, N163, N4597);
or OR2 (N4898, N4897, N4719);
nor NOR4 (N4899, N4898, N3943, N2646, N3002);
xor XOR2 (N4900, N4887, N4205);
xor XOR2 (N4901, N4900, N2001);
nand NAND2 (N4902, N4890, N1206);
nand NAND3 (N4903, N4859, N1734, N1513);
and AND2 (N4904, N4895, N9);
or OR4 (N4905, N4896, N2158, N4021, N2645);
or OR3 (N4906, N4893, N2486, N3612);
or OR4 (N4907, N4905, N3001, N14, N379);
nor NOR3 (N4908, N4891, N1996, N4664);
buf BUF1 (N4909, N4907);
or OR4 (N4910, N4909, N1570, N2203, N3433);
not NOT1 (N4911, N4903);
nand NAND2 (N4912, N4910, N2985);
or OR2 (N4913, N4892, N1649);
and AND4 (N4914, N4878, N2952, N1224, N386);
not NOT1 (N4915, N4906);
xor XOR2 (N4916, N4902, N2806);
nor NOR2 (N4917, N4901, N1698);
not NOT1 (N4918, N4916);
xor XOR2 (N4919, N4899, N234);
buf BUF1 (N4920, N4913);
or OR3 (N4921, N4920, N1889, N3265);
or OR4 (N4922, N4912, N796, N1025, N3417);
and AND2 (N4923, N4915, N4845);
and AND4 (N4924, N4911, N3174, N226, N4249);
nand NAND3 (N4925, N4904, N1120, N3020);
nand NAND2 (N4926, N4918, N777);
not NOT1 (N4927, N4919);
not NOT1 (N4928, N4925);
xor XOR2 (N4929, N4928, N797);
not NOT1 (N4930, N4914);
xor XOR2 (N4931, N4929, N2893);
nand NAND2 (N4932, N4921, N3832);
xor XOR2 (N4933, N4917, N767);
and AND4 (N4934, N4930, N4223, N449, N2623);
and AND3 (N4935, N4924, N127, N2243);
or OR3 (N4936, N4927, N1016, N3914);
or OR3 (N4937, N4934, N659, N466);
not NOT1 (N4938, N4935);
nor NOR4 (N4939, N4926, N1946, N3573, N657);
nand NAND3 (N4940, N4931, N2070, N2507);
nor NOR2 (N4941, N4908, N3238);
or OR2 (N4942, N4937, N2990);
or OR2 (N4943, N4936, N2517);
or OR2 (N4944, N4923, N212);
or OR4 (N4945, N4922, N3355, N4810, N3048);
nand NAND4 (N4946, N4944, N2490, N4203, N3932);
or OR3 (N4947, N4945, N4495, N1630);
not NOT1 (N4948, N4940);
buf BUF1 (N4949, N4939);
not NOT1 (N4950, N4942);
buf BUF1 (N4951, N4946);
xor XOR2 (N4952, N4951, N3039);
not NOT1 (N4953, N4948);
nor NOR3 (N4954, N4947, N393, N878);
and AND3 (N4955, N4938, N1590, N1550);
not NOT1 (N4956, N4932);
not NOT1 (N4957, N4954);
not NOT1 (N4958, N4949);
nand NAND4 (N4959, N4941, N718, N288, N3310);
xor XOR2 (N4960, N4952, N1185);
nand NAND3 (N4961, N4933, N1244, N4145);
and AND4 (N4962, N4961, N4136, N3948, N2805);
nor NOR2 (N4963, N4962, N3995);
nand NAND4 (N4964, N4950, N3319, N2935, N4040);
not NOT1 (N4965, N4958);
nor NOR4 (N4966, N4963, N1377, N4542, N3405);
xor XOR2 (N4967, N4960, N4606);
and AND3 (N4968, N4965, N4263, N2622);
or OR3 (N4969, N4955, N1552, N318);
and AND3 (N4970, N4957, N679, N3450);
buf BUF1 (N4971, N4966);
or OR3 (N4972, N4968, N4654, N2419);
nand NAND2 (N4973, N4956, N4313);
xor XOR2 (N4974, N4973, N3176);
buf BUF1 (N4975, N4967);
not NOT1 (N4976, N4970);
nand NAND3 (N4977, N4972, N1065, N3007);
xor XOR2 (N4978, N4953, N3538);
and AND2 (N4979, N4971, N3690);
nand NAND4 (N4980, N4943, N1159, N556, N632);
nand NAND2 (N4981, N4974, N4823);
xor XOR2 (N4982, N4977, N4527);
nor NOR3 (N4983, N4980, N2513, N4207);
nand NAND4 (N4984, N4981, N2375, N1252, N1983);
buf BUF1 (N4985, N4976);
or OR4 (N4986, N4979, N1273, N2876, N3201);
and AND4 (N4987, N4984, N4552, N622, N183);
xor XOR2 (N4988, N4975, N2090);
nor NOR3 (N4989, N4988, N1259, N3886);
not NOT1 (N4990, N4986);
xor XOR2 (N4991, N4983, N1418);
xor XOR2 (N4992, N4978, N3825);
and AND4 (N4993, N4964, N4770, N2010, N2329);
not NOT1 (N4994, N4993);
nor NOR4 (N4995, N4991, N3191, N1486, N3762);
and AND2 (N4996, N4995, N89);
nor NOR2 (N4997, N4992, N4853);
nand NAND3 (N4998, N4990, N2518, N4684);
nand NAND3 (N4999, N4994, N1125, N2092);
nor NOR2 (N5000, N4985, N1343);
nor NOR2 (N5001, N4997, N1565);
nor NOR4 (N5002, N5000, N1216, N1182, N3677);
not NOT1 (N5003, N5002);
xor XOR2 (N5004, N4959, N1720);
or OR3 (N5005, N4987, N3506, N4488);
nor NOR2 (N5006, N4999, N406);
nand NAND4 (N5007, N4969, N1625, N3351, N1151);
nand NAND2 (N5008, N5005, N4096);
buf BUF1 (N5009, N5008);
nor NOR2 (N5010, N5003, N461);
nand NAND3 (N5011, N5004, N2757, N3259);
buf BUF1 (N5012, N4996);
not NOT1 (N5013, N5010);
nor NOR2 (N5014, N4989, N3534);
or OR3 (N5015, N5013, N2127, N2129);
buf BUF1 (N5016, N4982);
not NOT1 (N5017, N4998);
or OR3 (N5018, N5016, N4112, N2405);
buf BUF1 (N5019, N5011);
nand NAND4 (N5020, N5006, N4559, N2457, N2925);
not NOT1 (N5021, N5012);
not NOT1 (N5022, N5014);
buf BUF1 (N5023, N5019);
not NOT1 (N5024, N5007);
nor NOR3 (N5025, N5018, N1514, N3782);
not NOT1 (N5026, N5015);
nor NOR4 (N5027, N5017, N3247, N289, N800);
buf BUF1 (N5028, N5001);
nor NOR4 (N5029, N5009, N3579, N3457, N4166);
not NOT1 (N5030, N5025);
nor NOR4 (N5031, N5030, N4233, N4137, N2450);
nand NAND2 (N5032, N5028, N3404);
buf BUF1 (N5033, N5024);
buf BUF1 (N5034, N5023);
xor XOR2 (N5035, N5022, N3876);
or OR4 (N5036, N5032, N4883, N2050, N3893);
not NOT1 (N5037, N5031);
not NOT1 (N5038, N5027);
nand NAND3 (N5039, N5033, N1515, N2847);
buf BUF1 (N5040, N5021);
xor XOR2 (N5041, N5020, N716);
nand NAND2 (N5042, N5040, N4140);
nand NAND2 (N5043, N5026, N85);
nand NAND3 (N5044, N5029, N1004, N4611);
not NOT1 (N5045, N5037);
buf BUF1 (N5046, N5042);
nor NOR4 (N5047, N5041, N1819, N987, N3459);
not NOT1 (N5048, N5036);
xor XOR2 (N5049, N5034, N4777);
xor XOR2 (N5050, N5043, N274);
and AND4 (N5051, N5050, N4330, N1482, N584);
buf BUF1 (N5052, N5047);
and AND3 (N5053, N5049, N5035, N4058);
xor XOR2 (N5054, N4311, N4362);
not NOT1 (N5055, N5039);
buf BUF1 (N5056, N5051);
and AND4 (N5057, N5054, N4048, N3569, N1060);
and AND3 (N5058, N5053, N4746, N1189);
not NOT1 (N5059, N5057);
and AND2 (N5060, N5044, N142);
nor NOR3 (N5061, N5038, N4506, N3134);
and AND2 (N5062, N5058, N1049);
or OR3 (N5063, N5062, N1453, N3287);
or OR3 (N5064, N5048, N1581, N1813);
and AND3 (N5065, N5056, N3429, N1603);
and AND3 (N5066, N5059, N2263, N2633);
not NOT1 (N5067, N5045);
xor XOR2 (N5068, N5063, N990);
buf BUF1 (N5069, N5055);
xor XOR2 (N5070, N5067, N2550);
nand NAND4 (N5071, N5065, N1663, N4086, N908);
nand NAND2 (N5072, N5060, N699);
xor XOR2 (N5073, N5071, N4153);
nor NOR4 (N5074, N5069, N3998, N3881, N3157);
nand NAND2 (N5075, N5070, N2526);
or OR3 (N5076, N5074, N683, N681);
not NOT1 (N5077, N5064);
nand NAND4 (N5078, N5061, N1050, N1137, N1136);
not NOT1 (N5079, N5046);
nor NOR2 (N5080, N5077, N3529);
or OR2 (N5081, N5078, N337);
nor NOR4 (N5082, N5076, N3056, N5071, N242);
or OR3 (N5083, N5066, N4308, N4794);
not NOT1 (N5084, N5068);
nand NAND3 (N5085, N5084, N3362, N3082);
not NOT1 (N5086, N5072);
and AND2 (N5087, N5052, N3369);
buf BUF1 (N5088, N5080);
nand NAND2 (N5089, N5088, N3139);
and AND2 (N5090, N5089, N4878);
or OR3 (N5091, N5087, N3960, N715);
nand NAND4 (N5092, N5090, N215, N3654, N3837);
nand NAND4 (N5093, N5073, N1300, N4552, N379);
nand NAND3 (N5094, N5075, N2827, N3216);
nor NOR3 (N5095, N5094, N836, N1745);
and AND2 (N5096, N5086, N996);
and AND2 (N5097, N5079, N1809);
nor NOR2 (N5098, N5092, N2984);
or OR4 (N5099, N5097, N2639, N2582, N1005);
nor NOR3 (N5100, N5081, N35, N2474);
nor NOR2 (N5101, N5095, N4491);
or OR4 (N5102, N5091, N32, N1570, N955);
nand NAND4 (N5103, N5093, N158, N3382, N4311);
buf BUF1 (N5104, N5098);
and AND3 (N5105, N5082, N3861, N62);
xor XOR2 (N5106, N5085, N2279);
not NOT1 (N5107, N5099);
nor NOR4 (N5108, N5102, N1836, N907, N3942);
or OR4 (N5109, N5107, N5020, N3126, N2695);
or OR4 (N5110, N5105, N3163, N1326, N732);
not NOT1 (N5111, N5103);
nor NOR2 (N5112, N5100, N4254);
nand NAND2 (N5113, N5096, N3677);
or OR4 (N5114, N5106, N1958, N3326, N1390);
or OR2 (N5115, N5108, N4612);
not NOT1 (N5116, N5111);
not NOT1 (N5117, N5109);
buf BUF1 (N5118, N5104);
or OR4 (N5119, N5117, N3045, N3809, N1704);
nor NOR2 (N5120, N5115, N3818);
nand NAND2 (N5121, N5118, N1768);
nor NOR4 (N5122, N5114, N128, N4681, N2845);
buf BUF1 (N5123, N5101);
buf BUF1 (N5124, N5121);
not NOT1 (N5125, N5110);
xor XOR2 (N5126, N5125, N3220);
not NOT1 (N5127, N5119);
xor XOR2 (N5128, N5124, N1777);
nand NAND2 (N5129, N5116, N990);
nand NAND4 (N5130, N5083, N5102, N3001, N4802);
and AND2 (N5131, N5122, N676);
not NOT1 (N5132, N5123);
buf BUF1 (N5133, N5112);
and AND2 (N5134, N5130, N3831);
not NOT1 (N5135, N5120);
nand NAND2 (N5136, N5131, N4046);
and AND4 (N5137, N5126, N2329, N4222, N1285);
and AND3 (N5138, N5113, N2457, N4019);
not NOT1 (N5139, N5137);
nor NOR4 (N5140, N5139, N4202, N5107, N2484);
nand NAND3 (N5141, N5140, N1211, N3955);
not NOT1 (N5142, N5134);
buf BUF1 (N5143, N5127);
nand NAND3 (N5144, N5142, N1886, N5060);
xor XOR2 (N5145, N5129, N1033);
nand NAND3 (N5146, N5136, N4742, N3448);
not NOT1 (N5147, N5138);
not NOT1 (N5148, N5143);
and AND4 (N5149, N5148, N1840, N3593, N1288);
xor XOR2 (N5150, N5145, N4953);
buf BUF1 (N5151, N5149);
or OR2 (N5152, N5141, N1010);
not NOT1 (N5153, N5151);
buf BUF1 (N5154, N5146);
nand NAND2 (N5155, N5128, N4314);
nand NAND4 (N5156, N5150, N4823, N3254, N2062);
buf BUF1 (N5157, N5153);
and AND2 (N5158, N5156, N951);
and AND2 (N5159, N5157, N2386);
nand NAND4 (N5160, N5135, N1843, N4983, N2237);
buf BUF1 (N5161, N5158);
and AND3 (N5162, N5160, N3574, N326);
xor XOR2 (N5163, N5159, N2769);
nand NAND4 (N5164, N5133, N3376, N3967, N2166);
and AND3 (N5165, N5152, N1614, N5124);
buf BUF1 (N5166, N5165);
nor NOR2 (N5167, N5161, N3307);
nand NAND2 (N5168, N5162, N1959);
xor XOR2 (N5169, N5163, N618);
and AND2 (N5170, N5144, N3329);
and AND2 (N5171, N5166, N2486);
or OR2 (N5172, N5170, N3786);
not NOT1 (N5173, N5164);
not NOT1 (N5174, N5154);
nand NAND4 (N5175, N5173, N3417, N3373, N545);
not NOT1 (N5176, N5171);
xor XOR2 (N5177, N5155, N3445);
buf BUF1 (N5178, N5147);
xor XOR2 (N5179, N5175, N3442);
or OR2 (N5180, N5172, N3402);
buf BUF1 (N5181, N5132);
buf BUF1 (N5182, N5181);
xor XOR2 (N5183, N5176, N4986);
and AND3 (N5184, N5168, N2546, N4061);
and AND4 (N5185, N5184, N390, N486, N3527);
nor NOR3 (N5186, N5174, N4789, N2843);
nand NAND3 (N5187, N5179, N3076, N3939);
not NOT1 (N5188, N5183);
buf BUF1 (N5189, N5167);
not NOT1 (N5190, N5188);
nor NOR2 (N5191, N5189, N3418);
buf BUF1 (N5192, N5177);
nor NOR4 (N5193, N5190, N901, N2803, N724);
or OR3 (N5194, N5178, N1281, N1268);
nor NOR2 (N5195, N5180, N2587);
xor XOR2 (N5196, N5186, N3253);
and AND3 (N5197, N5187, N1222, N3439);
buf BUF1 (N5198, N5191);
buf BUF1 (N5199, N5182);
not NOT1 (N5200, N5193);
or OR4 (N5201, N5196, N4066, N3011, N4517);
or OR4 (N5202, N5195, N1737, N1357, N2338);
nand NAND4 (N5203, N5169, N818, N2413, N3002);
not NOT1 (N5204, N5202);
and AND4 (N5205, N5197, N1741, N5185, N981);
buf BUF1 (N5206, N1608);
or OR2 (N5207, N5205, N1429);
or OR4 (N5208, N5203, N1415, N188, N211);
nand NAND3 (N5209, N5199, N3912, N244);
or OR3 (N5210, N5198, N4801, N3793);
buf BUF1 (N5211, N5208);
nor NOR3 (N5212, N5194, N471, N1788);
and AND4 (N5213, N5211, N420, N2826, N2920);
nand NAND3 (N5214, N5204, N460, N1104);
nand NAND3 (N5215, N5209, N1797, N1018);
not NOT1 (N5216, N5213);
buf BUF1 (N5217, N5201);
buf BUF1 (N5218, N5206);
or OR2 (N5219, N5192, N4112);
nor NOR2 (N5220, N5219, N2444);
not NOT1 (N5221, N5216);
nand NAND4 (N5222, N5217, N2733, N2334, N1564);
and AND4 (N5223, N5215, N4623, N2659, N1139);
or OR4 (N5224, N5223, N2029, N5138, N2531);
nor NOR3 (N5225, N5224, N1108, N5176);
xor XOR2 (N5226, N5218, N403);
xor XOR2 (N5227, N5212, N3801);
or OR2 (N5228, N5227, N1848);
xor XOR2 (N5229, N5200, N887);
nand NAND3 (N5230, N5225, N1772, N595);
or OR4 (N5231, N5220, N1515, N623, N698);
not NOT1 (N5232, N5214);
and AND4 (N5233, N5229, N1471, N2096, N2743);
or OR2 (N5234, N5230, N3557);
buf BUF1 (N5235, N5234);
buf BUF1 (N5236, N5222);
xor XOR2 (N5237, N5232, N2302);
xor XOR2 (N5238, N5226, N2015);
xor XOR2 (N5239, N5221, N4432);
xor XOR2 (N5240, N5235, N1287);
not NOT1 (N5241, N5240);
xor XOR2 (N5242, N5238, N1148);
nor NOR4 (N5243, N5207, N3585, N4236, N3096);
not NOT1 (N5244, N5228);
nand NAND2 (N5245, N5241, N4283);
nor NOR2 (N5246, N5239, N4027);
not NOT1 (N5247, N5231);
not NOT1 (N5248, N5244);
nor NOR2 (N5249, N5233, N4272);
or OR4 (N5250, N5249, N3561, N2856, N136);
buf BUF1 (N5251, N5247);
nand NAND2 (N5252, N5237, N4984);
xor XOR2 (N5253, N5250, N2189);
xor XOR2 (N5254, N5243, N1326);
nand NAND2 (N5255, N5253, N3558);
not NOT1 (N5256, N5248);
nor NOR2 (N5257, N5252, N3257);
nor NOR2 (N5258, N5251, N2531);
not NOT1 (N5259, N5246);
nor NOR4 (N5260, N5210, N3188, N617, N3540);
not NOT1 (N5261, N5256);
or OR4 (N5262, N5245, N2604, N563, N3880);
and AND2 (N5263, N5259, N1137);
and AND3 (N5264, N5257, N2204, N3026);
and AND2 (N5265, N5262, N3538);
xor XOR2 (N5266, N5261, N4266);
nor NOR3 (N5267, N5236, N1332, N1792);
and AND3 (N5268, N5264, N2043, N4518);
nand NAND3 (N5269, N5267, N5245, N1533);
nand NAND4 (N5270, N5269, N1277, N1859, N4639);
and AND3 (N5271, N5263, N5105, N2096);
nor NOR2 (N5272, N5255, N3220);
or OR4 (N5273, N5268, N2659, N376, N171);
nor NOR3 (N5274, N5265, N2363, N4483);
xor XOR2 (N5275, N5270, N1855);
not NOT1 (N5276, N5258);
nor NOR3 (N5277, N5272, N3033, N3168);
xor XOR2 (N5278, N5273, N2738);
nand NAND2 (N5279, N5260, N3533);
xor XOR2 (N5280, N5278, N857);
not NOT1 (N5281, N5275);
buf BUF1 (N5282, N5281);
and AND3 (N5283, N5254, N2788, N4362);
buf BUF1 (N5284, N5280);
and AND4 (N5285, N5274, N1113, N493, N2494);
or OR4 (N5286, N5271, N559, N4440, N3918);
not NOT1 (N5287, N5279);
nand NAND3 (N5288, N5282, N89, N3294);
and AND2 (N5289, N5287, N2990);
and AND4 (N5290, N5289, N4069, N4578, N1153);
xor XOR2 (N5291, N5283, N2197);
nand NAND3 (N5292, N5286, N5085, N3924);
and AND4 (N5293, N5285, N3791, N2045, N361);
and AND4 (N5294, N5293, N765, N2221, N4375);
nor NOR2 (N5295, N5290, N2698);
and AND2 (N5296, N5294, N630);
nor NOR4 (N5297, N5296, N1274, N1245, N3378);
xor XOR2 (N5298, N5242, N796);
nand NAND3 (N5299, N5291, N3059, N3798);
xor XOR2 (N5300, N5288, N3748);
not NOT1 (N5301, N5292);
nor NOR3 (N5302, N5284, N2849, N2194);
nor NOR3 (N5303, N5295, N318, N2999);
and AND4 (N5304, N5303, N4886, N2409, N1949);
and AND3 (N5305, N5304, N3936, N929);
buf BUF1 (N5306, N5298);
xor XOR2 (N5307, N5297, N2905);
nor NOR3 (N5308, N5277, N3259, N5260);
and AND4 (N5309, N5307, N148, N2184, N3742);
nand NAND4 (N5310, N5309, N4483, N4006, N4453);
not NOT1 (N5311, N5276);
buf BUF1 (N5312, N5308);
and AND2 (N5313, N5306, N2758);
nor NOR4 (N5314, N5302, N2981, N4747, N2406);
nor NOR2 (N5315, N5312, N572);
not NOT1 (N5316, N5299);
nor NOR4 (N5317, N5311, N5194, N4441, N3227);
or OR2 (N5318, N5315, N2001);
nand NAND4 (N5319, N5314, N3808, N1642, N1949);
or OR2 (N5320, N5319, N1166);
nand NAND3 (N5321, N5301, N5217, N1043);
and AND4 (N5322, N5318, N1941, N663, N1765);
nand NAND3 (N5323, N5317, N1442, N510);
nor NOR3 (N5324, N5313, N731, N3722);
buf BUF1 (N5325, N5316);
and AND4 (N5326, N5300, N690, N3724, N2133);
not NOT1 (N5327, N5322);
xor XOR2 (N5328, N5310, N1894);
xor XOR2 (N5329, N5328, N2721);
nand NAND3 (N5330, N5326, N2178, N132);
xor XOR2 (N5331, N5320, N4214);
nand NAND4 (N5332, N5325, N1927, N2165, N2600);
not NOT1 (N5333, N5323);
xor XOR2 (N5334, N5331, N272);
nand NAND3 (N5335, N5266, N4865, N4564);
not NOT1 (N5336, N5329);
not NOT1 (N5337, N5336);
buf BUF1 (N5338, N5321);
and AND4 (N5339, N5337, N3206, N4381, N2815);
nor NOR3 (N5340, N5334, N885, N6);
nand NAND2 (N5341, N5335, N2423);
buf BUF1 (N5342, N5324);
or OR4 (N5343, N5339, N4358, N2804, N1993);
and AND3 (N5344, N5343, N3566, N3850);
not NOT1 (N5345, N5305);
nand NAND3 (N5346, N5333, N5220, N2044);
xor XOR2 (N5347, N5345, N4790);
nor NOR2 (N5348, N5342, N650);
and AND4 (N5349, N5347, N3101, N4381, N4650);
buf BUF1 (N5350, N5341);
xor XOR2 (N5351, N5338, N5333);
nand NAND4 (N5352, N5350, N1948, N4937, N3217);
or OR4 (N5353, N5348, N1175, N3656, N1497);
buf BUF1 (N5354, N5351);
not NOT1 (N5355, N5354);
buf BUF1 (N5356, N5340);
nand NAND3 (N5357, N5355, N1947, N3085);
not NOT1 (N5358, N5327);
nor NOR4 (N5359, N5357, N3029, N505, N4896);
buf BUF1 (N5360, N5353);
xor XOR2 (N5361, N5359, N939);
or OR4 (N5362, N5346, N3882, N3334, N3888);
nand NAND4 (N5363, N5349, N2331, N4519, N372);
or OR4 (N5364, N5356, N5082, N1902, N3668);
or OR2 (N5365, N5330, N1756);
and AND2 (N5366, N5362, N5081);
xor XOR2 (N5367, N5360, N2684);
or OR2 (N5368, N5366, N1980);
not NOT1 (N5369, N5365);
not NOT1 (N5370, N5364);
nand NAND2 (N5371, N5332, N5337);
buf BUF1 (N5372, N5352);
nor NOR4 (N5373, N5363, N2833, N5182, N3081);
nor NOR3 (N5374, N5369, N4281, N990);
xor XOR2 (N5375, N5373, N3036);
buf BUF1 (N5376, N5370);
or OR2 (N5377, N5344, N4811);
nor NOR2 (N5378, N5368, N590);
buf BUF1 (N5379, N5378);
not NOT1 (N5380, N5375);
xor XOR2 (N5381, N5379, N1979);
not NOT1 (N5382, N5371);
xor XOR2 (N5383, N5372, N3123);
buf BUF1 (N5384, N5377);
buf BUF1 (N5385, N5358);
nor NOR2 (N5386, N5361, N1009);
xor XOR2 (N5387, N5384, N2487);
or OR4 (N5388, N5374, N613, N3856, N3925);
buf BUF1 (N5389, N5388);
nand NAND4 (N5390, N5385, N4282, N3928, N4012);
xor XOR2 (N5391, N5383, N2860);
not NOT1 (N5392, N5390);
xor XOR2 (N5393, N5391, N1311);
or OR4 (N5394, N5393, N1771, N1577, N4483);
nand NAND2 (N5395, N5367, N2985);
not NOT1 (N5396, N5387);
not NOT1 (N5397, N5389);
xor XOR2 (N5398, N5382, N1720);
not NOT1 (N5399, N5398);
nor NOR4 (N5400, N5386, N3539, N1857, N293);
xor XOR2 (N5401, N5396, N58);
and AND3 (N5402, N5400, N3828, N3986);
xor XOR2 (N5403, N5401, N4265);
xor XOR2 (N5404, N5402, N1321);
buf BUF1 (N5405, N5399);
and AND4 (N5406, N5403, N5064, N1834, N5371);
nor NOR3 (N5407, N5404, N5168, N1762);
nand NAND2 (N5408, N5405, N4671);
or OR3 (N5409, N5376, N1837, N2918);
buf BUF1 (N5410, N5394);
buf BUF1 (N5411, N5381);
nand NAND3 (N5412, N5410, N5151, N1088);
buf BUF1 (N5413, N5411);
nor NOR3 (N5414, N5408, N674, N1575);
or OR4 (N5415, N5413, N5406, N4992, N3973);
nor NOR3 (N5416, N1784, N4958, N2770);
not NOT1 (N5417, N5414);
or OR4 (N5418, N5397, N2271, N1415, N2195);
nand NAND4 (N5419, N5409, N3547, N1789, N2937);
nor NOR2 (N5420, N5419, N2738);
buf BUF1 (N5421, N5392);
or OR3 (N5422, N5420, N2869, N1149);
xor XOR2 (N5423, N5422, N4650);
nor NOR2 (N5424, N5380, N5411);
nor NOR3 (N5425, N5418, N3088, N1557);
nand NAND2 (N5426, N5425, N2397);
nor NOR3 (N5427, N5416, N2870, N2763);
buf BUF1 (N5428, N5407);
and AND3 (N5429, N5412, N789, N1580);
not NOT1 (N5430, N5426);
not NOT1 (N5431, N5430);
or OR2 (N5432, N5395, N4603);
not NOT1 (N5433, N5415);
and AND2 (N5434, N5429, N4824);
nand NAND3 (N5435, N5434, N3002, N3332);
nand NAND2 (N5436, N5424, N3457);
xor XOR2 (N5437, N5428, N1590);
nor NOR3 (N5438, N5423, N1043, N887);
and AND4 (N5439, N5436, N3108, N2680, N1085);
nor NOR4 (N5440, N5439, N2426, N2153, N2785);
and AND2 (N5441, N5435, N2866);
xor XOR2 (N5442, N5417, N771);
nor NOR4 (N5443, N5442, N3117, N1954, N3047);
or OR3 (N5444, N5438, N924, N4768);
and AND2 (N5445, N5441, N5044);
nor NOR2 (N5446, N5445, N1584);
not NOT1 (N5447, N5437);
and AND4 (N5448, N5427, N2497, N1115, N3040);
or OR3 (N5449, N5421, N1760, N3382);
buf BUF1 (N5450, N5443);
not NOT1 (N5451, N5444);
or OR4 (N5452, N5433, N4141, N3257, N3530);
buf BUF1 (N5453, N5432);
nor NOR4 (N5454, N5448, N2083, N3963, N1200);
nor NOR4 (N5455, N5454, N902, N1655, N4068);
or OR3 (N5456, N5451, N2132, N332);
or OR4 (N5457, N5456, N2244, N1160, N1102);
nand NAND3 (N5458, N5457, N2525, N4398);
not NOT1 (N5459, N5447);
or OR3 (N5460, N5458, N5041, N3721);
not NOT1 (N5461, N5452);
and AND3 (N5462, N5459, N2061, N4836);
not NOT1 (N5463, N5453);
xor XOR2 (N5464, N5449, N4450);
nor NOR4 (N5465, N5450, N1909, N3258, N534);
or OR4 (N5466, N5431, N3519, N2634, N3125);
nor NOR4 (N5467, N5461, N5110, N5, N4901);
buf BUF1 (N5468, N5440);
nor NOR2 (N5469, N5446, N4952);
not NOT1 (N5470, N5465);
nor NOR3 (N5471, N5467, N4641, N3878);
nand NAND4 (N5472, N5460, N5123, N4812, N4424);
buf BUF1 (N5473, N5464);
nor NOR3 (N5474, N5473, N3840, N2148);
not NOT1 (N5475, N5474);
nand NAND2 (N5476, N5469, N4720);
and AND3 (N5477, N5472, N5290, N4931);
or OR3 (N5478, N5477, N3871, N957);
and AND3 (N5479, N5470, N997, N3837);
not NOT1 (N5480, N5455);
or OR4 (N5481, N5478, N2991, N4033, N1026);
xor XOR2 (N5482, N5481, N2507);
nor NOR2 (N5483, N5462, N460);
not NOT1 (N5484, N5479);
nor NOR2 (N5485, N5466, N2287);
nor NOR4 (N5486, N5468, N992, N1258, N1435);
and AND3 (N5487, N5480, N2225, N2947);
xor XOR2 (N5488, N5483, N2596);
and AND4 (N5489, N5463, N1968, N320, N4043);
xor XOR2 (N5490, N5488, N2022);
buf BUF1 (N5491, N5482);
xor XOR2 (N5492, N5471, N3816);
or OR3 (N5493, N5486, N4332, N2603);
nor NOR3 (N5494, N5487, N1476, N149);
nand NAND3 (N5495, N5493, N1524, N3490);
xor XOR2 (N5496, N5489, N3147);
nand NAND2 (N5497, N5496, N380);
buf BUF1 (N5498, N5497);
not NOT1 (N5499, N5491);
or OR2 (N5500, N5484, N1622);
buf BUF1 (N5501, N5500);
buf BUF1 (N5502, N5485);
or OR2 (N5503, N5498, N959);
and AND2 (N5504, N5494, N3079);
and AND2 (N5505, N5502, N4837);
buf BUF1 (N5506, N5501);
xor XOR2 (N5507, N5492, N4260);
and AND4 (N5508, N5507, N3145, N3117, N426);
buf BUF1 (N5509, N5505);
nand NAND3 (N5510, N5503, N2627, N203);
and AND2 (N5511, N5504, N1768);
nor NOR2 (N5512, N5499, N2419);
and AND4 (N5513, N5476, N3593, N3998, N511);
or OR3 (N5514, N5490, N4911, N1648);
nand NAND3 (N5515, N5510, N1830, N569);
or OR4 (N5516, N5511, N5086, N4321, N902);
or OR4 (N5517, N5506, N1149, N2767, N2663);
buf BUF1 (N5518, N5509);
and AND3 (N5519, N5515, N2296, N3342);
not NOT1 (N5520, N5513);
not NOT1 (N5521, N5512);
nor NOR2 (N5522, N5520, N560);
nand NAND2 (N5523, N5518, N5362);
or OR2 (N5524, N5521, N3143);
nor NOR2 (N5525, N5495, N4378);
buf BUF1 (N5526, N5524);
and AND4 (N5527, N5508, N1375, N3097, N2014);
or OR3 (N5528, N5525, N3445, N85);
buf BUF1 (N5529, N5526);
and AND2 (N5530, N5517, N1144);
xor XOR2 (N5531, N5514, N1846);
not NOT1 (N5532, N5522);
and AND4 (N5533, N5528, N5401, N1302, N1223);
and AND3 (N5534, N5516, N251, N3343);
or OR4 (N5535, N5533, N941, N4091, N3462);
and AND4 (N5536, N5475, N1524, N2627, N4617);
xor XOR2 (N5537, N5519, N410);
nor NOR4 (N5538, N5537, N3173, N750, N241);
nor NOR3 (N5539, N5538, N2682, N2473);
nor NOR4 (N5540, N5535, N3355, N4542, N5226);
not NOT1 (N5541, N5527);
not NOT1 (N5542, N5529);
buf BUF1 (N5543, N5534);
or OR4 (N5544, N5530, N2107, N1593, N3844);
buf BUF1 (N5545, N5523);
and AND2 (N5546, N5542, N1609);
or OR3 (N5547, N5543, N1838, N5529);
xor XOR2 (N5548, N5546, N2925);
xor XOR2 (N5549, N5541, N179);
xor XOR2 (N5550, N5545, N1575);
nor NOR4 (N5551, N5544, N5521, N3348, N1172);
xor XOR2 (N5552, N5547, N628);
xor XOR2 (N5553, N5531, N2253);
buf BUF1 (N5554, N5540);
not NOT1 (N5555, N5548);
xor XOR2 (N5556, N5553, N2469);
xor XOR2 (N5557, N5536, N1836);
not NOT1 (N5558, N5555);
xor XOR2 (N5559, N5539, N3054);
nor NOR4 (N5560, N5557, N3935, N2740, N5411);
nand NAND3 (N5561, N5556, N1228, N5548);
buf BUF1 (N5562, N5532);
buf BUF1 (N5563, N5549);
xor XOR2 (N5564, N5562, N5553);
and AND2 (N5565, N5551, N3135);
buf BUF1 (N5566, N5564);
not NOT1 (N5567, N5565);
and AND3 (N5568, N5558, N2417, N1898);
nor NOR2 (N5569, N5561, N1558);
and AND2 (N5570, N5560, N4269);
and AND4 (N5571, N5554, N814, N1837, N5040);
nor NOR2 (N5572, N5569, N1203);
nand NAND3 (N5573, N5571, N2291, N2439);
not NOT1 (N5574, N5552);
nand NAND4 (N5575, N5566, N2109, N2719, N4326);
buf BUF1 (N5576, N5573);
buf BUF1 (N5577, N5567);
xor XOR2 (N5578, N5563, N568);
not NOT1 (N5579, N5574);
nor NOR4 (N5580, N5559, N2240, N4226, N3940);
nor NOR3 (N5581, N5580, N5413, N5125);
nor NOR4 (N5582, N5576, N656, N3862, N727);
not NOT1 (N5583, N5550);
nand NAND2 (N5584, N5577, N4314);
buf BUF1 (N5585, N5572);
or OR2 (N5586, N5585, N3881);
nand NAND2 (N5587, N5582, N951);
buf BUF1 (N5588, N5583);
nor NOR2 (N5589, N5586, N5353);
or OR4 (N5590, N5587, N2929, N2489, N4982);
or OR3 (N5591, N5589, N968, N4019);
not NOT1 (N5592, N5570);
not NOT1 (N5593, N5592);
nor NOR3 (N5594, N5575, N2430, N5096);
xor XOR2 (N5595, N5568, N1324);
and AND2 (N5596, N5591, N2093);
nor NOR3 (N5597, N5596, N2084, N5360);
or OR4 (N5598, N5594, N4000, N1974, N1341);
and AND4 (N5599, N5598, N3564, N1129, N227);
or OR2 (N5600, N5593, N3662);
and AND2 (N5601, N5588, N3950);
buf BUF1 (N5602, N5599);
nor NOR2 (N5603, N5584, N3790);
nor NOR3 (N5604, N5595, N1360, N4196);
nand NAND3 (N5605, N5590, N2, N519);
xor XOR2 (N5606, N5581, N2899);
or OR3 (N5607, N5578, N5156, N4316);
or OR3 (N5608, N5607, N2536, N2038);
not NOT1 (N5609, N5605);
xor XOR2 (N5610, N5601, N3992);
buf BUF1 (N5611, N5610);
or OR4 (N5612, N5600, N3198, N3440, N2748);
and AND4 (N5613, N5606, N481, N4210, N288);
xor XOR2 (N5614, N5609, N3719);
nor NOR4 (N5615, N5603, N5471, N4257, N3685);
nor NOR4 (N5616, N5613, N1599, N3479, N5202);
nand NAND2 (N5617, N5597, N4192);
and AND3 (N5618, N5617, N5295, N778);
buf BUF1 (N5619, N5614);
buf BUF1 (N5620, N5615);
xor XOR2 (N5621, N5616, N3583);
and AND3 (N5622, N5608, N5007, N5164);
and AND3 (N5623, N5620, N3198, N1445);
buf BUF1 (N5624, N5622);
buf BUF1 (N5625, N5619);
nor NOR4 (N5626, N5579, N3763, N5183, N221);
buf BUF1 (N5627, N5602);
nor NOR3 (N5628, N5627, N721, N3128);
or OR3 (N5629, N5604, N1636, N4620);
not NOT1 (N5630, N5612);
and AND4 (N5631, N5628, N868, N3508, N3662);
or OR3 (N5632, N5630, N3997, N3435);
buf BUF1 (N5633, N5631);
xor XOR2 (N5634, N5611, N3198);
and AND4 (N5635, N5623, N3937, N1601, N3757);
not NOT1 (N5636, N5624);
xor XOR2 (N5637, N5636, N3576);
xor XOR2 (N5638, N5626, N3632);
nand NAND4 (N5639, N5618, N1269, N4105, N4621);
or OR2 (N5640, N5625, N3282);
and AND3 (N5641, N5640, N2654, N242);
or OR2 (N5642, N5641, N4985);
xor XOR2 (N5643, N5632, N236);
not NOT1 (N5644, N5629);
nor NOR4 (N5645, N5638, N2197, N1047, N3097);
xor XOR2 (N5646, N5644, N2727);
nor NOR4 (N5647, N5633, N5618, N2211, N3108);
xor XOR2 (N5648, N5639, N1344);
not NOT1 (N5649, N5648);
nor NOR4 (N5650, N5649, N1172, N2391, N1115);
nand NAND3 (N5651, N5643, N418, N4811);
nor NOR4 (N5652, N5634, N182, N738, N4635);
nand NAND4 (N5653, N5621, N235, N3097, N823);
and AND3 (N5654, N5650, N1061, N2584);
not NOT1 (N5655, N5651);
nand NAND2 (N5656, N5635, N2058);
xor XOR2 (N5657, N5654, N4693);
or OR3 (N5658, N5646, N5563, N1862);
not NOT1 (N5659, N5656);
nor NOR2 (N5660, N5659, N3885);
nor NOR2 (N5661, N5655, N2144);
or OR4 (N5662, N5642, N1348, N4743, N3187);
xor XOR2 (N5663, N5661, N5183);
not NOT1 (N5664, N5653);
not NOT1 (N5665, N5652);
nor NOR4 (N5666, N5657, N201, N2129, N5591);
buf BUF1 (N5667, N5637);
and AND4 (N5668, N5663, N3300, N5564, N2894);
nand NAND4 (N5669, N5668, N2037, N4243, N493);
nor NOR3 (N5670, N5660, N4930, N2457);
nand NAND3 (N5671, N5670, N4816, N3027);
nand NAND3 (N5672, N5662, N341, N3622);
nand NAND2 (N5673, N5645, N5608);
and AND4 (N5674, N5664, N1436, N3775, N1837);
xor XOR2 (N5675, N5672, N1181);
xor XOR2 (N5676, N5666, N5295);
not NOT1 (N5677, N5647);
not NOT1 (N5678, N5667);
buf BUF1 (N5679, N5676);
or OR4 (N5680, N5671, N2563, N3829, N1705);
not NOT1 (N5681, N5658);
nand NAND2 (N5682, N5674, N4120);
xor XOR2 (N5683, N5678, N2223);
or OR3 (N5684, N5677, N4064, N497);
nand NAND3 (N5685, N5683, N4721, N3012);
nand NAND3 (N5686, N5685, N1282, N5029);
nor NOR4 (N5687, N5673, N2477, N2399, N1510);
and AND4 (N5688, N5687, N2323, N4739, N1418);
buf BUF1 (N5689, N5665);
and AND2 (N5690, N5675, N1103);
xor XOR2 (N5691, N5669, N93);
or OR4 (N5692, N5682, N3895, N3411, N1766);
nand NAND3 (N5693, N5690, N4480, N34);
or OR3 (N5694, N5681, N3901, N225);
nor NOR4 (N5695, N5688, N5454, N1868, N428);
or OR3 (N5696, N5693, N2041, N760);
or OR2 (N5697, N5691, N1979);
and AND4 (N5698, N5694, N4495, N942, N1802);
buf BUF1 (N5699, N5698);
not NOT1 (N5700, N5692);
nand NAND3 (N5701, N5684, N3583, N2799);
buf BUF1 (N5702, N5689);
nand NAND3 (N5703, N5679, N419, N1356);
or OR4 (N5704, N5696, N4448, N4850, N4257);
and AND4 (N5705, N5703, N2722, N1239, N3838);
xor XOR2 (N5706, N5701, N1024);
nor NOR2 (N5707, N5680, N1715);
xor XOR2 (N5708, N5700, N1709);
nor NOR4 (N5709, N5695, N5173, N1273, N4633);
or OR4 (N5710, N5702, N5661, N3817, N841);
xor XOR2 (N5711, N5710, N3163);
nor NOR3 (N5712, N5708, N3158, N3848);
nor NOR4 (N5713, N5712, N963, N5244, N4861);
not NOT1 (N5714, N5711);
nor NOR4 (N5715, N5686, N4386, N2466, N5556);
nor NOR2 (N5716, N5699, N2087);
buf BUF1 (N5717, N5713);
not NOT1 (N5718, N5714);
not NOT1 (N5719, N5717);
nand NAND2 (N5720, N5705, N521);
nor NOR3 (N5721, N5709, N1401, N3156);
nor NOR2 (N5722, N5704, N1035);
nor NOR4 (N5723, N5722, N3305, N2195, N1219);
not NOT1 (N5724, N5715);
or OR4 (N5725, N5706, N5698, N5451, N1665);
buf BUF1 (N5726, N5720);
xor XOR2 (N5727, N5707, N4857);
nor NOR2 (N5728, N5724, N738);
or OR3 (N5729, N5719, N752, N5092);
nand NAND2 (N5730, N5726, N782);
not NOT1 (N5731, N5728);
or OR4 (N5732, N5723, N4591, N950, N1080);
nand NAND3 (N5733, N5727, N5462, N382);
xor XOR2 (N5734, N5730, N729);
nand NAND4 (N5735, N5718, N4519, N3647, N3636);
nand NAND4 (N5736, N5733, N5469, N3730, N1595);
not NOT1 (N5737, N5731);
nor NOR4 (N5738, N5736, N4153, N1909, N5448);
and AND3 (N5739, N5716, N1681, N5497);
xor XOR2 (N5740, N5732, N677);
or OR3 (N5741, N5738, N4036, N3091);
xor XOR2 (N5742, N5741, N5146);
nor NOR3 (N5743, N5739, N2809, N1325);
buf BUF1 (N5744, N5743);
or OR4 (N5745, N5734, N5450, N5552, N548);
xor XOR2 (N5746, N5735, N4107);
and AND4 (N5747, N5746, N2598, N1009, N2824);
or OR4 (N5748, N5745, N2578, N1123, N5325);
buf BUF1 (N5749, N5747);
xor XOR2 (N5750, N5725, N5071);
not NOT1 (N5751, N5749);
buf BUF1 (N5752, N5751);
nor NOR2 (N5753, N5729, N3234);
nor NOR3 (N5754, N5753, N1730, N35);
nand NAND4 (N5755, N5752, N4190, N436, N5363);
buf BUF1 (N5756, N5740);
buf BUF1 (N5757, N5742);
or OR4 (N5758, N5754, N946, N5273, N4539);
and AND4 (N5759, N5757, N3838, N3232, N5486);
not NOT1 (N5760, N5758);
nand NAND3 (N5761, N5721, N4796, N1083);
buf BUF1 (N5762, N5759);
buf BUF1 (N5763, N5760);
nor NOR4 (N5764, N5697, N2793, N5458, N5430);
and AND2 (N5765, N5762, N3383);
not NOT1 (N5766, N5765);
xor XOR2 (N5767, N5748, N2782);
and AND3 (N5768, N5750, N2059, N624);
and AND2 (N5769, N5768, N3933);
nand NAND2 (N5770, N5763, N2);
and AND2 (N5771, N5764, N2414);
nor NOR2 (N5772, N5755, N5298);
xor XOR2 (N5773, N5766, N5267);
or OR3 (N5774, N5761, N4329, N560);
not NOT1 (N5775, N5773);
and AND2 (N5776, N5767, N3906);
and AND2 (N5777, N5769, N2064);
not NOT1 (N5778, N5744);
xor XOR2 (N5779, N5771, N434);
nor NOR2 (N5780, N5779, N3746);
not NOT1 (N5781, N5780);
nand NAND3 (N5782, N5775, N159, N4813);
and AND3 (N5783, N5770, N1068, N2678);
nor NOR2 (N5784, N5777, N4857);
nand NAND2 (N5785, N5774, N986);
or OR3 (N5786, N5737, N3478, N2789);
and AND2 (N5787, N5782, N4999);
not NOT1 (N5788, N5785);
xor XOR2 (N5789, N5784, N3805);
and AND2 (N5790, N5783, N775);
or OR4 (N5791, N5781, N4042, N3113, N726);
not NOT1 (N5792, N5772);
nand NAND4 (N5793, N5790, N5003, N3762, N861);
buf BUF1 (N5794, N5791);
and AND4 (N5795, N5756, N2660, N2000, N4207);
xor XOR2 (N5796, N5794, N3339);
nand NAND4 (N5797, N5786, N3248, N4728, N2061);
not NOT1 (N5798, N5789);
nand NAND4 (N5799, N5795, N949, N307, N1664);
nor NOR4 (N5800, N5793, N1651, N1937, N4942);
buf BUF1 (N5801, N5776);
nor NOR2 (N5802, N5792, N4358);
and AND2 (N5803, N5787, N4080);
xor XOR2 (N5804, N5778, N3231);
nor NOR4 (N5805, N5803, N4297, N555, N3956);
not NOT1 (N5806, N5802);
xor XOR2 (N5807, N5796, N5201);
and AND4 (N5808, N5799, N2758, N1106, N1135);
not NOT1 (N5809, N5800);
not NOT1 (N5810, N5788);
and AND2 (N5811, N5805, N628);
buf BUF1 (N5812, N5804);
or OR2 (N5813, N5810, N508);
and AND2 (N5814, N5798, N2019);
and AND3 (N5815, N5811, N5243, N3822);
nand NAND3 (N5816, N5815, N3219, N2011);
or OR4 (N5817, N5812, N170, N1981, N2321);
nand NAND2 (N5818, N5807, N3290);
and AND4 (N5819, N5814, N4353, N1043, N709);
xor XOR2 (N5820, N5809, N4950);
buf BUF1 (N5821, N5820);
buf BUF1 (N5822, N5816);
nor NOR3 (N5823, N5806, N3564, N4373);
or OR3 (N5824, N5801, N358, N257);
nand NAND3 (N5825, N5813, N3118, N2571);
not NOT1 (N5826, N5819);
nand NAND4 (N5827, N5823, N4957, N5541, N3911);
nor NOR2 (N5828, N5797, N652);
xor XOR2 (N5829, N5827, N4782);
nor NOR4 (N5830, N5825, N293, N4186, N2568);
and AND4 (N5831, N5821, N3574, N4910, N4707);
nand NAND2 (N5832, N5831, N283);
and AND4 (N5833, N5822, N2533, N4756, N2305);
and AND2 (N5834, N5833, N3206);
or OR4 (N5835, N5824, N1040, N3378, N212);
xor XOR2 (N5836, N5817, N3286);
not NOT1 (N5837, N5829);
nor NOR2 (N5838, N5834, N733);
xor XOR2 (N5839, N5837, N570);
not NOT1 (N5840, N5830);
and AND4 (N5841, N5839, N4044, N457, N5079);
not NOT1 (N5842, N5841);
nor NOR4 (N5843, N5818, N5158, N3437, N81);
nor NOR4 (N5844, N5843, N1080, N2861, N5755);
or OR4 (N5845, N5832, N3965, N3740, N2684);
or OR2 (N5846, N5840, N2427);
xor XOR2 (N5847, N5838, N4603);
xor XOR2 (N5848, N5842, N2350);
and AND2 (N5849, N5808, N3788);
buf BUF1 (N5850, N5845);
or OR2 (N5851, N5848, N5384);
or OR4 (N5852, N5836, N5683, N4021, N5311);
xor XOR2 (N5853, N5852, N3601);
not NOT1 (N5854, N5828);
nand NAND4 (N5855, N5854, N5342, N1150, N4250);
nand NAND2 (N5856, N5847, N3186);
nor NOR2 (N5857, N5853, N177);
buf BUF1 (N5858, N5856);
nand NAND2 (N5859, N5858, N711);
not NOT1 (N5860, N5850);
nand NAND3 (N5861, N5859, N5817, N4068);
or OR2 (N5862, N5851, N1518);
not NOT1 (N5863, N5857);
and AND3 (N5864, N5835, N3303, N5515);
or OR2 (N5865, N5861, N2571);
nand NAND4 (N5866, N5846, N1530, N1813, N3111);
or OR3 (N5867, N5862, N3792, N3245);
xor XOR2 (N5868, N5865, N3895);
and AND4 (N5869, N5860, N3437, N2729, N1117);
xor XOR2 (N5870, N5867, N5220);
nor NOR2 (N5871, N5866, N1975);
xor XOR2 (N5872, N5849, N4306);
buf BUF1 (N5873, N5826);
not NOT1 (N5874, N5863);
xor XOR2 (N5875, N5870, N406);
not NOT1 (N5876, N5869);
nand NAND3 (N5877, N5844, N2022, N5718);
or OR2 (N5878, N5871, N2082);
buf BUF1 (N5879, N5878);
or OR2 (N5880, N5868, N4812);
buf BUF1 (N5881, N5873);
buf BUF1 (N5882, N5874);
not NOT1 (N5883, N5880);
nand NAND3 (N5884, N5879, N1996, N4947);
buf BUF1 (N5885, N5872);
nand NAND3 (N5886, N5864, N1465, N217);
nor NOR4 (N5887, N5875, N2245, N1324, N4980);
not NOT1 (N5888, N5881);
nand NAND3 (N5889, N5886, N5426, N3411);
nor NOR2 (N5890, N5877, N764);
xor XOR2 (N5891, N5885, N2542);
or OR2 (N5892, N5855, N3584);
buf BUF1 (N5893, N5892);
xor XOR2 (N5894, N5890, N4944);
nor NOR4 (N5895, N5889, N5105, N3898, N4080);
not NOT1 (N5896, N5895);
not NOT1 (N5897, N5888);
nor NOR3 (N5898, N5891, N1286, N1759);
buf BUF1 (N5899, N5884);
nor NOR4 (N5900, N5893, N3090, N4667, N4728);
or OR2 (N5901, N5883, N1739);
not NOT1 (N5902, N5896);
or OR2 (N5903, N5900, N4613);
or OR3 (N5904, N5887, N5670, N3806);
and AND2 (N5905, N5902, N1558);
xor XOR2 (N5906, N5905, N3335);
nor NOR3 (N5907, N5897, N3931, N5705);
nand NAND4 (N5908, N5898, N5068, N1418, N2030);
not NOT1 (N5909, N5903);
not NOT1 (N5910, N5906);
nand NAND2 (N5911, N5908, N5314);
and AND3 (N5912, N5907, N3654, N2006);
not NOT1 (N5913, N5910);
nand NAND2 (N5914, N5911, N1353);
buf BUF1 (N5915, N5913);
or OR2 (N5916, N5882, N2279);
nand NAND4 (N5917, N5914, N2150, N2568, N3903);
buf BUF1 (N5918, N5917);
not NOT1 (N5919, N5915);
not NOT1 (N5920, N5899);
or OR4 (N5921, N5904, N1818, N3331, N5112);
or OR3 (N5922, N5876, N5447, N4476);
or OR4 (N5923, N5901, N833, N5603, N542);
and AND4 (N5924, N5894, N5211, N1016, N1435);
not NOT1 (N5925, N5923);
buf BUF1 (N5926, N5922);
or OR3 (N5927, N5924, N1213, N2608);
or OR4 (N5928, N5926, N371, N5744, N3453);
xor XOR2 (N5929, N5919, N3239);
nor NOR2 (N5930, N5927, N2796);
or OR4 (N5931, N5912, N3315, N5209, N1756);
xor XOR2 (N5932, N5916, N963);
xor XOR2 (N5933, N5932, N1846);
or OR3 (N5934, N5918, N4479, N5064);
xor XOR2 (N5935, N5920, N1138);
or OR3 (N5936, N5921, N4778, N3301);
xor XOR2 (N5937, N5931, N3362);
and AND2 (N5938, N5935, N3322);
xor XOR2 (N5939, N5938, N4196);
and AND4 (N5940, N5925, N5771, N1771, N4379);
xor XOR2 (N5941, N5928, N1677);
nand NAND2 (N5942, N5936, N2715);
xor XOR2 (N5943, N5939, N4513);
not NOT1 (N5944, N5933);
and AND2 (N5945, N5909, N401);
nor NOR2 (N5946, N5945, N3798);
not NOT1 (N5947, N5940);
or OR3 (N5948, N5941, N1477, N2925);
or OR4 (N5949, N5948, N3583, N3749, N958);
or OR2 (N5950, N5949, N5019);
or OR3 (N5951, N5934, N866, N5649);
buf BUF1 (N5952, N5950);
or OR2 (N5953, N5951, N3605);
and AND2 (N5954, N5953, N2313);
buf BUF1 (N5955, N5944);
and AND3 (N5956, N5952, N5451, N3692);
or OR4 (N5957, N5946, N2796, N3513, N4269);
not NOT1 (N5958, N5957);
xor XOR2 (N5959, N5954, N302);
nor NOR4 (N5960, N5937, N2725, N378, N3091);
nand NAND4 (N5961, N5942, N4943, N2320, N4746);
xor XOR2 (N5962, N5943, N3154);
or OR2 (N5963, N5959, N4612);
and AND4 (N5964, N5963, N2813, N4703, N575);
xor XOR2 (N5965, N5960, N5061);
and AND2 (N5966, N5955, N399);
buf BUF1 (N5967, N5930);
buf BUF1 (N5968, N5929);
xor XOR2 (N5969, N5947, N1355);
nand NAND3 (N5970, N5965, N1286, N1100);
xor XOR2 (N5971, N5958, N1136);
buf BUF1 (N5972, N5971);
nor NOR3 (N5973, N5967, N3042, N5572);
nand NAND2 (N5974, N5972, N1461);
or OR4 (N5975, N5966, N1216, N5695, N1172);
xor XOR2 (N5976, N5969, N5231);
and AND2 (N5977, N5970, N5710);
not NOT1 (N5978, N5968);
and AND3 (N5979, N5976, N954, N4993);
not NOT1 (N5980, N5978);
buf BUF1 (N5981, N5961);
not NOT1 (N5982, N5979);
and AND3 (N5983, N5964, N5937, N4695);
nor NOR3 (N5984, N5983, N4555, N113);
buf BUF1 (N5985, N5982);
and AND3 (N5986, N5980, N3604, N407);
or OR4 (N5987, N5962, N4963, N2365, N4081);
nand NAND3 (N5988, N5974, N1632, N3937);
nor NOR4 (N5989, N5985, N4193, N502, N5872);
or OR3 (N5990, N5984, N49, N4131);
xor XOR2 (N5991, N5987, N4374);
and AND2 (N5992, N5956, N1297);
nand NAND4 (N5993, N5992, N2201, N5582, N2056);
nor NOR2 (N5994, N5981, N2689);
xor XOR2 (N5995, N5994, N2009);
nand NAND3 (N5996, N5973, N1354, N2754);
buf BUF1 (N5997, N5975);
not NOT1 (N5998, N5990);
and AND2 (N5999, N5977, N3951);
and AND4 (N6000, N5998, N608, N1129, N4059);
not NOT1 (N6001, N5988);
nor NOR3 (N6002, N5989, N3776, N85);
or OR2 (N6003, N6000, N72);
nand NAND4 (N6004, N5986, N3307, N5398, N762);
nor NOR4 (N6005, N5996, N2092, N2913, N5951);
xor XOR2 (N6006, N5993, N3308);
nand NAND2 (N6007, N6004, N4703);
not NOT1 (N6008, N6005);
not NOT1 (N6009, N6007);
or OR4 (N6010, N5991, N635, N1735, N3013);
and AND4 (N6011, N6006, N3771, N111, N5370);
and AND4 (N6012, N6011, N3962, N759, N3066);
and AND2 (N6013, N6012, N5204);
and AND4 (N6014, N5997, N3025, N1815, N3450);
nor NOR3 (N6015, N6010, N2984, N3368);
buf BUF1 (N6016, N6001);
buf BUF1 (N6017, N6008);
nand NAND2 (N6018, N6002, N5037);
or OR4 (N6019, N5999, N4931, N1062, N468);
buf BUF1 (N6020, N6015);
nand NAND3 (N6021, N6016, N4672, N1739);
not NOT1 (N6022, N6003);
buf BUF1 (N6023, N6009);
or OR3 (N6024, N5995, N5407, N256);
not NOT1 (N6025, N6024);
nor NOR4 (N6026, N6022, N221, N925, N793);
or OR2 (N6027, N6026, N4507);
nand NAND2 (N6028, N6019, N1496);
not NOT1 (N6029, N6028);
and AND3 (N6030, N6017, N4211, N567);
nand NAND4 (N6031, N6023, N5667, N3539, N5554);
or OR2 (N6032, N6029, N2419);
buf BUF1 (N6033, N6021);
buf BUF1 (N6034, N6018);
not NOT1 (N6035, N6027);
or OR4 (N6036, N6020, N3244, N935, N2363);
or OR4 (N6037, N6033, N3102, N3155, N919);
buf BUF1 (N6038, N6013);
or OR2 (N6039, N6030, N3812);
nand NAND3 (N6040, N6014, N275, N3163);
buf BUF1 (N6041, N6038);
and AND3 (N6042, N6037, N4192, N1251);
xor XOR2 (N6043, N6036, N5716);
and AND3 (N6044, N6042, N3499, N4954);
and AND4 (N6045, N6044, N4981, N130, N654);
buf BUF1 (N6046, N6031);
and AND2 (N6047, N6043, N2226);
nand NAND2 (N6048, N6032, N2777);
nand NAND2 (N6049, N6040, N1647);
nand NAND3 (N6050, N6025, N2365, N4213);
nor NOR2 (N6051, N6048, N2605);
or OR4 (N6052, N6045, N1520, N423, N4777);
not NOT1 (N6053, N6039);
xor XOR2 (N6054, N6035, N2059);
xor XOR2 (N6055, N6054, N3405);
or OR3 (N6056, N6046, N639, N373);
xor XOR2 (N6057, N6041, N1132);
buf BUF1 (N6058, N6056);
or OR2 (N6059, N6051, N3418);
buf BUF1 (N6060, N6057);
buf BUF1 (N6061, N6059);
nor NOR2 (N6062, N6055, N6031);
xor XOR2 (N6063, N6062, N541);
or OR2 (N6064, N6049, N4737);
not NOT1 (N6065, N6052);
buf BUF1 (N6066, N6063);
buf BUF1 (N6067, N6058);
nor NOR3 (N6068, N6061, N4777, N2963);
xor XOR2 (N6069, N6047, N5089);
or OR2 (N6070, N6053, N2248);
buf BUF1 (N6071, N6068);
nor NOR2 (N6072, N6069, N4861);
nor NOR4 (N6073, N6034, N4018, N5391, N5604);
not NOT1 (N6074, N6065);
buf BUF1 (N6075, N6071);
not NOT1 (N6076, N6070);
xor XOR2 (N6077, N6060, N5647);
buf BUF1 (N6078, N6067);
nor NOR3 (N6079, N6073, N2392, N881);
xor XOR2 (N6080, N6050, N183);
or OR3 (N6081, N6074, N3654, N924);
nor NOR4 (N6082, N6064, N3762, N1856, N155);
nand NAND3 (N6083, N6076, N4493, N4648);
nand NAND2 (N6084, N6072, N551);
nor NOR4 (N6085, N6078, N5926, N5391, N4223);
and AND4 (N6086, N6081, N2983, N502, N51);
not NOT1 (N6087, N6075);
xor XOR2 (N6088, N6084, N5293);
and AND2 (N6089, N6088, N2028);
and AND4 (N6090, N6087, N1692, N2244, N4806);
buf BUF1 (N6091, N6083);
and AND2 (N6092, N6091, N3728);
nand NAND3 (N6093, N6080, N2555, N3499);
or OR3 (N6094, N6079, N5506, N5318);
or OR4 (N6095, N6089, N2557, N5914, N1588);
buf BUF1 (N6096, N6090);
and AND4 (N6097, N6085, N3816, N2209, N5030);
buf BUF1 (N6098, N6095);
nand NAND4 (N6099, N6066, N619, N5959, N5529);
xor XOR2 (N6100, N6094, N2981);
and AND2 (N6101, N6092, N1386);
not NOT1 (N6102, N6100);
nand NAND3 (N6103, N6099, N3890, N3731);
or OR2 (N6104, N6077, N1316);
and AND3 (N6105, N6104, N4761, N5931);
buf BUF1 (N6106, N6082);
or OR2 (N6107, N6103, N1226);
nor NOR4 (N6108, N6102, N3168, N2903, N5404);
xor XOR2 (N6109, N6096, N4193);
nor NOR4 (N6110, N6097, N4876, N3603, N5673);
or OR4 (N6111, N6105, N3965, N5308, N3524);
buf BUF1 (N6112, N6106);
xor XOR2 (N6113, N6109, N3278);
buf BUF1 (N6114, N6113);
not NOT1 (N6115, N6107);
buf BUF1 (N6116, N6114);
or OR2 (N6117, N6112, N4288);
and AND4 (N6118, N6108, N2568, N1687, N5295);
nand NAND3 (N6119, N6093, N5981, N5318);
xor XOR2 (N6120, N6117, N2479);
or OR4 (N6121, N6098, N3531, N2286, N5320);
buf BUF1 (N6122, N6110);
or OR2 (N6123, N6086, N393);
and AND3 (N6124, N6121, N2062, N531);
nor NOR3 (N6125, N6116, N4654, N5332);
buf BUF1 (N6126, N6118);
and AND4 (N6127, N6111, N5101, N12, N1341);
or OR2 (N6128, N6119, N5425);
buf BUF1 (N6129, N6126);
and AND3 (N6130, N6128, N2889, N64);
not NOT1 (N6131, N6122);
xor XOR2 (N6132, N6123, N1499);
xor XOR2 (N6133, N6131, N1707);
or OR3 (N6134, N6127, N5746, N5855);
xor XOR2 (N6135, N6129, N5751);
and AND4 (N6136, N6132, N4049, N1398, N1814);
buf BUF1 (N6137, N6101);
buf BUF1 (N6138, N6130);
or OR3 (N6139, N6120, N839, N3345);
nand NAND3 (N6140, N6138, N1548, N194);
not NOT1 (N6141, N6140);
buf BUF1 (N6142, N6133);
and AND2 (N6143, N6139, N3919);
xor XOR2 (N6144, N6141, N2693);
buf BUF1 (N6145, N6125);
nor NOR4 (N6146, N6145, N2754, N5746, N4974);
not NOT1 (N6147, N6137);
or OR4 (N6148, N6143, N3062, N816, N5878);
xor XOR2 (N6149, N6144, N5293);
xor XOR2 (N6150, N6135, N1267);
or OR2 (N6151, N6150, N2149);
or OR4 (N6152, N6147, N1030, N6050, N4162);
xor XOR2 (N6153, N6148, N5414);
nand NAND2 (N6154, N6134, N4110);
or OR3 (N6155, N6153, N2043, N3950);
not NOT1 (N6156, N6151);
or OR4 (N6157, N6149, N2633, N3105, N362);
nand NAND4 (N6158, N6155, N2142, N1686, N1818);
and AND4 (N6159, N6136, N4144, N5585, N1373);
not NOT1 (N6160, N6152);
nor NOR4 (N6161, N6146, N2328, N1385, N4205);
not NOT1 (N6162, N6154);
nand NAND4 (N6163, N6124, N831, N1544, N2187);
nor NOR2 (N6164, N6156, N17);
nor NOR2 (N6165, N6159, N10);
or OR4 (N6166, N6160, N5388, N1924, N4224);
xor XOR2 (N6167, N6165, N4195);
buf BUF1 (N6168, N6142);
buf BUF1 (N6169, N6161);
not NOT1 (N6170, N6115);
xor XOR2 (N6171, N6157, N2467);
or OR3 (N6172, N6168, N786, N1435);
nand NAND3 (N6173, N6169, N5474, N1159);
xor XOR2 (N6174, N6172, N383);
and AND3 (N6175, N6163, N3908, N3592);
and AND4 (N6176, N6167, N360, N3604, N3307);
and AND2 (N6177, N6174, N2499);
nand NAND3 (N6178, N6171, N436, N6055);
nand NAND3 (N6179, N6164, N4035, N5901);
and AND3 (N6180, N6175, N3363, N3123);
and AND4 (N6181, N6179, N3524, N82, N5749);
xor XOR2 (N6182, N6176, N1642);
buf BUF1 (N6183, N6158);
nand NAND3 (N6184, N6170, N1925, N1858);
nor NOR2 (N6185, N6184, N3110);
xor XOR2 (N6186, N6183, N3014);
nor NOR3 (N6187, N6166, N2517, N530);
nand NAND2 (N6188, N6162, N408);
not NOT1 (N6189, N6173);
buf BUF1 (N6190, N6185);
nand NAND2 (N6191, N6182, N1145);
not NOT1 (N6192, N6180);
nand NAND4 (N6193, N6191, N4527, N3829, N1008);
and AND3 (N6194, N6188, N3169, N334);
buf BUF1 (N6195, N6186);
not NOT1 (N6196, N6195);
nor NOR3 (N6197, N6194, N5393, N5275);
or OR4 (N6198, N6190, N1374, N2387, N117);
nand NAND3 (N6199, N6178, N1681, N2897);
xor XOR2 (N6200, N6181, N3477);
nor NOR4 (N6201, N6187, N2416, N3405, N1706);
nand NAND2 (N6202, N6197, N3938);
xor XOR2 (N6203, N6177, N2747);
buf BUF1 (N6204, N6200);
xor XOR2 (N6205, N6201, N4786);
not NOT1 (N6206, N6204);
not NOT1 (N6207, N6192);
buf BUF1 (N6208, N6193);
and AND3 (N6209, N6206, N105, N1105);
not NOT1 (N6210, N6203);
not NOT1 (N6211, N6210);
and AND3 (N6212, N6199, N2614, N4837);
or OR2 (N6213, N6211, N195);
buf BUF1 (N6214, N6202);
xor XOR2 (N6215, N6214, N5154);
xor XOR2 (N6216, N6212, N1770);
xor XOR2 (N6217, N6213, N2768);
nand NAND3 (N6218, N6207, N5737, N3375);
nor NOR4 (N6219, N6196, N6052, N3606, N5964);
buf BUF1 (N6220, N6209);
nand NAND4 (N6221, N6208, N442, N3073, N5722);
nor NOR4 (N6222, N6217, N2862, N3346, N1773);
or OR4 (N6223, N6221, N4800, N5113, N2319);
xor XOR2 (N6224, N6219, N2194);
or OR4 (N6225, N6223, N3334, N5508, N681);
nor NOR2 (N6226, N6222, N1392);
and AND3 (N6227, N6226, N3233, N2954);
or OR3 (N6228, N6216, N5829, N3342);
nand NAND3 (N6229, N6189, N3280, N540);
or OR2 (N6230, N6220, N5017);
or OR2 (N6231, N6230, N1876);
nand NAND3 (N6232, N6225, N1115, N3958);
buf BUF1 (N6233, N6215);
buf BUF1 (N6234, N6232);
buf BUF1 (N6235, N6218);
nand NAND2 (N6236, N6231, N5590);
or OR3 (N6237, N6228, N701, N334);
nor NOR3 (N6238, N6233, N5792, N2501);
buf BUF1 (N6239, N6224);
nor NOR4 (N6240, N6205, N2568, N4686, N3379);
nand NAND4 (N6241, N6235, N690, N5418, N752);
not NOT1 (N6242, N6238);
xor XOR2 (N6243, N6242, N1046);
nand NAND4 (N6244, N6240, N3828, N6024, N4544);
nand NAND2 (N6245, N6243, N4699);
nand NAND2 (N6246, N6227, N285);
or OR3 (N6247, N6241, N5884, N1038);
nand NAND3 (N6248, N6234, N4473, N5182);
buf BUF1 (N6249, N6229);
buf BUF1 (N6250, N6198);
or OR2 (N6251, N6244, N4596);
xor XOR2 (N6252, N6249, N1361);
nor NOR3 (N6253, N6250, N4029, N3089);
or OR4 (N6254, N6239, N3547, N237, N1473);
nor NOR3 (N6255, N6248, N2137, N6110);
nor NOR2 (N6256, N6252, N3741);
xor XOR2 (N6257, N6247, N618);
xor XOR2 (N6258, N6245, N5874);
nand NAND2 (N6259, N6236, N648);
buf BUF1 (N6260, N6246);
nor NOR3 (N6261, N6256, N2575, N800);
and AND3 (N6262, N6255, N4903, N568);
or OR2 (N6263, N6261, N5101);
xor XOR2 (N6264, N6237, N1500);
nor NOR4 (N6265, N6263, N875, N674, N4734);
buf BUF1 (N6266, N6253);
buf BUF1 (N6267, N6266);
nand NAND2 (N6268, N6267, N3195);
or OR2 (N6269, N6254, N451);
or OR4 (N6270, N6268, N4586, N4699, N153);
or OR3 (N6271, N6259, N5355, N2626);
not NOT1 (N6272, N6265);
not NOT1 (N6273, N6272);
buf BUF1 (N6274, N6262);
nand NAND3 (N6275, N6258, N2381, N648);
and AND3 (N6276, N6264, N5055, N202);
xor XOR2 (N6277, N6271, N731);
or OR3 (N6278, N6275, N1985, N3076);
nor NOR2 (N6279, N6274, N725);
buf BUF1 (N6280, N6276);
not NOT1 (N6281, N6280);
not NOT1 (N6282, N6260);
buf BUF1 (N6283, N6282);
nand NAND4 (N6284, N6270, N1732, N4639, N439);
not NOT1 (N6285, N6279);
and AND3 (N6286, N6257, N5162, N4284);
or OR2 (N6287, N6251, N856);
xor XOR2 (N6288, N6278, N2374);
xor XOR2 (N6289, N6285, N594);
and AND2 (N6290, N6281, N5558);
or OR3 (N6291, N6287, N2350, N47);
xor XOR2 (N6292, N6283, N5796);
buf BUF1 (N6293, N6269);
and AND4 (N6294, N6291, N2691, N1826, N2643);
xor XOR2 (N6295, N6277, N756);
xor XOR2 (N6296, N6284, N1193);
not NOT1 (N6297, N6296);
not NOT1 (N6298, N6289);
xor XOR2 (N6299, N6290, N3833);
not NOT1 (N6300, N6294);
and AND3 (N6301, N6298, N3666, N5447);
not NOT1 (N6302, N6288);
not NOT1 (N6303, N6297);
buf BUF1 (N6304, N6299);
not NOT1 (N6305, N6293);
not NOT1 (N6306, N6305);
nand NAND2 (N6307, N6304, N1013);
or OR4 (N6308, N6306, N5835, N1485, N5141);
buf BUF1 (N6309, N6302);
xor XOR2 (N6310, N6309, N3396);
not NOT1 (N6311, N6307);
nor NOR4 (N6312, N6311, N6310, N480, N312);
nor NOR4 (N6313, N3613, N6105, N3035, N1223);
nand NAND4 (N6314, N6286, N5911, N3685, N1717);
not NOT1 (N6315, N6314);
and AND3 (N6316, N6292, N5825, N4144);
not NOT1 (N6317, N6313);
not NOT1 (N6318, N6308);
not NOT1 (N6319, N6315);
not NOT1 (N6320, N6303);
buf BUF1 (N6321, N6300);
not NOT1 (N6322, N6320);
nor NOR3 (N6323, N6322, N3643, N5261);
and AND3 (N6324, N6323, N168, N4149);
buf BUF1 (N6325, N6273);
nor NOR3 (N6326, N6295, N4301, N4896);
and AND4 (N6327, N6318, N3640, N3646, N1091);
or OR2 (N6328, N6325, N2712);
buf BUF1 (N6329, N6327);
not NOT1 (N6330, N6319);
nand NAND2 (N6331, N6301, N3743);
or OR3 (N6332, N6321, N1521, N770);
buf BUF1 (N6333, N6331);
xor XOR2 (N6334, N6326, N5484);
and AND4 (N6335, N6329, N5601, N5716, N5675);
buf BUF1 (N6336, N6316);
or OR2 (N6337, N6335, N1600);
or OR3 (N6338, N6330, N700, N3219);
not NOT1 (N6339, N6338);
xor XOR2 (N6340, N6332, N5454);
nand NAND4 (N6341, N6336, N2213, N3247, N3122);
or OR2 (N6342, N6328, N724);
buf BUF1 (N6343, N6324);
nand NAND3 (N6344, N6342, N4588, N3973);
or OR3 (N6345, N6339, N5288, N2318);
and AND3 (N6346, N6312, N3842, N5172);
buf BUF1 (N6347, N6317);
xor XOR2 (N6348, N6343, N502);
buf BUF1 (N6349, N6345);
or OR4 (N6350, N6347, N483, N3749, N2750);
nand NAND2 (N6351, N6337, N1884);
nand NAND3 (N6352, N6350, N2758, N5243);
nand NAND2 (N6353, N6348, N3329);
buf BUF1 (N6354, N6353);
nor NOR2 (N6355, N6351, N3085);
and AND2 (N6356, N6354, N2573);
nor NOR3 (N6357, N6352, N757, N4196);
xor XOR2 (N6358, N6341, N5285);
xor XOR2 (N6359, N6355, N2575);
buf BUF1 (N6360, N6334);
xor XOR2 (N6361, N6360, N3289);
and AND3 (N6362, N6333, N3415, N3204);
and AND4 (N6363, N6362, N3787, N4969, N5013);
or OR2 (N6364, N6346, N4854);
or OR3 (N6365, N6359, N877, N4132);
nand NAND3 (N6366, N6365, N2618, N643);
nor NOR3 (N6367, N6356, N3439, N3827);
or OR2 (N6368, N6358, N680);
buf BUF1 (N6369, N6364);
nor NOR2 (N6370, N6340, N5372);
nor NOR3 (N6371, N6367, N3405, N2794);
not NOT1 (N6372, N6363);
buf BUF1 (N6373, N6371);
not NOT1 (N6374, N6366);
or OR3 (N6375, N6374, N1587, N4260);
xor XOR2 (N6376, N6373, N3439);
or OR4 (N6377, N6357, N5648, N2057, N2437);
not NOT1 (N6378, N6377);
or OR4 (N6379, N6378, N4062, N222, N1887);
not NOT1 (N6380, N6370);
nand NAND3 (N6381, N6349, N2513, N1160);
and AND3 (N6382, N6369, N5983, N115);
and AND4 (N6383, N6380, N3758, N1350, N350);
not NOT1 (N6384, N6382);
nand NAND3 (N6385, N6383, N2216, N6264);
or OR2 (N6386, N6372, N2722);
buf BUF1 (N6387, N6376);
nand NAND3 (N6388, N6368, N672, N4613);
and AND3 (N6389, N6381, N5789, N496);
nand NAND4 (N6390, N6384, N4589, N5683, N878);
buf BUF1 (N6391, N6386);
not NOT1 (N6392, N6375);
nor NOR2 (N6393, N6391, N5948);
not NOT1 (N6394, N6393);
not NOT1 (N6395, N6379);
or OR4 (N6396, N6389, N3079, N3274, N5572);
and AND2 (N6397, N6390, N3467);
and AND2 (N6398, N6395, N2025);
not NOT1 (N6399, N6361);
buf BUF1 (N6400, N6385);
and AND3 (N6401, N6387, N5808, N2452);
xor XOR2 (N6402, N6401, N3270);
or OR4 (N6403, N6394, N2362, N3426, N2747);
xor XOR2 (N6404, N6399, N3036);
not NOT1 (N6405, N6388);
and AND2 (N6406, N6403, N3123);
nand NAND4 (N6407, N6398, N3701, N4765, N693);
not NOT1 (N6408, N6396);
nand NAND4 (N6409, N6407, N1621, N3533, N5285);
or OR4 (N6410, N6404, N872, N2355, N5660);
buf BUF1 (N6411, N6402);
buf BUF1 (N6412, N6397);
not NOT1 (N6413, N6410);
xor XOR2 (N6414, N6344, N4803);
xor XOR2 (N6415, N6412, N860);
buf BUF1 (N6416, N6414);
buf BUF1 (N6417, N6408);
buf BUF1 (N6418, N6409);
buf BUF1 (N6419, N6416);
xor XOR2 (N6420, N6418, N430);
nand NAND4 (N6421, N6392, N470, N1429, N2503);
nor NOR2 (N6422, N6405, N5751);
buf BUF1 (N6423, N6419);
nand NAND3 (N6424, N6421, N387, N4537);
or OR3 (N6425, N6400, N366, N6179);
nand NAND2 (N6426, N6406, N5379);
nor NOR2 (N6427, N6413, N4729);
xor XOR2 (N6428, N6427, N3);
not NOT1 (N6429, N6417);
and AND4 (N6430, N6415, N2741, N529, N3155);
xor XOR2 (N6431, N6420, N1335);
and AND4 (N6432, N6424, N5373, N3771, N5185);
or OR4 (N6433, N6422, N319, N2646, N3051);
not NOT1 (N6434, N6429);
xor XOR2 (N6435, N6426, N5876);
nand NAND4 (N6436, N6435, N1613, N2738, N21);
buf BUF1 (N6437, N6432);
buf BUF1 (N6438, N6430);
nor NOR4 (N6439, N6433, N2059, N4192, N277);
nor NOR3 (N6440, N6439, N921, N3996);
nor NOR4 (N6441, N6411, N5727, N5885, N2161);
nor NOR3 (N6442, N6434, N1868, N4030);
not NOT1 (N6443, N6441);
or OR4 (N6444, N6437, N2749, N4230, N2639);
not NOT1 (N6445, N6444);
or OR3 (N6446, N6428, N4977, N2241);
nor NOR4 (N6447, N6431, N179, N6011, N5777);
xor XOR2 (N6448, N6423, N597);
not NOT1 (N6449, N6448);
or OR2 (N6450, N6425, N1881);
or OR4 (N6451, N6446, N664, N3810, N3239);
or OR4 (N6452, N6447, N5015, N5382, N2071);
or OR2 (N6453, N6452, N1472);
not NOT1 (N6454, N6449);
buf BUF1 (N6455, N6440);
and AND4 (N6456, N6450, N523, N2265, N2546);
not NOT1 (N6457, N6438);
nor NOR4 (N6458, N6451, N895, N4207, N1256);
xor XOR2 (N6459, N6443, N4664);
or OR3 (N6460, N6453, N4865, N788);
not NOT1 (N6461, N6455);
buf BUF1 (N6462, N6456);
xor XOR2 (N6463, N6460, N3716);
buf BUF1 (N6464, N6463);
and AND2 (N6465, N6454, N4157);
xor XOR2 (N6466, N6442, N2182);
and AND3 (N6467, N6461, N3747, N4067);
or OR2 (N6468, N6457, N2570);
buf BUF1 (N6469, N6436);
not NOT1 (N6470, N6458);
buf BUF1 (N6471, N6468);
nor NOR2 (N6472, N6465, N6415);
not NOT1 (N6473, N6459);
and AND3 (N6474, N6467, N3056, N5128);
and AND3 (N6475, N6469, N1895, N3414);
nand NAND2 (N6476, N6462, N1874);
or OR3 (N6477, N6470, N2079, N3263);
not NOT1 (N6478, N6466);
nor NOR4 (N6479, N6477, N5469, N3352, N3074);
not NOT1 (N6480, N6472);
not NOT1 (N6481, N6475);
or OR3 (N6482, N6480, N21, N2023);
not NOT1 (N6483, N6464);
nor NOR4 (N6484, N6482, N3150, N1054, N1848);
and AND4 (N6485, N6445, N5258, N2213, N5900);
nand NAND4 (N6486, N6478, N136, N1733, N2975);
or OR2 (N6487, N6473, N6373);
buf BUF1 (N6488, N6471);
or OR4 (N6489, N6479, N4429, N3682, N1175);
xor XOR2 (N6490, N6476, N5893);
nor NOR3 (N6491, N6489, N5095, N4087);
or OR3 (N6492, N6490, N5730, N5290);
nor NOR4 (N6493, N6481, N917, N2234, N1880);
or OR2 (N6494, N6491, N5946);
nor NOR2 (N6495, N6474, N1077);
nor NOR3 (N6496, N6483, N4771, N5692);
or OR3 (N6497, N6493, N6457, N4960);
nand NAND3 (N6498, N6492, N2762, N2872);
or OR3 (N6499, N6488, N2502, N6148);
and AND3 (N6500, N6498, N3610, N5190);
and AND3 (N6501, N6494, N1415, N6299);
buf BUF1 (N6502, N6485);
buf BUF1 (N6503, N6500);
buf BUF1 (N6504, N6497);
nor NOR4 (N6505, N6487, N1364, N4183, N3379);
nor NOR4 (N6506, N6496, N5666, N2064, N4594);
and AND2 (N6507, N6503, N1298);
buf BUF1 (N6508, N6504);
buf BUF1 (N6509, N6508);
buf BUF1 (N6510, N6499);
not NOT1 (N6511, N6510);
buf BUF1 (N6512, N6505);
nor NOR3 (N6513, N6506, N3585, N6012);
nand NAND4 (N6514, N6509, N2263, N1139, N640);
not NOT1 (N6515, N6507);
not NOT1 (N6516, N6502);
buf BUF1 (N6517, N6501);
not NOT1 (N6518, N6511);
xor XOR2 (N6519, N6513, N2490);
nor NOR4 (N6520, N6495, N3529, N5606, N5545);
nor NOR3 (N6521, N6517, N5057, N3544);
xor XOR2 (N6522, N6520, N1595);
nor NOR3 (N6523, N6515, N2735, N127);
nor NOR4 (N6524, N6484, N6413, N2874, N601);
xor XOR2 (N6525, N6514, N3858);
nor NOR3 (N6526, N6524, N4394, N1643);
and AND3 (N6527, N6519, N5429, N1071);
or OR3 (N6528, N6522, N2418, N4017);
nor NOR3 (N6529, N6486, N4840, N1284);
nand NAND3 (N6530, N6528, N719, N3233);
nand NAND3 (N6531, N6516, N418, N6008);
or OR2 (N6532, N6518, N6401);
or OR3 (N6533, N6531, N5458, N3311);
xor XOR2 (N6534, N6523, N1014);
nand NAND4 (N6535, N6512, N6182, N4249, N690);
nand NAND4 (N6536, N6532, N1847, N6499, N2013);
nand NAND2 (N6537, N6521, N4366);
buf BUF1 (N6538, N6527);
not NOT1 (N6539, N6536);
and AND3 (N6540, N6537, N3811, N4672);
buf BUF1 (N6541, N6525);
buf BUF1 (N6542, N6541);
nand NAND2 (N6543, N6542, N3906);
buf BUF1 (N6544, N6539);
and AND4 (N6545, N6538, N5837, N3246, N230);
nor NOR3 (N6546, N6535, N3949, N5216);
or OR4 (N6547, N6529, N1683, N2256, N2515);
nand NAND4 (N6548, N6526, N5813, N5651, N5804);
buf BUF1 (N6549, N6545);
and AND4 (N6550, N6533, N5074, N854, N1712);
not NOT1 (N6551, N6530);
and AND4 (N6552, N6546, N1535, N5767, N1500);
buf BUF1 (N6553, N6551);
or OR3 (N6554, N6544, N5130, N5741);
not NOT1 (N6555, N6549);
nor NOR4 (N6556, N6534, N5097, N4614, N4676);
not NOT1 (N6557, N6555);
and AND4 (N6558, N6557, N5048, N1764, N5596);
xor XOR2 (N6559, N6543, N2063);
buf BUF1 (N6560, N6553);
nand NAND3 (N6561, N6556, N1748, N1061);
nor NOR2 (N6562, N6547, N2967);
nor NOR4 (N6563, N6559, N3580, N5662, N5230);
buf BUF1 (N6564, N6552);
or OR4 (N6565, N6554, N3401, N6262, N1243);
or OR4 (N6566, N6562, N6465, N1894, N5771);
nor NOR3 (N6567, N6550, N4948, N745);
nand NAND3 (N6568, N6567, N3593, N4879);
and AND4 (N6569, N6564, N4843, N474, N2488);
not NOT1 (N6570, N6565);
buf BUF1 (N6571, N6558);
buf BUF1 (N6572, N6568);
not NOT1 (N6573, N6570);
xor XOR2 (N6574, N6572, N4283);
not NOT1 (N6575, N6571);
not NOT1 (N6576, N6560);
nor NOR2 (N6577, N6575, N1516);
xor XOR2 (N6578, N6548, N4699);
buf BUF1 (N6579, N6577);
buf BUF1 (N6580, N6576);
or OR4 (N6581, N6561, N846, N1207, N4452);
buf BUF1 (N6582, N6579);
not NOT1 (N6583, N6540);
buf BUF1 (N6584, N6569);
and AND3 (N6585, N6573, N5923, N4834);
and AND2 (N6586, N6578, N4288);
buf BUF1 (N6587, N6582);
buf BUF1 (N6588, N6566);
and AND3 (N6589, N6584, N2557, N2154);
buf BUF1 (N6590, N6580);
nor NOR2 (N6591, N6586, N220);
xor XOR2 (N6592, N6581, N305);
or OR3 (N6593, N6590, N633, N3776);
not NOT1 (N6594, N6591);
not NOT1 (N6595, N6589);
xor XOR2 (N6596, N6595, N3295);
not NOT1 (N6597, N6574);
and AND3 (N6598, N6588, N769, N2459);
nand NAND3 (N6599, N6594, N5199, N6581);
nor NOR3 (N6600, N6583, N1827, N543);
not NOT1 (N6601, N6599);
xor XOR2 (N6602, N6600, N2306);
or OR2 (N6603, N6563, N2567);
not NOT1 (N6604, N6602);
or OR3 (N6605, N6587, N5223, N2017);
or OR2 (N6606, N6585, N6377);
nand NAND3 (N6607, N6603, N5588, N5631);
nand NAND2 (N6608, N6592, N273);
buf BUF1 (N6609, N6596);
buf BUF1 (N6610, N6606);
nor NOR3 (N6611, N6605, N5796, N4260);
nor NOR3 (N6612, N6607, N4194, N1725);
nor NOR4 (N6613, N6612, N278, N2404, N5012);
xor XOR2 (N6614, N6601, N3944);
xor XOR2 (N6615, N6611, N2923);
and AND4 (N6616, N6614, N6562, N3074, N2205);
or OR4 (N6617, N6597, N1491, N5971, N4202);
not NOT1 (N6618, N6610);
not NOT1 (N6619, N6604);
nand NAND3 (N6620, N6598, N4671, N2969);
or OR4 (N6621, N6615, N54, N618, N3666);
not NOT1 (N6622, N6613);
xor XOR2 (N6623, N6619, N1315);
nand NAND2 (N6624, N6609, N3132);
nand NAND3 (N6625, N6623, N982, N1451);
xor XOR2 (N6626, N6617, N2223);
and AND2 (N6627, N6621, N1580);
or OR2 (N6628, N6627, N3656);
nand NAND4 (N6629, N6616, N1166, N3640, N2704);
nand NAND3 (N6630, N6624, N4236, N6586);
nor NOR4 (N6631, N6628, N1803, N89, N3391);
or OR4 (N6632, N6620, N3015, N2769, N762);
or OR4 (N6633, N6630, N4039, N4501, N1754);
nand NAND3 (N6634, N6625, N5921, N5037);
xor XOR2 (N6635, N6629, N607);
xor XOR2 (N6636, N6622, N1086);
and AND3 (N6637, N6608, N5670, N5495);
or OR3 (N6638, N6632, N4334, N556);
nor NOR4 (N6639, N6631, N2146, N876, N1692);
not NOT1 (N6640, N6639);
not NOT1 (N6641, N6640);
and AND3 (N6642, N6637, N6036, N1330);
or OR4 (N6643, N6638, N3147, N3213, N678);
buf BUF1 (N6644, N6642);
and AND3 (N6645, N6635, N756, N5319);
xor XOR2 (N6646, N6636, N574);
nand NAND2 (N6647, N6646, N2840);
buf BUF1 (N6648, N6647);
nor NOR2 (N6649, N6644, N1393);
buf BUF1 (N6650, N6645);
nand NAND4 (N6651, N6618, N4775, N178, N4150);
and AND2 (N6652, N6634, N314);
not NOT1 (N6653, N6650);
and AND4 (N6654, N6641, N4938, N1173, N5369);
and AND2 (N6655, N6648, N6395);
buf BUF1 (N6656, N6633);
nand NAND4 (N6657, N6651, N5450, N4135, N1351);
or OR4 (N6658, N6626, N2291, N1514, N6438);
nor NOR3 (N6659, N6643, N4091, N239);
or OR4 (N6660, N6653, N2365, N4411, N730);
and AND4 (N6661, N6649, N3887, N971, N2500);
xor XOR2 (N6662, N6659, N1587);
xor XOR2 (N6663, N6593, N3837);
nor NOR3 (N6664, N6660, N3508, N4040);
nand NAND3 (N6665, N6661, N6113, N4092);
or OR4 (N6666, N6657, N5136, N5392, N5504);
not NOT1 (N6667, N6666);
xor XOR2 (N6668, N6667, N5108);
not NOT1 (N6669, N6658);
buf BUF1 (N6670, N6669);
not NOT1 (N6671, N6663);
buf BUF1 (N6672, N6670);
and AND3 (N6673, N6656, N3178, N99);
or OR2 (N6674, N6665, N196);
buf BUF1 (N6675, N6674);
buf BUF1 (N6676, N6671);
or OR3 (N6677, N6662, N4813, N4141);
buf BUF1 (N6678, N6654);
and AND4 (N6679, N6655, N1062, N1363, N4932);
xor XOR2 (N6680, N6668, N5505);
nand NAND3 (N6681, N6675, N2152, N321);
buf BUF1 (N6682, N6652);
not NOT1 (N6683, N6672);
nand NAND2 (N6684, N6677, N4666);
nand NAND2 (N6685, N6684, N2168);
nand NAND2 (N6686, N6682, N6233);
nor NOR3 (N6687, N6679, N5278, N147);
xor XOR2 (N6688, N6685, N87);
buf BUF1 (N6689, N6686);
buf BUF1 (N6690, N6673);
buf BUF1 (N6691, N6680);
buf BUF1 (N6692, N6690);
not NOT1 (N6693, N6692);
not NOT1 (N6694, N6691);
nand NAND2 (N6695, N6664, N3620);
or OR3 (N6696, N6695, N326, N3216);
not NOT1 (N6697, N6676);
or OR3 (N6698, N6697, N5609, N4354);
nand NAND4 (N6699, N6683, N2340, N2861, N4723);
xor XOR2 (N6700, N6681, N756);
and AND4 (N6701, N6688, N3500, N773, N3852);
and AND2 (N6702, N6696, N2607);
or OR3 (N6703, N6687, N2268, N431);
buf BUF1 (N6704, N6678);
and AND3 (N6705, N6700, N1263, N1469);
nor NOR4 (N6706, N6693, N3379, N5739, N6199);
nor NOR2 (N6707, N6689, N1764);
buf BUF1 (N6708, N6704);
not NOT1 (N6709, N6701);
and AND3 (N6710, N6694, N958, N4282);
xor XOR2 (N6711, N6703, N6001);
nor NOR2 (N6712, N6699, N772);
or OR3 (N6713, N6711, N1508, N2236);
xor XOR2 (N6714, N6706, N6433);
nor NOR3 (N6715, N6713, N4230, N2434);
buf BUF1 (N6716, N6708);
and AND3 (N6717, N6716, N2940, N407);
not NOT1 (N6718, N6709);
or OR2 (N6719, N6705, N5536);
buf BUF1 (N6720, N6698);
xor XOR2 (N6721, N6719, N3192);
buf BUF1 (N6722, N6702);
not NOT1 (N6723, N6718);
and AND2 (N6724, N6707, N3087);
xor XOR2 (N6725, N6720, N6476);
xor XOR2 (N6726, N6723, N3915);
nand NAND3 (N6727, N6717, N6493, N3102);
nand NAND3 (N6728, N6721, N6005, N4778);
xor XOR2 (N6729, N6725, N6255);
buf BUF1 (N6730, N6728);
nor NOR3 (N6731, N6710, N2325, N6294);
nand NAND3 (N6732, N6715, N1692, N3859);
nor NOR2 (N6733, N6730, N2922);
xor XOR2 (N6734, N6733, N767);
nor NOR3 (N6735, N6734, N2042, N1491);
and AND3 (N6736, N6714, N2942, N6264);
buf BUF1 (N6737, N6727);
nand NAND3 (N6738, N6726, N3234, N5753);
nor NOR3 (N6739, N6732, N3708, N5262);
buf BUF1 (N6740, N6739);
not NOT1 (N6741, N6712);
nor NOR3 (N6742, N6731, N4228, N2280);
or OR3 (N6743, N6740, N3174, N2129);
xor XOR2 (N6744, N6743, N82);
or OR4 (N6745, N6736, N3253, N3483, N5391);
and AND4 (N6746, N6722, N5314, N3779, N6618);
or OR4 (N6747, N6741, N1051, N3196, N1830);
nor NOR3 (N6748, N6745, N1049, N3678);
buf BUF1 (N6749, N6738);
nor NOR4 (N6750, N6744, N5021, N5937, N2166);
nor NOR2 (N6751, N6737, N1763);
and AND4 (N6752, N6751, N6049, N1687, N2691);
nor NOR3 (N6753, N6748, N1299, N1688);
or OR3 (N6754, N6752, N5134, N6388);
buf BUF1 (N6755, N6735);
not NOT1 (N6756, N6746);
xor XOR2 (N6757, N6753, N2792);
buf BUF1 (N6758, N6750);
nand NAND3 (N6759, N6729, N231, N4854);
or OR3 (N6760, N6756, N2372, N4778);
or OR3 (N6761, N6760, N5150, N2752);
not NOT1 (N6762, N6747);
nand NAND3 (N6763, N6749, N5535, N5629);
and AND2 (N6764, N6724, N5264);
or OR2 (N6765, N6757, N6299);
not NOT1 (N6766, N6761);
nand NAND3 (N6767, N6763, N4083, N5229);
nor NOR3 (N6768, N6754, N6152, N973);
or OR4 (N6769, N6768, N357, N5234, N5359);
not NOT1 (N6770, N6764);
nor NOR4 (N6771, N6765, N4844, N1337, N1017);
and AND3 (N6772, N6755, N3319, N512);
nand NAND3 (N6773, N6762, N5355, N71);
and AND4 (N6774, N6770, N778, N5843, N4644);
nand NAND4 (N6775, N6767, N1561, N2009, N914);
or OR2 (N6776, N6773, N863);
nor NOR2 (N6777, N6771, N2556);
nand NAND4 (N6778, N6774, N6757, N6248, N3452);
and AND4 (N6779, N6766, N875, N5938, N682);
xor XOR2 (N6780, N6775, N1799);
xor XOR2 (N6781, N6772, N1976);
and AND2 (N6782, N6780, N1469);
nand NAND2 (N6783, N6776, N1156);
nand NAND2 (N6784, N6777, N4716);
nor NOR2 (N6785, N6742, N1517);
and AND3 (N6786, N6781, N6718, N679);
nand NAND4 (N6787, N6783, N33, N1838, N2111);
not NOT1 (N6788, N6782);
or OR2 (N6789, N6786, N878);
not NOT1 (N6790, N6778);
xor XOR2 (N6791, N6787, N1068);
nor NOR4 (N6792, N6759, N4292, N2866, N201);
nor NOR4 (N6793, N6791, N3625, N369, N2857);
nor NOR4 (N6794, N6788, N5895, N5935, N809);
xor XOR2 (N6795, N6785, N5844);
not NOT1 (N6796, N6794);
not NOT1 (N6797, N6795);
nor NOR4 (N6798, N6789, N5570, N3324, N650);
nor NOR4 (N6799, N6793, N4962, N5035, N3474);
and AND3 (N6800, N6792, N3465, N2597);
nor NOR2 (N6801, N6790, N457);
not NOT1 (N6802, N6779);
and AND3 (N6803, N6799, N1508, N749);
nand NAND2 (N6804, N6784, N1678);
buf BUF1 (N6805, N6758);
and AND3 (N6806, N6801, N3776, N4651);
nor NOR2 (N6807, N6805, N668);
or OR4 (N6808, N6769, N3188, N6039, N2043);
nand NAND4 (N6809, N6796, N4880, N4239, N6752);
and AND3 (N6810, N6802, N2322, N6021);
nand NAND4 (N6811, N6809, N4427, N1319, N88);
nand NAND2 (N6812, N6804, N2262);
xor XOR2 (N6813, N6806, N5314);
and AND2 (N6814, N6810, N194);
and AND3 (N6815, N6814, N2298, N3155);
xor XOR2 (N6816, N6808, N6638);
or OR2 (N6817, N6797, N5351);
nand NAND4 (N6818, N6807, N336, N2882, N26);
xor XOR2 (N6819, N6816, N2271);
nand NAND4 (N6820, N6813, N4511, N5621, N6157);
nor NOR4 (N6821, N6817, N1883, N2897, N3106);
and AND3 (N6822, N6812, N4680, N5569);
not NOT1 (N6823, N6819);
or OR4 (N6824, N6822, N2086, N4624, N5255);
xor XOR2 (N6825, N6824, N43);
nor NOR4 (N6826, N6820, N6479, N3547, N5508);
not NOT1 (N6827, N6798);
not NOT1 (N6828, N6826);
xor XOR2 (N6829, N6818, N2482);
nor NOR3 (N6830, N6829, N437, N351);
not NOT1 (N6831, N6800);
nand NAND4 (N6832, N6830, N1570, N6627, N6748);
or OR4 (N6833, N6821, N1051, N6797, N4865);
xor XOR2 (N6834, N6833, N3722);
buf BUF1 (N6835, N6827);
buf BUF1 (N6836, N6835);
nor NOR4 (N6837, N6803, N4506, N325, N3527);
nand NAND3 (N6838, N6828, N4840, N1192);
nor NOR3 (N6839, N6836, N2856, N4227);
or OR2 (N6840, N6838, N5223);
buf BUF1 (N6841, N6834);
or OR3 (N6842, N6825, N2379, N6691);
and AND3 (N6843, N6839, N2346, N542);
and AND2 (N6844, N6841, N331);
xor XOR2 (N6845, N6811, N199);
buf BUF1 (N6846, N6845);
nor NOR4 (N6847, N6844, N1787, N1137, N3195);
xor XOR2 (N6848, N6840, N1667);
and AND2 (N6849, N6843, N5944);
and AND2 (N6850, N6848, N6264);
or OR4 (N6851, N6846, N5420, N1894, N2507);
nor NOR2 (N6852, N6847, N2229);
buf BUF1 (N6853, N6831);
nand NAND3 (N6854, N6850, N3374, N4119);
nor NOR2 (N6855, N6815, N1643);
xor XOR2 (N6856, N6854, N3648);
nor NOR2 (N6857, N6853, N6153);
or OR2 (N6858, N6842, N1258);
and AND2 (N6859, N6852, N2071);
xor XOR2 (N6860, N6856, N3827);
nor NOR3 (N6861, N6857, N6332, N5470);
xor XOR2 (N6862, N6837, N3275);
buf BUF1 (N6863, N6858);
nor NOR3 (N6864, N6849, N1885, N262);
buf BUF1 (N6865, N6862);
nor NOR4 (N6866, N6861, N2472, N782, N5616);
nor NOR4 (N6867, N6855, N3954, N2225, N3304);
or OR4 (N6868, N6851, N6144, N6146, N1621);
or OR3 (N6869, N6863, N5164, N5367);
nor NOR4 (N6870, N6823, N1659, N4713, N5626);
or OR3 (N6871, N6869, N5597, N2608);
nand NAND3 (N6872, N6866, N4350, N4274);
or OR3 (N6873, N6870, N1321, N6502);
or OR2 (N6874, N6865, N2902);
or OR2 (N6875, N6873, N5085);
buf BUF1 (N6876, N6868);
nand NAND2 (N6877, N6867, N552);
not NOT1 (N6878, N6859);
nor NOR3 (N6879, N6860, N36, N3686);
and AND4 (N6880, N6871, N6078, N3319, N5629);
or OR2 (N6881, N6876, N3377);
buf BUF1 (N6882, N6877);
not NOT1 (N6883, N6878);
buf BUF1 (N6884, N6832);
nand NAND2 (N6885, N6875, N2043);
and AND3 (N6886, N6885, N3366, N4732);
buf BUF1 (N6887, N6880);
nand NAND3 (N6888, N6874, N1654, N5186);
nand NAND3 (N6889, N6872, N1761, N97);
xor XOR2 (N6890, N6881, N3113);
nand NAND2 (N6891, N6887, N2573);
and AND4 (N6892, N6882, N2614, N6041, N3268);
xor XOR2 (N6893, N6890, N4778);
nand NAND3 (N6894, N6879, N720, N1898);
xor XOR2 (N6895, N6886, N5572);
and AND2 (N6896, N6894, N6638);
and AND3 (N6897, N6888, N5399, N5612);
nand NAND2 (N6898, N6891, N4782);
xor XOR2 (N6899, N6898, N6688);
xor XOR2 (N6900, N6893, N6080);
nor NOR3 (N6901, N6884, N4035, N2528);
or OR3 (N6902, N6899, N4422, N1459);
nand NAND3 (N6903, N6897, N1607, N6598);
nand NAND3 (N6904, N6889, N5424, N5308);
or OR3 (N6905, N6904, N3175, N5618);
nand NAND4 (N6906, N6883, N5266, N4391, N1008);
xor XOR2 (N6907, N6895, N6267);
or OR3 (N6908, N6900, N6166, N2892);
or OR4 (N6909, N6896, N2756, N4991, N2647);
not NOT1 (N6910, N6909);
xor XOR2 (N6911, N6864, N3966);
nand NAND2 (N6912, N6910, N6253);
and AND4 (N6913, N6902, N1503, N577, N3868);
nand NAND3 (N6914, N6907, N5288, N222);
not NOT1 (N6915, N6905);
nor NOR2 (N6916, N6913, N3758);
nand NAND4 (N6917, N6914, N6054, N6089, N5148);
nand NAND4 (N6918, N6892, N2750, N375, N4470);
buf BUF1 (N6919, N6903);
not NOT1 (N6920, N6916);
or OR2 (N6921, N6911, N4935);
nand NAND3 (N6922, N6908, N557, N1927);
or OR3 (N6923, N6918, N2307, N306);
xor XOR2 (N6924, N6921, N2237);
nor NOR2 (N6925, N6919, N3571);
nand NAND3 (N6926, N6912, N473, N1403);
not NOT1 (N6927, N6915);
xor XOR2 (N6928, N6920, N6391);
nand NAND4 (N6929, N6926, N3969, N770, N1396);
or OR4 (N6930, N6901, N4941, N2040, N3186);
buf BUF1 (N6931, N6930);
and AND4 (N6932, N6924, N6395, N5919, N739);
xor XOR2 (N6933, N6929, N2339);
and AND2 (N6934, N6923, N4640);
nand NAND3 (N6935, N6934, N3037, N939);
or OR2 (N6936, N6917, N4343);
nor NOR2 (N6937, N6928, N6842);
nand NAND3 (N6938, N6925, N4746, N942);
nor NOR2 (N6939, N6922, N3355);
nand NAND4 (N6940, N6931, N5358, N437, N1775);
xor XOR2 (N6941, N6927, N3804);
nor NOR3 (N6942, N6906, N6286, N3320);
nor NOR2 (N6943, N6941, N1287);
nor NOR4 (N6944, N6935, N1250, N1426, N2623);
and AND2 (N6945, N6936, N2682);
and AND2 (N6946, N6939, N4477);
nor NOR4 (N6947, N6938, N5622, N355, N5326);
and AND2 (N6948, N6943, N6013);
nand NAND3 (N6949, N6947, N1260, N549);
xor XOR2 (N6950, N6933, N1579);
xor XOR2 (N6951, N6945, N3452);
nand NAND3 (N6952, N6951, N2806, N1171);
and AND3 (N6953, N6952, N5497, N6423);
or OR3 (N6954, N6949, N3332, N4688);
not NOT1 (N6955, N6954);
not NOT1 (N6956, N6944);
buf BUF1 (N6957, N6950);
or OR4 (N6958, N6953, N926, N2706, N1097);
buf BUF1 (N6959, N6958);
nor NOR2 (N6960, N6932, N3866);
xor XOR2 (N6961, N6955, N4555);
xor XOR2 (N6962, N6946, N3362);
or OR2 (N6963, N6960, N5984);
buf BUF1 (N6964, N6961);
or OR2 (N6965, N6937, N2327);
xor XOR2 (N6966, N6962, N1322);
and AND4 (N6967, N6940, N2050, N1444, N6870);
not NOT1 (N6968, N6956);
nand NAND3 (N6969, N6942, N6403, N4248);
xor XOR2 (N6970, N6963, N6556);
not NOT1 (N6971, N6948);
buf BUF1 (N6972, N6957);
and AND4 (N6973, N6959, N6494, N214, N2704);
buf BUF1 (N6974, N6966);
or OR4 (N6975, N6964, N5720, N3838, N6103);
nor NOR3 (N6976, N6973, N4743, N6471);
nand NAND3 (N6977, N6969, N3572, N4793);
and AND2 (N6978, N6971, N4230);
and AND2 (N6979, N6978, N2153);
not NOT1 (N6980, N6975);
or OR2 (N6981, N6968, N2476);
buf BUF1 (N6982, N6979);
nand NAND4 (N6983, N6982, N3776, N3714, N6440);
nor NOR4 (N6984, N6977, N3183, N962, N970);
or OR3 (N6985, N6976, N210, N3577);
xor XOR2 (N6986, N6967, N3713);
and AND3 (N6987, N6972, N4248, N2053);
nand NAND2 (N6988, N6974, N5309);
nor NOR3 (N6989, N6965, N6860, N3394);
not NOT1 (N6990, N6980);
xor XOR2 (N6991, N6990, N4028);
nor NOR3 (N6992, N6970, N6788, N3910);
xor XOR2 (N6993, N6984, N6915);
nand NAND2 (N6994, N6986, N148);
not NOT1 (N6995, N6994);
nand NAND3 (N6996, N6985, N131, N4505);
nand NAND2 (N6997, N6995, N6786);
not NOT1 (N6998, N6983);
buf BUF1 (N6999, N6993);
buf BUF1 (N7000, N6999);
not NOT1 (N7001, N6989);
nor NOR3 (N7002, N6987, N5806, N5330);
or OR2 (N7003, N7001, N6565);
and AND4 (N7004, N6988, N5840, N4457, N5668);
xor XOR2 (N7005, N6992, N2143);
nor NOR4 (N7006, N6998, N1208, N6237, N2932);
not NOT1 (N7007, N7003);
xor XOR2 (N7008, N7005, N3069);
or OR2 (N7009, N7007, N2792);
xor XOR2 (N7010, N7008, N6339);
xor XOR2 (N7011, N7009, N3727);
not NOT1 (N7012, N7000);
buf BUF1 (N7013, N7010);
xor XOR2 (N7014, N6981, N1209);
or OR4 (N7015, N7014, N5812, N2261, N388);
nor NOR3 (N7016, N6996, N3963, N1730);
nor NOR4 (N7017, N7006, N5481, N2871, N2236);
xor XOR2 (N7018, N7016, N1462);
not NOT1 (N7019, N6997);
nand NAND4 (N7020, N7019, N4154, N5557, N670);
and AND4 (N7021, N7017, N3242, N3774, N4021);
nor NOR4 (N7022, N7011, N5300, N4932, N507);
or OR4 (N7023, N7020, N1763, N4433, N3082);
xor XOR2 (N7024, N7015, N5548);
and AND2 (N7025, N7021, N736);
nor NOR4 (N7026, N7018, N5490, N1809, N3401);
not NOT1 (N7027, N7022);
xor XOR2 (N7028, N7012, N2550);
xor XOR2 (N7029, N7026, N813);
not NOT1 (N7030, N6991);
not NOT1 (N7031, N7023);
not NOT1 (N7032, N7002);
buf BUF1 (N7033, N7004);
or OR2 (N7034, N7032, N1000);
and AND3 (N7035, N7031, N3453, N6541);
nand NAND2 (N7036, N7027, N1552);
xor XOR2 (N7037, N7013, N2118);
nor NOR4 (N7038, N7034, N6039, N4410, N1190);
nand NAND2 (N7039, N7028, N3681);
and AND2 (N7040, N7039, N1192);
nor NOR3 (N7041, N7033, N4409, N2319);
xor XOR2 (N7042, N7036, N774);
not NOT1 (N7043, N7042);
xor XOR2 (N7044, N7024, N6216);
buf BUF1 (N7045, N7025);
xor XOR2 (N7046, N7035, N5690);
not NOT1 (N7047, N7045);
and AND4 (N7048, N7038, N5873, N1427, N4743);
and AND3 (N7049, N7043, N5363, N2890);
xor XOR2 (N7050, N7046, N2164);
and AND4 (N7051, N7040, N1737, N4923, N6135);
buf BUF1 (N7052, N7051);
and AND3 (N7053, N7052, N5099, N6173);
or OR3 (N7054, N7048, N5773, N211);
xor XOR2 (N7055, N7030, N5765);
xor XOR2 (N7056, N7050, N5353);
xor XOR2 (N7057, N7056, N5701);
not NOT1 (N7058, N7049);
or OR4 (N7059, N7055, N5173, N3189, N2118);
nor NOR2 (N7060, N7029, N389);
nand NAND2 (N7061, N7060, N4655);
xor XOR2 (N7062, N7058, N3667);
nand NAND4 (N7063, N7061, N5482, N819, N2364);
not NOT1 (N7064, N7062);
xor XOR2 (N7065, N7037, N2045);
buf BUF1 (N7066, N7041);
xor XOR2 (N7067, N7059, N7022);
nor NOR2 (N7068, N7054, N4704);
xor XOR2 (N7069, N7057, N5825);
and AND3 (N7070, N7066, N6782, N6622);
buf BUF1 (N7071, N7053);
not NOT1 (N7072, N7070);
not NOT1 (N7073, N7044);
and AND3 (N7074, N7071, N5519, N1363);
buf BUF1 (N7075, N7072);
xor XOR2 (N7076, N7069, N154);
nor NOR3 (N7077, N7067, N3513, N1533);
buf BUF1 (N7078, N7063);
and AND2 (N7079, N7077, N5977);
nand NAND2 (N7080, N7073, N652);
xor XOR2 (N7081, N7080, N6856);
not NOT1 (N7082, N7074);
nor NOR4 (N7083, N7076, N6836, N4810, N387);
nand NAND2 (N7084, N7078, N7073);
nor NOR3 (N7085, N7083, N4361, N595);
xor XOR2 (N7086, N7082, N122);
xor XOR2 (N7087, N7086, N1295);
not NOT1 (N7088, N7087);
not NOT1 (N7089, N7075);
nor NOR2 (N7090, N7089, N1423);
buf BUF1 (N7091, N7079);
and AND4 (N7092, N7091, N6508, N2602, N5028);
xor XOR2 (N7093, N7064, N7013);
or OR3 (N7094, N7068, N3805, N4147);
nand NAND3 (N7095, N7065, N4116, N2011);
nand NAND4 (N7096, N7094, N814, N4946, N5832);
buf BUF1 (N7097, N7095);
buf BUF1 (N7098, N7090);
and AND3 (N7099, N7047, N3751, N5179);
not NOT1 (N7100, N7093);
buf BUF1 (N7101, N7088);
not NOT1 (N7102, N7099);
and AND4 (N7103, N7100, N3634, N2907, N4077);
nor NOR2 (N7104, N7096, N6505);
xor XOR2 (N7105, N7098, N5556);
and AND2 (N7106, N7101, N4281);
or OR4 (N7107, N7104, N6836, N4218, N1111);
not NOT1 (N7108, N7097);
and AND3 (N7109, N7103, N1807, N5195);
buf BUF1 (N7110, N7109);
not NOT1 (N7111, N7105);
and AND4 (N7112, N7106, N5516, N599, N3839);
buf BUF1 (N7113, N7084);
nand NAND3 (N7114, N7113, N1117, N3746);
xor XOR2 (N7115, N7092, N2260);
nor NOR3 (N7116, N7114, N2421, N5630);
xor XOR2 (N7117, N7085, N1091);
or OR4 (N7118, N7108, N5712, N2664, N2945);
not NOT1 (N7119, N7116);
xor XOR2 (N7120, N7115, N548);
buf BUF1 (N7121, N7120);
xor XOR2 (N7122, N7118, N4020);
not NOT1 (N7123, N7081);
buf BUF1 (N7124, N7123);
buf BUF1 (N7125, N7117);
or OR3 (N7126, N7107, N4484, N1360);
and AND2 (N7127, N7124, N2369);
and AND2 (N7128, N7125, N5796);
not NOT1 (N7129, N7122);
and AND4 (N7130, N7126, N173, N6380, N6785);
xor XOR2 (N7131, N7111, N5204);
and AND3 (N7132, N7112, N6609, N2026);
or OR4 (N7133, N7128, N2546, N4724, N6310);
xor XOR2 (N7134, N7110, N426);
and AND2 (N7135, N7131, N4412);
buf BUF1 (N7136, N7129);
xor XOR2 (N7137, N7135, N6208);
and AND2 (N7138, N7102, N7099);
and AND4 (N7139, N7130, N5273, N6184, N2450);
nand NAND3 (N7140, N7133, N4651, N3833);
or OR3 (N7141, N7132, N2138, N51);
or OR3 (N7142, N7119, N5052, N352);
nand NAND2 (N7143, N7142, N3458);
and AND3 (N7144, N7127, N4560, N626);
nand NAND2 (N7145, N7137, N577);
or OR4 (N7146, N7145, N5333, N4510, N6715);
nand NAND2 (N7147, N7136, N2377);
not NOT1 (N7148, N7146);
or OR4 (N7149, N7121, N5604, N5314, N1954);
or OR2 (N7150, N7149, N4009);
xor XOR2 (N7151, N7148, N835);
buf BUF1 (N7152, N7140);
and AND4 (N7153, N7141, N1907, N1206, N3394);
buf BUF1 (N7154, N7139);
and AND2 (N7155, N7153, N5567);
not NOT1 (N7156, N7138);
buf BUF1 (N7157, N7152);
nand NAND3 (N7158, N7144, N5, N3452);
and AND2 (N7159, N7147, N2049);
nand NAND3 (N7160, N7150, N3494, N5144);
buf BUF1 (N7161, N7143);
nand NAND3 (N7162, N7160, N2679, N1281);
nand NAND4 (N7163, N7159, N127, N5992, N734);
xor XOR2 (N7164, N7154, N783);
nand NAND2 (N7165, N7162, N4918);
not NOT1 (N7166, N7158);
and AND3 (N7167, N7166, N4439, N6400);
or OR2 (N7168, N7161, N2233);
nand NAND4 (N7169, N7156, N6763, N3256, N3177);
xor XOR2 (N7170, N7164, N2855);
xor XOR2 (N7171, N7151, N2362);
or OR3 (N7172, N7168, N466, N928);
or OR2 (N7173, N7171, N6174);
and AND3 (N7174, N7172, N2204, N891);
nand NAND3 (N7175, N7155, N6478, N767);
or OR2 (N7176, N7157, N2855);
xor XOR2 (N7177, N7134, N209);
and AND2 (N7178, N7167, N2067);
not NOT1 (N7179, N7175);
and AND4 (N7180, N7179, N1662, N459, N5242);
buf BUF1 (N7181, N7165);
and AND4 (N7182, N7170, N836, N1913, N6837);
xor XOR2 (N7183, N7163, N4331);
buf BUF1 (N7184, N7174);
buf BUF1 (N7185, N7173);
or OR4 (N7186, N7177, N730, N1939, N6825);
nor NOR2 (N7187, N7169, N524);
nand NAND3 (N7188, N7180, N2256, N3753);
buf BUF1 (N7189, N7188);
nand NAND4 (N7190, N7182, N1052, N1588, N137);
or OR4 (N7191, N7185, N4762, N882, N4582);
not NOT1 (N7192, N7176);
xor XOR2 (N7193, N7184, N4145);
and AND3 (N7194, N7186, N1547, N5374);
and AND3 (N7195, N7187, N6016, N5010);
nor NOR4 (N7196, N7183, N7025, N3668, N4550);
xor XOR2 (N7197, N7190, N7007);
xor XOR2 (N7198, N7189, N2243);
nor NOR4 (N7199, N7196, N3005, N5385, N2667);
not NOT1 (N7200, N7178);
nand NAND2 (N7201, N7200, N6409);
and AND3 (N7202, N7199, N3539, N3943);
and AND3 (N7203, N7197, N4796, N1511);
xor XOR2 (N7204, N7193, N5988);
buf BUF1 (N7205, N7181);
or OR4 (N7206, N7194, N883, N1495, N3260);
and AND3 (N7207, N7192, N6544, N3847);
and AND2 (N7208, N7202, N3585);
nand NAND4 (N7209, N7205, N2223, N2228, N5833);
nor NOR4 (N7210, N7201, N2741, N3391, N6763);
nor NOR2 (N7211, N7206, N4545);
not NOT1 (N7212, N7203);
buf BUF1 (N7213, N7211);
xor XOR2 (N7214, N7209, N4733);
not NOT1 (N7215, N7208);
and AND4 (N7216, N7215, N5498, N4653, N4356);
not NOT1 (N7217, N7213);
xor XOR2 (N7218, N7216, N3030);
and AND2 (N7219, N7214, N3237);
or OR2 (N7220, N7218, N4322);
xor XOR2 (N7221, N7212, N367);
or OR3 (N7222, N7219, N1126, N5530);
and AND2 (N7223, N7191, N4106);
xor XOR2 (N7224, N7207, N6824);
nand NAND2 (N7225, N7198, N7056);
nand NAND2 (N7226, N7204, N6079);
xor XOR2 (N7227, N7210, N4247);
xor XOR2 (N7228, N7220, N3834);
not NOT1 (N7229, N7224);
buf BUF1 (N7230, N7221);
buf BUF1 (N7231, N7226);
xor XOR2 (N7232, N7222, N6666);
nand NAND2 (N7233, N7227, N1628);
not NOT1 (N7234, N7231);
nor NOR4 (N7235, N7225, N5154, N498, N2374);
nand NAND3 (N7236, N7232, N6799, N4484);
and AND3 (N7237, N7217, N5145, N3790);
or OR2 (N7238, N7235, N6624);
nand NAND4 (N7239, N7234, N4985, N3874, N2409);
xor XOR2 (N7240, N7239, N3920);
xor XOR2 (N7241, N7229, N4315);
or OR4 (N7242, N7228, N2388, N3554, N2703);
xor XOR2 (N7243, N7242, N5358);
buf BUF1 (N7244, N7243);
or OR3 (N7245, N7223, N6410, N5356);
buf BUF1 (N7246, N7230);
or OR3 (N7247, N7236, N2305, N53);
or OR4 (N7248, N7247, N1104, N3147, N1696);
or OR2 (N7249, N7245, N2212);
nand NAND4 (N7250, N7248, N867, N3284, N3082);
and AND2 (N7251, N7237, N6873);
buf BUF1 (N7252, N7233);
and AND4 (N7253, N7251, N1259, N3156, N3445);
and AND2 (N7254, N7250, N5059);
and AND2 (N7255, N7252, N4755);
buf BUF1 (N7256, N7246);
not NOT1 (N7257, N7254);
or OR2 (N7258, N7255, N5388);
buf BUF1 (N7259, N7258);
or OR3 (N7260, N7240, N4783, N639);
buf BUF1 (N7261, N7257);
nor NOR4 (N7262, N7260, N1087, N5751, N1006);
or OR2 (N7263, N7195, N2298);
not NOT1 (N7264, N7238);
not NOT1 (N7265, N7262);
xor XOR2 (N7266, N7265, N3545);
and AND4 (N7267, N7264, N3580, N6125, N5932);
nand NAND2 (N7268, N7241, N5886);
and AND2 (N7269, N7253, N4473);
nor NOR3 (N7270, N7268, N3480, N4741);
nor NOR2 (N7271, N7263, N5431);
nand NAND4 (N7272, N7270, N6632, N4472, N2058);
nand NAND4 (N7273, N7244, N6861, N4315, N5979);
buf BUF1 (N7274, N7249);
buf BUF1 (N7275, N7261);
nand NAND3 (N7276, N7273, N2758, N3824);
nor NOR4 (N7277, N7267, N1397, N5972, N5977);
xor XOR2 (N7278, N7266, N4410);
not NOT1 (N7279, N7278);
and AND4 (N7280, N7256, N3211, N271, N1346);
or OR3 (N7281, N7275, N2964, N1618);
nand NAND2 (N7282, N7269, N4742);
nand NAND4 (N7283, N7272, N248, N2979, N1475);
not NOT1 (N7284, N7279);
nor NOR3 (N7285, N7276, N5796, N5543);
buf BUF1 (N7286, N7285);
or OR4 (N7287, N7274, N2064, N6364, N537);
or OR3 (N7288, N7284, N847, N1243);
nand NAND2 (N7289, N7286, N5508);
not NOT1 (N7290, N7277);
not NOT1 (N7291, N7288);
xor XOR2 (N7292, N7290, N2147);
xor XOR2 (N7293, N7271, N7167);
nor NOR3 (N7294, N7283, N4156, N6434);
not NOT1 (N7295, N7289);
nor NOR3 (N7296, N7292, N59, N7182);
or OR2 (N7297, N7280, N1735);
or OR3 (N7298, N7297, N4635, N7195);
nand NAND2 (N7299, N7298, N4045);
buf BUF1 (N7300, N7299);
xor XOR2 (N7301, N7281, N2689);
buf BUF1 (N7302, N7287);
or OR3 (N7303, N7282, N1001, N6169);
not NOT1 (N7304, N7293);
xor XOR2 (N7305, N7302, N7216);
nor NOR4 (N7306, N7300, N758, N384, N4533);
buf BUF1 (N7307, N7259);
nor NOR3 (N7308, N7296, N512, N299);
and AND4 (N7309, N7308, N1472, N6555, N4551);
or OR3 (N7310, N7294, N6843, N3675);
nand NAND3 (N7311, N7309, N956, N4322);
nand NAND3 (N7312, N7304, N1951, N813);
or OR4 (N7313, N7295, N2248, N5592, N2712);
nor NOR4 (N7314, N7303, N1814, N3339, N7149);
not NOT1 (N7315, N7301);
nand NAND4 (N7316, N7314, N2339, N6005, N2685);
not NOT1 (N7317, N7315);
and AND4 (N7318, N7291, N2514, N4763, N5705);
nor NOR3 (N7319, N7311, N3038, N3328);
and AND3 (N7320, N7317, N3118, N1314);
not NOT1 (N7321, N7307);
nand NAND4 (N7322, N7320, N1994, N3704, N362);
and AND3 (N7323, N7306, N2993, N6730);
xor XOR2 (N7324, N7312, N3739);
nor NOR4 (N7325, N7310, N1279, N201, N1031);
xor XOR2 (N7326, N7319, N854);
nor NOR2 (N7327, N7313, N4758);
not NOT1 (N7328, N7318);
or OR3 (N7329, N7316, N1133, N716);
buf BUF1 (N7330, N7323);
and AND3 (N7331, N7321, N4509, N632);
not NOT1 (N7332, N7327);
buf BUF1 (N7333, N7329);
nand NAND2 (N7334, N7332, N5925);
nand NAND3 (N7335, N7322, N6742, N5881);
and AND2 (N7336, N7331, N3);
and AND2 (N7337, N7330, N7313);
buf BUF1 (N7338, N7335);
not NOT1 (N7339, N7338);
nand NAND2 (N7340, N7326, N825);
not NOT1 (N7341, N7336);
and AND4 (N7342, N7334, N2744, N74, N2796);
nand NAND4 (N7343, N7340, N1109, N2745, N3309);
buf BUF1 (N7344, N7305);
buf BUF1 (N7345, N7344);
and AND3 (N7346, N7328, N4051, N181);
nand NAND4 (N7347, N7346, N2146, N4264, N1086);
not NOT1 (N7348, N7339);
nor NOR2 (N7349, N7324, N1314);
nor NOR3 (N7350, N7343, N5023, N3067);
buf BUF1 (N7351, N7341);
nand NAND3 (N7352, N7342, N4784, N5832);
and AND4 (N7353, N7351, N3668, N3476, N1932);
buf BUF1 (N7354, N7352);
nand NAND4 (N7355, N7350, N2415, N4739, N1620);
xor XOR2 (N7356, N7333, N4337);
nor NOR4 (N7357, N7345, N700, N3222, N1686);
xor XOR2 (N7358, N7353, N822);
not NOT1 (N7359, N7354);
nor NOR2 (N7360, N7358, N5913);
and AND2 (N7361, N7347, N971);
buf BUF1 (N7362, N7356);
buf BUF1 (N7363, N7359);
buf BUF1 (N7364, N7362);
xor XOR2 (N7365, N7337, N4859);
not NOT1 (N7366, N7363);
or OR3 (N7367, N7349, N257, N6050);
nand NAND2 (N7368, N7364, N1228);
not NOT1 (N7369, N7365);
not NOT1 (N7370, N7357);
nand NAND4 (N7371, N7325, N940, N6400, N6650);
nor NOR3 (N7372, N7367, N2201, N1458);
and AND4 (N7373, N7360, N3647, N351, N7103);
not NOT1 (N7374, N7366);
buf BUF1 (N7375, N7373);
not NOT1 (N7376, N7374);
and AND3 (N7377, N7376, N454, N3332);
nor NOR3 (N7378, N7361, N489, N637);
or OR2 (N7379, N7377, N3174);
not NOT1 (N7380, N7348);
or OR2 (N7381, N7371, N2736);
nand NAND2 (N7382, N7378, N4163);
or OR4 (N7383, N7372, N5029, N5895, N3888);
and AND3 (N7384, N7379, N5949, N4876);
nand NAND2 (N7385, N7368, N6989);
not NOT1 (N7386, N7370);
nand NAND4 (N7387, N7385, N4091, N3794, N1385);
or OR3 (N7388, N7383, N3687, N6521);
nand NAND4 (N7389, N7355, N5699, N1768, N2273);
nor NOR2 (N7390, N7384, N1531);
or OR2 (N7391, N7387, N1967);
xor XOR2 (N7392, N7388, N3152);
nand NAND3 (N7393, N7375, N2932, N4870);
xor XOR2 (N7394, N7391, N4100);
buf BUF1 (N7395, N7369);
buf BUF1 (N7396, N7394);
or OR3 (N7397, N7382, N4888, N6424);
nor NOR3 (N7398, N7390, N1132, N3016);
nand NAND4 (N7399, N7398, N4490, N6942, N733);
xor XOR2 (N7400, N7381, N2075);
and AND2 (N7401, N7395, N3082);
or OR2 (N7402, N7389, N6872);
or OR3 (N7403, N7401, N4222, N6112);
and AND2 (N7404, N7397, N1618);
or OR3 (N7405, N7399, N26, N3066);
buf BUF1 (N7406, N7400);
or OR3 (N7407, N7393, N2533, N2811);
and AND2 (N7408, N7380, N5079);
nor NOR3 (N7409, N7405, N5108, N6400);
nand NAND3 (N7410, N7386, N4432, N2502);
not NOT1 (N7411, N7403);
or OR3 (N7412, N7396, N2623, N1573);
nor NOR3 (N7413, N7402, N4511, N6524);
nand NAND3 (N7414, N7412, N6610, N4641);
xor XOR2 (N7415, N7410, N575);
not NOT1 (N7416, N7414);
buf BUF1 (N7417, N7415);
xor XOR2 (N7418, N7409, N6045);
and AND4 (N7419, N7407, N452, N7261, N7187);
not NOT1 (N7420, N7417);
nand NAND4 (N7421, N7420, N4207, N6338, N3384);
nor NOR3 (N7422, N7418, N2607, N5440);
xor XOR2 (N7423, N7404, N7225);
or OR2 (N7424, N7416, N6047);
and AND3 (N7425, N7408, N46, N5747);
not NOT1 (N7426, N7419);
or OR4 (N7427, N7425, N3139, N3606, N6524);
and AND3 (N7428, N7406, N3668, N1372);
buf BUF1 (N7429, N7413);
not NOT1 (N7430, N7426);
xor XOR2 (N7431, N7421, N6407);
nor NOR2 (N7432, N7430, N826);
not NOT1 (N7433, N7428);
nor NOR3 (N7434, N7392, N4011, N7297);
or OR3 (N7435, N7422, N1482, N1445);
buf BUF1 (N7436, N7411);
or OR2 (N7437, N7436, N3204);
xor XOR2 (N7438, N7424, N3136);
nor NOR4 (N7439, N7435, N1738, N4862, N145);
and AND2 (N7440, N7423, N5921);
xor XOR2 (N7441, N7427, N101);
nor NOR3 (N7442, N7429, N6872, N7363);
and AND2 (N7443, N7438, N1927);
buf BUF1 (N7444, N7442);
not NOT1 (N7445, N7437);
buf BUF1 (N7446, N7431);
xor XOR2 (N7447, N7439, N6874);
nand NAND4 (N7448, N7443, N6545, N5070, N4991);
and AND3 (N7449, N7447, N5313, N4230);
and AND4 (N7450, N7445, N3881, N5079, N5358);
and AND3 (N7451, N7450, N6648, N6435);
nor NOR3 (N7452, N7446, N3078, N6094);
not NOT1 (N7453, N7440);
and AND4 (N7454, N7449, N5028, N3660, N711);
xor XOR2 (N7455, N7451, N3993);
buf BUF1 (N7456, N7432);
xor XOR2 (N7457, N7454, N5122);
and AND4 (N7458, N7455, N4540, N7423, N2917);
buf BUF1 (N7459, N7452);
nor NOR4 (N7460, N7448, N747, N6822, N6896);
nor NOR3 (N7461, N7444, N1132, N4598);
buf BUF1 (N7462, N7458);
or OR4 (N7463, N7441, N6878, N7334, N5810);
nor NOR3 (N7464, N7434, N2642, N1769);
xor XOR2 (N7465, N7463, N7303);
nand NAND4 (N7466, N7460, N3318, N3354, N3909);
buf BUF1 (N7467, N7462);
nand NAND4 (N7468, N7465, N1751, N1926, N3669);
and AND3 (N7469, N7461, N6147, N4220);
or OR3 (N7470, N7469, N2155, N2289);
buf BUF1 (N7471, N7456);
or OR3 (N7472, N7464, N2324, N2102);
nand NAND2 (N7473, N7472, N997);
buf BUF1 (N7474, N7433);
or OR3 (N7475, N7457, N5743, N3201);
not NOT1 (N7476, N7470);
xor XOR2 (N7477, N7466, N3882);
or OR3 (N7478, N7453, N6868, N617);
and AND2 (N7479, N7474, N453);
not NOT1 (N7480, N7467);
nor NOR2 (N7481, N7478, N4705);
and AND4 (N7482, N7476, N1968, N3187, N2617);
not NOT1 (N7483, N7482);
or OR4 (N7484, N7459, N3648, N5626, N4975);
or OR4 (N7485, N7479, N3236, N6648, N6008);
nor NOR4 (N7486, N7483, N2553, N172, N6588);
nor NOR3 (N7487, N7471, N2553, N3097);
nor NOR3 (N7488, N7481, N7101, N4526);
not NOT1 (N7489, N7480);
not NOT1 (N7490, N7468);
or OR4 (N7491, N7488, N3843, N587, N5827);
nand NAND2 (N7492, N7477, N2037);
xor XOR2 (N7493, N7484, N6924);
or OR4 (N7494, N7473, N46, N7101, N4391);
xor XOR2 (N7495, N7492, N1947);
nand NAND4 (N7496, N7485, N124, N6367, N6532);
nand NAND4 (N7497, N7475, N5531, N1352, N6611);
buf BUF1 (N7498, N7497);
buf BUF1 (N7499, N7489);
not NOT1 (N7500, N7487);
nand NAND3 (N7501, N7499, N6911, N6355);
nand NAND2 (N7502, N7491, N3850);
buf BUF1 (N7503, N7501);
buf BUF1 (N7504, N7503);
nand NAND3 (N7505, N7496, N226, N1950);
or OR2 (N7506, N7495, N1314);
xor XOR2 (N7507, N7490, N1292);
buf BUF1 (N7508, N7493);
buf BUF1 (N7509, N7498);
or OR4 (N7510, N7508, N6459, N7110, N4478);
nor NOR3 (N7511, N7506, N1243, N6820);
not NOT1 (N7512, N7500);
nor NOR3 (N7513, N7504, N2708, N1279);
buf BUF1 (N7514, N7486);
and AND4 (N7515, N7507, N6905, N3035, N1281);
xor XOR2 (N7516, N7511, N7419);
not NOT1 (N7517, N7494);
or OR2 (N7518, N7510, N5548);
buf BUF1 (N7519, N7518);
not NOT1 (N7520, N7519);
or OR3 (N7521, N7513, N5890, N4223);
nand NAND3 (N7522, N7520, N3653, N5242);
and AND2 (N7523, N7515, N738);
xor XOR2 (N7524, N7505, N12);
or OR4 (N7525, N7521, N2497, N5456, N4237);
or OR2 (N7526, N7524, N6813);
nor NOR2 (N7527, N7516, N3121);
and AND3 (N7528, N7502, N7497, N4202);
not NOT1 (N7529, N7525);
nor NOR4 (N7530, N7517, N1294, N4946, N6068);
and AND4 (N7531, N7526, N3518, N2871, N118);
nor NOR4 (N7532, N7527, N3025, N1598, N411);
nor NOR4 (N7533, N7529, N1613, N5180, N5084);
nand NAND4 (N7534, N7528, N375, N4641, N6206);
or OR2 (N7535, N7532, N4632);
nor NOR2 (N7536, N7514, N5777);
xor XOR2 (N7537, N7534, N6936);
or OR4 (N7538, N7509, N848, N3669, N2454);
buf BUF1 (N7539, N7535);
or OR3 (N7540, N7512, N1003, N2449);
nand NAND4 (N7541, N7536, N3375, N1230, N376);
buf BUF1 (N7542, N7522);
not NOT1 (N7543, N7539);
and AND3 (N7544, N7533, N299, N6479);
not NOT1 (N7545, N7537);
buf BUF1 (N7546, N7538);
nand NAND3 (N7547, N7523, N2463, N939);
nor NOR2 (N7548, N7531, N3738);
nand NAND2 (N7549, N7545, N436);
and AND2 (N7550, N7542, N2737);
xor XOR2 (N7551, N7541, N6756);
xor XOR2 (N7552, N7540, N4041);
buf BUF1 (N7553, N7544);
and AND2 (N7554, N7550, N6446);
nor NOR4 (N7555, N7543, N803, N250, N3398);
and AND2 (N7556, N7551, N6933);
xor XOR2 (N7557, N7530, N6829);
xor XOR2 (N7558, N7555, N5412);
xor XOR2 (N7559, N7546, N615);
nand NAND4 (N7560, N7557, N4601, N2370, N159);
xor XOR2 (N7561, N7549, N7075);
xor XOR2 (N7562, N7558, N3354);
xor XOR2 (N7563, N7553, N2800);
nor NOR3 (N7564, N7561, N4637, N6111);
or OR3 (N7565, N7556, N844, N1646);
not NOT1 (N7566, N7554);
and AND4 (N7567, N7559, N1359, N2717, N437);
buf BUF1 (N7568, N7560);
buf BUF1 (N7569, N7568);
xor XOR2 (N7570, N7567, N4852);
not NOT1 (N7571, N7570);
nand NAND2 (N7572, N7548, N2658);
or OR4 (N7573, N7562, N3572, N1637, N3737);
nand NAND4 (N7574, N7565, N5578, N1346, N3484);
not NOT1 (N7575, N7566);
not NOT1 (N7576, N7572);
xor XOR2 (N7577, N7571, N4437);
or OR4 (N7578, N7564, N7212, N3140, N4000);
buf BUF1 (N7579, N7569);
and AND3 (N7580, N7576, N4361, N6318);
nor NOR3 (N7581, N7578, N865, N89);
nor NOR4 (N7582, N7581, N3311, N670, N3675);
or OR2 (N7583, N7573, N235);
nor NOR3 (N7584, N7577, N5197, N5585);
not NOT1 (N7585, N7579);
nand NAND4 (N7586, N7563, N2903, N4237, N3390);
or OR4 (N7587, N7583, N303, N2068, N2637);
nor NOR4 (N7588, N7586, N545, N6699, N5387);
xor XOR2 (N7589, N7588, N377);
and AND2 (N7590, N7547, N7184);
not NOT1 (N7591, N7582);
nor NOR3 (N7592, N7574, N5398, N3914);
xor XOR2 (N7593, N7591, N826);
not NOT1 (N7594, N7575);
and AND4 (N7595, N7584, N2555, N4786, N2086);
and AND3 (N7596, N7587, N3699, N3679);
xor XOR2 (N7597, N7580, N2082);
nand NAND4 (N7598, N7592, N240, N3202, N5724);
not NOT1 (N7599, N7594);
or OR4 (N7600, N7585, N1670, N5397, N3040);
xor XOR2 (N7601, N7593, N6091);
buf BUF1 (N7602, N7589);
nand NAND2 (N7603, N7590, N2771);
and AND3 (N7604, N7596, N71, N5823);
or OR3 (N7605, N7597, N873, N282);
and AND3 (N7606, N7602, N616, N582);
nor NOR4 (N7607, N7604, N807, N4936, N4064);
not NOT1 (N7608, N7599);
nand NAND2 (N7609, N7595, N1528);
and AND2 (N7610, N7605, N1269);
nand NAND4 (N7611, N7607, N6701, N6795, N1206);
nand NAND2 (N7612, N7600, N4333);
xor XOR2 (N7613, N7603, N7024);
nand NAND3 (N7614, N7611, N4817, N2976);
nor NOR2 (N7615, N7614, N6391);
xor XOR2 (N7616, N7598, N312);
xor XOR2 (N7617, N7616, N2144);
nor NOR4 (N7618, N7610, N1819, N7005, N3730);
not NOT1 (N7619, N7552);
nand NAND2 (N7620, N7609, N7589);
not NOT1 (N7621, N7617);
and AND2 (N7622, N7601, N50);
nor NOR4 (N7623, N7618, N2775, N6961, N2011);
buf BUF1 (N7624, N7621);
or OR4 (N7625, N7613, N4401, N1744, N4306);
not NOT1 (N7626, N7608);
nand NAND4 (N7627, N7615, N7534, N3161, N3670);
nor NOR2 (N7628, N7620, N4271);
nor NOR3 (N7629, N7606, N1719, N4143);
nand NAND4 (N7630, N7625, N5143, N4498, N3730);
nand NAND4 (N7631, N7623, N2045, N1266, N1130);
not NOT1 (N7632, N7626);
xor XOR2 (N7633, N7629, N4872);
not NOT1 (N7634, N7632);
or OR2 (N7635, N7628, N1169);
nand NAND4 (N7636, N7633, N7477, N413, N5583);
nand NAND3 (N7637, N7636, N2467, N4048);
not NOT1 (N7638, N7624);
or OR4 (N7639, N7612, N2878, N44, N3680);
nand NAND3 (N7640, N7637, N7327, N6096);
or OR3 (N7641, N7639, N615, N4670);
nor NOR4 (N7642, N7622, N7460, N4349, N5430);
or OR3 (N7643, N7627, N239, N4136);
or OR2 (N7644, N7631, N3032);
buf BUF1 (N7645, N7634);
buf BUF1 (N7646, N7644);
not NOT1 (N7647, N7646);
and AND4 (N7648, N7635, N401, N2181, N5511);
nor NOR3 (N7649, N7643, N719, N7564);
buf BUF1 (N7650, N7630);
buf BUF1 (N7651, N7650);
xor XOR2 (N7652, N7638, N2261);
or OR4 (N7653, N7619, N1509, N4974, N575);
nand NAND2 (N7654, N7647, N4587);
not NOT1 (N7655, N7651);
nor NOR2 (N7656, N7653, N3323);
and AND3 (N7657, N7656, N6065, N1373);
xor XOR2 (N7658, N7657, N6191);
buf BUF1 (N7659, N7645);
buf BUF1 (N7660, N7659);
not NOT1 (N7661, N7648);
nor NOR2 (N7662, N7640, N2320);
buf BUF1 (N7663, N7649);
xor XOR2 (N7664, N7642, N6508);
nor NOR2 (N7665, N7641, N7343);
xor XOR2 (N7666, N7665, N6311);
or OR2 (N7667, N7660, N3757);
nand NAND2 (N7668, N7658, N95);
nand NAND4 (N7669, N7652, N4733, N925, N7216);
and AND3 (N7670, N7668, N1086, N3816);
nand NAND3 (N7671, N7664, N1197, N6046);
not NOT1 (N7672, N7662);
xor XOR2 (N7673, N7672, N5739);
nand NAND3 (N7674, N7669, N269, N7055);
xor XOR2 (N7675, N7671, N6213);
buf BUF1 (N7676, N7670);
not NOT1 (N7677, N7676);
and AND4 (N7678, N7654, N5965, N2846, N659);
nand NAND3 (N7679, N7666, N2683, N284);
or OR3 (N7680, N7661, N5360, N4517);
nand NAND3 (N7681, N7655, N1486, N2116);
not NOT1 (N7682, N7663);
buf BUF1 (N7683, N7679);
and AND3 (N7684, N7674, N4538, N1998);
or OR2 (N7685, N7682, N1103);
buf BUF1 (N7686, N7673);
buf BUF1 (N7687, N7677);
or OR4 (N7688, N7686, N3290, N7010, N3067);
or OR3 (N7689, N7688, N5318, N4952);
not NOT1 (N7690, N7678);
xor XOR2 (N7691, N7681, N2219);
nand NAND3 (N7692, N7680, N4843, N4322);
or OR4 (N7693, N7687, N1736, N550, N6865);
or OR3 (N7694, N7667, N7045, N1882);
nand NAND4 (N7695, N7685, N5343, N1129, N7492);
or OR4 (N7696, N7693, N1689, N6781, N6787);
nand NAND4 (N7697, N7695, N3597, N6642, N4025);
nor NOR2 (N7698, N7684, N1899);
or OR3 (N7699, N7689, N2489, N312);
xor XOR2 (N7700, N7696, N2298);
xor XOR2 (N7701, N7691, N194);
buf BUF1 (N7702, N7699);
and AND4 (N7703, N7701, N255, N7000, N3619);
nor NOR3 (N7704, N7694, N4753, N56);
and AND4 (N7705, N7702, N2159, N6738, N3628);
nand NAND3 (N7706, N7690, N5642, N5187);
xor XOR2 (N7707, N7675, N1170);
or OR4 (N7708, N7705, N4929, N2215, N4899);
not NOT1 (N7709, N7706);
nor NOR2 (N7710, N7708, N2966);
xor XOR2 (N7711, N7710, N7692);
nor NOR2 (N7712, N259, N4183);
xor XOR2 (N7713, N7703, N1670);
buf BUF1 (N7714, N7704);
buf BUF1 (N7715, N7713);
buf BUF1 (N7716, N7698);
nor NOR2 (N7717, N7712, N316);
and AND4 (N7718, N7707, N2046, N4727, N1713);
or OR2 (N7719, N7718, N3729);
nand NAND3 (N7720, N7715, N5287, N5175);
not NOT1 (N7721, N7697);
nand NAND3 (N7722, N7720, N4603, N1883);
buf BUF1 (N7723, N7716);
or OR4 (N7724, N7714, N5871, N7349, N7593);
buf BUF1 (N7725, N7721);
not NOT1 (N7726, N7709);
nand NAND3 (N7727, N7723, N1785, N6436);
and AND3 (N7728, N7726, N7496, N1607);
nand NAND4 (N7729, N7717, N3212, N4216, N1591);
or OR2 (N7730, N7683, N4704);
buf BUF1 (N7731, N7725);
not NOT1 (N7732, N7724);
not NOT1 (N7733, N7719);
xor XOR2 (N7734, N7728, N2943);
buf BUF1 (N7735, N7732);
not NOT1 (N7736, N7711);
buf BUF1 (N7737, N7722);
or OR3 (N7738, N7734, N5225, N6744);
or OR4 (N7739, N7737, N6357, N2907, N2614);
nor NOR4 (N7740, N7736, N1925, N155, N2083);
or OR2 (N7741, N7738, N4779);
xor XOR2 (N7742, N7741, N374);
nand NAND3 (N7743, N7735, N1892, N1769);
xor XOR2 (N7744, N7727, N6341);
nand NAND4 (N7745, N7739, N2183, N7613, N4672);
or OR3 (N7746, N7743, N5160, N1687);
xor XOR2 (N7747, N7729, N4682);
nor NOR2 (N7748, N7746, N3428);
nand NAND2 (N7749, N7748, N5147);
or OR4 (N7750, N7742, N7321, N1205, N1560);
and AND2 (N7751, N7730, N5616);
xor XOR2 (N7752, N7733, N6317);
or OR4 (N7753, N7745, N5842, N3701, N579);
nand NAND4 (N7754, N7731, N540, N2905, N5583);
or OR3 (N7755, N7753, N3821, N5395);
or OR3 (N7756, N7744, N1523, N1272);
not NOT1 (N7757, N7749);
buf BUF1 (N7758, N7752);
nand NAND4 (N7759, N7740, N4384, N4001, N3847);
nand NAND3 (N7760, N7758, N5477, N1850);
nor NOR3 (N7761, N7750, N5039, N23);
and AND4 (N7762, N7761, N1112, N3463, N4127);
nand NAND4 (N7763, N7747, N7135, N5279, N5115);
nand NAND4 (N7764, N7759, N2339, N5879, N4638);
buf BUF1 (N7765, N7762);
xor XOR2 (N7766, N7760, N4114);
buf BUF1 (N7767, N7754);
xor XOR2 (N7768, N7751, N4865);
nor NOR3 (N7769, N7755, N1872, N6305);
nor NOR2 (N7770, N7764, N7211);
nand NAND2 (N7771, N7767, N4188);
nand NAND2 (N7772, N7757, N7295);
nand NAND4 (N7773, N7768, N1944, N392, N6518);
buf BUF1 (N7774, N7700);
not NOT1 (N7775, N7756);
and AND4 (N7776, N7765, N2759, N186, N3342);
or OR4 (N7777, N7773, N4221, N7390, N2938);
and AND2 (N7778, N7766, N4478);
buf BUF1 (N7779, N7774);
buf BUF1 (N7780, N7777);
or OR4 (N7781, N7769, N2128, N1197, N3786);
and AND4 (N7782, N7763, N364, N3373, N2900);
and AND4 (N7783, N7778, N1101, N7075, N1322);
or OR3 (N7784, N7772, N5255, N6160);
nor NOR2 (N7785, N7784, N4641);
xor XOR2 (N7786, N7775, N6691);
nand NAND3 (N7787, N7781, N3343, N3483);
nor NOR3 (N7788, N7770, N2651, N1972);
nand NAND4 (N7789, N7771, N7756, N2693, N6173);
nor NOR4 (N7790, N7782, N6182, N5916, N6710);
not NOT1 (N7791, N7787);
not NOT1 (N7792, N7783);
and AND3 (N7793, N7789, N4916, N6893);
and AND4 (N7794, N7788, N1120, N1027, N6984);
nand NAND3 (N7795, N7785, N807, N2821);
nand NAND3 (N7796, N7786, N7268, N6375);
and AND2 (N7797, N7795, N624);
buf BUF1 (N7798, N7793);
and AND2 (N7799, N7790, N5618);
xor XOR2 (N7800, N7796, N2290);
and AND4 (N7801, N7780, N7346, N941, N1415);
nor NOR4 (N7802, N7794, N3955, N5659, N5751);
nand NAND4 (N7803, N7798, N3707, N5392, N6236);
nor NOR3 (N7804, N7800, N5985, N3181);
buf BUF1 (N7805, N7803);
nand NAND3 (N7806, N7791, N6288, N5954);
xor XOR2 (N7807, N7799, N6156);
and AND4 (N7808, N7805, N764, N2384, N3314);
buf BUF1 (N7809, N7797);
or OR3 (N7810, N7806, N6750, N6835);
buf BUF1 (N7811, N7776);
buf BUF1 (N7812, N7808);
buf BUF1 (N7813, N7807);
or OR4 (N7814, N7779, N6229, N6996, N4699);
buf BUF1 (N7815, N7813);
nand NAND4 (N7816, N7814, N342, N2028, N2770);
and AND4 (N7817, N7812, N7386, N1487, N5764);
and AND3 (N7818, N7810, N6577, N4148);
or OR2 (N7819, N7801, N1441);
nor NOR4 (N7820, N7792, N456, N1445, N6750);
and AND3 (N7821, N7816, N142, N6099);
and AND2 (N7822, N7809, N624);
nor NOR4 (N7823, N7822, N2989, N4169, N4979);
or OR2 (N7824, N7823, N5875);
nor NOR3 (N7825, N7802, N29, N2221);
or OR3 (N7826, N7815, N1413, N3615);
or OR4 (N7827, N7824, N3557, N102, N4155);
or OR2 (N7828, N7817, N6123);
or OR3 (N7829, N7820, N3215, N5229);
not NOT1 (N7830, N7827);
and AND3 (N7831, N7804, N5095, N346);
buf BUF1 (N7832, N7811);
nor NOR2 (N7833, N7831, N2619);
or OR2 (N7834, N7828, N2882);
and AND4 (N7835, N7825, N3963, N908, N253);
not NOT1 (N7836, N7832);
or OR4 (N7837, N7826, N5692, N3493, N3304);
or OR2 (N7838, N7830, N3051);
xor XOR2 (N7839, N7836, N4176);
buf BUF1 (N7840, N7838);
or OR4 (N7841, N7833, N7325, N6963, N5300);
nand NAND4 (N7842, N7837, N2169, N1488, N7715);
xor XOR2 (N7843, N7841, N7373);
nand NAND2 (N7844, N7842, N5232);
not NOT1 (N7845, N7835);
and AND4 (N7846, N7818, N4849, N5000, N679);
not NOT1 (N7847, N7845);
buf BUF1 (N7848, N7839);
buf BUF1 (N7849, N7847);
buf BUF1 (N7850, N7849);
buf BUF1 (N7851, N7850);
nor NOR2 (N7852, N7840, N1477);
buf BUF1 (N7853, N7846);
not NOT1 (N7854, N7843);
xor XOR2 (N7855, N7834, N6236);
nor NOR2 (N7856, N7829, N7546);
or OR4 (N7857, N7821, N7576, N5225, N5447);
or OR4 (N7858, N7853, N3581, N401, N3398);
buf BUF1 (N7859, N7855);
nor NOR4 (N7860, N7844, N4784, N296, N3213);
or OR4 (N7861, N7819, N4660, N3109, N7729);
buf BUF1 (N7862, N7851);
or OR2 (N7863, N7848, N1161);
nor NOR2 (N7864, N7856, N2623);
nor NOR2 (N7865, N7863, N3684);
nand NAND2 (N7866, N7857, N989);
nor NOR4 (N7867, N7861, N3439, N4051, N3143);
nor NOR3 (N7868, N7860, N5392, N840);
and AND4 (N7869, N7862, N854, N7662, N7428);
or OR4 (N7870, N7852, N814, N7750, N3491);
or OR4 (N7871, N7864, N719, N6809, N2545);
not NOT1 (N7872, N7871);
buf BUF1 (N7873, N7858);
or OR2 (N7874, N7870, N404);
nand NAND2 (N7875, N7867, N7444);
nor NOR4 (N7876, N7865, N6602, N2966, N1176);
not NOT1 (N7877, N7869);
and AND3 (N7878, N7859, N1827, N1212);
not NOT1 (N7879, N7875);
nand NAND4 (N7880, N7854, N7466, N3387, N6553);
nand NAND4 (N7881, N7868, N7079, N4652, N6557);
buf BUF1 (N7882, N7878);
xor XOR2 (N7883, N7881, N2928);
xor XOR2 (N7884, N7883, N5184);
xor XOR2 (N7885, N7879, N3217);
and AND2 (N7886, N7876, N2327);
xor XOR2 (N7887, N7874, N3039);
and AND4 (N7888, N7882, N701, N572, N4059);
xor XOR2 (N7889, N7888, N2647);
not NOT1 (N7890, N7889);
and AND3 (N7891, N7872, N413, N1309);
nor NOR4 (N7892, N7873, N254, N88, N7205);
nor NOR2 (N7893, N7866, N4985);
xor XOR2 (N7894, N7885, N2144);
nand NAND4 (N7895, N7891, N1329, N5027, N1777);
or OR2 (N7896, N7887, N713);
xor XOR2 (N7897, N7886, N1547);
or OR3 (N7898, N7880, N4274, N4821);
or OR3 (N7899, N7877, N4174, N5033);
xor XOR2 (N7900, N7897, N379);
not NOT1 (N7901, N7892);
not NOT1 (N7902, N7894);
nand NAND4 (N7903, N7899, N2181, N6691, N4963);
nor NOR4 (N7904, N7896, N518, N2863, N3382);
buf BUF1 (N7905, N7903);
xor XOR2 (N7906, N7898, N14);
or OR3 (N7907, N7890, N1866, N1598);
nand NAND3 (N7908, N7895, N3660, N2896);
or OR4 (N7909, N7893, N2741, N7425, N7773);
or OR4 (N7910, N7884, N7652, N1713, N2489);
not NOT1 (N7911, N7901);
or OR3 (N7912, N7910, N3781, N6004);
xor XOR2 (N7913, N7908, N4736);
nor NOR4 (N7914, N7909, N6253, N3803, N7088);
not NOT1 (N7915, N7912);
and AND3 (N7916, N7906, N192, N6533);
xor XOR2 (N7917, N7907, N3204);
buf BUF1 (N7918, N7914);
xor XOR2 (N7919, N7917, N531);
nand NAND3 (N7920, N7913, N2740, N3562);
nand NAND4 (N7921, N7919, N1440, N5512, N5722);
xor XOR2 (N7922, N7900, N4561);
xor XOR2 (N7923, N7920, N2394);
and AND2 (N7924, N7916, N1544);
or OR4 (N7925, N7923, N7533, N5767, N6710);
buf BUF1 (N7926, N7918);
or OR2 (N7927, N7921, N6327);
or OR2 (N7928, N7926, N550);
buf BUF1 (N7929, N7925);
nor NOR3 (N7930, N7927, N5219, N6447);
not NOT1 (N7931, N7930);
nand NAND3 (N7932, N7928, N926, N382);
nand NAND2 (N7933, N7929, N2733);
and AND2 (N7934, N7904, N6250);
buf BUF1 (N7935, N7932);
not NOT1 (N7936, N7924);
and AND3 (N7937, N7934, N6052, N2242);
or OR4 (N7938, N7931, N4570, N3760, N4630);
or OR2 (N7939, N7902, N1195);
nor NOR4 (N7940, N7933, N4478, N972, N5999);
and AND4 (N7941, N7915, N6202, N285, N4728);
buf BUF1 (N7942, N7938);
and AND3 (N7943, N7935, N7800, N5583);
not NOT1 (N7944, N7943);
nor NOR2 (N7945, N7944, N1035);
nor NOR4 (N7946, N7922, N2292, N6437, N6716);
buf BUF1 (N7947, N7911);
buf BUF1 (N7948, N7947);
buf BUF1 (N7949, N7939);
nor NOR3 (N7950, N7941, N2651, N7381);
xor XOR2 (N7951, N7942, N571);
not NOT1 (N7952, N7950);
and AND2 (N7953, N7945, N5310);
xor XOR2 (N7954, N7952, N3277);
and AND3 (N7955, N7954, N6738, N6570);
buf BUF1 (N7956, N7953);
nor NOR3 (N7957, N7946, N3122, N7950);
or OR3 (N7958, N7940, N4245, N3380);
or OR3 (N7959, N7951, N2368, N2561);
buf BUF1 (N7960, N7905);
nand NAND4 (N7961, N7955, N3831, N4417, N5547);
xor XOR2 (N7962, N7937, N1289);
nand NAND3 (N7963, N7962, N5887, N177);
xor XOR2 (N7964, N7948, N4093);
xor XOR2 (N7965, N7961, N7300);
and AND2 (N7966, N7956, N4072);
and AND2 (N7967, N7966, N3153);
buf BUF1 (N7968, N7967);
buf BUF1 (N7969, N7959);
and AND4 (N7970, N7964, N2776, N5481, N1996);
nor NOR2 (N7971, N7960, N4343);
xor XOR2 (N7972, N7949, N6878);
or OR3 (N7973, N7972, N3217, N6481);
xor XOR2 (N7974, N7971, N4873);
xor XOR2 (N7975, N7968, N3930);
xor XOR2 (N7976, N7963, N7064);
buf BUF1 (N7977, N7965);
or OR4 (N7978, N7974, N1296, N6742, N7562);
or OR3 (N7979, N7969, N763, N4119);
buf BUF1 (N7980, N7936);
xor XOR2 (N7981, N7957, N3195);
and AND4 (N7982, N7975, N2428, N678, N3537);
nand NAND2 (N7983, N7979, N991);
buf BUF1 (N7984, N7983);
or OR3 (N7985, N7980, N7231, N764);
buf BUF1 (N7986, N7984);
and AND4 (N7987, N7970, N1824, N5387, N7496);
and AND3 (N7988, N7978, N5148, N2533);
nand NAND4 (N7989, N7986, N1174, N751, N6894);
or OR4 (N7990, N7987, N2269, N6879, N6206);
or OR2 (N7991, N7973, N7046);
xor XOR2 (N7992, N7989, N877);
buf BUF1 (N7993, N7981);
nor NOR4 (N7994, N7985, N4860, N6327, N438);
nor NOR4 (N7995, N7958, N2988, N7725, N3380);
nor NOR2 (N7996, N7991, N1472);
not NOT1 (N7997, N7977);
xor XOR2 (N7998, N7992, N7828);
not NOT1 (N7999, N7994);
not NOT1 (N8000, N7990);
nand NAND3 (N8001, N7993, N5550, N7012);
nand NAND2 (N8002, N7998, N7417);
buf BUF1 (N8003, N8000);
or OR4 (N8004, N7976, N6553, N5713, N5371);
or OR4 (N8005, N8003, N7304, N5674, N1971);
nor NOR4 (N8006, N7988, N4822, N7309, N3126);
nor NOR2 (N8007, N7982, N2645);
nand NAND2 (N8008, N8002, N2824);
nand NAND4 (N8009, N7996, N1536, N2266, N5666);
nor NOR2 (N8010, N8006, N501);
or OR2 (N8011, N8001, N3263);
xor XOR2 (N8012, N7997, N6088);
xor XOR2 (N8013, N7999, N6110);
buf BUF1 (N8014, N8013);
nand NAND4 (N8015, N8010, N6865, N6865, N4626);
nor NOR3 (N8016, N8015, N3227, N3242);
not NOT1 (N8017, N8014);
or OR3 (N8018, N7995, N5645, N5143);
nand NAND4 (N8019, N8017, N3053, N6712, N7714);
not NOT1 (N8020, N8004);
and AND3 (N8021, N8007, N5448, N7400);
nor NOR4 (N8022, N8021, N3701, N6707, N7400);
not NOT1 (N8023, N8022);
or OR3 (N8024, N8012, N3482, N1652);
and AND3 (N8025, N8023, N2060, N2730);
xor XOR2 (N8026, N8024, N5045);
xor XOR2 (N8027, N8016, N5262);
or OR4 (N8028, N8026, N914, N5087, N4277);
nand NAND3 (N8029, N8011, N4947, N4685);
nand NAND2 (N8030, N8028, N7337);
not NOT1 (N8031, N8019);
nor NOR4 (N8032, N8020, N6595, N4250, N1494);
nor NOR2 (N8033, N8008, N3563);
xor XOR2 (N8034, N8027, N2692);
nor NOR2 (N8035, N8009, N5598);
nor NOR3 (N8036, N8033, N5323, N544);
buf BUF1 (N8037, N8034);
or OR4 (N8038, N8037, N4499, N1024, N6466);
not NOT1 (N8039, N8032);
nand NAND2 (N8040, N8005, N2764);
nor NOR2 (N8041, N8025, N6712);
and AND3 (N8042, N8031, N7888, N317);
nand NAND2 (N8043, N8039, N2713);
buf BUF1 (N8044, N8040);
buf BUF1 (N8045, N8018);
and AND3 (N8046, N8035, N985, N1210);
or OR3 (N8047, N8036, N7555, N4874);
and AND2 (N8048, N8041, N449);
or OR2 (N8049, N8044, N3828);
nand NAND2 (N8050, N8045, N4118);
not NOT1 (N8051, N8043);
or OR2 (N8052, N8049, N2989);
not NOT1 (N8053, N8048);
and AND4 (N8054, N8046, N4398, N5299, N2445);
not NOT1 (N8055, N8052);
not NOT1 (N8056, N8050);
and AND2 (N8057, N8055, N4867);
nand NAND2 (N8058, N8053, N3564);
not NOT1 (N8059, N8056);
nand NAND3 (N8060, N8058, N4034, N3112);
or OR2 (N8061, N8047, N6973);
not NOT1 (N8062, N8057);
not NOT1 (N8063, N8051);
nand NAND2 (N8064, N8059, N1535);
and AND2 (N8065, N8062, N2093);
and AND4 (N8066, N8030, N7081, N1339, N5327);
buf BUF1 (N8067, N8065);
not NOT1 (N8068, N8038);
nand NAND4 (N8069, N8063, N5420, N1530, N2893);
nor NOR2 (N8070, N8068, N3617);
and AND2 (N8071, N8066, N2071);
or OR2 (N8072, N8054, N5828);
or OR2 (N8073, N8060, N3591);
not NOT1 (N8074, N8067);
nand NAND4 (N8075, N8074, N2896, N7733, N3159);
or OR2 (N8076, N8029, N3412);
nand NAND2 (N8077, N8042, N6122);
not NOT1 (N8078, N8064);
nand NAND3 (N8079, N8072, N3002, N1557);
not NOT1 (N8080, N8075);
or OR2 (N8081, N8078, N6829);
nand NAND2 (N8082, N8080, N4808);
and AND2 (N8083, N8061, N3383);
xor XOR2 (N8084, N8069, N2217);
or OR4 (N8085, N8084, N7962, N6165, N4534);
xor XOR2 (N8086, N8085, N489);
buf BUF1 (N8087, N8070);
or OR4 (N8088, N8079, N4526, N1218, N854);
nor NOR4 (N8089, N8087, N5277, N1972, N2079);
not NOT1 (N8090, N8073);
and AND2 (N8091, N8076, N4127);
xor XOR2 (N8092, N8081, N5787);
buf BUF1 (N8093, N8071);
nand NAND2 (N8094, N8083, N3207);
xor XOR2 (N8095, N8088, N6627);
nand NAND2 (N8096, N8093, N234);
nand NAND3 (N8097, N8096, N5732, N2989);
buf BUF1 (N8098, N8086);
nand NAND3 (N8099, N8082, N985, N7612);
nor NOR2 (N8100, N8092, N4387);
xor XOR2 (N8101, N8097, N1399);
nand NAND3 (N8102, N8077, N4875, N7025);
or OR3 (N8103, N8094, N4586, N6015);
nor NOR2 (N8104, N8091, N730);
nand NAND2 (N8105, N8104, N4201);
buf BUF1 (N8106, N8105);
nor NOR3 (N8107, N8099, N294, N3764);
not NOT1 (N8108, N8107);
nor NOR3 (N8109, N8100, N3313, N172);
nor NOR2 (N8110, N8101, N2122);
or OR2 (N8111, N8102, N6750);
nor NOR2 (N8112, N8106, N6910);
buf BUF1 (N8113, N8090);
or OR4 (N8114, N8112, N7326, N3927, N4740);
buf BUF1 (N8115, N8111);
nand NAND3 (N8116, N8115, N2053, N801);
nand NAND3 (N8117, N8114, N5580, N8001);
or OR2 (N8118, N8113, N1576);
nor NOR3 (N8119, N8098, N3260, N1186);
buf BUF1 (N8120, N8117);
xor XOR2 (N8121, N8109, N7139);
buf BUF1 (N8122, N8121);
xor XOR2 (N8123, N8120, N3108);
or OR4 (N8124, N8089, N2611, N7530, N3762);
and AND2 (N8125, N8118, N5769);
nand NAND2 (N8126, N8116, N5953);
and AND4 (N8127, N8103, N5605, N4251, N5903);
buf BUF1 (N8128, N8124);
nor NOR3 (N8129, N8125, N5292, N7345);
or OR3 (N8130, N8119, N2715, N4879);
xor XOR2 (N8131, N8128, N1534);
xor XOR2 (N8132, N8127, N5601);
nand NAND4 (N8133, N8132, N2760, N1688, N326);
buf BUF1 (N8134, N8126);
nor NOR3 (N8135, N8110, N2012, N3745);
nand NAND4 (N8136, N8133, N5452, N1091, N4275);
nor NOR2 (N8137, N8134, N2220);
buf BUF1 (N8138, N8095);
or OR4 (N8139, N8108, N3203, N7123, N1051);
buf BUF1 (N8140, N8123);
not NOT1 (N8141, N8122);
xor XOR2 (N8142, N8136, N7142);
buf BUF1 (N8143, N8142);
not NOT1 (N8144, N8137);
xor XOR2 (N8145, N8138, N3916);
nor NOR3 (N8146, N8141, N6389, N915);
or OR2 (N8147, N8131, N4655);
xor XOR2 (N8148, N8147, N7986);
nor NOR3 (N8149, N8130, N2657, N1160);
or OR2 (N8150, N8140, N7013);
not NOT1 (N8151, N8135);
nand NAND3 (N8152, N8151, N3164, N937);
buf BUF1 (N8153, N8145);
and AND3 (N8154, N8150, N4530, N7596);
buf BUF1 (N8155, N8146);
and AND4 (N8156, N8153, N4584, N3076, N6705);
nor NOR2 (N8157, N8152, N2898);
nor NOR4 (N8158, N8157, N2780, N4311, N20);
buf BUF1 (N8159, N8154);
nand NAND3 (N8160, N8155, N2616, N2626);
xor XOR2 (N8161, N8156, N2537);
and AND3 (N8162, N8160, N332, N3280);
or OR2 (N8163, N8149, N6304);
nand NAND4 (N8164, N8129, N4106, N6183, N7825);
buf BUF1 (N8165, N8159);
xor XOR2 (N8166, N8158, N7675);
or OR2 (N8167, N8144, N6870);
and AND4 (N8168, N8166, N4261, N1763, N5253);
or OR2 (N8169, N8165, N5425);
nand NAND2 (N8170, N8148, N2452);
buf BUF1 (N8171, N8139);
nor NOR3 (N8172, N8171, N6651, N1511);
nand NAND3 (N8173, N8143, N3938, N6890);
buf BUF1 (N8174, N8169);
nand NAND3 (N8175, N8172, N6492, N201);
or OR2 (N8176, N8161, N1699);
not NOT1 (N8177, N8163);
buf BUF1 (N8178, N8177);
or OR4 (N8179, N8173, N2065, N4336, N6341);
buf BUF1 (N8180, N8168);
and AND4 (N8181, N8176, N4438, N4099, N4719);
xor XOR2 (N8182, N8181, N468);
nand NAND2 (N8183, N8182, N3681);
nand NAND2 (N8184, N8183, N7038);
buf BUF1 (N8185, N8178);
buf BUF1 (N8186, N8167);
nand NAND4 (N8187, N8184, N5213, N3581, N5903);
nor NOR2 (N8188, N8175, N6216);
not NOT1 (N8189, N8164);
nand NAND3 (N8190, N8174, N5527, N4670);
not NOT1 (N8191, N8170);
and AND4 (N8192, N8180, N501, N6165, N1793);
nor NOR4 (N8193, N8179, N6736, N496, N615);
nor NOR4 (N8194, N8186, N3413, N7298, N5113);
or OR4 (N8195, N8185, N4583, N3343, N5351);
not NOT1 (N8196, N8190);
and AND4 (N8197, N8196, N2940, N974, N4572);
and AND3 (N8198, N8192, N7985, N3205);
nor NOR4 (N8199, N8191, N5684, N4942, N417);
xor XOR2 (N8200, N8162, N4462);
buf BUF1 (N8201, N8198);
or OR4 (N8202, N8187, N6333, N4506, N7084);
buf BUF1 (N8203, N8200);
nor NOR2 (N8204, N8193, N855);
not NOT1 (N8205, N8203);
or OR3 (N8206, N8204, N4511, N1239);
nor NOR3 (N8207, N8199, N2315, N6732);
or OR3 (N8208, N8188, N259, N3103);
buf BUF1 (N8209, N8197);
buf BUF1 (N8210, N8207);
nand NAND3 (N8211, N8206, N2983, N4215);
xor XOR2 (N8212, N8210, N5120);
nor NOR2 (N8213, N8194, N1618);
buf BUF1 (N8214, N8205);
nor NOR4 (N8215, N8212, N2158, N8021, N7774);
not NOT1 (N8216, N8202);
or OR4 (N8217, N8215, N6568, N3191, N2451);
nand NAND4 (N8218, N8217, N5412, N5423, N7211);
nor NOR4 (N8219, N8209, N3487, N716, N1404);
and AND3 (N8220, N8208, N7673, N4822);
not NOT1 (N8221, N8189);
or OR2 (N8222, N8221, N5403);
and AND4 (N8223, N8195, N5448, N5212, N5183);
and AND2 (N8224, N8201, N3601);
and AND3 (N8225, N8220, N1667, N7198);
or OR4 (N8226, N8211, N3520, N4636, N6482);
xor XOR2 (N8227, N8224, N425);
xor XOR2 (N8228, N8222, N4408);
xor XOR2 (N8229, N8216, N1680);
buf BUF1 (N8230, N8213);
or OR4 (N8231, N8229, N3512, N1626, N5711);
or OR2 (N8232, N8231, N1137);
or OR2 (N8233, N8225, N5507);
nand NAND4 (N8234, N8226, N7284, N603, N2913);
not NOT1 (N8235, N8214);
nand NAND2 (N8236, N8233, N877);
not NOT1 (N8237, N8223);
nand NAND2 (N8238, N8219, N2211);
xor XOR2 (N8239, N8235, N3732);
not NOT1 (N8240, N8227);
xor XOR2 (N8241, N8237, N5815);
nand NAND4 (N8242, N8228, N341, N2271, N4635);
or OR3 (N8243, N8239, N3523, N1785);
xor XOR2 (N8244, N8230, N4800);
not NOT1 (N8245, N8241);
and AND4 (N8246, N8240, N4010, N4576, N1815);
xor XOR2 (N8247, N8243, N125);
buf BUF1 (N8248, N8245);
buf BUF1 (N8249, N8248);
and AND3 (N8250, N8232, N6327, N946);
buf BUF1 (N8251, N8244);
nor NOR2 (N8252, N8246, N3814);
buf BUF1 (N8253, N8252);
buf BUF1 (N8254, N8247);
buf BUF1 (N8255, N8251);
nor NOR3 (N8256, N8254, N5673, N3576);
nor NOR4 (N8257, N8238, N4701, N6909, N6073);
nand NAND3 (N8258, N8257, N4432, N218);
not NOT1 (N8259, N8258);
and AND3 (N8260, N8250, N6378, N1765);
or OR2 (N8261, N8259, N1117);
nor NOR4 (N8262, N8261, N3630, N4587, N405);
xor XOR2 (N8263, N8253, N4753);
and AND3 (N8264, N8236, N250, N6187);
or OR2 (N8265, N8255, N3622);
buf BUF1 (N8266, N8263);
xor XOR2 (N8267, N8242, N7601);
xor XOR2 (N8268, N8249, N4991);
nor NOR3 (N8269, N8262, N1938, N1541);
xor XOR2 (N8270, N8269, N5157);
not NOT1 (N8271, N8266);
nand NAND4 (N8272, N8234, N5656, N4681, N6700);
nor NOR2 (N8273, N8271, N2097);
nor NOR3 (N8274, N8260, N7242, N933);
buf BUF1 (N8275, N8272);
nand NAND3 (N8276, N8267, N691, N7568);
not NOT1 (N8277, N8264);
not NOT1 (N8278, N8270);
xor XOR2 (N8279, N8275, N399);
nand NAND4 (N8280, N8278, N1198, N6161, N4820);
nand NAND4 (N8281, N8256, N7789, N1145, N3244);
not NOT1 (N8282, N8280);
and AND3 (N8283, N8265, N5152, N2357);
or OR2 (N8284, N8268, N1408);
nand NAND2 (N8285, N8282, N4330);
or OR3 (N8286, N8281, N138, N6457);
and AND3 (N8287, N8279, N5043, N8283);
xor XOR2 (N8288, N5867, N3348);
nor NOR4 (N8289, N8218, N152, N6530, N4508);
not NOT1 (N8290, N8284);
and AND4 (N8291, N8286, N506, N3867, N5609);
or OR3 (N8292, N8291, N8193, N4605);
not NOT1 (N8293, N8290);
buf BUF1 (N8294, N8276);
or OR3 (N8295, N8289, N2975, N3301);
or OR3 (N8296, N8293, N5015, N6635);
xor XOR2 (N8297, N8296, N3535);
or OR3 (N8298, N8297, N8247, N6679);
and AND2 (N8299, N8298, N6791);
nor NOR3 (N8300, N8273, N1991, N1901);
xor XOR2 (N8301, N8285, N1189);
and AND4 (N8302, N8277, N7417, N7449, N92);
and AND3 (N8303, N8292, N4540, N4448);
and AND4 (N8304, N8295, N2169, N3138, N3526);
and AND4 (N8305, N8304, N6028, N5097, N7096);
nand NAND2 (N8306, N8288, N5564);
and AND2 (N8307, N8274, N6698);
not NOT1 (N8308, N8287);
buf BUF1 (N8309, N8294);
xor XOR2 (N8310, N8299, N5320);
nand NAND2 (N8311, N8300, N7258);
and AND2 (N8312, N8307, N5684);
nor NOR4 (N8313, N8311, N6691, N7258, N1829);
and AND2 (N8314, N8312, N8005);
nor NOR3 (N8315, N8314, N3267, N5407);
nor NOR3 (N8316, N8313, N481, N2888);
nor NOR4 (N8317, N8309, N1645, N1908, N707);
buf BUF1 (N8318, N8316);
nor NOR3 (N8319, N8301, N260, N6905);
or OR2 (N8320, N8315, N8029);
xor XOR2 (N8321, N8306, N707);
and AND4 (N8322, N8303, N7187, N2594, N4418);
buf BUF1 (N8323, N8321);
nand NAND4 (N8324, N8320, N4128, N77, N919);
buf BUF1 (N8325, N8318);
xor XOR2 (N8326, N8302, N8128);
and AND2 (N8327, N8325, N3789);
xor XOR2 (N8328, N8326, N6192);
buf BUF1 (N8329, N8327);
or OR2 (N8330, N8328, N1001);
or OR2 (N8331, N8329, N2769);
buf BUF1 (N8332, N8319);
buf BUF1 (N8333, N8322);
buf BUF1 (N8334, N8333);
xor XOR2 (N8335, N8323, N6774);
or OR3 (N8336, N8330, N2222, N6118);
not NOT1 (N8337, N8336);
or OR3 (N8338, N8334, N691, N7467);
or OR4 (N8339, N8305, N7103, N3725, N507);
nor NOR4 (N8340, N8337, N6106, N8260, N3532);
not NOT1 (N8341, N8331);
not NOT1 (N8342, N8338);
xor XOR2 (N8343, N8324, N6569);
xor XOR2 (N8344, N8341, N309);
and AND4 (N8345, N8332, N3198, N2083, N2410);
buf BUF1 (N8346, N8343);
nand NAND2 (N8347, N8308, N5429);
or OR4 (N8348, N8340, N4603, N2869, N3391);
nor NOR2 (N8349, N8339, N6650);
xor XOR2 (N8350, N8348, N6320);
nor NOR4 (N8351, N8342, N5526, N7356, N6573);
buf BUF1 (N8352, N8347);
nand NAND3 (N8353, N8344, N2532, N7736);
nand NAND4 (N8354, N8346, N7874, N2146, N3292);
and AND3 (N8355, N8353, N5500, N1315);
nand NAND2 (N8356, N8310, N4931);
buf BUF1 (N8357, N8355);
nand NAND4 (N8358, N8350, N411, N2654, N550);
buf BUF1 (N8359, N8351);
xor XOR2 (N8360, N8357, N2170);
not NOT1 (N8361, N8360);
not NOT1 (N8362, N8358);
nor NOR3 (N8363, N8359, N664, N2214);
not NOT1 (N8364, N8335);
or OR2 (N8365, N8352, N5002);
not NOT1 (N8366, N8356);
buf BUF1 (N8367, N8354);
and AND2 (N8368, N8367, N1988);
xor XOR2 (N8369, N8366, N4577);
or OR4 (N8370, N8368, N6732, N6051, N2029);
nor NOR4 (N8371, N8370, N1834, N5412, N399);
xor XOR2 (N8372, N8349, N8148);
nor NOR2 (N8373, N8371, N3928);
and AND3 (N8374, N8317, N1314, N1106);
nand NAND3 (N8375, N8345, N3872, N7266);
not NOT1 (N8376, N8361);
buf BUF1 (N8377, N8376);
or OR3 (N8378, N8363, N2353, N3476);
nand NAND4 (N8379, N8375, N2505, N557, N4466);
and AND3 (N8380, N8372, N300, N6941);
buf BUF1 (N8381, N8365);
not NOT1 (N8382, N8373);
nor NOR2 (N8383, N8378, N3042);
not NOT1 (N8384, N8380);
nand NAND4 (N8385, N8364, N586, N1198, N4658);
buf BUF1 (N8386, N8382);
not NOT1 (N8387, N8362);
or OR3 (N8388, N8386, N3258, N5516);
xor XOR2 (N8389, N8374, N7837);
xor XOR2 (N8390, N8383, N3587);
nor NOR3 (N8391, N8389, N5131, N4972);
buf BUF1 (N8392, N8377);
nor NOR3 (N8393, N8392, N1870, N8363);
not NOT1 (N8394, N8391);
nand NAND4 (N8395, N8381, N1717, N3591, N8393);
or OR4 (N8396, N1862, N6920, N6888, N3297);
nand NAND4 (N8397, N8385, N5905, N2500, N5115);
or OR4 (N8398, N8390, N325, N1639, N8102);
xor XOR2 (N8399, N8398, N4367);
xor XOR2 (N8400, N8394, N2141);
or OR4 (N8401, N8388, N6762, N8144, N6375);
not NOT1 (N8402, N8397);
not NOT1 (N8403, N8379);
xor XOR2 (N8404, N8401, N4746);
or OR3 (N8405, N8400, N4780, N5416);
nor NOR3 (N8406, N8405, N824, N8276);
not NOT1 (N8407, N8384);
and AND3 (N8408, N8399, N6097, N2122);
nand NAND2 (N8409, N8404, N3448);
not NOT1 (N8410, N8396);
buf BUF1 (N8411, N8403);
xor XOR2 (N8412, N8408, N3587);
nand NAND2 (N8413, N8402, N5062);
and AND4 (N8414, N8410, N8007, N2229, N1603);
nand NAND2 (N8415, N8413, N1594);
nor NOR2 (N8416, N8412, N7662);
xor XOR2 (N8417, N8411, N125);
not NOT1 (N8418, N8409);
not NOT1 (N8419, N8395);
and AND2 (N8420, N8417, N7299);
nor NOR4 (N8421, N8369, N8010, N2213, N63);
and AND4 (N8422, N8415, N475, N2365, N4255);
and AND4 (N8423, N8407, N5626, N6913, N3246);
and AND2 (N8424, N8418, N8250);
or OR4 (N8425, N8422, N7094, N4259, N6111);
or OR3 (N8426, N8420, N4106, N5498);
xor XOR2 (N8427, N8416, N7791);
or OR2 (N8428, N8421, N4489);
nor NOR3 (N8429, N8425, N7634, N7243);
and AND4 (N8430, N8423, N4250, N6240, N1004);
not NOT1 (N8431, N8428);
not NOT1 (N8432, N8419);
nor NOR3 (N8433, N8424, N5208, N4574);
nor NOR2 (N8434, N8414, N4910);
and AND4 (N8435, N8433, N3832, N1997, N6436);
xor XOR2 (N8436, N8387, N4088);
xor XOR2 (N8437, N8431, N6062);
nor NOR4 (N8438, N8426, N1392, N7026, N2179);
nor NOR2 (N8439, N8436, N6167);
nor NOR3 (N8440, N8406, N4248, N8336);
or OR3 (N8441, N8430, N7517, N2542);
xor XOR2 (N8442, N8437, N689);
buf BUF1 (N8443, N8442);
not NOT1 (N8444, N8435);
not NOT1 (N8445, N8429);
nand NAND4 (N8446, N8445, N6001, N2323, N8379);
xor XOR2 (N8447, N8434, N5817);
xor XOR2 (N8448, N8446, N4014);
buf BUF1 (N8449, N8447);
or OR2 (N8450, N8438, N4827);
and AND4 (N8451, N8439, N5924, N7579, N3771);
not NOT1 (N8452, N8441);
nor NOR4 (N8453, N8444, N5691, N1887, N7837);
or OR2 (N8454, N8452, N7443);
and AND4 (N8455, N8432, N4844, N5543, N3268);
nand NAND4 (N8456, N8455, N2295, N5839, N2611);
and AND2 (N8457, N8451, N1908);
not NOT1 (N8458, N8443);
nor NOR3 (N8459, N8449, N247, N5049);
or OR4 (N8460, N8456, N3065, N280, N1561);
or OR3 (N8461, N8459, N7999, N8019);
or OR2 (N8462, N8427, N967);
or OR4 (N8463, N8440, N8005, N3936, N177);
nor NOR4 (N8464, N8450, N3519, N6318, N4425);
buf BUF1 (N8465, N8457);
xor XOR2 (N8466, N8462, N3322);
xor XOR2 (N8467, N8448, N6550);
xor XOR2 (N8468, N8461, N4378);
not NOT1 (N8469, N8454);
nor NOR4 (N8470, N8467, N5871, N5716, N1590);
not NOT1 (N8471, N8466);
not NOT1 (N8472, N8469);
xor XOR2 (N8473, N8470, N5552);
nand NAND2 (N8474, N8458, N6712);
buf BUF1 (N8475, N8453);
or OR2 (N8476, N8464, N3525);
or OR2 (N8477, N8476, N2478);
not NOT1 (N8478, N8472);
or OR3 (N8479, N8475, N6651, N1929);
and AND3 (N8480, N8463, N5567, N1308);
nand NAND3 (N8481, N8465, N5933, N6475);
nand NAND3 (N8482, N8473, N7279, N1944);
not NOT1 (N8483, N8477);
xor XOR2 (N8484, N8481, N4732);
not NOT1 (N8485, N8483);
buf BUF1 (N8486, N8471);
nand NAND2 (N8487, N8468, N6218);
xor XOR2 (N8488, N8480, N4899);
and AND4 (N8489, N8478, N2057, N6154, N1320);
buf BUF1 (N8490, N8484);
nor NOR2 (N8491, N8487, N270);
nor NOR3 (N8492, N8490, N6610, N622);
nand NAND3 (N8493, N8486, N3446, N1962);
nand NAND3 (N8494, N8482, N2408, N3757);
not NOT1 (N8495, N8460);
not NOT1 (N8496, N8494);
or OR3 (N8497, N8491, N1876, N7041);
xor XOR2 (N8498, N8474, N7693);
buf BUF1 (N8499, N8493);
xor XOR2 (N8500, N8496, N6619);
nor NOR2 (N8501, N8497, N5448);
nor NOR4 (N8502, N8495, N1648, N2952, N2267);
and AND4 (N8503, N8501, N1744, N7123, N2948);
nor NOR3 (N8504, N8479, N2237, N4700);
or OR4 (N8505, N8503, N3425, N4848, N8429);
buf BUF1 (N8506, N8489);
nand NAND4 (N8507, N8505, N8505, N7891, N6042);
or OR3 (N8508, N8498, N4858, N3114);
and AND2 (N8509, N8492, N7845);
and AND2 (N8510, N8485, N4740);
and AND3 (N8511, N8499, N6565, N239);
buf BUF1 (N8512, N8508);
xor XOR2 (N8513, N8512, N4700);
not NOT1 (N8514, N8502);
nand NAND4 (N8515, N8511, N2905, N1853, N6445);
xor XOR2 (N8516, N8488, N2400);
and AND3 (N8517, N8504, N5162, N3775);
nor NOR3 (N8518, N8516, N7229, N4023);
xor XOR2 (N8519, N8507, N2435);
nor NOR2 (N8520, N8500, N1218);
nand NAND3 (N8521, N8514, N1099, N2322);
xor XOR2 (N8522, N8521, N8368);
nor NOR2 (N8523, N8506, N3833);
xor XOR2 (N8524, N8510, N75);
buf BUF1 (N8525, N8519);
and AND4 (N8526, N8517, N2453, N8062, N1436);
and AND3 (N8527, N8509, N4026, N2966);
nor NOR2 (N8528, N8518, N2524);
nand NAND2 (N8529, N8515, N177);
xor XOR2 (N8530, N8513, N2061);
buf BUF1 (N8531, N8523);
nand NAND4 (N8532, N8526, N4433, N2568, N3093);
nor NOR2 (N8533, N8529, N1650);
buf BUF1 (N8534, N8531);
or OR2 (N8535, N8525, N5349);
nand NAND3 (N8536, N8535, N6243, N2512);
not NOT1 (N8537, N8524);
xor XOR2 (N8538, N8533, N4839);
or OR4 (N8539, N8537, N7272, N1837, N80);
not NOT1 (N8540, N8539);
and AND4 (N8541, N8528, N5973, N387, N8445);
nand NAND3 (N8542, N8532, N7750, N3278);
or OR3 (N8543, N8520, N336, N7084);
not NOT1 (N8544, N8541);
and AND3 (N8545, N8544, N7486, N7418);
nand NAND3 (N8546, N8527, N1177, N4799);
and AND3 (N8547, N8536, N4395, N2069);
not NOT1 (N8548, N8543);
buf BUF1 (N8549, N8542);
not NOT1 (N8550, N8530);
buf BUF1 (N8551, N8545);
nand NAND4 (N8552, N8548, N6715, N3869, N6742);
xor XOR2 (N8553, N8550, N5498);
buf BUF1 (N8554, N8522);
buf BUF1 (N8555, N8553);
or OR4 (N8556, N8546, N6997, N2951, N2191);
and AND3 (N8557, N8555, N4606, N8023);
nor NOR4 (N8558, N8540, N4792, N4020, N3948);
xor XOR2 (N8559, N8549, N1988);
not NOT1 (N8560, N8551);
and AND3 (N8561, N8554, N3021, N3546);
xor XOR2 (N8562, N8552, N7559);
not NOT1 (N8563, N8538);
xor XOR2 (N8564, N8559, N3406);
and AND2 (N8565, N8561, N8063);
or OR3 (N8566, N8557, N2474, N386);
or OR4 (N8567, N8565, N5969, N6837, N1479);
and AND3 (N8568, N8563, N3401, N4705);
or OR4 (N8569, N8564, N3946, N6455, N6853);
and AND4 (N8570, N8560, N322, N4601, N8128);
nor NOR2 (N8571, N8547, N4367);
xor XOR2 (N8572, N8569, N5650);
nand NAND3 (N8573, N8572, N2410, N1010);
buf BUF1 (N8574, N8567);
xor XOR2 (N8575, N8562, N3006);
nand NAND3 (N8576, N8573, N3066, N7151);
not NOT1 (N8577, N8556);
not NOT1 (N8578, N8574);
not NOT1 (N8579, N8534);
xor XOR2 (N8580, N8579, N6830);
nand NAND3 (N8581, N8577, N213, N1454);
not NOT1 (N8582, N8578);
xor XOR2 (N8583, N8571, N455);
buf BUF1 (N8584, N8575);
buf BUF1 (N8585, N8558);
xor XOR2 (N8586, N8566, N5708);
nand NAND3 (N8587, N8580, N3134, N4977);
or OR3 (N8588, N8576, N5447, N3309);
and AND3 (N8589, N8583, N6887, N2229);
nor NOR3 (N8590, N8581, N336, N7750);
buf BUF1 (N8591, N8589);
nand NAND2 (N8592, N8568, N4113);
nand NAND2 (N8593, N8585, N2545);
not NOT1 (N8594, N8570);
xor XOR2 (N8595, N8586, N4472);
and AND3 (N8596, N8594, N551, N7208);
not NOT1 (N8597, N8595);
not NOT1 (N8598, N8587);
buf BUF1 (N8599, N8591);
xor XOR2 (N8600, N8599, N3725);
nand NAND2 (N8601, N8588, N2912);
or OR2 (N8602, N8598, N259);
and AND2 (N8603, N8593, N3396);
not NOT1 (N8604, N8590);
nand NAND4 (N8605, N8604, N4347, N6354, N7593);
or OR3 (N8606, N8605, N971, N5797);
xor XOR2 (N8607, N8602, N2732);
buf BUF1 (N8608, N8607);
and AND3 (N8609, N8606, N6131, N741);
nand NAND3 (N8610, N8600, N2817, N2476);
xor XOR2 (N8611, N8597, N715);
and AND3 (N8612, N8596, N7284, N8211);
and AND4 (N8613, N8582, N6394, N574, N4366);
or OR4 (N8614, N8609, N3412, N7670, N2716);
buf BUF1 (N8615, N8610);
and AND3 (N8616, N8601, N5600, N8113);
xor XOR2 (N8617, N8613, N4510);
and AND4 (N8618, N8612, N3785, N2915, N3960);
or OR3 (N8619, N8592, N841, N3823);
buf BUF1 (N8620, N8584);
or OR2 (N8621, N8620, N57);
or OR4 (N8622, N8616, N3003, N3744, N7734);
nand NAND4 (N8623, N8611, N7055, N4087, N1219);
or OR4 (N8624, N8608, N3585, N1227, N1045);
nor NOR3 (N8625, N8622, N4917, N4808);
nand NAND4 (N8626, N8623, N47, N7105, N8404);
nand NAND4 (N8627, N8615, N5100, N4011, N8477);
nand NAND4 (N8628, N8619, N6767, N2396, N2212);
not NOT1 (N8629, N8625);
buf BUF1 (N8630, N8621);
or OR3 (N8631, N8617, N1017, N2202);
nand NAND3 (N8632, N8624, N519, N171);
nand NAND2 (N8633, N8603, N807);
buf BUF1 (N8634, N8632);
or OR4 (N8635, N8614, N6863, N1151, N664);
and AND4 (N8636, N8626, N7722, N1072, N5332);
nor NOR2 (N8637, N8635, N683);
or OR4 (N8638, N8633, N7141, N3216, N8346);
not NOT1 (N8639, N8637);
not NOT1 (N8640, N8638);
nor NOR3 (N8641, N8627, N3169, N5160);
not NOT1 (N8642, N8631);
xor XOR2 (N8643, N8628, N5322);
xor XOR2 (N8644, N8642, N6196);
not NOT1 (N8645, N8641);
not NOT1 (N8646, N8643);
not NOT1 (N8647, N8644);
nor NOR4 (N8648, N8636, N3650, N7745, N6849);
not NOT1 (N8649, N8634);
or OR4 (N8650, N8629, N6440, N3454, N3181);
and AND4 (N8651, N8649, N4404, N4006, N7822);
buf BUF1 (N8652, N8646);
xor XOR2 (N8653, N8650, N7458);
not NOT1 (N8654, N8652);
nor NOR2 (N8655, N8630, N7591);
not NOT1 (N8656, N8645);
and AND2 (N8657, N8639, N8459);
not NOT1 (N8658, N8647);
or OR2 (N8659, N8656, N6879);
buf BUF1 (N8660, N8657);
buf BUF1 (N8661, N8653);
or OR2 (N8662, N8655, N6389);
nor NOR4 (N8663, N8654, N8067, N6267, N5296);
nor NOR2 (N8664, N8661, N5118);
or OR4 (N8665, N8640, N5258, N7825, N5702);
xor XOR2 (N8666, N8648, N3863);
not NOT1 (N8667, N8665);
or OR3 (N8668, N8663, N3362, N1359);
xor XOR2 (N8669, N8660, N5949);
buf BUF1 (N8670, N8666);
nor NOR2 (N8671, N8664, N2249);
xor XOR2 (N8672, N8659, N5755);
xor XOR2 (N8673, N8651, N8152);
nand NAND2 (N8674, N8658, N1521);
xor XOR2 (N8675, N8674, N2364);
buf BUF1 (N8676, N8669);
not NOT1 (N8677, N8670);
not NOT1 (N8678, N8662);
buf BUF1 (N8679, N8618);
nand NAND3 (N8680, N8668, N7619, N7558);
nor NOR2 (N8681, N8675, N6160);
nor NOR4 (N8682, N8672, N7576, N8418, N7240);
nand NAND3 (N8683, N8682, N8079, N2002);
buf BUF1 (N8684, N8667);
nor NOR4 (N8685, N8680, N5694, N6613, N4769);
not NOT1 (N8686, N8679);
nand NAND4 (N8687, N8671, N6831, N7420, N5959);
buf BUF1 (N8688, N8685);
nand NAND2 (N8689, N8673, N1540);
buf BUF1 (N8690, N8677);
xor XOR2 (N8691, N8686, N3085);
not NOT1 (N8692, N8678);
xor XOR2 (N8693, N8690, N7130);
xor XOR2 (N8694, N8692, N4140);
or OR3 (N8695, N8684, N7352, N8476);
buf BUF1 (N8696, N8676);
and AND4 (N8697, N8683, N7535, N2407, N728);
and AND3 (N8698, N8694, N2665, N8587);
or OR3 (N8699, N8691, N4442, N1945);
xor XOR2 (N8700, N8698, N7066);
nand NAND2 (N8701, N8700, N920);
nand NAND2 (N8702, N8688, N4530);
not NOT1 (N8703, N8695);
buf BUF1 (N8704, N8693);
nor NOR3 (N8705, N8681, N7546, N1867);
not NOT1 (N8706, N8687);
xor XOR2 (N8707, N8697, N2293);
nor NOR2 (N8708, N8706, N2034);
nand NAND2 (N8709, N8707, N136);
or OR3 (N8710, N8704, N7265, N3759);
or OR2 (N8711, N8689, N6950);
buf BUF1 (N8712, N8709);
buf BUF1 (N8713, N8703);
xor XOR2 (N8714, N8702, N8187);
and AND4 (N8715, N8712, N1837, N1658, N2397);
nand NAND2 (N8716, N8710, N6128);
buf BUF1 (N8717, N8696);
buf BUF1 (N8718, N8699);
nand NAND2 (N8719, N8701, N3338);
not NOT1 (N8720, N8713);
and AND4 (N8721, N8719, N2044, N6288, N645);
and AND2 (N8722, N8708, N6159);
or OR3 (N8723, N8716, N7381, N5385);
xor XOR2 (N8724, N8705, N3706);
nand NAND4 (N8725, N8722, N6790, N6843, N2080);
not NOT1 (N8726, N8724);
not NOT1 (N8727, N8718);
buf BUF1 (N8728, N8727);
nor NOR3 (N8729, N8711, N401, N7165);
not NOT1 (N8730, N8714);
xor XOR2 (N8731, N8721, N435);
nor NOR3 (N8732, N8731, N319, N7855);
xor XOR2 (N8733, N8732, N2384);
and AND4 (N8734, N8733, N1124, N5696, N689);
xor XOR2 (N8735, N8728, N1193);
and AND2 (N8736, N8726, N1805);
and AND3 (N8737, N8723, N901, N224);
or OR3 (N8738, N8734, N7820, N2934);
xor XOR2 (N8739, N8736, N1945);
and AND2 (N8740, N8715, N778);
nor NOR2 (N8741, N8725, N1221);
not NOT1 (N8742, N8739);
or OR2 (N8743, N8735, N4237);
or OR4 (N8744, N8741, N6667, N6330, N2345);
not NOT1 (N8745, N8729);
xor XOR2 (N8746, N8740, N5028);
nor NOR4 (N8747, N8743, N2260, N8019, N310);
not NOT1 (N8748, N8738);
not NOT1 (N8749, N8744);
buf BUF1 (N8750, N8730);
buf BUF1 (N8751, N8720);
and AND2 (N8752, N8751, N1543);
nor NOR2 (N8753, N8742, N2850);
or OR4 (N8754, N8749, N7928, N2916, N447);
nand NAND4 (N8755, N8752, N886, N6886, N517);
buf BUF1 (N8756, N8717);
nor NOR3 (N8757, N8753, N2872, N2765);
and AND3 (N8758, N8754, N8367, N99);
nand NAND3 (N8759, N8746, N7199, N2705);
or OR4 (N8760, N8745, N6098, N6322, N767);
or OR4 (N8761, N8756, N1995, N3158, N6636);
nor NOR4 (N8762, N8760, N3213, N8696, N5433);
not NOT1 (N8763, N8759);
or OR4 (N8764, N8761, N5181, N6188, N2650);
or OR4 (N8765, N8747, N1615, N1936, N6253);
or OR3 (N8766, N8757, N1043, N3343);
xor XOR2 (N8767, N8750, N788);
buf BUF1 (N8768, N8737);
not NOT1 (N8769, N8765);
buf BUF1 (N8770, N8766);
not NOT1 (N8771, N8768);
and AND4 (N8772, N8755, N5541, N3325, N5663);
nor NOR2 (N8773, N8758, N6815);
or OR3 (N8774, N8769, N8398, N4922);
buf BUF1 (N8775, N8771);
nand NAND2 (N8776, N8773, N3842);
buf BUF1 (N8777, N8762);
and AND2 (N8778, N8767, N5912);
and AND3 (N8779, N8777, N1105, N4585);
xor XOR2 (N8780, N8774, N620);
and AND2 (N8781, N8778, N1467);
or OR4 (N8782, N8763, N6245, N6526, N322);
xor XOR2 (N8783, N8770, N7546);
or OR3 (N8784, N8779, N5962, N7640);
or OR2 (N8785, N8764, N2504);
and AND4 (N8786, N8782, N1919, N879, N8470);
not NOT1 (N8787, N8776);
xor XOR2 (N8788, N8787, N3727);
nand NAND3 (N8789, N8788, N5229, N5921);
and AND4 (N8790, N8772, N6411, N5160, N3300);
buf BUF1 (N8791, N8789);
buf BUF1 (N8792, N8748);
not NOT1 (N8793, N8781);
xor XOR2 (N8794, N8780, N8700);
nand NAND4 (N8795, N8784, N1735, N495, N6786);
not NOT1 (N8796, N8775);
nand NAND4 (N8797, N8790, N1454, N8576, N4263);
and AND3 (N8798, N8786, N2055, N172);
nor NOR2 (N8799, N8795, N5248);
buf BUF1 (N8800, N8796);
and AND2 (N8801, N8783, N402);
or OR4 (N8802, N8785, N8746, N6486, N8515);
nand NAND2 (N8803, N8797, N5935);
nand NAND3 (N8804, N8792, N1146, N3942);
or OR3 (N8805, N8801, N3971, N7054);
xor XOR2 (N8806, N8798, N5994);
and AND4 (N8807, N8791, N23, N6121, N3726);
and AND2 (N8808, N8802, N753);
or OR2 (N8809, N8800, N3125);
nand NAND4 (N8810, N8794, N2918, N7960, N382);
or OR2 (N8811, N8807, N441);
and AND2 (N8812, N8808, N8681);
nor NOR4 (N8813, N8793, N2071, N2851, N2601);
or OR2 (N8814, N8806, N7566);
not NOT1 (N8815, N8810);
xor XOR2 (N8816, N8812, N5582);
buf BUF1 (N8817, N8809);
not NOT1 (N8818, N8804);
xor XOR2 (N8819, N8799, N3641);
nand NAND2 (N8820, N8803, N417);
or OR2 (N8821, N8814, N7276);
xor XOR2 (N8822, N8821, N7067);
nand NAND4 (N8823, N8805, N3424, N7783, N821);
not NOT1 (N8824, N8815);
xor XOR2 (N8825, N8824, N6661);
not NOT1 (N8826, N8813);
nor NOR3 (N8827, N8820, N2282, N4862);
nor NOR2 (N8828, N8825, N2165);
not NOT1 (N8829, N8818);
nor NOR4 (N8830, N8819, N3879, N3608, N6763);
nor NOR3 (N8831, N8823, N1473, N743);
buf BUF1 (N8832, N8829);
or OR2 (N8833, N8817, N8201);
and AND4 (N8834, N8822, N2592, N6479, N3179);
xor XOR2 (N8835, N8827, N2051);
or OR3 (N8836, N8816, N8409, N86);
nand NAND4 (N8837, N8830, N2337, N2349, N1241);
not NOT1 (N8838, N8828);
not NOT1 (N8839, N8831);
not NOT1 (N8840, N8834);
or OR4 (N8841, N8836, N4925, N6733, N810);
not NOT1 (N8842, N8838);
not NOT1 (N8843, N8837);
or OR4 (N8844, N8826, N1450, N344, N1312);
or OR3 (N8845, N8832, N8389, N542);
nor NOR4 (N8846, N8840, N4555, N1646, N6620);
nand NAND3 (N8847, N8839, N6882, N8628);
nor NOR2 (N8848, N8846, N726);
xor XOR2 (N8849, N8845, N1564);
xor XOR2 (N8850, N8844, N2932);
or OR4 (N8851, N8847, N3887, N5528, N7890);
xor XOR2 (N8852, N8835, N6310);
nand NAND2 (N8853, N8843, N7407);
buf BUF1 (N8854, N8848);
buf BUF1 (N8855, N8833);
not NOT1 (N8856, N8811);
not NOT1 (N8857, N8842);
or OR2 (N8858, N8857, N5805);
nand NAND4 (N8859, N8855, N5260, N7730, N5595);
or OR4 (N8860, N8854, N1256, N6066, N1068);
xor XOR2 (N8861, N8856, N7000);
and AND4 (N8862, N8851, N5058, N7944, N519);
buf BUF1 (N8863, N8849);
and AND4 (N8864, N8858, N3971, N645, N2963);
nand NAND3 (N8865, N8862, N8644, N6960);
buf BUF1 (N8866, N8850);
xor XOR2 (N8867, N8841, N4082);
not NOT1 (N8868, N8866);
and AND2 (N8869, N8852, N1520);
and AND2 (N8870, N8860, N3467);
not NOT1 (N8871, N8869);
and AND4 (N8872, N8870, N8231, N2637, N5172);
nand NAND4 (N8873, N8859, N5038, N4079, N5184);
or OR2 (N8874, N8853, N2197);
not NOT1 (N8875, N8868);
and AND4 (N8876, N8867, N3903, N4474, N6037);
nor NOR4 (N8877, N8874, N262, N3898, N4782);
or OR2 (N8878, N8873, N2352);
xor XOR2 (N8879, N8877, N3795);
or OR4 (N8880, N8865, N2556, N529, N8817);
or OR2 (N8881, N8863, N7715);
or OR3 (N8882, N8876, N887, N2017);
not NOT1 (N8883, N8881);
xor XOR2 (N8884, N8871, N2156);
nor NOR4 (N8885, N8875, N1794, N2358, N2356);
nand NAND4 (N8886, N8884, N4648, N1912, N5030);
not NOT1 (N8887, N8878);
not NOT1 (N8888, N8882);
nor NOR2 (N8889, N8880, N2403);
nor NOR2 (N8890, N8889, N985);
and AND2 (N8891, N8886, N6715);
and AND4 (N8892, N8891, N5664, N8876, N3346);
or OR4 (N8893, N8864, N6849, N2066, N5842);
nor NOR3 (N8894, N8893, N1427, N3332);
nand NAND4 (N8895, N8887, N147, N448, N3666);
xor XOR2 (N8896, N8892, N3702);
buf BUF1 (N8897, N8895);
not NOT1 (N8898, N8897);
xor XOR2 (N8899, N8872, N292);
or OR4 (N8900, N8883, N7152, N2424, N7421);
nor NOR2 (N8901, N8894, N5645);
or OR3 (N8902, N8879, N4329, N1596);
or OR2 (N8903, N8901, N4080);
nor NOR4 (N8904, N8896, N4580, N3896, N2948);
nor NOR2 (N8905, N8861, N8315);
and AND3 (N8906, N8900, N24, N2013);
not NOT1 (N8907, N8906);
xor XOR2 (N8908, N8888, N136);
buf BUF1 (N8909, N8902);
nand NAND3 (N8910, N8899, N6121, N8287);
or OR3 (N8911, N8908, N8665, N4362);
not NOT1 (N8912, N8911);
xor XOR2 (N8913, N8912, N1847);
nand NAND4 (N8914, N8909, N2911, N5870, N285);
xor XOR2 (N8915, N8913, N4946);
and AND4 (N8916, N8898, N5973, N1099, N6925);
or OR3 (N8917, N8916, N5143, N435);
nor NOR4 (N8918, N8915, N7795, N4359, N5292);
nand NAND4 (N8919, N8903, N6766, N2360, N8363);
and AND2 (N8920, N8885, N3371);
nor NOR4 (N8921, N8918, N536, N4753, N2378);
xor XOR2 (N8922, N8920, N4578);
buf BUF1 (N8923, N8907);
nor NOR4 (N8924, N8923, N6550, N760, N6975);
nor NOR2 (N8925, N8924, N4636);
xor XOR2 (N8926, N8910, N8657);
nor NOR3 (N8927, N8904, N2927, N3465);
buf BUF1 (N8928, N8925);
or OR3 (N8929, N8921, N4068, N7462);
and AND2 (N8930, N8917, N7632);
or OR4 (N8931, N8926, N6001, N8621, N256);
xor XOR2 (N8932, N8919, N256);
buf BUF1 (N8933, N8930);
buf BUF1 (N8934, N8933);
nor NOR3 (N8935, N8922, N4801, N1437);
nor NOR2 (N8936, N8927, N6031);
or OR3 (N8937, N8928, N7756, N2465);
or OR4 (N8938, N8931, N8585, N7954, N4845);
nor NOR3 (N8939, N8935, N478, N2706);
xor XOR2 (N8940, N8937, N7071);
or OR3 (N8941, N8932, N2251, N2533);
xor XOR2 (N8942, N8905, N5030);
nand NAND4 (N8943, N8938, N6151, N4395, N7581);
buf BUF1 (N8944, N8939);
buf BUF1 (N8945, N8943);
or OR3 (N8946, N8934, N584, N1892);
not NOT1 (N8947, N8914);
or OR2 (N8948, N8940, N5588);
nand NAND2 (N8949, N8936, N347);
nor NOR4 (N8950, N8948, N2129, N858, N7180);
xor XOR2 (N8951, N8929, N2716);
not NOT1 (N8952, N8947);
and AND3 (N8953, N8946, N22, N1312);
or OR3 (N8954, N8944, N2958, N6076);
or OR3 (N8955, N8954, N893, N7640);
nor NOR4 (N8956, N8952, N8352, N7945, N5995);
or OR2 (N8957, N8953, N1014);
or OR2 (N8958, N8951, N6819);
nand NAND3 (N8959, N8890, N1359, N5141);
nor NOR3 (N8960, N8945, N6957, N6407);
buf BUF1 (N8961, N8955);
or OR4 (N8962, N8941, N4391, N3788, N736);
nand NAND3 (N8963, N8957, N5088, N6140);
or OR2 (N8964, N8961, N2668);
not NOT1 (N8965, N8960);
or OR4 (N8966, N8942, N535, N495, N2902);
or OR2 (N8967, N8956, N1679);
buf BUF1 (N8968, N8950);
nand NAND3 (N8969, N8949, N6437, N8755);
xor XOR2 (N8970, N8967, N4551);
nand NAND4 (N8971, N8965, N3209, N4236, N7556);
buf BUF1 (N8972, N8964);
or OR3 (N8973, N8968, N8969, N3034);
and AND2 (N8974, N5251, N3313);
not NOT1 (N8975, N8958);
buf BUF1 (N8976, N8970);
nand NAND4 (N8977, N8971, N2673, N3061, N3617);
nor NOR4 (N8978, N8975, N7664, N6714, N7191);
nand NAND4 (N8979, N8959, N2020, N2553, N7978);
nand NAND3 (N8980, N8973, N7524, N7566);
nor NOR2 (N8981, N8962, N3536);
or OR2 (N8982, N8981, N3558);
nor NOR2 (N8983, N8972, N6631);
or OR3 (N8984, N8982, N895, N7923);
buf BUF1 (N8985, N8984);
nor NOR4 (N8986, N8977, N4310, N8874, N6640);
and AND2 (N8987, N8976, N5201);
and AND2 (N8988, N8986, N8576);
nand NAND4 (N8989, N8983, N6403, N30, N3612);
and AND4 (N8990, N8979, N3122, N7648, N1610);
buf BUF1 (N8991, N8980);
xor XOR2 (N8992, N8985, N123);
buf BUF1 (N8993, N8988);
xor XOR2 (N8994, N8991, N4526);
not NOT1 (N8995, N8966);
xor XOR2 (N8996, N8963, N618);
nand NAND4 (N8997, N8989, N2199, N6431, N7099);
xor XOR2 (N8998, N8996, N3418);
xor XOR2 (N8999, N8992, N5971);
not NOT1 (N9000, N8978);
not NOT1 (N9001, N8998);
nand NAND2 (N9002, N8987, N2534);
or OR4 (N9003, N8974, N4924, N7255, N7979);
not NOT1 (N9004, N9003);
xor XOR2 (N9005, N9001, N5631);
xor XOR2 (N9006, N9000, N3667);
nor NOR2 (N9007, N8999, N2734);
nor NOR4 (N9008, N9005, N2742, N8072, N6276);
or OR4 (N9009, N8994, N64, N157, N5421);
buf BUF1 (N9010, N8990);
or OR2 (N9011, N9002, N5559);
nand NAND2 (N9012, N9007, N2068);
and AND4 (N9013, N8995, N5929, N404, N8061);
nand NAND3 (N9014, N9006, N185, N4663);
not NOT1 (N9015, N8997);
xor XOR2 (N9016, N9015, N6019);
nor NOR2 (N9017, N8993, N362);
xor XOR2 (N9018, N9011, N2017);
or OR3 (N9019, N9012, N6023, N8575);
not NOT1 (N9020, N9009);
or OR4 (N9021, N9014, N2598, N4036, N5353);
buf BUF1 (N9022, N9020);
or OR4 (N9023, N9004, N2071, N6971, N5161);
not NOT1 (N9024, N9021);
nand NAND4 (N9025, N9013, N3686, N825, N5300);
nand NAND3 (N9026, N9017, N6518, N4531);
nand NAND3 (N9027, N9008, N1238, N461);
buf BUF1 (N9028, N9023);
xor XOR2 (N9029, N9026, N1926);
nor NOR2 (N9030, N9027, N1864);
xor XOR2 (N9031, N9018, N5858);
nor NOR3 (N9032, N9025, N4253, N3728);
nand NAND3 (N9033, N9029, N8094, N8825);
nand NAND2 (N9034, N9010, N5963);
not NOT1 (N9035, N9028);
xor XOR2 (N9036, N9035, N1862);
or OR3 (N9037, N9036, N2480, N3699);
not NOT1 (N9038, N9016);
and AND4 (N9039, N9022, N2989, N8239, N8925);
xor XOR2 (N9040, N9030, N1043);
and AND2 (N9041, N9037, N5579);
nand NAND3 (N9042, N9039, N8821, N6288);
xor XOR2 (N9043, N9019, N8432);
buf BUF1 (N9044, N9034);
buf BUF1 (N9045, N9032);
xor XOR2 (N9046, N9024, N6137);
or OR4 (N9047, N9042, N5213, N7715, N4537);
xor XOR2 (N9048, N9045, N1314);
and AND3 (N9049, N9033, N6798, N6211);
xor XOR2 (N9050, N9031, N1756);
xor XOR2 (N9051, N9043, N5187);
nand NAND3 (N9052, N9044, N2923, N7555);
nor NOR3 (N9053, N9051, N6103, N6859);
xor XOR2 (N9054, N9047, N6248);
nor NOR2 (N9055, N9052, N4533);
nand NAND3 (N9056, N9048, N1185, N1008);
nand NAND4 (N9057, N9040, N7390, N2333, N6308);
not NOT1 (N9058, N9054);
buf BUF1 (N9059, N9055);
and AND2 (N9060, N9038, N7621);
not NOT1 (N9061, N9041);
nor NOR3 (N9062, N9059, N8033, N1809);
nor NOR2 (N9063, N9053, N6007);
nor NOR4 (N9064, N9057, N8872, N249, N5390);
nor NOR4 (N9065, N9064, N2260, N8189, N6523);
not NOT1 (N9066, N9061);
and AND3 (N9067, N9056, N3726, N218);
nor NOR4 (N9068, N9050, N4744, N6368, N4381);
xor XOR2 (N9069, N9065, N3027);
nand NAND2 (N9070, N9067, N2460);
or OR2 (N9071, N9063, N86);
nand NAND2 (N9072, N9062, N4724);
and AND3 (N9073, N9049, N4727, N5555);
xor XOR2 (N9074, N9071, N8079);
not NOT1 (N9075, N9058);
buf BUF1 (N9076, N9072);
and AND3 (N9077, N9046, N8337, N4363);
buf BUF1 (N9078, N9066);
nor NOR3 (N9079, N9078, N1101, N1070);
buf BUF1 (N9080, N9073);
nor NOR2 (N9081, N9070, N3829);
or OR4 (N9082, N9076, N3234, N451, N2362);
xor XOR2 (N9083, N9077, N4249);
buf BUF1 (N9084, N9068);
or OR3 (N9085, N9081, N7703, N8547);
nor NOR2 (N9086, N9075, N4864);
nor NOR3 (N9087, N9082, N2671, N2962);
not NOT1 (N9088, N9079);
and AND3 (N9089, N9083, N4189, N2350);
buf BUF1 (N9090, N9084);
nand NAND3 (N9091, N9069, N1756, N8177);
and AND3 (N9092, N9074, N8673, N7291);
xor XOR2 (N9093, N9086, N2053);
xor XOR2 (N9094, N9089, N2129);
nor NOR2 (N9095, N9094, N3777);
xor XOR2 (N9096, N9087, N6328);
and AND4 (N9097, N9088, N4726, N1318, N604);
nor NOR3 (N9098, N9096, N8976, N6894);
nand NAND4 (N9099, N9091, N407, N2656, N2121);
or OR2 (N9100, N9080, N6288);
buf BUF1 (N9101, N9099);
nand NAND3 (N9102, N9101, N9052, N1081);
not NOT1 (N9103, N9098);
nand NAND4 (N9104, N9093, N2980, N5329, N72);
or OR4 (N9105, N9102, N5256, N2221, N8808);
and AND2 (N9106, N9097, N1745);
or OR2 (N9107, N9060, N6375);
nand NAND3 (N9108, N9095, N5449, N2466);
nand NAND3 (N9109, N9107, N8987, N773);
or OR2 (N9110, N9108, N4471);
buf BUF1 (N9111, N9085);
nor NOR4 (N9112, N9103, N6526, N1025, N2890);
not NOT1 (N9113, N9104);
nor NOR4 (N9114, N9090, N5594, N2491, N7311);
nand NAND3 (N9115, N9110, N3086, N6230);
nand NAND4 (N9116, N9109, N8927, N4472, N356);
or OR4 (N9117, N9106, N6539, N8225, N7413);
nor NOR3 (N9118, N9111, N8463, N2705);
and AND4 (N9119, N9112, N4838, N5927, N5258);
xor XOR2 (N9120, N9113, N3970);
or OR4 (N9121, N9117, N7113, N7539, N857);
nor NOR4 (N9122, N9119, N219, N4442, N8129);
or OR3 (N9123, N9105, N6939, N7992);
nor NOR2 (N9124, N9118, N6432);
xor XOR2 (N9125, N9121, N2852);
or OR4 (N9126, N9092, N8602, N4180, N831);
not NOT1 (N9127, N9123);
xor XOR2 (N9128, N9115, N5672);
and AND4 (N9129, N9125, N5296, N4669, N6963);
and AND4 (N9130, N9129, N7935, N4232, N190);
or OR3 (N9131, N9116, N5673, N4865);
nand NAND2 (N9132, N9126, N1897);
not NOT1 (N9133, N9122);
not NOT1 (N9134, N9114);
or OR3 (N9135, N9131, N6019, N7318);
buf BUF1 (N9136, N9135);
nor NOR2 (N9137, N9133, N9073);
xor XOR2 (N9138, N9128, N756);
or OR2 (N9139, N9120, N3893);
buf BUF1 (N9140, N9138);
xor XOR2 (N9141, N9136, N8508);
nand NAND2 (N9142, N9141, N8689);
nand NAND3 (N9143, N9134, N461, N6629);
buf BUF1 (N9144, N9142);
not NOT1 (N9145, N9130);
nor NOR3 (N9146, N9137, N7769, N3001);
xor XOR2 (N9147, N9140, N2016);
xor XOR2 (N9148, N9100, N2615);
buf BUF1 (N9149, N9124);
not NOT1 (N9150, N9148);
xor XOR2 (N9151, N9144, N7197);
buf BUF1 (N9152, N9143);
nand NAND2 (N9153, N9147, N5730);
not NOT1 (N9154, N9127);
or OR4 (N9155, N9132, N4051, N5796, N6617);
buf BUF1 (N9156, N9153);
or OR4 (N9157, N9139, N6080, N1295, N4541);
xor XOR2 (N9158, N9150, N2977);
and AND4 (N9159, N9158, N7120, N5301, N6834);
and AND3 (N9160, N9151, N5315, N1277);
xor XOR2 (N9161, N9156, N5087);
buf BUF1 (N9162, N9161);
or OR3 (N9163, N9162, N8730, N2997);
not NOT1 (N9164, N9160);
buf BUF1 (N9165, N9152);
buf BUF1 (N9166, N9155);
xor XOR2 (N9167, N9163, N6858);
not NOT1 (N9168, N9154);
buf BUF1 (N9169, N9165);
nor NOR4 (N9170, N9166, N1720, N2702, N4971);
not NOT1 (N9171, N9146);
nor NOR4 (N9172, N9149, N6601, N4893, N4620);
buf BUF1 (N9173, N9168);
not NOT1 (N9174, N9145);
not NOT1 (N9175, N9170);
xor XOR2 (N9176, N9174, N4699);
buf BUF1 (N9177, N9172);
nand NAND4 (N9178, N9164, N3931, N5798, N5694);
not NOT1 (N9179, N9159);
nand NAND4 (N9180, N9157, N9152, N1413, N2383);
or OR4 (N9181, N9173, N1438, N1937, N4530);
xor XOR2 (N9182, N9178, N5070);
xor XOR2 (N9183, N9181, N873);
and AND2 (N9184, N9183, N6108);
not NOT1 (N9185, N9177);
buf BUF1 (N9186, N9175);
not NOT1 (N9187, N9184);
buf BUF1 (N9188, N9171);
not NOT1 (N9189, N9182);
not NOT1 (N9190, N9187);
and AND4 (N9191, N9179, N1098, N6336, N7911);
nand NAND4 (N9192, N9176, N7010, N648, N3372);
not NOT1 (N9193, N9180);
nor NOR3 (N9194, N9169, N6573, N102);
nand NAND3 (N9195, N9193, N5460, N1469);
not NOT1 (N9196, N9186);
or OR4 (N9197, N9194, N2318, N4854, N9066);
not NOT1 (N9198, N9197);
or OR3 (N9199, N9192, N7924, N6030);
nand NAND2 (N9200, N9185, N3253);
buf BUF1 (N9201, N9199);
xor XOR2 (N9202, N9188, N5336);
nor NOR4 (N9203, N9167, N6661, N4956, N4494);
and AND2 (N9204, N9190, N3271);
buf BUF1 (N9205, N9201);
not NOT1 (N9206, N9198);
nand NAND3 (N9207, N9205, N4514, N3810);
not NOT1 (N9208, N9204);
nor NOR2 (N9209, N9202, N4994);
not NOT1 (N9210, N9208);
or OR4 (N9211, N9191, N2951, N2523, N8940);
buf BUF1 (N9212, N9189);
nor NOR2 (N9213, N9212, N5700);
or OR4 (N9214, N9210, N1113, N3468, N1217);
buf BUF1 (N9215, N9209);
buf BUF1 (N9216, N9206);
and AND4 (N9217, N9216, N3487, N8595, N89);
nor NOR3 (N9218, N9214, N9031, N7332);
and AND2 (N9219, N9207, N8868);
or OR4 (N9220, N9211, N6034, N783, N5450);
nand NAND2 (N9221, N9217, N1022);
nor NOR3 (N9222, N9213, N6766, N6873);
nand NAND4 (N9223, N9200, N3810, N6187, N8379);
nor NOR3 (N9224, N9195, N4039, N8523);
nand NAND2 (N9225, N9221, N8129);
buf BUF1 (N9226, N9225);
or OR3 (N9227, N9220, N6358, N5713);
not NOT1 (N9228, N9227);
nand NAND3 (N9229, N9196, N1777, N1021);
buf BUF1 (N9230, N9223);
not NOT1 (N9231, N9222);
buf BUF1 (N9232, N9215);
buf BUF1 (N9233, N9229);
or OR4 (N9234, N9233, N5586, N5809, N2672);
buf BUF1 (N9235, N9226);
and AND3 (N9236, N9234, N4483, N5251);
xor XOR2 (N9237, N9230, N1494);
or OR2 (N9238, N9232, N7961);
and AND2 (N9239, N9236, N6894);
buf BUF1 (N9240, N9218);
not NOT1 (N9241, N9219);
or OR2 (N9242, N9237, N8269);
and AND3 (N9243, N9235, N8062, N4667);
nor NOR3 (N9244, N9224, N7838, N8000);
and AND2 (N9245, N9243, N6826);
buf BUF1 (N9246, N9240);
nor NOR4 (N9247, N9203, N1453, N8334, N2054);
buf BUF1 (N9248, N9246);
and AND4 (N9249, N9244, N7681, N323, N7962);
nand NAND2 (N9250, N9248, N6917);
buf BUF1 (N9251, N9238);
nand NAND3 (N9252, N9239, N8677, N5318);
and AND2 (N9253, N9228, N312);
not NOT1 (N9254, N9250);
not NOT1 (N9255, N9231);
or OR3 (N9256, N9252, N6374, N6136);
xor XOR2 (N9257, N9256, N8650);
and AND2 (N9258, N9251, N1002);
or OR3 (N9259, N9242, N4317, N1316);
buf BUF1 (N9260, N9255);
not NOT1 (N9261, N9247);
or OR3 (N9262, N9260, N8985, N142);
not NOT1 (N9263, N9253);
buf BUF1 (N9264, N9241);
or OR4 (N9265, N9249, N4622, N5489, N5951);
xor XOR2 (N9266, N9259, N1016);
nor NOR4 (N9267, N9258, N3293, N5214, N516);
and AND3 (N9268, N9257, N4951, N3937);
xor XOR2 (N9269, N9262, N1657);
or OR2 (N9270, N9267, N5312);
nand NAND4 (N9271, N9254, N6983, N4241, N9106);
nand NAND2 (N9272, N9266, N5628);
not NOT1 (N9273, N9261);
nor NOR4 (N9274, N9245, N2542, N8024, N1149);
xor XOR2 (N9275, N9274, N9142);
xor XOR2 (N9276, N9275, N5693);
xor XOR2 (N9277, N9265, N1667);
nor NOR2 (N9278, N9276, N3776);
or OR2 (N9279, N9270, N2812);
buf BUF1 (N9280, N9277);
xor XOR2 (N9281, N9263, N6861);
nand NAND4 (N9282, N9273, N1969, N1187, N1298);
not NOT1 (N9283, N9278);
or OR2 (N9284, N9283, N8705);
and AND2 (N9285, N9269, N6524);
and AND3 (N9286, N9271, N1207, N2713);
and AND2 (N9287, N9286, N5891);
nand NAND3 (N9288, N9284, N1820, N230);
xor XOR2 (N9289, N9268, N1005);
or OR2 (N9290, N9289, N5705);
or OR2 (N9291, N9279, N8523);
xor XOR2 (N9292, N9282, N9190);
or OR4 (N9293, N9290, N4400, N3718, N6937);
not NOT1 (N9294, N9264);
nor NOR4 (N9295, N9280, N2690, N1645, N6212);
nand NAND3 (N9296, N9281, N7374, N4122);
nor NOR3 (N9297, N9293, N7575, N1859);
nand NAND4 (N9298, N9295, N7015, N8768, N3294);
nor NOR4 (N9299, N9298, N4649, N6542, N3812);
buf BUF1 (N9300, N9285);
or OR3 (N9301, N9300, N3999, N2339);
not NOT1 (N9302, N9288);
nand NAND4 (N9303, N9301, N5757, N978, N3758);
not NOT1 (N9304, N9272);
not NOT1 (N9305, N9292);
buf BUF1 (N9306, N9296);
nand NAND2 (N9307, N9306, N1543);
nand NAND2 (N9308, N9307, N7606);
or OR4 (N9309, N9308, N8809, N7441, N303);
xor XOR2 (N9310, N9291, N2071);
buf BUF1 (N9311, N9302);
or OR4 (N9312, N9303, N9132, N2339, N4451);
xor XOR2 (N9313, N9305, N4572);
not NOT1 (N9314, N9294);
xor XOR2 (N9315, N9314, N8774);
and AND4 (N9316, N9287, N4689, N1357, N7289);
buf BUF1 (N9317, N9297);
xor XOR2 (N9318, N9299, N6683);
xor XOR2 (N9319, N9315, N7897);
buf BUF1 (N9320, N9304);
or OR3 (N9321, N9320, N8676, N579);
not NOT1 (N9322, N9312);
xor XOR2 (N9323, N9310, N457);
not NOT1 (N9324, N9318);
nand NAND2 (N9325, N9322, N6059);
and AND4 (N9326, N9319, N4372, N8983, N6246);
nand NAND2 (N9327, N9311, N5338);
nor NOR3 (N9328, N9309, N6526, N7775);
not NOT1 (N9329, N9325);
nand NAND2 (N9330, N9326, N7998);
nand NAND4 (N9331, N9317, N7618, N6298, N1788);
nand NAND3 (N9332, N9321, N5029, N2734);
nor NOR2 (N9333, N9329, N812);
or OR3 (N9334, N9333, N3758, N8775);
xor XOR2 (N9335, N9332, N3471);
nor NOR3 (N9336, N9331, N6242, N4896);
or OR2 (N9337, N9330, N5200);
xor XOR2 (N9338, N9334, N3928);
nor NOR4 (N9339, N9316, N5315, N775, N7347);
xor XOR2 (N9340, N9337, N3005);
or OR4 (N9341, N9327, N2206, N3377, N1243);
buf BUF1 (N9342, N9323);
nand NAND3 (N9343, N9313, N3587, N4790);
or OR3 (N9344, N9336, N2402, N5769);
xor XOR2 (N9345, N9342, N2378);
nor NOR4 (N9346, N9324, N7970, N587, N3821);
nand NAND2 (N9347, N9343, N8518);
xor XOR2 (N9348, N9341, N9175);
nor NOR4 (N9349, N9344, N2387, N4080, N2494);
or OR4 (N9350, N9338, N6586, N5163, N4095);
or OR3 (N9351, N9340, N8415, N5633);
nand NAND4 (N9352, N9345, N8032, N860, N6476);
not NOT1 (N9353, N9352);
and AND4 (N9354, N9346, N1150, N472, N8292);
and AND3 (N9355, N9339, N3618, N5447);
and AND3 (N9356, N9353, N1227, N166);
xor XOR2 (N9357, N9355, N6147);
or OR4 (N9358, N9357, N6344, N5359, N2746);
and AND3 (N9359, N9348, N7340, N4028);
buf BUF1 (N9360, N9354);
buf BUF1 (N9361, N9359);
xor XOR2 (N9362, N9328, N8087);
or OR2 (N9363, N9358, N5978);
nor NOR3 (N9364, N9350, N7361, N5223);
and AND3 (N9365, N9349, N3332, N418);
and AND3 (N9366, N9364, N1429, N4659);
or OR3 (N9367, N9335, N8399, N2501);
or OR4 (N9368, N9351, N8230, N8172, N6431);
nor NOR3 (N9369, N9360, N1844, N6478);
buf BUF1 (N9370, N9347);
or OR3 (N9371, N9366, N7292, N6545);
nand NAND2 (N9372, N9365, N1446);
xor XOR2 (N9373, N9372, N3763);
buf BUF1 (N9374, N9361);
nand NAND4 (N9375, N9369, N8262, N1378, N2554);
not NOT1 (N9376, N9375);
xor XOR2 (N9377, N9362, N8724);
xor XOR2 (N9378, N9377, N7351);
and AND2 (N9379, N9356, N1440);
or OR4 (N9380, N9379, N4677, N7107, N5577);
xor XOR2 (N9381, N9374, N7498);
or OR3 (N9382, N9380, N8349, N3890);
or OR3 (N9383, N9371, N1217, N6027);
nor NOR4 (N9384, N9373, N8536, N8002, N5683);
not NOT1 (N9385, N9382);
nand NAND2 (N9386, N9384, N3928);
and AND2 (N9387, N9386, N1611);
or OR4 (N9388, N9385, N8024, N69, N4447);
nand NAND2 (N9389, N9378, N3612);
and AND3 (N9390, N9368, N9213, N2606);
not NOT1 (N9391, N9389);
and AND2 (N9392, N9388, N5382);
buf BUF1 (N9393, N9376);
and AND4 (N9394, N9383, N8572, N2415, N8902);
or OR4 (N9395, N9393, N5296, N2876, N7257);
and AND2 (N9396, N9390, N5721);
buf BUF1 (N9397, N9395);
nand NAND4 (N9398, N9367, N2213, N8878, N1157);
or OR4 (N9399, N9363, N6339, N7879, N2834);
buf BUF1 (N9400, N9396);
or OR4 (N9401, N9387, N5136, N4100, N4481);
buf BUF1 (N9402, N9381);
and AND2 (N9403, N9394, N7270);
xor XOR2 (N9404, N9401, N3826);
xor XOR2 (N9405, N9370, N4518);
and AND2 (N9406, N9403, N896);
xor XOR2 (N9407, N9397, N7911);
nor NOR4 (N9408, N9404, N169, N5119, N8299);
not NOT1 (N9409, N9406);
buf BUF1 (N9410, N9392);
xor XOR2 (N9411, N9410, N2498);
not NOT1 (N9412, N9408);
not NOT1 (N9413, N9391);
xor XOR2 (N9414, N9402, N7737);
or OR2 (N9415, N9405, N7182);
nand NAND2 (N9416, N9415, N5813);
nor NOR2 (N9417, N9412, N8668);
nor NOR4 (N9418, N9416, N5173, N3713, N5256);
not NOT1 (N9419, N9398);
and AND3 (N9420, N9414, N3078, N2084);
or OR3 (N9421, N9400, N8018, N2129);
nor NOR3 (N9422, N9420, N7275, N8746);
nand NAND2 (N9423, N9418, N817);
nor NOR3 (N9424, N9413, N6912, N2790);
and AND4 (N9425, N9399, N2575, N1823, N7005);
and AND4 (N9426, N9409, N1414, N6334, N8056);
buf BUF1 (N9427, N9425);
nand NAND2 (N9428, N9419, N5272);
or OR2 (N9429, N9417, N4314);
and AND4 (N9430, N9421, N8817, N7182, N1814);
not NOT1 (N9431, N9428);
or OR2 (N9432, N9427, N6542);
nand NAND2 (N9433, N9426, N604);
nor NOR4 (N9434, N9430, N9150, N5080, N7865);
and AND2 (N9435, N9431, N5192);
nor NOR2 (N9436, N9423, N4834);
not NOT1 (N9437, N9432);
or OR2 (N9438, N9435, N890);
nand NAND2 (N9439, N9436, N1867);
buf BUF1 (N9440, N9433);
buf BUF1 (N9441, N9434);
buf BUF1 (N9442, N9429);
or OR3 (N9443, N9411, N421, N3590);
and AND2 (N9444, N9438, N7857);
or OR3 (N9445, N9437, N5085, N1771);
nand NAND2 (N9446, N9440, N2891);
or OR2 (N9447, N9424, N424);
not NOT1 (N9448, N9407);
nor NOR2 (N9449, N9442, N9414);
or OR4 (N9450, N9449, N8985, N3848, N1990);
and AND2 (N9451, N9444, N8040);
xor XOR2 (N9452, N9441, N8139);
or OR2 (N9453, N9450, N8201);
or OR4 (N9454, N9443, N4671, N4913, N2175);
xor XOR2 (N9455, N9446, N339);
nand NAND3 (N9456, N9451, N1591, N9245);
nor NOR3 (N9457, N9447, N5641, N9348);
or OR2 (N9458, N9448, N443);
nor NOR2 (N9459, N9454, N5405);
buf BUF1 (N9460, N9457);
nand NAND3 (N9461, N9452, N3750, N1093);
nor NOR3 (N9462, N9422, N6950, N7634);
buf BUF1 (N9463, N9455);
not NOT1 (N9464, N9459);
and AND4 (N9465, N9462, N7775, N2165, N7537);
nor NOR2 (N9466, N9464, N2809);
and AND3 (N9467, N9458, N9240, N6549);
xor XOR2 (N9468, N9463, N6285);
xor XOR2 (N9469, N9456, N6593);
and AND2 (N9470, N9465, N817);
buf BUF1 (N9471, N9469);
buf BUF1 (N9472, N9439);
not NOT1 (N9473, N9460);
or OR3 (N9474, N9453, N3789, N1432);
not NOT1 (N9475, N9472);
and AND4 (N9476, N9475, N7052, N2891, N1071);
or OR4 (N9477, N9468, N4168, N5417, N9017);
buf BUF1 (N9478, N9477);
buf BUF1 (N9479, N9473);
xor XOR2 (N9480, N9445, N2462);
not NOT1 (N9481, N9479);
buf BUF1 (N9482, N9481);
xor XOR2 (N9483, N9467, N3987);
or OR3 (N9484, N9461, N8921, N2210);
buf BUF1 (N9485, N9466);
buf BUF1 (N9486, N9485);
not NOT1 (N9487, N9480);
not NOT1 (N9488, N9486);
buf BUF1 (N9489, N9476);
xor XOR2 (N9490, N9474, N3936);
nor NOR3 (N9491, N9482, N2818, N1945);
nand NAND3 (N9492, N9478, N8678, N1770);
buf BUF1 (N9493, N9492);
or OR3 (N9494, N9493, N8144, N2522);
buf BUF1 (N9495, N9489);
nor NOR4 (N9496, N9490, N7368, N6402, N3075);
and AND3 (N9497, N9471, N8534, N3155);
nor NOR4 (N9498, N9470, N6066, N4363, N327);
xor XOR2 (N9499, N9494, N761);
xor XOR2 (N9500, N9498, N4012);
or OR4 (N9501, N9491, N2000, N8965, N9093);
xor XOR2 (N9502, N9499, N3570);
and AND3 (N9503, N9483, N7982, N8675);
or OR4 (N9504, N9500, N8652, N5153, N4229);
and AND3 (N9505, N9487, N1314, N2205);
nor NOR4 (N9506, N9484, N8765, N8444, N2257);
or OR3 (N9507, N9496, N3426, N7864);
buf BUF1 (N9508, N9507);
nor NOR3 (N9509, N9505, N8421, N53);
and AND2 (N9510, N9497, N6679);
nor NOR4 (N9511, N9509, N8056, N6204, N2256);
xor XOR2 (N9512, N9502, N4380);
not NOT1 (N9513, N9503);
and AND4 (N9514, N9511, N1272, N7733, N2412);
xor XOR2 (N9515, N9512, N6515);
buf BUF1 (N9516, N9488);
or OR4 (N9517, N9515, N7596, N3820, N7914);
or OR4 (N9518, N9508, N3273, N6616, N1132);
or OR2 (N9519, N9510, N2448);
nor NOR4 (N9520, N9513, N125, N9095, N6194);
xor XOR2 (N9521, N9516, N7740);
not NOT1 (N9522, N9495);
buf BUF1 (N9523, N9520);
not NOT1 (N9524, N9504);
and AND2 (N9525, N9524, N1045);
not NOT1 (N9526, N9519);
or OR3 (N9527, N9525, N3461, N8859);
and AND3 (N9528, N9506, N9265, N4582);
and AND4 (N9529, N9517, N2085, N8699, N7455);
and AND4 (N9530, N9528, N6497, N606, N7943);
or OR2 (N9531, N9501, N9168);
xor XOR2 (N9532, N9531, N2129);
and AND3 (N9533, N9514, N8198, N7393);
xor XOR2 (N9534, N9523, N5458);
xor XOR2 (N9535, N9532, N6158);
buf BUF1 (N9536, N9521);
not NOT1 (N9537, N9526);
and AND3 (N9538, N9530, N6896, N4423);
nor NOR3 (N9539, N9534, N1124, N4286);
nand NAND2 (N9540, N9529, N2554);
nand NAND2 (N9541, N9539, N6727);
xor XOR2 (N9542, N9541, N988);
buf BUF1 (N9543, N9538);
not NOT1 (N9544, N9535);
not NOT1 (N9545, N9533);
not NOT1 (N9546, N9543);
not NOT1 (N9547, N9527);
and AND2 (N9548, N9540, N1093);
or OR2 (N9549, N9548, N7532);
and AND2 (N9550, N9549, N744);
xor XOR2 (N9551, N9522, N6055);
buf BUF1 (N9552, N9551);
not NOT1 (N9553, N9552);
nand NAND4 (N9554, N9544, N2135, N2075, N3414);
xor XOR2 (N9555, N9537, N7677);
or OR4 (N9556, N9547, N2265, N5274, N8676);
and AND4 (N9557, N9556, N2006, N5195, N8120);
nor NOR2 (N9558, N9550, N8117);
nor NOR3 (N9559, N9518, N4089, N1989);
nor NOR2 (N9560, N9536, N1674);
xor XOR2 (N9561, N9559, N1983);
or OR2 (N9562, N9560, N359);
buf BUF1 (N9563, N9546);
buf BUF1 (N9564, N9545);
nand NAND2 (N9565, N9542, N700);
nand NAND4 (N9566, N9554, N1086, N5582, N3153);
not NOT1 (N9567, N9555);
buf BUF1 (N9568, N9564);
buf BUF1 (N9569, N9565);
and AND3 (N9570, N9561, N6250, N6974);
or OR2 (N9571, N9569, N7955);
nand NAND4 (N9572, N9562, N6735, N1311, N1235);
buf BUF1 (N9573, N9571);
buf BUF1 (N9574, N9573);
nand NAND4 (N9575, N9557, N92, N6934, N9304);
buf BUF1 (N9576, N9572);
nand NAND4 (N9577, N9558, N7978, N1817, N1595);
or OR2 (N9578, N9568, N7600);
and AND3 (N9579, N9563, N2615, N430);
xor XOR2 (N9580, N9570, N1019);
nor NOR3 (N9581, N9567, N1588, N6953);
or OR2 (N9582, N9553, N1145);
not NOT1 (N9583, N9575);
and AND2 (N9584, N9576, N5354);
or OR4 (N9585, N9574, N29, N4068, N614);
not NOT1 (N9586, N9580);
or OR3 (N9587, N9582, N4858, N4079);
nand NAND4 (N9588, N9566, N4258, N609, N7958);
or OR2 (N9589, N9581, N246);
or OR3 (N9590, N9587, N1587, N1772);
and AND4 (N9591, N9590, N2273, N6813, N880);
xor XOR2 (N9592, N9585, N1778);
nor NOR3 (N9593, N9577, N1445, N4361);
buf BUF1 (N9594, N9578);
nor NOR2 (N9595, N9583, N5463);
xor XOR2 (N9596, N9594, N904);
nand NAND2 (N9597, N9592, N952);
xor XOR2 (N9598, N9586, N7311);
nor NOR4 (N9599, N9584, N4793, N1750, N9560);
xor XOR2 (N9600, N9599, N9355);
nor NOR3 (N9601, N9593, N1824, N5858);
and AND4 (N9602, N9588, N8723, N4857, N651);
xor XOR2 (N9603, N9602, N3100);
nor NOR2 (N9604, N9591, N4249);
and AND2 (N9605, N9604, N3817);
buf BUF1 (N9606, N9601);
buf BUF1 (N9607, N9589);
nand NAND4 (N9608, N9596, N1684, N4738, N6108);
nand NAND3 (N9609, N9605, N2114, N3047);
nand NAND4 (N9610, N9600, N244, N1827, N7221);
nand NAND2 (N9611, N9606, N4049);
or OR3 (N9612, N9607, N156, N1827);
nand NAND2 (N9613, N9611, N8606);
nand NAND3 (N9614, N9595, N5813, N9495);
nor NOR3 (N9615, N9579, N7845, N6702);
nand NAND3 (N9616, N9597, N1384, N9526);
nor NOR4 (N9617, N9612, N8031, N5763, N5203);
buf BUF1 (N9618, N9616);
nand NAND2 (N9619, N9598, N7208);
nand NAND2 (N9620, N9617, N8244);
nand NAND2 (N9621, N9609, N5673);
buf BUF1 (N9622, N9603);
and AND4 (N9623, N9621, N9284, N5154, N499);
not NOT1 (N9624, N9622);
nand NAND2 (N9625, N9615, N911);
xor XOR2 (N9626, N9625, N8574);
not NOT1 (N9627, N9619);
nand NAND4 (N9628, N9623, N1151, N1374, N9287);
buf BUF1 (N9629, N9628);
not NOT1 (N9630, N9610);
buf BUF1 (N9631, N9613);
nand NAND2 (N9632, N9614, N8157);
nor NOR2 (N9633, N9630, N3250);
buf BUF1 (N9634, N9633);
nand NAND2 (N9635, N9632, N6455);
xor XOR2 (N9636, N9618, N1494);
not NOT1 (N9637, N9627);
buf BUF1 (N9638, N9626);
buf BUF1 (N9639, N9624);
not NOT1 (N9640, N9608);
not NOT1 (N9641, N9640);
xor XOR2 (N9642, N9635, N2091);
or OR4 (N9643, N9634, N1192, N6989, N927);
nand NAND4 (N9644, N9638, N2812, N9100, N7786);
and AND3 (N9645, N9644, N8334, N3471);
not NOT1 (N9646, N9631);
and AND2 (N9647, N9641, N5092);
buf BUF1 (N9648, N9642);
buf BUF1 (N9649, N9647);
buf BUF1 (N9650, N9620);
nor NOR2 (N9651, N9636, N4507);
nor NOR3 (N9652, N9649, N3884, N1459);
nor NOR4 (N9653, N9652, N2094, N4460, N6064);
nand NAND2 (N9654, N9651, N3696);
and AND4 (N9655, N9654, N6323, N3147, N5257);
xor XOR2 (N9656, N9639, N1414);
buf BUF1 (N9657, N9645);
buf BUF1 (N9658, N9653);
nand NAND2 (N9659, N9658, N5032);
or OR2 (N9660, N9655, N3114);
and AND4 (N9661, N9657, N3657, N2144, N4576);
xor XOR2 (N9662, N9637, N2514);
not NOT1 (N9663, N9656);
xor XOR2 (N9664, N9663, N8442);
nor NOR2 (N9665, N9629, N8423);
not NOT1 (N9666, N9664);
or OR2 (N9667, N9659, N9414);
not NOT1 (N9668, N9661);
not NOT1 (N9669, N9666);
nand NAND2 (N9670, N9668, N6655);
xor XOR2 (N9671, N9667, N9142);
xor XOR2 (N9672, N9671, N7488);
nor NOR4 (N9673, N9648, N906, N3599, N5095);
or OR4 (N9674, N9662, N5368, N1534, N7820);
xor XOR2 (N9675, N9665, N2223);
and AND3 (N9676, N9650, N5322, N5638);
buf BUF1 (N9677, N9672);
nor NOR2 (N9678, N9677, N2080);
or OR2 (N9679, N9646, N6354);
nand NAND4 (N9680, N9670, N4680, N7463, N4008);
buf BUF1 (N9681, N9674);
or OR2 (N9682, N9681, N1187);
and AND2 (N9683, N9660, N6663);
xor XOR2 (N9684, N9643, N2123);
and AND2 (N9685, N9675, N3735);
not NOT1 (N9686, N9673);
buf BUF1 (N9687, N9683);
nand NAND4 (N9688, N9687, N8084, N8942, N9087);
or OR4 (N9689, N9686, N28, N3448, N4619);
or OR4 (N9690, N9679, N9675, N4178, N802);
xor XOR2 (N9691, N9676, N1174);
not NOT1 (N9692, N9669);
nor NOR3 (N9693, N9690, N1432, N549);
not NOT1 (N9694, N9691);
buf BUF1 (N9695, N9678);
nand NAND3 (N9696, N9694, N6915, N4950);
or OR3 (N9697, N9680, N9585, N1025);
buf BUF1 (N9698, N9684);
buf BUF1 (N9699, N9692);
and AND3 (N9700, N9697, N9199, N7302);
buf BUF1 (N9701, N9700);
and AND4 (N9702, N9695, N4405, N7209, N1063);
and AND2 (N9703, N9696, N6807);
nand NAND4 (N9704, N9682, N8377, N9218, N6809);
not NOT1 (N9705, N9703);
buf BUF1 (N9706, N9688);
xor XOR2 (N9707, N9701, N5000);
xor XOR2 (N9708, N9693, N2128);
nand NAND2 (N9709, N9706, N927);
nand NAND2 (N9710, N9705, N575);
xor XOR2 (N9711, N9710, N1876);
xor XOR2 (N9712, N9685, N6965);
or OR3 (N9713, N9708, N7275, N5125);
nor NOR4 (N9714, N9712, N595, N2123, N3577);
nor NOR3 (N9715, N9704, N9242, N9201);
xor XOR2 (N9716, N9702, N7079);
and AND3 (N9717, N9689, N1136, N2318);
nor NOR3 (N9718, N9709, N4649, N1668);
or OR2 (N9719, N9714, N7875);
and AND2 (N9720, N9719, N4180);
nor NOR2 (N9721, N9707, N1360);
and AND3 (N9722, N9715, N5756, N789);
or OR4 (N9723, N9699, N9299, N1873, N4867);
nor NOR2 (N9724, N9717, N246);
not NOT1 (N9725, N9711);
xor XOR2 (N9726, N9723, N9239);
or OR3 (N9727, N9722, N2847, N1596);
not NOT1 (N9728, N9727);
or OR2 (N9729, N9728, N7339);
nand NAND2 (N9730, N9724, N1211);
not NOT1 (N9731, N9729);
xor XOR2 (N9732, N9721, N6460);
buf BUF1 (N9733, N9718);
and AND3 (N9734, N9716, N3025, N8621);
not NOT1 (N9735, N9698);
buf BUF1 (N9736, N9731);
nand NAND2 (N9737, N9726, N8652);
and AND2 (N9738, N9736, N4011);
xor XOR2 (N9739, N9732, N3627);
buf BUF1 (N9740, N9713);
nor NOR4 (N9741, N9730, N5358, N519, N7291);
or OR4 (N9742, N9738, N4681, N1238, N6170);
not NOT1 (N9743, N9740);
nand NAND3 (N9744, N9737, N2746, N1460);
not NOT1 (N9745, N9720);
nand NAND2 (N9746, N9741, N2500);
or OR4 (N9747, N9743, N3343, N706, N195);
not NOT1 (N9748, N9745);
nand NAND2 (N9749, N9747, N6209);
buf BUF1 (N9750, N9725);
buf BUF1 (N9751, N9749);
and AND4 (N9752, N9746, N877, N3862, N8898);
nor NOR4 (N9753, N9744, N1889, N5433, N8135);
xor XOR2 (N9754, N9742, N5662);
and AND2 (N9755, N9752, N2024);
and AND4 (N9756, N9734, N1976, N1550, N8);
xor XOR2 (N9757, N9754, N6262);
buf BUF1 (N9758, N9733);
nand NAND3 (N9759, N9758, N6664, N671);
nor NOR2 (N9760, N9759, N135);
xor XOR2 (N9761, N9760, N9681);
xor XOR2 (N9762, N9750, N7264);
xor XOR2 (N9763, N9762, N7468);
or OR2 (N9764, N9753, N6793);
and AND3 (N9765, N9751, N9463, N5838);
nand NAND3 (N9766, N9748, N6593, N8780);
nor NOR3 (N9767, N9764, N508, N1862);
buf BUF1 (N9768, N9739);
nand NAND3 (N9769, N9757, N3059, N5658);
or OR2 (N9770, N9761, N1455);
buf BUF1 (N9771, N9735);
or OR2 (N9772, N9770, N4719);
nand NAND2 (N9773, N9772, N2113);
and AND4 (N9774, N9768, N3677, N872, N1389);
not NOT1 (N9775, N9763);
nand NAND3 (N9776, N9773, N7691, N8760);
buf BUF1 (N9777, N9775);
or OR3 (N9778, N9774, N9367, N3224);
xor XOR2 (N9779, N9766, N4037);
or OR3 (N9780, N9767, N5194, N2589);
not NOT1 (N9781, N9778);
xor XOR2 (N9782, N9777, N6488);
and AND4 (N9783, N9756, N735, N2154, N65);
nand NAND2 (N9784, N9779, N4581);
nor NOR2 (N9785, N9782, N2643);
buf BUF1 (N9786, N9785);
and AND4 (N9787, N9771, N5040, N3648, N1465);
nor NOR4 (N9788, N9769, N7178, N1746, N435);
nand NAND2 (N9789, N9776, N1903);
or OR3 (N9790, N9780, N2646, N7218);
nand NAND2 (N9791, N9788, N8597);
nand NAND2 (N9792, N9787, N143);
not NOT1 (N9793, N9765);
nor NOR3 (N9794, N9786, N1027, N4108);
or OR2 (N9795, N9790, N6098);
nor NOR4 (N9796, N9781, N3160, N1866, N3179);
and AND4 (N9797, N9789, N2307, N6084, N4507);
xor XOR2 (N9798, N9793, N3978);
xor XOR2 (N9799, N9791, N4956);
xor XOR2 (N9800, N9795, N9673);
not NOT1 (N9801, N9800);
buf BUF1 (N9802, N9794);
or OR2 (N9803, N9798, N2488);
xor XOR2 (N9804, N9783, N3724);
or OR3 (N9805, N9803, N3374, N7054);
not NOT1 (N9806, N9755);
not NOT1 (N9807, N9805);
not NOT1 (N9808, N9796);
not NOT1 (N9809, N9808);
nor NOR3 (N9810, N9809, N5252, N4860);
not NOT1 (N9811, N9804);
xor XOR2 (N9812, N9784, N9192);
and AND3 (N9813, N9802, N116, N2352);
not NOT1 (N9814, N9813);
xor XOR2 (N9815, N9814, N8103);
buf BUF1 (N9816, N9792);
not NOT1 (N9817, N9812);
not NOT1 (N9818, N9807);
and AND3 (N9819, N9817, N5138, N2960);
nand NAND3 (N9820, N9819, N1669, N156);
xor XOR2 (N9821, N9815, N8009);
or OR2 (N9822, N9816, N2950);
and AND4 (N9823, N9806, N3286, N7781, N7229);
and AND3 (N9824, N9818, N3789, N6179);
xor XOR2 (N9825, N9823, N1903);
nor NOR2 (N9826, N9801, N4932);
nand NAND2 (N9827, N9824, N1794);
and AND2 (N9828, N9822, N6564);
nor NOR3 (N9829, N9797, N6898, N4228);
not NOT1 (N9830, N9799);
or OR2 (N9831, N9828, N7538);
nor NOR4 (N9832, N9811, N7933, N6335, N2893);
not NOT1 (N9833, N9830);
nor NOR3 (N9834, N9825, N422, N8879);
and AND3 (N9835, N9833, N6334, N6430);
nor NOR2 (N9836, N9826, N9587);
buf BUF1 (N9837, N9835);
xor XOR2 (N9838, N9834, N2627);
xor XOR2 (N9839, N9836, N8693);
and AND2 (N9840, N9837, N6975);
nor NOR3 (N9841, N9838, N334, N4607);
xor XOR2 (N9842, N9839, N8151);
or OR3 (N9843, N9821, N140, N6441);
xor XOR2 (N9844, N9831, N724);
buf BUF1 (N9845, N9843);
xor XOR2 (N9846, N9840, N6000);
buf BUF1 (N9847, N9845);
not NOT1 (N9848, N9841);
buf BUF1 (N9849, N9847);
nor NOR3 (N9850, N9849, N3103, N2970);
xor XOR2 (N9851, N9810, N2892);
buf BUF1 (N9852, N9848);
nor NOR3 (N9853, N9846, N2512, N3605);
or OR4 (N9854, N9850, N6691, N3120, N6568);
not NOT1 (N9855, N9820);
or OR3 (N9856, N9851, N1602, N7596);
xor XOR2 (N9857, N9827, N65);
xor XOR2 (N9858, N9856, N1391);
and AND4 (N9859, N9858, N6108, N8891, N7150);
and AND2 (N9860, N9853, N6828);
xor XOR2 (N9861, N9855, N1070);
buf BUF1 (N9862, N9844);
nor NOR3 (N9863, N9857, N2427, N1264);
buf BUF1 (N9864, N9863);
and AND3 (N9865, N9852, N8812, N5550);
xor XOR2 (N9866, N9829, N7414);
xor XOR2 (N9867, N9860, N5992);
xor XOR2 (N9868, N9832, N5322);
and AND2 (N9869, N9866, N6031);
and AND3 (N9870, N9842, N7802, N5721);
xor XOR2 (N9871, N9862, N9142);
nand NAND3 (N9872, N9869, N4420, N712);
not NOT1 (N9873, N9872);
not NOT1 (N9874, N9867);
nor NOR3 (N9875, N9871, N7782, N8028);
and AND2 (N9876, N9870, N4492);
or OR4 (N9877, N9874, N8321, N4732, N5682);
nand NAND3 (N9878, N9865, N8892, N926);
or OR3 (N9879, N9873, N8520, N8900);
nor NOR4 (N9880, N9877, N9708, N4529, N9069);
nor NOR2 (N9881, N9864, N3908);
xor XOR2 (N9882, N9880, N5420);
not NOT1 (N9883, N9859);
and AND2 (N9884, N9861, N5591);
nand NAND2 (N9885, N9878, N9253);
nor NOR2 (N9886, N9883, N7979);
nand NAND2 (N9887, N9881, N5642);
xor XOR2 (N9888, N9875, N8923);
and AND4 (N9889, N9854, N145, N606, N9612);
xor XOR2 (N9890, N9886, N7793);
nor NOR3 (N9891, N9890, N9071, N5076);
buf BUF1 (N9892, N9876);
nor NOR3 (N9893, N9868, N9058, N3126);
not NOT1 (N9894, N9888);
and AND4 (N9895, N9893, N6335, N7905, N8355);
not NOT1 (N9896, N9882);
nor NOR4 (N9897, N9892, N5367, N152, N9381);
nor NOR3 (N9898, N9895, N7136, N2683);
nor NOR4 (N9899, N9891, N2564, N6239, N5228);
not NOT1 (N9900, N9885);
xor XOR2 (N9901, N9896, N3048);
nand NAND4 (N9902, N9887, N3850, N9515, N8754);
nand NAND2 (N9903, N9899, N6368);
not NOT1 (N9904, N9889);
not NOT1 (N9905, N9897);
buf BUF1 (N9906, N9905);
or OR3 (N9907, N9901, N7529, N8717);
or OR2 (N9908, N9907, N1952);
nor NOR4 (N9909, N9900, N565, N4141, N4409);
not NOT1 (N9910, N9894);
or OR4 (N9911, N9898, N6001, N1385, N3074);
buf BUF1 (N9912, N9909);
and AND2 (N9913, N9912, N8971);
xor XOR2 (N9914, N9902, N9391);
and AND3 (N9915, N9906, N2866, N8287);
nor NOR2 (N9916, N9914, N6196);
nand NAND3 (N9917, N9910, N4639, N231);
or OR2 (N9918, N9884, N5434);
xor XOR2 (N9919, N9916, N5120);
or OR2 (N9920, N9917, N1273);
nor NOR4 (N9921, N9903, N7275, N2252, N3624);
buf BUF1 (N9922, N9915);
buf BUF1 (N9923, N9920);
nand NAND3 (N9924, N9879, N8892, N2430);
and AND3 (N9925, N9918, N538, N1380);
not NOT1 (N9926, N9911);
nor NOR4 (N9927, N9926, N5522, N8476, N4183);
buf BUF1 (N9928, N9908);
and AND3 (N9929, N9913, N6950, N4618);
xor XOR2 (N9930, N9928, N1036);
not NOT1 (N9931, N9929);
and AND2 (N9932, N9919, N455);
buf BUF1 (N9933, N9932);
nand NAND4 (N9934, N9931, N7614, N2197, N1364);
or OR3 (N9935, N9930, N319, N6903);
not NOT1 (N9936, N9933);
nand NAND3 (N9937, N9924, N6807, N6135);
or OR3 (N9938, N9923, N3817, N5209);
nand NAND2 (N9939, N9934, N7656);
and AND3 (N9940, N9937, N7389, N3477);
buf BUF1 (N9941, N9940);
buf BUF1 (N9942, N9935);
nor NOR3 (N9943, N9941, N2421, N8442);
not NOT1 (N9944, N9927);
xor XOR2 (N9945, N9942, N7231);
not NOT1 (N9946, N9943);
not NOT1 (N9947, N9904);
and AND3 (N9948, N9945, N6874, N7331);
xor XOR2 (N9949, N9947, N9843);
not NOT1 (N9950, N9946);
and AND3 (N9951, N9922, N9759, N8479);
nor NOR4 (N9952, N9938, N6537, N4058, N9019);
nor NOR3 (N9953, N9948, N3679, N5359);
nand NAND4 (N9954, N9949, N8573, N4573, N2811);
or OR3 (N9955, N9952, N8063, N6145);
or OR3 (N9956, N9939, N128, N982);
or OR3 (N9957, N9936, N5241, N396);
buf BUF1 (N9958, N9951);
nor NOR3 (N9959, N9958, N2363, N4653);
not NOT1 (N9960, N9925);
nand NAND2 (N9961, N9957, N8156);
nand NAND3 (N9962, N9960, N9028, N7155);
buf BUF1 (N9963, N9956);
and AND2 (N9964, N9963, N5780);
buf BUF1 (N9965, N9961);
nand NAND4 (N9966, N9950, N1424, N3924, N1236);
and AND4 (N9967, N9954, N720, N2683, N4344);
nor NOR2 (N9968, N9966, N1926);
buf BUF1 (N9969, N9968);
not NOT1 (N9970, N9953);
or OR2 (N9971, N9967, N7908);
nand NAND4 (N9972, N9971, N5934, N8030, N5095);
nor NOR2 (N9973, N9955, N2758);
and AND3 (N9974, N9964, N2232, N1315);
not NOT1 (N9975, N9921);
or OR3 (N9976, N9970, N506, N7305);
nor NOR4 (N9977, N9969, N51, N4712, N4053);
nand NAND2 (N9978, N9973, N106);
and AND3 (N9979, N9972, N9265, N9173);
nor NOR2 (N9980, N9977, N625);
and AND3 (N9981, N9965, N1709, N7847);
nor NOR3 (N9982, N9959, N361, N1270);
not NOT1 (N9983, N9976);
or OR3 (N9984, N9982, N4259, N7204);
or OR4 (N9985, N9962, N1079, N2023, N1822);
buf BUF1 (N9986, N9974);
buf BUF1 (N9987, N9975);
or OR4 (N9988, N9944, N4062, N3620, N6741);
nand NAND3 (N9989, N9984, N5352, N6351);
nor NOR3 (N9990, N9988, N2448, N7010);
nand NAND2 (N9991, N9987, N4020);
nand NAND3 (N9992, N9981, N4011, N5418);
and AND4 (N9993, N9990, N5524, N5517, N908);
and AND3 (N9994, N9986, N7971, N2097);
not NOT1 (N9995, N9994);
not NOT1 (N9996, N9979);
buf BUF1 (N9997, N9993);
and AND2 (N9998, N9997, N8031);
nand NAND2 (N9999, N9991, N712);
xor XOR2 (N10000, N9980, N7108);
nand NAND4 (N10001, N9978, N8052, N9326, N8027);
not NOT1 (N10002, N9996);
and AND3 (N10003, N9992, N3397, N5919);
and AND2 (N10004, N10001, N8167);
nor NOR2 (N10005, N9983, N7699);
nor NOR2 (N10006, N9995, N9131);
xor XOR2 (N10007, N9998, N4742);
and AND2 (N10008, N10003, N7524);
nand NAND3 (N10009, N10008, N6485, N4058);
nor NOR2 (N10010, N10002, N86);
buf BUF1 (N10011, N9999);
not NOT1 (N10012, N9985);
xor XOR2 (N10013, N10007, N8146);
or OR3 (N10014, N10005, N5097, N9127);
xor XOR2 (N10015, N10011, N188);
buf BUF1 (N10016, N9989);
or OR3 (N10017, N10016, N3698, N1138);
and AND3 (N10018, N10013, N2800, N426);
buf BUF1 (N10019, N10015);
or OR2 (N10020, N10009, N4651);
nor NOR2 (N10021, N10010, N5897);
not NOT1 (N10022, N10012);
nand NAND2 (N10023, N10017, N4602);
and AND2 (N10024, N10022, N5872);
or OR3 (N10025, N10014, N2673, N3102);
and AND2 (N10026, N10004, N3699);
xor XOR2 (N10027, N10000, N9139);
xor XOR2 (N10028, N10025, N5174);
nand NAND3 (N10029, N10018, N3921, N2557);
and AND2 (N10030, N10020, N3956);
buf BUF1 (N10031, N10029);
nor NOR2 (N10032, N10019, N4472);
nor NOR4 (N10033, N10026, N2988, N8589, N2666);
or OR4 (N10034, N10032, N2819, N3817, N4071);
and AND2 (N10035, N10033, N2067);
xor XOR2 (N10036, N10031, N825);
nand NAND2 (N10037, N10036, N7091);
and AND2 (N10038, N10024, N6140);
or OR4 (N10039, N10038, N3795, N5623, N2413);
xor XOR2 (N10040, N10028, N2476);
nand NAND2 (N10041, N10027, N1648);
nand NAND3 (N10042, N10041, N7861, N7002);
not NOT1 (N10043, N10039);
nand NAND2 (N10044, N10035, N9325);
nor NOR4 (N10045, N10021, N7968, N7777, N5355);
nor NOR4 (N10046, N10006, N8103, N1264, N6689);
nor NOR3 (N10047, N10042, N9460, N10029);
xor XOR2 (N10048, N10043, N1210);
not NOT1 (N10049, N10044);
nand NAND4 (N10050, N10047, N9413, N9026, N8654);
buf BUF1 (N10051, N10049);
nor NOR4 (N10052, N10037, N4379, N8058, N7693);
and AND2 (N10053, N10045, N4088);
nor NOR3 (N10054, N10051, N4071, N3835);
or OR3 (N10055, N10054, N9663, N5116);
xor XOR2 (N10056, N10053, N9290);
and AND3 (N10057, N10050, N1579, N2805);
nor NOR4 (N10058, N10052, N8597, N1550, N9208);
or OR2 (N10059, N10046, N5);
not NOT1 (N10060, N10056);
xor XOR2 (N10061, N10048, N7544);
xor XOR2 (N10062, N10030, N1551);
or OR2 (N10063, N10061, N3657);
buf BUF1 (N10064, N10063);
not NOT1 (N10065, N10055);
and AND2 (N10066, N10060, N2122);
not NOT1 (N10067, N10023);
xor XOR2 (N10068, N10064, N9161);
buf BUF1 (N10069, N10067);
or OR3 (N10070, N10068, N5069, N5417);
not NOT1 (N10071, N10057);
or OR4 (N10072, N10069, N3250, N4311, N2702);
nor NOR3 (N10073, N10058, N309, N6923);
and AND2 (N10074, N10034, N1855);
buf BUF1 (N10075, N10070);
nand NAND2 (N10076, N10073, N8945);
buf BUF1 (N10077, N10071);
not NOT1 (N10078, N10066);
nand NAND3 (N10079, N10076, N5971, N2493);
or OR2 (N10080, N10062, N3605);
xor XOR2 (N10081, N10072, N6873);
not NOT1 (N10082, N10059);
xor XOR2 (N10083, N10078, N7266);
and AND4 (N10084, N10083, N3626, N2591, N8408);
or OR3 (N10085, N10084, N9293, N3527);
xor XOR2 (N10086, N10075, N8137);
nor NOR2 (N10087, N10065, N5550);
or OR3 (N10088, N10079, N6180, N1880);
or OR3 (N10089, N10074, N8333, N4209);
not NOT1 (N10090, N10077);
not NOT1 (N10091, N10088);
and AND3 (N10092, N10081, N8197, N2166);
nand NAND3 (N10093, N10091, N7103, N5785);
nor NOR3 (N10094, N10090, N8317, N7489);
and AND4 (N10095, N10082, N9121, N4362, N5227);
not NOT1 (N10096, N10095);
buf BUF1 (N10097, N10093);
nor NOR4 (N10098, N10096, N3848, N1977, N1434);
buf BUF1 (N10099, N10040);
nand NAND2 (N10100, N10086, N9986);
or OR2 (N10101, N10097, N7688);
xor XOR2 (N10102, N10089, N3366);
and AND4 (N10103, N10098, N2471, N1124, N4153);
nor NOR2 (N10104, N10100, N5791);
buf BUF1 (N10105, N10094);
xor XOR2 (N10106, N10102, N8447);
nand NAND3 (N10107, N10087, N8977, N307);
or OR2 (N10108, N10101, N3124);
and AND4 (N10109, N10107, N9570, N848, N5544);
nor NOR2 (N10110, N10092, N3372);
and AND4 (N10111, N10106, N6433, N6709, N555);
xor XOR2 (N10112, N10103, N6117);
or OR3 (N10113, N10112, N5970, N7249);
not NOT1 (N10114, N10108);
and AND4 (N10115, N10109, N5215, N1409, N7653);
buf BUF1 (N10116, N10104);
nor NOR2 (N10117, N10115, N4596);
nand NAND4 (N10118, N10085, N5276, N1915, N1389);
or OR2 (N10119, N10111, N4816);
nor NOR3 (N10120, N10099, N9430, N4913);
xor XOR2 (N10121, N10119, N9253);
xor XOR2 (N10122, N10117, N8132);
buf BUF1 (N10123, N10114);
buf BUF1 (N10124, N10120);
nor NOR3 (N10125, N10113, N8399, N255);
not NOT1 (N10126, N10124);
buf BUF1 (N10127, N10105);
and AND4 (N10128, N10118, N4071, N4280, N7232);
and AND3 (N10129, N10080, N7883, N5091);
and AND4 (N10130, N10122, N6181, N5268, N7629);
and AND2 (N10131, N10128, N9944);
nand NAND2 (N10132, N10123, N7466);
or OR2 (N10133, N10127, N1605);
not NOT1 (N10134, N10129);
xor XOR2 (N10135, N10131, N5896);
buf BUF1 (N10136, N10121);
xor XOR2 (N10137, N10110, N6311);
or OR4 (N10138, N10135, N4601, N7367, N8982);
and AND4 (N10139, N10116, N9189, N5364, N3822);
and AND4 (N10140, N10126, N10109, N1487, N1380);
and AND4 (N10141, N10134, N9949, N8967, N3047);
nor NOR4 (N10142, N10139, N2024, N9670, N7102);
buf BUF1 (N10143, N10136);
nand NAND2 (N10144, N10138, N1116);
not NOT1 (N10145, N10125);
not NOT1 (N10146, N10143);
nor NOR4 (N10147, N10146, N9767, N2927, N9539);
xor XOR2 (N10148, N10144, N1640);
and AND4 (N10149, N10145, N4183, N6267, N3402);
or OR2 (N10150, N10142, N2620);
nor NOR3 (N10151, N10137, N3272, N6435);
or OR2 (N10152, N10148, N3305);
nand NAND2 (N10153, N10149, N5388);
nand NAND2 (N10154, N10133, N8839);
xor XOR2 (N10155, N10152, N8099);
or OR4 (N10156, N10140, N5172, N6227, N1817);
xor XOR2 (N10157, N10132, N578);
nand NAND4 (N10158, N10156, N9898, N1870, N1389);
nor NOR4 (N10159, N10154, N5594, N5310, N9210);
xor XOR2 (N10160, N10159, N925);
nor NOR2 (N10161, N10141, N5023);
buf BUF1 (N10162, N10161);
buf BUF1 (N10163, N10155);
not NOT1 (N10164, N10150);
xor XOR2 (N10165, N10151, N548);
not NOT1 (N10166, N10165);
or OR3 (N10167, N10164, N728, N8670);
or OR3 (N10168, N10160, N4574, N8552);
not NOT1 (N10169, N10168);
nand NAND4 (N10170, N10166, N9514, N4486, N3059);
nand NAND4 (N10171, N10153, N4049, N18, N2377);
and AND3 (N10172, N10169, N434, N7963);
buf BUF1 (N10173, N10158);
nor NOR3 (N10174, N10147, N679, N6149);
buf BUF1 (N10175, N10163);
nand NAND4 (N10176, N10130, N8297, N3942, N3660);
or OR3 (N10177, N10171, N3164, N1215);
or OR4 (N10178, N10177, N9705, N10150, N2663);
and AND4 (N10179, N10157, N4341, N723, N138);
or OR2 (N10180, N10173, N5349);
nor NOR2 (N10181, N10179, N7681);
or OR3 (N10182, N10181, N8554, N6203);
or OR3 (N10183, N10167, N3302, N6678);
or OR3 (N10184, N10183, N2722, N9120);
nand NAND4 (N10185, N10184, N543, N8345, N7143);
or OR4 (N10186, N10174, N8090, N4590, N8579);
xor XOR2 (N10187, N10172, N6735);
and AND2 (N10188, N10178, N5182);
buf BUF1 (N10189, N10175);
and AND4 (N10190, N10162, N8012, N3522, N3051);
or OR3 (N10191, N10170, N4920, N329);
or OR3 (N10192, N10185, N4824, N2319);
nor NOR4 (N10193, N10186, N938, N686, N1621);
nor NOR2 (N10194, N10187, N8954);
not NOT1 (N10195, N10188);
nand NAND4 (N10196, N10180, N3468, N1677, N7778);
or OR2 (N10197, N10192, N1803);
nand NAND2 (N10198, N10182, N428);
nand NAND3 (N10199, N10193, N4242, N9136);
nor NOR2 (N10200, N10194, N6559);
xor XOR2 (N10201, N10176, N7362);
not NOT1 (N10202, N10191);
not NOT1 (N10203, N10199);
buf BUF1 (N10204, N10190);
buf BUF1 (N10205, N10204);
not NOT1 (N10206, N10198);
buf BUF1 (N10207, N10197);
xor XOR2 (N10208, N10202, N5367);
nor NOR4 (N10209, N10201, N8688, N7623, N6765);
not NOT1 (N10210, N10200);
buf BUF1 (N10211, N10206);
and AND4 (N10212, N10208, N1551, N4620, N3904);
or OR4 (N10213, N10205, N6388, N3932, N7790);
nand NAND3 (N10214, N10213, N5485, N1312);
nand NAND4 (N10215, N10210, N4681, N10186, N286);
xor XOR2 (N10216, N10211, N132);
buf BUF1 (N10217, N10207);
or OR4 (N10218, N10203, N6718, N7351, N3181);
xor XOR2 (N10219, N10218, N7568);
xor XOR2 (N10220, N10209, N8900);
not NOT1 (N10221, N10212);
nand NAND2 (N10222, N10221, N4618);
nand NAND2 (N10223, N10222, N7725);
nor NOR2 (N10224, N10223, N5588);
buf BUF1 (N10225, N10217);
and AND4 (N10226, N10215, N6504, N8920, N7132);
or OR4 (N10227, N10196, N4491, N9170, N2659);
nor NOR4 (N10228, N10189, N3767, N6726, N2415);
and AND3 (N10229, N10227, N4962, N9667);
not NOT1 (N10230, N10216);
buf BUF1 (N10231, N10224);
or OR2 (N10232, N10220, N7643);
xor XOR2 (N10233, N10219, N126);
or OR3 (N10234, N10228, N4067, N8347);
or OR2 (N10235, N10231, N2567);
and AND4 (N10236, N10232, N7220, N3406, N5990);
nand NAND3 (N10237, N10214, N7683, N8675);
buf BUF1 (N10238, N10235);
nand NAND3 (N10239, N10195, N9305, N9801);
and AND4 (N10240, N10236, N3691, N6525, N6853);
and AND2 (N10241, N10230, N3137);
or OR2 (N10242, N10237, N8863);
xor XOR2 (N10243, N10229, N4664);
and AND3 (N10244, N10233, N3829, N5924);
not NOT1 (N10245, N10226);
nor NOR2 (N10246, N10244, N4668);
nor NOR3 (N10247, N10239, N5350, N9423);
nor NOR3 (N10248, N10247, N1155, N5581);
and AND4 (N10249, N10238, N7959, N5219, N7178);
buf BUF1 (N10250, N10234);
not NOT1 (N10251, N10249);
nand NAND3 (N10252, N10243, N7673, N2162);
not NOT1 (N10253, N10252);
nand NAND3 (N10254, N10253, N4007, N3329);
and AND2 (N10255, N10254, N6411);
xor XOR2 (N10256, N10255, N6328);
or OR3 (N10257, N10240, N9923, N2696);
nor NOR2 (N10258, N10245, N4314);
nand NAND2 (N10259, N10225, N1241);
nand NAND3 (N10260, N10257, N228, N1003);
xor XOR2 (N10261, N10258, N3913);
nor NOR3 (N10262, N10256, N4435, N2886);
or OR4 (N10263, N10262, N7337, N9709, N9443);
and AND4 (N10264, N10251, N1984, N342, N4972);
and AND4 (N10265, N10241, N3448, N4521, N8661);
nor NOR3 (N10266, N10250, N6757, N9357);
not NOT1 (N10267, N10261);
and AND2 (N10268, N10260, N74);
buf BUF1 (N10269, N10259);
nor NOR2 (N10270, N10268, N9537);
and AND2 (N10271, N10263, N1430);
xor XOR2 (N10272, N10265, N5279);
buf BUF1 (N10273, N10264);
nand NAND3 (N10274, N10272, N3370, N9121);
and AND2 (N10275, N10271, N5040);
not NOT1 (N10276, N10270);
buf BUF1 (N10277, N10275);
or OR4 (N10278, N10276, N8704, N5545, N2483);
or OR2 (N10279, N10266, N374);
xor XOR2 (N10280, N10269, N5505);
buf BUF1 (N10281, N10279);
nand NAND3 (N10282, N10274, N989, N6844);
buf BUF1 (N10283, N10278);
or OR3 (N10284, N10267, N8961, N5039);
buf BUF1 (N10285, N10242);
buf BUF1 (N10286, N10248);
nor NOR4 (N10287, N10246, N2784, N8146, N2486);
buf BUF1 (N10288, N10286);
or OR2 (N10289, N10273, N248);
not NOT1 (N10290, N10288);
xor XOR2 (N10291, N10287, N9515);
nor NOR2 (N10292, N10277, N7919);
xor XOR2 (N10293, N10291, N3735);
or OR2 (N10294, N10290, N7230);
buf BUF1 (N10295, N10280);
or OR3 (N10296, N10294, N3152, N3375);
and AND2 (N10297, N10285, N8429);
or OR2 (N10298, N10282, N2498);
buf BUF1 (N10299, N10297);
or OR4 (N10300, N10296, N5099, N8098, N5120);
buf BUF1 (N10301, N10299);
not NOT1 (N10302, N10284);
not NOT1 (N10303, N10301);
and AND3 (N10304, N10283, N4000, N9368);
xor XOR2 (N10305, N10298, N3723);
nand NAND4 (N10306, N10303, N4928, N6876, N645);
not NOT1 (N10307, N10300);
not NOT1 (N10308, N10289);
or OR4 (N10309, N10308, N6650, N5579, N1553);
buf BUF1 (N10310, N10292);
buf BUF1 (N10311, N10295);
nor NOR4 (N10312, N10309, N215, N482, N7871);
not NOT1 (N10313, N10293);
not NOT1 (N10314, N10313);
buf BUF1 (N10315, N10281);
buf BUF1 (N10316, N10310);
or OR3 (N10317, N10314, N4221, N6429);
or OR3 (N10318, N10302, N5355, N373);
or OR2 (N10319, N10317, N3039);
nand NAND2 (N10320, N10305, N5907);
not NOT1 (N10321, N10304);
not NOT1 (N10322, N10315);
nand NAND3 (N10323, N10311, N5673, N2924);
nand NAND3 (N10324, N10306, N1689, N6852);
and AND4 (N10325, N10319, N4447, N2765, N1854);
nor NOR3 (N10326, N10325, N6372, N6556);
buf BUF1 (N10327, N10322);
buf BUF1 (N10328, N10327);
nor NOR3 (N10329, N10323, N9719, N2239);
or OR4 (N10330, N10320, N4730, N7437, N5148);
not NOT1 (N10331, N10329);
and AND2 (N10332, N10321, N4609);
nand NAND4 (N10333, N10318, N8062, N8661, N528);
or OR2 (N10334, N10331, N6517);
not NOT1 (N10335, N10330);
xor XOR2 (N10336, N10334, N7174);
or OR3 (N10337, N10312, N2027, N8406);
nand NAND3 (N10338, N10336, N1979, N483);
nor NOR2 (N10339, N10316, N3027);
buf BUF1 (N10340, N10328);
nand NAND3 (N10341, N10339, N7040, N2615);
nor NOR2 (N10342, N10340, N1917);
nor NOR3 (N10343, N10338, N1308, N5985);
or OR2 (N10344, N10337, N2874);
nand NAND2 (N10345, N10341, N9942);
not NOT1 (N10346, N10335);
or OR2 (N10347, N10333, N4298);
nor NOR4 (N10348, N10324, N1356, N6537, N9802);
not NOT1 (N10349, N10345);
nor NOR2 (N10350, N10344, N732);
nand NAND3 (N10351, N10347, N10125, N9490);
nand NAND3 (N10352, N10343, N2631, N5154);
nor NOR3 (N10353, N10346, N657, N2641);
or OR3 (N10354, N10352, N6054, N6692);
not NOT1 (N10355, N10342);
buf BUF1 (N10356, N10348);
or OR3 (N10357, N10351, N7594, N8631);
not NOT1 (N10358, N10355);
nor NOR2 (N10359, N10357, N7673);
nor NOR2 (N10360, N10358, N8359);
nor NOR3 (N10361, N10356, N574, N3483);
or OR4 (N10362, N10360, N5085, N567, N7230);
or OR4 (N10363, N10350, N10117, N4065, N4547);
buf BUF1 (N10364, N10332);
or OR2 (N10365, N10362, N5291);
and AND4 (N10366, N10354, N3316, N6720, N5926);
xor XOR2 (N10367, N10366, N2005);
nand NAND2 (N10368, N10361, N3636);
xor XOR2 (N10369, N10349, N3603);
xor XOR2 (N10370, N10368, N7471);
not NOT1 (N10371, N10367);
and AND3 (N10372, N10371, N5311, N2703);
or OR3 (N10373, N10363, N606, N6765);
xor XOR2 (N10374, N10326, N7077);
not NOT1 (N10375, N10370);
nand NAND2 (N10376, N10364, N5354);
and AND2 (N10377, N10359, N6257);
and AND2 (N10378, N10353, N6807);
nor NOR2 (N10379, N10378, N7552);
xor XOR2 (N10380, N10376, N9458);
or OR2 (N10381, N10372, N6048);
nor NOR2 (N10382, N10374, N7776);
not NOT1 (N10383, N10380);
and AND2 (N10384, N10381, N9090);
not NOT1 (N10385, N10369);
xor XOR2 (N10386, N10377, N6841);
and AND4 (N10387, N10379, N1687, N1201, N3576);
nor NOR2 (N10388, N10365, N1129);
buf BUF1 (N10389, N10307);
nor NOR2 (N10390, N10373, N3482);
and AND4 (N10391, N10388, N10076, N2306, N7488);
and AND3 (N10392, N10391, N3650, N8965);
xor XOR2 (N10393, N10384, N2473);
and AND4 (N10394, N10392, N6313, N364, N9877);
nor NOR2 (N10395, N10383, N1893);
xor XOR2 (N10396, N10385, N5108);
nor NOR2 (N10397, N10390, N1969);
and AND3 (N10398, N10395, N714, N4207);
nor NOR4 (N10399, N10394, N8190, N4597, N4263);
not NOT1 (N10400, N10393);
buf BUF1 (N10401, N10382);
xor XOR2 (N10402, N10401, N3723);
nand NAND3 (N10403, N10400, N9341, N630);
nor NOR3 (N10404, N10398, N9307, N1079);
nor NOR3 (N10405, N10403, N1335, N7097);
buf BUF1 (N10406, N10387);
and AND4 (N10407, N10404, N2984, N9109, N8287);
not NOT1 (N10408, N10399);
not NOT1 (N10409, N10386);
or OR4 (N10410, N10397, N901, N4353, N5931);
buf BUF1 (N10411, N10410);
nand NAND2 (N10412, N10402, N8049);
nand NAND3 (N10413, N10405, N6613, N7292);
xor XOR2 (N10414, N10411, N201);
nor NOR2 (N10415, N10396, N747);
or OR3 (N10416, N10412, N120, N5542);
nand NAND2 (N10417, N10415, N10393);
nor NOR2 (N10418, N10408, N9206);
buf BUF1 (N10419, N10418);
not NOT1 (N10420, N10375);
or OR3 (N10421, N10420, N8502, N4595);
and AND4 (N10422, N10406, N3817, N7483, N4648);
xor XOR2 (N10423, N10389, N1108);
nand NAND3 (N10424, N10414, N1480, N435);
xor XOR2 (N10425, N10422, N8422);
nor NOR3 (N10426, N10423, N2243, N2139);
xor XOR2 (N10427, N10424, N8034);
nor NOR4 (N10428, N10426, N4379, N6276, N1054);
and AND2 (N10429, N10427, N3638);
not NOT1 (N10430, N10421);
or OR4 (N10431, N10416, N3187, N3185, N8596);
nor NOR3 (N10432, N10413, N5955, N5882);
or OR3 (N10433, N10432, N9211, N406);
nand NAND4 (N10434, N10433, N614, N3311, N4609);
nand NAND3 (N10435, N10434, N6790, N10306);
buf BUF1 (N10436, N10435);
nor NOR4 (N10437, N10436, N6109, N5585, N7737);
nand NAND3 (N10438, N10431, N6559, N8377);
or OR4 (N10439, N10429, N2700, N3251, N7083);
or OR4 (N10440, N10437, N10349, N7611, N6433);
buf BUF1 (N10441, N10407);
xor XOR2 (N10442, N10438, N3492);
nor NOR2 (N10443, N10442, N2048);
xor XOR2 (N10444, N10439, N5790);
not NOT1 (N10445, N10417);
or OR3 (N10446, N10445, N3476, N262);
not NOT1 (N10447, N10444);
buf BUF1 (N10448, N10443);
or OR2 (N10449, N10447, N2655);
buf BUF1 (N10450, N10446);
buf BUF1 (N10451, N10450);
buf BUF1 (N10452, N10428);
nor NOR2 (N10453, N10441, N9537);
buf BUF1 (N10454, N10419);
or OR3 (N10455, N10449, N201, N6490);
nor NOR3 (N10456, N10452, N5651, N5400);
or OR2 (N10457, N10454, N6165);
nand NAND3 (N10458, N10448, N9554, N6515);
nor NOR4 (N10459, N10457, N575, N6740, N3199);
not NOT1 (N10460, N10459);
buf BUF1 (N10461, N10460);
and AND3 (N10462, N10461, N3447, N5186);
buf BUF1 (N10463, N10425);
xor XOR2 (N10464, N10451, N3313);
not NOT1 (N10465, N10409);
buf BUF1 (N10466, N10430);
buf BUF1 (N10467, N10458);
not NOT1 (N10468, N10455);
not NOT1 (N10469, N10464);
or OR2 (N10470, N10462, N2773);
or OR2 (N10471, N10469, N9995);
nand NAND2 (N10472, N10468, N2224);
nor NOR4 (N10473, N10463, N3195, N4197, N3421);
nand NAND2 (N10474, N10465, N3771);
and AND4 (N10475, N10473, N2091, N4306, N2411);
xor XOR2 (N10476, N10467, N8469);
xor XOR2 (N10477, N10476, N1475);
not NOT1 (N10478, N10453);
nor NOR2 (N10479, N10466, N2554);
not NOT1 (N10480, N10471);
and AND2 (N10481, N10472, N2503);
or OR3 (N10482, N10475, N5020, N3821);
nand NAND4 (N10483, N10470, N2340, N5916, N10221);
buf BUF1 (N10484, N10482);
or OR3 (N10485, N10484, N3355, N1041);
nor NOR4 (N10486, N10483, N3085, N333, N6151);
xor XOR2 (N10487, N10478, N1015);
nor NOR3 (N10488, N10479, N7201, N5869);
xor XOR2 (N10489, N10486, N7542);
xor XOR2 (N10490, N10488, N5931);
xor XOR2 (N10491, N10456, N7511);
buf BUF1 (N10492, N10474);
nor NOR4 (N10493, N10485, N3114, N1176, N3907);
nand NAND3 (N10494, N10481, N8397, N4032);
nand NAND2 (N10495, N10440, N4379);
and AND3 (N10496, N10495, N7186, N5814);
not NOT1 (N10497, N10492);
nand NAND4 (N10498, N10496, N9627, N4351, N3365);
not NOT1 (N10499, N10494);
and AND4 (N10500, N10493, N342, N3073, N6173);
nand NAND2 (N10501, N10500, N9293);
nand NAND4 (N10502, N10491, N4789, N6553, N4587);
or OR2 (N10503, N10502, N5552);
and AND4 (N10504, N10497, N9887, N2900, N3036);
xor XOR2 (N10505, N10490, N565);
xor XOR2 (N10506, N10504, N3089);
and AND3 (N10507, N10499, N2781, N5258);
nor NOR3 (N10508, N10501, N104, N7957);
or OR3 (N10509, N10487, N1860, N5277);
not NOT1 (N10510, N10498);
not NOT1 (N10511, N10489);
xor XOR2 (N10512, N10510, N1134);
not NOT1 (N10513, N10506);
nand NAND3 (N10514, N10511, N6796, N10296);
buf BUF1 (N10515, N10507);
nor NOR4 (N10516, N10513, N6427, N2942, N385);
and AND2 (N10517, N10477, N9426);
nor NOR3 (N10518, N10503, N6958, N5582);
buf BUF1 (N10519, N10512);
nor NOR4 (N10520, N10518, N8777, N5268, N6004);
buf BUF1 (N10521, N10515);
not NOT1 (N10522, N10514);
not NOT1 (N10523, N10520);
xor XOR2 (N10524, N10508, N3926);
xor XOR2 (N10525, N10509, N8942);
not NOT1 (N10526, N10505);
nor NOR3 (N10527, N10522, N9810, N7668);
xor XOR2 (N10528, N10525, N7623);
or OR2 (N10529, N10524, N2791);
or OR2 (N10530, N10516, N3037);
nor NOR4 (N10531, N10530, N6467, N10192, N4079);
or OR4 (N10532, N10521, N3307, N2162, N9481);
buf BUF1 (N10533, N10532);
or OR3 (N10534, N10533, N5129, N4786);
or OR3 (N10535, N10480, N9347, N5395);
nand NAND3 (N10536, N10535, N9225, N6514);
nor NOR3 (N10537, N10527, N2431, N10293);
not NOT1 (N10538, N10534);
nand NAND4 (N10539, N10536, N3065, N656, N5045);
nand NAND3 (N10540, N10537, N1479, N6363);
and AND3 (N10541, N10519, N9258, N6319);
not NOT1 (N10542, N10539);
xor XOR2 (N10543, N10523, N7544);
not NOT1 (N10544, N10529);
nand NAND3 (N10545, N10544, N3887, N3169);
nand NAND4 (N10546, N10545, N282, N2093, N61);
not NOT1 (N10547, N10546);
nand NAND4 (N10548, N10541, N5130, N2456, N2971);
nand NAND4 (N10549, N10528, N2318, N3859, N5238);
and AND4 (N10550, N10531, N10054, N8518, N6531);
nor NOR2 (N10551, N10550, N3152);
or OR3 (N10552, N10526, N4465, N4245);
not NOT1 (N10553, N10542);
not NOT1 (N10554, N10553);
and AND4 (N10555, N10517, N2194, N2265, N5358);
and AND3 (N10556, N10554, N6412, N2615);
buf BUF1 (N10557, N10549);
nor NOR2 (N10558, N10555, N4397);
and AND4 (N10559, N10552, N628, N3425, N4402);
and AND4 (N10560, N10556, N231, N3393, N8975);
buf BUF1 (N10561, N10543);
or OR2 (N10562, N10551, N8135);
nor NOR2 (N10563, N10560, N7506);
nand NAND2 (N10564, N10558, N7479);
nand NAND4 (N10565, N10559, N9389, N6533, N3199);
buf BUF1 (N10566, N10548);
buf BUF1 (N10567, N10562);
and AND3 (N10568, N10565, N4534, N7525);
nor NOR3 (N10569, N10540, N8387, N9038);
and AND4 (N10570, N10557, N7501, N6918, N1555);
or OR4 (N10571, N10570, N10521, N8794, N2772);
nor NOR2 (N10572, N10569, N5287);
and AND3 (N10573, N10568, N2647, N6304);
not NOT1 (N10574, N10561);
not NOT1 (N10575, N10538);
nand NAND2 (N10576, N10571, N7432);
or OR3 (N10577, N10574, N6362, N3920);
not NOT1 (N10578, N10563);
xor XOR2 (N10579, N10576, N828);
or OR4 (N10580, N10575, N7886, N5384, N9660);
or OR3 (N10581, N10573, N1951, N2202);
not NOT1 (N10582, N10547);
or OR3 (N10583, N10578, N1616, N197);
not NOT1 (N10584, N10579);
buf BUF1 (N10585, N10584);
not NOT1 (N10586, N10581);
nor NOR4 (N10587, N10586, N2390, N7795, N2717);
not NOT1 (N10588, N10583);
buf BUF1 (N10589, N10572);
buf BUF1 (N10590, N10567);
or OR4 (N10591, N10582, N704, N10004, N1731);
buf BUF1 (N10592, N10589);
buf BUF1 (N10593, N10591);
nor NOR2 (N10594, N10577, N6905);
and AND3 (N10595, N10593, N5562, N4232);
and AND4 (N10596, N10595, N3368, N2627, N3253);
buf BUF1 (N10597, N10566);
buf BUF1 (N10598, N10590);
xor XOR2 (N10599, N10592, N7197);
nand NAND4 (N10600, N10594, N2037, N939, N8922);
or OR2 (N10601, N10587, N4662);
and AND2 (N10602, N10597, N8319);
xor XOR2 (N10603, N10599, N9610);
nand NAND4 (N10604, N10588, N9948, N2242, N1958);
nor NOR2 (N10605, N10601, N7105);
xor XOR2 (N10606, N10603, N93);
not NOT1 (N10607, N10585);
xor XOR2 (N10608, N10604, N3524);
and AND3 (N10609, N10598, N760, N10003);
nand NAND4 (N10610, N10596, N5629, N1129, N1727);
buf BUF1 (N10611, N10608);
and AND4 (N10612, N10607, N3306, N2388, N9915);
not NOT1 (N10613, N10606);
and AND2 (N10614, N10600, N4390);
nand NAND3 (N10615, N10613, N7514, N5211);
buf BUF1 (N10616, N10615);
nand NAND4 (N10617, N10610, N5689, N5593, N2755);
nor NOR3 (N10618, N10609, N6522, N9953);
and AND4 (N10619, N10611, N3879, N6392, N7935);
nor NOR3 (N10620, N10564, N8712, N8177);
nand NAND3 (N10621, N10612, N4449, N10611);
xor XOR2 (N10622, N10621, N8526);
nand NAND4 (N10623, N10605, N3731, N6881, N1714);
and AND4 (N10624, N10622, N3866, N3453, N5075);
or OR2 (N10625, N10618, N140);
buf BUF1 (N10626, N10614);
not NOT1 (N10627, N10620);
nand NAND2 (N10628, N10626, N1965);
not NOT1 (N10629, N10624);
nor NOR4 (N10630, N10617, N5244, N6844, N2720);
not NOT1 (N10631, N10619);
and AND4 (N10632, N10629, N9474, N3773, N455);
nor NOR2 (N10633, N10580, N3195);
not NOT1 (N10634, N10628);
xor XOR2 (N10635, N10630, N8940);
buf BUF1 (N10636, N10616);
and AND2 (N10637, N10631, N10048);
or OR2 (N10638, N10633, N6175);
and AND2 (N10639, N10638, N6503);
buf BUF1 (N10640, N10637);
and AND2 (N10641, N10632, N3446);
buf BUF1 (N10642, N10602);
or OR2 (N10643, N10641, N3475);
nand NAND3 (N10644, N10643, N8595, N10052);
nor NOR3 (N10645, N10639, N7742, N533);
buf BUF1 (N10646, N10636);
and AND3 (N10647, N10634, N4293, N8206);
nand NAND4 (N10648, N10647, N9832, N848, N9025);
and AND3 (N10649, N10623, N5950, N5464);
or OR2 (N10650, N10644, N1857);
or OR2 (N10651, N10646, N5198);
nor NOR2 (N10652, N10625, N5180);
buf BUF1 (N10653, N10649);
nor NOR4 (N10654, N10645, N3412, N2547, N2285);
nor NOR3 (N10655, N10650, N5621, N205);
buf BUF1 (N10656, N10642);
not NOT1 (N10657, N10653);
or OR2 (N10658, N10657, N2320);
xor XOR2 (N10659, N10654, N3745);
or OR3 (N10660, N10658, N5980, N5187);
nand NAND2 (N10661, N10652, N3145);
or OR4 (N10662, N10660, N2635, N2974, N9886);
nor NOR3 (N10663, N10627, N8033, N10614);
nor NOR2 (N10664, N10659, N4414);
not NOT1 (N10665, N10648);
xor XOR2 (N10666, N10656, N10647);
nand NAND3 (N10667, N10651, N7785, N3840);
xor XOR2 (N10668, N10666, N6273);
nand NAND3 (N10669, N10665, N6776, N1930);
xor XOR2 (N10670, N10635, N1849);
or OR3 (N10671, N10640, N5223, N8371);
not NOT1 (N10672, N10670);
xor XOR2 (N10673, N10663, N163);
nand NAND2 (N10674, N10669, N767);
and AND4 (N10675, N10668, N6768, N10455, N4801);
not NOT1 (N10676, N10674);
buf BUF1 (N10677, N10676);
and AND3 (N10678, N10667, N8333, N2702);
not NOT1 (N10679, N10672);
not NOT1 (N10680, N10678);
not NOT1 (N10681, N10671);
nor NOR2 (N10682, N10661, N3248);
nor NOR2 (N10683, N10679, N5878);
nand NAND2 (N10684, N10680, N4930);
buf BUF1 (N10685, N10681);
nand NAND3 (N10686, N10682, N311, N5232);
nand NAND4 (N10687, N10685, N9601, N9424, N5300);
buf BUF1 (N10688, N10675);
and AND4 (N10689, N10684, N3316, N9379, N6567);
buf BUF1 (N10690, N10689);
xor XOR2 (N10691, N10664, N4304);
and AND3 (N10692, N10662, N2056, N3227);
and AND4 (N10693, N10688, N1126, N7477, N975);
or OR2 (N10694, N10655, N4789);
nor NOR3 (N10695, N10677, N6963, N5641);
nor NOR4 (N10696, N10683, N5872, N4980, N2812);
or OR2 (N10697, N10673, N10289);
not NOT1 (N10698, N10693);
not NOT1 (N10699, N10690);
nand NAND2 (N10700, N10696, N1740);
nor NOR4 (N10701, N10700, N5380, N7873, N8024);
and AND4 (N10702, N10697, N7574, N1807, N10516);
nand NAND2 (N10703, N10701, N9237);
or OR2 (N10704, N10699, N5351);
nand NAND3 (N10705, N10694, N7653, N2276);
and AND4 (N10706, N10705, N8401, N1601, N4518);
nor NOR3 (N10707, N10691, N8349, N7884);
nor NOR2 (N10708, N10687, N4075);
or OR4 (N10709, N10704, N7510, N1978, N8278);
not NOT1 (N10710, N10706);
nand NAND3 (N10711, N10702, N1147, N10168);
or OR4 (N10712, N10711, N3085, N3330, N282);
not NOT1 (N10713, N10709);
and AND2 (N10714, N10695, N3463);
xor XOR2 (N10715, N10710, N7570);
buf BUF1 (N10716, N10713);
nor NOR2 (N10717, N10703, N2455);
buf BUF1 (N10718, N10698);
nand NAND3 (N10719, N10692, N1235, N3008);
not NOT1 (N10720, N10716);
nor NOR2 (N10721, N10720, N10554);
nor NOR3 (N10722, N10686, N2635, N5588);
nand NAND2 (N10723, N10715, N10479);
and AND2 (N10724, N10712, N1576);
and AND2 (N10725, N10721, N9484);
nor NOR3 (N10726, N10707, N7897, N3747);
not NOT1 (N10727, N10726);
buf BUF1 (N10728, N10727);
xor XOR2 (N10729, N10719, N10473);
buf BUF1 (N10730, N10708);
nor NOR2 (N10731, N10728, N7795);
nand NAND3 (N10732, N10725, N4016, N5113);
buf BUF1 (N10733, N10731);
nor NOR4 (N10734, N10730, N2619, N7423, N7800);
xor XOR2 (N10735, N10722, N1304);
xor XOR2 (N10736, N10733, N1716);
and AND4 (N10737, N10732, N8456, N9508, N1131);
nor NOR4 (N10738, N10723, N8671, N4256, N10483);
nor NOR4 (N10739, N10738, N8821, N8337, N3244);
and AND4 (N10740, N10714, N1217, N6632, N8089);
nor NOR3 (N10741, N10737, N9588, N6412);
xor XOR2 (N10742, N10741, N1048);
xor XOR2 (N10743, N10724, N3855);
and AND4 (N10744, N10729, N5379, N8478, N3230);
buf BUF1 (N10745, N10742);
or OR2 (N10746, N10718, N7696);
or OR2 (N10747, N10739, N6328);
nor NOR2 (N10748, N10746, N9292);
nor NOR2 (N10749, N10745, N6018);
nor NOR3 (N10750, N10743, N8419, N182);
nor NOR3 (N10751, N10717, N2352, N5266);
xor XOR2 (N10752, N10735, N10553);
nand NAND3 (N10753, N10752, N10004, N2321);
buf BUF1 (N10754, N10740);
buf BUF1 (N10755, N10750);
not NOT1 (N10756, N10736);
and AND2 (N10757, N10754, N3608);
and AND2 (N10758, N10755, N1439);
buf BUF1 (N10759, N10747);
not NOT1 (N10760, N10757);
nor NOR3 (N10761, N10744, N5635, N8355);
and AND3 (N10762, N10749, N8377, N4466);
nand NAND3 (N10763, N10734, N258, N583);
nor NOR3 (N10764, N10760, N1562, N5331);
and AND4 (N10765, N10751, N7721, N9420, N3869);
or OR4 (N10766, N10756, N378, N2210, N4490);
xor XOR2 (N10767, N10753, N1491);
and AND3 (N10768, N10766, N6163, N1832);
or OR3 (N10769, N10758, N3674, N7514);
nand NAND2 (N10770, N10763, N4073);
not NOT1 (N10771, N10770);
not NOT1 (N10772, N10762);
xor XOR2 (N10773, N10768, N8363);
nor NOR2 (N10774, N10761, N2857);
and AND2 (N10775, N10774, N8531);
or OR2 (N10776, N10759, N3724);
not NOT1 (N10777, N10767);
or OR2 (N10778, N10775, N7135);
nand NAND2 (N10779, N10771, N608);
buf BUF1 (N10780, N10773);
nand NAND3 (N10781, N10779, N2303, N3901);
or OR3 (N10782, N10765, N151, N920);
and AND2 (N10783, N10776, N2309);
and AND2 (N10784, N10778, N3060);
nor NOR2 (N10785, N10769, N7447);
nor NOR2 (N10786, N10764, N5335);
buf BUF1 (N10787, N10748);
nor NOR2 (N10788, N10782, N3202);
and AND4 (N10789, N10777, N8877, N986, N7858);
not NOT1 (N10790, N10780);
not NOT1 (N10791, N10784);
and AND4 (N10792, N10789, N4295, N1219, N2708);
not NOT1 (N10793, N10785);
xor XOR2 (N10794, N10788, N4494);
or OR2 (N10795, N10793, N4015);
and AND4 (N10796, N10772, N8375, N1431, N9446);
nand NAND3 (N10797, N10792, N1328, N6319);
buf BUF1 (N10798, N10794);
and AND4 (N10799, N10791, N5341, N8252, N8537);
nor NOR2 (N10800, N10781, N5674);
and AND4 (N10801, N10799, N2545, N4959, N5395);
xor XOR2 (N10802, N10797, N6175);
xor XOR2 (N10803, N10787, N5548);
nor NOR3 (N10804, N10798, N9870, N9770);
xor XOR2 (N10805, N10786, N5580);
xor XOR2 (N10806, N10790, N4331);
nor NOR3 (N10807, N10801, N1038, N2881);
buf BUF1 (N10808, N10802);
or OR2 (N10809, N10796, N10686);
and AND2 (N10810, N10803, N7088);
and AND2 (N10811, N10800, N2427);
nor NOR4 (N10812, N10811, N4886, N2499, N1227);
buf BUF1 (N10813, N10805);
nor NOR4 (N10814, N10806, N3833, N432, N6508);
buf BUF1 (N10815, N10795);
not NOT1 (N10816, N10808);
or OR2 (N10817, N10783, N9437);
and AND3 (N10818, N10816, N7806, N5179);
buf BUF1 (N10819, N10817);
and AND3 (N10820, N10813, N4852, N1811);
nand NAND2 (N10821, N10815, N6808);
and AND4 (N10822, N10814, N9507, N5496, N1584);
nor NOR2 (N10823, N10822, N9323);
nand NAND2 (N10824, N10810, N9608);
and AND2 (N10825, N10807, N3541);
xor XOR2 (N10826, N10818, N4769);
or OR2 (N10827, N10821, N6852);
nand NAND4 (N10828, N10804, N4541, N5676, N4999);
nand NAND2 (N10829, N10812, N10710);
xor XOR2 (N10830, N10828, N118);
nor NOR2 (N10831, N10824, N3740);
nor NOR4 (N10832, N10820, N980, N2208, N10768);
and AND4 (N10833, N10830, N3419, N9633, N4504);
not NOT1 (N10834, N10825);
not NOT1 (N10835, N10833);
and AND4 (N10836, N10834, N4967, N271, N8890);
xor XOR2 (N10837, N10832, N2538);
and AND3 (N10838, N10835, N793, N7258);
and AND3 (N10839, N10837, N8566, N6904);
xor XOR2 (N10840, N10826, N197);
and AND4 (N10841, N10838, N10444, N10101, N3735);
buf BUF1 (N10842, N10827);
nor NOR2 (N10843, N10839, N3327);
not NOT1 (N10844, N10840);
and AND3 (N10845, N10819, N4084, N8076);
or OR4 (N10846, N10841, N2682, N5352, N5177);
and AND4 (N10847, N10842, N8163, N6754, N3780);
or OR2 (N10848, N10836, N4567);
or OR3 (N10849, N10831, N9745, N7063);
nand NAND4 (N10850, N10823, N8452, N6571, N9942);
xor XOR2 (N10851, N10846, N4511);
xor XOR2 (N10852, N10844, N10337);
not NOT1 (N10853, N10829);
or OR2 (N10854, N10851, N6068);
and AND2 (N10855, N10854, N8937);
and AND2 (N10856, N10850, N2310);
and AND3 (N10857, N10856, N6190, N3102);
and AND2 (N10858, N10847, N618);
nor NOR3 (N10859, N10858, N2645, N7835);
and AND3 (N10860, N10853, N8066, N10140);
nor NOR3 (N10861, N10849, N2391, N2849);
or OR3 (N10862, N10809, N8520, N9748);
nand NAND4 (N10863, N10861, N2803, N665, N6892);
and AND2 (N10864, N10860, N10581);
and AND2 (N10865, N10857, N7373);
nor NOR4 (N10866, N10864, N8110, N10319, N6858);
not NOT1 (N10867, N10863);
nor NOR2 (N10868, N10845, N5412);
nand NAND3 (N10869, N10867, N4844, N4505);
nor NOR3 (N10870, N10859, N9160, N10700);
xor XOR2 (N10871, N10848, N7508);
nor NOR2 (N10872, N10866, N10202);
nand NAND3 (N10873, N10871, N6440, N1757);
or OR2 (N10874, N10868, N4394);
nand NAND4 (N10875, N10872, N1741, N3738, N8543);
xor XOR2 (N10876, N10875, N7024);
and AND4 (N10877, N10869, N5856, N1514, N1551);
and AND3 (N10878, N10876, N676, N7413);
nor NOR2 (N10879, N10852, N4772);
nor NOR2 (N10880, N10877, N1066);
buf BUF1 (N10881, N10873);
or OR2 (N10882, N10865, N3900);
buf BUF1 (N10883, N10870);
nor NOR4 (N10884, N10881, N29, N4595, N6931);
nand NAND3 (N10885, N10843, N2682, N6493);
or OR3 (N10886, N10878, N1867, N4102);
not NOT1 (N10887, N10874);
not NOT1 (N10888, N10886);
and AND4 (N10889, N10855, N9092, N2178, N6380);
not NOT1 (N10890, N10879);
or OR4 (N10891, N10887, N6193, N9624, N6070);
nand NAND2 (N10892, N10890, N9103);
nand NAND4 (N10893, N10885, N6418, N2317, N1034);
not NOT1 (N10894, N10884);
nand NAND3 (N10895, N10892, N8805, N1070);
xor XOR2 (N10896, N10882, N2952);
and AND4 (N10897, N10880, N922, N9590, N1803);
nor NOR3 (N10898, N10889, N5672, N7284);
not NOT1 (N10899, N10897);
nand NAND4 (N10900, N10893, N6187, N9360, N8494);
nor NOR2 (N10901, N10891, N3370);
buf BUF1 (N10902, N10899);
xor XOR2 (N10903, N10862, N8359);
and AND2 (N10904, N10901, N5502);
nor NOR4 (N10905, N10904, N3187, N2462, N6806);
or OR2 (N10906, N10903, N7138);
not NOT1 (N10907, N10894);
not NOT1 (N10908, N10902);
nand NAND3 (N10909, N10895, N3223, N5395);
and AND2 (N10910, N10883, N10848);
xor XOR2 (N10911, N10900, N7495);
xor XOR2 (N10912, N10896, N7879);
or OR4 (N10913, N10909, N6737, N8889, N5835);
not NOT1 (N10914, N10905);
nand NAND4 (N10915, N10906, N7839, N564, N7438);
or OR4 (N10916, N10911, N9346, N1203, N3247);
nand NAND2 (N10917, N10908, N10079);
xor XOR2 (N10918, N10917, N8390);
nor NOR4 (N10919, N10915, N2702, N3658, N1621);
nor NOR2 (N10920, N10910, N7362);
nand NAND4 (N10921, N10912, N2279, N471, N311);
xor XOR2 (N10922, N10913, N10404);
nand NAND2 (N10923, N10918, N839);
and AND4 (N10924, N10914, N2544, N3323, N5958);
not NOT1 (N10925, N10907);
nand NAND4 (N10926, N10920, N10571, N434, N7987);
and AND4 (N10927, N10923, N5005, N2640, N1909);
or OR4 (N10928, N10888, N6696, N2526, N1876);
buf BUF1 (N10929, N10922);
and AND2 (N10930, N10927, N5753);
not NOT1 (N10931, N10926);
not NOT1 (N10932, N10928);
nand NAND2 (N10933, N10932, N6319);
not NOT1 (N10934, N10919);
buf BUF1 (N10935, N10898);
nor NOR3 (N10936, N10934, N3804, N4253);
nand NAND4 (N10937, N10930, N6548, N2843, N7983);
nor NOR4 (N10938, N10935, N10443, N2586, N5078);
xor XOR2 (N10939, N10929, N63);
nor NOR3 (N10940, N10938, N4357, N6049);
not NOT1 (N10941, N10931);
nor NOR4 (N10942, N10937, N8370, N10245, N3114);
xor XOR2 (N10943, N10940, N7798);
nor NOR4 (N10944, N10921, N7503, N447, N5600);
nand NAND2 (N10945, N10933, N1058);
and AND2 (N10946, N10939, N8137);
xor XOR2 (N10947, N10942, N9471);
nand NAND2 (N10948, N10947, N7217);
nand NAND2 (N10949, N10943, N10059);
buf BUF1 (N10950, N10948);
nand NAND2 (N10951, N10944, N3839);
not NOT1 (N10952, N10945);
nand NAND4 (N10953, N10950, N4779, N10546, N7878);
and AND4 (N10954, N10924, N9995, N7947, N10192);
not NOT1 (N10955, N10954);
nand NAND3 (N10956, N10925, N766, N2689);
not NOT1 (N10957, N10953);
nor NOR3 (N10958, N10916, N9477, N10039);
and AND2 (N10959, N10946, N9120);
or OR2 (N10960, N10941, N8075);
or OR2 (N10961, N10952, N6677);
and AND4 (N10962, N10936, N4444, N5676, N3953);
buf BUF1 (N10963, N10956);
xor XOR2 (N10964, N10958, N5896);
and AND4 (N10965, N10955, N4629, N8983, N8309);
nand NAND3 (N10966, N10964, N1582, N10161);
nor NOR3 (N10967, N10963, N1821, N9876);
xor XOR2 (N10968, N10957, N10652);
or OR3 (N10969, N10959, N6942, N7635);
and AND2 (N10970, N10951, N7222);
nor NOR4 (N10971, N10965, N6001, N8647, N3776);
buf BUF1 (N10972, N10968);
buf BUF1 (N10973, N10960);
xor XOR2 (N10974, N10962, N4774);
not NOT1 (N10975, N10961);
or OR2 (N10976, N10975, N7608);
not NOT1 (N10977, N10976);
or OR3 (N10978, N10973, N890, N3290);
nor NOR3 (N10979, N10971, N6714, N10836);
and AND2 (N10980, N10979, N4191);
buf BUF1 (N10981, N10949);
not NOT1 (N10982, N10970);
or OR4 (N10983, N10981, N545, N5989, N347);
nand NAND3 (N10984, N10972, N8311, N5451);
nand NAND2 (N10985, N10966, N4888);
and AND2 (N10986, N10977, N6590);
nand NAND4 (N10987, N10983, N5439, N1427, N20);
nor NOR3 (N10988, N10974, N8081, N4006);
not NOT1 (N10989, N10988);
and AND4 (N10990, N10989, N7070, N5441, N41);
or OR3 (N10991, N10978, N3625, N9654);
and AND3 (N10992, N10985, N3180, N2024);
and AND2 (N10993, N10967, N7581);
or OR2 (N10994, N10982, N431);
buf BUF1 (N10995, N10992);
nor NOR2 (N10996, N10995, N6312);
buf BUF1 (N10997, N10991);
nand NAND4 (N10998, N10986, N4581, N10968, N4523);
xor XOR2 (N10999, N10994, N61);
or OR3 (N11000, N10998, N5315, N3191);
and AND4 (N11001, N10980, N9898, N8009, N9247);
xor XOR2 (N11002, N10990, N1174);
nor NOR2 (N11003, N10984, N792);
nor NOR3 (N11004, N10993, N4101, N4825);
or OR3 (N11005, N11003, N5569, N10726);
nor NOR3 (N11006, N11001, N2914, N5570);
buf BUF1 (N11007, N11000);
or OR3 (N11008, N11007, N3205, N3384);
or OR4 (N11009, N10996, N7363, N8295, N1217);
buf BUF1 (N11010, N11006);
and AND4 (N11011, N11002, N1794, N2809, N7329);
nand NAND3 (N11012, N11009, N10457, N7746);
nand NAND4 (N11013, N10987, N5049, N10140, N9387);
or OR2 (N11014, N11013, N864);
and AND2 (N11015, N11012, N3294);
buf BUF1 (N11016, N11008);
buf BUF1 (N11017, N11005);
or OR2 (N11018, N10999, N8208);
and AND4 (N11019, N11018, N379, N10818, N7391);
nand NAND2 (N11020, N11014, N2780);
nand NAND4 (N11021, N11004, N1758, N341, N7272);
not NOT1 (N11022, N10997);
nor NOR3 (N11023, N11016, N8482, N314);
and AND2 (N11024, N11017, N7902);
not NOT1 (N11025, N11020);
not NOT1 (N11026, N11011);
xor XOR2 (N11027, N11022, N10091);
and AND3 (N11028, N11025, N2056, N1185);
nand NAND3 (N11029, N11028, N8190, N4061);
buf BUF1 (N11030, N11019);
xor XOR2 (N11031, N11024, N521);
and AND2 (N11032, N11026, N7273);
or OR4 (N11033, N11010, N6259, N3505, N10162);
or OR3 (N11034, N11027, N3316, N3613);
and AND2 (N11035, N11021, N2360);
nand NAND3 (N11036, N11015, N5455, N3415);
and AND2 (N11037, N11030, N691);
buf BUF1 (N11038, N11034);
xor XOR2 (N11039, N11033, N2369);
or OR4 (N11040, N11038, N25, N1618, N7946);
not NOT1 (N11041, N11039);
and AND3 (N11042, N11041, N2197, N9380);
buf BUF1 (N11043, N11031);
nand NAND3 (N11044, N11032, N9181, N4990);
and AND3 (N11045, N10969, N6670, N2284);
nand NAND2 (N11046, N11044, N3598);
buf BUF1 (N11047, N11023);
not NOT1 (N11048, N11029);
and AND4 (N11049, N11048, N9241, N125, N6944);
xor XOR2 (N11050, N11043, N6451);
and AND3 (N11051, N11049, N4800, N3837);
and AND3 (N11052, N11040, N7058, N9166);
nor NOR4 (N11053, N11042, N5027, N6271, N454);
and AND2 (N11054, N11045, N10502);
nand NAND4 (N11055, N11046, N9630, N4469, N6468);
buf BUF1 (N11056, N11047);
xor XOR2 (N11057, N11037, N5889);
not NOT1 (N11058, N11051);
not NOT1 (N11059, N11053);
buf BUF1 (N11060, N11059);
xor XOR2 (N11061, N11056, N6933);
or OR4 (N11062, N11054, N318, N1946, N836);
nand NAND3 (N11063, N11057, N8964, N8016);
buf BUF1 (N11064, N11035);
xor XOR2 (N11065, N11060, N10838);
not NOT1 (N11066, N11065);
nand NAND4 (N11067, N11058, N3198, N3389, N4783);
xor XOR2 (N11068, N11061, N3565);
and AND3 (N11069, N11036, N10088, N4200);
xor XOR2 (N11070, N11067, N2543);
nor NOR3 (N11071, N11050, N1967, N5173);
nor NOR2 (N11072, N11064, N8412);
nand NAND4 (N11073, N11063, N6132, N5937, N725);
buf BUF1 (N11074, N11052);
or OR2 (N11075, N11073, N3093);
nor NOR4 (N11076, N11071, N9459, N4455, N2078);
buf BUF1 (N11077, N11066);
and AND2 (N11078, N11072, N6328);
or OR4 (N11079, N11076, N10241, N4891, N3363);
and AND2 (N11080, N11069, N2506);
nor NOR2 (N11081, N11070, N2265);
nor NOR3 (N11082, N11055, N3625, N8412);
buf BUF1 (N11083, N11062);
not NOT1 (N11084, N11083);
or OR3 (N11085, N11078, N9750, N10879);
not NOT1 (N11086, N11077);
buf BUF1 (N11087, N11074);
buf BUF1 (N11088, N11082);
nor NOR4 (N11089, N11080, N5659, N8480, N3974);
nor NOR4 (N11090, N11089, N5116, N6540, N8573);
nor NOR2 (N11091, N11087, N4864);
buf BUF1 (N11092, N11085);
nor NOR2 (N11093, N11068, N4035);
nor NOR4 (N11094, N11093, N690, N4968, N7275);
buf BUF1 (N11095, N11079);
not NOT1 (N11096, N11081);
buf BUF1 (N11097, N11095);
nor NOR4 (N11098, N11086, N1014, N8134, N2379);
xor XOR2 (N11099, N11094, N6987);
xor XOR2 (N11100, N11096, N5101);
buf BUF1 (N11101, N11075);
nor NOR4 (N11102, N11097, N10038, N9628, N3256);
buf BUF1 (N11103, N11090);
not NOT1 (N11104, N11103);
nor NOR4 (N11105, N11101, N8867, N10539, N8755);
and AND3 (N11106, N11100, N221, N4281);
not NOT1 (N11107, N11084);
not NOT1 (N11108, N11088);
and AND4 (N11109, N11092, N7871, N6094, N2282);
or OR2 (N11110, N11102, N8928);
not NOT1 (N11111, N11091);
xor XOR2 (N11112, N11108, N6529);
or OR4 (N11113, N11112, N7652, N5425, N7733);
buf BUF1 (N11114, N11109);
xor XOR2 (N11115, N11104, N4355);
and AND4 (N11116, N11113, N8834, N1209, N4598);
or OR2 (N11117, N11105, N9955);
xor XOR2 (N11118, N11099, N5700);
and AND3 (N11119, N11118, N1288, N10286);
nand NAND4 (N11120, N11098, N9707, N344, N2595);
nor NOR4 (N11121, N11106, N11091, N7282, N10082);
and AND2 (N11122, N11117, N8636);
nand NAND2 (N11123, N11116, N5773);
nand NAND4 (N11124, N11110, N10993, N1021, N9356);
xor XOR2 (N11125, N11119, N9468);
not NOT1 (N11126, N11120);
buf BUF1 (N11127, N11126);
xor XOR2 (N11128, N11123, N9288);
nor NOR4 (N11129, N11122, N10134, N10589, N692);
nor NOR2 (N11130, N11111, N3071);
nor NOR3 (N11131, N11114, N7158, N6800);
nor NOR3 (N11132, N11130, N3631, N7299);
nor NOR3 (N11133, N11132, N8073, N4891);
buf BUF1 (N11134, N11131);
xor XOR2 (N11135, N11125, N9839);
and AND4 (N11136, N11124, N3526, N4911, N1443);
nor NOR3 (N11137, N11133, N1577, N7988);
or OR2 (N11138, N11135, N9336);
nor NOR2 (N11139, N11115, N1424);
and AND4 (N11140, N11129, N7744, N1970, N888);
buf BUF1 (N11141, N11128);
nor NOR3 (N11142, N11127, N615, N2097);
or OR2 (N11143, N11140, N9793);
or OR3 (N11144, N11107, N540, N6015);
and AND2 (N11145, N11143, N3516);
xor XOR2 (N11146, N11139, N4925);
xor XOR2 (N11147, N11145, N7171);
nand NAND2 (N11148, N11134, N1885);
nand NAND4 (N11149, N11144, N3015, N1806, N304);
buf BUF1 (N11150, N11146);
xor XOR2 (N11151, N11149, N9709);
and AND2 (N11152, N11147, N4203);
xor XOR2 (N11153, N11151, N2162);
xor XOR2 (N11154, N11137, N1538);
nand NAND4 (N11155, N11154, N5244, N9031, N6402);
buf BUF1 (N11156, N11142);
and AND4 (N11157, N11138, N5053, N4663, N8284);
xor XOR2 (N11158, N11121, N7417);
nor NOR4 (N11159, N11153, N1554, N7775, N973);
nand NAND4 (N11160, N11155, N2860, N871, N3751);
or OR3 (N11161, N11148, N8711, N5465);
xor XOR2 (N11162, N11150, N3368);
or OR4 (N11163, N11159, N4498, N9335, N11010);
buf BUF1 (N11164, N11152);
buf BUF1 (N11165, N11157);
not NOT1 (N11166, N11161);
and AND3 (N11167, N11160, N4766, N10814);
buf BUF1 (N11168, N11167);
nand NAND4 (N11169, N11165, N6153, N7990, N1967);
not NOT1 (N11170, N11156);
buf BUF1 (N11171, N11169);
not NOT1 (N11172, N11164);
buf BUF1 (N11173, N11172);
nor NOR4 (N11174, N11163, N6301, N7783, N6266);
xor XOR2 (N11175, N11158, N2915);
nand NAND3 (N11176, N11175, N4265, N8916);
not NOT1 (N11177, N11136);
or OR2 (N11178, N11176, N2004);
xor XOR2 (N11179, N11178, N1042);
and AND2 (N11180, N11162, N8483);
nand NAND2 (N11181, N11180, N10748);
nand NAND2 (N11182, N11181, N9303);
nand NAND4 (N11183, N11141, N3838, N9621, N7979);
nand NAND3 (N11184, N11173, N794, N6218);
not NOT1 (N11185, N11168);
nand NAND3 (N11186, N11182, N7431, N580);
xor XOR2 (N11187, N11166, N8633);
buf BUF1 (N11188, N11187);
or OR3 (N11189, N11174, N3439, N2274);
and AND2 (N11190, N11184, N10341);
or OR3 (N11191, N11177, N8566, N3225);
not NOT1 (N11192, N11188);
and AND4 (N11193, N11190, N7063, N5507, N10698);
buf BUF1 (N11194, N11185);
not NOT1 (N11195, N11183);
or OR2 (N11196, N11194, N11148);
not NOT1 (N11197, N11195);
not NOT1 (N11198, N11179);
not NOT1 (N11199, N11191);
xor XOR2 (N11200, N11189, N7352);
xor XOR2 (N11201, N11196, N7324);
not NOT1 (N11202, N11197);
xor XOR2 (N11203, N11192, N7899);
nor NOR4 (N11204, N11170, N8936, N10347, N5001);
and AND2 (N11205, N11186, N624);
nand NAND2 (N11206, N11200, N2847);
buf BUF1 (N11207, N11203);
xor XOR2 (N11208, N11207, N6036);
xor XOR2 (N11209, N11198, N6089);
xor XOR2 (N11210, N11204, N5634);
and AND3 (N11211, N11210, N1945, N9016);
not NOT1 (N11212, N11208);
xor XOR2 (N11213, N11209, N341);
buf BUF1 (N11214, N11212);
xor XOR2 (N11215, N11211, N5320);
and AND3 (N11216, N11171, N1830, N6803);
nand NAND4 (N11217, N11193, N6296, N7530, N7128);
nor NOR3 (N11218, N11216, N10030, N10923);
xor XOR2 (N11219, N11202, N10010);
xor XOR2 (N11220, N11217, N5084);
not NOT1 (N11221, N11220);
and AND2 (N11222, N11218, N3528);
not NOT1 (N11223, N11221);
xor XOR2 (N11224, N11215, N2610);
buf BUF1 (N11225, N11213);
and AND4 (N11226, N11222, N1712, N5467, N7109);
nand NAND2 (N11227, N11214, N1579);
nand NAND4 (N11228, N11219, N7959, N9579, N6168);
nor NOR2 (N11229, N11227, N6249);
xor XOR2 (N11230, N11223, N4290);
buf BUF1 (N11231, N11228);
or OR4 (N11232, N11231, N3672, N2043, N3088);
and AND2 (N11233, N11226, N5247);
and AND4 (N11234, N11201, N5672, N2037, N3117);
buf BUF1 (N11235, N11206);
not NOT1 (N11236, N11225);
or OR2 (N11237, N11233, N328);
buf BUF1 (N11238, N11230);
buf BUF1 (N11239, N11232);
buf BUF1 (N11240, N11234);
buf BUF1 (N11241, N11238);
buf BUF1 (N11242, N11237);
and AND2 (N11243, N11224, N2717);
nor NOR4 (N11244, N11239, N3249, N7060, N6329);
xor XOR2 (N11245, N11236, N2125);
not NOT1 (N11246, N11244);
buf BUF1 (N11247, N11243);
and AND3 (N11248, N11229, N7911, N7228);
nor NOR4 (N11249, N11245, N3250, N5302, N2174);
xor XOR2 (N11250, N11241, N10477);
xor XOR2 (N11251, N11242, N9444);
and AND4 (N11252, N11246, N6003, N2256, N3119);
nand NAND3 (N11253, N11247, N6747, N5924);
xor XOR2 (N11254, N11253, N1441);
and AND4 (N11255, N11254, N6295, N7729, N10489);
nand NAND4 (N11256, N11235, N4004, N8483, N11252);
buf BUF1 (N11257, N7081);
nand NAND3 (N11258, N11248, N5063, N6944);
not NOT1 (N11259, N11199);
and AND2 (N11260, N11250, N8525);
and AND4 (N11261, N11240, N1731, N6453, N4025);
nand NAND2 (N11262, N11251, N8042);
not NOT1 (N11263, N11249);
and AND4 (N11264, N11261, N9413, N5379, N2583);
and AND2 (N11265, N11263, N7430);
buf BUF1 (N11266, N11257);
nand NAND3 (N11267, N11264, N3359, N8739);
and AND2 (N11268, N11205, N10855);
not NOT1 (N11269, N11266);
or OR4 (N11270, N11267, N3349, N1715, N7771);
not NOT1 (N11271, N11265);
buf BUF1 (N11272, N11270);
buf BUF1 (N11273, N11269);
nand NAND4 (N11274, N11272, N7668, N4275, N9747);
xor XOR2 (N11275, N11274, N8429);
xor XOR2 (N11276, N11271, N11198);
or OR3 (N11277, N11256, N9890, N8026);
nor NOR3 (N11278, N11255, N1077, N1443);
buf BUF1 (N11279, N11262);
buf BUF1 (N11280, N11259);
nand NAND3 (N11281, N11277, N3175, N6016);
not NOT1 (N11282, N11273);
buf BUF1 (N11283, N11268);
nor NOR2 (N11284, N11283, N8672);
buf BUF1 (N11285, N11279);
buf BUF1 (N11286, N11284);
xor XOR2 (N11287, N11282, N3920);
nor NOR4 (N11288, N11258, N7187, N6826, N6291);
not NOT1 (N11289, N11287);
not NOT1 (N11290, N11288);
nand NAND3 (N11291, N11285, N4019, N7686);
nand NAND4 (N11292, N11280, N7394, N3322, N6190);
or OR4 (N11293, N11275, N6377, N7756, N4709);
nand NAND3 (N11294, N11278, N4789, N6255);
nand NAND2 (N11295, N11294, N8759);
nor NOR4 (N11296, N11286, N1308, N6216, N7024);
xor XOR2 (N11297, N11295, N747);
buf BUF1 (N11298, N11289);
and AND4 (N11299, N11290, N8584, N2433, N5435);
nand NAND3 (N11300, N11296, N8641, N2689);
and AND4 (N11301, N11299, N1067, N4044, N754);
nand NAND2 (N11302, N11260, N507);
nor NOR2 (N11303, N11276, N7629);
or OR3 (N11304, N11301, N6055, N8662);
nand NAND4 (N11305, N11292, N2962, N5722, N6997);
not NOT1 (N11306, N11304);
nand NAND2 (N11307, N11306, N11157);
not NOT1 (N11308, N11307);
or OR4 (N11309, N11281, N11188, N1767, N2966);
xor XOR2 (N11310, N11298, N5298);
or OR4 (N11311, N11308, N9017, N8939, N4382);
nor NOR3 (N11312, N11302, N3964, N6551);
and AND2 (N11313, N11303, N10081);
xor XOR2 (N11314, N11297, N9932);
not NOT1 (N11315, N11312);
xor XOR2 (N11316, N11293, N6566);
nor NOR3 (N11317, N11310, N9369, N7737);
xor XOR2 (N11318, N11317, N154);
xor XOR2 (N11319, N11311, N10497);
buf BUF1 (N11320, N11319);
and AND2 (N11321, N11309, N2960);
nand NAND2 (N11322, N11305, N4141);
xor XOR2 (N11323, N11291, N9901);
not NOT1 (N11324, N11321);
not NOT1 (N11325, N11315);
nand NAND3 (N11326, N11325, N965, N1439);
and AND3 (N11327, N11323, N10294, N3314);
or OR4 (N11328, N11318, N5958, N4666, N3964);
xor XOR2 (N11329, N11300, N3250);
nor NOR4 (N11330, N11328, N8593, N9283, N5088);
buf BUF1 (N11331, N11329);
nor NOR4 (N11332, N11316, N2488, N8940, N9539);
and AND3 (N11333, N11327, N8798, N7787);
and AND3 (N11334, N11332, N216, N4414);
buf BUF1 (N11335, N11331);
not NOT1 (N11336, N11320);
xor XOR2 (N11337, N11333, N9716);
buf BUF1 (N11338, N11322);
buf BUF1 (N11339, N11330);
xor XOR2 (N11340, N11337, N3836);
buf BUF1 (N11341, N11313);
xor XOR2 (N11342, N11335, N1203);
or OR3 (N11343, N11326, N1626, N3772);
xor XOR2 (N11344, N11340, N361);
or OR4 (N11345, N11338, N10563, N3976, N4353);
and AND2 (N11346, N11336, N7787);
not NOT1 (N11347, N11314);
nand NAND3 (N11348, N11345, N6235, N5199);
not NOT1 (N11349, N11334);
nor NOR4 (N11350, N11341, N2754, N5640, N2693);
xor XOR2 (N11351, N11346, N9514);
not NOT1 (N11352, N11349);
not NOT1 (N11353, N11324);
xor XOR2 (N11354, N11350, N10747);
xor XOR2 (N11355, N11342, N10926);
xor XOR2 (N11356, N11354, N9834);
or OR2 (N11357, N11339, N7760);
buf BUF1 (N11358, N11351);
nand NAND2 (N11359, N11343, N10982);
and AND4 (N11360, N11355, N10374, N1191, N4231);
or OR4 (N11361, N11359, N5071, N8529, N2829);
xor XOR2 (N11362, N11353, N7567);
xor XOR2 (N11363, N11360, N5907);
buf BUF1 (N11364, N11358);
and AND2 (N11365, N11362, N9351);
not NOT1 (N11366, N11364);
xor XOR2 (N11367, N11357, N8099);
nor NOR3 (N11368, N11363, N8215, N8636);
nand NAND2 (N11369, N11344, N8442);
buf BUF1 (N11370, N11366);
not NOT1 (N11371, N11348);
not NOT1 (N11372, N11347);
nand NAND4 (N11373, N11361, N11327, N6902, N6659);
nor NOR3 (N11374, N11370, N6100, N3419);
or OR2 (N11375, N11356, N7721);
xor XOR2 (N11376, N11365, N9245);
buf BUF1 (N11377, N11371);
xor XOR2 (N11378, N11352, N2723);
buf BUF1 (N11379, N11373);
nor NOR2 (N11380, N11378, N7271);
nand NAND4 (N11381, N11374, N8436, N8288, N7058);
xor XOR2 (N11382, N11376, N2195);
not NOT1 (N11383, N11377);
and AND4 (N11384, N11372, N673, N1193, N6500);
nand NAND3 (N11385, N11384, N8787, N5947);
buf BUF1 (N11386, N11381);
nor NOR2 (N11387, N11375, N5743);
buf BUF1 (N11388, N11386);
xor XOR2 (N11389, N11383, N6937);
nand NAND2 (N11390, N11382, N10472);
or OR2 (N11391, N11389, N5883);
not NOT1 (N11392, N11367);
xor XOR2 (N11393, N11387, N10400);
nand NAND4 (N11394, N11380, N575, N4947, N4544);
nand NAND3 (N11395, N11391, N10933, N8721);
xor XOR2 (N11396, N11379, N3612);
buf BUF1 (N11397, N11390);
nor NOR2 (N11398, N11394, N11371);
buf BUF1 (N11399, N11368);
and AND3 (N11400, N11393, N1843, N9592);
buf BUF1 (N11401, N11399);
and AND2 (N11402, N11398, N3810);
nand NAND3 (N11403, N11388, N9512, N10250);
or OR3 (N11404, N11397, N2910, N8064);
buf BUF1 (N11405, N11385);
buf BUF1 (N11406, N11400);
buf BUF1 (N11407, N11401);
nor NOR4 (N11408, N11403, N6092, N5412, N5687);
or OR4 (N11409, N11392, N7972, N5617, N6671);
or OR3 (N11410, N11404, N7926, N5812);
and AND2 (N11411, N11395, N3958);
nand NAND2 (N11412, N11402, N7023);
nor NOR4 (N11413, N11412, N8329, N6312, N497);
xor XOR2 (N11414, N11409, N153);
and AND3 (N11415, N11406, N2444, N2331);
xor XOR2 (N11416, N11396, N10594);
nor NOR3 (N11417, N11408, N1450, N1753);
not NOT1 (N11418, N11369);
nand NAND3 (N11419, N11410, N5929, N33);
not NOT1 (N11420, N11415);
not NOT1 (N11421, N11405);
nor NOR2 (N11422, N11416, N4523);
or OR2 (N11423, N11421, N2775);
nor NOR3 (N11424, N11417, N4606, N8238);
or OR4 (N11425, N11419, N1558, N4902, N4187);
xor XOR2 (N11426, N11414, N4931);
not NOT1 (N11427, N11425);
buf BUF1 (N11428, N11407);
xor XOR2 (N11429, N11422, N6450);
nor NOR4 (N11430, N11423, N1446, N2993, N1894);
xor XOR2 (N11431, N11427, N6156);
not NOT1 (N11432, N11429);
xor XOR2 (N11433, N11426, N2989);
nor NOR3 (N11434, N11413, N3551, N3054);
buf BUF1 (N11435, N11430);
and AND2 (N11436, N11411, N1406);
or OR2 (N11437, N11436, N8561);
buf BUF1 (N11438, N11432);
nand NAND4 (N11439, N11424, N4783, N5667, N4068);
nand NAND4 (N11440, N11437, N11001, N8842, N6424);
not NOT1 (N11441, N11420);
or OR2 (N11442, N11435, N6774);
nand NAND3 (N11443, N11441, N1223, N7900);
xor XOR2 (N11444, N11438, N9070);
and AND2 (N11445, N11440, N2437);
and AND4 (N11446, N11418, N6403, N9632, N6338);
buf BUF1 (N11447, N11442);
not NOT1 (N11448, N11434);
or OR2 (N11449, N11448, N7476);
nor NOR4 (N11450, N11447, N3112, N248, N8651);
xor XOR2 (N11451, N11433, N9580);
nand NAND3 (N11452, N11431, N4310, N5095);
and AND2 (N11453, N11439, N1707);
buf BUF1 (N11454, N11444);
and AND4 (N11455, N11454, N11398, N5899, N4454);
nor NOR2 (N11456, N11451, N9544);
xor XOR2 (N11457, N11428, N10683);
and AND3 (N11458, N11453, N3554, N1484);
and AND4 (N11459, N11457, N8563, N9704, N4716);
buf BUF1 (N11460, N11446);
or OR4 (N11461, N11459, N9291, N10753, N2827);
not NOT1 (N11462, N11445);
or OR3 (N11463, N11456, N10966, N10300);
xor XOR2 (N11464, N11455, N6838);
not NOT1 (N11465, N11443);
not NOT1 (N11466, N11449);
not NOT1 (N11467, N11461);
xor XOR2 (N11468, N11462, N1223);
buf BUF1 (N11469, N11467);
nand NAND4 (N11470, N11460, N710, N3865, N2380);
buf BUF1 (N11471, N11470);
buf BUF1 (N11472, N11458);
nor NOR2 (N11473, N11450, N6229);
xor XOR2 (N11474, N11452, N9777);
xor XOR2 (N11475, N11466, N4859);
not NOT1 (N11476, N11475);
xor XOR2 (N11477, N11464, N8934);
nand NAND4 (N11478, N11469, N1567, N5235, N10241);
nor NOR2 (N11479, N11473, N5796);
nor NOR4 (N11480, N11472, N2553, N3446, N3942);
nand NAND3 (N11481, N11477, N9073, N7886);
buf BUF1 (N11482, N11478);
not NOT1 (N11483, N11465);
and AND4 (N11484, N11468, N11363, N6297, N5935);
and AND2 (N11485, N11476, N1243);
buf BUF1 (N11486, N11484);
and AND3 (N11487, N11471, N3570, N1043);
nand NAND2 (N11488, N11482, N10326);
nor NOR2 (N11489, N11487, N1933);
and AND4 (N11490, N11483, N159, N3510, N7202);
or OR3 (N11491, N11485, N1388, N1050);
nand NAND4 (N11492, N11474, N8487, N2943, N479);
not NOT1 (N11493, N11481);
and AND3 (N11494, N11480, N6061, N874);
not NOT1 (N11495, N11489);
and AND4 (N11496, N11488, N6058, N11256, N2740);
buf BUF1 (N11497, N11493);
nor NOR2 (N11498, N11496, N3015);
or OR4 (N11499, N11498, N2907, N6412, N2269);
nor NOR3 (N11500, N11486, N7260, N2723);
not NOT1 (N11501, N11494);
nand NAND4 (N11502, N11495, N3686, N1331, N5293);
xor XOR2 (N11503, N11499, N7826);
nor NOR3 (N11504, N11500, N330, N2629);
nor NOR4 (N11505, N11497, N11189, N3077, N6192);
and AND2 (N11506, N11504, N3534);
nor NOR3 (N11507, N11503, N5600, N7771);
not NOT1 (N11508, N11505);
nand NAND4 (N11509, N11508, N6810, N10062, N4968);
or OR2 (N11510, N11509, N3696);
nor NOR4 (N11511, N11507, N4857, N6597, N8875);
xor XOR2 (N11512, N11492, N7101);
buf BUF1 (N11513, N11491);
xor XOR2 (N11514, N11501, N5963);
nand NAND2 (N11515, N11513, N4062);
xor XOR2 (N11516, N11512, N3314);
xor XOR2 (N11517, N11479, N1367);
or OR2 (N11518, N11511, N5577);
xor XOR2 (N11519, N11518, N7500);
nor NOR3 (N11520, N11510, N1473, N9323);
or OR2 (N11521, N11515, N1881);
and AND4 (N11522, N11516, N2660, N5897, N636);
not NOT1 (N11523, N11521);
and AND2 (N11524, N11520, N6743);
nand NAND3 (N11525, N11517, N5719, N902);
buf BUF1 (N11526, N11524);
nand NAND2 (N11527, N11463, N5839);
xor XOR2 (N11528, N11502, N2929);
and AND2 (N11529, N11506, N3089);
not NOT1 (N11530, N11522);
or OR3 (N11531, N11528, N7551, N10162);
or OR3 (N11532, N11527, N9700, N9365);
nor NOR4 (N11533, N11490, N1997, N8852, N2079);
and AND3 (N11534, N11525, N1277, N3482);
xor XOR2 (N11535, N11526, N6192);
and AND3 (N11536, N11531, N3560, N4568);
nor NOR2 (N11537, N11533, N8124);
and AND2 (N11538, N11537, N3175);
nor NOR3 (N11539, N11519, N4633, N8115);
nor NOR3 (N11540, N11535, N4828, N5594);
and AND4 (N11541, N11534, N7917, N5031, N3121);
not NOT1 (N11542, N11536);
and AND4 (N11543, N11523, N384, N6549, N11121);
nand NAND2 (N11544, N11541, N549);
nand NAND3 (N11545, N11542, N1879, N1021);
nor NOR2 (N11546, N11530, N2665);
or OR3 (N11547, N11532, N1299, N8553);
nand NAND4 (N11548, N11514, N7573, N2933, N1226);
or OR4 (N11549, N11546, N363, N6797, N10782);
or OR3 (N11550, N11544, N1423, N6645);
not NOT1 (N11551, N11529);
buf BUF1 (N11552, N11540);
nor NOR2 (N11553, N11552, N6773);
not NOT1 (N11554, N11545);
xor XOR2 (N11555, N11549, N6182);
buf BUF1 (N11556, N11551);
xor XOR2 (N11557, N11555, N5066);
and AND3 (N11558, N11539, N11060, N8860);
and AND3 (N11559, N11553, N1437, N5948);
and AND4 (N11560, N11548, N4569, N1247, N11390);
nand NAND2 (N11561, N11559, N4822);
nor NOR3 (N11562, N11554, N11433, N13);
and AND4 (N11563, N11562, N1430, N3318, N3720);
buf BUF1 (N11564, N11556);
or OR3 (N11565, N11538, N7990, N5798);
xor XOR2 (N11566, N11558, N2617);
xor XOR2 (N11567, N11547, N9329);
nand NAND4 (N11568, N11550, N7939, N10354, N4587);
not NOT1 (N11569, N11557);
buf BUF1 (N11570, N11566);
buf BUF1 (N11571, N11567);
not NOT1 (N11572, N11565);
xor XOR2 (N11573, N11572, N10362);
buf BUF1 (N11574, N11569);
and AND3 (N11575, N11564, N8899, N5441);
nor NOR2 (N11576, N11568, N8582);
and AND3 (N11577, N11571, N531, N10332);
not NOT1 (N11578, N11563);
nor NOR4 (N11579, N11578, N11001, N4035, N10929);
and AND3 (N11580, N11543, N8828, N258);
or OR3 (N11581, N11573, N4196, N908);
nand NAND3 (N11582, N11574, N2730, N3981);
nor NOR4 (N11583, N11579, N11290, N130, N8475);
nand NAND3 (N11584, N11570, N2953, N7987);
nand NAND4 (N11585, N11584, N382, N3824, N823);
nand NAND2 (N11586, N11561, N1759);
nand NAND4 (N11587, N11576, N5762, N7373, N9008);
nor NOR3 (N11588, N11587, N1680, N2285);
and AND2 (N11589, N11582, N5645);
nor NOR3 (N11590, N11586, N10895, N6565);
xor XOR2 (N11591, N11583, N8748);
nand NAND3 (N11592, N11581, N8665, N8159);
and AND2 (N11593, N11588, N6966);
nand NAND2 (N11594, N11575, N9675);
nand NAND3 (N11595, N11591, N1952, N7371);
nor NOR2 (N11596, N11577, N8800);
and AND3 (N11597, N11596, N3295, N7920);
or OR4 (N11598, N11592, N8087, N3755, N7072);
nor NOR2 (N11599, N11585, N1300);
nand NAND2 (N11600, N11595, N7744);
nand NAND2 (N11601, N11580, N3575);
buf BUF1 (N11602, N11593);
not NOT1 (N11603, N11601);
not NOT1 (N11604, N11599);
xor XOR2 (N11605, N11560, N664);
nor NOR3 (N11606, N11597, N7486, N6896);
and AND3 (N11607, N11589, N5755, N3863);
or OR2 (N11608, N11607, N4541);
and AND4 (N11609, N11590, N1822, N763, N4711);
not NOT1 (N11610, N11609);
not NOT1 (N11611, N11600);
buf BUF1 (N11612, N11602);
and AND4 (N11613, N11603, N3002, N6876, N796);
buf BUF1 (N11614, N11613);
not NOT1 (N11615, N11604);
nor NOR3 (N11616, N11608, N10428, N8035);
xor XOR2 (N11617, N11612, N1844);
buf BUF1 (N11618, N11606);
nand NAND4 (N11619, N11616, N9417, N3815, N3299);
nor NOR4 (N11620, N11619, N10927, N1031, N9627);
or OR4 (N11621, N11605, N6165, N5462, N8505);
nor NOR2 (N11622, N11614, N11508);
nor NOR4 (N11623, N11618, N10630, N5661, N1878);
not NOT1 (N11624, N11598);
buf BUF1 (N11625, N11620);
nand NAND4 (N11626, N11621, N1656, N6328, N9554);
nand NAND3 (N11627, N11615, N3068, N6975);
nor NOR2 (N11628, N11625, N3436);
nand NAND3 (N11629, N11626, N1228, N4080);
not NOT1 (N11630, N11627);
buf BUF1 (N11631, N11611);
and AND4 (N11632, N11594, N5461, N6161, N8241);
or OR2 (N11633, N11617, N2150);
buf BUF1 (N11634, N11623);
nand NAND2 (N11635, N11624, N4720);
xor XOR2 (N11636, N11622, N4967);
or OR4 (N11637, N11630, N3025, N5808, N4726);
and AND4 (N11638, N11629, N5425, N11384, N4441);
and AND3 (N11639, N11635, N9385, N7391);
and AND3 (N11640, N11637, N4975, N4321);
or OR3 (N11641, N11634, N7729, N9111);
nand NAND2 (N11642, N11639, N15);
not NOT1 (N11643, N11633);
or OR2 (N11644, N11640, N5553);
xor XOR2 (N11645, N11631, N8681);
or OR4 (N11646, N11642, N5970, N1147, N185);
and AND3 (N11647, N11632, N10724, N726);
nand NAND4 (N11648, N11646, N6335, N3117, N3176);
nor NOR4 (N11649, N11648, N8722, N6417, N7642);
not NOT1 (N11650, N11628);
and AND4 (N11651, N11643, N538, N491, N8085);
or OR3 (N11652, N11649, N7786, N9646);
buf BUF1 (N11653, N11647);
nor NOR3 (N11654, N11650, N8741, N9053);
not NOT1 (N11655, N11654);
not NOT1 (N11656, N11655);
nor NOR4 (N11657, N11653, N5782, N9240, N11427);
nand NAND4 (N11658, N11645, N2555, N10874, N450);
and AND4 (N11659, N11657, N6594, N9705, N7757);
nor NOR2 (N11660, N11641, N1317);
not NOT1 (N11661, N11658);
xor XOR2 (N11662, N11644, N3736);
buf BUF1 (N11663, N11638);
nand NAND4 (N11664, N11636, N4117, N4743, N3458);
nand NAND3 (N11665, N11663, N5874, N10487);
or OR3 (N11666, N11652, N3342, N11473);
not NOT1 (N11667, N11656);
xor XOR2 (N11668, N11659, N2139);
not NOT1 (N11669, N11651);
or OR3 (N11670, N11664, N1630, N9121);
buf BUF1 (N11671, N11666);
or OR2 (N11672, N11610, N7813);
buf BUF1 (N11673, N11672);
not NOT1 (N11674, N11660);
buf BUF1 (N11675, N11665);
xor XOR2 (N11676, N11662, N6192);
xor XOR2 (N11677, N11674, N2047);
nor NOR3 (N11678, N11667, N8311, N8418);
buf BUF1 (N11679, N11673);
nand NAND2 (N11680, N11679, N11182);
or OR3 (N11681, N11671, N1677, N11108);
nor NOR4 (N11682, N11670, N3883, N2489, N5653);
xor XOR2 (N11683, N11661, N9718);
or OR4 (N11684, N11669, N5749, N3914, N29);
nand NAND3 (N11685, N11681, N11414, N6769);
buf BUF1 (N11686, N11677);
nor NOR4 (N11687, N11685, N5246, N2290, N6829);
not NOT1 (N11688, N11668);
and AND4 (N11689, N11680, N4995, N7578, N5018);
and AND4 (N11690, N11675, N10268, N3223, N2981);
xor XOR2 (N11691, N11686, N5600);
nor NOR3 (N11692, N11678, N217, N2407);
and AND3 (N11693, N11690, N7434, N9484);
or OR3 (N11694, N11693, N7127, N7171);
or OR2 (N11695, N11684, N3780);
nor NOR2 (N11696, N11676, N3953);
not NOT1 (N11697, N11688);
and AND4 (N11698, N11682, N834, N3729, N7461);
not NOT1 (N11699, N11694);
or OR4 (N11700, N11692, N9861, N112, N2317);
nand NAND2 (N11701, N11683, N4921);
nand NAND4 (N11702, N11698, N4458, N4482, N2476);
and AND4 (N11703, N11691, N7779, N1984, N11139);
nand NAND4 (N11704, N11697, N5297, N4532, N3918);
and AND4 (N11705, N11703, N9446, N7557, N10313);
or OR4 (N11706, N11696, N5860, N2846, N1354);
nand NAND4 (N11707, N11705, N9247, N9130, N6148);
not NOT1 (N11708, N11695);
or OR3 (N11709, N11702, N75, N8921);
and AND4 (N11710, N11707, N8302, N5519, N8355);
nor NOR2 (N11711, N11704, N7069);
not NOT1 (N11712, N11699);
or OR2 (N11713, N11706, N11483);
and AND3 (N11714, N11700, N1087, N2215);
nand NAND3 (N11715, N11709, N7801, N304);
xor XOR2 (N11716, N11708, N4683);
xor XOR2 (N11717, N11687, N8737);
nand NAND3 (N11718, N11714, N9247, N667);
and AND3 (N11719, N11716, N112, N5920);
nand NAND2 (N11720, N11711, N9814);
nand NAND3 (N11721, N11715, N2300, N10218);
nor NOR2 (N11722, N11710, N913);
buf BUF1 (N11723, N11717);
xor XOR2 (N11724, N11720, N8791);
buf BUF1 (N11725, N11719);
buf BUF1 (N11726, N11724);
buf BUF1 (N11727, N11721);
xor XOR2 (N11728, N11713, N10737);
xor XOR2 (N11729, N11728, N4371);
and AND2 (N11730, N11722, N8686);
buf BUF1 (N11731, N11729);
or OR4 (N11732, N11701, N1741, N945, N8372);
nand NAND2 (N11733, N11725, N10111);
nand NAND3 (N11734, N11723, N10650, N9139);
nor NOR3 (N11735, N11731, N8083, N10842);
nand NAND4 (N11736, N11735, N7048, N4899, N6560);
buf BUF1 (N11737, N11736);
xor XOR2 (N11738, N11726, N7452);
xor XOR2 (N11739, N11738, N10389);
nand NAND3 (N11740, N11727, N3533, N11736);
buf BUF1 (N11741, N11734);
buf BUF1 (N11742, N11689);
or OR4 (N11743, N11739, N2816, N3382, N2471);
buf BUF1 (N11744, N11718);
and AND3 (N11745, N11730, N1238, N3799);
nand NAND2 (N11746, N11737, N11121);
and AND4 (N11747, N11740, N9635, N922, N2617);
or OR3 (N11748, N11741, N8387, N9368);
buf BUF1 (N11749, N11744);
and AND2 (N11750, N11742, N3614);
or OR4 (N11751, N11712, N2956, N4611, N10669);
and AND4 (N11752, N11748, N2728, N9340, N6384);
not NOT1 (N11753, N11743);
nand NAND3 (N11754, N11749, N4647, N4132);
or OR3 (N11755, N11732, N11688, N1910);
nand NAND2 (N11756, N11746, N10795);
xor XOR2 (N11757, N11753, N948);
buf BUF1 (N11758, N11752);
not NOT1 (N11759, N11758);
nor NOR2 (N11760, N11747, N107);
nor NOR4 (N11761, N11755, N5899, N9572, N6847);
buf BUF1 (N11762, N11761);
xor XOR2 (N11763, N11733, N8662);
xor XOR2 (N11764, N11756, N1718);
xor XOR2 (N11765, N11759, N9500);
nand NAND4 (N11766, N11745, N10153, N9034, N6706);
xor XOR2 (N11767, N11751, N1500);
and AND2 (N11768, N11762, N260);
nor NOR3 (N11769, N11766, N5597, N2559);
nor NOR2 (N11770, N11769, N10924);
or OR3 (N11771, N11767, N10282, N1913);
nand NAND3 (N11772, N11764, N9656, N8009);
and AND2 (N11773, N11772, N2378);
nand NAND4 (N11774, N11750, N3291, N2472, N11366);
not NOT1 (N11775, N11760);
nand NAND3 (N11776, N11765, N502, N9567);
not NOT1 (N11777, N11773);
not NOT1 (N11778, N11770);
nand NAND4 (N11779, N11776, N5088, N10519, N7262);
or OR3 (N11780, N11754, N7644, N5507);
or OR4 (N11781, N11777, N81, N10055, N10567);
nor NOR3 (N11782, N11768, N10096, N7743);
buf BUF1 (N11783, N11771);
nand NAND3 (N11784, N11774, N5733, N3664);
not NOT1 (N11785, N11780);
and AND2 (N11786, N11782, N4557);
buf BUF1 (N11787, N11783);
and AND4 (N11788, N11779, N9459, N4581, N1009);
xor XOR2 (N11789, N11784, N7044);
xor XOR2 (N11790, N11763, N9707);
nor NOR4 (N11791, N11775, N7278, N4685, N9405);
not NOT1 (N11792, N11757);
buf BUF1 (N11793, N11789);
xor XOR2 (N11794, N11781, N10265);
nor NOR3 (N11795, N11785, N3651, N3491);
xor XOR2 (N11796, N11786, N6564);
and AND2 (N11797, N11794, N3276);
nand NAND4 (N11798, N11778, N11795, N1909, N3493);
nor NOR3 (N11799, N631, N2418, N7235);
and AND2 (N11800, N11788, N9850);
and AND2 (N11801, N11796, N11380);
buf BUF1 (N11802, N11798);
not NOT1 (N11803, N11800);
or OR3 (N11804, N11787, N295, N8372);
buf BUF1 (N11805, N11802);
buf BUF1 (N11806, N11793);
or OR4 (N11807, N11806, N4757, N1, N4427);
nor NOR2 (N11808, N11799, N6069);
not NOT1 (N11809, N11804);
nand NAND4 (N11810, N11807, N1635, N4662, N796);
not NOT1 (N11811, N11803);
nand NAND3 (N11812, N11805, N55, N5775);
nor NOR2 (N11813, N11810, N4134);
not NOT1 (N11814, N11791);
buf BUF1 (N11815, N11792);
xor XOR2 (N11816, N11813, N3764);
nor NOR4 (N11817, N11801, N11791, N7686, N9211);
nand NAND4 (N11818, N11790, N5678, N8481, N2984);
nor NOR3 (N11819, N11816, N3891, N6030);
and AND2 (N11820, N11812, N3176);
xor XOR2 (N11821, N11814, N504);
xor XOR2 (N11822, N11809, N2405);
and AND4 (N11823, N11822, N73, N5582, N4586);
nor NOR2 (N11824, N11819, N76);
and AND4 (N11825, N11797, N8013, N4622, N8147);
nand NAND3 (N11826, N11818, N1595, N2990);
nand NAND4 (N11827, N11823, N519, N1966, N8682);
or OR4 (N11828, N11824, N2451, N9286, N6699);
or OR3 (N11829, N11827, N10481, N5433);
nor NOR3 (N11830, N11811, N4019, N1496);
xor XOR2 (N11831, N11829, N8981);
and AND3 (N11832, N11826, N1175, N4712);
not NOT1 (N11833, N11817);
nand NAND2 (N11834, N11831, N7852);
or OR3 (N11835, N11834, N6594, N306);
and AND4 (N11836, N11820, N1990, N10381, N9005);
not NOT1 (N11837, N11836);
or OR2 (N11838, N11833, N11049);
buf BUF1 (N11839, N11821);
or OR4 (N11840, N11825, N4113, N9060, N11223);
and AND4 (N11841, N11815, N3642, N2193, N1815);
xor XOR2 (N11842, N11837, N3503);
and AND2 (N11843, N11828, N7467);
buf BUF1 (N11844, N11808);
buf BUF1 (N11845, N11842);
nor NOR2 (N11846, N11830, N6792);
nor NOR3 (N11847, N11846, N9091, N4149);
buf BUF1 (N11848, N11841);
nor NOR3 (N11849, N11838, N799, N2128);
nor NOR3 (N11850, N11848, N9668, N6566);
or OR3 (N11851, N11832, N8406, N11752);
xor XOR2 (N11852, N11839, N8638);
nor NOR3 (N11853, N11851, N10615, N1472);
or OR4 (N11854, N11850, N9556, N965, N8226);
not NOT1 (N11855, N11853);
and AND3 (N11856, N11852, N8053, N7236);
not NOT1 (N11857, N11849);
or OR2 (N11858, N11855, N11770);
and AND4 (N11859, N11835, N10593, N9712, N7360);
xor XOR2 (N11860, N11859, N515);
not NOT1 (N11861, N11854);
xor XOR2 (N11862, N11856, N3933);
nand NAND2 (N11863, N11847, N3064);
buf BUF1 (N11864, N11860);
buf BUF1 (N11865, N11864);
nand NAND3 (N11866, N11844, N1309, N9285);
or OR4 (N11867, N11857, N9510, N2866, N5224);
or OR4 (N11868, N11863, N5136, N8166, N3534);
or OR4 (N11869, N11868, N1209, N8694, N833);
xor XOR2 (N11870, N11866, N3873);
or OR2 (N11871, N11870, N7760);
xor XOR2 (N11872, N11867, N7082);
not NOT1 (N11873, N11872);
not NOT1 (N11874, N11845);
nor NOR2 (N11875, N11843, N4222);
nor NOR2 (N11876, N11865, N8119);
and AND2 (N11877, N11873, N8783);
and AND3 (N11878, N11871, N7298, N10629);
nor NOR2 (N11879, N11869, N4901);
and AND3 (N11880, N11878, N5606, N2988);
xor XOR2 (N11881, N11840, N5295);
not NOT1 (N11882, N11862);
not NOT1 (N11883, N11875);
nand NAND2 (N11884, N11876, N9215);
not NOT1 (N11885, N11874);
buf BUF1 (N11886, N11879);
xor XOR2 (N11887, N11882, N1176);
buf BUF1 (N11888, N11885);
xor XOR2 (N11889, N11880, N11819);
xor XOR2 (N11890, N11887, N2834);
buf BUF1 (N11891, N11888);
not NOT1 (N11892, N11886);
not NOT1 (N11893, N11889);
buf BUF1 (N11894, N11881);
xor XOR2 (N11895, N11891, N4958);
buf BUF1 (N11896, N11894);
not NOT1 (N11897, N11858);
and AND2 (N11898, N11893, N2666);
nand NAND4 (N11899, N11883, N7371, N1729, N2342);
nor NOR4 (N11900, N11892, N811, N765, N7743);
nor NOR3 (N11901, N11896, N6041, N3102);
buf BUF1 (N11902, N11900);
nor NOR4 (N11903, N11890, N299, N4819, N11081);
buf BUF1 (N11904, N11902);
xor XOR2 (N11905, N11903, N7804);
xor XOR2 (N11906, N11905, N7620);
buf BUF1 (N11907, N11884);
or OR3 (N11908, N11901, N2835, N10014);
or OR3 (N11909, N11908, N5068, N3560);
and AND2 (N11910, N11907, N10331);
nor NOR2 (N11911, N11861, N8187);
nor NOR4 (N11912, N11877, N3840, N7526, N3940);
not NOT1 (N11913, N11911);
not NOT1 (N11914, N11912);
nor NOR4 (N11915, N11913, N3144, N6673, N4082);
nor NOR4 (N11916, N11899, N4612, N2946, N3440);
or OR2 (N11917, N11898, N485);
xor XOR2 (N11918, N11897, N9093);
or OR4 (N11919, N11917, N3062, N6471, N2273);
xor XOR2 (N11920, N11906, N11113);
nor NOR3 (N11921, N11909, N2582, N10969);
buf BUF1 (N11922, N11919);
buf BUF1 (N11923, N11904);
and AND2 (N11924, N11920, N2788);
or OR4 (N11925, N11915, N7874, N327, N2514);
xor XOR2 (N11926, N11895, N10629);
nor NOR4 (N11927, N11926, N5693, N7254, N9320);
not NOT1 (N11928, N11924);
nor NOR3 (N11929, N11928, N4512, N2511);
or OR3 (N11930, N11927, N10232, N2113);
not NOT1 (N11931, N11914);
not NOT1 (N11932, N11930);
or OR2 (N11933, N11918, N4229);
or OR4 (N11934, N11929, N1677, N2124, N7126);
nand NAND2 (N11935, N11932, N1355);
not NOT1 (N11936, N11931);
xor XOR2 (N11937, N11922, N7765);
or OR2 (N11938, N11936, N1696);
nand NAND2 (N11939, N11934, N4357);
nand NAND4 (N11940, N11925, N5670, N1032, N5306);
and AND2 (N11941, N11939, N6660);
nand NAND3 (N11942, N11935, N5061, N11544);
nand NAND2 (N11943, N11916, N10435);
buf BUF1 (N11944, N11921);
nand NAND3 (N11945, N11943, N11551, N890);
and AND4 (N11946, N11940, N3424, N5010, N6688);
xor XOR2 (N11947, N11923, N2778);
xor XOR2 (N11948, N11937, N1562);
buf BUF1 (N11949, N11910);
not NOT1 (N11950, N11944);
nor NOR4 (N11951, N11938, N8929, N7909, N9280);
nor NOR2 (N11952, N11947, N2583);
buf BUF1 (N11953, N11948);
xor XOR2 (N11954, N11951, N5784);
and AND4 (N11955, N11952, N15, N6316, N815);
and AND2 (N11956, N11955, N3551);
nor NOR2 (N11957, N11953, N7204);
nor NOR2 (N11958, N11957, N1312);
not NOT1 (N11959, N11949);
and AND4 (N11960, N11959, N9987, N11095, N6607);
nor NOR3 (N11961, N11946, N7793, N6057);
buf BUF1 (N11962, N11958);
buf BUF1 (N11963, N11942);
not NOT1 (N11964, N11954);
and AND2 (N11965, N11964, N4191);
xor XOR2 (N11966, N11963, N3783);
nand NAND4 (N11967, N11961, N9631, N6949, N7439);
nor NOR4 (N11968, N11933, N6974, N916, N5725);
buf BUF1 (N11969, N11967);
and AND2 (N11970, N11965, N7465);
and AND4 (N11971, N11969, N5806, N665, N5917);
not NOT1 (N11972, N11941);
xor XOR2 (N11973, N11945, N5567);
nand NAND4 (N11974, N11972, N3721, N7259, N2090);
and AND3 (N11975, N11970, N8027, N8158);
and AND2 (N11976, N11966, N1881);
or OR3 (N11977, N11968, N9498, N10985);
nor NOR3 (N11978, N11975, N2949, N8701);
or OR3 (N11979, N11950, N8328, N11515);
nor NOR2 (N11980, N11971, N228);
nand NAND2 (N11981, N11979, N11978);
nand NAND2 (N11982, N5069, N9357);
or OR3 (N11983, N11974, N7589, N1202);
and AND2 (N11984, N11976, N8288);
or OR2 (N11985, N11960, N1270);
buf BUF1 (N11986, N11980);
buf BUF1 (N11987, N11984);
and AND2 (N11988, N11986, N6306);
or OR4 (N11989, N11982, N8023, N4342, N3941);
xor XOR2 (N11990, N11985, N41);
and AND4 (N11991, N11962, N6081, N8930, N8175);
nand NAND3 (N11992, N11973, N3056, N2771);
xor XOR2 (N11993, N11983, N6639);
nand NAND3 (N11994, N11990, N8607, N582);
xor XOR2 (N11995, N11981, N11142);
not NOT1 (N11996, N11992);
nor NOR3 (N11997, N11977, N10339, N10017);
or OR4 (N11998, N11996, N4558, N3512, N11171);
or OR3 (N11999, N11995, N6361, N10671);
buf BUF1 (N12000, N11991);
and AND2 (N12001, N11987, N4435);
or OR3 (N12002, N11999, N11004, N178);
buf BUF1 (N12003, N11956);
nor NOR2 (N12004, N11997, N2661);
xor XOR2 (N12005, N11998, N4509);
or OR2 (N12006, N11988, N9007);
xor XOR2 (N12007, N12004, N10657);
nor NOR4 (N12008, N11989, N9108, N8931, N7316);
nand NAND3 (N12009, N11993, N4060, N8187);
buf BUF1 (N12010, N12006);
not NOT1 (N12011, N12000);
or OR3 (N12012, N12002, N10529, N5135);
not NOT1 (N12013, N12001);
not NOT1 (N12014, N12010);
nor NOR2 (N12015, N12009, N9862);
nand NAND4 (N12016, N12014, N11023, N2816, N1631);
xor XOR2 (N12017, N12016, N6779);
or OR2 (N12018, N12017, N3527);
not NOT1 (N12019, N12003);
nand NAND4 (N12020, N11994, N593, N3038, N2202);
nor NOR4 (N12021, N12008, N10694, N10150, N11926);
or OR3 (N12022, N12005, N3334, N11089);
xor XOR2 (N12023, N12012, N9558);
buf BUF1 (N12024, N12015);
and AND3 (N12025, N12019, N8166, N11949);
and AND4 (N12026, N12020, N8621, N1188, N11118);
nor NOR3 (N12027, N12021, N10175, N3585);
nor NOR4 (N12028, N12027, N2276, N2603, N1265);
xor XOR2 (N12029, N12011, N11909);
nand NAND3 (N12030, N12023, N3988, N11391);
not NOT1 (N12031, N12013);
not NOT1 (N12032, N12031);
nor NOR4 (N12033, N12028, N7399, N5467, N6693);
not NOT1 (N12034, N12026);
nor NOR4 (N12035, N12030, N8239, N3223, N5129);
nand NAND3 (N12036, N12033, N7101, N7658);
nand NAND4 (N12037, N12032, N9658, N8502, N10582);
or OR3 (N12038, N12025, N10231, N11639);
nor NOR4 (N12039, N12007, N2863, N5578, N657);
or OR4 (N12040, N12022, N6710, N5437, N9928);
nor NOR2 (N12041, N12035, N260);
buf BUF1 (N12042, N12041);
not NOT1 (N12043, N12024);
buf BUF1 (N12044, N12038);
nand NAND2 (N12045, N12043, N5973);
nor NOR4 (N12046, N12040, N3727, N11198, N4557);
and AND3 (N12047, N12044, N11879, N10619);
buf BUF1 (N12048, N12046);
buf BUF1 (N12049, N12037);
not NOT1 (N12050, N12036);
and AND4 (N12051, N12048, N2408, N10871, N5118);
and AND2 (N12052, N12042, N990);
nor NOR4 (N12053, N12018, N7669, N9342, N5380);
nor NOR3 (N12054, N12051, N9217, N8431);
nor NOR3 (N12055, N12053, N4105, N7082);
buf BUF1 (N12056, N12050);
buf BUF1 (N12057, N12052);
nand NAND3 (N12058, N12056, N3004, N3107);
not NOT1 (N12059, N12058);
buf BUF1 (N12060, N12054);
and AND2 (N12061, N12049, N8492);
buf BUF1 (N12062, N12060);
nand NAND4 (N12063, N12057, N3146, N4827, N6452);
xor XOR2 (N12064, N12062, N4093);
and AND3 (N12065, N12039, N3981, N10374);
or OR3 (N12066, N12065, N2562, N6249);
buf BUF1 (N12067, N12064);
nand NAND3 (N12068, N12061, N6311, N11804);
or OR4 (N12069, N12068, N8456, N1349, N9839);
buf BUF1 (N12070, N12047);
xor XOR2 (N12071, N12029, N11997);
nand NAND2 (N12072, N12063, N1701);
nand NAND4 (N12073, N12045, N9309, N9157, N1645);
xor XOR2 (N12074, N12034, N9874);
not NOT1 (N12075, N12073);
buf BUF1 (N12076, N12066);
buf BUF1 (N12077, N12069);
not NOT1 (N12078, N12076);
buf BUF1 (N12079, N12074);
xor XOR2 (N12080, N12075, N10828);
xor XOR2 (N12081, N12059, N8274);
or OR4 (N12082, N12081, N10789, N2853, N9346);
nand NAND3 (N12083, N12067, N3288, N9549);
and AND2 (N12084, N12072, N2067);
nor NOR2 (N12085, N12070, N6881);
nor NOR2 (N12086, N12085, N4698);
not NOT1 (N12087, N12078);
buf BUF1 (N12088, N12084);
buf BUF1 (N12089, N12079);
or OR3 (N12090, N12083, N10531, N11058);
buf BUF1 (N12091, N12071);
and AND3 (N12092, N12089, N979, N8755);
nor NOR3 (N12093, N12091, N6669, N11254);
xor XOR2 (N12094, N12090, N10461);
and AND4 (N12095, N12093, N6985, N8691, N9653);
and AND4 (N12096, N12087, N3143, N2251, N9431);
xor XOR2 (N12097, N12096, N4550);
not NOT1 (N12098, N12092);
nor NOR3 (N12099, N12055, N5102, N10011);
not NOT1 (N12100, N12095);
buf BUF1 (N12101, N12097);
buf BUF1 (N12102, N12098);
and AND4 (N12103, N12086, N809, N10904, N5183);
nand NAND3 (N12104, N12094, N7494, N6323);
nor NOR4 (N12105, N12088, N5740, N747, N10758);
nor NOR4 (N12106, N12104, N4531, N5682, N7202);
nor NOR2 (N12107, N12082, N6992);
nand NAND3 (N12108, N12100, N11550, N1252);
xor XOR2 (N12109, N12106, N4881);
xor XOR2 (N12110, N12109, N10468);
xor XOR2 (N12111, N12102, N9027);
buf BUF1 (N12112, N12105);
nor NOR3 (N12113, N12112, N11621, N9281);
or OR4 (N12114, N12101, N7787, N8900, N11009);
not NOT1 (N12115, N12103);
nor NOR2 (N12116, N12113, N10430);
buf BUF1 (N12117, N12077);
nor NOR2 (N12118, N12107, N9790);
xor XOR2 (N12119, N12117, N2574);
nor NOR3 (N12120, N12118, N3619, N12064);
nor NOR3 (N12121, N12114, N8021, N2345);
nand NAND4 (N12122, N12115, N2072, N11663, N7530);
nand NAND3 (N12123, N12111, N6857, N1838);
and AND4 (N12124, N12122, N11607, N9929, N9834);
and AND2 (N12125, N12108, N6463);
not NOT1 (N12126, N12119);
xor XOR2 (N12127, N12121, N2610);
or OR3 (N12128, N12126, N7279, N4363);
xor XOR2 (N12129, N12080, N5022);
nor NOR2 (N12130, N12099, N8416);
nand NAND3 (N12131, N12128, N8206, N1298);
and AND4 (N12132, N12124, N3234, N4280, N8482);
nor NOR3 (N12133, N12129, N4416, N5987);
buf BUF1 (N12134, N12110);
buf BUF1 (N12135, N12133);
nand NAND2 (N12136, N12134, N8753);
not NOT1 (N12137, N12127);
xor XOR2 (N12138, N12116, N9710);
and AND4 (N12139, N12123, N6046, N11398, N12062);
nor NOR2 (N12140, N12138, N11883);
buf BUF1 (N12141, N12132);
buf BUF1 (N12142, N12135);
nor NOR2 (N12143, N12120, N3860);
or OR3 (N12144, N12140, N5959, N3742);
nand NAND4 (N12145, N12137, N1012, N2135, N4336);
and AND2 (N12146, N12131, N8693);
or OR2 (N12147, N12143, N6244);
xor XOR2 (N12148, N12147, N4440);
or OR3 (N12149, N12146, N10095, N7312);
not NOT1 (N12150, N12125);
xor XOR2 (N12151, N12139, N10390);
or OR2 (N12152, N12142, N247);
not NOT1 (N12153, N12145);
not NOT1 (N12154, N12148);
nand NAND4 (N12155, N12154, N6579, N1303, N10095);
buf BUF1 (N12156, N12130);
not NOT1 (N12157, N12136);
xor XOR2 (N12158, N12157, N962);
xor XOR2 (N12159, N12151, N7355);
nor NOR4 (N12160, N12144, N6722, N12029, N867);
nand NAND2 (N12161, N12159, N1365);
xor XOR2 (N12162, N12160, N11022);
xor XOR2 (N12163, N12152, N4933);
and AND3 (N12164, N12153, N11075, N5930);
nand NAND4 (N12165, N12149, N10974, N3770, N2070);
nor NOR2 (N12166, N12156, N8741);
or OR2 (N12167, N12164, N6597);
nor NOR2 (N12168, N12162, N6216);
buf BUF1 (N12169, N12158);
nand NAND2 (N12170, N12166, N2095);
xor XOR2 (N12171, N12169, N1784);
nor NOR4 (N12172, N12170, N8239, N1011, N527);
not NOT1 (N12173, N12168);
not NOT1 (N12174, N12173);
or OR4 (N12175, N12174, N5597, N4920, N3987);
and AND3 (N12176, N12171, N9628, N9242);
nand NAND3 (N12177, N12167, N6480, N3421);
xor XOR2 (N12178, N12165, N11947);
nor NOR3 (N12179, N12150, N430, N2274);
or OR3 (N12180, N12161, N6947, N4605);
nand NAND3 (N12181, N12155, N1590, N316);
and AND3 (N12182, N12163, N3947, N5211);
and AND3 (N12183, N12179, N4579, N7281);
and AND3 (N12184, N12181, N6213, N11317);
xor XOR2 (N12185, N12180, N1071);
not NOT1 (N12186, N12185);
xor XOR2 (N12187, N12177, N5233);
not NOT1 (N12188, N12178);
buf BUF1 (N12189, N12176);
nor NOR4 (N12190, N12182, N2083, N8231, N9070);
nor NOR2 (N12191, N12172, N9375);
and AND3 (N12192, N12188, N1500, N7145);
and AND2 (N12193, N12187, N2362);
not NOT1 (N12194, N12183);
and AND3 (N12195, N12141, N1324, N7689);
or OR2 (N12196, N12190, N9464);
not NOT1 (N12197, N12196);
or OR3 (N12198, N12194, N5301, N116);
xor XOR2 (N12199, N12189, N7854);
xor XOR2 (N12200, N12191, N4977);
or OR2 (N12201, N12197, N6846);
nand NAND3 (N12202, N12192, N8838, N10211);
buf BUF1 (N12203, N12201);
nand NAND4 (N12204, N12175, N5086, N7685, N1205);
nor NOR3 (N12205, N12199, N10509, N388);
or OR2 (N12206, N12193, N11855);
and AND3 (N12207, N12204, N6509, N2074);
not NOT1 (N12208, N12186);
or OR3 (N12209, N12202, N12079, N10780);
xor XOR2 (N12210, N12198, N10087);
or OR4 (N12211, N12208, N9689, N3308, N9170);
or OR3 (N12212, N12207, N1493, N12189);
buf BUF1 (N12213, N12200);
nand NAND4 (N12214, N12195, N11469, N7116, N11646);
buf BUF1 (N12215, N12205);
and AND3 (N12216, N12215, N1520, N2791);
not NOT1 (N12217, N12184);
and AND4 (N12218, N12203, N4404, N10888, N2233);
nor NOR4 (N12219, N12211, N10877, N3346, N4745);
buf BUF1 (N12220, N12212);
or OR2 (N12221, N12216, N12165);
nand NAND2 (N12222, N12206, N666);
xor XOR2 (N12223, N12218, N10400);
nor NOR2 (N12224, N12223, N11488);
nand NAND4 (N12225, N12210, N9146, N6840, N8324);
xor XOR2 (N12226, N12221, N10115);
nand NAND3 (N12227, N12209, N5541, N1372);
and AND3 (N12228, N12226, N4730, N11913);
nor NOR2 (N12229, N12219, N5463);
or OR4 (N12230, N12222, N9973, N7864, N9188);
nand NAND3 (N12231, N12217, N2296, N7805);
and AND4 (N12232, N12230, N10262, N10689, N9992);
buf BUF1 (N12233, N12214);
nand NAND2 (N12234, N12227, N3320);
xor XOR2 (N12235, N12224, N7023);
not NOT1 (N12236, N12220);
and AND2 (N12237, N12235, N8123);
and AND2 (N12238, N12229, N9353);
not NOT1 (N12239, N12231);
nor NOR3 (N12240, N12236, N3257, N10739);
nor NOR2 (N12241, N12213, N10331);
buf BUF1 (N12242, N12237);
or OR2 (N12243, N12228, N31);
not NOT1 (N12244, N12240);
and AND3 (N12245, N12232, N5199, N1567);
nand NAND4 (N12246, N12234, N8731, N7149, N5698);
buf BUF1 (N12247, N12238);
buf BUF1 (N12248, N12246);
xor XOR2 (N12249, N12225, N8667);
not NOT1 (N12250, N12242);
and AND4 (N12251, N12241, N4829, N9534, N12043);
or OR4 (N12252, N12233, N716, N7680, N5047);
buf BUF1 (N12253, N12244);
and AND2 (N12254, N12252, N3675);
nor NOR4 (N12255, N12254, N11051, N6746, N6020);
or OR4 (N12256, N12243, N7975, N86, N4118);
nand NAND3 (N12257, N12245, N6473, N12222);
and AND2 (N12258, N12239, N9557);
not NOT1 (N12259, N12250);
nand NAND4 (N12260, N12255, N7713, N8884, N1230);
and AND3 (N12261, N12247, N2430, N92);
or OR4 (N12262, N12261, N8592, N8377, N1692);
xor XOR2 (N12263, N12259, N9319);
or OR2 (N12264, N12262, N1891);
nor NOR4 (N12265, N12249, N12055, N1768, N10131);
buf BUF1 (N12266, N12260);
buf BUF1 (N12267, N12248);
nor NOR2 (N12268, N12251, N9916);
buf BUF1 (N12269, N12266);
nor NOR3 (N12270, N12267, N408, N10574);
nand NAND3 (N12271, N12253, N7309, N4228);
not NOT1 (N12272, N12265);
or OR2 (N12273, N12263, N2943);
or OR2 (N12274, N12256, N9598);
not NOT1 (N12275, N12271);
nor NOR3 (N12276, N12269, N53, N11841);
buf BUF1 (N12277, N12268);
or OR3 (N12278, N12276, N3906, N3007);
buf BUF1 (N12279, N12275);
nor NOR2 (N12280, N12279, N2990);
and AND2 (N12281, N12272, N394);
nor NOR3 (N12282, N12264, N12267, N8554);
not NOT1 (N12283, N12274);
and AND3 (N12284, N12258, N133, N1494);
nand NAND3 (N12285, N12282, N75, N4052);
buf BUF1 (N12286, N12277);
or OR3 (N12287, N12257, N9895, N12182);
and AND2 (N12288, N12283, N5842);
buf BUF1 (N12289, N12278);
xor XOR2 (N12290, N12289, N12188);
nor NOR4 (N12291, N12273, N3326, N5982, N7905);
or OR2 (N12292, N12288, N4538);
nand NAND3 (N12293, N12292, N1393, N11075);
nor NOR2 (N12294, N12287, N7291);
and AND2 (N12295, N12291, N5063);
xor XOR2 (N12296, N12285, N8893);
nor NOR2 (N12297, N12295, N6837);
xor XOR2 (N12298, N12284, N9168);
xor XOR2 (N12299, N12286, N11034);
nor NOR2 (N12300, N12298, N4861);
or OR4 (N12301, N12281, N2201, N10966, N3542);
buf BUF1 (N12302, N12290);
nor NOR3 (N12303, N12296, N1000, N11750);
nand NAND4 (N12304, N12293, N5058, N807, N6155);
not NOT1 (N12305, N12303);
xor XOR2 (N12306, N12297, N10145);
not NOT1 (N12307, N12270);
and AND4 (N12308, N12307, N4771, N5448, N5123);
and AND2 (N12309, N12299, N10594);
nand NAND2 (N12310, N12301, N6751);
buf BUF1 (N12311, N12294);
or OR2 (N12312, N12304, N1330);
not NOT1 (N12313, N12300);
and AND3 (N12314, N12313, N7524, N2768);
nand NAND3 (N12315, N12305, N7147, N9748);
nand NAND3 (N12316, N12315, N1348, N1921);
nand NAND3 (N12317, N12310, N4447, N1821);
buf BUF1 (N12318, N12312);
xor XOR2 (N12319, N12311, N10039);
nor NOR3 (N12320, N12308, N7907, N11183);
xor XOR2 (N12321, N12306, N2518);
or OR2 (N12322, N12321, N7019);
or OR2 (N12323, N12317, N2351);
nand NAND2 (N12324, N12302, N5078);
not NOT1 (N12325, N12319);
and AND3 (N12326, N12323, N203, N11425);
not NOT1 (N12327, N12309);
or OR3 (N12328, N12316, N2650, N5207);
not NOT1 (N12329, N12328);
or OR3 (N12330, N12322, N709, N9690);
and AND3 (N12331, N12325, N5957, N10489);
nor NOR2 (N12332, N12327, N3261);
xor XOR2 (N12333, N12332, N974);
and AND4 (N12334, N12329, N430, N118, N9033);
nor NOR3 (N12335, N12334, N5157, N4628);
not NOT1 (N12336, N12331);
nand NAND2 (N12337, N12330, N10747);
or OR2 (N12338, N12333, N10102);
nand NAND4 (N12339, N12335, N1706, N5564, N1654);
nor NOR2 (N12340, N12326, N743);
nor NOR4 (N12341, N12324, N6673, N1968, N10144);
nor NOR2 (N12342, N12314, N7706);
and AND2 (N12343, N12341, N10314);
nand NAND2 (N12344, N12336, N10836);
nor NOR4 (N12345, N12337, N5146, N1209, N10170);
buf BUF1 (N12346, N12342);
and AND4 (N12347, N12339, N7375, N2590, N10141);
xor XOR2 (N12348, N12280, N6944);
not NOT1 (N12349, N12318);
xor XOR2 (N12350, N12344, N9479);
nor NOR4 (N12351, N12350, N799, N3799, N5991);
not NOT1 (N12352, N12340);
nand NAND4 (N12353, N12349, N6692, N6664, N6294);
and AND3 (N12354, N12345, N3085, N7962);
and AND4 (N12355, N12348, N3303, N4755, N4385);
not NOT1 (N12356, N12354);
buf BUF1 (N12357, N12320);
and AND4 (N12358, N12351, N11493, N12222, N756);
or OR3 (N12359, N12356, N11081, N8276);
xor XOR2 (N12360, N12343, N11249);
nand NAND3 (N12361, N12360, N4129, N8309);
and AND2 (N12362, N12338, N364);
or OR4 (N12363, N12362, N4038, N7824, N11074);
buf BUF1 (N12364, N12347);
buf BUF1 (N12365, N12361);
nand NAND4 (N12366, N12364, N1375, N9190, N1084);
nand NAND4 (N12367, N12355, N9695, N7304, N4781);
nand NAND2 (N12368, N12367, N9259);
buf BUF1 (N12369, N12359);
and AND4 (N12370, N12363, N3227, N9588, N3255);
xor XOR2 (N12371, N12357, N10085);
nor NOR3 (N12372, N12366, N6760, N9935);
nand NAND2 (N12373, N12365, N81);
or OR2 (N12374, N12368, N3810);
buf BUF1 (N12375, N12346);
or OR3 (N12376, N12374, N4503, N5704);
nor NOR3 (N12377, N12372, N5648, N4274);
not NOT1 (N12378, N12353);
or OR3 (N12379, N12358, N2371, N5530);
or OR3 (N12380, N12379, N6852, N7795);
and AND3 (N12381, N12378, N8638, N4661);
nand NAND2 (N12382, N12377, N4985);
nor NOR2 (N12383, N12375, N4293);
and AND4 (N12384, N12381, N11456, N5817, N4385);
nor NOR3 (N12385, N12382, N8344, N10726);
or OR2 (N12386, N12370, N11021);
and AND2 (N12387, N12376, N5392);
nor NOR4 (N12388, N12386, N8455, N9561, N2536);
nor NOR4 (N12389, N12388, N9762, N2395, N964);
or OR3 (N12390, N12369, N3437, N5581);
xor XOR2 (N12391, N12389, N7448);
or OR3 (N12392, N12371, N8809, N11684);
nand NAND3 (N12393, N12391, N8686, N2042);
nand NAND2 (N12394, N12393, N5978);
nand NAND2 (N12395, N12392, N3041);
nand NAND3 (N12396, N12383, N11927, N8958);
nand NAND4 (N12397, N12373, N5820, N6318, N7243);
or OR2 (N12398, N12395, N2676);
xor XOR2 (N12399, N12397, N3408);
or OR4 (N12400, N12385, N11346, N5678, N1545);
not NOT1 (N12401, N12390);
not NOT1 (N12402, N12398);
xor XOR2 (N12403, N12394, N1414);
or OR4 (N12404, N12384, N3146, N7498, N9151);
nand NAND4 (N12405, N12380, N43, N6459, N5510);
nand NAND3 (N12406, N12399, N4839, N6357);
nand NAND3 (N12407, N12402, N5373, N8924);
and AND2 (N12408, N12401, N36);
and AND4 (N12409, N12406, N7180, N4401, N8803);
buf BUF1 (N12410, N12408);
not NOT1 (N12411, N12409);
nor NOR4 (N12412, N12403, N5175, N10154, N3291);
not NOT1 (N12413, N12404);
nor NOR2 (N12414, N12410, N6608);
nor NOR2 (N12415, N12352, N10727);
not NOT1 (N12416, N12396);
nor NOR3 (N12417, N12411, N2835, N7902);
not NOT1 (N12418, N12414);
buf BUF1 (N12419, N12412);
or OR2 (N12420, N12417, N6474);
xor XOR2 (N12421, N12407, N7923);
buf BUF1 (N12422, N12387);
nor NOR2 (N12423, N12422, N6075);
nand NAND4 (N12424, N12421, N5461, N10863, N3307);
xor XOR2 (N12425, N12423, N4241);
nand NAND3 (N12426, N12420, N1363, N5637);
buf BUF1 (N12427, N12419);
xor XOR2 (N12428, N12427, N7686);
nand NAND4 (N12429, N12426, N11400, N947, N11553);
nor NOR2 (N12430, N12416, N11549);
nand NAND2 (N12431, N12428, N5384);
nor NOR2 (N12432, N12418, N6842);
nor NOR4 (N12433, N12432, N2663, N11080, N4388);
buf BUF1 (N12434, N12413);
nor NOR2 (N12435, N12431, N450);
not NOT1 (N12436, N12429);
not NOT1 (N12437, N12425);
xor XOR2 (N12438, N12434, N6155);
not NOT1 (N12439, N12424);
or OR3 (N12440, N12437, N8592, N2969);
not NOT1 (N12441, N12400);
and AND4 (N12442, N12430, N2203, N1096, N4452);
or OR2 (N12443, N12433, N1501);
and AND2 (N12444, N12439, N1911);
not NOT1 (N12445, N12436);
nand NAND4 (N12446, N12445, N1040, N11196, N3805);
not NOT1 (N12447, N12446);
and AND2 (N12448, N12415, N8371);
xor XOR2 (N12449, N12447, N1315);
nor NOR4 (N12450, N12449, N6201, N1222, N6090);
xor XOR2 (N12451, N12440, N9104);
nor NOR4 (N12452, N12442, N1012, N5074, N752);
nor NOR3 (N12453, N12441, N1863, N39);
nor NOR4 (N12454, N12450, N907, N7128, N9168);
nor NOR3 (N12455, N12443, N7, N4867);
and AND3 (N12456, N12438, N8956, N3760);
and AND3 (N12457, N12448, N6038, N2142);
nor NOR2 (N12458, N12444, N1066);
buf BUF1 (N12459, N12456);
not NOT1 (N12460, N12435);
or OR3 (N12461, N12458, N1215, N3851);
and AND3 (N12462, N12453, N12454, N37);
buf BUF1 (N12463, N9992);
not NOT1 (N12464, N12457);
and AND2 (N12465, N12462, N1240);
buf BUF1 (N12466, N12463);
and AND2 (N12467, N12466, N5941);
xor XOR2 (N12468, N12464, N6409);
nor NOR3 (N12469, N12468, N6340, N7900);
nand NAND3 (N12470, N12455, N9317, N6187);
or OR2 (N12471, N12470, N505);
or OR4 (N12472, N12452, N5273, N4207, N10655);
not NOT1 (N12473, N12465);
and AND4 (N12474, N12473, N4458, N3008, N5491);
nor NOR4 (N12475, N12405, N6022, N4216, N7005);
or OR3 (N12476, N12475, N7010, N5581);
xor XOR2 (N12477, N12474, N9881);
xor XOR2 (N12478, N12476, N1446);
buf BUF1 (N12479, N12478);
nand NAND3 (N12480, N12460, N12417, N10072);
not NOT1 (N12481, N12451);
buf BUF1 (N12482, N12477);
xor XOR2 (N12483, N12461, N7382);
buf BUF1 (N12484, N12467);
xor XOR2 (N12485, N12469, N4434);
nor NOR2 (N12486, N12484, N4998);
buf BUF1 (N12487, N12479);
buf BUF1 (N12488, N12486);
not NOT1 (N12489, N12487);
buf BUF1 (N12490, N12485);
buf BUF1 (N12491, N12483);
buf BUF1 (N12492, N12472);
xor XOR2 (N12493, N12490, N6877);
xor XOR2 (N12494, N12488, N11748);
buf BUF1 (N12495, N12480);
not NOT1 (N12496, N12492);
nand NAND4 (N12497, N12471, N1446, N2425, N3981);
not NOT1 (N12498, N12489);
not NOT1 (N12499, N12491);
buf BUF1 (N12500, N12482);
xor XOR2 (N12501, N12493, N6032);
nor NOR2 (N12502, N12498, N10411);
nor NOR4 (N12503, N12494, N250, N6812, N10389);
nand NAND2 (N12504, N12500, N7890);
and AND3 (N12505, N12481, N10185, N2225);
nand NAND3 (N12506, N12501, N5117, N7507);
nor NOR2 (N12507, N12502, N7574);
not NOT1 (N12508, N12496);
not NOT1 (N12509, N12503);
buf BUF1 (N12510, N12509);
not NOT1 (N12511, N12495);
nand NAND4 (N12512, N12505, N5464, N9687, N8342);
nor NOR2 (N12513, N12507, N4615);
buf BUF1 (N12514, N12508);
or OR4 (N12515, N12499, N4219, N1910, N9401);
or OR4 (N12516, N12504, N11314, N2473, N9991);
buf BUF1 (N12517, N12514);
and AND3 (N12518, N12497, N8562, N4110);
or OR4 (N12519, N12517, N10809, N2553, N6678);
or OR3 (N12520, N12518, N2001, N11569);
not NOT1 (N12521, N12510);
and AND4 (N12522, N12512, N12089, N4304, N8263);
xor XOR2 (N12523, N12459, N10650);
nand NAND4 (N12524, N12521, N12006, N11803, N5496);
not NOT1 (N12525, N12516);
not NOT1 (N12526, N12513);
or OR2 (N12527, N12520, N4528);
not NOT1 (N12528, N12522);
nand NAND3 (N12529, N12524, N12483, N7993);
or OR3 (N12530, N12511, N8068, N3529);
buf BUF1 (N12531, N12526);
nand NAND4 (N12532, N12523, N3374, N5885, N8121);
not NOT1 (N12533, N12525);
xor XOR2 (N12534, N12533, N3275);
nor NOR4 (N12535, N12529, N8220, N1881, N9610);
xor XOR2 (N12536, N12519, N4397);
xor XOR2 (N12537, N12536, N7526);
not NOT1 (N12538, N12535);
and AND4 (N12539, N12532, N340, N6053, N3318);
buf BUF1 (N12540, N12538);
or OR2 (N12541, N12528, N1755);
nor NOR2 (N12542, N12540, N8939);
or OR3 (N12543, N12541, N1227, N5927);
nand NAND3 (N12544, N12515, N11077, N11378);
not NOT1 (N12545, N12537);
nor NOR4 (N12546, N12534, N11632, N116, N4650);
or OR2 (N12547, N12506, N942);
and AND4 (N12548, N12539, N101, N5751, N8562);
nand NAND3 (N12549, N12527, N3400, N7597);
buf BUF1 (N12550, N12549);
xor XOR2 (N12551, N12548, N5135);
xor XOR2 (N12552, N12550, N4839);
xor XOR2 (N12553, N12552, N5447);
and AND3 (N12554, N12547, N3874, N335);
not NOT1 (N12555, N12531);
not NOT1 (N12556, N12543);
or OR2 (N12557, N12546, N12310);
or OR4 (N12558, N12555, N9803, N4312, N3145);
nor NOR3 (N12559, N12542, N5745, N9830);
buf BUF1 (N12560, N12559);
nor NOR3 (N12561, N12558, N8655, N11388);
buf BUF1 (N12562, N12560);
nand NAND3 (N12563, N12551, N307, N359);
nor NOR3 (N12564, N12530, N3625, N7445);
or OR3 (N12565, N12554, N17, N9799);
xor XOR2 (N12566, N12565, N559);
nand NAND2 (N12567, N12557, N6802);
xor XOR2 (N12568, N12544, N2608);
buf BUF1 (N12569, N12564);
buf BUF1 (N12570, N12561);
buf BUF1 (N12571, N12567);
buf BUF1 (N12572, N12553);
and AND2 (N12573, N12562, N5950);
or OR4 (N12574, N12545, N11800, N3717, N6220);
buf BUF1 (N12575, N12570);
xor XOR2 (N12576, N12572, N1112);
buf BUF1 (N12577, N12573);
and AND4 (N12578, N12575, N10193, N1438, N9037);
or OR4 (N12579, N12574, N1469, N11076, N8984);
or OR4 (N12580, N12568, N10016, N11799, N7145);
not NOT1 (N12581, N12569);
nand NAND4 (N12582, N12579, N4847, N2520, N8955);
nor NOR3 (N12583, N12578, N6867, N3800);
nand NAND3 (N12584, N12563, N11931, N4494);
and AND3 (N12585, N12556, N8049, N5377);
buf BUF1 (N12586, N12580);
not NOT1 (N12587, N12584);
and AND3 (N12588, N12587, N12034, N970);
nand NAND3 (N12589, N12582, N4898, N8694);
nor NOR2 (N12590, N12581, N9355);
nor NOR4 (N12591, N12566, N5866, N9010, N12107);
and AND2 (N12592, N12583, N2951);
not NOT1 (N12593, N12585);
or OR3 (N12594, N12588, N5993, N6641);
buf BUF1 (N12595, N12577);
nor NOR4 (N12596, N12595, N4374, N3105, N8112);
buf BUF1 (N12597, N12590);
buf BUF1 (N12598, N12586);
xor XOR2 (N12599, N12571, N4878);
nand NAND2 (N12600, N12597, N8363);
and AND4 (N12601, N12576, N1585, N10725, N9414);
or OR2 (N12602, N12600, N5378);
buf BUF1 (N12603, N12592);
nor NOR3 (N12604, N12603, N4717, N7140);
nand NAND3 (N12605, N12604, N7794, N6137);
buf BUF1 (N12606, N12601);
nand NAND4 (N12607, N12602, N2612, N1881, N11274);
nor NOR2 (N12608, N12598, N8246);
buf BUF1 (N12609, N12593);
nor NOR4 (N12610, N12608, N4562, N3883, N6472);
or OR2 (N12611, N12589, N9134);
buf BUF1 (N12612, N12611);
xor XOR2 (N12613, N12599, N7244);
xor XOR2 (N12614, N12607, N1441);
nor NOR3 (N12615, N12612, N11076, N11747);
not NOT1 (N12616, N12614);
nor NOR4 (N12617, N12605, N2181, N6387, N11462);
xor XOR2 (N12618, N12596, N10518);
xor XOR2 (N12619, N12594, N8620);
not NOT1 (N12620, N12609);
xor XOR2 (N12621, N12617, N9504);
not NOT1 (N12622, N12606);
nand NAND4 (N12623, N12622, N51, N8646, N8743);
buf BUF1 (N12624, N12616);
nor NOR4 (N12625, N12618, N9887, N3582, N5921);
xor XOR2 (N12626, N12623, N387);
not NOT1 (N12627, N12625);
nand NAND3 (N12628, N12626, N6869, N5479);
nand NAND3 (N12629, N12627, N1665, N6658);
or OR3 (N12630, N12610, N6876, N5411);
nor NOR2 (N12631, N12613, N10913);
buf BUF1 (N12632, N12619);
buf BUF1 (N12633, N12629);
buf BUF1 (N12634, N12620);
and AND3 (N12635, N12630, N9233, N6521);
or OR4 (N12636, N12615, N7346, N2618, N8201);
nor NOR4 (N12637, N12635, N3401, N10699, N9720);
not NOT1 (N12638, N12634);
nand NAND3 (N12639, N12591, N907, N4535);
or OR4 (N12640, N12633, N5056, N4903, N3439);
nor NOR4 (N12641, N12632, N2107, N5713, N3159);
or OR4 (N12642, N12640, N3852, N2047, N9143);
nor NOR4 (N12643, N12638, N11849, N12598, N10774);
buf BUF1 (N12644, N12637);
nand NAND2 (N12645, N12644, N417);
not NOT1 (N12646, N12636);
nor NOR2 (N12647, N12641, N2714);
or OR3 (N12648, N12624, N7962, N6924);
buf BUF1 (N12649, N12621);
or OR4 (N12650, N12646, N1623, N10972, N5177);
xor XOR2 (N12651, N12648, N432);
nor NOR2 (N12652, N12647, N9511);
buf BUF1 (N12653, N12651);
or OR4 (N12654, N12645, N5082, N11829, N5218);
nor NOR4 (N12655, N12654, N2936, N12161, N9654);
buf BUF1 (N12656, N12653);
or OR2 (N12657, N12639, N551);
buf BUF1 (N12658, N12631);
or OR4 (N12659, N12652, N9089, N12037, N10033);
not NOT1 (N12660, N12643);
nor NOR4 (N12661, N12642, N2919, N12047, N1867);
and AND2 (N12662, N12656, N2280);
or OR2 (N12663, N12628, N9259);
nor NOR4 (N12664, N12661, N10357, N4600, N3295);
or OR2 (N12665, N12664, N12569);
nand NAND4 (N12666, N12660, N905, N11847, N12284);
and AND3 (N12667, N12655, N6667, N10976);
and AND2 (N12668, N12665, N3199);
buf BUF1 (N12669, N12650);
nor NOR3 (N12670, N12659, N2094, N11325);
and AND3 (N12671, N12662, N11248, N3423);
buf BUF1 (N12672, N12671);
nor NOR2 (N12673, N12672, N4951);
or OR3 (N12674, N12669, N8932, N463);
buf BUF1 (N12675, N12674);
nor NOR4 (N12676, N12657, N4941, N9031, N3070);
buf BUF1 (N12677, N12667);
xor XOR2 (N12678, N12673, N2547);
nor NOR2 (N12679, N12670, N11961);
buf BUF1 (N12680, N12658);
and AND3 (N12681, N12679, N5607, N7534);
or OR2 (N12682, N12678, N8846);
not NOT1 (N12683, N12676);
or OR4 (N12684, N12681, N3172, N9910, N6886);
not NOT1 (N12685, N12680);
or OR2 (N12686, N12649, N5925);
not NOT1 (N12687, N12685);
buf BUF1 (N12688, N12682);
xor XOR2 (N12689, N12663, N11392);
xor XOR2 (N12690, N12677, N4899);
or OR2 (N12691, N12683, N9600);
nand NAND2 (N12692, N12687, N11746);
and AND2 (N12693, N12690, N9133);
nor NOR4 (N12694, N12688, N6019, N352, N2003);
xor XOR2 (N12695, N12686, N10434);
or OR3 (N12696, N12668, N11392, N2603);
nand NAND4 (N12697, N12689, N4776, N11745, N7195);
xor XOR2 (N12698, N12666, N12475);
not NOT1 (N12699, N12684);
and AND2 (N12700, N12675, N7007);
not NOT1 (N12701, N12694);
nand NAND3 (N12702, N12698, N11537, N10057);
xor XOR2 (N12703, N12702, N2919);
or OR2 (N12704, N12700, N5712);
xor XOR2 (N12705, N12691, N5132);
nor NOR4 (N12706, N12703, N7213, N3476, N3309);
nand NAND3 (N12707, N12705, N7868, N11400);
or OR4 (N12708, N12692, N9278, N8034, N11165);
nor NOR3 (N12709, N12699, N11777, N8647);
xor XOR2 (N12710, N12704, N3405);
or OR2 (N12711, N12709, N1410);
buf BUF1 (N12712, N12693);
buf BUF1 (N12713, N12710);
buf BUF1 (N12714, N12701);
nor NOR2 (N12715, N12707, N7134);
xor XOR2 (N12716, N12695, N1900);
nand NAND2 (N12717, N12697, N12673);
not NOT1 (N12718, N12713);
xor XOR2 (N12719, N12696, N562);
xor XOR2 (N12720, N12706, N10979);
or OR3 (N12721, N12712, N5785, N4910);
or OR4 (N12722, N12719, N7434, N11612, N8672);
xor XOR2 (N12723, N12720, N9279);
not NOT1 (N12724, N12715);
and AND4 (N12725, N12718, N9063, N4785, N10636);
xor XOR2 (N12726, N12711, N6393);
not NOT1 (N12727, N12721);
nor NOR4 (N12728, N12727, N12503, N8076, N2967);
nand NAND2 (N12729, N12723, N4411);
buf BUF1 (N12730, N12708);
or OR2 (N12731, N12716, N10542);
not NOT1 (N12732, N12725);
nand NAND3 (N12733, N12726, N4523, N9991);
or OR4 (N12734, N12730, N11178, N8213, N10983);
not NOT1 (N12735, N12728);
and AND2 (N12736, N12732, N10988);
buf BUF1 (N12737, N12722);
or OR4 (N12738, N12714, N11584, N94, N5914);
nand NAND3 (N12739, N12724, N9269, N2679);
not NOT1 (N12740, N12733);
nor NOR2 (N12741, N12737, N4795);
nand NAND4 (N12742, N12731, N7318, N312, N437);
and AND3 (N12743, N12739, N10726, N6981);
nor NOR2 (N12744, N12717, N3295);
and AND3 (N12745, N12741, N1605, N5717);
or OR3 (N12746, N12744, N9938, N3064);
not NOT1 (N12747, N12745);
nand NAND4 (N12748, N12746, N12261, N10217, N9503);
or OR2 (N12749, N12743, N2332);
not NOT1 (N12750, N12747);
xor XOR2 (N12751, N12750, N9507);
xor XOR2 (N12752, N12729, N9899);
xor XOR2 (N12753, N12736, N1964);
or OR4 (N12754, N12735, N12693, N3337, N10422);
or OR3 (N12755, N12751, N10654, N10857);
nor NOR4 (N12756, N12748, N5923, N5297, N6477);
and AND4 (N12757, N12755, N420, N10657, N3174);
nor NOR3 (N12758, N12738, N9768, N1568);
nor NOR4 (N12759, N12753, N7993, N2894, N3383);
and AND4 (N12760, N12742, N8096, N3720, N4838);
and AND4 (N12761, N12752, N4831, N1760, N105);
or OR2 (N12762, N12760, N11145);
or OR3 (N12763, N12758, N2515, N1027);
buf BUF1 (N12764, N12756);
and AND4 (N12765, N12763, N1338, N9527, N3921);
or OR3 (N12766, N12764, N12193, N7959);
nand NAND4 (N12767, N12749, N2282, N12105, N2527);
or OR4 (N12768, N12762, N9977, N4098, N8334);
not NOT1 (N12769, N12757);
buf BUF1 (N12770, N12761);
nor NOR4 (N12771, N12734, N12060, N1697, N12076);
buf BUF1 (N12772, N12759);
nor NOR4 (N12773, N12771, N1052, N287, N11262);
buf BUF1 (N12774, N12754);
and AND3 (N12775, N12774, N10313, N4741);
nor NOR2 (N12776, N12770, N3513);
nand NAND4 (N12777, N12766, N6261, N1530, N8968);
or OR4 (N12778, N12777, N11697, N609, N2836);
buf BUF1 (N12779, N12778);
buf BUF1 (N12780, N12740);
or OR4 (N12781, N12773, N7056, N2770, N682);
not NOT1 (N12782, N12765);
not NOT1 (N12783, N12772);
nand NAND3 (N12784, N12768, N10282, N3831);
nor NOR3 (N12785, N12783, N9798, N5743);
not NOT1 (N12786, N12781);
not NOT1 (N12787, N12779);
nor NOR4 (N12788, N12782, N9621, N6400, N5746);
nand NAND2 (N12789, N12776, N10095);
and AND2 (N12790, N12788, N6482);
buf BUF1 (N12791, N12786);
not NOT1 (N12792, N12767);
and AND2 (N12793, N12785, N11859);
nor NOR2 (N12794, N12789, N8158);
nor NOR3 (N12795, N12792, N4853, N7777);
not NOT1 (N12796, N12780);
buf BUF1 (N12797, N12784);
and AND4 (N12798, N12795, N3629, N6188, N4105);
nand NAND3 (N12799, N12796, N6454, N4214);
and AND3 (N12800, N12797, N8358, N9185);
xor XOR2 (N12801, N12787, N2443);
buf BUF1 (N12802, N12793);
buf BUF1 (N12803, N12798);
not NOT1 (N12804, N12802);
and AND4 (N12805, N12803, N7358, N4648, N1807);
or OR4 (N12806, N12805, N1088, N9086, N10784);
or OR2 (N12807, N12800, N4962);
xor XOR2 (N12808, N12801, N2220);
or OR2 (N12809, N12806, N10428);
xor XOR2 (N12810, N12769, N11421);
xor XOR2 (N12811, N12799, N6294);
not NOT1 (N12812, N12809);
or OR4 (N12813, N12808, N145, N5716, N1278);
and AND2 (N12814, N12812, N3665);
and AND2 (N12815, N12807, N11595);
or OR4 (N12816, N12813, N5849, N8890, N10205);
nand NAND4 (N12817, N12814, N1141, N1863, N11395);
nor NOR2 (N12818, N12794, N1226);
or OR2 (N12819, N12790, N7096);
nor NOR3 (N12820, N12816, N1192, N10136);
nor NOR4 (N12821, N12810, N6224, N1039, N8848);
nor NOR4 (N12822, N12804, N4196, N5666, N3991);
buf BUF1 (N12823, N12775);
nor NOR4 (N12824, N12823, N6917, N8814, N3975);
and AND3 (N12825, N12815, N897, N12605);
or OR3 (N12826, N12817, N9576, N4914);
or OR4 (N12827, N12811, N11357, N386, N6109);
buf BUF1 (N12828, N12822);
or OR4 (N12829, N12824, N4425, N4545, N3724);
and AND3 (N12830, N12828, N9764, N11417);
xor XOR2 (N12831, N12827, N254);
or OR3 (N12832, N12820, N2799, N5086);
nor NOR2 (N12833, N12831, N10101);
nor NOR4 (N12834, N12819, N3030, N9190, N2077);
or OR3 (N12835, N12818, N6874, N3399);
xor XOR2 (N12836, N12791, N6610);
nor NOR2 (N12837, N12830, N10532);
buf BUF1 (N12838, N12837);
nand NAND2 (N12839, N12821, N9576);
xor XOR2 (N12840, N12839, N10397);
xor XOR2 (N12841, N12829, N6534);
buf BUF1 (N12842, N12834);
nor NOR2 (N12843, N12838, N5149);
nand NAND4 (N12844, N12842, N2686, N12411, N12478);
buf BUF1 (N12845, N12840);
nor NOR4 (N12846, N12833, N7385, N4332, N1460);
buf BUF1 (N12847, N12826);
buf BUF1 (N12848, N12845);
or OR3 (N12849, N12846, N1324, N9031);
nor NOR2 (N12850, N12825, N10258);
nand NAND4 (N12851, N12843, N12546, N9420, N12087);
and AND3 (N12852, N12849, N503, N10267);
and AND2 (N12853, N12844, N5665);
nor NOR2 (N12854, N12847, N7633);
not NOT1 (N12855, N12852);
nand NAND4 (N12856, N12836, N7811, N11445, N11181);
buf BUF1 (N12857, N12854);
or OR4 (N12858, N12853, N7380, N1712, N447);
xor XOR2 (N12859, N12841, N10936);
buf BUF1 (N12860, N12856);
or OR2 (N12861, N12848, N3277);
nand NAND4 (N12862, N12857, N10670, N11063, N5926);
and AND2 (N12863, N12858, N4852);
or OR2 (N12864, N12851, N4091);
nor NOR4 (N12865, N12862, N3625, N9531, N2317);
or OR3 (N12866, N12864, N3778, N7909);
nand NAND3 (N12867, N12865, N2618, N3665);
nand NAND2 (N12868, N12860, N2262);
not NOT1 (N12869, N12863);
nor NOR4 (N12870, N12832, N228, N1620, N2550);
nand NAND4 (N12871, N12866, N7573, N9237, N8480);
and AND2 (N12872, N12835, N5465);
xor XOR2 (N12873, N12859, N1086);
xor XOR2 (N12874, N12855, N10176);
not NOT1 (N12875, N12873);
or OR2 (N12876, N12871, N12135);
and AND4 (N12877, N12870, N11856, N3056, N4826);
not NOT1 (N12878, N12875);
not NOT1 (N12879, N12878);
not NOT1 (N12880, N12867);
nand NAND3 (N12881, N12874, N1751, N8435);
nor NOR3 (N12882, N12877, N11339, N611);
xor XOR2 (N12883, N12876, N6499);
nand NAND4 (N12884, N12882, N4180, N5636, N5040);
nor NOR4 (N12885, N12881, N700, N11413, N5544);
and AND4 (N12886, N12883, N2527, N1879, N4445);
not NOT1 (N12887, N12884);
not NOT1 (N12888, N12887);
xor XOR2 (N12889, N12861, N9361);
not NOT1 (N12890, N12886);
and AND4 (N12891, N12869, N8855, N5346, N10618);
not NOT1 (N12892, N12868);
nand NAND3 (N12893, N12890, N12468, N3794);
or OR4 (N12894, N12850, N11834, N7595, N7339);
buf BUF1 (N12895, N12889);
nand NAND3 (N12896, N12880, N7759, N2336);
and AND3 (N12897, N12891, N12323, N12105);
nand NAND4 (N12898, N12879, N2262, N11686, N6782);
xor XOR2 (N12899, N12894, N2682);
and AND2 (N12900, N12872, N5714);
and AND3 (N12901, N12900, N2224, N12837);
and AND2 (N12902, N12885, N5856);
not NOT1 (N12903, N12896);
not NOT1 (N12904, N12893);
and AND2 (N12905, N12899, N3495);
buf BUF1 (N12906, N12892);
and AND3 (N12907, N12897, N3564, N9785);
or OR3 (N12908, N12901, N343, N11764);
or OR3 (N12909, N12895, N3655, N4402);
xor XOR2 (N12910, N12904, N154);
and AND2 (N12911, N12909, N9355);
and AND4 (N12912, N12898, N12879, N628, N3663);
not NOT1 (N12913, N12903);
buf BUF1 (N12914, N12902);
nor NOR4 (N12915, N12908, N12666, N4269, N7802);
or OR2 (N12916, N12912, N11688);
or OR2 (N12917, N12905, N662);
xor XOR2 (N12918, N12907, N8786);
xor XOR2 (N12919, N12918, N6113);
xor XOR2 (N12920, N12906, N4660);
not NOT1 (N12921, N12910);
xor XOR2 (N12922, N12913, N7334);
nor NOR2 (N12923, N12921, N4148);
and AND2 (N12924, N12923, N3531);
and AND2 (N12925, N12922, N10420);
and AND3 (N12926, N12920, N4250, N2849);
nand NAND3 (N12927, N12919, N3995, N3294);
not NOT1 (N12928, N12888);
or OR4 (N12929, N12926, N7024, N5849, N7287);
xor XOR2 (N12930, N12911, N3708);
not NOT1 (N12931, N12928);
buf BUF1 (N12932, N12931);
and AND2 (N12933, N12917, N4777);
nor NOR3 (N12934, N12925, N1066, N3390);
nand NAND4 (N12935, N12932, N9003, N4695, N1430);
nand NAND3 (N12936, N12924, N10372, N3141);
not NOT1 (N12937, N12934);
or OR2 (N12938, N12930, N5324);
and AND2 (N12939, N12914, N6755);
nor NOR2 (N12940, N12927, N11938);
nand NAND2 (N12941, N12937, N2538);
buf BUF1 (N12942, N12935);
and AND4 (N12943, N12929, N2292, N816, N8675);
nor NOR3 (N12944, N12936, N5869, N10392);
not NOT1 (N12945, N12944);
buf BUF1 (N12946, N12940);
nor NOR2 (N12947, N12941, N7038);
or OR3 (N12948, N12938, N186, N2547);
not NOT1 (N12949, N12916);
buf BUF1 (N12950, N12949);
not NOT1 (N12951, N12943);
buf BUF1 (N12952, N12945);
buf BUF1 (N12953, N12951);
or OR2 (N12954, N12946, N10086);
and AND2 (N12955, N12933, N12861);
nor NOR2 (N12956, N12915, N5710);
not NOT1 (N12957, N12939);
and AND3 (N12958, N12956, N2458, N12194);
xor XOR2 (N12959, N12952, N5739);
nand NAND2 (N12960, N12958, N9849);
nand NAND2 (N12961, N12948, N1781);
or OR2 (N12962, N12942, N1459);
nand NAND4 (N12963, N12955, N9415, N2438, N10981);
nor NOR4 (N12964, N12953, N4874, N2288, N4980);
not NOT1 (N12965, N12961);
or OR2 (N12966, N12957, N6724);
buf BUF1 (N12967, N12947);
or OR3 (N12968, N12960, N9017, N4850);
not NOT1 (N12969, N12959);
buf BUF1 (N12970, N12968);
nand NAND3 (N12971, N12970, N7077, N1848);
buf BUF1 (N12972, N12969);
xor XOR2 (N12973, N12964, N2442);
not NOT1 (N12974, N12962);
nand NAND2 (N12975, N12973, N7537);
nand NAND2 (N12976, N12965, N11426);
or OR4 (N12977, N12950, N4910, N4298, N10307);
not NOT1 (N12978, N12975);
or OR2 (N12979, N12974, N5779);
buf BUF1 (N12980, N12963);
not NOT1 (N12981, N12966);
or OR2 (N12982, N12972, N2235);
not NOT1 (N12983, N12980);
xor XOR2 (N12984, N12954, N3927);
and AND2 (N12985, N12983, N9095);
and AND3 (N12986, N12985, N171, N4709);
nand NAND3 (N12987, N12978, N9255, N9374);
nand NAND2 (N12988, N12986, N9506);
nor NOR2 (N12989, N12982, N8252);
xor XOR2 (N12990, N12977, N10839);
nor NOR2 (N12991, N12988, N11939);
xor XOR2 (N12992, N12990, N10416);
not NOT1 (N12993, N12992);
not NOT1 (N12994, N12991);
nand NAND4 (N12995, N12971, N2744, N3217, N8383);
and AND3 (N12996, N12995, N5850, N8418);
or OR2 (N12997, N12967, N9168);
nor NOR2 (N12998, N12987, N12905);
nor NOR2 (N12999, N12996, N3160);
nor NOR3 (N13000, N12993, N4322, N2542);
nor NOR3 (N13001, N12976, N6725, N1430);
not NOT1 (N13002, N12989);
not NOT1 (N13003, N12981);
and AND2 (N13004, N13002, N7761);
buf BUF1 (N13005, N12997);
not NOT1 (N13006, N13004);
or OR4 (N13007, N13000, N3590, N11795, N6566);
not NOT1 (N13008, N12999);
xor XOR2 (N13009, N13001, N12990);
and AND2 (N13010, N12984, N9309);
not NOT1 (N13011, N13006);
and AND2 (N13012, N12998, N9615);
xor XOR2 (N13013, N13007, N2862);
or OR3 (N13014, N13011, N1685, N11459);
or OR3 (N13015, N13014, N327, N9317);
or OR2 (N13016, N13009, N11678);
xor XOR2 (N13017, N13016, N11241);
not NOT1 (N13018, N13008);
xor XOR2 (N13019, N13012, N4689);
buf BUF1 (N13020, N13003);
not NOT1 (N13021, N13017);
buf BUF1 (N13022, N13013);
not NOT1 (N13023, N12979);
and AND2 (N13024, N13018, N24);
buf BUF1 (N13025, N12994);
nand NAND2 (N13026, N13015, N1845);
and AND4 (N13027, N13021, N8001, N1637, N9057);
not NOT1 (N13028, N13025);
nor NOR4 (N13029, N13023, N7168, N10671, N3738);
or OR3 (N13030, N13020, N3560, N8321);
xor XOR2 (N13031, N13019, N7336);
xor XOR2 (N13032, N13010, N7745);
xor XOR2 (N13033, N13005, N590);
or OR3 (N13034, N13027, N2658, N4421);
not NOT1 (N13035, N13033);
nor NOR2 (N13036, N13032, N9867);
xor XOR2 (N13037, N13024, N520);
xor XOR2 (N13038, N13036, N11317);
nor NOR3 (N13039, N13028, N3804, N5305);
or OR4 (N13040, N13035, N934, N6108, N5390);
or OR2 (N13041, N13034, N294);
xor XOR2 (N13042, N13037, N6036);
and AND2 (N13043, N13026, N2059);
nor NOR4 (N13044, N13022, N7375, N12820, N9634);
or OR4 (N13045, N13041, N8768, N5876, N13044);
nor NOR2 (N13046, N6431, N6066);
not NOT1 (N13047, N13039);
or OR3 (N13048, N13030, N10369, N601);
xor XOR2 (N13049, N13043, N7171);
nand NAND4 (N13050, N13045, N10047, N11427, N10287);
nor NOR2 (N13051, N13046, N10460);
and AND4 (N13052, N13051, N3173, N7279, N2042);
xor XOR2 (N13053, N13031, N3253);
and AND4 (N13054, N13048, N4895, N12620, N6351);
and AND4 (N13055, N13054, N12334, N10211, N6476);
xor XOR2 (N13056, N13029, N6334);
not NOT1 (N13057, N13049);
nor NOR2 (N13058, N13057, N9493);
buf BUF1 (N13059, N13056);
nand NAND3 (N13060, N13050, N8469, N11557);
nand NAND3 (N13061, N13055, N1086, N10253);
and AND4 (N13062, N13038, N2396, N1882, N3426);
or OR2 (N13063, N13058, N7883);
not NOT1 (N13064, N13059);
nand NAND4 (N13065, N13040, N1084, N8399, N3590);
nand NAND4 (N13066, N13047, N1109, N12569, N4057);
not NOT1 (N13067, N13042);
nor NOR2 (N13068, N13053, N9384);
not NOT1 (N13069, N13063);
or OR3 (N13070, N13067, N10210, N8762);
xor XOR2 (N13071, N13061, N494);
or OR4 (N13072, N13070, N1038, N1960, N6096);
buf BUF1 (N13073, N13072);
not NOT1 (N13074, N13071);
buf BUF1 (N13075, N13052);
nor NOR4 (N13076, N13073, N11845, N1301, N9122);
buf BUF1 (N13077, N13060);
nand NAND2 (N13078, N13066, N9324);
not NOT1 (N13079, N13064);
or OR4 (N13080, N13062, N9288, N5893, N12522);
xor XOR2 (N13081, N13077, N1834);
and AND2 (N13082, N13075, N2755);
not NOT1 (N13083, N13079);
nand NAND3 (N13084, N13065, N12265, N8171);
not NOT1 (N13085, N13076);
not NOT1 (N13086, N13068);
and AND4 (N13087, N13080, N7795, N11472, N7129);
nor NOR3 (N13088, N13078, N360, N1623);
not NOT1 (N13089, N13083);
and AND2 (N13090, N13082, N7184);
and AND2 (N13091, N13084, N7840);
not NOT1 (N13092, N13086);
buf BUF1 (N13093, N13074);
nand NAND3 (N13094, N13089, N6723, N9864);
nand NAND2 (N13095, N13091, N6488);
and AND4 (N13096, N13085, N7848, N12877, N7845);
or OR2 (N13097, N13069, N8971);
not NOT1 (N13098, N13088);
not NOT1 (N13099, N13096);
and AND3 (N13100, N13097, N947, N6837);
or OR4 (N13101, N13094, N6019, N3825, N2987);
or OR2 (N13102, N13092, N10907);
or OR2 (N13103, N13081, N7989);
nand NAND4 (N13104, N13095, N12191, N3358, N6057);
not NOT1 (N13105, N13087);
xor XOR2 (N13106, N13105, N100);
xor XOR2 (N13107, N13099, N12837);
xor XOR2 (N13108, N13103, N9194);
or OR4 (N13109, N13106, N2671, N1389, N12343);
xor XOR2 (N13110, N13102, N7054);
nand NAND4 (N13111, N13110, N11650, N6846, N7749);
not NOT1 (N13112, N13104);
and AND3 (N13113, N13093, N4226, N704);
or OR2 (N13114, N13107, N3025);
nand NAND4 (N13115, N13090, N4994, N10737, N3047);
or OR4 (N13116, N13113, N5329, N7187, N12378);
nand NAND2 (N13117, N13108, N11254);
nor NOR3 (N13118, N13100, N5918, N4707);
nor NOR2 (N13119, N13118, N8756);
buf BUF1 (N13120, N13114);
buf BUF1 (N13121, N13119);
nand NAND4 (N13122, N13120, N7948, N769, N8830);
xor XOR2 (N13123, N13101, N9352);
nand NAND4 (N13124, N13121, N6760, N8254, N2451);
xor XOR2 (N13125, N13122, N365);
buf BUF1 (N13126, N13111);
and AND3 (N13127, N13109, N7739, N8126);
xor XOR2 (N13128, N13112, N10599);
and AND4 (N13129, N13125, N670, N11548, N10715);
nand NAND2 (N13130, N13128, N3488);
or OR3 (N13131, N13098, N12919, N5542);
nor NOR4 (N13132, N13124, N6408, N495, N7374);
or OR4 (N13133, N13132, N3685, N6160, N3461);
and AND4 (N13134, N13116, N4568, N9035, N7380);
not NOT1 (N13135, N13129);
xor XOR2 (N13136, N13134, N9601);
nor NOR2 (N13137, N13117, N748);
buf BUF1 (N13138, N13133);
and AND3 (N13139, N13136, N4655, N8546);
nor NOR4 (N13140, N13123, N7745, N8369, N7537);
and AND3 (N13141, N13135, N8494, N5050);
xor XOR2 (N13142, N13126, N4562);
nand NAND4 (N13143, N13130, N9640, N7597, N3781);
xor XOR2 (N13144, N13139, N5624);
buf BUF1 (N13145, N13127);
xor XOR2 (N13146, N13131, N13027);
nand NAND2 (N13147, N13141, N8260);
not NOT1 (N13148, N13144);
nand NAND3 (N13149, N13137, N2735, N12373);
nand NAND2 (N13150, N13143, N5132);
and AND4 (N13151, N13150, N2159, N9309, N3751);
xor XOR2 (N13152, N13138, N4474);
not NOT1 (N13153, N13152);
nor NOR4 (N13154, N13147, N10951, N7865, N9158);
buf BUF1 (N13155, N13146);
nand NAND3 (N13156, N13148, N277, N8882);
not NOT1 (N13157, N13142);
buf BUF1 (N13158, N13154);
or OR3 (N13159, N13158, N12713, N5297);
xor XOR2 (N13160, N13115, N6270);
not NOT1 (N13161, N13159);
not NOT1 (N13162, N13155);
and AND2 (N13163, N13161, N9166);
or OR2 (N13164, N13153, N8247);
not NOT1 (N13165, N13162);
xor XOR2 (N13166, N13140, N5642);
xor XOR2 (N13167, N13166, N4209);
xor XOR2 (N13168, N13145, N8533);
not NOT1 (N13169, N13151);
nor NOR4 (N13170, N13169, N4875, N10708, N7637);
and AND4 (N13171, N13163, N4416, N6131, N1833);
nand NAND3 (N13172, N13160, N2370, N3203);
nand NAND2 (N13173, N13149, N7800);
and AND4 (N13174, N13168, N9984, N5924, N12755);
and AND4 (N13175, N13173, N214, N9418, N8415);
and AND4 (N13176, N13157, N3810, N7541, N11647);
or OR2 (N13177, N13174, N5706);
nand NAND3 (N13178, N13167, N2357, N4587);
not NOT1 (N13179, N13172);
nor NOR4 (N13180, N13176, N11550, N8397, N8636);
nor NOR3 (N13181, N13165, N6755, N9797);
or OR3 (N13182, N13180, N8444, N3584);
nand NAND3 (N13183, N13175, N24, N4323);
buf BUF1 (N13184, N13177);
nand NAND2 (N13185, N13164, N3891);
and AND4 (N13186, N13171, N3245, N7937, N5986);
and AND3 (N13187, N13186, N2217, N1583);
nand NAND4 (N13188, N13179, N11471, N8232, N2895);
not NOT1 (N13189, N13185);
nand NAND2 (N13190, N13181, N6015);
nor NOR3 (N13191, N13184, N6759, N1792);
and AND4 (N13192, N13170, N9583, N5321, N523);
and AND3 (N13193, N13191, N1055, N8624);
xor XOR2 (N13194, N13183, N7621);
nor NOR2 (N13195, N13178, N8858);
buf BUF1 (N13196, N13195);
buf BUF1 (N13197, N13190);
or OR2 (N13198, N13194, N3561);
buf BUF1 (N13199, N13156);
nand NAND2 (N13200, N13198, N1047);
and AND3 (N13201, N13188, N2957, N10633);
and AND4 (N13202, N13189, N7077, N2251, N10201);
buf BUF1 (N13203, N13187);
and AND3 (N13204, N13192, N8282, N4305);
xor XOR2 (N13205, N13196, N4649);
nor NOR3 (N13206, N13202, N9303, N6643);
not NOT1 (N13207, N13193);
xor XOR2 (N13208, N13182, N10301);
and AND4 (N13209, N13205, N3113, N10671, N12985);
not NOT1 (N13210, N13208);
nor NOR3 (N13211, N13201, N318, N4091);
or OR4 (N13212, N13197, N6609, N7632, N10973);
nand NAND3 (N13213, N13204, N11407, N5979);
nor NOR3 (N13214, N13213, N832, N1114);
buf BUF1 (N13215, N13200);
nand NAND4 (N13216, N13203, N11421, N6057, N9253);
or OR2 (N13217, N13211, N12443);
or OR2 (N13218, N13217, N508);
and AND2 (N13219, N13207, N11063);
and AND4 (N13220, N13219, N8834, N4078, N1308);
nand NAND2 (N13221, N13199, N2710);
nor NOR3 (N13222, N13210, N5293, N1267);
nand NAND4 (N13223, N13218, N7657, N5142, N12168);
nand NAND2 (N13224, N13214, N2967);
xor XOR2 (N13225, N13220, N7482);
buf BUF1 (N13226, N13206);
buf BUF1 (N13227, N13222);
nor NOR2 (N13228, N13209, N8159);
or OR4 (N13229, N13225, N4789, N7811, N10929);
not NOT1 (N13230, N13215);
and AND4 (N13231, N13224, N6940, N10711, N446);
or OR4 (N13232, N13221, N10234, N12356, N4575);
xor XOR2 (N13233, N13228, N6143);
and AND3 (N13234, N13226, N8536, N2942);
xor XOR2 (N13235, N13216, N9766);
nand NAND4 (N13236, N13232, N9053, N7960, N12598);
xor XOR2 (N13237, N13230, N949);
nand NAND2 (N13238, N13227, N13208);
nand NAND3 (N13239, N13234, N4591, N9003);
and AND2 (N13240, N13233, N11594);
nand NAND4 (N13241, N13223, N5299, N7637, N11200);
not NOT1 (N13242, N13236);
and AND3 (N13243, N13231, N3647, N12567);
xor XOR2 (N13244, N13240, N9280);
not NOT1 (N13245, N13242);
or OR2 (N13246, N13241, N6439);
xor XOR2 (N13247, N13243, N4937);
xor XOR2 (N13248, N13237, N5079);
xor XOR2 (N13249, N13229, N12255);
xor XOR2 (N13250, N13239, N11256);
xor XOR2 (N13251, N13238, N2201);
or OR3 (N13252, N13251, N69, N6206);
nor NOR3 (N13253, N13248, N968, N39);
nand NAND4 (N13254, N13244, N10514, N9805, N12152);
nand NAND3 (N13255, N13235, N9410, N12347);
xor XOR2 (N13256, N13245, N11997);
xor XOR2 (N13257, N13246, N10648);
and AND4 (N13258, N13253, N4334, N10708, N10584);
or OR4 (N13259, N13255, N1602, N12350, N7669);
or OR2 (N13260, N13252, N5542);
xor XOR2 (N13261, N13257, N5611);
nand NAND3 (N13262, N13254, N2011, N2423);
not NOT1 (N13263, N13212);
nand NAND3 (N13264, N13250, N2158, N7928);
nor NOR3 (N13265, N13264, N2900, N2460);
nor NOR2 (N13266, N13262, N13010);
not NOT1 (N13267, N13265);
buf BUF1 (N13268, N13261);
and AND2 (N13269, N13247, N5023);
nand NAND2 (N13270, N13268, N3028);
nor NOR3 (N13271, N13260, N1770, N11505);
not NOT1 (N13272, N13263);
buf BUF1 (N13273, N13272);
not NOT1 (N13274, N13270);
xor XOR2 (N13275, N13256, N3132);
xor XOR2 (N13276, N13258, N7014);
or OR3 (N13277, N13269, N12848, N1111);
buf BUF1 (N13278, N13275);
nand NAND3 (N13279, N13274, N8584, N8060);
nand NAND3 (N13280, N13267, N3528, N9595);
xor XOR2 (N13281, N13279, N8831);
not NOT1 (N13282, N13273);
nor NOR4 (N13283, N13278, N7180, N3017, N242);
or OR4 (N13284, N13259, N9879, N4274, N7274);
nand NAND2 (N13285, N13277, N6492);
buf BUF1 (N13286, N13276);
not NOT1 (N13287, N13286);
not NOT1 (N13288, N13271);
buf BUF1 (N13289, N13266);
nand NAND3 (N13290, N13282, N5310, N1366);
or OR3 (N13291, N13288, N7880, N3483);
buf BUF1 (N13292, N13283);
or OR4 (N13293, N13249, N9938, N11902, N10069);
nor NOR3 (N13294, N13292, N12586, N12411);
xor XOR2 (N13295, N13289, N3280);
buf BUF1 (N13296, N13291);
nand NAND4 (N13297, N13284, N9416, N155, N8994);
xor XOR2 (N13298, N13293, N6730);
and AND4 (N13299, N13290, N8792, N12682, N2725);
nand NAND2 (N13300, N13298, N7800);
or OR2 (N13301, N13296, N12996);
nand NAND3 (N13302, N13297, N2593, N7084);
nand NAND3 (N13303, N13302, N10002, N1298);
buf BUF1 (N13304, N13303);
or OR3 (N13305, N13287, N3187, N5223);
xor XOR2 (N13306, N13294, N8135);
xor XOR2 (N13307, N13301, N2951);
nand NAND4 (N13308, N13300, N3130, N6624, N1325);
nor NOR4 (N13309, N13308, N10474, N8141, N12735);
or OR2 (N13310, N13295, N6390);
xor XOR2 (N13311, N13305, N5227);
not NOT1 (N13312, N13306);
and AND2 (N13313, N13309, N9030);
xor XOR2 (N13314, N13311, N1251);
or OR2 (N13315, N13285, N7394);
buf BUF1 (N13316, N13312);
and AND2 (N13317, N13281, N2919);
and AND4 (N13318, N13317, N9957, N5467, N2602);
xor XOR2 (N13319, N13313, N2519);
not NOT1 (N13320, N13310);
xor XOR2 (N13321, N13315, N6741);
and AND4 (N13322, N13280, N9862, N6425, N6975);
and AND2 (N13323, N13299, N10163);
and AND4 (N13324, N13318, N10698, N635, N12713);
not NOT1 (N13325, N13316);
and AND4 (N13326, N13320, N1927, N5706, N2439);
or OR2 (N13327, N13307, N991);
not NOT1 (N13328, N13327);
xor XOR2 (N13329, N13314, N226);
or OR4 (N13330, N13329, N13086, N2405, N7080);
buf BUF1 (N13331, N13330);
buf BUF1 (N13332, N13321);
not NOT1 (N13333, N13332);
not NOT1 (N13334, N13319);
not NOT1 (N13335, N13333);
not NOT1 (N13336, N13304);
xor XOR2 (N13337, N13322, N2576);
not NOT1 (N13338, N13325);
nand NAND4 (N13339, N13334, N12708, N5540, N9394);
or OR4 (N13340, N13337, N8531, N5202, N8605);
nand NAND4 (N13341, N13328, N967, N2452, N8324);
not NOT1 (N13342, N13335);
or OR3 (N13343, N13331, N341, N960);
and AND2 (N13344, N13338, N12397);
and AND3 (N13345, N13344, N7020, N7251);
nand NAND3 (N13346, N13340, N8091, N3164);
buf BUF1 (N13347, N13339);
buf BUF1 (N13348, N13345);
xor XOR2 (N13349, N13326, N12898);
and AND3 (N13350, N13324, N5039, N13224);
nand NAND2 (N13351, N13350, N6734);
buf BUF1 (N13352, N13342);
nand NAND3 (N13353, N13341, N9312, N1785);
xor XOR2 (N13354, N13336, N417);
buf BUF1 (N13355, N13351);
xor XOR2 (N13356, N13347, N9934);
not NOT1 (N13357, N13349);
or OR3 (N13358, N13346, N1281, N8318);
buf BUF1 (N13359, N13343);
not NOT1 (N13360, N13359);
buf BUF1 (N13361, N13355);
not NOT1 (N13362, N13361);
or OR3 (N13363, N13353, N13122, N1637);
and AND3 (N13364, N13348, N9441, N7571);
or OR3 (N13365, N13364, N13276, N7858);
or OR4 (N13366, N13357, N7456, N3948, N1100);
not NOT1 (N13367, N13362);
or OR2 (N13368, N13358, N8821);
and AND2 (N13369, N13360, N11640);
nor NOR2 (N13370, N13363, N449);
or OR3 (N13371, N13365, N5821, N11981);
or OR2 (N13372, N13323, N8626);
xor XOR2 (N13373, N13370, N8888);
nor NOR3 (N13374, N13352, N4964, N10506);
not NOT1 (N13375, N13356);
buf BUF1 (N13376, N13371);
nor NOR3 (N13377, N13369, N10889, N3327);
not NOT1 (N13378, N13374);
buf BUF1 (N13379, N13354);
buf BUF1 (N13380, N13367);
not NOT1 (N13381, N13377);
and AND4 (N13382, N13376, N7873, N11532, N1761);
xor XOR2 (N13383, N13380, N186);
not NOT1 (N13384, N13375);
xor XOR2 (N13385, N13382, N830);
buf BUF1 (N13386, N13372);
nor NOR3 (N13387, N13368, N5048, N10214);
and AND4 (N13388, N13384, N7748, N12908, N11115);
not NOT1 (N13389, N13381);
and AND3 (N13390, N13383, N7902, N2892);
xor XOR2 (N13391, N13390, N12500);
nor NOR3 (N13392, N13379, N1389, N7171);
or OR2 (N13393, N13385, N10736);
nand NAND4 (N13394, N13393, N12360, N3314, N8104);
not NOT1 (N13395, N13378);
and AND2 (N13396, N13387, N7417);
nor NOR4 (N13397, N13396, N9867, N199, N10486);
xor XOR2 (N13398, N13373, N11446);
not NOT1 (N13399, N13394);
nor NOR2 (N13400, N13388, N2954);
nand NAND2 (N13401, N13389, N637);
nor NOR4 (N13402, N13395, N13252, N13265, N3951);
or OR4 (N13403, N13399, N4280, N2107, N12398);
nand NAND2 (N13404, N13401, N3506);
and AND4 (N13405, N13402, N10046, N5506, N10471);
buf BUF1 (N13406, N13397);
or OR4 (N13407, N13391, N6427, N13146, N6849);
or OR4 (N13408, N13386, N3604, N3571, N8265);
and AND4 (N13409, N13404, N9746, N10354, N3509);
or OR4 (N13410, N13406, N1865, N10158, N2320);
xor XOR2 (N13411, N13403, N13023);
or OR3 (N13412, N13405, N12199, N6098);
and AND4 (N13413, N13412, N562, N2837, N8430);
xor XOR2 (N13414, N13408, N5747);
and AND3 (N13415, N13398, N13101, N6654);
or OR4 (N13416, N13409, N8694, N9927, N8500);
buf BUF1 (N13417, N13415);
or OR2 (N13418, N13413, N7794);
nand NAND4 (N13419, N13410, N6664, N3753, N12067);
nor NOR3 (N13420, N13419, N10944, N11670);
nor NOR4 (N13421, N13407, N1282, N11940, N5664);
nand NAND2 (N13422, N13418, N1650);
nand NAND2 (N13423, N13366, N4911);
buf BUF1 (N13424, N13416);
xor XOR2 (N13425, N13422, N11607);
and AND3 (N13426, N13421, N5377, N6408);
buf BUF1 (N13427, N13411);
and AND2 (N13428, N13420, N10797);
nor NOR4 (N13429, N13392, N4197, N1938, N13010);
xor XOR2 (N13430, N13400, N7214);
nor NOR3 (N13431, N13428, N3837, N5654);
and AND3 (N13432, N13427, N8040, N534);
nor NOR3 (N13433, N13431, N8042, N11285);
xor XOR2 (N13434, N13426, N5744);
and AND4 (N13435, N13434, N10817, N188, N8466);
or OR3 (N13436, N13429, N12558, N2941);
nor NOR2 (N13437, N13424, N9729);
xor XOR2 (N13438, N13423, N8756);
and AND4 (N13439, N13430, N1090, N3029, N12156);
xor XOR2 (N13440, N13438, N2226);
xor XOR2 (N13441, N13440, N7642);
not NOT1 (N13442, N13435);
or OR2 (N13443, N13425, N7833);
xor XOR2 (N13444, N13436, N7229);
nor NOR3 (N13445, N13442, N12050, N6818);
buf BUF1 (N13446, N13444);
not NOT1 (N13447, N13433);
or OR3 (N13448, N13414, N9963, N6848);
not NOT1 (N13449, N13446);
and AND2 (N13450, N13417, N9855);
not NOT1 (N13451, N13441);
nor NOR4 (N13452, N13451, N12573, N11274, N2821);
and AND3 (N13453, N13452, N1879, N11387);
nor NOR3 (N13454, N13447, N7951, N10081);
buf BUF1 (N13455, N13439);
or OR2 (N13456, N13448, N9737);
not NOT1 (N13457, N13450);
not NOT1 (N13458, N13453);
not NOT1 (N13459, N13456);
nand NAND2 (N13460, N13457, N13420);
or OR3 (N13461, N13460, N250, N9091);
nor NOR3 (N13462, N13461, N3280, N10163);
nor NOR2 (N13463, N13462, N5030);
and AND2 (N13464, N13459, N8344);
or OR4 (N13465, N13445, N4827, N612, N7767);
or OR3 (N13466, N13449, N10966, N10677);
not NOT1 (N13467, N13458);
and AND3 (N13468, N13466, N602, N4303);
or OR4 (N13469, N13443, N5648, N5692, N7695);
or OR4 (N13470, N13464, N5828, N11953, N12147);
buf BUF1 (N13471, N13432);
or OR2 (N13472, N13471, N239);
not NOT1 (N13473, N13467);
xor XOR2 (N13474, N13468, N10825);
buf BUF1 (N13475, N13472);
buf BUF1 (N13476, N13475);
xor XOR2 (N13477, N13455, N2478);
nand NAND3 (N13478, N13465, N12067, N6982);
xor XOR2 (N13479, N13437, N3707);
not NOT1 (N13480, N13454);
buf BUF1 (N13481, N13480);
not NOT1 (N13482, N13478);
and AND2 (N13483, N13470, N187);
or OR2 (N13484, N13483, N1420);
or OR3 (N13485, N13479, N10622, N1835);
buf BUF1 (N13486, N13473);
nor NOR3 (N13487, N13485, N10970, N4800);
nand NAND2 (N13488, N13487, N7091);
xor XOR2 (N13489, N13488, N12258);
or OR3 (N13490, N13476, N10477, N3784);
not NOT1 (N13491, N13481);
and AND3 (N13492, N13490, N12138, N9162);
nor NOR3 (N13493, N13489, N10180, N5846);
xor XOR2 (N13494, N13482, N6641);
buf BUF1 (N13495, N13477);
or OR4 (N13496, N13474, N12507, N12832, N5892);
and AND2 (N13497, N13491, N3097);
not NOT1 (N13498, N13494);
buf BUF1 (N13499, N13484);
xor XOR2 (N13500, N13486, N10014);
and AND3 (N13501, N13463, N8859, N304);
nor NOR3 (N13502, N13497, N11758, N11233);
nand NAND2 (N13503, N13495, N8646);
or OR4 (N13504, N13493, N11819, N5087, N8130);
buf BUF1 (N13505, N13498);
or OR2 (N13506, N13496, N11750);
nor NOR2 (N13507, N13503, N13495);
not NOT1 (N13508, N13506);
xor XOR2 (N13509, N13492, N8931);
and AND2 (N13510, N13502, N10977);
or OR3 (N13511, N13504, N6941, N2266);
nand NAND3 (N13512, N13507, N11165, N10863);
not NOT1 (N13513, N13509);
and AND3 (N13514, N13508, N6648, N1411);
or OR3 (N13515, N13514, N4726, N8477);
and AND3 (N13516, N13511, N2062, N4667);
xor XOR2 (N13517, N13515, N4165);
nor NOR4 (N13518, N13516, N11115, N2186, N4989);
nand NAND4 (N13519, N13505, N8446, N12920, N11679);
or OR3 (N13520, N13469, N4401, N1394);
not NOT1 (N13521, N13520);
or OR3 (N13522, N13512, N5250, N8307);
nand NAND4 (N13523, N13499, N1400, N6519, N5610);
or OR4 (N13524, N13523, N1903, N4474, N6607);
buf BUF1 (N13525, N13500);
and AND4 (N13526, N13525, N991, N12856, N10979);
xor XOR2 (N13527, N13518, N3736);
buf BUF1 (N13528, N13517);
nand NAND3 (N13529, N13521, N10250, N11025);
and AND2 (N13530, N13524, N10995);
buf BUF1 (N13531, N13510);
nand NAND3 (N13532, N13519, N2656, N2);
xor XOR2 (N13533, N13532, N1179);
nor NOR2 (N13534, N13529, N12065);
buf BUF1 (N13535, N13527);
or OR3 (N13536, N13533, N11645, N10454);
buf BUF1 (N13537, N13530);
xor XOR2 (N13538, N13535, N13504);
not NOT1 (N13539, N13538);
xor XOR2 (N13540, N13531, N5861);
xor XOR2 (N13541, N13501, N3377);
or OR3 (N13542, N13522, N912, N6006);
nor NOR4 (N13543, N13542, N3506, N12844, N12078);
nor NOR2 (N13544, N13536, N7914);
and AND4 (N13545, N13541, N4383, N8530, N12076);
buf BUF1 (N13546, N13539);
not NOT1 (N13547, N13544);
or OR4 (N13548, N13545, N6456, N1919, N1161);
and AND4 (N13549, N13537, N531, N656, N1939);
buf BUF1 (N13550, N13526);
nor NOR3 (N13551, N13528, N5898, N11964);
nand NAND2 (N13552, N13550, N5469);
and AND2 (N13553, N13546, N7986);
buf BUF1 (N13554, N13540);
xor XOR2 (N13555, N13548, N8977);
buf BUF1 (N13556, N13555);
nor NOR3 (N13557, N13534, N13067, N2325);
buf BUF1 (N13558, N13551);
or OR3 (N13559, N13543, N8759, N4099);
xor XOR2 (N13560, N13559, N2172);
buf BUF1 (N13561, N13558);
or OR4 (N13562, N13513, N3286, N4596, N9504);
and AND3 (N13563, N13547, N13542, N6943);
nand NAND2 (N13564, N13561, N6885);
buf BUF1 (N13565, N13563);
nor NOR4 (N13566, N13557, N538, N2717, N9097);
nor NOR2 (N13567, N13549, N6092);
xor XOR2 (N13568, N13566, N6445);
or OR2 (N13569, N13564, N6196);
buf BUF1 (N13570, N13568);
and AND4 (N13571, N13560, N6773, N12093, N2309);
not NOT1 (N13572, N13562);
xor XOR2 (N13573, N13567, N8927);
and AND4 (N13574, N13565, N6320, N3755, N8076);
or OR4 (N13575, N13571, N10286, N11767, N660);
not NOT1 (N13576, N13556);
nand NAND2 (N13577, N13553, N11774);
xor XOR2 (N13578, N13574, N9618);
nor NOR4 (N13579, N13572, N10917, N12215, N7899);
and AND3 (N13580, N13578, N10421, N12951);
nand NAND3 (N13581, N13552, N12285, N1109);
buf BUF1 (N13582, N13580);
xor XOR2 (N13583, N13554, N2834);
or OR2 (N13584, N13582, N7301);
nor NOR2 (N13585, N13581, N39);
buf BUF1 (N13586, N13577);
nand NAND2 (N13587, N13573, N11820);
and AND2 (N13588, N13579, N11659);
buf BUF1 (N13589, N13586);
nor NOR3 (N13590, N13588, N5904, N12469);
nand NAND2 (N13591, N13590, N3584);
or OR2 (N13592, N13584, N8904);
xor XOR2 (N13593, N13570, N9559);
xor XOR2 (N13594, N13591, N11602);
nand NAND3 (N13595, N13593, N7946, N12982);
or OR4 (N13596, N13594, N3377, N13535, N6188);
nand NAND4 (N13597, N13587, N7705, N2965, N4837);
xor XOR2 (N13598, N13583, N1196);
xor XOR2 (N13599, N13595, N12734);
nand NAND3 (N13600, N13596, N3835, N4359);
nor NOR2 (N13601, N13569, N9608);
not NOT1 (N13602, N13585);
and AND4 (N13603, N13575, N5002, N5678, N12699);
buf BUF1 (N13604, N13603);
buf BUF1 (N13605, N13597);
or OR3 (N13606, N13589, N5174, N1507);
not NOT1 (N13607, N13605);
not NOT1 (N13608, N13606);
xor XOR2 (N13609, N13607, N7495);
nand NAND4 (N13610, N13592, N3595, N10203, N761);
buf BUF1 (N13611, N13601);
not NOT1 (N13612, N13610);
nor NOR2 (N13613, N13602, N6396);
buf BUF1 (N13614, N13613);
and AND3 (N13615, N13576, N874, N1603);
or OR3 (N13616, N13604, N8230, N3368);
nor NOR4 (N13617, N13599, N8032, N7650, N6908);
or OR4 (N13618, N13615, N6301, N4079, N5683);
and AND4 (N13619, N13612, N2868, N5255, N10695);
buf BUF1 (N13620, N13617);
not NOT1 (N13621, N13611);
nand NAND3 (N13622, N13616, N9913, N4442);
xor XOR2 (N13623, N13620, N13535);
buf BUF1 (N13624, N13622);
nor NOR3 (N13625, N13598, N12108, N4326);
or OR4 (N13626, N13618, N497, N10231, N9606);
xor XOR2 (N13627, N13600, N2568);
nand NAND4 (N13628, N13614, N9359, N10943, N6918);
nand NAND4 (N13629, N13626, N258, N13033, N5682);
or OR2 (N13630, N13619, N1675);
nor NOR3 (N13631, N13629, N9121, N13488);
and AND3 (N13632, N13608, N7456, N1129);
or OR3 (N13633, N13625, N10425, N12333);
xor XOR2 (N13634, N13627, N6676);
buf BUF1 (N13635, N13628);
and AND2 (N13636, N13623, N3389);
nor NOR4 (N13637, N13621, N12730, N3393, N4686);
and AND3 (N13638, N13634, N11393, N8133);
nand NAND2 (N13639, N13624, N7797);
and AND2 (N13640, N13635, N3913);
and AND2 (N13641, N13640, N11190);
nand NAND2 (N13642, N13609, N13373);
buf BUF1 (N13643, N13641);
nand NAND4 (N13644, N13643, N3197, N10107, N8243);
xor XOR2 (N13645, N13638, N5195);
nand NAND2 (N13646, N13632, N5377);
nand NAND3 (N13647, N13642, N11033, N13489);
nand NAND3 (N13648, N13630, N6966, N11585);
or OR3 (N13649, N13631, N10087, N9009);
or OR2 (N13650, N13636, N12144);
and AND2 (N13651, N13646, N4349);
not NOT1 (N13652, N13647);
or OR4 (N13653, N13650, N537, N11802, N8913);
buf BUF1 (N13654, N13645);
or OR4 (N13655, N13649, N11067, N11669, N6853);
nand NAND4 (N13656, N13648, N7597, N10066, N5341);
or OR4 (N13657, N13653, N2463, N9169, N5414);
nand NAND3 (N13658, N13639, N1824, N11559);
nor NOR4 (N13659, N13656, N11586, N1449, N5559);
xor XOR2 (N13660, N13657, N2685);
nand NAND2 (N13661, N13658, N12711);
not NOT1 (N13662, N13661);
not NOT1 (N13663, N13633);
nor NOR3 (N13664, N13659, N10430, N3886);
and AND4 (N13665, N13660, N8396, N5175, N1778);
nand NAND4 (N13666, N13665, N3847, N11673, N12066);
or OR3 (N13667, N13666, N5802, N4081);
nor NOR2 (N13668, N13652, N11076);
and AND3 (N13669, N13668, N5609, N6424);
and AND3 (N13670, N13663, N13091, N11732);
nor NOR4 (N13671, N13670, N13384, N2027, N5435);
buf BUF1 (N13672, N13654);
buf BUF1 (N13673, N13667);
and AND3 (N13674, N13672, N3759, N11618);
nor NOR2 (N13675, N13671, N6965);
or OR4 (N13676, N13662, N12773, N12067, N10609);
and AND3 (N13677, N13673, N5013, N13458);
buf BUF1 (N13678, N13674);
buf BUF1 (N13679, N13655);
nor NOR3 (N13680, N13637, N11750, N8932);
nor NOR3 (N13681, N13678, N3766, N13582);
not NOT1 (N13682, N13679);
buf BUF1 (N13683, N13680);
and AND4 (N13684, N13677, N4944, N13119, N4280);
xor XOR2 (N13685, N13675, N9906);
not NOT1 (N13686, N13651);
buf BUF1 (N13687, N13664);
or OR3 (N13688, N13686, N337, N4391);
not NOT1 (N13689, N13681);
buf BUF1 (N13690, N13644);
and AND3 (N13691, N13690, N12496, N4216);
nand NAND3 (N13692, N13685, N8821, N7650);
nor NOR3 (N13693, N13684, N3043, N5117);
nor NOR3 (N13694, N13689, N8381, N9226);
nor NOR4 (N13695, N13693, N1247, N8949, N8590);
xor XOR2 (N13696, N13682, N682);
xor XOR2 (N13697, N13687, N4425);
xor XOR2 (N13698, N13688, N10718);
or OR2 (N13699, N13692, N12679);
nor NOR2 (N13700, N13694, N7800);
nand NAND3 (N13701, N13696, N10053, N12264);
xor XOR2 (N13702, N13697, N2299);
and AND3 (N13703, N13683, N2429, N5213);
xor XOR2 (N13704, N13676, N3526);
nand NAND4 (N13705, N13703, N375, N2703, N11493);
and AND4 (N13706, N13702, N6582, N10951, N6203);
and AND3 (N13707, N13704, N5112, N12541);
xor XOR2 (N13708, N13691, N4598);
buf BUF1 (N13709, N13701);
nor NOR2 (N13710, N13698, N4268);
not NOT1 (N13711, N13695);
buf BUF1 (N13712, N13705);
and AND3 (N13713, N13706, N3521, N5831);
nor NOR2 (N13714, N13707, N13514);
xor XOR2 (N13715, N13712, N13318);
nand NAND2 (N13716, N13714, N8998);
and AND4 (N13717, N13709, N12468, N12610, N7291);
xor XOR2 (N13718, N13708, N3567);
buf BUF1 (N13719, N13699);
nor NOR4 (N13720, N13710, N10412, N169, N10097);
not NOT1 (N13721, N13716);
nand NAND3 (N13722, N13711, N13609, N1915);
buf BUF1 (N13723, N13717);
buf BUF1 (N13724, N13715);
nand NAND2 (N13725, N13719, N6726);
xor XOR2 (N13726, N13720, N9401);
buf BUF1 (N13727, N13669);
nand NAND2 (N13728, N13723, N10219);
buf BUF1 (N13729, N13728);
and AND2 (N13730, N13724, N9044);
not NOT1 (N13731, N13721);
or OR2 (N13732, N13725, N12934);
xor XOR2 (N13733, N13731, N8081);
buf BUF1 (N13734, N13713);
nand NAND3 (N13735, N13727, N4782, N9941);
or OR4 (N13736, N13700, N9996, N4617, N1341);
and AND3 (N13737, N13734, N637, N8399);
xor XOR2 (N13738, N13729, N7401);
xor XOR2 (N13739, N13730, N12638);
xor XOR2 (N13740, N13737, N10467);
not NOT1 (N13741, N13739);
and AND2 (N13742, N13736, N12714);
nor NOR3 (N13743, N13740, N12326, N3113);
nor NOR4 (N13744, N13733, N13230, N6160, N9083);
nand NAND3 (N13745, N13743, N4622, N3637);
or OR2 (N13746, N13735, N4438);
nor NOR2 (N13747, N13742, N6305);
or OR2 (N13748, N13741, N10467);
not NOT1 (N13749, N13745);
xor XOR2 (N13750, N13738, N3839);
nand NAND3 (N13751, N13744, N9515, N7906);
xor XOR2 (N13752, N13722, N8140);
nand NAND3 (N13753, N13726, N13523, N890);
xor XOR2 (N13754, N13747, N5894);
and AND4 (N13755, N13732, N12543, N7899, N6782);
or OR2 (N13756, N13752, N4820);
and AND2 (N13757, N13755, N8544);
and AND3 (N13758, N13750, N4692, N11240);
and AND3 (N13759, N13753, N886, N12147);
nand NAND3 (N13760, N13758, N11314, N4626);
not NOT1 (N13761, N13760);
or OR3 (N13762, N13754, N9950, N7514);
nand NAND2 (N13763, N13761, N8037);
buf BUF1 (N13764, N13756);
and AND4 (N13765, N13746, N13208, N2259, N3284);
xor XOR2 (N13766, N13759, N8505);
nand NAND3 (N13767, N13763, N12816, N3605);
xor XOR2 (N13768, N13748, N9649);
nand NAND4 (N13769, N13766, N4860, N8930, N3247);
nor NOR4 (N13770, N13757, N1524, N7195, N10253);
nand NAND4 (N13771, N13769, N1147, N12281, N8765);
buf BUF1 (N13772, N13765);
nand NAND2 (N13773, N13770, N5633);
or OR4 (N13774, N13768, N6168, N3851, N5719);
nand NAND4 (N13775, N13718, N3015, N11817, N11281);
buf BUF1 (N13776, N13751);
and AND2 (N13777, N13762, N8898);
xor XOR2 (N13778, N13776, N11035);
not NOT1 (N13779, N13778);
not NOT1 (N13780, N13771);
xor XOR2 (N13781, N13779, N11282);
buf BUF1 (N13782, N13772);
not NOT1 (N13783, N13782);
buf BUF1 (N13784, N13773);
not NOT1 (N13785, N13767);
and AND4 (N13786, N13781, N10262, N5048, N11764);
buf BUF1 (N13787, N13784);
not NOT1 (N13788, N13777);
not NOT1 (N13789, N13783);
not NOT1 (N13790, N13749);
not NOT1 (N13791, N13787);
and AND4 (N13792, N13785, N7801, N7940, N1183);
nand NAND2 (N13793, N13774, N2212);
and AND3 (N13794, N13790, N6065, N7774);
or OR3 (N13795, N13788, N987, N13133);
buf BUF1 (N13796, N13764);
and AND3 (N13797, N13789, N4220, N2260);
buf BUF1 (N13798, N13791);
or OR2 (N13799, N13792, N5540);
buf BUF1 (N13800, N13798);
and AND2 (N13801, N13775, N3118);
or OR3 (N13802, N13800, N8433, N9532);
buf BUF1 (N13803, N13801);
nor NOR4 (N13804, N13795, N9331, N10924, N12651);
not NOT1 (N13805, N13803);
and AND2 (N13806, N13797, N4638);
nand NAND3 (N13807, N13802, N5948, N2195);
or OR3 (N13808, N13807, N7663, N5997);
xor XOR2 (N13809, N13804, N7312);
buf BUF1 (N13810, N13780);
nor NOR2 (N13811, N13799, N7364);
nand NAND3 (N13812, N13809, N7786, N13383);
xor XOR2 (N13813, N13810, N7950);
not NOT1 (N13814, N13811);
nor NOR3 (N13815, N13793, N8069, N1228);
nor NOR2 (N13816, N13805, N845);
buf BUF1 (N13817, N13814);
buf BUF1 (N13818, N13794);
nor NOR4 (N13819, N13813, N13813, N5081, N1128);
and AND4 (N13820, N13817, N10728, N13429, N1786);
nor NOR4 (N13821, N13816, N3711, N6694, N10903);
nor NOR4 (N13822, N13815, N13558, N8429, N8181);
buf BUF1 (N13823, N13819);
xor XOR2 (N13824, N13821, N2454);
xor XOR2 (N13825, N13786, N7051);
not NOT1 (N13826, N13806);
nor NOR3 (N13827, N13824, N10201, N4884);
nand NAND3 (N13828, N13826, N4058, N10810);
nor NOR4 (N13829, N13822, N4918, N7985, N12904);
nand NAND2 (N13830, N13812, N11793);
nor NOR3 (N13831, N13823, N264, N4682);
buf BUF1 (N13832, N13828);
buf BUF1 (N13833, N13832);
nand NAND4 (N13834, N13818, N9521, N1218, N10032);
and AND2 (N13835, N13834, N11729);
nor NOR2 (N13836, N13833, N11571);
or OR4 (N13837, N13831, N7022, N2678, N944);
nand NAND4 (N13838, N13825, N1214, N4819, N5858);
nand NAND3 (N13839, N13820, N8399, N13817);
or OR2 (N13840, N13836, N7769);
buf BUF1 (N13841, N13796);
or OR3 (N13842, N13841, N5575, N8798);
or OR3 (N13843, N13808, N4719, N217);
and AND2 (N13844, N13843, N9478);
and AND3 (N13845, N13829, N7033, N6127);
and AND3 (N13846, N13840, N4660, N10833);
nor NOR4 (N13847, N13837, N10244, N9845, N6259);
xor XOR2 (N13848, N13839, N12726);
or OR2 (N13849, N13838, N13201);
buf BUF1 (N13850, N13842);
and AND3 (N13851, N13827, N8514, N11087);
and AND2 (N13852, N13848, N5926);
buf BUF1 (N13853, N13850);
buf BUF1 (N13854, N13852);
nor NOR3 (N13855, N13851, N1365, N1606);
buf BUF1 (N13856, N13847);
xor XOR2 (N13857, N13830, N13366);
buf BUF1 (N13858, N13846);
nand NAND2 (N13859, N13857, N5406);
nand NAND2 (N13860, N13856, N8942);
or OR2 (N13861, N13844, N5516);
xor XOR2 (N13862, N13861, N4827);
nand NAND3 (N13863, N13862, N3989, N735);
nor NOR2 (N13864, N13835, N7396);
xor XOR2 (N13865, N13858, N4916);
or OR2 (N13866, N13849, N1497);
nor NOR4 (N13867, N13865, N3291, N7289, N13668);
or OR3 (N13868, N13845, N6886, N5443);
and AND2 (N13869, N13864, N1958);
not NOT1 (N13870, N13855);
buf BUF1 (N13871, N13863);
or OR2 (N13872, N13868, N9935);
nor NOR2 (N13873, N13854, N2898);
or OR4 (N13874, N13860, N12308, N9932, N2640);
or OR2 (N13875, N13872, N9787);
nor NOR3 (N13876, N13866, N11945, N647);
nor NOR4 (N13877, N13870, N13040, N12462, N9204);
and AND3 (N13878, N13853, N9727, N6537);
and AND3 (N13879, N13867, N10185, N12121);
and AND2 (N13880, N13875, N3228);
or OR2 (N13881, N13859, N5409);
xor XOR2 (N13882, N13877, N6380);
nand NAND2 (N13883, N13871, N11752);
not NOT1 (N13884, N13881);
not NOT1 (N13885, N13882);
or OR2 (N13886, N13884, N13199);
nor NOR4 (N13887, N13869, N6265, N13270, N3165);
nor NOR3 (N13888, N13880, N9034, N2297);
and AND2 (N13889, N13888, N10961);
nor NOR3 (N13890, N13883, N1599, N10905);
buf BUF1 (N13891, N13887);
and AND2 (N13892, N13878, N9169);
xor XOR2 (N13893, N13879, N9011);
xor XOR2 (N13894, N13893, N4347);
and AND4 (N13895, N13889, N1973, N7503, N1323);
buf BUF1 (N13896, N13892);
nor NOR4 (N13897, N13874, N7278, N6937, N8536);
and AND2 (N13898, N13891, N13233);
and AND3 (N13899, N13886, N12335, N1082);
not NOT1 (N13900, N13890);
nand NAND2 (N13901, N13900, N9679);
or OR3 (N13902, N13873, N11080, N443);
xor XOR2 (N13903, N13898, N2954);
and AND3 (N13904, N13903, N10651, N7787);
and AND3 (N13905, N13895, N7312, N12632);
and AND2 (N13906, N13897, N11765);
or OR3 (N13907, N13899, N5891, N9947);
xor XOR2 (N13908, N13896, N1596);
or OR3 (N13909, N13904, N5230, N11907);
buf BUF1 (N13910, N13909);
nand NAND4 (N13911, N13902, N7041, N2572, N4882);
and AND4 (N13912, N13908, N1651, N8918, N1848);
or OR2 (N13913, N13894, N6014);
or OR3 (N13914, N13912, N7908, N2955);
nor NOR3 (N13915, N13907, N12153, N2316);
nor NOR4 (N13916, N13915, N2994, N7579, N2117);
nor NOR4 (N13917, N13910, N7788, N11539, N13168);
buf BUF1 (N13918, N13913);
nand NAND2 (N13919, N13914, N3214);
or OR4 (N13920, N13885, N6654, N355, N3798);
nor NOR2 (N13921, N13911, N8530);
nor NOR4 (N13922, N13916, N11313, N8852, N697);
buf BUF1 (N13923, N13922);
xor XOR2 (N13924, N13919, N5937);
and AND3 (N13925, N13876, N7146, N6622);
and AND3 (N13926, N13925, N6249, N37);
xor XOR2 (N13927, N13905, N1996);
nor NOR3 (N13928, N13924, N6200, N1435);
and AND3 (N13929, N13901, N10731, N13149);
not NOT1 (N13930, N13923);
nand NAND2 (N13931, N13927, N8312);
buf BUF1 (N13932, N13931);
buf BUF1 (N13933, N13926);
and AND4 (N13934, N13920, N8240, N7530, N3527);
not NOT1 (N13935, N13934);
and AND2 (N13936, N13935, N2304);
nor NOR3 (N13937, N13932, N10158, N324);
not NOT1 (N13938, N13930);
nor NOR4 (N13939, N13917, N1484, N12623, N12536);
xor XOR2 (N13940, N13918, N4548);
or OR3 (N13941, N13937, N5394, N9110);
not NOT1 (N13942, N13940);
nand NAND2 (N13943, N13936, N12989);
and AND4 (N13944, N13938, N4586, N11415, N6257);
and AND4 (N13945, N13939, N8532, N6822, N6556);
nand NAND3 (N13946, N13928, N1586, N1431);
or OR4 (N13947, N13942, N11941, N6974, N13115);
xor XOR2 (N13948, N13933, N3918);
or OR2 (N13949, N13944, N6524);
and AND3 (N13950, N13949, N7300, N10153);
and AND4 (N13951, N13906, N12229, N2552, N11227);
and AND4 (N13952, N13941, N11960, N6155, N3980);
nor NOR2 (N13953, N13946, N11164);
or OR3 (N13954, N13945, N1015, N3798);
nor NOR2 (N13955, N13929, N5268);
nor NOR3 (N13956, N13948, N3268, N7786);
nand NAND3 (N13957, N13950, N6090, N7267);
or OR4 (N13958, N13943, N5318, N3324, N12298);
nand NAND3 (N13959, N13956, N10008, N6336);
nor NOR4 (N13960, N13921, N5031, N13386, N8931);
buf BUF1 (N13961, N13953);
not NOT1 (N13962, N13954);
nor NOR4 (N13963, N13960, N11598, N3622, N11784);
not NOT1 (N13964, N13952);
or OR4 (N13965, N13963, N3312, N4109, N11771);
nand NAND2 (N13966, N13955, N12164);
not NOT1 (N13967, N13951);
xor XOR2 (N13968, N13966, N3682);
or OR2 (N13969, N13961, N11579);
or OR2 (N13970, N13962, N11848);
or OR3 (N13971, N13947, N9758, N1965);
nor NOR4 (N13972, N13957, N2656, N5917, N10301);
nor NOR3 (N13973, N13969, N12119, N1164);
buf BUF1 (N13974, N13965);
or OR4 (N13975, N13964, N3675, N4852, N6762);
not NOT1 (N13976, N13972);
nor NOR3 (N13977, N13958, N12674, N5910);
buf BUF1 (N13978, N13970);
and AND3 (N13979, N13974, N6627, N5831);
buf BUF1 (N13980, N13977);
xor XOR2 (N13981, N13976, N1465);
buf BUF1 (N13982, N13979);
or OR3 (N13983, N13973, N8253, N10058);
not NOT1 (N13984, N13978);
xor XOR2 (N13985, N13981, N9824);
not NOT1 (N13986, N13984);
nand NAND2 (N13987, N13971, N12440);
nor NOR4 (N13988, N13968, N9934, N4031, N1161);
buf BUF1 (N13989, N13983);
buf BUF1 (N13990, N13980);
or OR3 (N13991, N13959, N4005, N2655);
not NOT1 (N13992, N13986);
nor NOR4 (N13993, N13982, N333, N13599, N8785);
not NOT1 (N13994, N13987);
nor NOR2 (N13995, N13975, N4275);
and AND2 (N13996, N13992, N13463);
nand NAND2 (N13997, N13996, N2380);
not NOT1 (N13998, N13990);
or OR4 (N13999, N13994, N5317, N3487, N10590);
nor NOR4 (N14000, N13999, N11502, N12162, N3434);
and AND4 (N14001, N14000, N10003, N11637, N6127);
nor NOR3 (N14002, N13988, N368, N13700);
not NOT1 (N14003, N13998);
nor NOR2 (N14004, N14002, N3933);
nand NAND4 (N14005, N13985, N12090, N12652, N9161);
xor XOR2 (N14006, N14001, N1125);
nor NOR4 (N14007, N14005, N13082, N4383, N1408);
nor NOR3 (N14008, N14003, N267, N4975);
nor NOR4 (N14009, N14004, N8079, N1515, N12155);
xor XOR2 (N14010, N14008, N12932);
or OR2 (N14011, N13993, N13187);
nor NOR2 (N14012, N14011, N11424);
and AND2 (N14013, N13995, N2082);
xor XOR2 (N14014, N14013, N7848);
nand NAND4 (N14015, N13989, N7252, N13129, N9325);
xor XOR2 (N14016, N14006, N4166);
and AND3 (N14017, N14015, N652, N2530);
not NOT1 (N14018, N13991);
xor XOR2 (N14019, N13997, N3828);
xor XOR2 (N14020, N14014, N4537);
xor XOR2 (N14021, N14020, N5691);
nor NOR3 (N14022, N14018, N10550, N5868);
or OR4 (N14023, N14012, N8721, N5203, N7496);
xor XOR2 (N14024, N14022, N12947);
not NOT1 (N14025, N14009);
xor XOR2 (N14026, N14023, N3057);
or OR3 (N14027, N14021, N5673, N11594);
buf BUF1 (N14028, N14026);
nor NOR2 (N14029, N14025, N1844);
buf BUF1 (N14030, N14028);
nand NAND4 (N14031, N14007, N10424, N5100, N2514);
nand NAND2 (N14032, N14027, N4522);
xor XOR2 (N14033, N14016, N3037);
or OR2 (N14034, N14030, N4192);
not NOT1 (N14035, N14031);
nand NAND2 (N14036, N14019, N12444);
buf BUF1 (N14037, N14032);
nor NOR4 (N14038, N14035, N9213, N13873, N3759);
buf BUF1 (N14039, N14029);
not NOT1 (N14040, N14034);
not NOT1 (N14041, N13967);
buf BUF1 (N14042, N14040);
buf BUF1 (N14043, N14042);
and AND3 (N14044, N14043, N8253, N6510);
xor XOR2 (N14045, N14044, N12407);
or OR2 (N14046, N14010, N13161);
buf BUF1 (N14047, N14045);
xor XOR2 (N14048, N14047, N5776);
and AND3 (N14049, N14033, N5871, N4558);
nor NOR2 (N14050, N14049, N2937);
or OR3 (N14051, N14050, N175, N9018);
xor XOR2 (N14052, N14048, N12958);
and AND3 (N14053, N14046, N2453, N11185);
and AND4 (N14054, N14052, N11904, N4456, N13620);
and AND4 (N14055, N14054, N13869, N7164, N1136);
and AND4 (N14056, N14053, N7423, N1194, N11);
or OR2 (N14057, N14017, N7647);
and AND3 (N14058, N14037, N444, N2311);
and AND4 (N14059, N14036, N4750, N11570, N13184);
buf BUF1 (N14060, N14039);
or OR3 (N14061, N14060, N9717, N11658);
xor XOR2 (N14062, N14041, N11998);
or OR2 (N14063, N14055, N6720);
nor NOR2 (N14064, N14038, N7615);
nor NOR3 (N14065, N14051, N5230, N2824);
nand NAND3 (N14066, N14065, N11663, N1655);
and AND3 (N14067, N14063, N7993, N1439);
and AND3 (N14068, N14067, N2830, N13699);
or OR3 (N14069, N14059, N13253, N6898);
not NOT1 (N14070, N14058);
or OR2 (N14071, N14024, N12902);
xor XOR2 (N14072, N14066, N10871);
not NOT1 (N14073, N14057);
buf BUF1 (N14074, N14072);
nor NOR3 (N14075, N14056, N10643, N8744);
buf BUF1 (N14076, N14061);
nand NAND2 (N14077, N14062, N792);
not NOT1 (N14078, N14068);
buf BUF1 (N14079, N14078);
xor XOR2 (N14080, N14075, N6304);
xor XOR2 (N14081, N14070, N12705);
not NOT1 (N14082, N14064);
nand NAND2 (N14083, N14073, N12794);
and AND2 (N14084, N14077, N1345);
not NOT1 (N14085, N14081);
not NOT1 (N14086, N14079);
nand NAND3 (N14087, N14069, N12062, N528);
or OR2 (N14088, N14071, N13518);
xor XOR2 (N14089, N14082, N12471);
buf BUF1 (N14090, N14085);
or OR2 (N14091, N14087, N8199);
xor XOR2 (N14092, N14080, N12345);
xor XOR2 (N14093, N14089, N7980);
or OR4 (N14094, N14074, N8285, N3717, N503);
xor XOR2 (N14095, N14094, N9740);
buf BUF1 (N14096, N14092);
nor NOR2 (N14097, N14086, N11017);
or OR4 (N14098, N14084, N462, N3758, N7021);
nor NOR4 (N14099, N14091, N10028, N3263, N9753);
buf BUF1 (N14100, N14097);
nor NOR4 (N14101, N14100, N2353, N9097, N561);
not NOT1 (N14102, N14083);
nand NAND4 (N14103, N14095, N12218, N8102, N2823);
xor XOR2 (N14104, N14076, N838);
xor XOR2 (N14105, N14099, N3438);
nand NAND3 (N14106, N14096, N4990, N3260);
nor NOR2 (N14107, N14103, N11625);
buf BUF1 (N14108, N14102);
not NOT1 (N14109, N14106);
nor NOR3 (N14110, N14107, N11276, N12640);
not NOT1 (N14111, N14090);
and AND4 (N14112, N14110, N8015, N10748, N1811);
and AND3 (N14113, N14109, N11726, N5976);
nand NAND3 (N14114, N14105, N1060, N1219);
xor XOR2 (N14115, N14098, N12157);
not NOT1 (N14116, N14104);
and AND3 (N14117, N14093, N10662, N5093);
buf BUF1 (N14118, N14101);
not NOT1 (N14119, N14117);
and AND3 (N14120, N14116, N3565, N13062);
nor NOR3 (N14121, N14113, N10687, N4666);
nand NAND3 (N14122, N14121, N7776, N4479);
nor NOR4 (N14123, N14122, N9431, N3829, N5846);
nor NOR2 (N14124, N14111, N2839);
nor NOR4 (N14125, N14112, N4272, N1493, N7241);
xor XOR2 (N14126, N14125, N4310);
and AND3 (N14127, N14108, N12944, N7957);
not NOT1 (N14128, N14114);
not NOT1 (N14129, N14126);
xor XOR2 (N14130, N14088, N1179);
or OR4 (N14131, N14123, N8919, N5507, N2852);
xor XOR2 (N14132, N14128, N13330);
nor NOR4 (N14133, N14124, N8625, N2875, N5516);
nand NAND2 (N14134, N14132, N6889);
or OR3 (N14135, N14133, N13504, N14130);
not NOT1 (N14136, N3812);
and AND3 (N14137, N14131, N785, N11873);
nand NAND3 (N14138, N14136, N13625, N234);
not NOT1 (N14139, N14119);
buf BUF1 (N14140, N14129);
or OR2 (N14141, N14138, N6501);
not NOT1 (N14142, N14141);
not NOT1 (N14143, N14127);
not NOT1 (N14144, N14120);
and AND2 (N14145, N14144, N5912);
nand NAND3 (N14146, N14142, N5074, N1256);
xor XOR2 (N14147, N14146, N5085);
not NOT1 (N14148, N14137);
nor NOR4 (N14149, N14140, N4970, N9638, N11190);
xor XOR2 (N14150, N14147, N779);
not NOT1 (N14151, N14143);
not NOT1 (N14152, N14139);
buf BUF1 (N14153, N14145);
nand NAND2 (N14154, N14135, N3888);
buf BUF1 (N14155, N14115);
and AND3 (N14156, N14150, N7111, N6481);
and AND2 (N14157, N14149, N8399);
not NOT1 (N14158, N14154);
buf BUF1 (N14159, N14118);
and AND3 (N14160, N14158, N6418, N9725);
and AND3 (N14161, N14148, N13753, N5510);
and AND2 (N14162, N14155, N13779);
not NOT1 (N14163, N14153);
xor XOR2 (N14164, N14134, N9635);
buf BUF1 (N14165, N14164);
or OR2 (N14166, N14156, N13035);
nor NOR3 (N14167, N14162, N1258, N5769);
nand NAND4 (N14168, N14163, N6817, N2828, N11029);
buf BUF1 (N14169, N14157);
buf BUF1 (N14170, N14161);
xor XOR2 (N14171, N14168, N7924);
or OR4 (N14172, N14170, N12842, N7458, N8783);
and AND3 (N14173, N14171, N3675, N8943);
not NOT1 (N14174, N14172);
nand NAND3 (N14175, N14167, N8560, N2802);
or OR3 (N14176, N14166, N2781, N12933);
nand NAND3 (N14177, N14160, N12630, N8087);
and AND2 (N14178, N14169, N9169);
xor XOR2 (N14179, N14175, N1071);
xor XOR2 (N14180, N14176, N2598);
or OR4 (N14181, N14177, N4501, N7104, N5175);
xor XOR2 (N14182, N14151, N5488);
buf BUF1 (N14183, N14165);
not NOT1 (N14184, N14183);
nor NOR2 (N14185, N14152, N7096);
not NOT1 (N14186, N14185);
or OR3 (N14187, N14178, N2392, N1393);
and AND3 (N14188, N14159, N12123, N11871);
nand NAND2 (N14189, N14181, N6035);
nor NOR4 (N14190, N14180, N1481, N5825, N9704);
nor NOR4 (N14191, N14173, N3036, N5096, N7530);
nand NAND3 (N14192, N14179, N10531, N5468);
nand NAND3 (N14193, N14190, N9228, N8082);
or OR4 (N14194, N14182, N11280, N1941, N8370);
and AND3 (N14195, N14189, N693, N9399);
buf BUF1 (N14196, N14184);
xor XOR2 (N14197, N14194, N3182);
xor XOR2 (N14198, N14192, N11467);
xor XOR2 (N14199, N14188, N4836);
or OR2 (N14200, N14186, N8023);
nand NAND2 (N14201, N14198, N9081);
buf BUF1 (N14202, N14201);
nor NOR3 (N14203, N14191, N1220, N6821);
buf BUF1 (N14204, N14197);
and AND3 (N14205, N14196, N9687, N208);
buf BUF1 (N14206, N14199);
nor NOR2 (N14207, N14174, N13204);
nand NAND2 (N14208, N14187, N2386);
xor XOR2 (N14209, N14208, N481);
nand NAND2 (N14210, N14205, N11523);
nand NAND2 (N14211, N14203, N2284);
nand NAND4 (N14212, N14200, N6930, N8798, N13101);
buf BUF1 (N14213, N14206);
and AND4 (N14214, N14210, N7928, N10102, N13510);
not NOT1 (N14215, N14202);
buf BUF1 (N14216, N14214);
nand NAND3 (N14217, N14204, N1197, N12769);
or OR2 (N14218, N14207, N11521);
or OR2 (N14219, N14213, N8521);
not NOT1 (N14220, N14212);
buf BUF1 (N14221, N14218);
xor XOR2 (N14222, N14219, N11198);
nand NAND3 (N14223, N14221, N12155, N9647);
nand NAND4 (N14224, N14222, N647, N8374, N1805);
or OR2 (N14225, N14211, N1350);
or OR3 (N14226, N14209, N7408, N3537);
and AND4 (N14227, N14220, N2339, N106, N8327);
nand NAND3 (N14228, N14224, N8615, N1842);
or OR4 (N14229, N14225, N9238, N3144, N12762);
nand NAND4 (N14230, N14215, N12340, N8542, N4366);
xor XOR2 (N14231, N14223, N260);
not NOT1 (N14232, N14217);
nand NAND4 (N14233, N14193, N3426, N14084, N121);
buf BUF1 (N14234, N14232);
nand NAND3 (N14235, N14227, N7255, N5529);
and AND2 (N14236, N14235, N7849);
and AND2 (N14237, N14236, N12784);
and AND2 (N14238, N14228, N4517);
and AND4 (N14239, N14195, N7125, N8185, N13321);
and AND4 (N14240, N14233, N13158, N4135, N10883);
not NOT1 (N14241, N14226);
and AND2 (N14242, N14238, N1504);
nor NOR3 (N14243, N14216, N4878, N12122);
not NOT1 (N14244, N14231);
nand NAND3 (N14245, N14229, N10733, N1506);
not NOT1 (N14246, N14239);
and AND2 (N14247, N14240, N1443);
and AND2 (N14248, N14245, N11845);
or OR2 (N14249, N14230, N4332);
buf BUF1 (N14250, N14247);
or OR4 (N14251, N14246, N3637, N11410, N7064);
and AND2 (N14252, N14241, N14120);
or OR4 (N14253, N14249, N11568, N1129, N5211);
nor NOR3 (N14254, N14252, N2284, N5997);
xor XOR2 (N14255, N14254, N130);
or OR2 (N14256, N14237, N5212);
buf BUF1 (N14257, N14250);
xor XOR2 (N14258, N14251, N4834);
buf BUF1 (N14259, N14258);
nor NOR2 (N14260, N14253, N498);
or OR3 (N14261, N14248, N11253, N6093);
buf BUF1 (N14262, N14259);
or OR2 (N14263, N14243, N6524);
nor NOR3 (N14264, N14263, N13460, N14084);
not NOT1 (N14265, N14256);
buf BUF1 (N14266, N14255);
xor XOR2 (N14267, N14260, N2481);
buf BUF1 (N14268, N14262);
nor NOR2 (N14269, N14234, N6678);
and AND4 (N14270, N14244, N9024, N7482, N3267);
or OR3 (N14271, N14265, N7589, N6183);
nor NOR2 (N14272, N14266, N2475);
xor XOR2 (N14273, N14261, N4015);
nand NAND4 (N14274, N14268, N10070, N9391, N8937);
nor NOR3 (N14275, N14269, N2313, N10814);
nand NAND4 (N14276, N14257, N3052, N5382, N6461);
nor NOR2 (N14277, N14267, N9143);
xor XOR2 (N14278, N14270, N11885);
not NOT1 (N14279, N14277);
and AND3 (N14280, N14276, N4105, N12882);
xor XOR2 (N14281, N14278, N541);
buf BUF1 (N14282, N14281);
xor XOR2 (N14283, N14242, N9175);
or OR2 (N14284, N14275, N11753);
xor XOR2 (N14285, N14272, N12687);
nand NAND3 (N14286, N14273, N8955, N3438);
xor XOR2 (N14287, N14285, N4351);
nand NAND4 (N14288, N14280, N1873, N2461, N11825);
or OR3 (N14289, N14287, N14183, N12436);
or OR2 (N14290, N14279, N8298);
nor NOR4 (N14291, N14284, N11248, N5876, N13153);
nor NOR4 (N14292, N14283, N4799, N1870, N2712);
xor XOR2 (N14293, N14289, N393);
nand NAND3 (N14294, N14271, N3523, N14065);
nand NAND3 (N14295, N14292, N1731, N867);
xor XOR2 (N14296, N14295, N3981);
not NOT1 (N14297, N14274);
xor XOR2 (N14298, N14293, N9293);
buf BUF1 (N14299, N14296);
buf BUF1 (N14300, N14291);
xor XOR2 (N14301, N14297, N173);
nor NOR2 (N14302, N14299, N1045);
xor XOR2 (N14303, N14290, N6016);
buf BUF1 (N14304, N14298);
or OR3 (N14305, N14303, N7432, N8706);
nor NOR3 (N14306, N14302, N13784, N5645);
nor NOR4 (N14307, N14282, N4459, N1263, N254);
nand NAND4 (N14308, N14307, N4277, N2180, N6436);
and AND3 (N14309, N14308, N10027, N4883);
and AND3 (N14310, N14264, N12109, N4156);
buf BUF1 (N14311, N14294);
or OR3 (N14312, N14306, N7631, N4730);
xor XOR2 (N14313, N14310, N13912);
and AND2 (N14314, N14286, N2262);
nand NAND4 (N14315, N14305, N3022, N2395, N610);
not NOT1 (N14316, N14314);
and AND2 (N14317, N14288, N4973);
or OR3 (N14318, N14300, N188, N10259);
not NOT1 (N14319, N14311);
nor NOR2 (N14320, N14316, N1901);
buf BUF1 (N14321, N14309);
not NOT1 (N14322, N14321);
nor NOR4 (N14323, N14318, N9382, N8565, N10415);
or OR4 (N14324, N14319, N7215, N12948, N6587);
nor NOR3 (N14325, N14304, N7089, N7764);
xor XOR2 (N14326, N14322, N10549);
nor NOR3 (N14327, N14325, N5435, N1358);
or OR3 (N14328, N14317, N8862, N3293);
nor NOR3 (N14329, N14313, N5787, N2817);
or OR3 (N14330, N14323, N1361, N14084);
buf BUF1 (N14331, N14329);
xor XOR2 (N14332, N14330, N10982);
and AND2 (N14333, N14327, N11563);
not NOT1 (N14334, N14331);
nor NOR3 (N14335, N14315, N10311, N4295);
xor XOR2 (N14336, N14326, N9757);
nand NAND3 (N14337, N14333, N13355, N2291);
nor NOR4 (N14338, N14335, N2278, N2097, N712);
nor NOR2 (N14339, N14312, N6681);
and AND2 (N14340, N14338, N7591);
nand NAND4 (N14341, N14301, N4643, N8857, N10521);
nor NOR2 (N14342, N14339, N8270);
buf BUF1 (N14343, N14336);
or OR4 (N14344, N14340, N2414, N2461, N2984);
nand NAND2 (N14345, N14324, N13860);
and AND3 (N14346, N14342, N11639, N2717);
and AND2 (N14347, N14332, N150);
nor NOR3 (N14348, N14341, N6907, N2246);
and AND3 (N14349, N14343, N6052, N13947);
buf BUF1 (N14350, N14345);
nand NAND4 (N14351, N14328, N6452, N3481, N3105);
and AND3 (N14352, N14344, N6364, N2939);
not NOT1 (N14353, N14351);
nand NAND3 (N14354, N14346, N3209, N9527);
nand NAND3 (N14355, N14349, N4107, N1017);
xor XOR2 (N14356, N14352, N10554);
or OR3 (N14357, N14320, N3368, N1105);
buf BUF1 (N14358, N14350);
xor XOR2 (N14359, N14354, N9878);
buf BUF1 (N14360, N14358);
buf BUF1 (N14361, N14337);
and AND2 (N14362, N14361, N14359);
and AND2 (N14363, N4002, N8710);
nor NOR2 (N14364, N14356, N5406);
buf BUF1 (N14365, N14360);
not NOT1 (N14366, N14355);
or OR2 (N14367, N14362, N8374);
xor XOR2 (N14368, N14365, N12511);
xor XOR2 (N14369, N14367, N3905);
not NOT1 (N14370, N14364);
and AND3 (N14371, N14368, N1725, N8067);
and AND3 (N14372, N14357, N9832, N2883);
and AND2 (N14373, N14363, N7445);
nand NAND2 (N14374, N14369, N7136);
nand NAND3 (N14375, N14371, N5183, N11516);
not NOT1 (N14376, N14347);
nor NOR2 (N14377, N14334, N8488);
not NOT1 (N14378, N14377);
or OR3 (N14379, N14370, N13944, N6453);
or OR2 (N14380, N14373, N10673);
nand NAND4 (N14381, N14380, N6867, N8359, N8479);
nor NOR3 (N14382, N14378, N11626, N5969);
or OR2 (N14383, N14374, N2106);
or OR2 (N14384, N14379, N1777);
xor XOR2 (N14385, N14375, N797);
not NOT1 (N14386, N14372);
nor NOR3 (N14387, N14376, N6704, N11019);
not NOT1 (N14388, N14385);
not NOT1 (N14389, N14382);
buf BUF1 (N14390, N14353);
buf BUF1 (N14391, N14348);
buf BUF1 (N14392, N14383);
not NOT1 (N14393, N14381);
buf BUF1 (N14394, N14387);
xor XOR2 (N14395, N14394, N5193);
xor XOR2 (N14396, N14388, N78);
xor XOR2 (N14397, N14389, N5192);
xor XOR2 (N14398, N14396, N10393);
or OR3 (N14399, N14390, N12516, N3321);
not NOT1 (N14400, N14384);
not NOT1 (N14401, N14393);
xor XOR2 (N14402, N14391, N4708);
xor XOR2 (N14403, N14401, N182);
not NOT1 (N14404, N14399);
nand NAND2 (N14405, N14395, N2393);
and AND3 (N14406, N14403, N11661, N9569);
and AND3 (N14407, N14398, N13838, N13262);
buf BUF1 (N14408, N14392);
nor NOR2 (N14409, N14407, N2737);
xor XOR2 (N14410, N14397, N11150);
nor NOR3 (N14411, N14404, N875, N3093);
or OR3 (N14412, N14411, N7723, N10017);
buf BUF1 (N14413, N14366);
nand NAND2 (N14414, N14409, N5906);
and AND2 (N14415, N14400, N5827);
nand NAND4 (N14416, N14414, N2129, N5386, N8848);
nand NAND3 (N14417, N14408, N11520, N10421);
xor XOR2 (N14418, N14416, N11623);
nor NOR3 (N14419, N14413, N4919, N13041);
nand NAND3 (N14420, N14405, N13288, N12688);
buf BUF1 (N14421, N14410);
and AND4 (N14422, N14386, N1977, N4504, N13480);
xor XOR2 (N14423, N14422, N2738);
and AND4 (N14424, N14418, N2714, N85, N13348);
nand NAND2 (N14425, N14424, N4922);
nor NOR4 (N14426, N14415, N10724, N3110, N12765);
or OR2 (N14427, N14421, N11912);
nor NOR3 (N14428, N14420, N4845, N10237);
nand NAND2 (N14429, N14426, N12822);
buf BUF1 (N14430, N14402);
not NOT1 (N14431, N14427);
buf BUF1 (N14432, N14417);
or OR2 (N14433, N14428, N11884);
and AND4 (N14434, N14406, N14082, N14123, N1871);
and AND2 (N14435, N14419, N11226);
or OR4 (N14436, N14412, N6646, N13242, N4687);
not NOT1 (N14437, N14432);
xor XOR2 (N14438, N14435, N13041);
nor NOR4 (N14439, N14423, N13050, N5806, N5819);
xor XOR2 (N14440, N14436, N6099);
not NOT1 (N14441, N14437);
or OR3 (N14442, N14434, N4149, N9735);
not NOT1 (N14443, N14431);
nor NOR4 (N14444, N14433, N9481, N10723, N11344);
nand NAND4 (N14445, N14439, N9094, N870, N9991);
or OR2 (N14446, N14425, N14424);
and AND3 (N14447, N14440, N2105, N12492);
nand NAND3 (N14448, N14445, N2354, N9483);
nor NOR4 (N14449, N14446, N4138, N5701, N562);
nor NOR4 (N14450, N14449, N5023, N7818, N3050);
or OR2 (N14451, N14429, N14069);
nor NOR2 (N14452, N14444, N2433);
buf BUF1 (N14453, N14443);
not NOT1 (N14454, N14447);
xor XOR2 (N14455, N14441, N11103);
and AND4 (N14456, N14454, N10212, N7661, N12678);
nand NAND2 (N14457, N14450, N4676);
and AND3 (N14458, N14453, N1426, N13840);
nor NOR2 (N14459, N14430, N12581);
or OR3 (N14460, N14442, N1448, N3026);
nor NOR3 (N14461, N14451, N6127, N69);
nand NAND3 (N14462, N14457, N9264, N8340);
nand NAND4 (N14463, N14462, N6273, N5612, N8001);
not NOT1 (N14464, N14463);
nand NAND2 (N14465, N14464, N11460);
or OR4 (N14466, N14459, N11481, N11730, N560);
or OR4 (N14467, N14458, N5850, N6147, N13608);
xor XOR2 (N14468, N14455, N4163);
or OR2 (N14469, N14460, N4308);
and AND4 (N14470, N14456, N8206, N12150, N13167);
xor XOR2 (N14471, N14461, N2227);
buf BUF1 (N14472, N14470);
and AND4 (N14473, N14468, N13875, N1781, N9083);
nor NOR4 (N14474, N14448, N10714, N2258, N8215);
nor NOR3 (N14475, N14469, N4730, N14101);
buf BUF1 (N14476, N14474);
not NOT1 (N14477, N14471);
not NOT1 (N14478, N14452);
and AND3 (N14479, N14466, N6216, N123);
and AND2 (N14480, N14478, N10103);
xor XOR2 (N14481, N14477, N11910);
and AND4 (N14482, N14467, N9418, N3197, N3045);
nand NAND4 (N14483, N14475, N1219, N2251, N13873);
nand NAND3 (N14484, N14483, N7319, N14003);
not NOT1 (N14485, N14473);
or OR2 (N14486, N14465, N10764);
or OR3 (N14487, N14480, N1502, N3732);
xor XOR2 (N14488, N14476, N9147);
nor NOR4 (N14489, N14482, N4909, N11232, N8736);
nor NOR2 (N14490, N14488, N8813);
nor NOR2 (N14491, N14479, N6789);
and AND3 (N14492, N14485, N1583, N1345);
or OR4 (N14493, N14472, N7894, N14003, N7603);
xor XOR2 (N14494, N14484, N3385);
nor NOR3 (N14495, N14486, N5850, N3673);
or OR2 (N14496, N14438, N7415);
nor NOR3 (N14497, N14481, N10866, N2457);
and AND4 (N14498, N14487, N13315, N861, N12888);
xor XOR2 (N14499, N14491, N11049);
not NOT1 (N14500, N14497);
not NOT1 (N14501, N14490);
buf BUF1 (N14502, N14498);
or OR3 (N14503, N14492, N1697, N3323);
and AND3 (N14504, N14493, N5659, N10799);
nor NOR4 (N14505, N14500, N13879, N4209, N3604);
nor NOR2 (N14506, N14503, N7625);
not NOT1 (N14507, N14506);
not NOT1 (N14508, N14496);
nor NOR3 (N14509, N14502, N11722, N858);
or OR2 (N14510, N14507, N8332);
and AND3 (N14511, N14494, N7934, N481);
and AND3 (N14512, N14504, N10720, N2417);
not NOT1 (N14513, N14512);
and AND2 (N14514, N14501, N4719);
buf BUF1 (N14515, N14511);
not NOT1 (N14516, N14489);
nor NOR3 (N14517, N14514, N10378, N403);
nor NOR2 (N14518, N14513, N14230);
xor XOR2 (N14519, N14509, N4070);
xor XOR2 (N14520, N14510, N11090);
not NOT1 (N14521, N14495);
or OR2 (N14522, N14520, N12123);
buf BUF1 (N14523, N14508);
and AND4 (N14524, N14522, N9297, N4358, N4656);
xor XOR2 (N14525, N14517, N11650);
nand NAND3 (N14526, N14515, N7929, N330);
buf BUF1 (N14527, N14516);
or OR4 (N14528, N14499, N3328, N12341, N8841);
buf BUF1 (N14529, N14525);
not NOT1 (N14530, N14523);
nor NOR4 (N14531, N14518, N7288, N9744, N11864);
nand NAND2 (N14532, N14530, N9861);
not NOT1 (N14533, N14521);
nor NOR3 (N14534, N14529, N13472, N13750);
or OR4 (N14535, N14527, N268, N13336, N2275);
and AND3 (N14536, N14526, N11728, N7602);
nor NOR3 (N14537, N14528, N13591, N3677);
buf BUF1 (N14538, N14537);
xor XOR2 (N14539, N14536, N6557);
buf BUF1 (N14540, N14531);
nor NOR3 (N14541, N14539, N2031, N4137);
nor NOR3 (N14542, N14519, N9257, N10325);
nand NAND4 (N14543, N14541, N4277, N8435, N4666);
or OR2 (N14544, N14540, N5280);
nor NOR4 (N14545, N14543, N11733, N6476, N7700);
buf BUF1 (N14546, N14534);
buf BUF1 (N14547, N14542);
and AND4 (N14548, N14535, N3968, N9383, N1619);
nor NOR4 (N14549, N14524, N6900, N12899, N3782);
buf BUF1 (N14550, N14544);
not NOT1 (N14551, N14533);
and AND4 (N14552, N14505, N10778, N11038, N3191);
and AND4 (N14553, N14552, N10550, N5367, N11200);
not NOT1 (N14554, N14553);
not NOT1 (N14555, N14550);
nor NOR2 (N14556, N14548, N3857);
nor NOR3 (N14557, N14549, N5309, N13750);
buf BUF1 (N14558, N14532);
nand NAND2 (N14559, N14555, N8358);
and AND2 (N14560, N14546, N11880);
nand NAND3 (N14561, N14538, N5669, N2259);
nor NOR2 (N14562, N14561, N3942);
or OR4 (N14563, N14551, N1369, N456, N9035);
and AND4 (N14564, N14557, N10954, N2147, N1158);
or OR2 (N14565, N14545, N12869);
xor XOR2 (N14566, N14564, N6701);
nor NOR4 (N14567, N14556, N7670, N14353, N3548);
or OR2 (N14568, N14560, N14133);
xor XOR2 (N14569, N14566, N7416);
nor NOR3 (N14570, N14562, N5007, N3916);
nor NOR4 (N14571, N14570, N2244, N3614, N10917);
buf BUF1 (N14572, N14559);
buf BUF1 (N14573, N14569);
nor NOR2 (N14574, N14565, N11854);
nand NAND4 (N14575, N14571, N9346, N4629, N13799);
nand NAND3 (N14576, N14567, N14208, N5398);
nor NOR2 (N14577, N14573, N5465);
nor NOR3 (N14578, N14577, N14231, N9645);
nor NOR4 (N14579, N14574, N3997, N11897, N12689);
buf BUF1 (N14580, N14563);
and AND3 (N14581, N14558, N8631, N4228);
not NOT1 (N14582, N14581);
and AND3 (N14583, N14575, N9425, N5044);
not NOT1 (N14584, N14580);
buf BUF1 (N14585, N14554);
nand NAND4 (N14586, N14579, N7415, N9808, N12421);
nand NAND4 (N14587, N14586, N12333, N8991, N13582);
buf BUF1 (N14588, N14583);
nor NOR3 (N14589, N14547, N7396, N13005);
not NOT1 (N14590, N14589);
not NOT1 (N14591, N14578);
and AND3 (N14592, N14590, N13570, N12912);
or OR4 (N14593, N14582, N10710, N13679, N755);
buf BUF1 (N14594, N14584);
and AND3 (N14595, N14588, N14016, N11515);
xor XOR2 (N14596, N14594, N12987);
nor NOR3 (N14597, N14587, N5303, N11649);
xor XOR2 (N14598, N14572, N5027);
nand NAND2 (N14599, N14598, N14476);
nand NAND3 (N14600, N14585, N9035, N8837);
buf BUF1 (N14601, N14591);
buf BUF1 (N14602, N14595);
nor NOR3 (N14603, N14601, N6727, N12638);
xor XOR2 (N14604, N14576, N10619);
nor NOR4 (N14605, N14603, N11057, N9513, N9061);
buf BUF1 (N14606, N14596);
nor NOR3 (N14607, N14592, N3780, N782);
nor NOR2 (N14608, N14599, N8000);
xor XOR2 (N14609, N14604, N869);
nand NAND4 (N14610, N14597, N7743, N1788, N3627);
not NOT1 (N14611, N14610);
nor NOR4 (N14612, N14593, N9299, N7416, N11677);
or OR4 (N14613, N14611, N13769, N914, N13971);
xor XOR2 (N14614, N14606, N6183);
and AND3 (N14615, N14614, N7119, N696);
or OR2 (N14616, N14605, N2157);
not NOT1 (N14617, N14609);
not NOT1 (N14618, N14612);
xor XOR2 (N14619, N14607, N12647);
and AND4 (N14620, N14608, N11025, N5371, N5627);
or OR3 (N14621, N14602, N2038, N2185);
buf BUF1 (N14622, N14617);
nand NAND3 (N14623, N14600, N4315, N2124);
buf BUF1 (N14624, N14623);
xor XOR2 (N14625, N14620, N1766);
not NOT1 (N14626, N14616);
xor XOR2 (N14627, N14568, N5661);
and AND3 (N14628, N14619, N3387, N846);
and AND3 (N14629, N14613, N6375, N10153);
xor XOR2 (N14630, N14628, N8145);
nand NAND3 (N14631, N14630, N2620, N14454);
or OR4 (N14632, N14629, N9353, N11118, N10833);
or OR4 (N14633, N14631, N5365, N1591, N1378);
xor XOR2 (N14634, N14622, N4044);
and AND4 (N14635, N14627, N5000, N3084, N900);
xor XOR2 (N14636, N14632, N6932);
or OR4 (N14637, N14634, N4680, N3158, N2870);
nor NOR2 (N14638, N14624, N380);
nor NOR4 (N14639, N14633, N480, N10216, N7536);
xor XOR2 (N14640, N14618, N10467);
buf BUF1 (N14641, N14636);
not NOT1 (N14642, N14639);
or OR2 (N14643, N14637, N3628);
and AND3 (N14644, N14615, N13867, N11467);
buf BUF1 (N14645, N14644);
buf BUF1 (N14646, N14626);
buf BUF1 (N14647, N14641);
and AND4 (N14648, N14635, N3370, N2018, N7924);
xor XOR2 (N14649, N14642, N7201);
and AND3 (N14650, N14649, N9041, N8205);
not NOT1 (N14651, N14647);
not NOT1 (N14652, N14621);
and AND4 (N14653, N14643, N11592, N9940, N6379);
buf BUF1 (N14654, N14651);
xor XOR2 (N14655, N14654, N13439);
and AND4 (N14656, N14653, N10598, N7712, N7171);
and AND3 (N14657, N14645, N3368, N7788);
not NOT1 (N14658, N14656);
or OR2 (N14659, N14648, N7695);
or OR3 (N14660, N14640, N14131, N3397);
nand NAND3 (N14661, N14652, N14078, N6145);
and AND4 (N14662, N14625, N2209, N10549, N10427);
and AND2 (N14663, N14646, N104);
nor NOR3 (N14664, N14662, N5904, N14497);
buf BUF1 (N14665, N14650);
and AND3 (N14666, N14655, N4562, N8835);
and AND3 (N14667, N14657, N7437, N555);
and AND2 (N14668, N14659, N1032);
nand NAND2 (N14669, N14661, N7716);
not NOT1 (N14670, N14668);
or OR4 (N14671, N14665, N1835, N4337, N14127);
nand NAND3 (N14672, N14666, N7653, N8103);
nand NAND2 (N14673, N14667, N5286);
xor XOR2 (N14674, N14664, N7187);
buf BUF1 (N14675, N14669);
and AND4 (N14676, N14675, N1581, N5205, N2912);
or OR2 (N14677, N14671, N4685);
nor NOR4 (N14678, N14660, N400, N7272, N9807);
and AND4 (N14679, N14663, N9127, N1713, N11634);
not NOT1 (N14680, N14676);
xor XOR2 (N14681, N14680, N11909);
nor NOR3 (N14682, N14678, N6384, N4702);
not NOT1 (N14683, N14658);
not NOT1 (N14684, N14674);
and AND2 (N14685, N14684, N10382);
nor NOR4 (N14686, N14681, N7909, N7161, N10936);
and AND3 (N14687, N14638, N10656, N3088);
buf BUF1 (N14688, N14672);
buf BUF1 (N14689, N14679);
or OR4 (N14690, N14677, N1182, N8188, N8406);
nand NAND4 (N14691, N14686, N6854, N5509, N585);
and AND3 (N14692, N14688, N7103, N8286);
not NOT1 (N14693, N14689);
nand NAND3 (N14694, N14693, N5937, N13793);
xor XOR2 (N14695, N14673, N6867);
not NOT1 (N14696, N14695);
or OR3 (N14697, N14670, N2106, N3965);
buf BUF1 (N14698, N14692);
xor XOR2 (N14699, N14696, N1749);
buf BUF1 (N14700, N14697);
or OR3 (N14701, N14700, N8350, N14592);
not NOT1 (N14702, N14690);
buf BUF1 (N14703, N14682);
or OR4 (N14704, N14683, N2158, N1786, N13588);
xor XOR2 (N14705, N14698, N2731);
not NOT1 (N14706, N14701);
nand NAND2 (N14707, N14703, N4392);
nand NAND3 (N14708, N14691, N9083, N2702);
nor NOR3 (N14709, N14706, N7642, N9398);
not NOT1 (N14710, N14702);
nand NAND3 (N14711, N14705, N8742, N932);
and AND4 (N14712, N14694, N318, N12559, N5988);
xor XOR2 (N14713, N14704, N12982);
and AND2 (N14714, N14709, N11171);
and AND4 (N14715, N14712, N12648, N11753, N9038);
not NOT1 (N14716, N14713);
nor NOR2 (N14717, N14687, N5587);
xor XOR2 (N14718, N14715, N7114);
nand NAND2 (N14719, N14707, N12025);
xor XOR2 (N14720, N14710, N1845);
xor XOR2 (N14721, N14714, N13920);
and AND4 (N14722, N14716, N5732, N12546, N12227);
nand NAND2 (N14723, N14699, N4334);
or OR3 (N14724, N14721, N7241, N12227);
buf BUF1 (N14725, N14722);
and AND4 (N14726, N14718, N2365, N10709, N5332);
xor XOR2 (N14727, N14685, N2080);
nor NOR4 (N14728, N14711, N3070, N1910, N2359);
and AND3 (N14729, N14719, N11628, N14092);
xor XOR2 (N14730, N14729, N4195);
nor NOR3 (N14731, N14726, N5317, N1312);
nand NAND3 (N14732, N14730, N8521, N13091);
buf BUF1 (N14733, N14724);
nand NAND4 (N14734, N14732, N4526, N14257, N9815);
and AND2 (N14735, N14725, N7007);
nor NOR3 (N14736, N14708, N1133, N5089);
not NOT1 (N14737, N14720);
not NOT1 (N14738, N14728);
nor NOR4 (N14739, N14733, N11234, N6472, N10774);
buf BUF1 (N14740, N14737);
and AND3 (N14741, N14727, N4300, N1500);
not NOT1 (N14742, N14740);
xor XOR2 (N14743, N14734, N1022);
xor XOR2 (N14744, N14731, N8941);
and AND4 (N14745, N14736, N8462, N12310, N14328);
not NOT1 (N14746, N14735);
buf BUF1 (N14747, N14739);
buf BUF1 (N14748, N14744);
nor NOR4 (N14749, N14743, N3621, N338, N8488);
xor XOR2 (N14750, N14746, N841);
buf BUF1 (N14751, N14748);
or OR3 (N14752, N14751, N1528, N8051);
nand NAND3 (N14753, N14747, N4110, N231);
nand NAND3 (N14754, N14749, N983, N720);
xor XOR2 (N14755, N14738, N8348);
nand NAND2 (N14756, N14745, N13637);
and AND4 (N14757, N14753, N9764, N12274, N2499);
or OR3 (N14758, N14755, N6653, N10113);
and AND2 (N14759, N14717, N3968);
buf BUF1 (N14760, N14758);
or OR4 (N14761, N14757, N9198, N5884, N6753);
not NOT1 (N14762, N14752);
xor XOR2 (N14763, N14761, N14055);
or OR3 (N14764, N14760, N3105, N4525);
and AND4 (N14765, N14741, N1709, N9770, N11630);
or OR3 (N14766, N14742, N1394, N8357);
nand NAND2 (N14767, N14764, N6260);
and AND3 (N14768, N14756, N11036, N6915);
and AND3 (N14769, N14766, N73, N8483);
nand NAND2 (N14770, N14759, N4230);
and AND4 (N14771, N14754, N1957, N11582, N10675);
and AND2 (N14772, N14762, N10645);
and AND2 (N14773, N14769, N6895);
nor NOR2 (N14774, N14770, N5372);
nand NAND3 (N14775, N14767, N8250, N13876);
not NOT1 (N14776, N14763);
not NOT1 (N14777, N14765);
not NOT1 (N14778, N14750);
and AND4 (N14779, N14768, N9242, N8239, N7421);
nand NAND3 (N14780, N14774, N3197, N13238);
nor NOR4 (N14781, N14777, N212, N1314, N3791);
nor NOR4 (N14782, N14723, N11606, N12367, N7101);
xor XOR2 (N14783, N14772, N3304);
nor NOR3 (N14784, N14781, N9675, N9694);
not NOT1 (N14785, N14780);
or OR4 (N14786, N14776, N6608, N9639, N14544);
or OR4 (N14787, N14782, N4061, N6726, N4211);
nand NAND3 (N14788, N14775, N3348, N7920);
buf BUF1 (N14789, N14788);
xor XOR2 (N14790, N14771, N6958);
not NOT1 (N14791, N14779);
xor XOR2 (N14792, N14791, N7292);
nor NOR3 (N14793, N14787, N1855, N8015);
nor NOR3 (N14794, N14783, N4486, N908);
nand NAND4 (N14795, N14773, N7145, N2616, N6669);
xor XOR2 (N14796, N14785, N3459);
or OR4 (N14797, N14790, N3220, N8894, N7259);
buf BUF1 (N14798, N14796);
nor NOR2 (N14799, N14795, N151);
buf BUF1 (N14800, N14792);
xor XOR2 (N14801, N14784, N4513);
or OR3 (N14802, N14778, N8011, N1042);
xor XOR2 (N14803, N14800, N2890);
and AND3 (N14804, N14786, N4430, N13503);
nor NOR2 (N14805, N14789, N8587);
and AND2 (N14806, N14802, N14626);
and AND3 (N14807, N14805, N1711, N6438);
not NOT1 (N14808, N14797);
xor XOR2 (N14809, N14808, N2240);
buf BUF1 (N14810, N14809);
not NOT1 (N14811, N14803);
not NOT1 (N14812, N14794);
and AND3 (N14813, N14798, N3699, N13741);
xor XOR2 (N14814, N14807, N9042);
nor NOR2 (N14815, N14813, N1901);
not NOT1 (N14816, N14799);
not NOT1 (N14817, N14793);
buf BUF1 (N14818, N14811);
nor NOR4 (N14819, N14817, N10229, N12398, N11754);
buf BUF1 (N14820, N14806);
and AND4 (N14821, N14819, N6130, N1746, N10681);
xor XOR2 (N14822, N14816, N10809);
buf BUF1 (N14823, N14814);
xor XOR2 (N14824, N14801, N13256);
nand NAND2 (N14825, N14823, N3167);
nor NOR4 (N14826, N14812, N6491, N12977, N8051);
nor NOR2 (N14827, N14826, N14249);
or OR2 (N14828, N14824, N12675);
nor NOR4 (N14829, N14820, N786, N7430, N4573);
buf BUF1 (N14830, N14810);
and AND2 (N14831, N14827, N2644);
xor XOR2 (N14832, N14828, N8391);
not NOT1 (N14833, N14825);
nand NAND2 (N14834, N14831, N12681);
or OR2 (N14835, N14822, N1885);
xor XOR2 (N14836, N14834, N11000);
or OR2 (N14837, N14829, N12702);
and AND3 (N14838, N14832, N2018, N13174);
xor XOR2 (N14839, N14830, N2361);
not NOT1 (N14840, N14818);
and AND3 (N14841, N14835, N7408, N12490);
nor NOR4 (N14842, N14833, N13938, N7597, N7390);
nor NOR3 (N14843, N14842, N454, N7588);
or OR2 (N14844, N14839, N2227);
nor NOR3 (N14845, N14821, N14524, N85);
nand NAND3 (N14846, N14804, N7042, N912);
buf BUF1 (N14847, N14841);
or OR2 (N14848, N14836, N4385);
not NOT1 (N14849, N14840);
buf BUF1 (N14850, N14815);
or OR3 (N14851, N14837, N1442, N10496);
xor XOR2 (N14852, N14843, N10544);
nor NOR3 (N14853, N14849, N9218, N14349);
xor XOR2 (N14854, N14838, N433);
not NOT1 (N14855, N14851);
not NOT1 (N14856, N14844);
not NOT1 (N14857, N14855);
not NOT1 (N14858, N14846);
buf BUF1 (N14859, N14852);
nor NOR2 (N14860, N14850, N10699);
nand NAND3 (N14861, N14848, N9921, N3627);
xor XOR2 (N14862, N14853, N4099);
not NOT1 (N14863, N14857);
nor NOR4 (N14864, N14845, N4231, N5193, N6762);
and AND4 (N14865, N14854, N6686, N10158, N2477);
buf BUF1 (N14866, N14861);
nand NAND2 (N14867, N14847, N13639);
buf BUF1 (N14868, N14865);
buf BUF1 (N14869, N14864);
nand NAND4 (N14870, N14860, N6572, N1081, N714);
xor XOR2 (N14871, N14863, N3154);
nor NOR4 (N14872, N14858, N8735, N11199, N8286);
nor NOR2 (N14873, N14856, N9771);
and AND4 (N14874, N14868, N3239, N4910, N9397);
and AND2 (N14875, N14873, N1599);
nand NAND2 (N14876, N14867, N3030);
and AND3 (N14877, N14862, N6753, N2713);
nand NAND2 (N14878, N14871, N10165);
xor XOR2 (N14879, N14859, N869);
and AND2 (N14880, N14877, N11107);
or OR3 (N14881, N14874, N12436, N4675);
buf BUF1 (N14882, N14875);
nand NAND4 (N14883, N14880, N10631, N6957, N8289);
xor XOR2 (N14884, N14869, N5856);
not NOT1 (N14885, N14878);
xor XOR2 (N14886, N14885, N13830);
nor NOR4 (N14887, N14876, N1156, N4151, N4916);
and AND2 (N14888, N14887, N12557);
xor XOR2 (N14889, N14881, N8127);
xor XOR2 (N14890, N14872, N14252);
buf BUF1 (N14891, N14890);
or OR2 (N14892, N14891, N5513);
nor NOR3 (N14893, N14889, N13714, N845);
not NOT1 (N14894, N14870);
not NOT1 (N14895, N14884);
nand NAND3 (N14896, N14886, N9975, N53);
nand NAND4 (N14897, N14895, N7660, N7820, N13722);
or OR3 (N14898, N14897, N14861, N8166);
and AND4 (N14899, N14882, N9333, N3923, N127);
nor NOR4 (N14900, N14879, N12144, N6790, N1879);
and AND4 (N14901, N14893, N14024, N1248, N3226);
and AND4 (N14902, N14883, N13318, N5858, N10905);
and AND3 (N14903, N14898, N4382, N8030);
not NOT1 (N14904, N14892);
nor NOR4 (N14905, N14899, N2336, N6284, N1259);
nor NOR3 (N14906, N14896, N14209, N348);
not NOT1 (N14907, N14904);
nor NOR3 (N14908, N14866, N8245, N14444);
buf BUF1 (N14909, N14905);
or OR2 (N14910, N14908, N10891);
buf BUF1 (N14911, N14888);
not NOT1 (N14912, N14910);
buf BUF1 (N14913, N14907);
nand NAND2 (N14914, N14902, N7605);
nand NAND2 (N14915, N14900, N14284);
or OR4 (N14916, N14894, N12703, N8789, N8132);
nand NAND2 (N14917, N14906, N14698);
xor XOR2 (N14918, N14914, N13263);
nand NAND3 (N14919, N14911, N1225, N12991);
buf BUF1 (N14920, N14917);
nand NAND3 (N14921, N14913, N4672, N4666);
xor XOR2 (N14922, N14920, N9922);
not NOT1 (N14923, N14916);
and AND2 (N14924, N14909, N14338);
and AND2 (N14925, N14923, N9759);
xor XOR2 (N14926, N14921, N3998);
nand NAND2 (N14927, N14912, N1135);
xor XOR2 (N14928, N14903, N4399);
not NOT1 (N14929, N14924);
buf BUF1 (N14930, N14901);
buf BUF1 (N14931, N14925);
nand NAND2 (N14932, N14922, N13408);
or OR4 (N14933, N14918, N10574, N7157, N4422);
buf BUF1 (N14934, N14915);
xor XOR2 (N14935, N14926, N3643);
nand NAND2 (N14936, N14928, N10552);
and AND2 (N14937, N14929, N13806);
nor NOR4 (N14938, N14933, N12167, N10627, N2295);
nand NAND3 (N14939, N14927, N3489, N4478);
xor XOR2 (N14940, N14930, N6699);
buf BUF1 (N14941, N14932);
nor NOR3 (N14942, N14937, N9013, N13411);
buf BUF1 (N14943, N14919);
or OR2 (N14944, N14936, N9945);
and AND2 (N14945, N14931, N8303);
and AND4 (N14946, N14945, N2486, N761, N3824);
nor NOR3 (N14947, N14939, N14862, N11681);
nand NAND2 (N14948, N14934, N14774);
nand NAND3 (N14949, N14944, N3595, N10588);
or OR3 (N14950, N14949, N6792, N3827);
buf BUF1 (N14951, N14941);
nor NOR4 (N14952, N14948, N13928, N13200, N14559);
xor XOR2 (N14953, N14950, N6389);
nand NAND3 (N14954, N14952, N12550, N797);
nor NOR3 (N14955, N14946, N4141, N9844);
buf BUF1 (N14956, N14955);
nor NOR4 (N14957, N14942, N1438, N13941, N11113);
or OR4 (N14958, N14943, N6628, N8839, N14555);
or OR3 (N14959, N14947, N13781, N7345);
nand NAND4 (N14960, N14940, N1608, N3052, N1965);
buf BUF1 (N14961, N14959);
not NOT1 (N14962, N14935);
nor NOR4 (N14963, N14960, N3914, N13585, N6900);
and AND4 (N14964, N14954, N2875, N2331, N4624);
nand NAND2 (N14965, N14961, N5348);
buf BUF1 (N14966, N14963);
and AND2 (N14967, N14951, N6389);
not NOT1 (N14968, N14953);
nand NAND4 (N14969, N14967, N13717, N6222, N12426);
nand NAND3 (N14970, N14938, N6281, N10054);
xor XOR2 (N14971, N14964, N13676);
not NOT1 (N14972, N14962);
and AND3 (N14973, N14965, N4116, N10929);
or OR4 (N14974, N14973, N14151, N4305, N11796);
nand NAND3 (N14975, N14972, N7869, N8426);
or OR2 (N14976, N14957, N12061);
not NOT1 (N14977, N14968);
buf BUF1 (N14978, N14969);
nand NAND2 (N14979, N14974, N13825);
xor XOR2 (N14980, N14975, N7238);
xor XOR2 (N14981, N14970, N14961);
and AND3 (N14982, N14958, N3056, N5396);
nor NOR2 (N14983, N14977, N11249);
xor XOR2 (N14984, N14980, N802);
not NOT1 (N14985, N14971);
and AND4 (N14986, N14978, N5175, N3175, N1821);
or OR4 (N14987, N14966, N7818, N2085, N12586);
xor XOR2 (N14988, N14979, N10912);
or OR2 (N14989, N14987, N12065);
or OR3 (N14990, N14982, N6671, N2365);
or OR2 (N14991, N14976, N9970);
or OR4 (N14992, N14984, N10877, N2826, N278);
xor XOR2 (N14993, N14986, N14263);
xor XOR2 (N14994, N14988, N8870);
nand NAND2 (N14995, N14985, N13024);
not NOT1 (N14996, N14990);
buf BUF1 (N14997, N14956);
not NOT1 (N14998, N14996);
nor NOR4 (N14999, N14997, N11676, N10313, N5560);
nor NOR3 (N15000, N14993, N13996, N13809);
nand NAND4 (N15001, N14995, N12193, N10625, N14205);
nor NOR3 (N15002, N14998, N9546, N13808);
not NOT1 (N15003, N14983);
and AND4 (N15004, N14991, N3689, N12681, N7994);
nor NOR2 (N15005, N15000, N6972);
xor XOR2 (N15006, N15003, N6873);
buf BUF1 (N15007, N15005);
xor XOR2 (N15008, N15007, N4396);
nand NAND3 (N15009, N15004, N13176, N1708);
nand NAND4 (N15010, N15008, N3126, N1896, N2927);
buf BUF1 (N15011, N15001);
or OR4 (N15012, N14992, N6914, N14889, N9424);
not NOT1 (N15013, N14981);
buf BUF1 (N15014, N14989);
nand NAND3 (N15015, N15013, N10254, N1349);
nor NOR3 (N15016, N15006, N9175, N7011);
buf BUF1 (N15017, N15012);
not NOT1 (N15018, N15015);
xor XOR2 (N15019, N15010, N13321);
xor XOR2 (N15020, N15016, N1762);
and AND3 (N15021, N15019, N10805, N7090);
buf BUF1 (N15022, N15017);
nor NOR3 (N15023, N15020, N4857, N8600);
and AND4 (N15024, N15023, N10106, N268, N7518);
buf BUF1 (N15025, N15021);
xor XOR2 (N15026, N15002, N9381);
not NOT1 (N15027, N15022);
buf BUF1 (N15028, N14999);
not NOT1 (N15029, N15026);
nand NAND4 (N15030, N15028, N705, N2310, N13974);
buf BUF1 (N15031, N15029);
nand NAND4 (N15032, N15014, N10305, N1989, N7691);
not NOT1 (N15033, N14994);
nand NAND2 (N15034, N15027, N12797);
not NOT1 (N15035, N15030);
buf BUF1 (N15036, N15018);
buf BUF1 (N15037, N15033);
xor XOR2 (N15038, N15034, N10670);
and AND3 (N15039, N15025, N13030, N7116);
xor XOR2 (N15040, N15036, N3554);
or OR2 (N15041, N15009, N3763);
nor NOR4 (N15042, N15041, N8864, N2093, N8927);
nor NOR3 (N15043, N15035, N267, N5744);
nor NOR3 (N15044, N15011, N7878, N13163);
nand NAND3 (N15045, N15043, N5387, N3817);
buf BUF1 (N15046, N15031);
buf BUF1 (N15047, N15037);
buf BUF1 (N15048, N15040);
or OR2 (N15049, N15038, N4333);
nor NOR2 (N15050, N15049, N8080);
xor XOR2 (N15051, N15050, N11299);
not NOT1 (N15052, N15047);
buf BUF1 (N15053, N15048);
buf BUF1 (N15054, N15051);
buf BUF1 (N15055, N15045);
or OR3 (N15056, N15052, N10353, N8903);
nor NOR4 (N15057, N15046, N920, N12725, N4505);
nor NOR2 (N15058, N15044, N2772);
xor XOR2 (N15059, N15055, N784);
not NOT1 (N15060, N15057);
buf BUF1 (N15061, N15024);
buf BUF1 (N15062, N15032);
or OR2 (N15063, N15062, N9997);
nand NAND4 (N15064, N15059, N5058, N4760, N14642);
buf BUF1 (N15065, N15042);
nand NAND2 (N15066, N15039, N797);
nand NAND4 (N15067, N15066, N3672, N4911, N6364);
and AND4 (N15068, N15053, N11853, N6517, N10017);
and AND2 (N15069, N15068, N362);
nand NAND3 (N15070, N15065, N13317, N6985);
not NOT1 (N15071, N15056);
nand NAND3 (N15072, N15061, N10073, N13233);
nand NAND3 (N15073, N15064, N2659, N874);
nor NOR2 (N15074, N15073, N13350);
nor NOR4 (N15075, N15071, N2172, N7653, N14048);
and AND4 (N15076, N15060, N4613, N7165, N588);
and AND4 (N15077, N15058, N7555, N10102, N198);
not NOT1 (N15078, N15077);
and AND3 (N15079, N15067, N4596, N11631);
nor NOR2 (N15080, N15079, N5817);
nand NAND3 (N15081, N15069, N2439, N7357);
or OR4 (N15082, N15072, N9265, N12620, N6213);
nand NAND4 (N15083, N15081, N11775, N3334, N240);
nor NOR4 (N15084, N15075, N9993, N9174, N8958);
nor NOR4 (N15085, N15063, N598, N1665, N13968);
and AND2 (N15086, N15070, N866);
nor NOR2 (N15087, N15076, N5808);
nand NAND4 (N15088, N15080, N1151, N11196, N10749);
xor XOR2 (N15089, N15082, N1005);
xor XOR2 (N15090, N15083, N8204);
xor XOR2 (N15091, N15086, N8079);
not NOT1 (N15092, N15078);
or OR3 (N15093, N15091, N13822, N4275);
nand NAND4 (N15094, N15087, N9623, N13897, N2454);
and AND2 (N15095, N15092, N8618);
or OR3 (N15096, N15090, N705, N9767);
nand NAND4 (N15097, N15054, N3959, N6516, N5951);
not NOT1 (N15098, N15088);
xor XOR2 (N15099, N15098, N8575);
not NOT1 (N15100, N15095);
not NOT1 (N15101, N15094);
or OR2 (N15102, N15096, N415);
nand NAND4 (N15103, N15074, N11595, N3212, N10793);
nand NAND3 (N15104, N15084, N11032, N9990);
not NOT1 (N15105, N15104);
nand NAND4 (N15106, N15103, N7006, N13648, N14972);
buf BUF1 (N15107, N15101);
nand NAND4 (N15108, N15093, N11279, N11965, N12767);
not NOT1 (N15109, N15097);
buf BUF1 (N15110, N15108);
not NOT1 (N15111, N15107);
buf BUF1 (N15112, N15089);
nand NAND3 (N15113, N15105, N8070, N5908);
nand NAND2 (N15114, N15085, N8714);
nor NOR4 (N15115, N15099, N5669, N14472, N10500);
and AND2 (N15116, N15112, N7099);
and AND3 (N15117, N15115, N4176, N5952);
not NOT1 (N15118, N15110);
nand NAND2 (N15119, N15100, N5989);
or OR2 (N15120, N15109, N3725);
xor XOR2 (N15121, N15102, N871);
and AND4 (N15122, N15106, N5288, N7616, N889);
nor NOR4 (N15123, N15117, N9938, N4706, N10465);
nand NAND3 (N15124, N15114, N10889, N7992);
not NOT1 (N15125, N15118);
buf BUF1 (N15126, N15119);
or OR4 (N15127, N15116, N12679, N3482, N3798);
xor XOR2 (N15128, N15124, N1155);
or OR2 (N15129, N15127, N12649);
nand NAND3 (N15130, N15120, N2043, N1656);
nor NOR2 (N15131, N15123, N12311);
nand NAND3 (N15132, N15128, N321, N6431);
nand NAND3 (N15133, N15121, N8950, N7135);
nand NAND4 (N15134, N15129, N11349, N13033, N3071);
buf BUF1 (N15135, N15130);
and AND4 (N15136, N15125, N5437, N14919, N1991);
buf BUF1 (N15137, N15135);
nand NAND2 (N15138, N15113, N13884);
nand NAND3 (N15139, N15138, N6098, N14939);
xor XOR2 (N15140, N15136, N3441);
not NOT1 (N15141, N15137);
and AND4 (N15142, N15141, N11684, N2875, N11853);
buf BUF1 (N15143, N15122);
buf BUF1 (N15144, N15111);
not NOT1 (N15145, N15144);
buf BUF1 (N15146, N15145);
nor NOR4 (N15147, N15143, N7962, N7920, N7505);
nor NOR3 (N15148, N15126, N11131, N5784);
not NOT1 (N15149, N15140);
nand NAND2 (N15150, N15148, N7119);
xor XOR2 (N15151, N15142, N10588);
not NOT1 (N15152, N15139);
nand NAND4 (N15153, N15134, N5378, N9341, N12602);
xor XOR2 (N15154, N15133, N3708);
and AND2 (N15155, N15150, N13696);
or OR4 (N15156, N15154, N9966, N5908, N10271);
buf BUF1 (N15157, N15147);
not NOT1 (N15158, N15153);
xor XOR2 (N15159, N15156, N6117);
nor NOR2 (N15160, N15151, N13105);
and AND4 (N15161, N15159, N7269, N7008, N13010);
and AND2 (N15162, N15152, N9157);
buf BUF1 (N15163, N15157);
and AND4 (N15164, N15160, N15006, N12084, N3583);
not NOT1 (N15165, N15149);
or OR4 (N15166, N15131, N452, N1008, N14201);
buf BUF1 (N15167, N15161);
or OR4 (N15168, N15146, N15036, N9822, N10353);
buf BUF1 (N15169, N15162);
and AND4 (N15170, N15155, N10755, N10915, N3077);
nand NAND2 (N15171, N15158, N14610);
xor XOR2 (N15172, N15168, N1685);
or OR4 (N15173, N15163, N12780, N12904, N14188);
or OR3 (N15174, N15172, N10019, N11128);
or OR4 (N15175, N15174, N11040, N8155, N10281);
nand NAND4 (N15176, N15175, N980, N1148, N9622);
xor XOR2 (N15177, N15164, N687);
nand NAND4 (N15178, N15167, N11455, N12250, N1307);
nor NOR4 (N15179, N15132, N4985, N2046, N5724);
and AND2 (N15180, N15177, N6497);
or OR2 (N15181, N15170, N6097);
nor NOR3 (N15182, N15178, N4055, N12442);
xor XOR2 (N15183, N15165, N2502);
buf BUF1 (N15184, N15171);
xor XOR2 (N15185, N15183, N983);
xor XOR2 (N15186, N15180, N9803);
or OR3 (N15187, N15176, N7250, N13303);
nor NOR4 (N15188, N15173, N4428, N2215, N6849);
not NOT1 (N15189, N15184);
and AND3 (N15190, N15189, N10401, N4312);
not NOT1 (N15191, N15166);
buf BUF1 (N15192, N15181);
xor XOR2 (N15193, N15191, N7694);
and AND2 (N15194, N15182, N7360);
or OR2 (N15195, N15192, N5523);
nand NAND3 (N15196, N15185, N8864, N11998);
buf BUF1 (N15197, N15188);
xor XOR2 (N15198, N15193, N5469);
or OR4 (N15199, N15187, N3547, N11374, N6783);
and AND2 (N15200, N15199, N9240);
nor NOR3 (N15201, N15196, N5340, N9493);
nand NAND4 (N15202, N15194, N5495, N3479, N4525);
nor NOR3 (N15203, N15186, N14518, N5905);
xor XOR2 (N15204, N15198, N10048);
xor XOR2 (N15205, N15201, N1882);
not NOT1 (N15206, N15203);
nand NAND2 (N15207, N15204, N3144);
nand NAND3 (N15208, N15205, N1850, N435);
nor NOR2 (N15209, N15208, N12489);
or OR2 (N15210, N15209, N2614);
or OR2 (N15211, N15207, N4612);
not NOT1 (N15212, N15195);
or OR2 (N15213, N15179, N5780);
or OR4 (N15214, N15202, N12262, N12304, N14283);
or OR3 (N15215, N15213, N10938, N11293);
not NOT1 (N15216, N15206);
nor NOR2 (N15217, N15190, N9428);
and AND2 (N15218, N15215, N14064);
not NOT1 (N15219, N15169);
xor XOR2 (N15220, N15216, N4185);
nor NOR2 (N15221, N15217, N4839);
nand NAND4 (N15222, N15211, N8165, N7246, N7829);
nand NAND2 (N15223, N15210, N6409);
not NOT1 (N15224, N15212);
xor XOR2 (N15225, N15214, N3107);
and AND4 (N15226, N15218, N545, N13209, N4255);
buf BUF1 (N15227, N15223);
xor XOR2 (N15228, N15220, N3556);
nand NAND4 (N15229, N15227, N2732, N3989, N6740);
or OR2 (N15230, N15197, N11473);
or OR4 (N15231, N15226, N806, N13458, N11787);
xor XOR2 (N15232, N15230, N3485);
xor XOR2 (N15233, N15224, N12871);
or OR2 (N15234, N15229, N2962);
buf BUF1 (N15235, N15222);
xor XOR2 (N15236, N15219, N4728);
and AND3 (N15237, N15225, N10567, N4402);
or OR3 (N15238, N15237, N6804, N9952);
or OR2 (N15239, N15232, N6717);
xor XOR2 (N15240, N15234, N3332);
and AND3 (N15241, N15221, N14545, N6260);
nor NOR2 (N15242, N15235, N9254);
not NOT1 (N15243, N15228);
nor NOR4 (N15244, N15233, N15131, N2444, N7870);
not NOT1 (N15245, N15241);
buf BUF1 (N15246, N15243);
buf BUF1 (N15247, N15231);
and AND2 (N15248, N15240, N2158);
nand NAND4 (N15249, N15246, N10428, N13157, N3881);
buf BUF1 (N15250, N15236);
nor NOR4 (N15251, N15239, N1906, N5547, N15182);
not NOT1 (N15252, N15247);
nor NOR3 (N15253, N15238, N12266, N3581);
buf BUF1 (N15254, N15245);
buf BUF1 (N15255, N15252);
or OR2 (N15256, N15250, N15043);
buf BUF1 (N15257, N15200);
xor XOR2 (N15258, N15242, N14855);
not NOT1 (N15259, N15251);
nand NAND4 (N15260, N15256, N12272, N1180, N1023);
and AND4 (N15261, N15258, N4954, N9236, N8735);
nor NOR4 (N15262, N15255, N2128, N9985, N13529);
or OR2 (N15263, N15257, N3855);
or OR2 (N15264, N15259, N9269);
and AND3 (N15265, N15253, N2154, N14397);
nor NOR2 (N15266, N15249, N3687);
or OR2 (N15267, N15266, N14535);
xor XOR2 (N15268, N15260, N1836);
and AND4 (N15269, N15268, N13034, N10555, N4424);
nand NAND2 (N15270, N15261, N2372);
buf BUF1 (N15271, N15254);
not NOT1 (N15272, N15269);
buf BUF1 (N15273, N15263);
buf BUF1 (N15274, N15267);
nand NAND3 (N15275, N15272, N8291, N8893);
xor XOR2 (N15276, N15248, N9134);
not NOT1 (N15277, N15271);
not NOT1 (N15278, N15276);
or OR2 (N15279, N15277, N9954);
nor NOR4 (N15280, N15273, N14070, N10132, N8293);
or OR2 (N15281, N15264, N2567);
buf BUF1 (N15282, N15270);
xor XOR2 (N15283, N15280, N10001);
xor XOR2 (N15284, N15278, N5678);
and AND4 (N15285, N15281, N1335, N5709, N7058);
nor NOR3 (N15286, N15265, N7024, N3535);
nor NOR2 (N15287, N15283, N2961);
nor NOR4 (N15288, N15274, N14411, N12873, N7486);
nand NAND2 (N15289, N15288, N3738);
buf BUF1 (N15290, N15275);
and AND3 (N15291, N15289, N10757, N1577);
nand NAND4 (N15292, N15286, N1330, N10542, N9848);
buf BUF1 (N15293, N15262);
or OR2 (N15294, N15290, N528);
and AND2 (N15295, N15284, N13101);
or OR2 (N15296, N15285, N12125);
nor NOR2 (N15297, N15294, N3206);
nand NAND4 (N15298, N15293, N8945, N4142, N14547);
nand NAND4 (N15299, N15282, N8196, N11249, N4305);
buf BUF1 (N15300, N15279);
xor XOR2 (N15301, N15291, N5803);
or OR4 (N15302, N15292, N4741, N119, N12441);
buf BUF1 (N15303, N15302);
nand NAND3 (N15304, N15295, N8143, N7249);
nand NAND3 (N15305, N15297, N14830, N5984);
buf BUF1 (N15306, N15299);
nand NAND2 (N15307, N15304, N1091);
xor XOR2 (N15308, N15305, N11485);
not NOT1 (N15309, N15306);
not NOT1 (N15310, N15303);
nor NOR2 (N15311, N15287, N8138);
buf BUF1 (N15312, N15301);
xor XOR2 (N15313, N15310, N5667);
buf BUF1 (N15314, N15244);
not NOT1 (N15315, N15311);
not NOT1 (N15316, N15298);
buf BUF1 (N15317, N15309);
not NOT1 (N15318, N15313);
and AND3 (N15319, N15312, N14054, N15101);
nor NOR2 (N15320, N15319, N14503);
xor XOR2 (N15321, N15300, N7613);
not NOT1 (N15322, N15321);
nand NAND4 (N15323, N15322, N6533, N11514, N7236);
buf BUF1 (N15324, N15317);
or OR4 (N15325, N15324, N9573, N9134, N11377);
and AND3 (N15326, N15325, N8377, N10312);
and AND2 (N15327, N15326, N11751);
nand NAND2 (N15328, N15320, N8965);
nand NAND4 (N15329, N15314, N4361, N5494, N11507);
not NOT1 (N15330, N15316);
or OR3 (N15331, N15296, N732, N13190);
or OR3 (N15332, N15318, N13614, N4820);
nand NAND3 (N15333, N15328, N13862, N2279);
nor NOR2 (N15334, N15332, N5495);
buf BUF1 (N15335, N15323);
buf BUF1 (N15336, N15334);
and AND3 (N15337, N15329, N5448, N9992);
or OR3 (N15338, N15335, N13101, N10923);
and AND2 (N15339, N15336, N12703);
buf BUF1 (N15340, N15333);
or OR2 (N15341, N15307, N5830);
and AND3 (N15342, N15308, N4350, N14754);
not NOT1 (N15343, N15327);
nand NAND3 (N15344, N15338, N14382, N3204);
not NOT1 (N15345, N15340);
buf BUF1 (N15346, N15339);
buf BUF1 (N15347, N15346);
and AND3 (N15348, N15342, N4475, N1260);
nand NAND2 (N15349, N15345, N10685);
xor XOR2 (N15350, N15348, N1668);
nor NOR4 (N15351, N15341, N6397, N12741, N3733);
buf BUF1 (N15352, N15337);
xor XOR2 (N15353, N15347, N539);
not NOT1 (N15354, N15343);
or OR3 (N15355, N15353, N3547, N2653);
buf BUF1 (N15356, N15331);
xor XOR2 (N15357, N15355, N5553);
nand NAND4 (N15358, N15315, N4799, N5647, N10658);
nand NAND2 (N15359, N15351, N8152);
not NOT1 (N15360, N15354);
nand NAND4 (N15361, N15357, N6414, N12947, N612);
xor XOR2 (N15362, N15356, N9126);
and AND3 (N15363, N15360, N14837, N8572);
buf BUF1 (N15364, N15350);
and AND2 (N15365, N15330, N7253);
nand NAND4 (N15366, N15365, N2941, N9804, N2154);
or OR3 (N15367, N15362, N1280, N10159);
or OR4 (N15368, N15361, N4723, N9722, N5898);
buf BUF1 (N15369, N15358);
nor NOR4 (N15370, N15364, N12830, N10515, N1501);
xor XOR2 (N15371, N15352, N13629);
not NOT1 (N15372, N15344);
nor NOR2 (N15373, N15349, N11782);
not NOT1 (N15374, N15373);
and AND4 (N15375, N15374, N3019, N10721, N12341);
xor XOR2 (N15376, N15368, N1621);
buf BUF1 (N15377, N15370);
xor XOR2 (N15378, N15366, N2452);
buf BUF1 (N15379, N15363);
buf BUF1 (N15380, N15372);
xor XOR2 (N15381, N15371, N5114);
buf BUF1 (N15382, N15379);
nor NOR2 (N15383, N15369, N4820);
nand NAND2 (N15384, N15359, N2736);
nor NOR3 (N15385, N15380, N7774, N298);
nor NOR2 (N15386, N15383, N1802);
nand NAND4 (N15387, N15377, N11289, N12580, N8500);
buf BUF1 (N15388, N15387);
nand NAND3 (N15389, N15376, N1854, N15003);
nor NOR4 (N15390, N15389, N8273, N12010, N5130);
not NOT1 (N15391, N15381);
and AND2 (N15392, N15391, N10275);
nor NOR3 (N15393, N15375, N3346, N9036);
xor XOR2 (N15394, N15386, N6012);
xor XOR2 (N15395, N15382, N12438);
or OR4 (N15396, N15388, N12020, N6137, N7595);
buf BUF1 (N15397, N15395);
nor NOR2 (N15398, N15367, N7112);
nand NAND4 (N15399, N15384, N3815, N7786, N2573);
or OR2 (N15400, N15392, N12878);
and AND2 (N15401, N15378, N12575);
xor XOR2 (N15402, N15396, N6943);
and AND2 (N15403, N15385, N13860);
not NOT1 (N15404, N15399);
xor XOR2 (N15405, N15393, N8377);
nand NAND3 (N15406, N15402, N4602, N5388);
not NOT1 (N15407, N15400);
nor NOR2 (N15408, N15407, N10945);
nor NOR3 (N15409, N15390, N11158, N10100);
or OR2 (N15410, N15401, N13835);
and AND4 (N15411, N15394, N4723, N8581, N10853);
or OR2 (N15412, N15405, N14151);
not NOT1 (N15413, N15398);
not NOT1 (N15414, N15410);
and AND3 (N15415, N15404, N12721, N11994);
not NOT1 (N15416, N15406);
and AND4 (N15417, N15411, N1678, N9356, N4887);
not NOT1 (N15418, N15416);
xor XOR2 (N15419, N15417, N14624);
nand NAND2 (N15420, N15412, N13368);
nand NAND2 (N15421, N15414, N3467);
not NOT1 (N15422, N15419);
not NOT1 (N15423, N15403);
not NOT1 (N15424, N15413);
xor XOR2 (N15425, N15421, N11534);
or OR3 (N15426, N15423, N13473, N2059);
xor XOR2 (N15427, N15409, N7371);
nand NAND3 (N15428, N15418, N8393, N5790);
nand NAND3 (N15429, N15425, N911, N5231);
buf BUF1 (N15430, N15420);
not NOT1 (N15431, N15397);
and AND3 (N15432, N15431, N5571, N11325);
not NOT1 (N15433, N15424);
nand NAND4 (N15434, N15415, N6266, N4036, N12790);
nand NAND2 (N15435, N15426, N6237);
not NOT1 (N15436, N15408);
and AND2 (N15437, N15436, N10794);
nand NAND3 (N15438, N15433, N1592, N7203);
and AND3 (N15439, N15430, N6736, N402);
nor NOR4 (N15440, N15432, N983, N8432, N10291);
or OR2 (N15441, N15438, N2158);
nor NOR2 (N15442, N15434, N4224);
xor XOR2 (N15443, N15435, N7943);
buf BUF1 (N15444, N15429);
nand NAND2 (N15445, N15428, N1510);
not NOT1 (N15446, N15427);
nor NOR2 (N15447, N15446, N3153);
xor XOR2 (N15448, N15437, N11946);
and AND3 (N15449, N15440, N3735, N10501);
nor NOR3 (N15450, N15444, N15199, N3716);
buf BUF1 (N15451, N15449);
or OR4 (N15452, N15442, N5750, N11803, N5121);
not NOT1 (N15453, N15422);
or OR4 (N15454, N15448, N9800, N8836, N2123);
nor NOR4 (N15455, N15452, N6263, N8608, N12208);
and AND2 (N15456, N15447, N12839);
nor NOR3 (N15457, N15455, N6504, N2549);
or OR3 (N15458, N15441, N6772, N2953);
nor NOR2 (N15459, N15445, N8563);
nand NAND4 (N15460, N15458, N8962, N10234, N8230);
nand NAND3 (N15461, N15456, N1954, N11421);
xor XOR2 (N15462, N15439, N1139);
nand NAND2 (N15463, N15461, N929);
xor XOR2 (N15464, N15454, N13027);
buf BUF1 (N15465, N15457);
nand NAND2 (N15466, N15463, N2703);
xor XOR2 (N15467, N15465, N6058);
xor XOR2 (N15468, N15451, N4854);
and AND2 (N15469, N15466, N7093);
xor XOR2 (N15470, N15460, N13127);
nand NAND4 (N15471, N15443, N14577, N14394, N10324);
nor NOR2 (N15472, N15450, N11568);
not NOT1 (N15473, N15459);
not NOT1 (N15474, N15462);
not NOT1 (N15475, N15464);
buf BUF1 (N15476, N15470);
nor NOR3 (N15477, N15474, N9321, N28);
buf BUF1 (N15478, N15473);
xor XOR2 (N15479, N15475, N13826);
not NOT1 (N15480, N15469);
nand NAND4 (N15481, N15480, N3344, N13140, N2739);
buf BUF1 (N15482, N15471);
nand NAND3 (N15483, N15478, N1666, N11499);
and AND2 (N15484, N15472, N12855);
xor XOR2 (N15485, N15479, N1441);
or OR2 (N15486, N15467, N6052);
nor NOR3 (N15487, N15482, N2376, N5372);
not NOT1 (N15488, N15484);
or OR2 (N15489, N15483, N2670);
or OR4 (N15490, N15453, N11354, N7204, N4663);
xor XOR2 (N15491, N15477, N894);
or OR2 (N15492, N15491, N3556);
nand NAND2 (N15493, N15489, N12345);
nor NOR4 (N15494, N15468, N13068, N10586, N4623);
buf BUF1 (N15495, N15493);
or OR4 (N15496, N15494, N7611, N6889, N4822);
xor XOR2 (N15497, N15490, N6143);
xor XOR2 (N15498, N15485, N5080);
or OR3 (N15499, N15496, N11925, N1412);
nor NOR2 (N15500, N15495, N11146);
and AND2 (N15501, N15476, N6026);
nor NOR4 (N15502, N15498, N9486, N8387, N10265);
buf BUF1 (N15503, N15486);
nand NAND3 (N15504, N15502, N5209, N4435);
and AND3 (N15505, N15501, N1663, N3264);
nor NOR4 (N15506, N15500, N10388, N7498, N6011);
and AND3 (N15507, N15492, N8120, N10791);
or OR2 (N15508, N15499, N12284);
nand NAND2 (N15509, N15507, N10610);
or OR3 (N15510, N15481, N1177, N9895);
xor XOR2 (N15511, N15487, N8469);
nor NOR3 (N15512, N15510, N3686, N9537);
or OR3 (N15513, N15497, N3983, N14982);
or OR4 (N15514, N15503, N3662, N14180, N2561);
buf BUF1 (N15515, N15509);
not NOT1 (N15516, N15488);
or OR2 (N15517, N15514, N1365);
not NOT1 (N15518, N15511);
nand NAND4 (N15519, N15512, N7939, N12884, N7074);
nand NAND3 (N15520, N15506, N2547, N153);
buf BUF1 (N15521, N15520);
or OR2 (N15522, N15519, N14092);
nand NAND3 (N15523, N15516, N6695, N11582);
nor NOR4 (N15524, N15505, N4080, N9137, N7104);
nor NOR3 (N15525, N15515, N8219, N10152);
nand NAND4 (N15526, N15521, N15214, N12308, N11090);
xor XOR2 (N15527, N15518, N8453);
nand NAND2 (N15528, N15504, N5164);
or OR3 (N15529, N15522, N10059, N4962);
or OR3 (N15530, N15523, N6172, N219);
nand NAND4 (N15531, N15529, N14378, N8414, N10196);
not NOT1 (N15532, N15508);
or OR2 (N15533, N15528, N729);
nand NAND3 (N15534, N15531, N8697, N4054);
and AND3 (N15535, N15524, N5550, N5125);
nand NAND2 (N15536, N15533, N11057);
nand NAND2 (N15537, N15513, N7193);
not NOT1 (N15538, N15526);
nand NAND3 (N15539, N15525, N8548, N12809);
nand NAND3 (N15540, N15536, N14358, N2905);
buf BUF1 (N15541, N15537);
nor NOR3 (N15542, N15541, N644, N12275);
nor NOR4 (N15543, N15527, N3028, N28, N10568);
buf BUF1 (N15544, N15535);
not NOT1 (N15545, N15530);
buf BUF1 (N15546, N15534);
and AND2 (N15547, N15517, N11692);
and AND4 (N15548, N15542, N11188, N12554, N5736);
xor XOR2 (N15549, N15543, N2340);
or OR2 (N15550, N15545, N10051);
nand NAND4 (N15551, N15546, N10530, N4262, N175);
or OR3 (N15552, N15538, N8692, N4394);
nand NAND4 (N15553, N15552, N1891, N2953, N2141);
xor XOR2 (N15554, N15549, N15077);
and AND3 (N15555, N15539, N4846, N6097);
xor XOR2 (N15556, N15544, N11840);
not NOT1 (N15557, N15550);
and AND3 (N15558, N15532, N2879, N12895);
nor NOR2 (N15559, N15548, N10348);
or OR3 (N15560, N15557, N4549, N12477);
or OR4 (N15561, N15559, N1693, N13737, N8111);
nand NAND2 (N15562, N15547, N10926);
buf BUF1 (N15563, N15554);
nor NOR3 (N15564, N15556, N9365, N721);
buf BUF1 (N15565, N15562);
not NOT1 (N15566, N15560);
and AND2 (N15567, N15551, N7988);
xor XOR2 (N15568, N15553, N352);
nand NAND3 (N15569, N15540, N3455, N4065);
or OR4 (N15570, N15558, N13542, N981, N4050);
xor XOR2 (N15571, N15568, N8535);
nor NOR4 (N15572, N15566, N15509, N14431, N2975);
not NOT1 (N15573, N15555);
nor NOR4 (N15574, N15573, N2992, N15548, N9524);
xor XOR2 (N15575, N15565, N4493);
nor NOR4 (N15576, N15572, N5090, N10165, N8262);
xor XOR2 (N15577, N15561, N14303);
buf BUF1 (N15578, N15564);
or OR2 (N15579, N15575, N5343);
not NOT1 (N15580, N15574);
buf BUF1 (N15581, N15570);
nand NAND3 (N15582, N15581, N2578, N11305);
nand NAND2 (N15583, N15577, N3175);
or OR4 (N15584, N15582, N1899, N14720, N3872);
nor NOR3 (N15585, N15563, N6274, N9848);
and AND3 (N15586, N15580, N7987, N4825);
and AND2 (N15587, N15585, N8688);
nand NAND3 (N15588, N15567, N651, N8261);
nor NOR4 (N15589, N15584, N6511, N12751, N598);
nand NAND4 (N15590, N15587, N5377, N4374, N4534);
buf BUF1 (N15591, N15588);
and AND3 (N15592, N15578, N2361, N9560);
buf BUF1 (N15593, N15591);
or OR2 (N15594, N15569, N14215);
buf BUF1 (N15595, N15579);
nand NAND3 (N15596, N15590, N14982, N1652);
nand NAND3 (N15597, N15596, N7403, N12510);
nor NOR4 (N15598, N15592, N1523, N13747, N14907);
buf BUF1 (N15599, N15594);
not NOT1 (N15600, N15589);
xor XOR2 (N15601, N15583, N15523);
nor NOR3 (N15602, N15597, N10131, N11721);
nor NOR2 (N15603, N15599, N7014);
or OR2 (N15604, N15593, N3328);
buf BUF1 (N15605, N15603);
and AND4 (N15606, N15571, N2655, N5681, N5343);
buf BUF1 (N15607, N15601);
not NOT1 (N15608, N15602);
xor XOR2 (N15609, N15607, N3775);
nand NAND2 (N15610, N15586, N3481);
buf BUF1 (N15611, N15606);
nand NAND4 (N15612, N15604, N13774, N2874, N4977);
or OR4 (N15613, N15595, N5650, N7384, N7547);
and AND3 (N15614, N15611, N4786, N7311);
or OR2 (N15615, N15605, N6104);
buf BUF1 (N15616, N15612);
nand NAND4 (N15617, N15598, N9951, N6995, N14668);
not NOT1 (N15618, N15610);
buf BUF1 (N15619, N15618);
or OR3 (N15620, N15615, N10087, N15548);
buf BUF1 (N15621, N15619);
not NOT1 (N15622, N15614);
nand NAND4 (N15623, N15622, N11152, N6661, N3650);
nor NOR4 (N15624, N15600, N9253, N2590, N13636);
buf BUF1 (N15625, N15613);
not NOT1 (N15626, N15621);
nor NOR2 (N15627, N15620, N1413);
xor XOR2 (N15628, N15626, N6213);
xor XOR2 (N15629, N15624, N7736);
or OR4 (N15630, N15609, N1323, N9024, N4268);
xor XOR2 (N15631, N15625, N9967);
not NOT1 (N15632, N15628);
xor XOR2 (N15633, N15629, N7171);
nor NOR3 (N15634, N15631, N8502, N9515);
or OR2 (N15635, N15617, N3922);
nand NAND3 (N15636, N15627, N10938, N10636);
nand NAND3 (N15637, N15616, N13561, N4917);
buf BUF1 (N15638, N15630);
nand NAND3 (N15639, N15623, N12826, N542);
xor XOR2 (N15640, N15632, N2094);
xor XOR2 (N15641, N15633, N2135);
xor XOR2 (N15642, N15640, N8537);
and AND3 (N15643, N15641, N13506, N5068);
and AND2 (N15644, N15638, N12377);
buf BUF1 (N15645, N15576);
or OR4 (N15646, N15637, N7205, N15382, N6891);
or OR4 (N15647, N15639, N6271, N3296, N8945);
and AND3 (N15648, N15642, N1987, N8284);
xor XOR2 (N15649, N15646, N9573);
not NOT1 (N15650, N15643);
and AND4 (N15651, N15634, N13945, N14918, N6901);
and AND4 (N15652, N15648, N10002, N8329, N978);
buf BUF1 (N15653, N15652);
and AND2 (N15654, N15653, N1992);
nor NOR2 (N15655, N15651, N12303);
or OR3 (N15656, N15654, N1244, N9867);
buf BUF1 (N15657, N15655);
buf BUF1 (N15658, N15657);
nor NOR4 (N15659, N15635, N9641, N14082, N8150);
nand NAND3 (N15660, N15608, N8810, N283);
nor NOR2 (N15661, N15656, N10909);
nand NAND4 (N15662, N15645, N10133, N9477, N628);
nand NAND3 (N15663, N15647, N14276, N145);
nor NOR4 (N15664, N15658, N11338, N3215, N425);
xor XOR2 (N15665, N15662, N890);
nand NAND4 (N15666, N15650, N14423, N3982, N721);
nor NOR2 (N15667, N15665, N5721);
nor NOR2 (N15668, N15666, N4833);
and AND3 (N15669, N15660, N11511, N2717);
xor XOR2 (N15670, N15668, N13664);
xor XOR2 (N15671, N15670, N631);
and AND2 (N15672, N15659, N5392);
xor XOR2 (N15673, N15667, N5547);
or OR3 (N15674, N15661, N3696, N5836);
and AND3 (N15675, N15673, N15106, N2875);
nand NAND3 (N15676, N15664, N13485, N6272);
nor NOR3 (N15677, N15675, N5131, N11705);
not NOT1 (N15678, N15672);
or OR3 (N15679, N15678, N15306, N3116);
nand NAND3 (N15680, N15674, N2796, N11898);
or OR4 (N15681, N15663, N10351, N8461, N7366);
xor XOR2 (N15682, N15671, N3105);
and AND4 (N15683, N15681, N2940, N10181, N5399);
xor XOR2 (N15684, N15682, N12867);
xor XOR2 (N15685, N15636, N9873);
xor XOR2 (N15686, N15669, N15495);
nor NOR4 (N15687, N15649, N10762, N5547, N1326);
and AND3 (N15688, N15687, N12882, N2257);
and AND3 (N15689, N15685, N257, N10756);
not NOT1 (N15690, N15676);
not NOT1 (N15691, N15689);
or OR4 (N15692, N15683, N699, N13927, N690);
xor XOR2 (N15693, N15680, N14139);
xor XOR2 (N15694, N15679, N3169);
buf BUF1 (N15695, N15677);
xor XOR2 (N15696, N15688, N5245);
nor NOR3 (N15697, N15696, N2043, N7029);
or OR4 (N15698, N15695, N14082, N2804, N12300);
xor XOR2 (N15699, N15644, N11271);
buf BUF1 (N15700, N15694);
xor XOR2 (N15701, N15691, N12081);
xor XOR2 (N15702, N15686, N6111);
not NOT1 (N15703, N15702);
nor NOR4 (N15704, N15693, N3780, N8301, N7424);
nor NOR2 (N15705, N15699, N9487);
nand NAND2 (N15706, N15701, N3202);
xor XOR2 (N15707, N15706, N11015);
nor NOR3 (N15708, N15705, N3434, N14701);
not NOT1 (N15709, N15697);
nand NAND2 (N15710, N15692, N4502);
xor XOR2 (N15711, N15708, N14288);
not NOT1 (N15712, N15711);
nand NAND3 (N15713, N15703, N10583, N2231);
nor NOR3 (N15714, N15710, N8382, N5266);
not NOT1 (N15715, N15712);
buf BUF1 (N15716, N15713);
buf BUF1 (N15717, N15684);
nand NAND4 (N15718, N15700, N13220, N11404, N8897);
buf BUF1 (N15719, N15715);
or OR3 (N15720, N15714, N336, N2789);
buf BUF1 (N15721, N15707);
xor XOR2 (N15722, N15709, N6857);
not NOT1 (N15723, N15718);
or OR4 (N15724, N15723, N8114, N7074, N7951);
xor XOR2 (N15725, N15704, N6882);
nand NAND2 (N15726, N15725, N799);
buf BUF1 (N15727, N15719);
nand NAND4 (N15728, N15698, N10660, N2410, N5089);
and AND2 (N15729, N15722, N5607);
buf BUF1 (N15730, N15728);
not NOT1 (N15731, N15724);
nor NOR3 (N15732, N15729, N8195, N7603);
buf BUF1 (N15733, N15720);
or OR2 (N15734, N15717, N13144);
xor XOR2 (N15735, N15727, N13935);
nor NOR4 (N15736, N15690, N2159, N14287, N4140);
and AND3 (N15737, N15726, N3659, N4417);
and AND4 (N15738, N15734, N4665, N15260, N11804);
nor NOR4 (N15739, N15736, N10535, N8576, N4932);
and AND2 (N15740, N15737, N5282);
not NOT1 (N15741, N15716);
buf BUF1 (N15742, N15733);
or OR4 (N15743, N15740, N6174, N12135, N12395);
nor NOR2 (N15744, N15732, N8680);
buf BUF1 (N15745, N15738);
nor NOR4 (N15746, N15742, N14897, N2313, N11478);
nand NAND2 (N15747, N15741, N1941);
or OR4 (N15748, N15743, N6843, N3876, N2403);
nand NAND2 (N15749, N15731, N10630);
not NOT1 (N15750, N15730);
or OR2 (N15751, N15735, N14527);
nand NAND4 (N15752, N15721, N11656, N8285, N10897);
nor NOR3 (N15753, N15747, N6414, N5563);
nor NOR2 (N15754, N15753, N4546);
or OR2 (N15755, N15746, N5170);
and AND4 (N15756, N15739, N319, N8443, N3497);
buf BUF1 (N15757, N15745);
and AND3 (N15758, N15749, N7904, N208);
nand NAND4 (N15759, N15754, N12927, N1750, N15412);
or OR4 (N15760, N15756, N4579, N8716, N10315);
buf BUF1 (N15761, N15760);
xor XOR2 (N15762, N15761, N6946);
buf BUF1 (N15763, N15755);
nand NAND2 (N15764, N15751, N4510);
or OR3 (N15765, N15744, N15251, N1039);
and AND3 (N15766, N15752, N3040, N5090);
not NOT1 (N15767, N15758);
xor XOR2 (N15768, N15750, N12189);
or OR3 (N15769, N15768, N8048, N3353);
xor XOR2 (N15770, N15759, N13152);
xor XOR2 (N15771, N15765, N14182);
or OR3 (N15772, N15762, N14999, N3066);
not NOT1 (N15773, N15757);
or OR4 (N15774, N15763, N9599, N11564, N1989);
nor NOR3 (N15775, N15764, N11219, N7356);
not NOT1 (N15776, N15748);
nor NOR4 (N15777, N15773, N239, N13483, N12842);
or OR3 (N15778, N15767, N1127, N4545);
or OR4 (N15779, N15774, N9881, N10462, N9102);
not NOT1 (N15780, N15766);
not NOT1 (N15781, N15777);
or OR4 (N15782, N15771, N15004, N12111, N15152);
or OR3 (N15783, N15770, N15767, N10134);
buf BUF1 (N15784, N15776);
nor NOR2 (N15785, N15779, N8435);
buf BUF1 (N15786, N15783);
xor XOR2 (N15787, N15769, N3511);
xor XOR2 (N15788, N15780, N4106);
nor NOR4 (N15789, N15782, N4509, N5227, N15274);
or OR2 (N15790, N15786, N15719);
xor XOR2 (N15791, N15789, N424);
nand NAND2 (N15792, N15791, N5158);
and AND4 (N15793, N15790, N12155, N9186, N1911);
buf BUF1 (N15794, N15787);
not NOT1 (N15795, N15778);
xor XOR2 (N15796, N15785, N14202);
nand NAND2 (N15797, N15792, N12792);
xor XOR2 (N15798, N15796, N9837);
or OR2 (N15799, N15772, N13548);
and AND2 (N15800, N15799, N7572);
not NOT1 (N15801, N15800);
buf BUF1 (N15802, N15795);
not NOT1 (N15803, N15802);
xor XOR2 (N15804, N15781, N7825);
or OR2 (N15805, N15798, N15023);
not NOT1 (N15806, N15793);
not NOT1 (N15807, N15784);
xor XOR2 (N15808, N15775, N1449);
or OR3 (N15809, N15805, N7056, N3080);
buf BUF1 (N15810, N15803);
and AND2 (N15811, N15809, N10898);
nor NOR2 (N15812, N15811, N2439);
nand NAND3 (N15813, N15797, N11639, N12622);
or OR2 (N15814, N15806, N4393);
nor NOR2 (N15815, N15794, N14615);
not NOT1 (N15816, N15788);
xor XOR2 (N15817, N15813, N2907);
not NOT1 (N15818, N15810);
and AND4 (N15819, N15804, N217, N1128, N1643);
nor NOR4 (N15820, N15812, N12726, N8928, N2144);
or OR4 (N15821, N15818, N5381, N15601, N4081);
nor NOR4 (N15822, N15820, N2627, N15427, N15736);
or OR4 (N15823, N15816, N8569, N1120, N75);
or OR4 (N15824, N15807, N699, N7135, N2506);
xor XOR2 (N15825, N15823, N7140);
xor XOR2 (N15826, N15808, N5739);
nor NOR2 (N15827, N15824, N9295);
and AND4 (N15828, N15815, N1805, N4244, N4580);
not NOT1 (N15829, N15825);
or OR3 (N15830, N15819, N2495, N10323);
nand NAND4 (N15831, N15827, N1703, N8479, N14512);
xor XOR2 (N15832, N15817, N2852);
nand NAND2 (N15833, N15826, N2642);
nor NOR2 (N15834, N15829, N14071);
and AND2 (N15835, N15814, N4169);
not NOT1 (N15836, N15822);
xor XOR2 (N15837, N15801, N4080);
not NOT1 (N15838, N15821);
nand NAND2 (N15839, N15831, N13699);
buf BUF1 (N15840, N15832);
buf BUF1 (N15841, N15836);
and AND3 (N15842, N15834, N10358, N12433);
or OR4 (N15843, N15830, N1545, N4714, N7269);
xor XOR2 (N15844, N15839, N10450);
and AND3 (N15845, N15840, N737, N15547);
nand NAND4 (N15846, N15838, N8622, N4272, N10649);
nor NOR3 (N15847, N15833, N3273, N1941);
nor NOR4 (N15848, N15835, N1890, N9127, N8135);
nor NOR3 (N15849, N15848, N3133, N13729);
nand NAND4 (N15850, N15844, N8447, N15036, N1929);
buf BUF1 (N15851, N15850);
buf BUF1 (N15852, N15828);
and AND2 (N15853, N15837, N14532);
buf BUF1 (N15854, N15841);
nand NAND4 (N15855, N15853, N7244, N3734, N13495);
and AND3 (N15856, N15849, N9006, N6326);
and AND2 (N15857, N15852, N3080);
or OR4 (N15858, N15857, N2690, N14988, N1543);
or OR3 (N15859, N15856, N4566, N11404);
and AND4 (N15860, N15847, N14355, N5183, N9164);
nor NOR3 (N15861, N15845, N4497, N13051);
nor NOR3 (N15862, N15861, N10821, N8964);
or OR2 (N15863, N15855, N328);
not NOT1 (N15864, N15854);
buf BUF1 (N15865, N15843);
nand NAND3 (N15866, N15863, N13741, N7232);
or OR4 (N15867, N15865, N5881, N9571, N4419);
not NOT1 (N15868, N15864);
not NOT1 (N15869, N15866);
xor XOR2 (N15870, N15846, N8500);
or OR2 (N15871, N15858, N4251);
nand NAND2 (N15872, N15862, N11912);
nand NAND2 (N15873, N15870, N8277);
not NOT1 (N15874, N15873);
and AND4 (N15875, N15868, N11083, N1415, N10119);
buf BUF1 (N15876, N15851);
nand NAND2 (N15877, N15876, N13734);
nor NOR4 (N15878, N15877, N9088, N450, N1453);
xor XOR2 (N15879, N15872, N10215);
not NOT1 (N15880, N15860);
and AND2 (N15881, N15878, N14969);
not NOT1 (N15882, N15880);
nor NOR4 (N15883, N15881, N10808, N2807, N6988);
not NOT1 (N15884, N15859);
buf BUF1 (N15885, N15875);
not NOT1 (N15886, N15884);
and AND2 (N15887, N15869, N8426);
buf BUF1 (N15888, N15883);
not NOT1 (N15889, N15886);
nand NAND4 (N15890, N15867, N1240, N14654, N13283);
buf BUF1 (N15891, N15882);
nand NAND2 (N15892, N15871, N13593);
and AND3 (N15893, N15842, N2073, N8135);
nor NOR3 (N15894, N15888, N11445, N15119);
buf BUF1 (N15895, N15890);
not NOT1 (N15896, N15894);
and AND4 (N15897, N15889, N1270, N3678, N11594);
and AND2 (N15898, N15895, N9254);
nor NOR4 (N15899, N15896, N7944, N14431, N6015);
buf BUF1 (N15900, N15887);
or OR2 (N15901, N15885, N1587);
nand NAND2 (N15902, N15900, N4155);
xor XOR2 (N15903, N15893, N5820);
nor NOR4 (N15904, N15901, N15139, N10347, N5451);
xor XOR2 (N15905, N15897, N13258);
not NOT1 (N15906, N15904);
not NOT1 (N15907, N15902);
not NOT1 (N15908, N15899);
and AND2 (N15909, N15903, N3861);
xor XOR2 (N15910, N15906, N6134);
or OR2 (N15911, N15908, N4405);
not NOT1 (N15912, N15874);
nand NAND3 (N15913, N15905, N1939, N6709);
xor XOR2 (N15914, N15910, N7226);
and AND3 (N15915, N15911, N14381, N7293);
nand NAND4 (N15916, N15879, N14545, N5656, N10730);
or OR3 (N15917, N15916, N683, N12128);
xor XOR2 (N15918, N15898, N10577);
nor NOR3 (N15919, N15917, N3231, N9976);
nand NAND3 (N15920, N15919, N6926, N14305);
or OR4 (N15921, N15907, N10404, N5897, N5349);
nand NAND4 (N15922, N15892, N6729, N13599, N3295);
xor XOR2 (N15923, N15891, N8403);
buf BUF1 (N15924, N15909);
and AND4 (N15925, N15922, N4777, N6459, N14965);
nand NAND3 (N15926, N15918, N10247, N592);
or OR3 (N15927, N15921, N12023, N11361);
nor NOR2 (N15928, N15927, N5614);
or OR3 (N15929, N15925, N5767, N9879);
buf BUF1 (N15930, N15914);
nor NOR2 (N15931, N15915, N11413);
nand NAND2 (N15932, N15929, N4217);
nor NOR2 (N15933, N15913, N987);
xor XOR2 (N15934, N15931, N13086);
or OR2 (N15935, N15932, N10154);
buf BUF1 (N15936, N15930);
or OR4 (N15937, N15920, N12481, N15742, N13034);
or OR3 (N15938, N15937, N9924, N14394);
or OR2 (N15939, N15934, N5283);
nor NOR3 (N15940, N15912, N13973, N8140);
nor NOR3 (N15941, N15936, N2235, N5657);
buf BUF1 (N15942, N15926);
buf BUF1 (N15943, N15940);
not NOT1 (N15944, N15933);
nor NOR3 (N15945, N15944, N2429, N6401);
not NOT1 (N15946, N15943);
xor XOR2 (N15947, N15945, N11836);
or OR4 (N15948, N15935, N437, N2304, N7488);
buf BUF1 (N15949, N15946);
buf BUF1 (N15950, N15948);
or OR2 (N15951, N15923, N5842);
nor NOR4 (N15952, N15949, N122, N11509, N12693);
nand NAND3 (N15953, N15928, N3279, N8902);
and AND4 (N15954, N15942, N6949, N7716, N6924);
and AND4 (N15955, N15953, N12876, N11002, N3754);
buf BUF1 (N15956, N15950);
nor NOR3 (N15957, N15939, N2112, N5771);
and AND2 (N15958, N15924, N4257);
xor XOR2 (N15959, N15954, N1856);
not NOT1 (N15960, N15952);
buf BUF1 (N15961, N15951);
or OR4 (N15962, N15955, N5732, N1765, N12648);
and AND2 (N15963, N15962, N1145);
nand NAND2 (N15964, N15957, N8715);
and AND3 (N15965, N15964, N13947, N12116);
xor XOR2 (N15966, N15963, N10395);
not NOT1 (N15967, N15966);
nand NAND2 (N15968, N15967, N6782);
and AND2 (N15969, N15938, N14105);
buf BUF1 (N15970, N15959);
and AND4 (N15971, N15956, N599, N1626, N11835);
or OR4 (N15972, N15971, N1646, N7377, N7851);
and AND2 (N15973, N15961, N4221);
nand NAND4 (N15974, N15969, N15144, N1119, N340);
buf BUF1 (N15975, N15974);
or OR2 (N15976, N15960, N10630);
nand NAND3 (N15977, N15970, N12533, N12511);
xor XOR2 (N15978, N15977, N6961);
xor XOR2 (N15979, N15972, N5632);
buf BUF1 (N15980, N15941);
not NOT1 (N15981, N15979);
or OR3 (N15982, N15978, N1513, N1944);
and AND4 (N15983, N15976, N8370, N8966, N3930);
nand NAND3 (N15984, N15973, N10011, N7561);
not NOT1 (N15985, N15983);
and AND4 (N15986, N15984, N15822, N10971, N12386);
nand NAND4 (N15987, N15980, N298, N11074, N10183);
not NOT1 (N15988, N15982);
and AND4 (N15989, N15988, N15774, N9247, N14002);
xor XOR2 (N15990, N15986, N1773);
or OR4 (N15991, N15987, N10637, N2203, N2979);
xor XOR2 (N15992, N15990, N1410);
nor NOR3 (N15993, N15947, N15924, N4994);
xor XOR2 (N15994, N15968, N7965);
xor XOR2 (N15995, N15991, N14992);
nand NAND2 (N15996, N15989, N2224);
and AND4 (N15997, N15995, N6313, N11373, N8360);
and AND2 (N15998, N15985, N7452);
nor NOR4 (N15999, N15997, N14287, N8129, N6874);
or OR3 (N16000, N15992, N14041, N7708);
and AND4 (N16001, N15975, N6507, N6899, N917);
and AND4 (N16002, N16000, N5729, N11510, N3100);
not NOT1 (N16003, N15965);
and AND4 (N16004, N15994, N11824, N13309, N15257);
and AND2 (N16005, N15996, N3152);
and AND4 (N16006, N15998, N10268, N6589, N9540);
nand NAND2 (N16007, N15981, N2333);
buf BUF1 (N16008, N16007);
or OR3 (N16009, N16005, N12421, N8861);
and AND3 (N16010, N16004, N14304, N8417);
nor NOR2 (N16011, N16006, N8851);
endmodule