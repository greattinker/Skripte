// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N1523,N1514,N1521,N1512,N1522,N1519,N1520,N1508,N1517,N1524;

not NOT1 (N25, N15);
nand NAND3 (N26, N15, N3, N21);
xor XOR2 (N27, N15, N26);
xor XOR2 (N28, N22, N24);
nand NAND3 (N29, N26, N21, N2);
not NOT1 (N30, N7);
or OR2 (N31, N22, N17);
not NOT1 (N32, N9);
not NOT1 (N33, N7);
or OR2 (N34, N30, N22);
xor XOR2 (N35, N26, N2);
and AND3 (N36, N9, N10, N16);
nand NAND4 (N37, N33, N11, N4, N10);
not NOT1 (N38, N36);
and AND2 (N39, N37, N34);
nand NAND2 (N40, N19, N28);
nand NAND3 (N41, N23, N5, N25);
and AND4 (N42, N24, N2, N25, N31);
not NOT1 (N43, N6);
and AND3 (N44, N40, N27, N41);
xor XOR2 (N45, N17, N24);
not NOT1 (N46, N38);
or OR2 (N47, N46, N5);
buf BUF1 (N48, N15);
or OR4 (N49, N32, N26, N37, N15);
nor NOR3 (N50, N29, N36, N26);
nand NAND4 (N51, N49, N48, N19, N4);
nand NAND2 (N52, N37, N7);
not NOT1 (N53, N42);
or OR3 (N54, N53, N53, N14);
nand NAND2 (N55, N39, N36);
or OR4 (N56, N45, N3, N6, N21);
nor NOR3 (N57, N43, N13, N47);
nand NAND3 (N58, N38, N11, N29);
and AND4 (N59, N50, N10, N16, N14);
nand NAND2 (N60, N44, N1);
nor NOR2 (N61, N59, N51);
buf BUF1 (N62, N29);
xor XOR2 (N63, N55, N23);
nor NOR3 (N64, N54, N31, N41);
or OR4 (N65, N52, N19, N33, N29);
or OR4 (N66, N56, N4, N51, N18);
and AND2 (N67, N61, N1);
xor XOR2 (N68, N57, N38);
or OR2 (N69, N58, N10);
xor XOR2 (N70, N69, N34);
and AND4 (N71, N67, N54, N70, N10);
nor NOR3 (N72, N53, N71, N58);
and AND2 (N73, N23, N30);
or OR3 (N74, N72, N12, N40);
or OR4 (N75, N63, N14, N35, N46);
not NOT1 (N76, N11);
xor XOR2 (N77, N64, N38);
buf BUF1 (N78, N68);
and AND2 (N79, N62, N38);
xor XOR2 (N80, N65, N75);
or OR3 (N81, N35, N6, N18);
not NOT1 (N82, N66);
xor XOR2 (N83, N73, N67);
nand NAND3 (N84, N60, N51, N63);
not NOT1 (N85, N74);
not NOT1 (N86, N82);
nor NOR4 (N87, N83, N62, N11, N5);
nand NAND2 (N88, N86, N66);
nand NAND2 (N89, N80, N33);
not NOT1 (N90, N76);
xor XOR2 (N91, N79, N78);
xor XOR2 (N92, N39, N71);
and AND2 (N93, N88, N82);
xor XOR2 (N94, N77, N89);
and AND4 (N95, N15, N89, N72, N12);
nand NAND3 (N96, N84, N57, N89);
nand NAND4 (N97, N94, N59, N78, N72);
and AND3 (N98, N85, N7, N53);
and AND2 (N99, N95, N20);
xor XOR2 (N100, N92, N13);
nor NOR3 (N101, N90, N88, N44);
xor XOR2 (N102, N100, N61);
buf BUF1 (N103, N81);
or OR2 (N104, N98, N72);
nor NOR3 (N105, N101, N62, N35);
and AND3 (N106, N96, N35, N75);
buf BUF1 (N107, N93);
nand NAND3 (N108, N106, N77, N80);
nand NAND2 (N109, N91, N9);
nand NAND4 (N110, N107, N22, N48, N44);
and AND2 (N111, N105, N57);
not NOT1 (N112, N103);
or OR4 (N113, N112, N28, N82, N91);
not NOT1 (N114, N99);
nand NAND2 (N115, N114, N102);
buf BUF1 (N116, N97);
nand NAND2 (N117, N91, N100);
not NOT1 (N118, N108);
xor XOR2 (N119, N118, N104);
and AND3 (N120, N90, N52, N90);
or OR2 (N121, N116, N47);
buf BUF1 (N122, N109);
or OR2 (N123, N113, N58);
and AND4 (N124, N115, N93, N47, N101);
xor XOR2 (N125, N119, N110);
nor NOR3 (N126, N114, N83, N99);
and AND4 (N127, N120, N23, N105, N109);
nor NOR2 (N128, N123, N43);
xor XOR2 (N129, N121, N13);
buf BUF1 (N130, N117);
nor NOR4 (N131, N87, N1, N113, N114);
and AND3 (N132, N111, N60, N67);
or OR4 (N133, N131, N115, N82, N128);
buf BUF1 (N134, N38);
nand NAND3 (N135, N134, N78, N113);
nor NOR2 (N136, N125, N99);
not NOT1 (N137, N126);
nor NOR4 (N138, N136, N32, N71, N2);
buf BUF1 (N139, N133);
and AND3 (N140, N122, N84, N128);
and AND2 (N141, N130, N26);
xor XOR2 (N142, N135, N20);
buf BUF1 (N143, N132);
or OR4 (N144, N138, N34, N104, N125);
nand NAND4 (N145, N143, N43, N30, N5);
nor NOR2 (N146, N140, N134);
buf BUF1 (N147, N129);
or OR3 (N148, N146, N136, N18);
nand NAND2 (N149, N141, N69);
and AND4 (N150, N124, N37, N4, N55);
or OR2 (N151, N137, N106);
nor NOR4 (N152, N149, N67, N39, N39);
buf BUF1 (N153, N147);
not NOT1 (N154, N152);
nor NOR3 (N155, N142, N120, N48);
nor NOR4 (N156, N139, N56, N36, N148);
and AND2 (N157, N115, N32);
nand NAND3 (N158, N154, N88, N125);
nor NOR2 (N159, N150, N152);
and AND3 (N160, N159, N56, N129);
and AND3 (N161, N145, N57, N73);
xor XOR2 (N162, N160, N117);
buf BUF1 (N163, N157);
or OR2 (N164, N156, N106);
nand NAND4 (N165, N158, N14, N93, N156);
xor XOR2 (N166, N155, N107);
and AND2 (N167, N161, N36);
buf BUF1 (N168, N165);
not NOT1 (N169, N168);
buf BUF1 (N170, N151);
and AND3 (N171, N169, N37, N158);
or OR3 (N172, N164, N100, N170);
buf BUF1 (N173, N150);
and AND2 (N174, N153, N60);
not NOT1 (N175, N171);
nand NAND3 (N176, N172, N109, N134);
nor NOR4 (N177, N144, N1, N145, N112);
nor NOR4 (N178, N176, N131, N74, N109);
buf BUF1 (N179, N177);
nor NOR4 (N180, N175, N146, N45, N147);
or OR4 (N181, N174, N138, N151, N119);
buf BUF1 (N182, N179);
nand NAND4 (N183, N182, N49, N40, N134);
nor NOR4 (N184, N178, N110, N20, N33);
and AND2 (N185, N162, N7);
and AND3 (N186, N183, N68, N96);
and AND4 (N187, N163, N184, N176, N158);
or OR3 (N188, N75, N107, N133);
nor NOR2 (N189, N188, N77);
nand NAND2 (N190, N186, N154);
nor NOR3 (N191, N167, N61, N102);
nor NOR2 (N192, N187, N168);
nand NAND2 (N193, N166, N21);
nor NOR2 (N194, N181, N22);
xor XOR2 (N195, N173, N20);
buf BUF1 (N196, N195);
xor XOR2 (N197, N185, N74);
and AND2 (N198, N193, N32);
xor XOR2 (N199, N190, N115);
or OR3 (N200, N191, N159, N74);
or OR3 (N201, N200, N93, N154);
and AND2 (N202, N201, N103);
nand NAND4 (N203, N194, N32, N185, N87);
nand NAND4 (N204, N197, N99, N9, N134);
or OR2 (N205, N196, N124);
or OR4 (N206, N189, N31, N113, N75);
not NOT1 (N207, N202);
nand NAND2 (N208, N204, N47);
or OR3 (N209, N199, N207, N38);
nand NAND4 (N210, N158, N53, N41, N171);
nand NAND4 (N211, N208, N161, N98, N139);
buf BUF1 (N212, N127);
and AND4 (N213, N211, N151, N18, N7);
buf BUF1 (N214, N198);
buf BUF1 (N215, N180);
buf BUF1 (N216, N213);
and AND4 (N217, N210, N191, N182, N48);
and AND3 (N218, N217, N79, N45);
buf BUF1 (N219, N206);
xor XOR2 (N220, N216, N53);
nor NOR3 (N221, N220, N53, N131);
and AND3 (N222, N221, N190, N71);
buf BUF1 (N223, N203);
or OR3 (N224, N209, N68, N29);
nor NOR4 (N225, N223, N23, N29, N20);
nand NAND2 (N226, N219, N149);
buf BUF1 (N227, N222);
or OR2 (N228, N205, N161);
nand NAND2 (N229, N227, N215);
or OR2 (N230, N209, N15);
xor XOR2 (N231, N226, N116);
buf BUF1 (N232, N218);
nor NOR2 (N233, N228, N127);
xor XOR2 (N234, N214, N140);
not NOT1 (N235, N234);
or OR2 (N236, N231, N235);
and AND2 (N237, N86, N74);
or OR2 (N238, N230, N140);
nor NOR3 (N239, N229, N56, N194);
nand NAND4 (N240, N237, N52, N15, N216);
and AND2 (N241, N212, N91);
or OR4 (N242, N241, N71, N31, N52);
buf BUF1 (N243, N232);
nor NOR4 (N244, N242, N164, N37, N32);
and AND4 (N245, N243, N16, N204, N155);
not NOT1 (N246, N224);
not NOT1 (N247, N244);
nand NAND4 (N248, N233, N192, N231, N50);
not NOT1 (N249, N74);
nor NOR2 (N250, N236, N217);
xor XOR2 (N251, N238, N50);
not NOT1 (N252, N225);
and AND2 (N253, N246, N243);
nor NOR3 (N254, N248, N204, N201);
or OR3 (N255, N239, N246, N84);
buf BUF1 (N256, N245);
and AND3 (N257, N249, N187, N199);
nand NAND2 (N258, N254, N248);
xor XOR2 (N259, N253, N62);
buf BUF1 (N260, N250);
nand NAND4 (N261, N255, N92, N138, N4);
buf BUF1 (N262, N256);
nor NOR4 (N263, N247, N232, N89, N223);
not NOT1 (N264, N252);
or OR4 (N265, N263, N244, N232, N57);
and AND3 (N266, N260, N157, N13);
nor NOR3 (N267, N258, N117, N95);
buf BUF1 (N268, N267);
not NOT1 (N269, N257);
or OR2 (N270, N266, N185);
or OR3 (N271, N251, N234, N126);
or OR2 (N272, N261, N252);
and AND3 (N273, N265, N54, N26);
nor NOR3 (N274, N262, N89, N211);
and AND3 (N275, N269, N13, N170);
and AND2 (N276, N271, N24);
nor NOR2 (N277, N273, N68);
nor NOR3 (N278, N259, N260, N62);
or OR2 (N279, N278, N200);
or OR2 (N280, N268, N211);
nand NAND2 (N281, N279, N184);
nor NOR3 (N282, N276, N88, N46);
and AND4 (N283, N280, N207, N165, N258);
nor NOR4 (N284, N270, N16, N152, N224);
not NOT1 (N285, N281);
buf BUF1 (N286, N275);
nor NOR2 (N287, N283, N278);
nor NOR2 (N288, N240, N253);
buf BUF1 (N289, N285);
not NOT1 (N290, N272);
nor NOR2 (N291, N277, N69);
nor NOR2 (N292, N289, N284);
nor NOR2 (N293, N139, N68);
xor XOR2 (N294, N292, N242);
buf BUF1 (N295, N290);
nand NAND4 (N296, N274, N207, N177, N2);
buf BUF1 (N297, N282);
nor NOR2 (N298, N297, N91);
buf BUF1 (N299, N298);
not NOT1 (N300, N287);
nand NAND2 (N301, N288, N277);
nand NAND3 (N302, N299, N36, N150);
nand NAND3 (N303, N294, N134, N231);
xor XOR2 (N304, N300, N87);
or OR3 (N305, N302, N78, N254);
or OR2 (N306, N303, N221);
not NOT1 (N307, N295);
nor NOR2 (N308, N301, N210);
nand NAND2 (N309, N308, N164);
nor NOR2 (N310, N293, N146);
xor XOR2 (N311, N296, N66);
buf BUF1 (N312, N291);
buf BUF1 (N313, N306);
or OR3 (N314, N304, N234, N118);
and AND4 (N315, N313, N281, N215, N20);
buf BUF1 (N316, N311);
or OR3 (N317, N309, N85, N119);
nand NAND3 (N318, N315, N184, N225);
nor NOR3 (N319, N305, N55, N78);
or OR4 (N320, N307, N187, N135, N296);
or OR3 (N321, N319, N108, N227);
nand NAND4 (N322, N317, N317, N296, N114);
or OR3 (N323, N314, N29, N288);
nor NOR3 (N324, N310, N158, N82);
buf BUF1 (N325, N322);
and AND4 (N326, N286, N46, N235, N136);
buf BUF1 (N327, N264);
not NOT1 (N328, N326);
buf BUF1 (N329, N327);
not NOT1 (N330, N324);
xor XOR2 (N331, N321, N120);
xor XOR2 (N332, N328, N29);
or OR4 (N333, N316, N266, N230, N52);
buf BUF1 (N334, N332);
nor NOR2 (N335, N331, N295);
nor NOR2 (N336, N312, N327);
nand NAND2 (N337, N334, N243);
and AND2 (N338, N325, N324);
nand NAND3 (N339, N318, N279, N217);
nand NAND4 (N340, N337, N163, N323, N128);
not NOT1 (N341, N255);
nor NOR3 (N342, N333, N277, N191);
buf BUF1 (N343, N335);
nand NAND4 (N344, N341, N51, N205, N342);
buf BUF1 (N345, N282);
nand NAND3 (N346, N344, N159, N17);
buf BUF1 (N347, N338);
or OR4 (N348, N343, N7, N221, N336);
xor XOR2 (N349, N295, N282);
nand NAND3 (N350, N348, N182, N176);
nor NOR2 (N351, N350, N240);
nor NOR2 (N352, N339, N2);
xor XOR2 (N353, N329, N250);
buf BUF1 (N354, N320);
nor NOR2 (N355, N353, N22);
nand NAND3 (N356, N330, N273, N155);
not NOT1 (N357, N354);
buf BUF1 (N358, N347);
or OR2 (N359, N346, N158);
xor XOR2 (N360, N359, N22);
or OR4 (N361, N358, N33, N286, N89);
or OR3 (N362, N357, N227, N46);
or OR4 (N363, N355, N280, N199, N88);
xor XOR2 (N364, N360, N159);
not NOT1 (N365, N352);
and AND2 (N366, N363, N319);
and AND2 (N367, N364, N352);
or OR3 (N368, N349, N157, N2);
buf BUF1 (N369, N368);
nor NOR2 (N370, N340, N136);
or OR2 (N371, N366, N298);
buf BUF1 (N372, N351);
nand NAND4 (N373, N372, N261, N251, N163);
or OR2 (N374, N369, N33);
buf BUF1 (N375, N356);
buf BUF1 (N376, N362);
not NOT1 (N377, N367);
xor XOR2 (N378, N365, N182);
nand NAND3 (N379, N375, N94, N186);
and AND4 (N380, N371, N106, N338, N87);
nand NAND3 (N381, N374, N74, N358);
not NOT1 (N382, N361);
buf BUF1 (N383, N381);
buf BUF1 (N384, N378);
nand NAND3 (N385, N380, N134, N240);
buf BUF1 (N386, N370);
and AND4 (N387, N377, N156, N228, N318);
not NOT1 (N388, N385);
or OR2 (N389, N376, N46);
and AND4 (N390, N389, N14, N367, N83);
xor XOR2 (N391, N345, N226);
and AND4 (N392, N387, N391, N324, N144);
not NOT1 (N393, N380);
nand NAND2 (N394, N393, N74);
xor XOR2 (N395, N373, N355);
xor XOR2 (N396, N388, N101);
not NOT1 (N397, N396);
nand NAND3 (N398, N394, N119, N181);
nand NAND2 (N399, N395, N217);
xor XOR2 (N400, N383, N397);
not NOT1 (N401, N296);
not NOT1 (N402, N401);
and AND2 (N403, N382, N155);
nor NOR4 (N404, N400, N113, N380, N153);
nor NOR2 (N405, N384, N255);
or OR2 (N406, N392, N302);
xor XOR2 (N407, N402, N189);
and AND3 (N408, N386, N51, N226);
buf BUF1 (N409, N406);
xor XOR2 (N410, N379, N302);
xor XOR2 (N411, N399, N224);
or OR3 (N412, N408, N320, N150);
nand NAND4 (N413, N411, N104, N188, N238);
buf BUF1 (N414, N403);
nor NOR4 (N415, N390, N190, N301, N175);
not NOT1 (N416, N398);
nand NAND3 (N417, N412, N240, N111);
nor NOR3 (N418, N414, N247, N232);
xor XOR2 (N419, N415, N70);
not NOT1 (N420, N416);
or OR3 (N421, N407, N75, N165);
buf BUF1 (N422, N417);
buf BUF1 (N423, N404);
nor NOR2 (N424, N413, N305);
xor XOR2 (N425, N410, N403);
nand NAND4 (N426, N425, N158, N396, N240);
or OR4 (N427, N422, N117, N232, N5);
xor XOR2 (N428, N424, N408);
nor NOR3 (N429, N427, N323, N93);
not NOT1 (N430, N405);
or OR3 (N431, N429, N326, N26);
or OR2 (N432, N409, N234);
or OR3 (N433, N426, N386, N11);
nand NAND4 (N434, N420, N155, N232, N76);
xor XOR2 (N435, N428, N39);
nor NOR4 (N436, N418, N158, N269, N14);
nor NOR4 (N437, N435, N57, N130, N287);
and AND4 (N438, N431, N398, N207, N364);
not NOT1 (N439, N433);
nand NAND4 (N440, N438, N76, N101, N43);
buf BUF1 (N441, N421);
nor NOR2 (N442, N440, N231);
buf BUF1 (N443, N442);
and AND3 (N444, N432, N102, N62);
buf BUF1 (N445, N437);
or OR4 (N446, N443, N177, N210, N45);
not NOT1 (N447, N445);
not NOT1 (N448, N423);
not NOT1 (N449, N434);
xor XOR2 (N450, N419, N256);
xor XOR2 (N451, N441, N450);
or OR4 (N452, N406, N239, N317, N54);
xor XOR2 (N453, N439, N344);
xor XOR2 (N454, N430, N39);
or OR4 (N455, N449, N192, N192, N185);
buf BUF1 (N456, N448);
and AND4 (N457, N454, N389, N151, N401);
buf BUF1 (N458, N455);
nor NOR2 (N459, N451, N126);
buf BUF1 (N460, N459);
not NOT1 (N461, N456);
nor NOR4 (N462, N461, N227, N171, N182);
nand NAND3 (N463, N452, N99, N167);
or OR3 (N464, N463, N399, N421);
nor NOR2 (N465, N462, N60);
not NOT1 (N466, N460);
and AND2 (N467, N465, N266);
not NOT1 (N468, N466);
and AND2 (N469, N436, N146);
nand NAND3 (N470, N444, N136, N407);
and AND4 (N471, N464, N139, N360, N177);
nand NAND3 (N472, N458, N164, N67);
buf BUF1 (N473, N468);
buf BUF1 (N474, N457);
and AND2 (N475, N446, N19);
xor XOR2 (N476, N473, N342);
nor NOR3 (N477, N467, N429, N445);
buf BUF1 (N478, N476);
nor NOR4 (N479, N474, N346, N336, N62);
xor XOR2 (N480, N477, N202);
and AND3 (N481, N479, N61, N210);
and AND4 (N482, N447, N409, N455, N331);
nand NAND2 (N483, N480, N317);
xor XOR2 (N484, N470, N147);
nor NOR2 (N485, N478, N223);
buf BUF1 (N486, N472);
buf BUF1 (N487, N481);
nand NAND2 (N488, N483, N426);
and AND4 (N489, N486, N120, N26, N275);
xor XOR2 (N490, N482, N400);
buf BUF1 (N491, N485);
xor XOR2 (N492, N491, N43);
nand NAND4 (N493, N489, N339, N223, N67);
or OR4 (N494, N490, N135, N21, N448);
buf BUF1 (N495, N471);
xor XOR2 (N496, N493, N399);
or OR3 (N497, N469, N374, N468);
xor XOR2 (N498, N484, N141);
not NOT1 (N499, N495);
not NOT1 (N500, N488);
nor NOR3 (N501, N498, N276, N126);
xor XOR2 (N502, N494, N33);
nor NOR4 (N503, N487, N416, N26, N378);
or OR3 (N504, N501, N296, N259);
not NOT1 (N505, N502);
nor NOR3 (N506, N503, N241, N350);
xor XOR2 (N507, N500, N186);
or OR4 (N508, N499, N65, N481, N298);
and AND4 (N509, N475, N109, N403, N169);
buf BUF1 (N510, N492);
xor XOR2 (N511, N505, N101);
not NOT1 (N512, N507);
xor XOR2 (N513, N453, N471);
or OR3 (N514, N512, N388, N319);
or OR4 (N515, N497, N88, N90, N341);
xor XOR2 (N516, N511, N335);
nor NOR2 (N517, N513, N390);
not NOT1 (N518, N510);
xor XOR2 (N519, N514, N90);
nand NAND4 (N520, N506, N173, N482, N494);
nor NOR4 (N521, N516, N191, N316, N447);
nand NAND4 (N522, N496, N301, N257, N80);
nand NAND3 (N523, N521, N244, N283);
buf BUF1 (N524, N520);
buf BUF1 (N525, N524);
or OR3 (N526, N522, N234, N176);
and AND3 (N527, N523, N302, N474);
or OR4 (N528, N517, N274, N74, N219);
or OR4 (N529, N518, N226, N163, N45);
nand NAND3 (N530, N515, N408, N100);
nor NOR4 (N531, N530, N198, N178, N147);
and AND2 (N532, N526, N167);
nor NOR2 (N533, N532, N352);
and AND3 (N534, N519, N461, N149);
nand NAND2 (N535, N509, N202);
not NOT1 (N536, N525);
nor NOR4 (N537, N508, N396, N141, N154);
not NOT1 (N538, N537);
nand NAND4 (N539, N527, N237, N280, N71);
nor NOR4 (N540, N539, N114, N254, N330);
xor XOR2 (N541, N535, N522);
xor XOR2 (N542, N540, N216);
or OR3 (N543, N534, N522, N99);
xor XOR2 (N544, N528, N414);
nor NOR4 (N545, N538, N339, N242, N364);
not NOT1 (N546, N536);
xor XOR2 (N547, N545, N168);
xor XOR2 (N548, N531, N108);
xor XOR2 (N549, N533, N278);
nand NAND2 (N550, N542, N85);
nor NOR4 (N551, N543, N224, N135, N485);
nand NAND4 (N552, N551, N180, N97, N540);
nor NOR4 (N553, N544, N223, N473, N437);
or OR2 (N554, N529, N517);
nor NOR3 (N555, N541, N394, N499);
or OR3 (N556, N546, N536, N356);
and AND2 (N557, N550, N492);
and AND2 (N558, N548, N350);
nand NAND4 (N559, N553, N105, N250, N90);
xor XOR2 (N560, N559, N228);
buf BUF1 (N561, N560);
not NOT1 (N562, N561);
nor NOR3 (N563, N552, N336, N10);
xor XOR2 (N564, N554, N212);
or OR4 (N565, N563, N69, N549, N526);
or OR4 (N566, N404, N18, N561, N206);
and AND4 (N567, N565, N64, N165, N496);
xor XOR2 (N568, N567, N133);
nand NAND3 (N569, N504, N196, N342);
nand NAND3 (N570, N547, N64, N59);
and AND3 (N571, N558, N16, N541);
or OR2 (N572, N566, N423);
and AND3 (N573, N562, N345, N140);
or OR2 (N574, N556, N389);
xor XOR2 (N575, N564, N274);
not NOT1 (N576, N573);
and AND4 (N577, N574, N250, N232, N367);
or OR3 (N578, N576, N308, N292);
nand NAND3 (N579, N575, N491, N369);
nor NOR3 (N580, N568, N419, N15);
not NOT1 (N581, N572);
or OR3 (N582, N557, N264, N568);
and AND3 (N583, N570, N71, N247);
not NOT1 (N584, N583);
xor XOR2 (N585, N577, N270);
xor XOR2 (N586, N584, N571);
not NOT1 (N587, N53);
buf BUF1 (N588, N579);
nor NOR2 (N589, N581, N90);
nor NOR3 (N590, N580, N420, N463);
buf BUF1 (N591, N569);
xor XOR2 (N592, N589, N425);
not NOT1 (N593, N590);
and AND2 (N594, N593, N576);
nor NOR3 (N595, N591, N569, N375);
and AND3 (N596, N587, N476, N285);
xor XOR2 (N597, N596, N156);
or OR4 (N598, N555, N259, N147, N542);
nor NOR2 (N599, N586, N336);
or OR4 (N600, N592, N143, N245, N39);
and AND4 (N601, N598, N413, N527, N464);
xor XOR2 (N602, N597, N87);
nand NAND2 (N603, N599, N473);
nor NOR3 (N604, N582, N560, N382);
not NOT1 (N605, N585);
nand NAND3 (N606, N600, N593, N29);
and AND3 (N607, N602, N258, N112);
or OR3 (N608, N605, N436, N144);
buf BUF1 (N609, N607);
buf BUF1 (N610, N608);
not NOT1 (N611, N588);
buf BUF1 (N612, N601);
or OR2 (N613, N604, N594);
buf BUF1 (N614, N211);
and AND4 (N615, N610, N94, N41, N239);
not NOT1 (N616, N611);
or OR4 (N617, N606, N31, N478, N568);
nor NOR2 (N618, N603, N357);
not NOT1 (N619, N615);
and AND3 (N620, N595, N481, N584);
or OR3 (N621, N620, N63, N166);
nand NAND2 (N622, N617, N41);
not NOT1 (N623, N619);
or OR2 (N624, N622, N277);
or OR3 (N625, N616, N140, N82);
xor XOR2 (N626, N612, N219);
or OR4 (N627, N618, N102, N2, N520);
buf BUF1 (N628, N609);
and AND2 (N629, N578, N1);
not NOT1 (N630, N614);
or OR4 (N631, N621, N578, N334, N18);
and AND2 (N632, N630, N149);
buf BUF1 (N633, N632);
and AND4 (N634, N625, N246, N486, N492);
and AND2 (N635, N633, N265);
nor NOR4 (N636, N624, N535, N288, N158);
or OR2 (N637, N626, N286);
buf BUF1 (N638, N623);
nand NAND2 (N639, N637, N91);
nor NOR3 (N640, N627, N31, N337);
or OR4 (N641, N639, N427, N47, N226);
or OR2 (N642, N640, N336);
nor NOR4 (N643, N641, N213, N634, N417);
nand NAND4 (N644, N483, N422, N634, N146);
xor XOR2 (N645, N629, N550);
xor XOR2 (N646, N635, N523);
nor NOR2 (N647, N643, N236);
not NOT1 (N648, N642);
nor NOR3 (N649, N631, N148, N404);
nor NOR4 (N650, N646, N73, N424, N416);
and AND3 (N651, N644, N350, N325);
nand NAND3 (N652, N651, N364, N94);
buf BUF1 (N653, N647);
not NOT1 (N654, N645);
buf BUF1 (N655, N650);
nand NAND3 (N656, N648, N98, N316);
nor NOR3 (N657, N638, N101, N526);
nand NAND2 (N658, N636, N198);
nor NOR4 (N659, N654, N537, N393, N85);
or OR3 (N660, N657, N270, N295);
nor NOR2 (N661, N653, N27);
buf BUF1 (N662, N658);
and AND4 (N663, N652, N594, N90, N399);
nor NOR2 (N664, N661, N222);
buf BUF1 (N665, N628);
and AND4 (N666, N665, N277, N426, N15);
nor NOR4 (N667, N613, N30, N350, N352);
nor NOR2 (N668, N659, N340);
and AND2 (N669, N667, N194);
nand NAND4 (N670, N669, N110, N535, N478);
buf BUF1 (N671, N664);
or OR2 (N672, N662, N418);
or OR3 (N673, N656, N478, N472);
buf BUF1 (N674, N663);
nand NAND3 (N675, N649, N271, N267);
nor NOR4 (N676, N655, N471, N584, N303);
nand NAND3 (N677, N675, N218, N496);
or OR4 (N678, N660, N72, N618, N523);
not NOT1 (N679, N674);
or OR2 (N680, N678, N365);
and AND4 (N681, N677, N589, N467, N96);
xor XOR2 (N682, N671, N496);
nor NOR4 (N683, N668, N166, N123, N533);
not NOT1 (N684, N680);
nor NOR3 (N685, N682, N613, N660);
nor NOR2 (N686, N666, N298);
nand NAND2 (N687, N684, N210);
not NOT1 (N688, N686);
and AND4 (N689, N673, N668, N52, N453);
buf BUF1 (N690, N689);
and AND4 (N691, N670, N353, N465, N123);
and AND3 (N692, N683, N582, N149);
not NOT1 (N693, N690);
not NOT1 (N694, N687);
buf BUF1 (N695, N693);
nand NAND2 (N696, N676, N551);
xor XOR2 (N697, N679, N669);
and AND2 (N698, N691, N400);
buf BUF1 (N699, N672);
nor NOR3 (N700, N685, N681, N543);
nor NOR2 (N701, N654, N689);
nand NAND3 (N702, N688, N338, N609);
xor XOR2 (N703, N698, N340);
nor NOR2 (N704, N700, N92);
nor NOR4 (N705, N695, N168, N432, N445);
nand NAND2 (N706, N692, N660);
and AND4 (N707, N703, N488, N260, N34);
or OR2 (N708, N694, N593);
and AND3 (N709, N699, N445, N79);
buf BUF1 (N710, N708);
buf BUF1 (N711, N705);
buf BUF1 (N712, N704);
xor XOR2 (N713, N709, N378);
and AND4 (N714, N712, N132, N321, N516);
and AND4 (N715, N711, N105, N473, N126);
xor XOR2 (N716, N713, N667);
not NOT1 (N717, N707);
not NOT1 (N718, N714);
not NOT1 (N719, N710);
buf BUF1 (N720, N715);
not NOT1 (N721, N720);
and AND2 (N722, N701, N5);
and AND3 (N723, N718, N560, N369);
or OR4 (N724, N702, N178, N458, N89);
buf BUF1 (N725, N696);
nor NOR4 (N726, N724, N448, N128, N376);
xor XOR2 (N727, N721, N214);
or OR2 (N728, N725, N341);
not NOT1 (N729, N728);
nor NOR2 (N730, N722, N525);
or OR2 (N731, N716, N406);
and AND4 (N732, N717, N648, N132, N426);
or OR4 (N733, N719, N357, N561, N227);
and AND3 (N734, N727, N590, N228);
not NOT1 (N735, N732);
xor XOR2 (N736, N697, N200);
and AND3 (N737, N723, N245, N406);
and AND2 (N738, N734, N532);
nor NOR4 (N739, N736, N235, N140, N18);
nor NOR3 (N740, N731, N673, N595);
nand NAND3 (N741, N739, N213, N607);
nand NAND3 (N742, N733, N202, N727);
nor NOR4 (N743, N735, N48, N190, N534);
xor XOR2 (N744, N742, N309);
nand NAND2 (N745, N730, N697);
or OR4 (N746, N740, N415, N135, N1);
nor NOR4 (N747, N745, N368, N241, N13);
not NOT1 (N748, N743);
not NOT1 (N749, N741);
nand NAND2 (N750, N748, N28);
nor NOR3 (N751, N737, N126, N571);
or OR3 (N752, N750, N546, N527);
buf BUF1 (N753, N749);
nor NOR4 (N754, N752, N345, N678, N355);
or OR3 (N755, N729, N585, N484);
xor XOR2 (N756, N755, N403);
not NOT1 (N757, N756);
nand NAND3 (N758, N754, N571, N202);
not NOT1 (N759, N751);
xor XOR2 (N760, N759, N746);
and AND2 (N761, N27, N131);
and AND2 (N762, N761, N175);
or OR3 (N763, N706, N443, N358);
nor NOR3 (N764, N744, N180, N463);
not NOT1 (N765, N726);
not NOT1 (N766, N747);
nor NOR2 (N767, N764, N417);
or OR4 (N768, N762, N21, N254, N428);
nand NAND2 (N769, N757, N94);
nor NOR3 (N770, N765, N651, N10);
not NOT1 (N771, N767);
nand NAND3 (N772, N758, N708, N214);
buf BUF1 (N773, N763);
buf BUF1 (N774, N773);
nor NOR2 (N775, N774, N633);
nor NOR4 (N776, N768, N523, N686, N479);
xor XOR2 (N777, N771, N42);
nor NOR3 (N778, N760, N725, N538);
nor NOR3 (N779, N772, N423, N305);
and AND2 (N780, N778, N178);
and AND2 (N781, N775, N606);
nand NAND3 (N782, N769, N2, N30);
buf BUF1 (N783, N738);
nor NOR3 (N784, N766, N757, N253);
and AND2 (N785, N753, N124);
and AND3 (N786, N770, N436, N711);
buf BUF1 (N787, N780);
xor XOR2 (N788, N787, N381);
buf BUF1 (N789, N776);
and AND4 (N790, N779, N274, N763, N310);
nor NOR3 (N791, N788, N606, N312);
nand NAND3 (N792, N790, N228, N393);
nor NOR3 (N793, N782, N532, N103);
nand NAND3 (N794, N781, N73, N583);
not NOT1 (N795, N783);
nor NOR4 (N796, N777, N565, N613, N151);
and AND4 (N797, N785, N306, N623, N295);
xor XOR2 (N798, N791, N53);
buf BUF1 (N799, N794);
nor NOR3 (N800, N799, N278, N587);
not NOT1 (N801, N793);
xor XOR2 (N802, N789, N75);
and AND2 (N803, N795, N253);
and AND3 (N804, N803, N27, N576);
not NOT1 (N805, N792);
buf BUF1 (N806, N796);
not NOT1 (N807, N804);
xor XOR2 (N808, N806, N584);
or OR3 (N809, N784, N775, N544);
nand NAND3 (N810, N802, N447, N2);
or OR2 (N811, N797, N484);
and AND3 (N812, N800, N176, N277);
nor NOR4 (N813, N801, N110, N436, N225);
and AND2 (N814, N813, N587);
not NOT1 (N815, N798);
nor NOR4 (N816, N814, N1, N679, N511);
nor NOR3 (N817, N786, N189, N435);
not NOT1 (N818, N805);
not NOT1 (N819, N817);
xor XOR2 (N820, N819, N548);
or OR3 (N821, N816, N521, N517);
nor NOR2 (N822, N815, N600);
not NOT1 (N823, N811);
and AND2 (N824, N821, N562);
buf BUF1 (N825, N823);
nor NOR4 (N826, N809, N353, N154, N719);
xor XOR2 (N827, N807, N558);
nand NAND2 (N828, N825, N65);
or OR3 (N829, N822, N580, N183);
xor XOR2 (N830, N827, N360);
xor XOR2 (N831, N826, N23);
and AND2 (N832, N831, N68);
nor NOR4 (N833, N810, N548, N329, N506);
or OR2 (N834, N833, N162);
and AND4 (N835, N830, N522, N201, N390);
buf BUF1 (N836, N812);
or OR3 (N837, N829, N792, N216);
buf BUF1 (N838, N808);
nor NOR3 (N839, N818, N738, N660);
not NOT1 (N840, N835);
nand NAND4 (N841, N839, N355, N305, N513);
buf BUF1 (N842, N837);
nand NAND3 (N843, N836, N312, N473);
not NOT1 (N844, N832);
not NOT1 (N845, N844);
or OR3 (N846, N820, N383, N347);
nor NOR3 (N847, N838, N165, N241);
nand NAND2 (N848, N843, N282);
not NOT1 (N849, N842);
nand NAND3 (N850, N841, N125, N731);
or OR4 (N851, N846, N816, N86, N771);
not NOT1 (N852, N840);
buf BUF1 (N853, N851);
and AND2 (N854, N828, N131);
nand NAND3 (N855, N847, N449, N351);
not NOT1 (N856, N853);
or OR2 (N857, N855, N649);
or OR4 (N858, N854, N478, N543, N461);
nor NOR2 (N859, N848, N168);
buf BUF1 (N860, N859);
not NOT1 (N861, N849);
buf BUF1 (N862, N852);
and AND4 (N863, N858, N204, N491, N704);
not NOT1 (N864, N861);
and AND4 (N865, N864, N852, N773, N389);
nand NAND2 (N866, N856, N566);
buf BUF1 (N867, N863);
not NOT1 (N868, N865);
nor NOR2 (N869, N850, N386);
xor XOR2 (N870, N824, N82);
xor XOR2 (N871, N857, N115);
xor XOR2 (N872, N869, N417);
nand NAND2 (N873, N871, N209);
and AND4 (N874, N860, N597, N266, N161);
xor XOR2 (N875, N873, N183);
xor XOR2 (N876, N875, N94);
not NOT1 (N877, N868);
xor XOR2 (N878, N870, N506);
and AND3 (N879, N866, N439, N21);
nor NOR3 (N880, N834, N590, N561);
nor NOR4 (N881, N877, N332, N500, N547);
nand NAND3 (N882, N862, N76, N38);
buf BUF1 (N883, N880);
or OR3 (N884, N876, N848, N121);
or OR3 (N885, N867, N331, N849);
buf BUF1 (N886, N881);
not NOT1 (N887, N882);
xor XOR2 (N888, N886, N790);
or OR3 (N889, N883, N355, N318);
nor NOR3 (N890, N872, N871, N332);
not NOT1 (N891, N884);
nor NOR3 (N892, N888, N851, N52);
nor NOR3 (N893, N887, N185, N64);
xor XOR2 (N894, N893, N873);
or OR2 (N895, N845, N615);
nor NOR3 (N896, N892, N796, N429);
nand NAND2 (N897, N889, N486);
not NOT1 (N898, N879);
nand NAND4 (N899, N897, N708, N313, N844);
buf BUF1 (N900, N899);
not NOT1 (N901, N891);
not NOT1 (N902, N900);
nor NOR2 (N903, N898, N116);
nor NOR2 (N904, N902, N1);
or OR2 (N905, N885, N723);
and AND2 (N906, N904, N766);
xor XOR2 (N907, N903, N523);
buf BUF1 (N908, N894);
or OR3 (N909, N895, N765, N562);
xor XOR2 (N910, N890, N522);
buf BUF1 (N911, N910);
xor XOR2 (N912, N878, N734);
xor XOR2 (N913, N905, N338);
or OR4 (N914, N896, N287, N778, N62);
nor NOR4 (N915, N914, N462, N898, N60);
nor NOR2 (N916, N907, N707);
and AND3 (N917, N901, N333, N824);
nand NAND3 (N918, N874, N650, N493);
buf BUF1 (N919, N911);
and AND2 (N920, N906, N154);
or OR2 (N921, N909, N664);
buf BUF1 (N922, N921);
nor NOR4 (N923, N912, N292, N431, N273);
and AND4 (N924, N919, N449, N454, N903);
or OR4 (N925, N920, N455, N104, N223);
not NOT1 (N926, N908);
xor XOR2 (N927, N925, N27);
buf BUF1 (N928, N913);
nor NOR2 (N929, N923, N375);
not NOT1 (N930, N924);
not NOT1 (N931, N915);
not NOT1 (N932, N929);
buf BUF1 (N933, N922);
not NOT1 (N934, N928);
and AND4 (N935, N932, N40, N860, N463);
xor XOR2 (N936, N934, N39);
not NOT1 (N937, N916);
not NOT1 (N938, N933);
xor XOR2 (N939, N927, N121);
buf BUF1 (N940, N931);
and AND3 (N941, N935, N389, N834);
nor NOR3 (N942, N940, N932, N707);
and AND4 (N943, N918, N798, N793, N755);
and AND2 (N944, N937, N720);
xor XOR2 (N945, N943, N516);
not NOT1 (N946, N944);
or OR2 (N947, N938, N271);
buf BUF1 (N948, N942);
or OR2 (N949, N947, N379);
and AND4 (N950, N936, N129, N607, N519);
buf BUF1 (N951, N949);
not NOT1 (N952, N930);
not NOT1 (N953, N939);
buf BUF1 (N954, N951);
xor XOR2 (N955, N941, N86);
buf BUF1 (N956, N952);
buf BUF1 (N957, N954);
xor XOR2 (N958, N956, N718);
and AND2 (N959, N948, N766);
xor XOR2 (N960, N953, N571);
nor NOR2 (N961, N945, N438);
and AND2 (N962, N958, N559);
xor XOR2 (N963, N962, N204);
and AND2 (N964, N946, N51);
not NOT1 (N965, N964);
or OR4 (N966, N959, N525, N66, N421);
not NOT1 (N967, N957);
nor NOR2 (N968, N960, N757);
nor NOR3 (N969, N963, N531, N398);
buf BUF1 (N970, N917);
xor XOR2 (N971, N967, N773);
and AND2 (N972, N969, N306);
buf BUF1 (N973, N961);
nor NOR2 (N974, N968, N544);
or OR2 (N975, N971, N880);
nor NOR3 (N976, N955, N446, N162);
buf BUF1 (N977, N975);
or OR4 (N978, N973, N205, N792, N115);
nand NAND3 (N979, N978, N837, N367);
nand NAND3 (N980, N950, N952, N471);
not NOT1 (N981, N979);
not NOT1 (N982, N926);
nand NAND3 (N983, N974, N458, N914);
or OR4 (N984, N982, N722, N862, N510);
or OR2 (N985, N972, N493);
not NOT1 (N986, N977);
xor XOR2 (N987, N986, N133);
buf BUF1 (N988, N981);
or OR4 (N989, N976, N317, N669, N756);
xor XOR2 (N990, N984, N299);
buf BUF1 (N991, N988);
and AND4 (N992, N987, N929, N556, N752);
xor XOR2 (N993, N980, N850);
buf BUF1 (N994, N993);
or OR2 (N995, N983, N723);
nor NOR4 (N996, N965, N314, N14, N3);
xor XOR2 (N997, N992, N249);
buf BUF1 (N998, N970);
or OR3 (N999, N989, N517, N831);
buf BUF1 (N1000, N991);
buf BUF1 (N1001, N998);
nand NAND3 (N1002, N997, N646, N880);
nand NAND2 (N1003, N994, N438);
or OR3 (N1004, N1000, N728, N683);
buf BUF1 (N1005, N990);
or OR4 (N1006, N999, N839, N565, N354);
not NOT1 (N1007, N1005);
not NOT1 (N1008, N1003);
nor NOR3 (N1009, N966, N848, N241);
and AND2 (N1010, N1001, N131);
or OR4 (N1011, N995, N912, N507, N826);
or OR4 (N1012, N996, N671, N287, N906);
not NOT1 (N1013, N1006);
or OR4 (N1014, N985, N25, N843, N851);
not NOT1 (N1015, N1012);
and AND3 (N1016, N1004, N582, N434);
nand NAND3 (N1017, N1014, N634, N368);
nand NAND4 (N1018, N1002, N881, N158, N887);
buf BUF1 (N1019, N1007);
nand NAND4 (N1020, N1011, N310, N117, N832);
buf BUF1 (N1021, N1015);
not NOT1 (N1022, N1013);
nor NOR2 (N1023, N1020, N352);
and AND3 (N1024, N1023, N269, N870);
not NOT1 (N1025, N1008);
or OR3 (N1026, N1016, N669, N477);
nand NAND3 (N1027, N1017, N419, N55);
nor NOR3 (N1028, N1025, N500, N870);
not NOT1 (N1029, N1021);
nand NAND3 (N1030, N1010, N786, N930);
or OR2 (N1031, N1009, N695);
or OR2 (N1032, N1031, N73);
nand NAND2 (N1033, N1022, N554);
xor XOR2 (N1034, N1018, N638);
nor NOR2 (N1035, N1033, N931);
buf BUF1 (N1036, N1026);
nor NOR2 (N1037, N1035, N946);
not NOT1 (N1038, N1029);
nor NOR4 (N1039, N1019, N75, N721, N548);
xor XOR2 (N1040, N1028, N315);
not NOT1 (N1041, N1039);
nor NOR3 (N1042, N1036, N664, N393);
xor XOR2 (N1043, N1041, N909);
xor XOR2 (N1044, N1043, N798);
xor XOR2 (N1045, N1034, N112);
not NOT1 (N1046, N1027);
and AND2 (N1047, N1032, N51);
or OR3 (N1048, N1040, N349, N192);
buf BUF1 (N1049, N1048);
not NOT1 (N1050, N1045);
xor XOR2 (N1051, N1049, N490);
and AND3 (N1052, N1044, N133, N986);
nor NOR2 (N1053, N1038, N225);
and AND2 (N1054, N1030, N815);
or OR4 (N1055, N1024, N423, N985, N856);
buf BUF1 (N1056, N1037);
and AND3 (N1057, N1053, N87, N644);
nor NOR3 (N1058, N1054, N88, N110);
and AND4 (N1059, N1047, N470, N427, N353);
buf BUF1 (N1060, N1057);
or OR2 (N1061, N1059, N423);
not NOT1 (N1062, N1055);
not NOT1 (N1063, N1062);
and AND4 (N1064, N1051, N478, N556, N108);
not NOT1 (N1065, N1052);
or OR2 (N1066, N1060, N643);
nand NAND3 (N1067, N1056, N789, N377);
buf BUF1 (N1068, N1058);
or OR4 (N1069, N1067, N900, N58, N224);
not NOT1 (N1070, N1064);
xor XOR2 (N1071, N1066, N294);
xor XOR2 (N1072, N1063, N368);
xor XOR2 (N1073, N1046, N776);
nand NAND4 (N1074, N1073, N235, N139, N449);
nor NOR2 (N1075, N1072, N425);
nor NOR4 (N1076, N1068, N464, N473, N867);
xor XOR2 (N1077, N1071, N593);
nand NAND2 (N1078, N1061, N78);
not NOT1 (N1079, N1078);
and AND4 (N1080, N1076, N644, N677, N207);
or OR4 (N1081, N1070, N757, N382, N649);
nor NOR3 (N1082, N1050, N177, N873);
nand NAND3 (N1083, N1042, N541, N121);
buf BUF1 (N1084, N1074);
xor XOR2 (N1085, N1069, N125);
xor XOR2 (N1086, N1081, N264);
nand NAND4 (N1087, N1075, N364, N363, N885);
buf BUF1 (N1088, N1085);
or OR3 (N1089, N1082, N127, N960);
not NOT1 (N1090, N1086);
and AND2 (N1091, N1087, N162);
nand NAND4 (N1092, N1079, N808, N738, N805);
not NOT1 (N1093, N1084);
or OR3 (N1094, N1091, N506, N708);
buf BUF1 (N1095, N1083);
and AND2 (N1096, N1095, N342);
nor NOR2 (N1097, N1077, N417);
nor NOR3 (N1098, N1092, N806, N741);
nand NAND4 (N1099, N1065, N1018, N337, N518);
nand NAND3 (N1100, N1098, N488, N135);
and AND3 (N1101, N1096, N87, N264);
and AND2 (N1102, N1093, N284);
nor NOR2 (N1103, N1080, N535);
or OR2 (N1104, N1103, N888);
and AND4 (N1105, N1090, N119, N307, N282);
xor XOR2 (N1106, N1088, N931);
not NOT1 (N1107, N1102);
and AND2 (N1108, N1101, N904);
buf BUF1 (N1109, N1099);
and AND3 (N1110, N1106, N965, N518);
xor XOR2 (N1111, N1109, N711);
not NOT1 (N1112, N1105);
xor XOR2 (N1113, N1104, N390);
nor NOR2 (N1114, N1112, N341);
not NOT1 (N1115, N1089);
buf BUF1 (N1116, N1110);
nor NOR3 (N1117, N1111, N449, N142);
buf BUF1 (N1118, N1116);
nor NOR2 (N1119, N1115, N741);
and AND4 (N1120, N1114, N951, N1040, N719);
nor NOR4 (N1121, N1107, N293, N533, N699);
not NOT1 (N1122, N1120);
and AND2 (N1123, N1100, N343);
nand NAND3 (N1124, N1097, N762, N725);
xor XOR2 (N1125, N1118, N987);
nand NAND2 (N1126, N1117, N490);
xor XOR2 (N1127, N1122, N827);
buf BUF1 (N1128, N1119);
and AND4 (N1129, N1124, N244, N340, N961);
buf BUF1 (N1130, N1127);
nor NOR4 (N1131, N1123, N404, N767, N91);
nand NAND2 (N1132, N1129, N868);
and AND3 (N1133, N1131, N512, N133);
and AND2 (N1134, N1125, N672);
and AND3 (N1135, N1132, N64, N1067);
nor NOR4 (N1136, N1134, N311, N409, N323);
buf BUF1 (N1137, N1121);
buf BUF1 (N1138, N1135);
xor XOR2 (N1139, N1094, N70);
not NOT1 (N1140, N1133);
xor XOR2 (N1141, N1136, N741);
xor XOR2 (N1142, N1108, N991);
not NOT1 (N1143, N1128);
xor XOR2 (N1144, N1126, N1057);
and AND2 (N1145, N1113, N601);
and AND3 (N1146, N1138, N250, N1069);
buf BUF1 (N1147, N1137);
or OR4 (N1148, N1147, N420, N773, N898);
or OR4 (N1149, N1141, N375, N423, N372);
not NOT1 (N1150, N1130);
xor XOR2 (N1151, N1143, N932);
nand NAND2 (N1152, N1151, N789);
and AND4 (N1153, N1139, N12, N670, N1094);
nand NAND4 (N1154, N1150, N131, N1105, N926);
nor NOR4 (N1155, N1153, N327, N333, N589);
nand NAND3 (N1156, N1144, N860, N34);
nand NAND2 (N1157, N1145, N1090);
buf BUF1 (N1158, N1148);
nor NOR2 (N1159, N1146, N918);
and AND2 (N1160, N1157, N1081);
and AND2 (N1161, N1142, N14);
buf BUF1 (N1162, N1158);
buf BUF1 (N1163, N1140);
nor NOR3 (N1164, N1155, N277, N828);
not NOT1 (N1165, N1161);
nand NAND2 (N1166, N1159, N74);
and AND4 (N1167, N1154, N813, N244, N113);
nand NAND3 (N1168, N1160, N415, N611);
not NOT1 (N1169, N1164);
xor XOR2 (N1170, N1162, N46);
nor NOR2 (N1171, N1163, N1132);
not NOT1 (N1172, N1149);
or OR3 (N1173, N1172, N188, N1080);
or OR3 (N1174, N1167, N218, N718);
xor XOR2 (N1175, N1169, N1013);
xor XOR2 (N1176, N1156, N101);
buf BUF1 (N1177, N1152);
xor XOR2 (N1178, N1176, N974);
not NOT1 (N1179, N1166);
not NOT1 (N1180, N1173);
not NOT1 (N1181, N1175);
xor XOR2 (N1182, N1165, N1098);
nand NAND4 (N1183, N1170, N437, N1103, N164);
buf BUF1 (N1184, N1168);
not NOT1 (N1185, N1183);
or OR2 (N1186, N1178, N1181);
or OR4 (N1187, N221, N826, N971, N490);
not NOT1 (N1188, N1185);
not NOT1 (N1189, N1188);
not NOT1 (N1190, N1182);
and AND2 (N1191, N1179, N1030);
xor XOR2 (N1192, N1177, N634);
and AND4 (N1193, N1190, N697, N38, N185);
xor XOR2 (N1194, N1186, N1166);
xor XOR2 (N1195, N1171, N1189);
not NOT1 (N1196, N695);
buf BUF1 (N1197, N1194);
not NOT1 (N1198, N1197);
or OR2 (N1199, N1192, N365);
nand NAND4 (N1200, N1198, N529, N444, N366);
xor XOR2 (N1201, N1199, N490);
buf BUF1 (N1202, N1196);
nor NOR2 (N1203, N1195, N389);
or OR3 (N1204, N1200, N1100, N11);
and AND4 (N1205, N1191, N417, N663, N774);
or OR2 (N1206, N1187, N792);
xor XOR2 (N1207, N1202, N1033);
buf BUF1 (N1208, N1174);
nor NOR3 (N1209, N1180, N265, N709);
or OR3 (N1210, N1208, N552, N224);
or OR3 (N1211, N1201, N947, N1192);
not NOT1 (N1212, N1209);
and AND3 (N1213, N1193, N549, N410);
not NOT1 (N1214, N1207);
buf BUF1 (N1215, N1214);
xor XOR2 (N1216, N1211, N329);
nor NOR4 (N1217, N1216, N379, N73, N561);
or OR2 (N1218, N1210, N339);
buf BUF1 (N1219, N1184);
xor XOR2 (N1220, N1206, N320);
xor XOR2 (N1221, N1205, N141);
xor XOR2 (N1222, N1219, N434);
nor NOR2 (N1223, N1204, N13);
buf BUF1 (N1224, N1213);
or OR2 (N1225, N1215, N560);
xor XOR2 (N1226, N1225, N395);
buf BUF1 (N1227, N1217);
nor NOR2 (N1228, N1222, N654);
and AND3 (N1229, N1218, N642, N692);
nand NAND2 (N1230, N1212, N1099);
nand NAND2 (N1231, N1223, N621);
nand NAND3 (N1232, N1221, N304, N55);
and AND4 (N1233, N1230, N70, N38, N661);
or OR4 (N1234, N1226, N68, N1160, N544);
xor XOR2 (N1235, N1234, N225);
xor XOR2 (N1236, N1229, N2);
nor NOR2 (N1237, N1236, N488);
nand NAND3 (N1238, N1233, N959, N716);
nand NAND3 (N1239, N1235, N1052, N382);
or OR3 (N1240, N1238, N905, N502);
xor XOR2 (N1241, N1227, N39);
buf BUF1 (N1242, N1203);
and AND4 (N1243, N1239, N529, N725, N530);
not NOT1 (N1244, N1242);
and AND2 (N1245, N1224, N985);
xor XOR2 (N1246, N1244, N1123);
or OR2 (N1247, N1241, N1174);
nand NAND2 (N1248, N1228, N421);
xor XOR2 (N1249, N1248, N793);
or OR3 (N1250, N1232, N1099, N1031);
and AND4 (N1251, N1247, N9, N1066, N993);
nor NOR3 (N1252, N1250, N950, N558);
xor XOR2 (N1253, N1220, N1123);
and AND2 (N1254, N1237, N153);
and AND3 (N1255, N1245, N1170, N417);
xor XOR2 (N1256, N1253, N1039);
xor XOR2 (N1257, N1231, N873);
xor XOR2 (N1258, N1240, N696);
xor XOR2 (N1259, N1246, N230);
nor NOR4 (N1260, N1257, N155, N219, N412);
buf BUF1 (N1261, N1251);
xor XOR2 (N1262, N1261, N372);
or OR4 (N1263, N1255, N1197, N470, N437);
not NOT1 (N1264, N1263);
and AND4 (N1265, N1254, N585, N610, N974);
nand NAND4 (N1266, N1249, N806, N346, N1189);
buf BUF1 (N1267, N1260);
and AND3 (N1268, N1258, N106, N736);
or OR2 (N1269, N1266, N1133);
or OR3 (N1270, N1264, N781, N1224);
nand NAND4 (N1271, N1270, N1124, N521, N172);
and AND3 (N1272, N1256, N295, N928);
buf BUF1 (N1273, N1272);
nand NAND4 (N1274, N1265, N32, N315, N353);
buf BUF1 (N1275, N1243);
nor NOR2 (N1276, N1259, N839);
xor XOR2 (N1277, N1271, N1003);
buf BUF1 (N1278, N1276);
xor XOR2 (N1279, N1269, N902);
nand NAND4 (N1280, N1278, N778, N328, N2);
and AND3 (N1281, N1268, N920, N1244);
xor XOR2 (N1282, N1277, N937);
buf BUF1 (N1283, N1279);
not NOT1 (N1284, N1275);
or OR4 (N1285, N1281, N1209, N1189, N962);
xor XOR2 (N1286, N1267, N232);
xor XOR2 (N1287, N1285, N18);
or OR2 (N1288, N1284, N366);
nor NOR4 (N1289, N1252, N168, N939, N1174);
and AND4 (N1290, N1282, N1204, N1162, N512);
nand NAND2 (N1291, N1280, N834);
or OR3 (N1292, N1274, N763, N604);
buf BUF1 (N1293, N1292);
nand NAND3 (N1294, N1289, N48, N198);
nor NOR4 (N1295, N1294, N381, N664, N21);
or OR4 (N1296, N1295, N325, N469, N32);
and AND4 (N1297, N1262, N634, N603, N162);
nor NOR4 (N1298, N1296, N468, N789, N334);
nor NOR3 (N1299, N1297, N478, N400);
xor XOR2 (N1300, N1299, N239);
not NOT1 (N1301, N1287);
nor NOR4 (N1302, N1288, N404, N668, N774);
and AND3 (N1303, N1301, N455, N1062);
buf BUF1 (N1304, N1303);
and AND2 (N1305, N1286, N348);
xor XOR2 (N1306, N1290, N228);
nand NAND2 (N1307, N1305, N667);
nor NOR2 (N1308, N1283, N913);
or OR4 (N1309, N1306, N1130, N206, N671);
and AND4 (N1310, N1309, N1175, N734, N936);
and AND2 (N1311, N1302, N1307);
or OR2 (N1312, N936, N995);
buf BUF1 (N1313, N1300);
and AND2 (N1314, N1310, N1178);
and AND4 (N1315, N1304, N498, N125, N255);
xor XOR2 (N1316, N1308, N714);
not NOT1 (N1317, N1312);
nand NAND4 (N1318, N1273, N1297, N427, N1021);
or OR4 (N1319, N1317, N88, N526, N247);
nor NOR4 (N1320, N1313, N485, N182, N1193);
xor XOR2 (N1321, N1314, N468);
nor NOR3 (N1322, N1319, N360, N375);
buf BUF1 (N1323, N1320);
or OR3 (N1324, N1321, N1111, N187);
nor NOR4 (N1325, N1315, N742, N1150, N319);
not NOT1 (N1326, N1325);
and AND4 (N1327, N1293, N321, N1136, N1145);
or OR3 (N1328, N1316, N63, N1089);
xor XOR2 (N1329, N1323, N658);
and AND2 (N1330, N1298, N404);
not NOT1 (N1331, N1318);
or OR3 (N1332, N1328, N1061, N986);
buf BUF1 (N1333, N1326);
nand NAND2 (N1334, N1322, N198);
or OR4 (N1335, N1332, N587, N489, N724);
not NOT1 (N1336, N1329);
buf BUF1 (N1337, N1330);
and AND2 (N1338, N1331, N716);
xor XOR2 (N1339, N1327, N810);
xor XOR2 (N1340, N1333, N1296);
nand NAND3 (N1341, N1324, N1152, N357);
buf BUF1 (N1342, N1335);
not NOT1 (N1343, N1342);
or OR4 (N1344, N1291, N4, N232, N624);
xor XOR2 (N1345, N1340, N823);
and AND4 (N1346, N1345, N1220, N1184, N753);
not NOT1 (N1347, N1336);
or OR4 (N1348, N1343, N571, N1346, N651);
or OR3 (N1349, N613, N694, N1099);
xor XOR2 (N1350, N1338, N286);
and AND4 (N1351, N1348, N495, N929, N854);
nor NOR2 (N1352, N1347, N688);
or OR3 (N1353, N1349, N1044, N77);
xor XOR2 (N1354, N1341, N491);
nor NOR2 (N1355, N1353, N985);
nand NAND2 (N1356, N1311, N176);
nand NAND3 (N1357, N1339, N718, N616);
buf BUF1 (N1358, N1350);
or OR2 (N1359, N1356, N27);
buf BUF1 (N1360, N1358);
not NOT1 (N1361, N1357);
nand NAND4 (N1362, N1360, N646, N394, N137);
xor XOR2 (N1363, N1344, N1170);
or OR2 (N1364, N1351, N1094);
and AND4 (N1365, N1355, N1307, N571, N963);
xor XOR2 (N1366, N1334, N530);
or OR4 (N1367, N1352, N1216, N1249, N307);
buf BUF1 (N1368, N1359);
or OR3 (N1369, N1367, N315, N1182);
nand NAND2 (N1370, N1337, N2);
buf BUF1 (N1371, N1370);
nor NOR4 (N1372, N1371, N1284, N2, N1317);
nor NOR3 (N1373, N1363, N215, N955);
xor XOR2 (N1374, N1362, N366);
nor NOR4 (N1375, N1365, N339, N758, N1091);
nor NOR4 (N1376, N1374, N1208, N504, N369);
not NOT1 (N1377, N1373);
not NOT1 (N1378, N1364);
nand NAND3 (N1379, N1368, N528, N868);
or OR4 (N1380, N1375, N1015, N95, N641);
or OR2 (N1381, N1377, N392);
buf BUF1 (N1382, N1378);
xor XOR2 (N1383, N1382, N45);
nand NAND4 (N1384, N1381, N1200, N1277, N83);
and AND2 (N1385, N1383, N120);
nand NAND4 (N1386, N1372, N122, N1361, N1180);
and AND2 (N1387, N1180, N1060);
and AND3 (N1388, N1379, N118, N804);
or OR3 (N1389, N1388, N459, N1184);
xor XOR2 (N1390, N1366, N1269);
and AND3 (N1391, N1369, N429, N343);
xor XOR2 (N1392, N1380, N552);
and AND2 (N1393, N1385, N669);
nand NAND3 (N1394, N1390, N1372, N890);
or OR3 (N1395, N1386, N13, N1226);
nand NAND2 (N1396, N1394, N741);
or OR2 (N1397, N1376, N799);
and AND2 (N1398, N1396, N109);
xor XOR2 (N1399, N1354, N949);
and AND4 (N1400, N1399, N887, N843, N712);
nor NOR3 (N1401, N1395, N627, N856);
buf BUF1 (N1402, N1401);
xor XOR2 (N1403, N1400, N304);
or OR3 (N1404, N1384, N711, N2);
not NOT1 (N1405, N1398);
buf BUF1 (N1406, N1397);
and AND3 (N1407, N1403, N64, N475);
and AND3 (N1408, N1393, N1212, N891);
not NOT1 (N1409, N1405);
or OR3 (N1410, N1387, N72, N792);
and AND4 (N1411, N1406, N172, N1382, N321);
or OR3 (N1412, N1391, N1160, N399);
or OR4 (N1413, N1411, N1173, N397, N19);
and AND3 (N1414, N1409, N552, N416);
nor NOR4 (N1415, N1412, N919, N1067, N229);
buf BUF1 (N1416, N1408);
or OR2 (N1417, N1392, N100);
or OR2 (N1418, N1416, N237);
not NOT1 (N1419, N1418);
nor NOR4 (N1420, N1410, N86, N849, N859);
buf BUF1 (N1421, N1407);
and AND2 (N1422, N1419, N581);
or OR2 (N1423, N1420, N249);
or OR4 (N1424, N1402, N1322, N1322, N1144);
or OR4 (N1425, N1424, N152, N1270, N1251);
buf BUF1 (N1426, N1414);
or OR4 (N1427, N1404, N175, N1359, N423);
or OR3 (N1428, N1425, N1029, N1100);
buf BUF1 (N1429, N1426);
buf BUF1 (N1430, N1389);
buf BUF1 (N1431, N1413);
xor XOR2 (N1432, N1428, N514);
nor NOR4 (N1433, N1430, N635, N733, N876);
buf BUF1 (N1434, N1417);
not NOT1 (N1435, N1421);
or OR3 (N1436, N1434, N1432, N103);
xor XOR2 (N1437, N173, N1041);
or OR2 (N1438, N1437, N1076);
and AND2 (N1439, N1438, N1212);
not NOT1 (N1440, N1439);
nand NAND3 (N1441, N1429, N970, N1229);
xor XOR2 (N1442, N1433, N1313);
or OR4 (N1443, N1422, N1431, N837, N1219);
not NOT1 (N1444, N1157);
and AND2 (N1445, N1427, N182);
nand NAND4 (N1446, N1441, N426, N299, N477);
and AND3 (N1447, N1440, N351, N553);
not NOT1 (N1448, N1423);
nand NAND2 (N1449, N1435, N716);
or OR2 (N1450, N1442, N1273);
buf BUF1 (N1451, N1449);
buf BUF1 (N1452, N1450);
buf BUF1 (N1453, N1415);
or OR2 (N1454, N1443, N779);
xor XOR2 (N1455, N1436, N1364);
and AND2 (N1456, N1455, N779);
nand NAND2 (N1457, N1451, N407);
not NOT1 (N1458, N1448);
xor XOR2 (N1459, N1446, N1055);
and AND2 (N1460, N1458, N542);
buf BUF1 (N1461, N1457);
nor NOR3 (N1462, N1453, N1314, N708);
or OR2 (N1463, N1459, N142);
and AND2 (N1464, N1461, N1039);
or OR4 (N1465, N1462, N1414, N887, N1219);
xor XOR2 (N1466, N1445, N400);
buf BUF1 (N1467, N1447);
xor XOR2 (N1468, N1465, N947);
not NOT1 (N1469, N1456);
xor XOR2 (N1470, N1454, N75);
nand NAND3 (N1471, N1470, N1374, N211);
nand NAND4 (N1472, N1460, N1161, N1207, N1204);
nor NOR3 (N1473, N1468, N1185, N241);
and AND2 (N1474, N1467, N188);
nor NOR2 (N1475, N1463, N975);
nand NAND4 (N1476, N1473, N1115, N469, N206);
nor NOR2 (N1477, N1472, N1255);
and AND4 (N1478, N1477, N153, N667, N139);
and AND2 (N1479, N1444, N1465);
buf BUF1 (N1480, N1479);
and AND3 (N1481, N1452, N965, N1367);
or OR3 (N1482, N1481, N376, N142);
not NOT1 (N1483, N1476);
nand NAND2 (N1484, N1483, N297);
and AND2 (N1485, N1475, N308);
buf BUF1 (N1486, N1478);
nor NOR3 (N1487, N1485, N1042, N105);
and AND2 (N1488, N1474, N1069);
and AND2 (N1489, N1482, N1109);
buf BUF1 (N1490, N1469);
or OR3 (N1491, N1486, N1201, N658);
nand NAND2 (N1492, N1484, N1393);
or OR3 (N1493, N1491, N165, N925);
xor XOR2 (N1494, N1492, N561);
not NOT1 (N1495, N1464);
not NOT1 (N1496, N1489);
not NOT1 (N1497, N1471);
buf BUF1 (N1498, N1488);
nand NAND3 (N1499, N1495, N895, N1227);
nor NOR4 (N1500, N1498, N388, N715, N260);
buf BUF1 (N1501, N1490);
nand NAND2 (N1502, N1497, N150);
nor NOR4 (N1503, N1499, N974, N454, N540);
nor NOR2 (N1504, N1487, N843);
buf BUF1 (N1505, N1504);
and AND3 (N1506, N1503, N1067, N1313);
nand NAND2 (N1507, N1496, N1236);
nand NAND3 (N1508, N1501, N695, N457);
not NOT1 (N1509, N1507);
buf BUF1 (N1510, N1505);
nand NAND3 (N1511, N1509, N594, N1180);
buf BUF1 (N1512, N1480);
not NOT1 (N1513, N1500);
or OR4 (N1514, N1494, N80, N724, N385);
nor NOR4 (N1515, N1502, N757, N635, N1191);
nor NOR2 (N1516, N1515, N768);
xor XOR2 (N1517, N1511, N24);
not NOT1 (N1518, N1510);
nand NAND4 (N1519, N1506, N1298, N1036, N371);
buf BUF1 (N1520, N1518);
buf BUF1 (N1521, N1513);
nor NOR3 (N1522, N1516, N50, N1455);
nand NAND4 (N1523, N1466, N1057, N83, N949);
nor NOR3 (N1524, N1493, N1234, N203);
endmodule