// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N620,N609,N614,N618,N621,N611,N613,N607,N619,N622;

xor XOR2 (N23, N11, N9);
or OR2 (N24, N5, N3);
and AND2 (N25, N8, N24);
xor XOR2 (N26, N22, N14);
buf BUF1 (N27, N24);
not NOT1 (N28, N25);
xor XOR2 (N29, N22, N14);
xor XOR2 (N30, N1, N10);
buf BUF1 (N31, N3);
or OR4 (N32, N14, N31, N22, N13);
nand NAND4 (N33, N10, N31, N17, N23);
buf BUF1 (N34, N23);
not NOT1 (N35, N24);
buf BUF1 (N36, N5);
buf BUF1 (N37, N35);
and AND3 (N38, N33, N9, N23);
or OR3 (N39, N30, N8, N26);
xor XOR2 (N40, N12, N1);
xor XOR2 (N41, N28, N24);
and AND2 (N42, N27, N8);
xor XOR2 (N43, N41, N30);
nand NAND4 (N44, N43, N26, N12, N35);
nand NAND4 (N45, N37, N13, N12, N10);
not NOT1 (N46, N29);
nor NOR2 (N47, N36, N45);
buf BUF1 (N48, N22);
nor NOR2 (N49, N34, N41);
buf BUF1 (N50, N46);
or OR3 (N51, N38, N5, N7);
xor XOR2 (N52, N51, N29);
nor NOR3 (N53, N40, N37, N1);
not NOT1 (N54, N52);
nor NOR3 (N55, N53, N45, N30);
and AND2 (N56, N55, N31);
and AND2 (N57, N48, N51);
not NOT1 (N58, N49);
or OR3 (N59, N32, N29, N32);
buf BUF1 (N60, N47);
nor NOR3 (N61, N50, N3, N15);
nand NAND4 (N62, N42, N44, N13, N19);
buf BUF1 (N63, N10);
buf BUF1 (N64, N59);
not NOT1 (N65, N60);
xor XOR2 (N66, N39, N10);
nor NOR2 (N67, N56, N32);
nor NOR2 (N68, N64, N42);
or OR4 (N69, N62, N15, N25, N30);
buf BUF1 (N70, N58);
buf BUF1 (N71, N65);
not NOT1 (N72, N69);
buf BUF1 (N73, N57);
buf BUF1 (N74, N73);
or OR2 (N75, N71, N41);
buf BUF1 (N76, N54);
not NOT1 (N77, N76);
buf BUF1 (N78, N77);
nand NAND4 (N79, N75, N75, N10, N57);
xor XOR2 (N80, N70, N20);
nand NAND3 (N81, N68, N27, N71);
buf BUF1 (N82, N72);
or OR4 (N83, N80, N17, N45, N27);
buf BUF1 (N84, N81);
xor XOR2 (N85, N78, N37);
or OR4 (N86, N74, N57, N16, N3);
and AND4 (N87, N83, N66, N6, N68);
buf BUF1 (N88, N4);
nor NOR4 (N89, N86, N10, N20, N71);
nand NAND2 (N90, N63, N13);
or OR3 (N91, N67, N31, N25);
or OR2 (N92, N89, N91);
not NOT1 (N93, N62);
and AND4 (N94, N61, N17, N76, N40);
or OR4 (N95, N87, N47, N14, N48);
and AND4 (N96, N93, N44, N30, N30);
and AND3 (N97, N92, N56, N5);
xor XOR2 (N98, N84, N25);
buf BUF1 (N99, N79);
nor NOR3 (N100, N98, N5, N60);
or OR2 (N101, N82, N46);
buf BUF1 (N102, N85);
and AND4 (N103, N90, N27, N86, N40);
not NOT1 (N104, N103);
not NOT1 (N105, N96);
nor NOR2 (N106, N101, N88);
and AND3 (N107, N94, N96, N37);
not NOT1 (N108, N40);
not NOT1 (N109, N106);
or OR4 (N110, N102, N25, N36, N77);
and AND4 (N111, N109, N97, N92, N91);
nand NAND2 (N112, N99, N40);
nor NOR4 (N113, N94, N95, N75, N57);
and AND4 (N114, N42, N72, N90, N109);
buf BUF1 (N115, N108);
and AND3 (N116, N112, N72, N84);
or OR4 (N117, N116, N72, N17, N25);
nor NOR4 (N118, N104, N39, N60, N94);
and AND2 (N119, N114, N77);
nand NAND3 (N120, N117, N95, N24);
buf BUF1 (N121, N111);
nand NAND3 (N122, N100, N44, N39);
buf BUF1 (N123, N118);
xor XOR2 (N124, N115, N86);
not NOT1 (N125, N122);
nor NOR4 (N126, N107, N81, N20, N72);
nor NOR3 (N127, N119, N40, N6);
buf BUF1 (N128, N124);
not NOT1 (N129, N125);
xor XOR2 (N130, N121, N40);
xor XOR2 (N131, N129, N107);
xor XOR2 (N132, N131, N118);
xor XOR2 (N133, N126, N31);
or OR4 (N134, N128, N115, N101, N89);
nand NAND4 (N135, N130, N72, N117, N119);
or OR4 (N136, N134, N133, N30, N83);
buf BUF1 (N137, N34);
nor NOR4 (N138, N113, N3, N45, N83);
nor NOR4 (N139, N123, N138, N114, N125);
buf BUF1 (N140, N87);
or OR3 (N141, N135, N112, N102);
and AND2 (N142, N127, N49);
nor NOR4 (N143, N139, N116, N138, N61);
nor NOR3 (N144, N136, N49, N6);
or OR2 (N145, N132, N31);
not NOT1 (N146, N110);
nand NAND2 (N147, N141, N10);
nor NOR3 (N148, N144, N113, N145);
not NOT1 (N149, N39);
nand NAND4 (N150, N148, N125, N110, N133);
xor XOR2 (N151, N142, N92);
not NOT1 (N152, N120);
nand NAND2 (N153, N140, N48);
not NOT1 (N154, N105);
and AND4 (N155, N150, N101, N102, N53);
buf BUF1 (N156, N152);
nand NAND3 (N157, N137, N130, N33);
and AND4 (N158, N154, N59, N150, N116);
or OR3 (N159, N143, N86, N25);
not NOT1 (N160, N146);
and AND2 (N161, N147, N19);
and AND4 (N162, N160, N31, N137, N84);
nor NOR3 (N163, N151, N124, N87);
xor XOR2 (N164, N162, N46);
not NOT1 (N165, N153);
xor XOR2 (N166, N158, N146);
or OR2 (N167, N159, N155);
nand NAND4 (N168, N77, N24, N2, N22);
not NOT1 (N169, N157);
and AND2 (N170, N167, N61);
buf BUF1 (N171, N168);
nand NAND2 (N172, N149, N49);
nor NOR2 (N173, N166, N13);
nand NAND4 (N174, N169, N17, N47, N43);
xor XOR2 (N175, N161, N81);
nor NOR4 (N176, N174, N81, N102, N102);
nand NAND3 (N177, N176, N125, N166);
nor NOR3 (N178, N165, N70, N173);
or OR3 (N179, N88, N128, N95);
not NOT1 (N180, N170);
nand NAND4 (N181, N178, N18, N33, N128);
buf BUF1 (N182, N163);
buf BUF1 (N183, N182);
nor NOR2 (N184, N177, N39);
and AND3 (N185, N183, N34, N179);
nand NAND2 (N186, N69, N43);
nor NOR4 (N187, N175, N186, N181, N45);
and AND2 (N188, N134, N115);
or OR4 (N189, N105, N153, N177, N29);
buf BUF1 (N190, N188);
buf BUF1 (N191, N184);
xor XOR2 (N192, N191, N165);
buf BUF1 (N193, N185);
not NOT1 (N194, N156);
nand NAND2 (N195, N189, N149);
xor XOR2 (N196, N164, N50);
buf BUF1 (N197, N194);
xor XOR2 (N198, N171, N37);
nand NAND3 (N199, N198, N197, N59);
not NOT1 (N200, N65);
not NOT1 (N201, N199);
buf BUF1 (N202, N201);
nor NOR2 (N203, N192, N74);
nor NOR4 (N204, N202, N202, N167, N59);
nand NAND3 (N205, N204, N119, N27);
or OR2 (N206, N193, N186);
nor NOR3 (N207, N190, N127, N7);
and AND3 (N208, N207, N95, N105);
buf BUF1 (N209, N205);
nand NAND4 (N210, N206, N61, N34, N209);
nor NOR4 (N211, N36, N75, N86, N77);
and AND4 (N212, N172, N69, N6, N101);
and AND3 (N213, N208, N126, N111);
nor NOR2 (N214, N210, N98);
not NOT1 (N215, N195);
nand NAND4 (N216, N211, N214, N169, N192);
nor NOR2 (N217, N154, N3);
nor NOR4 (N218, N217, N34, N171, N162);
buf BUF1 (N219, N196);
nand NAND3 (N220, N200, N123, N38);
xor XOR2 (N221, N219, N74);
not NOT1 (N222, N213);
buf BUF1 (N223, N221);
xor XOR2 (N224, N212, N218);
nand NAND4 (N225, N45, N124, N80, N117);
nand NAND2 (N226, N222, N198);
not NOT1 (N227, N225);
nand NAND3 (N228, N227, N188, N130);
and AND4 (N229, N223, N135, N66, N174);
nor NOR3 (N230, N226, N181, N154);
and AND3 (N231, N187, N80, N5);
not NOT1 (N232, N180);
and AND4 (N233, N230, N42, N19, N89);
or OR4 (N234, N215, N141, N228, N93);
or OR3 (N235, N20, N55, N138);
not NOT1 (N236, N235);
not NOT1 (N237, N229);
xor XOR2 (N238, N236, N106);
or OR4 (N239, N224, N179, N118, N54);
buf BUF1 (N240, N216);
and AND4 (N241, N203, N205, N240, N160);
not NOT1 (N242, N7);
or OR4 (N243, N231, N70, N128, N112);
not NOT1 (N244, N243);
and AND4 (N245, N242, N91, N15, N90);
or OR2 (N246, N245, N214);
buf BUF1 (N247, N244);
xor XOR2 (N248, N239, N64);
nand NAND4 (N249, N246, N1, N75, N45);
xor XOR2 (N250, N232, N82);
not NOT1 (N251, N237);
nand NAND2 (N252, N248, N36);
nand NAND4 (N253, N249, N113, N128, N174);
or OR4 (N254, N234, N68, N8, N137);
buf BUF1 (N255, N238);
xor XOR2 (N256, N253, N221);
and AND3 (N257, N233, N77, N97);
and AND4 (N258, N220, N132, N162, N216);
and AND2 (N259, N254, N203);
nand NAND2 (N260, N257, N3);
xor XOR2 (N261, N258, N126);
or OR4 (N262, N260, N42, N175, N119);
and AND2 (N263, N247, N128);
xor XOR2 (N264, N250, N61);
buf BUF1 (N265, N263);
xor XOR2 (N266, N259, N15);
and AND3 (N267, N264, N123, N75);
buf BUF1 (N268, N261);
and AND2 (N269, N267, N225);
nor NOR4 (N270, N268, N234, N51, N116);
buf BUF1 (N271, N256);
buf BUF1 (N272, N270);
nand NAND2 (N273, N266, N135);
and AND3 (N274, N265, N143, N85);
buf BUF1 (N275, N252);
xor XOR2 (N276, N269, N69);
xor XOR2 (N277, N271, N37);
nand NAND2 (N278, N272, N170);
nor NOR2 (N279, N274, N166);
not NOT1 (N280, N273);
and AND2 (N281, N280, N242);
nor NOR2 (N282, N277, N279);
nor NOR2 (N283, N45, N92);
or OR3 (N284, N251, N108, N204);
nand NAND3 (N285, N276, N26, N262);
xor XOR2 (N286, N237, N170);
buf BUF1 (N287, N278);
xor XOR2 (N288, N275, N21);
xor XOR2 (N289, N282, N178);
and AND2 (N290, N285, N95);
and AND3 (N291, N255, N198, N276);
or OR3 (N292, N290, N205, N50);
not NOT1 (N293, N281);
and AND3 (N294, N293, N107, N102);
xor XOR2 (N295, N289, N17);
or OR3 (N296, N283, N86, N199);
and AND4 (N297, N287, N234, N138, N90);
buf BUF1 (N298, N295);
and AND3 (N299, N292, N294, N44);
buf BUF1 (N300, N151);
xor XOR2 (N301, N284, N262);
or OR4 (N302, N297, N243, N94, N233);
or OR3 (N303, N301, N163, N294);
xor XOR2 (N304, N291, N242);
not NOT1 (N305, N299);
nor NOR3 (N306, N303, N121, N278);
xor XOR2 (N307, N288, N284);
nand NAND3 (N308, N286, N131, N88);
not NOT1 (N309, N307);
or OR3 (N310, N302, N94, N155);
and AND4 (N311, N298, N5, N191, N69);
buf BUF1 (N312, N309);
or OR2 (N313, N311, N40);
and AND3 (N314, N312, N298, N152);
nand NAND4 (N315, N314, N184, N134, N296);
buf BUF1 (N316, N23);
not NOT1 (N317, N300);
not NOT1 (N318, N310);
nand NAND3 (N319, N241, N11, N151);
or OR3 (N320, N317, N185, N151);
not NOT1 (N321, N304);
buf BUF1 (N322, N315);
nor NOR2 (N323, N308, N138);
nor NOR2 (N324, N320, N266);
nor NOR4 (N325, N323, N316, N33, N116);
and AND2 (N326, N22, N110);
not NOT1 (N327, N321);
buf BUF1 (N328, N313);
nand NAND4 (N329, N318, N240, N145, N157);
or OR3 (N330, N305, N149, N194);
or OR3 (N331, N329, N145, N310);
nor NOR3 (N332, N306, N84, N231);
and AND2 (N333, N327, N80);
and AND4 (N334, N322, N24, N246, N225);
not NOT1 (N335, N331);
buf BUF1 (N336, N334);
nand NAND3 (N337, N333, N175, N253);
not NOT1 (N338, N324);
xor XOR2 (N339, N337, N1);
not NOT1 (N340, N335);
not NOT1 (N341, N340);
not NOT1 (N342, N338);
or OR4 (N343, N336, N305, N170, N294);
xor XOR2 (N344, N341, N334);
or OR2 (N345, N330, N112);
buf BUF1 (N346, N328);
buf BUF1 (N347, N326);
xor XOR2 (N348, N347, N298);
buf BUF1 (N349, N343);
nand NAND3 (N350, N319, N89, N161);
not NOT1 (N351, N345);
or OR4 (N352, N344, N328, N222, N348);
buf BUF1 (N353, N152);
buf BUF1 (N354, N325);
buf BUF1 (N355, N354);
xor XOR2 (N356, N349, N38);
not NOT1 (N357, N350);
xor XOR2 (N358, N353, N36);
xor XOR2 (N359, N351, N146);
not NOT1 (N360, N352);
nor NOR3 (N361, N357, N157, N260);
or OR3 (N362, N355, N218, N355);
xor XOR2 (N363, N332, N178);
nand NAND3 (N364, N342, N159, N99);
or OR4 (N365, N360, N99, N42, N316);
not NOT1 (N366, N339);
nand NAND3 (N367, N362, N259, N323);
buf BUF1 (N368, N363);
buf BUF1 (N369, N358);
or OR2 (N370, N368, N65);
or OR2 (N371, N359, N219);
xor XOR2 (N372, N366, N74);
xor XOR2 (N373, N361, N204);
or OR3 (N374, N372, N182, N26);
buf BUF1 (N375, N365);
buf BUF1 (N376, N367);
or OR2 (N377, N370, N315);
buf BUF1 (N378, N375);
nor NOR4 (N379, N373, N52, N109, N36);
xor XOR2 (N380, N369, N304);
or OR3 (N381, N379, N128, N130);
nor NOR4 (N382, N374, N139, N196, N43);
not NOT1 (N383, N371);
or OR4 (N384, N356, N97, N12, N95);
or OR4 (N385, N378, N157, N62, N206);
not NOT1 (N386, N381);
buf BUF1 (N387, N380);
nand NAND4 (N388, N376, N285, N211, N109);
and AND3 (N389, N386, N183, N42);
and AND2 (N390, N346, N320);
and AND3 (N391, N389, N212, N47);
nor NOR3 (N392, N390, N387, N388);
and AND3 (N393, N28, N264, N67);
nand NAND2 (N394, N97, N19);
buf BUF1 (N395, N382);
and AND2 (N396, N393, N267);
nand NAND2 (N397, N364, N57);
and AND4 (N398, N392, N34, N23, N162);
buf BUF1 (N399, N384);
nor NOR3 (N400, N391, N371, N227);
nor NOR4 (N401, N394, N271, N240, N352);
xor XOR2 (N402, N396, N373);
xor XOR2 (N403, N400, N150);
and AND2 (N404, N403, N77);
nand NAND2 (N405, N399, N334);
nor NOR2 (N406, N385, N79);
buf BUF1 (N407, N404);
buf BUF1 (N408, N407);
and AND3 (N409, N402, N201, N9);
nand NAND4 (N410, N409, N25, N98, N331);
not NOT1 (N411, N397);
nand NAND3 (N412, N383, N119, N321);
or OR3 (N413, N401, N231, N116);
buf BUF1 (N414, N395);
xor XOR2 (N415, N405, N253);
and AND3 (N416, N415, N175, N160);
xor XOR2 (N417, N413, N305);
buf BUF1 (N418, N406);
buf BUF1 (N419, N412);
buf BUF1 (N420, N410);
and AND2 (N421, N416, N297);
not NOT1 (N422, N414);
or OR3 (N423, N418, N277, N410);
xor XOR2 (N424, N408, N385);
buf BUF1 (N425, N422);
or OR2 (N426, N417, N102);
or OR2 (N427, N423, N2);
and AND2 (N428, N425, N309);
xor XOR2 (N429, N426, N111);
nand NAND4 (N430, N427, N189, N184, N122);
not NOT1 (N431, N420);
or OR2 (N432, N429, N345);
nor NOR2 (N433, N430, N416);
xor XOR2 (N434, N377, N351);
not NOT1 (N435, N398);
not NOT1 (N436, N419);
or OR2 (N437, N432, N256);
buf BUF1 (N438, N428);
nor NOR4 (N439, N424, N38, N66, N311);
or OR4 (N440, N439, N346, N358, N345);
nand NAND2 (N441, N431, N358);
xor XOR2 (N442, N437, N3);
xor XOR2 (N443, N421, N372);
buf BUF1 (N444, N443);
nand NAND3 (N445, N442, N290, N326);
nand NAND4 (N446, N435, N141, N387, N174);
not NOT1 (N447, N441);
nand NAND4 (N448, N446, N436, N367, N26);
buf BUF1 (N449, N256);
or OR4 (N450, N411, N411, N42, N284);
xor XOR2 (N451, N444, N219);
buf BUF1 (N452, N450);
xor XOR2 (N453, N452, N451);
or OR4 (N454, N422, N433, N99, N275);
and AND4 (N455, N383, N52, N350, N2);
nand NAND3 (N456, N448, N449, N413);
buf BUF1 (N457, N360);
or OR4 (N458, N440, N310, N312, N4);
and AND2 (N459, N454, N309);
and AND4 (N460, N459, N71, N50, N286);
xor XOR2 (N461, N434, N24);
or OR2 (N462, N438, N113);
buf BUF1 (N463, N445);
nor NOR4 (N464, N463, N174, N105, N355);
not NOT1 (N465, N457);
not NOT1 (N466, N447);
buf BUF1 (N467, N464);
and AND3 (N468, N458, N89, N354);
and AND2 (N469, N466, N255);
not NOT1 (N470, N467);
and AND4 (N471, N453, N205, N83, N307);
not NOT1 (N472, N456);
xor XOR2 (N473, N461, N461);
not NOT1 (N474, N455);
nor NOR2 (N475, N473, N108);
and AND2 (N476, N475, N352);
nand NAND3 (N477, N460, N392, N231);
not NOT1 (N478, N469);
nand NAND4 (N479, N476, N152, N180, N189);
and AND3 (N480, N479, N213, N13);
nor NOR2 (N481, N465, N113);
buf BUF1 (N482, N471);
not NOT1 (N483, N462);
or OR4 (N484, N474, N397, N324, N354);
not NOT1 (N485, N472);
not NOT1 (N486, N484);
nor NOR2 (N487, N470, N460);
nand NAND3 (N488, N478, N368, N296);
and AND3 (N489, N477, N267, N112);
xor XOR2 (N490, N485, N371);
and AND4 (N491, N486, N152, N201, N267);
xor XOR2 (N492, N480, N362);
xor XOR2 (N493, N468, N428);
nor NOR2 (N494, N493, N187);
xor XOR2 (N495, N492, N130);
xor XOR2 (N496, N495, N169);
not NOT1 (N497, N483);
and AND2 (N498, N489, N294);
not NOT1 (N499, N488);
nand NAND2 (N500, N482, N89);
nor NOR4 (N501, N499, N419, N216, N279);
and AND3 (N502, N500, N338, N86);
not NOT1 (N503, N490);
buf BUF1 (N504, N494);
xor XOR2 (N505, N504, N39);
or OR3 (N506, N481, N414, N420);
nor NOR4 (N507, N505, N399, N342, N105);
xor XOR2 (N508, N503, N244);
or OR4 (N509, N497, N130, N487, N22);
buf BUF1 (N510, N490);
not NOT1 (N511, N496);
not NOT1 (N512, N509);
not NOT1 (N513, N511);
and AND2 (N514, N506, N482);
not NOT1 (N515, N510);
or OR2 (N516, N512, N107);
xor XOR2 (N517, N507, N424);
xor XOR2 (N518, N515, N135);
not NOT1 (N519, N501);
nor NOR2 (N520, N517, N114);
and AND3 (N521, N508, N103, N168);
and AND2 (N522, N514, N400);
nor NOR3 (N523, N516, N475, N30);
and AND3 (N524, N521, N215, N93);
xor XOR2 (N525, N524, N300);
buf BUF1 (N526, N498);
or OR3 (N527, N526, N374, N300);
xor XOR2 (N528, N502, N468);
buf BUF1 (N529, N522);
buf BUF1 (N530, N527);
nand NAND4 (N531, N519, N124, N471, N202);
buf BUF1 (N532, N531);
and AND4 (N533, N513, N482, N23, N148);
not NOT1 (N534, N528);
not NOT1 (N535, N532);
or OR3 (N536, N520, N376, N214);
xor XOR2 (N537, N530, N45);
nand NAND2 (N538, N537, N389);
not NOT1 (N539, N534);
and AND3 (N540, N518, N386, N353);
nand NAND3 (N541, N523, N56, N45);
nand NAND4 (N542, N533, N48, N29, N360);
buf BUF1 (N543, N491);
or OR4 (N544, N539, N496, N97, N13);
and AND4 (N545, N536, N532, N282, N156);
or OR4 (N546, N541, N26, N368, N287);
or OR3 (N547, N542, N369, N464);
xor XOR2 (N548, N529, N94);
buf BUF1 (N549, N544);
nor NOR3 (N550, N543, N368, N477);
and AND3 (N551, N548, N501, N469);
xor XOR2 (N552, N546, N189);
nand NAND4 (N553, N552, N503, N143, N315);
nor NOR3 (N554, N550, N244, N287);
xor XOR2 (N555, N551, N537);
xor XOR2 (N556, N538, N102);
or OR3 (N557, N525, N11, N459);
nand NAND4 (N558, N555, N516, N385, N554);
and AND3 (N559, N274, N482, N448);
nand NAND2 (N560, N547, N277);
nand NAND4 (N561, N540, N88, N556, N322);
nor NOR4 (N562, N169, N462, N458, N553);
buf BUF1 (N563, N81);
or OR4 (N564, N557, N270, N94, N60);
buf BUF1 (N565, N545);
buf BUF1 (N566, N562);
not NOT1 (N567, N565);
nand NAND2 (N568, N564, N170);
not NOT1 (N569, N568);
not NOT1 (N570, N535);
nor NOR4 (N571, N561, N518, N468, N401);
not NOT1 (N572, N571);
or OR2 (N573, N558, N98);
and AND3 (N574, N560, N1, N182);
not NOT1 (N575, N570);
nand NAND2 (N576, N573, N109);
or OR3 (N577, N549, N148, N377);
nor NOR3 (N578, N559, N161, N200);
not NOT1 (N579, N567);
xor XOR2 (N580, N577, N315);
nand NAND2 (N581, N563, N77);
xor XOR2 (N582, N581, N158);
or OR3 (N583, N579, N271, N346);
or OR4 (N584, N578, N313, N153, N71);
nand NAND2 (N585, N572, N293);
not NOT1 (N586, N566);
buf BUF1 (N587, N576);
not NOT1 (N588, N574);
and AND4 (N589, N588, N283, N564, N53);
not NOT1 (N590, N584);
not NOT1 (N591, N582);
buf BUF1 (N592, N586);
xor XOR2 (N593, N587, N88);
and AND2 (N594, N591, N345);
xor XOR2 (N595, N593, N163);
xor XOR2 (N596, N589, N446);
not NOT1 (N597, N585);
and AND4 (N598, N590, N456, N91, N171);
not NOT1 (N599, N595);
or OR3 (N600, N597, N206, N115);
not NOT1 (N601, N592);
xor XOR2 (N602, N575, N309);
nor NOR4 (N603, N596, N160, N120, N241);
nor NOR4 (N604, N603, N463, N593, N345);
not NOT1 (N605, N599);
xor XOR2 (N606, N601, N108);
or OR4 (N607, N605, N412, N49, N150);
xor XOR2 (N608, N604, N346);
and AND4 (N609, N598, N504, N211, N608);
or OR4 (N610, N422, N600, N588, N288);
nor NOR3 (N611, N428, N81, N478);
xor XOR2 (N612, N610, N436);
nand NAND2 (N613, N602, N355);
xor XOR2 (N614, N594, N384);
nor NOR3 (N615, N612, N248, N332);
and AND3 (N616, N580, N452, N525);
or OR2 (N617, N616, N445);
buf BUF1 (N618, N583);
nand NAND2 (N619, N569, N459);
and AND2 (N620, N617, N429);
and AND2 (N621, N606, N186);
xor XOR2 (N622, N615, N242);
endmodule