// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N6406,N6416,N6418,N6421,N6414,N6408,N6402,N6419,N6420,N6422;

xor XOR2 (N23, N7, N3);
buf BUF1 (N24, N12);
buf BUF1 (N25, N7);
not NOT1 (N26, N25);
nor NOR3 (N27, N19, N15, N4);
not NOT1 (N28, N5);
nand NAND4 (N29, N13, N25, N10, N27);
not NOT1 (N30, N12);
not NOT1 (N31, N6);
and AND3 (N32, N11, N20, N17);
and AND2 (N33, N12, N5);
and AND3 (N34, N20, N1, N29);
not NOT1 (N35, N19);
nor NOR3 (N36, N32, N11, N14);
and AND4 (N37, N35, N19, N11, N26);
not NOT1 (N38, N13);
nand NAND4 (N39, N24, N2, N25, N37);
nor NOR3 (N40, N18, N32, N1);
or OR4 (N41, N39, N38, N18, N17);
nor NOR4 (N42, N14, N12, N8, N21);
not NOT1 (N43, N40);
nor NOR4 (N44, N33, N11, N36, N22);
and AND3 (N45, N25, N14, N2);
nor NOR4 (N46, N42, N3, N4, N14);
or OR3 (N47, N31, N42, N31);
or OR4 (N48, N23, N33, N10, N28);
not NOT1 (N49, N14);
nor NOR3 (N50, N45, N30, N15);
not NOT1 (N51, N39);
nor NOR3 (N52, N43, N26, N21);
and AND3 (N53, N50, N36, N36);
and AND3 (N54, N53, N2, N53);
nand NAND2 (N55, N54, N32);
nor NOR3 (N56, N55, N2, N40);
or OR4 (N57, N47, N19, N2, N32);
not NOT1 (N58, N44);
nor NOR4 (N59, N56, N32, N34, N20);
xor XOR2 (N60, N37, N22);
nor NOR2 (N61, N46, N32);
not NOT1 (N62, N60);
nand NAND4 (N63, N41, N33, N42, N46);
and AND2 (N64, N48, N58);
or OR3 (N65, N19, N6, N11);
and AND4 (N66, N52, N41, N61, N36);
buf BUF1 (N67, N29);
buf BUF1 (N68, N49);
buf BUF1 (N69, N62);
nand NAND4 (N70, N67, N47, N5, N63);
nor NOR3 (N71, N44, N69, N21);
or OR2 (N72, N40, N59);
not NOT1 (N73, N33);
nand NAND3 (N74, N51, N60, N43);
nand NAND2 (N75, N65, N15);
and AND2 (N76, N71, N13);
xor XOR2 (N77, N57, N47);
or OR3 (N78, N64, N69, N77);
buf BUF1 (N79, N25);
buf BUF1 (N80, N74);
and AND4 (N81, N66, N53, N66, N24);
not NOT1 (N82, N73);
not NOT1 (N83, N79);
nand NAND2 (N84, N75, N39);
nor NOR2 (N85, N80, N21);
buf BUF1 (N86, N76);
nor NOR2 (N87, N82, N85);
or OR4 (N88, N15, N58, N38, N12);
nor NOR3 (N89, N70, N50, N20);
buf BUF1 (N90, N78);
nand NAND4 (N91, N72, N44, N85, N72);
nor NOR4 (N92, N88, N80, N74, N76);
xor XOR2 (N93, N84, N23);
xor XOR2 (N94, N91, N78);
nand NAND4 (N95, N87, N6, N54, N40);
buf BUF1 (N96, N93);
nor NOR2 (N97, N81, N58);
not NOT1 (N98, N95);
buf BUF1 (N99, N90);
nor NOR4 (N100, N96, N62, N66, N99);
xor XOR2 (N101, N32, N88);
xor XOR2 (N102, N92, N51);
xor XOR2 (N103, N68, N68);
or OR4 (N104, N94, N85, N87, N62);
or OR2 (N105, N103, N84);
buf BUF1 (N106, N89);
or OR4 (N107, N97, N20, N31, N100);
nor NOR3 (N108, N35, N56, N6);
not NOT1 (N109, N104);
xor XOR2 (N110, N86, N60);
not NOT1 (N111, N109);
buf BUF1 (N112, N106);
and AND3 (N113, N83, N55, N36);
nor NOR2 (N114, N102, N97);
nor NOR2 (N115, N107, N78);
and AND2 (N116, N112, N77);
not NOT1 (N117, N101);
buf BUF1 (N118, N113);
and AND3 (N119, N118, N12, N31);
nand NAND2 (N120, N119, N19);
or OR2 (N121, N116, N116);
not NOT1 (N122, N115);
and AND2 (N123, N117, N100);
nand NAND4 (N124, N114, N26, N86, N56);
or OR2 (N125, N122, N42);
buf BUF1 (N126, N108);
nor NOR4 (N127, N105, N115, N73, N77);
nor NOR4 (N128, N110, N126, N106, N8);
and AND3 (N129, N63, N112, N92);
nor NOR4 (N130, N123, N62, N9, N15);
and AND2 (N131, N124, N21);
or OR4 (N132, N111, N29, N81, N59);
xor XOR2 (N133, N120, N91);
nor NOR2 (N134, N98, N12);
or OR4 (N135, N129, N120, N24, N32);
or OR2 (N136, N134, N116);
xor XOR2 (N137, N131, N91);
xor XOR2 (N138, N136, N126);
and AND4 (N139, N127, N88, N112, N58);
or OR4 (N140, N133, N114, N30, N108);
not NOT1 (N141, N130);
or OR2 (N142, N141, N74);
xor XOR2 (N143, N125, N87);
or OR4 (N144, N140, N99, N57, N70);
nor NOR3 (N145, N121, N46, N111);
and AND4 (N146, N128, N5, N11, N50);
nor NOR3 (N147, N145, N115, N28);
buf BUF1 (N148, N132);
or OR4 (N149, N138, N46, N66, N62);
nand NAND2 (N150, N144, N40);
buf BUF1 (N151, N149);
buf BUF1 (N152, N151);
nor NOR3 (N153, N143, N9, N145);
buf BUF1 (N154, N139);
nand NAND3 (N155, N137, N91, N140);
not NOT1 (N156, N148);
not NOT1 (N157, N142);
buf BUF1 (N158, N156);
or OR3 (N159, N135, N32, N137);
xor XOR2 (N160, N152, N45);
xor XOR2 (N161, N158, N58);
buf BUF1 (N162, N146);
or OR2 (N163, N161, N36);
and AND4 (N164, N153, N72, N158, N29);
nand NAND3 (N165, N160, N48, N70);
buf BUF1 (N166, N162);
buf BUF1 (N167, N166);
and AND2 (N168, N165, N159);
and AND4 (N169, N28, N146, N113, N162);
xor XOR2 (N170, N155, N149);
xor XOR2 (N171, N154, N53);
xor XOR2 (N172, N171, N92);
or OR4 (N173, N167, N119, N29, N64);
not NOT1 (N174, N172);
nor NOR4 (N175, N173, N45, N71, N105);
xor XOR2 (N176, N168, N107);
and AND2 (N177, N164, N152);
nand NAND2 (N178, N147, N171);
buf BUF1 (N179, N175);
nand NAND3 (N180, N176, N77, N66);
nand NAND3 (N181, N150, N60, N32);
xor XOR2 (N182, N170, N88);
nor NOR3 (N183, N174, N48, N153);
xor XOR2 (N184, N181, N154);
nor NOR3 (N185, N184, N54, N95);
buf BUF1 (N186, N182);
nor NOR2 (N187, N180, N71);
nor NOR4 (N188, N157, N13, N51, N140);
xor XOR2 (N189, N187, N160);
nand NAND2 (N190, N183, N28);
not NOT1 (N191, N189);
xor XOR2 (N192, N177, N174);
nor NOR4 (N193, N188, N86, N45, N186);
xor XOR2 (N194, N172, N97);
nor NOR3 (N195, N190, N4, N70);
xor XOR2 (N196, N179, N70);
xor XOR2 (N197, N194, N155);
xor XOR2 (N198, N197, N1);
not NOT1 (N199, N198);
or OR3 (N200, N192, N134, N163);
or OR4 (N201, N130, N134, N93, N115);
or OR3 (N202, N196, N158, N127);
or OR3 (N203, N178, N67, N194);
nor NOR2 (N204, N199, N30);
not NOT1 (N205, N200);
buf BUF1 (N206, N202);
nand NAND2 (N207, N205, N133);
xor XOR2 (N208, N207, N66);
not NOT1 (N209, N206);
not NOT1 (N210, N201);
buf BUF1 (N211, N191);
buf BUF1 (N212, N185);
or OR2 (N213, N193, N75);
nor NOR2 (N214, N210, N208);
nor NOR2 (N215, N147, N212);
buf BUF1 (N216, N212);
xor XOR2 (N217, N216, N111);
and AND3 (N218, N203, N24, N50);
or OR2 (N219, N217, N25);
and AND2 (N220, N218, N130);
nand NAND3 (N221, N213, N53, N125);
buf BUF1 (N222, N221);
or OR4 (N223, N195, N143, N161, N139);
and AND3 (N224, N223, N214, N24);
and AND4 (N225, N173, N18, N18, N5);
buf BUF1 (N226, N219);
xor XOR2 (N227, N211, N189);
nor NOR2 (N228, N224, N82);
nand NAND2 (N229, N204, N26);
xor XOR2 (N230, N229, N179);
nor NOR4 (N231, N209, N84, N78, N14);
and AND4 (N232, N220, N19, N171, N38);
not NOT1 (N233, N215);
nand NAND3 (N234, N228, N59, N35);
not NOT1 (N235, N231);
or OR4 (N236, N230, N227, N7, N72);
and AND4 (N237, N177, N55, N175, N166);
nand NAND4 (N238, N236, N224, N121, N219);
xor XOR2 (N239, N222, N181);
and AND2 (N240, N169, N202);
or OR3 (N241, N233, N121, N63);
nor NOR2 (N242, N241, N125);
not NOT1 (N243, N239);
nor NOR3 (N244, N240, N167, N202);
and AND3 (N245, N242, N193, N178);
buf BUF1 (N246, N232);
buf BUF1 (N247, N238);
nor NOR3 (N248, N247, N207, N221);
xor XOR2 (N249, N248, N67);
nand NAND4 (N250, N234, N48, N179, N16);
or OR2 (N251, N246, N55);
nor NOR2 (N252, N226, N141);
and AND3 (N253, N244, N137, N198);
nor NOR2 (N254, N253, N137);
buf BUF1 (N255, N225);
or OR4 (N256, N251, N78, N61, N173);
nand NAND4 (N257, N256, N149, N126, N174);
nor NOR2 (N258, N243, N110);
nor NOR2 (N259, N245, N156);
not NOT1 (N260, N257);
nor NOR3 (N261, N249, N133, N28);
nor NOR3 (N262, N258, N105, N47);
not NOT1 (N263, N260);
buf BUF1 (N264, N252);
buf BUF1 (N265, N254);
xor XOR2 (N266, N261, N144);
or OR4 (N267, N235, N92, N7, N136);
and AND2 (N268, N250, N116);
and AND4 (N269, N259, N265, N191, N74);
xor XOR2 (N270, N264, N221);
nand NAND3 (N271, N162, N82, N67);
nand NAND2 (N272, N267, N122);
xor XOR2 (N273, N263, N71);
nand NAND2 (N274, N270, N152);
xor XOR2 (N275, N255, N231);
or OR3 (N276, N272, N162, N145);
not NOT1 (N277, N266);
or OR2 (N278, N277, N194);
nor NOR2 (N279, N237, N49);
not NOT1 (N280, N269);
not NOT1 (N281, N274);
nor NOR2 (N282, N271, N72);
and AND3 (N283, N278, N100, N101);
nand NAND4 (N284, N280, N181, N82, N48);
or OR2 (N285, N273, N235);
nor NOR2 (N286, N283, N254);
xor XOR2 (N287, N281, N76);
nand NAND4 (N288, N285, N273, N119, N235);
nor NOR2 (N289, N287, N283);
not NOT1 (N290, N289);
not NOT1 (N291, N275);
nand NAND2 (N292, N262, N276);
and AND2 (N293, N263, N102);
and AND3 (N294, N286, N175, N277);
nor NOR2 (N295, N284, N234);
xor XOR2 (N296, N288, N23);
buf BUF1 (N297, N268);
not NOT1 (N298, N296);
nor NOR2 (N299, N295, N248);
or OR3 (N300, N297, N193, N150);
nor NOR4 (N301, N292, N249, N109, N3);
and AND3 (N302, N293, N146, N102);
and AND3 (N303, N298, N111, N181);
nand NAND2 (N304, N300, N30);
not NOT1 (N305, N290);
or OR4 (N306, N279, N149, N246, N245);
nor NOR2 (N307, N304, N243);
nand NAND3 (N308, N301, N225, N33);
nand NAND4 (N309, N305, N60, N136, N105);
or OR3 (N310, N299, N137, N131);
buf BUF1 (N311, N294);
and AND3 (N312, N310, N122, N14);
or OR4 (N313, N309, N307, N236, N287);
nor NOR3 (N314, N108, N177, N115);
buf BUF1 (N315, N311);
nand NAND3 (N316, N302, N226, N199);
not NOT1 (N317, N291);
buf BUF1 (N318, N312);
nor NOR4 (N319, N306, N161, N305, N72);
nor NOR2 (N320, N315, N261);
xor XOR2 (N321, N314, N286);
xor XOR2 (N322, N313, N317);
xor XOR2 (N323, N255, N80);
nand NAND3 (N324, N320, N187, N118);
and AND4 (N325, N324, N14, N71, N213);
nor NOR3 (N326, N325, N185, N282);
nand NAND4 (N327, N94, N42, N77, N10);
buf BUF1 (N328, N308);
buf BUF1 (N329, N328);
nor NOR2 (N330, N321, N305);
xor XOR2 (N331, N319, N195);
buf BUF1 (N332, N330);
buf BUF1 (N333, N327);
not NOT1 (N334, N329);
not NOT1 (N335, N316);
and AND2 (N336, N323, N33);
xor XOR2 (N337, N322, N141);
nor NOR3 (N338, N318, N231, N105);
xor XOR2 (N339, N326, N87);
nand NAND4 (N340, N336, N139, N238, N186);
not NOT1 (N341, N303);
nor NOR4 (N342, N340, N177, N120, N148);
xor XOR2 (N343, N332, N260);
not NOT1 (N344, N343);
nor NOR4 (N345, N334, N267, N8, N227);
xor XOR2 (N346, N331, N304);
not NOT1 (N347, N341);
xor XOR2 (N348, N345, N210);
nand NAND4 (N349, N338, N140, N50, N12);
nand NAND4 (N350, N333, N92, N66, N112);
and AND3 (N351, N344, N334, N83);
and AND2 (N352, N342, N290);
not NOT1 (N353, N350);
xor XOR2 (N354, N339, N128);
nand NAND2 (N355, N352, N322);
xor XOR2 (N356, N353, N75);
buf BUF1 (N357, N335);
and AND3 (N358, N349, N356, N343);
buf BUF1 (N359, N8);
xor XOR2 (N360, N337, N129);
and AND4 (N361, N348, N294, N186, N91);
nand NAND2 (N362, N351, N223);
nand NAND3 (N363, N357, N166, N321);
buf BUF1 (N364, N354);
and AND2 (N365, N360, N3);
buf BUF1 (N366, N361);
not NOT1 (N367, N346);
xor XOR2 (N368, N347, N245);
nor NOR4 (N369, N362, N11, N278, N16);
buf BUF1 (N370, N367);
nor NOR4 (N371, N369, N332, N342, N268);
buf BUF1 (N372, N359);
and AND4 (N373, N371, N279, N64, N262);
nor NOR3 (N374, N365, N366, N256);
xor XOR2 (N375, N243, N312);
nor NOR2 (N376, N368, N329);
nor NOR3 (N377, N374, N173, N251);
and AND3 (N378, N377, N261, N332);
nor NOR2 (N379, N358, N277);
xor XOR2 (N380, N363, N205);
and AND2 (N381, N378, N219);
buf BUF1 (N382, N372);
nor NOR2 (N383, N373, N312);
nor NOR4 (N384, N375, N51, N13, N328);
and AND2 (N385, N355, N125);
and AND4 (N386, N364, N104, N26, N378);
or OR3 (N387, N381, N275, N63);
nand NAND4 (N388, N387, N139, N173, N278);
or OR3 (N389, N385, N279, N276);
not NOT1 (N390, N389);
nor NOR4 (N391, N380, N46, N171, N304);
nand NAND4 (N392, N379, N23, N145, N165);
or OR4 (N393, N376, N163, N376, N44);
nand NAND2 (N394, N386, N199);
or OR2 (N395, N383, N112);
xor XOR2 (N396, N393, N163);
xor XOR2 (N397, N394, N363);
nand NAND2 (N398, N396, N88);
nand NAND4 (N399, N384, N372, N143, N72);
buf BUF1 (N400, N391);
or OR3 (N401, N370, N40, N199);
nand NAND2 (N402, N395, N173);
and AND3 (N403, N401, N58, N260);
nand NAND2 (N404, N403, N19);
not NOT1 (N405, N390);
and AND3 (N406, N388, N336, N173);
nor NOR4 (N407, N399, N279, N288, N102);
nand NAND4 (N408, N392, N1, N225, N389);
and AND3 (N409, N408, N82, N103);
nand NAND4 (N410, N400, N290, N256, N219);
nand NAND2 (N411, N407, N369);
nand NAND4 (N412, N402, N228, N313, N126);
xor XOR2 (N413, N404, N204);
xor XOR2 (N414, N398, N325);
xor XOR2 (N415, N406, N28);
xor XOR2 (N416, N382, N372);
not NOT1 (N417, N413);
nor NOR4 (N418, N416, N238, N57, N163);
buf BUF1 (N419, N411);
or OR4 (N420, N412, N216, N20, N356);
and AND2 (N421, N418, N22);
or OR4 (N422, N421, N24, N36, N356);
buf BUF1 (N423, N410);
and AND2 (N424, N414, N124);
or OR3 (N425, N419, N335, N132);
nand NAND3 (N426, N409, N229, N39);
and AND3 (N427, N422, N86, N409);
not NOT1 (N428, N420);
and AND4 (N429, N426, N106, N299, N202);
not NOT1 (N430, N428);
xor XOR2 (N431, N429, N30);
and AND3 (N432, N415, N310, N320);
and AND4 (N433, N423, N126, N379, N217);
nand NAND3 (N434, N405, N374, N321);
xor XOR2 (N435, N417, N232);
xor XOR2 (N436, N424, N228);
nor NOR3 (N437, N436, N24, N186);
nor NOR4 (N438, N427, N203, N390, N198);
not NOT1 (N439, N397);
buf BUF1 (N440, N439);
nand NAND2 (N441, N435, N324);
and AND4 (N442, N434, N243, N121, N68);
not NOT1 (N443, N437);
xor XOR2 (N444, N442, N403);
nor NOR4 (N445, N430, N27, N29, N295);
not NOT1 (N446, N441);
and AND4 (N447, N433, N182, N81, N142);
not NOT1 (N448, N443);
or OR2 (N449, N445, N75);
xor XOR2 (N450, N432, N147);
nand NAND4 (N451, N425, N113, N423, N217);
and AND3 (N452, N438, N235, N85);
and AND4 (N453, N444, N51, N105, N33);
or OR2 (N454, N440, N221);
nand NAND3 (N455, N446, N241, N73);
not NOT1 (N456, N448);
and AND4 (N457, N455, N51, N121, N376);
or OR4 (N458, N457, N143, N392, N357);
and AND3 (N459, N450, N353, N273);
nand NAND3 (N460, N453, N396, N213);
nand NAND3 (N461, N454, N448, N226);
not NOT1 (N462, N451);
and AND4 (N463, N449, N29, N326, N8);
or OR4 (N464, N459, N172, N456, N24);
or OR2 (N465, N35, N443);
or OR2 (N466, N462, N71);
nand NAND3 (N467, N463, N97, N278);
xor XOR2 (N468, N460, N70);
not NOT1 (N469, N465);
nor NOR4 (N470, N431, N148, N390, N245);
xor XOR2 (N471, N461, N4);
nand NAND4 (N472, N471, N278, N135, N22);
or OR2 (N473, N452, N19);
and AND4 (N474, N467, N347, N454, N87);
nor NOR3 (N475, N472, N99, N466);
and AND3 (N476, N267, N341, N321);
nand NAND4 (N477, N475, N3, N65, N260);
nor NOR4 (N478, N477, N31, N136, N437);
xor XOR2 (N479, N478, N146);
buf BUF1 (N480, N468);
or OR4 (N481, N474, N48, N153, N102);
buf BUF1 (N482, N479);
xor XOR2 (N483, N447, N67);
and AND2 (N484, N469, N317);
or OR3 (N485, N482, N425, N212);
and AND3 (N486, N480, N237, N260);
or OR3 (N487, N486, N388, N400);
buf BUF1 (N488, N473);
not NOT1 (N489, N481);
not NOT1 (N490, N476);
buf BUF1 (N491, N489);
xor XOR2 (N492, N491, N180);
xor XOR2 (N493, N464, N80);
or OR3 (N494, N487, N472, N323);
not NOT1 (N495, N492);
not NOT1 (N496, N483);
nand NAND3 (N497, N494, N127, N129);
and AND2 (N498, N490, N4);
and AND2 (N499, N495, N219);
xor XOR2 (N500, N493, N93);
xor XOR2 (N501, N470, N398);
and AND2 (N502, N496, N492);
and AND2 (N503, N498, N109);
buf BUF1 (N504, N501);
nor NOR4 (N505, N484, N290, N385, N172);
nand NAND3 (N506, N488, N187, N396);
nand NAND3 (N507, N506, N436, N387);
xor XOR2 (N508, N502, N2);
xor XOR2 (N509, N504, N203);
not NOT1 (N510, N509);
and AND4 (N511, N458, N151, N45, N332);
buf BUF1 (N512, N507);
xor XOR2 (N513, N511, N37);
nand NAND4 (N514, N503, N500, N208, N45);
buf BUF1 (N515, N279);
and AND4 (N516, N499, N456, N210, N228);
xor XOR2 (N517, N516, N429);
xor XOR2 (N518, N514, N26);
buf BUF1 (N519, N518);
and AND2 (N520, N497, N314);
buf BUF1 (N521, N519);
not NOT1 (N522, N513);
nand NAND4 (N523, N520, N279, N195, N176);
or OR3 (N524, N522, N162, N372);
xor XOR2 (N525, N523, N211);
and AND2 (N526, N512, N68);
or OR2 (N527, N521, N335);
xor XOR2 (N528, N485, N296);
not NOT1 (N529, N525);
buf BUF1 (N530, N510);
xor XOR2 (N531, N505, N519);
or OR2 (N532, N530, N269);
not NOT1 (N533, N527);
buf BUF1 (N534, N524);
and AND4 (N535, N531, N102, N283, N308);
xor XOR2 (N536, N534, N406);
xor XOR2 (N537, N533, N528);
nand NAND2 (N538, N147, N101);
nor NOR4 (N539, N535, N289, N189, N413);
not NOT1 (N540, N529);
buf BUF1 (N541, N532);
not NOT1 (N542, N536);
xor XOR2 (N543, N541, N40);
or OR3 (N544, N538, N531, N457);
nor NOR2 (N545, N517, N33);
or OR4 (N546, N540, N11, N167, N424);
buf BUF1 (N547, N543);
nor NOR4 (N548, N508, N265, N520, N178);
and AND4 (N549, N546, N346, N79, N56);
and AND4 (N550, N539, N528, N537, N157);
nand NAND4 (N551, N166, N119, N190, N292);
or OR2 (N552, N548, N388);
and AND3 (N553, N544, N537, N22);
nand NAND4 (N554, N547, N369, N322, N184);
or OR3 (N555, N551, N206, N443);
not NOT1 (N556, N553);
and AND3 (N557, N526, N230, N204);
nand NAND4 (N558, N554, N378, N544, N348);
buf BUF1 (N559, N542);
xor XOR2 (N560, N549, N200);
buf BUF1 (N561, N558);
nand NAND4 (N562, N556, N59, N548, N411);
nand NAND2 (N563, N560, N388);
and AND2 (N564, N563, N553);
not NOT1 (N565, N515);
nand NAND4 (N566, N555, N55, N429, N172);
and AND2 (N567, N552, N452);
nor NOR3 (N568, N562, N452, N213);
xor XOR2 (N569, N566, N217);
nand NAND4 (N570, N545, N345, N401, N100);
nand NAND3 (N571, N550, N562, N135);
and AND3 (N572, N571, N96, N116);
or OR2 (N573, N567, N525);
and AND2 (N574, N561, N193);
xor XOR2 (N575, N570, N366);
nand NAND2 (N576, N572, N2);
and AND2 (N577, N564, N312);
buf BUF1 (N578, N575);
buf BUF1 (N579, N559);
or OR2 (N580, N565, N139);
or OR3 (N581, N577, N74, N373);
xor XOR2 (N582, N579, N33);
nand NAND4 (N583, N568, N93, N462, N426);
nand NAND3 (N584, N576, N249, N220);
and AND4 (N585, N557, N570, N239, N453);
nand NAND2 (N586, N573, N249);
or OR4 (N587, N581, N508, N226, N465);
nand NAND2 (N588, N578, N306);
nand NAND3 (N589, N580, N499, N281);
buf BUF1 (N590, N587);
and AND2 (N591, N582, N257);
or OR3 (N592, N589, N393, N483);
buf BUF1 (N593, N590);
and AND4 (N594, N592, N379, N44, N483);
buf BUF1 (N595, N584);
and AND3 (N596, N588, N234, N434);
not NOT1 (N597, N583);
and AND3 (N598, N595, N244, N443);
not NOT1 (N599, N574);
nand NAND3 (N600, N597, N215, N497);
xor XOR2 (N601, N569, N28);
nor NOR4 (N602, N591, N86, N181, N529);
nor NOR4 (N603, N594, N508, N573, N306);
not NOT1 (N604, N598);
xor XOR2 (N605, N604, N533);
not NOT1 (N606, N596);
nand NAND2 (N607, N593, N116);
not NOT1 (N608, N586);
xor XOR2 (N609, N605, N253);
and AND3 (N610, N599, N525, N122);
not NOT1 (N611, N601);
nor NOR3 (N612, N585, N554, N178);
buf BUF1 (N613, N606);
xor XOR2 (N614, N613, N222);
not NOT1 (N615, N608);
not NOT1 (N616, N615);
nand NAND3 (N617, N600, N79, N296);
not NOT1 (N618, N602);
nor NOR4 (N619, N607, N265, N289, N603);
xor XOR2 (N620, N580, N251);
and AND2 (N621, N614, N607);
and AND2 (N622, N620, N537);
and AND3 (N623, N618, N408, N268);
and AND2 (N624, N611, N268);
and AND2 (N625, N624, N433);
and AND3 (N626, N610, N477, N130);
nand NAND2 (N627, N616, N389);
buf BUF1 (N628, N612);
nor NOR2 (N629, N617, N217);
not NOT1 (N630, N628);
or OR3 (N631, N609, N495, N595);
nor NOR4 (N632, N621, N244, N412, N139);
and AND2 (N633, N627, N583);
or OR4 (N634, N622, N322, N443, N614);
nand NAND2 (N635, N630, N129);
nor NOR3 (N636, N629, N495, N492);
xor XOR2 (N637, N631, N161);
or OR2 (N638, N633, N35);
nor NOR3 (N639, N634, N336, N440);
not NOT1 (N640, N638);
nand NAND3 (N641, N637, N482, N248);
nor NOR2 (N642, N635, N113);
nand NAND4 (N643, N632, N604, N614, N588);
or OR3 (N644, N623, N368, N26);
xor XOR2 (N645, N626, N288);
nand NAND3 (N646, N625, N393, N334);
nor NOR4 (N647, N639, N185, N218, N220);
and AND4 (N648, N644, N619, N540, N201);
buf BUF1 (N649, N239);
not NOT1 (N650, N640);
nor NOR2 (N651, N643, N591);
nand NAND2 (N652, N649, N201);
or OR3 (N653, N641, N257, N564);
nand NAND3 (N654, N651, N363, N441);
nand NAND3 (N655, N647, N607, N336);
and AND4 (N656, N636, N214, N113, N271);
or OR2 (N657, N653, N508);
xor XOR2 (N658, N648, N51);
and AND3 (N659, N646, N519, N286);
xor XOR2 (N660, N652, N256);
nor NOR2 (N661, N645, N514);
xor XOR2 (N662, N660, N539);
not NOT1 (N663, N662);
and AND3 (N664, N642, N409, N286);
xor XOR2 (N665, N664, N376);
nor NOR2 (N666, N665, N186);
or OR3 (N667, N654, N394, N98);
not NOT1 (N668, N663);
nor NOR2 (N669, N668, N189);
nor NOR4 (N670, N657, N303, N138, N281);
and AND4 (N671, N655, N101, N377, N383);
and AND4 (N672, N671, N162, N605, N44);
nand NAND4 (N673, N658, N154, N123, N560);
buf BUF1 (N674, N650);
nor NOR2 (N675, N666, N653);
not NOT1 (N676, N673);
and AND3 (N677, N669, N173, N117);
or OR4 (N678, N661, N207, N452, N377);
nand NAND2 (N679, N670, N341);
nor NOR2 (N680, N672, N678);
nor NOR2 (N681, N72, N550);
and AND3 (N682, N679, N49, N106);
xor XOR2 (N683, N675, N251);
or OR2 (N684, N682, N229);
xor XOR2 (N685, N683, N112);
nand NAND3 (N686, N676, N430, N400);
buf BUF1 (N687, N686);
xor XOR2 (N688, N667, N71);
nor NOR4 (N689, N674, N646, N623, N91);
not NOT1 (N690, N656);
or OR4 (N691, N685, N633, N123, N468);
or OR2 (N692, N687, N336);
buf BUF1 (N693, N681);
nor NOR3 (N694, N677, N129, N291);
buf BUF1 (N695, N691);
xor XOR2 (N696, N688, N330);
or OR3 (N697, N659, N263, N624);
and AND3 (N698, N693, N593, N422);
buf BUF1 (N699, N692);
nor NOR4 (N700, N699, N216, N579, N397);
not NOT1 (N701, N694);
nor NOR3 (N702, N684, N652, N664);
or OR4 (N703, N695, N368, N267, N388);
nor NOR4 (N704, N690, N89, N697, N245);
nand NAND2 (N705, N322, N469);
not NOT1 (N706, N700);
nor NOR2 (N707, N702, N220);
nand NAND4 (N708, N703, N576, N379, N546);
not NOT1 (N709, N705);
or OR4 (N710, N708, N73, N348, N34);
nor NOR3 (N711, N704, N85, N352);
xor XOR2 (N712, N707, N293);
nor NOR2 (N713, N712, N33);
or OR4 (N714, N680, N445, N181, N300);
nand NAND4 (N715, N706, N300, N671, N143);
xor XOR2 (N716, N701, N304);
or OR2 (N717, N696, N670);
or OR2 (N718, N698, N308);
or OR3 (N719, N689, N372, N705);
buf BUF1 (N720, N710);
nand NAND3 (N721, N716, N192, N274);
or OR4 (N722, N709, N407, N60, N120);
buf BUF1 (N723, N713);
xor XOR2 (N724, N723, N237);
buf BUF1 (N725, N718);
not NOT1 (N726, N724);
nand NAND3 (N727, N726, N635, N436);
nor NOR4 (N728, N715, N74, N519, N523);
and AND3 (N729, N714, N682, N267);
xor XOR2 (N730, N722, N231);
buf BUF1 (N731, N717);
nand NAND4 (N732, N730, N491, N584, N551);
xor XOR2 (N733, N711, N100);
and AND3 (N734, N727, N317, N510);
nand NAND3 (N735, N719, N189, N61);
xor XOR2 (N736, N735, N89);
nor NOR2 (N737, N720, N658);
buf BUF1 (N738, N729);
nor NOR4 (N739, N737, N90, N219, N318);
not NOT1 (N740, N732);
not NOT1 (N741, N740);
nor NOR3 (N742, N738, N616, N161);
buf BUF1 (N743, N728);
xor XOR2 (N744, N741, N57);
nor NOR4 (N745, N739, N138, N697, N326);
or OR3 (N746, N742, N298, N214);
nor NOR2 (N747, N746, N164);
or OR4 (N748, N721, N612, N77, N636);
or OR2 (N749, N733, N89);
nand NAND2 (N750, N744, N553);
xor XOR2 (N751, N748, N80);
not NOT1 (N752, N750);
not NOT1 (N753, N752);
and AND2 (N754, N725, N697);
buf BUF1 (N755, N731);
buf BUF1 (N756, N755);
nor NOR4 (N757, N745, N184, N469, N554);
not NOT1 (N758, N754);
nand NAND2 (N759, N734, N301);
nand NAND3 (N760, N749, N32, N280);
or OR4 (N761, N753, N599, N24, N720);
nor NOR4 (N762, N736, N640, N88, N504);
nand NAND4 (N763, N747, N12, N615, N52);
not NOT1 (N764, N751);
nor NOR2 (N765, N757, N423);
nand NAND3 (N766, N743, N46, N191);
or OR2 (N767, N762, N636);
xor XOR2 (N768, N756, N589);
and AND4 (N769, N760, N497, N417, N116);
not NOT1 (N770, N761);
buf BUF1 (N771, N767);
buf BUF1 (N772, N771);
not NOT1 (N773, N766);
xor XOR2 (N774, N769, N451);
or OR3 (N775, N774, N752, N628);
not NOT1 (N776, N770);
or OR4 (N777, N758, N771, N588, N615);
and AND3 (N778, N764, N464, N11);
nand NAND4 (N779, N763, N115, N13, N702);
and AND3 (N780, N776, N72, N730);
or OR3 (N781, N779, N358, N414);
not NOT1 (N782, N775);
and AND3 (N783, N782, N429, N586);
or OR4 (N784, N759, N720, N734, N127);
or OR2 (N785, N784, N770);
not NOT1 (N786, N783);
and AND2 (N787, N768, N370);
nand NAND4 (N788, N781, N189, N241, N113);
and AND3 (N789, N785, N773, N283);
nor NOR2 (N790, N135, N515);
buf BUF1 (N791, N765);
nor NOR4 (N792, N788, N760, N551, N3);
nor NOR4 (N793, N792, N723, N730, N673);
buf BUF1 (N794, N791);
and AND3 (N795, N786, N249, N691);
or OR2 (N796, N793, N489);
not NOT1 (N797, N772);
not NOT1 (N798, N778);
and AND4 (N799, N794, N29, N376, N559);
xor XOR2 (N800, N799, N76);
buf BUF1 (N801, N798);
nand NAND2 (N802, N780, N202);
nor NOR2 (N803, N789, N614);
not NOT1 (N804, N803);
nor NOR2 (N805, N795, N378);
nor NOR2 (N806, N790, N457);
buf BUF1 (N807, N787);
not NOT1 (N808, N806);
xor XOR2 (N809, N800, N786);
nor NOR4 (N810, N777, N669, N771, N253);
not NOT1 (N811, N807);
and AND2 (N812, N804, N418);
and AND3 (N813, N810, N62, N242);
nand NAND4 (N814, N796, N55, N120, N236);
and AND4 (N815, N811, N86, N43, N810);
nand NAND2 (N816, N797, N346);
not NOT1 (N817, N805);
xor XOR2 (N818, N813, N266);
and AND4 (N819, N812, N535, N158, N42);
not NOT1 (N820, N814);
buf BUF1 (N821, N820);
not NOT1 (N822, N809);
and AND3 (N823, N802, N772, N516);
nor NOR4 (N824, N819, N132, N60, N333);
not NOT1 (N825, N801);
or OR4 (N826, N823, N782, N161, N643);
nor NOR2 (N827, N815, N490);
nand NAND2 (N828, N818, N549);
or OR3 (N829, N822, N685, N238);
and AND3 (N830, N821, N272, N482);
and AND4 (N831, N824, N370, N447, N649);
buf BUF1 (N832, N826);
not NOT1 (N833, N828);
or OR3 (N834, N817, N221, N344);
buf BUF1 (N835, N816);
xor XOR2 (N836, N834, N227);
and AND4 (N837, N835, N413, N721, N577);
nor NOR4 (N838, N830, N82, N643, N684);
not NOT1 (N839, N827);
buf BUF1 (N840, N829);
xor XOR2 (N841, N836, N343);
and AND2 (N842, N837, N812);
and AND4 (N843, N840, N750, N458, N627);
buf BUF1 (N844, N838);
and AND3 (N845, N842, N440, N385);
buf BUF1 (N846, N832);
buf BUF1 (N847, N833);
xor XOR2 (N848, N831, N780);
nor NOR2 (N849, N839, N842);
not NOT1 (N850, N808);
nor NOR2 (N851, N844, N679);
or OR4 (N852, N841, N147, N277, N706);
buf BUF1 (N853, N846);
buf BUF1 (N854, N851);
nand NAND4 (N855, N854, N37, N199, N742);
xor XOR2 (N856, N853, N385);
or OR3 (N857, N848, N747, N847);
or OR2 (N858, N87, N546);
nor NOR2 (N859, N849, N465);
nand NAND2 (N860, N859, N244);
buf BUF1 (N861, N843);
buf BUF1 (N862, N861);
or OR2 (N863, N850, N490);
or OR2 (N864, N858, N804);
or OR2 (N865, N825, N276);
buf BUF1 (N866, N855);
xor XOR2 (N867, N857, N516);
or OR4 (N868, N863, N557, N200, N553);
nor NOR2 (N869, N862, N449);
nand NAND3 (N870, N868, N353, N326);
not NOT1 (N871, N864);
or OR2 (N872, N856, N769);
or OR3 (N873, N867, N560, N95);
nand NAND4 (N874, N865, N368, N150, N631);
or OR3 (N875, N874, N739, N805);
and AND4 (N876, N873, N772, N460, N670);
or OR3 (N877, N852, N379, N489);
not NOT1 (N878, N871);
and AND4 (N879, N866, N553, N354, N693);
nand NAND3 (N880, N875, N671, N341);
nor NOR2 (N881, N860, N620);
nor NOR3 (N882, N881, N480, N256);
or OR4 (N883, N872, N284, N797, N769);
xor XOR2 (N884, N877, N415);
nor NOR4 (N885, N883, N392, N612, N347);
nand NAND4 (N886, N880, N160, N286, N444);
nand NAND2 (N887, N870, N440);
buf BUF1 (N888, N878);
nand NAND4 (N889, N879, N617, N796, N760);
and AND3 (N890, N885, N449, N252);
buf BUF1 (N891, N884);
xor XOR2 (N892, N869, N61);
nor NOR4 (N893, N892, N510, N558, N647);
nor NOR3 (N894, N890, N595, N798);
or OR4 (N895, N845, N670, N507, N802);
buf BUF1 (N896, N876);
and AND3 (N897, N896, N209, N788);
or OR4 (N898, N882, N207, N571, N758);
buf BUF1 (N899, N893);
nand NAND3 (N900, N886, N627, N871);
or OR3 (N901, N900, N55, N394);
xor XOR2 (N902, N895, N75);
nand NAND4 (N903, N891, N512, N595, N712);
nand NAND3 (N904, N899, N307, N347);
nand NAND2 (N905, N898, N214);
buf BUF1 (N906, N904);
and AND3 (N907, N889, N119, N71);
xor XOR2 (N908, N894, N535);
nand NAND2 (N909, N905, N448);
or OR4 (N910, N907, N150, N183, N288);
buf BUF1 (N911, N888);
or OR2 (N912, N897, N218);
or OR4 (N913, N910, N363, N674, N509);
and AND4 (N914, N911, N596, N455, N376);
nand NAND2 (N915, N913, N612);
nor NOR3 (N916, N906, N200, N282);
nand NAND2 (N917, N887, N379);
or OR3 (N918, N912, N690, N463);
not NOT1 (N919, N903);
not NOT1 (N920, N915);
or OR4 (N921, N918, N639, N628, N30);
or OR4 (N922, N917, N868, N104, N663);
and AND2 (N923, N901, N744);
nand NAND4 (N924, N922, N671, N765, N181);
nand NAND3 (N925, N909, N616, N96);
nor NOR2 (N926, N920, N305);
buf BUF1 (N927, N924);
xor XOR2 (N928, N925, N321);
not NOT1 (N929, N921);
nor NOR4 (N930, N923, N440, N94, N248);
or OR3 (N931, N927, N474, N515);
not NOT1 (N932, N902);
buf BUF1 (N933, N926);
or OR3 (N934, N930, N603, N690);
not NOT1 (N935, N934);
nand NAND3 (N936, N908, N301, N501);
or OR4 (N937, N928, N818, N113, N540);
nor NOR2 (N938, N929, N530);
nand NAND2 (N939, N937, N358);
or OR2 (N940, N914, N389);
buf BUF1 (N941, N935);
buf BUF1 (N942, N933);
and AND3 (N943, N932, N324, N166);
xor XOR2 (N944, N936, N352);
not NOT1 (N945, N941);
nor NOR4 (N946, N943, N539, N197, N202);
nand NAND4 (N947, N940, N218, N723, N553);
nand NAND2 (N948, N942, N315);
nor NOR3 (N949, N939, N551, N492);
nor NOR3 (N950, N948, N827, N379);
buf BUF1 (N951, N947);
nand NAND3 (N952, N938, N385, N859);
and AND3 (N953, N945, N44, N575);
or OR3 (N954, N944, N668, N344);
not NOT1 (N955, N951);
xor XOR2 (N956, N955, N225);
and AND3 (N957, N952, N846, N735);
nand NAND3 (N958, N949, N311, N527);
not NOT1 (N959, N953);
not NOT1 (N960, N950);
buf BUF1 (N961, N931);
and AND2 (N962, N916, N567);
buf BUF1 (N963, N919);
not NOT1 (N964, N956);
xor XOR2 (N965, N962, N650);
or OR4 (N966, N954, N744, N178, N53);
nor NOR3 (N967, N960, N368, N925);
not NOT1 (N968, N961);
or OR4 (N969, N957, N65, N628, N610);
and AND4 (N970, N946, N437, N195, N88);
xor XOR2 (N971, N969, N713);
not NOT1 (N972, N959);
or OR3 (N973, N966, N491, N620);
or OR4 (N974, N965, N574, N332, N780);
xor XOR2 (N975, N963, N53);
nor NOR2 (N976, N968, N281);
and AND2 (N977, N971, N700);
not NOT1 (N978, N973);
nor NOR2 (N979, N975, N856);
nor NOR4 (N980, N967, N357, N693, N397);
buf BUF1 (N981, N978);
xor XOR2 (N982, N964, N45);
or OR2 (N983, N972, N517);
or OR3 (N984, N981, N292, N874);
xor XOR2 (N985, N970, N765);
nand NAND3 (N986, N983, N464, N306);
xor XOR2 (N987, N977, N503);
not NOT1 (N988, N980);
nand NAND3 (N989, N974, N773, N446);
and AND4 (N990, N976, N329, N709, N846);
not NOT1 (N991, N990);
xor XOR2 (N992, N989, N65);
and AND4 (N993, N987, N585, N109, N311);
nor NOR4 (N994, N985, N966, N99, N983);
or OR4 (N995, N982, N156, N451, N563);
buf BUF1 (N996, N979);
or OR3 (N997, N991, N152, N868);
or OR4 (N998, N994, N825, N710, N84);
not NOT1 (N999, N988);
buf BUF1 (N1000, N999);
xor XOR2 (N1001, N997, N823);
nor NOR4 (N1002, N958, N122, N431, N889);
xor XOR2 (N1003, N1002, N820);
and AND4 (N1004, N1003, N738, N653, N843);
and AND4 (N1005, N1001, N796, N476, N74);
not NOT1 (N1006, N993);
and AND3 (N1007, N1004, N622, N357);
nand NAND3 (N1008, N1007, N957, N703);
and AND2 (N1009, N1008, N969);
nand NAND3 (N1010, N1009, N525, N993);
buf BUF1 (N1011, N992);
nor NOR3 (N1012, N1010, N703, N895);
nand NAND2 (N1013, N996, N776);
and AND3 (N1014, N1005, N489, N978);
nand NAND3 (N1015, N986, N527, N332);
xor XOR2 (N1016, N1006, N222);
nand NAND4 (N1017, N1012, N975, N779, N434);
nor NOR2 (N1018, N995, N539);
nand NAND4 (N1019, N998, N236, N125, N727);
nor NOR2 (N1020, N984, N654);
and AND3 (N1021, N1011, N192, N887);
buf BUF1 (N1022, N1014);
nand NAND3 (N1023, N1022, N960, N118);
and AND2 (N1024, N1019, N776);
not NOT1 (N1025, N1023);
xor XOR2 (N1026, N1020, N566);
nor NOR2 (N1027, N1016, N836);
nand NAND2 (N1028, N1015, N235);
nand NAND2 (N1029, N1021, N547);
nand NAND3 (N1030, N1026, N485, N332);
and AND3 (N1031, N1000, N929, N30);
not NOT1 (N1032, N1028);
not NOT1 (N1033, N1032);
nand NAND4 (N1034, N1027, N220, N59, N118);
nand NAND3 (N1035, N1018, N439, N642);
not NOT1 (N1036, N1035);
nand NAND4 (N1037, N1033, N305, N682, N814);
xor XOR2 (N1038, N1013, N707);
buf BUF1 (N1039, N1030);
xor XOR2 (N1040, N1039, N775);
xor XOR2 (N1041, N1017, N793);
or OR4 (N1042, N1038, N869, N131, N665);
xor XOR2 (N1043, N1029, N1006);
nor NOR4 (N1044, N1041, N153, N951, N85);
not NOT1 (N1045, N1040);
or OR3 (N1046, N1044, N173, N657);
buf BUF1 (N1047, N1031);
buf BUF1 (N1048, N1036);
not NOT1 (N1049, N1024);
and AND3 (N1050, N1047, N635, N785);
buf BUF1 (N1051, N1045);
nor NOR3 (N1052, N1046, N654, N347);
not NOT1 (N1053, N1051);
nor NOR2 (N1054, N1043, N750);
nand NAND2 (N1055, N1025, N102);
nand NAND4 (N1056, N1048, N728, N205, N740);
buf BUF1 (N1057, N1056);
not NOT1 (N1058, N1037);
buf BUF1 (N1059, N1042);
xor XOR2 (N1060, N1058, N574);
and AND3 (N1061, N1054, N514, N119);
nor NOR4 (N1062, N1057, N375, N325, N388);
xor XOR2 (N1063, N1049, N892);
buf BUF1 (N1064, N1059);
nor NOR3 (N1065, N1055, N115, N712);
or OR3 (N1066, N1052, N28, N661);
nor NOR2 (N1067, N1066, N761);
or OR2 (N1068, N1064, N154);
xor XOR2 (N1069, N1061, N249);
nor NOR2 (N1070, N1068, N442);
not NOT1 (N1071, N1065);
nor NOR3 (N1072, N1067, N680, N279);
nor NOR3 (N1073, N1034, N604, N748);
or OR2 (N1074, N1072, N537);
buf BUF1 (N1075, N1050);
buf BUF1 (N1076, N1074);
not NOT1 (N1077, N1063);
nor NOR2 (N1078, N1073, N476);
buf BUF1 (N1079, N1075);
or OR4 (N1080, N1062, N746, N13, N956);
nand NAND2 (N1081, N1076, N259);
and AND3 (N1082, N1080, N686, N369);
and AND3 (N1083, N1082, N75, N681);
buf BUF1 (N1084, N1053);
not NOT1 (N1085, N1083);
nand NAND3 (N1086, N1079, N439, N754);
buf BUF1 (N1087, N1070);
buf BUF1 (N1088, N1060);
nor NOR4 (N1089, N1085, N163, N1062, N396);
nand NAND3 (N1090, N1084, N225, N192);
buf BUF1 (N1091, N1069);
not NOT1 (N1092, N1091);
and AND2 (N1093, N1078, N758);
not NOT1 (N1094, N1090);
or OR4 (N1095, N1081, N1042, N620, N803);
xor XOR2 (N1096, N1077, N847);
nor NOR4 (N1097, N1088, N132, N826, N249);
nand NAND3 (N1098, N1087, N779, N942);
or OR3 (N1099, N1089, N239, N612);
buf BUF1 (N1100, N1093);
and AND2 (N1101, N1098, N264);
or OR4 (N1102, N1071, N759, N217, N59);
nand NAND3 (N1103, N1086, N442, N286);
nand NAND4 (N1104, N1092, N203, N777, N717);
buf BUF1 (N1105, N1094);
nand NAND2 (N1106, N1095, N641);
buf BUF1 (N1107, N1102);
xor XOR2 (N1108, N1105, N258);
not NOT1 (N1109, N1107);
not NOT1 (N1110, N1106);
buf BUF1 (N1111, N1109);
not NOT1 (N1112, N1111);
nand NAND2 (N1113, N1101, N1010);
nor NOR2 (N1114, N1103, N686);
buf BUF1 (N1115, N1113);
not NOT1 (N1116, N1099);
not NOT1 (N1117, N1115);
nor NOR3 (N1118, N1116, N625, N152);
xor XOR2 (N1119, N1096, N211);
nor NOR2 (N1120, N1104, N657);
buf BUF1 (N1121, N1114);
nand NAND2 (N1122, N1112, N275);
and AND4 (N1123, N1100, N370, N1022, N308);
and AND3 (N1124, N1097, N942, N536);
xor XOR2 (N1125, N1118, N264);
buf BUF1 (N1126, N1110);
and AND4 (N1127, N1117, N37, N626, N404);
buf BUF1 (N1128, N1122);
buf BUF1 (N1129, N1127);
buf BUF1 (N1130, N1119);
nor NOR2 (N1131, N1129, N360);
xor XOR2 (N1132, N1125, N137);
xor XOR2 (N1133, N1120, N565);
nor NOR2 (N1134, N1123, N1074);
buf BUF1 (N1135, N1108);
or OR4 (N1136, N1124, N620, N809, N1006);
and AND2 (N1137, N1136, N214);
nand NAND4 (N1138, N1135, N831, N454, N50);
nand NAND3 (N1139, N1131, N924, N175);
nor NOR3 (N1140, N1132, N589, N334);
nor NOR3 (N1141, N1140, N926, N126);
nand NAND2 (N1142, N1130, N56);
buf BUF1 (N1143, N1133);
buf BUF1 (N1144, N1141);
or OR4 (N1145, N1134, N526, N726, N825);
buf BUF1 (N1146, N1138);
and AND4 (N1147, N1126, N928, N272, N497);
not NOT1 (N1148, N1139);
nand NAND4 (N1149, N1145, N252, N645, N778);
not NOT1 (N1150, N1149);
not NOT1 (N1151, N1137);
nor NOR3 (N1152, N1143, N1057, N791);
nor NOR2 (N1153, N1152, N1134);
not NOT1 (N1154, N1153);
not NOT1 (N1155, N1147);
or OR3 (N1156, N1121, N462, N432);
and AND2 (N1157, N1156, N1100);
buf BUF1 (N1158, N1128);
and AND4 (N1159, N1150, N94, N419, N1036);
nor NOR3 (N1160, N1157, N863, N1089);
buf BUF1 (N1161, N1151);
not NOT1 (N1162, N1154);
and AND2 (N1163, N1158, N1086);
not NOT1 (N1164, N1163);
buf BUF1 (N1165, N1144);
nor NOR4 (N1166, N1164, N981, N1099, N332);
not NOT1 (N1167, N1159);
xor XOR2 (N1168, N1162, N400);
and AND3 (N1169, N1142, N998, N182);
nor NOR4 (N1170, N1160, N359, N1143, N917);
nor NOR2 (N1171, N1168, N472);
xor XOR2 (N1172, N1161, N479);
or OR3 (N1173, N1172, N422, N183);
not NOT1 (N1174, N1146);
buf BUF1 (N1175, N1174);
nand NAND3 (N1176, N1175, N639, N822);
not NOT1 (N1177, N1171);
and AND2 (N1178, N1155, N462);
or OR3 (N1179, N1167, N1164, N536);
xor XOR2 (N1180, N1176, N856);
buf BUF1 (N1181, N1148);
buf BUF1 (N1182, N1180);
buf BUF1 (N1183, N1178);
buf BUF1 (N1184, N1183);
and AND4 (N1185, N1169, N181, N1063, N811);
buf BUF1 (N1186, N1170);
buf BUF1 (N1187, N1177);
buf BUF1 (N1188, N1173);
or OR3 (N1189, N1187, N825, N500);
nor NOR4 (N1190, N1185, N70, N463, N337);
nor NOR2 (N1191, N1188, N763);
not NOT1 (N1192, N1166);
or OR2 (N1193, N1192, N990);
buf BUF1 (N1194, N1189);
buf BUF1 (N1195, N1179);
buf BUF1 (N1196, N1193);
or OR3 (N1197, N1181, N342, N1069);
nand NAND3 (N1198, N1197, N133, N748);
nand NAND2 (N1199, N1194, N916);
not NOT1 (N1200, N1165);
nor NOR2 (N1201, N1184, N523);
and AND2 (N1202, N1191, N660);
or OR4 (N1203, N1198, N1089, N883, N164);
or OR3 (N1204, N1196, N728, N1098);
not NOT1 (N1205, N1201);
buf BUF1 (N1206, N1202);
buf BUF1 (N1207, N1195);
buf BUF1 (N1208, N1204);
and AND2 (N1209, N1203, N590);
and AND3 (N1210, N1209, N244, N550);
nand NAND3 (N1211, N1207, N492, N125);
not NOT1 (N1212, N1206);
buf BUF1 (N1213, N1199);
and AND3 (N1214, N1211, N222, N871);
not NOT1 (N1215, N1182);
xor XOR2 (N1216, N1190, N432);
not NOT1 (N1217, N1210);
xor XOR2 (N1218, N1213, N718);
buf BUF1 (N1219, N1216);
xor XOR2 (N1220, N1217, N1025);
nor NOR3 (N1221, N1186, N913, N1013);
buf BUF1 (N1222, N1221);
nand NAND4 (N1223, N1200, N180, N961, N1002);
nand NAND4 (N1224, N1222, N788, N1063, N108);
or OR4 (N1225, N1219, N979, N551, N1);
buf BUF1 (N1226, N1223);
nor NOR4 (N1227, N1224, N747, N400, N395);
nand NAND3 (N1228, N1227, N613, N798);
or OR4 (N1229, N1220, N1063, N654, N809);
nand NAND3 (N1230, N1225, N1007, N46);
or OR3 (N1231, N1205, N278, N244);
buf BUF1 (N1232, N1214);
nand NAND2 (N1233, N1230, N116);
and AND4 (N1234, N1229, N1143, N631, N309);
nor NOR2 (N1235, N1234, N246);
and AND3 (N1236, N1218, N1015, N644);
and AND4 (N1237, N1228, N1078, N89, N137);
or OR3 (N1238, N1231, N1076, N473);
not NOT1 (N1239, N1208);
nand NAND2 (N1240, N1239, N588);
nand NAND4 (N1241, N1215, N1080, N848, N606);
nand NAND4 (N1242, N1237, N258, N1082, N35);
not NOT1 (N1243, N1232);
not NOT1 (N1244, N1212);
not NOT1 (N1245, N1243);
and AND4 (N1246, N1241, N884, N1154, N1154);
not NOT1 (N1247, N1238);
xor XOR2 (N1248, N1246, N661);
or OR3 (N1249, N1240, N822, N778);
nand NAND3 (N1250, N1233, N149, N1158);
nand NAND2 (N1251, N1236, N360);
and AND4 (N1252, N1247, N564, N554, N480);
and AND2 (N1253, N1235, N601);
nand NAND2 (N1254, N1248, N700);
not NOT1 (N1255, N1250);
xor XOR2 (N1256, N1255, N727);
or OR3 (N1257, N1226, N210, N941);
xor XOR2 (N1258, N1251, N815);
nand NAND3 (N1259, N1253, N1059, N196);
not NOT1 (N1260, N1258);
buf BUF1 (N1261, N1242);
not NOT1 (N1262, N1254);
and AND2 (N1263, N1257, N346);
or OR3 (N1264, N1263, N329, N895);
xor XOR2 (N1265, N1262, N246);
buf BUF1 (N1266, N1265);
not NOT1 (N1267, N1266);
nand NAND2 (N1268, N1245, N280);
buf BUF1 (N1269, N1249);
buf BUF1 (N1270, N1259);
not NOT1 (N1271, N1268);
nand NAND2 (N1272, N1261, N123);
xor XOR2 (N1273, N1260, N776);
nand NAND2 (N1274, N1252, N436);
and AND4 (N1275, N1267, N1141, N449, N333);
and AND2 (N1276, N1273, N1038);
and AND3 (N1277, N1271, N683, N1217);
nand NAND3 (N1278, N1276, N813, N297);
or OR4 (N1279, N1278, N247, N752, N48);
xor XOR2 (N1280, N1270, N1132);
xor XOR2 (N1281, N1279, N696);
xor XOR2 (N1282, N1277, N541);
buf BUF1 (N1283, N1256);
xor XOR2 (N1284, N1264, N499);
or OR2 (N1285, N1283, N264);
nor NOR3 (N1286, N1280, N1150, N18);
and AND2 (N1287, N1274, N502);
and AND3 (N1288, N1286, N967, N967);
or OR2 (N1289, N1285, N375);
nand NAND2 (N1290, N1244, N512);
and AND2 (N1291, N1289, N175);
buf BUF1 (N1292, N1281);
or OR4 (N1293, N1291, N161, N443, N955);
and AND2 (N1294, N1288, N1136);
nand NAND2 (N1295, N1290, N1004);
buf BUF1 (N1296, N1287);
and AND3 (N1297, N1293, N986, N832);
or OR3 (N1298, N1275, N934, N518);
not NOT1 (N1299, N1294);
and AND4 (N1300, N1298, N234, N650, N820);
nand NAND4 (N1301, N1272, N1205, N456, N26);
not NOT1 (N1302, N1295);
nor NOR2 (N1303, N1282, N314);
buf BUF1 (N1304, N1301);
xor XOR2 (N1305, N1303, N783);
and AND3 (N1306, N1302, N472, N846);
and AND2 (N1307, N1300, N920);
or OR2 (N1308, N1296, N175);
nor NOR3 (N1309, N1306, N410, N729);
nand NAND4 (N1310, N1269, N85, N346, N619);
or OR4 (N1311, N1305, N945, N1092, N1023);
nand NAND4 (N1312, N1304, N299, N668, N877);
xor XOR2 (N1313, N1310, N290);
buf BUF1 (N1314, N1308);
and AND3 (N1315, N1312, N857, N1087);
buf BUF1 (N1316, N1299);
nand NAND3 (N1317, N1309, N1059, N856);
nand NAND4 (N1318, N1317, N321, N512, N1243);
xor XOR2 (N1319, N1316, N1242);
and AND2 (N1320, N1314, N956);
or OR3 (N1321, N1284, N776, N581);
nor NOR4 (N1322, N1311, N969, N314, N1178);
xor XOR2 (N1323, N1292, N681);
and AND3 (N1324, N1297, N1072, N193);
nand NAND3 (N1325, N1323, N1224, N811);
or OR4 (N1326, N1318, N249, N600, N1127);
buf BUF1 (N1327, N1321);
buf BUF1 (N1328, N1322);
buf BUF1 (N1329, N1325);
buf BUF1 (N1330, N1324);
nand NAND3 (N1331, N1319, N1300, N1304);
buf BUF1 (N1332, N1313);
nor NOR4 (N1333, N1328, N1323, N551, N464);
xor XOR2 (N1334, N1331, N153);
not NOT1 (N1335, N1332);
and AND3 (N1336, N1330, N1174, N1245);
nor NOR3 (N1337, N1333, N736, N969);
or OR2 (N1338, N1336, N857);
nand NAND2 (N1339, N1334, N1122);
xor XOR2 (N1340, N1335, N1271);
or OR3 (N1341, N1327, N225, N529);
buf BUF1 (N1342, N1341);
buf BUF1 (N1343, N1329);
nor NOR2 (N1344, N1315, N62);
nand NAND3 (N1345, N1340, N1140, N1138);
nor NOR3 (N1346, N1320, N966, N1146);
or OR4 (N1347, N1346, N345, N1050, N460);
nand NAND4 (N1348, N1307, N393, N620, N252);
buf BUF1 (N1349, N1339);
nor NOR2 (N1350, N1342, N704);
buf BUF1 (N1351, N1343);
nor NOR2 (N1352, N1347, N154);
buf BUF1 (N1353, N1350);
not NOT1 (N1354, N1349);
nor NOR4 (N1355, N1337, N263, N597, N969);
nor NOR2 (N1356, N1354, N172);
or OR2 (N1357, N1338, N792);
xor XOR2 (N1358, N1351, N402);
or OR3 (N1359, N1357, N299, N989);
or OR2 (N1360, N1356, N242);
buf BUF1 (N1361, N1360);
nor NOR2 (N1362, N1361, N918);
nand NAND2 (N1363, N1362, N899);
nor NOR3 (N1364, N1353, N1201, N680);
and AND3 (N1365, N1348, N311, N787);
not NOT1 (N1366, N1345);
xor XOR2 (N1367, N1352, N420);
not NOT1 (N1368, N1364);
xor XOR2 (N1369, N1363, N688);
buf BUF1 (N1370, N1368);
not NOT1 (N1371, N1355);
and AND3 (N1372, N1358, N743, N234);
nand NAND2 (N1373, N1344, N1310);
not NOT1 (N1374, N1367);
nor NOR4 (N1375, N1366, N638, N195, N223);
nand NAND2 (N1376, N1373, N358);
xor XOR2 (N1377, N1371, N1304);
or OR3 (N1378, N1374, N1197, N837);
nand NAND3 (N1379, N1326, N108, N807);
buf BUF1 (N1380, N1370);
xor XOR2 (N1381, N1378, N247);
nor NOR3 (N1382, N1380, N229, N351);
or OR4 (N1383, N1381, N317, N843, N511);
nand NAND4 (N1384, N1376, N248, N1101, N476);
xor XOR2 (N1385, N1384, N947);
buf BUF1 (N1386, N1375);
buf BUF1 (N1387, N1365);
xor XOR2 (N1388, N1383, N810);
buf BUF1 (N1389, N1372);
not NOT1 (N1390, N1377);
nand NAND2 (N1391, N1359, N565);
xor XOR2 (N1392, N1386, N342);
nor NOR3 (N1393, N1382, N141, N136);
or OR3 (N1394, N1393, N1109, N481);
xor XOR2 (N1395, N1387, N552);
nor NOR2 (N1396, N1385, N160);
nand NAND3 (N1397, N1388, N677, N762);
buf BUF1 (N1398, N1392);
or OR2 (N1399, N1369, N763);
or OR3 (N1400, N1395, N277, N360);
xor XOR2 (N1401, N1389, N434);
and AND4 (N1402, N1398, N1178, N1291, N964);
nand NAND2 (N1403, N1401, N424);
or OR3 (N1404, N1400, N667, N293);
not NOT1 (N1405, N1402);
nand NAND4 (N1406, N1405, N857, N768, N131);
nor NOR3 (N1407, N1379, N1074, N925);
buf BUF1 (N1408, N1399);
nand NAND4 (N1409, N1403, N511, N1100, N504);
and AND2 (N1410, N1407, N876);
and AND3 (N1411, N1409, N1006, N436);
not NOT1 (N1412, N1390);
nand NAND2 (N1413, N1412, N1196);
or OR2 (N1414, N1404, N1062);
or OR2 (N1415, N1410, N774);
or OR4 (N1416, N1414, N1228, N37, N985);
nor NOR2 (N1417, N1406, N395);
nor NOR3 (N1418, N1397, N721, N170);
nand NAND3 (N1419, N1413, N1214, N358);
buf BUF1 (N1420, N1417);
nand NAND4 (N1421, N1396, N1115, N1048, N225);
xor XOR2 (N1422, N1420, N1172);
buf BUF1 (N1423, N1419);
nand NAND2 (N1424, N1408, N1018);
and AND4 (N1425, N1391, N108, N1066, N968);
and AND3 (N1426, N1421, N1311, N711);
not NOT1 (N1427, N1411);
nor NOR4 (N1428, N1424, N1074, N822, N1173);
nand NAND4 (N1429, N1428, N1034, N1214, N1233);
not NOT1 (N1430, N1394);
not NOT1 (N1431, N1429);
nand NAND3 (N1432, N1426, N779, N448);
and AND3 (N1433, N1432, N199, N1186);
and AND2 (N1434, N1418, N826);
nor NOR3 (N1435, N1427, N273, N818);
buf BUF1 (N1436, N1423);
and AND4 (N1437, N1436, N757, N673, N629);
or OR4 (N1438, N1425, N1272, N1031, N855);
xor XOR2 (N1439, N1430, N1299);
and AND3 (N1440, N1439, N999, N1305);
or OR2 (N1441, N1416, N318);
or OR2 (N1442, N1437, N6);
nand NAND3 (N1443, N1431, N615, N594);
nand NAND2 (N1444, N1440, N591);
nand NAND2 (N1445, N1444, N185);
buf BUF1 (N1446, N1435);
nor NOR4 (N1447, N1446, N981, N806, N908);
or OR3 (N1448, N1433, N876, N568);
or OR2 (N1449, N1438, N679);
nor NOR3 (N1450, N1448, N107, N823);
nand NAND2 (N1451, N1445, N1104);
xor XOR2 (N1452, N1441, N889);
or OR2 (N1453, N1447, N966);
nor NOR3 (N1454, N1450, N355, N143);
or OR2 (N1455, N1453, N1363);
not NOT1 (N1456, N1449);
buf BUF1 (N1457, N1454);
or OR4 (N1458, N1442, N541, N390, N645);
and AND4 (N1459, N1456, N760, N1090, N1205);
xor XOR2 (N1460, N1452, N1000);
not NOT1 (N1461, N1451);
nand NAND4 (N1462, N1415, N1189, N142, N849);
or OR2 (N1463, N1459, N1140);
and AND2 (N1464, N1462, N418);
or OR2 (N1465, N1443, N669);
or OR4 (N1466, N1463, N242, N373, N792);
or OR4 (N1467, N1466, N226, N625, N549);
nand NAND3 (N1468, N1464, N1062, N175);
nand NAND3 (N1469, N1434, N301, N508);
buf BUF1 (N1470, N1458);
xor XOR2 (N1471, N1465, N468);
xor XOR2 (N1472, N1471, N170);
nand NAND4 (N1473, N1468, N1391, N465, N806);
buf BUF1 (N1474, N1461);
buf BUF1 (N1475, N1472);
and AND4 (N1476, N1475, N58, N653, N102);
and AND4 (N1477, N1467, N1008, N303, N872);
not NOT1 (N1478, N1474);
nand NAND4 (N1479, N1470, N1432, N587, N436);
buf BUF1 (N1480, N1478);
buf BUF1 (N1481, N1460);
and AND4 (N1482, N1479, N1150, N531, N703);
buf BUF1 (N1483, N1469);
or OR4 (N1484, N1422, N409, N417, N786);
or OR3 (N1485, N1483, N544, N428);
and AND2 (N1486, N1480, N921);
xor XOR2 (N1487, N1481, N131);
and AND4 (N1488, N1473, N3, N1375, N1235);
nor NOR4 (N1489, N1487, N601, N701, N110);
buf BUF1 (N1490, N1489);
buf BUF1 (N1491, N1484);
xor XOR2 (N1492, N1476, N176);
and AND4 (N1493, N1477, N1161, N325, N573);
buf BUF1 (N1494, N1485);
xor XOR2 (N1495, N1486, N1405);
xor XOR2 (N1496, N1482, N1176);
and AND3 (N1497, N1496, N949, N1089);
or OR3 (N1498, N1494, N599, N910);
buf BUF1 (N1499, N1490);
nand NAND4 (N1500, N1488, N555, N534, N732);
or OR3 (N1501, N1457, N1257, N918);
xor XOR2 (N1502, N1495, N456);
xor XOR2 (N1503, N1491, N612);
not NOT1 (N1504, N1502);
nand NAND2 (N1505, N1499, N1343);
and AND4 (N1506, N1497, N1258, N528, N1327);
nand NAND3 (N1507, N1504, N860, N985);
nand NAND2 (N1508, N1501, N1240);
buf BUF1 (N1509, N1506);
xor XOR2 (N1510, N1508, N1014);
or OR3 (N1511, N1507, N1323, N1266);
buf BUF1 (N1512, N1500);
nor NOR2 (N1513, N1509, N1312);
or OR2 (N1514, N1510, N715);
and AND2 (N1515, N1514, N1152);
nor NOR3 (N1516, N1505, N834, N348);
xor XOR2 (N1517, N1512, N405);
xor XOR2 (N1518, N1503, N724);
and AND2 (N1519, N1492, N1031);
nand NAND4 (N1520, N1519, N866, N358, N702);
nor NOR4 (N1521, N1498, N607, N1437, N637);
xor XOR2 (N1522, N1515, N477);
and AND3 (N1523, N1517, N1190, N333);
xor XOR2 (N1524, N1516, N821);
nor NOR2 (N1525, N1513, N161);
or OR2 (N1526, N1493, N151);
not NOT1 (N1527, N1518);
nor NOR4 (N1528, N1511, N1231, N98, N1431);
nand NAND4 (N1529, N1525, N734, N699, N970);
xor XOR2 (N1530, N1526, N553);
and AND4 (N1531, N1520, N1440, N750, N1466);
xor XOR2 (N1532, N1455, N1349);
not NOT1 (N1533, N1522);
buf BUF1 (N1534, N1530);
nand NAND2 (N1535, N1521, N1370);
not NOT1 (N1536, N1524);
and AND4 (N1537, N1528, N41, N196, N1243);
not NOT1 (N1538, N1523);
buf BUF1 (N1539, N1532);
buf BUF1 (N1540, N1533);
nand NAND2 (N1541, N1534, N1363);
or OR4 (N1542, N1536, N506, N278, N1190);
nand NAND3 (N1543, N1541, N465, N1268);
not NOT1 (N1544, N1527);
or OR2 (N1545, N1543, N174);
buf BUF1 (N1546, N1539);
not NOT1 (N1547, N1538);
or OR3 (N1548, N1542, N1077, N897);
nand NAND4 (N1549, N1545, N606, N1038, N1197);
buf BUF1 (N1550, N1529);
and AND3 (N1551, N1531, N2, N954);
buf BUF1 (N1552, N1547);
nor NOR2 (N1553, N1551, N302);
and AND3 (N1554, N1553, N1085, N181);
xor XOR2 (N1555, N1552, N695);
not NOT1 (N1556, N1535);
or OR2 (N1557, N1540, N1158);
or OR2 (N1558, N1555, N170);
buf BUF1 (N1559, N1550);
or OR4 (N1560, N1537, N793, N805, N1285);
nand NAND3 (N1561, N1544, N756, N1163);
or OR3 (N1562, N1546, N141, N779);
xor XOR2 (N1563, N1562, N80);
nand NAND4 (N1564, N1548, N1302, N1378, N1330);
and AND2 (N1565, N1549, N1136);
not NOT1 (N1566, N1556);
not NOT1 (N1567, N1560);
nand NAND3 (N1568, N1565, N1021, N439);
not NOT1 (N1569, N1561);
nand NAND4 (N1570, N1564, N404, N769, N1028);
xor XOR2 (N1571, N1568, N1155);
xor XOR2 (N1572, N1554, N862);
and AND4 (N1573, N1567, N346, N367, N651);
nand NAND3 (N1574, N1569, N382, N228);
buf BUF1 (N1575, N1563);
xor XOR2 (N1576, N1572, N855);
not NOT1 (N1577, N1557);
nor NOR2 (N1578, N1566, N857);
buf BUF1 (N1579, N1576);
buf BUF1 (N1580, N1577);
not NOT1 (N1581, N1575);
and AND2 (N1582, N1580, N251);
nor NOR4 (N1583, N1571, N1293, N1369, N65);
not NOT1 (N1584, N1574);
nand NAND3 (N1585, N1558, N1440, N1039);
xor XOR2 (N1586, N1585, N920);
or OR2 (N1587, N1559, N630);
nand NAND4 (N1588, N1583, N1251, N1177, N1577);
or OR4 (N1589, N1588, N614, N713, N836);
nor NOR4 (N1590, N1578, N519, N551, N1522);
nor NOR3 (N1591, N1589, N78, N45);
nand NAND4 (N1592, N1582, N777, N794, N686);
not NOT1 (N1593, N1587);
nor NOR3 (N1594, N1593, N1373, N1017);
and AND4 (N1595, N1579, N745, N1164, N332);
nor NOR2 (N1596, N1595, N1172);
nor NOR3 (N1597, N1592, N203, N1072);
not NOT1 (N1598, N1581);
not NOT1 (N1599, N1596);
xor XOR2 (N1600, N1590, N774);
nor NOR2 (N1601, N1584, N1033);
nand NAND2 (N1602, N1573, N1217);
buf BUF1 (N1603, N1586);
nand NAND3 (N1604, N1598, N743, N589);
xor XOR2 (N1605, N1604, N86);
buf BUF1 (N1606, N1603);
not NOT1 (N1607, N1600);
nand NAND3 (N1608, N1602, N1078, N390);
buf BUF1 (N1609, N1601);
not NOT1 (N1610, N1591);
nor NOR2 (N1611, N1594, N687);
nor NOR3 (N1612, N1570, N1460, N455);
not NOT1 (N1613, N1599);
nor NOR3 (N1614, N1609, N393, N1420);
xor XOR2 (N1615, N1610, N1384);
nor NOR2 (N1616, N1608, N704);
buf BUF1 (N1617, N1612);
nand NAND2 (N1618, N1607, N194);
xor XOR2 (N1619, N1615, N686);
or OR4 (N1620, N1617, N764, N818, N453);
nand NAND2 (N1621, N1605, N316);
nand NAND2 (N1622, N1597, N553);
xor XOR2 (N1623, N1618, N1537);
not NOT1 (N1624, N1606);
not NOT1 (N1625, N1611);
and AND3 (N1626, N1622, N1172, N177);
and AND3 (N1627, N1620, N224, N37);
nor NOR3 (N1628, N1616, N579, N1063);
and AND3 (N1629, N1619, N78, N24);
not NOT1 (N1630, N1628);
not NOT1 (N1631, N1627);
nor NOR2 (N1632, N1614, N331);
nor NOR3 (N1633, N1626, N1078, N1283);
or OR3 (N1634, N1631, N1431, N360);
nor NOR2 (N1635, N1630, N273);
buf BUF1 (N1636, N1621);
nor NOR3 (N1637, N1613, N45, N1636);
nor NOR3 (N1638, N623, N141, N1159);
or OR3 (N1639, N1637, N1630, N24);
and AND4 (N1640, N1625, N1559, N1215, N296);
or OR2 (N1641, N1633, N586);
nand NAND3 (N1642, N1629, N910, N747);
buf BUF1 (N1643, N1623);
or OR4 (N1644, N1624, N1099, N415, N69);
and AND3 (N1645, N1634, N660, N578);
not NOT1 (N1646, N1638);
xor XOR2 (N1647, N1641, N1091);
buf BUF1 (N1648, N1639);
xor XOR2 (N1649, N1640, N1318);
or OR2 (N1650, N1649, N832);
or OR2 (N1651, N1632, N1207);
not NOT1 (N1652, N1646);
or OR4 (N1653, N1645, N438, N950, N1365);
xor XOR2 (N1654, N1650, N675);
nor NOR2 (N1655, N1642, N961);
nand NAND3 (N1656, N1644, N1378, N823);
or OR3 (N1657, N1654, N1182, N723);
nand NAND3 (N1658, N1651, N1158, N708);
not NOT1 (N1659, N1652);
xor XOR2 (N1660, N1656, N90);
xor XOR2 (N1661, N1660, N1533);
not NOT1 (N1662, N1643);
and AND2 (N1663, N1648, N1117);
or OR4 (N1664, N1662, N1130, N1019, N227);
xor XOR2 (N1665, N1663, N1586);
or OR4 (N1666, N1657, N477, N1097, N1040);
xor XOR2 (N1667, N1635, N733);
and AND4 (N1668, N1667, N1182, N318, N1335);
and AND3 (N1669, N1661, N1320, N1384);
and AND2 (N1670, N1658, N1622);
and AND4 (N1671, N1670, N616, N220, N187);
buf BUF1 (N1672, N1671);
buf BUF1 (N1673, N1666);
not NOT1 (N1674, N1659);
xor XOR2 (N1675, N1673, N1562);
nor NOR2 (N1676, N1647, N655);
and AND3 (N1677, N1668, N1188, N774);
nand NAND4 (N1678, N1677, N381, N944, N609);
xor XOR2 (N1679, N1672, N933);
and AND2 (N1680, N1679, N1311);
nand NAND3 (N1681, N1674, N509, N1354);
not NOT1 (N1682, N1655);
and AND2 (N1683, N1678, N33);
nor NOR2 (N1684, N1680, N483);
xor XOR2 (N1685, N1682, N129);
buf BUF1 (N1686, N1681);
buf BUF1 (N1687, N1683);
or OR4 (N1688, N1669, N1363, N266, N1480);
nand NAND2 (N1689, N1653, N686);
nor NOR3 (N1690, N1664, N1200, N216);
nand NAND2 (N1691, N1685, N820);
buf BUF1 (N1692, N1688);
nand NAND2 (N1693, N1686, N1527);
not NOT1 (N1694, N1675);
nor NOR3 (N1695, N1693, N1683, N1294);
nand NAND4 (N1696, N1687, N693, N655, N905);
nand NAND4 (N1697, N1696, N1340, N1439, N1144);
nor NOR4 (N1698, N1676, N267, N580, N776);
buf BUF1 (N1699, N1692);
and AND4 (N1700, N1699, N460, N892, N322);
and AND3 (N1701, N1684, N1698, N790);
buf BUF1 (N1702, N48);
buf BUF1 (N1703, N1700);
buf BUF1 (N1704, N1703);
or OR4 (N1705, N1665, N1233, N56, N109);
not NOT1 (N1706, N1705);
xor XOR2 (N1707, N1690, N1073);
and AND2 (N1708, N1691, N1629);
nor NOR2 (N1709, N1695, N156);
nand NAND4 (N1710, N1689, N1576, N1343, N170);
nand NAND2 (N1711, N1707, N667);
xor XOR2 (N1712, N1697, N220);
nor NOR3 (N1713, N1694, N480, N1015);
not NOT1 (N1714, N1711);
buf BUF1 (N1715, N1709);
nand NAND2 (N1716, N1713, N380);
xor XOR2 (N1717, N1701, N564);
not NOT1 (N1718, N1714);
and AND4 (N1719, N1704, N121, N763, N1080);
buf BUF1 (N1720, N1718);
buf BUF1 (N1721, N1717);
or OR3 (N1722, N1710, N1675, N1055);
nor NOR4 (N1723, N1716, N199, N27, N1578);
not NOT1 (N1724, N1708);
nand NAND4 (N1725, N1721, N113, N882, N1121);
nand NAND4 (N1726, N1702, N1314, N1319, N142);
nor NOR2 (N1727, N1722, N1213);
or OR3 (N1728, N1715, N239, N1345);
not NOT1 (N1729, N1706);
xor XOR2 (N1730, N1723, N530);
xor XOR2 (N1731, N1728, N434);
and AND4 (N1732, N1719, N1026, N185, N777);
and AND3 (N1733, N1732, N1046, N47);
not NOT1 (N1734, N1727);
not NOT1 (N1735, N1712);
or OR2 (N1736, N1731, N210);
nand NAND3 (N1737, N1726, N1165, N1567);
xor XOR2 (N1738, N1735, N1121);
nand NAND3 (N1739, N1733, N684, N102);
buf BUF1 (N1740, N1737);
xor XOR2 (N1741, N1729, N995);
not NOT1 (N1742, N1720);
or OR3 (N1743, N1742, N1027, N1082);
and AND3 (N1744, N1741, N182, N1686);
and AND2 (N1745, N1740, N1061);
nor NOR2 (N1746, N1744, N58);
and AND3 (N1747, N1730, N1244, N275);
nor NOR4 (N1748, N1738, N511, N1638, N628);
or OR3 (N1749, N1748, N1195, N225);
not NOT1 (N1750, N1734);
nand NAND3 (N1751, N1750, N523, N20);
nor NOR4 (N1752, N1725, N1607, N1702, N87);
buf BUF1 (N1753, N1752);
not NOT1 (N1754, N1746);
xor XOR2 (N1755, N1754, N677);
xor XOR2 (N1756, N1749, N58);
xor XOR2 (N1757, N1753, N1253);
xor XOR2 (N1758, N1736, N12);
or OR2 (N1759, N1756, N395);
nand NAND3 (N1760, N1758, N1370, N27);
xor XOR2 (N1761, N1745, N1415);
not NOT1 (N1762, N1761);
buf BUF1 (N1763, N1747);
or OR4 (N1764, N1739, N719, N516, N1567);
nor NOR4 (N1765, N1762, N256, N549, N342);
or OR2 (N1766, N1757, N403);
nor NOR4 (N1767, N1751, N1377, N659, N1454);
and AND4 (N1768, N1724, N940, N636, N1331);
and AND3 (N1769, N1743, N647, N423);
not NOT1 (N1770, N1764);
buf BUF1 (N1771, N1766);
and AND2 (N1772, N1765, N282);
and AND3 (N1773, N1759, N857, N717);
or OR4 (N1774, N1767, N952, N260, N1090);
xor XOR2 (N1775, N1774, N1080);
xor XOR2 (N1776, N1755, N421);
buf BUF1 (N1777, N1770);
or OR4 (N1778, N1773, N1724, N1357, N1636);
and AND4 (N1779, N1769, N853, N1247, N358);
or OR4 (N1780, N1778, N651, N1265, N428);
nand NAND4 (N1781, N1775, N1608, N1072, N191);
and AND4 (N1782, N1779, N847, N1365, N579);
nand NAND4 (N1783, N1780, N1746, N630, N1494);
xor XOR2 (N1784, N1772, N775);
buf BUF1 (N1785, N1771);
or OR4 (N1786, N1782, N601, N1305, N1427);
nand NAND3 (N1787, N1785, N1114, N212);
buf BUF1 (N1788, N1781);
xor XOR2 (N1789, N1777, N1761);
or OR3 (N1790, N1776, N1332, N139);
xor XOR2 (N1791, N1788, N694);
or OR2 (N1792, N1786, N7);
buf BUF1 (N1793, N1789);
and AND3 (N1794, N1760, N1032, N1426);
nor NOR2 (N1795, N1787, N1352);
or OR2 (N1796, N1795, N101);
xor XOR2 (N1797, N1784, N1637);
or OR4 (N1798, N1783, N1790, N375, N205);
nand NAND4 (N1799, N872, N555, N1104, N1497);
not NOT1 (N1800, N1768);
buf BUF1 (N1801, N1797);
and AND3 (N1802, N1793, N275, N358);
nor NOR2 (N1803, N1802, N1771);
and AND4 (N1804, N1796, N1319, N1388, N1037);
buf BUF1 (N1805, N1801);
nor NOR4 (N1806, N1805, N1385, N185, N943);
nand NAND4 (N1807, N1798, N997, N555, N683);
nor NOR4 (N1808, N1806, N824, N973, N844);
buf BUF1 (N1809, N1791);
nor NOR2 (N1810, N1799, N734);
or OR3 (N1811, N1810, N763, N684);
xor XOR2 (N1812, N1804, N1650);
buf BUF1 (N1813, N1800);
nand NAND4 (N1814, N1763, N111, N541, N1173);
not NOT1 (N1815, N1792);
not NOT1 (N1816, N1808);
xor XOR2 (N1817, N1811, N1235);
and AND3 (N1818, N1813, N945, N536);
not NOT1 (N1819, N1809);
not NOT1 (N1820, N1817);
and AND4 (N1821, N1818, N236, N1745, N545);
nand NAND3 (N1822, N1815, N479, N231);
nor NOR2 (N1823, N1812, N1213);
nand NAND3 (N1824, N1814, N250, N334);
and AND4 (N1825, N1822, N1199, N1163, N1038);
not NOT1 (N1826, N1825);
xor XOR2 (N1827, N1824, N858);
and AND2 (N1828, N1821, N1752);
xor XOR2 (N1829, N1816, N393);
or OR4 (N1830, N1820, N1699, N1800, N474);
or OR4 (N1831, N1829, N503, N1457, N1165);
nand NAND4 (N1832, N1803, N668, N587, N675);
and AND2 (N1833, N1828, N341);
not NOT1 (N1834, N1819);
not NOT1 (N1835, N1833);
nand NAND2 (N1836, N1832, N1495);
nor NOR2 (N1837, N1826, N101);
and AND2 (N1838, N1837, N1430);
nand NAND2 (N1839, N1831, N1019);
buf BUF1 (N1840, N1834);
xor XOR2 (N1841, N1836, N784);
xor XOR2 (N1842, N1839, N1507);
buf BUF1 (N1843, N1807);
not NOT1 (N1844, N1841);
nand NAND2 (N1845, N1827, N491);
xor XOR2 (N1846, N1840, N308);
nor NOR2 (N1847, N1843, N99);
nor NOR2 (N1848, N1823, N1184);
nor NOR4 (N1849, N1845, N349, N15, N489);
and AND2 (N1850, N1848, N1149);
buf BUF1 (N1851, N1842);
or OR2 (N1852, N1835, N1413);
and AND3 (N1853, N1849, N1058, N254);
nand NAND4 (N1854, N1850, N869, N1850, N1325);
buf BUF1 (N1855, N1852);
or OR2 (N1856, N1830, N810);
not NOT1 (N1857, N1853);
nor NOR2 (N1858, N1847, N1040);
not NOT1 (N1859, N1854);
not NOT1 (N1860, N1844);
or OR4 (N1861, N1860, N1152, N1402, N542);
not NOT1 (N1862, N1859);
or OR2 (N1863, N1858, N1782);
nand NAND4 (N1864, N1838, N1124, N72, N833);
buf BUF1 (N1865, N1864);
xor XOR2 (N1866, N1846, N325);
not NOT1 (N1867, N1865);
nor NOR3 (N1868, N1856, N615, N147);
xor XOR2 (N1869, N1862, N374);
or OR2 (N1870, N1869, N671);
not NOT1 (N1871, N1857);
not NOT1 (N1872, N1868);
xor XOR2 (N1873, N1867, N1750);
and AND2 (N1874, N1873, N217);
or OR3 (N1875, N1863, N186, N1264);
and AND3 (N1876, N1872, N1363, N121);
or OR4 (N1877, N1855, N900, N1320, N649);
buf BUF1 (N1878, N1870);
xor XOR2 (N1879, N1874, N1777);
xor XOR2 (N1880, N1875, N596);
buf BUF1 (N1881, N1871);
and AND2 (N1882, N1879, N1233);
and AND4 (N1883, N1878, N833, N379, N867);
nor NOR4 (N1884, N1877, N1142, N89, N1308);
nand NAND4 (N1885, N1794, N1090, N333, N312);
xor XOR2 (N1886, N1884, N1502);
or OR4 (N1887, N1885, N152, N12, N1532);
or OR3 (N1888, N1851, N819, N566);
not NOT1 (N1889, N1882);
buf BUF1 (N1890, N1861);
or OR3 (N1891, N1880, N1155, N1582);
buf BUF1 (N1892, N1876);
not NOT1 (N1893, N1892);
buf BUF1 (N1894, N1886);
not NOT1 (N1895, N1893);
or OR3 (N1896, N1895, N975, N577);
buf BUF1 (N1897, N1866);
nor NOR3 (N1898, N1890, N1548, N1253);
nand NAND4 (N1899, N1894, N1102, N468, N632);
not NOT1 (N1900, N1887);
xor XOR2 (N1901, N1899, N1334);
nand NAND4 (N1902, N1897, N1293, N27, N539);
and AND2 (N1903, N1902, N1156);
nor NOR3 (N1904, N1900, N1880, N1163);
xor XOR2 (N1905, N1888, N824);
buf BUF1 (N1906, N1896);
buf BUF1 (N1907, N1905);
or OR2 (N1908, N1904, N1323);
and AND3 (N1909, N1891, N355, N1461);
or OR4 (N1910, N1906, N1424, N1571, N521);
nor NOR2 (N1911, N1909, N996);
nand NAND2 (N1912, N1907, N582);
or OR3 (N1913, N1911, N453, N1353);
and AND4 (N1914, N1908, N202, N1218, N1769);
buf BUF1 (N1915, N1913);
buf BUF1 (N1916, N1914);
nor NOR2 (N1917, N1915, N782);
not NOT1 (N1918, N1912);
buf BUF1 (N1919, N1881);
or OR4 (N1920, N1901, N1404, N430, N1828);
buf BUF1 (N1921, N1889);
and AND3 (N1922, N1918, N980, N694);
or OR2 (N1923, N1920, N1229);
xor XOR2 (N1924, N1910, N604);
nand NAND3 (N1925, N1919, N875, N251);
or OR3 (N1926, N1924, N1434, N729);
nor NOR4 (N1927, N1925, N452, N98, N851);
nor NOR4 (N1928, N1923, N1536, N957, N118);
buf BUF1 (N1929, N1928);
or OR4 (N1930, N1927, N474, N289, N51);
nand NAND4 (N1931, N1903, N1827, N509, N600);
and AND4 (N1932, N1926, N332, N29, N1856);
buf BUF1 (N1933, N1883);
nand NAND2 (N1934, N1921, N570);
nor NOR4 (N1935, N1922, N1591, N741, N411);
and AND2 (N1936, N1930, N449);
or OR4 (N1937, N1931, N1504, N53, N1753);
nor NOR4 (N1938, N1916, N1881, N895, N1407);
and AND3 (N1939, N1929, N525, N1508);
or OR4 (N1940, N1939, N959, N1316, N1179);
xor XOR2 (N1941, N1917, N1711);
nor NOR4 (N1942, N1936, N106, N448, N1052);
nor NOR2 (N1943, N1940, N1753);
xor XOR2 (N1944, N1898, N594);
nand NAND2 (N1945, N1943, N344);
not NOT1 (N1946, N1942);
or OR3 (N1947, N1945, N619, N1776);
nor NOR3 (N1948, N1941, N959, N1050);
buf BUF1 (N1949, N1948);
buf BUF1 (N1950, N1949);
nand NAND4 (N1951, N1950, N542, N1372, N182);
not NOT1 (N1952, N1944);
and AND2 (N1953, N1933, N1584);
nand NAND2 (N1954, N1953, N1496);
buf BUF1 (N1955, N1946);
buf BUF1 (N1956, N1937);
buf BUF1 (N1957, N1935);
buf BUF1 (N1958, N1947);
buf BUF1 (N1959, N1955);
buf BUF1 (N1960, N1952);
buf BUF1 (N1961, N1960);
or OR4 (N1962, N1961, N525, N1032, N1360);
nor NOR2 (N1963, N1934, N564);
buf BUF1 (N1964, N1963);
nor NOR3 (N1965, N1959, N893, N810);
xor XOR2 (N1966, N1932, N1443);
nor NOR3 (N1967, N1966, N205, N1017);
not NOT1 (N1968, N1965);
nand NAND4 (N1969, N1938, N263, N1780, N675);
nand NAND4 (N1970, N1969, N1849, N66, N587);
nor NOR4 (N1971, N1970, N143, N814, N988);
nand NAND4 (N1972, N1967, N310, N1862, N213);
nand NAND2 (N1973, N1958, N1641);
and AND4 (N1974, N1971, N161, N945, N607);
buf BUF1 (N1975, N1964);
nand NAND4 (N1976, N1973, N976, N1735, N1726);
buf BUF1 (N1977, N1972);
xor XOR2 (N1978, N1975, N1650);
buf BUF1 (N1979, N1977);
xor XOR2 (N1980, N1978, N1383);
nand NAND2 (N1981, N1957, N574);
and AND3 (N1982, N1976, N23, N142);
nand NAND4 (N1983, N1980, N293, N61, N872);
and AND2 (N1984, N1979, N163);
nor NOR4 (N1985, N1954, N612, N1778, N307);
buf BUF1 (N1986, N1962);
xor XOR2 (N1987, N1986, N1204);
and AND4 (N1988, N1981, N1650, N660, N1798);
buf BUF1 (N1989, N1988);
or OR3 (N1990, N1987, N1731, N1249);
nand NAND4 (N1991, N1983, N374, N685, N902);
nand NAND3 (N1992, N1985, N1504, N215);
not NOT1 (N1993, N1990);
or OR4 (N1994, N1982, N1316, N1465, N1241);
not NOT1 (N1995, N1991);
and AND2 (N1996, N1995, N1032);
and AND4 (N1997, N1956, N447, N1193, N471);
xor XOR2 (N1998, N1984, N326);
or OR3 (N1999, N1968, N548, N1910);
buf BUF1 (N2000, N1974);
or OR2 (N2001, N1992, N757);
not NOT1 (N2002, N1989);
not NOT1 (N2003, N2000);
nand NAND2 (N2004, N1994, N1933);
xor XOR2 (N2005, N2003, N1493);
or OR4 (N2006, N1998, N750, N727, N1678);
buf BUF1 (N2007, N2005);
and AND4 (N2008, N2004, N1006, N1056, N1013);
buf BUF1 (N2009, N1997);
nor NOR3 (N2010, N2006, N1601, N491);
buf BUF1 (N2011, N2002);
buf BUF1 (N2012, N2008);
buf BUF1 (N2013, N2001);
and AND2 (N2014, N2009, N502);
xor XOR2 (N2015, N1996, N1834);
and AND2 (N2016, N1993, N749);
buf BUF1 (N2017, N2016);
nor NOR4 (N2018, N1999, N1367, N1513, N1991);
xor XOR2 (N2019, N2015, N948);
not NOT1 (N2020, N2013);
nand NAND2 (N2021, N2019, N487);
not NOT1 (N2022, N1951);
nand NAND3 (N2023, N2020, N1691, N1543);
xor XOR2 (N2024, N2022, N1406);
or OR3 (N2025, N2010, N1480, N150);
xor XOR2 (N2026, N2017, N1727);
or OR3 (N2027, N2007, N1644, N316);
nand NAND2 (N2028, N2026, N493);
not NOT1 (N2029, N2014);
nor NOR2 (N2030, N2024, N1743);
nor NOR4 (N2031, N2011, N1150, N246, N679);
and AND2 (N2032, N2012, N929);
xor XOR2 (N2033, N2028, N1439);
nor NOR4 (N2034, N2021, N1933, N5, N434);
buf BUF1 (N2035, N2031);
or OR3 (N2036, N2030, N1427, N704);
nand NAND3 (N2037, N2025, N1512, N609);
not NOT1 (N2038, N2032);
xor XOR2 (N2039, N2023, N1315);
not NOT1 (N2040, N2037);
buf BUF1 (N2041, N2035);
not NOT1 (N2042, N2040);
xor XOR2 (N2043, N2029, N104);
nor NOR2 (N2044, N2018, N1762);
xor XOR2 (N2045, N2036, N84);
nand NAND4 (N2046, N2043, N199, N1167, N794);
not NOT1 (N2047, N2038);
buf BUF1 (N2048, N2041);
nor NOR4 (N2049, N2044, N981, N1219, N715);
nor NOR4 (N2050, N2039, N1320, N120, N395);
buf BUF1 (N2051, N2042);
nand NAND2 (N2052, N2046, N1600);
xor XOR2 (N2053, N2048, N1397);
nand NAND4 (N2054, N2053, N1620, N1372, N117);
nor NOR4 (N2055, N2034, N960, N1105, N1523);
nand NAND3 (N2056, N2054, N551, N101);
nor NOR4 (N2057, N2049, N482, N932, N72);
and AND2 (N2058, N2027, N1689);
xor XOR2 (N2059, N2057, N930);
nand NAND2 (N2060, N2052, N450);
or OR4 (N2061, N2050, N1955, N878, N637);
and AND4 (N2062, N2033, N72, N1322, N43);
not NOT1 (N2063, N2060);
not NOT1 (N2064, N2059);
or OR4 (N2065, N2047, N1757, N1764, N905);
nand NAND4 (N2066, N2065, N545, N1339, N971);
nor NOR2 (N2067, N2062, N1673);
nor NOR4 (N2068, N2067, N1870, N88, N225);
not NOT1 (N2069, N2051);
buf BUF1 (N2070, N2061);
nand NAND3 (N2071, N2058, N1723, N1940);
nor NOR3 (N2072, N2070, N905, N558);
xor XOR2 (N2073, N2045, N449);
nand NAND3 (N2074, N2071, N259, N2055);
xor XOR2 (N2075, N774, N339);
xor XOR2 (N2076, N2074, N2016);
nand NAND3 (N2077, N2064, N314, N1266);
buf BUF1 (N2078, N2063);
buf BUF1 (N2079, N2076);
not NOT1 (N2080, N2072);
nor NOR3 (N2081, N2080, N1005, N436);
nor NOR4 (N2082, N2068, N719, N980, N976);
or OR3 (N2083, N2081, N22, N927);
buf BUF1 (N2084, N2077);
nand NAND2 (N2085, N2073, N590);
or OR4 (N2086, N2078, N1737, N1794, N2058);
nor NOR3 (N2087, N2066, N154, N45);
buf BUF1 (N2088, N2069);
xor XOR2 (N2089, N2087, N1158);
buf BUF1 (N2090, N2056);
not NOT1 (N2091, N2089);
buf BUF1 (N2092, N2090);
and AND2 (N2093, N2092, N1873);
xor XOR2 (N2094, N2079, N935);
buf BUF1 (N2095, N2084);
nor NOR4 (N2096, N2085, N432, N920, N1308);
and AND4 (N2097, N2094, N1892, N2050, N758);
nor NOR4 (N2098, N2088, N490, N1219, N384);
or OR3 (N2099, N2096, N451, N290);
and AND3 (N2100, N2095, N954, N1885);
nor NOR3 (N2101, N2075, N1372, N39);
buf BUF1 (N2102, N2098);
and AND4 (N2103, N2093, N1495, N196, N1875);
xor XOR2 (N2104, N2100, N287);
and AND2 (N2105, N2097, N585);
buf BUF1 (N2106, N2103);
nand NAND4 (N2107, N2099, N1519, N1241, N982);
nand NAND3 (N2108, N2091, N1377, N1543);
and AND2 (N2109, N2107, N704);
nand NAND4 (N2110, N2105, N1726, N760, N439);
xor XOR2 (N2111, N2109, N210);
xor XOR2 (N2112, N2111, N1068);
nor NOR2 (N2113, N2086, N838);
buf BUF1 (N2114, N2110);
xor XOR2 (N2115, N2102, N293);
nor NOR4 (N2116, N2115, N1382, N887, N1082);
or OR2 (N2117, N2106, N7);
and AND3 (N2118, N2114, N111, N499);
xor XOR2 (N2119, N2101, N1561);
not NOT1 (N2120, N2108);
buf BUF1 (N2121, N2104);
xor XOR2 (N2122, N2118, N1931);
buf BUF1 (N2123, N2122);
and AND2 (N2124, N2121, N307);
and AND4 (N2125, N2083, N907, N546, N399);
nand NAND3 (N2126, N2116, N445, N240);
or OR3 (N2127, N2113, N1188, N1527);
not NOT1 (N2128, N2127);
nor NOR4 (N2129, N2128, N324, N772, N453);
or OR3 (N2130, N2124, N36, N1861);
or OR4 (N2131, N2117, N1430, N1884, N669);
and AND3 (N2132, N2112, N1456, N88);
and AND3 (N2133, N2123, N1858, N113);
not NOT1 (N2134, N2120);
or OR4 (N2135, N2126, N1075, N1724, N434);
not NOT1 (N2136, N2132);
and AND3 (N2137, N2133, N1569, N185);
not NOT1 (N2138, N2129);
nand NAND2 (N2139, N2082, N1158);
nand NAND4 (N2140, N2137, N1935, N954, N514);
xor XOR2 (N2141, N2131, N501);
buf BUF1 (N2142, N2136);
or OR4 (N2143, N2135, N245, N743, N398);
nor NOR3 (N2144, N2140, N1119, N1278);
not NOT1 (N2145, N2144);
not NOT1 (N2146, N2139);
buf BUF1 (N2147, N2141);
nor NOR3 (N2148, N2130, N698, N547);
buf BUF1 (N2149, N2146);
buf BUF1 (N2150, N2145);
xor XOR2 (N2151, N2148, N1625);
nand NAND3 (N2152, N2150, N2146, N788);
not NOT1 (N2153, N2151);
nor NOR3 (N2154, N2143, N1319, N811);
buf BUF1 (N2155, N2149);
or OR4 (N2156, N2154, N2009, N1989, N1929);
and AND2 (N2157, N2142, N1042);
nor NOR3 (N2158, N2153, N1423, N177);
xor XOR2 (N2159, N2152, N1628);
or OR4 (N2160, N2156, N2, N1631, N1427);
or OR2 (N2161, N2157, N2156);
or OR3 (N2162, N2134, N263, N2036);
and AND4 (N2163, N2155, N1479, N921, N1751);
or OR2 (N2164, N2138, N73);
nor NOR4 (N2165, N2160, N72, N4, N147);
or OR2 (N2166, N2165, N222);
nand NAND3 (N2167, N2161, N361, N1201);
nand NAND3 (N2168, N2163, N1685, N228);
xor XOR2 (N2169, N2119, N841);
or OR3 (N2170, N2164, N620, N431);
not NOT1 (N2171, N2158);
nand NAND3 (N2172, N2169, N2131, N302);
not NOT1 (N2173, N2172);
or OR4 (N2174, N2159, N407, N665, N2125);
or OR4 (N2175, N517, N1479, N130, N197);
buf BUF1 (N2176, N2171);
nand NAND3 (N2177, N2168, N550, N457);
not NOT1 (N2178, N2166);
xor XOR2 (N2179, N2147, N453);
nor NOR4 (N2180, N2173, N1090, N1259, N1877);
buf BUF1 (N2181, N2178);
and AND2 (N2182, N2181, N2045);
xor XOR2 (N2183, N2182, N78);
nand NAND2 (N2184, N2162, N508);
nor NOR2 (N2185, N2183, N675);
and AND4 (N2186, N2179, N158, N244, N561);
nor NOR3 (N2187, N2176, N595, N145);
xor XOR2 (N2188, N2174, N1099);
xor XOR2 (N2189, N2184, N1022);
nor NOR2 (N2190, N2180, N2059);
xor XOR2 (N2191, N2167, N666);
not NOT1 (N2192, N2170);
and AND3 (N2193, N2187, N991, N7);
not NOT1 (N2194, N2190);
or OR4 (N2195, N2175, N365, N1101, N814);
nor NOR2 (N2196, N2194, N934);
not NOT1 (N2197, N2191);
and AND3 (N2198, N2197, N1883, N1634);
and AND2 (N2199, N2189, N1434);
and AND2 (N2200, N2196, N844);
xor XOR2 (N2201, N2185, N666);
or OR4 (N2202, N2199, N929, N1695, N661);
buf BUF1 (N2203, N2193);
or OR4 (N2204, N2198, N1697, N88, N1874);
or OR3 (N2205, N2186, N1135, N385);
or OR4 (N2206, N2203, N391, N2198, N469);
and AND3 (N2207, N2192, N767, N1888);
xor XOR2 (N2208, N2200, N1415);
buf BUF1 (N2209, N2201);
buf BUF1 (N2210, N2207);
xor XOR2 (N2211, N2208, N1703);
and AND4 (N2212, N2205, N1954, N1565, N1608);
or OR3 (N2213, N2202, N1069, N1264);
nor NOR2 (N2214, N2177, N480);
xor XOR2 (N2215, N2195, N273);
nor NOR4 (N2216, N2209, N2076, N1717, N480);
nand NAND3 (N2217, N2214, N62, N399);
nand NAND4 (N2218, N2217, N1178, N1367, N487);
not NOT1 (N2219, N2218);
not NOT1 (N2220, N2204);
nand NAND4 (N2221, N2213, N305, N650, N2039);
or OR2 (N2222, N2211, N1291);
or OR4 (N2223, N2219, N22, N1981, N1181);
and AND3 (N2224, N2221, N1691, N1715);
not NOT1 (N2225, N2212);
buf BUF1 (N2226, N2224);
and AND2 (N2227, N2216, N2062);
nand NAND2 (N2228, N2222, N397);
or OR4 (N2229, N2215, N942, N71, N184);
xor XOR2 (N2230, N2229, N1088);
not NOT1 (N2231, N2223);
or OR2 (N2232, N2226, N1302);
not NOT1 (N2233, N2232);
or OR4 (N2234, N2231, N1342, N448, N567);
nand NAND2 (N2235, N2233, N1924);
xor XOR2 (N2236, N2220, N1429);
and AND2 (N2237, N2228, N1707);
not NOT1 (N2238, N2235);
and AND2 (N2239, N2236, N194);
nand NAND3 (N2240, N2238, N759, N1375);
or OR4 (N2241, N2237, N318, N309, N1786);
buf BUF1 (N2242, N2234);
not NOT1 (N2243, N2240);
or OR4 (N2244, N2188, N867, N663, N1323);
and AND2 (N2245, N2206, N1101);
and AND3 (N2246, N2230, N2145, N1702);
buf BUF1 (N2247, N2241);
xor XOR2 (N2248, N2210, N826);
xor XOR2 (N2249, N2225, N1017);
or OR3 (N2250, N2249, N2157, N2080);
or OR2 (N2251, N2227, N1149);
buf BUF1 (N2252, N2243);
xor XOR2 (N2253, N2239, N1531);
nand NAND4 (N2254, N2242, N2210, N2099, N434);
xor XOR2 (N2255, N2251, N927);
not NOT1 (N2256, N2253);
nor NOR3 (N2257, N2244, N1159, N2044);
not NOT1 (N2258, N2250);
nor NOR4 (N2259, N2247, N835, N697, N507);
and AND3 (N2260, N2259, N1616, N1667);
and AND3 (N2261, N2258, N1740, N1381);
or OR3 (N2262, N2257, N1405, N2253);
buf BUF1 (N2263, N2254);
xor XOR2 (N2264, N2248, N1215);
xor XOR2 (N2265, N2245, N2064);
nand NAND4 (N2266, N2264, N1859, N831, N854);
and AND3 (N2267, N2266, N1945, N2186);
xor XOR2 (N2268, N2263, N744);
nor NOR3 (N2269, N2256, N1655, N1786);
xor XOR2 (N2270, N2261, N804);
and AND3 (N2271, N2260, N1922, N1247);
not NOT1 (N2272, N2271);
nor NOR4 (N2273, N2255, N198, N1202, N2007);
nand NAND4 (N2274, N2273, N2115, N667, N1925);
nand NAND4 (N2275, N2246, N1080, N1546, N1937);
and AND4 (N2276, N2275, N646, N2067, N1048);
nor NOR3 (N2277, N2274, N1628, N1720);
nand NAND2 (N2278, N2270, N189);
xor XOR2 (N2279, N2278, N1589);
not NOT1 (N2280, N2269);
buf BUF1 (N2281, N2280);
not NOT1 (N2282, N2279);
buf BUF1 (N2283, N2272);
xor XOR2 (N2284, N2267, N1925);
nor NOR4 (N2285, N2282, N1992, N858, N828);
or OR3 (N2286, N2268, N167, N2097);
nand NAND3 (N2287, N2284, N1272, N109);
and AND2 (N2288, N2265, N1554);
and AND4 (N2289, N2281, N1122, N745, N1065);
nor NOR4 (N2290, N2262, N499, N44, N375);
or OR4 (N2291, N2277, N944, N34, N1510);
xor XOR2 (N2292, N2285, N1525);
not NOT1 (N2293, N2276);
not NOT1 (N2294, N2289);
not NOT1 (N2295, N2293);
or OR2 (N2296, N2283, N1404);
nand NAND3 (N2297, N2296, N1084, N1473);
and AND4 (N2298, N2288, N1635, N1805, N1366);
xor XOR2 (N2299, N2286, N1304);
buf BUF1 (N2300, N2294);
xor XOR2 (N2301, N2287, N494);
nor NOR4 (N2302, N2299, N451, N1974, N839);
and AND3 (N2303, N2291, N834, N1130);
xor XOR2 (N2304, N2252, N1115);
not NOT1 (N2305, N2298);
nand NAND3 (N2306, N2303, N1978, N993);
and AND4 (N2307, N2297, N27, N282, N2084);
xor XOR2 (N2308, N2290, N1903);
or OR3 (N2309, N2300, N1233, N122);
nor NOR4 (N2310, N2295, N1689, N117, N1175);
nor NOR3 (N2311, N2310, N1430, N570);
or OR4 (N2312, N2311, N224, N328, N1469);
not NOT1 (N2313, N2301);
nand NAND4 (N2314, N2304, N568, N897, N465);
and AND2 (N2315, N2302, N2011);
buf BUF1 (N2316, N2313);
xor XOR2 (N2317, N2305, N1084);
or OR2 (N2318, N2314, N2115);
and AND2 (N2319, N2309, N667);
xor XOR2 (N2320, N2319, N2128);
not NOT1 (N2321, N2315);
or OR2 (N2322, N2318, N5);
xor XOR2 (N2323, N2316, N612);
buf BUF1 (N2324, N2308);
nor NOR2 (N2325, N2321, N916);
and AND4 (N2326, N2322, N793, N1483, N1718);
nand NAND3 (N2327, N2292, N56, N67);
buf BUF1 (N2328, N2317);
buf BUF1 (N2329, N2320);
not NOT1 (N2330, N2327);
nor NOR4 (N2331, N2307, N101, N1281, N1505);
and AND3 (N2332, N2330, N1906, N495);
buf BUF1 (N2333, N2312);
nor NOR4 (N2334, N2331, N1615, N1528, N336);
not NOT1 (N2335, N2325);
and AND3 (N2336, N2326, N660, N649);
or OR2 (N2337, N2336, N305);
or OR4 (N2338, N2306, N1987, N1325, N2212);
xor XOR2 (N2339, N2324, N2061);
nand NAND2 (N2340, N2333, N1363);
nand NAND3 (N2341, N2340, N1554, N1754);
nor NOR2 (N2342, N2332, N869);
and AND2 (N2343, N2329, N310);
xor XOR2 (N2344, N2338, N938);
xor XOR2 (N2345, N2337, N2328);
not NOT1 (N2346, N661);
buf BUF1 (N2347, N2342);
or OR3 (N2348, N2347, N995, N2259);
or OR2 (N2349, N2343, N273);
or OR2 (N2350, N2348, N2024);
nand NAND2 (N2351, N2341, N594);
nor NOR3 (N2352, N2344, N1988, N789);
xor XOR2 (N2353, N2349, N2146);
xor XOR2 (N2354, N2346, N1265);
not NOT1 (N2355, N2352);
not NOT1 (N2356, N2351);
nor NOR3 (N2357, N2335, N359, N497);
xor XOR2 (N2358, N2345, N391);
buf BUF1 (N2359, N2323);
xor XOR2 (N2360, N2334, N968);
and AND2 (N2361, N2360, N525);
buf BUF1 (N2362, N2357);
and AND3 (N2363, N2339, N24, N1652);
nand NAND3 (N2364, N2362, N962, N300);
and AND3 (N2365, N2350, N1342, N2112);
buf BUF1 (N2366, N2354);
nand NAND3 (N2367, N2366, N959, N331);
nor NOR3 (N2368, N2365, N404, N1670);
buf BUF1 (N2369, N2363);
and AND2 (N2370, N2359, N1154);
nor NOR4 (N2371, N2370, N609, N1658, N1678);
or OR2 (N2372, N2367, N1412);
xor XOR2 (N2373, N2355, N2088);
xor XOR2 (N2374, N2361, N1885);
xor XOR2 (N2375, N2373, N1045);
not NOT1 (N2376, N2374);
and AND4 (N2377, N2371, N1782, N1059, N613);
nor NOR4 (N2378, N2353, N790, N1976, N1898);
buf BUF1 (N2379, N2358);
not NOT1 (N2380, N2378);
nor NOR3 (N2381, N2376, N973, N143);
nor NOR3 (N2382, N2380, N670, N1571);
not NOT1 (N2383, N2381);
xor XOR2 (N2384, N2382, N1688);
nor NOR3 (N2385, N2369, N2365, N430);
xor XOR2 (N2386, N2385, N626);
nor NOR2 (N2387, N2368, N896);
xor XOR2 (N2388, N2377, N1620);
nor NOR2 (N2389, N2356, N2353);
and AND3 (N2390, N2384, N2043, N1191);
and AND3 (N2391, N2379, N1121, N642);
buf BUF1 (N2392, N2390);
and AND4 (N2393, N2388, N2149, N615, N1420);
and AND4 (N2394, N2392, N2051, N1114, N1666);
nor NOR4 (N2395, N2391, N757, N850, N1117);
or OR3 (N2396, N2383, N1901, N761);
and AND3 (N2397, N2393, N1076, N2016);
and AND2 (N2398, N2394, N749);
nand NAND3 (N2399, N2386, N1968, N1920);
nand NAND3 (N2400, N2387, N433, N1342);
nor NOR3 (N2401, N2375, N1665, N163);
xor XOR2 (N2402, N2395, N1745);
nand NAND4 (N2403, N2396, N1513, N705, N312);
buf BUF1 (N2404, N2372);
nand NAND3 (N2405, N2403, N1151, N854);
or OR3 (N2406, N2401, N1563, N1444);
nor NOR4 (N2407, N2404, N635, N1076, N1710);
buf BUF1 (N2408, N2400);
and AND3 (N2409, N2402, N1339, N1501);
xor XOR2 (N2410, N2407, N2399);
nor NOR4 (N2411, N65, N893, N1536, N1130);
not NOT1 (N2412, N2389);
or OR4 (N2413, N2410, N1335, N1848, N775);
and AND3 (N2414, N2412, N1926, N2194);
buf BUF1 (N2415, N2364);
xor XOR2 (N2416, N2408, N564);
buf BUF1 (N2417, N2414);
nor NOR3 (N2418, N2411, N1438, N505);
nor NOR4 (N2419, N2405, N232, N2392, N1596);
not NOT1 (N2420, N2406);
xor XOR2 (N2421, N2420, N205);
xor XOR2 (N2422, N2409, N243);
nand NAND2 (N2423, N2417, N1303);
buf BUF1 (N2424, N2421);
not NOT1 (N2425, N2424);
xor XOR2 (N2426, N2419, N1643);
not NOT1 (N2427, N2425);
nand NAND2 (N2428, N2422, N217);
nor NOR3 (N2429, N2427, N2279, N1029);
nand NAND4 (N2430, N2397, N830, N2240, N121);
buf BUF1 (N2431, N2418);
not NOT1 (N2432, N2415);
or OR4 (N2433, N2423, N998, N1655, N2326);
not NOT1 (N2434, N2428);
xor XOR2 (N2435, N2434, N892);
not NOT1 (N2436, N2426);
xor XOR2 (N2437, N2430, N1643);
nor NOR2 (N2438, N2432, N1856);
buf BUF1 (N2439, N2431);
nor NOR2 (N2440, N2398, N2232);
buf BUF1 (N2441, N2438);
nor NOR2 (N2442, N2435, N996);
or OR2 (N2443, N2442, N1233);
nand NAND3 (N2444, N2429, N1738, N241);
and AND4 (N2445, N2439, N517, N409, N2274);
buf BUF1 (N2446, N2416);
and AND2 (N2447, N2446, N245);
not NOT1 (N2448, N2444);
and AND4 (N2449, N2443, N246, N1208, N1842);
and AND3 (N2450, N2440, N717, N1315);
nor NOR4 (N2451, N2441, N1911, N44, N1935);
or OR4 (N2452, N2451, N1706, N1375, N1025);
or OR4 (N2453, N2449, N2298, N481, N1942);
nor NOR2 (N2454, N2448, N71);
and AND3 (N2455, N2454, N169, N1768);
or OR4 (N2456, N2445, N205, N1548, N270);
xor XOR2 (N2457, N2447, N451);
and AND2 (N2458, N2437, N981);
or OR4 (N2459, N2458, N1756, N2133, N2087);
and AND3 (N2460, N2436, N1658, N48);
nand NAND4 (N2461, N2460, N2326, N419, N1801);
buf BUF1 (N2462, N2459);
or OR2 (N2463, N2461, N1296);
or OR4 (N2464, N2453, N742, N165, N1780);
nand NAND2 (N2465, N2433, N1344);
buf BUF1 (N2466, N2450);
or OR3 (N2467, N2452, N471, N1238);
xor XOR2 (N2468, N2463, N511);
nand NAND4 (N2469, N2464, N463, N2056, N449);
nand NAND2 (N2470, N2466, N1856);
nand NAND4 (N2471, N2462, N132, N1143, N212);
not NOT1 (N2472, N2413);
nor NOR3 (N2473, N2469, N830, N1383);
buf BUF1 (N2474, N2473);
nor NOR2 (N2475, N2472, N1512);
not NOT1 (N2476, N2467);
or OR3 (N2477, N2474, N2440, N2019);
nor NOR2 (N2478, N2468, N803);
buf BUF1 (N2479, N2456);
buf BUF1 (N2480, N2479);
and AND3 (N2481, N2477, N1396, N1509);
nor NOR2 (N2482, N2457, N1653);
and AND3 (N2483, N2455, N1371, N1011);
nand NAND3 (N2484, N2478, N1334, N536);
nor NOR3 (N2485, N2480, N13, N1739);
not NOT1 (N2486, N2465);
xor XOR2 (N2487, N2475, N1441);
nand NAND3 (N2488, N2476, N818, N785);
and AND2 (N2489, N2486, N2252);
and AND4 (N2490, N2482, N151, N779, N1078);
not NOT1 (N2491, N2485);
nor NOR2 (N2492, N2487, N2480);
xor XOR2 (N2493, N2492, N1624);
nand NAND4 (N2494, N2488, N384, N571, N1492);
nand NAND4 (N2495, N2484, N1492, N2172, N582);
nand NAND2 (N2496, N2494, N2186);
nand NAND4 (N2497, N2470, N197, N1915, N1906);
buf BUF1 (N2498, N2493);
xor XOR2 (N2499, N2498, N1151);
or OR4 (N2500, N2490, N41, N1261, N1670);
not NOT1 (N2501, N2471);
nor NOR4 (N2502, N2496, N671, N1501, N169);
buf BUF1 (N2503, N2501);
nand NAND2 (N2504, N2497, N421);
xor XOR2 (N2505, N2503, N842);
xor XOR2 (N2506, N2500, N839);
not NOT1 (N2507, N2495);
or OR4 (N2508, N2504, N433, N2039, N319);
nor NOR4 (N2509, N2502, N1564, N226, N881);
buf BUF1 (N2510, N2489);
and AND4 (N2511, N2481, N1012, N920, N2155);
not NOT1 (N2512, N2506);
buf BUF1 (N2513, N2483);
nor NOR2 (N2514, N2509, N78);
not NOT1 (N2515, N2499);
buf BUF1 (N2516, N2513);
nand NAND2 (N2517, N2507, N2357);
nor NOR4 (N2518, N2514, N1628, N2076, N2486);
buf BUF1 (N2519, N2515);
not NOT1 (N2520, N2491);
or OR2 (N2521, N2510, N1383);
buf BUF1 (N2522, N2508);
not NOT1 (N2523, N2505);
or OR4 (N2524, N2511, N2274, N978, N1326);
or OR4 (N2525, N2518, N125, N1748, N1512);
nand NAND2 (N2526, N2523, N1608);
xor XOR2 (N2527, N2524, N164);
not NOT1 (N2528, N2525);
xor XOR2 (N2529, N2520, N322);
and AND4 (N2530, N2522, N2052, N2417, N1395);
buf BUF1 (N2531, N2529);
nand NAND2 (N2532, N2527, N2286);
nand NAND3 (N2533, N2528, N784, N581);
nand NAND4 (N2534, N2526, N2347, N193, N2163);
nor NOR3 (N2535, N2531, N1033, N723);
xor XOR2 (N2536, N2534, N666);
and AND3 (N2537, N2512, N1948, N1361);
nand NAND4 (N2538, N2516, N156, N2084, N974);
not NOT1 (N2539, N2535);
and AND4 (N2540, N2538, N1788, N324, N1810);
not NOT1 (N2541, N2533);
nor NOR4 (N2542, N2532, N1864, N392, N539);
not NOT1 (N2543, N2540);
and AND3 (N2544, N2530, N1821, N1424);
nand NAND4 (N2545, N2536, N1110, N66, N1276);
xor XOR2 (N2546, N2517, N10);
buf BUF1 (N2547, N2541);
nand NAND4 (N2548, N2546, N1342, N2235, N1802);
and AND2 (N2549, N2521, N2475);
xor XOR2 (N2550, N2519, N930);
and AND3 (N2551, N2549, N1125, N238);
or OR4 (N2552, N2539, N429, N1756, N363);
nand NAND3 (N2553, N2552, N123, N1528);
buf BUF1 (N2554, N2550);
xor XOR2 (N2555, N2545, N1565);
buf BUF1 (N2556, N2548);
or OR2 (N2557, N2554, N508);
and AND3 (N2558, N2557, N1203, N156);
nand NAND2 (N2559, N2553, N2528);
xor XOR2 (N2560, N2551, N629);
nand NAND4 (N2561, N2547, N2238, N153, N367);
nand NAND3 (N2562, N2542, N1635, N2199);
buf BUF1 (N2563, N2561);
nor NOR4 (N2564, N2544, N2232, N165, N2158);
or OR4 (N2565, N2559, N1940, N1359, N2095);
buf BUF1 (N2566, N2564);
nand NAND3 (N2567, N2537, N324, N1532);
or OR3 (N2568, N2566, N1853, N736);
xor XOR2 (N2569, N2567, N1411);
or OR3 (N2570, N2568, N2462, N243);
not NOT1 (N2571, N2555);
nand NAND4 (N2572, N2569, N2550, N1271, N924);
and AND3 (N2573, N2571, N2043, N662);
or OR4 (N2574, N2563, N938, N313, N386);
not NOT1 (N2575, N2556);
not NOT1 (N2576, N2562);
and AND2 (N2577, N2565, N1846);
and AND4 (N2578, N2574, N2485, N1705, N505);
and AND4 (N2579, N2572, N2050, N1833, N753);
and AND3 (N2580, N2570, N1540, N1818);
nor NOR3 (N2581, N2578, N175, N1451);
buf BUF1 (N2582, N2581);
and AND3 (N2583, N2573, N2526, N1970);
nor NOR4 (N2584, N2583, N995, N2347, N963);
not NOT1 (N2585, N2584);
buf BUF1 (N2586, N2585);
or OR4 (N2587, N2543, N715, N2082, N1461);
not NOT1 (N2588, N2579);
or OR4 (N2589, N2580, N1996, N1948, N370);
buf BUF1 (N2590, N2587);
buf BUF1 (N2591, N2576);
or OR2 (N2592, N2575, N1630);
not NOT1 (N2593, N2592);
nand NAND4 (N2594, N2589, N2350, N1336, N870);
and AND3 (N2595, N2582, N2057, N722);
and AND2 (N2596, N2595, N1876);
xor XOR2 (N2597, N2560, N1559);
nor NOR2 (N2598, N2577, N1925);
nand NAND2 (N2599, N2597, N1779);
or OR3 (N2600, N2590, N1347, N1955);
nor NOR3 (N2601, N2600, N523, N1719);
and AND3 (N2602, N2591, N2493, N1615);
and AND3 (N2603, N2602, N976, N704);
nand NAND4 (N2604, N2586, N396, N2129, N2471);
and AND3 (N2605, N2594, N1034, N611);
nand NAND4 (N2606, N2598, N1185, N2558, N1180);
nor NOR2 (N2607, N811, N136);
and AND3 (N2608, N2593, N2124, N1995);
and AND4 (N2609, N2599, N2210, N2172, N1451);
or OR4 (N2610, N2608, N652, N612, N2520);
xor XOR2 (N2611, N2601, N174);
nor NOR2 (N2612, N2603, N2431);
or OR3 (N2613, N2606, N2305, N68);
and AND3 (N2614, N2605, N913, N2012);
buf BUF1 (N2615, N2611);
and AND3 (N2616, N2607, N120, N2589);
nor NOR4 (N2617, N2604, N2468, N999, N2012);
not NOT1 (N2618, N2613);
buf BUF1 (N2619, N2618);
not NOT1 (N2620, N2615);
nand NAND3 (N2621, N2612, N1331, N426);
buf BUF1 (N2622, N2596);
or OR4 (N2623, N2614, N273, N1494, N632);
buf BUF1 (N2624, N2621);
buf BUF1 (N2625, N2622);
nor NOR3 (N2626, N2610, N2536, N221);
nor NOR3 (N2627, N2626, N54, N653);
nand NAND2 (N2628, N2619, N234);
buf BUF1 (N2629, N2624);
not NOT1 (N2630, N2588);
buf BUF1 (N2631, N2628);
not NOT1 (N2632, N2625);
and AND2 (N2633, N2631, N1461);
nor NOR3 (N2634, N2620, N2230, N578);
or OR3 (N2635, N2630, N869, N2425);
not NOT1 (N2636, N2627);
not NOT1 (N2637, N2623);
or OR3 (N2638, N2629, N998, N2595);
nor NOR2 (N2639, N2638, N2051);
nand NAND2 (N2640, N2639, N2406);
and AND4 (N2641, N2637, N576, N880, N1979);
or OR2 (N2642, N2617, N2038);
buf BUF1 (N2643, N2634);
nand NAND4 (N2644, N2616, N1239, N2066, N391);
not NOT1 (N2645, N2640);
xor XOR2 (N2646, N2644, N1689);
or OR2 (N2647, N2636, N1893);
buf BUF1 (N2648, N2641);
xor XOR2 (N2649, N2645, N988);
or OR3 (N2650, N2646, N2299, N607);
and AND4 (N2651, N2609, N1708, N209, N1011);
nor NOR2 (N2652, N2635, N62);
and AND2 (N2653, N2642, N2526);
nor NOR3 (N2654, N2633, N976, N527);
xor XOR2 (N2655, N2651, N1689);
not NOT1 (N2656, N2649);
nor NOR3 (N2657, N2653, N1578, N306);
and AND2 (N2658, N2654, N95);
buf BUF1 (N2659, N2652);
buf BUF1 (N2660, N2659);
buf BUF1 (N2661, N2650);
nand NAND4 (N2662, N2632, N2535, N1940, N1626);
or OR3 (N2663, N2647, N1946, N258);
or OR4 (N2664, N2656, N1116, N175, N1448);
nor NOR3 (N2665, N2643, N1156, N1629);
nand NAND3 (N2666, N2657, N1539, N2288);
not NOT1 (N2667, N2660);
nand NAND2 (N2668, N2664, N2414);
xor XOR2 (N2669, N2655, N505);
nand NAND4 (N2670, N2668, N1555, N1230, N2419);
or OR4 (N2671, N2666, N322, N99, N1385);
or OR4 (N2672, N2648, N1712, N819, N972);
buf BUF1 (N2673, N2671);
nand NAND3 (N2674, N2672, N2158, N1971);
not NOT1 (N2675, N2667);
nand NAND2 (N2676, N2675, N2347);
nor NOR4 (N2677, N2658, N289, N1039, N824);
nand NAND2 (N2678, N2661, N278);
buf BUF1 (N2679, N2669);
nand NAND3 (N2680, N2670, N2613, N782);
buf BUF1 (N2681, N2676);
and AND2 (N2682, N2663, N1968);
nor NOR3 (N2683, N2681, N2055, N2304);
nand NAND3 (N2684, N2678, N1847, N1732);
buf BUF1 (N2685, N2673);
nand NAND3 (N2686, N2665, N2040, N2496);
or OR2 (N2687, N2684, N2507);
not NOT1 (N2688, N2683);
and AND4 (N2689, N2686, N2661, N2254, N630);
buf BUF1 (N2690, N2680);
not NOT1 (N2691, N2687);
nand NAND4 (N2692, N2674, N2243, N2308, N1965);
nand NAND4 (N2693, N2691, N517, N1480, N1915);
xor XOR2 (N2694, N2688, N1399);
xor XOR2 (N2695, N2693, N1389);
or OR4 (N2696, N2695, N794, N583, N2317);
nor NOR3 (N2697, N2696, N35, N1142);
not NOT1 (N2698, N2694);
xor XOR2 (N2699, N2697, N1470);
not NOT1 (N2700, N2692);
nor NOR2 (N2701, N2679, N1674);
buf BUF1 (N2702, N2689);
not NOT1 (N2703, N2662);
or OR3 (N2704, N2700, N1298, N304);
nor NOR4 (N2705, N2685, N1929, N2245, N1116);
xor XOR2 (N2706, N2704, N2658);
and AND4 (N2707, N2690, N2621, N995, N408);
or OR3 (N2708, N2698, N1880, N900);
nor NOR3 (N2709, N2707, N56, N1527);
or OR2 (N2710, N2702, N230);
xor XOR2 (N2711, N2710, N1332);
or OR2 (N2712, N2701, N308);
xor XOR2 (N2713, N2708, N856);
and AND2 (N2714, N2699, N1220);
nor NOR2 (N2715, N2677, N597);
not NOT1 (N2716, N2706);
buf BUF1 (N2717, N2715);
nor NOR4 (N2718, N2716, N2396, N127, N985);
not NOT1 (N2719, N2712);
nand NAND3 (N2720, N2718, N1689, N810);
buf BUF1 (N2721, N2709);
nor NOR3 (N2722, N2682, N54, N2419);
and AND4 (N2723, N2703, N932, N1147, N2001);
nand NAND2 (N2724, N2721, N2517);
xor XOR2 (N2725, N2720, N2046);
not NOT1 (N2726, N2724);
nor NOR3 (N2727, N2711, N415, N163);
or OR3 (N2728, N2727, N347, N1349);
buf BUF1 (N2729, N2717);
buf BUF1 (N2730, N2722);
buf BUF1 (N2731, N2714);
buf BUF1 (N2732, N2730);
or OR3 (N2733, N2729, N2140, N238);
nor NOR3 (N2734, N2731, N1421, N1804);
or OR3 (N2735, N2719, N2621, N271);
not NOT1 (N2736, N2705);
nor NOR3 (N2737, N2728, N939, N2055);
nand NAND3 (N2738, N2725, N2380, N2035);
nor NOR3 (N2739, N2735, N1559, N1114);
or OR2 (N2740, N2734, N1167);
not NOT1 (N2741, N2740);
xor XOR2 (N2742, N2736, N2183);
nor NOR2 (N2743, N2742, N1905);
nor NOR4 (N2744, N2741, N336, N2340, N901);
xor XOR2 (N2745, N2743, N2273);
buf BUF1 (N2746, N2745);
not NOT1 (N2747, N2732);
nand NAND3 (N2748, N2746, N165, N455);
nand NAND4 (N2749, N2747, N1238, N718, N60);
and AND3 (N2750, N2739, N765, N526);
nand NAND2 (N2751, N2737, N2173);
xor XOR2 (N2752, N2738, N534);
and AND3 (N2753, N2726, N2629, N1103);
nor NOR2 (N2754, N2752, N442);
and AND3 (N2755, N2713, N1754, N1836);
nor NOR3 (N2756, N2748, N1731, N1238);
not NOT1 (N2757, N2733);
nor NOR2 (N2758, N2757, N345);
nand NAND4 (N2759, N2723, N2160, N624, N1114);
nor NOR3 (N2760, N2749, N2640, N2263);
xor XOR2 (N2761, N2758, N26);
not NOT1 (N2762, N2761);
buf BUF1 (N2763, N2759);
buf BUF1 (N2764, N2751);
or OR4 (N2765, N2756, N1601, N1873, N511);
nand NAND3 (N2766, N2755, N2414, N1447);
xor XOR2 (N2767, N2760, N257);
not NOT1 (N2768, N2744);
nor NOR2 (N2769, N2753, N112);
or OR2 (N2770, N2762, N1269);
and AND2 (N2771, N2768, N36);
or OR3 (N2772, N2754, N1839, N2075);
or OR2 (N2773, N2770, N2301);
buf BUF1 (N2774, N2769);
and AND3 (N2775, N2774, N1925, N1335);
buf BUF1 (N2776, N2775);
nor NOR3 (N2777, N2776, N530, N2161);
not NOT1 (N2778, N2765);
nand NAND4 (N2779, N2773, N662, N73, N1529);
buf BUF1 (N2780, N2764);
nand NAND4 (N2781, N2780, N1633, N730, N348);
or OR2 (N2782, N2781, N1763);
not NOT1 (N2783, N2766);
or OR4 (N2784, N2777, N1613, N731, N1305);
xor XOR2 (N2785, N2772, N2499);
xor XOR2 (N2786, N2785, N1436);
nand NAND4 (N2787, N2783, N476, N1924, N424);
not NOT1 (N2788, N2782);
and AND3 (N2789, N2767, N1200, N1683);
not NOT1 (N2790, N2779);
not NOT1 (N2791, N2771);
and AND3 (N2792, N2750, N2419, N457);
and AND3 (N2793, N2789, N2674, N1705);
nor NOR2 (N2794, N2786, N1227);
not NOT1 (N2795, N2788);
nor NOR3 (N2796, N2763, N1006, N696);
nor NOR3 (N2797, N2796, N294, N2092);
and AND3 (N2798, N2790, N825, N368);
nor NOR3 (N2799, N2787, N1265, N952);
xor XOR2 (N2800, N2792, N2512);
and AND2 (N2801, N2784, N1804);
and AND4 (N2802, N2797, N2736, N880, N643);
xor XOR2 (N2803, N2802, N2034);
nand NAND2 (N2804, N2798, N224);
nor NOR4 (N2805, N2803, N2072, N91, N1055);
and AND4 (N2806, N2778, N722, N1191, N1919);
and AND2 (N2807, N2794, N2427);
nor NOR2 (N2808, N2791, N430);
xor XOR2 (N2809, N2800, N717);
xor XOR2 (N2810, N2804, N2329);
and AND2 (N2811, N2805, N1983);
nor NOR4 (N2812, N2801, N2632, N717, N1421);
nand NAND4 (N2813, N2807, N1698, N1100, N1095);
not NOT1 (N2814, N2806);
xor XOR2 (N2815, N2799, N1015);
nand NAND2 (N2816, N2795, N423);
buf BUF1 (N2817, N2808);
not NOT1 (N2818, N2814);
and AND3 (N2819, N2811, N111, N1562);
nand NAND4 (N2820, N2809, N843, N651, N2425);
or OR4 (N2821, N2810, N2775, N1462, N444);
nand NAND2 (N2822, N2816, N2100);
and AND2 (N2823, N2821, N1136);
and AND4 (N2824, N2813, N805, N1521, N227);
and AND4 (N2825, N2820, N568, N1576, N2335);
or OR3 (N2826, N2815, N2163, N1590);
and AND4 (N2827, N2823, N2320, N2612, N663);
not NOT1 (N2828, N2822);
not NOT1 (N2829, N2817);
or OR4 (N2830, N2827, N2692, N2312, N2583);
nor NOR2 (N2831, N2830, N1927);
nor NOR2 (N2832, N2824, N333);
buf BUF1 (N2833, N2818);
nand NAND3 (N2834, N2828, N1774, N309);
not NOT1 (N2835, N2832);
nand NAND2 (N2836, N2826, N265);
nand NAND4 (N2837, N2833, N2307, N2744, N376);
xor XOR2 (N2838, N2837, N1867);
and AND3 (N2839, N2835, N332, N1814);
buf BUF1 (N2840, N2793);
nor NOR4 (N2841, N2812, N319, N2558, N1685);
buf BUF1 (N2842, N2829);
not NOT1 (N2843, N2831);
buf BUF1 (N2844, N2838);
nor NOR4 (N2845, N2843, N1359, N2201, N1875);
or OR2 (N2846, N2845, N2570);
and AND4 (N2847, N2839, N875, N475, N869);
buf BUF1 (N2848, N2847);
or OR2 (N2849, N2840, N2752);
xor XOR2 (N2850, N2846, N1894);
nand NAND2 (N2851, N2841, N2810);
buf BUF1 (N2852, N2819);
or OR3 (N2853, N2844, N982, N2781);
buf BUF1 (N2854, N2849);
xor XOR2 (N2855, N2834, N2451);
or OR3 (N2856, N2850, N1669, N1861);
nor NOR2 (N2857, N2851, N2274);
or OR2 (N2858, N2836, N2014);
or OR4 (N2859, N2848, N140, N425, N2302);
nor NOR2 (N2860, N2852, N966);
nor NOR3 (N2861, N2860, N22, N1313);
nor NOR2 (N2862, N2859, N314);
buf BUF1 (N2863, N2857);
buf BUF1 (N2864, N2825);
buf BUF1 (N2865, N2855);
not NOT1 (N2866, N2861);
not NOT1 (N2867, N2854);
and AND3 (N2868, N2865, N923, N2243);
or OR3 (N2869, N2864, N1507, N2042);
buf BUF1 (N2870, N2856);
nor NOR4 (N2871, N2870, N663, N2096, N1461);
buf BUF1 (N2872, N2842);
xor XOR2 (N2873, N2871, N695);
xor XOR2 (N2874, N2872, N629);
not NOT1 (N2875, N2853);
and AND4 (N2876, N2866, N1855, N2381, N897);
nand NAND3 (N2877, N2876, N1610, N1543);
or OR4 (N2878, N2875, N2513, N980, N1957);
not NOT1 (N2879, N2874);
nor NOR3 (N2880, N2868, N96, N1191);
and AND2 (N2881, N2867, N1656);
nand NAND2 (N2882, N2881, N442);
xor XOR2 (N2883, N2877, N1477);
nand NAND4 (N2884, N2858, N1577, N350, N683);
not NOT1 (N2885, N2869);
not NOT1 (N2886, N2863);
buf BUF1 (N2887, N2880);
and AND3 (N2888, N2862, N680, N1399);
or OR3 (N2889, N2885, N709, N240);
and AND3 (N2890, N2889, N2809, N444);
nor NOR3 (N2891, N2873, N1575, N1298);
nor NOR3 (N2892, N2884, N2170, N2664);
not NOT1 (N2893, N2883);
nor NOR3 (N2894, N2879, N815, N1598);
not NOT1 (N2895, N2894);
nor NOR3 (N2896, N2887, N2579, N88);
nand NAND3 (N2897, N2888, N238, N957);
or OR2 (N2898, N2895, N1320);
nand NAND3 (N2899, N2897, N2422, N164);
nand NAND3 (N2900, N2882, N2824, N1310);
xor XOR2 (N2901, N2878, N2125);
xor XOR2 (N2902, N2899, N2881);
nor NOR4 (N2903, N2891, N1166, N732, N284);
buf BUF1 (N2904, N2886);
nor NOR2 (N2905, N2902, N1823);
not NOT1 (N2906, N2904);
not NOT1 (N2907, N2898);
nor NOR3 (N2908, N2893, N819, N2345);
nor NOR3 (N2909, N2896, N2812, N711);
buf BUF1 (N2910, N2905);
not NOT1 (N2911, N2892);
not NOT1 (N2912, N2890);
or OR2 (N2913, N2910, N577);
or OR4 (N2914, N2900, N411, N2551, N840);
not NOT1 (N2915, N2901);
buf BUF1 (N2916, N2907);
not NOT1 (N2917, N2911);
buf BUF1 (N2918, N2912);
not NOT1 (N2919, N2909);
buf BUF1 (N2920, N2908);
xor XOR2 (N2921, N2920, N2196);
and AND3 (N2922, N2914, N165, N1182);
or OR4 (N2923, N2906, N1889, N28, N2309);
xor XOR2 (N2924, N2916, N1123);
buf BUF1 (N2925, N2923);
not NOT1 (N2926, N2924);
nor NOR3 (N2927, N2922, N1214, N1039);
nand NAND2 (N2928, N2927, N1708);
nor NOR4 (N2929, N2917, N1366, N1593, N1442);
nand NAND4 (N2930, N2929, N1442, N2365, N91);
buf BUF1 (N2931, N2921);
buf BUF1 (N2932, N2915);
nand NAND3 (N2933, N2930, N1497, N142);
buf BUF1 (N2934, N2925);
or OR4 (N2935, N2903, N2301, N1990, N2308);
buf BUF1 (N2936, N2931);
nor NOR2 (N2937, N2933, N893);
nand NAND3 (N2938, N2928, N881, N1259);
buf BUF1 (N2939, N2926);
and AND3 (N2940, N2935, N1218, N2020);
or OR3 (N2941, N2913, N114, N2820);
nand NAND2 (N2942, N2934, N2626);
buf BUF1 (N2943, N2941);
buf BUF1 (N2944, N2937);
or OR3 (N2945, N2940, N193, N2319);
and AND3 (N2946, N2918, N404, N1587);
xor XOR2 (N2947, N2945, N519);
nand NAND2 (N2948, N2919, N245);
nand NAND4 (N2949, N2936, N1693, N2310, N2551);
and AND3 (N2950, N2946, N1750, N503);
nor NOR2 (N2951, N2950, N490);
not NOT1 (N2952, N2948);
not NOT1 (N2953, N2938);
and AND2 (N2954, N2944, N294);
nand NAND3 (N2955, N2943, N680, N2064);
and AND3 (N2956, N2947, N1176, N873);
not NOT1 (N2957, N2951);
nand NAND3 (N2958, N2957, N286, N230);
or OR3 (N2959, N2942, N2095, N1177);
nor NOR3 (N2960, N2932, N1357, N29);
nor NOR2 (N2961, N2952, N108);
not NOT1 (N2962, N2955);
not NOT1 (N2963, N2939);
buf BUF1 (N2964, N2960);
nor NOR4 (N2965, N2964, N1315, N2301, N2538);
buf BUF1 (N2966, N2963);
or OR2 (N2967, N2962, N1734);
and AND4 (N2968, N2961, N2492, N505, N314);
buf BUF1 (N2969, N2965);
not NOT1 (N2970, N2954);
not NOT1 (N2971, N2949);
and AND4 (N2972, N2968, N1265, N2814, N2292);
not NOT1 (N2973, N2970);
and AND4 (N2974, N2966, N754, N1324, N2396);
buf BUF1 (N2975, N2969);
nand NAND3 (N2976, N2956, N450, N530);
and AND2 (N2977, N2975, N858);
nand NAND2 (N2978, N2973, N1995);
buf BUF1 (N2979, N2977);
xor XOR2 (N2980, N2974, N1606);
and AND4 (N2981, N2959, N338, N338, N214);
nand NAND3 (N2982, N2978, N510, N2093);
and AND3 (N2983, N2981, N2008, N1626);
buf BUF1 (N2984, N2976);
nor NOR2 (N2985, N2984, N2894);
and AND2 (N2986, N2953, N2522);
buf BUF1 (N2987, N2958);
nand NAND4 (N2988, N2980, N2740, N2620, N2429);
or OR4 (N2989, N2983, N55, N1842, N2294);
buf BUF1 (N2990, N2971);
buf BUF1 (N2991, N2967);
xor XOR2 (N2992, N2990, N175);
not NOT1 (N2993, N2982);
buf BUF1 (N2994, N2972);
nor NOR3 (N2995, N2987, N1264, N2057);
or OR4 (N2996, N2988, N1695, N103, N914);
xor XOR2 (N2997, N2979, N892);
and AND2 (N2998, N2997, N2128);
and AND3 (N2999, N2991, N705, N2606);
buf BUF1 (N3000, N2996);
nand NAND4 (N3001, N2986, N2439, N2668, N945);
or OR3 (N3002, N2985, N1347, N901);
nand NAND2 (N3003, N2999, N2970);
and AND4 (N3004, N2998, N1921, N1446, N1808);
not NOT1 (N3005, N2994);
nor NOR3 (N3006, N3000, N1962, N537);
xor XOR2 (N3007, N3002, N515);
or OR3 (N3008, N3006, N705, N1456);
nand NAND4 (N3009, N3003, N2985, N2823, N2833);
nand NAND4 (N3010, N3005, N2820, N1318, N2204);
or OR2 (N3011, N3010, N1897);
and AND4 (N3012, N2993, N2539, N1152, N1502);
nor NOR3 (N3013, N3009, N815, N652);
nand NAND3 (N3014, N3004, N2336, N2726);
nand NAND4 (N3015, N3007, N2005, N985, N1833);
or OR4 (N3016, N3008, N948, N1076, N946);
nand NAND4 (N3017, N2995, N162, N2620, N39);
nand NAND4 (N3018, N3012, N389, N2768, N131);
not NOT1 (N3019, N3014);
buf BUF1 (N3020, N3015);
and AND4 (N3021, N3013, N548, N2844, N1546);
nor NOR4 (N3022, N2989, N2360, N209, N1724);
not NOT1 (N3023, N3001);
not NOT1 (N3024, N3016);
nand NAND2 (N3025, N3019, N76);
buf BUF1 (N3026, N3018);
nor NOR4 (N3027, N3020, N2969, N2734, N2223);
or OR3 (N3028, N2992, N377, N1739);
and AND4 (N3029, N3024, N145, N1429, N2626);
buf BUF1 (N3030, N3025);
or OR3 (N3031, N3011, N1228, N675);
and AND2 (N3032, N3022, N2605);
nand NAND2 (N3033, N3030, N1952);
xor XOR2 (N3034, N3033, N2214);
not NOT1 (N3035, N3027);
not NOT1 (N3036, N3028);
nor NOR2 (N3037, N3026, N1293);
buf BUF1 (N3038, N3035);
nand NAND2 (N3039, N3029, N2977);
nor NOR4 (N3040, N3034, N1120, N1224, N289);
nor NOR2 (N3041, N3037, N2337);
or OR4 (N3042, N3038, N1737, N1763, N467);
not NOT1 (N3043, N3031);
nand NAND3 (N3044, N3021, N1681, N1237);
nand NAND2 (N3045, N3040, N1619);
buf BUF1 (N3046, N3023);
not NOT1 (N3047, N3044);
nand NAND3 (N3048, N3046, N767, N2761);
and AND2 (N3049, N3045, N1612);
nand NAND4 (N3050, N3039, N1199, N1374, N1051);
xor XOR2 (N3051, N3050, N2023);
nand NAND4 (N3052, N3049, N2967, N961, N844);
xor XOR2 (N3053, N3042, N2406);
and AND4 (N3054, N3036, N1260, N2515, N64);
or OR4 (N3055, N3047, N647, N1210, N1600);
xor XOR2 (N3056, N3055, N2306);
nand NAND4 (N3057, N3051, N2840, N675, N1756);
not NOT1 (N3058, N3032);
nor NOR3 (N3059, N3052, N1429, N1618);
and AND2 (N3060, N3054, N1780);
nor NOR3 (N3061, N3053, N1081, N1760);
not NOT1 (N3062, N3017);
and AND2 (N3063, N3060, N2185);
xor XOR2 (N3064, N3061, N2080);
not NOT1 (N3065, N3041);
xor XOR2 (N3066, N3048, N1037);
xor XOR2 (N3067, N3066, N1439);
not NOT1 (N3068, N3043);
nand NAND4 (N3069, N3063, N340, N2992, N1712);
not NOT1 (N3070, N3062);
nor NOR2 (N3071, N3064, N285);
or OR2 (N3072, N3071, N2210);
nor NOR3 (N3073, N3056, N5, N470);
and AND4 (N3074, N3067, N346, N1405, N295);
or OR3 (N3075, N3059, N1576, N1752);
or OR2 (N3076, N3073, N2486);
nor NOR4 (N3077, N3074, N638, N2627, N2245);
nand NAND2 (N3078, N3058, N1488);
xor XOR2 (N3079, N3068, N505);
not NOT1 (N3080, N3072);
nor NOR2 (N3081, N3070, N1211);
and AND3 (N3082, N3080, N3005, N2950);
or OR4 (N3083, N3082, N2714, N2552, N2690);
not NOT1 (N3084, N3078);
nor NOR2 (N3085, N3077, N1195);
nor NOR2 (N3086, N3084, N2514);
and AND4 (N3087, N3076, N1743, N2127, N1019);
nor NOR4 (N3088, N3079, N1965, N1941, N1009);
not NOT1 (N3089, N3057);
nand NAND4 (N3090, N3081, N2317, N433, N472);
nand NAND4 (N3091, N3088, N1338, N795, N1174);
or OR2 (N3092, N3065, N2563);
not NOT1 (N3093, N3075);
buf BUF1 (N3094, N3092);
or OR4 (N3095, N3089, N1981, N269, N1958);
xor XOR2 (N3096, N3094, N647);
and AND4 (N3097, N3085, N610, N1757, N1466);
xor XOR2 (N3098, N3069, N3027);
nand NAND3 (N3099, N3097, N1065, N94);
xor XOR2 (N3100, N3098, N2232);
xor XOR2 (N3101, N3091, N330);
xor XOR2 (N3102, N3100, N2837);
or OR4 (N3103, N3093, N1528, N1326, N688);
buf BUF1 (N3104, N3101);
buf BUF1 (N3105, N3090);
not NOT1 (N3106, N3103);
and AND2 (N3107, N3087, N1673);
not NOT1 (N3108, N3096);
buf BUF1 (N3109, N3083);
and AND3 (N3110, N3108, N1733, N2972);
buf BUF1 (N3111, N3099);
xor XOR2 (N3112, N3111, N2360);
buf BUF1 (N3113, N3095);
nor NOR3 (N3114, N3107, N2271, N1690);
buf BUF1 (N3115, N3110);
nand NAND3 (N3116, N3112, N2676, N2248);
buf BUF1 (N3117, N3113);
and AND3 (N3118, N3115, N1636, N688);
xor XOR2 (N3119, N3104, N3039);
xor XOR2 (N3120, N3117, N3100);
nor NOR3 (N3121, N3086, N378, N45);
nand NAND4 (N3122, N3109, N375, N2852, N2412);
nor NOR4 (N3123, N3119, N1101, N1969, N2985);
buf BUF1 (N3124, N3123);
or OR2 (N3125, N3118, N3016);
not NOT1 (N3126, N3105);
buf BUF1 (N3127, N3126);
and AND3 (N3128, N3125, N51, N1768);
xor XOR2 (N3129, N3106, N671);
buf BUF1 (N3130, N3124);
not NOT1 (N3131, N3120);
buf BUF1 (N3132, N3127);
not NOT1 (N3133, N3130);
nor NOR4 (N3134, N3116, N2434, N2716, N1747);
xor XOR2 (N3135, N3133, N1290);
or OR4 (N3136, N3134, N282, N378, N1411);
nor NOR3 (N3137, N3114, N1974, N3059);
and AND4 (N3138, N3102, N2164, N2714, N153);
nor NOR4 (N3139, N3121, N158, N89, N1448);
buf BUF1 (N3140, N3128);
not NOT1 (N3141, N3131);
nand NAND4 (N3142, N3141, N1206, N2621, N1877);
nor NOR4 (N3143, N3122, N2801, N2283, N3036);
nand NAND4 (N3144, N3139, N1655, N25, N2912);
or OR3 (N3145, N3142, N119, N512);
not NOT1 (N3146, N3129);
buf BUF1 (N3147, N3132);
and AND3 (N3148, N3137, N2280, N1070);
not NOT1 (N3149, N3146);
or OR2 (N3150, N3149, N807);
xor XOR2 (N3151, N3144, N2790);
and AND3 (N3152, N3135, N2447, N113);
nand NAND2 (N3153, N3151, N603);
nor NOR3 (N3154, N3153, N2056, N2544);
xor XOR2 (N3155, N3150, N2359);
xor XOR2 (N3156, N3147, N1743);
nand NAND4 (N3157, N3143, N1525, N1989, N2382);
nor NOR3 (N3158, N3138, N2421, N1491);
xor XOR2 (N3159, N3158, N2817);
and AND2 (N3160, N3148, N1902);
and AND3 (N3161, N3159, N1421, N2959);
and AND4 (N3162, N3160, N2201, N2983, N919);
or OR4 (N3163, N3154, N45, N1628, N3027);
or OR3 (N3164, N3161, N2093, N941);
buf BUF1 (N3165, N3136);
and AND3 (N3166, N3155, N499, N1372);
nand NAND4 (N3167, N3140, N2355, N2342, N376);
or OR2 (N3168, N3165, N227);
not NOT1 (N3169, N3156);
nor NOR4 (N3170, N3145, N2595, N964, N2712);
not NOT1 (N3171, N3166);
nor NOR3 (N3172, N3170, N3158, N2001);
not NOT1 (N3173, N3169);
nand NAND4 (N3174, N3172, N784, N848, N1795);
not NOT1 (N3175, N3168);
xor XOR2 (N3176, N3174, N2606);
not NOT1 (N3177, N3171);
nand NAND4 (N3178, N3173, N543, N442, N244);
and AND4 (N3179, N3162, N2522, N1269, N3067);
and AND3 (N3180, N3152, N248, N2057);
nand NAND2 (N3181, N3177, N633);
buf BUF1 (N3182, N3175);
nor NOR3 (N3183, N3178, N1922, N705);
nand NAND2 (N3184, N3180, N798);
buf BUF1 (N3185, N3163);
nor NOR2 (N3186, N3164, N389);
xor XOR2 (N3187, N3184, N678);
nor NOR2 (N3188, N3187, N979);
nor NOR3 (N3189, N3176, N232, N3059);
and AND2 (N3190, N3181, N989);
nor NOR4 (N3191, N3183, N147, N2948, N2611);
nand NAND2 (N3192, N3191, N2578);
or OR4 (N3193, N3186, N3039, N2299, N1306);
and AND3 (N3194, N3189, N2303, N2478);
xor XOR2 (N3195, N3190, N2970);
buf BUF1 (N3196, N3194);
nand NAND3 (N3197, N3179, N2839, N163);
not NOT1 (N3198, N3182);
nand NAND2 (N3199, N3192, N1525);
xor XOR2 (N3200, N3198, N1931);
nand NAND3 (N3201, N3200, N661, N46);
nand NAND3 (N3202, N3188, N1109, N2130);
not NOT1 (N3203, N3185);
xor XOR2 (N3204, N3157, N2066);
and AND3 (N3205, N3196, N2162, N1929);
or OR4 (N3206, N3195, N3063, N2158, N994);
nand NAND3 (N3207, N3197, N3068, N1319);
nand NAND2 (N3208, N3202, N568);
buf BUF1 (N3209, N3204);
not NOT1 (N3210, N3209);
xor XOR2 (N3211, N3193, N2802);
nand NAND4 (N3212, N3201, N997, N836, N1963);
nor NOR4 (N3213, N3205, N749, N3101, N2786);
buf BUF1 (N3214, N3210);
and AND2 (N3215, N3208, N297);
and AND3 (N3216, N3212, N1798, N2288);
nor NOR3 (N3217, N3207, N2050, N2935);
buf BUF1 (N3218, N3214);
buf BUF1 (N3219, N3206);
buf BUF1 (N3220, N3199);
nand NAND3 (N3221, N3218, N1220, N1385);
buf BUF1 (N3222, N3216);
and AND4 (N3223, N3203, N2586, N2139, N979);
buf BUF1 (N3224, N3222);
xor XOR2 (N3225, N3213, N1541);
xor XOR2 (N3226, N3221, N1779);
nor NOR4 (N3227, N3219, N2081, N2668, N240);
nand NAND4 (N3228, N3224, N1700, N2434, N1146);
not NOT1 (N3229, N3167);
not NOT1 (N3230, N3211);
xor XOR2 (N3231, N3225, N2546);
buf BUF1 (N3232, N3228);
nor NOR2 (N3233, N3217, N3166);
nand NAND4 (N3234, N3226, N1853, N654, N1833);
xor XOR2 (N3235, N3229, N2451);
not NOT1 (N3236, N3230);
nor NOR4 (N3237, N3231, N2925, N1603, N661);
or OR3 (N3238, N3234, N1193, N2473);
not NOT1 (N3239, N3220);
nand NAND2 (N3240, N3236, N213);
or OR2 (N3241, N3227, N2233);
or OR2 (N3242, N3237, N1476);
not NOT1 (N3243, N3241);
and AND3 (N3244, N3235, N566, N1883);
nor NOR4 (N3245, N3244, N2054, N1957, N1599);
nor NOR3 (N3246, N3223, N1399, N1682);
buf BUF1 (N3247, N3246);
buf BUF1 (N3248, N3233);
or OR4 (N3249, N3245, N524, N2608, N2304);
nor NOR4 (N3250, N3249, N479, N978, N859);
not NOT1 (N3251, N3247);
not NOT1 (N3252, N3215);
xor XOR2 (N3253, N3250, N1592);
and AND3 (N3254, N3252, N255, N2083);
not NOT1 (N3255, N3232);
xor XOR2 (N3256, N3238, N1503);
or OR4 (N3257, N3256, N300, N141, N2581);
nor NOR2 (N3258, N3248, N2177);
not NOT1 (N3259, N3251);
and AND2 (N3260, N3240, N2711);
or OR4 (N3261, N3254, N1908, N3110, N895);
or OR2 (N3262, N3259, N2388);
and AND4 (N3263, N3260, N1116, N1848, N1063);
nand NAND4 (N3264, N3262, N517, N3211, N2041);
xor XOR2 (N3265, N3257, N1392);
or OR3 (N3266, N3264, N984, N1963);
buf BUF1 (N3267, N3242);
buf BUF1 (N3268, N3267);
xor XOR2 (N3269, N3268, N906);
not NOT1 (N3270, N3266);
xor XOR2 (N3271, N3239, N2093);
or OR4 (N3272, N3258, N2168, N2954, N566);
and AND2 (N3273, N3243, N944);
nor NOR3 (N3274, N3261, N842, N1575);
and AND4 (N3275, N3269, N2133, N1874, N1322);
buf BUF1 (N3276, N3271);
nand NAND3 (N3277, N3270, N1784, N1542);
nand NAND4 (N3278, N3263, N75, N1504, N802);
buf BUF1 (N3279, N3255);
buf BUF1 (N3280, N3276);
and AND2 (N3281, N3280, N710);
nor NOR3 (N3282, N3275, N3266, N721);
nor NOR2 (N3283, N3265, N3032);
not NOT1 (N3284, N3282);
buf BUF1 (N3285, N3281);
or OR3 (N3286, N3253, N900, N967);
not NOT1 (N3287, N3277);
nand NAND3 (N3288, N3283, N599, N1613);
not NOT1 (N3289, N3279);
buf BUF1 (N3290, N3287);
buf BUF1 (N3291, N3290);
buf BUF1 (N3292, N3278);
nand NAND4 (N3293, N3272, N2447, N827, N377);
or OR4 (N3294, N3274, N2525, N1327, N2718);
not NOT1 (N3295, N3288);
buf BUF1 (N3296, N3284);
or OR3 (N3297, N3285, N2476, N801);
and AND3 (N3298, N3289, N800, N1884);
or OR3 (N3299, N3293, N379, N770);
xor XOR2 (N3300, N3298, N900);
and AND4 (N3301, N3294, N1701, N3084, N513);
buf BUF1 (N3302, N3273);
not NOT1 (N3303, N3286);
not NOT1 (N3304, N3302);
or OR4 (N3305, N3301, N151, N2453, N1709);
buf BUF1 (N3306, N3297);
buf BUF1 (N3307, N3295);
or OR4 (N3308, N3300, N712, N2894, N903);
buf BUF1 (N3309, N3299);
nand NAND2 (N3310, N3306, N1409);
and AND4 (N3311, N3291, N699, N1369, N2448);
not NOT1 (N3312, N3307);
not NOT1 (N3313, N3296);
or OR4 (N3314, N3292, N1637, N1677, N2853);
xor XOR2 (N3315, N3310, N1711);
or OR4 (N3316, N3304, N2753, N1265, N2900);
nand NAND3 (N3317, N3303, N2413, N1230);
buf BUF1 (N3318, N3316);
and AND4 (N3319, N3317, N1566, N1502, N2562);
nor NOR3 (N3320, N3313, N2017, N1754);
not NOT1 (N3321, N3320);
nor NOR4 (N3322, N3321, N2254, N2613, N1213);
nand NAND3 (N3323, N3318, N514, N48);
nor NOR4 (N3324, N3319, N3110, N3292, N359);
and AND2 (N3325, N3312, N1298);
not NOT1 (N3326, N3315);
or OR2 (N3327, N3326, N3176);
nor NOR2 (N3328, N3322, N721);
xor XOR2 (N3329, N3305, N714);
not NOT1 (N3330, N3328);
and AND4 (N3331, N3327, N3270, N232, N3316);
nor NOR3 (N3332, N3329, N339, N2100);
buf BUF1 (N3333, N3324);
not NOT1 (N3334, N3333);
xor XOR2 (N3335, N3308, N55);
not NOT1 (N3336, N3334);
buf BUF1 (N3337, N3335);
nor NOR4 (N3338, N3309, N3103, N3091, N415);
or OR4 (N3339, N3323, N285, N1710, N1751);
nand NAND3 (N3340, N3332, N2997, N3004);
xor XOR2 (N3341, N3311, N2458);
buf BUF1 (N3342, N3336);
not NOT1 (N3343, N3340);
nand NAND2 (N3344, N3314, N1692);
buf BUF1 (N3345, N3341);
nor NOR2 (N3346, N3344, N36);
or OR4 (N3347, N3338, N1364, N3023, N3074);
nand NAND4 (N3348, N3343, N1443, N610, N845);
nor NOR2 (N3349, N3331, N568);
and AND2 (N3350, N3349, N274);
nand NAND4 (N3351, N3347, N797, N2217, N2176);
buf BUF1 (N3352, N3346);
and AND3 (N3353, N3342, N225, N1774);
nor NOR3 (N3354, N3353, N77, N2826);
nor NOR2 (N3355, N3351, N728);
nand NAND3 (N3356, N3350, N1237, N2175);
and AND4 (N3357, N3330, N105, N3119, N2394);
or OR2 (N3358, N3354, N2938);
nand NAND4 (N3359, N3357, N3047, N1279, N2493);
nor NOR3 (N3360, N3339, N1709, N328);
nor NOR3 (N3361, N3356, N3030, N2732);
or OR4 (N3362, N3358, N764, N3154, N551);
buf BUF1 (N3363, N3361);
buf BUF1 (N3364, N3325);
and AND2 (N3365, N3363, N1991);
xor XOR2 (N3366, N3364, N873);
not NOT1 (N3367, N3345);
or OR4 (N3368, N3348, N763, N1190, N1451);
buf BUF1 (N3369, N3360);
or OR2 (N3370, N3355, N3215);
not NOT1 (N3371, N3367);
or OR3 (N3372, N3362, N1109, N1811);
nor NOR3 (N3373, N3366, N503, N3239);
nand NAND3 (N3374, N3373, N1829, N2710);
and AND3 (N3375, N3337, N651, N192);
not NOT1 (N3376, N3372);
buf BUF1 (N3377, N3365);
not NOT1 (N3378, N3352);
nor NOR4 (N3379, N3375, N238, N1743, N1256);
nand NAND4 (N3380, N3369, N423, N3061, N546);
buf BUF1 (N3381, N3376);
xor XOR2 (N3382, N3370, N1662);
nand NAND4 (N3383, N3378, N2669, N1673, N1085);
or OR2 (N3384, N3381, N111);
xor XOR2 (N3385, N3379, N3077);
xor XOR2 (N3386, N3385, N411);
and AND3 (N3387, N3377, N20, N1294);
xor XOR2 (N3388, N3383, N2656);
nor NOR4 (N3389, N3384, N3188, N591, N2906);
or OR2 (N3390, N3380, N2684);
xor XOR2 (N3391, N3386, N71);
nor NOR4 (N3392, N3391, N1295, N2943, N1003);
nor NOR2 (N3393, N3359, N2467);
nand NAND4 (N3394, N3388, N2276, N328, N2645);
xor XOR2 (N3395, N3389, N1330);
nand NAND2 (N3396, N3387, N3287);
buf BUF1 (N3397, N3374);
buf BUF1 (N3398, N3394);
not NOT1 (N3399, N3371);
nor NOR4 (N3400, N3395, N2932, N1931, N1197);
and AND3 (N3401, N3382, N1559, N3090);
xor XOR2 (N3402, N3399, N740);
or OR3 (N3403, N3402, N2774, N190);
and AND4 (N3404, N3401, N1991, N171, N1773);
not NOT1 (N3405, N3403);
not NOT1 (N3406, N3368);
or OR3 (N3407, N3397, N3372, N1656);
or OR3 (N3408, N3406, N2073, N1587);
nand NAND2 (N3409, N3396, N2951);
nand NAND3 (N3410, N3390, N3193, N3270);
or OR2 (N3411, N3409, N1426);
nand NAND4 (N3412, N3398, N623, N2025, N119);
nor NOR2 (N3413, N3404, N551);
nor NOR4 (N3414, N3411, N359, N981, N1339);
not NOT1 (N3415, N3392);
not NOT1 (N3416, N3413);
and AND2 (N3417, N3408, N531);
and AND4 (N3418, N3405, N2899, N3187, N735);
buf BUF1 (N3419, N3400);
and AND3 (N3420, N3407, N2648, N3384);
xor XOR2 (N3421, N3412, N2757);
xor XOR2 (N3422, N3415, N1471);
and AND3 (N3423, N3410, N2976, N170);
or OR4 (N3424, N3416, N815, N3422, N488);
buf BUF1 (N3425, N529);
or OR2 (N3426, N3425, N2816);
not NOT1 (N3427, N3418);
and AND4 (N3428, N3426, N439, N586, N2046);
xor XOR2 (N3429, N3420, N2155);
buf BUF1 (N3430, N3414);
and AND3 (N3431, N3428, N1679, N2353);
nand NAND2 (N3432, N3427, N3391);
nand NAND2 (N3433, N3421, N204);
and AND4 (N3434, N3393, N887, N2227, N2536);
not NOT1 (N3435, N3419);
nand NAND2 (N3436, N3433, N597);
not NOT1 (N3437, N3431);
buf BUF1 (N3438, N3424);
buf BUF1 (N3439, N3435);
and AND3 (N3440, N3438, N2365, N2994);
buf BUF1 (N3441, N3439);
nor NOR4 (N3442, N3417, N2484, N2422, N783);
xor XOR2 (N3443, N3436, N2702);
nand NAND3 (N3444, N3437, N2591, N2942);
not NOT1 (N3445, N3432);
or OR3 (N3446, N3429, N65, N1672);
buf BUF1 (N3447, N3445);
xor XOR2 (N3448, N3443, N1206);
buf BUF1 (N3449, N3430);
nor NOR4 (N3450, N3441, N3344, N2929, N151);
nand NAND3 (N3451, N3442, N1658, N119);
buf BUF1 (N3452, N3423);
and AND2 (N3453, N3448, N561);
not NOT1 (N3454, N3452);
nand NAND4 (N3455, N3447, N2255, N2988, N1585);
not NOT1 (N3456, N3455);
or OR2 (N3457, N3434, N177);
not NOT1 (N3458, N3457);
and AND2 (N3459, N3446, N1822);
buf BUF1 (N3460, N3449);
xor XOR2 (N3461, N3450, N2952);
nand NAND4 (N3462, N3459, N2786, N2747, N1397);
nor NOR4 (N3463, N3458, N1363, N2036, N1114);
xor XOR2 (N3464, N3463, N811);
not NOT1 (N3465, N3454);
nor NOR3 (N3466, N3460, N891, N396);
and AND3 (N3467, N3464, N1904, N3011);
nand NAND3 (N3468, N3440, N3141, N1241);
buf BUF1 (N3469, N3456);
or OR4 (N3470, N3453, N3059, N1829, N143);
and AND3 (N3471, N3465, N70, N2250);
nor NOR4 (N3472, N3461, N802, N1087, N1899);
xor XOR2 (N3473, N3467, N2689);
or OR3 (N3474, N3469, N2192, N2260);
xor XOR2 (N3475, N3474, N3421);
not NOT1 (N3476, N3462);
nand NAND3 (N3477, N3476, N2722, N1460);
not NOT1 (N3478, N3470);
and AND4 (N3479, N3475, N2857, N3350, N51);
or OR4 (N3480, N3466, N2213, N384, N987);
not NOT1 (N3481, N3477);
and AND3 (N3482, N3444, N346, N1598);
and AND3 (N3483, N3478, N2718, N1246);
xor XOR2 (N3484, N3483, N1958);
xor XOR2 (N3485, N3471, N110);
nor NOR3 (N3486, N3481, N22, N426);
and AND2 (N3487, N3486, N1945);
xor XOR2 (N3488, N3472, N1285);
xor XOR2 (N3489, N3451, N2296);
xor XOR2 (N3490, N3484, N928);
and AND4 (N3491, N3468, N189, N447, N1571);
not NOT1 (N3492, N3489);
and AND4 (N3493, N3479, N668, N1570, N1806);
xor XOR2 (N3494, N3487, N1506);
xor XOR2 (N3495, N3480, N2740);
xor XOR2 (N3496, N3482, N2188);
or OR2 (N3497, N3492, N3460);
or OR2 (N3498, N3485, N1895);
or OR3 (N3499, N3498, N69, N620);
or OR3 (N3500, N3499, N775, N3333);
or OR2 (N3501, N3500, N760);
nor NOR2 (N3502, N3473, N646);
nor NOR2 (N3503, N3495, N2930);
nand NAND4 (N3504, N3501, N1243, N2182, N2934);
or OR2 (N3505, N3502, N436);
buf BUF1 (N3506, N3504);
buf BUF1 (N3507, N3490);
buf BUF1 (N3508, N3488);
xor XOR2 (N3509, N3496, N2022);
not NOT1 (N3510, N3505);
or OR3 (N3511, N3508, N61, N1331);
buf BUF1 (N3512, N3510);
or OR4 (N3513, N3512, N1797, N3313, N1876);
xor XOR2 (N3514, N3497, N1992);
nand NAND3 (N3515, N3511, N380, N2104);
and AND2 (N3516, N3514, N1159);
nor NOR2 (N3517, N3513, N1680);
and AND4 (N3518, N3491, N1392, N2005, N27);
or OR2 (N3519, N3517, N2344);
and AND3 (N3520, N3493, N3142, N1608);
nor NOR3 (N3521, N3516, N2819, N3237);
and AND4 (N3522, N3494, N1903, N732, N1698);
and AND3 (N3523, N3509, N2068, N950);
buf BUF1 (N3524, N3523);
nand NAND4 (N3525, N3518, N2564, N605, N1868);
nand NAND3 (N3526, N3520, N1575, N858);
xor XOR2 (N3527, N3524, N908);
or OR2 (N3528, N3526, N784);
xor XOR2 (N3529, N3519, N2079);
and AND4 (N3530, N3503, N62, N359, N1565);
and AND4 (N3531, N3525, N1517, N580, N1055);
and AND4 (N3532, N3528, N164, N2875, N1699);
buf BUF1 (N3533, N3507);
nand NAND3 (N3534, N3532, N2931, N1266);
buf BUF1 (N3535, N3530);
buf BUF1 (N3536, N3534);
nand NAND4 (N3537, N3515, N2282, N80, N2988);
not NOT1 (N3538, N3506);
nand NAND3 (N3539, N3533, N3247, N2216);
nand NAND2 (N3540, N3538, N1692);
xor XOR2 (N3541, N3531, N1887);
nand NAND3 (N3542, N3529, N2719, N822);
and AND4 (N3543, N3537, N1534, N2479, N1562);
not NOT1 (N3544, N3539);
nor NOR4 (N3545, N3544, N940, N1584, N3021);
xor XOR2 (N3546, N3541, N253);
xor XOR2 (N3547, N3545, N1866);
nor NOR3 (N3548, N3527, N2837, N2108);
buf BUF1 (N3549, N3548);
nand NAND2 (N3550, N3547, N2698);
buf BUF1 (N3551, N3535);
nand NAND2 (N3552, N3550, N2557);
nand NAND2 (N3553, N3521, N3128);
xor XOR2 (N3554, N3536, N2416);
xor XOR2 (N3555, N3551, N1619);
or OR2 (N3556, N3552, N3204);
and AND2 (N3557, N3540, N2379);
buf BUF1 (N3558, N3554);
nand NAND2 (N3559, N3549, N67);
or OR2 (N3560, N3559, N2941);
nand NAND4 (N3561, N3555, N1769, N426, N3193);
and AND2 (N3562, N3557, N3305);
buf BUF1 (N3563, N3562);
not NOT1 (N3564, N3558);
not NOT1 (N3565, N3522);
buf BUF1 (N3566, N3564);
or OR4 (N3567, N3543, N1860, N2633, N1265);
buf BUF1 (N3568, N3567);
or OR2 (N3569, N3561, N2644);
or OR2 (N3570, N3566, N1433);
or OR4 (N3571, N3570, N1303, N1725, N2);
nor NOR2 (N3572, N3546, N191);
and AND3 (N3573, N3542, N308, N377);
or OR4 (N3574, N3565, N998, N3249, N754);
or OR2 (N3575, N3553, N3248);
xor XOR2 (N3576, N3556, N2693);
buf BUF1 (N3577, N3574);
nand NAND4 (N3578, N3571, N956, N825, N79);
buf BUF1 (N3579, N3578);
not NOT1 (N3580, N3573);
nand NAND2 (N3581, N3568, N2534);
nand NAND3 (N3582, N3560, N313, N1267);
nor NOR3 (N3583, N3569, N1656, N2002);
or OR4 (N3584, N3581, N2318, N3064, N629);
xor XOR2 (N3585, N3572, N2487);
nor NOR2 (N3586, N3579, N418);
and AND3 (N3587, N3563, N1587, N2365);
or OR3 (N3588, N3582, N675, N488);
buf BUF1 (N3589, N3588);
buf BUF1 (N3590, N3575);
and AND2 (N3591, N3584, N3087);
and AND2 (N3592, N3590, N2971);
nor NOR4 (N3593, N3589, N180, N3251, N1316);
not NOT1 (N3594, N3576);
or OR3 (N3595, N3592, N954, N1335);
and AND4 (N3596, N3577, N3538, N3190, N114);
not NOT1 (N3597, N3594);
nand NAND3 (N3598, N3580, N411, N927);
or OR2 (N3599, N3585, N4);
not NOT1 (N3600, N3586);
and AND4 (N3601, N3593, N2100, N662, N3447);
buf BUF1 (N3602, N3600);
nand NAND2 (N3603, N3597, N3114);
nor NOR2 (N3604, N3601, N2739);
nor NOR4 (N3605, N3587, N3422, N542, N2167);
buf BUF1 (N3606, N3583);
not NOT1 (N3607, N3596);
nor NOR4 (N3608, N3607, N2236, N1043, N100);
nand NAND4 (N3609, N3602, N304, N454, N1158);
xor XOR2 (N3610, N3598, N2123);
or OR4 (N3611, N3604, N1172, N3547, N2116);
or OR4 (N3612, N3603, N3600, N9, N107);
not NOT1 (N3613, N3599);
nor NOR4 (N3614, N3591, N1698, N1024, N1567);
or OR3 (N3615, N3605, N2122, N2673);
nand NAND2 (N3616, N3615, N1633);
or OR4 (N3617, N3611, N2889, N960, N70);
and AND4 (N3618, N3609, N455, N1263, N688);
and AND2 (N3619, N3613, N969);
buf BUF1 (N3620, N3614);
buf BUF1 (N3621, N3612);
nor NOR3 (N3622, N3617, N1700, N2362);
xor XOR2 (N3623, N3610, N1234);
buf BUF1 (N3624, N3608);
buf BUF1 (N3625, N3618);
nand NAND3 (N3626, N3595, N2916, N3448);
nand NAND2 (N3627, N3622, N3624);
or OR3 (N3628, N2938, N1854, N388);
or OR2 (N3629, N3616, N2944);
nand NAND2 (N3630, N3629, N3615);
and AND4 (N3631, N3630, N761, N1278, N2032);
nor NOR3 (N3632, N3628, N1120, N1135);
not NOT1 (N3633, N3627);
xor XOR2 (N3634, N3623, N319);
buf BUF1 (N3635, N3631);
nand NAND2 (N3636, N3619, N621);
or OR2 (N3637, N3636, N631);
and AND4 (N3638, N3634, N546, N3406, N203);
and AND3 (N3639, N3621, N2455, N3124);
xor XOR2 (N3640, N3633, N3016);
xor XOR2 (N3641, N3637, N1374);
not NOT1 (N3642, N3639);
not NOT1 (N3643, N3606);
nor NOR4 (N3644, N3632, N2637, N2116, N732);
xor XOR2 (N3645, N3640, N3176);
or OR4 (N3646, N3620, N2075, N2763, N1475);
nand NAND2 (N3647, N3638, N651);
nor NOR2 (N3648, N3626, N2455);
or OR4 (N3649, N3644, N219, N2329, N1319);
not NOT1 (N3650, N3646);
buf BUF1 (N3651, N3650);
nand NAND2 (N3652, N3625, N622);
not NOT1 (N3653, N3652);
and AND4 (N3654, N3647, N2623, N1541, N1220);
buf BUF1 (N3655, N3654);
and AND4 (N3656, N3635, N3149, N2006, N1758);
not NOT1 (N3657, N3655);
not NOT1 (N3658, N3651);
xor XOR2 (N3659, N3643, N1007);
buf BUF1 (N3660, N3659);
nand NAND2 (N3661, N3656, N2191);
nand NAND4 (N3662, N3641, N2165, N2636, N2069);
nor NOR4 (N3663, N3653, N1977, N1765, N2281);
xor XOR2 (N3664, N3648, N2385);
xor XOR2 (N3665, N3663, N2975);
xor XOR2 (N3666, N3662, N3651);
and AND2 (N3667, N3665, N1803);
nor NOR2 (N3668, N3660, N2767);
and AND2 (N3669, N3661, N1400);
and AND3 (N3670, N3645, N462, N3197);
or OR4 (N3671, N3658, N1786, N740, N1381);
or OR2 (N3672, N3664, N909);
nand NAND3 (N3673, N3668, N2716, N3178);
and AND3 (N3674, N3673, N900, N298);
buf BUF1 (N3675, N3667);
nor NOR4 (N3676, N3674, N2528, N3592, N125);
not NOT1 (N3677, N3669);
and AND3 (N3678, N3649, N760, N782);
and AND2 (N3679, N3657, N1479);
or OR4 (N3680, N3679, N2780, N3087, N1585);
and AND4 (N3681, N3680, N1990, N3235, N1179);
and AND3 (N3682, N3681, N3361, N1322);
or OR2 (N3683, N3678, N810);
not NOT1 (N3684, N3682);
nand NAND4 (N3685, N3676, N2277, N1853, N1118);
not NOT1 (N3686, N3683);
buf BUF1 (N3687, N3671);
not NOT1 (N3688, N3684);
and AND3 (N3689, N3675, N576, N1663);
and AND4 (N3690, N3687, N3576, N933, N2043);
and AND3 (N3691, N3666, N314, N2588);
nand NAND3 (N3692, N3672, N2888, N1040);
and AND2 (N3693, N3688, N2190);
and AND2 (N3694, N3642, N968);
or OR4 (N3695, N3693, N950, N2242, N1483);
nand NAND3 (N3696, N3689, N923, N296);
buf BUF1 (N3697, N3695);
or OR4 (N3698, N3685, N2307, N2185, N3661);
nor NOR2 (N3699, N3694, N464);
or OR2 (N3700, N3692, N576);
nor NOR3 (N3701, N3690, N3282, N1215);
not NOT1 (N3702, N3670);
not NOT1 (N3703, N3701);
nor NOR4 (N3704, N3703, N730, N3277, N2367);
not NOT1 (N3705, N3702);
or OR3 (N3706, N3696, N1359, N923);
buf BUF1 (N3707, N3700);
nor NOR3 (N3708, N3706, N3321, N1166);
and AND4 (N3709, N3691, N654, N1934, N1594);
not NOT1 (N3710, N3707);
and AND2 (N3711, N3709, N2711);
and AND3 (N3712, N3698, N2182, N2795);
buf BUF1 (N3713, N3711);
and AND4 (N3714, N3697, N3651, N3414, N539);
nand NAND3 (N3715, N3714, N1942, N173);
nand NAND3 (N3716, N3712, N2040, N1997);
and AND2 (N3717, N3713, N432);
and AND4 (N3718, N3716, N2269, N840, N3455);
and AND3 (N3719, N3677, N575, N2790);
or OR3 (N3720, N3705, N1468, N168);
and AND2 (N3721, N3717, N2299);
nor NOR4 (N3722, N3708, N688, N2015, N2420);
or OR2 (N3723, N3720, N2828);
buf BUF1 (N3724, N3710);
xor XOR2 (N3725, N3719, N1424);
xor XOR2 (N3726, N3723, N2167);
nor NOR2 (N3727, N3724, N558);
not NOT1 (N3728, N3718);
nor NOR2 (N3729, N3715, N3237);
and AND4 (N3730, N3686, N2698, N3511, N2894);
and AND2 (N3731, N3729, N2150);
buf BUF1 (N3732, N3722);
or OR2 (N3733, N3721, N2187);
and AND2 (N3734, N3726, N3045);
and AND3 (N3735, N3733, N695, N2251);
nand NAND4 (N3736, N3735, N2506, N2518, N1878);
nand NAND3 (N3737, N3734, N3287, N2501);
nand NAND2 (N3738, N3730, N3704);
and AND2 (N3739, N592, N3718);
nor NOR2 (N3740, N3728, N1322);
or OR4 (N3741, N3725, N2856, N116, N2698);
and AND3 (N3742, N3736, N2685, N167);
and AND3 (N3743, N3737, N732, N3554);
and AND4 (N3744, N3741, N3663, N1251, N3732);
nor NOR3 (N3745, N1749, N2103, N2060);
and AND2 (N3746, N3739, N3563);
xor XOR2 (N3747, N3742, N2049);
or OR4 (N3748, N3727, N1780, N3687, N1438);
and AND2 (N3749, N3748, N1327);
or OR3 (N3750, N3743, N2184, N1156);
xor XOR2 (N3751, N3731, N2071);
buf BUF1 (N3752, N3746);
and AND4 (N3753, N3699, N1111, N3339, N3169);
xor XOR2 (N3754, N3740, N1848);
nand NAND4 (N3755, N3754, N2074, N2061, N2003);
not NOT1 (N3756, N3745);
nor NOR3 (N3757, N3751, N1690, N762);
nand NAND3 (N3758, N3744, N2567, N533);
nand NAND3 (N3759, N3747, N1321, N585);
and AND4 (N3760, N3738, N2750, N2084, N3708);
not NOT1 (N3761, N3758);
and AND3 (N3762, N3753, N2636, N114);
nor NOR4 (N3763, N3755, N1313, N472, N2413);
nor NOR4 (N3764, N3752, N1375, N3291, N3429);
xor XOR2 (N3765, N3759, N3424);
or OR3 (N3766, N3761, N1505, N2082);
nand NAND4 (N3767, N3765, N1559, N2822, N2329);
nand NAND2 (N3768, N3756, N1542);
not NOT1 (N3769, N3750);
nor NOR3 (N3770, N3767, N2101, N2011);
nor NOR4 (N3771, N3757, N3377, N1443, N1597);
buf BUF1 (N3772, N3749);
nand NAND4 (N3773, N3768, N3210, N1304, N1719);
nor NOR3 (N3774, N3760, N3189, N2414);
nand NAND2 (N3775, N3766, N710);
buf BUF1 (N3776, N3764);
or OR4 (N3777, N3763, N2642, N3318, N2500);
nor NOR2 (N3778, N3762, N528);
buf BUF1 (N3779, N3777);
or OR4 (N3780, N3770, N699, N2374, N3201);
buf BUF1 (N3781, N3778);
nor NOR3 (N3782, N3771, N2440, N496);
buf BUF1 (N3783, N3781);
nand NAND4 (N3784, N3783, N81, N192, N1871);
not NOT1 (N3785, N3784);
xor XOR2 (N3786, N3775, N1044);
xor XOR2 (N3787, N3774, N204);
nand NAND4 (N3788, N3773, N1024, N2713, N253);
buf BUF1 (N3789, N3776);
nand NAND4 (N3790, N3769, N3104, N2904, N3115);
or OR3 (N3791, N3780, N790, N354);
not NOT1 (N3792, N3788);
xor XOR2 (N3793, N3779, N2313);
xor XOR2 (N3794, N3790, N1410);
or OR2 (N3795, N3793, N1047);
not NOT1 (N3796, N3787);
xor XOR2 (N3797, N3789, N3224);
and AND2 (N3798, N3797, N2318);
nor NOR3 (N3799, N3772, N1046, N3307);
xor XOR2 (N3800, N3796, N3462);
xor XOR2 (N3801, N3798, N605);
or OR4 (N3802, N3795, N31, N2342, N2323);
or OR4 (N3803, N3802, N1695, N1247, N1481);
or OR4 (N3804, N3782, N1980, N3710, N3701);
xor XOR2 (N3805, N3794, N3756);
not NOT1 (N3806, N3786);
buf BUF1 (N3807, N3806);
nand NAND4 (N3808, N3801, N2981, N1421, N2600);
and AND3 (N3809, N3800, N1920, N3283);
nand NAND4 (N3810, N3807, N3627, N2246, N302);
buf BUF1 (N3811, N3804);
nor NOR2 (N3812, N3810, N1362);
nand NAND4 (N3813, N3805, N1647, N3346, N1408);
and AND4 (N3814, N3785, N1684, N2445, N479);
not NOT1 (N3815, N3791);
buf BUF1 (N3816, N3809);
buf BUF1 (N3817, N3799);
xor XOR2 (N3818, N3816, N148);
xor XOR2 (N3819, N3817, N3578);
nor NOR3 (N3820, N3812, N2243, N3146);
buf BUF1 (N3821, N3792);
buf BUF1 (N3822, N3811);
nand NAND2 (N3823, N3813, N2733);
not NOT1 (N3824, N3814);
nor NOR3 (N3825, N3815, N259, N1660);
xor XOR2 (N3826, N3808, N1387);
nor NOR4 (N3827, N3818, N373, N2763, N1030);
not NOT1 (N3828, N3824);
not NOT1 (N3829, N3823);
nor NOR3 (N3830, N3820, N51, N2165);
or OR3 (N3831, N3825, N300, N848);
or OR3 (N3832, N3822, N551, N2805);
nor NOR2 (N3833, N3832, N2123);
or OR4 (N3834, N3821, N1174, N3208, N560);
nor NOR4 (N3835, N3826, N1278, N3557, N3792);
nand NAND3 (N3836, N3833, N2304, N1959);
and AND3 (N3837, N3830, N2503, N1365);
buf BUF1 (N3838, N3831);
not NOT1 (N3839, N3838);
not NOT1 (N3840, N3803);
nand NAND2 (N3841, N3819, N3592);
xor XOR2 (N3842, N3834, N1289);
and AND4 (N3843, N3841, N1404, N2329, N3690);
or OR3 (N3844, N3828, N2171, N3100);
and AND4 (N3845, N3842, N1182, N334, N2284);
and AND4 (N3846, N3843, N873, N3627, N2299);
or OR2 (N3847, N3846, N1705);
buf BUF1 (N3848, N3835);
xor XOR2 (N3849, N3839, N2745);
xor XOR2 (N3850, N3837, N1376);
or OR3 (N3851, N3847, N3602, N3840);
not NOT1 (N3852, N2738);
not NOT1 (N3853, N3852);
not NOT1 (N3854, N3848);
not NOT1 (N3855, N3853);
nand NAND4 (N3856, N3829, N2617, N999, N1889);
nand NAND2 (N3857, N3854, N2183);
and AND4 (N3858, N3856, N3267, N93, N2838);
not NOT1 (N3859, N3836);
xor XOR2 (N3860, N3851, N1580);
nand NAND2 (N3861, N3857, N3166);
not NOT1 (N3862, N3859);
xor XOR2 (N3863, N3850, N1158);
nand NAND4 (N3864, N3862, N1061, N859, N2790);
nand NAND3 (N3865, N3855, N923, N2740);
nor NOR4 (N3866, N3845, N2891, N138, N3512);
and AND3 (N3867, N3844, N302, N3288);
and AND2 (N3868, N3866, N214);
nand NAND3 (N3869, N3860, N2410, N2386);
nand NAND2 (N3870, N3863, N1559);
or OR2 (N3871, N3864, N3103);
nand NAND3 (N3872, N3871, N3701, N195);
xor XOR2 (N3873, N3858, N3828);
or OR2 (N3874, N3849, N2043);
xor XOR2 (N3875, N3865, N2868);
and AND3 (N3876, N3867, N2221, N1146);
buf BUF1 (N3877, N3872);
not NOT1 (N3878, N3869);
not NOT1 (N3879, N3875);
buf BUF1 (N3880, N3877);
nand NAND2 (N3881, N3827, N2009);
xor XOR2 (N3882, N3878, N2424);
nor NOR2 (N3883, N3876, N3457);
xor XOR2 (N3884, N3879, N2968);
buf BUF1 (N3885, N3883);
not NOT1 (N3886, N3868);
and AND3 (N3887, N3881, N1425, N3264);
xor XOR2 (N3888, N3886, N2911);
xor XOR2 (N3889, N3873, N1019);
not NOT1 (N3890, N3884);
buf BUF1 (N3891, N3882);
not NOT1 (N3892, N3874);
nor NOR3 (N3893, N3880, N2936, N3405);
or OR4 (N3894, N3893, N679, N1386, N498);
or OR2 (N3895, N3887, N3516);
nand NAND3 (N3896, N3890, N1692, N1257);
buf BUF1 (N3897, N3861);
or OR3 (N3898, N3894, N680, N2144);
and AND2 (N3899, N3895, N1180);
buf BUF1 (N3900, N3898);
nand NAND4 (N3901, N3889, N1832, N2208, N528);
and AND4 (N3902, N3891, N2061, N776, N2489);
nand NAND4 (N3903, N3870, N3880, N97, N1916);
nand NAND3 (N3904, N3902, N988, N1173);
and AND2 (N3905, N3904, N2133);
or OR4 (N3906, N3888, N3798, N2265, N1683);
not NOT1 (N3907, N3892);
or OR3 (N3908, N3906, N1239, N1231);
not NOT1 (N3909, N3905);
not NOT1 (N3910, N3908);
buf BUF1 (N3911, N3885);
nor NOR4 (N3912, N3909, N3465, N1007, N865);
buf BUF1 (N3913, N3910);
not NOT1 (N3914, N3911);
buf BUF1 (N3915, N3896);
nor NOR4 (N3916, N3897, N3752, N311, N3748);
nand NAND3 (N3917, N3903, N475, N3389);
and AND4 (N3918, N3899, N929, N1303, N811);
and AND4 (N3919, N3901, N3130, N2276, N1681);
buf BUF1 (N3920, N3917);
nor NOR3 (N3921, N3907, N257, N2666);
not NOT1 (N3922, N3921);
and AND3 (N3923, N3912, N1910, N2076);
xor XOR2 (N3924, N3915, N2232);
buf BUF1 (N3925, N3919);
or OR4 (N3926, N3920, N576, N638, N1820);
or OR4 (N3927, N3913, N3144, N1984, N2347);
xor XOR2 (N3928, N3924, N339);
and AND3 (N3929, N3914, N359, N1185);
buf BUF1 (N3930, N3918);
not NOT1 (N3931, N3926);
or OR2 (N3932, N3922, N762);
xor XOR2 (N3933, N3928, N24);
or OR3 (N3934, N3923, N2071, N384);
xor XOR2 (N3935, N3929, N3191);
xor XOR2 (N3936, N3925, N3889);
nand NAND4 (N3937, N3935, N3766, N1521, N2087);
xor XOR2 (N3938, N3900, N472);
and AND3 (N3939, N3916, N205, N2940);
nor NOR4 (N3940, N3936, N3020, N1086, N140);
not NOT1 (N3941, N3927);
and AND2 (N3942, N3937, N3819);
not NOT1 (N3943, N3939);
and AND4 (N3944, N3933, N1036, N1057, N1882);
xor XOR2 (N3945, N3941, N634);
buf BUF1 (N3946, N3930);
and AND4 (N3947, N3934, N1106, N583, N374);
buf BUF1 (N3948, N3943);
not NOT1 (N3949, N3932);
or OR3 (N3950, N3947, N3483, N3716);
xor XOR2 (N3951, N3950, N1272);
not NOT1 (N3952, N3948);
xor XOR2 (N3953, N3938, N2466);
not NOT1 (N3954, N3931);
xor XOR2 (N3955, N3953, N3475);
xor XOR2 (N3956, N3949, N1293);
xor XOR2 (N3957, N3946, N2435);
or OR4 (N3958, N3942, N152, N2460, N3892);
not NOT1 (N3959, N3952);
not NOT1 (N3960, N3944);
buf BUF1 (N3961, N3957);
or OR4 (N3962, N3940, N462, N644, N347);
nor NOR4 (N3963, N3956, N2677, N143, N1192);
nand NAND4 (N3964, N3958, N647, N2157, N2340);
nand NAND2 (N3965, N3960, N2950);
buf BUF1 (N3966, N3954);
xor XOR2 (N3967, N3962, N3163);
nand NAND4 (N3968, N3966, N3628, N2113, N3615);
nor NOR3 (N3969, N3945, N318, N3838);
or OR2 (N3970, N3965, N1926);
nor NOR3 (N3971, N3963, N3368, N2961);
nor NOR4 (N3972, N3969, N3201, N2843, N30);
nand NAND3 (N3973, N3959, N2524, N956);
and AND2 (N3974, N3964, N3932);
not NOT1 (N3975, N3968);
or OR4 (N3976, N3970, N2653, N2065, N577);
and AND4 (N3977, N3955, N50, N318, N1863);
nor NOR3 (N3978, N3973, N2439, N3548);
nor NOR4 (N3979, N3972, N763, N2435, N300);
xor XOR2 (N3980, N3951, N609);
nor NOR3 (N3981, N3976, N2128, N1418);
or OR4 (N3982, N3974, N107, N1853, N2476);
xor XOR2 (N3983, N3977, N2442);
buf BUF1 (N3984, N3975);
buf BUF1 (N3985, N3984);
nor NOR2 (N3986, N3985, N2870);
not NOT1 (N3987, N3980);
or OR4 (N3988, N3967, N338, N2006, N2589);
or OR2 (N3989, N3983, N3203);
nand NAND3 (N3990, N3989, N1883, N1756);
nor NOR2 (N3991, N3978, N3475);
buf BUF1 (N3992, N3991);
nand NAND2 (N3993, N3961, N2951);
not NOT1 (N3994, N3986);
xor XOR2 (N3995, N3993, N385);
and AND4 (N3996, N3990, N1221, N1694, N2883);
and AND2 (N3997, N3979, N3391);
not NOT1 (N3998, N3971);
buf BUF1 (N3999, N3987);
and AND3 (N4000, N3992, N1190, N1166);
nand NAND4 (N4001, N3997, N3217, N395, N225);
and AND2 (N4002, N3998, N222);
buf BUF1 (N4003, N3996);
and AND3 (N4004, N4002, N2564, N2951);
nor NOR3 (N4005, N3988, N907, N508);
buf BUF1 (N4006, N4004);
nor NOR4 (N4007, N3982, N44, N1196, N2241);
nor NOR4 (N4008, N4000, N3485, N3116, N2947);
buf BUF1 (N4009, N3994);
and AND4 (N4010, N4009, N2406, N2991, N1711);
buf BUF1 (N4011, N4003);
nand NAND2 (N4012, N3995, N45);
nor NOR2 (N4013, N4012, N1901);
not NOT1 (N4014, N4013);
or OR4 (N4015, N4006, N812, N2960, N315);
or OR2 (N4016, N4010, N1194);
buf BUF1 (N4017, N3999);
xor XOR2 (N4018, N4016, N55);
nand NAND2 (N4019, N4001, N3447);
nand NAND2 (N4020, N4011, N3483);
nand NAND3 (N4021, N4019, N3348, N2290);
buf BUF1 (N4022, N4020);
nor NOR4 (N4023, N4008, N2772, N1727, N3895);
nor NOR4 (N4024, N4023, N282, N3125, N281);
and AND3 (N4025, N4017, N3407, N3748);
buf BUF1 (N4026, N4007);
xor XOR2 (N4027, N4025, N495);
buf BUF1 (N4028, N4022);
buf BUF1 (N4029, N4021);
xor XOR2 (N4030, N3981, N485);
and AND3 (N4031, N4014, N1658, N361);
buf BUF1 (N4032, N4030);
not NOT1 (N4033, N4018);
not NOT1 (N4034, N4032);
buf BUF1 (N4035, N4028);
nand NAND3 (N4036, N4015, N1266, N855);
nor NOR3 (N4037, N4027, N1033, N1734);
nor NOR2 (N4038, N4005, N1143);
nor NOR2 (N4039, N4034, N3438);
nor NOR4 (N4040, N4033, N3616, N2155, N3816);
or OR4 (N4041, N4026, N1930, N356, N1244);
nand NAND4 (N4042, N4024, N2920, N3417, N3523);
nor NOR4 (N4043, N4038, N2065, N958, N555);
nor NOR4 (N4044, N4035, N1003, N3253, N3116);
or OR2 (N4045, N4042, N2823);
nand NAND2 (N4046, N4029, N565);
nor NOR3 (N4047, N4041, N3070, N1192);
not NOT1 (N4048, N4039);
nor NOR2 (N4049, N4040, N1749);
not NOT1 (N4050, N4036);
buf BUF1 (N4051, N4044);
or OR2 (N4052, N4048, N1883);
or OR4 (N4053, N4043, N3293, N884, N1622);
nand NAND2 (N4054, N4053, N1236);
not NOT1 (N4055, N4031);
nand NAND3 (N4056, N4046, N691, N3513);
not NOT1 (N4057, N4054);
or OR3 (N4058, N4050, N2117, N842);
not NOT1 (N4059, N4051);
or OR4 (N4060, N4055, N3132, N2226, N324);
or OR3 (N4061, N4052, N2884, N2002);
buf BUF1 (N4062, N4056);
nor NOR3 (N4063, N4061, N2106, N3199);
and AND3 (N4064, N4060, N3963, N3560);
nor NOR2 (N4065, N4045, N1145);
buf BUF1 (N4066, N4064);
nand NAND2 (N4067, N4063, N1592);
buf BUF1 (N4068, N4057);
or OR3 (N4069, N4059, N1021, N1514);
xor XOR2 (N4070, N4068, N460);
not NOT1 (N4071, N4070);
nor NOR2 (N4072, N4065, N2929);
xor XOR2 (N4073, N4049, N3259);
buf BUF1 (N4074, N4058);
nand NAND2 (N4075, N4071, N4040);
not NOT1 (N4076, N4073);
or OR4 (N4077, N4067, N3789, N1255, N1140);
and AND4 (N4078, N4076, N1525, N1951, N3117);
not NOT1 (N4079, N4069);
not NOT1 (N4080, N4047);
buf BUF1 (N4081, N4077);
buf BUF1 (N4082, N4080);
and AND3 (N4083, N4062, N1384, N4076);
nor NOR4 (N4084, N4082, N3076, N515, N562);
nand NAND4 (N4085, N4074, N2438, N1094, N3113);
or OR3 (N4086, N4072, N2035, N1221);
and AND3 (N4087, N4078, N2318, N3175);
nor NOR3 (N4088, N4066, N106, N2544);
nor NOR4 (N4089, N4079, N3566, N738, N1369);
and AND2 (N4090, N4085, N2638);
nor NOR2 (N4091, N4037, N3940);
buf BUF1 (N4092, N4090);
and AND4 (N4093, N4089, N2218, N3327, N1580);
xor XOR2 (N4094, N4084, N751);
nand NAND2 (N4095, N4083, N3732);
not NOT1 (N4096, N4093);
buf BUF1 (N4097, N4086);
nand NAND3 (N4098, N4091, N3481, N1482);
not NOT1 (N4099, N4092);
and AND2 (N4100, N4098, N1366);
or OR3 (N4101, N4095, N776, N3282);
xor XOR2 (N4102, N4099, N787);
buf BUF1 (N4103, N4096);
not NOT1 (N4104, N4100);
not NOT1 (N4105, N4088);
not NOT1 (N4106, N4104);
not NOT1 (N4107, N4097);
not NOT1 (N4108, N4075);
nor NOR2 (N4109, N4087, N1087);
nand NAND4 (N4110, N4102, N1393, N2107, N1883);
not NOT1 (N4111, N4105);
nor NOR3 (N4112, N4103, N2212, N1640);
nand NAND3 (N4113, N4106, N2548, N2038);
nor NOR4 (N4114, N4094, N192, N2092, N58);
nand NAND4 (N4115, N4113, N3933, N814, N3628);
xor XOR2 (N4116, N4114, N2714);
buf BUF1 (N4117, N4107);
and AND2 (N4118, N4117, N411);
nor NOR4 (N4119, N4118, N284, N2306, N2806);
not NOT1 (N4120, N4115);
buf BUF1 (N4121, N4119);
or OR4 (N4122, N4121, N3349, N1372, N2384);
nand NAND3 (N4123, N4101, N3142, N1676);
nand NAND2 (N4124, N4108, N2756);
or OR4 (N4125, N4122, N3548, N2155, N119);
and AND2 (N4126, N4109, N2324);
nor NOR3 (N4127, N4120, N2987, N777);
not NOT1 (N4128, N4123);
not NOT1 (N4129, N4128);
and AND2 (N4130, N4129, N3123);
or OR3 (N4131, N4130, N3140, N1861);
xor XOR2 (N4132, N4124, N3606);
nor NOR3 (N4133, N4125, N21, N1840);
and AND2 (N4134, N4133, N830);
and AND3 (N4135, N4111, N2756, N2338);
or OR3 (N4136, N4131, N1555, N2340);
and AND3 (N4137, N4132, N881, N1506);
not NOT1 (N4138, N4136);
xor XOR2 (N4139, N4110, N3899);
nand NAND4 (N4140, N4137, N14, N2883, N1892);
or OR3 (N4141, N4081, N3219, N4002);
not NOT1 (N4142, N4135);
and AND3 (N4143, N4127, N2456, N1448);
or OR2 (N4144, N4112, N1140);
xor XOR2 (N4145, N4141, N2306);
buf BUF1 (N4146, N4134);
and AND2 (N4147, N4126, N128);
nor NOR3 (N4148, N4146, N2951, N3325);
buf BUF1 (N4149, N4140);
or OR3 (N4150, N4139, N4032, N3198);
nand NAND2 (N4151, N4143, N1589);
not NOT1 (N4152, N4142);
nor NOR4 (N4153, N4151, N1621, N613, N2738);
or OR3 (N4154, N4149, N1919, N3679);
nor NOR2 (N4155, N4154, N2511);
or OR2 (N4156, N4138, N3034);
xor XOR2 (N4157, N4145, N2371);
not NOT1 (N4158, N4155);
or OR3 (N4159, N4116, N7, N1836);
xor XOR2 (N4160, N4159, N1554);
nor NOR2 (N4161, N4157, N4063);
xor XOR2 (N4162, N4153, N3622);
and AND2 (N4163, N4158, N3390);
xor XOR2 (N4164, N4147, N57);
xor XOR2 (N4165, N4163, N2644);
not NOT1 (N4166, N4160);
buf BUF1 (N4167, N4162);
nand NAND4 (N4168, N4167, N3990, N2826, N1743);
and AND4 (N4169, N4165, N2990, N1943, N2213);
nand NAND2 (N4170, N4148, N3772);
buf BUF1 (N4171, N4150);
nor NOR2 (N4172, N4171, N4139);
or OR4 (N4173, N4164, N2956, N2784, N4087);
or OR3 (N4174, N4152, N2146, N2477);
nor NOR4 (N4175, N4174, N3371, N2997, N3923);
or OR3 (N4176, N4169, N214, N2696);
nand NAND3 (N4177, N4176, N2128, N1496);
and AND4 (N4178, N4175, N1871, N2998, N2397);
buf BUF1 (N4179, N4170);
xor XOR2 (N4180, N4156, N4118);
xor XOR2 (N4181, N4177, N2315);
xor XOR2 (N4182, N4178, N2539);
or OR3 (N4183, N4179, N89, N988);
or OR4 (N4184, N4144, N3934, N3924, N3876);
or OR3 (N4185, N4183, N2076, N2228);
and AND4 (N4186, N4185, N788, N1572, N4033);
buf BUF1 (N4187, N4184);
or OR4 (N4188, N4180, N185, N649, N2508);
buf BUF1 (N4189, N4187);
xor XOR2 (N4190, N4181, N3230);
nor NOR4 (N4191, N4173, N702, N2517, N2232);
buf BUF1 (N4192, N4168);
nand NAND3 (N4193, N4186, N2780, N4146);
and AND3 (N4194, N4188, N176, N3938);
nand NAND4 (N4195, N4192, N173, N251, N2270);
or OR2 (N4196, N4191, N2164);
not NOT1 (N4197, N4172);
or OR2 (N4198, N4190, N3138);
not NOT1 (N4199, N4198);
or OR4 (N4200, N4196, N3192, N126, N3924);
and AND3 (N4201, N4199, N503, N1425);
nor NOR4 (N4202, N4161, N3203, N2871, N2077);
buf BUF1 (N4203, N4182);
or OR2 (N4204, N4189, N2458);
nor NOR3 (N4205, N4203, N1818, N2009);
nand NAND3 (N4206, N4202, N1825, N1529);
not NOT1 (N4207, N4166);
buf BUF1 (N4208, N4206);
nand NAND4 (N4209, N4197, N864, N3361, N2912);
nand NAND3 (N4210, N4207, N505, N3255);
nor NOR4 (N4211, N4194, N819, N4084, N2348);
xor XOR2 (N4212, N4211, N3764);
nand NAND3 (N4213, N4212, N461, N4112);
not NOT1 (N4214, N4195);
and AND3 (N4215, N4200, N1130, N1916);
nor NOR3 (N4216, N4213, N2440, N3799);
buf BUF1 (N4217, N4205);
buf BUF1 (N4218, N4204);
and AND2 (N4219, N4208, N1676);
and AND3 (N4220, N4193, N1442, N303);
xor XOR2 (N4221, N4215, N1880);
not NOT1 (N4222, N4209);
not NOT1 (N4223, N4219);
buf BUF1 (N4224, N4218);
not NOT1 (N4225, N4210);
buf BUF1 (N4226, N4216);
not NOT1 (N4227, N4222);
nand NAND2 (N4228, N4220, N4099);
and AND3 (N4229, N4224, N1026, N2149);
xor XOR2 (N4230, N4201, N1365);
buf BUF1 (N4231, N4227);
nand NAND2 (N4232, N4223, N2058);
nand NAND4 (N4233, N4231, N795, N2315, N2955);
or OR4 (N4234, N4214, N552, N2034, N3390);
nand NAND4 (N4235, N4234, N3410, N1270, N1524);
nor NOR3 (N4236, N4226, N3103, N2616);
xor XOR2 (N4237, N4217, N1740);
not NOT1 (N4238, N4229);
not NOT1 (N4239, N4236);
not NOT1 (N4240, N4230);
buf BUF1 (N4241, N4235);
buf BUF1 (N4242, N4228);
xor XOR2 (N4243, N4225, N1335);
xor XOR2 (N4244, N4232, N1952);
and AND3 (N4245, N4240, N3087, N3020);
buf BUF1 (N4246, N4237);
not NOT1 (N4247, N4233);
or OR3 (N4248, N4246, N2113, N4225);
or OR2 (N4249, N4243, N1448);
and AND2 (N4250, N4249, N2218);
nand NAND2 (N4251, N4248, N3621);
and AND4 (N4252, N4238, N2346, N1003, N1324);
nor NOR3 (N4253, N4239, N2858, N2147);
nor NOR4 (N4254, N4242, N3326, N948, N2642);
nand NAND4 (N4255, N4253, N950, N1451, N2020);
or OR2 (N4256, N4241, N1259);
not NOT1 (N4257, N4255);
nand NAND2 (N4258, N4245, N2917);
nor NOR3 (N4259, N4257, N3887, N3687);
or OR3 (N4260, N4244, N2694, N2644);
xor XOR2 (N4261, N4221, N1681);
not NOT1 (N4262, N4251);
nor NOR3 (N4263, N4259, N2024, N3493);
or OR2 (N4264, N4256, N3829);
buf BUF1 (N4265, N4263);
or OR2 (N4266, N4265, N1354);
xor XOR2 (N4267, N4252, N544);
and AND3 (N4268, N4254, N1712, N952);
or OR4 (N4269, N4247, N3239, N1376, N3571);
xor XOR2 (N4270, N4260, N397);
nor NOR4 (N4271, N4267, N2446, N1873, N3818);
nand NAND2 (N4272, N4268, N3444);
not NOT1 (N4273, N4266);
nor NOR4 (N4274, N4272, N2447, N1759, N4121);
nor NOR4 (N4275, N4262, N1620, N2599, N4232);
nand NAND3 (N4276, N4274, N24, N3527);
or OR3 (N4277, N4261, N2036, N1668);
not NOT1 (N4278, N4264);
or OR4 (N4279, N4250, N2598, N271, N1693);
xor XOR2 (N4280, N4276, N2406);
not NOT1 (N4281, N4280);
nand NAND3 (N4282, N4279, N2293, N1163);
xor XOR2 (N4283, N4281, N1593);
nor NOR2 (N4284, N4269, N4025);
nand NAND4 (N4285, N4258, N900, N3878, N4251);
nor NOR2 (N4286, N4273, N3635);
buf BUF1 (N4287, N4271);
buf BUF1 (N4288, N4275);
not NOT1 (N4289, N4270);
or OR4 (N4290, N4284, N1661, N1874, N590);
nor NOR4 (N4291, N4282, N360, N760, N1301);
and AND4 (N4292, N4283, N3062, N1032, N2750);
buf BUF1 (N4293, N4287);
nand NAND2 (N4294, N4288, N621);
buf BUF1 (N4295, N4291);
xor XOR2 (N4296, N4290, N2023);
nor NOR3 (N4297, N4292, N2112, N2320);
and AND3 (N4298, N4285, N2077, N3967);
and AND3 (N4299, N4286, N3568, N316);
xor XOR2 (N4300, N4293, N3008);
xor XOR2 (N4301, N4295, N49);
xor XOR2 (N4302, N4289, N669);
xor XOR2 (N4303, N4277, N4109);
nor NOR4 (N4304, N4278, N2581, N1354, N2247);
not NOT1 (N4305, N4302);
or OR4 (N4306, N4304, N3748, N4234, N3118);
not NOT1 (N4307, N4296);
not NOT1 (N4308, N4301);
buf BUF1 (N4309, N4307);
xor XOR2 (N4310, N4298, N3897);
nor NOR4 (N4311, N4297, N4025, N1547, N188);
or OR2 (N4312, N4311, N3147);
buf BUF1 (N4313, N4294);
buf BUF1 (N4314, N4310);
and AND4 (N4315, N4299, N1243, N652, N20);
nand NAND3 (N4316, N4312, N1677, N1445);
or OR2 (N4317, N4309, N965);
xor XOR2 (N4318, N4316, N2491);
nor NOR3 (N4319, N4306, N2486, N2507);
nor NOR2 (N4320, N4318, N1567);
xor XOR2 (N4321, N4313, N31);
and AND4 (N4322, N4317, N532, N1529, N2893);
nor NOR2 (N4323, N4303, N2237);
and AND3 (N4324, N4321, N4179, N645);
nor NOR2 (N4325, N4315, N1800);
buf BUF1 (N4326, N4308);
nor NOR4 (N4327, N4322, N2464, N408, N3600);
or OR3 (N4328, N4319, N3977, N1627);
not NOT1 (N4329, N4300);
buf BUF1 (N4330, N4324);
not NOT1 (N4331, N4325);
or OR3 (N4332, N4328, N2463, N708);
nor NOR2 (N4333, N4323, N1829);
or OR2 (N4334, N4320, N133);
buf BUF1 (N4335, N4331);
nand NAND2 (N4336, N4333, N2497);
nand NAND2 (N4337, N4305, N3462);
nand NAND2 (N4338, N4335, N1845);
and AND4 (N4339, N4327, N1822, N354, N2579);
nand NAND2 (N4340, N4336, N402);
and AND4 (N4341, N4340, N205, N842, N2632);
nand NAND4 (N4342, N4330, N4086, N4325, N3508);
or OR3 (N4343, N4339, N1104, N2288);
not NOT1 (N4344, N4342);
and AND3 (N4345, N4314, N3537, N344);
and AND4 (N4346, N4326, N757, N3989, N1559);
nor NOR4 (N4347, N4345, N1567, N2527, N3930);
and AND3 (N4348, N4344, N2334, N1965);
nor NOR3 (N4349, N4343, N1679, N1272);
nor NOR3 (N4350, N4334, N3767, N2590);
nor NOR4 (N4351, N4349, N1437, N409, N3001);
not NOT1 (N4352, N4341);
or OR4 (N4353, N4329, N949, N2186, N4342);
buf BUF1 (N4354, N4350);
or OR3 (N4355, N4348, N1132, N1467);
buf BUF1 (N4356, N4354);
buf BUF1 (N4357, N4356);
xor XOR2 (N4358, N4338, N4150);
and AND3 (N4359, N4352, N358, N2773);
and AND2 (N4360, N4355, N3423);
and AND2 (N4361, N4332, N2149);
nand NAND3 (N4362, N4359, N718, N1889);
and AND3 (N4363, N4361, N586, N1641);
nor NOR3 (N4364, N4346, N1967, N1625);
or OR3 (N4365, N4363, N1441, N2090);
nand NAND3 (N4366, N4365, N21, N4300);
nor NOR3 (N4367, N4366, N1350, N1041);
nor NOR3 (N4368, N4367, N2697, N867);
nor NOR4 (N4369, N4353, N3922, N3236, N1838);
nand NAND2 (N4370, N4357, N111);
xor XOR2 (N4371, N4370, N684);
not NOT1 (N4372, N4347);
xor XOR2 (N4373, N4371, N3796);
nor NOR3 (N4374, N4351, N143, N3468);
xor XOR2 (N4375, N4372, N1394);
buf BUF1 (N4376, N4375);
nand NAND2 (N4377, N4358, N916);
nand NAND2 (N4378, N4369, N2284);
xor XOR2 (N4379, N4374, N3812);
xor XOR2 (N4380, N4368, N780);
not NOT1 (N4381, N4380);
xor XOR2 (N4382, N4377, N4154);
xor XOR2 (N4383, N4337, N1173);
nor NOR3 (N4384, N4376, N1185, N2625);
or OR3 (N4385, N4383, N4197, N715);
or OR4 (N4386, N4379, N1108, N3494, N1172);
or OR4 (N4387, N4360, N1259, N277, N1330);
not NOT1 (N4388, N4378);
nand NAND4 (N4389, N4384, N3956, N3491, N2477);
not NOT1 (N4390, N4381);
nor NOR3 (N4391, N4389, N2712, N4059);
xor XOR2 (N4392, N4364, N2092);
buf BUF1 (N4393, N4387);
nor NOR2 (N4394, N4385, N3572);
and AND4 (N4395, N4390, N1935, N2426, N696);
nand NAND4 (N4396, N4386, N703, N105, N1609);
and AND2 (N4397, N4388, N4359);
or OR2 (N4398, N4396, N2074);
or OR3 (N4399, N4395, N1251, N2303);
not NOT1 (N4400, N4382);
xor XOR2 (N4401, N4362, N1101);
nor NOR2 (N4402, N4373, N2957);
or OR4 (N4403, N4400, N1996, N294, N2379);
xor XOR2 (N4404, N4393, N235);
nand NAND3 (N4405, N4397, N1107, N1491);
not NOT1 (N4406, N4391);
nor NOR4 (N4407, N4405, N2759, N3227, N1478);
and AND2 (N4408, N4398, N762);
nand NAND3 (N4409, N4404, N3466, N1892);
xor XOR2 (N4410, N4409, N2577);
buf BUF1 (N4411, N4399);
xor XOR2 (N4412, N4392, N849);
and AND3 (N4413, N4410, N2085, N3150);
nor NOR4 (N4414, N4394, N3370, N4056, N3441);
xor XOR2 (N4415, N4411, N2326);
nand NAND3 (N4416, N4407, N663, N1766);
nand NAND2 (N4417, N4403, N962);
buf BUF1 (N4418, N4416);
xor XOR2 (N4419, N4413, N533);
not NOT1 (N4420, N4408);
nand NAND2 (N4421, N4401, N1060);
buf BUF1 (N4422, N4421);
nand NAND4 (N4423, N4422, N2519, N2965, N3605);
xor XOR2 (N4424, N4414, N2007);
nor NOR2 (N4425, N4402, N524);
nand NAND2 (N4426, N4419, N1092);
nor NOR2 (N4427, N4406, N1341);
nand NAND3 (N4428, N4426, N1753, N1274);
buf BUF1 (N4429, N4415);
and AND3 (N4430, N4428, N924, N1703);
buf BUF1 (N4431, N4429);
nor NOR4 (N4432, N4418, N4063, N3215, N2932);
not NOT1 (N4433, N4417);
not NOT1 (N4434, N4425);
nor NOR3 (N4435, N4420, N947, N949);
buf BUF1 (N4436, N4432);
or OR4 (N4437, N4435, N4198, N403, N992);
and AND4 (N4438, N4433, N2667, N1679, N2359);
not NOT1 (N4439, N4434);
nor NOR3 (N4440, N4436, N2079, N3561);
and AND2 (N4441, N4430, N1723);
and AND4 (N4442, N4424, N572, N2751, N377);
or OR3 (N4443, N4412, N2883, N3782);
nor NOR3 (N4444, N4443, N3295, N1100);
or OR3 (N4445, N4431, N1899, N1243);
and AND3 (N4446, N4440, N1286, N4404);
buf BUF1 (N4447, N4439);
nor NOR3 (N4448, N4423, N3609, N1935);
buf BUF1 (N4449, N4427);
buf BUF1 (N4450, N4442);
nand NAND4 (N4451, N4438, N3145, N4354, N82);
not NOT1 (N4452, N4446);
not NOT1 (N4453, N4447);
xor XOR2 (N4454, N4451, N2703);
and AND3 (N4455, N4452, N1495, N355);
buf BUF1 (N4456, N4448);
not NOT1 (N4457, N4445);
or OR4 (N4458, N4454, N699, N1570, N3378);
xor XOR2 (N4459, N4449, N1659);
nand NAND4 (N4460, N4457, N3005, N726, N2506);
not NOT1 (N4461, N4453);
nand NAND2 (N4462, N4437, N3901);
nand NAND4 (N4463, N4441, N3871, N3629, N1971);
nor NOR4 (N4464, N4463, N4136, N2600, N464);
xor XOR2 (N4465, N4459, N1288);
buf BUF1 (N4466, N4465);
nand NAND2 (N4467, N4460, N2383);
xor XOR2 (N4468, N4466, N3546);
buf BUF1 (N4469, N4456);
nor NOR2 (N4470, N4468, N2974);
nand NAND3 (N4471, N4455, N1354, N393);
and AND2 (N4472, N4471, N888);
nand NAND3 (N4473, N4444, N3297, N2545);
nor NOR4 (N4474, N4472, N2385, N1559, N3187);
buf BUF1 (N4475, N4458);
not NOT1 (N4476, N4469);
nor NOR3 (N4477, N4467, N2080, N1034);
not NOT1 (N4478, N4464);
or OR4 (N4479, N4474, N706, N3385, N2925);
not NOT1 (N4480, N4478);
nand NAND2 (N4481, N4462, N2408);
or OR4 (N4482, N4477, N1539, N483, N1110);
or OR2 (N4483, N4476, N1686);
nand NAND4 (N4484, N4475, N3950, N3073, N826);
not NOT1 (N4485, N4450);
nand NAND3 (N4486, N4473, N3627, N2005);
nand NAND2 (N4487, N4486, N3896);
not NOT1 (N4488, N4487);
not NOT1 (N4489, N4470);
nand NAND2 (N4490, N4484, N295);
or OR2 (N4491, N4488, N2059);
nand NAND2 (N4492, N4482, N13);
and AND2 (N4493, N4491, N2660);
nor NOR2 (N4494, N4485, N2322);
not NOT1 (N4495, N4461);
or OR2 (N4496, N4492, N2555);
xor XOR2 (N4497, N4483, N3443);
and AND4 (N4498, N4493, N4211, N3681, N228);
xor XOR2 (N4499, N4479, N4371);
buf BUF1 (N4500, N4481);
nand NAND3 (N4501, N4500, N4065, N1761);
not NOT1 (N4502, N4501);
or OR3 (N4503, N4499, N3093, N3995);
nand NAND2 (N4504, N4480, N3876);
nand NAND2 (N4505, N4495, N1578);
buf BUF1 (N4506, N4502);
nand NAND4 (N4507, N4498, N2426, N3449, N1041);
nand NAND3 (N4508, N4506, N3908, N2222);
buf BUF1 (N4509, N4497);
nand NAND3 (N4510, N4504, N3813, N1938);
nor NOR2 (N4511, N4489, N2914);
buf BUF1 (N4512, N4490);
buf BUF1 (N4513, N4508);
not NOT1 (N4514, N4505);
nor NOR4 (N4515, N4509, N2330, N4200, N4019);
xor XOR2 (N4516, N4503, N2393);
or OR3 (N4517, N4511, N2247, N3724);
and AND4 (N4518, N4513, N4087, N2586, N2335);
nor NOR2 (N4519, N4518, N1441);
and AND4 (N4520, N4514, N2772, N147, N2024);
xor XOR2 (N4521, N4496, N1009);
and AND3 (N4522, N4512, N4178, N2386);
and AND3 (N4523, N4521, N1221, N718);
not NOT1 (N4524, N4519);
nand NAND2 (N4525, N4523, N2030);
nand NAND2 (N4526, N4524, N4366);
or OR4 (N4527, N4525, N1767, N2184, N2560);
nor NOR3 (N4528, N4526, N3400, N2188);
xor XOR2 (N4529, N4507, N3087);
not NOT1 (N4530, N4494);
or OR2 (N4531, N4516, N650);
xor XOR2 (N4532, N4510, N4042);
and AND2 (N4533, N4520, N1332);
buf BUF1 (N4534, N4533);
xor XOR2 (N4535, N4530, N2588);
and AND3 (N4536, N4522, N1644, N4182);
and AND3 (N4537, N4535, N42, N1034);
and AND2 (N4538, N4517, N870);
buf BUF1 (N4539, N4527);
or OR3 (N4540, N4529, N3455, N3520);
xor XOR2 (N4541, N4532, N2340);
not NOT1 (N4542, N4537);
xor XOR2 (N4543, N4536, N4138);
or OR4 (N4544, N4539, N3895, N906, N1368);
not NOT1 (N4545, N4538);
xor XOR2 (N4546, N4531, N2697);
and AND2 (N4547, N4541, N4410);
xor XOR2 (N4548, N4547, N4105);
buf BUF1 (N4549, N4543);
or OR4 (N4550, N4544, N3883, N2130, N307);
and AND4 (N4551, N4542, N3701, N3266, N4467);
and AND2 (N4552, N4515, N247);
buf BUF1 (N4553, N4552);
buf BUF1 (N4554, N4553);
nor NOR3 (N4555, N4528, N1143, N3095);
and AND4 (N4556, N4545, N3869, N3104, N850);
nand NAND2 (N4557, N4549, N1401);
nand NAND2 (N4558, N4540, N1254);
nand NAND3 (N4559, N4555, N2715, N1013);
not NOT1 (N4560, N4557);
not NOT1 (N4561, N4534);
not NOT1 (N4562, N4546);
nand NAND2 (N4563, N4559, N1270);
nor NOR2 (N4564, N4558, N667);
nand NAND4 (N4565, N4562, N3238, N3226, N1263);
nor NOR3 (N4566, N4551, N234, N500);
nor NOR2 (N4567, N4550, N914);
buf BUF1 (N4568, N4563);
xor XOR2 (N4569, N4566, N1335);
nand NAND2 (N4570, N4560, N415);
nor NOR4 (N4571, N4569, N814, N4237, N2937);
nand NAND4 (N4572, N4564, N4313, N886, N4546);
or OR3 (N4573, N4565, N1968, N2014);
not NOT1 (N4574, N4548);
not NOT1 (N4575, N4556);
buf BUF1 (N4576, N4554);
buf BUF1 (N4577, N4573);
and AND4 (N4578, N4574, N4163, N27, N505);
and AND2 (N4579, N4567, N640);
or OR2 (N4580, N4579, N3648);
or OR4 (N4581, N4580, N4026, N2331, N4080);
not NOT1 (N4582, N4572);
buf BUF1 (N4583, N4578);
not NOT1 (N4584, N4575);
xor XOR2 (N4585, N4568, N1776);
xor XOR2 (N4586, N4585, N2162);
xor XOR2 (N4587, N4561, N4180);
nand NAND4 (N4588, N4584, N3526, N3532, N1037);
xor XOR2 (N4589, N4582, N3802);
nand NAND3 (N4590, N4571, N2694, N1667);
nor NOR2 (N4591, N4583, N269);
xor XOR2 (N4592, N4570, N2818);
nand NAND2 (N4593, N4581, N463);
nand NAND4 (N4594, N4587, N3204, N4496, N2795);
or OR2 (N4595, N4589, N1589);
buf BUF1 (N4596, N4588);
nand NAND4 (N4597, N4596, N821, N2981, N2047);
nor NOR3 (N4598, N4594, N332, N679);
not NOT1 (N4599, N4590);
and AND2 (N4600, N4598, N2854);
buf BUF1 (N4601, N4592);
buf BUF1 (N4602, N4600);
xor XOR2 (N4603, N4586, N1879);
buf BUF1 (N4604, N4593);
and AND4 (N4605, N4603, N1144, N2091, N1395);
not NOT1 (N4606, N4577);
or OR2 (N4607, N4599, N956);
not NOT1 (N4608, N4607);
and AND2 (N4609, N4604, N3482);
xor XOR2 (N4610, N4605, N220);
or OR2 (N4611, N4576, N406);
xor XOR2 (N4612, N4602, N2616);
nand NAND4 (N4613, N4595, N2256, N288, N4449);
not NOT1 (N4614, N4591);
xor XOR2 (N4615, N4601, N3649);
xor XOR2 (N4616, N4614, N785);
not NOT1 (N4617, N4615);
nor NOR4 (N4618, N4612, N553, N1935, N4611);
not NOT1 (N4619, N2232);
buf BUF1 (N4620, N4597);
nand NAND4 (N4621, N4620, N3262, N3775, N2818);
xor XOR2 (N4622, N4616, N241);
buf BUF1 (N4623, N4622);
nand NAND2 (N4624, N4621, N3523);
nor NOR4 (N4625, N4606, N2651, N2182, N3210);
or OR3 (N4626, N4613, N2184, N3710);
and AND4 (N4627, N4609, N2122, N4005, N2397);
buf BUF1 (N4628, N4623);
nor NOR3 (N4629, N4619, N3930, N2095);
not NOT1 (N4630, N4610);
buf BUF1 (N4631, N4627);
nand NAND3 (N4632, N4630, N642, N3558);
buf BUF1 (N4633, N4624);
or OR3 (N4634, N4632, N277, N4234);
and AND4 (N4635, N4626, N3070, N1536, N36);
nor NOR3 (N4636, N4618, N2408, N1843);
not NOT1 (N4637, N4633);
and AND4 (N4638, N4631, N1374, N2900, N319);
nor NOR4 (N4639, N4637, N104, N1040, N703);
xor XOR2 (N4640, N4608, N383);
or OR4 (N4641, N4629, N608, N2475, N3325);
not NOT1 (N4642, N4641);
nand NAND2 (N4643, N4638, N4498);
or OR4 (N4644, N4634, N4447, N1706, N936);
nand NAND3 (N4645, N4635, N3514, N1230);
and AND3 (N4646, N4640, N3408, N2493);
nand NAND4 (N4647, N4625, N1264, N4, N2546);
or OR2 (N4648, N4643, N4053);
buf BUF1 (N4649, N4642);
and AND3 (N4650, N4644, N2898, N3421);
xor XOR2 (N4651, N4649, N1453);
nor NOR2 (N4652, N4650, N2271);
nor NOR4 (N4653, N4639, N3086, N615, N3431);
nand NAND2 (N4654, N4648, N3553);
not NOT1 (N4655, N4653);
xor XOR2 (N4656, N4647, N1548);
or OR3 (N4657, N4628, N7, N811);
not NOT1 (N4658, N4646);
or OR4 (N4659, N4617, N3373, N1492, N4475);
nand NAND3 (N4660, N4636, N725, N1558);
or OR3 (N4661, N4655, N3734, N4080);
buf BUF1 (N4662, N4645);
or OR2 (N4663, N4657, N4457);
buf BUF1 (N4664, N4656);
or OR3 (N4665, N4652, N1895, N2257);
nor NOR4 (N4666, N4660, N2947, N764, N608);
nor NOR4 (N4667, N4665, N838, N2771, N2496);
xor XOR2 (N4668, N4667, N2641);
buf BUF1 (N4669, N4662);
xor XOR2 (N4670, N4651, N314);
xor XOR2 (N4671, N4664, N1002);
and AND2 (N4672, N4666, N1934);
xor XOR2 (N4673, N4663, N4648);
nand NAND4 (N4674, N4672, N1961, N4518, N3464);
nand NAND4 (N4675, N4654, N1812, N1585, N2534);
nor NOR2 (N4676, N4659, N1749);
nor NOR3 (N4677, N4669, N386, N1880);
and AND4 (N4678, N4661, N4610, N3274, N2175);
xor XOR2 (N4679, N4678, N2047);
and AND4 (N4680, N4658, N3622, N3348, N618);
xor XOR2 (N4681, N4675, N874);
buf BUF1 (N4682, N4677);
or OR2 (N4683, N4674, N2490);
nor NOR3 (N4684, N4681, N4669, N143);
xor XOR2 (N4685, N4683, N4460);
nor NOR2 (N4686, N4682, N1178);
buf BUF1 (N4687, N4684);
nor NOR3 (N4688, N4679, N732, N828);
nand NAND3 (N4689, N4680, N3515, N3190);
xor XOR2 (N4690, N4687, N374);
buf BUF1 (N4691, N4689);
not NOT1 (N4692, N4671);
and AND2 (N4693, N4690, N3858);
nor NOR2 (N4694, N4670, N255);
buf BUF1 (N4695, N4685);
and AND4 (N4696, N4692, N204, N2059, N3649);
nand NAND2 (N4697, N4676, N4415);
nor NOR4 (N4698, N4668, N1979, N3335, N3699);
not NOT1 (N4699, N4698);
not NOT1 (N4700, N4688);
not NOT1 (N4701, N4700);
or OR2 (N4702, N4701, N4328);
xor XOR2 (N4703, N4693, N153);
and AND4 (N4704, N4686, N3885, N717, N1835);
or OR3 (N4705, N4704, N3619, N3355);
not NOT1 (N4706, N4699);
nand NAND3 (N4707, N4705, N2904, N2470);
buf BUF1 (N4708, N4695);
nand NAND3 (N4709, N4691, N1851, N131);
buf BUF1 (N4710, N4694);
nor NOR2 (N4711, N4702, N178);
nand NAND2 (N4712, N4697, N3112);
nand NAND4 (N4713, N4710, N4648, N2815, N413);
nor NOR2 (N4714, N4713, N4412);
and AND3 (N4715, N4714, N903, N2863);
and AND2 (N4716, N4703, N3606);
not NOT1 (N4717, N4707);
not NOT1 (N4718, N4716);
or OR4 (N4719, N4712, N2079, N1610, N46);
and AND4 (N4720, N4717, N7, N1985, N2145);
buf BUF1 (N4721, N4719);
and AND2 (N4722, N4720, N3509);
and AND2 (N4723, N4673, N3927);
xor XOR2 (N4724, N4709, N4522);
and AND3 (N4725, N4722, N245, N2796);
or OR2 (N4726, N4715, N2041);
xor XOR2 (N4727, N4706, N917);
or OR4 (N4728, N4708, N2225, N1203, N116);
nor NOR2 (N4729, N4726, N3608);
and AND4 (N4730, N4696, N4713, N664, N2451);
nand NAND2 (N4731, N4727, N4005);
buf BUF1 (N4732, N4728);
buf BUF1 (N4733, N4730);
xor XOR2 (N4734, N4729, N2117);
nor NOR3 (N4735, N4725, N1599, N183);
not NOT1 (N4736, N4734);
and AND3 (N4737, N4723, N1325, N268);
or OR4 (N4738, N4731, N3649, N1193, N4512);
nand NAND3 (N4739, N4711, N4622, N2126);
xor XOR2 (N4740, N4718, N2243);
xor XOR2 (N4741, N4739, N3282);
buf BUF1 (N4742, N4733);
xor XOR2 (N4743, N4732, N2249);
nor NOR2 (N4744, N4743, N1018);
nor NOR2 (N4745, N4735, N3037);
nor NOR3 (N4746, N4742, N2939, N4656);
buf BUF1 (N4747, N4744);
not NOT1 (N4748, N4741);
nand NAND4 (N4749, N4737, N2081, N2360, N1826);
and AND4 (N4750, N4724, N2553, N1726, N2156);
not NOT1 (N4751, N4749);
not NOT1 (N4752, N4738);
nand NAND3 (N4753, N4750, N4385, N2359);
nand NAND3 (N4754, N4721, N572, N3895);
nor NOR2 (N4755, N4746, N3324);
nor NOR4 (N4756, N4753, N2047, N3220, N1225);
and AND3 (N4757, N4736, N3934, N804);
nand NAND3 (N4758, N4754, N2612, N1137);
nor NOR4 (N4759, N4740, N4450, N2301, N2754);
xor XOR2 (N4760, N4747, N4259);
and AND2 (N4761, N4751, N2504);
and AND2 (N4762, N4748, N3407);
xor XOR2 (N4763, N4755, N864);
nand NAND2 (N4764, N4752, N4339);
buf BUF1 (N4765, N4757);
buf BUF1 (N4766, N4764);
xor XOR2 (N4767, N4765, N2747);
and AND3 (N4768, N4756, N4586, N601);
and AND3 (N4769, N4763, N1971, N2481);
buf BUF1 (N4770, N4767);
xor XOR2 (N4771, N4760, N3643);
buf BUF1 (N4772, N4758);
nand NAND3 (N4773, N4768, N1526, N3907);
nor NOR4 (N4774, N4769, N1549, N4496, N3204);
and AND4 (N4775, N4771, N1883, N2485, N240);
not NOT1 (N4776, N4773);
buf BUF1 (N4777, N4775);
buf BUF1 (N4778, N4745);
buf BUF1 (N4779, N4770);
nand NAND3 (N4780, N4778, N634, N2921);
nor NOR3 (N4781, N4762, N1551, N2928);
nor NOR2 (N4782, N4777, N2124);
not NOT1 (N4783, N4774);
or OR4 (N4784, N4772, N2309, N434, N976);
xor XOR2 (N4785, N4776, N360);
nor NOR4 (N4786, N4784, N455, N1701, N403);
or OR2 (N4787, N4785, N1046);
nor NOR4 (N4788, N4766, N4272, N4762, N2717);
nand NAND4 (N4789, N4779, N1270, N885, N327);
buf BUF1 (N4790, N4761);
nand NAND3 (N4791, N4782, N4727, N972);
xor XOR2 (N4792, N4790, N3079);
xor XOR2 (N4793, N4791, N2298);
buf BUF1 (N4794, N4781);
xor XOR2 (N4795, N4793, N2906);
not NOT1 (N4796, N4759);
not NOT1 (N4797, N4787);
nand NAND2 (N4798, N4788, N3624);
or OR3 (N4799, N4792, N4221, N3212);
or OR4 (N4800, N4786, N3609, N1164, N4433);
not NOT1 (N4801, N4797);
nand NAND3 (N4802, N4783, N2480, N2291);
nand NAND2 (N4803, N4780, N4566);
or OR4 (N4804, N4795, N2117, N82, N1732);
buf BUF1 (N4805, N4803);
not NOT1 (N4806, N4796);
buf BUF1 (N4807, N4801);
buf BUF1 (N4808, N4789);
buf BUF1 (N4809, N4798);
nand NAND2 (N4810, N4799, N2416);
or OR3 (N4811, N4794, N3202, N735);
and AND4 (N4812, N4810, N462, N3527, N3269);
not NOT1 (N4813, N4806);
xor XOR2 (N4814, N4808, N2246);
or OR2 (N4815, N4805, N4441);
nand NAND3 (N4816, N4800, N471, N1880);
xor XOR2 (N4817, N4811, N2968);
nand NAND3 (N4818, N4804, N336, N4280);
or OR2 (N4819, N4802, N2643);
or OR3 (N4820, N4818, N1580, N126);
nor NOR4 (N4821, N4809, N4070, N154, N831);
or OR2 (N4822, N4813, N2080);
buf BUF1 (N4823, N4822);
not NOT1 (N4824, N4812);
nand NAND2 (N4825, N4816, N739);
or OR4 (N4826, N4807, N3748, N2895, N1503);
xor XOR2 (N4827, N4814, N2873);
not NOT1 (N4828, N4820);
not NOT1 (N4829, N4823);
nand NAND3 (N4830, N4828, N1571, N1397);
nor NOR4 (N4831, N4819, N540, N4653, N1944);
xor XOR2 (N4832, N4830, N3724);
or OR4 (N4833, N4829, N4431, N813, N159);
xor XOR2 (N4834, N4815, N3455);
or OR2 (N4835, N4833, N882);
nor NOR4 (N4836, N4821, N4368, N2534, N1849);
not NOT1 (N4837, N4834);
and AND3 (N4838, N4825, N4544, N2867);
nor NOR2 (N4839, N4836, N1442);
not NOT1 (N4840, N4839);
and AND2 (N4841, N4838, N598);
not NOT1 (N4842, N4824);
xor XOR2 (N4843, N4831, N3429);
nor NOR3 (N4844, N4827, N1168, N907);
nor NOR4 (N4845, N4837, N3395, N3900, N1423);
and AND2 (N4846, N4817, N2662);
not NOT1 (N4847, N4844);
or OR3 (N4848, N4832, N2864, N93);
or OR4 (N4849, N4841, N1418, N523, N2892);
nor NOR2 (N4850, N4846, N430);
and AND4 (N4851, N4826, N4365, N4678, N1180);
xor XOR2 (N4852, N4843, N4156);
nand NAND2 (N4853, N4850, N3061);
and AND2 (N4854, N4835, N1488);
or OR3 (N4855, N4845, N1531, N3232);
nand NAND3 (N4856, N4853, N3286, N3412);
nand NAND3 (N4857, N4847, N1938, N1405);
xor XOR2 (N4858, N4851, N3630);
not NOT1 (N4859, N4840);
and AND4 (N4860, N4848, N600, N955, N2041);
nand NAND3 (N4861, N4855, N3819, N2199);
not NOT1 (N4862, N4842);
nor NOR4 (N4863, N4858, N2608, N127, N3758);
and AND2 (N4864, N4856, N3086);
not NOT1 (N4865, N4859);
buf BUF1 (N4866, N4864);
or OR3 (N4867, N4861, N3154, N3739);
and AND4 (N4868, N4860, N944, N2796, N3189);
nor NOR2 (N4869, N4849, N1237);
not NOT1 (N4870, N4854);
nor NOR4 (N4871, N4865, N1312, N3265, N535);
nand NAND2 (N4872, N4857, N3052);
and AND4 (N4873, N4870, N3610, N2030, N1961);
and AND3 (N4874, N4863, N4820, N125);
xor XOR2 (N4875, N4866, N420);
nand NAND4 (N4876, N4875, N928, N1166, N806);
buf BUF1 (N4877, N4867);
nor NOR4 (N4878, N4852, N3347, N2160, N4489);
or OR4 (N4879, N4877, N2575, N1494, N3050);
nor NOR3 (N4880, N4874, N1700, N1553);
xor XOR2 (N4881, N4880, N337);
nand NAND4 (N4882, N4868, N3321, N3720, N1509);
not NOT1 (N4883, N4882);
buf BUF1 (N4884, N4872);
or OR3 (N4885, N4884, N1502, N2668);
nand NAND4 (N4886, N4883, N3945, N2740, N4264);
or OR2 (N4887, N4886, N570);
buf BUF1 (N4888, N4878);
nand NAND4 (N4889, N4888, N4243, N1923, N3317);
and AND4 (N4890, N4879, N677, N4121, N2148);
and AND3 (N4891, N4862, N929, N3844);
xor XOR2 (N4892, N4891, N539);
or OR4 (N4893, N4873, N2776, N3465, N3183);
nand NAND2 (N4894, N4893, N1832);
and AND2 (N4895, N4890, N2620);
nor NOR2 (N4896, N4892, N3897);
or OR3 (N4897, N4871, N4123, N2119);
not NOT1 (N4898, N4897);
buf BUF1 (N4899, N4889);
nand NAND2 (N4900, N4895, N2900);
xor XOR2 (N4901, N4898, N3599);
xor XOR2 (N4902, N4896, N924);
buf BUF1 (N4903, N4902);
buf BUF1 (N4904, N4887);
nand NAND3 (N4905, N4901, N526, N3460);
or OR2 (N4906, N4869, N3998);
xor XOR2 (N4907, N4885, N4215);
and AND4 (N4908, N4903, N2687, N2451, N3730);
nand NAND4 (N4909, N4906, N177, N2616, N3097);
buf BUF1 (N4910, N4904);
nor NOR3 (N4911, N4876, N1287, N4158);
or OR3 (N4912, N4905, N2638, N1331);
buf BUF1 (N4913, N4909);
xor XOR2 (N4914, N4899, N2914);
nand NAND2 (N4915, N4907, N989);
buf BUF1 (N4916, N4912);
nor NOR3 (N4917, N4916, N282, N4615);
not NOT1 (N4918, N4917);
not NOT1 (N4919, N4894);
not NOT1 (N4920, N4915);
nor NOR2 (N4921, N4900, N2365);
not NOT1 (N4922, N4919);
xor XOR2 (N4923, N4921, N3493);
not NOT1 (N4924, N4881);
buf BUF1 (N4925, N4908);
buf BUF1 (N4926, N4914);
not NOT1 (N4927, N4913);
buf BUF1 (N4928, N4926);
or OR3 (N4929, N4927, N829, N3237);
and AND2 (N4930, N4925, N2308);
or OR3 (N4931, N4928, N2041, N914);
buf BUF1 (N4932, N4931);
buf BUF1 (N4933, N4924);
buf BUF1 (N4934, N4911);
buf BUF1 (N4935, N4920);
buf BUF1 (N4936, N4933);
nor NOR4 (N4937, N4922, N992, N1293, N2333);
not NOT1 (N4938, N4934);
or OR2 (N4939, N4932, N1632);
not NOT1 (N4940, N4936);
nor NOR3 (N4941, N4940, N3771, N3568);
nand NAND3 (N4942, N4910, N1483, N3015);
xor XOR2 (N4943, N4941, N1477);
not NOT1 (N4944, N4938);
nor NOR3 (N4945, N4930, N4702, N439);
and AND3 (N4946, N4929, N1064, N1585);
not NOT1 (N4947, N4939);
nor NOR3 (N4948, N4918, N2612, N1318);
nand NAND4 (N4949, N4946, N2400, N993, N1694);
nand NAND3 (N4950, N4947, N4754, N1501);
nand NAND4 (N4951, N4942, N4472, N2678, N2235);
or OR4 (N4952, N4950, N272, N1852, N3088);
xor XOR2 (N4953, N4935, N74);
nand NAND2 (N4954, N4943, N628);
and AND3 (N4955, N4948, N2248, N233);
nand NAND4 (N4956, N4937, N2513, N4110, N4108);
and AND4 (N4957, N4955, N2694, N4278, N2093);
nand NAND3 (N4958, N4957, N198, N2306);
nor NOR2 (N4959, N4923, N1187);
nor NOR3 (N4960, N4958, N1683, N3664);
nor NOR2 (N4961, N4945, N2709);
nand NAND2 (N4962, N4961, N4205);
nor NOR4 (N4963, N4962, N4861, N3277, N3840);
xor XOR2 (N4964, N4953, N2781);
or OR4 (N4965, N4954, N548, N3422, N3376);
and AND2 (N4966, N4951, N3474);
or OR4 (N4967, N4952, N1297, N965, N3068);
not NOT1 (N4968, N4966);
xor XOR2 (N4969, N4949, N2637);
not NOT1 (N4970, N4967);
nand NAND3 (N4971, N4960, N4563, N2548);
nor NOR4 (N4972, N4944, N718, N1298, N2474);
buf BUF1 (N4973, N4968);
not NOT1 (N4974, N4956);
and AND2 (N4975, N4964, N4526);
or OR3 (N4976, N4965, N1760, N2751);
and AND3 (N4977, N4973, N394, N308);
nand NAND3 (N4978, N4977, N871, N720);
or OR3 (N4979, N4974, N4337, N557);
nor NOR4 (N4980, N4969, N2494, N1703, N1821);
buf BUF1 (N4981, N4971);
or OR2 (N4982, N4981, N3051);
not NOT1 (N4983, N4975);
nand NAND4 (N4984, N4980, N4820, N4648, N4612);
or OR3 (N4985, N4972, N3298, N2012);
or OR3 (N4986, N4979, N361, N1932);
and AND2 (N4987, N4976, N2444);
nor NOR4 (N4988, N4984, N2987, N945, N82);
not NOT1 (N4989, N4959);
and AND2 (N4990, N4986, N1850);
and AND3 (N4991, N4987, N456, N4799);
buf BUF1 (N4992, N4978);
xor XOR2 (N4993, N4992, N136);
buf BUF1 (N4994, N4993);
nand NAND2 (N4995, N4985, N4962);
buf BUF1 (N4996, N4988);
buf BUF1 (N4997, N4982);
nor NOR4 (N4998, N4989, N781, N1613, N615);
not NOT1 (N4999, N4983);
xor XOR2 (N5000, N4995, N2005);
buf BUF1 (N5001, N4997);
not NOT1 (N5002, N4991);
or OR4 (N5003, N4998, N2823, N1779, N4777);
nand NAND3 (N5004, N4994, N2278, N3310);
buf BUF1 (N5005, N4963);
and AND3 (N5006, N5005, N173, N1115);
not NOT1 (N5007, N4999);
nand NAND2 (N5008, N5006, N1124);
and AND3 (N5009, N4970, N3794, N3771);
buf BUF1 (N5010, N5007);
xor XOR2 (N5011, N5009, N1944);
nand NAND4 (N5012, N5003, N1593, N699, N225);
nor NOR2 (N5013, N5011, N2497);
not NOT1 (N5014, N5012);
buf BUF1 (N5015, N5004);
buf BUF1 (N5016, N5014);
nor NOR2 (N5017, N5016, N263);
buf BUF1 (N5018, N5013);
not NOT1 (N5019, N4990);
and AND3 (N5020, N5002, N1725, N450);
xor XOR2 (N5021, N5020, N2331);
nand NAND3 (N5022, N5018, N2277, N4279);
and AND2 (N5023, N5008, N1891);
xor XOR2 (N5024, N5017, N1986);
and AND4 (N5025, N5023, N4359, N3163, N4243);
not NOT1 (N5026, N5000);
and AND3 (N5027, N5001, N1012, N4343);
buf BUF1 (N5028, N5027);
nand NAND4 (N5029, N5026, N4855, N2630, N1700);
or OR3 (N5030, N5015, N1172, N1104);
buf BUF1 (N5031, N5022);
buf BUF1 (N5032, N5029);
xor XOR2 (N5033, N5032, N189);
or OR4 (N5034, N5025, N4208, N2454, N1415);
or OR2 (N5035, N5030, N1570);
or OR4 (N5036, N4996, N2944, N1328, N3135);
and AND4 (N5037, N5033, N3891, N3016, N3854);
not NOT1 (N5038, N5019);
buf BUF1 (N5039, N5037);
and AND3 (N5040, N5035, N4472, N2878);
nor NOR4 (N5041, N5021, N3400, N1731, N302);
and AND2 (N5042, N5028, N1519);
nor NOR4 (N5043, N5039, N520, N17, N3059);
and AND4 (N5044, N5024, N1345, N188, N278);
xor XOR2 (N5045, N5034, N3174);
nor NOR2 (N5046, N5038, N97);
not NOT1 (N5047, N5010);
buf BUF1 (N5048, N5040);
or OR4 (N5049, N5044, N3161, N1350, N4500);
xor XOR2 (N5050, N5041, N3462);
or OR2 (N5051, N5042, N3478);
nor NOR2 (N5052, N5049, N4763);
xor XOR2 (N5053, N5050, N4177);
and AND4 (N5054, N5036, N2059, N3880, N2561);
buf BUF1 (N5055, N5046);
not NOT1 (N5056, N5031);
nand NAND2 (N5057, N5045, N2332);
not NOT1 (N5058, N5043);
nand NAND3 (N5059, N5055, N95, N1477);
and AND4 (N5060, N5048, N2035, N2389, N4935);
nor NOR2 (N5061, N5047, N816);
xor XOR2 (N5062, N5054, N1557);
and AND2 (N5063, N5061, N4047);
and AND2 (N5064, N5053, N4768);
buf BUF1 (N5065, N5062);
nor NOR2 (N5066, N5065, N2756);
xor XOR2 (N5067, N5059, N4610);
or OR2 (N5068, N5064, N568);
buf BUF1 (N5069, N5051);
buf BUF1 (N5070, N5058);
and AND3 (N5071, N5060, N1929, N1625);
nand NAND3 (N5072, N5063, N201, N457);
nand NAND2 (N5073, N5069, N135);
or OR2 (N5074, N5052, N2562);
or OR2 (N5075, N5066, N1791);
and AND3 (N5076, N5067, N1934, N3099);
buf BUF1 (N5077, N5070);
and AND4 (N5078, N5077, N2415, N2686, N2517);
not NOT1 (N5079, N5057);
not NOT1 (N5080, N5073);
not NOT1 (N5081, N5074);
buf BUF1 (N5082, N5080);
buf BUF1 (N5083, N5078);
not NOT1 (N5084, N5071);
nor NOR2 (N5085, N5081, N2789);
not NOT1 (N5086, N5075);
buf BUF1 (N5087, N5056);
or OR4 (N5088, N5072, N2271, N1754, N3888);
xor XOR2 (N5089, N5084, N352);
or OR2 (N5090, N5083, N980);
buf BUF1 (N5091, N5085);
xor XOR2 (N5092, N5086, N2577);
nand NAND4 (N5093, N5091, N3194, N4023, N815);
or OR4 (N5094, N5092, N2439, N4663, N1198);
nor NOR4 (N5095, N5090, N1237, N2615, N4246);
buf BUF1 (N5096, N5093);
or OR3 (N5097, N5088, N379, N651);
buf BUF1 (N5098, N5082);
nor NOR3 (N5099, N5076, N3049, N2907);
or OR2 (N5100, N5098, N1988);
nor NOR4 (N5101, N5079, N4468, N1566, N3840);
not NOT1 (N5102, N5100);
buf BUF1 (N5103, N5102);
not NOT1 (N5104, N5103);
nor NOR2 (N5105, N5087, N3433);
not NOT1 (N5106, N5068);
and AND2 (N5107, N5099, N2969);
buf BUF1 (N5108, N5104);
nor NOR4 (N5109, N5101, N4843, N4343, N3872);
buf BUF1 (N5110, N5095);
xor XOR2 (N5111, N5097, N3954);
buf BUF1 (N5112, N5094);
xor XOR2 (N5113, N5107, N971);
nor NOR3 (N5114, N5105, N1834, N1694);
or OR2 (N5115, N5111, N1248);
not NOT1 (N5116, N5108);
nor NOR4 (N5117, N5109, N4065, N478, N2597);
buf BUF1 (N5118, N5115);
nor NOR2 (N5119, N5116, N1362);
and AND4 (N5120, N5119, N3687, N1375, N1485);
buf BUF1 (N5121, N5089);
nand NAND2 (N5122, N5113, N169);
not NOT1 (N5123, N5120);
nor NOR2 (N5124, N5118, N83);
not NOT1 (N5125, N5096);
nor NOR2 (N5126, N5121, N1554);
buf BUF1 (N5127, N5110);
not NOT1 (N5128, N5106);
xor XOR2 (N5129, N5126, N2581);
and AND3 (N5130, N5128, N2713, N608);
nor NOR4 (N5131, N5127, N1974, N3510, N274);
buf BUF1 (N5132, N5117);
nand NAND2 (N5133, N5123, N4272);
not NOT1 (N5134, N5131);
or OR2 (N5135, N5132, N1129);
nand NAND3 (N5136, N5134, N2254, N4301);
and AND4 (N5137, N5122, N3796, N4318, N348);
not NOT1 (N5138, N5130);
buf BUF1 (N5139, N5114);
xor XOR2 (N5140, N5136, N2072);
and AND2 (N5141, N5140, N3856);
or OR3 (N5142, N5129, N4235, N3088);
nor NOR4 (N5143, N5112, N224, N915, N3087);
xor XOR2 (N5144, N5137, N272);
not NOT1 (N5145, N5142);
xor XOR2 (N5146, N5144, N3291);
and AND4 (N5147, N5139, N2388, N3213, N712);
and AND4 (N5148, N5138, N2964, N3340, N3930);
xor XOR2 (N5149, N5141, N3114);
and AND2 (N5150, N5133, N2210);
nand NAND4 (N5151, N5148, N3190, N3563, N966);
nor NOR2 (N5152, N5150, N1084);
not NOT1 (N5153, N5149);
nor NOR3 (N5154, N5124, N3069, N1969);
nor NOR4 (N5155, N5135, N1659, N1385, N4927);
nand NAND3 (N5156, N5147, N3674, N2845);
nor NOR4 (N5157, N5146, N4845, N4997, N2245);
xor XOR2 (N5158, N5151, N4955);
not NOT1 (N5159, N5143);
or OR2 (N5160, N5157, N4122);
xor XOR2 (N5161, N5125, N4737);
nand NAND2 (N5162, N5152, N4175);
nand NAND2 (N5163, N5159, N3697);
xor XOR2 (N5164, N5161, N2300);
and AND2 (N5165, N5154, N2153);
xor XOR2 (N5166, N5145, N4397);
buf BUF1 (N5167, N5156);
nand NAND3 (N5168, N5165, N2090, N5161);
or OR4 (N5169, N5153, N1236, N3050, N1987);
and AND4 (N5170, N5164, N3363, N5129, N2602);
xor XOR2 (N5171, N5169, N3982);
nand NAND3 (N5172, N5166, N2899, N1119);
or OR2 (N5173, N5171, N1688);
and AND4 (N5174, N5158, N4093, N4604, N4426);
buf BUF1 (N5175, N5163);
and AND2 (N5176, N5172, N252);
not NOT1 (N5177, N5162);
nor NOR3 (N5178, N5167, N3281, N1337);
and AND3 (N5179, N5173, N4592, N2197);
or OR2 (N5180, N5178, N5081);
and AND4 (N5181, N5177, N3567, N2727, N1371);
nand NAND2 (N5182, N5176, N1028);
and AND3 (N5183, N5179, N1674, N4286);
not NOT1 (N5184, N5168);
and AND2 (N5185, N5155, N843);
nand NAND2 (N5186, N5175, N4664);
xor XOR2 (N5187, N5184, N3136);
nor NOR4 (N5188, N5187, N3957, N3878, N1406);
nand NAND3 (N5189, N5180, N2831, N3010);
not NOT1 (N5190, N5160);
nor NOR4 (N5191, N5182, N147, N373, N3186);
not NOT1 (N5192, N5189);
nor NOR2 (N5193, N5183, N1146);
and AND4 (N5194, N5188, N473, N1925, N3971);
or OR3 (N5195, N5194, N3799, N234);
buf BUF1 (N5196, N5181);
or OR3 (N5197, N5186, N4278, N4680);
not NOT1 (N5198, N5170);
xor XOR2 (N5199, N5174, N3847);
nor NOR2 (N5200, N5196, N4421);
not NOT1 (N5201, N5197);
buf BUF1 (N5202, N5199);
nor NOR3 (N5203, N5191, N1208, N188);
or OR2 (N5204, N5192, N824);
or OR4 (N5205, N5190, N3274, N2698, N1861);
nand NAND3 (N5206, N5203, N567, N4920);
nor NOR4 (N5207, N5201, N1269, N1900, N206);
xor XOR2 (N5208, N5185, N979);
nor NOR2 (N5209, N5193, N734);
buf BUF1 (N5210, N5198);
xor XOR2 (N5211, N5195, N3130);
not NOT1 (N5212, N5206);
nor NOR3 (N5213, N5200, N1297, N2053);
and AND4 (N5214, N5213, N4431, N824, N330);
xor XOR2 (N5215, N5207, N2480);
not NOT1 (N5216, N5208);
and AND3 (N5217, N5210, N1349, N4747);
xor XOR2 (N5218, N5214, N3016);
xor XOR2 (N5219, N5218, N2641);
not NOT1 (N5220, N5215);
and AND2 (N5221, N5216, N1682);
nand NAND3 (N5222, N5205, N747, N5128);
or OR2 (N5223, N5222, N380);
buf BUF1 (N5224, N5211);
buf BUF1 (N5225, N5217);
or OR4 (N5226, N5220, N1826, N3389, N2206);
nand NAND4 (N5227, N5204, N2570, N2424, N274);
and AND4 (N5228, N5225, N2943, N74, N3093);
or OR3 (N5229, N5227, N4115, N825);
nor NOR4 (N5230, N5209, N4940, N3343, N517);
nor NOR4 (N5231, N5202, N3441, N910, N1095);
nand NAND4 (N5232, N5219, N4966, N3266, N4391);
nand NAND2 (N5233, N5231, N5178);
or OR3 (N5234, N5229, N3216, N2115);
not NOT1 (N5235, N5223);
nor NOR4 (N5236, N5230, N1605, N1007, N3515);
xor XOR2 (N5237, N5234, N148);
nand NAND2 (N5238, N5237, N156);
nor NOR3 (N5239, N5232, N4097, N3185);
nor NOR2 (N5240, N5224, N3432);
nor NOR2 (N5241, N5238, N4955);
not NOT1 (N5242, N5233);
xor XOR2 (N5243, N5221, N2526);
buf BUF1 (N5244, N5239);
buf BUF1 (N5245, N5212);
or OR3 (N5246, N5228, N3514, N1217);
or OR3 (N5247, N5236, N4163, N2531);
not NOT1 (N5248, N5247);
nor NOR3 (N5249, N5226, N3194, N2076);
or OR2 (N5250, N5249, N2059);
xor XOR2 (N5251, N5235, N4755);
and AND2 (N5252, N5241, N3350);
or OR4 (N5253, N5244, N2470, N2729, N1634);
xor XOR2 (N5254, N5252, N2243);
nor NOR4 (N5255, N5242, N1036, N2230, N5039);
nor NOR3 (N5256, N5254, N3404, N1880);
nor NOR4 (N5257, N5253, N639, N4230, N2437);
nor NOR3 (N5258, N5240, N3640, N3736);
buf BUF1 (N5259, N5243);
nor NOR2 (N5260, N5250, N2808);
not NOT1 (N5261, N5251);
nor NOR2 (N5262, N5245, N4281);
nand NAND4 (N5263, N5262, N2942, N873, N5161);
xor XOR2 (N5264, N5248, N4627);
nor NOR2 (N5265, N5259, N1281);
and AND3 (N5266, N5264, N13, N2268);
buf BUF1 (N5267, N5257);
nand NAND3 (N5268, N5261, N1655, N1240);
xor XOR2 (N5269, N5268, N3285);
not NOT1 (N5270, N5265);
nor NOR2 (N5271, N5270, N4521);
buf BUF1 (N5272, N5263);
buf BUF1 (N5273, N5266);
nor NOR3 (N5274, N5269, N4644, N344);
nor NOR2 (N5275, N5256, N3055);
nand NAND3 (N5276, N5246, N449, N2161);
or OR3 (N5277, N5273, N2992, N958);
nand NAND3 (N5278, N5277, N1110, N1137);
not NOT1 (N5279, N5255);
xor XOR2 (N5280, N5267, N3996);
nor NOR4 (N5281, N5271, N3508, N430, N2743);
not NOT1 (N5282, N5280);
or OR3 (N5283, N5276, N290, N1160);
xor XOR2 (N5284, N5278, N1627);
or OR4 (N5285, N5283, N449, N163, N2404);
nand NAND4 (N5286, N5260, N672, N3900, N5108);
xor XOR2 (N5287, N5279, N2729);
xor XOR2 (N5288, N5272, N1741);
not NOT1 (N5289, N5281);
not NOT1 (N5290, N5258);
or OR2 (N5291, N5285, N4702);
and AND3 (N5292, N5282, N1315, N741);
not NOT1 (N5293, N5290);
or OR3 (N5294, N5293, N730, N3824);
nor NOR2 (N5295, N5284, N3811);
or OR3 (N5296, N5288, N4296, N4233);
xor XOR2 (N5297, N5289, N5031);
buf BUF1 (N5298, N5287);
nand NAND4 (N5299, N5298, N43, N1214, N1932);
nand NAND3 (N5300, N5292, N1093, N5135);
buf BUF1 (N5301, N5297);
not NOT1 (N5302, N5301);
and AND4 (N5303, N5294, N1122, N76, N876);
not NOT1 (N5304, N5295);
not NOT1 (N5305, N5275);
not NOT1 (N5306, N5296);
or OR2 (N5307, N5299, N2426);
xor XOR2 (N5308, N5291, N436);
or OR2 (N5309, N5303, N2609);
buf BUF1 (N5310, N5274);
or OR4 (N5311, N5304, N4542, N1753, N4325);
buf BUF1 (N5312, N5286);
and AND2 (N5313, N5302, N3130);
xor XOR2 (N5314, N5308, N4124);
xor XOR2 (N5315, N5312, N2372);
not NOT1 (N5316, N5300);
not NOT1 (N5317, N5310);
nand NAND3 (N5318, N5306, N1158, N3850);
and AND2 (N5319, N5314, N442);
xor XOR2 (N5320, N5317, N453);
or OR4 (N5321, N5307, N3530, N1921, N1511);
xor XOR2 (N5322, N5311, N1705);
xor XOR2 (N5323, N5316, N2977);
not NOT1 (N5324, N5315);
buf BUF1 (N5325, N5313);
not NOT1 (N5326, N5325);
nand NAND2 (N5327, N5321, N3774);
or OR3 (N5328, N5305, N554, N754);
xor XOR2 (N5329, N5309, N2775);
or OR3 (N5330, N5327, N2143, N2232);
nand NAND3 (N5331, N5326, N329, N3894);
and AND3 (N5332, N5320, N2673, N3473);
nand NAND4 (N5333, N5319, N282, N3960, N4584);
and AND4 (N5334, N5333, N964, N3921, N317);
or OR2 (N5335, N5330, N1197);
nand NAND4 (N5336, N5329, N1958, N2063, N3925);
and AND4 (N5337, N5336, N2109, N4139, N3594);
and AND4 (N5338, N5318, N1769, N1634, N1064);
and AND4 (N5339, N5337, N700, N1278, N3554);
nor NOR4 (N5340, N5334, N3567, N3311, N1026);
not NOT1 (N5341, N5322);
not NOT1 (N5342, N5339);
nand NAND3 (N5343, N5332, N2507, N2385);
nand NAND2 (N5344, N5323, N257);
xor XOR2 (N5345, N5324, N2547);
xor XOR2 (N5346, N5343, N3119);
and AND2 (N5347, N5345, N1217);
nor NOR3 (N5348, N5341, N1492, N321);
or OR3 (N5349, N5347, N3950, N5226);
buf BUF1 (N5350, N5349);
nand NAND2 (N5351, N5344, N3448);
buf BUF1 (N5352, N5328);
and AND4 (N5353, N5338, N1906, N3106, N4798);
nand NAND2 (N5354, N5348, N4);
xor XOR2 (N5355, N5346, N537);
or OR2 (N5356, N5342, N3359);
not NOT1 (N5357, N5335);
buf BUF1 (N5358, N5350);
and AND4 (N5359, N5331, N413, N2308, N2860);
nor NOR3 (N5360, N5359, N800, N1444);
and AND4 (N5361, N5354, N3423, N4182, N1089);
not NOT1 (N5362, N5352);
buf BUF1 (N5363, N5351);
or OR2 (N5364, N5356, N894);
or OR2 (N5365, N5353, N3520);
xor XOR2 (N5366, N5360, N2870);
nor NOR3 (N5367, N5357, N2373, N2727);
nor NOR2 (N5368, N5355, N838);
nor NOR2 (N5369, N5340, N410);
not NOT1 (N5370, N5364);
and AND3 (N5371, N5366, N3853, N4924);
nor NOR2 (N5372, N5365, N475);
not NOT1 (N5373, N5372);
nor NOR4 (N5374, N5368, N1055, N2839, N1564);
nor NOR4 (N5375, N5371, N3457, N4437, N4884);
or OR2 (N5376, N5373, N5271);
or OR2 (N5377, N5358, N4871);
and AND2 (N5378, N5370, N2375);
buf BUF1 (N5379, N5377);
or OR3 (N5380, N5369, N1478, N308);
xor XOR2 (N5381, N5363, N2532);
buf BUF1 (N5382, N5362);
buf BUF1 (N5383, N5382);
nand NAND4 (N5384, N5381, N3295, N513, N5368);
and AND4 (N5385, N5376, N1297, N1305, N3331);
nor NOR2 (N5386, N5385, N2676);
not NOT1 (N5387, N5386);
and AND4 (N5388, N5374, N681, N2994, N4869);
and AND2 (N5389, N5367, N1444);
not NOT1 (N5390, N5375);
xor XOR2 (N5391, N5383, N4102);
or OR4 (N5392, N5389, N5351, N4860, N119);
and AND4 (N5393, N5388, N835, N2617, N3586);
nor NOR4 (N5394, N5379, N757, N924, N3074);
buf BUF1 (N5395, N5393);
nand NAND3 (N5396, N5390, N1732, N2743);
or OR3 (N5397, N5394, N122, N2589);
not NOT1 (N5398, N5380);
or OR2 (N5399, N5391, N2192);
or OR2 (N5400, N5399, N4735);
or OR4 (N5401, N5400, N3261, N5173, N2876);
or OR4 (N5402, N5396, N5023, N28, N2708);
and AND4 (N5403, N5402, N1341, N521, N4574);
xor XOR2 (N5404, N5387, N1889);
not NOT1 (N5405, N5401);
nor NOR3 (N5406, N5398, N1876, N1128);
xor XOR2 (N5407, N5406, N3123);
xor XOR2 (N5408, N5405, N2247);
nor NOR3 (N5409, N5403, N4990, N4597);
nor NOR3 (N5410, N5408, N555, N2887);
xor XOR2 (N5411, N5407, N1397);
or OR4 (N5412, N5410, N333, N4757, N552);
buf BUF1 (N5413, N5411);
not NOT1 (N5414, N5397);
buf BUF1 (N5415, N5404);
buf BUF1 (N5416, N5414);
nor NOR3 (N5417, N5412, N4046, N3122);
and AND3 (N5418, N5395, N3604, N3469);
or OR4 (N5419, N5418, N1653, N2988, N4805);
buf BUF1 (N5420, N5415);
xor XOR2 (N5421, N5409, N1636);
buf BUF1 (N5422, N5419);
xor XOR2 (N5423, N5421, N3121);
or OR3 (N5424, N5422, N3869, N2468);
nor NOR2 (N5425, N5384, N444);
nor NOR2 (N5426, N5417, N3553);
and AND4 (N5427, N5423, N1462, N2221, N136);
not NOT1 (N5428, N5392);
or OR2 (N5429, N5413, N3496);
xor XOR2 (N5430, N5361, N380);
buf BUF1 (N5431, N5429);
or OR3 (N5432, N5430, N4902, N4856);
buf BUF1 (N5433, N5428);
not NOT1 (N5434, N5432);
buf BUF1 (N5435, N5424);
and AND4 (N5436, N5416, N1570, N5214, N263);
not NOT1 (N5437, N5427);
or OR3 (N5438, N5420, N5360, N4756);
and AND4 (N5439, N5434, N3731, N4071, N3592);
or OR4 (N5440, N5439, N2571, N1435, N448);
nor NOR2 (N5441, N5438, N1609);
nand NAND2 (N5442, N5436, N3311);
buf BUF1 (N5443, N5442);
xor XOR2 (N5444, N5443, N3220);
or OR2 (N5445, N5426, N1419);
or OR2 (N5446, N5441, N2503);
not NOT1 (N5447, N5440);
and AND2 (N5448, N5378, N2786);
nor NOR3 (N5449, N5425, N2299, N4888);
or OR4 (N5450, N5449, N936, N2537, N3517);
xor XOR2 (N5451, N5435, N935);
or OR4 (N5452, N5433, N3434, N4337, N3297);
xor XOR2 (N5453, N5437, N1459);
nor NOR2 (N5454, N5444, N5208);
xor XOR2 (N5455, N5450, N3138);
xor XOR2 (N5456, N5452, N3357);
and AND4 (N5457, N5445, N3234, N3284, N378);
or OR4 (N5458, N5453, N2338, N1126, N3689);
or OR4 (N5459, N5458, N3934, N3920, N4343);
xor XOR2 (N5460, N5448, N2901);
nand NAND2 (N5461, N5431, N2667);
buf BUF1 (N5462, N5454);
nor NOR2 (N5463, N5459, N2347);
not NOT1 (N5464, N5460);
or OR2 (N5465, N5455, N3831);
buf BUF1 (N5466, N5461);
nor NOR2 (N5467, N5447, N5240);
xor XOR2 (N5468, N5467, N1125);
buf BUF1 (N5469, N5466);
and AND4 (N5470, N5457, N4882, N399, N3892);
xor XOR2 (N5471, N5465, N3587);
xor XOR2 (N5472, N5456, N2810);
and AND3 (N5473, N5446, N2642, N632);
buf BUF1 (N5474, N5468);
not NOT1 (N5475, N5473);
and AND3 (N5476, N5471, N985, N3796);
nand NAND3 (N5477, N5469, N4014, N864);
nand NAND4 (N5478, N5451, N4118, N1294, N3092);
buf BUF1 (N5479, N5474);
nand NAND4 (N5480, N5462, N1745, N2495, N4373);
not NOT1 (N5481, N5470);
and AND4 (N5482, N5479, N108, N1, N1762);
nand NAND2 (N5483, N5477, N3081);
nand NAND4 (N5484, N5483, N2714, N4148, N160);
nand NAND3 (N5485, N5481, N4362, N571);
and AND2 (N5486, N5482, N3782);
and AND3 (N5487, N5472, N5069, N1839);
nand NAND3 (N5488, N5464, N3336, N2996);
buf BUF1 (N5489, N5478);
nor NOR2 (N5490, N5476, N1439);
or OR3 (N5491, N5475, N2396, N941);
xor XOR2 (N5492, N5480, N3383);
xor XOR2 (N5493, N5484, N240);
nor NOR3 (N5494, N5463, N5454, N4225);
nor NOR4 (N5495, N5487, N4874, N356, N608);
nand NAND3 (N5496, N5492, N4154, N5119);
buf BUF1 (N5497, N5485);
buf BUF1 (N5498, N5489);
xor XOR2 (N5499, N5493, N1306);
nor NOR2 (N5500, N5496, N408);
nand NAND3 (N5501, N5498, N4821, N362);
nand NAND3 (N5502, N5494, N1796, N3836);
and AND4 (N5503, N5491, N552, N1986, N2032);
not NOT1 (N5504, N5495);
buf BUF1 (N5505, N5503);
nor NOR3 (N5506, N5501, N589, N791);
nand NAND3 (N5507, N5505, N3010, N5343);
and AND3 (N5508, N5490, N5479, N5479);
buf BUF1 (N5509, N5506);
buf BUF1 (N5510, N5486);
or OR2 (N5511, N5508, N1231);
buf BUF1 (N5512, N5500);
not NOT1 (N5513, N5497);
buf BUF1 (N5514, N5512);
xor XOR2 (N5515, N5507, N246);
nor NOR3 (N5516, N5514, N4355, N1008);
buf BUF1 (N5517, N5509);
or OR3 (N5518, N5488, N4932, N3492);
buf BUF1 (N5519, N5511);
nor NOR2 (N5520, N5518, N3361);
not NOT1 (N5521, N5510);
and AND2 (N5522, N5499, N2024);
not NOT1 (N5523, N5513);
or OR2 (N5524, N5522, N3793);
buf BUF1 (N5525, N5519);
nand NAND4 (N5526, N5521, N5154, N1479, N4574);
nand NAND4 (N5527, N5504, N2828, N3440, N1888);
not NOT1 (N5528, N5517);
nor NOR4 (N5529, N5524, N3622, N4040, N1730);
xor XOR2 (N5530, N5515, N238);
buf BUF1 (N5531, N5530);
not NOT1 (N5532, N5523);
xor XOR2 (N5533, N5520, N2029);
xor XOR2 (N5534, N5532, N2568);
and AND3 (N5535, N5526, N1725, N4261);
nand NAND2 (N5536, N5531, N2525);
and AND2 (N5537, N5527, N163);
nor NOR4 (N5538, N5529, N3357, N912, N4404);
nand NAND2 (N5539, N5534, N1873);
not NOT1 (N5540, N5528);
or OR3 (N5541, N5516, N788, N4089);
nor NOR2 (N5542, N5536, N741);
nor NOR4 (N5543, N5537, N3568, N1633, N3648);
buf BUF1 (N5544, N5502);
nand NAND2 (N5545, N5540, N875);
nand NAND3 (N5546, N5525, N1827, N4177);
and AND3 (N5547, N5542, N994, N2774);
nor NOR2 (N5548, N5539, N1891);
xor XOR2 (N5549, N5546, N3113);
or OR4 (N5550, N5548, N2842, N2515, N1937);
nand NAND3 (N5551, N5545, N2317, N226);
nand NAND4 (N5552, N5535, N386, N4385, N4613);
or OR2 (N5553, N5541, N764);
nand NAND3 (N5554, N5533, N4694, N1964);
nand NAND3 (N5555, N5549, N4594, N3825);
buf BUF1 (N5556, N5555);
not NOT1 (N5557, N5556);
nor NOR4 (N5558, N5557, N536, N4498, N2143);
and AND4 (N5559, N5543, N1906, N734, N3688);
or OR2 (N5560, N5558, N3613);
xor XOR2 (N5561, N5552, N4654);
buf BUF1 (N5562, N5544);
nand NAND3 (N5563, N5547, N4740, N5254);
or OR2 (N5564, N5563, N1120);
xor XOR2 (N5565, N5564, N5159);
xor XOR2 (N5566, N5551, N3185);
and AND4 (N5567, N5538, N4239, N4403, N2714);
or OR4 (N5568, N5567, N5431, N4911, N5530);
not NOT1 (N5569, N5553);
and AND3 (N5570, N5566, N3863, N1899);
xor XOR2 (N5571, N5570, N2664);
not NOT1 (N5572, N5569);
or OR3 (N5573, N5568, N970, N1036);
nor NOR3 (N5574, N5573, N1024, N5347);
buf BUF1 (N5575, N5574);
xor XOR2 (N5576, N5550, N193);
nand NAND4 (N5577, N5572, N3171, N2276, N4649);
xor XOR2 (N5578, N5565, N2068);
not NOT1 (N5579, N5561);
nand NAND4 (N5580, N5560, N4321, N432, N1096);
buf BUF1 (N5581, N5562);
xor XOR2 (N5582, N5575, N36);
or OR3 (N5583, N5581, N620, N5375);
not NOT1 (N5584, N5580);
not NOT1 (N5585, N5559);
and AND4 (N5586, N5577, N298, N4070, N4759);
nor NOR2 (N5587, N5579, N1544);
xor XOR2 (N5588, N5583, N5312);
or OR4 (N5589, N5578, N1743, N3743, N194);
nor NOR4 (N5590, N5554, N1505, N819, N3977);
or OR2 (N5591, N5587, N5103);
buf BUF1 (N5592, N5589);
nor NOR3 (N5593, N5582, N3221, N2174);
xor XOR2 (N5594, N5591, N920);
buf BUF1 (N5595, N5592);
and AND4 (N5596, N5571, N1849, N2917, N4149);
and AND2 (N5597, N5585, N4708);
nor NOR2 (N5598, N5586, N1965);
xor XOR2 (N5599, N5594, N2548);
or OR3 (N5600, N5576, N84, N2951);
nor NOR2 (N5601, N5590, N1990);
and AND2 (N5602, N5593, N750);
nand NAND3 (N5603, N5595, N2857, N851);
and AND4 (N5604, N5603, N3582, N2180, N458);
nand NAND3 (N5605, N5601, N527, N3541);
nand NAND3 (N5606, N5600, N4068, N3757);
nor NOR2 (N5607, N5599, N2224);
nor NOR2 (N5608, N5602, N356);
nor NOR2 (N5609, N5596, N377);
xor XOR2 (N5610, N5597, N5063);
nand NAND4 (N5611, N5588, N2123, N5125, N2594);
and AND4 (N5612, N5604, N194, N4615, N2332);
and AND4 (N5613, N5612, N5130, N1460, N799);
nand NAND2 (N5614, N5607, N3793);
nand NAND4 (N5615, N5613, N296, N3480, N4507);
nand NAND2 (N5616, N5609, N4029);
or OR4 (N5617, N5598, N2952, N2361, N4202);
nor NOR3 (N5618, N5616, N453, N1681);
buf BUF1 (N5619, N5615);
xor XOR2 (N5620, N5614, N4386);
xor XOR2 (N5621, N5605, N2888);
nand NAND4 (N5622, N5584, N1538, N1844, N2587);
and AND3 (N5623, N5621, N1629, N4586);
and AND2 (N5624, N5617, N903);
not NOT1 (N5625, N5610);
not NOT1 (N5626, N5611);
nor NOR3 (N5627, N5624, N2919, N3364);
buf BUF1 (N5628, N5618);
nand NAND3 (N5629, N5626, N1208, N1393);
and AND2 (N5630, N5619, N5538);
or OR4 (N5631, N5627, N2785, N1255, N1328);
or OR3 (N5632, N5630, N5389, N1394);
not NOT1 (N5633, N5632);
buf BUF1 (N5634, N5628);
xor XOR2 (N5635, N5633, N5245);
and AND3 (N5636, N5606, N3348, N3779);
nand NAND3 (N5637, N5623, N4516, N5019);
buf BUF1 (N5638, N5636);
xor XOR2 (N5639, N5629, N3288);
or OR2 (N5640, N5620, N2651);
xor XOR2 (N5641, N5608, N4540);
not NOT1 (N5642, N5634);
not NOT1 (N5643, N5631);
nand NAND4 (N5644, N5637, N1063, N707, N959);
not NOT1 (N5645, N5639);
and AND2 (N5646, N5638, N4120);
not NOT1 (N5647, N5641);
buf BUF1 (N5648, N5622);
and AND3 (N5649, N5645, N4415, N2986);
not NOT1 (N5650, N5647);
or OR3 (N5651, N5649, N4074, N4608);
buf BUF1 (N5652, N5648);
nor NOR2 (N5653, N5643, N3099);
xor XOR2 (N5654, N5642, N4297);
buf BUF1 (N5655, N5651);
not NOT1 (N5656, N5646);
nand NAND2 (N5657, N5635, N2570);
and AND4 (N5658, N5625, N132, N2516, N2121);
xor XOR2 (N5659, N5653, N2820);
and AND3 (N5660, N5656, N3993, N417);
xor XOR2 (N5661, N5644, N2554);
nand NAND4 (N5662, N5657, N3883, N2182, N40);
nor NOR4 (N5663, N5659, N3641, N1715, N124);
nor NOR3 (N5664, N5654, N3638, N2225);
and AND2 (N5665, N5662, N315);
nor NOR3 (N5666, N5640, N2033, N1032);
and AND3 (N5667, N5658, N437, N711);
or OR4 (N5668, N5655, N2636, N5170, N1098);
or OR4 (N5669, N5650, N5294, N3377, N1945);
or OR2 (N5670, N5667, N833);
nor NOR3 (N5671, N5665, N3577, N121);
nand NAND4 (N5672, N5666, N4826, N163, N3287);
not NOT1 (N5673, N5664);
nor NOR2 (N5674, N5661, N60);
nand NAND2 (N5675, N5670, N161);
buf BUF1 (N5676, N5669);
xor XOR2 (N5677, N5672, N4397);
xor XOR2 (N5678, N5668, N1196);
nand NAND2 (N5679, N5678, N2134);
nand NAND4 (N5680, N5671, N843, N2368, N2839);
buf BUF1 (N5681, N5663);
and AND4 (N5682, N5676, N3343, N1721, N5214);
not NOT1 (N5683, N5679);
and AND2 (N5684, N5683, N3128);
nand NAND2 (N5685, N5684, N2566);
not NOT1 (N5686, N5680);
nor NOR4 (N5687, N5652, N872, N4205, N2669);
nand NAND3 (N5688, N5682, N464, N4404);
and AND3 (N5689, N5681, N2390, N4682);
nand NAND3 (N5690, N5689, N3419, N4538);
and AND2 (N5691, N5660, N1935);
nand NAND2 (N5692, N5673, N5608);
xor XOR2 (N5693, N5674, N4290);
nand NAND2 (N5694, N5688, N2241);
nand NAND4 (N5695, N5685, N4022, N3400, N930);
or OR3 (N5696, N5692, N2062, N4851);
nand NAND3 (N5697, N5690, N2646, N5607);
buf BUF1 (N5698, N5675);
not NOT1 (N5699, N5695);
or OR4 (N5700, N5699, N1441, N3779, N4609);
or OR4 (N5701, N5693, N5408, N2907, N3673);
xor XOR2 (N5702, N5691, N90);
nand NAND2 (N5703, N5677, N618);
not NOT1 (N5704, N5702);
nand NAND2 (N5705, N5687, N576);
and AND2 (N5706, N5686, N2325);
not NOT1 (N5707, N5706);
xor XOR2 (N5708, N5707, N4613);
nand NAND4 (N5709, N5698, N3011, N5193, N981);
or OR2 (N5710, N5701, N2414);
or OR3 (N5711, N5703, N5271, N2458);
nor NOR2 (N5712, N5709, N1315);
nand NAND3 (N5713, N5700, N1240, N97);
not NOT1 (N5714, N5708);
nor NOR4 (N5715, N5696, N409, N4109, N3564);
nand NAND3 (N5716, N5713, N3483, N5014);
or OR3 (N5717, N5710, N2634, N5585);
nand NAND2 (N5718, N5705, N625);
not NOT1 (N5719, N5704);
or OR2 (N5720, N5694, N3630);
buf BUF1 (N5721, N5697);
and AND2 (N5722, N5719, N5493);
nor NOR2 (N5723, N5720, N3519);
not NOT1 (N5724, N5718);
buf BUF1 (N5725, N5715);
or OR3 (N5726, N5725, N4811, N2866);
or OR3 (N5727, N5721, N3993, N3600);
nor NOR3 (N5728, N5711, N1764, N1462);
nor NOR3 (N5729, N5724, N4996, N975);
not NOT1 (N5730, N5717);
xor XOR2 (N5731, N5726, N1219);
or OR2 (N5732, N5730, N2075);
buf BUF1 (N5733, N5727);
nor NOR2 (N5734, N5733, N917);
not NOT1 (N5735, N5732);
nor NOR3 (N5736, N5731, N4546, N3115);
or OR2 (N5737, N5729, N1709);
xor XOR2 (N5738, N5723, N5442);
xor XOR2 (N5739, N5716, N2606);
nand NAND3 (N5740, N5735, N5703, N2382);
buf BUF1 (N5741, N5714);
nand NAND2 (N5742, N5741, N873);
or OR3 (N5743, N5736, N1333, N5464);
buf BUF1 (N5744, N5743);
xor XOR2 (N5745, N5738, N1816);
nand NAND2 (N5746, N5737, N5137);
xor XOR2 (N5747, N5712, N4707);
nand NAND2 (N5748, N5722, N1284);
and AND4 (N5749, N5742, N4522, N923, N4917);
buf BUF1 (N5750, N5728);
and AND4 (N5751, N5744, N1958, N2634, N5552);
nor NOR4 (N5752, N5739, N2654, N676, N3466);
nand NAND3 (N5753, N5747, N2657, N5057);
nand NAND4 (N5754, N5740, N89, N1978, N1250);
not NOT1 (N5755, N5746);
nor NOR2 (N5756, N5754, N4397);
not NOT1 (N5757, N5750);
and AND3 (N5758, N5753, N1053, N601);
nand NAND4 (N5759, N5758, N4120, N2008, N5447);
nor NOR3 (N5760, N5752, N4184, N5504);
not NOT1 (N5761, N5751);
or OR2 (N5762, N5749, N2599);
or OR4 (N5763, N5762, N1802, N2087, N3639);
xor XOR2 (N5764, N5761, N2700);
nand NAND3 (N5765, N5763, N1442, N3138);
not NOT1 (N5766, N5757);
nand NAND4 (N5767, N5760, N298, N5512, N2474);
nand NAND4 (N5768, N5767, N2456, N3818, N5160);
nand NAND2 (N5769, N5755, N1968);
nor NOR4 (N5770, N5756, N5221, N5180, N5325);
nand NAND2 (N5771, N5770, N2817);
not NOT1 (N5772, N5759);
not NOT1 (N5773, N5769);
buf BUF1 (N5774, N5771);
nor NOR2 (N5775, N5768, N4861);
buf BUF1 (N5776, N5766);
or OR2 (N5777, N5745, N1991);
not NOT1 (N5778, N5765);
nor NOR2 (N5779, N5773, N5120);
nor NOR3 (N5780, N5734, N3498, N3673);
buf BUF1 (N5781, N5764);
not NOT1 (N5782, N5780);
buf BUF1 (N5783, N5772);
nand NAND2 (N5784, N5783, N4457);
nand NAND3 (N5785, N5775, N3989, N3200);
nand NAND3 (N5786, N5778, N2429, N2983);
xor XOR2 (N5787, N5774, N4024);
nand NAND2 (N5788, N5779, N3346);
nor NOR2 (N5789, N5788, N1953);
buf BUF1 (N5790, N5787);
or OR3 (N5791, N5748, N777, N227);
nand NAND2 (N5792, N5790, N1450);
nor NOR2 (N5793, N5789, N924);
buf BUF1 (N5794, N5777);
not NOT1 (N5795, N5786);
buf BUF1 (N5796, N5792);
xor XOR2 (N5797, N5796, N5631);
not NOT1 (N5798, N5784);
not NOT1 (N5799, N5795);
nand NAND2 (N5800, N5799, N5126);
or OR3 (N5801, N5793, N2910, N4208);
xor XOR2 (N5802, N5801, N5441);
buf BUF1 (N5803, N5798);
nand NAND2 (N5804, N5803, N1168);
not NOT1 (N5805, N5802);
buf BUF1 (N5806, N5805);
and AND2 (N5807, N5806, N4015);
buf BUF1 (N5808, N5800);
buf BUF1 (N5809, N5804);
nand NAND4 (N5810, N5781, N233, N2747, N2924);
xor XOR2 (N5811, N5807, N5420);
nand NAND2 (N5812, N5809, N4087);
nor NOR3 (N5813, N5808, N832, N5007);
xor XOR2 (N5814, N5791, N4964);
buf BUF1 (N5815, N5794);
buf BUF1 (N5816, N5776);
not NOT1 (N5817, N5815);
buf BUF1 (N5818, N5811);
nand NAND4 (N5819, N5797, N1921, N1894, N2051);
or OR4 (N5820, N5814, N1831, N3569, N4968);
nand NAND2 (N5821, N5816, N39);
and AND2 (N5822, N5818, N2900);
and AND2 (N5823, N5782, N1624);
xor XOR2 (N5824, N5813, N153);
nand NAND3 (N5825, N5824, N2373, N4824);
buf BUF1 (N5826, N5819);
xor XOR2 (N5827, N5812, N1482);
nand NAND2 (N5828, N5821, N2742);
nand NAND2 (N5829, N5785, N4842);
nor NOR3 (N5830, N5825, N305, N1317);
buf BUF1 (N5831, N5828);
nor NOR2 (N5832, N5831, N1995);
not NOT1 (N5833, N5829);
nor NOR3 (N5834, N5827, N3820, N2869);
buf BUF1 (N5835, N5822);
not NOT1 (N5836, N5826);
nand NAND4 (N5837, N5823, N5556, N3206, N2783);
nand NAND2 (N5838, N5837, N4681);
not NOT1 (N5839, N5817);
not NOT1 (N5840, N5834);
or OR4 (N5841, N5832, N3203, N1241, N3281);
nand NAND2 (N5842, N5830, N5759);
or OR4 (N5843, N5842, N2576, N292, N2351);
or OR3 (N5844, N5838, N3795, N3408);
not NOT1 (N5845, N5844);
xor XOR2 (N5846, N5835, N5355);
and AND2 (N5847, N5839, N3618);
nor NOR4 (N5848, N5847, N5572, N2007, N2106);
nor NOR4 (N5849, N5820, N2617, N5030, N1112);
and AND2 (N5850, N5810, N5243);
xor XOR2 (N5851, N5840, N3913);
nand NAND2 (N5852, N5843, N1041);
nor NOR4 (N5853, N5845, N1219, N5111, N3864);
buf BUF1 (N5854, N5846);
not NOT1 (N5855, N5849);
and AND2 (N5856, N5850, N462);
and AND3 (N5857, N5854, N3803, N5493);
and AND4 (N5858, N5833, N5521, N4026, N5118);
buf BUF1 (N5859, N5858);
or OR3 (N5860, N5856, N1625, N4387);
buf BUF1 (N5861, N5848);
xor XOR2 (N5862, N5853, N2212);
buf BUF1 (N5863, N5836);
nand NAND4 (N5864, N5859, N4982, N763, N4900);
xor XOR2 (N5865, N5862, N4525);
or OR3 (N5866, N5855, N2530, N4597);
not NOT1 (N5867, N5866);
xor XOR2 (N5868, N5867, N5527);
xor XOR2 (N5869, N5860, N5676);
nand NAND2 (N5870, N5868, N5551);
buf BUF1 (N5871, N5863);
buf BUF1 (N5872, N5869);
buf BUF1 (N5873, N5841);
or OR4 (N5874, N5870, N1703, N1605, N3746);
nand NAND2 (N5875, N5873, N756);
not NOT1 (N5876, N5851);
not NOT1 (N5877, N5876);
or OR3 (N5878, N5865, N5200, N4875);
nor NOR3 (N5879, N5861, N4726, N3262);
nand NAND3 (N5880, N5864, N4372, N5053);
or OR3 (N5881, N5877, N256, N3533);
buf BUF1 (N5882, N5857);
and AND3 (N5883, N5882, N5255, N4521);
not NOT1 (N5884, N5872);
not NOT1 (N5885, N5880);
xor XOR2 (N5886, N5879, N1837);
xor XOR2 (N5887, N5878, N3173);
not NOT1 (N5888, N5881);
xor XOR2 (N5889, N5852, N4471);
nor NOR3 (N5890, N5889, N4241, N2671);
or OR3 (N5891, N5883, N2144, N1870);
not NOT1 (N5892, N5890);
nor NOR3 (N5893, N5875, N2238, N1730);
not NOT1 (N5894, N5892);
nand NAND2 (N5895, N5894, N2801);
buf BUF1 (N5896, N5895);
or OR3 (N5897, N5884, N611, N5807);
not NOT1 (N5898, N5888);
or OR2 (N5899, N5891, N5060);
buf BUF1 (N5900, N5896);
xor XOR2 (N5901, N5900, N2603);
not NOT1 (N5902, N5893);
and AND2 (N5903, N5874, N3475);
buf BUF1 (N5904, N5902);
nand NAND4 (N5905, N5904, N4615, N1101, N5103);
and AND2 (N5906, N5901, N4401);
nor NOR2 (N5907, N5897, N1182);
xor XOR2 (N5908, N5906, N2911);
nand NAND3 (N5909, N5907, N4830, N687);
buf BUF1 (N5910, N5905);
buf BUF1 (N5911, N5871);
and AND4 (N5912, N5898, N4039, N4118, N1489);
buf BUF1 (N5913, N5899);
nand NAND4 (N5914, N5885, N5348, N4268, N2820);
not NOT1 (N5915, N5912);
not NOT1 (N5916, N5910);
buf BUF1 (N5917, N5915);
nor NOR3 (N5918, N5887, N2842, N5351);
and AND3 (N5919, N5913, N715, N2235);
not NOT1 (N5920, N5886);
or OR3 (N5921, N5909, N5203, N5069);
xor XOR2 (N5922, N5908, N2833);
xor XOR2 (N5923, N5903, N3565);
not NOT1 (N5924, N5921);
nor NOR4 (N5925, N5916, N2927, N2461, N4358);
xor XOR2 (N5926, N5919, N1809);
nand NAND4 (N5927, N5922, N4265, N1014, N3227);
xor XOR2 (N5928, N5926, N5667);
xor XOR2 (N5929, N5925, N4725);
xor XOR2 (N5930, N5923, N3598);
and AND4 (N5931, N5930, N3367, N3000, N1732);
not NOT1 (N5932, N5927);
and AND4 (N5933, N5911, N763, N5124, N2202);
and AND2 (N5934, N5933, N5246);
buf BUF1 (N5935, N5934);
not NOT1 (N5936, N5929);
xor XOR2 (N5937, N5924, N2825);
xor XOR2 (N5938, N5917, N5877);
and AND2 (N5939, N5937, N3795);
not NOT1 (N5940, N5918);
nand NAND3 (N5941, N5940, N818, N4984);
and AND3 (N5942, N5932, N2991, N2707);
xor XOR2 (N5943, N5931, N2069);
not NOT1 (N5944, N5935);
or OR3 (N5945, N5914, N3545, N3476);
buf BUF1 (N5946, N5944);
xor XOR2 (N5947, N5920, N2456);
xor XOR2 (N5948, N5945, N5147);
buf BUF1 (N5949, N5948);
nor NOR2 (N5950, N5941, N3027);
or OR4 (N5951, N5943, N321, N3032, N1881);
not NOT1 (N5952, N5950);
nand NAND3 (N5953, N5946, N1259, N1483);
nor NOR4 (N5954, N5942, N2994, N2790, N3347);
nor NOR3 (N5955, N5951, N4850, N3651);
and AND4 (N5956, N5939, N2006, N684, N3648);
not NOT1 (N5957, N5955);
buf BUF1 (N5958, N5928);
and AND3 (N5959, N5936, N5589, N1410);
not NOT1 (N5960, N5938);
and AND4 (N5961, N5960, N5535, N2148, N5919);
not NOT1 (N5962, N5952);
not NOT1 (N5963, N5959);
buf BUF1 (N5964, N5962);
and AND2 (N5965, N5956, N2657);
nand NAND3 (N5966, N5947, N4923, N2158);
or OR3 (N5967, N5963, N4934, N4553);
or OR3 (N5968, N5953, N3683, N5904);
and AND2 (N5969, N5961, N4616);
or OR3 (N5970, N5968, N5699, N1072);
xor XOR2 (N5971, N5966, N5775);
and AND3 (N5972, N5957, N1287, N563);
xor XOR2 (N5973, N5949, N1519);
and AND2 (N5974, N5969, N4014);
buf BUF1 (N5975, N5972);
and AND2 (N5976, N5958, N4520);
or OR4 (N5977, N5954, N889, N1538, N2315);
nand NAND2 (N5978, N5973, N5440);
not NOT1 (N5979, N5970);
nand NAND4 (N5980, N5978, N2578, N1106, N5398);
buf BUF1 (N5981, N5964);
or OR3 (N5982, N5974, N4838, N3159);
nand NAND3 (N5983, N5965, N5466, N5292);
and AND4 (N5984, N5981, N4178, N4569, N4983);
xor XOR2 (N5985, N5984, N5118);
xor XOR2 (N5986, N5979, N2296);
not NOT1 (N5987, N5971);
or OR2 (N5988, N5982, N4475);
nor NOR3 (N5989, N5986, N3573, N4192);
xor XOR2 (N5990, N5988, N2451);
not NOT1 (N5991, N5975);
or OR2 (N5992, N5989, N3029);
or OR4 (N5993, N5980, N2916, N3610, N5774);
and AND2 (N5994, N5967, N870);
and AND3 (N5995, N5990, N5877, N1322);
nand NAND4 (N5996, N5985, N444, N1636, N3);
nor NOR3 (N5997, N5992, N4838, N3787);
buf BUF1 (N5998, N5991);
not NOT1 (N5999, N5995);
nand NAND3 (N6000, N5977, N1256, N2208);
not NOT1 (N6001, N5993);
and AND2 (N6002, N5997, N226);
buf BUF1 (N6003, N5976);
nand NAND2 (N6004, N6002, N285);
buf BUF1 (N6005, N5994);
nor NOR2 (N6006, N6003, N4140);
nor NOR2 (N6007, N6006, N898);
buf BUF1 (N6008, N6000);
not NOT1 (N6009, N5999);
or OR3 (N6010, N6005, N5440, N1804);
buf BUF1 (N6011, N5998);
xor XOR2 (N6012, N6004, N3732);
or OR4 (N6013, N6011, N2971, N832, N2293);
or OR3 (N6014, N6012, N5577, N1011);
and AND3 (N6015, N6008, N653, N934);
buf BUF1 (N6016, N5983);
nor NOR3 (N6017, N6007, N3751, N3392);
xor XOR2 (N6018, N6017, N3810);
xor XOR2 (N6019, N6015, N3021);
and AND2 (N6020, N6013, N5648);
buf BUF1 (N6021, N5996);
xor XOR2 (N6022, N6018, N5952);
buf BUF1 (N6023, N6016);
buf BUF1 (N6024, N6020);
and AND3 (N6025, N6023, N1328, N5436);
and AND4 (N6026, N5987, N4488, N3827, N2159);
xor XOR2 (N6027, N6001, N4358);
nand NAND4 (N6028, N6022, N5045, N2045, N632);
or OR2 (N6029, N6024, N3543);
xor XOR2 (N6030, N6028, N6024);
nor NOR2 (N6031, N6010, N1861);
or OR4 (N6032, N6021, N2070, N5823, N1954);
xor XOR2 (N6033, N6030, N1542);
buf BUF1 (N6034, N6014);
not NOT1 (N6035, N6027);
not NOT1 (N6036, N6026);
nand NAND3 (N6037, N6035, N4508, N1154);
and AND3 (N6038, N6032, N4321, N3736);
not NOT1 (N6039, N6034);
not NOT1 (N6040, N6036);
nand NAND4 (N6041, N6009, N462, N4241, N409);
nor NOR3 (N6042, N6038, N3285, N2273);
xor XOR2 (N6043, N6031, N3042);
and AND3 (N6044, N6019, N2175, N5502);
nor NOR4 (N6045, N6040, N4444, N818, N3174);
and AND2 (N6046, N6041, N2012);
or OR3 (N6047, N6033, N4087, N1453);
and AND4 (N6048, N6025, N3961, N1168, N1548);
not NOT1 (N6049, N6029);
not NOT1 (N6050, N6047);
buf BUF1 (N6051, N6044);
nand NAND2 (N6052, N6051, N2804);
nand NAND2 (N6053, N6052, N1259);
nand NAND3 (N6054, N6043, N1818, N3648);
nand NAND3 (N6055, N6054, N1990, N4286);
or OR2 (N6056, N6050, N2313);
nor NOR3 (N6057, N6048, N5701, N228);
nor NOR4 (N6058, N6049, N4504, N2677, N1242);
buf BUF1 (N6059, N6058);
nand NAND2 (N6060, N6037, N513);
nor NOR4 (N6061, N6055, N4939, N2973, N425);
xor XOR2 (N6062, N6053, N1127);
not NOT1 (N6063, N6060);
buf BUF1 (N6064, N6056);
nand NAND3 (N6065, N6042, N868, N2537);
and AND2 (N6066, N6064, N4016);
nand NAND3 (N6067, N6065, N1617, N3270);
not NOT1 (N6068, N6061);
nor NOR2 (N6069, N6059, N3319);
nor NOR3 (N6070, N6057, N6036, N4869);
nor NOR4 (N6071, N6063, N796, N5373, N3524);
xor XOR2 (N6072, N6039, N1820);
and AND2 (N6073, N6062, N3121);
nand NAND4 (N6074, N6072, N4409, N4013, N1595);
not NOT1 (N6075, N6073);
nand NAND4 (N6076, N6071, N4953, N2031, N4353);
nand NAND3 (N6077, N6069, N188, N253);
xor XOR2 (N6078, N6045, N4573);
buf BUF1 (N6079, N6077);
buf BUF1 (N6080, N6075);
and AND4 (N6081, N6067, N2240, N758, N1238);
and AND2 (N6082, N6068, N1280);
xor XOR2 (N6083, N6074, N2461);
not NOT1 (N6084, N6083);
not NOT1 (N6085, N6076);
xor XOR2 (N6086, N6079, N2213);
xor XOR2 (N6087, N6078, N5796);
buf BUF1 (N6088, N6070);
xor XOR2 (N6089, N6081, N1239);
and AND4 (N6090, N6085, N5637, N2260, N4127);
or OR3 (N6091, N6080, N5913, N5388);
or OR4 (N6092, N6088, N1986, N2828, N4723);
nor NOR4 (N6093, N6089, N4249, N1364, N4291);
buf BUF1 (N6094, N6087);
or OR3 (N6095, N6082, N4236, N1662);
buf BUF1 (N6096, N6084);
nor NOR2 (N6097, N6096, N5822);
or OR3 (N6098, N6090, N2272, N961);
buf BUF1 (N6099, N6046);
buf BUF1 (N6100, N6066);
nor NOR4 (N6101, N6099, N1500, N5663, N467);
or OR3 (N6102, N6100, N873, N4202);
not NOT1 (N6103, N6097);
nor NOR3 (N6104, N6095, N1118, N5269);
nand NAND3 (N6105, N6092, N2083, N4685);
buf BUF1 (N6106, N6101);
nand NAND3 (N6107, N6093, N5932, N557);
not NOT1 (N6108, N6106);
and AND4 (N6109, N6094, N164, N4175, N4779);
and AND4 (N6110, N6107, N4837, N2998, N5848);
not NOT1 (N6111, N6109);
or OR2 (N6112, N6091, N3969);
buf BUF1 (N6113, N6111);
or OR2 (N6114, N6104, N3741);
buf BUF1 (N6115, N6112);
xor XOR2 (N6116, N6102, N394);
xor XOR2 (N6117, N6114, N4041);
and AND2 (N6118, N6115, N5113);
nand NAND4 (N6119, N6116, N5941, N4988, N5544);
nand NAND2 (N6120, N6110, N2098);
not NOT1 (N6121, N6086);
nor NOR4 (N6122, N6118, N3836, N116, N2792);
xor XOR2 (N6123, N6120, N4981);
not NOT1 (N6124, N6108);
buf BUF1 (N6125, N6117);
buf BUF1 (N6126, N6121);
xor XOR2 (N6127, N6113, N921);
not NOT1 (N6128, N6119);
xor XOR2 (N6129, N6126, N3176);
buf BUF1 (N6130, N6098);
or OR4 (N6131, N6124, N2498, N1849, N3825);
not NOT1 (N6132, N6129);
xor XOR2 (N6133, N6123, N4661);
not NOT1 (N6134, N6127);
not NOT1 (N6135, N6133);
buf BUF1 (N6136, N6132);
or OR2 (N6137, N6135, N1255);
or OR4 (N6138, N6137, N2507, N5728, N3006);
not NOT1 (N6139, N6125);
buf BUF1 (N6140, N6136);
xor XOR2 (N6141, N6139, N2686);
nand NAND4 (N6142, N6122, N3516, N4551, N6135);
or OR3 (N6143, N6130, N3239, N2845);
xor XOR2 (N6144, N6142, N3868);
xor XOR2 (N6145, N6134, N1424);
buf BUF1 (N6146, N6128);
nor NOR4 (N6147, N6145, N2908, N6064, N1810);
or OR4 (N6148, N6144, N2693, N4801, N1274);
nand NAND3 (N6149, N6103, N2005, N5323);
nor NOR3 (N6150, N6143, N2651, N3765);
and AND2 (N6151, N6141, N3973);
xor XOR2 (N6152, N6148, N60);
xor XOR2 (N6153, N6151, N4663);
buf BUF1 (N6154, N6105);
and AND2 (N6155, N6149, N5974);
not NOT1 (N6156, N6152);
and AND2 (N6157, N6140, N6066);
buf BUF1 (N6158, N6131);
nor NOR4 (N6159, N6153, N1060, N1416, N5656);
or OR2 (N6160, N6159, N4555);
or OR2 (N6161, N6138, N352);
or OR3 (N6162, N6161, N1989, N3295);
not NOT1 (N6163, N6156);
nor NOR3 (N6164, N6163, N5934, N3536);
buf BUF1 (N6165, N6155);
not NOT1 (N6166, N6165);
nand NAND2 (N6167, N6158, N3809);
or OR4 (N6168, N6146, N5001, N3714, N4904);
or OR3 (N6169, N6157, N1308, N4356);
and AND2 (N6170, N6150, N603);
or OR3 (N6171, N6166, N519, N1155);
or OR4 (N6172, N6171, N5022, N4794, N3351);
nor NOR2 (N6173, N6164, N3294);
nand NAND2 (N6174, N6169, N4451);
and AND4 (N6175, N6173, N517, N986, N1088);
or OR3 (N6176, N6172, N5305, N835);
and AND2 (N6177, N6174, N3035);
buf BUF1 (N6178, N6175);
nor NOR4 (N6179, N6178, N3127, N4140, N643);
buf BUF1 (N6180, N6179);
nor NOR2 (N6181, N6177, N4597);
xor XOR2 (N6182, N6176, N2882);
nor NOR4 (N6183, N6181, N3737, N6099, N5044);
nand NAND4 (N6184, N6160, N4576, N4118, N2570);
xor XOR2 (N6185, N6182, N573);
or OR2 (N6186, N6180, N3410);
nand NAND2 (N6187, N6154, N2926);
nor NOR2 (N6188, N6168, N67);
nor NOR4 (N6189, N6170, N250, N3903, N3139);
not NOT1 (N6190, N6185);
buf BUF1 (N6191, N6167);
and AND2 (N6192, N6184, N1304);
xor XOR2 (N6193, N6188, N1962);
xor XOR2 (N6194, N6187, N1233);
xor XOR2 (N6195, N6191, N1702);
and AND4 (N6196, N6162, N4810, N1792, N5627);
or OR3 (N6197, N6186, N5835, N746);
or OR2 (N6198, N6147, N1849);
and AND2 (N6199, N6197, N2323);
and AND4 (N6200, N6192, N4036, N1341, N3898);
buf BUF1 (N6201, N6194);
xor XOR2 (N6202, N6183, N2711);
xor XOR2 (N6203, N6196, N4255);
and AND2 (N6204, N6202, N4629);
nor NOR2 (N6205, N6203, N5470);
or OR2 (N6206, N6201, N3081);
xor XOR2 (N6207, N6195, N2197);
nor NOR2 (N6208, N6205, N4637);
buf BUF1 (N6209, N6200);
xor XOR2 (N6210, N6189, N3766);
and AND3 (N6211, N6198, N4580, N1243);
nand NAND2 (N6212, N6193, N2439);
not NOT1 (N6213, N6209);
nand NAND3 (N6214, N6199, N818, N2330);
or OR4 (N6215, N6211, N1585, N1746, N5086);
xor XOR2 (N6216, N6212, N5016);
xor XOR2 (N6217, N6207, N4699);
and AND4 (N6218, N6213, N4305, N4226, N1986);
nand NAND4 (N6219, N6208, N256, N5478, N2515);
or OR4 (N6220, N6190, N1740, N3502, N4239);
not NOT1 (N6221, N6210);
nand NAND4 (N6222, N6220, N1446, N5936, N3371);
nand NAND3 (N6223, N6221, N2107, N5182);
nor NOR3 (N6224, N6215, N4513, N5305);
or OR4 (N6225, N6206, N3283, N2498, N3434);
not NOT1 (N6226, N6204);
not NOT1 (N6227, N6219);
or OR2 (N6228, N6224, N1610);
and AND2 (N6229, N6227, N2913);
nand NAND3 (N6230, N6218, N59, N886);
or OR4 (N6231, N6216, N587, N4951, N4944);
xor XOR2 (N6232, N6222, N5150);
not NOT1 (N6233, N6226);
or OR3 (N6234, N6214, N4085, N4387);
xor XOR2 (N6235, N6231, N2630);
buf BUF1 (N6236, N6232);
buf BUF1 (N6237, N6235);
not NOT1 (N6238, N6233);
xor XOR2 (N6239, N6238, N2421);
or OR2 (N6240, N6234, N5452);
or OR2 (N6241, N6228, N638);
and AND3 (N6242, N6240, N2249, N5272);
or OR4 (N6243, N6223, N703, N1777, N4909);
nand NAND3 (N6244, N6241, N3425, N1342);
buf BUF1 (N6245, N6237);
nand NAND4 (N6246, N6244, N5346, N4932, N5119);
or OR3 (N6247, N6229, N1240, N6124);
xor XOR2 (N6248, N6239, N2962);
nand NAND2 (N6249, N6242, N1628);
xor XOR2 (N6250, N6225, N5928);
xor XOR2 (N6251, N6248, N2911);
xor XOR2 (N6252, N6247, N2386);
nand NAND3 (N6253, N6243, N2251, N1150);
nor NOR4 (N6254, N6253, N888, N1993, N1158);
and AND3 (N6255, N6230, N4990, N1191);
and AND2 (N6256, N6252, N4203);
buf BUF1 (N6257, N6245);
not NOT1 (N6258, N6249);
not NOT1 (N6259, N6236);
and AND3 (N6260, N6256, N4618, N2333);
not NOT1 (N6261, N6246);
buf BUF1 (N6262, N6250);
xor XOR2 (N6263, N6261, N4638);
or OR2 (N6264, N6260, N1615);
xor XOR2 (N6265, N6258, N902);
and AND3 (N6266, N6259, N5205, N1749);
not NOT1 (N6267, N6257);
nor NOR3 (N6268, N6262, N1676, N1544);
nor NOR4 (N6269, N6267, N4512, N1519, N26);
xor XOR2 (N6270, N6266, N1705);
not NOT1 (N6271, N6251);
and AND4 (N6272, N6270, N5671, N4169, N5853);
buf BUF1 (N6273, N6255);
nand NAND2 (N6274, N6264, N1409);
xor XOR2 (N6275, N6217, N850);
xor XOR2 (N6276, N6269, N855);
nand NAND4 (N6277, N6265, N3160, N3934, N1029);
and AND3 (N6278, N6268, N2216, N1798);
or OR3 (N6279, N6277, N5289, N2530);
not NOT1 (N6280, N6278);
nor NOR3 (N6281, N6272, N826, N1505);
xor XOR2 (N6282, N6254, N3427);
buf BUF1 (N6283, N6275);
buf BUF1 (N6284, N6273);
nor NOR2 (N6285, N6281, N2342);
and AND2 (N6286, N6279, N4128);
and AND4 (N6287, N6274, N5391, N5836, N4999);
not NOT1 (N6288, N6283);
or OR2 (N6289, N6280, N1243);
or OR4 (N6290, N6284, N3909, N4234, N5246);
or OR3 (N6291, N6287, N279, N2321);
not NOT1 (N6292, N6276);
not NOT1 (N6293, N6286);
and AND2 (N6294, N6289, N5248);
nand NAND2 (N6295, N6282, N3950);
nor NOR2 (N6296, N6291, N2312);
buf BUF1 (N6297, N6271);
nand NAND4 (N6298, N6295, N197, N4988, N962);
not NOT1 (N6299, N6290);
or OR4 (N6300, N6294, N144, N3733, N5037);
nor NOR3 (N6301, N6293, N4807, N1273);
nor NOR4 (N6302, N6298, N4831, N2730, N2357);
nand NAND2 (N6303, N6302, N6134);
or OR3 (N6304, N6300, N3826, N4811);
nor NOR3 (N6305, N6263, N2380, N3860);
and AND2 (N6306, N6303, N930);
not NOT1 (N6307, N6305);
nand NAND2 (N6308, N6297, N3690);
nor NOR2 (N6309, N6299, N2326);
buf BUF1 (N6310, N6301);
nor NOR2 (N6311, N6296, N626);
xor XOR2 (N6312, N6304, N1293);
xor XOR2 (N6313, N6310, N2751);
buf BUF1 (N6314, N6306);
or OR2 (N6315, N6288, N3080);
buf BUF1 (N6316, N6315);
or OR4 (N6317, N6311, N6063, N4465, N3568);
not NOT1 (N6318, N6314);
nand NAND2 (N6319, N6307, N786);
nand NAND4 (N6320, N6285, N2066, N3624, N1930);
nor NOR3 (N6321, N6318, N2012, N4328);
nand NAND2 (N6322, N6316, N560);
nand NAND4 (N6323, N6322, N1999, N3131, N1356);
xor XOR2 (N6324, N6308, N5113);
xor XOR2 (N6325, N6317, N4084);
and AND3 (N6326, N6323, N6308, N4566);
buf BUF1 (N6327, N6326);
nand NAND3 (N6328, N6321, N1568, N5233);
not NOT1 (N6329, N6309);
not NOT1 (N6330, N6327);
nor NOR3 (N6331, N6292, N5993, N2180);
buf BUF1 (N6332, N6320);
xor XOR2 (N6333, N6319, N3007);
buf BUF1 (N6334, N6329);
xor XOR2 (N6335, N6324, N2018);
not NOT1 (N6336, N6313);
buf BUF1 (N6337, N6335);
xor XOR2 (N6338, N6336, N3698);
or OR4 (N6339, N6325, N2709, N2585, N3152);
nand NAND2 (N6340, N6332, N3846);
or OR4 (N6341, N6339, N6271, N3438, N3321);
or OR4 (N6342, N6333, N2842, N3816, N741);
and AND3 (N6343, N6338, N4003, N6339);
or OR3 (N6344, N6331, N5740, N2402);
nand NAND4 (N6345, N6334, N758, N5145, N4241);
and AND4 (N6346, N6343, N4816, N2285, N1641);
nor NOR4 (N6347, N6342, N247, N3861, N1016);
xor XOR2 (N6348, N6340, N540);
xor XOR2 (N6349, N6337, N5154);
not NOT1 (N6350, N6349);
nand NAND3 (N6351, N6312, N3243, N1298);
or OR2 (N6352, N6345, N2340);
nor NOR2 (N6353, N6348, N1281);
nand NAND3 (N6354, N6352, N79, N5968);
buf BUF1 (N6355, N6347);
and AND3 (N6356, N6346, N532, N995);
nor NOR3 (N6357, N6354, N4168, N2886);
nand NAND4 (N6358, N6351, N983, N3973, N5086);
nand NAND2 (N6359, N6328, N2485);
not NOT1 (N6360, N6357);
nor NOR2 (N6361, N6353, N4277);
buf BUF1 (N6362, N6355);
and AND4 (N6363, N6361, N255, N4600, N6252);
nor NOR2 (N6364, N6344, N5151);
buf BUF1 (N6365, N6362);
and AND3 (N6366, N6330, N5082, N6209);
not NOT1 (N6367, N6360);
not NOT1 (N6368, N6366);
nor NOR3 (N6369, N6367, N1151, N1771);
buf BUF1 (N6370, N6359);
not NOT1 (N6371, N6363);
nand NAND4 (N6372, N6370, N4361, N4157, N5715);
xor XOR2 (N6373, N6358, N4033);
buf BUF1 (N6374, N6368);
xor XOR2 (N6375, N6350, N2641);
and AND2 (N6376, N6341, N588);
or OR3 (N6377, N6371, N1845, N4975);
or OR2 (N6378, N6356, N4679);
buf BUF1 (N6379, N6373);
not NOT1 (N6380, N6379);
and AND2 (N6381, N6374, N6267);
and AND3 (N6382, N6364, N1878, N938);
not NOT1 (N6383, N6382);
buf BUF1 (N6384, N6381);
xor XOR2 (N6385, N6372, N4194);
nor NOR4 (N6386, N6384, N5605, N1661, N5051);
nand NAND2 (N6387, N6375, N6271);
or OR2 (N6388, N6383, N1744);
nor NOR3 (N6389, N6385, N5708, N112);
or OR2 (N6390, N6386, N471);
buf BUF1 (N6391, N6389);
nand NAND2 (N6392, N6377, N4058);
xor XOR2 (N6393, N6391, N3679);
or OR2 (N6394, N6369, N5530);
xor XOR2 (N6395, N6392, N4048);
xor XOR2 (N6396, N6388, N534);
nor NOR3 (N6397, N6396, N1405, N3559);
nand NAND3 (N6398, N6390, N795, N5765);
and AND3 (N6399, N6393, N5077, N5637);
buf BUF1 (N6400, N6376);
not NOT1 (N6401, N6380);
buf BUF1 (N6402, N6400);
not NOT1 (N6403, N6399);
or OR3 (N6404, N6395, N3058, N837);
buf BUF1 (N6405, N6398);
xor XOR2 (N6406, N6378, N3425);
buf BUF1 (N6407, N6403);
and AND2 (N6408, N6394, N1723);
nand NAND3 (N6409, N6401, N4727, N402);
and AND4 (N6410, N6365, N5244, N813, N1962);
buf BUF1 (N6411, N6404);
not NOT1 (N6412, N6411);
nand NAND3 (N6413, N6409, N4090, N2630);
not NOT1 (N6414, N6397);
buf BUF1 (N6415, N6407);
xor XOR2 (N6416, N6405, N2052);
nor NOR4 (N6417, N6410, N6349, N4757, N3744);
and AND2 (N6418, N6417, N4983);
or OR2 (N6419, N6412, N1581);
and AND4 (N6420, N6415, N627, N1043, N5925);
xor XOR2 (N6421, N6413, N5120);
nand NAND4 (N6422, N6387, N3871, N2489, N3589);
endmodule