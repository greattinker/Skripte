// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N3219,N3216,N3214,N3218,N3220,N3208,N3211,N3213,N3210,N3221;

and AND2 (N22, N21, N18);
xor XOR2 (N23, N18, N12);
xor XOR2 (N24, N7, N10);
xor XOR2 (N25, N5, N22);
xor XOR2 (N26, N23, N25);
nor NOR4 (N27, N17, N3, N9, N3);
and AND2 (N28, N12, N24);
or OR4 (N29, N21, N2, N10, N26);
buf BUF1 (N30, N10);
xor XOR2 (N31, N2, N12);
nor NOR2 (N32, N6, N26);
xor XOR2 (N33, N30, N8);
buf BUF1 (N34, N16);
and AND4 (N35, N5, N12, N12, N19);
nor NOR4 (N36, N26, N29, N3, N15);
or OR4 (N37, N10, N27, N23, N25);
nand NAND2 (N38, N4, N16);
nor NOR4 (N39, N14, N19, N25, N12);
nand NAND4 (N40, N35, N34, N16, N13);
and AND4 (N41, N27, N22, N40, N31);
nor NOR3 (N42, N13, N2, N41);
or OR4 (N43, N21, N19, N41, N22);
and AND2 (N44, N39, N7);
not NOT1 (N45, N18);
not NOT1 (N46, N37);
not NOT1 (N47, N38);
xor XOR2 (N48, N45, N37);
or OR3 (N49, N32, N44, N20);
buf BUF1 (N50, N42);
not NOT1 (N51, N24);
not NOT1 (N52, N49);
and AND4 (N53, N52, N23, N1, N32);
buf BUF1 (N54, N28);
xor XOR2 (N55, N48, N25);
buf BUF1 (N56, N43);
and AND4 (N57, N47, N1, N32, N35);
xor XOR2 (N58, N50, N47);
nand NAND3 (N59, N58, N23, N58);
and AND3 (N60, N51, N47, N39);
buf BUF1 (N61, N59);
and AND2 (N62, N55, N28);
not NOT1 (N63, N36);
nand NAND3 (N64, N53, N42, N42);
nor NOR4 (N65, N64, N4, N18, N18);
buf BUF1 (N66, N46);
not NOT1 (N67, N54);
xor XOR2 (N68, N33, N46);
nand NAND4 (N69, N67, N25, N52, N57);
or OR4 (N70, N59, N38, N55, N15);
xor XOR2 (N71, N61, N51);
and AND2 (N72, N69, N44);
and AND4 (N73, N63, N37, N57, N42);
xor XOR2 (N74, N60, N33);
and AND3 (N75, N74, N20, N25);
or OR3 (N76, N66, N73, N29);
and AND3 (N77, N74, N50, N61);
nor NOR4 (N78, N76, N58, N76, N74);
or OR3 (N79, N72, N45, N53);
nor NOR2 (N80, N68, N30);
buf BUF1 (N81, N77);
or OR3 (N82, N62, N47, N72);
not NOT1 (N83, N56);
or OR4 (N84, N82, N36, N68, N58);
buf BUF1 (N85, N65);
nand NAND3 (N86, N75, N12, N43);
not NOT1 (N87, N81);
buf BUF1 (N88, N70);
buf BUF1 (N89, N83);
not NOT1 (N90, N89);
not NOT1 (N91, N84);
and AND2 (N92, N71, N87);
not NOT1 (N93, N55);
nor NOR3 (N94, N80, N69, N35);
or OR4 (N95, N85, N24, N12, N51);
nand NAND2 (N96, N79, N66);
buf BUF1 (N97, N93);
and AND4 (N98, N90, N16, N42, N26);
buf BUF1 (N99, N94);
xor XOR2 (N100, N91, N75);
xor XOR2 (N101, N100, N20);
buf BUF1 (N102, N78);
nor NOR4 (N103, N86, N55, N90, N35);
nor NOR4 (N104, N92, N2, N2, N15);
nand NAND3 (N105, N101, N104, N41);
not NOT1 (N106, N101);
and AND4 (N107, N99, N65, N72, N13);
buf BUF1 (N108, N96);
and AND3 (N109, N107, N92, N15);
and AND3 (N110, N97, N103, N107);
nand NAND3 (N111, N74, N13, N41);
or OR3 (N112, N98, N15, N91);
or OR2 (N113, N88, N52);
nor NOR4 (N114, N106, N53, N3, N40);
xor XOR2 (N115, N110, N108);
nor NOR3 (N116, N47, N52, N33);
nand NAND3 (N117, N111, N76, N32);
or OR4 (N118, N105, N117, N103, N10);
nand NAND2 (N119, N110, N76);
buf BUF1 (N120, N119);
xor XOR2 (N121, N115, N94);
xor XOR2 (N122, N102, N116);
buf BUF1 (N123, N19);
or OR4 (N124, N114, N100, N113, N74);
nor NOR2 (N125, N46, N114);
and AND4 (N126, N109, N123, N7, N23);
or OR2 (N127, N33, N4);
buf BUF1 (N128, N125);
buf BUF1 (N129, N126);
buf BUF1 (N130, N121);
and AND3 (N131, N122, N100, N36);
and AND3 (N132, N124, N70, N29);
or OR3 (N133, N128, N90, N45);
and AND2 (N134, N133, N24);
buf BUF1 (N135, N118);
xor XOR2 (N136, N112, N129);
nor NOR3 (N137, N132, N93, N38);
not NOT1 (N138, N108);
and AND4 (N139, N127, N31, N89, N23);
xor XOR2 (N140, N134, N20);
and AND3 (N141, N95, N107, N89);
buf BUF1 (N142, N138);
and AND3 (N143, N141, N114, N117);
buf BUF1 (N144, N135);
xor XOR2 (N145, N131, N105);
nand NAND2 (N146, N143, N112);
nor NOR4 (N147, N130, N121, N145, N45);
not NOT1 (N148, N138);
not NOT1 (N149, N136);
nor NOR3 (N150, N144, N148, N76);
buf BUF1 (N151, N126);
and AND3 (N152, N147, N16, N31);
not NOT1 (N153, N149);
and AND4 (N154, N151, N62, N52, N54);
and AND2 (N155, N140, N129);
nand NAND2 (N156, N154, N45);
or OR3 (N157, N156, N74, N93);
buf BUF1 (N158, N120);
nand NAND3 (N159, N158, N58, N45);
nand NAND4 (N160, N137, N36, N117, N102);
not NOT1 (N161, N142);
or OR2 (N162, N139, N9);
or OR4 (N163, N160, N3, N99, N145);
nand NAND2 (N164, N159, N15);
not NOT1 (N165, N163);
and AND4 (N166, N155, N100, N67, N29);
not NOT1 (N167, N150);
or OR3 (N168, N165, N106, N3);
nor NOR4 (N169, N153, N30, N25, N69);
or OR4 (N170, N152, N60, N37, N151);
or OR3 (N171, N162, N12, N16);
or OR2 (N172, N166, N143);
nand NAND2 (N173, N157, N67);
and AND2 (N174, N170, N127);
nand NAND4 (N175, N171, N48, N142, N97);
nor NOR2 (N176, N167, N144);
and AND3 (N177, N173, N109, N92);
or OR4 (N178, N174, N51, N98, N92);
or OR4 (N179, N164, N82, N50, N156);
xor XOR2 (N180, N169, N102);
nand NAND4 (N181, N175, N43, N37, N2);
or OR4 (N182, N179, N26, N140, N26);
buf BUF1 (N183, N178);
or OR3 (N184, N176, N21, N102);
and AND2 (N185, N183, N120);
nand NAND3 (N186, N185, N108, N44);
nand NAND3 (N187, N181, N12, N39);
xor XOR2 (N188, N184, N23);
buf BUF1 (N189, N177);
not NOT1 (N190, N188);
and AND3 (N191, N180, N9, N14);
nand NAND2 (N192, N168, N52);
xor XOR2 (N193, N192, N100);
or OR3 (N194, N146, N125, N31);
xor XOR2 (N195, N190, N75);
or OR2 (N196, N195, N189);
and AND2 (N197, N169, N62);
and AND2 (N198, N196, N186);
xor XOR2 (N199, N152, N29);
nor NOR3 (N200, N194, N166, N189);
nand NAND2 (N201, N200, N82);
not NOT1 (N202, N187);
or OR3 (N203, N193, N76, N84);
or OR3 (N204, N198, N98, N20);
nor NOR3 (N205, N203, N204, N25);
or OR4 (N206, N199, N61, N190, N153);
or OR2 (N207, N206, N110);
nor NOR2 (N208, N59, N130);
xor XOR2 (N209, N201, N146);
nand NAND3 (N210, N191, N140, N100);
nor NOR4 (N211, N161, N144, N84, N185);
buf BUF1 (N212, N172);
nand NAND4 (N213, N182, N154, N68, N147);
buf BUF1 (N214, N213);
nand NAND3 (N215, N207, N159, N170);
xor XOR2 (N216, N208, N32);
nor NOR3 (N217, N209, N189, N84);
nor NOR2 (N218, N197, N73);
not NOT1 (N219, N210);
nand NAND4 (N220, N216, N29, N156, N149);
xor XOR2 (N221, N205, N40);
nand NAND4 (N222, N217, N130, N88, N109);
not NOT1 (N223, N221);
nor NOR3 (N224, N222, N162, N107);
nor NOR2 (N225, N223, N32);
xor XOR2 (N226, N211, N48);
and AND2 (N227, N202, N39);
nor NOR4 (N228, N224, N28, N124, N34);
and AND2 (N229, N225, N125);
nor NOR3 (N230, N226, N147, N117);
nand NAND4 (N231, N229, N107, N110, N86);
or OR3 (N232, N230, N209, N34);
not NOT1 (N233, N215);
nand NAND3 (N234, N227, N40, N9);
or OR3 (N235, N233, N191, N61);
buf BUF1 (N236, N228);
and AND4 (N237, N214, N162, N221, N17);
nand NAND2 (N238, N235, N231);
nand NAND4 (N239, N26, N92, N207, N137);
and AND2 (N240, N218, N185);
nor NOR2 (N241, N220, N49);
xor XOR2 (N242, N239, N211);
and AND4 (N243, N241, N182, N183, N92);
not NOT1 (N244, N237);
buf BUF1 (N245, N243);
nand NAND3 (N246, N232, N170, N121);
and AND2 (N247, N242, N3);
buf BUF1 (N248, N236);
xor XOR2 (N249, N248, N75);
not NOT1 (N250, N245);
nand NAND2 (N251, N247, N87);
not NOT1 (N252, N246);
xor XOR2 (N253, N250, N234);
or OR3 (N254, N189, N226, N76);
nand NAND4 (N255, N219, N177, N251, N14);
and AND2 (N256, N220, N119);
and AND2 (N257, N212, N56);
or OR4 (N258, N252, N169, N145, N140);
buf BUF1 (N259, N240);
nor NOR3 (N260, N253, N54, N237);
and AND4 (N261, N259, N50, N14, N77);
nor NOR4 (N262, N249, N30, N153, N205);
nor NOR2 (N263, N255, N149);
xor XOR2 (N264, N244, N195);
and AND4 (N265, N256, N202, N155, N250);
or OR2 (N266, N265, N217);
not NOT1 (N267, N264);
nand NAND2 (N268, N262, N45);
nand NAND2 (N269, N267, N115);
buf BUF1 (N270, N257);
xor XOR2 (N271, N261, N207);
nor NOR4 (N272, N266, N48, N78, N63);
or OR2 (N273, N269, N240);
xor XOR2 (N274, N271, N92);
not NOT1 (N275, N263);
nor NOR2 (N276, N272, N36);
not NOT1 (N277, N270);
nor NOR2 (N278, N274, N23);
not NOT1 (N279, N254);
xor XOR2 (N280, N276, N203);
nand NAND2 (N281, N277, N229);
buf BUF1 (N282, N238);
and AND4 (N283, N280, N171, N110, N188);
buf BUF1 (N284, N258);
xor XOR2 (N285, N281, N131);
nand NAND3 (N286, N273, N118, N125);
not NOT1 (N287, N268);
or OR4 (N288, N260, N252, N58, N60);
buf BUF1 (N289, N284);
xor XOR2 (N290, N289, N89);
xor XOR2 (N291, N282, N26);
xor XOR2 (N292, N285, N284);
not NOT1 (N293, N292);
and AND2 (N294, N288, N87);
not NOT1 (N295, N287);
nand NAND3 (N296, N283, N58, N9);
xor XOR2 (N297, N293, N56);
xor XOR2 (N298, N286, N190);
nand NAND3 (N299, N295, N240, N213);
and AND3 (N300, N290, N60, N261);
buf BUF1 (N301, N297);
nor NOR2 (N302, N298, N17);
nand NAND3 (N303, N294, N4, N297);
or OR3 (N304, N302, N284, N209);
and AND2 (N305, N304, N302);
or OR3 (N306, N303, N77, N245);
xor XOR2 (N307, N291, N246);
xor XOR2 (N308, N275, N92);
nor NOR4 (N309, N301, N85, N211, N234);
nor NOR3 (N310, N279, N228, N162);
or OR2 (N311, N307, N217);
buf BUF1 (N312, N311);
xor XOR2 (N313, N309, N105);
buf BUF1 (N314, N308);
nor NOR4 (N315, N305, N145, N149, N275);
buf BUF1 (N316, N314);
not NOT1 (N317, N310);
nand NAND4 (N318, N278, N79, N160, N110);
not NOT1 (N319, N318);
nor NOR4 (N320, N296, N64, N296, N60);
or OR3 (N321, N306, N174, N264);
not NOT1 (N322, N299);
and AND3 (N323, N320, N212, N18);
buf BUF1 (N324, N315);
xor XOR2 (N325, N313, N190);
or OR4 (N326, N317, N40, N294, N263);
or OR4 (N327, N325, N20, N249, N150);
not NOT1 (N328, N326);
nor NOR4 (N329, N328, N213, N200, N60);
nand NAND2 (N330, N312, N151);
not NOT1 (N331, N300);
nand NAND2 (N332, N324, N221);
xor XOR2 (N333, N330, N109);
not NOT1 (N334, N332);
nand NAND4 (N335, N327, N123, N136, N70);
nor NOR4 (N336, N319, N187, N255, N47);
not NOT1 (N337, N336);
xor XOR2 (N338, N333, N170);
or OR4 (N339, N338, N227, N31, N278);
or OR3 (N340, N331, N117, N289);
nor NOR3 (N341, N339, N329, N165);
nand NAND4 (N342, N168, N277, N163, N244);
or OR3 (N343, N335, N52, N122);
and AND4 (N344, N343, N117, N13, N318);
buf BUF1 (N345, N341);
not NOT1 (N346, N337);
not NOT1 (N347, N344);
xor XOR2 (N348, N345, N94);
xor XOR2 (N349, N321, N183);
xor XOR2 (N350, N323, N198);
nand NAND2 (N351, N334, N293);
and AND4 (N352, N351, N350, N24, N58);
not NOT1 (N353, N144);
or OR2 (N354, N349, N286);
nand NAND3 (N355, N348, N174, N251);
xor XOR2 (N356, N322, N45);
nand NAND2 (N357, N354, N344);
xor XOR2 (N358, N356, N210);
nor NOR3 (N359, N353, N155, N40);
buf BUF1 (N360, N357);
or OR4 (N361, N358, N161, N30, N38);
not NOT1 (N362, N316);
buf BUF1 (N363, N346);
nor NOR4 (N364, N361, N201, N320, N128);
buf BUF1 (N365, N340);
not NOT1 (N366, N355);
xor XOR2 (N367, N366, N301);
nor NOR4 (N368, N367, N338, N81, N317);
not NOT1 (N369, N368);
nand NAND3 (N370, N347, N315, N284);
xor XOR2 (N371, N352, N163);
nor NOR3 (N372, N363, N35, N370);
nor NOR2 (N373, N209, N355);
nor NOR3 (N374, N359, N345, N98);
or OR2 (N375, N362, N283);
xor XOR2 (N376, N360, N193);
nor NOR3 (N377, N364, N376, N304);
xor XOR2 (N378, N337, N365);
buf BUF1 (N379, N290);
or OR2 (N380, N372, N265);
xor XOR2 (N381, N374, N128);
nand NAND4 (N382, N381, N123, N266, N120);
and AND4 (N383, N377, N83, N146, N124);
not NOT1 (N384, N380);
nor NOR4 (N385, N379, N53, N106, N145);
nand NAND3 (N386, N369, N312, N316);
or OR4 (N387, N382, N2, N5, N300);
buf BUF1 (N388, N342);
nand NAND3 (N389, N378, N267, N61);
nand NAND3 (N390, N387, N360, N370);
buf BUF1 (N391, N375);
xor XOR2 (N392, N384, N175);
buf BUF1 (N393, N388);
buf BUF1 (N394, N391);
nand NAND2 (N395, N394, N390);
buf BUF1 (N396, N269);
not NOT1 (N397, N386);
and AND4 (N398, N389, N25, N131, N76);
not NOT1 (N399, N393);
and AND2 (N400, N385, N226);
and AND3 (N401, N392, N110, N100);
nand NAND4 (N402, N396, N315, N57, N395);
and AND3 (N403, N193, N44, N292);
xor XOR2 (N404, N402, N149);
nor NOR2 (N405, N398, N29);
or OR2 (N406, N371, N73);
xor XOR2 (N407, N403, N335);
buf BUF1 (N408, N405);
not NOT1 (N409, N399);
and AND2 (N410, N400, N98);
not NOT1 (N411, N406);
xor XOR2 (N412, N410, N309);
nand NAND4 (N413, N407, N397, N130, N85);
not NOT1 (N414, N12);
xor XOR2 (N415, N373, N232);
buf BUF1 (N416, N413);
or OR2 (N417, N408, N215);
and AND4 (N418, N411, N388, N333, N388);
or OR3 (N419, N415, N143, N383);
nand NAND4 (N420, N230, N289, N227, N9);
nor NOR3 (N421, N414, N308, N336);
nand NAND4 (N422, N420, N106, N23, N191);
buf BUF1 (N423, N401);
nor NOR3 (N424, N422, N138, N257);
xor XOR2 (N425, N417, N124);
buf BUF1 (N426, N424);
or OR3 (N427, N423, N17, N211);
buf BUF1 (N428, N416);
buf BUF1 (N429, N412);
buf BUF1 (N430, N421);
xor XOR2 (N431, N418, N365);
not NOT1 (N432, N431);
not NOT1 (N433, N427);
xor XOR2 (N434, N432, N45);
nor NOR2 (N435, N429, N63);
or OR4 (N436, N426, N282, N410, N26);
xor XOR2 (N437, N433, N16);
and AND2 (N438, N436, N163);
nor NOR3 (N439, N430, N88, N313);
not NOT1 (N440, N428);
nor NOR3 (N441, N404, N439, N238);
buf BUF1 (N442, N111);
xor XOR2 (N443, N441, N15);
nand NAND4 (N444, N440, N39, N191, N180);
or OR4 (N445, N425, N280, N362, N364);
nor NOR3 (N446, N445, N274, N99);
not NOT1 (N447, N444);
xor XOR2 (N448, N442, N339);
and AND3 (N449, N435, N55, N389);
and AND2 (N450, N409, N166);
buf BUF1 (N451, N448);
or OR4 (N452, N449, N428, N331, N257);
or OR2 (N453, N451, N293);
and AND4 (N454, N443, N270, N248, N49);
not NOT1 (N455, N447);
not NOT1 (N456, N454);
xor XOR2 (N457, N452, N11);
and AND2 (N458, N437, N310);
nand NAND3 (N459, N453, N58, N282);
or OR2 (N460, N419, N410);
not NOT1 (N461, N455);
or OR2 (N462, N461, N193);
nand NAND4 (N463, N462, N231, N150, N111);
nor NOR2 (N464, N438, N402);
buf BUF1 (N465, N456);
buf BUF1 (N466, N458);
nor NOR2 (N467, N465, N210);
and AND2 (N468, N450, N70);
buf BUF1 (N469, N466);
xor XOR2 (N470, N459, N281);
nand NAND3 (N471, N467, N46, N326);
nor NOR2 (N472, N463, N278);
nand NAND3 (N473, N469, N206, N349);
or OR2 (N474, N473, N366);
and AND2 (N475, N464, N77);
nand NAND4 (N476, N470, N308, N364, N147);
not NOT1 (N477, N434);
nor NOR4 (N478, N477, N181, N254, N477);
not NOT1 (N479, N475);
or OR4 (N480, N446, N213, N467, N228);
and AND2 (N481, N460, N178);
nor NOR4 (N482, N468, N453, N401, N161);
nor NOR3 (N483, N472, N313, N454);
or OR3 (N484, N474, N236, N479);
nor NOR2 (N485, N372, N103);
nand NAND4 (N486, N476, N313, N436, N89);
or OR2 (N487, N484, N331);
buf BUF1 (N488, N483);
xor XOR2 (N489, N481, N442);
xor XOR2 (N490, N489, N38);
xor XOR2 (N491, N486, N483);
and AND4 (N492, N485, N292, N152, N387);
not NOT1 (N493, N480);
buf BUF1 (N494, N491);
or OR4 (N495, N492, N231, N383, N135);
nor NOR2 (N496, N457, N185);
and AND3 (N497, N482, N344, N131);
not NOT1 (N498, N497);
or OR2 (N499, N498, N179);
nand NAND2 (N500, N499, N257);
nand NAND2 (N501, N494, N459);
nor NOR3 (N502, N478, N482, N325);
nor NOR2 (N503, N488, N105);
nand NAND3 (N504, N500, N410, N217);
xor XOR2 (N505, N496, N17);
xor XOR2 (N506, N495, N22);
or OR4 (N507, N471, N167, N290, N186);
and AND4 (N508, N493, N202, N218, N447);
buf BUF1 (N509, N503);
or OR2 (N510, N505, N6);
nor NOR3 (N511, N506, N413, N289);
nor NOR3 (N512, N508, N213, N13);
or OR4 (N513, N487, N304, N94, N253);
nor NOR4 (N514, N513, N365, N135, N204);
nor NOR3 (N515, N502, N173, N41);
and AND3 (N516, N504, N10, N67);
not NOT1 (N517, N515);
not NOT1 (N518, N516);
not NOT1 (N519, N509);
xor XOR2 (N520, N519, N464);
and AND3 (N521, N490, N391, N60);
nor NOR2 (N522, N514, N386);
buf BUF1 (N523, N507);
nor NOR2 (N524, N501, N196);
or OR4 (N525, N521, N11, N488, N429);
or OR3 (N526, N522, N252, N369);
and AND3 (N527, N510, N171, N426);
buf BUF1 (N528, N511);
buf BUF1 (N529, N512);
xor XOR2 (N530, N523, N299);
buf BUF1 (N531, N518);
or OR4 (N532, N520, N383, N205, N509);
buf BUF1 (N533, N524);
nand NAND4 (N534, N530, N85, N242, N99);
nand NAND4 (N535, N525, N3, N286, N483);
buf BUF1 (N536, N535);
and AND3 (N537, N517, N242, N484);
or OR2 (N538, N537, N439);
or OR3 (N539, N527, N14, N371);
and AND2 (N540, N526, N366);
xor XOR2 (N541, N538, N168);
nand NAND4 (N542, N532, N142, N200, N374);
buf BUF1 (N543, N539);
not NOT1 (N544, N529);
nand NAND3 (N545, N540, N305, N239);
buf BUF1 (N546, N542);
nor NOR3 (N547, N534, N219, N302);
and AND3 (N548, N536, N276, N144);
xor XOR2 (N549, N544, N18);
nor NOR4 (N550, N533, N27, N498, N130);
not NOT1 (N551, N546);
nand NAND2 (N552, N549, N452);
buf BUF1 (N553, N541);
nand NAND2 (N554, N552, N374);
and AND3 (N555, N531, N246, N514);
buf BUF1 (N556, N545);
nand NAND2 (N557, N551, N235);
or OR3 (N558, N550, N153, N434);
not NOT1 (N559, N555);
not NOT1 (N560, N554);
nor NOR4 (N561, N557, N487, N175, N546);
not NOT1 (N562, N528);
or OR4 (N563, N556, N196, N430, N552);
or OR2 (N564, N558, N141);
and AND2 (N565, N562, N548);
and AND2 (N566, N8, N447);
nand NAND2 (N567, N561, N34);
xor XOR2 (N568, N559, N540);
not NOT1 (N569, N566);
or OR4 (N570, N553, N129, N301, N199);
buf BUF1 (N571, N547);
nand NAND4 (N572, N565, N476, N101, N191);
nor NOR2 (N573, N570, N380);
not NOT1 (N574, N563);
and AND4 (N575, N572, N205, N76, N228);
nor NOR2 (N576, N569, N134);
xor XOR2 (N577, N564, N16);
or OR2 (N578, N573, N245);
nand NAND3 (N579, N575, N568, N560);
nor NOR4 (N580, N165, N252, N98, N98);
or OR2 (N581, N250, N548);
xor XOR2 (N582, N543, N423);
not NOT1 (N583, N567);
and AND4 (N584, N582, N6, N62, N100);
nand NAND4 (N585, N574, N183, N534, N40);
and AND4 (N586, N585, N379, N200, N376);
xor XOR2 (N587, N580, N4);
xor XOR2 (N588, N576, N584);
not NOT1 (N589, N139);
and AND3 (N590, N571, N558, N84);
not NOT1 (N591, N577);
not NOT1 (N592, N581);
not NOT1 (N593, N592);
not NOT1 (N594, N588);
nor NOR3 (N595, N586, N371, N419);
xor XOR2 (N596, N583, N127);
not NOT1 (N597, N594);
or OR2 (N598, N595, N186);
and AND2 (N599, N578, N224);
nor NOR2 (N600, N589, N402);
not NOT1 (N601, N597);
or OR4 (N602, N601, N244, N592, N51);
and AND4 (N603, N593, N303, N560, N477);
or OR3 (N604, N591, N191, N443);
buf BUF1 (N605, N587);
xor XOR2 (N606, N579, N553);
nand NAND2 (N607, N590, N445);
xor XOR2 (N608, N599, N144);
nor NOR4 (N609, N605, N450, N533, N17);
nor NOR2 (N610, N604, N371);
nand NAND4 (N611, N607, N27, N389, N246);
nand NAND4 (N612, N598, N278, N448, N114);
buf BUF1 (N613, N596);
buf BUF1 (N614, N611);
nand NAND4 (N615, N609, N557, N250, N28);
xor XOR2 (N616, N613, N388);
or OR3 (N617, N610, N340, N274);
buf BUF1 (N618, N612);
buf BUF1 (N619, N602);
xor XOR2 (N620, N608, N199);
nand NAND4 (N621, N616, N527, N31, N206);
not NOT1 (N622, N617);
nand NAND2 (N623, N619, N346);
not NOT1 (N624, N621);
and AND2 (N625, N606, N396);
or OR2 (N626, N622, N427);
buf BUF1 (N627, N624);
and AND2 (N628, N623, N5);
xor XOR2 (N629, N620, N574);
not NOT1 (N630, N618);
xor XOR2 (N631, N626, N434);
nor NOR3 (N632, N629, N290, N470);
not NOT1 (N633, N625);
xor XOR2 (N634, N631, N436);
xor XOR2 (N635, N633, N60);
buf BUF1 (N636, N615);
buf BUF1 (N637, N603);
or OR3 (N638, N630, N29, N460);
nand NAND3 (N639, N627, N412, N358);
and AND2 (N640, N614, N68);
or OR3 (N641, N640, N265, N402);
nand NAND3 (N642, N634, N107, N65);
nand NAND4 (N643, N636, N308, N508, N432);
xor XOR2 (N644, N600, N97);
or OR2 (N645, N632, N460);
nor NOR2 (N646, N628, N124);
and AND2 (N647, N641, N16);
and AND4 (N648, N642, N516, N604, N583);
nor NOR4 (N649, N646, N101, N425, N188);
xor XOR2 (N650, N639, N226);
or OR4 (N651, N645, N123, N404, N416);
nor NOR4 (N652, N647, N422, N149, N78);
or OR2 (N653, N652, N413);
nand NAND4 (N654, N653, N366, N49, N588);
nand NAND4 (N655, N644, N208, N399, N276);
not NOT1 (N656, N649);
not NOT1 (N657, N651);
not NOT1 (N658, N655);
buf BUF1 (N659, N650);
nor NOR4 (N660, N648, N368, N128, N412);
buf BUF1 (N661, N635);
or OR3 (N662, N656, N658, N86);
and AND2 (N663, N61, N585);
buf BUF1 (N664, N654);
nand NAND3 (N665, N660, N417, N58);
nand NAND2 (N666, N643, N233);
buf BUF1 (N667, N661);
or OR3 (N668, N666, N198, N469);
nand NAND4 (N669, N663, N321, N444, N79);
nor NOR3 (N670, N667, N186, N140);
nand NAND3 (N671, N669, N389, N194);
nand NAND3 (N672, N659, N372, N154);
nor NOR3 (N673, N662, N559, N463);
nor NOR3 (N674, N657, N143, N24);
nand NAND3 (N675, N670, N86, N612);
buf BUF1 (N676, N673);
buf BUF1 (N677, N671);
xor XOR2 (N678, N672, N188);
nand NAND3 (N679, N665, N570, N536);
nor NOR2 (N680, N678, N611);
not NOT1 (N681, N677);
nand NAND2 (N682, N675, N467);
nor NOR4 (N683, N664, N513, N354, N626);
xor XOR2 (N684, N637, N281);
buf BUF1 (N685, N683);
xor XOR2 (N686, N679, N355);
buf BUF1 (N687, N680);
not NOT1 (N688, N674);
xor XOR2 (N689, N688, N30);
xor XOR2 (N690, N684, N67);
nand NAND4 (N691, N689, N24, N184, N405);
and AND3 (N692, N682, N335, N99);
and AND2 (N693, N676, N368);
nand NAND4 (N694, N638, N272, N285, N445);
nor NOR3 (N695, N692, N73, N130);
or OR2 (N696, N687, N183);
buf BUF1 (N697, N695);
nor NOR2 (N698, N668, N213);
nor NOR3 (N699, N693, N63, N182);
xor XOR2 (N700, N694, N465);
and AND4 (N701, N698, N434, N172, N389);
not NOT1 (N702, N699);
nor NOR4 (N703, N685, N439, N190, N673);
or OR4 (N704, N686, N603, N2, N444);
xor XOR2 (N705, N681, N407);
nor NOR2 (N706, N690, N545);
not NOT1 (N707, N702);
buf BUF1 (N708, N704);
xor XOR2 (N709, N703, N143);
buf BUF1 (N710, N696);
or OR2 (N711, N710, N436);
nor NOR4 (N712, N706, N204, N213, N26);
and AND4 (N713, N712, N462, N323, N472);
and AND3 (N714, N709, N355, N536);
and AND4 (N715, N700, N610, N382, N636);
or OR3 (N716, N701, N472, N315);
xor XOR2 (N717, N713, N402);
not NOT1 (N718, N705);
and AND4 (N719, N718, N494, N665, N331);
or OR2 (N720, N711, N51);
and AND3 (N721, N716, N268, N88);
or OR2 (N722, N720, N322);
nand NAND3 (N723, N697, N126, N522);
or OR4 (N724, N723, N515, N656, N284);
buf BUF1 (N725, N714);
not NOT1 (N726, N715);
not NOT1 (N727, N719);
buf BUF1 (N728, N724);
buf BUF1 (N729, N721);
not NOT1 (N730, N722);
buf BUF1 (N731, N691);
not NOT1 (N732, N727);
or OR2 (N733, N726, N13);
or OR3 (N734, N729, N694, N107);
xor XOR2 (N735, N734, N489);
and AND2 (N736, N730, N313);
nand NAND4 (N737, N731, N730, N734, N659);
nor NOR3 (N738, N708, N267, N122);
xor XOR2 (N739, N736, N20);
not NOT1 (N740, N733);
not NOT1 (N741, N725);
xor XOR2 (N742, N738, N41);
or OR2 (N743, N717, N426);
xor XOR2 (N744, N728, N651);
xor XOR2 (N745, N737, N361);
buf BUF1 (N746, N740);
or OR2 (N747, N742, N107);
nor NOR2 (N748, N707, N665);
nor NOR3 (N749, N744, N46, N89);
buf BUF1 (N750, N732);
not NOT1 (N751, N735);
buf BUF1 (N752, N751);
and AND2 (N753, N750, N581);
nor NOR3 (N754, N753, N661, N13);
and AND3 (N755, N745, N374, N329);
not NOT1 (N756, N746);
xor XOR2 (N757, N754, N55);
nor NOR4 (N758, N743, N675, N130, N308);
buf BUF1 (N759, N747);
not NOT1 (N760, N758);
nand NAND4 (N761, N760, N606, N68, N78);
and AND2 (N762, N741, N150);
nand NAND4 (N763, N739, N205, N230, N627);
not NOT1 (N764, N748);
xor XOR2 (N765, N763, N310);
nor NOR3 (N766, N762, N395, N525);
not NOT1 (N767, N752);
xor XOR2 (N768, N749, N540);
nand NAND3 (N769, N766, N474, N701);
and AND3 (N770, N757, N436, N440);
nand NAND4 (N771, N770, N214, N97, N264);
nand NAND2 (N772, N755, N63);
nand NAND3 (N773, N759, N276, N496);
nand NAND2 (N774, N756, N132);
and AND4 (N775, N765, N587, N124, N237);
nand NAND4 (N776, N775, N633, N141, N380);
or OR3 (N777, N774, N275, N14);
xor XOR2 (N778, N768, N614);
and AND2 (N779, N776, N419);
buf BUF1 (N780, N773);
and AND3 (N781, N761, N67, N143);
and AND4 (N782, N779, N553, N408, N771);
nand NAND3 (N783, N706, N668, N69);
nor NOR2 (N784, N780, N309);
buf BUF1 (N785, N782);
xor XOR2 (N786, N778, N466);
buf BUF1 (N787, N764);
or OR3 (N788, N767, N140, N17);
nor NOR4 (N789, N785, N403, N90, N453);
not NOT1 (N790, N781);
nand NAND3 (N791, N789, N644, N628);
xor XOR2 (N792, N786, N620);
nor NOR2 (N793, N787, N686);
or OR4 (N794, N793, N192, N582, N556);
or OR4 (N795, N792, N763, N651, N337);
buf BUF1 (N796, N794);
or OR3 (N797, N796, N515, N57);
and AND2 (N798, N790, N713);
nor NOR3 (N799, N788, N532, N293);
nand NAND3 (N800, N772, N166, N137);
or OR4 (N801, N777, N549, N89, N370);
not NOT1 (N802, N783);
xor XOR2 (N803, N799, N216);
nand NAND4 (N804, N791, N365, N38, N542);
buf BUF1 (N805, N804);
not NOT1 (N806, N769);
or OR3 (N807, N806, N118, N24);
nand NAND4 (N808, N795, N157, N557, N453);
xor XOR2 (N809, N801, N12);
and AND2 (N810, N807, N84);
not NOT1 (N811, N802);
or OR2 (N812, N797, N156);
nor NOR3 (N813, N784, N336, N751);
nor NOR3 (N814, N812, N721, N324);
xor XOR2 (N815, N800, N96);
not NOT1 (N816, N815);
not NOT1 (N817, N803);
nand NAND4 (N818, N809, N174, N265, N551);
nor NOR2 (N819, N798, N2);
and AND3 (N820, N813, N654, N497);
nand NAND4 (N821, N810, N379, N697, N728);
buf BUF1 (N822, N811);
nor NOR2 (N823, N822, N784);
nor NOR2 (N824, N823, N281);
nor NOR3 (N825, N819, N674, N202);
and AND2 (N826, N814, N620);
xor XOR2 (N827, N826, N596);
nor NOR3 (N828, N816, N219, N193);
or OR3 (N829, N808, N382, N83);
buf BUF1 (N830, N828);
and AND4 (N831, N824, N470, N717, N357);
buf BUF1 (N832, N827);
nand NAND4 (N833, N831, N455, N687, N799);
nand NAND2 (N834, N821, N6);
or OR4 (N835, N830, N172, N707, N633);
nor NOR4 (N836, N820, N412, N624, N283);
xor XOR2 (N837, N835, N324);
and AND4 (N838, N836, N409, N255, N530);
or OR4 (N839, N817, N659, N240, N795);
xor XOR2 (N840, N838, N559);
not NOT1 (N841, N825);
not NOT1 (N842, N841);
buf BUF1 (N843, N834);
and AND3 (N844, N840, N313, N556);
and AND2 (N845, N805, N161);
nor NOR2 (N846, N839, N837);
not NOT1 (N847, N555);
not NOT1 (N848, N843);
buf BUF1 (N849, N842);
nor NOR2 (N850, N818, N154);
xor XOR2 (N851, N832, N8);
buf BUF1 (N852, N833);
or OR2 (N853, N849, N806);
not NOT1 (N854, N829);
xor XOR2 (N855, N852, N352);
buf BUF1 (N856, N851);
nand NAND2 (N857, N845, N481);
nor NOR4 (N858, N856, N830, N181, N33);
nor NOR2 (N859, N854, N824);
not NOT1 (N860, N858);
or OR4 (N861, N850, N814, N535, N170);
and AND2 (N862, N859, N26);
nor NOR4 (N863, N857, N59, N699, N451);
or OR3 (N864, N862, N616, N357);
not NOT1 (N865, N863);
not NOT1 (N866, N848);
nor NOR2 (N867, N855, N133);
and AND4 (N868, N867, N493, N243, N460);
buf BUF1 (N869, N860);
xor XOR2 (N870, N853, N31);
or OR4 (N871, N870, N606, N826, N116);
and AND3 (N872, N844, N260, N780);
nor NOR2 (N873, N861, N305);
and AND3 (N874, N873, N77, N425);
buf BUF1 (N875, N869);
nand NAND3 (N876, N866, N235, N546);
and AND2 (N877, N864, N259);
nor NOR4 (N878, N846, N136, N506, N874);
nand NAND2 (N879, N610, N699);
nand NAND4 (N880, N875, N745, N376, N170);
not NOT1 (N881, N871);
not NOT1 (N882, N872);
nor NOR3 (N883, N847, N683, N754);
not NOT1 (N884, N878);
nand NAND4 (N885, N881, N131, N779, N537);
or OR4 (N886, N885, N196, N843, N116);
or OR4 (N887, N865, N68, N437, N458);
buf BUF1 (N888, N876);
buf BUF1 (N889, N883);
and AND2 (N890, N879, N339);
xor XOR2 (N891, N887, N173);
or OR2 (N892, N877, N241);
and AND4 (N893, N882, N272, N476, N333);
nor NOR4 (N894, N886, N206, N110, N114);
nor NOR3 (N895, N880, N113, N715);
nand NAND4 (N896, N895, N835, N781, N257);
xor XOR2 (N897, N894, N272);
nand NAND2 (N898, N889, N60);
nor NOR4 (N899, N891, N745, N156, N111);
not NOT1 (N900, N892);
xor XOR2 (N901, N884, N546);
nor NOR4 (N902, N888, N611, N255, N248);
buf BUF1 (N903, N902);
nor NOR4 (N904, N900, N259, N895, N801);
buf BUF1 (N905, N901);
buf BUF1 (N906, N896);
nor NOR3 (N907, N903, N78, N823);
not NOT1 (N908, N898);
and AND4 (N909, N907, N382, N743, N879);
nand NAND2 (N910, N909, N151);
nand NAND4 (N911, N893, N296, N279, N739);
not NOT1 (N912, N904);
not NOT1 (N913, N908);
and AND4 (N914, N913, N818, N766, N892);
buf BUF1 (N915, N899);
nor NOR2 (N916, N915, N596);
buf BUF1 (N917, N910);
not NOT1 (N918, N897);
xor XOR2 (N919, N917, N868);
and AND3 (N920, N831, N8, N513);
buf BUF1 (N921, N911);
nand NAND3 (N922, N918, N257, N191);
and AND3 (N923, N905, N456, N529);
not NOT1 (N924, N921);
nand NAND3 (N925, N890, N118, N618);
not NOT1 (N926, N925);
or OR4 (N927, N916, N653, N786, N554);
and AND2 (N928, N920, N745);
not NOT1 (N929, N922);
or OR3 (N930, N906, N336, N910);
nor NOR3 (N931, N924, N534, N610);
buf BUF1 (N932, N926);
xor XOR2 (N933, N929, N802);
buf BUF1 (N934, N912);
xor XOR2 (N935, N914, N673);
nor NOR4 (N936, N919, N34, N683, N859);
nand NAND2 (N937, N936, N870);
nand NAND4 (N938, N935, N891, N533, N184);
and AND3 (N939, N931, N841, N584);
nand NAND3 (N940, N939, N434, N254);
xor XOR2 (N941, N927, N441);
buf BUF1 (N942, N940);
nand NAND2 (N943, N933, N729);
and AND3 (N944, N943, N77, N942);
xor XOR2 (N945, N429, N914);
and AND2 (N946, N938, N368);
nor NOR3 (N947, N930, N84, N481);
buf BUF1 (N948, N941);
or OR2 (N949, N923, N307);
and AND3 (N950, N934, N817, N205);
nor NOR3 (N951, N937, N77, N941);
nand NAND4 (N952, N945, N45, N896, N666);
xor XOR2 (N953, N932, N593);
nand NAND3 (N954, N944, N806, N67);
buf BUF1 (N955, N950);
xor XOR2 (N956, N953, N35);
nand NAND3 (N957, N928, N944, N297);
buf BUF1 (N958, N952);
buf BUF1 (N959, N951);
xor XOR2 (N960, N949, N336);
buf BUF1 (N961, N955);
not NOT1 (N962, N961);
nor NOR4 (N963, N946, N767, N862, N236);
nand NAND2 (N964, N959, N259);
not NOT1 (N965, N956);
xor XOR2 (N966, N963, N439);
buf BUF1 (N967, N964);
nor NOR3 (N968, N966, N186, N830);
not NOT1 (N969, N947);
or OR2 (N970, N967, N291);
or OR2 (N971, N962, N426);
or OR3 (N972, N970, N638, N21);
xor XOR2 (N973, N948, N730);
not NOT1 (N974, N954);
xor XOR2 (N975, N957, N422);
nor NOR3 (N976, N969, N125, N82);
or OR2 (N977, N965, N255);
buf BUF1 (N978, N968);
nand NAND4 (N979, N974, N111, N329, N570);
buf BUF1 (N980, N972);
nand NAND4 (N981, N976, N175, N231, N797);
and AND3 (N982, N960, N879, N243);
or OR2 (N983, N980, N243);
not NOT1 (N984, N975);
nand NAND4 (N985, N958, N977, N258, N927);
not NOT1 (N986, N900);
and AND4 (N987, N982, N937, N317, N923);
or OR4 (N988, N971, N460, N226, N986);
nand NAND4 (N989, N933, N86, N869, N447);
nand NAND3 (N990, N984, N556, N26);
and AND4 (N991, N978, N971, N134, N861);
nor NOR3 (N992, N987, N927, N980);
xor XOR2 (N993, N990, N864);
buf BUF1 (N994, N992);
nor NOR3 (N995, N983, N62, N680);
xor XOR2 (N996, N993, N103);
not NOT1 (N997, N991);
xor XOR2 (N998, N985, N703);
buf BUF1 (N999, N995);
buf BUF1 (N1000, N981);
buf BUF1 (N1001, N1000);
buf BUF1 (N1002, N999);
buf BUF1 (N1003, N996);
or OR3 (N1004, N994, N895, N555);
xor XOR2 (N1005, N998, N898);
nand NAND4 (N1006, N1001, N36, N751, N316);
or OR4 (N1007, N973, N774, N212, N630);
nor NOR4 (N1008, N979, N102, N698, N906);
and AND2 (N1009, N997, N805);
xor XOR2 (N1010, N1004, N665);
xor XOR2 (N1011, N1009, N17);
buf BUF1 (N1012, N1005);
nor NOR3 (N1013, N1011, N158, N32);
and AND3 (N1014, N989, N656, N578);
xor XOR2 (N1015, N1012, N934);
nor NOR4 (N1016, N1006, N1006, N140, N859);
buf BUF1 (N1017, N988);
or OR3 (N1018, N1002, N523, N39);
not NOT1 (N1019, N1018);
and AND4 (N1020, N1008, N612, N112, N403);
not NOT1 (N1021, N1010);
nor NOR2 (N1022, N1021, N761);
xor XOR2 (N1023, N1022, N461);
nor NOR2 (N1024, N1017, N914);
buf BUF1 (N1025, N1019);
and AND2 (N1026, N1025, N808);
or OR2 (N1027, N1013, N485);
and AND3 (N1028, N1016, N843, N203);
nand NAND3 (N1029, N1003, N1015, N805);
and AND2 (N1030, N862, N505);
or OR2 (N1031, N1029, N720);
not NOT1 (N1032, N1030);
or OR4 (N1033, N1027, N988, N116, N347);
nand NAND3 (N1034, N1020, N832, N498);
nor NOR3 (N1035, N1023, N1019, N1016);
buf BUF1 (N1036, N1035);
or OR2 (N1037, N1024, N711);
nor NOR3 (N1038, N1014, N135, N334);
and AND2 (N1039, N1031, N35);
and AND4 (N1040, N1037, N29, N23, N19);
and AND3 (N1041, N1038, N697, N451);
and AND3 (N1042, N1034, N436, N628);
buf BUF1 (N1043, N1028);
and AND4 (N1044, N1036, N936, N900, N10);
or OR3 (N1045, N1042, N825, N349);
not NOT1 (N1046, N1026);
buf BUF1 (N1047, N1044);
xor XOR2 (N1048, N1041, N8);
not NOT1 (N1049, N1047);
or OR3 (N1050, N1040, N338, N111);
not NOT1 (N1051, N1043);
nor NOR2 (N1052, N1045, N578);
buf BUF1 (N1053, N1051);
not NOT1 (N1054, N1007);
or OR2 (N1055, N1032, N464);
nor NOR4 (N1056, N1050, N25, N517, N120);
and AND3 (N1057, N1054, N911, N676);
not NOT1 (N1058, N1055);
and AND2 (N1059, N1048, N480);
nor NOR4 (N1060, N1049, N570, N592, N200);
nor NOR4 (N1061, N1060, N185, N104, N632);
or OR2 (N1062, N1052, N454);
or OR2 (N1063, N1033, N679);
buf BUF1 (N1064, N1061);
or OR4 (N1065, N1046, N1018, N870, N777);
nor NOR4 (N1066, N1062, N593, N896, N821);
and AND2 (N1067, N1039, N794);
and AND2 (N1068, N1057, N57);
and AND4 (N1069, N1058, N841, N194, N555);
nand NAND3 (N1070, N1068, N538, N588);
nor NOR4 (N1071, N1063, N118, N400, N82);
or OR2 (N1072, N1056, N466);
nand NAND3 (N1073, N1066, N878, N228);
and AND3 (N1074, N1064, N180, N43);
buf BUF1 (N1075, N1070);
nor NOR3 (N1076, N1075, N1023, N988);
nor NOR4 (N1077, N1071, N267, N863, N951);
nor NOR2 (N1078, N1076, N313);
nand NAND4 (N1079, N1065, N113, N546, N816);
nor NOR4 (N1080, N1072, N433, N688, N445);
xor XOR2 (N1081, N1079, N200);
not NOT1 (N1082, N1067);
and AND4 (N1083, N1073, N37, N607, N1001);
buf BUF1 (N1084, N1082);
nor NOR3 (N1085, N1081, N569, N896);
buf BUF1 (N1086, N1074);
nor NOR2 (N1087, N1086, N634);
nand NAND4 (N1088, N1053, N193, N875, N585);
nand NAND3 (N1089, N1088, N1014, N285);
or OR2 (N1090, N1083, N72);
xor XOR2 (N1091, N1084, N485);
nand NAND4 (N1092, N1059, N194, N520, N1066);
and AND4 (N1093, N1069, N749, N347, N519);
xor XOR2 (N1094, N1085, N828);
nor NOR2 (N1095, N1078, N1073);
nand NAND3 (N1096, N1094, N946, N288);
nand NAND3 (N1097, N1090, N273, N798);
nand NAND4 (N1098, N1077, N45, N194, N706);
and AND2 (N1099, N1080, N516);
or OR2 (N1100, N1087, N315);
buf BUF1 (N1101, N1089);
nand NAND3 (N1102, N1099, N183, N544);
buf BUF1 (N1103, N1095);
xor XOR2 (N1104, N1100, N181);
or OR4 (N1105, N1103, N776, N464, N132);
xor XOR2 (N1106, N1104, N582);
nor NOR4 (N1107, N1096, N123, N543, N150);
and AND3 (N1108, N1101, N922, N1094);
not NOT1 (N1109, N1092);
not NOT1 (N1110, N1108);
xor XOR2 (N1111, N1098, N121);
nand NAND3 (N1112, N1109, N1007, N941);
nor NOR2 (N1113, N1111, N485);
nor NOR4 (N1114, N1110, N674, N379, N156);
nor NOR4 (N1115, N1097, N783, N496, N214);
not NOT1 (N1116, N1102);
nand NAND4 (N1117, N1113, N98, N1106, N177);
not NOT1 (N1118, N125);
buf BUF1 (N1119, N1114);
not NOT1 (N1120, N1115);
nand NAND4 (N1121, N1119, N996, N973, N218);
xor XOR2 (N1122, N1118, N556);
or OR4 (N1123, N1093, N282, N968, N659);
buf BUF1 (N1124, N1123);
not NOT1 (N1125, N1116);
buf BUF1 (N1126, N1124);
nor NOR2 (N1127, N1120, N317);
or OR4 (N1128, N1121, N641, N214, N142);
not NOT1 (N1129, N1117);
nor NOR4 (N1130, N1125, N166, N602, N65);
or OR4 (N1131, N1128, N102, N487, N964);
or OR3 (N1132, N1107, N353, N61);
buf BUF1 (N1133, N1130);
nor NOR3 (N1134, N1133, N202, N630);
nand NAND3 (N1135, N1131, N532, N53);
buf BUF1 (N1136, N1112);
or OR3 (N1137, N1136, N925, N1033);
nand NAND4 (N1138, N1122, N860, N296, N500);
buf BUF1 (N1139, N1126);
buf BUF1 (N1140, N1091);
not NOT1 (N1141, N1105);
nand NAND2 (N1142, N1137, N776);
or OR4 (N1143, N1138, N983, N769, N747);
or OR3 (N1144, N1141, N647, N481);
not NOT1 (N1145, N1134);
nand NAND2 (N1146, N1145, N802);
or OR2 (N1147, N1146, N802);
nor NOR4 (N1148, N1142, N275, N568, N116);
or OR4 (N1149, N1139, N1070, N913, N1061);
xor XOR2 (N1150, N1140, N194);
not NOT1 (N1151, N1148);
xor XOR2 (N1152, N1147, N306);
nor NOR4 (N1153, N1150, N824, N422, N996);
and AND4 (N1154, N1152, N1119, N1019, N1026);
buf BUF1 (N1155, N1149);
xor XOR2 (N1156, N1151, N660);
not NOT1 (N1157, N1153);
not NOT1 (N1158, N1135);
or OR3 (N1159, N1132, N53, N501);
or OR2 (N1160, N1155, N846);
or OR2 (N1161, N1144, N1037);
and AND4 (N1162, N1156, N713, N212, N403);
not NOT1 (N1163, N1127);
and AND3 (N1164, N1163, N722, N525);
or OR3 (N1165, N1154, N578, N550);
xor XOR2 (N1166, N1164, N1076);
and AND3 (N1167, N1165, N845, N826);
nand NAND4 (N1168, N1162, N307, N36, N604);
buf BUF1 (N1169, N1157);
and AND4 (N1170, N1158, N835, N883, N668);
nor NOR3 (N1171, N1166, N343, N979);
xor XOR2 (N1172, N1168, N1147);
nor NOR2 (N1173, N1129, N557);
not NOT1 (N1174, N1170);
nor NOR2 (N1175, N1174, N945);
xor XOR2 (N1176, N1172, N357);
and AND3 (N1177, N1160, N1109, N880);
nand NAND2 (N1178, N1143, N1177);
not NOT1 (N1179, N959);
and AND2 (N1180, N1176, N1052);
nor NOR2 (N1181, N1173, N272);
not NOT1 (N1182, N1180);
nand NAND4 (N1183, N1161, N957, N241, N1065);
nand NAND2 (N1184, N1182, N588);
nand NAND2 (N1185, N1175, N148);
xor XOR2 (N1186, N1167, N1081);
nor NOR2 (N1187, N1181, N176);
nand NAND2 (N1188, N1169, N1082);
nand NAND2 (N1189, N1183, N866);
and AND4 (N1190, N1159, N115, N491, N783);
and AND4 (N1191, N1187, N727, N459, N353);
and AND4 (N1192, N1188, N137, N222, N710);
nor NOR4 (N1193, N1186, N373, N71, N581);
and AND3 (N1194, N1185, N6, N137);
nand NAND3 (N1195, N1193, N481, N731);
nor NOR4 (N1196, N1189, N554, N789, N403);
or OR2 (N1197, N1195, N883);
nor NOR4 (N1198, N1171, N317, N55, N60);
buf BUF1 (N1199, N1198);
nand NAND4 (N1200, N1197, N402, N844, N1146);
nor NOR2 (N1201, N1196, N429);
or OR2 (N1202, N1191, N505);
xor XOR2 (N1203, N1201, N784);
not NOT1 (N1204, N1190);
not NOT1 (N1205, N1203);
not NOT1 (N1206, N1200);
nand NAND3 (N1207, N1179, N414, N1059);
not NOT1 (N1208, N1178);
buf BUF1 (N1209, N1207);
buf BUF1 (N1210, N1184);
not NOT1 (N1211, N1204);
or OR2 (N1212, N1210, N897);
xor XOR2 (N1213, N1212, N1182);
nand NAND4 (N1214, N1199, N296, N876, N204);
nor NOR3 (N1215, N1213, N963, N759);
xor XOR2 (N1216, N1206, N669);
nor NOR2 (N1217, N1205, N1178);
and AND4 (N1218, N1216, N138, N560, N882);
xor XOR2 (N1219, N1209, N1099);
and AND3 (N1220, N1219, N384, N1210);
and AND4 (N1221, N1218, N1137, N977, N236);
nand NAND2 (N1222, N1221, N403);
and AND4 (N1223, N1192, N539, N862, N316);
and AND4 (N1224, N1215, N655, N1020, N1155);
nor NOR3 (N1225, N1220, N950, N178);
nand NAND4 (N1226, N1202, N1084, N661, N454);
and AND3 (N1227, N1226, N272, N1096);
not NOT1 (N1228, N1194);
xor XOR2 (N1229, N1228, N757);
nor NOR3 (N1230, N1211, N1118, N1076);
nand NAND3 (N1231, N1222, N757, N377);
nor NOR3 (N1232, N1217, N102, N290);
and AND3 (N1233, N1232, N1037, N1100);
or OR4 (N1234, N1230, N1218, N378, N727);
nand NAND4 (N1235, N1227, N981, N47, N373);
or OR3 (N1236, N1223, N356, N29);
not NOT1 (N1237, N1234);
buf BUF1 (N1238, N1237);
xor XOR2 (N1239, N1224, N284);
nand NAND2 (N1240, N1233, N278);
nor NOR3 (N1241, N1235, N1000, N54);
nand NAND4 (N1242, N1240, N1030, N735, N949);
nor NOR4 (N1243, N1231, N729, N10, N918);
or OR4 (N1244, N1242, N1142, N725, N1057);
not NOT1 (N1245, N1208);
not NOT1 (N1246, N1229);
and AND2 (N1247, N1246, N620);
nor NOR4 (N1248, N1238, N249, N655, N163);
buf BUF1 (N1249, N1243);
not NOT1 (N1250, N1241);
nand NAND2 (N1251, N1236, N19);
and AND2 (N1252, N1249, N358);
and AND4 (N1253, N1244, N354, N987, N12);
or OR4 (N1254, N1214, N329, N118, N1023);
or OR4 (N1255, N1225, N1106, N1223, N330);
and AND2 (N1256, N1255, N106);
nor NOR2 (N1257, N1256, N850);
or OR4 (N1258, N1247, N92, N319, N1050);
buf BUF1 (N1259, N1250);
or OR4 (N1260, N1248, N1024, N1034, N177);
xor XOR2 (N1261, N1258, N694);
and AND3 (N1262, N1239, N797, N303);
or OR2 (N1263, N1259, N279);
nor NOR2 (N1264, N1261, N812);
nor NOR4 (N1265, N1252, N643, N786, N1169);
nor NOR4 (N1266, N1253, N1126, N142, N25);
xor XOR2 (N1267, N1245, N533);
or OR4 (N1268, N1265, N847, N469, N821);
or OR3 (N1269, N1262, N1138, N724);
buf BUF1 (N1270, N1268);
or OR3 (N1271, N1264, N882, N20);
or OR2 (N1272, N1271, N894);
nor NOR3 (N1273, N1270, N388, N1129);
nand NAND3 (N1274, N1254, N616, N892);
nor NOR2 (N1275, N1251, N998);
or OR2 (N1276, N1267, N398);
nand NAND2 (N1277, N1276, N939);
not NOT1 (N1278, N1260);
not NOT1 (N1279, N1272);
nor NOR3 (N1280, N1269, N1040, N351);
xor XOR2 (N1281, N1263, N1124);
and AND2 (N1282, N1281, N203);
nor NOR4 (N1283, N1282, N308, N309, N111);
and AND3 (N1284, N1279, N1190, N783);
xor XOR2 (N1285, N1274, N1160);
not NOT1 (N1286, N1275);
xor XOR2 (N1287, N1284, N385);
xor XOR2 (N1288, N1285, N407);
or OR2 (N1289, N1283, N720);
buf BUF1 (N1290, N1289);
buf BUF1 (N1291, N1287);
nand NAND2 (N1292, N1273, N191);
nor NOR3 (N1293, N1288, N324, N1050);
buf BUF1 (N1294, N1278);
buf BUF1 (N1295, N1266);
not NOT1 (N1296, N1294);
nand NAND3 (N1297, N1280, N205, N293);
not NOT1 (N1298, N1293);
or OR3 (N1299, N1290, N1093, N619);
nand NAND4 (N1300, N1277, N1138, N1251, N944);
buf BUF1 (N1301, N1300);
not NOT1 (N1302, N1299);
and AND4 (N1303, N1301, N501, N500, N159);
and AND4 (N1304, N1298, N714, N910, N850);
xor XOR2 (N1305, N1295, N1269);
and AND2 (N1306, N1291, N1118);
and AND4 (N1307, N1304, N343, N1066, N617);
buf BUF1 (N1308, N1307);
nor NOR4 (N1309, N1257, N1084, N318, N972);
xor XOR2 (N1310, N1306, N334);
not NOT1 (N1311, N1305);
not NOT1 (N1312, N1309);
or OR2 (N1313, N1292, N677);
xor XOR2 (N1314, N1302, N928);
or OR2 (N1315, N1313, N52);
xor XOR2 (N1316, N1312, N1);
and AND2 (N1317, N1316, N1035);
nand NAND3 (N1318, N1317, N750, N600);
nand NAND4 (N1319, N1286, N1150, N440, N261);
and AND2 (N1320, N1311, N937);
nor NOR4 (N1321, N1310, N477, N818, N1255);
xor XOR2 (N1322, N1319, N41);
xor XOR2 (N1323, N1318, N1205);
nor NOR2 (N1324, N1308, N670);
nand NAND3 (N1325, N1303, N906, N1250);
xor XOR2 (N1326, N1297, N714);
nand NAND2 (N1327, N1326, N1066);
xor XOR2 (N1328, N1314, N592);
nor NOR2 (N1329, N1325, N523);
nor NOR2 (N1330, N1320, N922);
or OR4 (N1331, N1324, N1137, N32, N124);
buf BUF1 (N1332, N1322);
nand NAND2 (N1333, N1315, N1080);
and AND2 (N1334, N1329, N1280);
not NOT1 (N1335, N1327);
nor NOR4 (N1336, N1330, N1118, N1245, N1140);
not NOT1 (N1337, N1336);
buf BUF1 (N1338, N1323);
xor XOR2 (N1339, N1321, N742);
buf BUF1 (N1340, N1331);
and AND3 (N1341, N1333, N889, N906);
and AND3 (N1342, N1334, N866, N1156);
nand NAND4 (N1343, N1342, N803, N117, N1302);
nand NAND4 (N1344, N1335, N1304, N835, N605);
xor XOR2 (N1345, N1332, N1253);
not NOT1 (N1346, N1343);
or OR2 (N1347, N1341, N784);
nand NAND4 (N1348, N1346, N668, N361, N674);
xor XOR2 (N1349, N1296, N645);
xor XOR2 (N1350, N1339, N714);
xor XOR2 (N1351, N1338, N1181);
and AND4 (N1352, N1349, N1033, N324, N129);
or OR2 (N1353, N1328, N504);
xor XOR2 (N1354, N1352, N262);
buf BUF1 (N1355, N1347);
nor NOR3 (N1356, N1340, N370, N217);
nand NAND2 (N1357, N1354, N984);
and AND4 (N1358, N1357, N992, N890, N501);
not NOT1 (N1359, N1344);
buf BUF1 (N1360, N1353);
buf BUF1 (N1361, N1360);
and AND3 (N1362, N1355, N1008, N99);
xor XOR2 (N1363, N1351, N400);
and AND3 (N1364, N1350, N551, N488);
xor XOR2 (N1365, N1337, N1179);
nand NAND2 (N1366, N1359, N421);
and AND4 (N1367, N1363, N422, N241, N221);
xor XOR2 (N1368, N1345, N769);
nand NAND2 (N1369, N1368, N947);
and AND3 (N1370, N1364, N246, N84);
buf BUF1 (N1371, N1356);
nand NAND4 (N1372, N1348, N457, N1198, N997);
buf BUF1 (N1373, N1371);
or OR4 (N1374, N1367, N221, N233, N98);
nor NOR4 (N1375, N1374, N1082, N645, N758);
not NOT1 (N1376, N1362);
nor NOR2 (N1377, N1376, N66);
or OR3 (N1378, N1358, N490, N803);
and AND2 (N1379, N1361, N492);
xor XOR2 (N1380, N1369, N461);
buf BUF1 (N1381, N1373);
or OR2 (N1382, N1370, N533);
nand NAND4 (N1383, N1379, N870, N935, N1121);
or OR2 (N1384, N1380, N807);
and AND4 (N1385, N1384, N960, N626, N1052);
and AND2 (N1386, N1366, N1012);
xor XOR2 (N1387, N1378, N443);
and AND2 (N1388, N1372, N326);
xor XOR2 (N1389, N1383, N184);
xor XOR2 (N1390, N1365, N1372);
and AND4 (N1391, N1388, N1107, N138, N1114);
nand NAND2 (N1392, N1381, N950);
nor NOR4 (N1393, N1391, N1047, N770, N567);
nand NAND4 (N1394, N1385, N432, N477, N334);
or OR4 (N1395, N1390, N58, N1185, N1069);
buf BUF1 (N1396, N1393);
xor XOR2 (N1397, N1375, N625);
nand NAND3 (N1398, N1397, N1158, N861);
nor NOR2 (N1399, N1398, N357);
or OR4 (N1400, N1396, N165, N12, N399);
or OR3 (N1401, N1392, N1364, N972);
nand NAND2 (N1402, N1386, N59);
not NOT1 (N1403, N1377);
xor XOR2 (N1404, N1400, N9);
nor NOR4 (N1405, N1389, N230, N829, N42);
nor NOR4 (N1406, N1401, N993, N909, N1134);
nor NOR4 (N1407, N1394, N58, N93, N1069);
buf BUF1 (N1408, N1407);
not NOT1 (N1409, N1402);
or OR3 (N1410, N1409, N838, N679);
nor NOR3 (N1411, N1403, N767, N1371);
buf BUF1 (N1412, N1410);
buf BUF1 (N1413, N1412);
or OR3 (N1414, N1408, N570, N27);
buf BUF1 (N1415, N1399);
xor XOR2 (N1416, N1404, N428);
nor NOR2 (N1417, N1416, N1116);
xor XOR2 (N1418, N1405, N898);
or OR4 (N1419, N1415, N990, N1056, N191);
nor NOR2 (N1420, N1417, N500);
buf BUF1 (N1421, N1413);
or OR2 (N1422, N1421, N1069);
nand NAND3 (N1423, N1411, N1261, N598);
buf BUF1 (N1424, N1382);
or OR3 (N1425, N1406, N86, N270);
or OR3 (N1426, N1419, N1370, N207);
buf BUF1 (N1427, N1423);
nand NAND2 (N1428, N1414, N546);
and AND2 (N1429, N1427, N1186);
not NOT1 (N1430, N1424);
buf BUF1 (N1431, N1425);
nor NOR3 (N1432, N1387, N464, N236);
or OR2 (N1433, N1429, N86);
not NOT1 (N1434, N1426);
and AND3 (N1435, N1428, N734, N705);
or OR2 (N1436, N1430, N960);
or OR2 (N1437, N1436, N1062);
not NOT1 (N1438, N1433);
buf BUF1 (N1439, N1438);
xor XOR2 (N1440, N1422, N710);
nand NAND2 (N1441, N1439, N418);
xor XOR2 (N1442, N1418, N1080);
not NOT1 (N1443, N1440);
xor XOR2 (N1444, N1395, N890);
xor XOR2 (N1445, N1443, N224);
nor NOR4 (N1446, N1445, N964, N1365, N829);
nand NAND3 (N1447, N1437, N761, N335);
nor NOR2 (N1448, N1434, N12);
nand NAND4 (N1449, N1431, N966, N204, N990);
not NOT1 (N1450, N1442);
xor XOR2 (N1451, N1435, N1202);
or OR3 (N1452, N1448, N231, N592);
not NOT1 (N1453, N1451);
not NOT1 (N1454, N1444);
or OR2 (N1455, N1420, N1120);
not NOT1 (N1456, N1453);
buf BUF1 (N1457, N1441);
nor NOR4 (N1458, N1452, N8, N34, N307);
buf BUF1 (N1459, N1458);
buf BUF1 (N1460, N1459);
and AND4 (N1461, N1456, N1293, N242, N274);
nand NAND4 (N1462, N1461, N194, N1452, N1110);
buf BUF1 (N1463, N1449);
buf BUF1 (N1464, N1447);
buf BUF1 (N1465, N1450);
not NOT1 (N1466, N1457);
not NOT1 (N1467, N1463);
not NOT1 (N1468, N1464);
buf BUF1 (N1469, N1468);
and AND4 (N1470, N1466, N1069, N860, N861);
nor NOR3 (N1471, N1467, N600, N102);
or OR2 (N1472, N1455, N506);
nand NAND2 (N1473, N1469, N111);
or OR4 (N1474, N1470, N138, N1053, N133);
xor XOR2 (N1475, N1446, N13);
xor XOR2 (N1476, N1473, N883);
nand NAND4 (N1477, N1465, N492, N219, N256);
xor XOR2 (N1478, N1476, N546);
xor XOR2 (N1479, N1477, N98);
xor XOR2 (N1480, N1479, N1168);
nor NOR3 (N1481, N1474, N890, N654);
buf BUF1 (N1482, N1454);
and AND4 (N1483, N1481, N667, N1241, N1227);
buf BUF1 (N1484, N1475);
nor NOR3 (N1485, N1480, N570, N697);
nor NOR2 (N1486, N1485, N322);
nor NOR4 (N1487, N1484, N230, N388, N1337);
nand NAND4 (N1488, N1482, N1285, N1371, N463);
buf BUF1 (N1489, N1486);
nand NAND2 (N1490, N1432, N1391);
or OR4 (N1491, N1472, N439, N1446, N676);
not NOT1 (N1492, N1462);
nor NOR3 (N1493, N1488, N931, N718);
buf BUF1 (N1494, N1460);
xor XOR2 (N1495, N1492, N462);
or OR3 (N1496, N1493, N1200, N1032);
or OR3 (N1497, N1490, N509, N1460);
not NOT1 (N1498, N1489);
or OR4 (N1499, N1494, N859, N353, N332);
buf BUF1 (N1500, N1491);
not NOT1 (N1501, N1498);
nor NOR4 (N1502, N1497, N992, N878, N931);
xor XOR2 (N1503, N1500, N281);
and AND2 (N1504, N1483, N240);
or OR3 (N1505, N1487, N591, N410);
not NOT1 (N1506, N1503);
nor NOR2 (N1507, N1506, N1046);
and AND4 (N1508, N1499, N726, N1214, N404);
xor XOR2 (N1509, N1507, N381);
or OR2 (N1510, N1496, N1289);
nand NAND3 (N1511, N1502, N1446, N474);
not NOT1 (N1512, N1504);
nand NAND3 (N1513, N1512, N1079, N1112);
nor NOR4 (N1514, N1510, N1449, N1310, N1258);
not NOT1 (N1515, N1514);
buf BUF1 (N1516, N1513);
buf BUF1 (N1517, N1508);
nand NAND3 (N1518, N1471, N647, N1252);
nand NAND4 (N1519, N1501, N162, N602, N544);
nand NAND2 (N1520, N1519, N399);
and AND2 (N1521, N1515, N730);
nor NOR3 (N1522, N1516, N1136, N506);
buf BUF1 (N1523, N1520);
xor XOR2 (N1524, N1521, N1126);
not NOT1 (N1525, N1505);
nor NOR4 (N1526, N1522, N670, N225, N209);
xor XOR2 (N1527, N1524, N933);
xor XOR2 (N1528, N1478, N18);
nor NOR2 (N1529, N1517, N521);
not NOT1 (N1530, N1523);
nor NOR3 (N1531, N1525, N618, N513);
nor NOR4 (N1532, N1526, N937, N725, N901);
xor XOR2 (N1533, N1529, N186);
and AND4 (N1534, N1495, N1098, N848, N337);
or OR4 (N1535, N1533, N599, N921, N591);
buf BUF1 (N1536, N1511);
not NOT1 (N1537, N1535);
buf BUF1 (N1538, N1530);
not NOT1 (N1539, N1532);
not NOT1 (N1540, N1518);
nand NAND3 (N1541, N1539, N1509, N476);
not NOT1 (N1542, N621);
not NOT1 (N1543, N1531);
and AND4 (N1544, N1538, N611, N265, N719);
nor NOR3 (N1545, N1537, N402, N956);
nand NAND3 (N1546, N1534, N49, N1397);
or OR4 (N1547, N1544, N765, N1225, N1165);
not NOT1 (N1548, N1547);
buf BUF1 (N1549, N1546);
nand NAND4 (N1550, N1548, N670, N453, N968);
or OR2 (N1551, N1545, N960);
and AND2 (N1552, N1551, N1293);
nand NAND3 (N1553, N1543, N317, N490);
nand NAND3 (N1554, N1540, N959, N1163);
xor XOR2 (N1555, N1541, N1185);
nand NAND4 (N1556, N1528, N329, N837, N1414);
nor NOR2 (N1557, N1552, N464);
buf BUF1 (N1558, N1527);
xor XOR2 (N1559, N1549, N1023);
nand NAND4 (N1560, N1556, N757, N1385, N1006);
not NOT1 (N1561, N1554);
nand NAND2 (N1562, N1536, N1282);
or OR2 (N1563, N1559, N419);
nor NOR2 (N1564, N1550, N347);
xor XOR2 (N1565, N1563, N1094);
or OR3 (N1566, N1553, N561, N927);
or OR2 (N1567, N1542, N1211);
nand NAND3 (N1568, N1564, N172, N712);
and AND3 (N1569, N1558, N602, N1211);
not NOT1 (N1570, N1565);
nor NOR4 (N1571, N1568, N808, N494, N276);
nor NOR3 (N1572, N1561, N1101, N76);
and AND4 (N1573, N1557, N457, N499, N182);
and AND3 (N1574, N1566, N750, N1158);
not NOT1 (N1575, N1560);
xor XOR2 (N1576, N1555, N791);
nor NOR4 (N1577, N1570, N1274, N1376, N1525);
and AND4 (N1578, N1562, N296, N1040, N1252);
nand NAND4 (N1579, N1573, N281, N1236, N1340);
nand NAND3 (N1580, N1577, N402, N650);
and AND2 (N1581, N1576, N206);
or OR4 (N1582, N1569, N395, N1271, N281);
and AND2 (N1583, N1581, N1574);
or OR2 (N1584, N657, N785);
xor XOR2 (N1585, N1571, N752);
or OR3 (N1586, N1582, N1080, N324);
and AND4 (N1587, N1583, N975, N1250, N907);
xor XOR2 (N1588, N1586, N491);
or OR4 (N1589, N1575, N1008, N598, N607);
and AND3 (N1590, N1572, N476, N861);
xor XOR2 (N1591, N1590, N727);
buf BUF1 (N1592, N1578);
nor NOR2 (N1593, N1579, N622);
buf BUF1 (N1594, N1589);
xor XOR2 (N1595, N1592, N1592);
or OR3 (N1596, N1594, N996, N382);
not NOT1 (N1597, N1584);
and AND3 (N1598, N1567, N1557, N418);
buf BUF1 (N1599, N1587);
or OR2 (N1600, N1588, N1265);
buf BUF1 (N1601, N1591);
and AND2 (N1602, N1601, N666);
buf BUF1 (N1603, N1593);
nor NOR2 (N1604, N1599, N1092);
nor NOR3 (N1605, N1598, N1516, N1382);
xor XOR2 (N1606, N1604, N1347);
and AND3 (N1607, N1596, N128, N424);
xor XOR2 (N1608, N1605, N1018);
and AND3 (N1609, N1608, N245, N82);
or OR4 (N1610, N1607, N62, N953, N1358);
nor NOR4 (N1611, N1595, N84, N253, N1133);
buf BUF1 (N1612, N1602);
not NOT1 (N1613, N1609);
nor NOR4 (N1614, N1603, N1068, N1286, N1003);
nor NOR4 (N1615, N1580, N1152, N1312, N1200);
nor NOR4 (N1616, N1606, N675, N316, N1505);
or OR4 (N1617, N1610, N57, N1189, N1333);
nand NAND2 (N1618, N1600, N630);
xor XOR2 (N1619, N1585, N708);
not NOT1 (N1620, N1614);
nor NOR2 (N1621, N1612, N305);
nand NAND3 (N1622, N1619, N1371, N334);
nor NOR4 (N1623, N1613, N137, N823, N3);
nand NAND2 (N1624, N1623, N234);
not NOT1 (N1625, N1618);
nor NOR4 (N1626, N1625, N351, N730, N272);
and AND2 (N1627, N1617, N134);
and AND2 (N1628, N1621, N1453);
or OR4 (N1629, N1597, N101, N682, N1151);
nor NOR2 (N1630, N1627, N47);
not NOT1 (N1631, N1629);
buf BUF1 (N1632, N1620);
not NOT1 (N1633, N1630);
nand NAND4 (N1634, N1631, N281, N728, N423);
and AND3 (N1635, N1633, N184, N74);
nand NAND3 (N1636, N1622, N1580, N815);
not NOT1 (N1637, N1634);
xor XOR2 (N1638, N1637, N179);
nand NAND4 (N1639, N1624, N714, N1455, N728);
or OR3 (N1640, N1615, N690, N1179);
xor XOR2 (N1641, N1628, N569);
or OR3 (N1642, N1611, N1494, N635);
buf BUF1 (N1643, N1639);
nor NOR3 (N1644, N1643, N966, N1189);
nand NAND3 (N1645, N1640, N101, N450);
or OR3 (N1646, N1635, N439, N387);
or OR4 (N1647, N1642, N467, N1552, N886);
xor XOR2 (N1648, N1647, N971);
and AND4 (N1649, N1648, N618, N58, N99);
nand NAND2 (N1650, N1649, N1066);
nor NOR2 (N1651, N1626, N110);
and AND2 (N1652, N1651, N618);
and AND3 (N1653, N1645, N1219, N155);
not NOT1 (N1654, N1638);
nor NOR4 (N1655, N1641, N493, N196, N1342);
and AND3 (N1656, N1616, N335, N117);
nand NAND4 (N1657, N1632, N452, N1649, N683);
and AND3 (N1658, N1653, N1180, N693);
xor XOR2 (N1659, N1658, N1223);
and AND3 (N1660, N1654, N615, N1101);
nor NOR4 (N1661, N1650, N204, N62, N586);
or OR4 (N1662, N1659, N730, N529, N1334);
buf BUF1 (N1663, N1644);
not NOT1 (N1664, N1656);
not NOT1 (N1665, N1657);
not NOT1 (N1666, N1660);
and AND3 (N1667, N1666, N191, N456);
buf BUF1 (N1668, N1646);
or OR3 (N1669, N1665, N90, N972);
or OR2 (N1670, N1652, N1152);
buf BUF1 (N1671, N1662);
or OR3 (N1672, N1655, N42, N532);
or OR3 (N1673, N1669, N1477, N91);
not NOT1 (N1674, N1664);
buf BUF1 (N1675, N1672);
buf BUF1 (N1676, N1636);
buf BUF1 (N1677, N1667);
buf BUF1 (N1678, N1675);
and AND4 (N1679, N1678, N275, N263, N1098);
and AND3 (N1680, N1677, N880, N556);
nand NAND2 (N1681, N1679, N614);
buf BUF1 (N1682, N1676);
xor XOR2 (N1683, N1670, N1116);
nand NAND3 (N1684, N1674, N1599, N328);
nor NOR2 (N1685, N1681, N82);
xor XOR2 (N1686, N1685, N1627);
and AND2 (N1687, N1671, N1253);
not NOT1 (N1688, N1682);
buf BUF1 (N1689, N1680);
nand NAND4 (N1690, N1686, N1287, N946, N939);
xor XOR2 (N1691, N1673, N1108);
and AND2 (N1692, N1687, N1104);
xor XOR2 (N1693, N1683, N1054);
buf BUF1 (N1694, N1693);
buf BUF1 (N1695, N1688);
buf BUF1 (N1696, N1692);
not NOT1 (N1697, N1689);
nor NOR2 (N1698, N1697, N47);
nor NOR2 (N1699, N1684, N21);
and AND2 (N1700, N1695, N1694);
or OR3 (N1701, N491, N1406, N1262);
not NOT1 (N1702, N1661);
nand NAND4 (N1703, N1701, N8, N329, N931);
and AND2 (N1704, N1663, N1216);
buf BUF1 (N1705, N1698);
or OR4 (N1706, N1705, N1338, N309, N1148);
buf BUF1 (N1707, N1703);
and AND3 (N1708, N1702, N42, N890);
nor NOR3 (N1709, N1699, N946, N1053);
or OR2 (N1710, N1691, N1582);
not NOT1 (N1711, N1700);
nand NAND3 (N1712, N1704, N54, N580);
buf BUF1 (N1713, N1712);
nor NOR2 (N1714, N1706, N1467);
buf BUF1 (N1715, N1714);
not NOT1 (N1716, N1710);
or OR3 (N1717, N1696, N1688, N1347);
nand NAND3 (N1718, N1668, N1562, N764);
xor XOR2 (N1719, N1713, N177);
buf BUF1 (N1720, N1719);
and AND3 (N1721, N1708, N1393, N1123);
xor XOR2 (N1722, N1716, N443);
xor XOR2 (N1723, N1721, N1381);
buf BUF1 (N1724, N1709);
or OR2 (N1725, N1720, N1539);
xor XOR2 (N1726, N1717, N564);
buf BUF1 (N1727, N1690);
xor XOR2 (N1728, N1718, N866);
not NOT1 (N1729, N1715);
xor XOR2 (N1730, N1722, N1190);
and AND3 (N1731, N1725, N725, N278);
xor XOR2 (N1732, N1723, N606);
and AND3 (N1733, N1711, N200, N172);
and AND3 (N1734, N1729, N110, N1697);
and AND3 (N1735, N1728, N491, N1414);
and AND4 (N1736, N1735, N192, N1360, N325);
and AND3 (N1737, N1707, N1671, N1691);
not NOT1 (N1738, N1724);
buf BUF1 (N1739, N1736);
not NOT1 (N1740, N1727);
buf BUF1 (N1741, N1740);
xor XOR2 (N1742, N1734, N1280);
not NOT1 (N1743, N1732);
xor XOR2 (N1744, N1726, N628);
buf BUF1 (N1745, N1737);
nor NOR2 (N1746, N1731, N904);
nor NOR2 (N1747, N1730, N297);
and AND4 (N1748, N1745, N1023, N1640, N920);
and AND3 (N1749, N1744, N1415, N1512);
nor NOR2 (N1750, N1748, N804);
buf BUF1 (N1751, N1750);
and AND4 (N1752, N1738, N1016, N1486, N152);
buf BUF1 (N1753, N1751);
and AND4 (N1754, N1753, N957, N205, N1746);
nand NAND4 (N1755, N1489, N1303, N250, N796);
nand NAND3 (N1756, N1747, N949, N1665);
nand NAND3 (N1757, N1749, N382, N372);
nand NAND2 (N1758, N1743, N311);
nand NAND2 (N1759, N1733, N491);
nor NOR3 (N1760, N1741, N424, N464);
buf BUF1 (N1761, N1757);
nand NAND4 (N1762, N1754, N1421, N979, N750);
nor NOR4 (N1763, N1759, N345, N748, N102);
not NOT1 (N1764, N1755);
not NOT1 (N1765, N1764);
nor NOR2 (N1766, N1752, N42);
xor XOR2 (N1767, N1739, N1010);
xor XOR2 (N1768, N1763, N1053);
xor XOR2 (N1769, N1768, N1651);
buf BUF1 (N1770, N1766);
nor NOR4 (N1771, N1761, N1574, N1130, N1066);
buf BUF1 (N1772, N1762);
or OR4 (N1773, N1769, N1607, N1135, N70);
nor NOR4 (N1774, N1742, N964, N1658, N335);
or OR4 (N1775, N1756, N1213, N1363, N311);
xor XOR2 (N1776, N1774, N741);
nor NOR2 (N1777, N1760, N951);
and AND3 (N1778, N1775, N257, N1581);
nand NAND4 (N1779, N1773, N1681, N406, N742);
and AND4 (N1780, N1777, N1602, N977, N605);
nor NOR3 (N1781, N1770, N393, N42);
nand NAND2 (N1782, N1767, N371);
and AND4 (N1783, N1779, N55, N1535, N1219);
nor NOR3 (N1784, N1782, N52, N838);
or OR4 (N1785, N1765, N1457, N1296, N584);
nor NOR3 (N1786, N1778, N212, N1315);
buf BUF1 (N1787, N1780);
not NOT1 (N1788, N1786);
or OR4 (N1789, N1771, N81, N1750, N1457);
not NOT1 (N1790, N1784);
or OR2 (N1791, N1772, N269);
or OR4 (N1792, N1758, N1589, N1598, N1148);
or OR2 (N1793, N1781, N1282);
buf BUF1 (N1794, N1789);
buf BUF1 (N1795, N1791);
not NOT1 (N1796, N1785);
not NOT1 (N1797, N1796);
not NOT1 (N1798, N1792);
and AND4 (N1799, N1797, N765, N191, N1591);
xor XOR2 (N1800, N1798, N453);
and AND2 (N1801, N1787, N117);
and AND2 (N1802, N1801, N304);
or OR2 (N1803, N1790, N282);
nand NAND3 (N1804, N1776, N1643, N134);
xor XOR2 (N1805, N1794, N1576);
nor NOR2 (N1806, N1795, N1566);
and AND4 (N1807, N1806, N837, N1196, N1145);
and AND2 (N1808, N1799, N1423);
or OR3 (N1809, N1788, N1546, N1572);
not NOT1 (N1810, N1804);
not NOT1 (N1811, N1807);
nor NOR4 (N1812, N1805, N715, N17, N1100);
and AND2 (N1813, N1808, N573);
or OR4 (N1814, N1800, N1464, N1810, N739);
or OR3 (N1815, N1633, N90, N819);
nand NAND3 (N1816, N1803, N1022, N609);
and AND2 (N1817, N1812, N1752);
or OR2 (N1818, N1809, N759);
nor NOR3 (N1819, N1783, N1288, N1720);
and AND2 (N1820, N1815, N977);
and AND2 (N1821, N1819, N1632);
not NOT1 (N1822, N1802);
nand NAND2 (N1823, N1818, N918);
nand NAND2 (N1824, N1793, N1022);
xor XOR2 (N1825, N1813, N869);
or OR3 (N1826, N1814, N1022, N195);
xor XOR2 (N1827, N1820, N525);
xor XOR2 (N1828, N1817, N528);
and AND3 (N1829, N1816, N1212, N938);
nor NOR4 (N1830, N1811, N591, N139, N81);
nor NOR2 (N1831, N1826, N220);
and AND4 (N1832, N1827, N855, N200, N998);
or OR3 (N1833, N1831, N1443, N1646);
and AND2 (N1834, N1824, N365);
or OR2 (N1835, N1822, N1386);
nor NOR3 (N1836, N1829, N931, N631);
buf BUF1 (N1837, N1828);
not NOT1 (N1838, N1836);
or OR3 (N1839, N1838, N369, N348);
xor XOR2 (N1840, N1835, N1070);
or OR3 (N1841, N1834, N1289, N1254);
xor XOR2 (N1842, N1830, N962);
xor XOR2 (N1843, N1839, N1367);
xor XOR2 (N1844, N1825, N1042);
nand NAND3 (N1845, N1823, N1411, N1435);
nor NOR4 (N1846, N1843, N772, N871, N696);
buf BUF1 (N1847, N1845);
buf BUF1 (N1848, N1840);
not NOT1 (N1849, N1847);
buf BUF1 (N1850, N1832);
nand NAND4 (N1851, N1842, N495, N1659, N654);
nand NAND4 (N1852, N1833, N1556, N761, N200);
buf BUF1 (N1853, N1852);
buf BUF1 (N1854, N1846);
or OR4 (N1855, N1844, N1769, N700, N43);
buf BUF1 (N1856, N1848);
or OR4 (N1857, N1853, N486, N1090, N970);
or OR4 (N1858, N1855, N1114, N477, N516);
or OR4 (N1859, N1837, N594, N376, N1149);
buf BUF1 (N1860, N1859);
not NOT1 (N1861, N1841);
xor XOR2 (N1862, N1849, N758);
xor XOR2 (N1863, N1850, N1274);
and AND2 (N1864, N1851, N1624);
nor NOR2 (N1865, N1857, N1210);
nor NOR2 (N1866, N1864, N753);
and AND4 (N1867, N1866, N1763, N616, N1695);
or OR2 (N1868, N1854, N539);
nor NOR2 (N1869, N1856, N1138);
or OR2 (N1870, N1863, N482);
or OR2 (N1871, N1861, N1699);
or OR2 (N1872, N1868, N609);
or OR2 (N1873, N1862, N875);
buf BUF1 (N1874, N1870);
and AND2 (N1875, N1869, N1602);
and AND3 (N1876, N1875, N1862, N657);
and AND3 (N1877, N1876, N1201, N1337);
and AND4 (N1878, N1867, N627, N693, N1768);
buf BUF1 (N1879, N1858);
or OR3 (N1880, N1871, N1441, N632);
and AND2 (N1881, N1874, N493);
nand NAND3 (N1882, N1877, N1646, N1770);
buf BUF1 (N1883, N1879);
not NOT1 (N1884, N1882);
nor NOR4 (N1885, N1873, N1593, N700, N693);
and AND3 (N1886, N1885, N437, N493);
or OR3 (N1887, N1884, N1540, N318);
buf BUF1 (N1888, N1878);
nor NOR4 (N1889, N1880, N1313, N1512, N749);
nor NOR4 (N1890, N1888, N1396, N256, N1032);
not NOT1 (N1891, N1889);
nand NAND3 (N1892, N1886, N846, N1447);
xor XOR2 (N1893, N1821, N416);
and AND2 (N1894, N1891, N955);
buf BUF1 (N1895, N1890);
buf BUF1 (N1896, N1892);
xor XOR2 (N1897, N1860, N1669);
not NOT1 (N1898, N1895);
or OR2 (N1899, N1893, N866);
and AND2 (N1900, N1887, N1173);
not NOT1 (N1901, N1897);
nor NOR2 (N1902, N1894, N1761);
or OR3 (N1903, N1898, N1104, N182);
xor XOR2 (N1904, N1883, N1331);
and AND3 (N1905, N1865, N199, N1341);
or OR2 (N1906, N1901, N1370);
xor XOR2 (N1907, N1900, N1340);
and AND2 (N1908, N1903, N1879);
nor NOR2 (N1909, N1896, N903);
nor NOR4 (N1910, N1902, N567, N1184, N417);
or OR2 (N1911, N1906, N292);
xor XOR2 (N1912, N1872, N61);
or OR3 (N1913, N1909, N1159, N1183);
nor NOR2 (N1914, N1881, N1900);
nor NOR2 (N1915, N1908, N116);
and AND3 (N1916, N1915, N1068, N481);
xor XOR2 (N1917, N1916, N527);
not NOT1 (N1918, N1917);
buf BUF1 (N1919, N1911);
nand NAND3 (N1920, N1899, N347, N770);
xor XOR2 (N1921, N1918, N1623);
buf BUF1 (N1922, N1905);
nor NOR2 (N1923, N1920, N1449);
or OR4 (N1924, N1921, N1233, N419, N125);
xor XOR2 (N1925, N1923, N1736);
and AND2 (N1926, N1922, N567);
and AND3 (N1927, N1914, N948, N1341);
and AND3 (N1928, N1924, N721, N1893);
buf BUF1 (N1929, N1913);
not NOT1 (N1930, N1927);
or OR3 (N1931, N1919, N1356, N931);
or OR2 (N1932, N1912, N1833);
buf BUF1 (N1933, N1904);
and AND2 (N1934, N1910, N886);
or OR2 (N1935, N1934, N249);
nand NAND4 (N1936, N1907, N1562, N1210, N1087);
not NOT1 (N1937, N1936);
xor XOR2 (N1938, N1926, N976);
not NOT1 (N1939, N1935);
buf BUF1 (N1940, N1931);
xor XOR2 (N1941, N1925, N313);
and AND4 (N1942, N1929, N1683, N1657, N1444);
or OR2 (N1943, N1933, N1686);
or OR4 (N1944, N1939, N234, N1073, N359);
xor XOR2 (N1945, N1941, N1177);
or OR2 (N1946, N1932, N1921);
xor XOR2 (N1947, N1944, N534);
buf BUF1 (N1948, N1937);
xor XOR2 (N1949, N1938, N547);
or OR2 (N1950, N1949, N171);
buf BUF1 (N1951, N1943);
or OR2 (N1952, N1951, N1553);
nor NOR2 (N1953, N1950, N1905);
buf BUF1 (N1954, N1946);
and AND4 (N1955, N1930, N1627, N1643, N794);
buf BUF1 (N1956, N1928);
nor NOR4 (N1957, N1948, N1189, N10, N685);
nand NAND2 (N1958, N1957, N286);
not NOT1 (N1959, N1956);
and AND2 (N1960, N1954, N610);
and AND3 (N1961, N1955, N469, N869);
not NOT1 (N1962, N1959);
and AND4 (N1963, N1945, N1356, N1188, N195);
nand NAND2 (N1964, N1942, N1117);
buf BUF1 (N1965, N1958);
and AND2 (N1966, N1963, N1580);
or OR4 (N1967, N1964, N1806, N1651, N1622);
nand NAND2 (N1968, N1965, N1953);
buf BUF1 (N1969, N918);
and AND2 (N1970, N1961, N1820);
xor XOR2 (N1971, N1947, N1677);
and AND4 (N1972, N1952, N686, N1794, N1326);
nor NOR3 (N1973, N1970, N1133, N1384);
not NOT1 (N1974, N1972);
xor XOR2 (N1975, N1962, N1467);
not NOT1 (N1976, N1974);
nand NAND2 (N1977, N1960, N757);
and AND3 (N1978, N1940, N778, N217);
buf BUF1 (N1979, N1969);
nand NAND4 (N1980, N1966, N1028, N1185, N1541);
buf BUF1 (N1981, N1980);
and AND2 (N1982, N1973, N287);
nand NAND3 (N1983, N1976, N711, N1192);
or OR2 (N1984, N1982, N557);
or OR3 (N1985, N1967, N1977, N457);
nand NAND3 (N1986, N744, N151, N1395);
not NOT1 (N1987, N1978);
xor XOR2 (N1988, N1986, N1215);
or OR3 (N1989, N1984, N514, N282);
nand NAND3 (N1990, N1971, N1489, N801);
xor XOR2 (N1991, N1988, N1120);
buf BUF1 (N1992, N1990);
nand NAND3 (N1993, N1983, N1900, N150);
not NOT1 (N1994, N1981);
nor NOR3 (N1995, N1975, N101, N545);
buf BUF1 (N1996, N1993);
or OR4 (N1997, N1987, N1226, N969, N1048);
buf BUF1 (N1998, N1997);
nand NAND3 (N1999, N1992, N1484, N745);
xor XOR2 (N2000, N1996, N1099);
nand NAND4 (N2001, N1979, N1920, N1774, N644);
buf BUF1 (N2002, N1985);
buf BUF1 (N2003, N1995);
or OR4 (N2004, N2000, N1386, N259, N1267);
and AND3 (N2005, N1968, N1995, N710);
nand NAND2 (N2006, N2002, N1967);
nor NOR3 (N2007, N1999, N610, N309);
xor XOR2 (N2008, N2001, N1943);
or OR2 (N2009, N1998, N464);
nand NAND4 (N2010, N2004, N1722, N725, N255);
or OR3 (N2011, N1989, N1926, N1561);
and AND3 (N2012, N2005, N647, N304);
and AND4 (N2013, N2011, N506, N1965, N1822);
nor NOR3 (N2014, N1994, N116, N1044);
xor XOR2 (N2015, N2013, N1047);
or OR3 (N2016, N2007, N1287, N1893);
nand NAND2 (N2017, N2012, N1196);
and AND2 (N2018, N2015, N1934);
or OR4 (N2019, N2006, N603, N1198, N906);
xor XOR2 (N2020, N2016, N1710);
and AND3 (N2021, N2014, N419, N258);
not NOT1 (N2022, N2009);
nor NOR3 (N2023, N2008, N811, N380);
nand NAND3 (N2024, N2021, N1120, N1320);
buf BUF1 (N2025, N2017);
buf BUF1 (N2026, N2020);
not NOT1 (N2027, N2023);
not NOT1 (N2028, N1991);
buf BUF1 (N2029, N2028);
nor NOR4 (N2030, N2019, N1862, N1459, N1559);
nor NOR2 (N2031, N2029, N1135);
or OR3 (N2032, N2026, N1162, N515);
buf BUF1 (N2033, N2027);
not NOT1 (N2034, N2003);
xor XOR2 (N2035, N2018, N1380);
nand NAND4 (N2036, N2024, N935, N20, N717);
not NOT1 (N2037, N2036);
or OR2 (N2038, N2034, N1702);
xor XOR2 (N2039, N2037, N850);
nand NAND2 (N2040, N2022, N647);
nor NOR4 (N2041, N2030, N706, N2006, N1144);
or OR2 (N2042, N2031, N692);
or OR4 (N2043, N2039, N163, N1215, N427);
xor XOR2 (N2044, N2025, N813);
and AND2 (N2045, N2010, N1441);
and AND3 (N2046, N2042, N420, N340);
not NOT1 (N2047, N2046);
not NOT1 (N2048, N2045);
and AND3 (N2049, N2041, N1139, N1851);
buf BUF1 (N2050, N2038);
xor XOR2 (N2051, N2043, N1543);
and AND2 (N2052, N2047, N802);
or OR2 (N2053, N2032, N896);
and AND4 (N2054, N2050, N49, N358, N758);
and AND3 (N2055, N2049, N1825, N541);
buf BUF1 (N2056, N2048);
buf BUF1 (N2057, N2033);
nor NOR4 (N2058, N2054, N804, N26, N529);
nor NOR3 (N2059, N2052, N786, N805);
or OR3 (N2060, N2035, N985, N1030);
xor XOR2 (N2061, N2040, N1685);
nor NOR2 (N2062, N2058, N1367);
and AND2 (N2063, N2044, N369);
or OR3 (N2064, N2061, N822, N902);
nor NOR4 (N2065, N2053, N625, N1719, N1910);
xor XOR2 (N2066, N2059, N297);
xor XOR2 (N2067, N2057, N1990);
buf BUF1 (N2068, N2051);
and AND3 (N2069, N2055, N373, N287);
not NOT1 (N2070, N2062);
xor XOR2 (N2071, N2060, N203);
nor NOR2 (N2072, N2065, N743);
buf BUF1 (N2073, N2067);
and AND2 (N2074, N2071, N2037);
nand NAND3 (N2075, N2073, N1407, N1685);
and AND2 (N2076, N2072, N222);
nand NAND4 (N2077, N2074, N1640, N928, N1123);
and AND3 (N2078, N2066, N914, N156);
xor XOR2 (N2079, N2063, N110);
nand NAND4 (N2080, N2075, N514, N1921, N921);
buf BUF1 (N2081, N2069);
buf BUF1 (N2082, N2070);
nor NOR2 (N2083, N2068, N656);
or OR2 (N2084, N2056, N414);
xor XOR2 (N2085, N2082, N1650);
xor XOR2 (N2086, N2084, N1306);
buf BUF1 (N2087, N2085);
xor XOR2 (N2088, N2064, N2004);
xor XOR2 (N2089, N2081, N1952);
or OR3 (N2090, N2079, N276, N2085);
xor XOR2 (N2091, N2083, N1519);
not NOT1 (N2092, N2090);
nor NOR4 (N2093, N2080, N830, N1788, N294);
nor NOR3 (N2094, N2092, N1355, N489);
or OR4 (N2095, N2089, N428, N533, N234);
nand NAND2 (N2096, N2076, N2041);
not NOT1 (N2097, N2087);
not NOT1 (N2098, N2078);
not NOT1 (N2099, N2088);
xor XOR2 (N2100, N2077, N570);
buf BUF1 (N2101, N2091);
or OR3 (N2102, N2093, N1280, N717);
buf BUF1 (N2103, N2100);
or OR3 (N2104, N2094, N149, N129);
nand NAND4 (N2105, N2098, N1353, N44, N1807);
xor XOR2 (N2106, N2086, N635);
nand NAND4 (N2107, N2097, N1921, N1126, N91);
nand NAND3 (N2108, N2104, N406, N1231);
nor NOR4 (N2109, N2102, N1261, N687, N1250);
and AND2 (N2110, N2103, N1441);
or OR3 (N2111, N2107, N1668, N2070);
and AND2 (N2112, N2108, N1443);
or OR2 (N2113, N2105, N1305);
and AND3 (N2114, N2111, N1745, N1790);
nand NAND3 (N2115, N2109, N888, N1436);
nand NAND4 (N2116, N2114, N1338, N606, N790);
buf BUF1 (N2117, N2106);
xor XOR2 (N2118, N2112, N1390);
not NOT1 (N2119, N2115);
nand NAND4 (N2120, N2099, N1622, N493, N40);
nand NAND4 (N2121, N2117, N849, N768, N1135);
nand NAND4 (N2122, N2121, N1158, N471, N1158);
xor XOR2 (N2123, N2116, N683);
nor NOR3 (N2124, N2095, N1110, N169);
not NOT1 (N2125, N2119);
nor NOR3 (N2126, N2123, N409, N1416);
buf BUF1 (N2127, N2122);
or OR3 (N2128, N2124, N2112, N1197);
buf BUF1 (N2129, N2127);
nor NOR4 (N2130, N2125, N1482, N1199, N1950);
or OR4 (N2131, N2110, N1747, N2032, N545);
buf BUF1 (N2132, N2131);
nor NOR3 (N2133, N2113, N1385, N138);
and AND2 (N2134, N2126, N1872);
buf BUF1 (N2135, N2101);
buf BUF1 (N2136, N2120);
and AND4 (N2137, N2136, N1020, N928, N1909);
xor XOR2 (N2138, N2132, N861);
not NOT1 (N2139, N2135);
buf BUF1 (N2140, N2096);
nand NAND4 (N2141, N2134, N293, N1602, N2053);
nand NAND3 (N2142, N2139, N76, N1293);
and AND2 (N2143, N2138, N703);
xor XOR2 (N2144, N2142, N1503);
or OR2 (N2145, N2129, N1870);
and AND3 (N2146, N2140, N1147, N373);
not NOT1 (N2147, N2128);
nor NOR3 (N2148, N2118, N267, N987);
xor XOR2 (N2149, N2143, N1322);
nor NOR4 (N2150, N2141, N610, N994, N1651);
xor XOR2 (N2151, N2144, N1851);
nor NOR4 (N2152, N2150, N811, N1728, N568);
xor XOR2 (N2153, N2130, N1956);
nor NOR3 (N2154, N2147, N35, N1853);
nand NAND2 (N2155, N2137, N281);
or OR3 (N2156, N2146, N1351, N232);
xor XOR2 (N2157, N2154, N601);
or OR4 (N2158, N2133, N583, N844, N880);
and AND3 (N2159, N2157, N1843, N1532);
or OR3 (N2160, N2159, N1860, N260);
and AND2 (N2161, N2148, N31);
nor NOR3 (N2162, N2156, N1752, N432);
nand NAND3 (N2163, N2161, N1413, N1875);
nor NOR4 (N2164, N2151, N1458, N608, N1638);
xor XOR2 (N2165, N2145, N1788);
nand NAND4 (N2166, N2164, N1945, N1439, N456);
not NOT1 (N2167, N2153);
buf BUF1 (N2168, N2152);
and AND2 (N2169, N2162, N438);
nor NOR2 (N2170, N2160, N1606);
not NOT1 (N2171, N2149);
buf BUF1 (N2172, N2167);
xor XOR2 (N2173, N2171, N2028);
not NOT1 (N2174, N2169);
xor XOR2 (N2175, N2158, N1960);
buf BUF1 (N2176, N2168);
buf BUF1 (N2177, N2163);
buf BUF1 (N2178, N2177);
nand NAND2 (N2179, N2166, N1984);
nor NOR2 (N2180, N2165, N1383);
or OR3 (N2181, N2174, N1229, N1262);
xor XOR2 (N2182, N2172, N1062);
buf BUF1 (N2183, N2180);
xor XOR2 (N2184, N2176, N780);
and AND3 (N2185, N2175, N1676, N1529);
and AND4 (N2186, N2170, N1570, N1257, N413);
and AND2 (N2187, N2181, N1856);
xor XOR2 (N2188, N2184, N340);
xor XOR2 (N2189, N2182, N1086);
nor NOR2 (N2190, N2178, N1473);
and AND2 (N2191, N2183, N781);
nor NOR2 (N2192, N2189, N1205);
nor NOR4 (N2193, N2190, N1277, N341, N1767);
or OR4 (N2194, N2155, N1561, N158, N1154);
or OR2 (N2195, N2193, N1514);
nand NAND3 (N2196, N2187, N795, N441);
buf BUF1 (N2197, N2188);
not NOT1 (N2198, N2173);
buf BUF1 (N2199, N2185);
buf BUF1 (N2200, N2192);
or OR3 (N2201, N2194, N882, N123);
or OR4 (N2202, N2199, N923, N876, N1730);
buf BUF1 (N2203, N2186);
and AND4 (N2204, N2197, N826, N652, N1241);
and AND2 (N2205, N2179, N61);
nor NOR3 (N2206, N2203, N586, N1878);
and AND2 (N2207, N2205, N1003);
not NOT1 (N2208, N2196);
or OR3 (N2209, N2204, N771, N1866);
buf BUF1 (N2210, N2202);
nor NOR3 (N2211, N2207, N1945, N1673);
xor XOR2 (N2212, N2200, N1635);
buf BUF1 (N2213, N2210);
buf BUF1 (N2214, N2201);
or OR2 (N2215, N2213, N1123);
nor NOR4 (N2216, N2208, N308, N1888, N2087);
buf BUF1 (N2217, N2215);
nand NAND4 (N2218, N2212, N1870, N1078, N626);
or OR4 (N2219, N2211, N1143, N1787, N609);
or OR2 (N2220, N2217, N374);
or OR2 (N2221, N2206, N673);
nand NAND2 (N2222, N2220, N422);
or OR2 (N2223, N2222, N446);
buf BUF1 (N2224, N2191);
and AND4 (N2225, N2198, N1286, N1411, N1453);
buf BUF1 (N2226, N2214);
and AND4 (N2227, N2219, N2043, N172, N995);
not NOT1 (N2228, N2218);
xor XOR2 (N2229, N2228, N466);
not NOT1 (N2230, N2229);
not NOT1 (N2231, N2224);
not NOT1 (N2232, N2226);
nor NOR2 (N2233, N2225, N641);
not NOT1 (N2234, N2232);
nor NOR3 (N2235, N2234, N2045, N666);
nor NOR2 (N2236, N2231, N1576);
and AND3 (N2237, N2195, N657, N1709);
nor NOR2 (N2238, N2221, N227);
or OR3 (N2239, N2209, N357, N256);
and AND4 (N2240, N2230, N691, N14, N1666);
and AND4 (N2241, N2236, N1153, N1813, N1143);
nand NAND3 (N2242, N2241, N927, N1922);
nand NAND2 (N2243, N2223, N1439);
nor NOR2 (N2244, N2239, N733);
nand NAND4 (N2245, N2243, N1809, N1316, N693);
not NOT1 (N2246, N2242);
xor XOR2 (N2247, N2216, N2002);
not NOT1 (N2248, N2233);
buf BUF1 (N2249, N2235);
nor NOR2 (N2250, N2247, N1959);
or OR2 (N2251, N2238, N601);
and AND2 (N2252, N2240, N998);
and AND2 (N2253, N2252, N2141);
nor NOR4 (N2254, N2248, N1452, N275, N1396);
xor XOR2 (N2255, N2237, N550);
nor NOR3 (N2256, N2245, N13, N105);
not NOT1 (N2257, N2246);
xor XOR2 (N2258, N2250, N977);
and AND3 (N2259, N2249, N365, N1592);
nor NOR2 (N2260, N2244, N1712);
xor XOR2 (N2261, N2257, N1625);
xor XOR2 (N2262, N2256, N29);
or OR4 (N2263, N2258, N873, N1186, N1153);
or OR2 (N2264, N2261, N234);
buf BUF1 (N2265, N2264);
buf BUF1 (N2266, N2265);
and AND2 (N2267, N2255, N234);
not NOT1 (N2268, N2267);
or OR4 (N2269, N2227, N1971, N428, N1915);
xor XOR2 (N2270, N2269, N1152);
or OR3 (N2271, N2251, N565, N1087);
nand NAND2 (N2272, N2254, N1985);
or OR3 (N2273, N2260, N2160, N1621);
nor NOR3 (N2274, N2271, N956, N1886);
xor XOR2 (N2275, N2266, N466);
not NOT1 (N2276, N2253);
or OR3 (N2277, N2274, N887, N1863);
xor XOR2 (N2278, N2263, N1555);
nor NOR3 (N2279, N2259, N365, N363);
buf BUF1 (N2280, N2270);
and AND2 (N2281, N2262, N983);
nand NAND2 (N2282, N2273, N1112);
xor XOR2 (N2283, N2277, N1810);
buf BUF1 (N2284, N2283);
nor NOR3 (N2285, N2284, N611, N1084);
nor NOR3 (N2286, N2282, N1567, N1899);
not NOT1 (N2287, N2275);
or OR2 (N2288, N2286, N1377);
buf BUF1 (N2289, N2288);
and AND3 (N2290, N2279, N11, N616);
not NOT1 (N2291, N2285);
or OR3 (N2292, N2272, N1903, N2276);
xor XOR2 (N2293, N1126, N440);
not NOT1 (N2294, N2280);
xor XOR2 (N2295, N2278, N793);
xor XOR2 (N2296, N2291, N1920);
nand NAND2 (N2297, N2293, N967);
not NOT1 (N2298, N2268);
xor XOR2 (N2299, N2294, N169);
nand NAND3 (N2300, N2289, N1039, N303);
nor NOR2 (N2301, N2298, N2093);
nor NOR3 (N2302, N2281, N1885, N1451);
nand NAND4 (N2303, N2302, N456, N891, N2103);
nor NOR2 (N2304, N2299, N496);
or OR3 (N2305, N2290, N2178, N1598);
xor XOR2 (N2306, N2292, N1907);
or OR2 (N2307, N2297, N2236);
and AND4 (N2308, N2295, N1709, N2044, N1227);
buf BUF1 (N2309, N2287);
not NOT1 (N2310, N2307);
nand NAND2 (N2311, N2309, N2242);
buf BUF1 (N2312, N2308);
xor XOR2 (N2313, N2300, N1966);
or OR4 (N2314, N2305, N1570, N2255, N1704);
buf BUF1 (N2315, N2311);
buf BUF1 (N2316, N2301);
and AND3 (N2317, N2310, N154, N75);
not NOT1 (N2318, N2315);
or OR3 (N2319, N2313, N83, N1976);
nor NOR3 (N2320, N2314, N1003, N1386);
xor XOR2 (N2321, N2316, N1711);
nand NAND3 (N2322, N2303, N680, N1874);
buf BUF1 (N2323, N2322);
nor NOR4 (N2324, N2304, N334, N1156, N1779);
or OR3 (N2325, N2324, N291, N98);
not NOT1 (N2326, N2321);
not NOT1 (N2327, N2317);
nand NAND4 (N2328, N2312, N242, N1167, N658);
not NOT1 (N2329, N2326);
not NOT1 (N2330, N2306);
not NOT1 (N2331, N2325);
not NOT1 (N2332, N2327);
xor XOR2 (N2333, N2296, N408);
and AND4 (N2334, N2332, N521, N1901, N1108);
nand NAND4 (N2335, N2334, N462, N436, N1368);
not NOT1 (N2336, N2329);
buf BUF1 (N2337, N2328);
xor XOR2 (N2338, N2318, N803);
buf BUF1 (N2339, N2333);
xor XOR2 (N2340, N2330, N1796);
nor NOR4 (N2341, N2338, N720, N1367, N1713);
xor XOR2 (N2342, N2336, N1541);
and AND3 (N2343, N2339, N204, N849);
nor NOR2 (N2344, N2320, N714);
xor XOR2 (N2345, N2337, N1917);
or OR4 (N2346, N2343, N766, N2298, N1850);
buf BUF1 (N2347, N2319);
xor XOR2 (N2348, N2335, N536);
not NOT1 (N2349, N2347);
xor XOR2 (N2350, N2345, N2318);
not NOT1 (N2351, N2341);
buf BUF1 (N2352, N2331);
xor XOR2 (N2353, N2344, N1298);
xor XOR2 (N2354, N2353, N453);
not NOT1 (N2355, N2354);
or OR3 (N2356, N2342, N1154, N431);
buf BUF1 (N2357, N2351);
buf BUF1 (N2358, N2357);
or OR3 (N2359, N2340, N1923, N1230);
or OR4 (N2360, N2352, N1821, N2026, N1901);
nor NOR3 (N2361, N2348, N633, N904);
buf BUF1 (N2362, N2323);
nand NAND3 (N2363, N2358, N802, N1488);
and AND2 (N2364, N2355, N418);
nor NOR4 (N2365, N2349, N993, N1999, N1663);
buf BUF1 (N2366, N2359);
and AND2 (N2367, N2365, N782);
buf BUF1 (N2368, N2346);
or OR4 (N2369, N2368, N1337, N1973, N232);
buf BUF1 (N2370, N2350);
and AND2 (N2371, N2366, N1335);
or OR4 (N2372, N2363, N208, N1419, N688);
xor XOR2 (N2373, N2362, N2114);
xor XOR2 (N2374, N2356, N1114);
and AND4 (N2375, N2364, N1019, N847, N883);
or OR2 (N2376, N2374, N1826);
or OR2 (N2377, N2369, N81);
nand NAND2 (N2378, N2370, N596);
nor NOR3 (N2379, N2378, N1112, N1262);
not NOT1 (N2380, N2367);
xor XOR2 (N2381, N2360, N1848);
xor XOR2 (N2382, N2377, N249);
buf BUF1 (N2383, N2371);
nor NOR3 (N2384, N2372, N1159, N285);
and AND3 (N2385, N2380, N1658, N1315);
and AND4 (N2386, N2384, N1819, N999, N1067);
not NOT1 (N2387, N2375);
and AND3 (N2388, N2385, N792, N1518);
nor NOR3 (N2389, N2382, N2027, N734);
and AND4 (N2390, N2389, N2208, N2113, N870);
nand NAND4 (N2391, N2390, N895, N10, N294);
nor NOR4 (N2392, N2373, N990, N2208, N1803);
xor XOR2 (N2393, N2387, N2134);
and AND2 (N2394, N2386, N1695);
and AND4 (N2395, N2379, N880, N517, N812);
xor XOR2 (N2396, N2381, N833);
or OR3 (N2397, N2393, N283, N644);
nor NOR3 (N2398, N2392, N2023, N892);
nand NAND3 (N2399, N2361, N1916, N517);
xor XOR2 (N2400, N2391, N2172);
nand NAND3 (N2401, N2398, N2331, N2389);
buf BUF1 (N2402, N2397);
not NOT1 (N2403, N2376);
nand NAND2 (N2404, N2395, N1220);
buf BUF1 (N2405, N2394);
or OR2 (N2406, N2396, N2108);
or OR4 (N2407, N2400, N532, N1720, N567);
not NOT1 (N2408, N2405);
buf BUF1 (N2409, N2399);
not NOT1 (N2410, N2408);
nand NAND3 (N2411, N2409, N907, N2154);
and AND2 (N2412, N2406, N1781);
nand NAND4 (N2413, N2407, N1459, N497, N1660);
nand NAND3 (N2414, N2404, N709, N2198);
not NOT1 (N2415, N2410);
nand NAND4 (N2416, N2413, N1906, N1143, N1882);
nor NOR3 (N2417, N2383, N572, N1017);
nand NAND2 (N2418, N2415, N245);
buf BUF1 (N2419, N2418);
buf BUF1 (N2420, N2388);
or OR4 (N2421, N2414, N81, N1661, N59);
buf BUF1 (N2422, N2419);
or OR2 (N2423, N2402, N1117);
not NOT1 (N2424, N2417);
not NOT1 (N2425, N2403);
and AND3 (N2426, N2401, N631, N1968);
not NOT1 (N2427, N2420);
nand NAND2 (N2428, N2421, N868);
not NOT1 (N2429, N2427);
not NOT1 (N2430, N2411);
and AND4 (N2431, N2429, N1102, N1455, N585);
or OR4 (N2432, N2430, N1718, N772, N812);
and AND4 (N2433, N2423, N718, N1902, N974);
or OR3 (N2434, N2432, N55, N1501);
or OR3 (N2435, N2416, N873, N124);
xor XOR2 (N2436, N2424, N1879);
or OR3 (N2437, N2428, N2362, N2300);
not NOT1 (N2438, N2422);
or OR2 (N2439, N2435, N1136);
buf BUF1 (N2440, N2412);
or OR2 (N2441, N2433, N2327);
not NOT1 (N2442, N2434);
and AND3 (N2443, N2431, N841, N463);
nor NOR3 (N2444, N2441, N2273, N1126);
nor NOR2 (N2445, N2439, N1115);
nand NAND4 (N2446, N2445, N2193, N578, N305);
nor NOR4 (N2447, N2446, N306, N513, N1389);
buf BUF1 (N2448, N2436);
or OR2 (N2449, N2447, N1158);
buf BUF1 (N2450, N2426);
nor NOR2 (N2451, N2440, N1350);
not NOT1 (N2452, N2450);
not NOT1 (N2453, N2425);
buf BUF1 (N2454, N2448);
buf BUF1 (N2455, N2453);
and AND4 (N2456, N2443, N1189, N1723, N1368);
not NOT1 (N2457, N2452);
and AND4 (N2458, N2438, N842, N924, N1495);
or OR2 (N2459, N2451, N701);
xor XOR2 (N2460, N2454, N267);
xor XOR2 (N2461, N2455, N1922);
not NOT1 (N2462, N2444);
nor NOR3 (N2463, N2459, N1542, N1220);
nand NAND3 (N2464, N2462, N673, N1701);
nand NAND4 (N2465, N2457, N1137, N1670, N540);
and AND2 (N2466, N2442, N141);
or OR4 (N2467, N2463, N1753, N81, N1243);
not NOT1 (N2468, N2466);
xor XOR2 (N2469, N2465, N2081);
not NOT1 (N2470, N2469);
nor NOR4 (N2471, N2467, N2139, N706, N1551);
not NOT1 (N2472, N2458);
nor NOR3 (N2473, N2468, N1987, N1450);
or OR2 (N2474, N2456, N1701);
xor XOR2 (N2475, N2471, N787);
or OR3 (N2476, N2475, N621, N1666);
nor NOR3 (N2477, N2449, N1011, N1821);
xor XOR2 (N2478, N2474, N1756);
buf BUF1 (N2479, N2473);
nand NAND2 (N2480, N2472, N1567);
and AND3 (N2481, N2478, N232, N1156);
nor NOR2 (N2482, N2437, N1029);
buf BUF1 (N2483, N2477);
buf BUF1 (N2484, N2470);
xor XOR2 (N2485, N2464, N1841);
and AND4 (N2486, N2479, N1274, N534, N1641);
or OR4 (N2487, N2461, N1411, N1713, N2038);
or OR3 (N2488, N2480, N909, N1507);
not NOT1 (N2489, N2486);
or OR3 (N2490, N2487, N1165, N365);
buf BUF1 (N2491, N2482);
or OR3 (N2492, N2483, N2200, N1664);
nor NOR2 (N2493, N2476, N2341);
nor NOR2 (N2494, N2460, N1526);
and AND3 (N2495, N2484, N1973, N488);
nand NAND3 (N2496, N2492, N272, N1074);
nor NOR2 (N2497, N2488, N57);
nand NAND4 (N2498, N2489, N1873, N1907, N1590);
buf BUF1 (N2499, N2497);
nor NOR2 (N2500, N2495, N2055);
nor NOR4 (N2501, N2490, N2317, N1769, N1179);
nand NAND2 (N2502, N2499, N596);
or OR2 (N2503, N2501, N1716);
xor XOR2 (N2504, N2494, N1476);
or OR2 (N2505, N2485, N863);
or OR2 (N2506, N2493, N955);
nand NAND3 (N2507, N2505, N706, N1783);
and AND4 (N2508, N2507, N1750, N2006, N2475);
nand NAND2 (N2509, N2481, N1483);
buf BUF1 (N2510, N2502);
nor NOR2 (N2511, N2498, N2127);
nor NOR3 (N2512, N2506, N484, N1479);
xor XOR2 (N2513, N2496, N1564);
and AND3 (N2514, N2510, N1037, N2281);
xor XOR2 (N2515, N2509, N849);
xor XOR2 (N2516, N2503, N694);
and AND4 (N2517, N2491, N1829, N1802, N2398);
nand NAND4 (N2518, N2517, N673, N535, N1125);
xor XOR2 (N2519, N2512, N1926);
buf BUF1 (N2520, N2518);
nand NAND3 (N2521, N2513, N1438, N1541);
and AND4 (N2522, N2519, N264, N2088, N2155);
nor NOR3 (N2523, N2522, N1861, N53);
or OR3 (N2524, N2500, N2011, N2069);
nor NOR4 (N2525, N2524, N346, N932, N2034);
xor XOR2 (N2526, N2525, N653);
xor XOR2 (N2527, N2514, N1554);
xor XOR2 (N2528, N2526, N776);
nand NAND3 (N2529, N2523, N1177, N56);
nor NOR2 (N2530, N2515, N491);
buf BUF1 (N2531, N2527);
and AND2 (N2532, N2520, N2194);
nor NOR4 (N2533, N2516, N1990, N1285, N524);
nand NAND4 (N2534, N2521, N1230, N236, N1540);
and AND3 (N2535, N2534, N1949, N2268);
not NOT1 (N2536, N2533);
or OR3 (N2537, N2528, N175, N158);
and AND2 (N2538, N2536, N731);
or OR4 (N2539, N2504, N73, N55, N2512);
not NOT1 (N2540, N2539);
and AND3 (N2541, N2538, N264, N725);
and AND3 (N2542, N2537, N464, N671);
and AND3 (N2543, N2542, N362, N441);
buf BUF1 (N2544, N2540);
nand NAND3 (N2545, N2531, N396, N1243);
or OR4 (N2546, N2535, N444, N1921, N1658);
nand NAND3 (N2547, N2508, N465, N1514);
or OR4 (N2548, N2541, N1635, N470, N633);
nor NOR4 (N2549, N2545, N1588, N2154, N1302);
and AND4 (N2550, N2546, N2042, N2510, N1025);
nor NOR4 (N2551, N2547, N1017, N747, N2369);
buf BUF1 (N2552, N2548);
nand NAND3 (N2553, N2530, N1818, N121);
not NOT1 (N2554, N2549);
and AND4 (N2555, N2551, N534, N802, N2367);
xor XOR2 (N2556, N2529, N1340);
buf BUF1 (N2557, N2511);
and AND4 (N2558, N2550, N1073, N2038, N762);
and AND3 (N2559, N2557, N1779, N1134);
nor NOR3 (N2560, N2559, N699, N1702);
not NOT1 (N2561, N2560);
and AND3 (N2562, N2553, N116, N2207);
xor XOR2 (N2563, N2556, N1083);
and AND3 (N2564, N2543, N1863, N510);
and AND2 (N2565, N2555, N1630);
buf BUF1 (N2566, N2561);
nand NAND4 (N2567, N2544, N1261, N925, N1269);
buf BUF1 (N2568, N2565);
nand NAND4 (N2569, N2564, N384, N56, N2477);
nor NOR3 (N2570, N2562, N352, N2355);
and AND3 (N2571, N2552, N1979, N1731);
nand NAND2 (N2572, N2554, N433);
nor NOR4 (N2573, N2571, N2077, N590, N840);
xor XOR2 (N2574, N2567, N734);
or OR3 (N2575, N2568, N868, N1921);
nor NOR4 (N2576, N2573, N2307, N2284, N621);
buf BUF1 (N2577, N2572);
not NOT1 (N2578, N2576);
buf BUF1 (N2579, N2577);
buf BUF1 (N2580, N2570);
not NOT1 (N2581, N2563);
xor XOR2 (N2582, N2578, N28);
and AND4 (N2583, N2581, N2153, N1064, N2155);
and AND4 (N2584, N2575, N696, N1797, N1160);
nand NAND2 (N2585, N2569, N804);
not NOT1 (N2586, N2584);
buf BUF1 (N2587, N2583);
or OR4 (N2588, N2558, N1784, N795, N928);
xor XOR2 (N2589, N2566, N1214);
xor XOR2 (N2590, N2574, N1819);
xor XOR2 (N2591, N2582, N1655);
nand NAND2 (N2592, N2580, N440);
nor NOR3 (N2593, N2579, N2031, N2326);
buf BUF1 (N2594, N2588);
and AND3 (N2595, N2591, N572, N1497);
and AND4 (N2596, N2593, N10, N370, N2029);
not NOT1 (N2597, N2587);
or OR4 (N2598, N2594, N2047, N1922, N2341);
or OR4 (N2599, N2597, N178, N476, N443);
xor XOR2 (N2600, N2585, N815);
xor XOR2 (N2601, N2589, N2100);
buf BUF1 (N2602, N2596);
buf BUF1 (N2603, N2586);
nor NOR4 (N2604, N2532, N591, N1114, N1226);
nor NOR4 (N2605, N2595, N1083, N1078, N2456);
or OR2 (N2606, N2604, N1309);
nor NOR3 (N2607, N2590, N2011, N403);
not NOT1 (N2608, N2603);
not NOT1 (N2609, N2599);
or OR3 (N2610, N2602, N2136, N2051);
and AND3 (N2611, N2592, N1878, N2010);
and AND2 (N2612, N2598, N2149);
and AND4 (N2613, N2611, N1233, N354, N1799);
not NOT1 (N2614, N2610);
not NOT1 (N2615, N2613);
nand NAND3 (N2616, N2614, N2304, N1648);
xor XOR2 (N2617, N2605, N2385);
nor NOR4 (N2618, N2609, N1685, N983, N2110);
nor NOR3 (N2619, N2618, N2589, N1352);
nand NAND4 (N2620, N2617, N806, N321, N1161);
buf BUF1 (N2621, N2607);
xor XOR2 (N2622, N2620, N2148);
and AND3 (N2623, N2606, N1257, N1093);
buf BUF1 (N2624, N2621);
not NOT1 (N2625, N2623);
nor NOR3 (N2626, N2625, N2364, N526);
not NOT1 (N2627, N2622);
nor NOR3 (N2628, N2624, N137, N2597);
buf BUF1 (N2629, N2619);
buf BUF1 (N2630, N2600);
not NOT1 (N2631, N2626);
and AND3 (N2632, N2601, N2216, N1796);
or OR3 (N2633, N2616, N2241, N1984);
not NOT1 (N2634, N2632);
xor XOR2 (N2635, N2631, N295);
nand NAND2 (N2636, N2635, N1387);
nor NOR3 (N2637, N2634, N415, N636);
and AND4 (N2638, N2630, N480, N2150, N1067);
nor NOR4 (N2639, N2615, N53, N1927, N260);
buf BUF1 (N2640, N2629);
or OR4 (N2641, N2612, N888, N826, N1679);
and AND4 (N2642, N2627, N922, N2417, N2248);
buf BUF1 (N2643, N2640);
xor XOR2 (N2644, N2628, N925);
nand NAND3 (N2645, N2641, N2223, N2570);
buf BUF1 (N2646, N2633);
buf BUF1 (N2647, N2646);
not NOT1 (N2648, N2636);
and AND2 (N2649, N2643, N2203);
or OR4 (N2650, N2644, N1753, N1421, N1217);
or OR2 (N2651, N2637, N506);
and AND3 (N2652, N2638, N893, N2371);
xor XOR2 (N2653, N2648, N153);
nand NAND3 (N2654, N2653, N1272, N630);
nand NAND3 (N2655, N2649, N2371, N791);
nand NAND4 (N2656, N2650, N1090, N2551, N1620);
xor XOR2 (N2657, N2656, N1190);
not NOT1 (N2658, N2657);
nor NOR4 (N2659, N2655, N1120, N214, N2422);
or OR3 (N2660, N2642, N1275, N1113);
nand NAND3 (N2661, N2658, N1921, N1489);
not NOT1 (N2662, N2639);
not NOT1 (N2663, N2647);
buf BUF1 (N2664, N2608);
and AND3 (N2665, N2661, N465, N150);
nand NAND3 (N2666, N2652, N1371, N869);
nand NAND2 (N2667, N2666, N1192);
buf BUF1 (N2668, N2664);
or OR2 (N2669, N2645, N269);
nand NAND2 (N2670, N2663, N313);
and AND3 (N2671, N2669, N1249, N2239);
or OR4 (N2672, N2670, N1288, N2620, N2612);
and AND3 (N2673, N2668, N255, N2192);
or OR3 (N2674, N2667, N857, N2569);
buf BUF1 (N2675, N2651);
or OR2 (N2676, N2675, N706);
and AND4 (N2677, N2659, N2187, N1163, N818);
xor XOR2 (N2678, N2672, N1680);
xor XOR2 (N2679, N2676, N606);
nand NAND4 (N2680, N2673, N897, N1579, N2442);
or OR4 (N2681, N2678, N2152, N1390, N1371);
not NOT1 (N2682, N2660);
and AND3 (N2683, N2674, N758, N2236);
and AND2 (N2684, N2654, N1371);
not NOT1 (N2685, N2665);
or OR2 (N2686, N2662, N1468);
and AND3 (N2687, N2684, N54, N2530);
and AND4 (N2688, N2685, N1537, N1045, N473);
xor XOR2 (N2689, N2682, N576);
not NOT1 (N2690, N2689);
and AND2 (N2691, N2686, N1387);
nor NOR4 (N2692, N2680, N446, N662, N2568);
xor XOR2 (N2693, N2691, N258);
and AND4 (N2694, N2692, N252, N636, N1253);
not NOT1 (N2695, N2679);
xor XOR2 (N2696, N2694, N1511);
or OR2 (N2697, N2677, N1189);
or OR3 (N2698, N2681, N772, N2402);
nor NOR4 (N2699, N2690, N931, N2421, N747);
buf BUF1 (N2700, N2699);
nand NAND4 (N2701, N2697, N887, N137, N1125);
and AND2 (N2702, N2698, N1075);
and AND3 (N2703, N2671, N2251, N1760);
and AND2 (N2704, N2687, N1781);
nand NAND4 (N2705, N2696, N779, N688, N843);
nand NAND2 (N2706, N2702, N876);
buf BUF1 (N2707, N2706);
nor NOR4 (N2708, N2683, N1023, N2555, N958);
xor XOR2 (N2709, N2704, N117);
buf BUF1 (N2710, N2709);
nand NAND3 (N2711, N2710, N1673, N2354);
buf BUF1 (N2712, N2701);
nand NAND2 (N2713, N2688, N1993);
nor NOR3 (N2714, N2693, N2020, N2617);
nand NAND3 (N2715, N2705, N295, N354);
xor XOR2 (N2716, N2715, N2193);
xor XOR2 (N2717, N2716, N218);
nand NAND3 (N2718, N2700, N1552, N1742);
and AND3 (N2719, N2714, N325, N906);
and AND4 (N2720, N2711, N1322, N2174, N298);
and AND2 (N2721, N2719, N2128);
and AND4 (N2722, N2708, N1204, N910, N1472);
nand NAND4 (N2723, N2695, N1362, N2467, N100);
or OR3 (N2724, N2713, N543, N1750);
or OR4 (N2725, N2723, N2420, N1586, N1207);
or OR2 (N2726, N2717, N1845);
not NOT1 (N2727, N2707);
nor NOR3 (N2728, N2703, N1592, N1875);
and AND4 (N2729, N2725, N2332, N256, N2121);
or OR4 (N2730, N2722, N2280, N1482, N1868);
nor NOR3 (N2731, N2721, N996, N2256);
xor XOR2 (N2732, N2731, N188);
nand NAND4 (N2733, N2732, N896, N1606, N1078);
nor NOR2 (N2734, N2712, N606);
or OR3 (N2735, N2726, N1572, N2595);
or OR4 (N2736, N2733, N616, N2648, N1953);
not NOT1 (N2737, N2724);
nor NOR2 (N2738, N2735, N241);
and AND2 (N2739, N2718, N214);
xor XOR2 (N2740, N2737, N573);
buf BUF1 (N2741, N2740);
nor NOR2 (N2742, N2730, N1675);
buf BUF1 (N2743, N2736);
and AND2 (N2744, N2738, N2103);
nor NOR2 (N2745, N2744, N2282);
nand NAND2 (N2746, N2745, N767);
nor NOR3 (N2747, N2727, N2116, N666);
not NOT1 (N2748, N2729);
nor NOR2 (N2749, N2747, N1323);
not NOT1 (N2750, N2739);
buf BUF1 (N2751, N2742);
and AND3 (N2752, N2748, N1647, N2471);
and AND3 (N2753, N2750, N1087, N624);
nand NAND2 (N2754, N2752, N2182);
buf BUF1 (N2755, N2754);
nand NAND2 (N2756, N2720, N1592);
or OR4 (N2757, N2753, N106, N2224, N2139);
not NOT1 (N2758, N2749);
buf BUF1 (N2759, N2746);
not NOT1 (N2760, N2759);
xor XOR2 (N2761, N2756, N2754);
not NOT1 (N2762, N2761);
or OR4 (N2763, N2758, N185, N1434, N2110);
or OR4 (N2764, N2728, N1118, N2462, N813);
buf BUF1 (N2765, N2762);
nor NOR4 (N2766, N2734, N1633, N2272, N1321);
buf BUF1 (N2767, N2741);
and AND2 (N2768, N2743, N1538);
not NOT1 (N2769, N2751);
xor XOR2 (N2770, N2755, N18);
or OR3 (N2771, N2767, N89, N1337);
or OR2 (N2772, N2760, N410);
xor XOR2 (N2773, N2771, N1426);
xor XOR2 (N2774, N2770, N1118);
not NOT1 (N2775, N2768);
and AND2 (N2776, N2764, N313);
buf BUF1 (N2777, N2763);
nor NOR2 (N2778, N2773, N1961);
and AND4 (N2779, N2766, N2387, N1906, N912);
not NOT1 (N2780, N2776);
not NOT1 (N2781, N2775);
nor NOR2 (N2782, N2765, N581);
nand NAND4 (N2783, N2772, N2660, N2618, N2441);
nand NAND2 (N2784, N2777, N294);
buf BUF1 (N2785, N2783);
xor XOR2 (N2786, N2778, N438);
or OR2 (N2787, N2782, N2077);
or OR2 (N2788, N2780, N827);
xor XOR2 (N2789, N2757, N2033);
nand NAND4 (N2790, N2784, N1709, N947, N154);
nor NOR2 (N2791, N2785, N273);
xor XOR2 (N2792, N2790, N553);
nand NAND3 (N2793, N2774, N865, N2276);
and AND2 (N2794, N2781, N2264);
or OR2 (N2795, N2794, N2058);
and AND4 (N2796, N2795, N106, N1221, N141);
buf BUF1 (N2797, N2788);
and AND3 (N2798, N2791, N329, N1596);
buf BUF1 (N2799, N2769);
and AND2 (N2800, N2789, N1412);
not NOT1 (N2801, N2799);
or OR3 (N2802, N2787, N2769, N2528);
and AND4 (N2803, N2797, N1748, N2774, N896);
nand NAND3 (N2804, N2786, N625, N440);
nor NOR3 (N2805, N2796, N847, N987);
buf BUF1 (N2806, N2804);
nand NAND3 (N2807, N2798, N2722, N985);
buf BUF1 (N2808, N2805);
nor NOR3 (N2809, N2806, N454, N1868);
or OR3 (N2810, N2809, N166, N1873);
xor XOR2 (N2811, N2801, N1885);
or OR2 (N2812, N2803, N498);
xor XOR2 (N2813, N2811, N1865);
nor NOR4 (N2814, N2808, N1491, N2400, N1868);
and AND3 (N2815, N2812, N1849, N1118);
nor NOR2 (N2816, N2779, N173);
nand NAND2 (N2817, N2816, N1589);
xor XOR2 (N2818, N2807, N303);
xor XOR2 (N2819, N2815, N1786);
nand NAND4 (N2820, N2818, N1341, N2095, N201);
nor NOR3 (N2821, N2793, N323, N133);
buf BUF1 (N2822, N2800);
buf BUF1 (N2823, N2817);
buf BUF1 (N2824, N2810);
and AND4 (N2825, N2792, N2604, N1973, N376);
and AND2 (N2826, N2824, N942);
xor XOR2 (N2827, N2820, N1705);
xor XOR2 (N2828, N2822, N379);
and AND2 (N2829, N2802, N1556);
and AND2 (N2830, N2827, N1100);
nor NOR2 (N2831, N2828, N1781);
and AND3 (N2832, N2825, N2133, N1373);
not NOT1 (N2833, N2826);
xor XOR2 (N2834, N2833, N1614);
xor XOR2 (N2835, N2819, N2278);
xor XOR2 (N2836, N2829, N1762);
buf BUF1 (N2837, N2831);
buf BUF1 (N2838, N2823);
nand NAND3 (N2839, N2836, N332, N176);
nor NOR4 (N2840, N2834, N2004, N112, N58);
nand NAND4 (N2841, N2839, N1429, N1467, N2356);
not NOT1 (N2842, N2837);
and AND4 (N2843, N2832, N1019, N2351, N1339);
buf BUF1 (N2844, N2838);
buf BUF1 (N2845, N2813);
buf BUF1 (N2846, N2840);
and AND3 (N2847, N2821, N1876, N2639);
and AND3 (N2848, N2830, N1683, N672);
nand NAND2 (N2849, N2814, N1620);
nand NAND4 (N2850, N2849, N1907, N69, N1404);
and AND2 (N2851, N2835, N1181);
not NOT1 (N2852, N2847);
not NOT1 (N2853, N2850);
not NOT1 (N2854, N2843);
nor NOR4 (N2855, N2846, N804, N1701, N2838);
nand NAND3 (N2856, N2852, N1236, N2514);
nor NOR2 (N2857, N2841, N1548);
xor XOR2 (N2858, N2857, N2775);
xor XOR2 (N2859, N2856, N2278);
or OR3 (N2860, N2844, N1969, N1967);
and AND4 (N2861, N2845, N594, N2647, N2066);
or OR3 (N2862, N2861, N1525, N2765);
or OR3 (N2863, N2858, N1334, N2842);
nand NAND2 (N2864, N1546, N1075);
not NOT1 (N2865, N2864);
xor XOR2 (N2866, N2863, N2416);
nand NAND2 (N2867, N2853, N595);
not NOT1 (N2868, N2848);
or OR3 (N2869, N2868, N2396, N235);
and AND2 (N2870, N2865, N2296);
and AND2 (N2871, N2851, N2323);
buf BUF1 (N2872, N2869);
and AND3 (N2873, N2855, N532, N1137);
xor XOR2 (N2874, N2866, N2035);
nand NAND3 (N2875, N2870, N820, N2031);
xor XOR2 (N2876, N2860, N2095);
not NOT1 (N2877, N2871);
not NOT1 (N2878, N2854);
or OR4 (N2879, N2867, N2117, N1974, N2257);
xor XOR2 (N2880, N2872, N2844);
nand NAND3 (N2881, N2874, N2319, N1781);
nand NAND4 (N2882, N2862, N2254, N972, N1763);
nor NOR3 (N2883, N2879, N1564, N2134);
or OR3 (N2884, N2883, N120, N2542);
xor XOR2 (N2885, N2875, N2444);
xor XOR2 (N2886, N2882, N884);
nand NAND2 (N2887, N2886, N1101);
and AND4 (N2888, N2880, N549, N1001, N1972);
xor XOR2 (N2889, N2881, N1415);
buf BUF1 (N2890, N2888);
not NOT1 (N2891, N2877);
or OR3 (N2892, N2876, N642, N843);
nand NAND2 (N2893, N2859, N2627);
nand NAND4 (N2894, N2889, N2602, N789, N1578);
or OR4 (N2895, N2890, N330, N1961, N1172);
or OR2 (N2896, N2893, N953);
or OR4 (N2897, N2873, N2104, N1392, N1370);
or OR4 (N2898, N2885, N2390, N333, N767);
or OR3 (N2899, N2897, N1235, N616);
buf BUF1 (N2900, N2894);
xor XOR2 (N2901, N2887, N2280);
or OR2 (N2902, N2895, N2226);
nor NOR2 (N2903, N2899, N1765);
or OR2 (N2904, N2902, N948);
nor NOR2 (N2905, N2896, N2047);
nand NAND3 (N2906, N2884, N2125, N1700);
buf BUF1 (N2907, N2892);
nand NAND2 (N2908, N2904, N1653);
xor XOR2 (N2909, N2907, N2771);
nor NOR3 (N2910, N2898, N1409, N886);
not NOT1 (N2911, N2906);
buf BUF1 (N2912, N2903);
nor NOR2 (N2913, N2912, N1838);
not NOT1 (N2914, N2905);
nor NOR4 (N2915, N2878, N977, N445, N2139);
or OR4 (N2916, N2901, N378, N632, N2679);
or OR4 (N2917, N2915, N2063, N1768, N2593);
nor NOR4 (N2918, N2914, N2793, N1539, N48);
nor NOR3 (N2919, N2909, N2825, N2243);
nor NOR3 (N2920, N2917, N18, N2730);
nor NOR3 (N2921, N2910, N2362, N2809);
not NOT1 (N2922, N2921);
xor XOR2 (N2923, N2913, N714);
nor NOR2 (N2924, N2916, N2029);
xor XOR2 (N2925, N2908, N1578);
nor NOR4 (N2926, N2891, N1549, N290, N2174);
nor NOR4 (N2927, N2911, N937, N2760, N2076);
not NOT1 (N2928, N2900);
nor NOR2 (N2929, N2923, N1538);
xor XOR2 (N2930, N2918, N253);
buf BUF1 (N2931, N2922);
buf BUF1 (N2932, N2925);
nand NAND2 (N2933, N2928, N1575);
not NOT1 (N2934, N2924);
nand NAND2 (N2935, N2926, N2404);
and AND4 (N2936, N2919, N2418, N1569, N881);
or OR2 (N2937, N2931, N118);
xor XOR2 (N2938, N2935, N1982);
buf BUF1 (N2939, N2927);
nand NAND4 (N2940, N2938, N1874, N1407, N1721);
or OR3 (N2941, N2939, N1613, N1783);
xor XOR2 (N2942, N2920, N2774);
xor XOR2 (N2943, N2934, N2357);
nand NAND4 (N2944, N2929, N2865, N1328, N2512);
nor NOR4 (N2945, N2943, N2333, N477, N2359);
or OR2 (N2946, N2937, N1627);
and AND4 (N2947, N2933, N2591, N1221, N2397);
xor XOR2 (N2948, N2947, N1047);
nand NAND3 (N2949, N2940, N1074, N989);
nor NOR2 (N2950, N2945, N2413);
nand NAND3 (N2951, N2936, N2459, N548);
buf BUF1 (N2952, N2950);
not NOT1 (N2953, N2941);
nor NOR2 (N2954, N2942, N2925);
not NOT1 (N2955, N2954);
xor XOR2 (N2956, N2952, N2518);
buf BUF1 (N2957, N2951);
and AND4 (N2958, N2949, N1197, N1689, N1392);
and AND4 (N2959, N2932, N418, N1087, N2268);
not NOT1 (N2960, N2959);
nand NAND3 (N2961, N2956, N649, N2861);
and AND2 (N2962, N2930, N749);
buf BUF1 (N2963, N2962);
nand NAND3 (N2964, N2944, N1384, N66);
or OR3 (N2965, N2955, N288, N1606);
nor NOR3 (N2966, N2964, N880, N2356);
xor XOR2 (N2967, N2948, N1802);
or OR3 (N2968, N2966, N587, N386);
not NOT1 (N2969, N2961);
xor XOR2 (N2970, N2963, N907);
xor XOR2 (N2971, N2970, N71);
xor XOR2 (N2972, N2960, N560);
nor NOR2 (N2973, N2965, N967);
not NOT1 (N2974, N2958);
not NOT1 (N2975, N2973);
buf BUF1 (N2976, N2974);
nor NOR3 (N2977, N2953, N1197, N328);
xor XOR2 (N2978, N2968, N2387);
or OR4 (N2979, N2957, N1248, N2223, N2777);
buf BUF1 (N2980, N2975);
nand NAND3 (N2981, N2979, N1199, N359);
nand NAND4 (N2982, N2977, N2736, N1443, N1053);
nand NAND3 (N2983, N2980, N2262, N1397);
nand NAND4 (N2984, N2982, N689, N180, N2361);
nand NAND2 (N2985, N2976, N2023);
buf BUF1 (N2986, N2984);
nor NOR4 (N2987, N2971, N846, N2144, N1843);
not NOT1 (N2988, N2969);
not NOT1 (N2989, N2972);
buf BUF1 (N2990, N2988);
not NOT1 (N2991, N2981);
nor NOR4 (N2992, N2991, N2252, N331, N2521);
nor NOR3 (N2993, N2946, N2846, N841);
nor NOR4 (N2994, N2992, N2353, N711, N92);
and AND4 (N2995, N2967, N520, N1924, N1340);
nand NAND2 (N2996, N2993, N2086);
not NOT1 (N2997, N2994);
nand NAND3 (N2998, N2989, N903, N410);
xor XOR2 (N2999, N2997, N2512);
buf BUF1 (N3000, N2990);
or OR4 (N3001, N2998, N48, N2898, N1917);
and AND3 (N3002, N2995, N471, N1487);
or OR4 (N3003, N3002, N348, N1701, N335);
buf BUF1 (N3004, N2986);
xor XOR2 (N3005, N2978, N2529);
not NOT1 (N3006, N3004);
buf BUF1 (N3007, N3006);
or OR4 (N3008, N3000, N2590, N2045, N1809);
nand NAND3 (N3009, N2985, N2102, N16);
nor NOR3 (N3010, N3009, N1162, N2672);
not NOT1 (N3011, N2983);
or OR3 (N3012, N3003, N287, N1587);
or OR4 (N3013, N3001, N2261, N1490, N2025);
xor XOR2 (N3014, N2987, N702);
nor NOR3 (N3015, N2996, N2053, N9);
xor XOR2 (N3016, N3008, N1160);
buf BUF1 (N3017, N3012);
and AND4 (N3018, N3014, N1795, N2831, N632);
not NOT1 (N3019, N3015);
nand NAND2 (N3020, N3011, N2517);
and AND2 (N3021, N3013, N73);
nor NOR3 (N3022, N3010, N528, N2542);
and AND3 (N3023, N3020, N213, N171);
nor NOR2 (N3024, N3018, N901);
and AND2 (N3025, N3024, N2066);
nand NAND2 (N3026, N3022, N2757);
buf BUF1 (N3027, N3017);
or OR4 (N3028, N3027, N2557, N2342, N292);
buf BUF1 (N3029, N3023);
not NOT1 (N3030, N3005);
or OR3 (N3031, N3030, N2422, N2822);
buf BUF1 (N3032, N3025);
or OR2 (N3033, N3016, N2882);
or OR4 (N3034, N3026, N1401, N2883, N157);
not NOT1 (N3035, N2999);
not NOT1 (N3036, N3019);
buf BUF1 (N3037, N3007);
not NOT1 (N3038, N3035);
nor NOR3 (N3039, N3034, N1553, N1580);
and AND2 (N3040, N3032, N2765);
and AND4 (N3041, N3036, N751, N762, N1213);
or OR4 (N3042, N3021, N1705, N2314, N1768);
or OR2 (N3043, N3038, N1955);
nor NOR4 (N3044, N3042, N34, N249, N1693);
or OR4 (N3045, N3043, N1495, N1378, N836);
not NOT1 (N3046, N3040);
nand NAND4 (N3047, N3037, N335, N2387, N559);
nand NAND2 (N3048, N3031, N20);
and AND2 (N3049, N3033, N1777);
not NOT1 (N3050, N3049);
and AND2 (N3051, N3039, N269);
and AND2 (N3052, N3048, N108);
nand NAND3 (N3053, N3052, N2856, N153);
not NOT1 (N3054, N3028);
nand NAND4 (N3055, N3045, N2080, N2894, N67);
buf BUF1 (N3056, N3044);
buf BUF1 (N3057, N3051);
buf BUF1 (N3058, N3056);
xor XOR2 (N3059, N3055, N1273);
xor XOR2 (N3060, N3059, N1928);
xor XOR2 (N3061, N3047, N149);
nand NAND3 (N3062, N3060, N1314, N2934);
not NOT1 (N3063, N3054);
or OR4 (N3064, N3029, N2241, N222, N2402);
or OR2 (N3065, N3064, N715);
buf BUF1 (N3066, N3062);
nor NOR3 (N3067, N3053, N670, N1469);
not NOT1 (N3068, N3065);
nand NAND4 (N3069, N3058, N363, N469, N214);
nand NAND4 (N3070, N3063, N2668, N2578, N451);
buf BUF1 (N3071, N3041);
nor NOR4 (N3072, N3068, N1825, N427, N133);
nor NOR3 (N3073, N3057, N1563, N2799);
nand NAND2 (N3074, N3073, N2834);
nand NAND3 (N3075, N3061, N1387, N907);
buf BUF1 (N3076, N3072);
xor XOR2 (N3077, N3066, N376);
xor XOR2 (N3078, N3067, N1237);
or OR4 (N3079, N3075, N1804, N813, N2573);
buf BUF1 (N3080, N3070);
not NOT1 (N3081, N3050);
and AND2 (N3082, N3076, N600);
xor XOR2 (N3083, N3071, N2933);
nor NOR3 (N3084, N3046, N1308, N2250);
nor NOR2 (N3085, N3079, N2616);
nand NAND3 (N3086, N3069, N1273, N59);
buf BUF1 (N3087, N3080);
nand NAND3 (N3088, N3085, N772, N2887);
and AND4 (N3089, N3084, N1161, N481, N838);
buf BUF1 (N3090, N3074);
nand NAND3 (N3091, N3082, N2291, N711);
nand NAND3 (N3092, N3089, N1581, N1843);
nor NOR2 (N3093, N3083, N1317);
and AND3 (N3094, N3086, N23, N128);
nand NAND4 (N3095, N3088, N2949, N1530, N2027);
xor XOR2 (N3096, N3092, N2011);
and AND4 (N3097, N3091, N429, N1907, N797);
buf BUF1 (N3098, N3097);
and AND4 (N3099, N3087, N1355, N1081, N1912);
or OR4 (N3100, N3094, N1862, N2835, N1881);
not NOT1 (N3101, N3096);
not NOT1 (N3102, N3077);
nor NOR2 (N3103, N3090, N448);
not NOT1 (N3104, N3099);
or OR4 (N3105, N3100, N121, N1808, N167);
nor NOR3 (N3106, N3102, N3092, N1608);
nor NOR2 (N3107, N3101, N682);
and AND4 (N3108, N3104, N1846, N2988, N2571);
and AND3 (N3109, N3105, N1194, N1935);
nand NAND3 (N3110, N3081, N2093, N552);
nor NOR4 (N3111, N3095, N1105, N2208, N1025);
not NOT1 (N3112, N3098);
not NOT1 (N3113, N3093);
not NOT1 (N3114, N3112);
not NOT1 (N3115, N3114);
and AND3 (N3116, N3108, N2603, N2524);
and AND3 (N3117, N3115, N2554, N2473);
xor XOR2 (N3118, N3111, N2170);
buf BUF1 (N3119, N3110);
nor NOR4 (N3120, N3118, N2510, N834, N424);
nand NAND4 (N3121, N3119, N2484, N2653, N1299);
or OR3 (N3122, N3113, N2030, N1371);
not NOT1 (N3123, N3107);
nor NOR3 (N3124, N3120, N1399, N171);
or OR4 (N3125, N3117, N41, N3005, N2000);
and AND4 (N3126, N3121, N2550, N3058, N2033);
or OR3 (N3127, N3125, N431, N2453);
or OR3 (N3128, N3123, N593, N2959);
not NOT1 (N3129, N3127);
or OR3 (N3130, N3103, N374, N2150);
or OR2 (N3131, N3126, N385);
buf BUF1 (N3132, N3078);
nor NOR4 (N3133, N3116, N2309, N2046, N2891);
and AND3 (N3134, N3124, N181, N1958);
xor XOR2 (N3135, N3128, N663);
xor XOR2 (N3136, N3133, N613);
buf BUF1 (N3137, N3109);
xor XOR2 (N3138, N3106, N1310);
or OR4 (N3139, N3129, N1510, N1013, N286);
or OR4 (N3140, N3132, N1354, N3011, N115);
xor XOR2 (N3141, N3138, N247);
or OR2 (N3142, N3139, N1545);
and AND2 (N3143, N3141, N894);
xor XOR2 (N3144, N3131, N2578);
not NOT1 (N3145, N3122);
buf BUF1 (N3146, N3135);
and AND2 (N3147, N3143, N1723);
nand NAND3 (N3148, N3134, N182, N2357);
nor NOR4 (N3149, N3140, N2825, N1220, N2840);
buf BUF1 (N3150, N3136);
not NOT1 (N3151, N3142);
and AND2 (N3152, N3144, N180);
nand NAND2 (N3153, N3151, N1326);
not NOT1 (N3154, N3152);
nand NAND2 (N3155, N3145, N997);
not NOT1 (N3156, N3149);
nor NOR4 (N3157, N3156, N2478, N1862, N843);
nor NOR2 (N3158, N3130, N1734);
nand NAND3 (N3159, N3146, N1329, N1316);
or OR4 (N3160, N3158, N2271, N1130, N125);
buf BUF1 (N3161, N3147);
buf BUF1 (N3162, N3153);
nor NOR4 (N3163, N3150, N1814, N2445, N1532);
or OR4 (N3164, N3157, N2336, N2843, N1017);
and AND4 (N3165, N3159, N236, N188, N782);
nor NOR3 (N3166, N3163, N1564, N2578);
buf BUF1 (N3167, N3161);
not NOT1 (N3168, N3137);
and AND4 (N3169, N3167, N1545, N3029, N2033);
nand NAND4 (N3170, N3160, N715, N254, N2021);
or OR4 (N3171, N3170, N2008, N513, N2649);
buf BUF1 (N3172, N3168);
and AND2 (N3173, N3155, N410);
not NOT1 (N3174, N3162);
xor XOR2 (N3175, N3164, N1309);
not NOT1 (N3176, N3165);
xor XOR2 (N3177, N3169, N272);
not NOT1 (N3178, N3171);
buf BUF1 (N3179, N3175);
nor NOR2 (N3180, N3178, N813);
xor XOR2 (N3181, N3179, N1500);
nor NOR2 (N3182, N3174, N2117);
nand NAND2 (N3183, N3181, N3010);
nand NAND3 (N3184, N3176, N551, N3080);
or OR3 (N3185, N3177, N2134, N877);
nor NOR3 (N3186, N3172, N2112, N2924);
not NOT1 (N3187, N3148);
xor XOR2 (N3188, N3184, N35);
not NOT1 (N3189, N3180);
and AND3 (N3190, N3183, N1843, N2908);
and AND2 (N3191, N3173, N1925);
xor XOR2 (N3192, N3186, N1649);
and AND2 (N3193, N3188, N1955);
nor NOR2 (N3194, N3154, N1086);
nor NOR2 (N3195, N3193, N2879);
and AND2 (N3196, N3185, N2493);
nand NAND3 (N3197, N3195, N1895, N2191);
buf BUF1 (N3198, N3192);
nor NOR3 (N3199, N3187, N124, N2503);
nor NOR2 (N3200, N3196, N3099);
or OR4 (N3201, N3200, N573, N947, N2456);
nand NAND2 (N3202, N3198, N1701);
buf BUF1 (N3203, N3182);
not NOT1 (N3204, N3189);
or OR2 (N3205, N3204, N4);
not NOT1 (N3206, N3197);
and AND4 (N3207, N3194, N1019, N2885, N2678);
and AND4 (N3208, N3203, N1679, N2051, N2228);
not NOT1 (N3209, N3202);
xor XOR2 (N3210, N3166, N2644);
nand NAND3 (N3211, N3205, N1063, N3126);
xor XOR2 (N3212, N3191, N538);
nor NOR2 (N3213, N3209, N1591);
buf BUF1 (N3214, N3190);
or OR4 (N3215, N3201, N1234, N722, N2194);
nand NAND2 (N3216, N3212, N2487);
buf BUF1 (N3217, N3207);
nand NAND2 (N3218, N3215, N2700);
xor XOR2 (N3219, N3217, N350);
not NOT1 (N3220, N3206);
nor NOR4 (N3221, N3199, N1323, N1143, N2209);
endmodule