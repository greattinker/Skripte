// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N3218,N3211,N3212,N3215,N3217,N3202,N3209,N3197,N3210,N3219;

and AND4 (N20, N8, N13, N16, N18);
xor XOR2 (N21, N15, N18);
or OR4 (N22, N16, N20, N9, N3);
xor XOR2 (N23, N9, N21);
or OR2 (N24, N4, N2);
nor NOR3 (N25, N7, N10, N7);
nor NOR2 (N26, N18, N1);
buf BUF1 (N27, N25);
not NOT1 (N28, N1);
and AND4 (N29, N23, N25, N24, N15);
nor NOR2 (N30, N28, N15);
or OR4 (N31, N29, N10, N17, N1);
nor NOR4 (N32, N17, N31, N3, N3);
buf BUF1 (N33, N3);
or OR2 (N34, N25, N18);
nand NAND4 (N35, N9, N23, N7, N10);
xor XOR2 (N36, N2, N4);
nand NAND3 (N37, N29, N15, N6);
and AND3 (N38, N30, N13, N9);
not NOT1 (N39, N27);
not NOT1 (N40, N34);
buf BUF1 (N41, N32);
nand NAND3 (N42, N39, N38, N41);
or OR2 (N43, N20, N31);
nor NOR4 (N44, N31, N21, N28, N9);
nand NAND2 (N45, N36, N4);
buf BUF1 (N46, N45);
nor NOR3 (N47, N42, N27, N43);
not NOT1 (N48, N5);
nor NOR4 (N49, N26, N9, N4, N33);
buf BUF1 (N50, N31);
and AND4 (N51, N48, N1, N20, N30);
nand NAND4 (N52, N37, N26, N51, N37);
nor NOR3 (N53, N8, N7, N1);
not NOT1 (N54, N22);
xor XOR2 (N55, N40, N53);
and AND3 (N56, N34, N22, N23);
buf BUF1 (N57, N35);
nand NAND2 (N58, N47, N33);
buf BUF1 (N59, N57);
or OR3 (N60, N56, N2, N14);
or OR3 (N61, N46, N49, N44);
buf BUF1 (N62, N38);
and AND2 (N63, N38, N18);
buf BUF1 (N64, N61);
buf BUF1 (N65, N54);
nand NAND2 (N66, N65, N56);
and AND4 (N67, N50, N43, N42, N39);
or OR4 (N68, N60, N2, N28, N47);
buf BUF1 (N69, N52);
nand NAND3 (N70, N64, N32, N42);
nor NOR2 (N71, N66, N34);
buf BUF1 (N72, N63);
not NOT1 (N73, N68);
not NOT1 (N74, N71);
xor XOR2 (N75, N73, N4);
buf BUF1 (N76, N72);
and AND3 (N77, N74, N50, N36);
or OR2 (N78, N75, N33);
nor NOR2 (N79, N58, N69);
not NOT1 (N80, N58);
nor NOR3 (N81, N77, N4, N50);
and AND4 (N82, N62, N66, N35, N71);
nand NAND2 (N83, N82, N10);
nor NOR3 (N84, N67, N20, N39);
buf BUF1 (N85, N84);
buf BUF1 (N86, N80);
not NOT1 (N87, N55);
nor NOR3 (N88, N59, N33, N12);
buf BUF1 (N89, N86);
or OR3 (N90, N70, N6, N89);
and AND4 (N91, N20, N34, N48, N85);
not NOT1 (N92, N74);
nor NOR4 (N93, N87, N35, N20, N50);
or OR2 (N94, N92, N28);
buf BUF1 (N95, N76);
nand NAND2 (N96, N95, N75);
xor XOR2 (N97, N96, N42);
nand NAND2 (N98, N90, N29);
xor XOR2 (N99, N91, N48);
not NOT1 (N100, N97);
and AND4 (N101, N88, N22, N12, N15);
and AND4 (N102, N99, N11, N38, N73);
nand NAND3 (N103, N83, N38, N6);
or OR4 (N104, N94, N47, N30, N57);
not NOT1 (N105, N102);
or OR3 (N106, N78, N22, N9);
nor NOR4 (N107, N81, N4, N83, N28);
and AND4 (N108, N104, N92, N67, N94);
and AND2 (N109, N106, N46);
xor XOR2 (N110, N93, N47);
xor XOR2 (N111, N103, N85);
nand NAND3 (N112, N107, N40, N109);
and AND4 (N113, N97, N106, N106, N45);
buf BUF1 (N114, N105);
not NOT1 (N115, N110);
and AND2 (N116, N108, N69);
xor XOR2 (N117, N115, N44);
buf BUF1 (N118, N116);
nand NAND4 (N119, N114, N95, N116, N44);
and AND2 (N120, N100, N70);
xor XOR2 (N121, N112, N87);
not NOT1 (N122, N113);
and AND2 (N123, N98, N105);
nor NOR3 (N124, N117, N39, N15);
or OR2 (N125, N121, N106);
and AND2 (N126, N119, N48);
nand NAND3 (N127, N79, N103, N30);
nand NAND2 (N128, N101, N11);
not NOT1 (N129, N118);
not NOT1 (N130, N127);
nand NAND3 (N131, N128, N118, N45);
buf BUF1 (N132, N125);
buf BUF1 (N133, N123);
or OR3 (N134, N124, N61, N96);
nand NAND2 (N135, N133, N38);
nor NOR2 (N136, N132, N85);
nand NAND3 (N137, N129, N91, N29);
nor NOR2 (N138, N134, N107);
or OR4 (N139, N122, N49, N5, N92);
and AND3 (N140, N135, N88, N119);
nand NAND3 (N141, N138, N106, N139);
xor XOR2 (N142, N47, N100);
nor NOR2 (N143, N111, N123);
or OR3 (N144, N120, N60, N14);
buf BUF1 (N145, N140);
xor XOR2 (N146, N130, N95);
and AND3 (N147, N145, N29, N70);
not NOT1 (N148, N142);
and AND3 (N149, N136, N22, N13);
nand NAND3 (N150, N148, N57, N146);
and AND3 (N151, N125, N146, N23);
nor NOR3 (N152, N143, N104, N79);
or OR2 (N153, N150, N62);
xor XOR2 (N154, N137, N69);
and AND3 (N155, N152, N135, N11);
nor NOR3 (N156, N144, N90, N32);
buf BUF1 (N157, N149);
or OR2 (N158, N154, N23);
xor XOR2 (N159, N153, N43);
or OR3 (N160, N147, N92, N159);
and AND4 (N161, N157, N10, N57, N115);
xor XOR2 (N162, N90, N147);
nand NAND2 (N163, N126, N47);
buf BUF1 (N164, N131);
buf BUF1 (N165, N160);
xor XOR2 (N166, N165, N146);
buf BUF1 (N167, N162);
buf BUF1 (N168, N163);
buf BUF1 (N169, N151);
buf BUF1 (N170, N156);
buf BUF1 (N171, N158);
not NOT1 (N172, N171);
nand NAND4 (N173, N172, N44, N5, N53);
nand NAND2 (N174, N166, N87);
buf BUF1 (N175, N167);
or OR3 (N176, N161, N67, N101);
xor XOR2 (N177, N164, N38);
buf BUF1 (N178, N177);
or OR3 (N179, N168, N152, N34);
or OR3 (N180, N169, N61, N6);
or OR2 (N181, N141, N90);
nor NOR3 (N182, N178, N165, N78);
and AND4 (N183, N174, N137, N101, N103);
nor NOR4 (N184, N173, N174, N95, N98);
nor NOR2 (N185, N176, N73);
and AND2 (N186, N170, N137);
not NOT1 (N187, N183);
nand NAND3 (N188, N181, N172, N72);
nand NAND3 (N189, N179, N60, N142);
nand NAND2 (N190, N188, N189);
nor NOR2 (N191, N28, N4);
or OR2 (N192, N175, N133);
nand NAND2 (N193, N184, N120);
buf BUF1 (N194, N186);
xor XOR2 (N195, N192, N86);
xor XOR2 (N196, N187, N11);
xor XOR2 (N197, N196, N189);
not NOT1 (N198, N191);
nor NOR2 (N199, N182, N60);
nor NOR2 (N200, N198, N61);
and AND3 (N201, N190, N70, N6);
not NOT1 (N202, N200);
buf BUF1 (N203, N185);
not NOT1 (N204, N195);
not NOT1 (N205, N204);
or OR4 (N206, N194, N141, N15, N165);
or OR2 (N207, N203, N13);
buf BUF1 (N208, N207);
buf BUF1 (N209, N155);
buf BUF1 (N210, N197);
nor NOR4 (N211, N209, N67, N176, N138);
buf BUF1 (N212, N193);
not NOT1 (N213, N210);
not NOT1 (N214, N201);
or OR3 (N215, N180, N107, N12);
not NOT1 (N216, N205);
buf BUF1 (N217, N214);
buf BUF1 (N218, N206);
nor NOR2 (N219, N217, N43);
nand NAND4 (N220, N215, N62, N151, N44);
not NOT1 (N221, N202);
nand NAND4 (N222, N220, N197, N171, N189);
nand NAND4 (N223, N208, N74, N167, N94);
xor XOR2 (N224, N223, N212);
or OR3 (N225, N2, N77, N100);
buf BUF1 (N226, N222);
or OR2 (N227, N213, N95);
not NOT1 (N228, N225);
xor XOR2 (N229, N227, N115);
nor NOR3 (N230, N226, N97, N8);
and AND4 (N231, N221, N37, N212, N137);
and AND3 (N232, N216, N222, N169);
xor XOR2 (N233, N218, N160);
not NOT1 (N234, N224);
and AND2 (N235, N229, N153);
not NOT1 (N236, N232);
or OR3 (N237, N219, N10, N8);
nand NAND2 (N238, N233, N196);
nor NOR2 (N239, N211, N170);
nor NOR3 (N240, N228, N237, N98);
nand NAND2 (N241, N134, N150);
buf BUF1 (N242, N241);
xor XOR2 (N243, N236, N126);
nor NOR4 (N244, N239, N236, N71, N72);
not NOT1 (N245, N243);
xor XOR2 (N246, N238, N231);
not NOT1 (N247, N43);
or OR2 (N248, N244, N31);
buf BUF1 (N249, N235);
not NOT1 (N250, N246);
nor NOR4 (N251, N249, N78, N169, N81);
nor NOR3 (N252, N251, N46, N239);
nor NOR3 (N253, N199, N28, N213);
and AND3 (N254, N240, N3, N204);
or OR3 (N255, N254, N175, N143);
or OR2 (N256, N253, N89);
and AND4 (N257, N256, N130, N186, N71);
buf BUF1 (N258, N250);
not NOT1 (N259, N252);
or OR3 (N260, N248, N117, N105);
xor XOR2 (N261, N255, N101);
xor XOR2 (N262, N245, N18);
nor NOR3 (N263, N230, N87, N128);
or OR3 (N264, N242, N30, N192);
buf BUF1 (N265, N264);
or OR3 (N266, N257, N135, N201);
or OR2 (N267, N262, N46);
xor XOR2 (N268, N258, N170);
xor XOR2 (N269, N247, N116);
xor XOR2 (N270, N268, N186);
or OR4 (N271, N269, N150, N123, N134);
and AND3 (N272, N270, N122, N237);
not NOT1 (N273, N263);
and AND2 (N274, N260, N119);
buf BUF1 (N275, N273);
nand NAND2 (N276, N271, N97);
or OR2 (N277, N234, N242);
not NOT1 (N278, N266);
xor XOR2 (N279, N267, N59);
nor NOR3 (N280, N276, N172, N129);
nor NOR4 (N281, N265, N249, N113, N129);
nor NOR2 (N282, N278, N129);
and AND2 (N283, N261, N46);
or OR3 (N284, N282, N230, N40);
buf BUF1 (N285, N279);
or OR3 (N286, N275, N155, N185);
xor XOR2 (N287, N281, N58);
nand NAND3 (N288, N259, N115, N39);
or OR4 (N289, N277, N113, N13, N33);
nand NAND3 (N290, N272, N173, N219);
not NOT1 (N291, N284);
nor NOR4 (N292, N288, N225, N81, N189);
or OR2 (N293, N283, N97);
nand NAND3 (N294, N292, N232, N290);
xor XOR2 (N295, N200, N273);
and AND3 (N296, N285, N59, N208);
and AND4 (N297, N287, N125, N165, N7);
and AND4 (N298, N291, N217, N282, N280);
nor NOR3 (N299, N68, N173, N50);
xor XOR2 (N300, N295, N30);
buf BUF1 (N301, N289);
nand NAND2 (N302, N298, N269);
nor NOR4 (N303, N301, N195, N60, N110);
nand NAND2 (N304, N293, N97);
nor NOR4 (N305, N274, N196, N46, N215);
not NOT1 (N306, N297);
xor XOR2 (N307, N299, N134);
buf BUF1 (N308, N303);
buf BUF1 (N309, N302);
and AND3 (N310, N307, N225, N82);
buf BUF1 (N311, N286);
xor XOR2 (N312, N304, N73);
nand NAND2 (N313, N309, N31);
or OR4 (N314, N306, N191, N243, N90);
and AND3 (N315, N308, N35, N158);
nand NAND2 (N316, N313, N246);
nor NOR4 (N317, N315, N44, N180, N152);
xor XOR2 (N318, N300, N270);
nand NAND4 (N319, N317, N298, N262, N315);
buf BUF1 (N320, N294);
or OR2 (N321, N314, N55);
or OR2 (N322, N310, N90);
buf BUF1 (N323, N311);
not NOT1 (N324, N316);
and AND3 (N325, N322, N45, N149);
xor XOR2 (N326, N312, N164);
or OR4 (N327, N321, N259, N137, N304);
xor XOR2 (N328, N319, N172);
xor XOR2 (N329, N323, N303);
xor XOR2 (N330, N324, N112);
and AND2 (N331, N320, N14);
or OR2 (N332, N296, N62);
and AND3 (N333, N328, N178, N122);
or OR3 (N334, N305, N237, N137);
buf BUF1 (N335, N327);
or OR2 (N336, N318, N287);
xor XOR2 (N337, N333, N280);
not NOT1 (N338, N326);
and AND3 (N339, N329, N235, N96);
not NOT1 (N340, N334);
or OR2 (N341, N332, N183);
nor NOR2 (N342, N336, N153);
buf BUF1 (N343, N331);
nor NOR4 (N344, N338, N130, N324, N162);
and AND2 (N345, N335, N248);
not NOT1 (N346, N337);
buf BUF1 (N347, N346);
not NOT1 (N348, N347);
buf BUF1 (N349, N345);
buf BUF1 (N350, N339);
and AND3 (N351, N341, N146, N215);
and AND4 (N352, N350, N309, N174, N326);
and AND2 (N353, N351, N254);
nand NAND4 (N354, N330, N298, N212, N216);
buf BUF1 (N355, N353);
or OR3 (N356, N352, N97, N305);
and AND2 (N357, N344, N247);
buf BUF1 (N358, N325);
buf BUF1 (N359, N356);
nor NOR3 (N360, N349, N87, N102);
xor XOR2 (N361, N357, N332);
xor XOR2 (N362, N340, N340);
nand NAND3 (N363, N361, N60, N192);
not NOT1 (N364, N355);
xor XOR2 (N365, N348, N226);
not NOT1 (N366, N364);
xor XOR2 (N367, N342, N258);
nand NAND4 (N368, N343, N156, N270, N311);
xor XOR2 (N369, N366, N366);
nand NAND4 (N370, N367, N258, N9, N40);
buf BUF1 (N371, N368);
buf BUF1 (N372, N362);
nand NAND3 (N373, N371, N12, N28);
or OR2 (N374, N370, N137);
buf BUF1 (N375, N374);
xor XOR2 (N376, N369, N304);
nand NAND3 (N377, N365, N116, N68);
xor XOR2 (N378, N375, N45);
xor XOR2 (N379, N358, N124);
and AND3 (N380, N376, N82, N180);
and AND4 (N381, N354, N26, N54, N155);
not NOT1 (N382, N360);
not NOT1 (N383, N380);
and AND2 (N384, N383, N51);
not NOT1 (N385, N363);
nor NOR2 (N386, N384, N290);
nor NOR3 (N387, N381, N364, N269);
buf BUF1 (N388, N386);
or OR4 (N389, N388, N286, N56, N357);
nor NOR2 (N390, N387, N131);
not NOT1 (N391, N359);
and AND3 (N392, N378, N330, N334);
nor NOR4 (N393, N373, N212, N244, N162);
xor XOR2 (N394, N391, N8);
not NOT1 (N395, N394);
buf BUF1 (N396, N372);
buf BUF1 (N397, N396);
or OR2 (N398, N385, N234);
buf BUF1 (N399, N392);
buf BUF1 (N400, N398);
buf BUF1 (N401, N395);
buf BUF1 (N402, N390);
nand NAND3 (N403, N397, N124, N53);
xor XOR2 (N404, N402, N227);
and AND4 (N405, N404, N353, N270, N342);
xor XOR2 (N406, N393, N248);
nor NOR3 (N407, N401, N78, N396);
nor NOR4 (N408, N403, N141, N346, N397);
nor NOR3 (N409, N382, N316, N335);
not NOT1 (N410, N406);
xor XOR2 (N411, N377, N232);
buf BUF1 (N412, N409);
nor NOR4 (N413, N412, N322, N216, N191);
xor XOR2 (N414, N405, N98);
not NOT1 (N415, N411);
not NOT1 (N416, N400);
xor XOR2 (N417, N408, N407);
buf BUF1 (N418, N55);
nor NOR3 (N419, N414, N251, N216);
nand NAND2 (N420, N389, N139);
nand NAND2 (N421, N420, N269);
or OR3 (N422, N415, N18, N141);
buf BUF1 (N423, N379);
nand NAND3 (N424, N417, N31, N215);
xor XOR2 (N425, N421, N280);
and AND3 (N426, N399, N102, N394);
xor XOR2 (N427, N426, N186);
nand NAND2 (N428, N424, N98);
and AND2 (N429, N425, N388);
nor NOR4 (N430, N410, N429, N143, N261);
or OR2 (N431, N78, N27);
not NOT1 (N432, N413);
xor XOR2 (N433, N416, N199);
nor NOR2 (N434, N432, N362);
xor XOR2 (N435, N428, N20);
and AND4 (N436, N433, N386, N47, N47);
not NOT1 (N437, N419);
nor NOR2 (N438, N436, N350);
or OR2 (N439, N430, N423);
xor XOR2 (N440, N28, N266);
or OR3 (N441, N437, N119, N140);
nand NAND2 (N442, N440, N258);
nor NOR2 (N443, N418, N372);
buf BUF1 (N444, N443);
nor NOR4 (N445, N438, N424, N136, N26);
and AND2 (N446, N445, N60);
or OR3 (N447, N446, N445, N132);
not NOT1 (N448, N442);
not NOT1 (N449, N441);
nand NAND3 (N450, N431, N13, N150);
nor NOR3 (N451, N439, N349, N382);
and AND2 (N452, N447, N26);
xor XOR2 (N453, N444, N156);
buf BUF1 (N454, N453);
or OR3 (N455, N422, N248, N396);
nand NAND4 (N456, N448, N184, N2, N398);
xor XOR2 (N457, N452, N17);
nor NOR2 (N458, N457, N305);
xor XOR2 (N459, N434, N424);
xor XOR2 (N460, N454, N73);
nand NAND3 (N461, N459, N210, N200);
nor NOR4 (N462, N449, N13, N148, N441);
nand NAND2 (N463, N462, N175);
not NOT1 (N464, N450);
buf BUF1 (N465, N458);
xor XOR2 (N466, N456, N295);
or OR2 (N467, N427, N411);
not NOT1 (N468, N464);
buf BUF1 (N469, N465);
or OR3 (N470, N467, N375, N83);
xor XOR2 (N471, N463, N291);
and AND3 (N472, N469, N341, N425);
and AND2 (N473, N461, N60);
buf BUF1 (N474, N460);
not NOT1 (N475, N473);
nand NAND3 (N476, N470, N252, N299);
and AND4 (N477, N476, N399, N135, N133);
or OR2 (N478, N477, N243);
or OR2 (N479, N468, N119);
xor XOR2 (N480, N478, N339);
and AND3 (N481, N455, N105, N106);
buf BUF1 (N482, N466);
or OR2 (N483, N481, N209);
and AND3 (N484, N472, N28, N344);
or OR3 (N485, N471, N130, N354);
not NOT1 (N486, N479);
buf BUF1 (N487, N485);
xor XOR2 (N488, N475, N397);
nor NOR4 (N489, N487, N108, N228, N333);
or OR2 (N490, N480, N87);
and AND2 (N491, N486, N159);
xor XOR2 (N492, N451, N39);
or OR4 (N493, N489, N469, N94, N139);
buf BUF1 (N494, N484);
buf BUF1 (N495, N435);
nor NOR4 (N496, N488, N246, N272, N86);
xor XOR2 (N497, N474, N394);
and AND4 (N498, N491, N334, N334, N31);
nand NAND4 (N499, N495, N174, N55, N328);
buf BUF1 (N500, N499);
not NOT1 (N501, N498);
xor XOR2 (N502, N497, N413);
nand NAND2 (N503, N502, N40);
nand NAND2 (N504, N501, N293);
or OR3 (N505, N504, N461, N98);
and AND4 (N506, N490, N373, N215, N311);
or OR4 (N507, N503, N321, N288, N421);
buf BUF1 (N508, N483);
nand NAND4 (N509, N505, N314, N157, N86);
nor NOR3 (N510, N482, N168, N326);
nand NAND3 (N511, N494, N120, N154);
not NOT1 (N512, N496);
or OR4 (N513, N506, N84, N84, N113);
nor NOR2 (N514, N511, N79);
xor XOR2 (N515, N493, N267);
and AND2 (N516, N507, N81);
or OR2 (N517, N515, N82);
nand NAND2 (N518, N500, N330);
or OR2 (N519, N508, N470);
and AND4 (N520, N519, N341, N507, N99);
or OR3 (N521, N510, N1, N35);
and AND3 (N522, N512, N373, N473);
not NOT1 (N523, N514);
buf BUF1 (N524, N509);
nor NOR3 (N525, N521, N322, N65);
xor XOR2 (N526, N516, N132);
nor NOR2 (N527, N524, N218);
not NOT1 (N528, N492);
not NOT1 (N529, N518);
not NOT1 (N530, N526);
or OR4 (N531, N527, N288, N133, N335);
or OR2 (N532, N531, N418);
not NOT1 (N533, N517);
buf BUF1 (N534, N533);
or OR3 (N535, N522, N164, N104);
nor NOR4 (N536, N523, N54, N446, N101);
and AND2 (N537, N535, N156);
buf BUF1 (N538, N513);
and AND4 (N539, N520, N34, N290, N288);
and AND4 (N540, N525, N515, N17, N468);
buf BUF1 (N541, N534);
or OR4 (N542, N541, N14, N176, N111);
not NOT1 (N543, N529);
nor NOR4 (N544, N528, N227, N330, N4);
xor XOR2 (N545, N536, N97);
and AND3 (N546, N539, N306, N166);
nand NAND4 (N547, N545, N506, N434, N257);
nor NOR4 (N548, N544, N319, N272, N76);
not NOT1 (N549, N537);
nand NAND4 (N550, N547, N315, N24, N275);
buf BUF1 (N551, N548);
or OR2 (N552, N530, N388);
and AND4 (N553, N538, N150, N40, N351);
or OR3 (N554, N551, N456, N340);
xor XOR2 (N555, N550, N24);
nand NAND4 (N556, N553, N223, N529, N34);
and AND4 (N557, N542, N69, N75, N428);
or OR4 (N558, N546, N64, N141, N50);
xor XOR2 (N559, N543, N38);
xor XOR2 (N560, N552, N279);
and AND3 (N561, N556, N266, N225);
nand NAND2 (N562, N559, N348);
or OR2 (N563, N532, N365);
xor XOR2 (N564, N561, N562);
and AND2 (N565, N337, N391);
and AND3 (N566, N565, N20, N307);
or OR2 (N567, N560, N201);
or OR3 (N568, N557, N379, N134);
or OR4 (N569, N564, N212, N504, N533);
and AND3 (N570, N563, N231, N56);
and AND4 (N571, N567, N107, N190, N191);
nor NOR2 (N572, N566, N423);
buf BUF1 (N573, N540);
and AND4 (N574, N572, N361, N136, N537);
nor NOR2 (N575, N571, N83);
not NOT1 (N576, N568);
and AND2 (N577, N555, N458);
nand NAND4 (N578, N570, N553, N344, N58);
buf BUF1 (N579, N573);
nand NAND2 (N580, N558, N419);
and AND4 (N581, N580, N223, N45, N141);
nor NOR2 (N582, N569, N71);
buf BUF1 (N583, N574);
not NOT1 (N584, N579);
nor NOR2 (N585, N578, N70);
and AND4 (N586, N549, N456, N377, N251);
nand NAND2 (N587, N554, N256);
or OR2 (N588, N581, N485);
or OR4 (N589, N588, N343, N123, N422);
or OR4 (N590, N583, N538, N44, N495);
or OR4 (N591, N585, N421, N281, N471);
and AND2 (N592, N575, N13);
nor NOR4 (N593, N591, N248, N178, N338);
and AND2 (N594, N577, N369);
buf BUF1 (N595, N576);
xor XOR2 (N596, N582, N320);
or OR3 (N597, N584, N567, N139);
xor XOR2 (N598, N597, N285);
and AND3 (N599, N587, N166, N529);
or OR3 (N600, N589, N272, N586);
and AND2 (N601, N358, N312);
nand NAND4 (N602, N593, N128, N273, N101);
nor NOR4 (N603, N598, N250, N489, N499);
buf BUF1 (N604, N592);
nor NOR4 (N605, N590, N5, N406, N15);
or OR3 (N606, N596, N469, N185);
nand NAND4 (N607, N606, N293, N223, N385);
and AND3 (N608, N605, N386, N497);
nor NOR3 (N609, N599, N392, N281);
nor NOR4 (N610, N608, N133, N526, N487);
nand NAND4 (N611, N604, N310, N605, N32);
or OR3 (N612, N602, N555, N320);
nand NAND4 (N613, N595, N563, N86, N581);
xor XOR2 (N614, N600, N454);
nand NAND3 (N615, N609, N73, N128);
xor XOR2 (N616, N610, N294);
or OR2 (N617, N614, N107);
buf BUF1 (N618, N611);
buf BUF1 (N619, N613);
nor NOR2 (N620, N619, N389);
or OR3 (N621, N603, N553, N65);
not NOT1 (N622, N607);
or OR2 (N623, N621, N174);
or OR3 (N624, N617, N282, N615);
not NOT1 (N625, N287);
not NOT1 (N626, N622);
nand NAND2 (N627, N623, N239);
xor XOR2 (N628, N627, N555);
buf BUF1 (N629, N594);
xor XOR2 (N630, N618, N396);
xor XOR2 (N631, N601, N499);
nor NOR2 (N632, N624, N229);
xor XOR2 (N633, N612, N73);
or OR4 (N634, N632, N387, N396, N392);
nand NAND3 (N635, N616, N40, N115);
not NOT1 (N636, N628);
xor XOR2 (N637, N636, N321);
nand NAND4 (N638, N625, N405, N469, N326);
nand NAND4 (N639, N638, N441, N182, N373);
xor XOR2 (N640, N626, N515);
not NOT1 (N641, N635);
nor NOR2 (N642, N637, N555);
nand NAND4 (N643, N639, N401, N291, N404);
buf BUF1 (N644, N640);
xor XOR2 (N645, N634, N488);
and AND2 (N646, N630, N507);
buf BUF1 (N647, N644);
buf BUF1 (N648, N647);
xor XOR2 (N649, N645, N281);
xor XOR2 (N650, N649, N639);
or OR4 (N651, N633, N427, N508, N83);
not NOT1 (N652, N631);
not NOT1 (N653, N620);
nor NOR4 (N654, N652, N104, N470, N526);
and AND4 (N655, N629, N322, N236, N9);
nand NAND3 (N656, N654, N161, N327);
not NOT1 (N657, N656);
nand NAND3 (N658, N657, N561, N210);
and AND2 (N659, N651, N249);
or OR3 (N660, N659, N467, N139);
nor NOR4 (N661, N655, N588, N145, N96);
or OR3 (N662, N653, N73, N208);
or OR2 (N663, N658, N11);
nand NAND3 (N664, N646, N95, N396);
nand NAND4 (N665, N662, N426, N565, N586);
nor NOR4 (N666, N642, N422, N378, N515);
xor XOR2 (N667, N660, N459);
xor XOR2 (N668, N641, N156);
not NOT1 (N669, N668);
and AND3 (N670, N669, N441, N433);
xor XOR2 (N671, N661, N83);
not NOT1 (N672, N671);
nand NAND4 (N673, N665, N412, N205, N604);
or OR3 (N674, N670, N510, N140);
not NOT1 (N675, N650);
or OR4 (N676, N667, N86, N65, N109);
and AND3 (N677, N643, N12, N333);
nand NAND4 (N678, N674, N293, N101, N165);
xor XOR2 (N679, N663, N135);
nor NOR4 (N680, N672, N68, N146, N381);
and AND2 (N681, N664, N9);
xor XOR2 (N682, N679, N63);
not NOT1 (N683, N676);
nor NOR3 (N684, N682, N154, N62);
and AND4 (N685, N677, N172, N269, N500);
nor NOR2 (N686, N673, N128);
xor XOR2 (N687, N648, N416);
nor NOR4 (N688, N666, N122, N258, N313);
and AND2 (N689, N684, N68);
or OR2 (N690, N675, N438);
or OR3 (N691, N690, N359, N138);
nand NAND3 (N692, N691, N526, N283);
nor NOR4 (N693, N689, N337, N45, N539);
not NOT1 (N694, N688);
xor XOR2 (N695, N681, N599);
or OR2 (N696, N687, N682);
and AND3 (N697, N683, N323, N183);
or OR2 (N698, N697, N433);
xor XOR2 (N699, N696, N14);
not NOT1 (N700, N678);
xor XOR2 (N701, N699, N4);
and AND3 (N702, N693, N45, N593);
buf BUF1 (N703, N701);
not NOT1 (N704, N685);
xor XOR2 (N705, N702, N124);
buf BUF1 (N706, N705);
nand NAND3 (N707, N704, N492, N343);
or OR4 (N708, N692, N100, N330, N550);
or OR2 (N709, N703, N691);
xor XOR2 (N710, N707, N49);
or OR3 (N711, N708, N494, N609);
nor NOR2 (N712, N709, N393);
buf BUF1 (N713, N695);
nand NAND3 (N714, N711, N587, N266);
and AND4 (N715, N686, N273, N196, N80);
nand NAND4 (N716, N712, N397, N390, N512);
not NOT1 (N717, N715);
buf BUF1 (N718, N717);
buf BUF1 (N719, N713);
buf BUF1 (N720, N714);
or OR4 (N721, N680, N200, N674, N203);
nor NOR3 (N722, N720, N44, N86);
not NOT1 (N723, N719);
or OR3 (N724, N721, N283, N597);
nand NAND3 (N725, N698, N239, N229);
nand NAND3 (N726, N722, N154, N320);
not NOT1 (N727, N725);
nand NAND3 (N728, N726, N2, N324);
buf BUF1 (N729, N723);
not NOT1 (N730, N716);
and AND2 (N731, N727, N196);
xor XOR2 (N732, N728, N96);
and AND3 (N733, N700, N446, N447);
xor XOR2 (N734, N724, N40);
nor NOR2 (N735, N731, N342);
nand NAND4 (N736, N733, N577, N568, N683);
nor NOR3 (N737, N718, N212, N593);
nor NOR2 (N738, N694, N410);
nand NAND2 (N739, N730, N154);
nor NOR3 (N740, N734, N308, N12);
nand NAND4 (N741, N732, N64, N200, N281);
xor XOR2 (N742, N735, N226);
not NOT1 (N743, N710);
nor NOR2 (N744, N741, N93);
nor NOR2 (N745, N739, N606);
nand NAND2 (N746, N744, N347);
or OR2 (N747, N740, N334);
buf BUF1 (N748, N747);
buf BUF1 (N749, N748);
nor NOR3 (N750, N737, N114, N725);
nand NAND3 (N751, N706, N396, N405);
nor NOR3 (N752, N729, N509, N21);
buf BUF1 (N753, N752);
buf BUF1 (N754, N750);
nand NAND4 (N755, N749, N507, N679, N225);
nor NOR4 (N756, N753, N366, N515, N730);
nor NOR3 (N757, N736, N160, N563);
buf BUF1 (N758, N745);
not NOT1 (N759, N738);
not NOT1 (N760, N751);
nand NAND2 (N761, N757, N666);
not NOT1 (N762, N758);
not NOT1 (N763, N760);
buf BUF1 (N764, N761);
and AND4 (N765, N756, N676, N483, N211);
xor XOR2 (N766, N762, N454);
not NOT1 (N767, N754);
xor XOR2 (N768, N765, N339);
buf BUF1 (N769, N743);
nor NOR3 (N770, N759, N603, N406);
xor XOR2 (N771, N769, N323);
nand NAND2 (N772, N746, N623);
nand NAND4 (N773, N767, N692, N303, N518);
or OR2 (N774, N772, N561);
not NOT1 (N775, N763);
buf BUF1 (N776, N768);
xor XOR2 (N777, N775, N189);
nand NAND3 (N778, N773, N492, N509);
and AND4 (N779, N777, N414, N410, N100);
or OR2 (N780, N776, N166);
nand NAND3 (N781, N742, N489, N182);
or OR3 (N782, N771, N690, N289);
not NOT1 (N783, N755);
or OR3 (N784, N783, N352, N658);
buf BUF1 (N785, N778);
xor XOR2 (N786, N764, N553);
nand NAND4 (N787, N782, N748, N545, N598);
nand NAND4 (N788, N780, N594, N378, N102);
not NOT1 (N789, N784);
xor XOR2 (N790, N789, N476);
and AND2 (N791, N770, N285);
xor XOR2 (N792, N766, N407);
buf BUF1 (N793, N787);
and AND4 (N794, N781, N623, N647, N125);
nor NOR3 (N795, N793, N141, N709);
nand NAND3 (N796, N779, N362, N27);
and AND2 (N797, N796, N103);
not NOT1 (N798, N786);
nand NAND4 (N799, N788, N574, N660, N672);
or OR2 (N800, N785, N604);
nand NAND3 (N801, N797, N263, N220);
not NOT1 (N802, N774);
not NOT1 (N803, N800);
or OR2 (N804, N794, N372);
nor NOR2 (N805, N802, N675);
nand NAND2 (N806, N803, N491);
buf BUF1 (N807, N795);
not NOT1 (N808, N791);
or OR4 (N809, N808, N409, N319, N484);
buf BUF1 (N810, N792);
buf BUF1 (N811, N810);
and AND4 (N812, N806, N679, N173, N114);
not NOT1 (N813, N809);
and AND4 (N814, N805, N211, N654, N61);
xor XOR2 (N815, N801, N130);
not NOT1 (N816, N815);
or OR2 (N817, N807, N583);
or OR3 (N818, N814, N38, N651);
nand NAND4 (N819, N798, N116, N572, N163);
not NOT1 (N820, N812);
not NOT1 (N821, N819);
or OR2 (N822, N821, N34);
and AND2 (N823, N804, N597);
and AND4 (N824, N813, N707, N33, N338);
xor XOR2 (N825, N822, N371);
xor XOR2 (N826, N816, N357);
or OR3 (N827, N825, N594, N192);
and AND4 (N828, N818, N128, N27, N655);
not NOT1 (N829, N811);
xor XOR2 (N830, N820, N599);
or OR2 (N831, N827, N209);
nor NOR4 (N832, N824, N522, N183, N602);
nand NAND4 (N833, N829, N290, N21, N357);
or OR4 (N834, N830, N316, N812, N730);
nand NAND3 (N835, N817, N694, N443);
buf BUF1 (N836, N834);
buf BUF1 (N837, N836);
buf BUF1 (N838, N835);
buf BUF1 (N839, N823);
or OR4 (N840, N837, N34, N288, N420);
or OR3 (N841, N833, N554, N202);
and AND2 (N842, N838, N360);
buf BUF1 (N843, N828);
or OR4 (N844, N839, N703, N695, N33);
buf BUF1 (N845, N840);
and AND4 (N846, N844, N633, N60, N789);
nor NOR2 (N847, N845, N177);
nand NAND2 (N848, N847, N475);
buf BUF1 (N849, N848);
or OR2 (N850, N790, N112);
nand NAND4 (N851, N831, N810, N31, N94);
nor NOR2 (N852, N843, N403);
buf BUF1 (N853, N799);
nor NOR3 (N854, N832, N819, N792);
and AND2 (N855, N841, N687);
buf BUF1 (N856, N852);
buf BUF1 (N857, N855);
nor NOR4 (N858, N850, N724, N308, N371);
or OR3 (N859, N846, N684, N675);
buf BUF1 (N860, N854);
buf BUF1 (N861, N851);
not NOT1 (N862, N853);
nor NOR4 (N863, N857, N497, N538, N524);
or OR2 (N864, N842, N402);
nand NAND3 (N865, N860, N776, N735);
buf BUF1 (N866, N862);
xor XOR2 (N867, N866, N429);
xor XOR2 (N868, N856, N618);
xor XOR2 (N869, N863, N57);
nor NOR4 (N870, N864, N804, N359, N718);
not NOT1 (N871, N859);
buf BUF1 (N872, N868);
and AND4 (N873, N861, N643, N304, N750);
buf BUF1 (N874, N858);
nand NAND3 (N875, N869, N568, N265);
or OR3 (N876, N873, N274, N575);
or OR4 (N877, N872, N864, N712, N603);
xor XOR2 (N878, N871, N326);
nand NAND2 (N879, N849, N206);
xor XOR2 (N880, N877, N870);
not NOT1 (N881, N532);
nor NOR4 (N882, N879, N596, N502, N594);
or OR2 (N883, N875, N700);
and AND3 (N884, N881, N317, N366);
or OR4 (N885, N878, N717, N283, N125);
xor XOR2 (N886, N883, N515);
nand NAND4 (N887, N884, N93, N369, N171);
or OR2 (N888, N826, N738);
xor XOR2 (N889, N865, N188);
not NOT1 (N890, N867);
or OR4 (N891, N890, N837, N565, N374);
buf BUF1 (N892, N876);
and AND3 (N893, N886, N543, N851);
xor XOR2 (N894, N887, N822);
or OR3 (N895, N885, N705, N74);
nand NAND3 (N896, N895, N618, N350);
buf BUF1 (N897, N896);
buf BUF1 (N898, N880);
and AND2 (N899, N888, N659);
nand NAND2 (N900, N898, N293);
xor XOR2 (N901, N893, N178);
not NOT1 (N902, N900);
xor XOR2 (N903, N874, N544);
buf BUF1 (N904, N889);
nand NAND3 (N905, N882, N492, N769);
nor NOR4 (N906, N905, N859, N311, N331);
buf BUF1 (N907, N902);
and AND3 (N908, N897, N777, N70);
nand NAND4 (N909, N906, N686, N868, N495);
buf BUF1 (N910, N904);
buf BUF1 (N911, N903);
xor XOR2 (N912, N910, N857);
nand NAND2 (N913, N907, N226);
and AND3 (N914, N913, N208, N214);
not NOT1 (N915, N891);
and AND2 (N916, N915, N907);
not NOT1 (N917, N909);
not NOT1 (N918, N916);
xor XOR2 (N919, N917, N52);
buf BUF1 (N920, N892);
nand NAND4 (N921, N911, N184, N742, N328);
nand NAND2 (N922, N899, N800);
nor NOR3 (N923, N921, N431, N785);
nor NOR4 (N924, N918, N413, N510, N749);
not NOT1 (N925, N901);
not NOT1 (N926, N922);
or OR3 (N927, N926, N676, N714);
or OR4 (N928, N924, N73, N293, N688);
and AND4 (N929, N919, N246, N211, N167);
nor NOR2 (N930, N908, N489);
not NOT1 (N931, N894);
nor NOR4 (N932, N931, N836, N372, N850);
or OR2 (N933, N914, N191);
nand NAND3 (N934, N920, N857, N571);
buf BUF1 (N935, N927);
or OR3 (N936, N912, N582, N166);
xor XOR2 (N937, N929, N932);
nand NAND3 (N938, N399, N866, N361);
or OR3 (N939, N923, N864, N724);
or OR4 (N940, N933, N923, N481, N260);
xor XOR2 (N941, N934, N421);
xor XOR2 (N942, N939, N714);
nand NAND4 (N943, N935, N309, N26, N241);
or OR3 (N944, N938, N637, N851);
buf BUF1 (N945, N943);
xor XOR2 (N946, N925, N292);
nor NOR4 (N947, N937, N902, N938, N421);
or OR3 (N948, N942, N885, N712);
xor XOR2 (N949, N946, N825);
xor XOR2 (N950, N944, N268);
or OR4 (N951, N948, N619, N776, N546);
or OR3 (N952, N951, N743, N769);
nor NOR4 (N953, N952, N568, N510, N415);
buf BUF1 (N954, N941);
and AND2 (N955, N940, N297);
xor XOR2 (N956, N928, N899);
and AND3 (N957, N956, N935, N766);
nand NAND4 (N958, N930, N784, N413, N858);
xor XOR2 (N959, N945, N674);
and AND2 (N960, N947, N820);
not NOT1 (N961, N958);
nand NAND3 (N962, N960, N931, N940);
not NOT1 (N963, N953);
buf BUF1 (N964, N962);
or OR3 (N965, N957, N53, N775);
and AND3 (N966, N963, N704, N136);
nand NAND3 (N967, N955, N815, N175);
and AND3 (N968, N936, N271, N670);
or OR2 (N969, N968, N20);
not NOT1 (N970, N964);
not NOT1 (N971, N966);
not NOT1 (N972, N949);
not NOT1 (N973, N959);
not NOT1 (N974, N970);
not NOT1 (N975, N972);
nand NAND3 (N976, N954, N349, N432);
not NOT1 (N977, N971);
or OR2 (N978, N950, N579);
and AND3 (N979, N975, N18, N975);
buf BUF1 (N980, N969);
and AND4 (N981, N967, N369, N301, N83);
buf BUF1 (N982, N976);
not NOT1 (N983, N965);
and AND2 (N984, N973, N425);
or OR4 (N985, N961, N876, N155, N67);
not NOT1 (N986, N983);
or OR4 (N987, N984, N477, N671, N246);
buf BUF1 (N988, N979);
buf BUF1 (N989, N987);
or OR2 (N990, N974, N421);
buf BUF1 (N991, N985);
not NOT1 (N992, N991);
or OR3 (N993, N989, N944, N90);
nand NAND3 (N994, N988, N330, N941);
nand NAND2 (N995, N980, N897);
or OR4 (N996, N994, N677, N903, N858);
buf BUF1 (N997, N982);
xor XOR2 (N998, N981, N947);
buf BUF1 (N999, N992);
and AND3 (N1000, N999, N967, N580);
and AND2 (N1001, N990, N545);
and AND2 (N1002, N977, N572);
nand NAND3 (N1003, N1001, N775, N186);
not NOT1 (N1004, N978);
buf BUF1 (N1005, N1004);
nor NOR4 (N1006, N1003, N155, N192, N809);
nand NAND3 (N1007, N986, N657, N229);
nor NOR2 (N1008, N1005, N299);
nor NOR3 (N1009, N1008, N957, N240);
nand NAND3 (N1010, N1006, N417, N998);
and AND2 (N1011, N641, N839);
buf BUF1 (N1012, N997);
or OR2 (N1013, N1011, N89);
or OR3 (N1014, N1007, N589, N287);
xor XOR2 (N1015, N996, N595);
buf BUF1 (N1016, N1013);
or OR4 (N1017, N1000, N144, N949, N513);
or OR4 (N1018, N993, N532, N817, N352);
buf BUF1 (N1019, N1017);
xor XOR2 (N1020, N1016, N856);
nor NOR2 (N1021, N1015, N686);
nor NOR4 (N1022, N1012, N841, N785, N224);
and AND3 (N1023, N1018, N738, N708);
buf BUF1 (N1024, N1021);
nand NAND3 (N1025, N1022, N812, N443);
buf BUF1 (N1026, N1009);
buf BUF1 (N1027, N1025);
nand NAND2 (N1028, N1020, N367);
not NOT1 (N1029, N1027);
nand NAND3 (N1030, N1028, N5, N943);
xor XOR2 (N1031, N1030, N434);
and AND4 (N1032, N1031, N530, N289, N449);
nand NAND4 (N1033, N1014, N973, N448, N144);
and AND2 (N1034, N1023, N298);
xor XOR2 (N1035, N1002, N961);
nand NAND2 (N1036, N1026, N708);
xor XOR2 (N1037, N1033, N455);
nor NOR3 (N1038, N1019, N615, N868);
buf BUF1 (N1039, N1029);
nand NAND4 (N1040, N995, N690, N676, N30);
xor XOR2 (N1041, N1035, N738);
xor XOR2 (N1042, N1038, N235);
buf BUF1 (N1043, N1041);
not NOT1 (N1044, N1039);
xor XOR2 (N1045, N1044, N597);
nor NOR4 (N1046, N1037, N9, N864, N931);
nand NAND2 (N1047, N1034, N204);
buf BUF1 (N1048, N1024);
and AND4 (N1049, N1036, N266, N396, N952);
not NOT1 (N1050, N1049);
nand NAND3 (N1051, N1045, N38, N395);
nor NOR3 (N1052, N1040, N588, N199);
buf BUF1 (N1053, N1046);
not NOT1 (N1054, N1010);
nor NOR3 (N1055, N1051, N468, N291);
nand NAND2 (N1056, N1054, N942);
nor NOR4 (N1057, N1042, N721, N699, N271);
and AND2 (N1058, N1056, N238);
buf BUF1 (N1059, N1057);
xor XOR2 (N1060, N1048, N35);
xor XOR2 (N1061, N1059, N445);
xor XOR2 (N1062, N1053, N987);
nand NAND3 (N1063, N1032, N6, N682);
nand NAND4 (N1064, N1052, N319, N163, N1013);
xor XOR2 (N1065, N1063, N32);
or OR3 (N1066, N1065, N776, N600);
nand NAND4 (N1067, N1064, N359, N93, N147);
and AND2 (N1068, N1047, N239);
and AND3 (N1069, N1058, N78, N382);
and AND2 (N1070, N1066, N506);
xor XOR2 (N1071, N1061, N848);
and AND4 (N1072, N1050, N365, N60, N242);
nand NAND4 (N1073, N1043, N945, N132, N565);
nor NOR2 (N1074, N1073, N382);
or OR4 (N1075, N1070, N75, N281, N152);
xor XOR2 (N1076, N1055, N303);
and AND4 (N1077, N1062, N42, N465, N1053);
and AND3 (N1078, N1071, N824, N1065);
or OR4 (N1079, N1074, N632, N738, N574);
and AND3 (N1080, N1078, N1053, N159);
buf BUF1 (N1081, N1075);
or OR4 (N1082, N1072, N301, N125, N1069);
xor XOR2 (N1083, N835, N578);
nor NOR2 (N1084, N1082, N80);
xor XOR2 (N1085, N1079, N31);
and AND2 (N1086, N1067, N298);
or OR3 (N1087, N1083, N977, N51);
buf BUF1 (N1088, N1084);
xor XOR2 (N1089, N1076, N279);
xor XOR2 (N1090, N1080, N145);
and AND2 (N1091, N1090, N767);
buf BUF1 (N1092, N1086);
buf BUF1 (N1093, N1089);
or OR2 (N1094, N1060, N999);
buf BUF1 (N1095, N1081);
xor XOR2 (N1096, N1095, N230);
xor XOR2 (N1097, N1087, N954);
or OR3 (N1098, N1068, N677, N75);
or OR4 (N1099, N1096, N294, N561, N1009);
and AND4 (N1100, N1092, N263, N171, N407);
nor NOR4 (N1101, N1098, N1053, N250, N620);
or OR3 (N1102, N1091, N478, N705);
buf BUF1 (N1103, N1094);
xor XOR2 (N1104, N1103, N18);
buf BUF1 (N1105, N1097);
xor XOR2 (N1106, N1085, N739);
xor XOR2 (N1107, N1088, N1060);
nor NOR2 (N1108, N1077, N332);
and AND3 (N1109, N1107, N322, N847);
not NOT1 (N1110, N1106);
nand NAND4 (N1111, N1110, N66, N125, N475);
nor NOR4 (N1112, N1102, N973, N192, N516);
or OR3 (N1113, N1100, N1047, N365);
or OR2 (N1114, N1099, N237);
or OR3 (N1115, N1101, N910, N166);
xor XOR2 (N1116, N1115, N194);
not NOT1 (N1117, N1113);
not NOT1 (N1118, N1105);
nand NAND4 (N1119, N1093, N752, N384, N966);
not NOT1 (N1120, N1114);
or OR2 (N1121, N1109, N690);
not NOT1 (N1122, N1111);
and AND3 (N1123, N1122, N420, N998);
or OR2 (N1124, N1117, N1014);
nor NOR2 (N1125, N1112, N409);
buf BUF1 (N1126, N1118);
or OR2 (N1127, N1124, N311);
nand NAND3 (N1128, N1125, N278, N1001);
nand NAND3 (N1129, N1121, N383, N272);
or OR4 (N1130, N1129, N571, N1011, N527);
not NOT1 (N1131, N1130);
buf BUF1 (N1132, N1131);
buf BUF1 (N1133, N1116);
buf BUF1 (N1134, N1126);
not NOT1 (N1135, N1120);
nand NAND2 (N1136, N1134, N412);
or OR3 (N1137, N1119, N1047, N853);
and AND4 (N1138, N1133, N897, N15, N204);
not NOT1 (N1139, N1135);
buf BUF1 (N1140, N1138);
xor XOR2 (N1141, N1123, N215);
xor XOR2 (N1142, N1104, N508);
nand NAND4 (N1143, N1136, N854, N318, N1027);
or OR3 (N1144, N1108, N597, N471);
not NOT1 (N1145, N1127);
not NOT1 (N1146, N1137);
not NOT1 (N1147, N1140);
nor NOR2 (N1148, N1146, N1098);
and AND3 (N1149, N1147, N202, N883);
not NOT1 (N1150, N1143);
not NOT1 (N1151, N1144);
buf BUF1 (N1152, N1141);
buf BUF1 (N1153, N1149);
nand NAND4 (N1154, N1150, N412, N81, N18);
xor XOR2 (N1155, N1152, N1107);
or OR3 (N1156, N1153, N445, N211);
nand NAND3 (N1157, N1151, N812, N401);
nor NOR4 (N1158, N1148, N679, N814, N838);
not NOT1 (N1159, N1157);
or OR2 (N1160, N1158, N640);
or OR4 (N1161, N1145, N962, N870, N282);
xor XOR2 (N1162, N1155, N64);
and AND4 (N1163, N1128, N675, N326, N1137);
nor NOR4 (N1164, N1139, N974, N276, N82);
nor NOR4 (N1165, N1161, N468, N510, N361);
not NOT1 (N1166, N1154);
xor XOR2 (N1167, N1163, N1165);
nand NAND4 (N1168, N1026, N109, N503, N80);
not NOT1 (N1169, N1132);
not NOT1 (N1170, N1166);
xor XOR2 (N1171, N1170, N470);
nor NOR4 (N1172, N1171, N1098, N1032, N1111);
not NOT1 (N1173, N1156);
not NOT1 (N1174, N1159);
nand NAND4 (N1175, N1173, N1008, N976, N1076);
buf BUF1 (N1176, N1172);
buf BUF1 (N1177, N1162);
xor XOR2 (N1178, N1167, N276);
nand NAND4 (N1179, N1175, N741, N366, N688);
xor XOR2 (N1180, N1179, N875);
buf BUF1 (N1181, N1174);
nor NOR3 (N1182, N1160, N456, N729);
not NOT1 (N1183, N1182);
or OR2 (N1184, N1164, N590);
nor NOR4 (N1185, N1168, N296, N344, N598);
not NOT1 (N1186, N1176);
and AND2 (N1187, N1183, N119);
buf BUF1 (N1188, N1177);
buf BUF1 (N1189, N1184);
nand NAND2 (N1190, N1178, N336);
or OR3 (N1191, N1142, N803, N843);
not NOT1 (N1192, N1189);
or OR3 (N1193, N1185, N218, N837);
nor NOR2 (N1194, N1187, N902);
or OR3 (N1195, N1193, N1131, N915);
or OR2 (N1196, N1169, N487);
or OR2 (N1197, N1181, N1037);
xor XOR2 (N1198, N1195, N918);
nand NAND2 (N1199, N1194, N658);
xor XOR2 (N1200, N1196, N788);
and AND3 (N1201, N1200, N504, N394);
not NOT1 (N1202, N1191);
xor XOR2 (N1203, N1192, N741);
buf BUF1 (N1204, N1201);
xor XOR2 (N1205, N1188, N542);
buf BUF1 (N1206, N1180);
or OR4 (N1207, N1197, N338, N681, N900);
nor NOR3 (N1208, N1207, N544, N852);
buf BUF1 (N1209, N1199);
or OR2 (N1210, N1190, N560);
xor XOR2 (N1211, N1205, N328);
and AND3 (N1212, N1202, N331, N923);
buf BUF1 (N1213, N1186);
and AND2 (N1214, N1213, N170);
and AND4 (N1215, N1210, N1106, N652, N923);
or OR2 (N1216, N1204, N622);
nor NOR3 (N1217, N1212, N1058, N245);
or OR4 (N1218, N1206, N1080, N933, N1116);
buf BUF1 (N1219, N1198);
buf BUF1 (N1220, N1215);
not NOT1 (N1221, N1203);
or OR4 (N1222, N1217, N674, N404, N449);
nor NOR2 (N1223, N1209, N437);
not NOT1 (N1224, N1208);
or OR2 (N1225, N1223, N804);
not NOT1 (N1226, N1222);
buf BUF1 (N1227, N1214);
and AND2 (N1228, N1216, N1007);
nand NAND4 (N1229, N1211, N360, N69, N434);
nand NAND3 (N1230, N1229, N17, N578);
buf BUF1 (N1231, N1230);
and AND2 (N1232, N1224, N515);
not NOT1 (N1233, N1219);
nor NOR4 (N1234, N1221, N208, N844, N572);
buf BUF1 (N1235, N1218);
buf BUF1 (N1236, N1220);
buf BUF1 (N1237, N1228);
and AND4 (N1238, N1232, N432, N479, N824);
nand NAND3 (N1239, N1233, N689, N515);
nor NOR4 (N1240, N1226, N188, N48, N587);
buf BUF1 (N1241, N1240);
nand NAND2 (N1242, N1227, N291);
and AND2 (N1243, N1236, N25);
and AND3 (N1244, N1231, N25, N609);
not NOT1 (N1245, N1239);
not NOT1 (N1246, N1242);
and AND3 (N1247, N1244, N34, N832);
nand NAND4 (N1248, N1225, N1117, N490, N1207);
xor XOR2 (N1249, N1241, N267);
xor XOR2 (N1250, N1238, N1188);
buf BUF1 (N1251, N1234);
not NOT1 (N1252, N1250);
or OR3 (N1253, N1251, N455, N431);
or OR2 (N1254, N1235, N329);
not NOT1 (N1255, N1245);
nor NOR4 (N1256, N1246, N630, N1093, N441);
nor NOR4 (N1257, N1252, N216, N356, N461);
nand NAND2 (N1258, N1257, N54);
not NOT1 (N1259, N1237);
nand NAND2 (N1260, N1243, N795);
not NOT1 (N1261, N1260);
buf BUF1 (N1262, N1261);
nand NAND2 (N1263, N1247, N508);
xor XOR2 (N1264, N1255, N660);
xor XOR2 (N1265, N1259, N406);
xor XOR2 (N1266, N1263, N159);
xor XOR2 (N1267, N1256, N855);
xor XOR2 (N1268, N1264, N296);
or OR2 (N1269, N1248, N1204);
and AND3 (N1270, N1254, N424, N980);
buf BUF1 (N1271, N1265);
nor NOR3 (N1272, N1269, N1043, N1054);
and AND4 (N1273, N1272, N458, N211, N493);
xor XOR2 (N1274, N1253, N1124);
or OR3 (N1275, N1273, N1082, N331);
nor NOR3 (N1276, N1258, N139, N1137);
buf BUF1 (N1277, N1262);
and AND3 (N1278, N1267, N539, N722);
xor XOR2 (N1279, N1266, N1076);
nand NAND3 (N1280, N1277, N126, N317);
nor NOR2 (N1281, N1275, N171);
buf BUF1 (N1282, N1278);
buf BUF1 (N1283, N1271);
not NOT1 (N1284, N1279);
nor NOR3 (N1285, N1281, N945, N905);
buf BUF1 (N1286, N1268);
or OR3 (N1287, N1284, N844, N1057);
nand NAND2 (N1288, N1283, N1257);
nand NAND3 (N1289, N1249, N411, N468);
buf BUF1 (N1290, N1274);
not NOT1 (N1291, N1276);
or OR2 (N1292, N1286, N553);
and AND2 (N1293, N1292, N63);
buf BUF1 (N1294, N1291);
or OR3 (N1295, N1280, N113, N896);
or OR4 (N1296, N1293, N168, N1154, N18);
xor XOR2 (N1297, N1282, N619);
or OR3 (N1298, N1294, N56, N1193);
xor XOR2 (N1299, N1270, N871);
nand NAND2 (N1300, N1288, N333);
nor NOR3 (N1301, N1287, N1047, N1273);
or OR2 (N1302, N1295, N697);
xor XOR2 (N1303, N1296, N468);
not NOT1 (N1304, N1290);
nor NOR2 (N1305, N1300, N305);
xor XOR2 (N1306, N1305, N382);
xor XOR2 (N1307, N1298, N748);
and AND4 (N1308, N1297, N57, N969, N542);
or OR4 (N1309, N1289, N539, N411, N1037);
buf BUF1 (N1310, N1307);
not NOT1 (N1311, N1285);
nor NOR4 (N1312, N1302, N1155, N1031, N41);
nand NAND4 (N1313, N1311, N653, N1191, N592);
not NOT1 (N1314, N1313);
buf BUF1 (N1315, N1303);
xor XOR2 (N1316, N1306, N306);
nand NAND2 (N1317, N1308, N140);
or OR2 (N1318, N1304, N60);
not NOT1 (N1319, N1314);
nand NAND4 (N1320, N1312, N963, N1204, N1313);
nor NOR4 (N1321, N1319, N31, N1057, N913);
nor NOR2 (N1322, N1321, N212);
and AND4 (N1323, N1315, N16, N367, N1158);
xor XOR2 (N1324, N1309, N151);
and AND2 (N1325, N1323, N158);
not NOT1 (N1326, N1301);
buf BUF1 (N1327, N1320);
nor NOR3 (N1328, N1316, N1034, N629);
xor XOR2 (N1329, N1325, N515);
not NOT1 (N1330, N1326);
not NOT1 (N1331, N1317);
nand NAND2 (N1332, N1318, N870);
nand NAND2 (N1333, N1332, N1048);
nor NOR3 (N1334, N1327, N762, N518);
nor NOR2 (N1335, N1330, N942);
xor XOR2 (N1336, N1334, N368);
nor NOR3 (N1337, N1331, N717, N554);
or OR2 (N1338, N1335, N363);
and AND2 (N1339, N1336, N1063);
buf BUF1 (N1340, N1338);
nand NAND2 (N1341, N1328, N19);
buf BUF1 (N1342, N1310);
xor XOR2 (N1343, N1322, N1154);
buf BUF1 (N1344, N1333);
xor XOR2 (N1345, N1342, N547);
or OR4 (N1346, N1343, N589, N55, N524);
not NOT1 (N1347, N1344);
nand NAND2 (N1348, N1337, N1027);
not NOT1 (N1349, N1324);
or OR4 (N1350, N1349, N396, N859, N703);
buf BUF1 (N1351, N1341);
nor NOR3 (N1352, N1340, N899, N1082);
and AND2 (N1353, N1347, N58);
nor NOR3 (N1354, N1329, N750, N1299);
or OR2 (N1355, N545, N825);
nor NOR3 (N1356, N1355, N1246, N66);
nand NAND4 (N1357, N1354, N461, N624, N1119);
buf BUF1 (N1358, N1356);
xor XOR2 (N1359, N1345, N1213);
nor NOR4 (N1360, N1339, N864, N209, N1159);
nand NAND3 (N1361, N1348, N1135, N629);
and AND4 (N1362, N1346, N203, N838, N236);
buf BUF1 (N1363, N1359);
and AND4 (N1364, N1363, N92, N1098, N1033);
xor XOR2 (N1365, N1353, N35);
or OR4 (N1366, N1358, N255, N1097, N531);
nor NOR2 (N1367, N1352, N1190);
or OR3 (N1368, N1361, N696, N867);
nand NAND4 (N1369, N1362, N452, N1116, N1078);
nor NOR2 (N1370, N1350, N732);
buf BUF1 (N1371, N1357);
xor XOR2 (N1372, N1367, N639);
nor NOR4 (N1373, N1370, N1243, N1346, N223);
and AND4 (N1374, N1371, N1223, N842, N793);
xor XOR2 (N1375, N1368, N630);
and AND3 (N1376, N1372, N439, N613);
and AND2 (N1377, N1369, N626);
nor NOR4 (N1378, N1376, N323, N1059, N197);
or OR3 (N1379, N1373, N245, N209);
and AND2 (N1380, N1364, N1143);
xor XOR2 (N1381, N1351, N1046);
or OR4 (N1382, N1365, N274, N1375, N326);
not NOT1 (N1383, N507);
or OR2 (N1384, N1366, N476);
xor XOR2 (N1385, N1381, N574);
nor NOR4 (N1386, N1382, N1242, N927, N1196);
buf BUF1 (N1387, N1379);
and AND3 (N1388, N1385, N923, N1204);
or OR4 (N1389, N1374, N291, N1338, N1290);
nor NOR2 (N1390, N1384, N1008);
or OR4 (N1391, N1387, N357, N783, N199);
xor XOR2 (N1392, N1386, N1276);
nor NOR4 (N1393, N1390, N615, N400, N957);
buf BUF1 (N1394, N1391);
and AND4 (N1395, N1392, N355, N92, N1271);
and AND2 (N1396, N1393, N752);
nand NAND4 (N1397, N1377, N1168, N808, N375);
not NOT1 (N1398, N1394);
or OR3 (N1399, N1389, N232, N136);
or OR2 (N1400, N1380, N433);
not NOT1 (N1401, N1399);
nor NOR4 (N1402, N1383, N320, N609, N587);
not NOT1 (N1403, N1395);
and AND4 (N1404, N1397, N1240, N503, N946);
not NOT1 (N1405, N1396);
xor XOR2 (N1406, N1403, N1358);
xor XOR2 (N1407, N1405, N298);
or OR3 (N1408, N1360, N661, N191);
not NOT1 (N1409, N1408);
buf BUF1 (N1410, N1407);
nand NAND4 (N1411, N1401, N387, N738, N954);
or OR4 (N1412, N1409, N735, N1386, N196);
buf BUF1 (N1413, N1412);
or OR4 (N1414, N1411, N1348, N1162, N509);
and AND2 (N1415, N1398, N1386);
or OR4 (N1416, N1378, N357, N325, N326);
nor NOR3 (N1417, N1410, N302, N970);
buf BUF1 (N1418, N1406);
not NOT1 (N1419, N1416);
buf BUF1 (N1420, N1419);
nand NAND4 (N1421, N1415, N211, N393, N720);
nor NOR3 (N1422, N1421, N222, N439);
and AND2 (N1423, N1388, N756);
nand NAND4 (N1424, N1414, N963, N411, N793);
nor NOR4 (N1425, N1422, N1303, N1279, N125);
xor XOR2 (N1426, N1420, N1011);
or OR3 (N1427, N1402, N137, N1064);
not NOT1 (N1428, N1418);
nand NAND4 (N1429, N1404, N303, N1329, N885);
or OR3 (N1430, N1413, N1054, N233);
or OR2 (N1431, N1429, N137);
not NOT1 (N1432, N1431);
not NOT1 (N1433, N1427);
and AND3 (N1434, N1432, N196, N362);
and AND3 (N1435, N1434, N1398, N470);
xor XOR2 (N1436, N1426, N212);
and AND3 (N1437, N1425, N881, N404);
and AND2 (N1438, N1437, N226);
xor XOR2 (N1439, N1428, N523);
nand NAND3 (N1440, N1435, N20, N619);
buf BUF1 (N1441, N1417);
buf BUF1 (N1442, N1439);
nand NAND2 (N1443, N1440, N509);
or OR4 (N1444, N1441, N323, N1219, N412);
nor NOR4 (N1445, N1433, N892, N28, N649);
or OR3 (N1446, N1443, N1311, N885);
nor NOR4 (N1447, N1436, N663, N188, N667);
nor NOR4 (N1448, N1430, N869, N442, N197);
xor XOR2 (N1449, N1400, N108);
and AND3 (N1450, N1445, N1312, N981);
not NOT1 (N1451, N1438);
nand NAND3 (N1452, N1448, N1356, N493);
or OR2 (N1453, N1442, N819);
not NOT1 (N1454, N1452);
xor XOR2 (N1455, N1450, N1235);
nor NOR2 (N1456, N1446, N947);
or OR2 (N1457, N1447, N1229);
and AND2 (N1458, N1457, N282);
or OR4 (N1459, N1444, N267, N1002, N563);
buf BUF1 (N1460, N1455);
nor NOR2 (N1461, N1453, N764);
and AND2 (N1462, N1456, N736);
xor XOR2 (N1463, N1454, N832);
buf BUF1 (N1464, N1463);
not NOT1 (N1465, N1460);
nor NOR3 (N1466, N1462, N942, N658);
nor NOR2 (N1467, N1459, N1318);
buf BUF1 (N1468, N1466);
or OR3 (N1469, N1451, N166, N1011);
nand NAND3 (N1470, N1465, N123, N1139);
nand NAND3 (N1471, N1470, N1299, N1005);
or OR4 (N1472, N1424, N51, N1128, N363);
nand NAND2 (N1473, N1467, N762);
xor XOR2 (N1474, N1468, N236);
or OR4 (N1475, N1472, N786, N1150, N64);
and AND3 (N1476, N1469, N293, N1372);
not NOT1 (N1477, N1461);
xor XOR2 (N1478, N1464, N269);
not NOT1 (N1479, N1471);
not NOT1 (N1480, N1476);
and AND3 (N1481, N1473, N964, N283);
or OR4 (N1482, N1478, N196, N419, N668);
buf BUF1 (N1483, N1481);
or OR4 (N1484, N1449, N686, N47, N473);
nand NAND2 (N1485, N1480, N805);
xor XOR2 (N1486, N1475, N394);
or OR2 (N1487, N1485, N603);
xor XOR2 (N1488, N1484, N1106);
nor NOR3 (N1489, N1477, N77, N395);
and AND4 (N1490, N1482, N828, N934, N55);
nand NAND3 (N1491, N1486, N228, N104);
not NOT1 (N1492, N1474);
or OR3 (N1493, N1489, N501, N476);
xor XOR2 (N1494, N1423, N245);
or OR4 (N1495, N1494, N601, N69, N1180);
nor NOR4 (N1496, N1488, N498, N345, N1336);
or OR2 (N1497, N1492, N18);
buf BUF1 (N1498, N1496);
or OR3 (N1499, N1458, N928, N1433);
buf BUF1 (N1500, N1493);
buf BUF1 (N1501, N1483);
xor XOR2 (N1502, N1490, N210);
xor XOR2 (N1503, N1499, N651);
nand NAND3 (N1504, N1500, N519, N1110);
nor NOR4 (N1505, N1487, N912, N1472, N1242);
or OR3 (N1506, N1498, N744, N231);
not NOT1 (N1507, N1479);
and AND3 (N1508, N1507, N423, N1346);
nor NOR4 (N1509, N1503, N994, N249, N29);
nor NOR3 (N1510, N1504, N522, N814);
nand NAND2 (N1511, N1501, N1464);
nor NOR3 (N1512, N1502, N344, N347);
xor XOR2 (N1513, N1512, N1368);
nand NAND3 (N1514, N1513, N970, N776);
not NOT1 (N1515, N1505);
nand NAND4 (N1516, N1510, N1234, N342, N1370);
not NOT1 (N1517, N1495);
not NOT1 (N1518, N1514);
and AND2 (N1519, N1508, N549);
not NOT1 (N1520, N1519);
buf BUF1 (N1521, N1516);
and AND4 (N1522, N1497, N1467, N1395, N977);
buf BUF1 (N1523, N1515);
buf BUF1 (N1524, N1517);
nand NAND4 (N1525, N1520, N479, N765, N1113);
or OR4 (N1526, N1524, N761, N1408, N1139);
nand NAND2 (N1527, N1518, N871);
nor NOR2 (N1528, N1511, N25);
xor XOR2 (N1529, N1523, N674);
buf BUF1 (N1530, N1522);
nand NAND4 (N1531, N1509, N725, N335, N620);
nand NAND4 (N1532, N1529, N861, N441, N701);
not NOT1 (N1533, N1528);
nand NAND2 (N1534, N1521, N923);
not NOT1 (N1535, N1506);
and AND4 (N1536, N1534, N662, N1422, N1190);
xor XOR2 (N1537, N1536, N336);
or OR4 (N1538, N1535, N399, N398, N1380);
and AND3 (N1539, N1537, N1302, N659);
or OR4 (N1540, N1539, N1404, N144, N1079);
nor NOR2 (N1541, N1533, N496);
or OR4 (N1542, N1541, N1026, N1174, N1251);
and AND4 (N1543, N1525, N732, N252, N18);
and AND3 (N1544, N1532, N142, N64);
not NOT1 (N1545, N1527);
and AND2 (N1546, N1540, N773);
buf BUF1 (N1547, N1545);
not NOT1 (N1548, N1546);
and AND4 (N1549, N1531, N838, N79, N1406);
or OR4 (N1550, N1544, N1136, N1277, N23);
not NOT1 (N1551, N1530);
buf BUF1 (N1552, N1549);
nor NOR4 (N1553, N1491, N1499, N422, N300);
buf BUF1 (N1554, N1553);
xor XOR2 (N1555, N1547, N1550);
xor XOR2 (N1556, N1373, N828);
not NOT1 (N1557, N1543);
buf BUF1 (N1558, N1551);
nand NAND2 (N1559, N1557, N1354);
or OR2 (N1560, N1526, N999);
nand NAND2 (N1561, N1559, N653);
nor NOR2 (N1562, N1556, N623);
not NOT1 (N1563, N1542);
nor NOR3 (N1564, N1560, N791, N1338);
nand NAND3 (N1565, N1554, N1355, N319);
xor XOR2 (N1566, N1558, N665);
and AND3 (N1567, N1555, N200, N205);
nand NAND4 (N1568, N1561, N491, N362, N1225);
nand NAND3 (N1569, N1552, N1027, N893);
or OR2 (N1570, N1569, N794);
buf BUF1 (N1571, N1538);
nand NAND4 (N1572, N1562, N1536, N898, N813);
and AND2 (N1573, N1572, N738);
and AND3 (N1574, N1563, N43, N824);
nand NAND2 (N1575, N1568, N1434);
buf BUF1 (N1576, N1548);
or OR3 (N1577, N1574, N1202, N952);
buf BUF1 (N1578, N1566);
not NOT1 (N1579, N1575);
or OR4 (N1580, N1567, N1480, N627, N1336);
nand NAND2 (N1581, N1573, N1565);
and AND2 (N1582, N1111, N986);
and AND4 (N1583, N1576, N942, N813, N613);
not NOT1 (N1584, N1579);
nor NOR3 (N1585, N1571, N689, N106);
and AND4 (N1586, N1564, N36, N1511, N1059);
nor NOR2 (N1587, N1581, N1103);
xor XOR2 (N1588, N1580, N72);
nor NOR2 (N1589, N1577, N98);
xor XOR2 (N1590, N1587, N1057);
or OR2 (N1591, N1586, N843);
nor NOR2 (N1592, N1588, N1257);
and AND2 (N1593, N1570, N638);
or OR3 (N1594, N1589, N910, N539);
xor XOR2 (N1595, N1578, N533);
nand NAND2 (N1596, N1590, N902);
buf BUF1 (N1597, N1596);
buf BUF1 (N1598, N1585);
or OR2 (N1599, N1583, N1559);
buf BUF1 (N1600, N1598);
buf BUF1 (N1601, N1599);
buf BUF1 (N1602, N1582);
not NOT1 (N1603, N1600);
xor XOR2 (N1604, N1602, N583);
nand NAND3 (N1605, N1584, N239, N490);
nand NAND2 (N1606, N1597, N1420);
nor NOR3 (N1607, N1603, N628, N1415);
xor XOR2 (N1608, N1594, N633);
nor NOR3 (N1609, N1601, N1017, N1293);
nor NOR2 (N1610, N1607, N488);
buf BUF1 (N1611, N1595);
xor XOR2 (N1612, N1604, N1553);
and AND2 (N1613, N1608, N1416);
buf BUF1 (N1614, N1605);
or OR4 (N1615, N1592, N1318, N152, N899);
nand NAND3 (N1616, N1611, N744, N1367);
buf BUF1 (N1617, N1591);
nand NAND2 (N1618, N1606, N165);
nand NAND2 (N1619, N1613, N1403);
nor NOR2 (N1620, N1619, N1153);
or OR2 (N1621, N1618, N650);
nand NAND2 (N1622, N1609, N725);
or OR3 (N1623, N1593, N791, N1197);
and AND3 (N1624, N1622, N66, N386);
nand NAND3 (N1625, N1610, N1517, N1488);
not NOT1 (N1626, N1615);
nand NAND2 (N1627, N1614, N1046);
xor XOR2 (N1628, N1623, N1498);
nor NOR4 (N1629, N1612, N1029, N212, N1327);
buf BUF1 (N1630, N1617);
xor XOR2 (N1631, N1627, N1085);
and AND4 (N1632, N1631, N1411, N562, N264);
buf BUF1 (N1633, N1624);
not NOT1 (N1634, N1630);
nor NOR3 (N1635, N1633, N1548, N1313);
buf BUF1 (N1636, N1620);
buf BUF1 (N1637, N1632);
not NOT1 (N1638, N1635);
nand NAND2 (N1639, N1628, N1499);
buf BUF1 (N1640, N1629);
xor XOR2 (N1641, N1625, N712);
nor NOR3 (N1642, N1637, N263, N797);
xor XOR2 (N1643, N1636, N1605);
nand NAND2 (N1644, N1639, N86);
xor XOR2 (N1645, N1638, N1484);
nand NAND4 (N1646, N1616, N1165, N1632, N581);
not NOT1 (N1647, N1640);
buf BUF1 (N1648, N1626);
nand NAND3 (N1649, N1644, N957, N33);
or OR2 (N1650, N1643, N115);
nor NOR3 (N1651, N1646, N1525, N1068);
buf BUF1 (N1652, N1645);
nand NAND2 (N1653, N1652, N279);
or OR3 (N1654, N1653, N1521, N1144);
and AND3 (N1655, N1650, N1028, N1092);
not NOT1 (N1656, N1655);
xor XOR2 (N1657, N1654, N1017);
nor NOR4 (N1658, N1651, N680, N94, N575);
not NOT1 (N1659, N1647);
nand NAND4 (N1660, N1634, N228, N301, N1185);
or OR3 (N1661, N1621, N626, N315);
nor NOR2 (N1662, N1661, N707);
xor XOR2 (N1663, N1662, N898);
or OR3 (N1664, N1657, N1164, N514);
and AND3 (N1665, N1659, N1365, N1051);
buf BUF1 (N1666, N1658);
and AND4 (N1667, N1649, N673, N1042, N1168);
or OR4 (N1668, N1660, N91, N604, N1094);
nor NOR2 (N1669, N1642, N749);
buf BUF1 (N1670, N1663);
or OR3 (N1671, N1669, N1568, N227);
and AND3 (N1672, N1666, N761, N530);
nand NAND3 (N1673, N1665, N742, N1537);
buf BUF1 (N1674, N1648);
nand NAND2 (N1675, N1656, N1429);
buf BUF1 (N1676, N1670);
buf BUF1 (N1677, N1668);
xor XOR2 (N1678, N1641, N333);
xor XOR2 (N1679, N1673, N276);
and AND4 (N1680, N1679, N113, N304, N1186);
xor XOR2 (N1681, N1677, N149);
nand NAND3 (N1682, N1678, N1186, N1370);
nand NAND4 (N1683, N1676, N1271, N1343, N1417);
or OR4 (N1684, N1680, N1100, N899, N504);
nor NOR2 (N1685, N1672, N224);
or OR4 (N1686, N1682, N1538, N1425, N247);
xor XOR2 (N1687, N1684, N1026);
nand NAND2 (N1688, N1686, N605);
and AND4 (N1689, N1667, N249, N1332, N721);
not NOT1 (N1690, N1671);
and AND4 (N1691, N1683, N1016, N1602, N300);
or OR4 (N1692, N1687, N1430, N309, N976);
buf BUF1 (N1693, N1688);
not NOT1 (N1694, N1674);
nor NOR4 (N1695, N1681, N239, N229, N680);
buf BUF1 (N1696, N1685);
and AND4 (N1697, N1694, N1491, N1343, N281);
xor XOR2 (N1698, N1696, N420);
or OR3 (N1699, N1698, N1158, N449);
xor XOR2 (N1700, N1699, N443);
and AND3 (N1701, N1675, N1604, N7);
buf BUF1 (N1702, N1690);
xor XOR2 (N1703, N1700, N1037);
nand NAND3 (N1704, N1691, N284, N197);
not NOT1 (N1705, N1692);
xor XOR2 (N1706, N1703, N1675);
or OR4 (N1707, N1693, N1037, N532, N905);
nand NAND3 (N1708, N1704, N354, N1283);
or OR2 (N1709, N1697, N1244);
nand NAND2 (N1710, N1702, N1397);
xor XOR2 (N1711, N1701, N644);
nand NAND3 (N1712, N1710, N818, N1363);
xor XOR2 (N1713, N1708, N630);
nand NAND4 (N1714, N1709, N1669, N492, N661);
nand NAND2 (N1715, N1705, N1711);
not NOT1 (N1716, N32);
or OR2 (N1717, N1695, N828);
nor NOR4 (N1718, N1716, N904, N1497, N739);
buf BUF1 (N1719, N1714);
or OR4 (N1720, N1664, N372, N1301, N1442);
not NOT1 (N1721, N1717);
nor NOR3 (N1722, N1720, N1354, N413);
buf BUF1 (N1723, N1712);
and AND4 (N1724, N1718, N780, N615, N454);
buf BUF1 (N1725, N1707);
xor XOR2 (N1726, N1723, N53);
buf BUF1 (N1727, N1726);
nand NAND4 (N1728, N1722, N1035, N74, N213);
not NOT1 (N1729, N1713);
nand NAND4 (N1730, N1727, N974, N136, N939);
nand NAND4 (N1731, N1689, N1448, N506, N1676);
nor NOR2 (N1732, N1729, N268);
buf BUF1 (N1733, N1731);
nand NAND4 (N1734, N1725, N41, N259, N218);
buf BUF1 (N1735, N1724);
nor NOR2 (N1736, N1733, N11);
xor XOR2 (N1737, N1734, N203);
not NOT1 (N1738, N1728);
xor XOR2 (N1739, N1738, N460);
xor XOR2 (N1740, N1715, N1117);
not NOT1 (N1741, N1739);
xor XOR2 (N1742, N1706, N60);
not NOT1 (N1743, N1732);
buf BUF1 (N1744, N1741);
nor NOR2 (N1745, N1742, N249);
xor XOR2 (N1746, N1740, N1166);
nor NOR4 (N1747, N1735, N1605, N1066, N1672);
not NOT1 (N1748, N1745);
nor NOR2 (N1749, N1746, N732);
nand NAND2 (N1750, N1719, N511);
not NOT1 (N1751, N1743);
xor XOR2 (N1752, N1721, N98);
xor XOR2 (N1753, N1736, N272);
nor NOR3 (N1754, N1730, N1163, N1260);
xor XOR2 (N1755, N1737, N282);
nor NOR3 (N1756, N1752, N337, N623);
not NOT1 (N1757, N1748);
or OR2 (N1758, N1755, N1309);
and AND2 (N1759, N1757, N772);
nand NAND3 (N1760, N1753, N1423, N794);
nor NOR3 (N1761, N1750, N1267, N519);
nand NAND2 (N1762, N1747, N1741);
not NOT1 (N1763, N1762);
and AND2 (N1764, N1763, N357);
buf BUF1 (N1765, N1760);
xor XOR2 (N1766, N1749, N132);
buf BUF1 (N1767, N1754);
nor NOR2 (N1768, N1764, N1146);
nor NOR4 (N1769, N1751, N1761, N509, N1496);
not NOT1 (N1770, N543);
buf BUF1 (N1771, N1768);
buf BUF1 (N1772, N1771);
not NOT1 (N1773, N1766);
and AND4 (N1774, N1770, N555, N540, N1129);
not NOT1 (N1775, N1769);
xor XOR2 (N1776, N1772, N1053);
buf BUF1 (N1777, N1774);
nor NOR4 (N1778, N1759, N331, N1675, N148);
buf BUF1 (N1779, N1765);
nand NAND3 (N1780, N1773, N663, N421);
not NOT1 (N1781, N1777);
not NOT1 (N1782, N1779);
and AND3 (N1783, N1756, N1768, N135);
or OR4 (N1784, N1780, N1327, N1061, N1061);
not NOT1 (N1785, N1758);
not NOT1 (N1786, N1767);
xor XOR2 (N1787, N1786, N660);
nor NOR4 (N1788, N1785, N626, N1406, N1278);
and AND4 (N1789, N1787, N1779, N1171, N1316);
xor XOR2 (N1790, N1776, N747);
and AND3 (N1791, N1788, N7, N1428);
or OR2 (N1792, N1744, N1129);
xor XOR2 (N1793, N1791, N131);
nor NOR4 (N1794, N1782, N1709, N413, N772);
and AND2 (N1795, N1775, N295);
nand NAND3 (N1796, N1783, N1292, N680);
nand NAND2 (N1797, N1784, N685);
nor NOR4 (N1798, N1792, N1398, N691, N361);
nand NAND4 (N1799, N1781, N1550, N422, N622);
nor NOR2 (N1800, N1794, N1697);
nor NOR4 (N1801, N1789, N1403, N78, N224);
buf BUF1 (N1802, N1801);
buf BUF1 (N1803, N1798);
buf BUF1 (N1804, N1793);
xor XOR2 (N1805, N1802, N1454);
xor XOR2 (N1806, N1796, N681);
nor NOR3 (N1807, N1806, N246, N862);
nand NAND2 (N1808, N1803, N306);
not NOT1 (N1809, N1778);
nor NOR2 (N1810, N1808, N1464);
or OR4 (N1811, N1790, N1049, N959, N1446);
nand NAND4 (N1812, N1799, N547, N1724, N1571);
xor XOR2 (N1813, N1811, N1272);
nor NOR4 (N1814, N1795, N1003, N1812, N1738);
not NOT1 (N1815, N1735);
buf BUF1 (N1816, N1814);
nor NOR4 (N1817, N1804, N1675, N27, N1277);
or OR4 (N1818, N1810, N802, N849, N1156);
or OR4 (N1819, N1817, N426, N834, N129);
nand NAND2 (N1820, N1819, N1103);
and AND2 (N1821, N1800, N972);
or OR2 (N1822, N1816, N719);
buf BUF1 (N1823, N1805);
and AND3 (N1824, N1797, N795, N111);
xor XOR2 (N1825, N1813, N842);
nand NAND3 (N1826, N1824, N1565, N1745);
nor NOR2 (N1827, N1820, N1515);
and AND4 (N1828, N1807, N1151, N122, N1262);
nand NAND4 (N1829, N1826, N148, N686, N1600);
nand NAND3 (N1830, N1825, N666, N996);
nand NAND4 (N1831, N1821, N729, N860, N180);
nor NOR4 (N1832, N1828, N366, N361, N106);
and AND4 (N1833, N1832, N1320, N668, N606);
buf BUF1 (N1834, N1833);
nor NOR2 (N1835, N1823, N1520);
xor XOR2 (N1836, N1818, N728);
buf BUF1 (N1837, N1836);
not NOT1 (N1838, N1829);
nand NAND3 (N1839, N1837, N1433, N1474);
or OR3 (N1840, N1830, N377, N433);
nand NAND2 (N1841, N1822, N71);
nor NOR2 (N1842, N1839, N1119);
buf BUF1 (N1843, N1831);
nor NOR2 (N1844, N1835, N504);
or OR2 (N1845, N1841, N1758);
buf BUF1 (N1846, N1842);
nand NAND4 (N1847, N1840, N128, N1829, N1466);
xor XOR2 (N1848, N1846, N233);
buf BUF1 (N1849, N1809);
nor NOR3 (N1850, N1827, N306, N1378);
nand NAND3 (N1851, N1815, N1609, N206);
not NOT1 (N1852, N1843);
xor XOR2 (N1853, N1847, N1684);
buf BUF1 (N1854, N1848);
not NOT1 (N1855, N1853);
buf BUF1 (N1856, N1850);
buf BUF1 (N1857, N1849);
or OR4 (N1858, N1851, N1507, N1698, N401);
and AND2 (N1859, N1857, N977);
nor NOR4 (N1860, N1845, N327, N1197, N870);
or OR2 (N1861, N1838, N695);
nor NOR2 (N1862, N1861, N915);
and AND3 (N1863, N1852, N450, N1298);
nor NOR4 (N1864, N1844, N374, N1684, N1264);
nor NOR3 (N1865, N1859, N1418, N1018);
and AND2 (N1866, N1865, N1139);
buf BUF1 (N1867, N1858);
buf BUF1 (N1868, N1866);
nor NOR4 (N1869, N1864, N304, N1504, N824);
not NOT1 (N1870, N1856);
not NOT1 (N1871, N1834);
and AND2 (N1872, N1870, N1714);
nand NAND3 (N1873, N1868, N476, N1838);
buf BUF1 (N1874, N1869);
xor XOR2 (N1875, N1874, N723);
xor XOR2 (N1876, N1873, N1755);
nor NOR2 (N1877, N1872, N495);
nand NAND2 (N1878, N1871, N771);
nand NAND2 (N1879, N1862, N1633);
not NOT1 (N1880, N1877);
xor XOR2 (N1881, N1876, N30);
nand NAND4 (N1882, N1878, N1254, N284, N719);
and AND2 (N1883, N1854, N441);
nand NAND4 (N1884, N1881, N1798, N1473, N1241);
buf BUF1 (N1885, N1867);
nor NOR2 (N1886, N1855, N829);
xor XOR2 (N1887, N1883, N697);
nor NOR3 (N1888, N1863, N825, N1877);
nor NOR4 (N1889, N1882, N174, N435, N837);
xor XOR2 (N1890, N1886, N6);
nor NOR2 (N1891, N1889, N881);
buf BUF1 (N1892, N1885);
buf BUF1 (N1893, N1891);
or OR4 (N1894, N1890, N1588, N1576, N881);
buf BUF1 (N1895, N1884);
and AND2 (N1896, N1879, N269);
buf BUF1 (N1897, N1894);
buf BUF1 (N1898, N1895);
nand NAND4 (N1899, N1875, N641, N388, N1147);
nand NAND2 (N1900, N1892, N574);
not NOT1 (N1901, N1888);
nor NOR4 (N1902, N1860, N351, N1343, N921);
xor XOR2 (N1903, N1897, N715);
buf BUF1 (N1904, N1898);
nor NOR4 (N1905, N1901, N844, N1188, N1272);
nand NAND4 (N1906, N1893, N465, N1820, N127);
not NOT1 (N1907, N1900);
nand NAND2 (N1908, N1907, N1711);
and AND3 (N1909, N1899, N391, N252);
or OR3 (N1910, N1903, N1762, N635);
nor NOR2 (N1911, N1908, N1525);
nand NAND2 (N1912, N1902, N1288);
nor NOR2 (N1913, N1880, N1794);
buf BUF1 (N1914, N1904);
buf BUF1 (N1915, N1912);
and AND2 (N1916, N1914, N613);
or OR2 (N1917, N1906, N1417);
and AND4 (N1918, N1915, N12, N1055, N108);
not NOT1 (N1919, N1913);
and AND2 (N1920, N1909, N309);
nand NAND4 (N1921, N1917, N1410, N1153, N937);
nor NOR3 (N1922, N1896, N769, N962);
nor NOR2 (N1923, N1910, N1317);
and AND2 (N1924, N1905, N1249);
nand NAND4 (N1925, N1921, N269, N959, N1353);
nor NOR4 (N1926, N1916, N259, N1323, N1891);
nor NOR3 (N1927, N1924, N277, N709);
buf BUF1 (N1928, N1918);
not NOT1 (N1929, N1923);
nand NAND3 (N1930, N1925, N1274, N1418);
nand NAND4 (N1931, N1887, N1656, N1657, N451);
or OR2 (N1932, N1930, N1567);
or OR4 (N1933, N1920, N897, N1271, N1860);
not NOT1 (N1934, N1922);
buf BUF1 (N1935, N1928);
nor NOR2 (N1936, N1935, N479);
buf BUF1 (N1937, N1911);
nor NOR4 (N1938, N1936, N1770, N1597, N1058);
or OR4 (N1939, N1934, N690, N557, N1396);
buf BUF1 (N1940, N1931);
xor XOR2 (N1941, N1937, N352);
not NOT1 (N1942, N1929);
xor XOR2 (N1943, N1919, N20);
nor NOR4 (N1944, N1942, N209, N1803, N168);
or OR2 (N1945, N1938, N46);
buf BUF1 (N1946, N1943);
xor XOR2 (N1947, N1944, N274);
nand NAND2 (N1948, N1947, N380);
not NOT1 (N1949, N1945);
nor NOR2 (N1950, N1948, N1070);
buf BUF1 (N1951, N1926);
nor NOR4 (N1952, N1941, N1634, N642, N1055);
nor NOR3 (N1953, N1950, N1251, N1177);
buf BUF1 (N1954, N1940);
not NOT1 (N1955, N1939);
not NOT1 (N1956, N1933);
or OR4 (N1957, N1953, N1590, N102, N194);
not NOT1 (N1958, N1951);
and AND3 (N1959, N1932, N1327, N719);
or OR2 (N1960, N1955, N1707);
nor NOR4 (N1961, N1927, N1904, N1302, N1666);
nor NOR4 (N1962, N1949, N439, N86, N1067);
xor XOR2 (N1963, N1962, N309);
buf BUF1 (N1964, N1963);
buf BUF1 (N1965, N1957);
or OR2 (N1966, N1965, N238);
xor XOR2 (N1967, N1946, N62);
and AND4 (N1968, N1966, N2, N1652, N708);
buf BUF1 (N1969, N1960);
and AND2 (N1970, N1969, N275);
nor NOR2 (N1971, N1967, N1041);
nand NAND2 (N1972, N1956, N1492);
and AND4 (N1973, N1968, N1573, N204, N1900);
xor XOR2 (N1974, N1952, N49);
or OR2 (N1975, N1971, N982);
or OR3 (N1976, N1964, N1903, N143);
xor XOR2 (N1977, N1954, N351);
xor XOR2 (N1978, N1973, N1132);
nor NOR4 (N1979, N1978, N691, N1257, N398);
xor XOR2 (N1980, N1979, N1440);
xor XOR2 (N1981, N1974, N303);
xor XOR2 (N1982, N1961, N63);
buf BUF1 (N1983, N1970);
and AND4 (N1984, N1975, N1379, N1213, N554);
xor XOR2 (N1985, N1981, N835);
nand NAND2 (N1986, N1959, N1884);
xor XOR2 (N1987, N1972, N1263);
buf BUF1 (N1988, N1983);
xor XOR2 (N1989, N1977, N319);
not NOT1 (N1990, N1986);
xor XOR2 (N1991, N1958, N1237);
buf BUF1 (N1992, N1985);
nor NOR2 (N1993, N1980, N1314);
nand NAND2 (N1994, N1991, N379);
nor NOR3 (N1995, N1982, N1957, N514);
and AND3 (N1996, N1992, N889, N946);
and AND3 (N1997, N1988, N788, N1732);
nand NAND2 (N1998, N1995, N1587);
or OR4 (N1999, N1994, N1706, N1562, N151);
and AND3 (N2000, N1998, N1484, N1976);
and AND2 (N2001, N436, N1972);
nor NOR4 (N2002, N1987, N559, N1748, N377);
or OR4 (N2003, N1984, N1288, N686, N971);
nand NAND3 (N2004, N1999, N6, N457);
or OR4 (N2005, N2000, N88, N1904, N418);
buf BUF1 (N2006, N1990);
buf BUF1 (N2007, N1993);
nand NAND4 (N2008, N2003, N1651, N240, N981);
nor NOR3 (N2009, N2007, N1103, N1893);
and AND3 (N2010, N1996, N661, N1878);
or OR3 (N2011, N2002, N254, N477);
nand NAND2 (N2012, N1989, N1165);
buf BUF1 (N2013, N2010);
or OR2 (N2014, N1997, N812);
and AND2 (N2015, N2009, N1909);
and AND4 (N2016, N2005, N1298, N1, N1205);
nor NOR4 (N2017, N2014, N919, N622, N1574);
not NOT1 (N2018, N2011);
buf BUF1 (N2019, N2017);
xor XOR2 (N2020, N2001, N457);
xor XOR2 (N2021, N2004, N558);
buf BUF1 (N2022, N2013);
not NOT1 (N2023, N2016);
and AND4 (N2024, N2006, N211, N214, N473);
not NOT1 (N2025, N2021);
not NOT1 (N2026, N2022);
not NOT1 (N2027, N2023);
buf BUF1 (N2028, N2019);
nand NAND2 (N2029, N2012, N937);
not NOT1 (N2030, N2025);
not NOT1 (N2031, N2020);
not NOT1 (N2032, N2027);
or OR3 (N2033, N2015, N257, N445);
xor XOR2 (N2034, N2018, N1832);
or OR4 (N2035, N2008, N541, N1899, N279);
nand NAND2 (N2036, N2026, N118);
xor XOR2 (N2037, N2030, N1728);
nor NOR2 (N2038, N2028, N815);
not NOT1 (N2039, N2032);
nor NOR3 (N2040, N2033, N943, N1844);
nor NOR3 (N2041, N2037, N1919, N1309);
or OR3 (N2042, N2038, N1787, N416);
nand NAND4 (N2043, N2036, N1379, N189, N317);
buf BUF1 (N2044, N2035);
not NOT1 (N2045, N2034);
nand NAND2 (N2046, N2029, N907);
xor XOR2 (N2047, N2046, N1688);
buf BUF1 (N2048, N2031);
not NOT1 (N2049, N2047);
nand NAND3 (N2050, N2044, N1879, N1888);
and AND4 (N2051, N2024, N299, N1736, N1726);
xor XOR2 (N2052, N2048, N1155);
nand NAND3 (N2053, N2039, N933, N207);
or OR4 (N2054, N2041, N1950, N932, N525);
xor XOR2 (N2055, N2043, N620);
xor XOR2 (N2056, N2054, N1783);
nand NAND4 (N2057, N2055, N1577, N613, N784);
and AND4 (N2058, N2050, N1532, N1769, N1886);
and AND4 (N2059, N2040, N580, N578, N1745);
xor XOR2 (N2060, N2053, N1437);
and AND4 (N2061, N2060, N426, N58, N2046);
nor NOR4 (N2062, N2056, N1317, N346, N1380);
nand NAND3 (N2063, N2057, N1053, N597);
nor NOR2 (N2064, N2058, N607);
xor XOR2 (N2065, N2045, N618);
or OR4 (N2066, N2064, N1555, N836, N1872);
or OR2 (N2067, N2051, N596);
not NOT1 (N2068, N2067);
and AND3 (N2069, N2062, N1813, N1217);
xor XOR2 (N2070, N2052, N2);
and AND3 (N2071, N2065, N834, N540);
and AND3 (N2072, N2063, N1934, N1603);
buf BUF1 (N2073, N2059);
buf BUF1 (N2074, N2061);
and AND2 (N2075, N2049, N916);
xor XOR2 (N2076, N2042, N896);
nor NOR2 (N2077, N2073, N563);
nand NAND4 (N2078, N2070, N71, N166, N1635);
and AND4 (N2079, N2066, N597, N550, N1850);
not NOT1 (N2080, N2071);
nor NOR2 (N2081, N2074, N1829);
not NOT1 (N2082, N2075);
or OR4 (N2083, N2076, N1480, N1015, N1625);
nor NOR2 (N2084, N2082, N1455);
nor NOR3 (N2085, N2081, N1029, N417);
or OR4 (N2086, N2080, N1334, N550, N919);
and AND3 (N2087, N2083, N1209, N734);
nor NOR3 (N2088, N2079, N653, N93);
not NOT1 (N2089, N2085);
nand NAND3 (N2090, N2086, N1316, N1437);
buf BUF1 (N2091, N2084);
and AND4 (N2092, N2068, N185, N714, N1693);
nor NOR2 (N2093, N2078, N65);
xor XOR2 (N2094, N2090, N1827);
xor XOR2 (N2095, N2087, N2011);
xor XOR2 (N2096, N2077, N367);
not NOT1 (N2097, N2091);
buf BUF1 (N2098, N2094);
nand NAND3 (N2099, N2072, N932, N2064);
or OR3 (N2100, N2069, N433, N411);
xor XOR2 (N2101, N2100, N2083);
nand NAND3 (N2102, N2089, N1089, N617);
nand NAND2 (N2103, N2101, N637);
nand NAND4 (N2104, N2088, N1068, N1122, N2084);
and AND2 (N2105, N2097, N720);
buf BUF1 (N2106, N2092);
or OR4 (N2107, N2102, N274, N48, N2088);
or OR2 (N2108, N2098, N1987);
nor NOR4 (N2109, N2096, N1495, N381, N1992);
and AND3 (N2110, N2107, N661, N1065);
or OR4 (N2111, N2104, N1792, N1425, N1672);
not NOT1 (N2112, N2108);
and AND2 (N2113, N2099, N38);
buf BUF1 (N2114, N2109);
buf BUF1 (N2115, N2103);
buf BUF1 (N2116, N2105);
not NOT1 (N2117, N2093);
and AND3 (N2118, N2110, N27, N1627);
not NOT1 (N2119, N2117);
nor NOR2 (N2120, N2095, N1789);
and AND3 (N2121, N2120, N858, N988);
not NOT1 (N2122, N2118);
buf BUF1 (N2123, N2115);
xor XOR2 (N2124, N2122, N1960);
buf BUF1 (N2125, N2119);
buf BUF1 (N2126, N2113);
and AND2 (N2127, N2121, N738);
not NOT1 (N2128, N2112);
not NOT1 (N2129, N2111);
not NOT1 (N2130, N2126);
not NOT1 (N2131, N2124);
and AND2 (N2132, N2116, N1383);
buf BUF1 (N2133, N2125);
and AND4 (N2134, N2129, N1191, N1081, N1300);
not NOT1 (N2135, N2133);
not NOT1 (N2136, N2114);
not NOT1 (N2137, N2132);
nand NAND2 (N2138, N2130, N1055);
xor XOR2 (N2139, N2123, N1689);
and AND2 (N2140, N2137, N1935);
or OR2 (N2141, N2135, N1933);
nor NOR2 (N2142, N2127, N651);
nand NAND4 (N2143, N2128, N1150, N1336, N72);
or OR3 (N2144, N2140, N1864, N1332);
nor NOR3 (N2145, N2134, N1206, N731);
not NOT1 (N2146, N2142);
and AND2 (N2147, N2144, N702);
nor NOR3 (N2148, N2138, N787, N844);
buf BUF1 (N2149, N2136);
buf BUF1 (N2150, N2143);
xor XOR2 (N2151, N2145, N1821);
buf BUF1 (N2152, N2141);
and AND3 (N2153, N2151, N72, N1534);
buf BUF1 (N2154, N2148);
and AND4 (N2155, N2139, N1452, N1341, N1461);
buf BUF1 (N2156, N2152);
nand NAND4 (N2157, N2154, N1494, N1221, N1587);
or OR4 (N2158, N2157, N975, N1132, N677);
not NOT1 (N2159, N2149);
xor XOR2 (N2160, N2106, N551);
nand NAND2 (N2161, N2150, N236);
nor NOR4 (N2162, N2153, N1824, N1739, N703);
and AND3 (N2163, N2161, N1007, N496);
or OR2 (N2164, N2159, N1278);
not NOT1 (N2165, N2164);
xor XOR2 (N2166, N2162, N1781);
nor NOR2 (N2167, N2131, N843);
or OR3 (N2168, N2166, N747, N1073);
not NOT1 (N2169, N2156);
xor XOR2 (N2170, N2146, N638);
or OR4 (N2171, N2169, N662, N1964, N1894);
and AND3 (N2172, N2163, N960, N446);
buf BUF1 (N2173, N2147);
or OR3 (N2174, N2155, N1382, N851);
or OR3 (N2175, N2173, N1817, N157);
or OR3 (N2176, N2172, N2155, N2149);
not NOT1 (N2177, N2168);
xor XOR2 (N2178, N2158, N2076);
buf BUF1 (N2179, N2167);
xor XOR2 (N2180, N2179, N1168);
nor NOR4 (N2181, N2171, N518, N934, N1006);
or OR4 (N2182, N2174, N1484, N149, N772);
nand NAND4 (N2183, N2181, N1709, N1866, N616);
nand NAND3 (N2184, N2176, N2115, N1257);
xor XOR2 (N2185, N2170, N18);
or OR3 (N2186, N2184, N1976, N130);
and AND3 (N2187, N2178, N1744, N1378);
buf BUF1 (N2188, N2175);
not NOT1 (N2189, N2165);
and AND4 (N2190, N2160, N777, N2086, N2105);
buf BUF1 (N2191, N2186);
xor XOR2 (N2192, N2177, N839);
and AND2 (N2193, N2183, N740);
or OR3 (N2194, N2191, N1896, N876);
and AND2 (N2195, N2182, N961);
or OR3 (N2196, N2187, N72, N1051);
and AND3 (N2197, N2196, N1324, N195);
xor XOR2 (N2198, N2189, N886);
nand NAND3 (N2199, N2195, N812, N1013);
and AND4 (N2200, N2193, N111, N18, N501);
xor XOR2 (N2201, N2198, N2011);
nand NAND3 (N2202, N2194, N1265, N1289);
and AND2 (N2203, N2199, N740);
or OR2 (N2204, N2188, N2078);
nand NAND2 (N2205, N2197, N1967);
not NOT1 (N2206, N2205);
and AND2 (N2207, N2206, N674);
not NOT1 (N2208, N2200);
not NOT1 (N2209, N2203);
nand NAND4 (N2210, N2190, N1029, N3, N2062);
nand NAND2 (N2211, N2180, N1342);
not NOT1 (N2212, N2210);
not NOT1 (N2213, N2212);
buf BUF1 (N2214, N2209);
and AND3 (N2215, N2211, N1661, N1549);
nor NOR3 (N2216, N2215, N349, N1518);
nand NAND3 (N2217, N2201, N1581, N390);
nand NAND4 (N2218, N2216, N621, N1942, N359);
not NOT1 (N2219, N2204);
xor XOR2 (N2220, N2219, N1380);
nor NOR2 (N2221, N2214, N1112);
not NOT1 (N2222, N2218);
xor XOR2 (N2223, N2217, N2030);
or OR3 (N2224, N2223, N1420, N1850);
and AND4 (N2225, N2213, N133, N1836, N881);
or OR4 (N2226, N2192, N387, N1386, N232);
or OR4 (N2227, N2185, N576, N358, N129);
and AND3 (N2228, N2202, N194, N1842);
not NOT1 (N2229, N2227);
or OR3 (N2230, N2225, N1676, N871);
nand NAND3 (N2231, N2220, N1283, N2064);
and AND4 (N2232, N2208, N1178, N379, N918);
nor NOR4 (N2233, N2224, N2001, N1881, N2016);
not NOT1 (N2234, N2228);
not NOT1 (N2235, N2230);
and AND2 (N2236, N2226, N1482);
or OR2 (N2237, N2235, N1552);
nor NOR2 (N2238, N2236, N1876);
or OR2 (N2239, N2238, N255);
or OR4 (N2240, N2234, N1083, N713, N742);
buf BUF1 (N2241, N2239);
and AND4 (N2242, N2229, N1876, N953, N1040);
nand NAND4 (N2243, N2240, N1059, N1334, N2112);
nand NAND4 (N2244, N2231, N2133, N713, N1121);
buf BUF1 (N2245, N2232);
nand NAND2 (N2246, N2242, N1554);
and AND2 (N2247, N2237, N10);
not NOT1 (N2248, N2246);
nor NOR3 (N2249, N2221, N1279, N1778);
nor NOR2 (N2250, N2243, N997);
not NOT1 (N2251, N2248);
xor XOR2 (N2252, N2250, N2008);
xor XOR2 (N2253, N2222, N325);
buf BUF1 (N2254, N2249);
xor XOR2 (N2255, N2247, N1962);
not NOT1 (N2256, N2241);
buf BUF1 (N2257, N2254);
or OR4 (N2258, N2251, N730, N666, N1723);
nor NOR2 (N2259, N2256, N626);
not NOT1 (N2260, N2258);
nor NOR2 (N2261, N2252, N773);
nor NOR4 (N2262, N2257, N910, N1639, N1242);
and AND2 (N2263, N2253, N210);
nor NOR4 (N2264, N2261, N399, N1950, N1373);
nor NOR4 (N2265, N2264, N1333, N1745, N1660);
not NOT1 (N2266, N2262);
not NOT1 (N2267, N2244);
xor XOR2 (N2268, N2266, N487);
nand NAND4 (N2269, N2233, N2181, N1646, N443);
nor NOR4 (N2270, N2207, N1089, N1963, N1594);
and AND3 (N2271, N2260, N1783, N203);
or OR4 (N2272, N2245, N489, N771, N1459);
not NOT1 (N2273, N2270);
nand NAND4 (N2274, N2265, N1718, N1340, N1244);
nand NAND3 (N2275, N2273, N527, N12);
xor XOR2 (N2276, N2259, N238);
nand NAND2 (N2277, N2263, N267);
buf BUF1 (N2278, N2272);
nor NOR3 (N2279, N2268, N1845, N2131);
not NOT1 (N2280, N2255);
and AND2 (N2281, N2269, N1145);
and AND4 (N2282, N2277, N6, N1324, N446);
not NOT1 (N2283, N2278);
buf BUF1 (N2284, N2271);
not NOT1 (N2285, N2281);
or OR2 (N2286, N2285, N1598);
buf BUF1 (N2287, N2280);
not NOT1 (N2288, N2286);
and AND4 (N2289, N2279, N302, N1018, N367);
and AND2 (N2290, N2283, N2150);
buf BUF1 (N2291, N2290);
nor NOR2 (N2292, N2274, N838);
nand NAND3 (N2293, N2282, N999, N231);
and AND3 (N2294, N2293, N253, N334);
buf BUF1 (N2295, N2288);
and AND3 (N2296, N2267, N1569, N2125);
nor NOR3 (N2297, N2284, N752, N1061);
nand NAND2 (N2298, N2287, N938);
nand NAND4 (N2299, N2291, N411, N2136, N170);
not NOT1 (N2300, N2297);
nor NOR3 (N2301, N2276, N1599, N581);
or OR2 (N2302, N2294, N2175);
nand NAND3 (N2303, N2292, N2015, N300);
xor XOR2 (N2304, N2295, N123);
xor XOR2 (N2305, N2289, N1192);
nand NAND3 (N2306, N2298, N428, N1435);
not NOT1 (N2307, N2303);
or OR2 (N2308, N2306, N1187);
buf BUF1 (N2309, N2302);
and AND2 (N2310, N2299, N856);
xor XOR2 (N2311, N2300, N1844);
nor NOR2 (N2312, N2296, N87);
or OR3 (N2313, N2311, N76, N1996);
nand NAND3 (N2314, N2309, N1983, N242);
and AND4 (N2315, N2312, N1003, N1226, N2117);
nor NOR3 (N2316, N2305, N363, N1202);
buf BUF1 (N2317, N2316);
and AND2 (N2318, N2315, N2149);
nor NOR3 (N2319, N2307, N1459, N1910);
buf BUF1 (N2320, N2317);
nor NOR2 (N2321, N2308, N1076);
nor NOR3 (N2322, N2301, N2165, N2115);
or OR3 (N2323, N2310, N325, N1218);
not NOT1 (N2324, N2275);
nand NAND4 (N2325, N2318, N1146, N305, N1135);
or OR4 (N2326, N2304, N2006, N712, N1610);
and AND4 (N2327, N2323, N1506, N909, N201);
and AND2 (N2328, N2324, N1441);
and AND3 (N2329, N2325, N906, N1229);
and AND2 (N2330, N2313, N341);
buf BUF1 (N2331, N2328);
nand NAND3 (N2332, N2327, N1441, N423);
nand NAND3 (N2333, N2320, N2088, N1460);
not NOT1 (N2334, N2326);
xor XOR2 (N2335, N2319, N1995);
or OR3 (N2336, N2314, N60, N1372);
nor NOR2 (N2337, N2321, N1035);
xor XOR2 (N2338, N2334, N190);
nand NAND4 (N2339, N2329, N87, N479, N173);
nand NAND4 (N2340, N2330, N967, N878, N1870);
xor XOR2 (N2341, N2340, N1874);
nor NOR2 (N2342, N2336, N558);
xor XOR2 (N2343, N2335, N1924);
buf BUF1 (N2344, N2341);
or OR4 (N2345, N2333, N284, N1020, N1956);
nand NAND3 (N2346, N2337, N684, N925);
nand NAND3 (N2347, N2344, N1122, N540);
not NOT1 (N2348, N2339);
or OR2 (N2349, N2346, N1744);
or OR3 (N2350, N2343, N1357, N2182);
buf BUF1 (N2351, N2338);
nor NOR4 (N2352, N2348, N1693, N2270, N1896);
nor NOR3 (N2353, N2351, N2223, N1044);
or OR4 (N2354, N2322, N1587, N2349, N341);
and AND2 (N2355, N1651, N1435);
buf BUF1 (N2356, N2354);
and AND4 (N2357, N2332, N177, N1079, N25);
and AND2 (N2358, N2352, N2011);
buf BUF1 (N2359, N2355);
and AND4 (N2360, N2331, N350, N1070, N1191);
buf BUF1 (N2361, N2358);
not NOT1 (N2362, N2350);
nand NAND2 (N2363, N2359, N59);
nand NAND4 (N2364, N2360, N1047, N1211, N1933);
xor XOR2 (N2365, N2356, N1880);
nor NOR3 (N2366, N2353, N449, N2158);
xor XOR2 (N2367, N2365, N1423);
and AND4 (N2368, N2362, N1232, N1551, N1159);
nor NOR4 (N2369, N2345, N1191, N1614, N160);
or OR2 (N2370, N2367, N862);
nand NAND3 (N2371, N2370, N2252, N996);
xor XOR2 (N2372, N2369, N355);
nand NAND3 (N2373, N2342, N2093, N622);
nor NOR2 (N2374, N2347, N545);
or OR2 (N2375, N2373, N326);
xor XOR2 (N2376, N2361, N1481);
not NOT1 (N2377, N2372);
or OR2 (N2378, N2376, N1068);
nand NAND4 (N2379, N2368, N365, N1663, N620);
and AND4 (N2380, N2366, N1629, N491, N1977);
nor NOR3 (N2381, N2363, N1147, N743);
buf BUF1 (N2382, N2371);
not NOT1 (N2383, N2379);
and AND4 (N2384, N2357, N1196, N309, N2348);
buf BUF1 (N2385, N2380);
buf BUF1 (N2386, N2385);
buf BUF1 (N2387, N2384);
and AND4 (N2388, N2378, N1929, N865, N2339);
nand NAND3 (N2389, N2377, N2101, N311);
or OR2 (N2390, N2375, N1867);
or OR3 (N2391, N2386, N734, N1923);
not NOT1 (N2392, N2364);
buf BUF1 (N2393, N2374);
nor NOR4 (N2394, N2383, N2040, N1173, N965);
xor XOR2 (N2395, N2394, N1483);
xor XOR2 (N2396, N2382, N1447);
not NOT1 (N2397, N2387);
nor NOR3 (N2398, N2381, N611, N2385);
nor NOR4 (N2399, N2397, N848, N289, N2388);
xor XOR2 (N2400, N927, N1282);
not NOT1 (N2401, N2392);
buf BUF1 (N2402, N2400);
nor NOR2 (N2403, N2396, N1629);
xor XOR2 (N2404, N2393, N1962);
nor NOR2 (N2405, N2401, N1743);
nor NOR3 (N2406, N2403, N1149, N549);
xor XOR2 (N2407, N2406, N807);
buf BUF1 (N2408, N2398);
nand NAND4 (N2409, N2389, N1845, N802, N66);
nand NAND4 (N2410, N2409, N1782, N409, N1939);
buf BUF1 (N2411, N2391);
nand NAND3 (N2412, N2395, N76, N329);
xor XOR2 (N2413, N2412, N1619);
nand NAND2 (N2414, N2413, N1043);
and AND4 (N2415, N2411, N2373, N358, N1133);
nand NAND2 (N2416, N2399, N1570);
nand NAND3 (N2417, N2407, N805, N955);
or OR4 (N2418, N2390, N1590, N377, N284);
nor NOR2 (N2419, N2417, N444);
nand NAND4 (N2420, N2415, N786, N187, N1554);
or OR4 (N2421, N2416, N2203, N2269, N616);
or OR3 (N2422, N2419, N2401, N1369);
buf BUF1 (N2423, N2420);
nand NAND3 (N2424, N2414, N249, N607);
or OR2 (N2425, N2408, N368);
and AND4 (N2426, N2418, N1581, N747, N2399);
and AND4 (N2427, N2421, N1820, N1060, N2096);
and AND2 (N2428, N2402, N2072);
nand NAND4 (N2429, N2410, N674, N1951, N1242);
or OR3 (N2430, N2425, N1330, N1096);
nor NOR2 (N2431, N2429, N1359);
nor NOR4 (N2432, N2423, N1955, N1128, N45);
and AND2 (N2433, N2430, N1383);
not NOT1 (N2434, N2432);
not NOT1 (N2435, N2422);
nand NAND3 (N2436, N2426, N32, N663);
not NOT1 (N2437, N2431);
or OR2 (N2438, N2405, N2207);
buf BUF1 (N2439, N2434);
not NOT1 (N2440, N2436);
xor XOR2 (N2441, N2424, N2182);
buf BUF1 (N2442, N2441);
buf BUF1 (N2443, N2437);
and AND3 (N2444, N2440, N1209, N1486);
xor XOR2 (N2445, N2439, N1300);
nor NOR4 (N2446, N2435, N1780, N336, N206);
not NOT1 (N2447, N2438);
and AND3 (N2448, N2447, N559, N1610);
nor NOR4 (N2449, N2404, N948, N1588, N1377);
xor XOR2 (N2450, N2449, N493);
xor XOR2 (N2451, N2446, N1874);
buf BUF1 (N2452, N2445);
nor NOR3 (N2453, N2451, N169, N55);
not NOT1 (N2454, N2453);
and AND3 (N2455, N2433, N324, N968);
nand NAND3 (N2456, N2455, N871, N1745);
buf BUF1 (N2457, N2450);
or OR2 (N2458, N2452, N1639);
not NOT1 (N2459, N2454);
nand NAND4 (N2460, N2444, N787, N1775, N1672);
or OR4 (N2461, N2456, N1529, N1386, N365);
or OR4 (N2462, N2442, N1960, N1068, N746);
xor XOR2 (N2463, N2458, N184);
nand NAND3 (N2464, N2459, N1158, N2176);
nor NOR4 (N2465, N2462, N2451, N1835, N2391);
xor XOR2 (N2466, N2427, N713);
xor XOR2 (N2467, N2428, N1862);
nor NOR3 (N2468, N2461, N694, N1407);
nand NAND3 (N2469, N2443, N1863, N486);
nor NOR4 (N2470, N2457, N2375, N1673, N279);
nor NOR2 (N2471, N2469, N1830);
or OR2 (N2472, N2467, N754);
and AND2 (N2473, N2460, N631);
and AND3 (N2474, N2470, N519, N2356);
or OR4 (N2475, N2468, N240, N2404, N1021);
and AND3 (N2476, N2471, N930, N1710);
nand NAND2 (N2477, N2474, N522);
and AND2 (N2478, N2472, N754);
not NOT1 (N2479, N2475);
nor NOR3 (N2480, N2477, N1765, N1362);
xor XOR2 (N2481, N2480, N1238);
nor NOR4 (N2482, N2478, N1656, N844, N1346);
nor NOR2 (N2483, N2448, N1285);
not NOT1 (N2484, N2481);
and AND3 (N2485, N2482, N1890, N852);
and AND4 (N2486, N2466, N446, N446, N425);
nand NAND4 (N2487, N2485, N449, N138, N1661);
nand NAND3 (N2488, N2464, N1629, N2384);
and AND3 (N2489, N2463, N16, N1314);
xor XOR2 (N2490, N2488, N775);
xor XOR2 (N2491, N2484, N1770);
or OR3 (N2492, N2490, N439, N1727);
and AND3 (N2493, N2486, N1590, N983);
and AND4 (N2494, N2491, N2259, N225, N1892);
nor NOR2 (N2495, N2492, N55);
or OR2 (N2496, N2493, N1295);
xor XOR2 (N2497, N2496, N739);
nor NOR4 (N2498, N2473, N129, N1026, N393);
nor NOR2 (N2499, N2497, N314);
xor XOR2 (N2500, N2494, N1086);
not NOT1 (N2501, N2499);
not NOT1 (N2502, N2498);
xor XOR2 (N2503, N2502, N540);
buf BUF1 (N2504, N2495);
and AND2 (N2505, N2487, N2495);
nor NOR2 (N2506, N2476, N1208);
xor XOR2 (N2507, N2501, N2006);
nand NAND4 (N2508, N2483, N1227, N2107, N1079);
not NOT1 (N2509, N2489);
xor XOR2 (N2510, N2479, N1595);
not NOT1 (N2511, N2505);
nor NOR2 (N2512, N2510, N1754);
or OR3 (N2513, N2500, N2316, N1455);
not NOT1 (N2514, N2508);
and AND3 (N2515, N2509, N2063, N629);
xor XOR2 (N2516, N2511, N928);
nor NOR2 (N2517, N2465, N2353);
nand NAND4 (N2518, N2513, N1822, N1761, N1431);
buf BUF1 (N2519, N2516);
buf BUF1 (N2520, N2517);
xor XOR2 (N2521, N2503, N77);
nor NOR3 (N2522, N2514, N1583, N162);
nand NAND3 (N2523, N2512, N1130, N1343);
nor NOR2 (N2524, N2521, N1694);
nand NAND2 (N2525, N2523, N432);
nor NOR4 (N2526, N2524, N20, N1694, N287);
buf BUF1 (N2527, N2526);
nand NAND4 (N2528, N2518, N2300, N152, N2342);
xor XOR2 (N2529, N2527, N409);
not NOT1 (N2530, N2520);
buf BUF1 (N2531, N2522);
and AND2 (N2532, N2519, N2136);
or OR3 (N2533, N2506, N1804, N1328);
not NOT1 (N2534, N2533);
nand NAND3 (N2535, N2528, N1968, N855);
xor XOR2 (N2536, N2534, N499);
nor NOR4 (N2537, N2515, N2051, N1040, N324);
buf BUF1 (N2538, N2536);
nand NAND4 (N2539, N2525, N16, N301, N495);
buf BUF1 (N2540, N2529);
buf BUF1 (N2541, N2538);
xor XOR2 (N2542, N2507, N1092);
not NOT1 (N2543, N2539);
and AND3 (N2544, N2540, N1679, N2268);
or OR2 (N2545, N2544, N2158);
xor XOR2 (N2546, N2543, N299);
nand NAND3 (N2547, N2542, N1047, N988);
nand NAND2 (N2548, N2546, N67);
and AND4 (N2549, N2545, N176, N1858, N756);
nor NOR3 (N2550, N2532, N2076, N435);
or OR3 (N2551, N2549, N950, N2332);
nor NOR2 (N2552, N2541, N1550);
nor NOR3 (N2553, N2531, N1101, N735);
nand NAND2 (N2554, N2504, N1725);
or OR4 (N2555, N2537, N1816, N2063, N279);
buf BUF1 (N2556, N2548);
and AND4 (N2557, N2556, N1498, N1150, N99);
not NOT1 (N2558, N2535);
or OR2 (N2559, N2557, N734);
xor XOR2 (N2560, N2559, N2161);
nand NAND4 (N2561, N2558, N1996, N1909, N1491);
xor XOR2 (N2562, N2551, N1992);
nand NAND2 (N2563, N2530, N357);
nor NOR3 (N2564, N2547, N1822, N608);
or OR3 (N2565, N2552, N67, N1341);
or OR4 (N2566, N2564, N916, N2527, N7);
or OR4 (N2567, N2553, N2101, N1948, N2344);
or OR3 (N2568, N2563, N440, N44);
not NOT1 (N2569, N2567);
and AND2 (N2570, N2561, N288);
or OR2 (N2571, N2570, N2410);
not NOT1 (N2572, N2560);
xor XOR2 (N2573, N2565, N182);
not NOT1 (N2574, N2571);
and AND4 (N2575, N2569, N363, N608, N2410);
not NOT1 (N2576, N2568);
or OR2 (N2577, N2550, N1817);
and AND4 (N2578, N2562, N2425, N363, N1312);
and AND3 (N2579, N2574, N1322, N2298);
or OR3 (N2580, N2572, N1398, N502);
buf BUF1 (N2581, N2575);
xor XOR2 (N2582, N2577, N4);
and AND4 (N2583, N2582, N1476, N621, N1770);
buf BUF1 (N2584, N2576);
nand NAND3 (N2585, N2578, N963, N95);
and AND3 (N2586, N2579, N2228, N2275);
or OR3 (N2587, N2583, N1713, N2512);
and AND4 (N2588, N2580, N1996, N1562, N2459);
nand NAND3 (N2589, N2585, N1422, N408);
or OR2 (N2590, N2586, N356);
buf BUF1 (N2591, N2590);
buf BUF1 (N2592, N2588);
and AND3 (N2593, N2587, N1832, N1683);
or OR2 (N2594, N2584, N814);
not NOT1 (N2595, N2566);
nand NAND3 (N2596, N2591, N2564, N807);
buf BUF1 (N2597, N2592);
xor XOR2 (N2598, N2593, N2137);
xor XOR2 (N2599, N2598, N1871);
buf BUF1 (N2600, N2595);
and AND3 (N2601, N2573, N433, N364);
nor NOR3 (N2602, N2555, N530, N1842);
nand NAND4 (N2603, N2602, N2338, N1856, N443);
nand NAND2 (N2604, N2601, N1708);
or OR2 (N2605, N2599, N9);
xor XOR2 (N2606, N2581, N378);
not NOT1 (N2607, N2604);
buf BUF1 (N2608, N2597);
buf BUF1 (N2609, N2596);
not NOT1 (N2610, N2594);
buf BUF1 (N2611, N2606);
nand NAND3 (N2612, N2605, N1950, N2454);
nand NAND4 (N2613, N2607, N1679, N2542, N897);
nor NOR3 (N2614, N2554, N604, N794);
nor NOR3 (N2615, N2603, N18, N1952);
or OR2 (N2616, N2612, N709);
nand NAND3 (N2617, N2610, N168, N2290);
buf BUF1 (N2618, N2616);
and AND2 (N2619, N2608, N310);
and AND2 (N2620, N2614, N1152);
or OR4 (N2621, N2615, N287, N1849, N1712);
not NOT1 (N2622, N2589);
or OR4 (N2623, N2609, N1184, N2451, N667);
nand NAND2 (N2624, N2619, N714);
not NOT1 (N2625, N2623);
xor XOR2 (N2626, N2622, N2612);
or OR2 (N2627, N2613, N2172);
buf BUF1 (N2628, N2600);
and AND4 (N2629, N2624, N1332, N1752, N1444);
not NOT1 (N2630, N2621);
buf BUF1 (N2631, N2626);
nor NOR3 (N2632, N2629, N2288, N2391);
or OR2 (N2633, N2617, N1523);
nor NOR4 (N2634, N2625, N2245, N2242, N1236);
or OR4 (N2635, N2620, N2225, N959, N167);
not NOT1 (N2636, N2630);
nor NOR3 (N2637, N2634, N1776, N2307);
xor XOR2 (N2638, N2611, N2369);
buf BUF1 (N2639, N2636);
nand NAND2 (N2640, N2627, N1709);
nand NAND2 (N2641, N2618, N1997);
nor NOR2 (N2642, N2635, N1760);
nand NAND3 (N2643, N2639, N185, N2241);
or OR2 (N2644, N2631, N1149);
and AND4 (N2645, N2632, N870, N231, N1879);
not NOT1 (N2646, N2628);
and AND3 (N2647, N2641, N2447, N1247);
and AND2 (N2648, N2647, N1884);
nor NOR4 (N2649, N2642, N1228, N2094, N2471);
or OR4 (N2650, N2648, N2643, N1287, N2503);
or OR2 (N2651, N1349, N2330);
or OR4 (N2652, N2644, N1580, N800, N945);
and AND4 (N2653, N2651, N2337, N2108, N2622);
not NOT1 (N2654, N2638);
nor NOR3 (N2655, N2640, N1086, N186);
or OR4 (N2656, N2649, N504, N833, N1606);
or OR4 (N2657, N2633, N611, N1141, N1936);
xor XOR2 (N2658, N2657, N408);
and AND4 (N2659, N2650, N1810, N247, N1094);
or OR2 (N2660, N2656, N1775);
or OR2 (N2661, N2654, N948);
or OR4 (N2662, N2653, N1688, N2554, N444);
not NOT1 (N2663, N2659);
xor XOR2 (N2664, N2658, N1476);
buf BUF1 (N2665, N2645);
nand NAND2 (N2666, N2663, N1368);
and AND4 (N2667, N2664, N1873, N377, N2621);
buf BUF1 (N2668, N2655);
xor XOR2 (N2669, N2667, N2594);
or OR4 (N2670, N2669, N706, N513, N869);
and AND4 (N2671, N2652, N288, N1580, N2649);
or OR2 (N2672, N2661, N2407);
xor XOR2 (N2673, N2665, N697);
or OR4 (N2674, N2672, N2351, N1965, N1710);
buf BUF1 (N2675, N2670);
nor NOR4 (N2676, N2675, N2172, N342, N1416);
and AND2 (N2677, N2662, N1224);
xor XOR2 (N2678, N2666, N2132);
or OR4 (N2679, N2677, N857, N720, N997);
buf BUF1 (N2680, N2668);
xor XOR2 (N2681, N2646, N1721);
or OR2 (N2682, N2678, N1671);
xor XOR2 (N2683, N2660, N1460);
or OR3 (N2684, N2676, N777, N1408);
buf BUF1 (N2685, N2674);
buf BUF1 (N2686, N2683);
not NOT1 (N2687, N2686);
or OR2 (N2688, N2685, N696);
nor NOR3 (N2689, N2671, N87, N813);
and AND4 (N2690, N2688, N53, N375, N2458);
xor XOR2 (N2691, N2673, N713);
xor XOR2 (N2692, N2687, N2588);
not NOT1 (N2693, N2680);
buf BUF1 (N2694, N2692);
and AND2 (N2695, N2689, N2352);
nor NOR4 (N2696, N2690, N2176, N897, N2205);
and AND4 (N2697, N2681, N647, N561, N1058);
and AND4 (N2698, N2696, N433, N1451, N1272);
not NOT1 (N2699, N2697);
nand NAND4 (N2700, N2694, N962, N2520, N763);
not NOT1 (N2701, N2693);
xor XOR2 (N2702, N2682, N1397);
and AND4 (N2703, N2701, N1319, N594, N591);
and AND2 (N2704, N2700, N399);
or OR2 (N2705, N2702, N2671);
nor NOR2 (N2706, N2695, N548);
nand NAND3 (N2707, N2637, N2277, N1944);
xor XOR2 (N2708, N2679, N2340);
or OR3 (N2709, N2707, N660, N1770);
not NOT1 (N2710, N2704);
nor NOR3 (N2711, N2691, N171, N10);
and AND2 (N2712, N2711, N975);
nor NOR3 (N2713, N2710, N433, N2630);
not NOT1 (N2714, N2703);
buf BUF1 (N2715, N2714);
buf BUF1 (N2716, N2713);
nor NOR3 (N2717, N2709, N443, N540);
not NOT1 (N2718, N2712);
xor XOR2 (N2719, N2715, N1964);
buf BUF1 (N2720, N2699);
nand NAND4 (N2721, N2719, N1314, N1613, N1502);
buf BUF1 (N2722, N2716);
and AND4 (N2723, N2721, N1900, N2628, N241);
xor XOR2 (N2724, N2722, N2483);
xor XOR2 (N2725, N2708, N1206);
nand NAND2 (N2726, N2723, N808);
or OR4 (N2727, N2725, N837, N652, N2270);
xor XOR2 (N2728, N2724, N2618);
not NOT1 (N2729, N2717);
nor NOR3 (N2730, N2705, N375, N1528);
nor NOR4 (N2731, N2684, N873, N939, N1094);
or OR2 (N2732, N2718, N2325);
buf BUF1 (N2733, N2728);
buf BUF1 (N2734, N2729);
not NOT1 (N2735, N2698);
xor XOR2 (N2736, N2720, N669);
buf BUF1 (N2737, N2706);
buf BUF1 (N2738, N2730);
or OR3 (N2739, N2726, N1543, N2105);
xor XOR2 (N2740, N2736, N2616);
nor NOR2 (N2741, N2740, N501);
or OR3 (N2742, N2741, N1438, N2025);
buf BUF1 (N2743, N2735);
nand NAND4 (N2744, N2734, N2404, N449, N613);
xor XOR2 (N2745, N2731, N2533);
buf BUF1 (N2746, N2742);
or OR4 (N2747, N2739, N247, N2414, N659);
nor NOR3 (N2748, N2743, N81, N2356);
buf BUF1 (N2749, N2744);
buf BUF1 (N2750, N2727);
not NOT1 (N2751, N2745);
nand NAND4 (N2752, N2751, N841, N557, N2023);
buf BUF1 (N2753, N2750);
nand NAND3 (N2754, N2748, N771, N1514);
or OR3 (N2755, N2747, N1924, N486);
nor NOR4 (N2756, N2754, N1278, N2209, N1520);
and AND4 (N2757, N2753, N1138, N2210, N265);
not NOT1 (N2758, N2732);
xor XOR2 (N2759, N2755, N1718);
buf BUF1 (N2760, N2733);
buf BUF1 (N2761, N2746);
buf BUF1 (N2762, N2761);
buf BUF1 (N2763, N2752);
buf BUF1 (N2764, N2759);
xor XOR2 (N2765, N2762, N2035);
nand NAND3 (N2766, N2765, N1356, N654);
and AND2 (N2767, N2757, N1426);
or OR3 (N2768, N2760, N2424, N507);
nor NOR4 (N2769, N2738, N536, N2096, N978);
xor XOR2 (N2770, N2758, N2198);
not NOT1 (N2771, N2764);
and AND3 (N2772, N2756, N2137, N2363);
or OR2 (N2773, N2737, N396);
or OR3 (N2774, N2749, N2131, N1012);
xor XOR2 (N2775, N2774, N463);
nand NAND2 (N2776, N2769, N2069);
nand NAND4 (N2777, N2771, N532, N678, N431);
nand NAND4 (N2778, N2767, N318, N2159, N178);
not NOT1 (N2779, N2773);
and AND2 (N2780, N2768, N1205);
and AND4 (N2781, N2777, N1722, N2158, N1843);
nand NAND3 (N2782, N2778, N95, N1834);
not NOT1 (N2783, N2763);
or OR3 (N2784, N2776, N659, N141);
xor XOR2 (N2785, N2784, N1424);
nor NOR2 (N2786, N2770, N2298);
nor NOR2 (N2787, N2766, N743);
xor XOR2 (N2788, N2775, N527);
nor NOR2 (N2789, N2783, N1507);
xor XOR2 (N2790, N2789, N1334);
nand NAND2 (N2791, N2790, N820);
xor XOR2 (N2792, N2772, N967);
not NOT1 (N2793, N2779);
xor XOR2 (N2794, N2788, N191);
nor NOR4 (N2795, N2780, N1708, N1081, N552);
or OR2 (N2796, N2794, N705);
xor XOR2 (N2797, N2781, N1189);
not NOT1 (N2798, N2786);
buf BUF1 (N2799, N2797);
xor XOR2 (N2800, N2782, N965);
buf BUF1 (N2801, N2791);
or OR3 (N2802, N2796, N1264, N332);
not NOT1 (N2803, N2802);
nand NAND2 (N2804, N2785, N2353);
or OR3 (N2805, N2787, N2717, N1780);
or OR2 (N2806, N2805, N2291);
not NOT1 (N2807, N2799);
xor XOR2 (N2808, N2800, N1790);
nand NAND3 (N2809, N2804, N653, N2348);
and AND4 (N2810, N2803, N2767, N1115, N785);
nand NAND3 (N2811, N2801, N839, N2183);
or OR4 (N2812, N2793, N2190, N633, N2223);
nand NAND3 (N2813, N2795, N2613, N2808);
or OR4 (N2814, N90, N1206, N177, N1958);
xor XOR2 (N2815, N2807, N1984);
not NOT1 (N2816, N2806);
nand NAND3 (N2817, N2813, N2382, N332);
nand NAND3 (N2818, N2798, N397, N572);
buf BUF1 (N2819, N2817);
not NOT1 (N2820, N2816);
xor XOR2 (N2821, N2811, N756);
and AND2 (N2822, N2821, N2819);
and AND4 (N2823, N1668, N1414, N2234, N6);
not NOT1 (N2824, N2818);
and AND2 (N2825, N2815, N2622);
nand NAND4 (N2826, N2823, N828, N1510, N1066);
and AND3 (N2827, N2792, N329, N2615);
xor XOR2 (N2828, N2826, N1103);
or OR2 (N2829, N2825, N534);
nand NAND3 (N2830, N2812, N294, N1063);
buf BUF1 (N2831, N2822);
nand NAND4 (N2832, N2830, N1877, N2070, N2156);
xor XOR2 (N2833, N2824, N2041);
nand NAND3 (N2834, N2832, N443, N877);
xor XOR2 (N2835, N2814, N154);
nand NAND2 (N2836, N2833, N71);
not NOT1 (N2837, N2828);
and AND4 (N2838, N2835, N973, N2780, N1703);
nor NOR3 (N2839, N2837, N913, N237);
not NOT1 (N2840, N2809);
and AND3 (N2841, N2810, N475, N1962);
nor NOR3 (N2842, N2836, N1413, N1617);
nand NAND4 (N2843, N2838, N802, N1834, N2481);
nor NOR3 (N2844, N2840, N1252, N1663);
nor NOR4 (N2845, N2834, N2554, N2006, N1572);
buf BUF1 (N2846, N2844);
nand NAND2 (N2847, N2841, N718);
not NOT1 (N2848, N2839);
buf BUF1 (N2849, N2827);
buf BUF1 (N2850, N2820);
and AND2 (N2851, N2846, N2104);
not NOT1 (N2852, N2850);
not NOT1 (N2853, N2831);
or OR3 (N2854, N2847, N1152, N1140);
and AND3 (N2855, N2829, N2761, N1174);
xor XOR2 (N2856, N2843, N209);
buf BUF1 (N2857, N2856);
nand NAND4 (N2858, N2852, N1344, N373, N1931);
nor NOR4 (N2859, N2848, N1771, N331, N673);
and AND3 (N2860, N2845, N2716, N2045);
buf BUF1 (N2861, N2842);
or OR3 (N2862, N2849, N1049, N2833);
and AND3 (N2863, N2861, N2109, N1970);
nand NAND2 (N2864, N2851, N1198);
not NOT1 (N2865, N2864);
nand NAND4 (N2866, N2857, N128, N1864, N586);
nor NOR4 (N2867, N2866, N2317, N574, N2300);
nand NAND2 (N2868, N2865, N2706);
not NOT1 (N2869, N2863);
xor XOR2 (N2870, N2855, N1629);
and AND2 (N2871, N2870, N775);
nor NOR3 (N2872, N2871, N765, N1534);
nand NAND4 (N2873, N2868, N2516, N1036, N653);
nand NAND2 (N2874, N2853, N544);
xor XOR2 (N2875, N2867, N2341);
not NOT1 (N2876, N2858);
nor NOR2 (N2877, N2854, N118);
xor XOR2 (N2878, N2869, N1886);
xor XOR2 (N2879, N2872, N1869);
buf BUF1 (N2880, N2874);
nand NAND2 (N2881, N2878, N648);
or OR4 (N2882, N2875, N676, N2817, N1324);
not NOT1 (N2883, N2882);
nor NOR3 (N2884, N2862, N1305, N2350);
buf BUF1 (N2885, N2876);
nand NAND2 (N2886, N2859, N2606);
nor NOR4 (N2887, N2885, N249, N1409, N1119);
and AND2 (N2888, N2880, N2833);
and AND4 (N2889, N2881, N2687, N2471, N1229);
xor XOR2 (N2890, N2888, N915);
xor XOR2 (N2891, N2884, N2214);
buf BUF1 (N2892, N2887);
buf BUF1 (N2893, N2860);
nand NAND2 (N2894, N2889, N75);
nand NAND3 (N2895, N2883, N1529, N2318);
not NOT1 (N2896, N2873);
and AND3 (N2897, N2891, N2639, N2473);
and AND3 (N2898, N2886, N973, N285);
or OR4 (N2899, N2892, N2567, N1057, N2728);
or OR4 (N2900, N2895, N2106, N1315, N1341);
buf BUF1 (N2901, N2898);
not NOT1 (N2902, N2899);
nor NOR2 (N2903, N2902, N984);
nand NAND2 (N2904, N2879, N1994);
or OR4 (N2905, N2877, N517, N1370, N1199);
and AND4 (N2906, N2896, N2441, N74, N2184);
nor NOR3 (N2907, N2893, N313, N441);
buf BUF1 (N2908, N2890);
not NOT1 (N2909, N2905);
buf BUF1 (N2910, N2901);
or OR2 (N2911, N2907, N297);
not NOT1 (N2912, N2903);
or OR4 (N2913, N2906, N1118, N956, N514);
and AND4 (N2914, N2913, N2040, N2303, N1220);
and AND4 (N2915, N2897, N973, N922, N244);
not NOT1 (N2916, N2915);
nand NAND2 (N2917, N2916, N1955);
xor XOR2 (N2918, N2911, N1890);
nand NAND3 (N2919, N2914, N1752, N967);
buf BUF1 (N2920, N2918);
nor NOR3 (N2921, N2917, N643, N1196);
buf BUF1 (N2922, N2912);
nor NOR2 (N2923, N2900, N2139);
nand NAND2 (N2924, N2919, N855);
or OR4 (N2925, N2920, N2740, N546, N2036);
nor NOR2 (N2926, N2925, N584);
and AND3 (N2927, N2904, N2589, N338);
and AND4 (N2928, N2909, N85, N2209, N438);
or OR3 (N2929, N2924, N1303, N1734);
or OR2 (N2930, N2923, N1575);
nand NAND4 (N2931, N2922, N1727, N1054, N1286);
and AND2 (N2932, N2921, N1424);
buf BUF1 (N2933, N2929);
and AND2 (N2934, N2910, N1327);
nor NOR3 (N2935, N2931, N631, N1762);
nand NAND4 (N2936, N2894, N778, N841, N1127);
xor XOR2 (N2937, N2930, N600);
not NOT1 (N2938, N2934);
xor XOR2 (N2939, N2928, N1757);
nor NOR2 (N2940, N2938, N470);
or OR3 (N2941, N2933, N1260, N273);
or OR3 (N2942, N2937, N780, N2649);
and AND2 (N2943, N2926, N1279);
and AND3 (N2944, N2939, N2912, N201);
not NOT1 (N2945, N2936);
nor NOR4 (N2946, N2944, N2513, N1159, N1334);
or OR3 (N2947, N2946, N193, N2174);
nor NOR4 (N2948, N2943, N2899, N2004, N1075);
nor NOR3 (N2949, N2932, N2077, N1820);
nand NAND2 (N2950, N2942, N1490);
nand NAND2 (N2951, N2927, N169);
or OR2 (N2952, N2940, N2566);
and AND2 (N2953, N2945, N1307);
nor NOR3 (N2954, N2953, N2021, N907);
nor NOR2 (N2955, N2951, N2656);
xor XOR2 (N2956, N2947, N752);
nor NOR4 (N2957, N2950, N1718, N2759, N1711);
xor XOR2 (N2958, N2952, N220);
nand NAND2 (N2959, N2954, N759);
or OR3 (N2960, N2908, N1035, N2793);
not NOT1 (N2961, N2948);
nand NAND3 (N2962, N2949, N1068, N628);
nor NOR4 (N2963, N2959, N1571, N56, N1184);
xor XOR2 (N2964, N2962, N177);
or OR4 (N2965, N2958, N909, N1557, N211);
not NOT1 (N2966, N2955);
buf BUF1 (N2967, N2966);
and AND2 (N2968, N2957, N1751);
not NOT1 (N2969, N2968);
xor XOR2 (N2970, N2963, N1773);
and AND2 (N2971, N2970, N1400);
buf BUF1 (N2972, N2960);
buf BUF1 (N2973, N2941);
or OR3 (N2974, N2969, N1351, N2097);
and AND2 (N2975, N2965, N2533);
nor NOR2 (N2976, N2961, N925);
not NOT1 (N2977, N2976);
not NOT1 (N2978, N2956);
nor NOR4 (N2979, N2971, N1686, N629, N558);
nor NOR2 (N2980, N2964, N1336);
or OR4 (N2981, N2978, N1171, N2523, N2228);
not NOT1 (N2982, N2975);
buf BUF1 (N2983, N2982);
nor NOR3 (N2984, N2974, N343, N196);
and AND3 (N2985, N2983, N624, N2424);
nor NOR2 (N2986, N2984, N2943);
nor NOR4 (N2987, N2967, N2654, N2624, N1640);
and AND2 (N2988, N2987, N193);
or OR2 (N2989, N2986, N878);
and AND2 (N2990, N2935, N1542);
and AND4 (N2991, N2973, N2068, N1764, N233);
nor NOR2 (N2992, N2988, N2834);
xor XOR2 (N2993, N2980, N429);
nand NAND3 (N2994, N2989, N2000, N2370);
nand NAND2 (N2995, N2992, N632);
or OR4 (N2996, N2993, N2016, N322, N304);
not NOT1 (N2997, N2995);
and AND2 (N2998, N2981, N791);
not NOT1 (N2999, N2994);
not NOT1 (N3000, N2972);
buf BUF1 (N3001, N2999);
nand NAND2 (N3002, N2985, N1526);
xor XOR2 (N3003, N2996, N801);
nand NAND3 (N3004, N2990, N1222, N2297);
or OR2 (N3005, N2979, N2148);
or OR2 (N3006, N3003, N2693);
not NOT1 (N3007, N2997);
xor XOR2 (N3008, N3006, N2523);
buf BUF1 (N3009, N2991);
nand NAND2 (N3010, N3008, N367);
buf BUF1 (N3011, N3000);
buf BUF1 (N3012, N3009);
and AND3 (N3013, N2998, N818, N2350);
nand NAND3 (N3014, N3012, N1834, N1908);
not NOT1 (N3015, N3002);
and AND4 (N3016, N3001, N2864, N2069, N1354);
buf BUF1 (N3017, N3014);
not NOT1 (N3018, N2977);
not NOT1 (N3019, N3015);
or OR3 (N3020, N3013, N2721, N1943);
or OR2 (N3021, N3010, N93);
not NOT1 (N3022, N3005);
nor NOR2 (N3023, N3004, N1858);
xor XOR2 (N3024, N3023, N754);
not NOT1 (N3025, N3016);
buf BUF1 (N3026, N3007);
nor NOR2 (N3027, N3020, N3016);
buf BUF1 (N3028, N3019);
not NOT1 (N3029, N3026);
buf BUF1 (N3030, N3028);
buf BUF1 (N3031, N3022);
buf BUF1 (N3032, N3018);
nor NOR2 (N3033, N3030, N2590);
or OR4 (N3034, N3025, N332, N2669, N777);
xor XOR2 (N3035, N3031, N1840);
nor NOR4 (N3036, N3021, N871, N2998, N2240);
and AND3 (N3037, N3034, N602, N1408);
not NOT1 (N3038, N3029);
xor XOR2 (N3039, N3017, N894);
nor NOR4 (N3040, N3032, N2588, N216, N1977);
xor XOR2 (N3041, N3011, N2006);
buf BUF1 (N3042, N3037);
not NOT1 (N3043, N3039);
nand NAND3 (N3044, N3041, N2631, N292);
not NOT1 (N3045, N3035);
nand NAND2 (N3046, N3044, N149);
nand NAND3 (N3047, N3027, N1491, N2350);
or OR4 (N3048, N3042, N828, N1070, N2863);
and AND3 (N3049, N3045, N422, N1264);
nand NAND3 (N3050, N3049, N2373, N2711);
buf BUF1 (N3051, N3046);
nor NOR2 (N3052, N3038, N211);
buf BUF1 (N3053, N3040);
or OR2 (N3054, N3048, N303);
nor NOR2 (N3055, N3047, N1327);
nand NAND2 (N3056, N3053, N148);
and AND3 (N3057, N3051, N878, N412);
nor NOR2 (N3058, N3054, N752);
and AND3 (N3059, N3057, N186, N2677);
not NOT1 (N3060, N3052);
nor NOR2 (N3061, N3024, N972);
buf BUF1 (N3062, N3061);
not NOT1 (N3063, N3033);
nand NAND2 (N3064, N3060, N79);
nand NAND4 (N3065, N3055, N2200, N1973, N2324);
or OR3 (N3066, N3036, N3010, N2259);
nor NOR4 (N3067, N3064, N2519, N148, N499);
buf BUF1 (N3068, N3059);
buf BUF1 (N3069, N3067);
not NOT1 (N3070, N3063);
xor XOR2 (N3071, N3066, N829);
nand NAND4 (N3072, N3043, N1462, N2995, N2308);
nand NAND3 (N3073, N3062, N2566, N1108);
xor XOR2 (N3074, N3058, N1843);
not NOT1 (N3075, N3069);
nand NAND3 (N3076, N3056, N1738, N2507);
xor XOR2 (N3077, N3072, N2836);
or OR4 (N3078, N3076, N2133, N1079, N2186);
nor NOR3 (N3079, N3078, N403, N1748);
not NOT1 (N3080, N3075);
nand NAND4 (N3081, N3070, N1558, N1241, N523);
or OR2 (N3082, N3073, N1224);
or OR2 (N3083, N3074, N3001);
not NOT1 (N3084, N3081);
nor NOR4 (N3085, N3080, N1741, N2317, N2677);
not NOT1 (N3086, N3079);
nand NAND4 (N3087, N3068, N2391, N2220, N1172);
nand NAND2 (N3088, N3087, N2027);
not NOT1 (N3089, N3077);
nand NAND4 (N3090, N3086, N1644, N805, N1885);
not NOT1 (N3091, N3089);
not NOT1 (N3092, N3084);
nand NAND2 (N3093, N3085, N2725);
nand NAND4 (N3094, N3050, N308, N2353, N1442);
not NOT1 (N3095, N3083);
and AND2 (N3096, N3082, N1456);
or OR3 (N3097, N3065, N3034, N2729);
and AND3 (N3098, N3097, N1420, N90);
or OR3 (N3099, N3092, N1824, N2259);
nand NAND4 (N3100, N3091, N661, N368, N2789);
xor XOR2 (N3101, N3098, N2533);
or OR2 (N3102, N3093, N1913);
and AND2 (N3103, N3099, N2860);
nor NOR2 (N3104, N3102, N255);
not NOT1 (N3105, N3100);
or OR4 (N3106, N3071, N2167, N2787, N829);
not NOT1 (N3107, N3088);
buf BUF1 (N3108, N3105);
nor NOR2 (N3109, N3108, N720);
or OR2 (N3110, N3101, N767);
buf BUF1 (N3111, N3104);
xor XOR2 (N3112, N3095, N607);
xor XOR2 (N3113, N3103, N640);
or OR2 (N3114, N3107, N2208);
xor XOR2 (N3115, N3111, N2605);
nor NOR3 (N3116, N3096, N2526, N408);
nor NOR4 (N3117, N3094, N408, N1137, N1893);
nand NAND4 (N3118, N3112, N1710, N1815, N2079);
nand NAND4 (N3119, N3118, N2934, N2330, N2537);
xor XOR2 (N3120, N3115, N998);
and AND4 (N3121, N3114, N1269, N2716, N484);
nand NAND2 (N3122, N3120, N2638);
nor NOR4 (N3123, N3117, N694, N2375, N1902);
xor XOR2 (N3124, N3121, N2240);
nor NOR4 (N3125, N3119, N2424, N19, N302);
nand NAND4 (N3126, N3090, N1306, N2172, N1253);
nand NAND3 (N3127, N3123, N1271, N434);
or OR2 (N3128, N3126, N2278);
not NOT1 (N3129, N3124);
nor NOR3 (N3130, N3110, N2052, N2406);
or OR3 (N3131, N3122, N1293, N2394);
xor XOR2 (N3132, N3128, N270);
nand NAND2 (N3133, N3130, N1881);
and AND3 (N3134, N3132, N2986, N1396);
and AND2 (N3135, N3109, N979);
xor XOR2 (N3136, N3125, N2556);
or OR3 (N3137, N3133, N1313, N200);
nor NOR2 (N3138, N3137, N769);
or OR4 (N3139, N3136, N2060, N1058, N190);
xor XOR2 (N3140, N3113, N2036);
buf BUF1 (N3141, N3135);
and AND4 (N3142, N3129, N1004, N2565, N2058);
not NOT1 (N3143, N3134);
buf BUF1 (N3144, N3116);
nand NAND3 (N3145, N3141, N866, N2121);
nand NAND3 (N3146, N3144, N3009, N1895);
or OR3 (N3147, N3139, N959, N932);
xor XOR2 (N3148, N3138, N1056);
nand NAND3 (N3149, N3106, N530, N2687);
nand NAND4 (N3150, N3127, N1124, N1463, N92);
xor XOR2 (N3151, N3143, N2661);
nand NAND4 (N3152, N3147, N842, N1496, N2372);
xor XOR2 (N3153, N3142, N1073);
nor NOR3 (N3154, N3145, N117, N1821);
xor XOR2 (N3155, N3152, N3152);
nor NOR4 (N3156, N3146, N3020, N1422, N3013);
not NOT1 (N3157, N3156);
or OR3 (N3158, N3140, N543, N3019);
nand NAND2 (N3159, N3150, N1739);
buf BUF1 (N3160, N3149);
or OR2 (N3161, N3158, N284);
or OR4 (N3162, N3151, N1844, N929, N1211);
or OR4 (N3163, N3154, N2926, N3052, N2123);
nand NAND4 (N3164, N3159, N1206, N1938, N315);
nor NOR2 (N3165, N3153, N80);
nand NAND2 (N3166, N3164, N1506);
and AND3 (N3167, N3161, N689, N440);
xor XOR2 (N3168, N3167, N2031);
nor NOR3 (N3169, N3168, N1913, N2886);
not NOT1 (N3170, N3155);
nor NOR4 (N3171, N3131, N615, N2029, N1351);
nand NAND3 (N3172, N3162, N2858, N1004);
xor XOR2 (N3173, N3157, N449);
nor NOR4 (N3174, N3166, N212, N1933, N110);
nor NOR3 (N3175, N3165, N694, N317);
nand NAND2 (N3176, N3171, N2715);
nor NOR3 (N3177, N3176, N810, N1815);
or OR3 (N3178, N3175, N1828, N854);
nand NAND3 (N3179, N3148, N678, N1375);
nor NOR4 (N3180, N3170, N2113, N2310, N2560);
buf BUF1 (N3181, N3174);
not NOT1 (N3182, N3163);
nand NAND3 (N3183, N3181, N857, N1099);
xor XOR2 (N3184, N3172, N383);
nor NOR3 (N3185, N3178, N2236, N1891);
buf BUF1 (N3186, N3173);
nand NAND4 (N3187, N3180, N3028, N1188, N2964);
not NOT1 (N3188, N3183);
or OR2 (N3189, N3184, N2224);
nand NAND3 (N3190, N3185, N2962, N1263);
nand NAND4 (N3191, N3190, N1415, N777, N2237);
not NOT1 (N3192, N3182);
xor XOR2 (N3193, N3187, N455);
xor XOR2 (N3194, N3188, N764);
xor XOR2 (N3195, N3191, N3008);
buf BUF1 (N3196, N3194);
not NOT1 (N3197, N3193);
nor NOR2 (N3198, N3192, N2205);
not NOT1 (N3199, N3195);
nand NAND4 (N3200, N3186, N2853, N152, N122);
nor NOR2 (N3201, N3200, N2194);
buf BUF1 (N3202, N3199);
or OR2 (N3203, N3198, N1188);
nor NOR3 (N3204, N3203, N390, N1829);
or OR2 (N3205, N3177, N691);
not NOT1 (N3206, N3205);
or OR2 (N3207, N3179, N831);
buf BUF1 (N3208, N3207);
buf BUF1 (N3209, N3189);
buf BUF1 (N3210, N3206);
not NOT1 (N3211, N3201);
nor NOR2 (N3212, N3204, N1614);
not NOT1 (N3213, N3208);
xor XOR2 (N3214, N3213, N248);
and AND3 (N3215, N3169, N1638, N2794);
or OR3 (N3216, N3196, N660, N2927);
nand NAND3 (N3217, N3216, N251, N1807);
not NOT1 (N3218, N3160);
and AND4 (N3219, N3214, N638, N361, N2548);
endmodule