// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N209,N206,N201,N205,N208,N200,N210,N204,N192,N211;

nor NOR4 (N12, N3, N1, N6, N4);
nand NAND3 (N13, N9, N12, N11);
not NOT1 (N14, N8);
nor NOR3 (N15, N12, N4, N11);
xor XOR2 (N16, N8, N7);
or OR4 (N17, N8, N8, N6, N8);
nor NOR4 (N18, N14, N8, N5, N15);
nor NOR4 (N19, N17, N13, N10, N17);
nand NAND2 (N20, N1, N12);
and AND3 (N21, N12, N5, N4);
nor NOR4 (N22, N20, N20, N15, N17);
nor NOR4 (N23, N8, N4, N15, N11);
nand NAND2 (N24, N21, N11);
nor NOR3 (N25, N10, N20, N11);
xor XOR2 (N26, N16, N24);
buf BUF1 (N27, N26);
not NOT1 (N28, N21);
not NOT1 (N29, N20);
nand NAND2 (N30, N1, N2);
nor NOR4 (N31, N22, N13, N6, N9);
or OR2 (N32, N17, N14);
and AND4 (N33, N31, N10, N13, N27);
nor NOR4 (N34, N26, N2, N7, N19);
not NOT1 (N35, N15);
and AND4 (N36, N25, N32, N18, N34);
nand NAND4 (N37, N26, N19, N31, N33);
xor XOR2 (N38, N3, N14);
buf BUF1 (N39, N7);
buf BUF1 (N40, N3);
and AND2 (N41, N37, N36);
buf BUF1 (N42, N40);
and AND4 (N43, N15, N17, N16, N16);
nor NOR3 (N44, N23, N1, N18);
nor NOR2 (N45, N44, N36);
buf BUF1 (N46, N28);
or OR4 (N47, N35, N27, N8, N16);
xor XOR2 (N48, N29, N46);
or OR3 (N49, N47, N12, N26);
buf BUF1 (N50, N20);
and AND4 (N51, N43, N23, N31, N40);
nand NAND2 (N52, N30, N38);
buf BUF1 (N53, N23);
buf BUF1 (N54, N53);
xor XOR2 (N55, N48, N21);
nor NOR3 (N56, N41, N24, N33);
and AND2 (N57, N56, N25);
buf BUF1 (N58, N51);
nand NAND4 (N59, N49, N25, N41, N43);
not NOT1 (N60, N45);
nand NAND2 (N61, N59, N10);
buf BUF1 (N62, N39);
not NOT1 (N63, N58);
nor NOR3 (N64, N62, N29, N3);
buf BUF1 (N65, N50);
and AND2 (N66, N65, N31);
nand NAND2 (N67, N55, N39);
nor NOR4 (N68, N54, N30, N41, N46);
nor NOR3 (N69, N63, N47, N2);
nand NAND3 (N70, N52, N39, N26);
nor NOR4 (N71, N68, N39, N46, N66);
not NOT1 (N72, N53);
xor XOR2 (N73, N69, N15);
xor XOR2 (N74, N42, N60);
and AND2 (N75, N64, N64);
nand NAND2 (N76, N65, N36);
or OR2 (N77, N73, N50);
nand NAND4 (N78, N57, N5, N76, N32);
not NOT1 (N79, N49);
and AND2 (N80, N78, N5);
nor NOR2 (N81, N80, N16);
not NOT1 (N82, N72);
nand NAND4 (N83, N77, N33, N17, N19);
or OR3 (N84, N61, N4, N79);
and AND4 (N85, N27, N61, N71, N23);
buf BUF1 (N86, N21);
nor NOR3 (N87, N84, N49, N11);
and AND4 (N88, N67, N20, N43, N79);
or OR4 (N89, N88, N84, N37, N74);
buf BUF1 (N90, N65);
not NOT1 (N91, N81);
not NOT1 (N92, N83);
nand NAND3 (N93, N85, N69, N91);
nor NOR2 (N94, N51, N30);
nand NAND4 (N95, N82, N75, N51, N84);
nand NAND2 (N96, N82, N46);
or OR4 (N97, N87, N57, N3, N48);
or OR2 (N98, N94, N41);
and AND4 (N99, N89, N4, N27, N48);
and AND4 (N100, N99, N95, N45, N46);
not NOT1 (N101, N53);
nor NOR4 (N102, N96, N40, N37, N32);
and AND4 (N103, N101, N64, N102, N42);
buf BUF1 (N104, N52);
xor XOR2 (N105, N86, N52);
or OR3 (N106, N90, N72, N14);
nand NAND2 (N107, N92, N1);
or OR2 (N108, N97, N40);
not NOT1 (N109, N93);
and AND4 (N110, N108, N46, N34, N47);
nand NAND3 (N111, N105, N96, N21);
and AND4 (N112, N98, N35, N9, N11);
or OR3 (N113, N100, N35, N102);
nand NAND2 (N114, N104, N63);
xor XOR2 (N115, N114, N24);
xor XOR2 (N116, N112, N24);
nand NAND2 (N117, N110, N116);
nor NOR4 (N118, N33, N30, N100, N32);
nand NAND2 (N119, N103, N37);
xor XOR2 (N120, N106, N116);
buf BUF1 (N121, N115);
nor NOR3 (N122, N121, N22, N67);
and AND3 (N123, N118, N2, N17);
nand NAND4 (N124, N109, N10, N97, N39);
nor NOR3 (N125, N70, N16, N81);
buf BUF1 (N126, N107);
nand NAND2 (N127, N125, N119);
not NOT1 (N128, N11);
buf BUF1 (N129, N111);
buf BUF1 (N130, N120);
not NOT1 (N131, N127);
nor NOR3 (N132, N117, N70, N41);
not NOT1 (N133, N131);
xor XOR2 (N134, N132, N102);
and AND3 (N135, N134, N87, N133);
nor NOR4 (N136, N109, N41, N33, N59);
and AND3 (N137, N124, N11, N93);
or OR4 (N138, N137, N102, N73, N82);
and AND3 (N139, N138, N116, N38);
nand NAND2 (N140, N128, N49);
and AND4 (N141, N136, N27, N110, N50);
nor NOR2 (N142, N130, N64);
and AND4 (N143, N122, N56, N38, N127);
xor XOR2 (N144, N142, N6);
nand NAND2 (N145, N139, N84);
buf BUF1 (N146, N143);
not NOT1 (N147, N146);
and AND2 (N148, N147, N118);
or OR4 (N149, N148, N58, N144, N106);
nand NAND4 (N150, N125, N115, N74, N1);
nand NAND3 (N151, N129, N93, N105);
buf BUF1 (N152, N140);
not NOT1 (N153, N149);
nand NAND3 (N154, N153, N119, N72);
or OR2 (N155, N154, N82);
nand NAND3 (N156, N152, N4, N67);
xor XOR2 (N157, N156, N50);
and AND3 (N158, N155, N99, N130);
and AND2 (N159, N123, N102);
or OR2 (N160, N145, N78);
nand NAND2 (N161, N160, N66);
or OR4 (N162, N113, N120, N82, N57);
xor XOR2 (N163, N161, N70);
buf BUF1 (N164, N162);
buf BUF1 (N165, N159);
nor NOR2 (N166, N165, N5);
nor NOR4 (N167, N163, N88, N80, N46);
or OR2 (N168, N151, N30);
xor XOR2 (N169, N168, N158);
xor XOR2 (N170, N133, N156);
nand NAND3 (N171, N150, N48, N121);
buf BUF1 (N172, N135);
and AND4 (N173, N126, N91, N136, N48);
buf BUF1 (N174, N170);
nor NOR2 (N175, N172, N49);
or OR2 (N176, N169, N55);
not NOT1 (N177, N175);
or OR4 (N178, N157, N30, N173, N177);
nand NAND4 (N179, N67, N29, N88, N174);
xor XOR2 (N180, N80, N19);
not NOT1 (N181, N6);
xor XOR2 (N182, N179, N168);
nand NAND3 (N183, N178, N6, N179);
nor NOR2 (N184, N176, N151);
nor NOR2 (N185, N184, N179);
nand NAND2 (N186, N164, N134);
and AND2 (N187, N181, N75);
xor XOR2 (N188, N186, N66);
not NOT1 (N189, N187);
not NOT1 (N190, N180);
and AND3 (N191, N185, N46, N37);
nand NAND3 (N192, N167, N62, N182);
xor XOR2 (N193, N51, N159);
not NOT1 (N194, N141);
not NOT1 (N195, N194);
and AND4 (N196, N190, N23, N144, N61);
xor XOR2 (N197, N183, N93);
nor NOR2 (N198, N171, N27);
xor XOR2 (N199, N198, N14);
not NOT1 (N200, N193);
xor XOR2 (N201, N195, N96);
nand NAND3 (N202, N166, N161, N93);
nand NAND2 (N203, N189, N15);
xor XOR2 (N204, N196, N136);
and AND4 (N205, N197, N153, N88, N125);
buf BUF1 (N206, N191);
and AND2 (N207, N188, N175);
nand NAND2 (N208, N202, N23);
buf BUF1 (N209, N203);
or OR2 (N210, N199, N134);
and AND4 (N211, N207, N33, N33, N182);
endmodule