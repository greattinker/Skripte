// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N112,N114,N116,N115,N110,N117,N113,N118,N119,N120;

or OR4 (N21, N9, N10, N11, N15);
nand NAND3 (N22, N21, N3, N12);
and AND3 (N23, N5, N14, N12);
or OR3 (N24, N22, N7, N14);
buf BUF1 (N25, N4);
nor NOR4 (N26, N19, N7, N23, N25);
xor XOR2 (N27, N3, N5);
not NOT1 (N28, N3);
or OR2 (N29, N24, N20);
not NOT1 (N30, N28);
or OR4 (N31, N8, N22, N27, N22);
buf BUF1 (N32, N13);
xor XOR2 (N33, N7, N13);
and AND2 (N34, N1, N15);
nand NAND4 (N35, N24, N4, N34, N32);
not NOT1 (N36, N13);
or OR4 (N37, N33, N28, N4, N36);
nor NOR4 (N38, N24, N26, N18, N25);
and AND2 (N39, N27, N33);
and AND3 (N40, N29, N5, N17);
xor XOR2 (N41, N29, N17);
xor XOR2 (N42, N21, N30);
not NOT1 (N43, N22);
not NOT1 (N44, N3);
and AND2 (N45, N37, N27);
nor NOR4 (N46, N41, N32, N21, N18);
and AND2 (N47, N44, N33);
not NOT1 (N48, N42);
or OR3 (N49, N40, N33, N1);
nor NOR3 (N50, N48, N38, N24);
or OR3 (N51, N37, N40, N12);
and AND3 (N52, N39, N30, N11);
buf BUF1 (N53, N50);
nor NOR4 (N54, N45, N11, N24, N7);
xor XOR2 (N55, N43, N6);
buf BUF1 (N56, N47);
buf BUF1 (N57, N52);
not NOT1 (N58, N54);
nand NAND4 (N59, N46, N27, N53, N1);
xor XOR2 (N60, N14, N46);
nor NOR2 (N61, N55, N42);
not NOT1 (N62, N35);
buf BUF1 (N63, N59);
not NOT1 (N64, N57);
and AND2 (N65, N60, N27);
not NOT1 (N66, N62);
nor NOR4 (N67, N61, N4, N42, N61);
xor XOR2 (N68, N64, N53);
xor XOR2 (N69, N63, N24);
xor XOR2 (N70, N58, N12);
not NOT1 (N71, N51);
or OR3 (N72, N56, N52, N12);
xor XOR2 (N73, N72, N10);
or OR2 (N74, N69, N55);
nand NAND2 (N75, N65, N63);
and AND2 (N76, N31, N73);
buf BUF1 (N77, N49);
and AND3 (N78, N26, N63, N32);
nand NAND4 (N79, N67, N3, N10, N35);
or OR4 (N80, N68, N73, N42, N9);
xor XOR2 (N81, N71, N6);
not NOT1 (N82, N77);
nand NAND3 (N83, N75, N5, N57);
not NOT1 (N84, N74);
nor NOR3 (N85, N66, N56, N67);
or OR2 (N86, N84, N62);
xor XOR2 (N87, N85, N1);
or OR3 (N88, N79, N85, N62);
nor NOR3 (N89, N70, N52, N33);
nand NAND3 (N90, N86, N65, N29);
or OR2 (N91, N81, N70);
buf BUF1 (N92, N83);
buf BUF1 (N93, N76);
nor NOR3 (N94, N93, N19, N40);
not NOT1 (N95, N94);
not NOT1 (N96, N87);
nor NOR3 (N97, N88, N55, N17);
or OR4 (N98, N97, N27, N97, N63);
xor XOR2 (N99, N95, N85);
and AND4 (N100, N96, N92, N49, N52);
and AND2 (N101, N26, N80);
not NOT1 (N102, N85);
nor NOR3 (N103, N82, N24, N97);
not NOT1 (N104, N102);
nand NAND2 (N105, N103, N20);
and AND3 (N106, N101, N22, N74);
and AND3 (N107, N104, N61, N37);
nand NAND2 (N108, N91, N107);
and AND2 (N109, N108, N27);
buf BUF1 (N110, N105);
nor NOR4 (N111, N25, N53, N80, N25);
and AND3 (N112, N98, N27, N76);
or OR4 (N113, N99, N79, N91, N1);
not NOT1 (N114, N100);
and AND3 (N115, N90, N12, N55);
or OR4 (N116, N78, N24, N106, N107);
xor XOR2 (N117, N61, N12);
or OR4 (N118, N109, N89, N62, N34);
nor NOR3 (N119, N87, N23, N111);
xor XOR2 (N120, N111, N83);
endmodule