// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N715,N709,N710,N714,N717,N701,N718,N716,N713,N719;

and AND3 (N20, N19, N18, N17);
buf BUF1 (N21, N5);
not NOT1 (N22, N14);
and AND3 (N23, N5, N13, N4);
nor NOR4 (N24, N19, N18, N2, N14);
or OR4 (N25, N16, N14, N17, N12);
buf BUF1 (N26, N25);
nand NAND4 (N27, N14, N17, N13, N2);
and AND4 (N28, N24, N1, N22, N24);
or OR4 (N29, N7, N9, N2, N27);
or OR3 (N30, N15, N8, N1);
not NOT1 (N31, N9);
and AND4 (N32, N1, N19, N2, N6);
nand NAND3 (N33, N18, N1, N22);
and AND3 (N34, N23, N14, N4);
or OR4 (N35, N26, N18, N32, N15);
buf BUF1 (N36, N31);
not NOT1 (N37, N15);
buf BUF1 (N38, N37);
not NOT1 (N39, N29);
buf BUF1 (N40, N39);
buf BUF1 (N41, N36);
nor NOR4 (N42, N33, N34, N9, N5);
nor NOR2 (N43, N38, N35);
nor NOR4 (N44, N17, N11, N22, N39);
or OR4 (N45, N13, N40, N25, N13);
not NOT1 (N46, N11);
buf BUF1 (N47, N42);
xor XOR2 (N48, N45, N30);
not NOT1 (N49, N16);
not NOT1 (N50, N46);
nand NAND4 (N51, N47, N36, N15, N31);
not NOT1 (N52, N20);
not NOT1 (N53, N41);
buf BUF1 (N54, N50);
and AND4 (N55, N43, N4, N31, N39);
xor XOR2 (N56, N44, N27);
or OR2 (N57, N56, N47);
not NOT1 (N58, N52);
nand NAND3 (N59, N48, N45, N15);
nand NAND4 (N60, N51, N43, N39, N14);
or OR2 (N61, N58, N19);
or OR4 (N62, N54, N7, N57, N50);
and AND3 (N63, N10, N40, N2);
nor NOR3 (N64, N61, N38, N59);
nor NOR3 (N65, N56, N24, N20);
and AND4 (N66, N64, N50, N49, N5);
not NOT1 (N67, N58);
not NOT1 (N68, N62);
not NOT1 (N69, N55);
or OR4 (N70, N68, N2, N40, N48);
buf BUF1 (N71, N65);
xor XOR2 (N72, N63, N59);
and AND2 (N73, N53, N46);
or OR3 (N74, N71, N57, N4);
nand NAND2 (N75, N72, N10);
buf BUF1 (N76, N60);
nor NOR2 (N77, N74, N19);
or OR3 (N78, N21, N47, N12);
nand NAND3 (N79, N70, N60, N74);
and AND2 (N80, N78, N77);
not NOT1 (N81, N74);
nor NOR4 (N82, N81, N11, N63, N28);
not NOT1 (N83, N27);
buf BUF1 (N84, N80);
xor XOR2 (N85, N83, N71);
buf BUF1 (N86, N69);
or OR3 (N87, N84, N16, N1);
not NOT1 (N88, N76);
nor NOR2 (N89, N88, N59);
nor NOR3 (N90, N87, N7, N45);
nand NAND2 (N91, N90, N52);
xor XOR2 (N92, N82, N58);
or OR2 (N93, N73, N12);
or OR2 (N94, N67, N13);
and AND3 (N95, N75, N9, N32);
not NOT1 (N96, N93);
nor NOR4 (N97, N96, N96, N20, N35);
or OR4 (N98, N66, N96, N57, N57);
and AND4 (N99, N89, N26, N64, N51);
nor NOR2 (N100, N91, N78);
or OR3 (N101, N98, N99, N95);
not NOT1 (N102, N19);
buf BUF1 (N103, N3);
or OR2 (N104, N102, N79);
or OR2 (N105, N39, N58);
and AND4 (N106, N105, N72, N39, N70);
not NOT1 (N107, N100);
nor NOR4 (N108, N92, N62, N86, N55);
and AND2 (N109, N16, N34);
xor XOR2 (N110, N106, N42);
nor NOR2 (N111, N104, N74);
nand NAND3 (N112, N109, N1, N4);
or OR4 (N113, N85, N3, N49, N15);
xor XOR2 (N114, N97, N66);
not NOT1 (N115, N112);
nand NAND4 (N116, N103, N98, N17, N35);
nor NOR2 (N117, N107, N21);
and AND3 (N118, N116, N109, N36);
xor XOR2 (N119, N117, N50);
and AND3 (N120, N108, N113, N85);
xor XOR2 (N121, N33, N104);
or OR2 (N122, N115, N26);
nand NAND3 (N123, N122, N81, N91);
nand NAND3 (N124, N123, N39, N118);
nor NOR2 (N125, N95, N110);
nand NAND3 (N126, N18, N6, N74);
nand NAND2 (N127, N101, N114);
not NOT1 (N128, N51);
and AND3 (N129, N126, N65, N116);
and AND4 (N130, N120, N12, N40, N91);
and AND3 (N131, N130, N85, N37);
or OR3 (N132, N127, N106, N4);
buf BUF1 (N133, N119);
nand NAND2 (N134, N132, N126);
xor XOR2 (N135, N133, N64);
nor NOR4 (N136, N121, N9, N34, N43);
or OR2 (N137, N131, N10);
or OR3 (N138, N94, N62, N39);
not NOT1 (N139, N136);
and AND4 (N140, N135, N134, N78, N54);
xor XOR2 (N141, N77, N61);
nand NAND3 (N142, N129, N28, N24);
xor XOR2 (N143, N128, N39);
or OR2 (N144, N125, N98);
and AND2 (N145, N124, N95);
nand NAND4 (N146, N141, N142, N131, N127);
and AND2 (N147, N54, N58);
nand NAND4 (N148, N137, N75, N66, N145);
buf BUF1 (N149, N100);
not NOT1 (N150, N111);
or OR4 (N151, N139, N35, N22, N52);
buf BUF1 (N152, N143);
nand NAND2 (N153, N144, N117);
buf BUF1 (N154, N140);
and AND4 (N155, N138, N50, N98, N102);
not NOT1 (N156, N155);
and AND4 (N157, N151, N83, N90, N77);
nand NAND3 (N158, N152, N140, N25);
nor NOR4 (N159, N157, N74, N132, N6);
and AND3 (N160, N148, N142, N42);
xor XOR2 (N161, N156, N148);
nor NOR2 (N162, N146, N44);
and AND2 (N163, N149, N3);
and AND4 (N164, N159, N102, N134, N87);
buf BUF1 (N165, N147);
nor NOR4 (N166, N161, N147, N125, N132);
not NOT1 (N167, N163);
nand NAND4 (N168, N160, N141, N39, N66);
or OR2 (N169, N167, N50);
and AND3 (N170, N150, N58, N99);
not NOT1 (N171, N166);
or OR4 (N172, N164, N148, N60, N126);
or OR4 (N173, N154, N110, N81, N147);
and AND4 (N174, N170, N69, N170, N66);
or OR4 (N175, N168, N61, N43, N72);
nand NAND2 (N176, N171, N117);
buf BUF1 (N177, N176);
or OR4 (N178, N169, N168, N113, N143);
and AND2 (N179, N175, N134);
and AND3 (N180, N165, N89, N90);
or OR2 (N181, N162, N55);
nor NOR3 (N182, N180, N41, N180);
nand NAND2 (N183, N181, N72);
and AND4 (N184, N178, N78, N131, N182);
nor NOR4 (N185, N23, N33, N113, N154);
nand NAND4 (N186, N153, N95, N79, N31);
or OR2 (N187, N177, N16);
and AND4 (N188, N186, N72, N145, N117);
nor NOR4 (N189, N185, N84, N23, N86);
xor XOR2 (N190, N179, N10);
and AND2 (N191, N174, N140);
nand NAND4 (N192, N189, N164, N55, N39);
xor XOR2 (N193, N190, N162);
or OR2 (N194, N193, N51);
buf BUF1 (N195, N172);
nor NOR2 (N196, N184, N24);
not NOT1 (N197, N158);
nor NOR3 (N198, N183, N14, N187);
not NOT1 (N199, N36);
nand NAND4 (N200, N196, N80, N30, N5);
or OR4 (N201, N192, N152, N28, N78);
not NOT1 (N202, N198);
not NOT1 (N203, N191);
buf BUF1 (N204, N199);
not NOT1 (N205, N194);
buf BUF1 (N206, N205);
xor XOR2 (N207, N201, N107);
and AND3 (N208, N207, N82, N24);
buf BUF1 (N209, N202);
xor XOR2 (N210, N197, N200);
nand NAND3 (N211, N139, N77, N181);
xor XOR2 (N212, N210, N93);
nand NAND2 (N213, N173, N73);
nand NAND3 (N214, N206, N186, N188);
buf BUF1 (N215, N199);
buf BUF1 (N216, N214);
not NOT1 (N217, N208);
nor NOR3 (N218, N209, N106, N140);
nand NAND4 (N219, N213, N160, N154, N202);
buf BUF1 (N220, N204);
and AND4 (N221, N203, N186, N113, N206);
xor XOR2 (N222, N219, N22);
not NOT1 (N223, N216);
and AND2 (N224, N195, N164);
not NOT1 (N225, N218);
xor XOR2 (N226, N220, N217);
nor NOR2 (N227, N98, N13);
buf BUF1 (N228, N221);
nor NOR2 (N229, N228, N115);
nand NAND4 (N230, N227, N228, N217, N145);
xor XOR2 (N231, N230, N186);
not NOT1 (N232, N212);
not NOT1 (N233, N223);
not NOT1 (N234, N215);
xor XOR2 (N235, N231, N139);
xor XOR2 (N236, N235, N153);
not NOT1 (N237, N229);
and AND4 (N238, N232, N16, N6, N185);
nand NAND2 (N239, N224, N90);
or OR4 (N240, N239, N179, N70, N176);
nand NAND4 (N241, N237, N118, N224, N153);
nor NOR3 (N242, N226, N166, N44);
nand NAND4 (N243, N240, N105, N112, N101);
nor NOR4 (N244, N225, N143, N148, N132);
or OR4 (N245, N234, N48, N25, N105);
not NOT1 (N246, N211);
nand NAND2 (N247, N238, N22);
or OR2 (N248, N247, N68);
and AND2 (N249, N236, N189);
xor XOR2 (N250, N248, N193);
nor NOR3 (N251, N222, N196, N154);
nand NAND4 (N252, N243, N31, N2, N100);
not NOT1 (N253, N245);
xor XOR2 (N254, N242, N205);
nand NAND4 (N255, N252, N72, N110, N30);
xor XOR2 (N256, N254, N221);
buf BUF1 (N257, N246);
or OR2 (N258, N256, N213);
xor XOR2 (N259, N244, N216);
nor NOR4 (N260, N249, N94, N166, N99);
and AND4 (N261, N250, N186, N124, N209);
not NOT1 (N262, N258);
buf BUF1 (N263, N262);
and AND3 (N264, N261, N64, N82);
or OR2 (N265, N257, N236);
not NOT1 (N266, N251);
not NOT1 (N267, N253);
or OR2 (N268, N266, N35);
and AND4 (N269, N233, N116, N142, N133);
not NOT1 (N270, N259);
not NOT1 (N271, N241);
or OR3 (N272, N260, N84, N106);
or OR3 (N273, N272, N221, N207);
nand NAND4 (N274, N267, N140, N173, N266);
xor XOR2 (N275, N273, N18);
nand NAND4 (N276, N264, N52, N47, N255);
xor XOR2 (N277, N76, N9);
nor NOR3 (N278, N269, N31, N229);
and AND3 (N279, N268, N263, N15);
not NOT1 (N280, N105);
xor XOR2 (N281, N265, N257);
nand NAND4 (N282, N277, N241, N216, N81);
or OR2 (N283, N282, N240);
buf BUF1 (N284, N276);
or OR3 (N285, N275, N204, N261);
and AND3 (N286, N284, N106, N217);
nor NOR2 (N287, N271, N129);
nor NOR2 (N288, N283, N169);
and AND2 (N289, N281, N102);
or OR2 (N290, N270, N111);
or OR4 (N291, N285, N226, N276, N172);
nand NAND2 (N292, N288, N62);
nor NOR4 (N293, N274, N13, N101, N223);
not NOT1 (N294, N287);
not NOT1 (N295, N292);
nor NOR2 (N296, N294, N44);
xor XOR2 (N297, N295, N38);
not NOT1 (N298, N290);
nor NOR4 (N299, N280, N194, N231, N144);
nor NOR2 (N300, N299, N156);
nor NOR3 (N301, N293, N118, N68);
nand NAND2 (N302, N301, N34);
xor XOR2 (N303, N296, N228);
and AND2 (N304, N278, N294);
and AND2 (N305, N304, N49);
not NOT1 (N306, N289);
nor NOR2 (N307, N306, N300);
xor XOR2 (N308, N192, N128);
not NOT1 (N309, N298);
and AND4 (N310, N279, N252, N275, N166);
nand NAND4 (N311, N310, N154, N281, N233);
not NOT1 (N312, N297);
not NOT1 (N313, N286);
not NOT1 (N314, N313);
xor XOR2 (N315, N302, N311);
or OR2 (N316, N309, N111);
or OR2 (N317, N126, N79);
xor XOR2 (N318, N308, N285);
and AND3 (N319, N307, N128, N96);
and AND2 (N320, N305, N54);
buf BUF1 (N321, N319);
and AND4 (N322, N320, N173, N97, N312);
or OR4 (N323, N171, N307, N15, N125);
xor XOR2 (N324, N314, N101);
or OR4 (N325, N303, N60, N243, N157);
and AND2 (N326, N322, N200);
nor NOR4 (N327, N321, N78, N11, N162);
not NOT1 (N328, N326);
and AND3 (N329, N318, N141, N325);
nor NOR2 (N330, N301, N15);
nor NOR3 (N331, N330, N135, N18);
xor XOR2 (N332, N315, N139);
xor XOR2 (N333, N329, N221);
xor XOR2 (N334, N333, N8);
xor XOR2 (N335, N334, N167);
xor XOR2 (N336, N331, N201);
nand NAND3 (N337, N336, N171, N299);
buf BUF1 (N338, N337);
and AND2 (N339, N291, N130);
or OR2 (N340, N339, N257);
or OR3 (N341, N338, N19, N79);
or OR4 (N342, N340, N224, N8, N277);
buf BUF1 (N343, N317);
and AND2 (N344, N327, N173);
or OR4 (N345, N342, N307, N173, N216);
nor NOR2 (N346, N316, N335);
or OR2 (N347, N328, N1);
or OR2 (N348, N204, N63);
or OR3 (N349, N332, N332, N99);
and AND2 (N350, N344, N227);
buf BUF1 (N351, N348);
nor NOR4 (N352, N347, N153, N22, N152);
nand NAND2 (N353, N345, N182);
buf BUF1 (N354, N324);
or OR3 (N355, N343, N70, N152);
nand NAND3 (N356, N350, N225, N105);
nand NAND3 (N357, N351, N354, N54);
nor NOR3 (N358, N110, N36, N347);
buf BUF1 (N359, N341);
xor XOR2 (N360, N359, N311);
not NOT1 (N361, N353);
xor XOR2 (N362, N352, N96);
or OR2 (N363, N362, N17);
and AND4 (N364, N346, N217, N51, N211);
or OR2 (N365, N356, N157);
nand NAND4 (N366, N365, N76, N170, N187);
or OR2 (N367, N357, N121);
not NOT1 (N368, N366);
buf BUF1 (N369, N360);
nor NOR2 (N370, N358, N269);
or OR4 (N371, N364, N330, N239, N194);
not NOT1 (N372, N368);
buf BUF1 (N373, N361);
buf BUF1 (N374, N323);
nand NAND2 (N375, N367, N327);
xor XOR2 (N376, N374, N249);
and AND2 (N377, N372, N327);
nor NOR2 (N378, N349, N49);
nand NAND2 (N379, N371, N180);
not NOT1 (N380, N369);
nand NAND4 (N381, N375, N221, N240, N117);
and AND4 (N382, N380, N311, N373, N136);
xor XOR2 (N383, N304, N346);
nor NOR3 (N384, N383, N299, N37);
xor XOR2 (N385, N379, N85);
not NOT1 (N386, N376);
xor XOR2 (N387, N370, N312);
xor XOR2 (N388, N381, N294);
or OR4 (N389, N363, N51, N28, N379);
nand NAND3 (N390, N385, N341, N200);
xor XOR2 (N391, N388, N248);
nor NOR4 (N392, N384, N281, N125, N101);
and AND4 (N393, N387, N249, N77, N370);
nor NOR4 (N394, N392, N247, N365, N7);
and AND4 (N395, N393, N251, N128, N374);
and AND3 (N396, N391, N36, N36);
nor NOR2 (N397, N396, N197);
nor NOR3 (N398, N397, N380, N282);
and AND4 (N399, N395, N58, N150, N97);
not NOT1 (N400, N394);
nand NAND2 (N401, N389, N2);
not NOT1 (N402, N386);
or OR3 (N403, N400, N307, N388);
or OR3 (N404, N403, N160, N275);
nand NAND4 (N405, N398, N156, N86, N294);
buf BUF1 (N406, N404);
buf BUF1 (N407, N390);
nor NOR2 (N408, N402, N171);
not NOT1 (N409, N405);
xor XOR2 (N410, N378, N204);
xor XOR2 (N411, N407, N176);
and AND2 (N412, N355, N163);
xor XOR2 (N413, N409, N186);
nor NOR3 (N414, N401, N167, N4);
or OR4 (N415, N412, N148, N159, N373);
not NOT1 (N416, N399);
not NOT1 (N417, N406);
xor XOR2 (N418, N408, N235);
nand NAND4 (N419, N382, N37, N247, N306);
not NOT1 (N420, N410);
xor XOR2 (N421, N414, N214);
nand NAND3 (N422, N420, N114, N114);
nor NOR3 (N423, N377, N69, N200);
nor NOR3 (N424, N417, N277, N181);
nor NOR2 (N425, N413, N299);
buf BUF1 (N426, N423);
xor XOR2 (N427, N424, N274);
or OR4 (N428, N421, N1, N208, N357);
and AND4 (N429, N425, N34, N117, N369);
nand NAND3 (N430, N428, N428, N392);
xor XOR2 (N431, N422, N326);
and AND4 (N432, N430, N343, N386, N367);
xor XOR2 (N433, N418, N305);
xor XOR2 (N434, N433, N257);
and AND4 (N435, N419, N36, N138, N168);
or OR4 (N436, N415, N41, N131, N20);
and AND2 (N437, N426, N275);
nand NAND4 (N438, N416, N105, N188, N387);
nor NOR2 (N439, N432, N30);
nand NAND2 (N440, N434, N8);
and AND2 (N441, N429, N70);
buf BUF1 (N442, N439);
not NOT1 (N443, N436);
nand NAND3 (N444, N427, N116, N327);
nand NAND4 (N445, N441, N140, N410, N347);
or OR2 (N446, N443, N323);
nor NOR3 (N447, N431, N209, N272);
nor NOR4 (N448, N445, N268, N69, N406);
not NOT1 (N449, N447);
xor XOR2 (N450, N442, N6);
not NOT1 (N451, N440);
not NOT1 (N452, N449);
and AND3 (N453, N452, N247, N272);
nand NAND4 (N454, N446, N53, N209, N445);
buf BUF1 (N455, N435);
buf BUF1 (N456, N444);
nand NAND2 (N457, N454, N96);
nand NAND3 (N458, N437, N2, N65);
buf BUF1 (N459, N438);
or OR2 (N460, N448, N124);
and AND4 (N461, N459, N38, N44, N345);
buf BUF1 (N462, N461);
buf BUF1 (N463, N411);
xor XOR2 (N464, N450, N24);
and AND4 (N465, N453, N127, N325, N388);
nand NAND4 (N466, N457, N2, N435, N193);
xor XOR2 (N467, N451, N123);
nand NAND4 (N468, N462, N435, N329, N207);
not NOT1 (N469, N460);
nand NAND4 (N470, N466, N215, N239, N69);
or OR2 (N471, N469, N234);
or OR3 (N472, N458, N275, N37);
nand NAND3 (N473, N456, N273, N7);
xor XOR2 (N474, N473, N417);
nor NOR4 (N475, N474, N407, N453, N56);
xor XOR2 (N476, N472, N471);
nand NAND3 (N477, N84, N109, N199);
or OR2 (N478, N463, N458);
xor XOR2 (N479, N467, N459);
or OR2 (N480, N479, N359);
and AND2 (N481, N465, N154);
or OR4 (N482, N478, N330, N229, N45);
not NOT1 (N483, N470);
nor NOR3 (N484, N480, N294, N131);
nor NOR3 (N485, N483, N145, N80);
not NOT1 (N486, N482);
and AND2 (N487, N476, N135);
not NOT1 (N488, N484);
or OR3 (N489, N477, N406, N444);
or OR4 (N490, N475, N427, N271, N340);
nor NOR2 (N491, N455, N56);
and AND3 (N492, N491, N50, N247);
or OR4 (N493, N488, N214, N486, N144);
not NOT1 (N494, N117);
nand NAND2 (N495, N468, N331);
xor XOR2 (N496, N492, N285);
nor NOR4 (N497, N494, N450, N454, N283);
nand NAND2 (N498, N487, N477);
nor NOR2 (N499, N489, N120);
nor NOR3 (N500, N490, N319, N100);
and AND4 (N501, N464, N450, N52, N343);
nand NAND4 (N502, N481, N13, N59, N257);
buf BUF1 (N503, N499);
xor XOR2 (N504, N496, N73);
not NOT1 (N505, N504);
not NOT1 (N506, N498);
nand NAND3 (N507, N495, N110, N402);
not NOT1 (N508, N502);
xor XOR2 (N509, N501, N77);
not NOT1 (N510, N493);
or OR4 (N511, N506, N361, N385, N146);
buf BUF1 (N512, N503);
xor XOR2 (N513, N500, N237);
nand NAND4 (N514, N505, N229, N472, N81);
nand NAND3 (N515, N513, N224, N30);
and AND3 (N516, N510, N426, N395);
xor XOR2 (N517, N485, N355);
not NOT1 (N518, N511);
or OR3 (N519, N508, N358, N327);
not NOT1 (N520, N509);
and AND3 (N521, N518, N43, N518);
not NOT1 (N522, N497);
not NOT1 (N523, N522);
nand NAND2 (N524, N514, N230);
buf BUF1 (N525, N523);
buf BUF1 (N526, N521);
buf BUF1 (N527, N519);
buf BUF1 (N528, N512);
and AND3 (N529, N524, N129, N1);
not NOT1 (N530, N529);
nand NAND2 (N531, N527, N446);
or OR3 (N532, N517, N454, N530);
nor NOR2 (N533, N480, N331);
nor NOR2 (N534, N528, N222);
xor XOR2 (N535, N531, N362);
nor NOR4 (N536, N516, N69, N204, N202);
buf BUF1 (N537, N536);
nand NAND3 (N538, N533, N409, N25);
nor NOR3 (N539, N525, N442, N137);
nand NAND3 (N540, N539, N232, N159);
nor NOR3 (N541, N540, N511, N378);
buf BUF1 (N542, N537);
and AND4 (N543, N535, N235, N35, N264);
buf BUF1 (N544, N542);
and AND2 (N545, N532, N382);
nor NOR4 (N546, N526, N189, N211, N2);
nor NOR4 (N547, N534, N346, N393, N447);
xor XOR2 (N548, N538, N338);
and AND2 (N549, N507, N385);
nand NAND3 (N550, N546, N204, N325);
nor NOR3 (N551, N547, N207, N411);
buf BUF1 (N552, N541);
buf BUF1 (N553, N545);
xor XOR2 (N554, N550, N484);
and AND3 (N555, N520, N402, N144);
or OR3 (N556, N548, N415, N187);
nor NOR4 (N557, N543, N412, N313, N230);
xor XOR2 (N558, N554, N340);
not NOT1 (N559, N553);
nor NOR4 (N560, N559, N208, N74, N131);
not NOT1 (N561, N515);
nand NAND3 (N562, N552, N484, N520);
not NOT1 (N563, N555);
not NOT1 (N564, N549);
xor XOR2 (N565, N558, N222);
nand NAND3 (N566, N561, N444, N190);
xor XOR2 (N567, N565, N535);
buf BUF1 (N568, N557);
xor XOR2 (N569, N563, N251);
nor NOR4 (N570, N568, N227, N456, N535);
nand NAND2 (N571, N560, N411);
not NOT1 (N572, N566);
not NOT1 (N573, N564);
xor XOR2 (N574, N551, N214);
and AND4 (N575, N544, N457, N372, N465);
not NOT1 (N576, N574);
nor NOR3 (N577, N562, N229, N291);
or OR4 (N578, N576, N183, N35, N468);
nor NOR4 (N579, N577, N566, N27, N398);
or OR3 (N580, N571, N492, N563);
nand NAND2 (N581, N567, N129);
buf BUF1 (N582, N572);
xor XOR2 (N583, N579, N129);
buf BUF1 (N584, N582);
or OR3 (N585, N580, N495, N422);
not NOT1 (N586, N556);
or OR3 (N587, N581, N37, N18);
buf BUF1 (N588, N573);
and AND2 (N589, N578, N468);
xor XOR2 (N590, N585, N33);
nand NAND3 (N591, N584, N427, N75);
not NOT1 (N592, N570);
or OR2 (N593, N588, N65);
and AND2 (N594, N591, N508);
nand NAND4 (N595, N590, N452, N581, N553);
or OR3 (N596, N594, N118, N35);
nand NAND4 (N597, N596, N533, N186, N321);
nand NAND2 (N598, N575, N101);
xor XOR2 (N599, N593, N359);
nor NOR2 (N600, N586, N207);
buf BUF1 (N601, N587);
not NOT1 (N602, N589);
xor XOR2 (N603, N569, N165);
or OR4 (N604, N603, N429, N236, N590);
xor XOR2 (N605, N583, N215);
buf BUF1 (N606, N597);
or OR4 (N607, N602, N18, N401, N268);
nand NAND4 (N608, N601, N524, N476, N158);
not NOT1 (N609, N595);
not NOT1 (N610, N605);
nand NAND2 (N611, N606, N93);
or OR4 (N612, N600, N438, N464, N243);
and AND3 (N613, N592, N544, N206);
or OR3 (N614, N599, N553, N438);
nor NOR3 (N615, N613, N570, N200);
nand NAND3 (N616, N614, N256, N89);
xor XOR2 (N617, N610, N490);
nor NOR2 (N618, N615, N17);
or OR3 (N619, N616, N283, N566);
and AND4 (N620, N609, N106, N611, N268);
not NOT1 (N621, N412);
xor XOR2 (N622, N612, N498);
not NOT1 (N623, N617);
nor NOR3 (N624, N619, N51, N511);
nor NOR3 (N625, N618, N385, N153);
or OR4 (N626, N604, N521, N34, N9);
xor XOR2 (N627, N620, N137);
nand NAND2 (N628, N625, N237);
nand NAND4 (N629, N623, N318, N612, N285);
not NOT1 (N630, N626);
or OR4 (N631, N621, N519, N247, N470);
or OR2 (N632, N608, N408);
xor XOR2 (N633, N630, N491);
nor NOR4 (N634, N632, N380, N206, N14);
and AND3 (N635, N633, N325, N251);
not NOT1 (N636, N628);
nor NOR3 (N637, N624, N586, N412);
xor XOR2 (N638, N634, N130);
buf BUF1 (N639, N635);
nor NOR4 (N640, N639, N412, N630, N302);
nand NAND2 (N641, N629, N277);
not NOT1 (N642, N641);
and AND2 (N643, N607, N195);
nor NOR3 (N644, N642, N193, N431);
or OR4 (N645, N643, N256, N441, N618);
nand NAND4 (N646, N627, N257, N224, N20);
not NOT1 (N647, N640);
nand NAND2 (N648, N646, N277);
or OR3 (N649, N638, N29, N112);
xor XOR2 (N650, N647, N429);
and AND3 (N651, N649, N194, N507);
nor NOR3 (N652, N631, N425, N98);
nor NOR2 (N653, N636, N593);
not NOT1 (N654, N622);
or OR3 (N655, N653, N576, N433);
or OR2 (N656, N655, N53);
buf BUF1 (N657, N648);
buf BUF1 (N658, N657);
and AND3 (N659, N644, N466, N127);
xor XOR2 (N660, N650, N347);
or OR4 (N661, N598, N641, N247, N258);
nand NAND4 (N662, N656, N306, N374, N264);
nor NOR4 (N663, N651, N196, N131, N524);
buf BUF1 (N664, N660);
or OR2 (N665, N645, N388);
nor NOR2 (N666, N658, N396);
and AND2 (N667, N659, N392);
not NOT1 (N668, N637);
buf BUF1 (N669, N665);
nand NAND3 (N670, N661, N300, N668);
xor XOR2 (N671, N495, N517);
nor NOR2 (N672, N666, N332);
and AND4 (N673, N652, N103, N540, N62);
nand NAND2 (N674, N662, N162);
nor NOR3 (N675, N670, N612, N108);
or OR4 (N676, N667, N260, N120, N158);
nor NOR3 (N677, N654, N565, N400);
buf BUF1 (N678, N671);
and AND4 (N679, N677, N249, N72, N179);
and AND3 (N680, N669, N61, N322);
xor XOR2 (N681, N679, N263);
or OR2 (N682, N674, N336);
not NOT1 (N683, N676);
or OR2 (N684, N682, N348);
or OR4 (N685, N673, N136, N32, N682);
and AND2 (N686, N664, N268);
buf BUF1 (N687, N675);
not NOT1 (N688, N683);
nor NOR3 (N689, N678, N71, N655);
xor XOR2 (N690, N686, N575);
and AND4 (N691, N685, N165, N22, N450);
nand NAND2 (N692, N672, N649);
nor NOR4 (N693, N692, N393, N347, N523);
xor XOR2 (N694, N687, N347);
or OR2 (N695, N688, N589);
buf BUF1 (N696, N691);
xor XOR2 (N697, N680, N390);
nor NOR3 (N698, N693, N109, N575);
buf BUF1 (N699, N684);
nor NOR2 (N700, N698, N154);
xor XOR2 (N701, N697, N387);
or OR2 (N702, N699, N145);
buf BUF1 (N703, N695);
buf BUF1 (N704, N703);
xor XOR2 (N705, N696, N125);
nor NOR4 (N706, N663, N603, N269, N201);
and AND2 (N707, N689, N609);
xor XOR2 (N708, N707, N610);
and AND3 (N709, N702, N79, N642);
nor NOR3 (N710, N708, N524, N197);
or OR3 (N711, N700, N298, N101);
or OR2 (N712, N681, N525);
nor NOR4 (N713, N694, N289, N497, N362);
or OR2 (N714, N704, N86);
nand NAND2 (N715, N712, N273);
and AND2 (N716, N711, N658);
nor NOR3 (N717, N705, N558, N439);
not NOT1 (N718, N690);
xor XOR2 (N719, N706, N107);
endmodule