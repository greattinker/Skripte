// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N25614,N25609,N25616,N25600,N25621,N25615,N25623,N25619,N25622,N25624;

not NOT1 (N25, N4);
nand NAND3 (N26, N10, N7, N23);
xor XOR2 (N27, N9, N25);
or OR2 (N28, N23, N12);
or OR3 (N29, N16, N6, N11);
not NOT1 (N30, N22);
or OR4 (N31, N9, N6, N29, N10);
buf BUF1 (N32, N13);
or OR2 (N33, N8, N25);
buf BUF1 (N34, N24);
buf BUF1 (N35, N26);
buf BUF1 (N36, N4);
buf BUF1 (N37, N19);
not NOT1 (N38, N27);
xor XOR2 (N39, N30, N27);
or OR4 (N40, N34, N18, N39, N21);
and AND2 (N41, N23, N28);
buf BUF1 (N42, N1);
not NOT1 (N43, N42);
nand NAND4 (N44, N40, N25, N31, N25);
buf BUF1 (N45, N25);
and AND3 (N46, N41, N20, N18);
nand NAND2 (N47, N32, N35);
or OR4 (N48, N19, N31, N28, N40);
and AND4 (N49, N46, N48, N47, N31);
or OR4 (N50, N2, N12, N28, N40);
nand NAND3 (N51, N32, N5, N20);
nand NAND2 (N52, N37, N2);
buf BUF1 (N53, N36);
buf BUF1 (N54, N45);
nand NAND2 (N55, N51, N49);
and AND3 (N56, N7, N8, N10);
xor XOR2 (N57, N38, N50);
and AND4 (N58, N11, N37, N35, N48);
or OR4 (N59, N58, N30, N33, N31);
xor XOR2 (N60, N31, N57);
or OR3 (N61, N23, N5, N11);
or OR4 (N62, N61, N32, N32, N59);
xor XOR2 (N63, N28, N17);
nand NAND2 (N64, N54, N4);
buf BUF1 (N65, N60);
nor NOR4 (N66, N55, N14, N57, N53);
xor XOR2 (N67, N30, N10);
xor XOR2 (N68, N67, N19);
nand NAND4 (N69, N64, N59, N21, N30);
nor NOR3 (N70, N44, N16, N8);
buf BUF1 (N71, N56);
xor XOR2 (N72, N52, N64);
or OR3 (N73, N68, N47, N39);
not NOT1 (N74, N63);
or OR2 (N75, N65, N6);
xor XOR2 (N76, N72, N70);
nand NAND3 (N77, N33, N2, N56);
buf BUF1 (N78, N62);
buf BUF1 (N79, N71);
nor NOR4 (N80, N78, N21, N27, N65);
not NOT1 (N81, N74);
xor XOR2 (N82, N43, N68);
or OR2 (N83, N75, N52);
nand NAND4 (N84, N82, N16, N54, N25);
not NOT1 (N85, N76);
xor XOR2 (N86, N69, N23);
nand NAND3 (N87, N83, N11, N34);
not NOT1 (N88, N86);
buf BUF1 (N89, N81);
buf BUF1 (N90, N73);
or OR3 (N91, N80, N6, N47);
nor NOR3 (N92, N85, N29, N12);
xor XOR2 (N93, N87, N3);
nand NAND4 (N94, N92, N14, N48, N8);
nor NOR3 (N95, N91, N81, N57);
xor XOR2 (N96, N89, N87);
not NOT1 (N97, N77);
or OR2 (N98, N79, N17);
or OR4 (N99, N88, N71, N8, N63);
and AND3 (N100, N94, N26, N49);
buf BUF1 (N101, N95);
or OR4 (N102, N84, N10, N54, N6);
nand NAND2 (N103, N96, N59);
and AND4 (N104, N102, N27, N89, N94);
xor XOR2 (N105, N93, N41);
nor NOR4 (N106, N100, N76, N32, N14);
or OR4 (N107, N105, N9, N68, N79);
xor XOR2 (N108, N99, N90);
nor NOR3 (N109, N92, N41, N92);
buf BUF1 (N110, N98);
nor NOR4 (N111, N109, N12, N14, N39);
xor XOR2 (N112, N110, N29);
nor NOR3 (N113, N104, N3, N59);
nor NOR2 (N114, N112, N2);
buf BUF1 (N115, N114);
nand NAND4 (N116, N111, N96, N52, N94);
nor NOR3 (N117, N108, N82, N47);
xor XOR2 (N118, N97, N79);
or OR3 (N119, N103, N58, N45);
buf BUF1 (N120, N101);
xor XOR2 (N121, N116, N50);
and AND2 (N122, N121, N4);
xor XOR2 (N123, N115, N23);
buf BUF1 (N124, N123);
nand NAND4 (N125, N117, N122, N23, N99);
not NOT1 (N126, N44);
nor NOR2 (N127, N118, N65);
buf BUF1 (N128, N113);
and AND4 (N129, N124, N6, N79, N55);
nand NAND2 (N130, N107, N51);
nor NOR2 (N131, N120, N43);
or OR4 (N132, N131, N57, N130, N17);
nor NOR3 (N133, N20, N48, N111);
buf BUF1 (N134, N128);
nor NOR2 (N135, N126, N74);
xor XOR2 (N136, N132, N104);
buf BUF1 (N137, N136);
or OR2 (N138, N137, N2);
nand NAND2 (N139, N138, N133);
not NOT1 (N140, N93);
or OR4 (N141, N140, N70, N137, N127);
or OR4 (N142, N86, N44, N96, N50);
nor NOR3 (N143, N125, N53, N55);
or OR3 (N144, N119, N53, N96);
buf BUF1 (N145, N134);
not NOT1 (N146, N141);
and AND4 (N147, N129, N90, N84, N99);
nor NOR4 (N148, N147, N117, N43, N119);
and AND3 (N149, N106, N123, N88);
or OR3 (N150, N135, N64, N126);
buf BUF1 (N151, N144);
nand NAND2 (N152, N66, N132);
or OR2 (N153, N151, N79);
and AND3 (N154, N153, N88, N121);
not NOT1 (N155, N145);
xor XOR2 (N156, N146, N29);
nand NAND2 (N157, N142, N71);
and AND4 (N158, N148, N26, N67, N147);
not NOT1 (N159, N158);
or OR4 (N160, N156, N54, N39, N19);
or OR2 (N161, N150, N14);
xor XOR2 (N162, N161, N41);
buf BUF1 (N163, N154);
buf BUF1 (N164, N149);
and AND2 (N165, N160, N129);
nor NOR2 (N166, N165, N48);
nor NOR3 (N167, N139, N127, N147);
nand NAND2 (N168, N163, N164);
xor XOR2 (N169, N116, N143);
nand NAND2 (N170, N17, N113);
and AND4 (N171, N168, N32, N14, N67);
not NOT1 (N172, N166);
xor XOR2 (N173, N169, N127);
or OR2 (N174, N170, N29);
and AND3 (N175, N157, N122, N145);
buf BUF1 (N176, N173);
nor NOR4 (N177, N159, N153, N133, N118);
buf BUF1 (N178, N162);
not NOT1 (N179, N175);
xor XOR2 (N180, N177, N109);
nor NOR4 (N181, N176, N72, N180, N150);
nor NOR2 (N182, N1, N62);
nand NAND2 (N183, N152, N93);
buf BUF1 (N184, N179);
nor NOR2 (N185, N171, N13);
and AND2 (N186, N167, N92);
nand NAND2 (N187, N182, N46);
and AND3 (N188, N183, N78, N185);
or OR2 (N189, N76, N112);
nand NAND2 (N190, N155, N56);
and AND2 (N191, N187, N5);
not NOT1 (N192, N188);
nor NOR4 (N193, N181, N4, N188, N99);
nor NOR4 (N194, N192, N175, N158, N61);
or OR4 (N195, N189, N180, N120, N14);
or OR4 (N196, N193, N191, N53, N113);
or OR2 (N197, N90, N57);
buf BUF1 (N198, N172);
nor NOR2 (N199, N198, N8);
nand NAND2 (N200, N178, N111);
nand NAND4 (N201, N186, N130, N187, N121);
buf BUF1 (N202, N174);
nor NOR3 (N203, N200, N9, N120);
not NOT1 (N204, N203);
or OR4 (N205, N194, N117, N102, N71);
and AND3 (N206, N204, N85, N198);
or OR4 (N207, N206, N197, N108, N92);
and AND3 (N208, N68, N91, N99);
or OR3 (N209, N208, N165, N190);
nor NOR3 (N210, N197, N93, N77);
and AND3 (N211, N196, N138, N167);
nand NAND4 (N212, N199, N49, N45, N3);
or OR3 (N213, N195, N197, N82);
buf BUF1 (N214, N209);
not NOT1 (N215, N212);
buf BUF1 (N216, N211);
nand NAND3 (N217, N210, N7, N102);
xor XOR2 (N218, N202, N177);
xor XOR2 (N219, N217, N9);
not NOT1 (N220, N201);
not NOT1 (N221, N205);
nand NAND3 (N222, N207, N106, N96);
and AND4 (N223, N218, N155, N205, N215);
and AND3 (N224, N38, N87, N19);
not NOT1 (N225, N223);
xor XOR2 (N226, N221, N31);
or OR4 (N227, N184, N68, N138, N147);
xor XOR2 (N228, N214, N200);
or OR3 (N229, N222, N173, N43);
xor XOR2 (N230, N229, N115);
nor NOR4 (N231, N225, N186, N23, N147);
xor XOR2 (N232, N219, N122);
not NOT1 (N233, N226);
or OR2 (N234, N233, N119);
nor NOR3 (N235, N224, N139, N10);
buf BUF1 (N236, N220);
nor NOR4 (N237, N216, N44, N64, N107);
xor XOR2 (N238, N230, N109);
or OR2 (N239, N235, N176);
nor NOR4 (N240, N227, N85, N127, N116);
nand NAND2 (N241, N231, N172);
nand NAND4 (N242, N234, N6, N55, N208);
not NOT1 (N243, N213);
buf BUF1 (N244, N241);
not NOT1 (N245, N239);
not NOT1 (N246, N228);
nor NOR2 (N247, N238, N47);
or OR3 (N248, N237, N190, N96);
and AND2 (N249, N246, N40);
nand NAND4 (N250, N240, N88, N157, N168);
not NOT1 (N251, N236);
nand NAND4 (N252, N243, N48, N63, N11);
not NOT1 (N253, N248);
and AND3 (N254, N232, N234, N90);
or OR3 (N255, N252, N34, N217);
buf BUF1 (N256, N254);
xor XOR2 (N257, N244, N82);
and AND4 (N258, N256, N50, N192, N232);
or OR4 (N259, N245, N77, N23, N20);
nand NAND3 (N260, N250, N106, N108);
not NOT1 (N261, N259);
and AND4 (N262, N255, N84, N18, N254);
or OR4 (N263, N251, N5, N51, N204);
buf BUF1 (N264, N242);
not NOT1 (N265, N249);
not NOT1 (N266, N265);
nor NOR4 (N267, N262, N183, N167, N221);
or OR3 (N268, N261, N262, N5);
nor NOR3 (N269, N266, N56, N64);
xor XOR2 (N270, N257, N61);
nor NOR4 (N271, N268, N236, N198, N95);
and AND2 (N272, N258, N254);
buf BUF1 (N273, N270);
not NOT1 (N274, N273);
or OR2 (N275, N271, N231);
nand NAND3 (N276, N269, N3, N267);
and AND3 (N277, N151, N132, N122);
not NOT1 (N278, N260);
not NOT1 (N279, N277);
and AND3 (N280, N279, N99, N79);
buf BUF1 (N281, N276);
buf BUF1 (N282, N264);
xor XOR2 (N283, N282, N123);
nand NAND4 (N284, N275, N117, N191, N100);
nor NOR2 (N285, N284, N72);
and AND4 (N286, N281, N86, N271, N196);
buf BUF1 (N287, N263);
xor XOR2 (N288, N287, N238);
or OR4 (N289, N288, N170, N227, N279);
not NOT1 (N290, N286);
xor XOR2 (N291, N280, N106);
not NOT1 (N292, N272);
not NOT1 (N293, N291);
nor NOR3 (N294, N293, N116, N202);
buf BUF1 (N295, N285);
and AND4 (N296, N247, N246, N130, N137);
xor XOR2 (N297, N296, N183);
nor NOR4 (N298, N292, N247, N61, N99);
or OR2 (N299, N289, N31);
xor XOR2 (N300, N299, N235);
or OR3 (N301, N294, N65, N31);
xor XOR2 (N302, N295, N186);
nor NOR2 (N303, N290, N171);
xor XOR2 (N304, N283, N296);
xor XOR2 (N305, N298, N8);
not NOT1 (N306, N253);
and AND3 (N307, N306, N154, N273);
nor NOR3 (N308, N297, N211, N55);
or OR2 (N309, N307, N168);
not NOT1 (N310, N305);
buf BUF1 (N311, N308);
and AND3 (N312, N301, N62, N182);
xor XOR2 (N313, N309, N102);
and AND4 (N314, N311, N262, N177, N20);
xor XOR2 (N315, N303, N143);
xor XOR2 (N316, N300, N164);
buf BUF1 (N317, N310);
buf BUF1 (N318, N315);
nand NAND3 (N319, N316, N67, N47);
xor XOR2 (N320, N319, N15);
xor XOR2 (N321, N278, N55);
nor NOR4 (N322, N274, N74, N316, N26);
and AND3 (N323, N313, N179, N49);
buf BUF1 (N324, N314);
not NOT1 (N325, N318);
nand NAND3 (N326, N312, N223, N37);
nor NOR4 (N327, N326, N254, N303, N245);
and AND4 (N328, N304, N74, N131, N307);
xor XOR2 (N329, N320, N267);
nand NAND3 (N330, N302, N204, N316);
buf BUF1 (N331, N317);
and AND4 (N332, N323, N187, N131, N182);
nor NOR4 (N333, N327, N52, N56, N249);
nor NOR2 (N334, N322, N127);
xor XOR2 (N335, N331, N324);
and AND3 (N336, N288, N267, N29);
nor NOR3 (N337, N332, N293, N4);
xor XOR2 (N338, N329, N328);
xor XOR2 (N339, N98, N198);
or OR3 (N340, N321, N242, N15);
and AND4 (N341, N330, N130, N41, N271);
or OR2 (N342, N335, N134);
buf BUF1 (N343, N338);
not NOT1 (N344, N334);
and AND3 (N345, N333, N21, N304);
not NOT1 (N346, N340);
not NOT1 (N347, N346);
buf BUF1 (N348, N347);
or OR2 (N349, N344, N3);
nor NOR4 (N350, N345, N321, N319, N98);
and AND2 (N351, N348, N113);
nor NOR3 (N352, N325, N287, N327);
xor XOR2 (N353, N337, N99);
xor XOR2 (N354, N353, N23);
or OR3 (N355, N349, N278, N224);
and AND3 (N356, N343, N100, N199);
nand NAND3 (N357, N352, N79, N211);
nor NOR4 (N358, N339, N306, N296, N116);
buf BUF1 (N359, N350);
xor XOR2 (N360, N341, N234);
nand NAND2 (N361, N351, N291);
xor XOR2 (N362, N342, N206);
buf BUF1 (N363, N360);
not NOT1 (N364, N336);
nand NAND4 (N365, N361, N159, N266, N162);
not NOT1 (N366, N355);
not NOT1 (N367, N363);
not NOT1 (N368, N358);
buf BUF1 (N369, N365);
or OR4 (N370, N369, N19, N202, N27);
or OR3 (N371, N359, N217, N47);
xor XOR2 (N372, N356, N201);
or OR2 (N373, N367, N151);
not NOT1 (N374, N366);
buf BUF1 (N375, N357);
xor XOR2 (N376, N372, N50);
or OR4 (N377, N375, N277, N114, N58);
and AND3 (N378, N371, N285, N245);
nor NOR3 (N379, N368, N173, N270);
and AND2 (N380, N374, N17);
not NOT1 (N381, N373);
nor NOR2 (N382, N377, N284);
xor XOR2 (N383, N378, N358);
buf BUF1 (N384, N362);
xor XOR2 (N385, N383, N19);
xor XOR2 (N386, N384, N29);
not NOT1 (N387, N370);
nor NOR3 (N388, N386, N222, N270);
xor XOR2 (N389, N388, N222);
and AND4 (N390, N389, N237, N378, N329);
buf BUF1 (N391, N390);
or OR2 (N392, N387, N240);
and AND2 (N393, N391, N28);
nand NAND4 (N394, N376, N53, N7, N77);
buf BUF1 (N395, N354);
and AND3 (N396, N382, N381, N312);
not NOT1 (N397, N289);
nor NOR3 (N398, N395, N234, N234);
nand NAND4 (N399, N392, N41, N157, N278);
nor NOR4 (N400, N380, N185, N63, N87);
xor XOR2 (N401, N393, N96);
nand NAND2 (N402, N399, N77);
or OR2 (N403, N401, N89);
buf BUF1 (N404, N396);
xor XOR2 (N405, N403, N156);
or OR3 (N406, N364, N169, N282);
not NOT1 (N407, N405);
nand NAND4 (N408, N397, N257, N298, N271);
or OR4 (N409, N406, N315, N197, N59);
nor NOR2 (N410, N379, N84);
or OR3 (N411, N404, N344, N115);
xor XOR2 (N412, N385, N146);
not NOT1 (N413, N408);
nand NAND2 (N414, N410, N81);
xor XOR2 (N415, N414, N333);
nand NAND2 (N416, N407, N227);
buf BUF1 (N417, N409);
or OR2 (N418, N415, N202);
nor NOR3 (N419, N413, N79, N352);
nor NOR3 (N420, N402, N144, N37);
nor NOR2 (N421, N418, N55);
nand NAND3 (N422, N398, N230, N44);
buf BUF1 (N423, N420);
or OR4 (N424, N417, N276, N122, N39);
or OR3 (N425, N422, N173, N229);
or OR3 (N426, N411, N93, N193);
or OR2 (N427, N426, N193);
not NOT1 (N428, N412);
nor NOR3 (N429, N425, N179, N180);
not NOT1 (N430, N424);
buf BUF1 (N431, N430);
not NOT1 (N432, N428);
nand NAND3 (N433, N423, N261, N290);
not NOT1 (N434, N431);
and AND3 (N435, N433, N52, N279);
and AND3 (N436, N416, N275, N275);
not NOT1 (N437, N400);
or OR3 (N438, N437, N237, N102);
xor XOR2 (N439, N434, N292);
buf BUF1 (N440, N421);
and AND4 (N441, N438, N337, N51, N147);
xor XOR2 (N442, N441, N180);
not NOT1 (N443, N429);
or OR4 (N444, N439, N67, N9, N257);
nand NAND4 (N445, N436, N144, N196, N99);
nor NOR2 (N446, N445, N343);
nor NOR2 (N447, N432, N232);
and AND4 (N448, N447, N139, N345, N410);
not NOT1 (N449, N427);
nand NAND3 (N450, N443, N120, N45);
not NOT1 (N451, N450);
xor XOR2 (N452, N444, N111);
nand NAND2 (N453, N442, N293);
xor XOR2 (N454, N453, N207);
and AND2 (N455, N449, N212);
not NOT1 (N456, N454);
buf BUF1 (N457, N448);
nor NOR4 (N458, N456, N250, N58, N10);
and AND3 (N459, N435, N38, N278);
nor NOR2 (N460, N452, N89);
buf BUF1 (N461, N419);
nand NAND4 (N462, N457, N5, N55, N414);
nand NAND3 (N463, N459, N145, N121);
or OR2 (N464, N463, N109);
nand NAND2 (N465, N446, N293);
xor XOR2 (N466, N461, N110);
buf BUF1 (N467, N458);
and AND3 (N468, N440, N155, N283);
or OR4 (N469, N394, N398, N154, N158);
xor XOR2 (N470, N451, N365);
xor XOR2 (N471, N464, N351);
buf BUF1 (N472, N465);
xor XOR2 (N473, N460, N137);
or OR4 (N474, N471, N133, N221, N459);
xor XOR2 (N475, N462, N214);
not NOT1 (N476, N474);
and AND4 (N477, N470, N356, N466, N434);
not NOT1 (N478, N3);
nor NOR2 (N479, N475, N388);
xor XOR2 (N480, N476, N296);
not NOT1 (N481, N473);
buf BUF1 (N482, N468);
not NOT1 (N483, N481);
nand NAND3 (N484, N482, N220, N109);
nor NOR3 (N485, N472, N75, N329);
not NOT1 (N486, N484);
not NOT1 (N487, N486);
and AND2 (N488, N477, N311);
and AND4 (N489, N483, N349, N402, N403);
not NOT1 (N490, N485);
or OR4 (N491, N469, N9, N18, N365);
not NOT1 (N492, N487);
nor NOR4 (N493, N491, N456, N277, N87);
or OR3 (N494, N488, N114, N198);
xor XOR2 (N495, N478, N418);
buf BUF1 (N496, N479);
or OR3 (N497, N489, N405, N369);
nand NAND4 (N498, N455, N144, N378, N12);
buf BUF1 (N499, N480);
and AND3 (N500, N495, N203, N128);
buf BUF1 (N501, N467);
xor XOR2 (N502, N500, N428);
nand NAND4 (N503, N494, N274, N62, N416);
or OR3 (N504, N503, N348, N15);
buf BUF1 (N505, N499);
xor XOR2 (N506, N501, N93);
and AND4 (N507, N506, N332, N288, N418);
nor NOR4 (N508, N498, N277, N396, N292);
xor XOR2 (N509, N504, N469);
nor NOR3 (N510, N502, N421, N30);
not NOT1 (N511, N490);
and AND2 (N512, N497, N414);
or OR3 (N513, N493, N169, N347);
or OR3 (N514, N513, N88, N299);
buf BUF1 (N515, N514);
nor NOR3 (N516, N509, N183, N79);
buf BUF1 (N517, N496);
not NOT1 (N518, N512);
nand NAND2 (N519, N515, N54);
not NOT1 (N520, N507);
xor XOR2 (N521, N508, N108);
not NOT1 (N522, N510);
nand NAND3 (N523, N505, N303, N442);
not NOT1 (N524, N519);
buf BUF1 (N525, N523);
and AND4 (N526, N517, N268, N511, N18);
xor XOR2 (N527, N453, N53);
nand NAND4 (N528, N527, N75, N45, N174);
nor NOR2 (N529, N518, N344);
xor XOR2 (N530, N524, N226);
or OR3 (N531, N529, N441, N124);
buf BUF1 (N532, N528);
nor NOR3 (N533, N522, N527, N124);
or OR2 (N534, N531, N420);
not NOT1 (N535, N526);
nand NAND3 (N536, N492, N58, N316);
and AND2 (N537, N536, N418);
xor XOR2 (N538, N535, N299);
and AND4 (N539, N521, N493, N209, N411);
xor XOR2 (N540, N539, N471);
or OR2 (N541, N537, N279);
xor XOR2 (N542, N534, N2);
nand NAND4 (N543, N520, N537, N43, N186);
nand NAND4 (N544, N541, N51, N34, N82);
buf BUF1 (N545, N540);
nor NOR3 (N546, N545, N293, N148);
buf BUF1 (N547, N532);
or OR4 (N548, N516, N506, N29, N210);
nand NAND3 (N549, N530, N442, N192);
xor XOR2 (N550, N544, N187);
or OR3 (N551, N538, N529, N435);
and AND2 (N552, N547, N194);
nor NOR3 (N553, N552, N349, N452);
and AND3 (N554, N549, N159, N365);
nand NAND3 (N555, N548, N545, N90);
nand NAND4 (N556, N542, N345, N75, N90);
and AND4 (N557, N551, N191, N113, N86);
nand NAND2 (N558, N546, N22);
or OR2 (N559, N554, N300);
not NOT1 (N560, N525);
and AND3 (N561, N543, N508, N50);
and AND3 (N562, N533, N449, N257);
or OR2 (N563, N555, N312);
not NOT1 (N564, N563);
xor XOR2 (N565, N557, N560);
nand NAND2 (N566, N449, N231);
or OR4 (N567, N561, N388, N190, N37);
and AND3 (N568, N566, N391, N248);
buf BUF1 (N569, N559);
and AND4 (N570, N550, N56, N155, N235);
xor XOR2 (N571, N556, N514);
or OR4 (N572, N553, N168, N94, N64);
nor NOR2 (N573, N571, N326);
buf BUF1 (N574, N570);
xor XOR2 (N575, N558, N394);
xor XOR2 (N576, N575, N157);
buf BUF1 (N577, N568);
buf BUF1 (N578, N569);
not NOT1 (N579, N577);
or OR2 (N580, N562, N268);
not NOT1 (N581, N579);
nand NAND3 (N582, N574, N260, N312);
nor NOR3 (N583, N582, N218, N415);
or OR4 (N584, N578, N556, N87, N318);
nand NAND4 (N585, N584, N93, N428, N209);
nor NOR2 (N586, N585, N179);
xor XOR2 (N587, N581, N437);
nand NAND3 (N588, N572, N305, N500);
nor NOR3 (N589, N583, N518, N17);
nor NOR4 (N590, N565, N490, N266, N293);
not NOT1 (N591, N567);
nand NAND2 (N592, N573, N360);
and AND2 (N593, N576, N58);
nand NAND3 (N594, N587, N380, N483);
or OR3 (N595, N591, N493, N105);
or OR2 (N596, N593, N503);
not NOT1 (N597, N592);
not NOT1 (N598, N586);
buf BUF1 (N599, N598);
not NOT1 (N600, N588);
nor NOR4 (N601, N589, N2, N155, N313);
nor NOR3 (N602, N596, N583, N187);
and AND2 (N603, N590, N405);
buf BUF1 (N604, N599);
nor NOR4 (N605, N602, N70, N222, N190);
not NOT1 (N606, N594);
not NOT1 (N607, N595);
xor XOR2 (N608, N605, N43);
nand NAND3 (N609, N603, N466, N231);
nand NAND4 (N610, N606, N275, N422, N221);
nand NAND3 (N611, N607, N83, N241);
nand NAND4 (N612, N601, N264, N366, N156);
and AND3 (N613, N597, N60, N562);
nor NOR3 (N614, N609, N104, N350);
and AND3 (N615, N614, N417, N459);
not NOT1 (N616, N600);
nand NAND2 (N617, N613, N471);
nand NAND4 (N618, N610, N362, N599, N357);
buf BUF1 (N619, N611);
nor NOR2 (N620, N612, N281);
and AND3 (N621, N616, N516, N490);
or OR4 (N622, N620, N354, N71, N410);
nor NOR2 (N623, N621, N74);
nand NAND3 (N624, N623, N9, N128);
and AND4 (N625, N580, N291, N563, N465);
buf BUF1 (N626, N622);
or OR2 (N627, N625, N177);
and AND3 (N628, N564, N407, N549);
or OR2 (N629, N626, N98);
nor NOR3 (N630, N617, N456, N338);
xor XOR2 (N631, N604, N578);
and AND2 (N632, N608, N627);
xor XOR2 (N633, N529, N543);
or OR2 (N634, N619, N457);
and AND2 (N635, N624, N113);
nor NOR3 (N636, N634, N297, N361);
buf BUF1 (N637, N632);
nand NAND2 (N638, N615, N548);
buf BUF1 (N639, N618);
not NOT1 (N640, N635);
xor XOR2 (N641, N629, N389);
xor XOR2 (N642, N628, N443);
nor NOR2 (N643, N639, N211);
nor NOR3 (N644, N630, N128, N463);
or OR3 (N645, N641, N297, N369);
nor NOR4 (N646, N644, N101, N85, N38);
nand NAND2 (N647, N637, N363);
nor NOR3 (N648, N646, N18, N23);
and AND2 (N649, N640, N256);
and AND3 (N650, N642, N68, N273);
not NOT1 (N651, N647);
not NOT1 (N652, N636);
nand NAND2 (N653, N651, N10);
nor NOR4 (N654, N648, N552, N398, N566);
nand NAND2 (N655, N649, N257);
buf BUF1 (N656, N643);
xor XOR2 (N657, N650, N431);
or OR2 (N658, N657, N11);
xor XOR2 (N659, N652, N566);
nand NAND4 (N660, N631, N149, N303, N22);
buf BUF1 (N661, N655);
and AND4 (N662, N638, N588, N358, N566);
buf BUF1 (N663, N654);
or OR2 (N664, N645, N502);
nor NOR4 (N665, N633, N181, N398, N622);
and AND4 (N666, N658, N292, N312, N155);
xor XOR2 (N667, N666, N37);
nor NOR4 (N668, N665, N454, N432, N451);
buf BUF1 (N669, N664);
xor XOR2 (N670, N661, N236);
and AND3 (N671, N669, N391, N198);
nor NOR3 (N672, N668, N632, N253);
nor NOR3 (N673, N670, N471, N500);
or OR3 (N674, N663, N64, N325);
and AND4 (N675, N667, N285, N91, N609);
buf BUF1 (N676, N673);
not NOT1 (N677, N671);
or OR3 (N678, N656, N357, N392);
or OR4 (N679, N678, N599, N143, N296);
not NOT1 (N680, N653);
nor NOR4 (N681, N672, N72, N130, N75);
buf BUF1 (N682, N675);
buf BUF1 (N683, N680);
nor NOR2 (N684, N679, N386);
xor XOR2 (N685, N676, N31);
nand NAND2 (N686, N684, N326);
and AND3 (N687, N677, N128, N367);
xor XOR2 (N688, N682, N263);
nand NAND4 (N689, N681, N288, N547, N610);
not NOT1 (N690, N660);
not NOT1 (N691, N662);
not NOT1 (N692, N686);
buf BUF1 (N693, N685);
and AND4 (N694, N688, N601, N598, N587);
nor NOR4 (N695, N692, N249, N587, N591);
buf BUF1 (N696, N695);
or OR3 (N697, N683, N212, N55);
xor XOR2 (N698, N689, N140);
and AND2 (N699, N696, N152);
and AND3 (N700, N697, N381, N517);
xor XOR2 (N701, N674, N319);
nand NAND4 (N702, N659, N589, N524, N259);
and AND4 (N703, N687, N657, N294, N694);
buf BUF1 (N704, N522);
nand NAND2 (N705, N700, N4);
nor NOR4 (N706, N690, N127, N614, N334);
nand NAND3 (N707, N705, N316, N19);
and AND3 (N708, N704, N390, N644);
xor XOR2 (N709, N708, N69);
xor XOR2 (N710, N709, N653);
nor NOR2 (N711, N699, N682);
xor XOR2 (N712, N707, N470);
not NOT1 (N713, N702);
nor NOR3 (N714, N710, N700, N429);
and AND3 (N715, N712, N308, N165);
nand NAND4 (N716, N714, N91, N39, N6);
nor NOR2 (N717, N711, N127);
buf BUF1 (N718, N701);
buf BUF1 (N719, N718);
not NOT1 (N720, N719);
buf BUF1 (N721, N716);
buf BUF1 (N722, N720);
xor XOR2 (N723, N713, N464);
buf BUF1 (N724, N703);
not NOT1 (N725, N723);
nand NAND2 (N726, N717, N178);
not NOT1 (N727, N706);
nor NOR4 (N728, N693, N86, N415, N712);
or OR4 (N729, N722, N527, N330, N660);
not NOT1 (N730, N727);
or OR3 (N731, N726, N140, N419);
buf BUF1 (N732, N728);
buf BUF1 (N733, N691);
not NOT1 (N734, N730);
not NOT1 (N735, N731);
buf BUF1 (N736, N729);
or OR4 (N737, N724, N487, N500, N71);
nand NAND3 (N738, N732, N69, N369);
nand NAND2 (N739, N715, N155);
not NOT1 (N740, N725);
not NOT1 (N741, N735);
and AND2 (N742, N733, N403);
xor XOR2 (N743, N740, N479);
nor NOR3 (N744, N698, N616, N440);
xor XOR2 (N745, N744, N412);
not NOT1 (N746, N737);
or OR2 (N747, N741, N524);
xor XOR2 (N748, N736, N374);
not NOT1 (N749, N738);
and AND2 (N750, N745, N431);
and AND3 (N751, N739, N101, N666);
not NOT1 (N752, N743);
nand NAND2 (N753, N749, N73);
not NOT1 (N754, N747);
or OR2 (N755, N750, N229);
xor XOR2 (N756, N742, N733);
buf BUF1 (N757, N752);
not NOT1 (N758, N748);
or OR4 (N759, N753, N468, N636, N184);
not NOT1 (N760, N754);
nand NAND3 (N761, N758, N6, N492);
nor NOR2 (N762, N751, N307);
nand NAND4 (N763, N756, N703, N607, N90);
xor XOR2 (N764, N734, N155);
nand NAND3 (N765, N759, N291, N385);
not NOT1 (N766, N757);
buf BUF1 (N767, N763);
and AND4 (N768, N762, N164, N703, N722);
xor XOR2 (N769, N765, N704);
and AND3 (N770, N769, N686, N630);
nand NAND3 (N771, N767, N173, N460);
nand NAND2 (N772, N768, N411);
buf BUF1 (N773, N770);
or OR3 (N774, N721, N737, N670);
and AND3 (N775, N774, N524, N405);
and AND3 (N776, N766, N196, N128);
buf BUF1 (N777, N746);
nand NAND2 (N778, N775, N378);
nor NOR3 (N779, N777, N728, N3);
or OR3 (N780, N764, N388, N472);
buf BUF1 (N781, N760);
buf BUF1 (N782, N781);
not NOT1 (N783, N772);
xor XOR2 (N784, N779, N189);
nand NAND4 (N785, N761, N395, N202, N154);
nor NOR4 (N786, N773, N277, N353, N78);
and AND3 (N787, N755, N378, N184);
nand NAND2 (N788, N780, N262);
not NOT1 (N789, N786);
or OR4 (N790, N788, N69, N756, N464);
xor XOR2 (N791, N784, N381);
nand NAND3 (N792, N787, N233, N428);
buf BUF1 (N793, N790);
or OR2 (N794, N789, N79);
or OR2 (N795, N778, N441);
nor NOR4 (N796, N776, N700, N219, N426);
nand NAND2 (N797, N794, N742);
nor NOR3 (N798, N782, N68, N184);
or OR2 (N799, N793, N503);
or OR4 (N800, N796, N778, N80, N419);
or OR2 (N801, N797, N595);
nand NAND2 (N802, N785, N459);
xor XOR2 (N803, N795, N420);
nand NAND2 (N804, N801, N255);
buf BUF1 (N805, N783);
not NOT1 (N806, N802);
buf BUF1 (N807, N805);
or OR4 (N808, N803, N345, N565, N740);
xor XOR2 (N809, N771, N214);
nand NAND3 (N810, N807, N326, N273);
and AND3 (N811, N792, N46, N585);
nand NAND2 (N812, N806, N697);
or OR3 (N813, N810, N8, N446);
or OR3 (N814, N798, N797, N223);
xor XOR2 (N815, N811, N600);
not NOT1 (N816, N815);
buf BUF1 (N817, N808);
xor XOR2 (N818, N814, N336);
or OR4 (N819, N809, N362, N430, N400);
nor NOR2 (N820, N819, N800);
xor XOR2 (N821, N94, N452);
nor NOR2 (N822, N818, N195);
buf BUF1 (N823, N820);
nor NOR2 (N824, N791, N731);
buf BUF1 (N825, N804);
nor NOR4 (N826, N812, N143, N718, N388);
buf BUF1 (N827, N821);
buf BUF1 (N828, N822);
xor XOR2 (N829, N813, N59);
and AND2 (N830, N799, N384);
nand NAND4 (N831, N817, N634, N638, N18);
nor NOR3 (N832, N830, N81, N303);
nor NOR2 (N833, N823, N157);
and AND3 (N834, N829, N789, N187);
buf BUF1 (N835, N831);
nor NOR3 (N836, N828, N549, N594);
nor NOR2 (N837, N833, N549);
xor XOR2 (N838, N825, N802);
nor NOR3 (N839, N832, N664, N605);
xor XOR2 (N840, N826, N159);
and AND2 (N841, N837, N276);
nand NAND2 (N842, N838, N125);
buf BUF1 (N843, N827);
nand NAND2 (N844, N816, N337);
nor NOR2 (N845, N835, N491);
nand NAND2 (N846, N843, N484);
nand NAND2 (N847, N834, N563);
buf BUF1 (N848, N840);
nand NAND3 (N849, N848, N124, N490);
and AND4 (N850, N849, N712, N501, N194);
and AND4 (N851, N850, N372, N31, N32);
nand NAND2 (N852, N844, N56);
and AND2 (N853, N845, N529);
nand NAND4 (N854, N851, N463, N671, N285);
xor XOR2 (N855, N852, N353);
not NOT1 (N856, N824);
buf BUF1 (N857, N839);
not NOT1 (N858, N855);
not NOT1 (N859, N858);
not NOT1 (N860, N854);
nand NAND3 (N861, N847, N161, N296);
not NOT1 (N862, N856);
nor NOR2 (N863, N859, N111);
and AND4 (N864, N836, N533, N615, N693);
and AND3 (N865, N841, N804, N290);
buf BUF1 (N866, N865);
nor NOR4 (N867, N842, N295, N23, N56);
buf BUF1 (N868, N857);
nand NAND4 (N869, N863, N229, N111, N117);
not NOT1 (N870, N868);
not NOT1 (N871, N846);
xor XOR2 (N872, N866, N279);
or OR4 (N873, N861, N129, N684, N733);
buf BUF1 (N874, N862);
and AND3 (N875, N853, N257, N775);
not NOT1 (N876, N875);
or OR2 (N877, N860, N816);
and AND2 (N878, N871, N71);
not NOT1 (N879, N877);
and AND2 (N880, N872, N486);
nor NOR4 (N881, N864, N293, N776, N235);
nand NAND3 (N882, N870, N152, N64);
and AND2 (N883, N873, N669);
not NOT1 (N884, N869);
nor NOR3 (N885, N878, N63, N775);
or OR3 (N886, N885, N534, N838);
nor NOR4 (N887, N881, N106, N321, N774);
xor XOR2 (N888, N880, N789);
nor NOR4 (N889, N867, N306, N251, N627);
or OR2 (N890, N882, N108);
buf BUF1 (N891, N874);
xor XOR2 (N892, N888, N353);
buf BUF1 (N893, N889);
and AND2 (N894, N886, N715);
or OR3 (N895, N884, N382, N266);
buf BUF1 (N896, N891);
and AND4 (N897, N876, N373, N572, N250);
or OR3 (N898, N890, N378, N891);
buf BUF1 (N899, N879);
not NOT1 (N900, N896);
buf BUF1 (N901, N893);
nor NOR2 (N902, N883, N57);
not NOT1 (N903, N898);
nor NOR3 (N904, N901, N543, N218);
not NOT1 (N905, N892);
or OR4 (N906, N900, N380, N647, N626);
buf BUF1 (N907, N904);
buf BUF1 (N908, N899);
buf BUF1 (N909, N908);
and AND3 (N910, N887, N555, N793);
not NOT1 (N911, N902);
not NOT1 (N912, N905);
and AND4 (N913, N897, N189, N554, N163);
and AND2 (N914, N911, N401);
nor NOR2 (N915, N894, N159);
or OR3 (N916, N903, N240, N617);
nand NAND3 (N917, N910, N402, N709);
nand NAND4 (N918, N916, N673, N721, N181);
buf BUF1 (N919, N913);
or OR2 (N920, N909, N264);
nand NAND4 (N921, N895, N249, N154, N557);
and AND4 (N922, N920, N692, N529, N414);
xor XOR2 (N923, N915, N429);
buf BUF1 (N924, N907);
xor XOR2 (N925, N912, N730);
nor NOR4 (N926, N914, N180, N458, N142);
and AND2 (N927, N925, N861);
nand NAND3 (N928, N922, N275, N851);
xor XOR2 (N929, N919, N809);
not NOT1 (N930, N929);
nand NAND3 (N931, N928, N315, N293);
not NOT1 (N932, N917);
nor NOR3 (N933, N924, N158, N421);
not NOT1 (N934, N933);
nand NAND4 (N935, N906, N215, N89, N745);
nand NAND2 (N936, N934, N247);
or OR4 (N937, N931, N594, N107, N201);
or OR4 (N938, N923, N546, N382, N649);
buf BUF1 (N939, N930);
nor NOR3 (N940, N936, N61, N498);
nand NAND3 (N941, N926, N353, N769);
or OR3 (N942, N921, N464, N692);
buf BUF1 (N943, N941);
nand NAND3 (N944, N940, N558, N466);
xor XOR2 (N945, N927, N86);
not NOT1 (N946, N943);
xor XOR2 (N947, N942, N75);
nor NOR3 (N948, N939, N264, N225);
and AND2 (N949, N932, N393);
xor XOR2 (N950, N935, N211);
and AND3 (N951, N938, N356, N171);
nor NOR2 (N952, N944, N422);
nor NOR4 (N953, N937, N297, N762, N712);
nand NAND3 (N954, N949, N118, N177);
buf BUF1 (N955, N954);
not NOT1 (N956, N945);
and AND3 (N957, N918, N10, N439);
xor XOR2 (N958, N952, N626);
buf BUF1 (N959, N950);
nor NOR2 (N960, N959, N221);
buf BUF1 (N961, N955);
not NOT1 (N962, N951);
nor NOR2 (N963, N961, N147);
or OR3 (N964, N947, N859, N219);
and AND4 (N965, N963, N326, N744, N683);
buf BUF1 (N966, N948);
nand NAND4 (N967, N965, N409, N431, N124);
not NOT1 (N968, N960);
or OR2 (N969, N967, N911);
or OR4 (N970, N958, N465, N942, N131);
and AND4 (N971, N956, N97, N87, N773);
and AND4 (N972, N953, N545, N235, N579);
and AND4 (N973, N970, N437, N314, N111);
or OR3 (N974, N966, N566, N698);
not NOT1 (N975, N968);
and AND3 (N976, N973, N728, N879);
xor XOR2 (N977, N957, N885);
or OR3 (N978, N969, N439, N672);
buf BUF1 (N979, N972);
nand NAND4 (N980, N976, N72, N523, N921);
or OR2 (N981, N978, N766);
xor XOR2 (N982, N946, N204);
or OR2 (N983, N971, N583);
and AND3 (N984, N983, N855, N809);
buf BUF1 (N985, N964);
not NOT1 (N986, N979);
buf BUF1 (N987, N984);
nor NOR3 (N988, N981, N117, N879);
xor XOR2 (N989, N988, N753);
or OR3 (N990, N986, N471, N477);
nand NAND3 (N991, N982, N892, N737);
xor XOR2 (N992, N962, N841);
or OR4 (N993, N980, N330, N132, N833);
nor NOR3 (N994, N985, N312, N194);
nor NOR2 (N995, N990, N4);
buf BUF1 (N996, N977);
nand NAND2 (N997, N974, N212);
xor XOR2 (N998, N996, N18);
nor NOR3 (N999, N994, N391, N954);
or OR4 (N1000, N991, N407, N189, N570);
nor NOR4 (N1001, N993, N747, N416, N825);
buf BUF1 (N1002, N1000);
not NOT1 (N1003, N989);
xor XOR2 (N1004, N992, N72);
not NOT1 (N1005, N995);
nor NOR3 (N1006, N1005, N42, N455);
not NOT1 (N1007, N1003);
nand NAND2 (N1008, N987, N25);
and AND3 (N1009, N1001, N931, N370);
nor NOR3 (N1010, N1002, N538, N442);
nand NAND3 (N1011, N1007, N266, N349);
or OR3 (N1012, N1009, N431, N131);
not NOT1 (N1013, N1006);
nand NAND2 (N1014, N1012, N213);
buf BUF1 (N1015, N1004);
and AND2 (N1016, N997, N437);
nor NOR2 (N1017, N1011, N598);
nand NAND3 (N1018, N1013, N991, N442);
xor XOR2 (N1019, N1018, N262);
buf BUF1 (N1020, N1016);
and AND3 (N1021, N1014, N628, N299);
xor XOR2 (N1022, N1019, N157);
or OR2 (N1023, N999, N173);
not NOT1 (N1024, N1023);
nor NOR3 (N1025, N1015, N671, N711);
nor NOR3 (N1026, N1008, N513, N577);
or OR3 (N1027, N1017, N34, N785);
buf BUF1 (N1028, N1021);
nand NAND4 (N1029, N1025, N392, N219, N90);
and AND4 (N1030, N1026, N746, N416, N94);
nor NOR3 (N1031, N998, N1009, N166);
nor NOR3 (N1032, N1030, N763, N318);
nand NAND3 (N1033, N1010, N780, N417);
or OR2 (N1034, N1032, N393);
nand NAND4 (N1035, N1033, N455, N659, N135);
or OR4 (N1036, N1020, N648, N596, N311);
nor NOR3 (N1037, N1035, N899, N50);
or OR2 (N1038, N975, N646);
and AND2 (N1039, N1028, N119);
nor NOR3 (N1040, N1038, N593, N192);
buf BUF1 (N1041, N1024);
not NOT1 (N1042, N1039);
xor XOR2 (N1043, N1034, N1025);
or OR2 (N1044, N1022, N36);
or OR2 (N1045, N1027, N426);
buf BUF1 (N1046, N1044);
or OR3 (N1047, N1031, N334, N375);
nand NAND3 (N1048, N1045, N566, N465);
or OR4 (N1049, N1046, N659, N31, N227);
xor XOR2 (N1050, N1049, N989);
nand NAND2 (N1051, N1036, N757);
buf BUF1 (N1052, N1043);
xor XOR2 (N1053, N1037, N886);
or OR2 (N1054, N1042, N920);
not NOT1 (N1055, N1029);
nand NAND3 (N1056, N1051, N332, N941);
and AND2 (N1057, N1055, N520);
and AND3 (N1058, N1052, N181, N54);
not NOT1 (N1059, N1056);
and AND3 (N1060, N1057, N449, N550);
not NOT1 (N1061, N1048);
not NOT1 (N1062, N1040);
xor XOR2 (N1063, N1053, N638);
xor XOR2 (N1064, N1050, N969);
and AND4 (N1065, N1060, N19, N216, N77);
nand NAND2 (N1066, N1061, N561);
or OR3 (N1067, N1066, N998, N400);
buf BUF1 (N1068, N1054);
xor XOR2 (N1069, N1065, N361);
and AND4 (N1070, N1041, N566, N801, N117);
not NOT1 (N1071, N1058);
nand NAND3 (N1072, N1047, N114, N573);
or OR4 (N1073, N1069, N526, N137, N595);
xor XOR2 (N1074, N1071, N306);
nand NAND4 (N1075, N1063, N148, N938, N76);
nor NOR3 (N1076, N1070, N145, N76);
and AND2 (N1077, N1076, N807);
nand NAND4 (N1078, N1062, N18, N618, N1014);
not NOT1 (N1079, N1075);
buf BUF1 (N1080, N1068);
or OR4 (N1081, N1064, N81, N392, N333);
or OR2 (N1082, N1080, N696);
and AND3 (N1083, N1072, N487, N831);
nor NOR3 (N1084, N1079, N801, N762);
nor NOR4 (N1085, N1081, N1040, N401, N871);
xor XOR2 (N1086, N1067, N6);
or OR4 (N1087, N1083, N597, N790, N234);
and AND4 (N1088, N1078, N328, N921, N80);
nand NAND3 (N1089, N1077, N250, N1062);
or OR4 (N1090, N1087, N661, N1051, N306);
xor XOR2 (N1091, N1073, N8);
or OR3 (N1092, N1084, N235, N46);
xor XOR2 (N1093, N1090, N501);
and AND3 (N1094, N1074, N668, N159);
or OR2 (N1095, N1092, N900);
buf BUF1 (N1096, N1089);
nand NAND2 (N1097, N1059, N816);
xor XOR2 (N1098, N1095, N105);
not NOT1 (N1099, N1096);
nor NOR2 (N1100, N1093, N860);
or OR2 (N1101, N1082, N55);
or OR4 (N1102, N1094, N447, N1011, N614);
and AND3 (N1103, N1086, N57, N262);
nand NAND2 (N1104, N1098, N673);
not NOT1 (N1105, N1085);
xor XOR2 (N1106, N1102, N236);
nand NAND4 (N1107, N1097, N65, N774, N233);
and AND4 (N1108, N1088, N1055, N777, N1038);
or OR4 (N1109, N1099, N873, N137, N860);
not NOT1 (N1110, N1106);
buf BUF1 (N1111, N1104);
nand NAND4 (N1112, N1105, N842, N626, N673);
not NOT1 (N1113, N1108);
nor NOR4 (N1114, N1101, N310, N1095, N642);
not NOT1 (N1115, N1110);
or OR3 (N1116, N1115, N1028, N1010);
not NOT1 (N1117, N1107);
not NOT1 (N1118, N1114);
buf BUF1 (N1119, N1118);
or OR4 (N1120, N1111, N348, N310, N527);
and AND3 (N1121, N1116, N418, N67);
xor XOR2 (N1122, N1112, N1060);
or OR3 (N1123, N1119, N274, N123);
and AND2 (N1124, N1100, N1108);
not NOT1 (N1125, N1120);
and AND4 (N1126, N1121, N820, N537, N548);
and AND4 (N1127, N1091, N423, N111, N578);
or OR4 (N1128, N1123, N1083, N853, N768);
not NOT1 (N1129, N1113);
and AND3 (N1130, N1109, N391, N946);
not NOT1 (N1131, N1127);
xor XOR2 (N1132, N1130, N886);
nor NOR2 (N1133, N1124, N887);
and AND3 (N1134, N1126, N218, N560);
xor XOR2 (N1135, N1131, N1034);
and AND4 (N1136, N1125, N69, N234, N524);
and AND3 (N1137, N1134, N845, N178);
or OR4 (N1138, N1133, N440, N42, N907);
not NOT1 (N1139, N1137);
buf BUF1 (N1140, N1128);
not NOT1 (N1141, N1122);
not NOT1 (N1142, N1141);
nand NAND2 (N1143, N1135, N736);
and AND2 (N1144, N1129, N699);
buf BUF1 (N1145, N1136);
or OR2 (N1146, N1139, N1140);
xor XOR2 (N1147, N849, N233);
or OR2 (N1148, N1138, N544);
and AND4 (N1149, N1146, N64, N1136, N518);
and AND3 (N1150, N1143, N1082, N314);
nand NAND4 (N1151, N1150, N1102, N831, N300);
nand NAND2 (N1152, N1144, N94);
nor NOR3 (N1153, N1145, N985, N987);
nor NOR2 (N1154, N1103, N652);
buf BUF1 (N1155, N1148);
nor NOR4 (N1156, N1152, N192, N375, N594);
nand NAND3 (N1157, N1149, N721, N427);
nor NOR2 (N1158, N1156, N580);
not NOT1 (N1159, N1154);
nor NOR2 (N1160, N1153, N329);
and AND3 (N1161, N1132, N112, N1099);
xor XOR2 (N1162, N1160, N57);
xor XOR2 (N1163, N1161, N283);
and AND2 (N1164, N1142, N151);
and AND2 (N1165, N1155, N75);
nand NAND4 (N1166, N1165, N509, N763, N446);
or OR3 (N1167, N1157, N790, N514);
or OR4 (N1168, N1151, N822, N554, N151);
and AND3 (N1169, N1163, N176, N171);
xor XOR2 (N1170, N1164, N650);
buf BUF1 (N1171, N1167);
nor NOR3 (N1172, N1117, N514, N809);
xor XOR2 (N1173, N1171, N736);
not NOT1 (N1174, N1170);
not NOT1 (N1175, N1173);
nor NOR4 (N1176, N1168, N848, N504, N325);
buf BUF1 (N1177, N1174);
not NOT1 (N1178, N1166);
nand NAND2 (N1179, N1162, N923);
and AND3 (N1180, N1159, N232, N649);
and AND2 (N1181, N1178, N745);
nor NOR4 (N1182, N1169, N738, N379, N616);
or OR2 (N1183, N1172, N820);
nor NOR3 (N1184, N1181, N40, N697);
nor NOR4 (N1185, N1182, N940, N201, N639);
or OR3 (N1186, N1177, N165, N25);
nor NOR2 (N1187, N1186, N925);
xor XOR2 (N1188, N1179, N655);
or OR4 (N1189, N1183, N664, N60, N142);
nand NAND2 (N1190, N1176, N1062);
and AND4 (N1191, N1189, N165, N499, N966);
nor NOR2 (N1192, N1175, N1000);
or OR3 (N1193, N1147, N365, N109);
xor XOR2 (N1194, N1158, N1007);
xor XOR2 (N1195, N1180, N121);
and AND4 (N1196, N1190, N872, N619, N805);
or OR2 (N1197, N1188, N759);
and AND3 (N1198, N1191, N744, N847);
or OR3 (N1199, N1198, N944, N647);
or OR4 (N1200, N1196, N958, N476, N598);
and AND4 (N1201, N1194, N58, N1092, N197);
or OR3 (N1202, N1185, N356, N171);
and AND3 (N1203, N1201, N1013, N868);
or OR2 (N1204, N1187, N761);
and AND4 (N1205, N1197, N1063, N459, N164);
or OR2 (N1206, N1204, N379);
nor NOR2 (N1207, N1195, N932);
nor NOR4 (N1208, N1184, N235, N220, N306);
buf BUF1 (N1209, N1193);
and AND2 (N1210, N1199, N860);
nor NOR2 (N1211, N1205, N1088);
not NOT1 (N1212, N1209);
buf BUF1 (N1213, N1192);
nor NOR4 (N1214, N1206, N533, N482, N345);
or OR4 (N1215, N1213, N918, N611, N501);
not NOT1 (N1216, N1212);
xor XOR2 (N1217, N1200, N997);
buf BUF1 (N1218, N1214);
buf BUF1 (N1219, N1203);
not NOT1 (N1220, N1217);
or OR2 (N1221, N1211, N881);
not NOT1 (N1222, N1202);
nand NAND4 (N1223, N1207, N1124, N1090, N207);
xor XOR2 (N1224, N1218, N479);
nor NOR3 (N1225, N1208, N159, N644);
nor NOR4 (N1226, N1223, N443, N330, N1122);
nor NOR2 (N1227, N1220, N1193);
nand NAND3 (N1228, N1222, N1190, N395);
or OR4 (N1229, N1225, N758, N51, N201);
and AND2 (N1230, N1210, N569);
and AND4 (N1231, N1229, N1023, N26, N672);
buf BUF1 (N1232, N1227);
xor XOR2 (N1233, N1231, N189);
xor XOR2 (N1234, N1228, N864);
xor XOR2 (N1235, N1216, N1015);
nor NOR2 (N1236, N1226, N870);
nor NOR3 (N1237, N1234, N616, N238);
and AND3 (N1238, N1235, N1082, N999);
nand NAND4 (N1239, N1230, N463, N578, N612);
and AND4 (N1240, N1224, N700, N878, N1021);
nand NAND3 (N1241, N1240, N899, N1144);
buf BUF1 (N1242, N1233);
xor XOR2 (N1243, N1236, N623);
buf BUF1 (N1244, N1215);
nor NOR2 (N1245, N1241, N1104);
nand NAND3 (N1246, N1221, N1022, N535);
or OR3 (N1247, N1243, N709, N692);
buf BUF1 (N1248, N1237);
nand NAND2 (N1249, N1245, N602);
nor NOR3 (N1250, N1249, N433, N878);
buf BUF1 (N1251, N1238);
and AND3 (N1252, N1246, N521, N916);
and AND3 (N1253, N1250, N870, N242);
nand NAND4 (N1254, N1253, N1233, N1031, N92);
xor XOR2 (N1255, N1251, N507);
xor XOR2 (N1256, N1247, N1042);
and AND2 (N1257, N1255, N502);
not NOT1 (N1258, N1244);
not NOT1 (N1259, N1232);
nor NOR4 (N1260, N1239, N266, N5, N676);
nand NAND3 (N1261, N1260, N935, N38);
nand NAND4 (N1262, N1261, N94, N687, N1006);
not NOT1 (N1263, N1252);
xor XOR2 (N1264, N1263, N19);
xor XOR2 (N1265, N1259, N488);
and AND3 (N1266, N1258, N96, N684);
or OR3 (N1267, N1248, N1250, N802);
and AND3 (N1268, N1254, N832, N463);
nand NAND4 (N1269, N1267, N35, N312, N182);
nand NAND4 (N1270, N1262, N217, N1175, N1030);
nor NOR3 (N1271, N1269, N696, N404);
and AND3 (N1272, N1271, N1162, N142);
nor NOR3 (N1273, N1266, N3, N488);
not NOT1 (N1274, N1256);
xor XOR2 (N1275, N1274, N1067);
buf BUF1 (N1276, N1264);
or OR2 (N1277, N1273, N525);
not NOT1 (N1278, N1277);
xor XOR2 (N1279, N1242, N105);
and AND2 (N1280, N1270, N1121);
buf BUF1 (N1281, N1272);
or OR2 (N1282, N1265, N31);
not NOT1 (N1283, N1276);
and AND4 (N1284, N1279, N908, N9, N109);
nor NOR2 (N1285, N1275, N59);
or OR4 (N1286, N1281, N750, N1241, N409);
nor NOR2 (N1287, N1280, N843);
and AND3 (N1288, N1282, N35, N524);
or OR2 (N1289, N1268, N971);
buf BUF1 (N1290, N1285);
nand NAND2 (N1291, N1219, N366);
not NOT1 (N1292, N1278);
xor XOR2 (N1293, N1284, N781);
and AND4 (N1294, N1257, N102, N376, N1241);
nor NOR3 (N1295, N1287, N61, N1279);
nand NAND3 (N1296, N1283, N1091, N760);
and AND2 (N1297, N1294, N416);
nand NAND3 (N1298, N1295, N1163, N1097);
buf BUF1 (N1299, N1286);
buf BUF1 (N1300, N1298);
buf BUF1 (N1301, N1289);
nand NAND2 (N1302, N1288, N137);
nand NAND3 (N1303, N1300, N480, N883);
or OR4 (N1304, N1302, N895, N1015, N927);
nor NOR4 (N1305, N1301, N929, N367, N106);
or OR2 (N1306, N1305, N51);
nand NAND2 (N1307, N1293, N669);
nand NAND3 (N1308, N1299, N481, N995);
and AND3 (N1309, N1296, N495, N1159);
and AND2 (N1310, N1297, N850);
nor NOR2 (N1311, N1308, N1064);
nor NOR3 (N1312, N1291, N27, N1299);
or OR4 (N1313, N1304, N1199, N1215, N102);
and AND2 (N1314, N1307, N598);
not NOT1 (N1315, N1306);
nand NAND3 (N1316, N1303, N659, N369);
nor NOR2 (N1317, N1313, N1148);
nand NAND4 (N1318, N1309, N1034, N436, N1295);
or OR2 (N1319, N1312, N1037);
buf BUF1 (N1320, N1316);
xor XOR2 (N1321, N1310, N930);
nand NAND3 (N1322, N1321, N687, N645);
or OR4 (N1323, N1320, N18, N284, N341);
nor NOR4 (N1324, N1290, N481, N1314, N366);
xor XOR2 (N1325, N316, N703);
or OR4 (N1326, N1318, N584, N1208, N1282);
xor XOR2 (N1327, N1315, N729);
xor XOR2 (N1328, N1326, N1255);
not NOT1 (N1329, N1328);
or OR3 (N1330, N1323, N154, N384);
not NOT1 (N1331, N1311);
or OR2 (N1332, N1325, N278);
nand NAND2 (N1333, N1322, N375);
buf BUF1 (N1334, N1329);
buf BUF1 (N1335, N1330);
or OR3 (N1336, N1332, N1302, N207);
or OR2 (N1337, N1334, N194);
and AND3 (N1338, N1335, N727, N1124);
xor XOR2 (N1339, N1319, N1093);
nand NAND3 (N1340, N1333, N19, N952);
not NOT1 (N1341, N1340);
and AND4 (N1342, N1317, N765, N746, N175);
nor NOR3 (N1343, N1292, N1169, N783);
or OR2 (N1344, N1343, N338);
nand NAND3 (N1345, N1342, N423, N946);
xor XOR2 (N1346, N1327, N230);
nand NAND2 (N1347, N1331, N1143);
not NOT1 (N1348, N1339);
or OR3 (N1349, N1336, N633, N1337);
not NOT1 (N1350, N222);
buf BUF1 (N1351, N1349);
not NOT1 (N1352, N1345);
buf BUF1 (N1353, N1352);
nor NOR2 (N1354, N1347, N1232);
nor NOR2 (N1355, N1353, N97);
buf BUF1 (N1356, N1341);
buf BUF1 (N1357, N1344);
nor NOR2 (N1358, N1355, N1217);
buf BUF1 (N1359, N1338);
nand NAND2 (N1360, N1351, N631);
buf BUF1 (N1361, N1356);
xor XOR2 (N1362, N1348, N1208);
or OR3 (N1363, N1358, N479, N861);
and AND4 (N1364, N1361, N1114, N1174, N300);
buf BUF1 (N1365, N1360);
nor NOR4 (N1366, N1346, N579, N707, N191);
and AND2 (N1367, N1354, N474);
or OR3 (N1368, N1359, N437, N230);
nor NOR2 (N1369, N1357, N371);
xor XOR2 (N1370, N1368, N1187);
nand NAND2 (N1371, N1363, N698);
xor XOR2 (N1372, N1365, N1028);
nand NAND2 (N1373, N1364, N1285);
and AND3 (N1374, N1372, N964, N1197);
not NOT1 (N1375, N1362);
nand NAND3 (N1376, N1366, N1284, N643);
nor NOR3 (N1377, N1374, N1113, N1169);
nand NAND2 (N1378, N1369, N901);
xor XOR2 (N1379, N1376, N486);
xor XOR2 (N1380, N1373, N86);
buf BUF1 (N1381, N1371);
buf BUF1 (N1382, N1324);
or OR4 (N1383, N1382, N606, N899, N856);
and AND3 (N1384, N1367, N766, N1176);
nand NAND2 (N1385, N1380, N357);
not NOT1 (N1386, N1379);
nand NAND2 (N1387, N1383, N282);
and AND2 (N1388, N1381, N173);
buf BUF1 (N1389, N1378);
or OR2 (N1390, N1389, N157);
buf BUF1 (N1391, N1386);
nor NOR4 (N1392, N1390, N950, N1070, N935);
xor XOR2 (N1393, N1370, N249);
buf BUF1 (N1394, N1377);
not NOT1 (N1395, N1394);
and AND4 (N1396, N1385, N816, N176, N237);
xor XOR2 (N1397, N1388, N87);
xor XOR2 (N1398, N1393, N990);
or OR4 (N1399, N1395, N485, N1070, N433);
and AND4 (N1400, N1392, N1163, N560, N739);
buf BUF1 (N1401, N1375);
and AND4 (N1402, N1400, N976, N785, N881);
and AND4 (N1403, N1399, N139, N1004, N654);
and AND2 (N1404, N1403, N1219);
nor NOR3 (N1405, N1387, N494, N1206);
and AND4 (N1406, N1398, N745, N705, N1323);
or OR3 (N1407, N1397, N756, N16);
nand NAND2 (N1408, N1401, N610);
nand NAND4 (N1409, N1406, N580, N108, N873);
nor NOR4 (N1410, N1402, N276, N84, N109);
nor NOR2 (N1411, N1350, N1310);
nand NAND3 (N1412, N1411, N86, N1040);
nand NAND3 (N1413, N1410, N568, N215);
or OR2 (N1414, N1407, N1270);
xor XOR2 (N1415, N1412, N959);
nor NOR3 (N1416, N1391, N155, N1089);
nor NOR3 (N1417, N1408, N924, N7);
buf BUF1 (N1418, N1414);
and AND4 (N1419, N1418, N21, N544, N819);
nor NOR3 (N1420, N1409, N59, N618);
nand NAND3 (N1421, N1419, N360, N1012);
xor XOR2 (N1422, N1396, N1009);
and AND3 (N1423, N1413, N616, N188);
nand NAND3 (N1424, N1405, N190, N561);
xor XOR2 (N1425, N1424, N196);
not NOT1 (N1426, N1384);
buf BUF1 (N1427, N1420);
xor XOR2 (N1428, N1423, N23);
and AND3 (N1429, N1416, N116, N233);
buf BUF1 (N1430, N1428);
not NOT1 (N1431, N1415);
xor XOR2 (N1432, N1429, N728);
not NOT1 (N1433, N1421);
xor XOR2 (N1434, N1404, N22);
nand NAND4 (N1435, N1430, N947, N315, N204);
or OR3 (N1436, N1432, N415, N229);
xor XOR2 (N1437, N1425, N197);
or OR3 (N1438, N1436, N631, N51);
buf BUF1 (N1439, N1427);
buf BUF1 (N1440, N1437);
xor XOR2 (N1441, N1439, N469);
not NOT1 (N1442, N1438);
nand NAND4 (N1443, N1422, N919, N242, N208);
buf BUF1 (N1444, N1426);
nand NAND2 (N1445, N1443, N1383);
not NOT1 (N1446, N1434);
not NOT1 (N1447, N1445);
or OR3 (N1448, N1417, N653, N621);
buf BUF1 (N1449, N1444);
buf BUF1 (N1450, N1433);
xor XOR2 (N1451, N1441, N760);
or OR4 (N1452, N1440, N36, N619, N221);
or OR2 (N1453, N1448, N918);
nand NAND4 (N1454, N1449, N896, N1409, N998);
nor NOR4 (N1455, N1452, N853, N544, N1188);
xor XOR2 (N1456, N1453, N974);
and AND2 (N1457, N1456, N1126);
not NOT1 (N1458, N1451);
buf BUF1 (N1459, N1450);
not NOT1 (N1460, N1447);
not NOT1 (N1461, N1457);
nand NAND4 (N1462, N1460, N1245, N233, N1044);
or OR3 (N1463, N1458, N263, N247);
buf BUF1 (N1464, N1454);
and AND4 (N1465, N1461, N907, N1055, N723);
not NOT1 (N1466, N1465);
nor NOR4 (N1467, N1463, N1042, N705, N1398);
nor NOR3 (N1468, N1431, N102, N313);
nand NAND4 (N1469, N1462, N185, N975, N99);
and AND4 (N1470, N1459, N220, N671, N701);
not NOT1 (N1471, N1468);
nor NOR2 (N1472, N1455, N1075);
and AND4 (N1473, N1469, N772, N215, N422);
nor NOR3 (N1474, N1446, N64, N1065);
nand NAND2 (N1475, N1464, N414);
buf BUF1 (N1476, N1475);
buf BUF1 (N1477, N1474);
nor NOR3 (N1478, N1466, N544, N662);
buf BUF1 (N1479, N1470);
not NOT1 (N1480, N1473);
or OR4 (N1481, N1472, N718, N623, N1260);
xor XOR2 (N1482, N1442, N1415);
not NOT1 (N1483, N1477);
nor NOR4 (N1484, N1482, N11, N861, N253);
buf BUF1 (N1485, N1478);
nand NAND4 (N1486, N1435, N990, N18, N1372);
buf BUF1 (N1487, N1481);
buf BUF1 (N1488, N1485);
and AND2 (N1489, N1471, N1344);
xor XOR2 (N1490, N1483, N738);
and AND2 (N1491, N1487, N1436);
nand NAND3 (N1492, N1490, N311, N1337);
xor XOR2 (N1493, N1479, N766);
and AND4 (N1494, N1489, N679, N227, N855);
not NOT1 (N1495, N1493);
not NOT1 (N1496, N1476);
xor XOR2 (N1497, N1495, N1426);
nor NOR3 (N1498, N1484, N59, N1147);
nand NAND2 (N1499, N1486, N1187);
nor NOR3 (N1500, N1492, N264, N320);
or OR2 (N1501, N1496, N1308);
nor NOR3 (N1502, N1500, N166, N105);
and AND2 (N1503, N1502, N1469);
xor XOR2 (N1504, N1501, N732);
xor XOR2 (N1505, N1499, N846);
or OR4 (N1506, N1467, N774, N1443, N150);
buf BUF1 (N1507, N1503);
and AND3 (N1508, N1491, N1483, N1368);
buf BUF1 (N1509, N1504);
buf BUF1 (N1510, N1508);
nor NOR3 (N1511, N1510, N526, N566);
xor XOR2 (N1512, N1511, N312);
nor NOR2 (N1513, N1497, N1347);
or OR3 (N1514, N1506, N1044, N597);
or OR4 (N1515, N1480, N970, N708, N1336);
buf BUF1 (N1516, N1505);
or OR4 (N1517, N1498, N251, N890, N966);
xor XOR2 (N1518, N1512, N1397);
nor NOR4 (N1519, N1488, N57, N1250, N1084);
and AND4 (N1520, N1507, N536, N775, N79);
nand NAND2 (N1521, N1517, N809);
xor XOR2 (N1522, N1494, N502);
not NOT1 (N1523, N1518);
or OR3 (N1524, N1515, N1389, N1100);
or OR2 (N1525, N1516, N431);
and AND4 (N1526, N1519, N133, N1319, N1182);
or OR4 (N1527, N1523, N833, N591, N309);
and AND3 (N1528, N1520, N1073, N1152);
nand NAND2 (N1529, N1528, N1461);
buf BUF1 (N1530, N1524);
xor XOR2 (N1531, N1522, N507);
not NOT1 (N1532, N1514);
not NOT1 (N1533, N1521);
nand NAND2 (N1534, N1530, N1201);
nand NAND2 (N1535, N1531, N548);
not NOT1 (N1536, N1529);
not NOT1 (N1537, N1533);
or OR2 (N1538, N1534, N485);
nand NAND3 (N1539, N1535, N735, N604);
nor NOR4 (N1540, N1513, N1168, N556, N1267);
nand NAND3 (N1541, N1536, N776, N1434);
xor XOR2 (N1542, N1509, N1395);
nor NOR4 (N1543, N1525, N256, N1521, N277);
and AND4 (N1544, N1542, N86, N238, N1066);
or OR2 (N1545, N1532, N1497);
nor NOR4 (N1546, N1538, N1179, N100, N1487);
xor XOR2 (N1547, N1526, N192);
not NOT1 (N1548, N1544);
xor XOR2 (N1549, N1541, N799);
and AND3 (N1550, N1546, N1453, N1163);
and AND4 (N1551, N1548, N42, N708, N353);
and AND4 (N1552, N1539, N537, N1530, N1435);
xor XOR2 (N1553, N1543, N12);
not NOT1 (N1554, N1553);
nor NOR4 (N1555, N1551, N1297, N1421, N156);
and AND3 (N1556, N1527, N468, N947);
and AND2 (N1557, N1555, N1508);
or OR3 (N1558, N1557, N1076, N1100);
or OR3 (N1559, N1545, N1005, N1541);
or OR3 (N1560, N1552, N693, N93);
buf BUF1 (N1561, N1554);
xor XOR2 (N1562, N1559, N34);
buf BUF1 (N1563, N1540);
nor NOR3 (N1564, N1558, N268, N1371);
and AND2 (N1565, N1561, N774);
nand NAND2 (N1566, N1556, N1560);
nor NOR4 (N1567, N1257, N988, N404, N840);
not NOT1 (N1568, N1565);
nor NOR4 (N1569, N1562, N1369, N328, N1499);
nand NAND4 (N1570, N1547, N1105, N230, N38);
not NOT1 (N1571, N1569);
nor NOR4 (N1572, N1550, N1484, N572, N84);
xor XOR2 (N1573, N1572, N986);
buf BUF1 (N1574, N1567);
or OR3 (N1575, N1564, N1160, N876);
buf BUF1 (N1576, N1537);
buf BUF1 (N1577, N1575);
xor XOR2 (N1578, N1566, N1568);
buf BUF1 (N1579, N1335);
and AND3 (N1580, N1563, N884, N1058);
and AND3 (N1581, N1579, N1201, N1411);
buf BUF1 (N1582, N1571);
or OR4 (N1583, N1570, N689, N1503, N673);
and AND2 (N1584, N1577, N1343);
nor NOR4 (N1585, N1583, N1563, N1256, N1118);
xor XOR2 (N1586, N1576, N1571);
nand NAND3 (N1587, N1574, N1306, N68);
and AND4 (N1588, N1586, N881, N766, N1381);
nor NOR3 (N1589, N1584, N1179, N566);
nand NAND4 (N1590, N1587, N94, N982, N118);
xor XOR2 (N1591, N1588, N1453);
not NOT1 (N1592, N1591);
nor NOR4 (N1593, N1549, N1202, N975, N120);
and AND2 (N1594, N1580, N287);
or OR3 (N1595, N1592, N1243, N1538);
xor XOR2 (N1596, N1578, N1357);
and AND3 (N1597, N1582, N259, N1274);
nor NOR2 (N1598, N1596, N480);
nand NAND3 (N1599, N1598, N1283, N861);
nor NOR3 (N1600, N1573, N849, N741);
and AND3 (N1601, N1590, N237, N317);
buf BUF1 (N1602, N1601);
nand NAND4 (N1603, N1593, N777, N1406, N1166);
xor XOR2 (N1604, N1589, N475);
nand NAND4 (N1605, N1603, N1376, N1437, N650);
not NOT1 (N1606, N1599);
xor XOR2 (N1607, N1606, N706);
buf BUF1 (N1608, N1594);
and AND2 (N1609, N1595, N1463);
xor XOR2 (N1610, N1607, N1467);
nor NOR4 (N1611, N1602, N839, N596, N1296);
not NOT1 (N1612, N1604);
xor XOR2 (N1613, N1610, N97);
and AND4 (N1614, N1611, N1369, N1132, N1425);
nand NAND4 (N1615, N1614, N799, N1156, N507);
or OR2 (N1616, N1600, N687);
not NOT1 (N1617, N1609);
not NOT1 (N1618, N1617);
or OR3 (N1619, N1618, N602, N996);
xor XOR2 (N1620, N1581, N1075);
or OR3 (N1621, N1585, N868, N539);
buf BUF1 (N1622, N1616);
or OR3 (N1623, N1597, N1242, N87);
or OR2 (N1624, N1613, N591);
xor XOR2 (N1625, N1622, N965);
and AND2 (N1626, N1621, N518);
nor NOR4 (N1627, N1612, N788, N1194, N588);
or OR4 (N1628, N1624, N1129, N1553, N1198);
and AND4 (N1629, N1619, N887, N1286, N68);
and AND2 (N1630, N1608, N101);
not NOT1 (N1631, N1630);
or OR4 (N1632, N1605, N1095, N500, N269);
nor NOR3 (N1633, N1632, N1176, N1491);
not NOT1 (N1634, N1629);
or OR2 (N1635, N1615, N1010);
nand NAND3 (N1636, N1633, N812, N1381);
not NOT1 (N1637, N1620);
or OR2 (N1638, N1627, N1323);
nand NAND2 (N1639, N1626, N167);
nor NOR3 (N1640, N1625, N1490, N579);
nand NAND2 (N1641, N1638, N1286);
or OR3 (N1642, N1636, N1419, N1363);
nor NOR2 (N1643, N1635, N734);
xor XOR2 (N1644, N1640, N481);
nand NAND2 (N1645, N1639, N560);
xor XOR2 (N1646, N1634, N1174);
and AND4 (N1647, N1642, N116, N763, N1332);
or OR3 (N1648, N1623, N245, N847);
and AND3 (N1649, N1631, N267, N450);
xor XOR2 (N1650, N1646, N1489);
buf BUF1 (N1651, N1637);
and AND4 (N1652, N1650, N106, N104, N14);
nand NAND3 (N1653, N1628, N1001, N1375);
nand NAND4 (N1654, N1649, N544, N687, N1363);
xor XOR2 (N1655, N1654, N215);
nand NAND2 (N1656, N1647, N620);
nand NAND4 (N1657, N1648, N610, N1314, N1612);
and AND2 (N1658, N1641, N596);
buf BUF1 (N1659, N1643);
nor NOR2 (N1660, N1658, N104);
or OR2 (N1661, N1645, N215);
xor XOR2 (N1662, N1661, N591);
and AND4 (N1663, N1660, N375, N1627, N255);
or OR2 (N1664, N1652, N660);
and AND3 (N1665, N1664, N75, N1335);
nand NAND4 (N1666, N1663, N623, N486, N361);
xor XOR2 (N1667, N1655, N634);
nor NOR4 (N1668, N1651, N547, N1409, N1656);
or OR3 (N1669, N832, N247, N1207);
nand NAND4 (N1670, N1653, N479, N145, N1467);
nor NOR4 (N1671, N1668, N233, N689, N786);
buf BUF1 (N1672, N1666);
buf BUF1 (N1673, N1667);
xor XOR2 (N1674, N1657, N1215);
nor NOR4 (N1675, N1670, N1067, N165, N1435);
or OR2 (N1676, N1659, N345);
buf BUF1 (N1677, N1672);
not NOT1 (N1678, N1665);
nand NAND4 (N1679, N1669, N816, N1469, N1170);
not NOT1 (N1680, N1644);
buf BUF1 (N1681, N1673);
or OR4 (N1682, N1681, N382, N1370, N1122);
not NOT1 (N1683, N1679);
not NOT1 (N1684, N1682);
xor XOR2 (N1685, N1674, N841);
nor NOR2 (N1686, N1677, N699);
nand NAND3 (N1687, N1683, N1041, N1685);
buf BUF1 (N1688, N252);
nand NAND4 (N1689, N1676, N1620, N668, N924);
or OR2 (N1690, N1686, N1129);
and AND2 (N1691, N1671, N1585);
buf BUF1 (N1692, N1691);
nor NOR3 (N1693, N1692, N1683, N1322);
not NOT1 (N1694, N1662);
buf BUF1 (N1695, N1689);
xor XOR2 (N1696, N1694, N843);
nand NAND3 (N1697, N1688, N20, N268);
and AND3 (N1698, N1680, N1231, N1172);
and AND2 (N1699, N1675, N1429);
or OR4 (N1700, N1690, N1068, N605, N865);
or OR2 (N1701, N1699, N529);
xor XOR2 (N1702, N1693, N1221);
nand NAND4 (N1703, N1696, N38, N1465, N1410);
xor XOR2 (N1704, N1687, N1328);
nand NAND2 (N1705, N1702, N888);
xor XOR2 (N1706, N1698, N718);
nor NOR3 (N1707, N1700, N1493, N142);
nand NAND3 (N1708, N1704, N641, N330);
and AND4 (N1709, N1708, N23, N59, N503);
not NOT1 (N1710, N1707);
nand NAND4 (N1711, N1701, N800, N986, N531);
not NOT1 (N1712, N1697);
not NOT1 (N1713, N1678);
and AND3 (N1714, N1695, N1636, N653);
xor XOR2 (N1715, N1684, N800);
or OR3 (N1716, N1706, N324, N1074);
xor XOR2 (N1717, N1716, N943);
nand NAND3 (N1718, N1705, N979, N1438);
nand NAND4 (N1719, N1712, N82, N1009, N1198);
buf BUF1 (N1720, N1717);
nor NOR2 (N1721, N1713, N300);
xor XOR2 (N1722, N1710, N1354);
xor XOR2 (N1723, N1711, N1708);
nor NOR2 (N1724, N1718, N189);
and AND3 (N1725, N1722, N802, N505);
buf BUF1 (N1726, N1723);
not NOT1 (N1727, N1709);
and AND3 (N1728, N1724, N256, N137);
and AND4 (N1729, N1720, N904, N1628, N1370);
and AND3 (N1730, N1719, N1139, N58);
nand NAND4 (N1731, N1726, N177, N914, N1563);
nor NOR4 (N1732, N1721, N1443, N523, N203);
buf BUF1 (N1733, N1727);
or OR3 (N1734, N1732, N79, N196);
or OR2 (N1735, N1714, N990);
and AND2 (N1736, N1703, N273);
not NOT1 (N1737, N1733);
buf BUF1 (N1738, N1729);
xor XOR2 (N1739, N1736, N1299);
nor NOR3 (N1740, N1735, N1631, N1099);
buf BUF1 (N1741, N1740);
buf BUF1 (N1742, N1715);
or OR4 (N1743, N1737, N1375, N789, N219);
not NOT1 (N1744, N1731);
xor XOR2 (N1745, N1728, N410);
not NOT1 (N1746, N1743);
buf BUF1 (N1747, N1746);
and AND2 (N1748, N1725, N97);
not NOT1 (N1749, N1739);
not NOT1 (N1750, N1745);
nand NAND2 (N1751, N1747, N748);
xor XOR2 (N1752, N1750, N1279);
not NOT1 (N1753, N1748);
buf BUF1 (N1754, N1742);
buf BUF1 (N1755, N1753);
nor NOR2 (N1756, N1730, N287);
nand NAND2 (N1757, N1754, N50);
and AND4 (N1758, N1744, N186, N1054, N608);
xor XOR2 (N1759, N1758, N1382);
buf BUF1 (N1760, N1751);
xor XOR2 (N1761, N1757, N1627);
buf BUF1 (N1762, N1734);
and AND3 (N1763, N1752, N539, N658);
xor XOR2 (N1764, N1738, N1679);
nand NAND2 (N1765, N1761, N1392);
nand NAND2 (N1766, N1762, N242);
buf BUF1 (N1767, N1749);
or OR2 (N1768, N1741, N649);
xor XOR2 (N1769, N1766, N109);
not NOT1 (N1770, N1759);
nand NAND3 (N1771, N1770, N959, N674);
nor NOR2 (N1772, N1771, N600);
or OR4 (N1773, N1769, N900, N1108, N285);
xor XOR2 (N1774, N1763, N1480);
nor NOR4 (N1775, N1772, N148, N811, N1543);
or OR3 (N1776, N1765, N402, N165);
or OR3 (N1777, N1760, N107, N499);
nand NAND3 (N1778, N1773, N741, N696);
nor NOR2 (N1779, N1775, N304);
nor NOR2 (N1780, N1768, N422);
and AND4 (N1781, N1774, N1514, N1008, N414);
nand NAND4 (N1782, N1779, N274, N1745, N1714);
nor NOR4 (N1783, N1756, N516, N1566, N366);
nor NOR3 (N1784, N1776, N377, N1737);
not NOT1 (N1785, N1767);
and AND3 (N1786, N1755, N213, N1506);
not NOT1 (N1787, N1784);
nand NAND4 (N1788, N1780, N1472, N714, N948);
buf BUF1 (N1789, N1787);
xor XOR2 (N1790, N1781, N1326);
buf BUF1 (N1791, N1777);
nand NAND3 (N1792, N1782, N1273, N1128);
nor NOR3 (N1793, N1786, N340, N119);
buf BUF1 (N1794, N1783);
nand NAND2 (N1795, N1785, N1734);
nor NOR2 (N1796, N1791, N488);
buf BUF1 (N1797, N1796);
not NOT1 (N1798, N1793);
buf BUF1 (N1799, N1764);
not NOT1 (N1800, N1795);
buf BUF1 (N1801, N1797);
not NOT1 (N1802, N1788);
not NOT1 (N1803, N1801);
nor NOR3 (N1804, N1803, N738, N1408);
and AND4 (N1805, N1778, N298, N608, N828);
nor NOR4 (N1806, N1800, N1726, N579, N369);
nor NOR2 (N1807, N1790, N1061);
buf BUF1 (N1808, N1804);
nand NAND4 (N1809, N1789, N1306, N957, N906);
nor NOR3 (N1810, N1798, N1280, N1197);
nand NAND2 (N1811, N1806, N316);
or OR4 (N1812, N1802, N504, N1077, N331);
xor XOR2 (N1813, N1811, N1103);
buf BUF1 (N1814, N1807);
not NOT1 (N1815, N1794);
nand NAND4 (N1816, N1792, N434, N1053, N1056);
xor XOR2 (N1817, N1810, N303);
nand NAND2 (N1818, N1815, N1150);
and AND4 (N1819, N1816, N515, N369, N932);
and AND3 (N1820, N1808, N1040, N227);
buf BUF1 (N1821, N1817);
buf BUF1 (N1822, N1809);
not NOT1 (N1823, N1822);
xor XOR2 (N1824, N1814, N127);
not NOT1 (N1825, N1823);
not NOT1 (N1826, N1813);
not NOT1 (N1827, N1824);
nand NAND2 (N1828, N1805, N1414);
and AND3 (N1829, N1820, N1509, N1767);
buf BUF1 (N1830, N1818);
and AND3 (N1831, N1828, N832, N735);
nor NOR3 (N1832, N1825, N209, N1602);
nand NAND4 (N1833, N1799, N1341, N1680, N582);
not NOT1 (N1834, N1833);
nand NAND2 (N1835, N1827, N165);
or OR3 (N1836, N1826, N1517, N1369);
not NOT1 (N1837, N1829);
and AND3 (N1838, N1821, N1388, N916);
nor NOR3 (N1839, N1836, N829, N164);
nand NAND3 (N1840, N1832, N593, N748);
xor XOR2 (N1841, N1831, N1028);
nor NOR2 (N1842, N1835, N1555);
and AND4 (N1843, N1838, N168, N84, N637);
nor NOR3 (N1844, N1837, N636, N1727);
nand NAND3 (N1845, N1839, N1663, N130);
or OR4 (N1846, N1830, N1308, N166, N358);
and AND2 (N1847, N1846, N622);
or OR2 (N1848, N1841, N24);
not NOT1 (N1849, N1812);
or OR4 (N1850, N1834, N324, N1631, N1155);
buf BUF1 (N1851, N1840);
nand NAND2 (N1852, N1842, N916);
xor XOR2 (N1853, N1844, N10);
and AND3 (N1854, N1851, N580, N1106);
not NOT1 (N1855, N1845);
and AND3 (N1856, N1852, N1583, N960);
nor NOR2 (N1857, N1819, N259);
and AND2 (N1858, N1855, N1067);
xor XOR2 (N1859, N1850, N160);
nor NOR4 (N1860, N1859, N57, N1096, N1158);
and AND3 (N1861, N1843, N1647, N701);
nor NOR4 (N1862, N1848, N107, N382, N277);
not NOT1 (N1863, N1861);
buf BUF1 (N1864, N1856);
and AND4 (N1865, N1864, N746, N1202, N1525);
nor NOR2 (N1866, N1858, N1783);
and AND3 (N1867, N1847, N195, N511);
or OR3 (N1868, N1862, N1228, N1284);
xor XOR2 (N1869, N1868, N979);
or OR2 (N1870, N1863, N1148);
nand NAND3 (N1871, N1866, N1812, N1732);
or OR4 (N1872, N1870, N1508, N655, N888);
buf BUF1 (N1873, N1871);
and AND4 (N1874, N1869, N280, N775, N1451);
or OR2 (N1875, N1853, N46);
not NOT1 (N1876, N1849);
not NOT1 (N1877, N1875);
and AND4 (N1878, N1865, N895, N569, N94);
nand NAND4 (N1879, N1874, N441, N1650, N1302);
xor XOR2 (N1880, N1867, N832);
and AND4 (N1881, N1854, N729, N1679, N1305);
or OR3 (N1882, N1876, N233, N435);
nor NOR2 (N1883, N1882, N1592);
buf BUF1 (N1884, N1879);
buf BUF1 (N1885, N1880);
buf BUF1 (N1886, N1884);
not NOT1 (N1887, N1860);
not NOT1 (N1888, N1872);
not NOT1 (N1889, N1877);
not NOT1 (N1890, N1886);
buf BUF1 (N1891, N1890);
xor XOR2 (N1892, N1878, N1531);
xor XOR2 (N1893, N1887, N261);
nand NAND4 (N1894, N1881, N100, N1184, N1778);
nor NOR3 (N1895, N1885, N186, N393);
buf BUF1 (N1896, N1894);
nor NOR4 (N1897, N1888, N728, N1598, N1875);
buf BUF1 (N1898, N1873);
nand NAND3 (N1899, N1898, N797, N1321);
not NOT1 (N1900, N1889);
buf BUF1 (N1901, N1857);
and AND3 (N1902, N1901, N134, N1554);
xor XOR2 (N1903, N1899, N92);
or OR4 (N1904, N1900, N1847, N530, N1613);
and AND4 (N1905, N1904, N1004, N573, N1058);
nor NOR3 (N1906, N1895, N1138, N668);
buf BUF1 (N1907, N1897);
or OR3 (N1908, N1906, N1833, N139);
not NOT1 (N1909, N1905);
nor NOR2 (N1910, N1902, N1007);
nand NAND4 (N1911, N1908, N627, N1080, N1804);
or OR2 (N1912, N1911, N762);
nand NAND2 (N1913, N1909, N795);
xor XOR2 (N1914, N1896, N1595);
not NOT1 (N1915, N1892);
not NOT1 (N1916, N1912);
buf BUF1 (N1917, N1910);
xor XOR2 (N1918, N1893, N1502);
not NOT1 (N1919, N1907);
or OR4 (N1920, N1903, N433, N360, N70);
or OR4 (N1921, N1919, N172, N1286, N427);
nor NOR2 (N1922, N1883, N1063);
and AND3 (N1923, N1917, N770, N692);
nor NOR4 (N1924, N1914, N805, N816, N1029);
nand NAND3 (N1925, N1924, N1075, N602);
nand NAND3 (N1926, N1920, N389, N393);
buf BUF1 (N1927, N1915);
or OR3 (N1928, N1922, N1414, N1646);
nor NOR3 (N1929, N1921, N1662, N1655);
nor NOR3 (N1930, N1927, N836, N1609);
nor NOR4 (N1931, N1926, N74, N104, N883);
xor XOR2 (N1932, N1930, N834);
not NOT1 (N1933, N1929);
buf BUF1 (N1934, N1923);
or OR3 (N1935, N1891, N350, N1660);
not NOT1 (N1936, N1925);
xor XOR2 (N1937, N1936, N1492);
or OR4 (N1938, N1928, N1695, N957, N1644);
buf BUF1 (N1939, N1916);
nand NAND3 (N1940, N1918, N1019, N257);
xor XOR2 (N1941, N1933, N1309);
xor XOR2 (N1942, N1941, N1918);
and AND2 (N1943, N1939, N68);
buf BUF1 (N1944, N1937);
not NOT1 (N1945, N1944);
nor NOR2 (N1946, N1913, N1643);
not NOT1 (N1947, N1942);
nor NOR4 (N1948, N1932, N1713, N5, N1300);
buf BUF1 (N1949, N1938);
and AND2 (N1950, N1940, N1135);
xor XOR2 (N1951, N1935, N1377);
and AND3 (N1952, N1949, N725, N1230);
xor XOR2 (N1953, N1934, N2);
and AND4 (N1954, N1931, N1676, N177, N1756);
xor XOR2 (N1955, N1950, N815);
buf BUF1 (N1956, N1948);
not NOT1 (N1957, N1954);
or OR4 (N1958, N1951, N753, N1629, N1597);
or OR4 (N1959, N1955, N217, N1767, N682);
buf BUF1 (N1960, N1947);
xor XOR2 (N1961, N1960, N1514);
not NOT1 (N1962, N1958);
not NOT1 (N1963, N1945);
buf BUF1 (N1964, N1961);
buf BUF1 (N1965, N1964);
xor XOR2 (N1966, N1956, N583);
nand NAND2 (N1967, N1952, N901);
nor NOR4 (N1968, N1963, N1500, N1826, N642);
xor XOR2 (N1969, N1965, N1329);
nand NAND2 (N1970, N1957, N1477);
not NOT1 (N1971, N1970);
nor NOR4 (N1972, N1946, N1028, N1413, N1970);
or OR4 (N1973, N1971, N977, N1307, N1078);
or OR2 (N1974, N1966, N1418);
xor XOR2 (N1975, N1968, N1812);
or OR3 (N1976, N1973, N661, N1502);
nand NAND2 (N1977, N1962, N1334);
nand NAND4 (N1978, N1967, N1514, N1324, N41);
not NOT1 (N1979, N1976);
buf BUF1 (N1980, N1953);
buf BUF1 (N1981, N1978);
nand NAND4 (N1982, N1977, N1243, N1781, N366);
not NOT1 (N1983, N1969);
nand NAND4 (N1984, N1959, N753, N333, N1436);
nand NAND2 (N1985, N1980, N515);
buf BUF1 (N1986, N1984);
nor NOR3 (N1987, N1986, N249, N513);
and AND2 (N1988, N1985, N1350);
nor NOR2 (N1989, N1943, N765);
and AND4 (N1990, N1988, N1740, N582, N1940);
nor NOR3 (N1991, N1981, N1861, N706);
buf BUF1 (N1992, N1979);
and AND4 (N1993, N1992, N1066, N1327, N1841);
nor NOR2 (N1994, N1990, N617);
not NOT1 (N1995, N1983);
and AND2 (N1996, N1972, N1001);
buf BUF1 (N1997, N1987);
nand NAND2 (N1998, N1974, N1097);
buf BUF1 (N1999, N1994);
xor XOR2 (N2000, N1995, N1339);
nand NAND4 (N2001, N1998, N937, N1892, N1872);
xor XOR2 (N2002, N1996, N1081);
not NOT1 (N2003, N2000);
nor NOR2 (N2004, N1993, N1789);
nor NOR2 (N2005, N2002, N1175);
nor NOR2 (N2006, N2001, N722);
nor NOR4 (N2007, N1982, N1356, N936, N184);
nor NOR4 (N2008, N2006, N453, N444, N1092);
and AND3 (N2009, N2005, N291, N1464);
buf BUF1 (N2010, N2003);
xor XOR2 (N2011, N2004, N640);
buf BUF1 (N2012, N2011);
xor XOR2 (N2013, N2012, N1768);
and AND3 (N2014, N1997, N389, N1556);
buf BUF1 (N2015, N2009);
and AND4 (N2016, N2008, N571, N1345, N245);
xor XOR2 (N2017, N2010, N1432);
and AND3 (N2018, N2015, N1275, N893);
buf BUF1 (N2019, N2017);
nand NAND4 (N2020, N2013, N19, N1764, N712);
not NOT1 (N2021, N2007);
not NOT1 (N2022, N2018);
or OR4 (N2023, N1989, N776, N188, N1040);
and AND4 (N2024, N1991, N1563, N1121, N1869);
or OR4 (N2025, N2016, N1778, N778, N1246);
or OR3 (N2026, N2025, N1997, N1243);
nor NOR3 (N2027, N2020, N958, N1902);
xor XOR2 (N2028, N2026, N1221);
not NOT1 (N2029, N2024);
not NOT1 (N2030, N2021);
and AND2 (N2031, N2023, N929);
nand NAND2 (N2032, N2027, N1568);
xor XOR2 (N2033, N2014, N1341);
and AND3 (N2034, N2031, N405, N172);
nand NAND3 (N2035, N1975, N1724, N1792);
or OR4 (N2036, N2030, N545, N1033, N295);
and AND3 (N2037, N2034, N721, N1871);
xor XOR2 (N2038, N2036, N1553);
or OR3 (N2039, N2033, N472, N2036);
buf BUF1 (N2040, N2037);
or OR3 (N2041, N2039, N77, N1666);
buf BUF1 (N2042, N2035);
xor XOR2 (N2043, N2019, N392);
buf BUF1 (N2044, N2043);
xor XOR2 (N2045, N2032, N1445);
not NOT1 (N2046, N1999);
xor XOR2 (N2047, N2038, N1918);
nor NOR4 (N2048, N2046, N789, N1050, N966);
or OR2 (N2049, N2022, N1388);
or OR3 (N2050, N2044, N660, N1758);
or OR3 (N2051, N2045, N777, N18);
not NOT1 (N2052, N2029);
or OR4 (N2053, N2051, N463, N232, N278);
not NOT1 (N2054, N2040);
not NOT1 (N2055, N2054);
nor NOR2 (N2056, N2048, N612);
nand NAND3 (N2057, N2055, N315, N181);
or OR3 (N2058, N2050, N1712, N1733);
and AND3 (N2059, N2058, N1836, N1707);
not NOT1 (N2060, N2028);
and AND3 (N2061, N2041, N279, N815);
nand NAND2 (N2062, N2061, N1487);
nor NOR3 (N2063, N2047, N1962, N897);
nand NAND3 (N2064, N2062, N250, N1407);
nor NOR2 (N2065, N2049, N1982);
not NOT1 (N2066, N2059);
or OR3 (N2067, N2063, N1996, N1067);
nand NAND4 (N2068, N2064, N35, N1778, N681);
and AND2 (N2069, N2066, N1341);
or OR4 (N2070, N2057, N2049, N1380, N560);
not NOT1 (N2071, N2053);
xor XOR2 (N2072, N2067, N1429);
nand NAND3 (N2073, N2052, N1114, N1586);
nand NAND2 (N2074, N2060, N1821);
nand NAND2 (N2075, N2069, N1874);
buf BUF1 (N2076, N2075);
and AND4 (N2077, N2072, N477, N1592, N1520);
buf BUF1 (N2078, N2071);
not NOT1 (N2079, N2042);
and AND4 (N2080, N2070, N1352, N366, N1520);
not NOT1 (N2081, N2065);
nand NAND2 (N2082, N2073, N683);
or OR3 (N2083, N2079, N1976, N2009);
nand NAND3 (N2084, N2076, N807, N344);
xor XOR2 (N2085, N2074, N804);
and AND2 (N2086, N2056, N186);
not NOT1 (N2087, N2081);
and AND4 (N2088, N2080, N1606, N1673, N393);
and AND3 (N2089, N2083, N269, N97);
buf BUF1 (N2090, N2087);
nor NOR2 (N2091, N2078, N1368);
or OR3 (N2092, N2088, N1185, N213);
or OR3 (N2093, N2068, N3, N854);
xor XOR2 (N2094, N2093, N1456);
nand NAND3 (N2095, N2091, N56, N1725);
xor XOR2 (N2096, N2090, N987);
nand NAND2 (N2097, N2089, N1820);
not NOT1 (N2098, N2095);
or OR4 (N2099, N2097, N932, N805, N803);
buf BUF1 (N2100, N2098);
or OR4 (N2101, N2099, N1952, N474, N907);
nor NOR3 (N2102, N2100, N489, N782);
or OR4 (N2103, N2094, N1097, N2047, N2048);
or OR2 (N2104, N2084, N1776);
buf BUF1 (N2105, N2086);
xor XOR2 (N2106, N2104, N1024);
nand NAND2 (N2107, N2101, N393);
nand NAND3 (N2108, N2106, N32, N2007);
or OR2 (N2109, N2108, N1130);
not NOT1 (N2110, N2092);
and AND4 (N2111, N2110, N1399, N1208, N1052);
nor NOR3 (N2112, N2085, N101, N659);
nor NOR3 (N2113, N2102, N550, N1617);
not NOT1 (N2114, N2109);
or OR3 (N2115, N2113, N2022, N697);
and AND2 (N2116, N2111, N1244);
and AND3 (N2117, N2114, N859, N2005);
xor XOR2 (N2118, N2105, N730);
nand NAND3 (N2119, N2117, N1341, N1725);
buf BUF1 (N2120, N2116);
and AND3 (N2121, N2082, N1263, N622);
nor NOR4 (N2122, N2121, N1638, N1917, N186);
buf BUF1 (N2123, N2119);
and AND2 (N2124, N2123, N1608);
not NOT1 (N2125, N2107);
buf BUF1 (N2126, N2118);
and AND2 (N2127, N2115, N119);
buf BUF1 (N2128, N2096);
and AND2 (N2129, N2103, N1262);
and AND4 (N2130, N2125, N728, N1371, N2117);
buf BUF1 (N2131, N2122);
buf BUF1 (N2132, N2129);
not NOT1 (N2133, N2120);
xor XOR2 (N2134, N2132, N933);
or OR3 (N2135, N2134, N159, N1935);
or OR4 (N2136, N2124, N1312, N1213, N586);
xor XOR2 (N2137, N2077, N1925);
not NOT1 (N2138, N2133);
xor XOR2 (N2139, N2130, N1375);
xor XOR2 (N2140, N2126, N781);
buf BUF1 (N2141, N2139);
not NOT1 (N2142, N2140);
xor XOR2 (N2143, N2138, N540);
nand NAND4 (N2144, N2127, N310, N179, N1782);
nor NOR3 (N2145, N2142, N951, N1086);
xor XOR2 (N2146, N2128, N1575);
or OR2 (N2147, N2136, N340);
and AND2 (N2148, N2112, N172);
buf BUF1 (N2149, N2147);
buf BUF1 (N2150, N2141);
or OR2 (N2151, N2149, N1367);
not NOT1 (N2152, N2146);
and AND3 (N2153, N2148, N1297, N247);
or OR3 (N2154, N2135, N533, N1579);
buf BUF1 (N2155, N2137);
and AND4 (N2156, N2150, N2139, N296, N1293);
buf BUF1 (N2157, N2145);
buf BUF1 (N2158, N2143);
or OR2 (N2159, N2156, N1787);
or OR4 (N2160, N2154, N1465, N21, N1772);
xor XOR2 (N2161, N2144, N87);
nor NOR4 (N2162, N2161, N1325, N667, N784);
buf BUF1 (N2163, N2131);
nand NAND4 (N2164, N2158, N776, N246, N2031);
or OR3 (N2165, N2164, N415, N1327);
nor NOR4 (N2166, N2163, N472, N1406, N716);
and AND2 (N2167, N2165, N1337);
xor XOR2 (N2168, N2155, N1714);
xor XOR2 (N2169, N2152, N591);
and AND2 (N2170, N2153, N903);
and AND4 (N2171, N2170, N1866, N144, N311);
not NOT1 (N2172, N2157);
buf BUF1 (N2173, N2151);
nor NOR4 (N2174, N2162, N98, N964, N1265);
xor XOR2 (N2175, N2159, N874);
xor XOR2 (N2176, N2166, N456);
nor NOR4 (N2177, N2160, N1351, N1689, N236);
nand NAND4 (N2178, N2167, N1109, N1375, N916);
and AND4 (N2179, N2174, N2173, N855, N132);
nor NOR2 (N2180, N1681, N1485);
not NOT1 (N2181, N2179);
and AND3 (N2182, N2178, N1621, N27);
not NOT1 (N2183, N2171);
nor NOR4 (N2184, N2169, N2183, N454, N784);
xor XOR2 (N2185, N362, N674);
or OR4 (N2186, N2177, N618, N92, N289);
buf BUF1 (N2187, N2182);
buf BUF1 (N2188, N2168);
and AND2 (N2189, N2180, N7);
nor NOR2 (N2190, N2172, N271);
nor NOR4 (N2191, N2188, N200, N1094, N539);
nand NAND2 (N2192, N2189, N1418);
nor NOR2 (N2193, N2181, N461);
and AND4 (N2194, N2192, N749, N1558, N244);
xor XOR2 (N2195, N2190, N597);
xor XOR2 (N2196, N2187, N1530);
nand NAND4 (N2197, N2195, N1642, N1155, N459);
buf BUF1 (N2198, N2176);
nand NAND2 (N2199, N2175, N1078);
xor XOR2 (N2200, N2193, N970);
xor XOR2 (N2201, N2191, N136);
and AND2 (N2202, N2184, N1024);
nor NOR2 (N2203, N2197, N734);
nand NAND3 (N2204, N2201, N715, N2058);
or OR4 (N2205, N2203, N1924, N441, N348);
nand NAND2 (N2206, N2194, N1181);
not NOT1 (N2207, N2185);
or OR4 (N2208, N2196, N1612, N511, N689);
xor XOR2 (N2209, N2199, N413);
nand NAND3 (N2210, N2198, N408, N1729);
and AND3 (N2211, N2186, N990, N1662);
nand NAND2 (N2212, N2210, N1150);
buf BUF1 (N2213, N2200);
or OR2 (N2214, N2204, N723);
nand NAND3 (N2215, N2213, N1947, N837);
xor XOR2 (N2216, N2207, N141);
or OR4 (N2217, N2208, N1703, N620, N1028);
and AND4 (N2218, N2205, N998, N1920, N205);
not NOT1 (N2219, N2211);
nand NAND4 (N2220, N2215, N1335, N233, N221);
buf BUF1 (N2221, N2214);
xor XOR2 (N2222, N2209, N446);
nand NAND2 (N2223, N2222, N1408);
or OR4 (N2224, N2206, N1163, N1870, N160);
or OR3 (N2225, N2220, N1023, N2079);
nor NOR2 (N2226, N2217, N229);
and AND3 (N2227, N2216, N1053, N593);
xor XOR2 (N2228, N2212, N460);
buf BUF1 (N2229, N2219);
buf BUF1 (N2230, N2223);
and AND4 (N2231, N2218, N266, N1479, N1787);
or OR2 (N2232, N2224, N613);
and AND2 (N2233, N2230, N1904);
buf BUF1 (N2234, N2226);
nor NOR2 (N2235, N2229, N66);
not NOT1 (N2236, N2228);
nor NOR4 (N2237, N2221, N153, N1461, N1754);
buf BUF1 (N2238, N2237);
nand NAND3 (N2239, N2225, N1031, N1260);
buf BUF1 (N2240, N2231);
and AND3 (N2241, N2240, N824, N1903);
or OR2 (N2242, N2232, N974);
xor XOR2 (N2243, N2233, N1773);
nand NAND2 (N2244, N2234, N1999);
xor XOR2 (N2245, N2243, N1779);
or OR3 (N2246, N2227, N1195, N190);
nand NAND4 (N2247, N2235, N350, N173, N2127);
xor XOR2 (N2248, N2244, N1746);
not NOT1 (N2249, N2239);
buf BUF1 (N2250, N2249);
not NOT1 (N2251, N2202);
buf BUF1 (N2252, N2248);
and AND3 (N2253, N2252, N955, N1942);
xor XOR2 (N2254, N2238, N279);
or OR4 (N2255, N2245, N167, N89, N818);
and AND2 (N2256, N2246, N856);
or OR2 (N2257, N2254, N1281);
buf BUF1 (N2258, N2241);
and AND2 (N2259, N2256, N763);
xor XOR2 (N2260, N2247, N1634);
nand NAND4 (N2261, N2236, N954, N66, N2249);
and AND3 (N2262, N2259, N2185, N1194);
buf BUF1 (N2263, N2255);
buf BUF1 (N2264, N2258);
nand NAND2 (N2265, N2251, N1860);
or OR4 (N2266, N2265, N549, N877, N505);
or OR2 (N2267, N2263, N1759);
nand NAND3 (N2268, N2257, N157, N841);
not NOT1 (N2269, N2268);
and AND3 (N2270, N2242, N130, N560);
xor XOR2 (N2271, N2264, N1434);
or OR4 (N2272, N2267, N1334, N1088, N1064);
not NOT1 (N2273, N2272);
nor NOR3 (N2274, N2266, N777, N1943);
buf BUF1 (N2275, N2274);
nand NAND2 (N2276, N2270, N2067);
nor NOR2 (N2277, N2262, N705);
xor XOR2 (N2278, N2271, N1697);
and AND3 (N2279, N2250, N715, N335);
or OR4 (N2280, N2279, N2192, N1346, N1517);
and AND3 (N2281, N2269, N279, N2072);
nand NAND2 (N2282, N2281, N281);
or OR3 (N2283, N2260, N746, N2055);
buf BUF1 (N2284, N2282);
xor XOR2 (N2285, N2275, N934);
nor NOR4 (N2286, N2276, N1803, N1052, N1246);
buf BUF1 (N2287, N2283);
buf BUF1 (N2288, N2280);
xor XOR2 (N2289, N2253, N716);
nor NOR4 (N2290, N2284, N1992, N1973, N519);
and AND3 (N2291, N2288, N1244, N162);
and AND4 (N2292, N2261, N1716, N11, N938);
nor NOR2 (N2293, N2277, N347);
xor XOR2 (N2294, N2291, N290);
xor XOR2 (N2295, N2285, N486);
and AND3 (N2296, N2278, N974, N191);
nand NAND2 (N2297, N2287, N925);
and AND3 (N2298, N2289, N2182, N1575);
buf BUF1 (N2299, N2293);
nand NAND2 (N2300, N2290, N1035);
nor NOR3 (N2301, N2273, N97, N519);
and AND4 (N2302, N2298, N2268, N730, N612);
buf BUF1 (N2303, N2296);
nor NOR3 (N2304, N2300, N686, N411);
and AND3 (N2305, N2302, N292, N2186);
nor NOR3 (N2306, N2292, N2255, N2082);
and AND3 (N2307, N2304, N428, N2001);
or OR2 (N2308, N2307, N1009);
nand NAND4 (N2309, N2295, N1731, N1862, N119);
buf BUF1 (N2310, N2286);
nand NAND2 (N2311, N2301, N995);
or OR3 (N2312, N2306, N226, N1805);
and AND4 (N2313, N2309, N1853, N889, N1514);
nand NAND2 (N2314, N2311, N1947);
nor NOR4 (N2315, N2313, N685, N2048, N1446);
and AND4 (N2316, N2299, N1663, N1591, N575);
buf BUF1 (N2317, N2294);
not NOT1 (N2318, N2303);
or OR3 (N2319, N2314, N617, N1382);
nand NAND3 (N2320, N2316, N1919, N463);
buf BUF1 (N2321, N2297);
not NOT1 (N2322, N2305);
nor NOR2 (N2323, N2315, N1903);
not NOT1 (N2324, N2320);
not NOT1 (N2325, N2322);
nor NOR2 (N2326, N2324, N1694);
nor NOR2 (N2327, N2317, N2022);
or OR2 (N2328, N2318, N2293);
not NOT1 (N2329, N2308);
nor NOR3 (N2330, N2328, N2045, N486);
xor XOR2 (N2331, N2310, N907);
not NOT1 (N2332, N2326);
nor NOR4 (N2333, N2312, N1995, N1735, N1916);
nor NOR4 (N2334, N2333, N1099, N1917, N184);
xor XOR2 (N2335, N2331, N265);
xor XOR2 (N2336, N2330, N783);
xor XOR2 (N2337, N2321, N2214);
and AND4 (N2338, N2335, N1837, N1071, N403);
nor NOR2 (N2339, N2337, N1723);
xor XOR2 (N2340, N2329, N1155);
xor XOR2 (N2341, N2340, N920);
nor NOR2 (N2342, N2341, N1118);
nor NOR3 (N2343, N2336, N1141, N1855);
and AND3 (N2344, N2325, N899, N1525);
xor XOR2 (N2345, N2319, N644);
buf BUF1 (N2346, N2338);
not NOT1 (N2347, N2334);
not NOT1 (N2348, N2344);
nand NAND2 (N2349, N2346, N610);
xor XOR2 (N2350, N2342, N475);
or OR2 (N2351, N2332, N1815);
and AND3 (N2352, N2349, N742, N460);
nor NOR4 (N2353, N2352, N1339, N1510, N853);
buf BUF1 (N2354, N2339);
nand NAND4 (N2355, N2348, N1262, N2021, N369);
nand NAND4 (N2356, N2351, N1927, N1537, N540);
xor XOR2 (N2357, N2343, N1650);
nor NOR4 (N2358, N2356, N701, N662, N2237);
or OR3 (N2359, N2347, N2342, N1428);
nor NOR3 (N2360, N2353, N817, N2300);
or OR4 (N2361, N2360, N141, N381, N449);
or OR2 (N2362, N2350, N1682);
nand NAND2 (N2363, N2355, N368);
nand NAND3 (N2364, N2358, N1833, N209);
buf BUF1 (N2365, N2327);
xor XOR2 (N2366, N2323, N1739);
or OR4 (N2367, N2366, N1624, N327, N1917);
not NOT1 (N2368, N2361);
or OR2 (N2369, N2345, N1007);
nand NAND2 (N2370, N2369, N2190);
nor NOR4 (N2371, N2359, N577, N600, N2281);
nand NAND2 (N2372, N2354, N2328);
nor NOR3 (N2373, N2365, N1676, N264);
nand NAND4 (N2374, N2364, N1976, N1850, N2120);
nand NAND2 (N2375, N2357, N415);
not NOT1 (N2376, N2375);
and AND3 (N2377, N2368, N1845, N636);
xor XOR2 (N2378, N2377, N348);
buf BUF1 (N2379, N2363);
and AND3 (N2380, N2379, N1389, N829);
buf BUF1 (N2381, N2380);
xor XOR2 (N2382, N2381, N414);
and AND2 (N2383, N2378, N166);
xor XOR2 (N2384, N2370, N457);
or OR2 (N2385, N2376, N229);
and AND2 (N2386, N2382, N2299);
buf BUF1 (N2387, N2362);
and AND4 (N2388, N2386, N1991, N36, N157);
or OR3 (N2389, N2374, N402, N1601);
not NOT1 (N2390, N2373);
nor NOR4 (N2391, N2384, N1343, N1849, N670);
buf BUF1 (N2392, N2391);
and AND3 (N2393, N2372, N1727, N63);
buf BUF1 (N2394, N2393);
xor XOR2 (N2395, N2389, N1509);
not NOT1 (N2396, N2383);
and AND3 (N2397, N2394, N201, N2340);
nor NOR2 (N2398, N2388, N1219);
buf BUF1 (N2399, N2387);
nand NAND3 (N2400, N2395, N1776, N1906);
not NOT1 (N2401, N2371);
or OR3 (N2402, N2398, N1186, N1259);
not NOT1 (N2403, N2400);
and AND3 (N2404, N2401, N2251, N2036);
buf BUF1 (N2405, N2397);
xor XOR2 (N2406, N2405, N2319);
and AND2 (N2407, N2406, N1552);
or OR2 (N2408, N2402, N575);
nand NAND3 (N2409, N2367, N756, N678);
xor XOR2 (N2410, N2407, N142);
nand NAND3 (N2411, N2409, N1672, N1920);
xor XOR2 (N2412, N2411, N958);
or OR4 (N2413, N2408, N870, N371, N1198);
not NOT1 (N2414, N2410);
xor XOR2 (N2415, N2399, N446);
nand NAND3 (N2416, N2413, N1471, N1803);
xor XOR2 (N2417, N2403, N2057);
nand NAND4 (N2418, N2396, N1731, N1179, N836);
not NOT1 (N2419, N2415);
buf BUF1 (N2420, N2416);
nand NAND2 (N2421, N2404, N2365);
nand NAND4 (N2422, N2390, N2209, N741, N2228);
or OR2 (N2423, N2412, N620);
xor XOR2 (N2424, N2392, N1785);
not NOT1 (N2425, N2422);
or OR4 (N2426, N2417, N2401, N864, N631);
buf BUF1 (N2427, N2424);
or OR2 (N2428, N2420, N1268);
not NOT1 (N2429, N2414);
not NOT1 (N2430, N2385);
nand NAND2 (N2431, N2418, N1882);
nor NOR3 (N2432, N2427, N2339, N843);
nor NOR3 (N2433, N2425, N2019, N699);
or OR2 (N2434, N2421, N1250);
nand NAND4 (N2435, N2431, N443, N2378, N71);
and AND4 (N2436, N2419, N279, N1188, N2243);
or OR2 (N2437, N2423, N198);
not NOT1 (N2438, N2432);
nand NAND2 (N2439, N2430, N1522);
or OR4 (N2440, N2435, N1310, N981, N374);
nor NOR4 (N2441, N2440, N51, N182, N106);
xor XOR2 (N2442, N2436, N980);
or OR4 (N2443, N2442, N227, N2, N2154);
and AND3 (N2444, N2438, N1011, N1536);
xor XOR2 (N2445, N2443, N837);
not NOT1 (N2446, N2426);
nand NAND3 (N2447, N2444, N2350, N415);
or OR4 (N2448, N2433, N1529, N1814, N1598);
and AND2 (N2449, N2437, N2299);
or OR4 (N2450, N2449, N1922, N1273, N1688);
or OR3 (N2451, N2448, N1785, N998);
not NOT1 (N2452, N2441);
xor XOR2 (N2453, N2451, N1838);
nor NOR3 (N2454, N2447, N453, N2043);
and AND2 (N2455, N2429, N2283);
and AND2 (N2456, N2450, N2358);
xor XOR2 (N2457, N2434, N707);
buf BUF1 (N2458, N2455);
buf BUF1 (N2459, N2456);
and AND3 (N2460, N2459, N504, N818);
not NOT1 (N2461, N2452);
buf BUF1 (N2462, N2460);
nor NOR4 (N2463, N2453, N159, N311, N2330);
and AND2 (N2464, N2439, N608);
nand NAND3 (N2465, N2457, N2035, N1828);
not NOT1 (N2466, N2458);
nor NOR4 (N2467, N2464, N1131, N1186, N1819);
or OR3 (N2468, N2445, N602, N1713);
nor NOR3 (N2469, N2466, N1948, N2360);
buf BUF1 (N2470, N2467);
nor NOR2 (N2471, N2462, N120);
xor XOR2 (N2472, N2465, N1079);
or OR4 (N2473, N2469, N685, N1255, N1943);
nor NOR2 (N2474, N2468, N2024);
and AND4 (N2475, N2454, N237, N559, N2366);
nand NAND4 (N2476, N2463, N1603, N1308, N467);
buf BUF1 (N2477, N2474);
nor NOR4 (N2478, N2428, N702, N2445, N419);
nand NAND2 (N2479, N2478, N1809);
or OR4 (N2480, N2471, N1473, N1727, N1386);
not NOT1 (N2481, N2446);
xor XOR2 (N2482, N2480, N2473);
and AND4 (N2483, N2372, N1798, N1671, N2015);
buf BUF1 (N2484, N2476);
nor NOR3 (N2485, N2483, N1229, N1393);
buf BUF1 (N2486, N2482);
and AND3 (N2487, N2481, N2438, N2294);
xor XOR2 (N2488, N2472, N1895);
xor XOR2 (N2489, N2485, N1479);
and AND4 (N2490, N2479, N1199, N272, N2226);
xor XOR2 (N2491, N2477, N1508);
xor XOR2 (N2492, N2490, N237);
or OR4 (N2493, N2470, N2371, N2147, N228);
nand NAND2 (N2494, N2493, N619);
not NOT1 (N2495, N2494);
nand NAND2 (N2496, N2495, N2478);
nor NOR3 (N2497, N2475, N1466, N2295);
nand NAND4 (N2498, N2491, N2126, N2120, N297);
not NOT1 (N2499, N2488);
nor NOR2 (N2500, N2489, N1676);
buf BUF1 (N2501, N2499);
not NOT1 (N2502, N2500);
buf BUF1 (N2503, N2486);
nor NOR4 (N2504, N2492, N1561, N1331, N54);
buf BUF1 (N2505, N2496);
xor XOR2 (N2506, N2497, N1277);
nand NAND3 (N2507, N2505, N1118, N2475);
not NOT1 (N2508, N2506);
nand NAND3 (N2509, N2504, N1597, N1580);
and AND4 (N2510, N2498, N1427, N2005, N772);
not NOT1 (N2511, N2509);
buf BUF1 (N2512, N2503);
nand NAND4 (N2513, N2512, N1310, N436, N1459);
and AND2 (N2514, N2502, N2371);
nand NAND4 (N2515, N2508, N792, N1786, N121);
and AND3 (N2516, N2487, N145, N958);
not NOT1 (N2517, N2513);
nor NOR4 (N2518, N2484, N232, N1663, N2273);
nor NOR2 (N2519, N2516, N1008);
xor XOR2 (N2520, N2518, N1460);
nand NAND2 (N2521, N2461, N821);
buf BUF1 (N2522, N2517);
and AND4 (N2523, N2511, N262, N597, N639);
nor NOR4 (N2524, N2523, N94, N1402, N554);
or OR2 (N2525, N2510, N392);
and AND3 (N2526, N2520, N784, N1573);
and AND2 (N2527, N2514, N424);
nor NOR4 (N2528, N2525, N938, N1499, N2360);
not NOT1 (N2529, N2528);
buf BUF1 (N2530, N2527);
nand NAND2 (N2531, N2529, N1989);
buf BUF1 (N2532, N2507);
and AND2 (N2533, N2524, N2374);
buf BUF1 (N2534, N2519);
xor XOR2 (N2535, N2530, N1339);
or OR3 (N2536, N2526, N2532, N2469);
and AND4 (N2537, N1988, N1148, N344, N380);
buf BUF1 (N2538, N2536);
xor XOR2 (N2539, N2533, N2487);
xor XOR2 (N2540, N2537, N25);
buf BUF1 (N2541, N2535);
not NOT1 (N2542, N2531);
buf BUF1 (N2543, N2521);
buf BUF1 (N2544, N2543);
xor XOR2 (N2545, N2540, N2394);
not NOT1 (N2546, N2545);
and AND2 (N2547, N2539, N591);
or OR4 (N2548, N2544, N1534, N1993, N1883);
or OR3 (N2549, N2522, N1322, N786);
nand NAND2 (N2550, N2542, N2419);
and AND4 (N2551, N2538, N1279, N2294, N1723);
xor XOR2 (N2552, N2548, N1180);
buf BUF1 (N2553, N2547);
or OR4 (N2554, N2515, N467, N2464, N2444);
not NOT1 (N2555, N2541);
and AND4 (N2556, N2534, N1723, N578, N1420);
xor XOR2 (N2557, N2553, N946);
or OR4 (N2558, N2550, N1640, N2325, N1033);
or OR4 (N2559, N2558, N2490, N816, N243);
nand NAND4 (N2560, N2554, N1923, N2065, N85);
or OR3 (N2561, N2549, N1708, N550);
nand NAND4 (N2562, N2546, N1741, N2130, N2013);
not NOT1 (N2563, N2562);
and AND2 (N2564, N2560, N781);
buf BUF1 (N2565, N2563);
not NOT1 (N2566, N2564);
buf BUF1 (N2567, N2552);
buf BUF1 (N2568, N2559);
and AND4 (N2569, N2568, N2340, N1785, N2402);
and AND3 (N2570, N2501, N940, N1307);
not NOT1 (N2571, N2555);
buf BUF1 (N2572, N2556);
xor XOR2 (N2573, N2551, N1957);
or OR3 (N2574, N2561, N2345, N1187);
nand NAND2 (N2575, N2557, N191);
xor XOR2 (N2576, N2567, N2571);
buf BUF1 (N2577, N1929);
nor NOR4 (N2578, N2572, N446, N1072, N2128);
xor XOR2 (N2579, N2578, N1910);
nand NAND2 (N2580, N2573, N2115);
buf BUF1 (N2581, N2577);
or OR2 (N2582, N2570, N1391);
and AND2 (N2583, N2582, N2144);
and AND3 (N2584, N2574, N1958, N1151);
not NOT1 (N2585, N2579);
nor NOR2 (N2586, N2583, N1463);
and AND4 (N2587, N2584, N2095, N212, N1397);
buf BUF1 (N2588, N2575);
buf BUF1 (N2589, N2576);
xor XOR2 (N2590, N2589, N1567);
nor NOR3 (N2591, N2587, N2274, N192);
and AND2 (N2592, N2569, N1029);
not NOT1 (N2593, N2586);
and AND2 (N2594, N2580, N2288);
nor NOR2 (N2595, N2585, N1519);
nor NOR3 (N2596, N2566, N1030, N801);
nor NOR3 (N2597, N2592, N1342, N1019);
or OR2 (N2598, N2596, N2303);
not NOT1 (N2599, N2593);
and AND4 (N2600, N2599, N1668, N1444, N1950);
xor XOR2 (N2601, N2598, N1569);
not NOT1 (N2602, N2588);
buf BUF1 (N2603, N2601);
nand NAND3 (N2604, N2565, N2071, N37);
not NOT1 (N2605, N2603);
not NOT1 (N2606, N2604);
buf BUF1 (N2607, N2594);
or OR2 (N2608, N2606, N1038);
buf BUF1 (N2609, N2595);
not NOT1 (N2610, N2590);
xor XOR2 (N2611, N2610, N329);
not NOT1 (N2612, N2597);
or OR4 (N2613, N2600, N1900, N2415, N2234);
xor XOR2 (N2614, N2608, N33);
xor XOR2 (N2615, N2581, N471);
nor NOR4 (N2616, N2607, N873, N839, N1075);
or OR4 (N2617, N2614, N1641, N729, N311);
and AND3 (N2618, N2602, N99, N347);
not NOT1 (N2619, N2618);
not NOT1 (N2620, N2617);
nand NAND4 (N2621, N2613, N2200, N2605, N2022);
or OR4 (N2622, N2057, N853, N1172, N2557);
xor XOR2 (N2623, N2616, N1270);
not NOT1 (N2624, N2620);
and AND4 (N2625, N2611, N1894, N2440, N269);
nand NAND4 (N2626, N2621, N133, N2198, N305);
not NOT1 (N2627, N2623);
nor NOR3 (N2628, N2626, N696, N1951);
not NOT1 (N2629, N2615);
not NOT1 (N2630, N2628);
buf BUF1 (N2631, N2624);
or OR4 (N2632, N2631, N1408, N1341, N1052);
and AND2 (N2633, N2625, N1626);
nand NAND4 (N2634, N2629, N1541, N2421, N1107);
or OR3 (N2635, N2619, N1523, N1849);
not NOT1 (N2636, N2630);
xor XOR2 (N2637, N2612, N2503);
and AND2 (N2638, N2633, N1493);
xor XOR2 (N2639, N2638, N985);
nor NOR4 (N2640, N2591, N841, N2326, N481);
not NOT1 (N2641, N2622);
and AND3 (N2642, N2609, N2119, N1307);
not NOT1 (N2643, N2642);
or OR4 (N2644, N2636, N1388, N33, N2023);
or OR2 (N2645, N2637, N1619);
buf BUF1 (N2646, N2634);
and AND3 (N2647, N2632, N966, N152);
nand NAND3 (N2648, N2641, N20, N181);
nand NAND4 (N2649, N2646, N759, N1526, N766);
buf BUF1 (N2650, N2635);
and AND4 (N2651, N2640, N898, N2286, N1994);
buf BUF1 (N2652, N2649);
buf BUF1 (N2653, N2648);
and AND3 (N2654, N2645, N74, N1415);
not NOT1 (N2655, N2654);
nand NAND2 (N2656, N2652, N933);
buf BUF1 (N2657, N2651);
and AND4 (N2658, N2657, N263, N1599, N1645);
buf BUF1 (N2659, N2650);
or OR4 (N2660, N2643, N142, N161, N961);
nand NAND2 (N2661, N2639, N125);
not NOT1 (N2662, N2644);
nand NAND4 (N2663, N2662, N2226, N1101, N504);
not NOT1 (N2664, N2653);
nor NOR4 (N2665, N2663, N1803, N501, N1034);
or OR4 (N2666, N2665, N256, N780, N1376);
xor XOR2 (N2667, N2661, N1324);
nand NAND2 (N2668, N2647, N668);
or OR2 (N2669, N2667, N365);
or OR3 (N2670, N2664, N244, N1300);
nor NOR2 (N2671, N2668, N607);
nand NAND2 (N2672, N2670, N2059);
xor XOR2 (N2673, N2669, N1015);
or OR2 (N2674, N2658, N1972);
not NOT1 (N2675, N2673);
and AND3 (N2676, N2659, N1764, N1528);
nor NOR3 (N2677, N2671, N2408, N477);
or OR4 (N2678, N2660, N1019, N1466, N2564);
not NOT1 (N2679, N2677);
nand NAND3 (N2680, N2679, N734, N1912);
not NOT1 (N2681, N2674);
and AND4 (N2682, N2680, N2538, N204, N2078);
buf BUF1 (N2683, N2656);
nand NAND4 (N2684, N2682, N1855, N2185, N1218);
nor NOR3 (N2685, N2672, N2030, N2582);
or OR2 (N2686, N2676, N1483);
and AND3 (N2687, N2681, N2456, N691);
not NOT1 (N2688, N2678);
xor XOR2 (N2689, N2627, N831);
nor NOR2 (N2690, N2683, N922);
or OR4 (N2691, N2675, N1322, N1121, N607);
xor XOR2 (N2692, N2691, N187);
and AND2 (N2693, N2688, N2623);
nor NOR2 (N2694, N2690, N338);
nor NOR3 (N2695, N2685, N2188, N2531);
xor XOR2 (N2696, N2655, N2112);
nand NAND2 (N2697, N2692, N2554);
nand NAND3 (N2698, N2684, N1153, N223);
not NOT1 (N2699, N2686);
and AND4 (N2700, N2687, N1656, N1595, N1535);
and AND4 (N2701, N2666, N933, N2167, N59);
xor XOR2 (N2702, N2698, N1000);
xor XOR2 (N2703, N2700, N953);
buf BUF1 (N2704, N2701);
nand NAND4 (N2705, N2702, N424, N1281, N2568);
buf BUF1 (N2706, N2705);
not NOT1 (N2707, N2694);
buf BUF1 (N2708, N2693);
and AND2 (N2709, N2707, N1566);
not NOT1 (N2710, N2695);
nor NOR3 (N2711, N2709, N1253, N2509);
xor XOR2 (N2712, N2699, N16);
or OR2 (N2713, N2689, N2259);
or OR2 (N2714, N2711, N664);
and AND2 (N2715, N2703, N2064);
or OR2 (N2716, N2704, N2693);
buf BUF1 (N2717, N2712);
nor NOR3 (N2718, N2710, N139, N1322);
buf BUF1 (N2719, N2706);
or OR2 (N2720, N2697, N2668);
nand NAND3 (N2721, N2717, N1767, N2108);
buf BUF1 (N2722, N2713);
not NOT1 (N2723, N2720);
nand NAND4 (N2724, N2719, N2338, N2404, N2606);
nand NAND3 (N2725, N2716, N2347, N2714);
nand NAND4 (N2726, N2486, N2614, N2369, N1746);
and AND3 (N2727, N2722, N175, N1771);
not NOT1 (N2728, N2708);
not NOT1 (N2729, N2718);
buf BUF1 (N2730, N2727);
or OR3 (N2731, N2726, N2060, N1397);
nor NOR3 (N2732, N2723, N2541, N1380);
nand NAND2 (N2733, N2715, N1012);
nor NOR4 (N2734, N2732, N315, N2144, N1523);
not NOT1 (N2735, N2696);
nor NOR4 (N2736, N2730, N2649, N2215, N342);
and AND3 (N2737, N2721, N1816, N45);
nand NAND3 (N2738, N2735, N2422, N363);
nand NAND4 (N2739, N2724, N2522, N8, N1062);
not NOT1 (N2740, N2738);
nor NOR2 (N2741, N2737, N1842);
or OR3 (N2742, N2739, N2222, N1654);
and AND2 (N2743, N2734, N841);
buf BUF1 (N2744, N2729);
buf BUF1 (N2745, N2733);
nor NOR3 (N2746, N2736, N1375, N2135);
nand NAND2 (N2747, N2742, N53);
or OR4 (N2748, N2744, N2044, N413, N808);
not NOT1 (N2749, N2731);
nand NAND4 (N2750, N2728, N1260, N703, N2001);
xor XOR2 (N2751, N2747, N384);
not NOT1 (N2752, N2745);
xor XOR2 (N2753, N2749, N1077);
not NOT1 (N2754, N2753);
nor NOR2 (N2755, N2741, N1533);
not NOT1 (N2756, N2752);
or OR4 (N2757, N2754, N1304, N334, N1138);
nor NOR4 (N2758, N2757, N2618, N562, N2348);
not NOT1 (N2759, N2758);
nor NOR2 (N2760, N2751, N2552);
nor NOR2 (N2761, N2750, N2557);
not NOT1 (N2762, N2756);
buf BUF1 (N2763, N2740);
or OR2 (N2764, N2760, N1049);
and AND3 (N2765, N2763, N2337, N1938);
and AND4 (N2766, N2746, N1966, N1356, N495);
buf BUF1 (N2767, N2725);
or OR3 (N2768, N2762, N231, N235);
or OR3 (N2769, N2764, N1253, N1239);
or OR4 (N2770, N2755, N929, N2115, N354);
or OR2 (N2771, N2766, N1);
nand NAND2 (N2772, N2768, N1133);
or OR4 (N2773, N2748, N2507, N2082, N152);
or OR3 (N2774, N2765, N2026, N652);
not NOT1 (N2775, N2774);
nor NOR3 (N2776, N2767, N2190, N1196);
and AND3 (N2777, N2743, N50, N1787);
nand NAND4 (N2778, N2761, N1589, N1941, N1656);
nand NAND3 (N2779, N2773, N2065, N2693);
nor NOR4 (N2780, N2772, N1331, N938, N29);
nand NAND3 (N2781, N2771, N973, N881);
xor XOR2 (N2782, N2781, N626);
and AND4 (N2783, N2775, N1642, N703, N1676);
nor NOR2 (N2784, N2769, N2325);
buf BUF1 (N2785, N2770);
or OR3 (N2786, N2785, N769, N1275);
buf BUF1 (N2787, N2759);
and AND2 (N2788, N2786, N881);
nand NAND4 (N2789, N2777, N1470, N2047, N567);
nand NAND4 (N2790, N2782, N2639, N2597, N2338);
nor NOR3 (N2791, N2790, N2640, N1461);
not NOT1 (N2792, N2788);
and AND2 (N2793, N2779, N2052);
xor XOR2 (N2794, N2778, N1479);
and AND4 (N2795, N2791, N322, N168, N2637);
not NOT1 (N2796, N2793);
not NOT1 (N2797, N2789);
not NOT1 (N2798, N2797);
buf BUF1 (N2799, N2776);
nand NAND2 (N2800, N2792, N1411);
not NOT1 (N2801, N2794);
not NOT1 (N2802, N2795);
nand NAND3 (N2803, N2802, N1167, N217);
not NOT1 (N2804, N2800);
not NOT1 (N2805, N2799);
buf BUF1 (N2806, N2804);
xor XOR2 (N2807, N2798, N2764);
and AND2 (N2808, N2806, N918);
nor NOR3 (N2809, N2780, N1194, N1096);
and AND3 (N2810, N2784, N958, N1430);
xor XOR2 (N2811, N2801, N614);
nor NOR3 (N2812, N2811, N916, N472);
not NOT1 (N2813, N2810);
xor XOR2 (N2814, N2805, N413);
and AND3 (N2815, N2814, N2428, N2097);
not NOT1 (N2816, N2796);
not NOT1 (N2817, N2808);
nor NOR2 (N2818, N2809, N1609);
nor NOR4 (N2819, N2818, N593, N98, N317);
and AND3 (N2820, N2787, N1591, N829);
not NOT1 (N2821, N2817);
nor NOR4 (N2822, N2820, N848, N626, N1147);
xor XOR2 (N2823, N2816, N2510);
xor XOR2 (N2824, N2783, N816);
or OR3 (N2825, N2819, N1000, N2365);
xor XOR2 (N2826, N2824, N2286);
not NOT1 (N2827, N2822);
not NOT1 (N2828, N2815);
buf BUF1 (N2829, N2812);
nand NAND2 (N2830, N2823, N1112);
not NOT1 (N2831, N2830);
and AND3 (N2832, N2831, N2560, N1417);
or OR2 (N2833, N2832, N1590);
nor NOR4 (N2834, N2807, N197, N811, N1014);
buf BUF1 (N2835, N2833);
not NOT1 (N2836, N2821);
buf BUF1 (N2837, N2826);
not NOT1 (N2838, N2835);
buf BUF1 (N2839, N2834);
nor NOR3 (N2840, N2828, N356, N2120);
and AND2 (N2841, N2840, N225);
xor XOR2 (N2842, N2838, N2236);
buf BUF1 (N2843, N2837);
not NOT1 (N2844, N2843);
and AND2 (N2845, N2836, N1060);
nor NOR4 (N2846, N2803, N974, N1826, N2811);
not NOT1 (N2847, N2827);
or OR3 (N2848, N2844, N190, N758);
or OR3 (N2849, N2839, N1979, N7);
buf BUF1 (N2850, N2845);
and AND2 (N2851, N2842, N2143);
xor XOR2 (N2852, N2846, N1236);
and AND4 (N2853, N2848, N386, N2461, N1663);
xor XOR2 (N2854, N2850, N2593);
buf BUF1 (N2855, N2825);
nor NOR3 (N2856, N2855, N119, N2399);
nor NOR3 (N2857, N2856, N57, N2555);
xor XOR2 (N2858, N2852, N592);
xor XOR2 (N2859, N2841, N1564);
nor NOR4 (N2860, N2853, N1294, N2034, N476);
xor XOR2 (N2861, N2849, N2116);
and AND2 (N2862, N2851, N1391);
and AND4 (N2863, N2858, N1759, N479, N1830);
buf BUF1 (N2864, N2859);
not NOT1 (N2865, N2857);
or OR4 (N2866, N2863, N1143, N1299, N1456);
buf BUF1 (N2867, N2865);
nand NAND3 (N2868, N2862, N66, N2385);
not NOT1 (N2869, N2847);
nand NAND4 (N2870, N2869, N520, N2057, N1636);
xor XOR2 (N2871, N2813, N1464);
not NOT1 (N2872, N2854);
xor XOR2 (N2873, N2868, N439);
nor NOR2 (N2874, N2866, N765);
nand NAND2 (N2875, N2873, N1549);
buf BUF1 (N2876, N2860);
and AND2 (N2877, N2829, N1459);
not NOT1 (N2878, N2875);
xor XOR2 (N2879, N2878, N1764);
or OR4 (N2880, N2879, N1851, N440, N276);
and AND3 (N2881, N2877, N2832, N1961);
buf BUF1 (N2882, N2876);
xor XOR2 (N2883, N2881, N891);
or OR3 (N2884, N2883, N1150, N1253);
or OR3 (N2885, N2872, N598, N2663);
nand NAND4 (N2886, N2867, N329, N1771, N1823);
buf BUF1 (N2887, N2870);
or OR3 (N2888, N2885, N1949, N2320);
nand NAND4 (N2889, N2880, N2735, N356, N813);
buf BUF1 (N2890, N2861);
or OR2 (N2891, N2889, N2884);
nand NAND2 (N2892, N1384, N2405);
and AND3 (N2893, N2887, N1977, N1319);
nand NAND2 (N2894, N2886, N384);
nand NAND2 (N2895, N2864, N2133);
or OR4 (N2896, N2890, N1432, N989, N2384);
or OR3 (N2897, N2888, N2536, N120);
nor NOR2 (N2898, N2897, N2509);
nor NOR4 (N2899, N2898, N1421, N1674, N1333);
nor NOR4 (N2900, N2895, N2865, N1629, N1929);
and AND4 (N2901, N2899, N1044, N2070, N1767);
xor XOR2 (N2902, N2892, N1307);
nand NAND4 (N2903, N2871, N2403, N1042, N1563);
buf BUF1 (N2904, N2900);
nand NAND2 (N2905, N2894, N2651);
nand NAND2 (N2906, N2901, N731);
xor XOR2 (N2907, N2893, N453);
xor XOR2 (N2908, N2907, N696);
or OR4 (N2909, N2882, N1978, N237, N800);
or OR3 (N2910, N2874, N1954, N51);
nand NAND3 (N2911, N2906, N1892, N2617);
buf BUF1 (N2912, N2909);
or OR4 (N2913, N2912, N2313, N969, N140);
nand NAND3 (N2914, N2913, N183, N2263);
xor XOR2 (N2915, N2910, N180);
nor NOR2 (N2916, N2902, N2829);
nor NOR2 (N2917, N2903, N494);
and AND4 (N2918, N2915, N2713, N1631, N810);
nor NOR4 (N2919, N2918, N1574, N2738, N1626);
nand NAND4 (N2920, N2919, N1665, N323, N1949);
nor NOR4 (N2921, N2904, N1564, N857, N2742);
or OR3 (N2922, N2896, N1729, N1822);
nor NOR4 (N2923, N2911, N1584, N1780, N2774);
xor XOR2 (N2924, N2908, N372);
nor NOR4 (N2925, N2921, N1625, N2390, N2514);
and AND4 (N2926, N2905, N1279, N1714, N2854);
and AND3 (N2927, N2926, N806, N2490);
buf BUF1 (N2928, N2925);
or OR2 (N2929, N2922, N2830);
buf BUF1 (N2930, N2924);
and AND2 (N2931, N2914, N1380);
buf BUF1 (N2932, N2917);
buf BUF1 (N2933, N2891);
nor NOR2 (N2934, N2929, N699);
xor XOR2 (N2935, N2930, N2442);
nor NOR4 (N2936, N2928, N902, N2319, N1831);
buf BUF1 (N2937, N2923);
nor NOR4 (N2938, N2935, N1943, N530, N1901);
nor NOR2 (N2939, N2934, N1358);
xor XOR2 (N2940, N2920, N2029);
nand NAND2 (N2941, N2931, N2235);
and AND3 (N2942, N2936, N549, N2536);
xor XOR2 (N2943, N2927, N1639);
not NOT1 (N2944, N2940);
or OR3 (N2945, N2944, N2854, N59);
nor NOR3 (N2946, N2939, N1426, N2024);
nand NAND4 (N2947, N2916, N2329, N1945, N721);
and AND2 (N2948, N2945, N2730);
or OR3 (N2949, N2938, N198, N2321);
not NOT1 (N2950, N2932);
not NOT1 (N2951, N2948);
nand NAND2 (N2952, N2942, N1586);
xor XOR2 (N2953, N2950, N2589);
nand NAND3 (N2954, N2946, N2025, N1011);
buf BUF1 (N2955, N2954);
nor NOR2 (N2956, N2937, N1180);
nand NAND4 (N2957, N2952, N4, N937, N2789);
nand NAND4 (N2958, N2953, N2184, N1239, N2535);
or OR4 (N2959, N2956, N1921, N1846, N620);
not NOT1 (N2960, N2959);
and AND2 (N2961, N2955, N2703);
not NOT1 (N2962, N2949);
and AND3 (N2963, N2947, N1750, N760);
buf BUF1 (N2964, N2961);
and AND3 (N2965, N2957, N1375, N337);
nor NOR4 (N2966, N2964, N661, N989, N2056);
and AND3 (N2967, N2965, N51, N2900);
not NOT1 (N2968, N2967);
or OR3 (N2969, N2962, N2022, N582);
buf BUF1 (N2970, N2943);
xor XOR2 (N2971, N2958, N12);
xor XOR2 (N2972, N2933, N820);
nand NAND2 (N2973, N2972, N1585);
buf BUF1 (N2974, N2963);
nor NOR2 (N2975, N2966, N2311);
buf BUF1 (N2976, N2973);
xor XOR2 (N2977, N2951, N855);
nand NAND2 (N2978, N2971, N2746);
xor XOR2 (N2979, N2941, N2689);
and AND2 (N2980, N2974, N333);
nand NAND3 (N2981, N2975, N1432, N53);
or OR4 (N2982, N2978, N1350, N2644, N1318);
nor NOR2 (N2983, N2970, N2556);
not NOT1 (N2984, N2977);
not NOT1 (N2985, N2979);
not NOT1 (N2986, N2969);
and AND4 (N2987, N2980, N1, N2013, N2378);
and AND2 (N2988, N2982, N1005);
nand NAND3 (N2989, N2983, N1629, N644);
xor XOR2 (N2990, N2986, N6);
not NOT1 (N2991, N2988);
or OR3 (N2992, N2985, N999, N1445);
nand NAND3 (N2993, N2991, N953, N4);
nand NAND4 (N2994, N2993, N378, N2492, N1022);
or OR2 (N2995, N2968, N821);
or OR4 (N2996, N2994, N2247, N2272, N1408);
not NOT1 (N2997, N2992);
buf BUF1 (N2998, N2976);
nand NAND3 (N2999, N2989, N2138, N2901);
buf BUF1 (N3000, N2981);
buf BUF1 (N3001, N2987);
not NOT1 (N3002, N3001);
nand NAND3 (N3003, N3002, N2827, N2107);
or OR3 (N3004, N2960, N1585, N49);
xor XOR2 (N3005, N2998, N2037);
nor NOR2 (N3006, N3004, N1999);
buf BUF1 (N3007, N2997);
nor NOR4 (N3008, N3003, N2423, N2954, N1198);
not NOT1 (N3009, N3000);
or OR2 (N3010, N3008, N221);
nand NAND2 (N3011, N3009, N1739);
and AND2 (N3012, N2999, N579);
not NOT1 (N3013, N3005);
buf BUF1 (N3014, N3010);
and AND4 (N3015, N3014, N2817, N2055, N763);
or OR4 (N3016, N3013, N647, N1107, N2192);
nor NOR2 (N3017, N3012, N1704);
or OR4 (N3018, N3016, N436, N2237, N1713);
xor XOR2 (N3019, N3015, N846);
and AND3 (N3020, N2990, N2854, N2599);
xor XOR2 (N3021, N3019, N2957);
or OR2 (N3022, N2995, N1323);
buf BUF1 (N3023, N3018);
buf BUF1 (N3024, N3021);
not NOT1 (N3025, N3006);
and AND2 (N3026, N3025, N2499);
nor NOR2 (N3027, N3007, N1162);
buf BUF1 (N3028, N3027);
or OR2 (N3029, N3011, N1778);
buf BUF1 (N3030, N2996);
buf BUF1 (N3031, N3024);
not NOT1 (N3032, N3022);
buf BUF1 (N3033, N3017);
xor XOR2 (N3034, N3023, N454);
and AND2 (N3035, N3028, N1911);
buf BUF1 (N3036, N3034);
buf BUF1 (N3037, N3031);
xor XOR2 (N3038, N3029, N1712);
and AND4 (N3039, N3026, N1631, N1824, N1085);
or OR4 (N3040, N3020, N1447, N1183, N871);
xor XOR2 (N3041, N3039, N1273);
or OR2 (N3042, N3036, N1602);
and AND4 (N3043, N3042, N2453, N630, N1728);
nand NAND3 (N3044, N3035, N2177, N737);
buf BUF1 (N3045, N3032);
not NOT1 (N3046, N3033);
nor NOR4 (N3047, N3044, N1055, N281, N1363);
and AND3 (N3048, N3040, N2706, N1991);
nor NOR4 (N3049, N3030, N2121, N1820, N970);
xor XOR2 (N3050, N3043, N2837);
nand NAND4 (N3051, N3041, N1558, N2440, N393);
buf BUF1 (N3052, N3049);
nand NAND4 (N3053, N3048, N1300, N1760, N2876);
nor NOR3 (N3054, N2984, N947, N2407);
or OR3 (N3055, N3050, N746, N1286);
and AND2 (N3056, N3047, N1924);
buf BUF1 (N3057, N3053);
or OR2 (N3058, N3051, N2039);
and AND2 (N3059, N3057, N479);
not NOT1 (N3060, N3054);
and AND3 (N3061, N3046, N1896, N963);
nor NOR4 (N3062, N3060, N1791, N157, N497);
not NOT1 (N3063, N3058);
and AND2 (N3064, N3062, N749);
and AND2 (N3065, N3038, N1008);
not NOT1 (N3066, N3056);
nand NAND2 (N3067, N3065, N1050);
buf BUF1 (N3068, N3064);
xor XOR2 (N3069, N3052, N2682);
and AND4 (N3070, N3066, N990, N2735, N2438);
nand NAND2 (N3071, N3059, N48);
or OR3 (N3072, N3055, N1884, N602);
not NOT1 (N3073, N3067);
or OR3 (N3074, N3037, N2522, N632);
or OR2 (N3075, N3045, N94);
and AND2 (N3076, N3075, N1925);
nand NAND2 (N3077, N3069, N1371);
or OR3 (N3078, N3061, N1040, N852);
nor NOR4 (N3079, N3063, N434, N2265, N629);
or OR4 (N3080, N3074, N50, N1502, N2817);
and AND4 (N3081, N3078, N1221, N2507, N1062);
or OR4 (N3082, N3068, N466, N306, N2159);
xor XOR2 (N3083, N3072, N2688);
buf BUF1 (N3084, N3076);
not NOT1 (N3085, N3080);
nor NOR4 (N3086, N3083, N2402, N1326, N688);
xor XOR2 (N3087, N3084, N2166);
buf BUF1 (N3088, N3070);
xor XOR2 (N3089, N3073, N1281);
or OR2 (N3090, N3081, N2727);
not NOT1 (N3091, N3071);
and AND2 (N3092, N3090, N555);
nor NOR2 (N3093, N3086, N687);
xor XOR2 (N3094, N3091, N1599);
nand NAND3 (N3095, N3082, N2848, N1939);
nor NOR4 (N3096, N3095, N2308, N1894, N759);
and AND3 (N3097, N3089, N1686, N1496);
or OR3 (N3098, N3093, N1301, N2731);
xor XOR2 (N3099, N3097, N893);
and AND2 (N3100, N3079, N2790);
xor XOR2 (N3101, N3100, N349);
buf BUF1 (N3102, N3101);
and AND4 (N3103, N3094, N1173, N1167, N2821);
buf BUF1 (N3104, N3087);
and AND3 (N3105, N3103, N2675, N883);
buf BUF1 (N3106, N3099);
nand NAND4 (N3107, N3098, N1529, N2406, N75);
and AND3 (N3108, N3106, N1071, N193);
buf BUF1 (N3109, N3085);
nor NOR2 (N3110, N3088, N2762);
nor NOR2 (N3111, N3105, N1759);
and AND4 (N3112, N3102, N1637, N2334, N2894);
nor NOR2 (N3113, N3109, N2881);
not NOT1 (N3114, N3111);
nor NOR4 (N3115, N3077, N1363, N1338, N159);
buf BUF1 (N3116, N3108);
nand NAND3 (N3117, N3107, N2130, N960);
or OR4 (N3118, N3113, N536, N71, N2074);
buf BUF1 (N3119, N3114);
xor XOR2 (N3120, N3096, N57);
nand NAND2 (N3121, N3119, N2431);
buf BUF1 (N3122, N3115);
or OR4 (N3123, N3120, N2707, N2892, N64);
nand NAND4 (N3124, N3092, N992, N898, N1234);
nor NOR2 (N3125, N3123, N2857);
xor XOR2 (N3126, N3118, N2324);
nand NAND3 (N3127, N3116, N388, N1707);
nor NOR3 (N3128, N3125, N351, N2306);
nor NOR2 (N3129, N3124, N2853);
buf BUF1 (N3130, N3110);
or OR3 (N3131, N3129, N2537, N2421);
or OR4 (N3132, N3122, N1553, N1073, N944);
nand NAND2 (N3133, N3127, N2176);
nand NAND2 (N3134, N3104, N2038);
buf BUF1 (N3135, N3117);
and AND2 (N3136, N3121, N617);
and AND4 (N3137, N3126, N2398, N3053, N1199);
xor XOR2 (N3138, N3134, N2149);
xor XOR2 (N3139, N3131, N944);
buf BUF1 (N3140, N3135);
not NOT1 (N3141, N3136);
nor NOR3 (N3142, N3137, N3003, N2143);
or OR4 (N3143, N3133, N3069, N2758, N919);
nand NAND3 (N3144, N3138, N2138, N879);
buf BUF1 (N3145, N3140);
or OR3 (N3146, N3141, N2009, N813);
nand NAND3 (N3147, N3130, N2127, N291);
or OR4 (N3148, N3146, N1731, N906, N728);
xor XOR2 (N3149, N3142, N155);
not NOT1 (N3150, N3147);
and AND4 (N3151, N3144, N1737, N1096, N445);
nor NOR3 (N3152, N3139, N1977, N358);
nor NOR4 (N3153, N3149, N1416, N675, N2513);
buf BUF1 (N3154, N3128);
nor NOR3 (N3155, N3112, N1223, N1393);
buf BUF1 (N3156, N3154);
nor NOR2 (N3157, N3152, N134);
not NOT1 (N3158, N3156);
nor NOR3 (N3159, N3157, N1670, N1572);
xor XOR2 (N3160, N3143, N2991);
not NOT1 (N3161, N3155);
and AND3 (N3162, N3158, N1357, N3113);
or OR2 (N3163, N3153, N1812);
and AND3 (N3164, N3161, N93, N3085);
buf BUF1 (N3165, N3160);
or OR2 (N3166, N3132, N406);
buf BUF1 (N3167, N3150);
and AND3 (N3168, N3163, N835, N2516);
or OR2 (N3169, N3162, N2452);
nor NOR4 (N3170, N3159, N2618, N1368, N1937);
and AND4 (N3171, N3165, N2621, N2456, N2954);
buf BUF1 (N3172, N3145);
or OR2 (N3173, N3151, N1760);
and AND2 (N3174, N3170, N496);
xor XOR2 (N3175, N3168, N2620);
and AND2 (N3176, N3166, N141);
nand NAND2 (N3177, N3176, N1474);
xor XOR2 (N3178, N3172, N2521);
or OR3 (N3179, N3164, N2499, N2523);
and AND2 (N3180, N3171, N2168);
or OR4 (N3181, N3167, N2249, N1476, N466);
xor XOR2 (N3182, N3179, N1090);
buf BUF1 (N3183, N3174);
buf BUF1 (N3184, N3175);
nor NOR3 (N3185, N3180, N1965, N437);
not NOT1 (N3186, N3182);
nor NOR2 (N3187, N3177, N443);
nor NOR2 (N3188, N3183, N1358);
xor XOR2 (N3189, N3173, N1203);
not NOT1 (N3190, N3148);
and AND3 (N3191, N3185, N545, N1778);
nor NOR2 (N3192, N3191, N1686);
buf BUF1 (N3193, N3192);
not NOT1 (N3194, N3193);
nand NAND2 (N3195, N3186, N2449);
xor XOR2 (N3196, N3188, N753);
and AND4 (N3197, N3196, N1781, N1804, N1560);
buf BUF1 (N3198, N3178);
xor XOR2 (N3199, N3184, N738);
nor NOR2 (N3200, N3195, N3069);
nand NAND2 (N3201, N3187, N164);
nand NAND4 (N3202, N3194, N656, N50, N2056);
xor XOR2 (N3203, N3169, N1982);
xor XOR2 (N3204, N3197, N2971);
or OR2 (N3205, N3199, N2169);
buf BUF1 (N3206, N3181);
nor NOR3 (N3207, N3202, N1880, N1624);
and AND4 (N3208, N3206, N309, N698, N701);
and AND3 (N3209, N3189, N425, N365);
not NOT1 (N3210, N3204);
not NOT1 (N3211, N3208);
or OR3 (N3212, N3203, N2078, N1670);
buf BUF1 (N3213, N3209);
nand NAND3 (N3214, N3205, N322, N567);
nor NOR4 (N3215, N3198, N1592, N2123, N2821);
xor XOR2 (N3216, N3212, N3124);
nor NOR3 (N3217, N3200, N1337, N3038);
not NOT1 (N3218, N3210);
buf BUF1 (N3219, N3201);
nand NAND4 (N3220, N3214, N1145, N2493, N2860);
and AND3 (N3221, N3207, N2087, N671);
xor XOR2 (N3222, N3220, N1894);
nand NAND4 (N3223, N3213, N689, N386, N786);
and AND4 (N3224, N3215, N1346, N876, N1125);
or OR3 (N3225, N3211, N1449, N1378);
buf BUF1 (N3226, N3219);
or OR2 (N3227, N3226, N2117);
buf BUF1 (N3228, N3216);
and AND4 (N3229, N3190, N1835, N1213, N1383);
buf BUF1 (N3230, N3223);
and AND3 (N3231, N3228, N2202, N2800);
nor NOR3 (N3232, N3217, N2330, N548);
nand NAND4 (N3233, N3222, N2307, N3061, N2258);
buf BUF1 (N3234, N3232);
nand NAND4 (N3235, N3230, N331, N2327, N2460);
and AND4 (N3236, N3224, N1306, N272, N1523);
buf BUF1 (N3237, N3231);
nor NOR3 (N3238, N3229, N3022, N1323);
xor XOR2 (N3239, N3233, N457);
and AND4 (N3240, N3235, N2458, N1986, N1933);
xor XOR2 (N3241, N3238, N736);
nand NAND3 (N3242, N3221, N33, N641);
or OR2 (N3243, N3234, N2003);
not NOT1 (N3244, N3240);
nand NAND3 (N3245, N3242, N3200, N3127);
or OR3 (N3246, N3245, N171, N3077);
not NOT1 (N3247, N3244);
xor XOR2 (N3248, N3246, N1176);
nand NAND3 (N3249, N3247, N1794, N138);
not NOT1 (N3250, N3237);
and AND2 (N3251, N3250, N1839);
buf BUF1 (N3252, N3239);
nor NOR3 (N3253, N3251, N186, N2266);
or OR4 (N3254, N3253, N1218, N2485, N1181);
nor NOR2 (N3255, N3227, N1142);
nand NAND2 (N3256, N3255, N2532);
not NOT1 (N3257, N3225);
nor NOR4 (N3258, N3252, N1977, N928, N3242);
and AND3 (N3259, N3257, N2471, N824);
not NOT1 (N3260, N3218);
buf BUF1 (N3261, N3260);
nor NOR4 (N3262, N3258, N2185, N2878, N1031);
nor NOR2 (N3263, N3249, N3148);
and AND4 (N3264, N3236, N2296, N3127, N3210);
nand NAND2 (N3265, N3261, N2194);
and AND4 (N3266, N3262, N1886, N2333, N505);
nand NAND2 (N3267, N3263, N2861);
nand NAND3 (N3268, N3266, N3254, N700);
xor XOR2 (N3269, N3243, N2830);
nor NOR3 (N3270, N2121, N2435, N828);
buf BUF1 (N3271, N3269);
nor NOR3 (N3272, N3259, N1909, N2208);
and AND3 (N3273, N3248, N1372, N1478);
or OR3 (N3274, N3268, N2757, N3013);
buf BUF1 (N3275, N3270);
xor XOR2 (N3276, N3264, N481);
not NOT1 (N3277, N3256);
and AND4 (N3278, N3265, N1132, N658, N1308);
nand NAND3 (N3279, N3278, N5, N1061);
buf BUF1 (N3280, N3277);
not NOT1 (N3281, N3273);
nand NAND3 (N3282, N3279, N44, N1808);
nand NAND3 (N3283, N3272, N1044, N790);
or OR3 (N3284, N3282, N2532, N1402);
xor XOR2 (N3285, N3274, N2376);
buf BUF1 (N3286, N3283);
nand NAND4 (N3287, N3280, N1528, N828, N1815);
nand NAND4 (N3288, N3285, N1304, N207, N1057);
nor NOR2 (N3289, N3241, N2381);
nand NAND3 (N3290, N3275, N2016, N2679);
xor XOR2 (N3291, N3281, N1037);
and AND4 (N3292, N3267, N1074, N3074, N3157);
nand NAND4 (N3293, N3284, N1322, N2265, N1141);
buf BUF1 (N3294, N3287);
nor NOR4 (N3295, N3291, N2150, N2618, N1231);
not NOT1 (N3296, N3293);
not NOT1 (N3297, N3288);
and AND2 (N3298, N3294, N2810);
and AND2 (N3299, N3290, N1768);
nand NAND3 (N3300, N3296, N2836, N1671);
nor NOR3 (N3301, N3299, N86, N2398);
not NOT1 (N3302, N3289);
nor NOR4 (N3303, N3302, N3022, N2414, N1941);
buf BUF1 (N3304, N3301);
or OR4 (N3305, N3292, N2272, N2940, N1071);
nor NOR4 (N3306, N3303, N16, N3022, N1321);
nor NOR3 (N3307, N3305, N2902, N3190);
or OR2 (N3308, N3271, N1435);
nor NOR4 (N3309, N3304, N203, N2844, N570);
or OR3 (N3310, N3309, N2437, N2284);
xor XOR2 (N3311, N3286, N721);
nand NAND2 (N3312, N3300, N1937);
buf BUF1 (N3313, N3276);
or OR2 (N3314, N3308, N1781);
nand NAND3 (N3315, N3311, N1386, N1100);
nor NOR3 (N3316, N3312, N1611, N2053);
or OR3 (N3317, N3307, N1642, N1448);
not NOT1 (N3318, N3297);
not NOT1 (N3319, N3310);
xor XOR2 (N3320, N3314, N3177);
xor XOR2 (N3321, N3320, N2814);
xor XOR2 (N3322, N3317, N1929);
nor NOR4 (N3323, N3319, N1475, N1489, N588);
buf BUF1 (N3324, N3315);
buf BUF1 (N3325, N3298);
buf BUF1 (N3326, N3322);
not NOT1 (N3327, N3323);
buf BUF1 (N3328, N3318);
buf BUF1 (N3329, N3295);
nand NAND3 (N3330, N3328, N61, N2158);
buf BUF1 (N3331, N3321);
not NOT1 (N3332, N3329);
nand NAND2 (N3333, N3313, N272);
nand NAND2 (N3334, N3306, N449);
or OR3 (N3335, N3334, N1601, N1256);
nand NAND2 (N3336, N3332, N2203);
buf BUF1 (N3337, N3336);
xor XOR2 (N3338, N3335, N3251);
buf BUF1 (N3339, N3316);
buf BUF1 (N3340, N3326);
not NOT1 (N3341, N3340);
and AND3 (N3342, N3330, N1176, N1377);
and AND2 (N3343, N3337, N2148);
nand NAND2 (N3344, N3338, N2926);
nor NOR4 (N3345, N3333, N114, N1039, N2819);
and AND4 (N3346, N3325, N999, N619, N3289);
and AND4 (N3347, N3331, N173, N190, N1337);
nand NAND4 (N3348, N3341, N1598, N467, N1701);
nand NAND4 (N3349, N3348, N1521, N2605, N608);
nor NOR2 (N3350, N3345, N1687);
or OR3 (N3351, N3343, N550, N1879);
or OR2 (N3352, N3339, N1993);
nand NAND2 (N3353, N3342, N2717);
xor XOR2 (N3354, N3344, N2648);
and AND4 (N3355, N3354, N1974, N716, N2316);
nor NOR4 (N3356, N3355, N410, N2678, N170);
nor NOR2 (N3357, N3352, N740);
xor XOR2 (N3358, N3346, N2928);
or OR2 (N3359, N3357, N909);
or OR2 (N3360, N3358, N296);
or OR4 (N3361, N3324, N1442, N2535, N2409);
and AND2 (N3362, N3349, N1728);
nand NAND3 (N3363, N3356, N3292, N1946);
nor NOR3 (N3364, N3360, N700, N1030);
or OR2 (N3365, N3347, N427);
nor NOR2 (N3366, N3364, N2143);
and AND2 (N3367, N3350, N2087);
not NOT1 (N3368, N3363);
not NOT1 (N3369, N3351);
nor NOR2 (N3370, N3367, N66);
nor NOR2 (N3371, N3365, N2915);
xor XOR2 (N3372, N3366, N1527);
or OR4 (N3373, N3362, N78, N1533, N1778);
buf BUF1 (N3374, N3327);
and AND4 (N3375, N3369, N2284, N2669, N2769);
nand NAND3 (N3376, N3373, N2483, N1584);
xor XOR2 (N3377, N3368, N991);
nor NOR3 (N3378, N3370, N1365, N1189);
and AND2 (N3379, N3378, N1866);
xor XOR2 (N3380, N3353, N2167);
xor XOR2 (N3381, N3371, N2245);
and AND3 (N3382, N3377, N1026, N3093);
nor NOR2 (N3383, N3361, N2845);
xor XOR2 (N3384, N3372, N1279);
or OR4 (N3385, N3382, N929, N3161, N3272);
and AND2 (N3386, N3359, N2083);
buf BUF1 (N3387, N3375);
and AND3 (N3388, N3381, N360, N3216);
nor NOR4 (N3389, N3376, N1317, N265, N1158);
or OR3 (N3390, N3388, N1586, N1203);
nor NOR4 (N3391, N3390, N2884, N3296, N3257);
and AND4 (N3392, N3389, N2065, N347, N781);
not NOT1 (N3393, N3392);
buf BUF1 (N3394, N3384);
or OR4 (N3395, N3391, N2611, N631, N2614);
nor NOR2 (N3396, N3385, N2517);
nor NOR3 (N3397, N3387, N1827, N1128);
not NOT1 (N3398, N3374);
nor NOR4 (N3399, N3398, N2352, N2440, N1316);
xor XOR2 (N3400, N3394, N2208);
xor XOR2 (N3401, N3393, N2831);
buf BUF1 (N3402, N3383);
buf BUF1 (N3403, N3379);
buf BUF1 (N3404, N3399);
not NOT1 (N3405, N3380);
buf BUF1 (N3406, N3397);
buf BUF1 (N3407, N3400);
nor NOR2 (N3408, N3395, N127);
and AND2 (N3409, N3406, N2049);
not NOT1 (N3410, N3404);
nand NAND4 (N3411, N3409, N1064, N2797, N11);
nand NAND2 (N3412, N3410, N2035);
buf BUF1 (N3413, N3402);
not NOT1 (N3414, N3411);
buf BUF1 (N3415, N3401);
not NOT1 (N3416, N3405);
nor NOR3 (N3417, N3412, N1347, N895);
or OR3 (N3418, N3415, N2172, N883);
nand NAND2 (N3419, N3418, N2017);
not NOT1 (N3420, N3413);
nand NAND3 (N3421, N3416, N1442, N3293);
not NOT1 (N3422, N3408);
nand NAND2 (N3423, N3386, N2202);
or OR4 (N3424, N3421, N1849, N1623, N2466);
not NOT1 (N3425, N3423);
nand NAND4 (N3426, N3420, N2548, N3156, N1386);
or OR4 (N3427, N3403, N1072, N1647, N1579);
buf BUF1 (N3428, N3407);
and AND3 (N3429, N3422, N2191, N2782);
nand NAND4 (N3430, N3424, N2888, N1511, N546);
xor XOR2 (N3431, N3428, N526);
nor NOR3 (N3432, N3429, N2118, N2946);
and AND2 (N3433, N3430, N2721);
nor NOR2 (N3434, N3414, N2362);
or OR3 (N3435, N3433, N165, N474);
not NOT1 (N3436, N3431);
xor XOR2 (N3437, N3432, N3160);
buf BUF1 (N3438, N3435);
nand NAND4 (N3439, N3434, N1587, N1720, N1164);
buf BUF1 (N3440, N3439);
nand NAND3 (N3441, N3417, N1012, N184);
xor XOR2 (N3442, N3437, N3092);
xor XOR2 (N3443, N3440, N2331);
not NOT1 (N3444, N3396);
not NOT1 (N3445, N3443);
xor XOR2 (N3446, N3419, N3058);
nor NOR3 (N3447, N3446, N3086, N198);
xor XOR2 (N3448, N3427, N1233);
nand NAND2 (N3449, N3448, N1617);
not NOT1 (N3450, N3445);
not NOT1 (N3451, N3450);
or OR3 (N3452, N3426, N3237, N1049);
nand NAND3 (N3453, N3441, N1836, N2120);
nand NAND4 (N3454, N3451, N2036, N3245, N3057);
or OR4 (N3455, N3452, N2990, N3189, N989);
buf BUF1 (N3456, N3444);
or OR2 (N3457, N3447, N2470);
nand NAND2 (N3458, N3438, N2755);
xor XOR2 (N3459, N3457, N2721);
not NOT1 (N3460, N3455);
nor NOR2 (N3461, N3460, N2035);
buf BUF1 (N3462, N3436);
xor XOR2 (N3463, N3459, N693);
nand NAND3 (N3464, N3458, N41, N962);
nor NOR3 (N3465, N3464, N2907, N1389);
buf BUF1 (N3466, N3465);
and AND2 (N3467, N3449, N2323);
buf BUF1 (N3468, N3462);
buf BUF1 (N3469, N3461);
nor NOR2 (N3470, N3453, N2580);
buf BUF1 (N3471, N3466);
buf BUF1 (N3472, N3454);
nor NOR3 (N3473, N3472, N3213, N570);
or OR4 (N3474, N3442, N982, N1720, N1687);
nor NOR2 (N3475, N3469, N3092);
nand NAND4 (N3476, N3467, N1122, N3354, N870);
and AND2 (N3477, N3470, N928);
nand NAND4 (N3478, N3476, N2837, N1655, N2979);
buf BUF1 (N3479, N3475);
xor XOR2 (N3480, N3425, N1131);
nand NAND3 (N3481, N3480, N2355, N2485);
nor NOR3 (N3482, N3477, N960, N2398);
buf BUF1 (N3483, N3482);
buf BUF1 (N3484, N3483);
xor XOR2 (N3485, N3468, N2376);
buf BUF1 (N3486, N3479);
and AND2 (N3487, N3471, N3335);
or OR3 (N3488, N3463, N2393, N852);
xor XOR2 (N3489, N3484, N1750);
xor XOR2 (N3490, N3481, N3179);
or OR2 (N3491, N3456, N2143);
or OR3 (N3492, N3485, N2173, N1312);
nor NOR4 (N3493, N3491, N2048, N3461, N84);
nor NOR3 (N3494, N3478, N1394, N1531);
buf BUF1 (N3495, N3488);
nand NAND4 (N3496, N3473, N3386, N2375, N2122);
and AND4 (N3497, N3493, N1231, N2542, N2523);
buf BUF1 (N3498, N3494);
xor XOR2 (N3499, N3498, N156);
xor XOR2 (N3500, N3499, N1913);
buf BUF1 (N3501, N3487);
not NOT1 (N3502, N3495);
nand NAND3 (N3503, N3486, N2732, N2009);
nand NAND3 (N3504, N3502, N2142, N2558);
or OR2 (N3505, N3474, N1554);
not NOT1 (N3506, N3501);
nor NOR3 (N3507, N3503, N1731, N3417);
not NOT1 (N3508, N3496);
and AND2 (N3509, N3508, N2472);
xor XOR2 (N3510, N3490, N2235);
xor XOR2 (N3511, N3497, N2305);
or OR2 (N3512, N3509, N2698);
not NOT1 (N3513, N3489);
nor NOR4 (N3514, N3505, N1865, N3344, N1910);
not NOT1 (N3515, N3504);
buf BUF1 (N3516, N3500);
or OR4 (N3517, N3506, N2340, N1454, N2765);
or OR3 (N3518, N3507, N3092, N1847);
and AND4 (N3519, N3516, N549, N1454, N454);
buf BUF1 (N3520, N3511);
buf BUF1 (N3521, N3520);
or OR4 (N3522, N3512, N1891, N3162, N3145);
nand NAND3 (N3523, N3518, N3097, N2720);
or OR3 (N3524, N3515, N3137, N3007);
nor NOR4 (N3525, N3519, N1513, N303, N90);
nor NOR4 (N3526, N3514, N418, N1330, N1116);
and AND3 (N3527, N3510, N2739, N80);
and AND4 (N3528, N3521, N1105, N1486, N1508);
or OR3 (N3529, N3525, N2465, N3398);
buf BUF1 (N3530, N3524);
and AND3 (N3531, N3517, N2545, N364);
buf BUF1 (N3532, N3526);
nand NAND4 (N3533, N3529, N3492, N995, N1958);
or OR4 (N3534, N1672, N2411, N3056, N1471);
or OR2 (N3535, N3513, N2077);
xor XOR2 (N3536, N3522, N184);
nor NOR3 (N3537, N3527, N2768, N2202);
buf BUF1 (N3538, N3528);
not NOT1 (N3539, N3538);
and AND4 (N3540, N3530, N664, N3245, N1037);
buf BUF1 (N3541, N3523);
buf BUF1 (N3542, N3536);
xor XOR2 (N3543, N3539, N1051);
buf BUF1 (N3544, N3541);
buf BUF1 (N3545, N3540);
buf BUF1 (N3546, N3531);
buf BUF1 (N3547, N3534);
xor XOR2 (N3548, N3543, N1144);
buf BUF1 (N3549, N3533);
or OR3 (N3550, N3545, N3503, N2574);
and AND2 (N3551, N3535, N425);
nand NAND3 (N3552, N3542, N783, N2877);
and AND2 (N3553, N3532, N794);
xor XOR2 (N3554, N3547, N3321);
buf BUF1 (N3555, N3544);
buf BUF1 (N3556, N3537);
xor XOR2 (N3557, N3553, N164);
nor NOR3 (N3558, N3555, N2768, N2516);
buf BUF1 (N3559, N3549);
nor NOR3 (N3560, N3551, N578, N2673);
nor NOR2 (N3561, N3559, N61);
buf BUF1 (N3562, N3548);
not NOT1 (N3563, N3552);
xor XOR2 (N3564, N3558, N799);
nand NAND4 (N3565, N3564, N188, N3531, N3031);
not NOT1 (N3566, N3550);
nor NOR2 (N3567, N3560, N1209);
nand NAND4 (N3568, N3557, N1394, N173, N1117);
nor NOR3 (N3569, N3546, N504, N238);
and AND2 (N3570, N3562, N1072);
not NOT1 (N3571, N3563);
nand NAND3 (N3572, N3565, N1959, N2988);
xor XOR2 (N3573, N3572, N1785);
and AND2 (N3574, N3568, N2175);
xor XOR2 (N3575, N3573, N2345);
and AND3 (N3576, N3556, N42, N751);
or OR4 (N3577, N3554, N1695, N79, N1057);
xor XOR2 (N3578, N3570, N115);
not NOT1 (N3579, N3561);
nor NOR3 (N3580, N3567, N2414, N120);
buf BUF1 (N3581, N3576);
xor XOR2 (N3582, N3574, N223);
not NOT1 (N3583, N3569);
nor NOR2 (N3584, N3575, N108);
or OR4 (N3585, N3577, N3145, N3046, N313);
nand NAND3 (N3586, N3584, N356, N158);
and AND2 (N3587, N3586, N2441);
nor NOR4 (N3588, N3585, N1737, N1844, N1162);
xor XOR2 (N3589, N3579, N1603);
and AND4 (N3590, N3588, N2395, N3250, N1292);
not NOT1 (N3591, N3583);
not NOT1 (N3592, N3591);
nand NAND3 (N3593, N3571, N269, N2097);
or OR2 (N3594, N3582, N253);
not NOT1 (N3595, N3581);
or OR4 (N3596, N3566, N1196, N451, N882);
not NOT1 (N3597, N3593);
and AND4 (N3598, N3597, N617, N1065, N1730);
and AND3 (N3599, N3595, N1879, N937);
not NOT1 (N3600, N3596);
xor XOR2 (N3601, N3580, N3536);
not NOT1 (N3602, N3598);
not NOT1 (N3603, N3587);
and AND2 (N3604, N3603, N131);
xor XOR2 (N3605, N3602, N3538);
xor XOR2 (N3606, N3590, N2902);
and AND2 (N3607, N3606, N754);
nand NAND2 (N3608, N3604, N2216);
nor NOR2 (N3609, N3605, N3296);
nor NOR4 (N3610, N3601, N3246, N37, N1702);
not NOT1 (N3611, N3607);
and AND3 (N3612, N3589, N190, N431);
not NOT1 (N3613, N3594);
or OR4 (N3614, N3592, N2543, N2048, N859);
nand NAND2 (N3615, N3600, N3287);
xor XOR2 (N3616, N3610, N2811);
nor NOR2 (N3617, N3599, N220);
nand NAND3 (N3618, N3617, N2700, N2899);
nor NOR2 (N3619, N3618, N1907);
nor NOR4 (N3620, N3615, N1201, N435, N2993);
buf BUF1 (N3621, N3608);
not NOT1 (N3622, N3619);
not NOT1 (N3623, N3614);
nand NAND4 (N3624, N3623, N643, N1431, N3467);
nor NOR3 (N3625, N3611, N2510, N2108);
nor NOR3 (N3626, N3624, N1304, N982);
not NOT1 (N3627, N3612);
or OR4 (N3628, N3616, N2560, N3142, N2178);
and AND3 (N3629, N3621, N2277, N1026);
xor XOR2 (N3630, N3626, N2238);
or OR3 (N3631, N3629, N2872, N2187);
xor XOR2 (N3632, N3625, N1539);
xor XOR2 (N3633, N3620, N1273);
buf BUF1 (N3634, N3628);
nand NAND2 (N3635, N3578, N697);
xor XOR2 (N3636, N3630, N1181);
nor NOR2 (N3637, N3633, N1620);
not NOT1 (N3638, N3635);
nor NOR4 (N3639, N3634, N2948, N3461, N1981);
and AND3 (N3640, N3632, N733, N3007);
not NOT1 (N3641, N3636);
buf BUF1 (N3642, N3609);
not NOT1 (N3643, N3640);
xor XOR2 (N3644, N3643, N232);
xor XOR2 (N3645, N3613, N2169);
nand NAND3 (N3646, N3637, N2535, N137);
buf BUF1 (N3647, N3641);
nand NAND2 (N3648, N3627, N3135);
and AND3 (N3649, N3646, N3134, N2404);
nand NAND2 (N3650, N3647, N1219);
not NOT1 (N3651, N3645);
or OR2 (N3652, N3650, N2225);
not NOT1 (N3653, N3638);
xor XOR2 (N3654, N3642, N2550);
nor NOR2 (N3655, N3654, N2188);
or OR2 (N3656, N3649, N2262);
buf BUF1 (N3657, N3622);
or OR2 (N3658, N3631, N2454);
nor NOR3 (N3659, N3657, N2951, N701);
nand NAND2 (N3660, N3653, N2445);
or OR4 (N3661, N3658, N3072, N288, N2476);
nor NOR3 (N3662, N3661, N1590, N2654);
nor NOR2 (N3663, N3659, N2380);
or OR2 (N3664, N3652, N3548);
or OR2 (N3665, N3656, N610);
xor XOR2 (N3666, N3664, N2184);
and AND3 (N3667, N3655, N569, N3242);
buf BUF1 (N3668, N3660);
and AND4 (N3669, N3651, N2747, N3386, N1801);
nand NAND2 (N3670, N3667, N2294);
xor XOR2 (N3671, N3644, N159);
nand NAND3 (N3672, N3666, N1430, N551);
and AND4 (N3673, N3662, N2744, N2039, N1809);
and AND4 (N3674, N3668, N2342, N2395, N232);
nand NAND3 (N3675, N3648, N2969, N796);
nand NAND2 (N3676, N3669, N1371);
nand NAND2 (N3677, N3676, N2324);
not NOT1 (N3678, N3674);
or OR4 (N3679, N3672, N1550, N3440, N675);
and AND4 (N3680, N3639, N753, N3417, N2090);
not NOT1 (N3681, N3670);
buf BUF1 (N3682, N3678);
buf BUF1 (N3683, N3665);
xor XOR2 (N3684, N3663, N3331);
or OR3 (N3685, N3682, N1073, N2329);
buf BUF1 (N3686, N3680);
nor NOR2 (N3687, N3686, N3073);
nand NAND4 (N3688, N3681, N2546, N68, N2220);
or OR3 (N3689, N3673, N662, N3286);
buf BUF1 (N3690, N3677);
and AND4 (N3691, N3683, N1401, N1508, N1333);
xor XOR2 (N3692, N3689, N2294);
nor NOR3 (N3693, N3671, N1749, N3232);
and AND3 (N3694, N3693, N1401, N3622);
nor NOR3 (N3695, N3679, N2145, N2602);
or OR4 (N3696, N3687, N352, N2652, N2256);
nand NAND4 (N3697, N3684, N1456, N2487, N3422);
nor NOR2 (N3698, N3690, N2516);
not NOT1 (N3699, N3685);
or OR2 (N3700, N3675, N3684);
and AND2 (N3701, N3697, N2233);
xor XOR2 (N3702, N3688, N55);
or OR3 (N3703, N3698, N2485, N3679);
not NOT1 (N3704, N3703);
nor NOR2 (N3705, N3696, N2469);
xor XOR2 (N3706, N3700, N2404);
and AND3 (N3707, N3701, N1112, N759);
not NOT1 (N3708, N3704);
nor NOR2 (N3709, N3692, N1370);
not NOT1 (N3710, N3707);
xor XOR2 (N3711, N3709, N638);
not NOT1 (N3712, N3710);
buf BUF1 (N3713, N3711);
or OR3 (N3714, N3691, N3687, N2617);
nor NOR2 (N3715, N3699, N1401);
nand NAND2 (N3716, N3713, N476);
and AND4 (N3717, N3714, N1719, N1115, N2824);
nand NAND4 (N3718, N3712, N1971, N1111, N1556);
xor XOR2 (N3719, N3706, N1662);
nor NOR2 (N3720, N3715, N1301);
xor XOR2 (N3721, N3695, N2522);
nor NOR2 (N3722, N3720, N2984);
nor NOR2 (N3723, N3721, N3716);
not NOT1 (N3724, N2965);
buf BUF1 (N3725, N3705);
buf BUF1 (N3726, N3708);
buf BUF1 (N3727, N3723);
or OR2 (N3728, N3718, N2534);
or OR4 (N3729, N3724, N745, N3238, N2823);
buf BUF1 (N3730, N3729);
nand NAND3 (N3731, N3702, N2930, N1602);
or OR4 (N3732, N3719, N3534, N1800, N527);
nand NAND4 (N3733, N3730, N2922, N1111, N1323);
or OR2 (N3734, N3728, N104);
nand NAND3 (N3735, N3732, N2901, N619);
nand NAND3 (N3736, N3727, N2774, N279);
xor XOR2 (N3737, N3725, N385);
and AND4 (N3738, N3717, N1402, N1544, N2560);
xor XOR2 (N3739, N3733, N3482);
nor NOR3 (N3740, N3739, N2322, N2401);
xor XOR2 (N3741, N3722, N1433);
xor XOR2 (N3742, N3734, N3317);
or OR4 (N3743, N3742, N1105, N2442, N639);
nand NAND4 (N3744, N3737, N293, N1254, N765);
nand NAND2 (N3745, N3694, N1538);
or OR3 (N3746, N3744, N2275, N3299);
and AND2 (N3747, N3736, N2183);
not NOT1 (N3748, N3731);
xor XOR2 (N3749, N3747, N709);
or OR3 (N3750, N3726, N2611, N2885);
xor XOR2 (N3751, N3750, N3029);
and AND3 (N3752, N3751, N2042, N895);
buf BUF1 (N3753, N3748);
or OR4 (N3754, N3741, N1155, N2637, N830);
buf BUF1 (N3755, N3735);
xor XOR2 (N3756, N3743, N1545);
and AND4 (N3757, N3752, N800, N3373, N1042);
nand NAND2 (N3758, N3754, N3466);
buf BUF1 (N3759, N3738);
or OR3 (N3760, N3756, N933, N2589);
not NOT1 (N3761, N3753);
or OR2 (N3762, N3746, N1371);
buf BUF1 (N3763, N3761);
xor XOR2 (N3764, N3755, N2506);
not NOT1 (N3765, N3749);
or OR2 (N3766, N3757, N1430);
nor NOR2 (N3767, N3766, N3540);
nand NAND4 (N3768, N3759, N898, N2006, N630);
or OR4 (N3769, N3745, N2191, N2814, N753);
nand NAND2 (N3770, N3763, N517);
buf BUF1 (N3771, N3760);
xor XOR2 (N3772, N3769, N308);
xor XOR2 (N3773, N3770, N353);
xor XOR2 (N3774, N3767, N3304);
nand NAND2 (N3775, N3762, N2351);
buf BUF1 (N3776, N3774);
not NOT1 (N3777, N3768);
buf BUF1 (N3778, N3765);
nand NAND4 (N3779, N3764, N2124, N2349, N3657);
nand NAND2 (N3780, N3777, N1734);
buf BUF1 (N3781, N3772);
nand NAND4 (N3782, N3780, N14, N1919, N2667);
buf BUF1 (N3783, N3758);
nand NAND3 (N3784, N3783, N3599, N2550);
and AND2 (N3785, N3771, N2955);
xor XOR2 (N3786, N3773, N3498);
buf BUF1 (N3787, N3775);
nand NAND4 (N3788, N3786, N2288, N2769, N1324);
nor NOR2 (N3789, N3788, N1384);
and AND3 (N3790, N3776, N746, N2301);
buf BUF1 (N3791, N3790);
or OR4 (N3792, N3782, N2703, N3109, N649);
not NOT1 (N3793, N3792);
and AND4 (N3794, N3779, N591, N405, N1526);
nand NAND2 (N3795, N3787, N744);
and AND4 (N3796, N3778, N3144, N2487, N1028);
nor NOR2 (N3797, N3740, N1408);
not NOT1 (N3798, N3784);
nand NAND4 (N3799, N3785, N1598, N2140, N2733);
nor NOR3 (N3800, N3789, N1839, N352);
or OR4 (N3801, N3800, N1437, N873, N3739);
nand NAND4 (N3802, N3795, N1200, N2496, N2155);
buf BUF1 (N3803, N3781);
xor XOR2 (N3804, N3801, N2987);
or OR2 (N3805, N3802, N1588);
nand NAND4 (N3806, N3805, N2778, N2545, N1363);
nor NOR3 (N3807, N3803, N2788, N3323);
and AND3 (N3808, N3791, N818, N425);
buf BUF1 (N3809, N3796);
not NOT1 (N3810, N3799);
or OR3 (N3811, N3798, N1734, N2241);
xor XOR2 (N3812, N3811, N3398);
nor NOR2 (N3813, N3793, N2011);
xor XOR2 (N3814, N3806, N979);
or OR4 (N3815, N3804, N2111, N679, N2997);
buf BUF1 (N3816, N3814);
or OR2 (N3817, N3816, N3427);
not NOT1 (N3818, N3794);
buf BUF1 (N3819, N3809);
buf BUF1 (N3820, N3807);
buf BUF1 (N3821, N3819);
or OR3 (N3822, N3821, N2175, N2302);
or OR3 (N3823, N3818, N219, N785);
buf BUF1 (N3824, N3822);
or OR2 (N3825, N3824, N3462);
nand NAND2 (N3826, N3823, N1979);
or OR2 (N3827, N3825, N1685);
not NOT1 (N3828, N3820);
xor XOR2 (N3829, N3828, N3518);
not NOT1 (N3830, N3813);
or OR4 (N3831, N3797, N1852, N2297, N2188);
not NOT1 (N3832, N3815);
buf BUF1 (N3833, N3832);
or OR2 (N3834, N3808, N2533);
nor NOR3 (N3835, N3834, N1034, N557);
nand NAND4 (N3836, N3827, N548, N3188, N3703);
or OR4 (N3837, N3826, N3700, N270, N2279);
not NOT1 (N3838, N3817);
not NOT1 (N3839, N3830);
or OR2 (N3840, N3835, N1777);
or OR4 (N3841, N3838, N2802, N286, N3663);
nor NOR2 (N3842, N3810, N1241);
and AND3 (N3843, N3836, N3831, N1646);
or OR3 (N3844, N3129, N100, N2597);
xor XOR2 (N3845, N3844, N660);
nor NOR4 (N3846, N3837, N1899, N1255, N472);
nand NAND4 (N3847, N3846, N326, N1157, N64);
not NOT1 (N3848, N3829);
not NOT1 (N3849, N3847);
nor NOR2 (N3850, N3842, N2663);
not NOT1 (N3851, N3833);
xor XOR2 (N3852, N3841, N2769);
not NOT1 (N3853, N3839);
nand NAND4 (N3854, N3845, N3163, N1053, N438);
xor XOR2 (N3855, N3851, N3775);
not NOT1 (N3856, N3848);
not NOT1 (N3857, N3840);
buf BUF1 (N3858, N3852);
and AND2 (N3859, N3812, N3137);
or OR4 (N3860, N3849, N121, N3391, N1558);
nor NOR2 (N3861, N3860, N2165);
and AND2 (N3862, N3843, N391);
buf BUF1 (N3863, N3855);
nor NOR4 (N3864, N3854, N428, N3236, N776);
xor XOR2 (N3865, N3863, N1045);
and AND4 (N3866, N3862, N828, N1207, N3046);
not NOT1 (N3867, N3865);
not NOT1 (N3868, N3861);
nand NAND4 (N3869, N3864, N874, N1768, N1042);
or OR3 (N3870, N3869, N1386, N1959);
nand NAND4 (N3871, N3856, N1384, N3478, N2729);
not NOT1 (N3872, N3857);
buf BUF1 (N3873, N3853);
buf BUF1 (N3874, N3871);
nor NOR3 (N3875, N3873, N2740, N3252);
xor XOR2 (N3876, N3866, N3519);
buf BUF1 (N3877, N3868);
nor NOR3 (N3878, N3874, N2636, N1256);
or OR4 (N3879, N3876, N2798, N3457, N1201);
not NOT1 (N3880, N3867);
xor XOR2 (N3881, N3870, N743);
or OR4 (N3882, N3881, N431, N128, N1674);
and AND2 (N3883, N3859, N1601);
nand NAND4 (N3884, N3875, N1018, N228, N3188);
nor NOR3 (N3885, N3878, N2892, N3305);
and AND3 (N3886, N3858, N2528, N1849);
xor XOR2 (N3887, N3884, N3220);
and AND2 (N3888, N3850, N1306);
buf BUF1 (N3889, N3879);
and AND2 (N3890, N3887, N2967);
buf BUF1 (N3891, N3885);
nor NOR2 (N3892, N3891, N415);
or OR3 (N3893, N3888, N92, N2746);
or OR3 (N3894, N3893, N1266, N1203);
not NOT1 (N3895, N3872);
nand NAND3 (N3896, N3886, N2380, N2225);
not NOT1 (N3897, N3896);
nor NOR3 (N3898, N3880, N2684, N66);
buf BUF1 (N3899, N3890);
or OR2 (N3900, N3877, N49);
not NOT1 (N3901, N3898);
buf BUF1 (N3902, N3899);
buf BUF1 (N3903, N3882);
and AND2 (N3904, N3897, N1738);
nor NOR2 (N3905, N3903, N2342);
xor XOR2 (N3906, N3889, N1774);
nor NOR4 (N3907, N3894, N2879, N3015, N1788);
nor NOR4 (N3908, N3901, N424, N3195, N2851);
xor XOR2 (N3909, N3900, N33);
or OR2 (N3910, N3902, N3231);
not NOT1 (N3911, N3883);
nor NOR4 (N3912, N3907, N2228, N3873, N3432);
xor XOR2 (N3913, N3909, N3242);
buf BUF1 (N3914, N3912);
nor NOR4 (N3915, N3911, N9, N944, N1557);
or OR3 (N3916, N3910, N392, N3673);
not NOT1 (N3917, N3916);
nor NOR3 (N3918, N3917, N162, N2482);
not NOT1 (N3919, N3904);
or OR3 (N3920, N3905, N405, N1196);
not NOT1 (N3921, N3892);
xor XOR2 (N3922, N3914, N3899);
xor XOR2 (N3923, N3915, N3885);
buf BUF1 (N3924, N3913);
nand NAND4 (N3925, N3924, N538, N124, N2411);
or OR4 (N3926, N3922, N1998, N3029, N2877);
and AND2 (N3927, N3908, N3099);
nand NAND3 (N3928, N3918, N2390, N557);
buf BUF1 (N3929, N3895);
or OR2 (N3930, N3925, N1658);
or OR4 (N3931, N3919, N34, N2456, N723);
xor XOR2 (N3932, N3931, N2387);
buf BUF1 (N3933, N3921);
xor XOR2 (N3934, N3932, N3157);
nor NOR4 (N3935, N3927, N697, N536, N2564);
xor XOR2 (N3936, N3934, N1163);
not NOT1 (N3937, N3936);
xor XOR2 (N3938, N3923, N1363);
or OR3 (N3939, N3937, N336, N2794);
nand NAND2 (N3940, N3928, N2382);
and AND2 (N3941, N3938, N2290);
and AND3 (N3942, N3906, N3426, N2407);
nor NOR2 (N3943, N3933, N3396);
nand NAND3 (N3944, N3943, N728, N798);
buf BUF1 (N3945, N3944);
buf BUF1 (N3946, N3935);
xor XOR2 (N3947, N3926, N1944);
not NOT1 (N3948, N3920);
or OR3 (N3949, N3939, N704, N1756);
buf BUF1 (N3950, N3945);
or OR2 (N3951, N3946, N3425);
or OR4 (N3952, N3948, N356, N2230, N3355);
nand NAND4 (N3953, N3941, N960, N2876, N3038);
nor NOR3 (N3954, N3952, N600, N897);
not NOT1 (N3955, N3940);
nand NAND3 (N3956, N3947, N3410, N1373);
not NOT1 (N3957, N3942);
buf BUF1 (N3958, N3954);
xor XOR2 (N3959, N3955, N2335);
or OR4 (N3960, N3953, N3725, N2754, N1484);
not NOT1 (N3961, N3949);
nand NAND3 (N3962, N3951, N1389, N2657);
xor XOR2 (N3963, N3950, N2722);
not NOT1 (N3964, N3956);
and AND3 (N3965, N3960, N1767, N2980);
not NOT1 (N3966, N3963);
buf BUF1 (N3967, N3961);
nand NAND4 (N3968, N3965, N3761, N1777, N968);
nand NAND3 (N3969, N3930, N1734, N2129);
nor NOR2 (N3970, N3967, N1183);
xor XOR2 (N3971, N3968, N3535);
and AND2 (N3972, N3958, N2910);
and AND3 (N3973, N3964, N2859, N2761);
xor XOR2 (N3974, N3971, N185);
not NOT1 (N3975, N3929);
nand NAND4 (N3976, N3973, N1894, N2046, N3008);
not NOT1 (N3977, N3970);
nor NOR2 (N3978, N3966, N2869);
nor NOR4 (N3979, N3977, N1416, N3695, N870);
not NOT1 (N3980, N3959);
nor NOR4 (N3981, N3975, N1861, N2099, N3047);
and AND3 (N3982, N3979, N2543, N2308);
xor XOR2 (N3983, N3969, N368);
xor XOR2 (N3984, N3957, N2485);
xor XOR2 (N3985, N3974, N3087);
xor XOR2 (N3986, N3962, N2842);
or OR4 (N3987, N3982, N678, N592, N2612);
not NOT1 (N3988, N3972);
and AND4 (N3989, N3986, N619, N3060, N3199);
buf BUF1 (N3990, N3989);
nor NOR2 (N3991, N3988, N3804);
nor NOR4 (N3992, N3976, N725, N2334, N1467);
buf BUF1 (N3993, N3987);
buf BUF1 (N3994, N3985);
nor NOR2 (N3995, N3980, N622);
and AND2 (N3996, N3993, N2766);
nor NOR2 (N3997, N3981, N827);
buf BUF1 (N3998, N3983);
nand NAND3 (N3999, N3994, N1864, N1646);
buf BUF1 (N4000, N3998);
not NOT1 (N4001, N3996);
nor NOR3 (N4002, N3984, N1842, N2149);
nand NAND4 (N4003, N3991, N434, N2378, N2969);
not NOT1 (N4004, N3990);
nor NOR3 (N4005, N4003, N3193, N1057);
xor XOR2 (N4006, N3978, N2124);
and AND3 (N4007, N3992, N1802, N126);
and AND2 (N4008, N3999, N3406);
and AND3 (N4009, N4004, N641, N1409);
or OR4 (N4010, N4008, N2237, N3053, N2131);
xor XOR2 (N4011, N4002, N2561);
xor XOR2 (N4012, N4010, N3591);
and AND4 (N4013, N4009, N8, N3463, N3051);
not NOT1 (N4014, N4011);
buf BUF1 (N4015, N4005);
nand NAND2 (N4016, N4015, N3191);
or OR3 (N4017, N4016, N1007, N2436);
or OR4 (N4018, N4012, N3, N2697, N1430);
xor XOR2 (N4019, N3995, N731);
and AND2 (N4020, N4006, N2437);
nand NAND2 (N4021, N4017, N1379);
nor NOR2 (N4022, N4019, N1808);
nor NOR3 (N4023, N4020, N2810, N1911);
buf BUF1 (N4024, N4018);
xor XOR2 (N4025, N4000, N3740);
not NOT1 (N4026, N4001);
nand NAND2 (N4027, N4014, N3507);
not NOT1 (N4028, N4024);
not NOT1 (N4029, N4007);
or OR3 (N4030, N4029, N2, N2157);
not NOT1 (N4031, N4013);
or OR2 (N4032, N4026, N2317);
or OR3 (N4033, N4032, N3485, N879);
or OR2 (N4034, N4021, N715);
nand NAND2 (N4035, N4028, N416);
not NOT1 (N4036, N4035);
nand NAND4 (N4037, N4036, N1562, N206, N1537);
xor XOR2 (N4038, N4034, N4036);
not NOT1 (N4039, N4031);
xor XOR2 (N4040, N4039, N1386);
nand NAND3 (N4041, N4022, N712, N1257);
and AND3 (N4042, N4023, N2319, N2386);
and AND2 (N4043, N4042, N2615);
nand NAND2 (N4044, N4033, N3);
nor NOR3 (N4045, N4030, N3329, N390);
nor NOR3 (N4046, N3997, N291, N2857);
not NOT1 (N4047, N4037);
buf BUF1 (N4048, N4025);
buf BUF1 (N4049, N4047);
nand NAND4 (N4050, N4041, N2225, N2181, N2470);
nand NAND4 (N4051, N4027, N618, N2694, N644);
nand NAND2 (N4052, N4050, N2046);
not NOT1 (N4053, N4051);
not NOT1 (N4054, N4045);
xor XOR2 (N4055, N4048, N1008);
not NOT1 (N4056, N4054);
buf BUF1 (N4057, N4043);
or OR2 (N4058, N4057, N1089);
or OR2 (N4059, N4044, N3052);
and AND4 (N4060, N4049, N1479, N2449, N1618);
nand NAND3 (N4061, N4052, N1073, N1888);
or OR2 (N4062, N4055, N1353);
xor XOR2 (N4063, N4062, N1920);
nor NOR3 (N4064, N4058, N1214, N2540);
or OR2 (N4065, N4064, N1194);
not NOT1 (N4066, N4060);
nand NAND3 (N4067, N4066, N2730, N1741);
xor XOR2 (N4068, N4056, N3505);
nor NOR4 (N4069, N4068, N2998, N3804, N3459);
xor XOR2 (N4070, N4067, N943);
not NOT1 (N4071, N4070);
xor XOR2 (N4072, N4069, N326);
nand NAND2 (N4073, N4061, N192);
buf BUF1 (N4074, N4046);
xor XOR2 (N4075, N4040, N1448);
or OR2 (N4076, N4074, N827);
nand NAND4 (N4077, N4071, N720, N1697, N2313);
buf BUF1 (N4078, N4038);
xor XOR2 (N4079, N4063, N1893);
nor NOR4 (N4080, N4078, N1044, N1856, N2003);
xor XOR2 (N4081, N4077, N1602);
nor NOR2 (N4082, N4075, N803);
and AND4 (N4083, N4053, N100, N1178, N1027);
and AND2 (N4084, N4080, N680);
nor NOR3 (N4085, N4082, N1831, N2428);
or OR2 (N4086, N4072, N1519);
or OR4 (N4087, N4084, N1858, N1057, N3180);
xor XOR2 (N4088, N4083, N2333);
nand NAND4 (N4089, N4081, N2896, N2847, N3552);
nor NOR3 (N4090, N4089, N588, N2928);
and AND3 (N4091, N4090, N1017, N1260);
or OR4 (N4092, N4076, N645, N2009, N1540);
buf BUF1 (N4093, N4091);
not NOT1 (N4094, N4059);
nand NAND2 (N4095, N4073, N324);
and AND4 (N4096, N4087, N214, N2230, N939);
nor NOR2 (N4097, N4096, N3895);
xor XOR2 (N4098, N4079, N3613);
buf BUF1 (N4099, N4088);
nand NAND2 (N4100, N4095, N50);
nor NOR4 (N4101, N4092, N192, N2730, N4095);
not NOT1 (N4102, N4097);
buf BUF1 (N4103, N4101);
or OR3 (N4104, N4086, N3523, N1906);
or OR4 (N4105, N4065, N2635, N162, N914);
buf BUF1 (N4106, N4100);
nand NAND4 (N4107, N4085, N2967, N3399, N2856);
or OR2 (N4108, N4107, N3334);
nor NOR3 (N4109, N4094, N1654, N933);
xor XOR2 (N4110, N4098, N215);
nor NOR3 (N4111, N4103, N454, N3412);
nand NAND3 (N4112, N4111, N4034, N424);
nor NOR3 (N4113, N4108, N1070, N2649);
buf BUF1 (N4114, N4105);
nand NAND4 (N4115, N4104, N3027, N3057, N4110);
or OR3 (N4116, N2409, N1302, N2276);
and AND3 (N4117, N4093, N1040, N2120);
and AND2 (N4118, N4109, N1847);
nor NOR2 (N4119, N4112, N1652);
nand NAND3 (N4120, N4113, N1743, N1527);
nand NAND3 (N4121, N4114, N1940, N565);
nor NOR2 (N4122, N4099, N1018);
buf BUF1 (N4123, N4121);
or OR3 (N4124, N4102, N1888, N1208);
xor XOR2 (N4125, N4123, N3159);
buf BUF1 (N4126, N4118);
nand NAND4 (N4127, N4116, N3801, N455, N3818);
nor NOR3 (N4128, N4124, N2350, N1153);
or OR2 (N4129, N4127, N597);
nor NOR4 (N4130, N4128, N2098, N1252, N213);
and AND3 (N4131, N4119, N3630, N373);
nand NAND4 (N4132, N4126, N1851, N2239, N3465);
or OR4 (N4133, N4125, N1274, N1507, N1824);
nor NOR3 (N4134, N4122, N953, N1233);
not NOT1 (N4135, N4117);
and AND4 (N4136, N4134, N277, N575, N2584);
nor NOR4 (N4137, N4131, N846, N1884, N1214);
nor NOR4 (N4138, N4120, N1079, N905, N167);
xor XOR2 (N4139, N4132, N740);
and AND3 (N4140, N4135, N2947, N2885);
or OR2 (N4141, N4139, N2656);
buf BUF1 (N4142, N4129);
xor XOR2 (N4143, N4130, N3106);
and AND4 (N4144, N4136, N601, N3886, N2095);
not NOT1 (N4145, N4144);
not NOT1 (N4146, N4115);
nand NAND3 (N4147, N4106, N946, N1087);
nor NOR2 (N4148, N4141, N442);
nand NAND2 (N4149, N4133, N2660);
and AND2 (N4150, N4143, N1806);
or OR4 (N4151, N4140, N2232, N2198, N1062);
and AND4 (N4152, N4149, N4127, N40, N2803);
not NOT1 (N4153, N4151);
nand NAND3 (N4154, N4137, N3627, N1353);
buf BUF1 (N4155, N4150);
or OR2 (N4156, N4153, N1260);
nor NOR4 (N4157, N4138, N611, N1692, N376);
buf BUF1 (N4158, N4155);
and AND4 (N4159, N4147, N1618, N2141, N3401);
nand NAND4 (N4160, N4154, N3987, N2214, N3002);
xor XOR2 (N4161, N4160, N947);
buf BUF1 (N4162, N4161);
nand NAND2 (N4163, N4158, N1861);
nand NAND2 (N4164, N4163, N2670);
xor XOR2 (N4165, N4146, N1455);
nor NOR3 (N4166, N4157, N2917, N1547);
and AND4 (N4167, N4164, N2315, N922, N2728);
nor NOR2 (N4168, N4159, N4031);
nand NAND4 (N4169, N4145, N3934, N1039, N489);
not NOT1 (N4170, N4148);
not NOT1 (N4171, N4167);
nor NOR3 (N4172, N4169, N3676, N2579);
and AND4 (N4173, N4170, N1928, N2539, N2523);
nand NAND3 (N4174, N4162, N4001, N4010);
not NOT1 (N4175, N4172);
not NOT1 (N4176, N4156);
not NOT1 (N4177, N4176);
nand NAND2 (N4178, N4165, N2713);
and AND2 (N4179, N4173, N4150);
not NOT1 (N4180, N4175);
and AND4 (N4181, N4177, N3103, N2739, N674);
nor NOR2 (N4182, N4171, N2799);
nor NOR4 (N4183, N4180, N1717, N3500, N1199);
nand NAND3 (N4184, N4142, N4152, N1129);
or OR3 (N4185, N902, N2532, N3232);
buf BUF1 (N4186, N4182);
nor NOR3 (N4187, N4185, N3389, N2865);
buf BUF1 (N4188, N4181);
and AND3 (N4189, N4184, N905, N2590);
nor NOR2 (N4190, N4174, N3215);
nor NOR2 (N4191, N4190, N3325);
and AND3 (N4192, N4178, N3940, N3333);
nand NAND4 (N4193, N4188, N107, N1953, N2763);
or OR4 (N4194, N4186, N92, N2999, N1043);
not NOT1 (N4195, N4189);
nand NAND3 (N4196, N4179, N3596, N1450);
xor XOR2 (N4197, N4187, N3902);
or OR4 (N4198, N4183, N107, N3603, N1032);
buf BUF1 (N4199, N4168);
not NOT1 (N4200, N4193);
buf BUF1 (N4201, N4199);
xor XOR2 (N4202, N4195, N395);
not NOT1 (N4203, N4194);
xor XOR2 (N4204, N4192, N1686);
or OR4 (N4205, N4197, N2349, N1824, N1975);
and AND4 (N4206, N4196, N1120, N537, N3877);
nand NAND4 (N4207, N4198, N3346, N215, N702);
nor NOR3 (N4208, N4207, N2661, N3805);
not NOT1 (N4209, N4203);
nor NOR2 (N4210, N4166, N847);
xor XOR2 (N4211, N4202, N1659);
nand NAND3 (N4212, N4191, N2875, N2806);
and AND3 (N4213, N4201, N922, N255);
xor XOR2 (N4214, N4200, N1669);
xor XOR2 (N4215, N4206, N1217);
nor NOR3 (N4216, N4213, N3558, N506);
buf BUF1 (N4217, N4208);
nand NAND3 (N4218, N4211, N3762, N3594);
nand NAND2 (N4219, N4204, N1132);
not NOT1 (N4220, N4210);
or OR4 (N4221, N4215, N2342, N498, N1210);
nor NOR2 (N4222, N4219, N1489);
nor NOR4 (N4223, N4214, N1839, N596, N2763);
buf BUF1 (N4224, N4212);
nand NAND4 (N4225, N4218, N3635, N1486, N1906);
xor XOR2 (N4226, N4205, N2088);
and AND3 (N4227, N4225, N2605, N3556);
and AND2 (N4228, N4222, N3997);
nand NAND3 (N4229, N4226, N3157, N1713);
xor XOR2 (N4230, N4224, N3655);
not NOT1 (N4231, N4223);
and AND3 (N4232, N4221, N1324, N543);
nand NAND4 (N4233, N4217, N3478, N958, N3513);
not NOT1 (N4234, N4227);
nor NOR2 (N4235, N4234, N2518);
buf BUF1 (N4236, N4231);
buf BUF1 (N4237, N4235);
nor NOR4 (N4238, N4233, N16, N3178, N972);
nor NOR2 (N4239, N4237, N3243);
not NOT1 (N4240, N4239);
buf BUF1 (N4241, N4229);
not NOT1 (N4242, N4238);
xor XOR2 (N4243, N4242, N1153);
not NOT1 (N4244, N4232);
or OR2 (N4245, N4216, N3405);
not NOT1 (N4246, N4240);
nand NAND3 (N4247, N4243, N422, N2326);
nand NAND4 (N4248, N4244, N574, N1644, N1758);
not NOT1 (N4249, N4220);
nor NOR4 (N4250, N4247, N3407, N2149, N2376);
xor XOR2 (N4251, N4246, N2273);
xor XOR2 (N4252, N4241, N1672);
and AND3 (N4253, N4236, N1683, N2033);
buf BUF1 (N4254, N4249);
and AND4 (N4255, N4230, N92, N2409, N2553);
and AND3 (N4256, N4228, N3233, N480);
and AND3 (N4257, N4256, N1991, N3098);
xor XOR2 (N4258, N4257, N1600);
nand NAND4 (N4259, N4250, N3096, N3542, N3853);
not NOT1 (N4260, N4255);
not NOT1 (N4261, N4258);
nand NAND4 (N4262, N4248, N1214, N1439, N4105);
nand NAND3 (N4263, N4209, N1750, N186);
xor XOR2 (N4264, N4260, N1705);
nor NOR2 (N4265, N4245, N473);
nand NAND4 (N4266, N4263, N184, N3766, N177);
and AND4 (N4267, N4262, N3881, N754, N3487);
nand NAND3 (N4268, N4251, N2406, N1891);
xor XOR2 (N4269, N4267, N3196);
nand NAND2 (N4270, N4269, N3152);
nor NOR2 (N4271, N4254, N2030);
nor NOR3 (N4272, N4253, N1279, N2304);
not NOT1 (N4273, N4252);
not NOT1 (N4274, N4266);
or OR2 (N4275, N4274, N2982);
xor XOR2 (N4276, N4265, N275);
nor NOR2 (N4277, N4261, N2684);
and AND2 (N4278, N4276, N2174);
not NOT1 (N4279, N4268);
nor NOR3 (N4280, N4272, N2126, N1830);
xor XOR2 (N4281, N4275, N2212);
nor NOR3 (N4282, N4270, N3264, N3135);
nor NOR4 (N4283, N4259, N874, N4182, N2514);
and AND4 (N4284, N4279, N1382, N1920, N4098);
or OR3 (N4285, N4284, N3650, N2333);
nor NOR2 (N4286, N4285, N553);
nand NAND2 (N4287, N4277, N2355);
not NOT1 (N4288, N4282);
xor XOR2 (N4289, N4264, N4067);
xor XOR2 (N4290, N4286, N2493);
not NOT1 (N4291, N4288);
xor XOR2 (N4292, N4287, N1362);
xor XOR2 (N4293, N4289, N1323);
or OR2 (N4294, N4283, N2807);
xor XOR2 (N4295, N4292, N3205);
and AND3 (N4296, N4293, N895, N3889);
nand NAND4 (N4297, N4271, N4094, N4237, N3623);
nor NOR4 (N4298, N4294, N4137, N3263, N3632);
nor NOR4 (N4299, N4291, N1256, N2718, N2628);
and AND2 (N4300, N4295, N4217);
buf BUF1 (N4301, N4300);
nand NAND2 (N4302, N4298, N742);
nor NOR3 (N4303, N4290, N1231, N2464);
nand NAND2 (N4304, N4302, N2144);
nor NOR3 (N4305, N4281, N2243, N2749);
xor XOR2 (N4306, N4273, N3408);
nand NAND3 (N4307, N4304, N18, N3322);
nand NAND2 (N4308, N4303, N2834);
and AND3 (N4309, N4305, N3956, N1956);
or OR4 (N4310, N4309, N3584, N954, N2633);
buf BUF1 (N4311, N4299);
nand NAND2 (N4312, N4278, N83);
or OR3 (N4313, N4306, N2162, N36);
nand NAND2 (N4314, N4312, N1866);
nor NOR2 (N4315, N4310, N3521);
buf BUF1 (N4316, N4313);
or OR4 (N4317, N4308, N1983, N699, N1313);
not NOT1 (N4318, N4317);
and AND4 (N4319, N4296, N1770, N3819, N2776);
nor NOR4 (N4320, N4318, N3192, N57, N207);
or OR2 (N4321, N4315, N3817);
and AND3 (N4322, N4314, N2404, N1392);
and AND4 (N4323, N4321, N1575, N2035, N2105);
not NOT1 (N4324, N4311);
nor NOR3 (N4325, N4323, N2027, N380);
not NOT1 (N4326, N4325);
or OR3 (N4327, N4319, N3060, N3258);
and AND3 (N4328, N4280, N2317, N2212);
nand NAND4 (N4329, N4328, N2657, N226, N3202);
not NOT1 (N4330, N4326);
buf BUF1 (N4331, N4330);
buf BUF1 (N4332, N4301);
xor XOR2 (N4333, N4329, N4279);
and AND4 (N4334, N4331, N247, N680, N240);
buf BUF1 (N4335, N4324);
and AND3 (N4336, N4316, N1878, N2590);
or OR3 (N4337, N4333, N3480, N2118);
nor NOR4 (N4338, N4332, N525, N2346, N1886);
nand NAND2 (N4339, N4322, N2136);
and AND2 (N4340, N4334, N3918);
and AND3 (N4341, N4339, N2673, N2790);
nand NAND4 (N4342, N4338, N912, N3316, N2374);
xor XOR2 (N4343, N4337, N3326);
nand NAND3 (N4344, N4336, N220, N2421);
nor NOR4 (N4345, N4335, N2054, N4018, N2761);
nor NOR3 (N4346, N4342, N295, N2528);
nand NAND4 (N4347, N4343, N730, N1727, N3515);
or OR4 (N4348, N4297, N719, N3789, N1992);
or OR2 (N4349, N4346, N2043);
buf BUF1 (N4350, N4345);
xor XOR2 (N4351, N4347, N3250);
nand NAND4 (N4352, N4327, N3093, N530, N785);
xor XOR2 (N4353, N4344, N473);
xor XOR2 (N4354, N4320, N3729);
and AND2 (N4355, N4351, N282);
or OR4 (N4356, N4354, N4036, N4136, N2693);
not NOT1 (N4357, N4350);
or OR4 (N4358, N4355, N4233, N317, N3489);
or OR3 (N4359, N4357, N145, N440);
xor XOR2 (N4360, N4353, N75);
or OR3 (N4361, N4340, N2310, N1751);
buf BUF1 (N4362, N4349);
not NOT1 (N4363, N4362);
or OR3 (N4364, N4361, N3738, N1080);
nor NOR3 (N4365, N4358, N2728, N3199);
and AND3 (N4366, N4359, N31, N2426);
xor XOR2 (N4367, N4363, N38);
xor XOR2 (N4368, N4365, N1548);
buf BUF1 (N4369, N4366);
not NOT1 (N4370, N4341);
and AND2 (N4371, N4368, N256);
nand NAND2 (N4372, N4356, N467);
and AND2 (N4373, N4370, N2016);
buf BUF1 (N4374, N4364);
xor XOR2 (N4375, N4374, N2040);
and AND2 (N4376, N4373, N2756);
and AND2 (N4377, N4352, N375);
or OR4 (N4378, N4376, N196, N2336, N4289);
and AND2 (N4379, N4307, N3283);
or OR4 (N4380, N4375, N1696, N3828, N4001);
not NOT1 (N4381, N4380);
nand NAND3 (N4382, N4367, N3514, N1636);
not NOT1 (N4383, N4348);
buf BUF1 (N4384, N4360);
not NOT1 (N4385, N4371);
nor NOR2 (N4386, N4379, N40);
and AND2 (N4387, N4372, N2911);
and AND2 (N4388, N4369, N1492);
nor NOR2 (N4389, N4382, N2266);
and AND2 (N4390, N4389, N961);
or OR2 (N4391, N4387, N732);
nor NOR2 (N4392, N4388, N980);
or OR4 (N4393, N4392, N3244, N3302, N2353);
xor XOR2 (N4394, N4377, N3114);
nor NOR4 (N4395, N4386, N178, N1667, N2577);
not NOT1 (N4396, N4383);
nand NAND2 (N4397, N4378, N823);
nor NOR2 (N4398, N4394, N761);
not NOT1 (N4399, N4398);
or OR3 (N4400, N4385, N2212, N760);
or OR4 (N4401, N4393, N2702, N1907, N582);
nor NOR2 (N4402, N4391, N107);
nand NAND2 (N4403, N4381, N8);
xor XOR2 (N4404, N4399, N3324);
or OR2 (N4405, N4402, N3671);
not NOT1 (N4406, N4395);
xor XOR2 (N4407, N4400, N21);
and AND3 (N4408, N4401, N2475, N2908);
nand NAND2 (N4409, N4397, N685);
nor NOR2 (N4410, N4406, N4330);
or OR3 (N4411, N4409, N1522, N2872);
buf BUF1 (N4412, N4403);
or OR2 (N4413, N4408, N3671);
nor NOR2 (N4414, N4413, N878);
xor XOR2 (N4415, N4390, N3382);
and AND4 (N4416, N4412, N3667, N2652, N3048);
not NOT1 (N4417, N4404);
nor NOR2 (N4418, N4411, N3971);
nand NAND3 (N4419, N4414, N625, N823);
nand NAND3 (N4420, N4405, N159, N687);
not NOT1 (N4421, N4384);
or OR4 (N4422, N4421, N2703, N3074, N934);
buf BUF1 (N4423, N4418);
nor NOR4 (N4424, N4410, N2895, N3091, N2063);
and AND3 (N4425, N4396, N2850, N1082);
buf BUF1 (N4426, N4423);
and AND3 (N4427, N4424, N4383, N2493);
buf BUF1 (N4428, N4419);
nor NOR3 (N4429, N4415, N40, N1429);
nor NOR2 (N4430, N4417, N3435);
or OR2 (N4431, N4422, N2079);
xor XOR2 (N4432, N4429, N4357);
nor NOR4 (N4433, N4416, N2118, N3507, N2622);
and AND2 (N4434, N4433, N2803);
nand NAND2 (N4435, N4428, N3276);
xor XOR2 (N4436, N4425, N1846);
buf BUF1 (N4437, N4436);
xor XOR2 (N4438, N4431, N1375);
buf BUF1 (N4439, N4420);
xor XOR2 (N4440, N4434, N2169);
nand NAND4 (N4441, N4439, N890, N279, N2178);
or OR2 (N4442, N4427, N2879);
and AND3 (N4443, N4441, N959, N3919);
not NOT1 (N4444, N4443);
not NOT1 (N4445, N4407);
not NOT1 (N4446, N4426);
xor XOR2 (N4447, N4430, N1773);
not NOT1 (N4448, N4446);
buf BUF1 (N4449, N4432);
or OR2 (N4450, N4440, N3284);
xor XOR2 (N4451, N4435, N2089);
nor NOR3 (N4452, N4444, N332, N787);
and AND2 (N4453, N4445, N3425);
nor NOR3 (N4454, N4453, N451, N1284);
and AND3 (N4455, N4454, N2675, N3998);
nor NOR2 (N4456, N4448, N1086);
xor XOR2 (N4457, N4437, N1871);
nor NOR3 (N4458, N4450, N566, N3542);
nand NAND2 (N4459, N4451, N1037);
and AND4 (N4460, N4459, N1400, N1687, N2093);
buf BUF1 (N4461, N4438);
xor XOR2 (N4462, N4449, N1723);
buf BUF1 (N4463, N4461);
and AND4 (N4464, N4442, N2374, N3368, N545);
xor XOR2 (N4465, N4463, N2336);
nand NAND2 (N4466, N4465, N350);
nor NOR3 (N4467, N4464, N725, N1885);
and AND2 (N4468, N4456, N2826);
and AND2 (N4469, N4457, N3226);
or OR3 (N4470, N4452, N3701, N4006);
or OR2 (N4471, N4468, N2445);
and AND3 (N4472, N4469, N2162, N3739);
nor NOR2 (N4473, N4455, N3786);
nor NOR2 (N4474, N4473, N3698);
nor NOR3 (N4475, N4470, N392, N2326);
buf BUF1 (N4476, N4460);
buf BUF1 (N4477, N4466);
nand NAND4 (N4478, N4447, N4074, N365, N2931);
and AND2 (N4479, N4476, N2411);
nor NOR4 (N4480, N4462, N1231, N2688, N891);
xor XOR2 (N4481, N4467, N443);
xor XOR2 (N4482, N4475, N1462);
nor NOR4 (N4483, N4481, N4419, N4067, N3876);
buf BUF1 (N4484, N4480);
nor NOR2 (N4485, N4472, N2699);
xor XOR2 (N4486, N4485, N3020);
nand NAND2 (N4487, N4483, N458);
and AND2 (N4488, N4478, N659);
or OR2 (N4489, N4484, N2787);
not NOT1 (N4490, N4458);
not NOT1 (N4491, N4489);
or OR4 (N4492, N4479, N811, N4131, N1884);
not NOT1 (N4493, N4490);
buf BUF1 (N4494, N4487);
or OR2 (N4495, N4471, N4277);
and AND2 (N4496, N4488, N3083);
nand NAND3 (N4497, N4495, N1006, N3977);
nor NOR3 (N4498, N4482, N413, N1315);
not NOT1 (N4499, N4494);
nor NOR4 (N4500, N4497, N1431, N1234, N1424);
nand NAND3 (N4501, N4486, N2647, N1496);
buf BUF1 (N4502, N4474);
nor NOR2 (N4503, N4499, N3282);
not NOT1 (N4504, N4501);
or OR3 (N4505, N4500, N1745, N2579);
nor NOR3 (N4506, N4496, N417, N4145);
xor XOR2 (N4507, N4506, N4132);
buf BUF1 (N4508, N4493);
not NOT1 (N4509, N4498);
not NOT1 (N4510, N4505);
buf BUF1 (N4511, N4509);
buf BUF1 (N4512, N4492);
nor NOR3 (N4513, N4477, N3844, N4043);
buf BUF1 (N4514, N4512);
not NOT1 (N4515, N4504);
and AND3 (N4516, N4508, N589, N39);
and AND3 (N4517, N4511, N2104, N1474);
not NOT1 (N4518, N4517);
nand NAND4 (N4519, N4502, N4038, N256, N1204);
nor NOR4 (N4520, N4510, N2535, N2268, N950);
or OR3 (N4521, N4513, N839, N3500);
nand NAND4 (N4522, N4520, N3169, N521, N582);
nand NAND2 (N4523, N4518, N4079);
xor XOR2 (N4524, N4515, N1914);
and AND2 (N4525, N4507, N1690);
buf BUF1 (N4526, N4519);
xor XOR2 (N4527, N4524, N2819);
buf BUF1 (N4528, N4523);
and AND3 (N4529, N4527, N19, N1965);
buf BUF1 (N4530, N4526);
nor NOR3 (N4531, N4521, N3907, N1513);
nor NOR3 (N4532, N4514, N3267, N2333);
nor NOR4 (N4533, N4530, N2429, N512, N2558);
not NOT1 (N4534, N4516);
or OR3 (N4535, N4529, N4300, N2876);
or OR4 (N4536, N4531, N952, N3201, N417);
nand NAND3 (N4537, N4535, N1779, N2338);
nand NAND3 (N4538, N4503, N3241, N2288);
buf BUF1 (N4539, N4534);
and AND2 (N4540, N4533, N2617);
not NOT1 (N4541, N4536);
nand NAND4 (N4542, N4491, N3254, N111, N1301);
buf BUF1 (N4543, N4525);
nor NOR2 (N4544, N4538, N2589);
not NOT1 (N4545, N4537);
and AND4 (N4546, N4528, N4228, N3443, N3465);
nand NAND4 (N4547, N4532, N2813, N398, N3121);
nand NAND3 (N4548, N4546, N770, N2961);
nor NOR4 (N4549, N4545, N3718, N1461, N435);
nand NAND2 (N4550, N4541, N869);
buf BUF1 (N4551, N4549);
xor XOR2 (N4552, N4550, N573);
not NOT1 (N4553, N4539);
and AND2 (N4554, N4551, N1813);
and AND3 (N4555, N4554, N4064, N1443);
xor XOR2 (N4556, N4522, N3448);
nor NOR3 (N4557, N4555, N2611, N4454);
xor XOR2 (N4558, N4552, N2998);
buf BUF1 (N4559, N4543);
nand NAND2 (N4560, N4557, N4089);
not NOT1 (N4561, N4547);
nor NOR4 (N4562, N4540, N555, N3608, N1285);
nand NAND2 (N4563, N4556, N3449);
or OR4 (N4564, N4558, N775, N3480, N3221);
xor XOR2 (N4565, N4564, N1123);
and AND4 (N4566, N4560, N604, N4003, N2164);
not NOT1 (N4567, N4561);
or OR4 (N4568, N4548, N2011, N1162, N2013);
and AND4 (N4569, N4568, N1812, N719, N732);
or OR3 (N4570, N4563, N2849, N3546);
nor NOR2 (N4571, N4562, N1913);
or OR2 (N4572, N4566, N866);
xor XOR2 (N4573, N4565, N540);
and AND2 (N4574, N4571, N1502);
xor XOR2 (N4575, N4559, N3670);
nor NOR4 (N4576, N4553, N2199, N1134, N4183);
nor NOR3 (N4577, N4576, N1305, N480);
nor NOR4 (N4578, N4572, N449, N3006, N2341);
not NOT1 (N4579, N4578);
buf BUF1 (N4580, N4573);
not NOT1 (N4581, N4575);
not NOT1 (N4582, N4542);
and AND4 (N4583, N4574, N3247, N2060, N635);
xor XOR2 (N4584, N4582, N65);
buf BUF1 (N4585, N4570);
xor XOR2 (N4586, N4584, N3175);
and AND2 (N4587, N4581, N1276);
buf BUF1 (N4588, N4585);
xor XOR2 (N4589, N4586, N2174);
not NOT1 (N4590, N4583);
not NOT1 (N4591, N4544);
or OR4 (N4592, N4569, N2531, N780, N1654);
not NOT1 (N4593, N4592);
and AND3 (N4594, N4593, N3584, N1719);
or OR3 (N4595, N4580, N3048, N3487);
not NOT1 (N4596, N4579);
or OR3 (N4597, N4587, N759, N2246);
buf BUF1 (N4598, N4595);
or OR3 (N4599, N4596, N74, N3787);
buf BUF1 (N4600, N4577);
nor NOR3 (N4601, N4598, N2998, N2142);
nor NOR2 (N4602, N4588, N4125);
and AND4 (N4603, N4590, N1465, N3366, N2673);
xor XOR2 (N4604, N4600, N1302);
nand NAND4 (N4605, N4589, N4391, N49, N3168);
and AND2 (N4606, N4604, N2100);
buf BUF1 (N4607, N4591);
nand NAND3 (N4608, N4603, N3185, N3970);
buf BUF1 (N4609, N4567);
buf BUF1 (N4610, N4594);
nor NOR2 (N4611, N4605, N406);
xor XOR2 (N4612, N4610, N4219);
nor NOR3 (N4613, N4611, N768, N3764);
nand NAND2 (N4614, N4607, N3797);
xor XOR2 (N4615, N4609, N4431);
nand NAND2 (N4616, N4615, N3754);
or OR4 (N4617, N4612, N4512, N2922, N4552);
not NOT1 (N4618, N4606);
nand NAND2 (N4619, N4617, N2692);
or OR3 (N4620, N4602, N2290, N1927);
nand NAND2 (N4621, N4620, N3704);
not NOT1 (N4622, N4614);
nand NAND3 (N4623, N4616, N145, N4086);
nand NAND4 (N4624, N4608, N1131, N3201, N4320);
buf BUF1 (N4625, N4601);
xor XOR2 (N4626, N4597, N1153);
not NOT1 (N4627, N4624);
buf BUF1 (N4628, N4599);
and AND4 (N4629, N4625, N3010, N605, N955);
nor NOR4 (N4630, N4618, N2949, N2254, N1938);
or OR2 (N4631, N4622, N3177);
xor XOR2 (N4632, N4626, N1082);
nor NOR2 (N4633, N4630, N1800);
and AND3 (N4634, N4627, N1419, N875);
nand NAND3 (N4635, N4633, N269, N434);
buf BUF1 (N4636, N4629);
xor XOR2 (N4637, N4628, N2059);
nor NOR3 (N4638, N4619, N4362, N1599);
buf BUF1 (N4639, N4631);
xor XOR2 (N4640, N4623, N1117);
xor XOR2 (N4641, N4637, N2977);
or OR3 (N4642, N4635, N1267, N990);
nand NAND4 (N4643, N4613, N1117, N1198, N1076);
not NOT1 (N4644, N4643);
buf BUF1 (N4645, N4639);
nor NOR3 (N4646, N4621, N3335, N2556);
xor XOR2 (N4647, N4642, N2592);
nand NAND3 (N4648, N4644, N2627, N3270);
or OR2 (N4649, N4645, N3122);
not NOT1 (N4650, N4649);
xor XOR2 (N4651, N4636, N912);
or OR2 (N4652, N4638, N4350);
nand NAND3 (N4653, N4641, N1018, N3472);
nand NAND3 (N4654, N4634, N3980, N2706);
buf BUF1 (N4655, N4640);
buf BUF1 (N4656, N4654);
nand NAND2 (N4657, N4651, N4197);
nor NOR3 (N4658, N4656, N4433, N3294);
nor NOR3 (N4659, N4655, N2084, N1611);
and AND2 (N4660, N4658, N3669);
nor NOR3 (N4661, N4632, N2885, N58);
nand NAND2 (N4662, N4652, N3310);
nand NAND2 (N4663, N4646, N2983);
not NOT1 (N4664, N4661);
nand NAND4 (N4665, N4664, N2214, N1293, N1381);
nor NOR4 (N4666, N4662, N2769, N2969, N1039);
or OR3 (N4667, N4648, N1025, N2295);
or OR3 (N4668, N4647, N2360, N1451);
and AND4 (N4669, N4657, N827, N2099, N90);
not NOT1 (N4670, N4665);
not NOT1 (N4671, N4650);
not NOT1 (N4672, N4660);
nand NAND4 (N4673, N4659, N4541, N4160, N4005);
and AND3 (N4674, N4671, N1590, N2635);
nor NOR2 (N4675, N4653, N2076);
and AND2 (N4676, N4668, N337);
nand NAND3 (N4677, N4673, N2300, N4468);
xor XOR2 (N4678, N4676, N820);
nor NOR2 (N4679, N4663, N3732);
buf BUF1 (N4680, N4678);
not NOT1 (N4681, N4675);
buf BUF1 (N4682, N4666);
and AND4 (N4683, N4667, N4264, N2825, N1459);
nor NOR2 (N4684, N4683, N2255);
nand NAND2 (N4685, N4681, N3847);
nand NAND4 (N4686, N4677, N2459, N3274, N462);
nand NAND3 (N4687, N4682, N2280, N3605);
and AND2 (N4688, N4684, N2696);
or OR4 (N4689, N4674, N3671, N1783, N2146);
buf BUF1 (N4690, N4679);
not NOT1 (N4691, N4680);
or OR2 (N4692, N4690, N1155);
xor XOR2 (N4693, N4670, N2866);
not NOT1 (N4694, N4669);
and AND2 (N4695, N4687, N2517);
nor NOR2 (N4696, N4691, N7);
xor XOR2 (N4697, N4685, N1516);
or OR2 (N4698, N4694, N653);
not NOT1 (N4699, N4692);
nor NOR4 (N4700, N4686, N3259, N4321, N2855);
or OR4 (N4701, N4688, N750, N4043, N480);
xor XOR2 (N4702, N4701, N1670);
not NOT1 (N4703, N4697);
nand NAND2 (N4704, N4700, N2200);
nor NOR2 (N4705, N4702, N4491);
buf BUF1 (N4706, N4693);
buf BUF1 (N4707, N4703);
nand NAND3 (N4708, N4706, N2486, N3226);
not NOT1 (N4709, N4699);
nor NOR4 (N4710, N4672, N2713, N2399, N4654);
buf BUF1 (N4711, N4696);
or OR4 (N4712, N4689, N242, N2159, N1257);
xor XOR2 (N4713, N4704, N621);
xor XOR2 (N4714, N4713, N1993);
nand NAND4 (N4715, N4705, N1589, N4151, N1212);
buf BUF1 (N4716, N4711);
or OR3 (N4717, N4715, N1022, N4544);
or OR2 (N4718, N4714, N2931);
nor NOR3 (N4719, N4717, N324, N3381);
nor NOR2 (N4720, N4716, N334);
buf BUF1 (N4721, N4710);
or OR3 (N4722, N4712, N4217, N3905);
buf BUF1 (N4723, N4698);
nand NAND3 (N4724, N4719, N2086, N1092);
not NOT1 (N4725, N4721);
not NOT1 (N4726, N4724);
nand NAND4 (N4727, N4708, N851, N4649, N2369);
xor XOR2 (N4728, N4722, N2721);
nor NOR3 (N4729, N4707, N1486, N3874);
and AND2 (N4730, N4709, N830);
or OR2 (N4731, N4723, N1967);
nand NAND4 (N4732, N4726, N3217, N4602, N4382);
buf BUF1 (N4733, N4732);
or OR2 (N4734, N4727, N3656);
buf BUF1 (N4735, N4718);
nand NAND3 (N4736, N4733, N4563, N318);
nor NOR2 (N4737, N4720, N1580);
xor XOR2 (N4738, N4736, N3702);
xor XOR2 (N4739, N4729, N626);
xor XOR2 (N4740, N4731, N3744);
nor NOR4 (N4741, N4734, N1629, N2700, N1193);
nand NAND3 (N4742, N4735, N3426, N2568);
or OR3 (N4743, N4741, N1064, N976);
buf BUF1 (N4744, N4743);
or OR2 (N4745, N4738, N4037);
buf BUF1 (N4746, N4739);
or OR2 (N4747, N4737, N1680);
nand NAND2 (N4748, N4740, N2872);
nand NAND3 (N4749, N4742, N2295, N1927);
or OR2 (N4750, N4744, N4687);
nor NOR3 (N4751, N4728, N346, N3036);
nor NOR2 (N4752, N4751, N3954);
buf BUF1 (N4753, N4746);
or OR2 (N4754, N4725, N4506);
buf BUF1 (N4755, N4753);
or OR3 (N4756, N4752, N4523, N1863);
nor NOR2 (N4757, N4695, N2344);
nor NOR2 (N4758, N4756, N3682);
and AND3 (N4759, N4730, N4149, N2192);
and AND3 (N4760, N4748, N1891, N3481);
or OR2 (N4761, N4750, N3737);
nor NOR4 (N4762, N4758, N4417, N629, N1797);
and AND4 (N4763, N4760, N3477, N1276, N2568);
not NOT1 (N4764, N4754);
nand NAND4 (N4765, N4764, N1566, N237, N3870);
xor XOR2 (N4766, N4745, N3607);
not NOT1 (N4767, N4766);
xor XOR2 (N4768, N4755, N886);
or OR3 (N4769, N4762, N4038, N4292);
nand NAND3 (N4770, N4761, N161, N1935);
nand NAND2 (N4771, N4768, N2002);
xor XOR2 (N4772, N4769, N85);
and AND4 (N4773, N4765, N4008, N1323, N1543);
and AND3 (N4774, N4770, N1851, N2894);
nand NAND2 (N4775, N4774, N2854);
xor XOR2 (N4776, N4772, N241);
xor XOR2 (N4777, N4757, N1577);
buf BUF1 (N4778, N4759);
or OR2 (N4779, N4747, N4480);
nor NOR3 (N4780, N4776, N1168, N4498);
xor XOR2 (N4781, N4773, N1089);
not NOT1 (N4782, N4771);
not NOT1 (N4783, N4749);
xor XOR2 (N4784, N4767, N1074);
buf BUF1 (N4785, N4781);
nand NAND3 (N4786, N4763, N2861, N2384);
or OR4 (N4787, N4775, N1338, N355, N1912);
nand NAND2 (N4788, N4785, N641);
nand NAND2 (N4789, N4779, N3026);
nand NAND4 (N4790, N4784, N2034, N4131, N2386);
or OR3 (N4791, N4790, N1734, N1130);
buf BUF1 (N4792, N4789);
and AND4 (N4793, N4792, N1642, N849, N3797);
xor XOR2 (N4794, N4777, N1888);
buf BUF1 (N4795, N4786);
and AND4 (N4796, N4782, N1905, N3420, N4530);
nor NOR2 (N4797, N4787, N1746);
xor XOR2 (N4798, N4794, N1177);
or OR3 (N4799, N4778, N2768, N1950);
buf BUF1 (N4800, N4788);
or OR2 (N4801, N4798, N1360);
not NOT1 (N4802, N4800);
not NOT1 (N4803, N4795);
not NOT1 (N4804, N4797);
and AND2 (N4805, N4796, N753);
or OR4 (N4806, N4783, N529, N931, N3359);
not NOT1 (N4807, N4806);
xor XOR2 (N4808, N4807, N3699);
or OR4 (N4809, N4801, N2457, N4121, N4271);
and AND2 (N4810, N4805, N364);
nor NOR4 (N4811, N4810, N4652, N1215, N3505);
buf BUF1 (N4812, N4802);
nor NOR4 (N4813, N4804, N4006, N1774, N3524);
buf BUF1 (N4814, N4812);
nand NAND4 (N4815, N4811, N23, N1053, N496);
nand NAND3 (N4816, N4780, N1739, N1380);
buf BUF1 (N4817, N4814);
and AND3 (N4818, N4817, N2103, N4621);
nand NAND4 (N4819, N4809, N4395, N46, N3558);
and AND4 (N4820, N4818, N1939, N4772, N2128);
not NOT1 (N4821, N4803);
nor NOR2 (N4822, N4820, N29);
buf BUF1 (N4823, N4822);
or OR4 (N4824, N4821, N3055, N4775, N3199);
nor NOR3 (N4825, N4823, N662, N2287);
xor XOR2 (N4826, N4793, N3773);
and AND3 (N4827, N4791, N1806, N3843);
nand NAND2 (N4828, N4816, N2074);
xor XOR2 (N4829, N4826, N1419);
buf BUF1 (N4830, N4819);
or OR2 (N4831, N4825, N3898);
and AND2 (N4832, N4824, N3766);
buf BUF1 (N4833, N4813);
buf BUF1 (N4834, N4827);
and AND2 (N4835, N4833, N1367);
and AND4 (N4836, N4834, N3744, N1294, N1317);
xor XOR2 (N4837, N4829, N1289);
or OR4 (N4838, N4835, N123, N4370, N3549);
nor NOR2 (N4839, N4828, N2977);
buf BUF1 (N4840, N4830);
nand NAND2 (N4841, N4840, N3303);
xor XOR2 (N4842, N4815, N2401);
and AND4 (N4843, N4831, N448, N4336, N1468);
buf BUF1 (N4844, N4837);
and AND4 (N4845, N4836, N1784, N2327, N2345);
xor XOR2 (N4846, N4841, N2256);
or OR3 (N4847, N4843, N3116, N60);
xor XOR2 (N4848, N4844, N181);
nand NAND2 (N4849, N4832, N4085);
xor XOR2 (N4850, N4849, N98);
nand NAND3 (N4851, N4850, N3015, N117);
nand NAND2 (N4852, N4845, N3017);
buf BUF1 (N4853, N4838);
buf BUF1 (N4854, N4851);
and AND2 (N4855, N4847, N1195);
and AND3 (N4856, N4853, N2051, N4721);
nor NOR3 (N4857, N4848, N1943, N2798);
and AND2 (N4858, N4852, N3476);
not NOT1 (N4859, N4856);
xor XOR2 (N4860, N4799, N2603);
nor NOR2 (N4861, N4839, N4084);
xor XOR2 (N4862, N4808, N4617);
nand NAND3 (N4863, N4861, N3397, N1249);
xor XOR2 (N4864, N4855, N1813);
and AND4 (N4865, N4864, N3015, N2084, N2480);
nor NOR4 (N4866, N4842, N2325, N3498, N4492);
not NOT1 (N4867, N4859);
nand NAND3 (N4868, N4858, N1631, N3637);
nor NOR2 (N4869, N4868, N2206);
not NOT1 (N4870, N4846);
and AND3 (N4871, N4870, N501, N3112);
nor NOR4 (N4872, N4857, N2996, N4732, N2015);
nor NOR4 (N4873, N4869, N1713, N1273, N2085);
buf BUF1 (N4874, N4873);
not NOT1 (N4875, N4854);
nor NOR4 (N4876, N4875, N6, N1279, N989);
and AND2 (N4877, N4860, N2319);
and AND4 (N4878, N4865, N2189, N880, N1075);
and AND4 (N4879, N4876, N3576, N958, N2370);
buf BUF1 (N4880, N4872);
and AND2 (N4881, N4862, N3798);
nand NAND3 (N4882, N4877, N468, N4391);
xor XOR2 (N4883, N4878, N4855);
nor NOR2 (N4884, N4866, N134);
not NOT1 (N4885, N4871);
nand NAND2 (N4886, N4879, N4864);
buf BUF1 (N4887, N4881);
and AND2 (N4888, N4887, N2718);
not NOT1 (N4889, N4885);
xor XOR2 (N4890, N4886, N3209);
nand NAND4 (N4891, N4880, N4673, N3619, N2693);
nand NAND2 (N4892, N4884, N2407);
buf BUF1 (N4893, N4888);
not NOT1 (N4894, N4892);
nor NOR3 (N4895, N4890, N1134, N2851);
or OR4 (N4896, N4874, N2243, N2746, N1320);
and AND3 (N4897, N4889, N4763, N4413);
nor NOR2 (N4898, N4883, N1822);
nand NAND4 (N4899, N4882, N2344, N900, N4354);
nor NOR2 (N4900, N4899, N4659);
nor NOR3 (N4901, N4867, N3405, N2960);
nor NOR3 (N4902, N4900, N2816, N2708);
or OR2 (N4903, N4891, N2119);
xor XOR2 (N4904, N4898, N4325);
or OR2 (N4905, N4903, N3177);
xor XOR2 (N4906, N4894, N879);
xor XOR2 (N4907, N4897, N3352);
or OR3 (N4908, N4907, N3102, N93);
nand NAND2 (N4909, N4902, N3039);
nor NOR3 (N4910, N4904, N4157, N2928);
and AND2 (N4911, N4910, N2682);
or OR4 (N4912, N4901, N1353, N2934, N484);
and AND3 (N4913, N4906, N4415, N2665);
buf BUF1 (N4914, N4896);
not NOT1 (N4915, N4863);
nor NOR2 (N4916, N4908, N4813);
or OR3 (N4917, N4911, N4148, N1732);
buf BUF1 (N4918, N4895);
buf BUF1 (N4919, N4912);
and AND4 (N4920, N4919, N4578, N315, N91);
nand NAND2 (N4921, N4920, N2139);
and AND4 (N4922, N4914, N582, N1457, N4921);
or OR2 (N4923, N920, N1899);
not NOT1 (N4924, N4909);
or OR3 (N4925, N4924, N2019, N1140);
or OR4 (N4926, N4913, N4472, N1672, N3228);
and AND2 (N4927, N4905, N3508);
nor NOR4 (N4928, N4918, N4003, N2886, N3406);
xor XOR2 (N4929, N4922, N3593);
nor NOR3 (N4930, N4926, N1128, N4511);
buf BUF1 (N4931, N4930);
xor XOR2 (N4932, N4893, N2066);
nor NOR4 (N4933, N4916, N442, N1476, N538);
or OR4 (N4934, N4915, N1754, N2862, N4439);
nand NAND4 (N4935, N4923, N1460, N737, N1773);
not NOT1 (N4936, N4929);
nand NAND2 (N4937, N4928, N2399);
nand NAND3 (N4938, N4927, N1545, N3999);
not NOT1 (N4939, N4933);
and AND3 (N4940, N4917, N174, N235);
nand NAND4 (N4941, N4938, N134, N2222, N2898);
buf BUF1 (N4942, N4925);
nand NAND3 (N4943, N4932, N3798, N2102);
nor NOR2 (N4944, N4940, N2158);
not NOT1 (N4945, N4937);
or OR4 (N4946, N4939, N1391, N1889, N2066);
nand NAND2 (N4947, N4945, N3963);
buf BUF1 (N4948, N4936);
nor NOR3 (N4949, N4943, N386, N3663);
nor NOR3 (N4950, N4941, N3916, N3406);
nand NAND4 (N4951, N4946, N2282, N3460, N4210);
nor NOR4 (N4952, N4935, N2689, N3872, N1677);
xor XOR2 (N4953, N4949, N1511);
buf BUF1 (N4954, N4931);
nand NAND3 (N4955, N4950, N3738, N2542);
xor XOR2 (N4956, N4947, N2958);
or OR3 (N4957, N4956, N3675, N1693);
and AND4 (N4958, N4957, N2849, N2212, N3230);
or OR4 (N4959, N4944, N4885, N4387, N4800);
or OR4 (N4960, N4948, N2325, N2528, N138);
or OR4 (N4961, N4959, N3816, N3050, N2676);
nor NOR3 (N4962, N4942, N7, N3385);
buf BUF1 (N4963, N4953);
nor NOR2 (N4964, N4952, N3705);
buf BUF1 (N4965, N4962);
nand NAND2 (N4966, N4963, N268);
buf BUF1 (N4967, N4958);
nor NOR2 (N4968, N4955, N200);
not NOT1 (N4969, N4961);
xor XOR2 (N4970, N4965, N349);
not NOT1 (N4971, N4966);
xor XOR2 (N4972, N4934, N3023);
not NOT1 (N4973, N4964);
buf BUF1 (N4974, N4968);
nand NAND3 (N4975, N4973, N2948, N1842);
nor NOR3 (N4976, N4951, N582, N2667);
and AND3 (N4977, N4972, N4647, N1944);
or OR3 (N4978, N4960, N4168, N3490);
nand NAND4 (N4979, N4977, N2155, N3019, N3388);
xor XOR2 (N4980, N4975, N4299);
not NOT1 (N4981, N4976);
nor NOR2 (N4982, N4971, N1722);
buf BUF1 (N4983, N4967);
nor NOR3 (N4984, N4980, N357, N987);
buf BUF1 (N4985, N4954);
nor NOR2 (N4986, N4970, N636);
not NOT1 (N4987, N4979);
and AND4 (N4988, N4984, N997, N4137, N3941);
or OR2 (N4989, N4985, N3585);
and AND3 (N4990, N4969, N2283, N729);
or OR4 (N4991, N4987, N2044, N1723, N4245);
or OR4 (N4992, N4989, N3533, N4609, N2709);
not NOT1 (N4993, N4982);
nor NOR2 (N4994, N4988, N4797);
or OR2 (N4995, N4993, N4021);
xor XOR2 (N4996, N4978, N670);
xor XOR2 (N4997, N4981, N2308);
and AND3 (N4998, N4991, N4752, N4256);
and AND4 (N4999, N4990, N2831, N3755, N3979);
and AND3 (N5000, N4986, N3535, N3144);
not NOT1 (N5001, N4983);
or OR2 (N5002, N4999, N2579);
buf BUF1 (N5003, N4998);
xor XOR2 (N5004, N4997, N826);
and AND4 (N5005, N4996, N2531, N2810, N1127);
or OR3 (N5006, N4995, N2965, N3578);
buf BUF1 (N5007, N5002);
nor NOR3 (N5008, N5001, N142, N50);
or OR4 (N5009, N5008, N2255, N4191, N4720);
nand NAND2 (N5010, N5007, N2460);
nand NAND2 (N5011, N5004, N2597);
xor XOR2 (N5012, N4974, N2678);
buf BUF1 (N5013, N5006);
and AND4 (N5014, N5013, N4904, N4793, N4449);
and AND4 (N5015, N4992, N2404, N3259, N1076);
not NOT1 (N5016, N4994);
nand NAND4 (N5017, N5000, N4808, N4782, N1992);
and AND4 (N5018, N5017, N3704, N622, N3821);
and AND3 (N5019, N5015, N3330, N743);
not NOT1 (N5020, N5016);
or OR2 (N5021, N5009, N1611);
nand NAND2 (N5022, N5020, N3426);
and AND4 (N5023, N5018, N2051, N3711, N4493);
or OR4 (N5024, N5010, N2623, N3015, N1);
xor XOR2 (N5025, N5003, N1866);
buf BUF1 (N5026, N5011);
xor XOR2 (N5027, N5025, N3777);
xor XOR2 (N5028, N5022, N3737);
xor XOR2 (N5029, N5005, N1804);
buf BUF1 (N5030, N5029);
or OR4 (N5031, N5023, N2562, N1349, N2435);
buf BUF1 (N5032, N5030);
buf BUF1 (N5033, N5027);
not NOT1 (N5034, N5032);
nor NOR3 (N5035, N5019, N441, N3923);
xor XOR2 (N5036, N5026, N3661);
nor NOR3 (N5037, N5034, N585, N4590);
xor XOR2 (N5038, N5037, N699);
nand NAND2 (N5039, N5021, N2154);
not NOT1 (N5040, N5036);
not NOT1 (N5041, N5033);
buf BUF1 (N5042, N5035);
buf BUF1 (N5043, N5012);
nand NAND3 (N5044, N5031, N3859, N4439);
or OR4 (N5045, N5039, N3520, N956, N1183);
xor XOR2 (N5046, N5045, N2782);
not NOT1 (N5047, N5040);
and AND3 (N5048, N5046, N4916, N2857);
xor XOR2 (N5049, N5024, N4161);
xor XOR2 (N5050, N5014, N1239);
xor XOR2 (N5051, N5043, N518);
xor XOR2 (N5052, N5048, N537);
xor XOR2 (N5053, N5047, N3863);
xor XOR2 (N5054, N5028, N2753);
or OR4 (N5055, N5042, N4115, N4793, N4399);
not NOT1 (N5056, N5053);
and AND3 (N5057, N5055, N4145, N4843);
or OR3 (N5058, N5038, N4177, N2468);
buf BUF1 (N5059, N5054);
or OR4 (N5060, N5057, N4665, N802, N3128);
nand NAND3 (N5061, N5052, N1468, N4391);
and AND4 (N5062, N5059, N4769, N4799, N751);
or OR4 (N5063, N5044, N1963, N3512, N1522);
or OR3 (N5064, N5056, N860, N1709);
nor NOR4 (N5065, N5050, N220, N3450, N2255);
not NOT1 (N5066, N5060);
nand NAND4 (N5067, N5058, N3373, N3704, N2296);
nand NAND2 (N5068, N5049, N534);
and AND4 (N5069, N5041, N5035, N2361, N3194);
nor NOR3 (N5070, N5064, N1458, N1936);
not NOT1 (N5071, N5069);
and AND4 (N5072, N5051, N2187, N4377, N563);
buf BUF1 (N5073, N5066);
nand NAND4 (N5074, N5073, N4894, N2928, N1015);
nand NAND2 (N5075, N5072, N402);
and AND3 (N5076, N5063, N475, N2359);
and AND4 (N5077, N5070, N1494, N2896, N4964);
and AND2 (N5078, N5062, N2269);
not NOT1 (N5079, N5077);
xor XOR2 (N5080, N5079, N2053);
or OR4 (N5081, N5078, N1571, N4911, N5046);
not NOT1 (N5082, N5080);
nand NAND2 (N5083, N5061, N3522);
nand NAND4 (N5084, N5071, N2750, N1640, N3374);
nor NOR2 (N5085, N5083, N1595);
buf BUF1 (N5086, N5085);
and AND2 (N5087, N5074, N3047);
or OR2 (N5088, N5086, N4439);
xor XOR2 (N5089, N5075, N4439);
buf BUF1 (N5090, N5087);
buf BUF1 (N5091, N5089);
not NOT1 (N5092, N5090);
buf BUF1 (N5093, N5068);
not NOT1 (N5094, N5076);
nor NOR4 (N5095, N5084, N4984, N1489, N476);
not NOT1 (N5096, N5093);
or OR2 (N5097, N5091, N1569);
or OR2 (N5098, N5097, N2634);
and AND4 (N5099, N5065, N2361, N3635, N4086);
nor NOR3 (N5100, N5094, N1746, N1853);
xor XOR2 (N5101, N5100, N1097);
nand NAND3 (N5102, N5067, N742, N2939);
not NOT1 (N5103, N5099);
or OR3 (N5104, N5095, N1610, N222);
nand NAND4 (N5105, N5104, N1506, N2909, N1442);
or OR2 (N5106, N5092, N359);
nor NOR4 (N5107, N5102, N1823, N4200, N128);
nand NAND4 (N5108, N5081, N4606, N4154, N3985);
xor XOR2 (N5109, N5088, N543);
and AND3 (N5110, N5096, N475, N3258);
or OR2 (N5111, N5107, N1017);
or OR4 (N5112, N5101, N1462, N2433, N749);
nor NOR3 (N5113, N5106, N250, N3159);
nor NOR2 (N5114, N5105, N4744);
buf BUF1 (N5115, N5103);
xor XOR2 (N5116, N5115, N2961);
nor NOR4 (N5117, N5112, N921, N503, N2277);
xor XOR2 (N5118, N5098, N193);
not NOT1 (N5119, N5113);
buf BUF1 (N5120, N5111);
xor XOR2 (N5121, N5119, N113);
nand NAND3 (N5122, N5120, N68, N1346);
nand NAND2 (N5123, N5117, N2251);
xor XOR2 (N5124, N5122, N4317);
and AND4 (N5125, N5110, N439, N4807, N1343);
buf BUF1 (N5126, N5082);
not NOT1 (N5127, N5124);
or OR3 (N5128, N5118, N2226, N345);
or OR4 (N5129, N5125, N83, N2988, N1189);
and AND4 (N5130, N5109, N193, N477, N1081);
xor XOR2 (N5131, N5126, N626);
xor XOR2 (N5132, N5121, N438);
buf BUF1 (N5133, N5114);
buf BUF1 (N5134, N5131);
and AND3 (N5135, N5129, N4960, N3363);
not NOT1 (N5136, N5135);
nor NOR4 (N5137, N5116, N3519, N4376, N2018);
and AND3 (N5138, N5132, N581, N4667);
xor XOR2 (N5139, N5108, N4433);
buf BUF1 (N5140, N5139);
xor XOR2 (N5141, N5137, N3713);
buf BUF1 (N5142, N5138);
and AND4 (N5143, N5134, N403, N3374, N75);
and AND4 (N5144, N5130, N3506, N1828, N4416);
and AND2 (N5145, N5140, N1814);
buf BUF1 (N5146, N5142);
not NOT1 (N5147, N5143);
nand NAND2 (N5148, N5144, N3681);
nor NOR4 (N5149, N5127, N1111, N1624, N4973);
buf BUF1 (N5150, N5128);
nand NAND2 (N5151, N5147, N5127);
nand NAND2 (N5152, N5136, N1326);
nor NOR2 (N5153, N5145, N3173);
or OR2 (N5154, N5133, N2168);
nand NAND3 (N5155, N5151, N3487, N4080);
nand NAND3 (N5156, N5123, N3442, N7);
and AND4 (N5157, N5141, N3237, N4121, N4008);
xor XOR2 (N5158, N5146, N1390);
or OR2 (N5159, N5149, N3164);
not NOT1 (N5160, N5154);
or OR3 (N5161, N5155, N1611, N1130);
or OR2 (N5162, N5150, N1516);
nor NOR3 (N5163, N5157, N1875, N1428);
not NOT1 (N5164, N5156);
buf BUF1 (N5165, N5160);
not NOT1 (N5166, N5165);
or OR4 (N5167, N5164, N4339, N2302, N46);
nand NAND4 (N5168, N5153, N4925, N1103, N3290);
xor XOR2 (N5169, N5158, N3779);
buf BUF1 (N5170, N5163);
xor XOR2 (N5171, N5167, N3802);
not NOT1 (N5172, N5148);
not NOT1 (N5173, N5166);
nand NAND3 (N5174, N5162, N2257, N2124);
not NOT1 (N5175, N5168);
or OR4 (N5176, N5169, N3240, N3361, N2303);
or OR3 (N5177, N5161, N705, N3250);
xor XOR2 (N5178, N5176, N2371);
not NOT1 (N5179, N5177);
or OR3 (N5180, N5172, N4073, N982);
nor NOR4 (N5181, N5179, N668, N332, N3337);
or OR4 (N5182, N5178, N1957, N1634, N3906);
not NOT1 (N5183, N5159);
buf BUF1 (N5184, N5175);
nand NAND4 (N5185, N5181, N2959, N1039, N1428);
nor NOR3 (N5186, N5173, N4677, N2889);
and AND4 (N5187, N5183, N4029, N2462, N1101);
buf BUF1 (N5188, N5186);
nand NAND4 (N5189, N5185, N108, N3633, N2895);
nand NAND3 (N5190, N5171, N1263, N4149);
not NOT1 (N5191, N5182);
xor XOR2 (N5192, N5180, N261);
not NOT1 (N5193, N5188);
nand NAND4 (N5194, N5193, N1331, N4048, N4095);
and AND4 (N5195, N5192, N188, N1891, N2780);
nand NAND4 (N5196, N5152, N206, N1837, N193);
xor XOR2 (N5197, N5196, N4109);
nor NOR4 (N5198, N5191, N1492, N4943, N1167);
xor XOR2 (N5199, N5197, N2059);
xor XOR2 (N5200, N5189, N3354);
or OR3 (N5201, N5187, N3788, N1012);
and AND4 (N5202, N5170, N656, N595, N4689);
buf BUF1 (N5203, N5195);
not NOT1 (N5204, N5199);
xor XOR2 (N5205, N5174, N2611);
or OR2 (N5206, N5200, N598);
xor XOR2 (N5207, N5206, N3626);
buf BUF1 (N5208, N5207);
nand NAND2 (N5209, N5203, N3760);
xor XOR2 (N5210, N5205, N3274);
nor NOR3 (N5211, N5190, N2862, N1267);
and AND2 (N5212, N5198, N4516);
and AND4 (N5213, N5212, N1444, N1713, N3442);
xor XOR2 (N5214, N5204, N4990);
xor XOR2 (N5215, N5210, N2941);
nand NAND4 (N5216, N5209, N2933, N326, N413);
xor XOR2 (N5217, N5214, N1111);
nand NAND4 (N5218, N5208, N3639, N2841, N673);
nand NAND4 (N5219, N5217, N1205, N5027, N2318);
and AND3 (N5220, N5211, N2309, N4362);
not NOT1 (N5221, N5213);
and AND2 (N5222, N5215, N527);
not NOT1 (N5223, N5221);
nand NAND4 (N5224, N5201, N1444, N1171, N2247);
buf BUF1 (N5225, N5219);
buf BUF1 (N5226, N5216);
or OR2 (N5227, N5224, N2833);
buf BUF1 (N5228, N5226);
and AND2 (N5229, N5194, N3591);
nor NOR4 (N5230, N5227, N2099, N2314, N204);
buf BUF1 (N5231, N5228);
nor NOR4 (N5232, N5223, N311, N5045, N3771);
nor NOR2 (N5233, N5225, N4383);
nor NOR2 (N5234, N5218, N2232);
xor XOR2 (N5235, N5231, N3710);
nand NAND3 (N5236, N5229, N4222, N1449);
nand NAND4 (N5237, N5236, N1697, N2319, N125);
nand NAND3 (N5238, N5220, N2614, N1198);
and AND2 (N5239, N5237, N237);
xor XOR2 (N5240, N5202, N597);
xor XOR2 (N5241, N5240, N4057);
nor NOR3 (N5242, N5230, N3978, N5096);
buf BUF1 (N5243, N5241);
not NOT1 (N5244, N5233);
and AND4 (N5245, N5239, N4911, N2172, N2305);
and AND2 (N5246, N5184, N3263);
nor NOR3 (N5247, N5242, N156, N3820);
and AND3 (N5248, N5232, N3934, N3601);
buf BUF1 (N5249, N5247);
nor NOR3 (N5250, N5249, N810, N3951);
nor NOR4 (N5251, N5222, N5205, N5121, N4661);
nand NAND2 (N5252, N5245, N2205);
or OR4 (N5253, N5235, N2047, N4644, N292);
xor XOR2 (N5254, N5243, N2635);
nand NAND2 (N5255, N5254, N2022);
or OR2 (N5256, N5238, N2732);
and AND3 (N5257, N5253, N4647, N2774);
xor XOR2 (N5258, N5234, N5079);
xor XOR2 (N5259, N5244, N1509);
nor NOR4 (N5260, N5251, N3493, N1042, N3038);
xor XOR2 (N5261, N5260, N1301);
or OR4 (N5262, N5250, N3948, N744, N1676);
xor XOR2 (N5263, N5255, N3078);
buf BUF1 (N5264, N5248);
nand NAND4 (N5265, N5258, N1903, N948, N462);
nand NAND4 (N5266, N5259, N4436, N527, N3911);
or OR4 (N5267, N5264, N492, N2071, N2877);
nand NAND4 (N5268, N5246, N395, N4520, N2114);
nor NOR4 (N5269, N5266, N4019, N1144, N3200);
xor XOR2 (N5270, N5269, N1858);
buf BUF1 (N5271, N5263);
buf BUF1 (N5272, N5252);
nor NOR3 (N5273, N5256, N2870, N417);
buf BUF1 (N5274, N5271);
xor XOR2 (N5275, N5262, N452);
not NOT1 (N5276, N5275);
and AND2 (N5277, N5257, N1184);
not NOT1 (N5278, N5273);
nor NOR2 (N5279, N5277, N903);
nand NAND2 (N5280, N5270, N3472);
not NOT1 (N5281, N5265);
buf BUF1 (N5282, N5278);
buf BUF1 (N5283, N5280);
xor XOR2 (N5284, N5281, N1945);
not NOT1 (N5285, N5267);
nor NOR3 (N5286, N5261, N4781, N2147);
or OR3 (N5287, N5279, N2573, N1910);
or OR2 (N5288, N5282, N4038);
xor XOR2 (N5289, N5274, N1389);
and AND4 (N5290, N5288, N1860, N2016, N1559);
not NOT1 (N5291, N5272);
nand NAND3 (N5292, N5284, N4563, N3832);
xor XOR2 (N5293, N5287, N3751);
nand NAND4 (N5294, N5285, N3568, N2778, N1865);
buf BUF1 (N5295, N5276);
xor XOR2 (N5296, N5293, N5119);
nand NAND2 (N5297, N5289, N4418);
and AND4 (N5298, N5283, N724, N237, N4966);
nand NAND3 (N5299, N5298, N3471, N2223);
not NOT1 (N5300, N5292);
not NOT1 (N5301, N5290);
or OR3 (N5302, N5297, N2487, N3065);
xor XOR2 (N5303, N5302, N1599);
buf BUF1 (N5304, N5303);
buf BUF1 (N5305, N5299);
not NOT1 (N5306, N5304);
xor XOR2 (N5307, N5295, N4484);
or OR3 (N5308, N5307, N4387, N1824);
and AND4 (N5309, N5294, N3783, N4142, N4273);
not NOT1 (N5310, N5309);
or OR2 (N5311, N5300, N1700);
buf BUF1 (N5312, N5268);
not NOT1 (N5313, N5312);
nand NAND3 (N5314, N5311, N3196, N3591);
and AND4 (N5315, N5306, N1491, N485, N4559);
or OR4 (N5316, N5286, N2809, N2542, N1825);
nor NOR2 (N5317, N5291, N809);
not NOT1 (N5318, N5314);
nor NOR4 (N5319, N5317, N2578, N1284, N1353);
nor NOR4 (N5320, N5319, N679, N3066, N704);
buf BUF1 (N5321, N5308);
nand NAND4 (N5322, N5301, N3654, N2847, N2248);
xor XOR2 (N5323, N5316, N1693);
or OR3 (N5324, N5321, N4096, N4377);
xor XOR2 (N5325, N5310, N4923);
nor NOR3 (N5326, N5313, N1636, N3160);
xor XOR2 (N5327, N5315, N4809);
or OR4 (N5328, N5322, N3987, N377, N1263);
not NOT1 (N5329, N5325);
xor XOR2 (N5330, N5327, N4186);
nor NOR2 (N5331, N5318, N772);
or OR3 (N5332, N5305, N1917, N186);
nand NAND3 (N5333, N5332, N4105, N2587);
buf BUF1 (N5334, N5296);
not NOT1 (N5335, N5330);
xor XOR2 (N5336, N5324, N737);
nor NOR3 (N5337, N5335, N3547, N18);
nor NOR3 (N5338, N5328, N1249, N2455);
buf BUF1 (N5339, N5323);
xor XOR2 (N5340, N5337, N3284);
or OR2 (N5341, N5326, N3695);
nand NAND2 (N5342, N5334, N58);
nor NOR4 (N5343, N5339, N4652, N3181, N4011);
or OR4 (N5344, N5342, N1190, N941, N2350);
nand NAND2 (N5345, N5338, N988);
and AND3 (N5346, N5343, N3088, N2032);
not NOT1 (N5347, N5345);
and AND2 (N5348, N5347, N1161);
xor XOR2 (N5349, N5329, N2735);
and AND4 (N5350, N5333, N964, N311, N2364);
and AND4 (N5351, N5340, N2275, N5215, N959);
or OR2 (N5352, N5346, N3854);
or OR2 (N5353, N5331, N5227);
nor NOR2 (N5354, N5353, N1491);
and AND4 (N5355, N5336, N1890, N387, N3818);
nand NAND3 (N5356, N5341, N3242, N2648);
xor XOR2 (N5357, N5350, N4558);
or OR3 (N5358, N5351, N2934, N1786);
nor NOR2 (N5359, N5357, N1788);
nor NOR3 (N5360, N5356, N4315, N1103);
xor XOR2 (N5361, N5320, N2293);
buf BUF1 (N5362, N5344);
nor NOR3 (N5363, N5362, N199, N485);
xor XOR2 (N5364, N5354, N4394);
and AND2 (N5365, N5359, N1897);
xor XOR2 (N5366, N5355, N583);
not NOT1 (N5367, N5358);
not NOT1 (N5368, N5363);
and AND4 (N5369, N5367, N5355, N4293, N2011);
nand NAND4 (N5370, N5361, N1536, N1611, N3963);
not NOT1 (N5371, N5364);
nand NAND3 (N5372, N5352, N5255, N2598);
nor NOR2 (N5373, N5372, N681);
and AND2 (N5374, N5360, N1094);
not NOT1 (N5375, N5371);
buf BUF1 (N5376, N5370);
and AND3 (N5377, N5369, N4398, N3829);
or OR4 (N5378, N5373, N1737, N1043, N3580);
not NOT1 (N5379, N5374);
not NOT1 (N5380, N5368);
and AND4 (N5381, N5376, N4091, N3900, N2220);
nor NOR2 (N5382, N5375, N2156);
not NOT1 (N5383, N5380);
buf BUF1 (N5384, N5378);
nand NAND4 (N5385, N5384, N397, N2835, N2536);
or OR4 (N5386, N5385, N3032, N4877, N1460);
buf BUF1 (N5387, N5348);
or OR2 (N5388, N5381, N2869);
buf BUF1 (N5389, N5388);
and AND4 (N5390, N5386, N3785, N133, N399);
and AND3 (N5391, N5365, N4006, N3608);
not NOT1 (N5392, N5377);
and AND3 (N5393, N5390, N3796, N3292);
or OR4 (N5394, N5349, N100, N4483, N5329);
xor XOR2 (N5395, N5393, N1756);
not NOT1 (N5396, N5387);
nand NAND2 (N5397, N5382, N1645);
or OR2 (N5398, N5389, N5381);
and AND4 (N5399, N5398, N1188, N1301, N644);
nand NAND2 (N5400, N5383, N3257);
xor XOR2 (N5401, N5366, N3589);
nand NAND3 (N5402, N5401, N1181, N5054);
not NOT1 (N5403, N5402);
and AND4 (N5404, N5400, N596, N1975, N4406);
buf BUF1 (N5405, N5399);
and AND2 (N5406, N5392, N918);
or OR3 (N5407, N5404, N1069, N5368);
nor NOR4 (N5408, N5391, N5378, N1240, N1821);
nor NOR2 (N5409, N5394, N810);
nand NAND2 (N5410, N5407, N1005);
xor XOR2 (N5411, N5408, N1576);
nor NOR3 (N5412, N5397, N4874, N4038);
or OR3 (N5413, N5396, N2340, N2341);
not NOT1 (N5414, N5413);
xor XOR2 (N5415, N5406, N1093);
nor NOR4 (N5416, N5412, N4210, N3174, N5311);
buf BUF1 (N5417, N5409);
not NOT1 (N5418, N5416);
not NOT1 (N5419, N5379);
nor NOR2 (N5420, N5410, N1911);
xor XOR2 (N5421, N5420, N576);
not NOT1 (N5422, N5405);
buf BUF1 (N5423, N5403);
or OR2 (N5424, N5411, N455);
not NOT1 (N5425, N5423);
nand NAND3 (N5426, N5425, N2334, N2139);
buf BUF1 (N5427, N5414);
nand NAND3 (N5428, N5417, N855, N3163);
nand NAND4 (N5429, N5395, N2410, N4160, N215);
or OR3 (N5430, N5422, N4453, N4745);
nand NAND2 (N5431, N5419, N2092);
not NOT1 (N5432, N5415);
nand NAND2 (N5433, N5424, N5001);
and AND3 (N5434, N5433, N1261, N899);
and AND3 (N5435, N5428, N4058, N3650);
or OR3 (N5436, N5431, N335, N3501);
not NOT1 (N5437, N5418);
nor NOR3 (N5438, N5430, N1417, N3266);
xor XOR2 (N5439, N5427, N1144);
and AND2 (N5440, N5435, N3428);
and AND2 (N5441, N5426, N676);
or OR4 (N5442, N5439, N1570, N2424, N1560);
nor NOR4 (N5443, N5441, N1536, N820, N2551);
nand NAND4 (N5444, N5443, N3597, N3006, N3816);
or OR3 (N5445, N5440, N990, N3276);
not NOT1 (N5446, N5429);
or OR3 (N5447, N5442, N1786, N3611);
and AND2 (N5448, N5445, N356);
and AND3 (N5449, N5447, N3145, N1704);
buf BUF1 (N5450, N5434);
nand NAND4 (N5451, N5448, N4360, N301, N3973);
or OR2 (N5452, N5446, N2949);
xor XOR2 (N5453, N5452, N3468);
nand NAND3 (N5454, N5436, N4544, N2879);
not NOT1 (N5455, N5444);
and AND3 (N5456, N5438, N1410, N3330);
nand NAND2 (N5457, N5454, N1572);
and AND2 (N5458, N5455, N5417);
not NOT1 (N5459, N5451);
nand NAND3 (N5460, N5432, N4170, N2047);
not NOT1 (N5461, N5450);
nor NOR3 (N5462, N5453, N2147, N903);
and AND2 (N5463, N5459, N4703);
nor NOR4 (N5464, N5437, N4032, N2375, N3575);
nand NAND4 (N5465, N5461, N867, N5369, N347);
and AND3 (N5466, N5464, N4079, N4110);
and AND2 (N5467, N5462, N3107);
nor NOR2 (N5468, N5467, N5214);
or OR4 (N5469, N5468, N637, N1075, N3650);
buf BUF1 (N5470, N5449);
nor NOR2 (N5471, N5458, N5448);
xor XOR2 (N5472, N5465, N3960);
nor NOR2 (N5473, N5463, N2145);
not NOT1 (N5474, N5473);
or OR4 (N5475, N5469, N4015, N1000, N3778);
nor NOR4 (N5476, N5475, N4616, N4997, N799);
or OR2 (N5477, N5456, N3937);
nor NOR3 (N5478, N5471, N3015, N1330);
buf BUF1 (N5479, N5472);
and AND3 (N5480, N5460, N3647, N1340);
xor XOR2 (N5481, N5470, N3980);
or OR2 (N5482, N5457, N5318);
xor XOR2 (N5483, N5481, N523);
and AND2 (N5484, N5474, N376);
or OR3 (N5485, N5478, N54, N3023);
and AND2 (N5486, N5466, N3919);
and AND3 (N5487, N5476, N4735, N5106);
not NOT1 (N5488, N5487);
nand NAND2 (N5489, N5477, N4036);
and AND2 (N5490, N5483, N1792);
and AND4 (N5491, N5484, N3809, N3676, N1351);
or OR4 (N5492, N5482, N2896, N3147, N3118);
nor NOR3 (N5493, N5490, N3002, N2768);
nand NAND4 (N5494, N5492, N3637, N3966, N2536);
nor NOR2 (N5495, N5489, N5349);
not NOT1 (N5496, N5491);
not NOT1 (N5497, N5486);
xor XOR2 (N5498, N5494, N2585);
buf BUF1 (N5499, N5498);
buf BUF1 (N5500, N5493);
not NOT1 (N5501, N5485);
buf BUF1 (N5502, N5497);
nor NOR4 (N5503, N5495, N5482, N1214, N2238);
nand NAND2 (N5504, N5480, N5053);
nor NOR3 (N5505, N5503, N4912, N210);
nor NOR2 (N5506, N5479, N550);
or OR3 (N5507, N5502, N2112, N2127);
and AND2 (N5508, N5507, N154);
nor NOR4 (N5509, N5508, N3270, N2623, N3162);
buf BUF1 (N5510, N5499);
or OR3 (N5511, N5506, N612, N438);
buf BUF1 (N5512, N5504);
and AND4 (N5513, N5509, N4127, N3111, N931);
not NOT1 (N5514, N5513);
or OR3 (N5515, N5511, N5449, N3934);
or OR2 (N5516, N5514, N1929);
nor NOR2 (N5517, N5512, N1111);
xor XOR2 (N5518, N5488, N908);
nor NOR3 (N5519, N5516, N273, N4988);
nand NAND3 (N5520, N5518, N4520, N944);
and AND2 (N5521, N5519, N3660);
nor NOR3 (N5522, N5521, N2615, N1012);
nand NAND2 (N5523, N5496, N5021);
nand NAND3 (N5524, N5510, N5011, N4172);
nor NOR4 (N5525, N5500, N3211, N4974, N4154);
nand NAND2 (N5526, N5524, N4479);
not NOT1 (N5527, N5505);
buf BUF1 (N5528, N5527);
xor XOR2 (N5529, N5520, N1882);
not NOT1 (N5530, N5501);
nor NOR3 (N5531, N5528, N5184, N4055);
and AND4 (N5532, N5522, N684, N5066, N4605);
not NOT1 (N5533, N5530);
xor XOR2 (N5534, N5529, N384);
nor NOR3 (N5535, N5523, N4724, N4784);
and AND4 (N5536, N5533, N2228, N1734, N3590);
xor XOR2 (N5537, N5526, N5031);
nor NOR3 (N5538, N5535, N4542, N593);
xor XOR2 (N5539, N5536, N1536);
xor XOR2 (N5540, N5532, N2120);
and AND4 (N5541, N5540, N2178, N2761, N430);
xor XOR2 (N5542, N5537, N1653);
or OR2 (N5543, N5539, N4471);
buf BUF1 (N5544, N5525);
buf BUF1 (N5545, N5515);
or OR3 (N5546, N5534, N2551, N5004);
not NOT1 (N5547, N5545);
and AND4 (N5548, N5543, N3349, N3214, N2431);
nand NAND4 (N5549, N5546, N541, N5180, N238);
xor XOR2 (N5550, N5542, N5269);
xor XOR2 (N5551, N5547, N4012);
buf BUF1 (N5552, N5531);
or OR2 (N5553, N5551, N5346);
not NOT1 (N5554, N5538);
nand NAND2 (N5555, N5421, N3571);
and AND3 (N5556, N5544, N5263, N2173);
and AND4 (N5557, N5548, N4969, N109, N2763);
nand NAND2 (N5558, N5550, N5300);
nand NAND3 (N5559, N5555, N523, N3918);
buf BUF1 (N5560, N5553);
and AND2 (N5561, N5560, N4003);
xor XOR2 (N5562, N5559, N5395);
buf BUF1 (N5563, N5552);
nand NAND3 (N5564, N5556, N679, N4086);
nor NOR2 (N5565, N5557, N5265);
not NOT1 (N5566, N5541);
nand NAND2 (N5567, N5565, N4821);
nor NOR3 (N5568, N5561, N4573, N4071);
buf BUF1 (N5569, N5566);
nand NAND2 (N5570, N5549, N3657);
nand NAND4 (N5571, N5554, N238, N508, N377);
xor XOR2 (N5572, N5568, N3247);
nor NOR2 (N5573, N5563, N593);
and AND4 (N5574, N5570, N1451, N1777, N5360);
nand NAND2 (N5575, N5572, N5122);
xor XOR2 (N5576, N5569, N2672);
buf BUF1 (N5577, N5575);
nand NAND2 (N5578, N5576, N1146);
nand NAND2 (N5579, N5574, N2158);
and AND2 (N5580, N5562, N966);
and AND4 (N5581, N5573, N480, N2925, N4706);
and AND4 (N5582, N5558, N3678, N487, N123);
and AND4 (N5583, N5579, N5043, N4640, N721);
or OR2 (N5584, N5571, N627);
nand NAND2 (N5585, N5578, N1591);
not NOT1 (N5586, N5580);
nor NOR4 (N5587, N5585, N2175, N4622, N4154);
not NOT1 (N5588, N5586);
not NOT1 (N5589, N5584);
or OR3 (N5590, N5567, N1848, N4056);
buf BUF1 (N5591, N5589);
and AND2 (N5592, N5581, N4030);
buf BUF1 (N5593, N5517);
or OR4 (N5594, N5590, N635, N4887, N1601);
or OR4 (N5595, N5583, N129, N228, N3297);
buf BUF1 (N5596, N5592);
nand NAND4 (N5597, N5593, N2769, N2671, N1900);
or OR3 (N5598, N5596, N4417, N82);
buf BUF1 (N5599, N5595);
or OR3 (N5600, N5591, N4476, N533);
nand NAND3 (N5601, N5599, N1777, N1664);
not NOT1 (N5602, N5588);
buf BUF1 (N5603, N5598);
and AND4 (N5604, N5564, N3127, N1220, N2688);
not NOT1 (N5605, N5577);
xor XOR2 (N5606, N5594, N2645);
xor XOR2 (N5607, N5606, N1883);
nor NOR3 (N5608, N5607, N4511, N1336);
nand NAND3 (N5609, N5582, N739, N3234);
xor XOR2 (N5610, N5603, N1163);
and AND3 (N5611, N5609, N3441, N1695);
or OR3 (N5612, N5605, N901, N2538);
buf BUF1 (N5613, N5602);
or OR4 (N5614, N5613, N3093, N4308, N4248);
or OR3 (N5615, N5614, N5416, N220);
nor NOR3 (N5616, N5611, N3140, N1694);
xor XOR2 (N5617, N5608, N4593);
and AND3 (N5618, N5587, N5064, N2567);
and AND4 (N5619, N5615, N1630, N1305, N1360);
not NOT1 (N5620, N5616);
buf BUF1 (N5621, N5601);
or OR3 (N5622, N5618, N5175, N2959);
not NOT1 (N5623, N5622);
xor XOR2 (N5624, N5623, N592);
and AND3 (N5625, N5617, N835, N583);
nand NAND3 (N5626, N5621, N4232, N964);
or OR2 (N5627, N5620, N1294);
nand NAND2 (N5628, N5619, N623);
and AND4 (N5629, N5612, N2724, N5183, N4937);
and AND4 (N5630, N5597, N5220, N4514, N4143);
nand NAND4 (N5631, N5610, N1662, N2483, N2738);
buf BUF1 (N5632, N5628);
nand NAND4 (N5633, N5604, N1326, N2775, N3583);
nand NAND2 (N5634, N5631, N2049);
nor NOR4 (N5635, N5633, N4434, N294, N1856);
or OR3 (N5636, N5629, N2257, N980);
nor NOR3 (N5637, N5626, N2744, N5508);
nand NAND4 (N5638, N5627, N3482, N2709, N5379);
xor XOR2 (N5639, N5634, N305);
xor XOR2 (N5640, N5637, N3573);
xor XOR2 (N5641, N5639, N1507);
nand NAND2 (N5642, N5624, N3032);
nor NOR2 (N5643, N5630, N3056);
buf BUF1 (N5644, N5638);
buf BUF1 (N5645, N5640);
buf BUF1 (N5646, N5642);
and AND4 (N5647, N5646, N536, N5504, N5158);
buf BUF1 (N5648, N5641);
xor XOR2 (N5649, N5636, N4994);
nand NAND2 (N5650, N5600, N3757);
nand NAND3 (N5651, N5649, N3145, N3309);
not NOT1 (N5652, N5632);
or OR3 (N5653, N5650, N3118, N2633);
nor NOR2 (N5654, N5643, N1205);
not NOT1 (N5655, N5652);
and AND4 (N5656, N5648, N785, N1692, N5273);
not NOT1 (N5657, N5653);
and AND3 (N5658, N5647, N986, N1313);
xor XOR2 (N5659, N5635, N2532);
not NOT1 (N5660, N5625);
and AND4 (N5661, N5660, N1205, N4810, N2200);
and AND4 (N5662, N5654, N4808, N1387, N1656);
xor XOR2 (N5663, N5656, N3179);
xor XOR2 (N5664, N5663, N5404);
xor XOR2 (N5665, N5655, N139);
not NOT1 (N5666, N5664);
or OR3 (N5667, N5659, N4163, N2709);
buf BUF1 (N5668, N5667);
xor XOR2 (N5669, N5644, N3887);
and AND4 (N5670, N5645, N1050, N172, N5305);
buf BUF1 (N5671, N5651);
nand NAND3 (N5672, N5665, N4998, N1672);
nor NOR3 (N5673, N5666, N1199, N3667);
or OR4 (N5674, N5669, N2530, N2711, N3304);
or OR4 (N5675, N5658, N177, N554, N2167);
or OR3 (N5676, N5672, N3054, N354);
xor XOR2 (N5677, N5671, N2650);
buf BUF1 (N5678, N5673);
nor NOR3 (N5679, N5662, N3910, N1726);
not NOT1 (N5680, N5679);
buf BUF1 (N5681, N5676);
nand NAND2 (N5682, N5677, N3996);
buf BUF1 (N5683, N5657);
nor NOR2 (N5684, N5670, N4549);
and AND3 (N5685, N5681, N2890, N5139);
nor NOR2 (N5686, N5680, N5271);
nand NAND3 (N5687, N5661, N2549, N3866);
nand NAND3 (N5688, N5686, N1427, N599);
xor XOR2 (N5689, N5688, N1721);
nand NAND4 (N5690, N5682, N4497, N4183, N25);
or OR2 (N5691, N5668, N832);
or OR3 (N5692, N5687, N3721, N4726);
nor NOR2 (N5693, N5685, N1689);
nand NAND3 (N5694, N5693, N2539, N5318);
nor NOR2 (N5695, N5694, N2936);
buf BUF1 (N5696, N5692);
nand NAND2 (N5697, N5696, N4126);
and AND4 (N5698, N5683, N2726, N5026, N2348);
xor XOR2 (N5699, N5691, N471);
nor NOR2 (N5700, N5675, N3091);
buf BUF1 (N5701, N5697);
nor NOR3 (N5702, N5684, N5342, N2288);
not NOT1 (N5703, N5689);
nand NAND4 (N5704, N5703, N2081, N4157, N411);
xor XOR2 (N5705, N5699, N1009);
xor XOR2 (N5706, N5674, N2688);
not NOT1 (N5707, N5695);
buf BUF1 (N5708, N5690);
nand NAND4 (N5709, N5706, N2514, N3304, N508);
nand NAND3 (N5710, N5678, N2812, N3200);
xor XOR2 (N5711, N5710, N2717);
or OR2 (N5712, N5711, N5245);
and AND4 (N5713, N5702, N5171, N3412, N2546);
or OR4 (N5714, N5713, N4803, N1260, N5432);
or OR2 (N5715, N5709, N2892);
xor XOR2 (N5716, N5707, N3240);
xor XOR2 (N5717, N5705, N3699);
nor NOR3 (N5718, N5700, N1216, N5432);
nand NAND3 (N5719, N5714, N64, N567);
or OR4 (N5720, N5716, N3708, N3878, N2329);
buf BUF1 (N5721, N5704);
xor XOR2 (N5722, N5717, N4319);
buf BUF1 (N5723, N5708);
and AND4 (N5724, N5712, N5464, N938, N4291);
buf BUF1 (N5725, N5720);
not NOT1 (N5726, N5698);
or OR4 (N5727, N5725, N2449, N1690, N3912);
and AND4 (N5728, N5723, N2120, N2205, N3901);
not NOT1 (N5729, N5718);
xor XOR2 (N5730, N5728, N1480);
buf BUF1 (N5731, N5726);
nor NOR2 (N5732, N5730, N2062);
nor NOR4 (N5733, N5727, N2023, N1064, N3574);
nor NOR4 (N5734, N5731, N3130, N1087, N2810);
xor XOR2 (N5735, N5724, N142);
and AND2 (N5736, N5719, N3605);
or OR3 (N5737, N5736, N1718, N4907);
not NOT1 (N5738, N5733);
not NOT1 (N5739, N5722);
buf BUF1 (N5740, N5735);
buf BUF1 (N5741, N5701);
or OR3 (N5742, N5739, N288, N215);
xor XOR2 (N5743, N5732, N2286);
nor NOR4 (N5744, N5741, N4075, N1436, N1553);
or OR4 (N5745, N5729, N4179, N5558, N272);
not NOT1 (N5746, N5742);
or OR4 (N5747, N5740, N3599, N4699, N3816);
not NOT1 (N5748, N5747);
or OR3 (N5749, N5715, N3808, N368);
buf BUF1 (N5750, N5737);
nand NAND3 (N5751, N5721, N779, N451);
xor XOR2 (N5752, N5748, N1323);
buf BUF1 (N5753, N5746);
or OR2 (N5754, N5750, N4713);
or OR4 (N5755, N5743, N4439, N2242, N2246);
buf BUF1 (N5756, N5752);
buf BUF1 (N5757, N5749);
xor XOR2 (N5758, N5754, N4646);
xor XOR2 (N5759, N5751, N3614);
xor XOR2 (N5760, N5745, N5473);
buf BUF1 (N5761, N5757);
or OR3 (N5762, N5755, N887, N1675);
buf BUF1 (N5763, N5744);
or OR2 (N5764, N5763, N5671);
xor XOR2 (N5765, N5760, N5219);
xor XOR2 (N5766, N5758, N867);
nor NOR2 (N5767, N5766, N1946);
or OR4 (N5768, N5761, N3383, N1987, N5592);
not NOT1 (N5769, N5764);
or OR4 (N5770, N5756, N4762, N1461, N5076);
xor XOR2 (N5771, N5759, N1476);
or OR2 (N5772, N5771, N257);
buf BUF1 (N5773, N5768);
or OR4 (N5774, N5773, N4935, N2779, N3209);
xor XOR2 (N5775, N5765, N5460);
or OR2 (N5776, N5734, N4804);
nand NAND2 (N5777, N5776, N3201);
xor XOR2 (N5778, N5753, N117);
nor NOR4 (N5779, N5770, N591, N4562, N4188);
xor XOR2 (N5780, N5777, N2002);
nor NOR3 (N5781, N5767, N4681, N1173);
xor XOR2 (N5782, N5778, N4608);
not NOT1 (N5783, N5769);
nand NAND3 (N5784, N5781, N4111, N1894);
and AND2 (N5785, N5774, N3815);
not NOT1 (N5786, N5780);
or OR4 (N5787, N5738, N5399, N4971, N920);
and AND2 (N5788, N5787, N5371);
and AND3 (N5789, N5779, N3560, N330);
buf BUF1 (N5790, N5782);
not NOT1 (N5791, N5762);
nor NOR2 (N5792, N5775, N4379);
or OR4 (N5793, N5783, N3693, N77, N5718);
nand NAND3 (N5794, N5790, N3786, N644);
xor XOR2 (N5795, N5789, N3514);
nor NOR3 (N5796, N5788, N5715, N4632);
buf BUF1 (N5797, N5794);
or OR2 (N5798, N5792, N4538);
not NOT1 (N5799, N5791);
or OR2 (N5800, N5793, N2758);
nor NOR2 (N5801, N5795, N2491);
not NOT1 (N5802, N5785);
not NOT1 (N5803, N5797);
nand NAND2 (N5804, N5786, N2110);
and AND4 (N5805, N5796, N679, N5202, N2245);
xor XOR2 (N5806, N5800, N1165);
and AND3 (N5807, N5804, N4865, N1543);
and AND3 (N5808, N5803, N4128, N1979);
xor XOR2 (N5809, N5808, N890);
nor NOR2 (N5810, N5807, N4740);
buf BUF1 (N5811, N5799);
xor XOR2 (N5812, N5801, N474);
buf BUF1 (N5813, N5798);
and AND2 (N5814, N5802, N2241);
nand NAND3 (N5815, N5812, N5414, N4023);
buf BUF1 (N5816, N5810);
nand NAND3 (N5817, N5816, N5067, N5003);
not NOT1 (N5818, N5817);
xor XOR2 (N5819, N5814, N5336);
xor XOR2 (N5820, N5809, N1100);
buf BUF1 (N5821, N5784);
and AND3 (N5822, N5819, N3962, N1714);
nand NAND4 (N5823, N5806, N493, N1786, N3125);
buf BUF1 (N5824, N5822);
xor XOR2 (N5825, N5813, N4057);
nor NOR2 (N5826, N5818, N4760);
not NOT1 (N5827, N5805);
nand NAND3 (N5828, N5772, N5617, N2221);
buf BUF1 (N5829, N5824);
xor XOR2 (N5830, N5815, N5068);
buf BUF1 (N5831, N5811);
and AND2 (N5832, N5820, N5638);
or OR4 (N5833, N5831, N3838, N402, N2745);
xor XOR2 (N5834, N5826, N5062);
nand NAND4 (N5835, N5827, N698, N3185, N3557);
and AND3 (N5836, N5835, N5282, N428);
and AND3 (N5837, N5828, N4060, N1670);
or OR4 (N5838, N5821, N4234, N4150, N4711);
not NOT1 (N5839, N5836);
not NOT1 (N5840, N5834);
nand NAND2 (N5841, N5825, N1223);
xor XOR2 (N5842, N5832, N5207);
not NOT1 (N5843, N5833);
and AND4 (N5844, N5839, N911, N4119, N5062);
nor NOR3 (N5845, N5830, N4291, N4110);
buf BUF1 (N5846, N5841);
and AND3 (N5847, N5838, N4397, N1751);
nor NOR2 (N5848, N5844, N3275);
and AND3 (N5849, N5823, N1273, N1836);
or OR3 (N5850, N5848, N1095, N155);
and AND4 (N5851, N5840, N393, N3989, N4428);
or OR3 (N5852, N5847, N2978, N1306);
not NOT1 (N5853, N5843);
nand NAND2 (N5854, N5846, N1763);
nand NAND2 (N5855, N5837, N4710);
nand NAND4 (N5856, N5851, N1294, N3395, N1989);
nor NOR3 (N5857, N5845, N5139, N1535);
nor NOR3 (N5858, N5842, N2291, N972);
not NOT1 (N5859, N5855);
or OR2 (N5860, N5858, N1469);
or OR2 (N5861, N5829, N3099);
nor NOR2 (N5862, N5859, N3219);
not NOT1 (N5863, N5862);
or OR2 (N5864, N5853, N5052);
nor NOR2 (N5865, N5852, N1040);
xor XOR2 (N5866, N5857, N3947);
nand NAND3 (N5867, N5854, N4379, N2562);
nand NAND2 (N5868, N5860, N4439);
buf BUF1 (N5869, N5867);
nand NAND4 (N5870, N5868, N5643, N4107, N1759);
and AND3 (N5871, N5850, N49, N2136);
not NOT1 (N5872, N5871);
buf BUF1 (N5873, N5856);
and AND3 (N5874, N5849, N140, N2760);
not NOT1 (N5875, N5864);
not NOT1 (N5876, N5865);
not NOT1 (N5877, N5866);
and AND4 (N5878, N5876, N4664, N3241, N5486);
buf BUF1 (N5879, N5873);
and AND2 (N5880, N5870, N4708);
nor NOR4 (N5881, N5872, N3757, N3045, N2366);
or OR2 (N5882, N5861, N2918);
nor NOR3 (N5883, N5869, N5104, N3822);
xor XOR2 (N5884, N5877, N3604);
xor XOR2 (N5885, N5863, N4220);
not NOT1 (N5886, N5880);
buf BUF1 (N5887, N5882);
or OR2 (N5888, N5883, N5338);
or OR4 (N5889, N5885, N1084, N4807, N3215);
buf BUF1 (N5890, N5887);
or OR4 (N5891, N5881, N3047, N2728, N5590);
nand NAND4 (N5892, N5875, N4512, N3924, N5144);
not NOT1 (N5893, N5892);
nand NAND2 (N5894, N5893, N2496);
xor XOR2 (N5895, N5879, N2202);
xor XOR2 (N5896, N5890, N5292);
nand NAND4 (N5897, N5884, N2808, N5198, N4797);
buf BUF1 (N5898, N5891);
and AND4 (N5899, N5894, N4958, N2299, N3067);
xor XOR2 (N5900, N5886, N4605);
nor NOR3 (N5901, N5878, N3740, N1685);
nand NAND2 (N5902, N5898, N4071);
nand NAND3 (N5903, N5902, N1006, N1120);
nor NOR2 (N5904, N5900, N4824);
nor NOR4 (N5905, N5903, N3900, N5208, N3920);
xor XOR2 (N5906, N5897, N4216);
or OR2 (N5907, N5874, N4579);
and AND2 (N5908, N5888, N572);
nor NOR3 (N5909, N5896, N2643, N2170);
nand NAND4 (N5910, N5901, N1482, N5000, N4708);
nand NAND2 (N5911, N5895, N1739);
not NOT1 (N5912, N5906);
buf BUF1 (N5913, N5909);
xor XOR2 (N5914, N5910, N5580);
xor XOR2 (N5915, N5905, N4674);
xor XOR2 (N5916, N5914, N2722);
not NOT1 (N5917, N5899);
buf BUF1 (N5918, N5916);
and AND4 (N5919, N5911, N1495, N5731, N4833);
not NOT1 (N5920, N5917);
and AND4 (N5921, N5912, N36, N1035, N1710);
nand NAND4 (N5922, N5904, N2538, N3482, N1034);
xor XOR2 (N5923, N5921, N5488);
and AND2 (N5924, N5889, N2759);
nor NOR4 (N5925, N5922, N5134, N5595, N5849);
and AND4 (N5926, N5919, N5667, N261, N2121);
buf BUF1 (N5927, N5918);
nor NOR4 (N5928, N5927, N4618, N4468, N3369);
buf BUF1 (N5929, N5928);
or OR2 (N5930, N5929, N541);
and AND2 (N5931, N5926, N1969);
xor XOR2 (N5932, N5907, N1406);
and AND4 (N5933, N5932, N2663, N4653, N5110);
buf BUF1 (N5934, N5923);
nor NOR3 (N5935, N5908, N4977, N1472);
buf BUF1 (N5936, N5935);
buf BUF1 (N5937, N5915);
buf BUF1 (N5938, N5924);
buf BUF1 (N5939, N5930);
or OR4 (N5940, N5936, N3262, N5720, N1995);
and AND3 (N5941, N5913, N1133, N5327);
buf BUF1 (N5942, N5925);
and AND2 (N5943, N5933, N4471);
or OR4 (N5944, N5940, N4775, N4442, N4554);
nand NAND2 (N5945, N5937, N3626);
nor NOR2 (N5946, N5931, N740);
buf BUF1 (N5947, N5920);
buf BUF1 (N5948, N5934);
nand NAND2 (N5949, N5943, N5144);
or OR2 (N5950, N5946, N5059);
or OR3 (N5951, N5944, N1943, N1852);
buf BUF1 (N5952, N5941);
buf BUF1 (N5953, N5939);
not NOT1 (N5954, N5952);
nand NAND3 (N5955, N5938, N2903, N655);
or OR2 (N5956, N5947, N1757);
nand NAND3 (N5957, N5951, N5785, N3151);
and AND4 (N5958, N5948, N2395, N1268, N3081);
xor XOR2 (N5959, N5949, N3299);
nor NOR3 (N5960, N5958, N1994, N2590);
or OR4 (N5961, N5945, N698, N1457, N5357);
buf BUF1 (N5962, N5954);
nor NOR4 (N5963, N5950, N4254, N3219, N701);
not NOT1 (N5964, N5960);
buf BUF1 (N5965, N5953);
nand NAND2 (N5966, N5956, N5892);
or OR4 (N5967, N5966, N2095, N2927, N3365);
buf BUF1 (N5968, N5965);
nor NOR3 (N5969, N5955, N1135, N5963);
or OR4 (N5970, N1914, N3521, N5545, N5284);
xor XOR2 (N5971, N5962, N5672);
or OR3 (N5972, N5942, N2487, N1857);
buf BUF1 (N5973, N5967);
not NOT1 (N5974, N5964);
not NOT1 (N5975, N5974);
nand NAND2 (N5976, N5970, N378);
nor NOR3 (N5977, N5959, N3007, N4311);
not NOT1 (N5978, N5961);
not NOT1 (N5979, N5976);
nor NOR3 (N5980, N5957, N2940, N3911);
nor NOR4 (N5981, N5968, N1841, N5518, N876);
nand NAND3 (N5982, N5978, N613, N1874);
and AND3 (N5983, N5971, N4762, N4558);
buf BUF1 (N5984, N5975);
buf BUF1 (N5985, N5980);
not NOT1 (N5986, N5972);
nor NOR4 (N5987, N5985, N496, N2439, N5245);
xor XOR2 (N5988, N5987, N5798);
and AND3 (N5989, N5979, N3115, N1161);
nand NAND2 (N5990, N5986, N3427);
not NOT1 (N5991, N5984);
or OR4 (N5992, N5990, N4379, N5394, N3835);
nor NOR4 (N5993, N5988, N5069, N1851, N2205);
and AND2 (N5994, N5981, N1355);
buf BUF1 (N5995, N5994);
buf BUF1 (N5996, N5995);
buf BUF1 (N5997, N5991);
or OR4 (N5998, N5973, N1364, N3704, N5401);
not NOT1 (N5999, N5993);
not NOT1 (N6000, N5969);
buf BUF1 (N6001, N6000);
nand NAND4 (N6002, N5982, N1316, N3175, N3067);
and AND3 (N6003, N6002, N85, N2177);
buf BUF1 (N6004, N5989);
nor NOR2 (N6005, N5977, N375);
not NOT1 (N6006, N5997);
not NOT1 (N6007, N5998);
nand NAND2 (N6008, N6001, N4997);
nor NOR2 (N6009, N5983, N1422);
buf BUF1 (N6010, N6004);
nor NOR2 (N6011, N6003, N4683);
and AND4 (N6012, N6011, N2955, N3887, N5812);
or OR4 (N6013, N6007, N3482, N3788, N1105);
buf BUF1 (N6014, N6012);
not NOT1 (N6015, N6010);
or OR3 (N6016, N6013, N1492, N935);
nor NOR4 (N6017, N6015, N355, N5613, N520);
buf BUF1 (N6018, N6016);
buf BUF1 (N6019, N6018);
and AND3 (N6020, N6019, N1663, N5366);
or OR2 (N6021, N5996, N2769);
nor NOR2 (N6022, N6020, N154);
or OR3 (N6023, N6005, N5348, N5005);
and AND3 (N6024, N6022, N5920, N5370);
not NOT1 (N6025, N6009);
and AND2 (N6026, N6021, N1956);
and AND2 (N6027, N5999, N4184);
buf BUF1 (N6028, N6023);
nor NOR3 (N6029, N6028, N2348, N2928);
or OR2 (N6030, N5992, N5240);
or OR3 (N6031, N6006, N52, N2024);
nor NOR2 (N6032, N6027, N2796);
nand NAND2 (N6033, N6025, N3092);
nand NAND3 (N6034, N6024, N4565, N2957);
not NOT1 (N6035, N6026);
not NOT1 (N6036, N6017);
nor NOR3 (N6037, N6029, N4065, N5239);
xor XOR2 (N6038, N6036, N3627);
and AND3 (N6039, N6035, N5566, N4987);
or OR3 (N6040, N6033, N5667, N3756);
buf BUF1 (N6041, N6031);
nor NOR4 (N6042, N6034, N5477, N136, N5427);
nand NAND4 (N6043, N6038, N2183, N3773, N5371);
xor XOR2 (N6044, N6039, N5259);
and AND2 (N6045, N6014, N1266);
buf BUF1 (N6046, N6042);
nand NAND4 (N6047, N6044, N2119, N5896, N4002);
not NOT1 (N6048, N6045);
buf BUF1 (N6049, N6048);
buf BUF1 (N6050, N6049);
and AND4 (N6051, N6032, N2358, N2011, N3462);
not NOT1 (N6052, N6046);
and AND4 (N6053, N6047, N408, N2192, N4346);
buf BUF1 (N6054, N6050);
or OR2 (N6055, N6040, N1292);
or OR2 (N6056, N6008, N3617);
not NOT1 (N6057, N6056);
xor XOR2 (N6058, N6055, N2421);
nand NAND3 (N6059, N6043, N2199, N1534);
or OR4 (N6060, N6041, N2134, N5237, N5847);
and AND2 (N6061, N6051, N1073);
not NOT1 (N6062, N6053);
nand NAND2 (N6063, N6059, N1680);
not NOT1 (N6064, N6054);
not NOT1 (N6065, N6061);
or OR2 (N6066, N6064, N5277);
buf BUF1 (N6067, N6066);
or OR4 (N6068, N6067, N139, N3262, N1757);
nand NAND4 (N6069, N6060, N3407, N1835, N567);
and AND4 (N6070, N6052, N5787, N2580, N1524);
or OR3 (N6071, N6030, N5036, N2281);
nor NOR3 (N6072, N6057, N1904, N673);
nand NAND4 (N6073, N6070, N5635, N5657, N3505);
xor XOR2 (N6074, N6073, N1669);
and AND4 (N6075, N6058, N1196, N3042, N3116);
not NOT1 (N6076, N6065);
xor XOR2 (N6077, N6062, N4939);
nand NAND2 (N6078, N6069, N544);
or OR2 (N6079, N6068, N4583);
xor XOR2 (N6080, N6077, N5032);
not NOT1 (N6081, N6074);
xor XOR2 (N6082, N6072, N2850);
or OR2 (N6083, N6080, N1645);
not NOT1 (N6084, N6079);
not NOT1 (N6085, N6076);
and AND4 (N6086, N6083, N453, N2211, N3813);
and AND2 (N6087, N6081, N4912);
xor XOR2 (N6088, N6082, N1459);
nand NAND3 (N6089, N6075, N5119, N4886);
and AND2 (N6090, N6078, N3037);
or OR4 (N6091, N6063, N2068, N2147, N245);
xor XOR2 (N6092, N6089, N841);
nor NOR4 (N6093, N6088, N5233, N4047, N4903);
and AND4 (N6094, N6093, N3004, N90, N1246);
buf BUF1 (N6095, N6071);
and AND2 (N6096, N6086, N3989);
and AND3 (N6097, N6037, N3116, N4207);
not NOT1 (N6098, N6094);
xor XOR2 (N6099, N6090, N5396);
nand NAND3 (N6100, N6092, N4849, N712);
nand NAND2 (N6101, N6099, N2756);
xor XOR2 (N6102, N6085, N5561);
not NOT1 (N6103, N6102);
or OR3 (N6104, N6098, N3869, N5029);
nand NAND2 (N6105, N6095, N2875);
and AND2 (N6106, N6097, N2033);
and AND3 (N6107, N6105, N326, N3891);
buf BUF1 (N6108, N6084);
nand NAND4 (N6109, N6107, N1912, N3444, N1558);
nor NOR4 (N6110, N6108, N2324, N4064, N2452);
or OR2 (N6111, N6100, N4494);
xor XOR2 (N6112, N6101, N2251);
nand NAND2 (N6113, N6096, N2462);
xor XOR2 (N6114, N6113, N3653);
or OR4 (N6115, N6112, N4806, N1774, N2554);
xor XOR2 (N6116, N6115, N1300);
nor NOR4 (N6117, N6109, N4816, N5814, N3233);
buf BUF1 (N6118, N6116);
or OR2 (N6119, N6118, N3466);
nor NOR2 (N6120, N6117, N2005);
and AND4 (N6121, N6104, N728, N3535, N1694);
xor XOR2 (N6122, N6106, N59);
xor XOR2 (N6123, N6091, N1194);
not NOT1 (N6124, N6111);
or OR2 (N6125, N6122, N6002);
not NOT1 (N6126, N6124);
xor XOR2 (N6127, N6123, N5312);
or OR3 (N6128, N6114, N757, N873);
nor NOR4 (N6129, N6125, N2068, N3748, N2312);
or OR3 (N6130, N6120, N1213, N1651);
nor NOR3 (N6131, N6103, N1618, N4506);
buf BUF1 (N6132, N6121);
nand NAND4 (N6133, N6129, N1027, N1174, N2391);
nand NAND4 (N6134, N6110, N6027, N1443, N2566);
or OR2 (N6135, N6133, N3798);
buf BUF1 (N6136, N6127);
not NOT1 (N6137, N6119);
buf BUF1 (N6138, N6134);
nor NOR3 (N6139, N6138, N3871, N2335);
nor NOR4 (N6140, N6128, N4210, N2634, N3767);
nand NAND4 (N6141, N6126, N2854, N4394, N2219);
and AND2 (N6142, N6141, N5913);
and AND3 (N6143, N6137, N1669, N3287);
nor NOR4 (N6144, N6136, N5744, N815, N1909);
nor NOR2 (N6145, N6132, N3096);
not NOT1 (N6146, N6131);
xor XOR2 (N6147, N6135, N3549);
nor NOR4 (N6148, N6143, N5726, N5493, N827);
or OR3 (N6149, N6139, N5095, N2336);
xor XOR2 (N6150, N6142, N826);
and AND2 (N6151, N6150, N298);
or OR2 (N6152, N6145, N1679);
or OR2 (N6153, N6087, N728);
nor NOR2 (N6154, N6146, N5649);
buf BUF1 (N6155, N6130);
or OR4 (N6156, N6153, N2847, N2051, N761);
buf BUF1 (N6157, N6156);
not NOT1 (N6158, N6148);
nor NOR3 (N6159, N6152, N2769, N2784);
nand NAND3 (N6160, N6157, N197, N1612);
and AND2 (N6161, N6151, N2651);
not NOT1 (N6162, N6158);
nor NOR4 (N6163, N6160, N536, N5938, N2872);
nand NAND3 (N6164, N6161, N532, N5497);
and AND2 (N6165, N6147, N3604);
not NOT1 (N6166, N6165);
not NOT1 (N6167, N6159);
and AND4 (N6168, N6164, N5463, N5509, N2496);
nand NAND2 (N6169, N6144, N2847);
buf BUF1 (N6170, N6163);
not NOT1 (N6171, N6166);
buf BUF1 (N6172, N6162);
buf BUF1 (N6173, N6169);
nand NAND2 (N6174, N6168, N5781);
buf BUF1 (N6175, N6149);
xor XOR2 (N6176, N6167, N501);
and AND2 (N6177, N6172, N3226);
nand NAND4 (N6178, N6155, N766, N4424, N4200);
xor XOR2 (N6179, N6177, N865);
xor XOR2 (N6180, N6140, N5007);
buf BUF1 (N6181, N6179);
or OR2 (N6182, N6181, N3119);
buf BUF1 (N6183, N6154);
and AND2 (N6184, N6176, N1650);
or OR4 (N6185, N6184, N3816, N2858, N4850);
or OR2 (N6186, N6173, N5643);
and AND4 (N6187, N6185, N630, N2934, N5478);
and AND3 (N6188, N6178, N1573, N4648);
buf BUF1 (N6189, N6171);
nand NAND4 (N6190, N6174, N406, N2741, N4304);
nor NOR2 (N6191, N6182, N524);
not NOT1 (N6192, N6186);
buf BUF1 (N6193, N6187);
nand NAND4 (N6194, N6188, N3130, N4213, N157);
nand NAND3 (N6195, N6192, N1603, N991);
and AND3 (N6196, N6193, N5872, N1268);
nor NOR2 (N6197, N6190, N4920);
xor XOR2 (N6198, N6183, N774);
not NOT1 (N6199, N6194);
buf BUF1 (N6200, N6175);
nor NOR3 (N6201, N6195, N5863, N5492);
and AND3 (N6202, N6199, N5951, N5029);
buf BUF1 (N6203, N6196);
and AND2 (N6204, N6198, N1907);
nor NOR3 (N6205, N6189, N1036, N1429);
not NOT1 (N6206, N6201);
buf BUF1 (N6207, N6170);
xor XOR2 (N6208, N6203, N3770);
and AND2 (N6209, N6204, N3096);
and AND4 (N6210, N6202, N1470, N2836, N4354);
xor XOR2 (N6211, N6206, N1346);
not NOT1 (N6212, N6208);
xor XOR2 (N6213, N6211, N3031);
and AND4 (N6214, N6207, N2547, N3239, N4439);
buf BUF1 (N6215, N6209);
nand NAND4 (N6216, N6213, N2950, N167, N2600);
nor NOR2 (N6217, N6197, N2399);
buf BUF1 (N6218, N6212);
buf BUF1 (N6219, N6216);
xor XOR2 (N6220, N6205, N3159);
xor XOR2 (N6221, N6191, N1289);
nand NAND2 (N6222, N6219, N209);
not NOT1 (N6223, N6210);
or OR2 (N6224, N6221, N2041);
and AND4 (N6225, N6223, N5906, N2840, N4187);
or OR2 (N6226, N6200, N4031);
nor NOR3 (N6227, N6217, N5442, N3960);
buf BUF1 (N6228, N6218);
or OR4 (N6229, N6224, N3095, N4529, N2996);
and AND3 (N6230, N6222, N968, N3527);
nand NAND3 (N6231, N6215, N2907, N5302);
not NOT1 (N6232, N6225);
and AND3 (N6233, N6227, N3161, N4200);
buf BUF1 (N6234, N6226);
buf BUF1 (N6235, N6234);
nor NOR3 (N6236, N6220, N2422, N4227);
or OR4 (N6237, N6180, N4028, N2483, N849);
or OR2 (N6238, N6233, N4164);
and AND3 (N6239, N6231, N927, N2011);
or OR3 (N6240, N6230, N3724, N3510);
buf BUF1 (N6241, N6228);
and AND2 (N6242, N6237, N1413);
or OR2 (N6243, N6242, N430);
or OR2 (N6244, N6236, N5492);
or OR3 (N6245, N6235, N3425, N5236);
buf BUF1 (N6246, N6245);
or OR3 (N6247, N6240, N5931, N1598);
xor XOR2 (N6248, N6246, N1088);
nor NOR2 (N6249, N6232, N146);
buf BUF1 (N6250, N6239);
nand NAND4 (N6251, N6249, N2032, N494, N5364);
buf BUF1 (N6252, N6229);
xor XOR2 (N6253, N6248, N4377);
nand NAND4 (N6254, N6253, N3235, N2580, N866);
xor XOR2 (N6255, N6243, N4537);
and AND3 (N6256, N6244, N3526, N5271);
not NOT1 (N6257, N6250);
buf BUF1 (N6258, N6254);
nand NAND4 (N6259, N6247, N4215, N1454, N3977);
buf BUF1 (N6260, N6256);
nand NAND3 (N6261, N6238, N5828, N2875);
buf BUF1 (N6262, N6259);
nand NAND3 (N6263, N6262, N2326, N3991);
not NOT1 (N6264, N6241);
nor NOR3 (N6265, N6261, N1679, N1454);
nor NOR3 (N6266, N6252, N527, N733);
nand NAND2 (N6267, N6258, N4161);
nor NOR4 (N6268, N6214, N1594, N5517, N2286);
nor NOR3 (N6269, N6267, N4363, N5383);
not NOT1 (N6270, N6265);
and AND3 (N6271, N6260, N4621, N2731);
not NOT1 (N6272, N6269);
nor NOR4 (N6273, N6270, N65, N2059, N22);
xor XOR2 (N6274, N6263, N5794);
not NOT1 (N6275, N6273);
nand NAND2 (N6276, N6268, N4763);
xor XOR2 (N6277, N6257, N4967);
nand NAND4 (N6278, N6255, N1730, N2019, N44);
and AND3 (N6279, N6276, N1878, N1915);
xor XOR2 (N6280, N6277, N39);
and AND2 (N6281, N6279, N736);
and AND2 (N6282, N6266, N5503);
not NOT1 (N6283, N6278);
nor NOR2 (N6284, N6272, N4376);
not NOT1 (N6285, N6282);
buf BUF1 (N6286, N6283);
nand NAND2 (N6287, N6264, N5558);
nand NAND2 (N6288, N6284, N727);
or OR3 (N6289, N6281, N978, N4216);
buf BUF1 (N6290, N6287);
xor XOR2 (N6291, N6280, N4043);
nor NOR2 (N6292, N6290, N4853);
buf BUF1 (N6293, N6288);
not NOT1 (N6294, N6285);
or OR2 (N6295, N6291, N3695);
nand NAND2 (N6296, N6251, N2798);
and AND4 (N6297, N6286, N699, N5900, N4048);
xor XOR2 (N6298, N6295, N3973);
buf BUF1 (N6299, N6294);
nand NAND2 (N6300, N6274, N5193);
nor NOR2 (N6301, N6293, N3800);
xor XOR2 (N6302, N6292, N2243);
not NOT1 (N6303, N6302);
nor NOR3 (N6304, N6289, N3861, N812);
or OR4 (N6305, N6300, N961, N4572, N22);
not NOT1 (N6306, N6299);
or OR4 (N6307, N6304, N2350, N6090, N4217);
not NOT1 (N6308, N6296);
nand NAND3 (N6309, N6297, N5694, N3597);
not NOT1 (N6310, N6298);
not NOT1 (N6311, N6305);
or OR4 (N6312, N6307, N5526, N3707, N2812);
nand NAND4 (N6313, N6310, N2116, N2610, N6277);
and AND2 (N6314, N6308, N5714);
or OR3 (N6315, N6313, N3683, N4906);
xor XOR2 (N6316, N6301, N6076);
not NOT1 (N6317, N6303);
and AND4 (N6318, N6311, N3381, N155, N5029);
buf BUF1 (N6319, N6318);
or OR3 (N6320, N6315, N1931, N168);
or OR2 (N6321, N6319, N6016);
buf BUF1 (N6322, N6320);
nor NOR4 (N6323, N6306, N4131, N6122, N95);
nand NAND4 (N6324, N6271, N615, N6103, N425);
buf BUF1 (N6325, N6309);
nor NOR3 (N6326, N6316, N3143, N589);
and AND2 (N6327, N6275, N2356);
or OR3 (N6328, N6323, N3204, N1815);
not NOT1 (N6329, N6322);
and AND4 (N6330, N6325, N408, N3597, N1485);
not NOT1 (N6331, N6329);
buf BUF1 (N6332, N6321);
nor NOR3 (N6333, N6317, N135, N2446);
nor NOR3 (N6334, N6333, N1263, N4769);
xor XOR2 (N6335, N6326, N750);
not NOT1 (N6336, N6324);
xor XOR2 (N6337, N6327, N1482);
buf BUF1 (N6338, N6312);
nand NAND3 (N6339, N6337, N1628, N1981);
nor NOR3 (N6340, N6335, N3390, N1239);
nand NAND4 (N6341, N6331, N1638, N4198, N2454);
nor NOR4 (N6342, N6328, N5549, N5768, N5279);
not NOT1 (N6343, N6339);
or OR2 (N6344, N6336, N3169);
nor NOR4 (N6345, N6330, N5187, N5717, N5997);
buf BUF1 (N6346, N6332);
nand NAND4 (N6347, N6345, N1360, N187, N853);
not NOT1 (N6348, N6346);
and AND2 (N6349, N6334, N3141);
or OR4 (N6350, N6347, N248, N4823, N5364);
not NOT1 (N6351, N6350);
and AND4 (N6352, N6351, N1761, N6130, N2311);
not NOT1 (N6353, N6342);
not NOT1 (N6354, N6341);
or OR3 (N6355, N6340, N4105, N1381);
not NOT1 (N6356, N6353);
or OR4 (N6357, N6352, N4234, N3114, N4227);
and AND4 (N6358, N6356, N5888, N5627, N578);
buf BUF1 (N6359, N6338);
or OR3 (N6360, N6357, N2953, N5538);
xor XOR2 (N6361, N6360, N5159);
nand NAND3 (N6362, N6314, N4532, N2775);
nor NOR2 (N6363, N6362, N1603);
nand NAND4 (N6364, N6344, N1950, N3144, N1497);
and AND4 (N6365, N6349, N3121, N1526, N5404);
and AND4 (N6366, N6355, N5531, N3809, N1164);
buf BUF1 (N6367, N6354);
or OR2 (N6368, N6361, N1652);
buf BUF1 (N6369, N6368);
not NOT1 (N6370, N6358);
nand NAND2 (N6371, N6343, N2949);
xor XOR2 (N6372, N6371, N822);
nor NOR3 (N6373, N6363, N4773, N3268);
nand NAND4 (N6374, N6366, N3376, N1680, N3309);
xor XOR2 (N6375, N6373, N5863);
or OR3 (N6376, N6375, N1440, N3267);
nor NOR4 (N6377, N6364, N2424, N6343, N638);
xor XOR2 (N6378, N6377, N4240);
nor NOR4 (N6379, N6376, N2081, N5017, N1509);
xor XOR2 (N6380, N6365, N926);
nand NAND3 (N6381, N6348, N2294, N4106);
nor NOR3 (N6382, N6378, N441, N1416);
or OR4 (N6383, N6380, N436, N2384, N533);
nand NAND2 (N6384, N6374, N3435);
nand NAND3 (N6385, N6384, N4782, N2807);
nand NAND2 (N6386, N6385, N4079);
xor XOR2 (N6387, N6369, N3407);
nor NOR4 (N6388, N6387, N2002, N3244, N338);
xor XOR2 (N6389, N6381, N5109);
xor XOR2 (N6390, N6370, N4780);
or OR4 (N6391, N6389, N944, N6376, N1105);
xor XOR2 (N6392, N6386, N2464);
buf BUF1 (N6393, N6391);
or OR2 (N6394, N6367, N5913);
xor XOR2 (N6395, N6359, N1284);
or OR3 (N6396, N6379, N1718, N2221);
xor XOR2 (N6397, N6388, N5599);
buf BUF1 (N6398, N6397);
nor NOR3 (N6399, N6383, N2234, N5354);
or OR2 (N6400, N6372, N83);
buf BUF1 (N6401, N6382);
nand NAND4 (N6402, N6400, N3983, N2485, N5431);
or OR3 (N6403, N6393, N6031, N4233);
and AND4 (N6404, N6390, N576, N1854, N4805);
and AND3 (N6405, N6404, N607, N3592);
not NOT1 (N6406, N6405);
nand NAND2 (N6407, N6401, N5895);
nand NAND3 (N6408, N6392, N4181, N849);
and AND2 (N6409, N6396, N6263);
nand NAND3 (N6410, N6407, N4154, N2444);
nand NAND3 (N6411, N6406, N4848, N5970);
nand NAND2 (N6412, N6394, N2850);
or OR2 (N6413, N6409, N2208);
nor NOR2 (N6414, N6403, N3552);
xor XOR2 (N6415, N6414, N3390);
xor XOR2 (N6416, N6412, N68);
or OR3 (N6417, N6411, N3391, N5795);
not NOT1 (N6418, N6413);
buf BUF1 (N6419, N6410);
not NOT1 (N6420, N6415);
not NOT1 (N6421, N6420);
xor XOR2 (N6422, N6398, N2002);
or OR2 (N6423, N6402, N1372);
and AND2 (N6424, N6423, N4701);
buf BUF1 (N6425, N6408);
and AND2 (N6426, N6417, N5335);
or OR2 (N6427, N6395, N1161);
buf BUF1 (N6428, N6426);
xor XOR2 (N6429, N6416, N346);
xor XOR2 (N6430, N6418, N3501);
not NOT1 (N6431, N6399);
not NOT1 (N6432, N6424);
xor XOR2 (N6433, N6428, N4175);
xor XOR2 (N6434, N6419, N688);
or OR3 (N6435, N6431, N2543, N910);
xor XOR2 (N6436, N6430, N456);
nand NAND3 (N6437, N6435, N723, N2102);
not NOT1 (N6438, N6421);
not NOT1 (N6439, N6427);
not NOT1 (N6440, N6432);
or OR4 (N6441, N6433, N4393, N251, N1568);
not NOT1 (N6442, N6439);
not NOT1 (N6443, N6442);
xor XOR2 (N6444, N6422, N917);
not NOT1 (N6445, N6441);
nand NAND3 (N6446, N6443, N5814, N4310);
nor NOR3 (N6447, N6429, N141, N1889);
and AND2 (N6448, N6437, N3198);
not NOT1 (N6449, N6446);
nor NOR4 (N6450, N6444, N4700, N5473, N4688);
or OR3 (N6451, N6449, N3801, N3424);
nor NOR4 (N6452, N6438, N5686, N1218, N1554);
nor NOR2 (N6453, N6434, N2177);
and AND3 (N6454, N6452, N6359, N5231);
and AND3 (N6455, N6436, N5464, N4538);
buf BUF1 (N6456, N6445);
nor NOR4 (N6457, N6440, N2636, N1249, N1814);
buf BUF1 (N6458, N6453);
xor XOR2 (N6459, N6447, N5160);
nor NOR3 (N6460, N6450, N5795, N5306);
xor XOR2 (N6461, N6459, N424);
or OR4 (N6462, N6425, N1875, N190, N176);
nor NOR3 (N6463, N6460, N6259, N2966);
xor XOR2 (N6464, N6461, N5832);
buf BUF1 (N6465, N6454);
xor XOR2 (N6466, N6456, N4173);
not NOT1 (N6467, N6466);
buf BUF1 (N6468, N6455);
and AND3 (N6469, N6458, N6329, N4647);
nand NAND3 (N6470, N6462, N4053, N4626);
buf BUF1 (N6471, N6463);
nand NAND2 (N6472, N6469, N1965);
or OR4 (N6473, N6465, N4804, N2772, N1376);
not NOT1 (N6474, N6467);
nor NOR4 (N6475, N6464, N3148, N3947, N2953);
or OR3 (N6476, N6475, N819, N6393);
and AND2 (N6477, N6471, N2980);
nor NOR4 (N6478, N6470, N4572, N4967, N5080);
or OR4 (N6479, N6468, N1311, N70, N642);
not NOT1 (N6480, N6457);
nor NOR3 (N6481, N6448, N3001, N3989);
and AND3 (N6482, N6477, N4875, N1958);
nor NOR4 (N6483, N6474, N872, N1758, N1841);
xor XOR2 (N6484, N6479, N1341);
xor XOR2 (N6485, N6473, N360);
or OR2 (N6486, N6485, N1819);
or OR2 (N6487, N6478, N3013);
not NOT1 (N6488, N6481);
and AND3 (N6489, N6472, N2677, N4808);
buf BUF1 (N6490, N6480);
xor XOR2 (N6491, N6487, N4939);
xor XOR2 (N6492, N6482, N1697);
or OR3 (N6493, N6491, N1758, N1252);
and AND3 (N6494, N6451, N5100, N441);
not NOT1 (N6495, N6486);
xor XOR2 (N6496, N6483, N3988);
xor XOR2 (N6497, N6484, N427);
xor XOR2 (N6498, N6493, N1876);
not NOT1 (N6499, N6496);
buf BUF1 (N6500, N6497);
and AND2 (N6501, N6494, N2099);
not NOT1 (N6502, N6501);
nor NOR2 (N6503, N6488, N3772);
not NOT1 (N6504, N6489);
nand NAND4 (N6505, N6499, N4747, N4776, N5542);
or OR3 (N6506, N6503, N1047, N319);
not NOT1 (N6507, N6492);
nor NOR3 (N6508, N6504, N2124, N1292);
not NOT1 (N6509, N6508);
nand NAND3 (N6510, N6498, N2168, N5149);
and AND3 (N6511, N6510, N5847, N5701);
not NOT1 (N6512, N6500);
nand NAND4 (N6513, N6511, N3804, N6412, N6022);
xor XOR2 (N6514, N6505, N5229);
not NOT1 (N6515, N6512);
and AND3 (N6516, N6507, N2042, N976);
or OR2 (N6517, N6516, N4608);
buf BUF1 (N6518, N6517);
or OR4 (N6519, N6502, N5750, N3710, N6181);
or OR4 (N6520, N6490, N4325, N329, N2584);
nand NAND2 (N6521, N6520, N5887);
nand NAND2 (N6522, N6515, N286);
nand NAND3 (N6523, N6476, N6108, N2298);
buf BUF1 (N6524, N6513);
and AND2 (N6525, N6522, N6065);
buf BUF1 (N6526, N6519);
xor XOR2 (N6527, N6523, N3842);
buf BUF1 (N6528, N6526);
not NOT1 (N6529, N6514);
not NOT1 (N6530, N6528);
nand NAND3 (N6531, N6518, N206, N1074);
or OR4 (N6532, N6531, N5096, N4682, N1611);
and AND4 (N6533, N6495, N1907, N3633, N5317);
or OR4 (N6534, N6530, N5242, N60, N1969);
not NOT1 (N6535, N6525);
buf BUF1 (N6536, N6533);
buf BUF1 (N6537, N6527);
and AND3 (N6538, N6532, N5781, N1028);
buf BUF1 (N6539, N6524);
nand NAND4 (N6540, N6529, N3726, N5041, N1891);
nand NAND2 (N6541, N6537, N5804);
nor NOR2 (N6542, N6538, N5833);
nor NOR2 (N6543, N6539, N5834);
not NOT1 (N6544, N6542);
and AND4 (N6545, N6544, N6068, N758, N4789);
xor XOR2 (N6546, N6535, N5306);
buf BUF1 (N6547, N6546);
nor NOR3 (N6548, N6534, N6199, N507);
nor NOR2 (N6549, N6548, N5138);
or OR3 (N6550, N6547, N1288, N3086);
and AND4 (N6551, N6545, N6132, N4238, N627);
buf BUF1 (N6552, N6509);
or OR3 (N6553, N6551, N3994, N1457);
nand NAND3 (N6554, N6536, N1691, N6066);
nor NOR3 (N6555, N6549, N5681, N3243);
xor XOR2 (N6556, N6506, N1672);
not NOT1 (N6557, N6521);
or OR2 (N6558, N6541, N3365);
not NOT1 (N6559, N6558);
nand NAND2 (N6560, N6550, N1937);
and AND3 (N6561, N6552, N2116, N2358);
nand NAND2 (N6562, N6555, N468);
nand NAND2 (N6563, N6554, N3143);
not NOT1 (N6564, N6557);
nand NAND4 (N6565, N6564, N2789, N515, N4619);
not NOT1 (N6566, N6562);
not NOT1 (N6567, N6560);
or OR4 (N6568, N6567, N1099, N6366, N5388);
xor XOR2 (N6569, N6563, N6455);
buf BUF1 (N6570, N6561);
or OR4 (N6571, N6568, N2655, N5689, N110);
nand NAND4 (N6572, N6553, N2935, N1239, N4343);
or OR2 (N6573, N6565, N628);
xor XOR2 (N6574, N6559, N5642);
nor NOR2 (N6575, N6570, N3971);
or OR4 (N6576, N6571, N1696, N2775, N1441);
and AND4 (N6577, N6573, N2334, N844, N4516);
not NOT1 (N6578, N6577);
and AND3 (N6579, N6569, N5815, N1105);
not NOT1 (N6580, N6578);
and AND2 (N6581, N6580, N3734);
xor XOR2 (N6582, N6576, N783);
or OR3 (N6583, N6575, N1355, N3658);
and AND2 (N6584, N6583, N4823);
or OR4 (N6585, N6543, N1609, N538, N6301);
xor XOR2 (N6586, N6579, N2296);
buf BUF1 (N6587, N6585);
or OR4 (N6588, N6587, N5523, N1579, N3383);
nor NOR3 (N6589, N6588, N3338, N5053);
not NOT1 (N6590, N6540);
and AND4 (N6591, N6586, N5969, N2517, N1335);
not NOT1 (N6592, N6582);
or OR3 (N6593, N6589, N3726, N887);
and AND2 (N6594, N6556, N5654);
nor NOR4 (N6595, N6590, N4146, N3982, N1893);
nand NAND2 (N6596, N6591, N572);
nor NOR2 (N6597, N6592, N5998);
nor NOR3 (N6598, N6566, N2131, N1205);
xor XOR2 (N6599, N6574, N4776);
not NOT1 (N6600, N6595);
buf BUF1 (N6601, N6572);
and AND2 (N6602, N6581, N1852);
xor XOR2 (N6603, N6601, N4680);
not NOT1 (N6604, N6599);
and AND2 (N6605, N6600, N4881);
xor XOR2 (N6606, N6605, N2017);
buf BUF1 (N6607, N6597);
or OR3 (N6608, N6602, N967, N55);
nand NAND4 (N6609, N6596, N3704, N1250, N330);
nor NOR3 (N6610, N6607, N1428, N1857);
xor XOR2 (N6611, N6606, N3966);
and AND2 (N6612, N6598, N3968);
buf BUF1 (N6613, N6611);
not NOT1 (N6614, N6604);
and AND2 (N6615, N6594, N2612);
and AND3 (N6616, N6615, N3137, N1374);
and AND4 (N6617, N6614, N1405, N4837, N5304);
xor XOR2 (N6618, N6612, N5669);
or OR2 (N6619, N6609, N5379);
xor XOR2 (N6620, N6618, N3450);
and AND4 (N6621, N6616, N1145, N290, N1541);
nor NOR4 (N6622, N6603, N4557, N5905, N1243);
and AND4 (N6623, N6608, N1399, N3314, N1617);
and AND2 (N6624, N6619, N4902);
nand NAND4 (N6625, N6584, N3749, N2737, N1602);
xor XOR2 (N6626, N6593, N2275);
xor XOR2 (N6627, N6613, N529);
nor NOR3 (N6628, N6626, N508, N228);
or OR2 (N6629, N6624, N5337);
buf BUF1 (N6630, N6623);
and AND2 (N6631, N6629, N3774);
and AND4 (N6632, N6617, N5969, N3583, N1978);
nand NAND3 (N6633, N6630, N6188, N5943);
or OR4 (N6634, N6621, N2063, N5607, N890);
xor XOR2 (N6635, N6610, N4116);
buf BUF1 (N6636, N6634);
and AND2 (N6637, N6627, N3605);
or OR4 (N6638, N6636, N2143, N646, N1500);
or OR4 (N6639, N6635, N1186, N1245, N966);
and AND4 (N6640, N6632, N1215, N1828, N4046);
nand NAND2 (N6641, N6628, N2520);
nand NAND2 (N6642, N6620, N601);
nor NOR4 (N6643, N6622, N415, N3666, N526);
buf BUF1 (N6644, N6625);
nor NOR2 (N6645, N6643, N5762);
not NOT1 (N6646, N6641);
nor NOR2 (N6647, N6640, N1742);
nor NOR3 (N6648, N6644, N4934, N5394);
nand NAND2 (N6649, N6638, N4613);
and AND4 (N6650, N6642, N4270, N3746, N5912);
or OR4 (N6651, N6647, N4402, N4882, N3898);
not NOT1 (N6652, N6645);
xor XOR2 (N6653, N6648, N1990);
nand NAND4 (N6654, N6633, N3230, N1638, N985);
nor NOR3 (N6655, N6637, N3345, N3801);
nor NOR3 (N6656, N6651, N3979, N3168);
or OR4 (N6657, N6650, N2335, N202, N1881);
xor XOR2 (N6658, N6655, N1557);
nor NOR3 (N6659, N6653, N6151, N3667);
nor NOR2 (N6660, N6654, N5195);
buf BUF1 (N6661, N6660);
buf BUF1 (N6662, N6656);
not NOT1 (N6663, N6646);
buf BUF1 (N6664, N6657);
and AND4 (N6665, N6639, N2134, N4785, N654);
xor XOR2 (N6666, N6661, N6658);
or OR3 (N6667, N112, N6278, N1938);
or OR3 (N6668, N6631, N6060, N6613);
and AND4 (N6669, N6663, N3579, N5020, N3175);
buf BUF1 (N6670, N6652);
nand NAND2 (N6671, N6670, N3374);
or OR2 (N6672, N6666, N5265);
buf BUF1 (N6673, N6662);
and AND3 (N6674, N6667, N5614, N2085);
xor XOR2 (N6675, N6649, N403);
nand NAND4 (N6676, N6665, N2018, N355, N6669);
nand NAND2 (N6677, N1518, N3623);
nand NAND4 (N6678, N6675, N5875, N4979, N4620);
xor XOR2 (N6679, N6672, N491);
or OR2 (N6680, N6671, N4321);
xor XOR2 (N6681, N6679, N6092);
buf BUF1 (N6682, N6681);
or OR2 (N6683, N6673, N4118);
nand NAND3 (N6684, N6680, N3101, N2156);
or OR3 (N6685, N6674, N2844, N4115);
xor XOR2 (N6686, N6668, N1948);
buf BUF1 (N6687, N6664);
buf BUF1 (N6688, N6686);
or OR2 (N6689, N6682, N3447);
nand NAND2 (N6690, N6688, N5264);
xor XOR2 (N6691, N6678, N3475);
or OR3 (N6692, N6685, N4334, N4178);
not NOT1 (N6693, N6683);
buf BUF1 (N6694, N6693);
or OR4 (N6695, N6689, N2698, N5197, N6089);
xor XOR2 (N6696, N6694, N1389);
buf BUF1 (N6697, N6695);
and AND2 (N6698, N6697, N5057);
or OR2 (N6699, N6677, N4594);
and AND3 (N6700, N6687, N3567, N618);
not NOT1 (N6701, N6699);
xor XOR2 (N6702, N6684, N296);
or OR4 (N6703, N6696, N3633, N3068, N5202);
not NOT1 (N6704, N6700);
xor XOR2 (N6705, N6702, N6293);
xor XOR2 (N6706, N6705, N750);
buf BUF1 (N6707, N6691);
xor XOR2 (N6708, N6698, N4564);
and AND4 (N6709, N6704, N2105, N911, N3382);
xor XOR2 (N6710, N6690, N1170);
xor XOR2 (N6711, N6707, N314);
nor NOR4 (N6712, N6659, N1904, N667, N6316);
buf BUF1 (N6713, N6709);
or OR3 (N6714, N6676, N869, N2354);
nand NAND2 (N6715, N6712, N6071);
and AND4 (N6716, N6715, N3638, N312, N2491);
or OR2 (N6717, N6710, N2491);
not NOT1 (N6718, N6703);
buf BUF1 (N6719, N6708);
buf BUF1 (N6720, N6713);
nand NAND2 (N6721, N6714, N568);
xor XOR2 (N6722, N6701, N2615);
nor NOR4 (N6723, N6711, N2965, N2780, N2067);
nand NAND2 (N6724, N6692, N5376);
xor XOR2 (N6725, N6720, N6011);
or OR2 (N6726, N6719, N6560);
buf BUF1 (N6727, N6722);
buf BUF1 (N6728, N6727);
or OR3 (N6729, N6718, N4106, N1948);
buf BUF1 (N6730, N6716);
and AND2 (N6731, N6717, N5367);
buf BUF1 (N6732, N6706);
or OR2 (N6733, N6728, N3023);
nor NOR2 (N6734, N6724, N2374);
nand NAND3 (N6735, N6732, N2150, N6649);
nand NAND3 (N6736, N6733, N6669, N4422);
and AND2 (N6737, N6725, N592);
not NOT1 (N6738, N6735);
or OR3 (N6739, N6736, N4910, N1577);
nand NAND3 (N6740, N6734, N1630, N1856);
buf BUF1 (N6741, N6723);
xor XOR2 (N6742, N6731, N897);
or OR2 (N6743, N6740, N1522);
nand NAND2 (N6744, N6738, N441);
not NOT1 (N6745, N6726);
or OR2 (N6746, N6744, N6196);
or OR4 (N6747, N6746, N5497, N3745, N6053);
and AND3 (N6748, N6741, N3603, N2788);
not NOT1 (N6749, N6747);
not NOT1 (N6750, N6730);
nor NOR4 (N6751, N6729, N4639, N3755, N3984);
not NOT1 (N6752, N6743);
not NOT1 (N6753, N6721);
nor NOR3 (N6754, N6753, N5908, N5223);
nor NOR3 (N6755, N6745, N265, N733);
or OR2 (N6756, N6750, N2);
or OR4 (N6757, N6754, N6059, N4698, N3203);
and AND4 (N6758, N6755, N197, N922, N6149);
xor XOR2 (N6759, N6752, N6463);
not NOT1 (N6760, N6737);
nand NAND4 (N6761, N6756, N2776, N609, N1610);
nor NOR4 (N6762, N6739, N3525, N4213, N3289);
buf BUF1 (N6763, N6762);
buf BUF1 (N6764, N6757);
not NOT1 (N6765, N6751);
not NOT1 (N6766, N6763);
or OR2 (N6767, N6764, N1444);
or OR3 (N6768, N6759, N2148, N6119);
or OR3 (N6769, N6758, N2988, N5453);
not NOT1 (N6770, N6768);
xor XOR2 (N6771, N6761, N3730);
nor NOR3 (N6772, N6769, N1973, N3957);
or OR4 (N6773, N6765, N6682, N3922, N4354);
and AND4 (N6774, N6760, N540, N3270, N1474);
buf BUF1 (N6775, N6771);
nor NOR2 (N6776, N6773, N801);
and AND2 (N6777, N6742, N2081);
buf BUF1 (N6778, N6767);
nor NOR2 (N6779, N6749, N6723);
not NOT1 (N6780, N6774);
nor NOR2 (N6781, N6779, N6207);
not NOT1 (N6782, N6781);
nor NOR3 (N6783, N6775, N5477, N3225);
not NOT1 (N6784, N6780);
nand NAND3 (N6785, N6783, N2914, N2639);
xor XOR2 (N6786, N6777, N2303);
not NOT1 (N6787, N6772);
xor XOR2 (N6788, N6776, N6409);
and AND2 (N6789, N6785, N4699);
and AND2 (N6790, N6787, N2628);
nand NAND2 (N6791, N6778, N111);
nand NAND3 (N6792, N6790, N6399, N2040);
nand NAND3 (N6793, N6786, N6638, N6179);
not NOT1 (N6794, N6791);
or OR3 (N6795, N6788, N3360, N2511);
or OR3 (N6796, N6770, N2175, N3526);
and AND3 (N6797, N6789, N6197, N5280);
xor XOR2 (N6798, N6794, N5151);
not NOT1 (N6799, N6792);
buf BUF1 (N6800, N6748);
nor NOR4 (N6801, N6766, N5420, N4440, N3943);
buf BUF1 (N6802, N6798);
nand NAND4 (N6803, N6799, N6586, N4420, N6052);
not NOT1 (N6804, N6784);
nor NOR2 (N6805, N6800, N5432);
or OR2 (N6806, N6801, N5322);
buf BUF1 (N6807, N6797);
nand NAND4 (N6808, N6806, N2755, N4262, N6326);
nor NOR2 (N6809, N6807, N1396);
buf BUF1 (N6810, N6796);
buf BUF1 (N6811, N6793);
nor NOR3 (N6812, N6809, N795, N2447);
not NOT1 (N6813, N6803);
nand NAND3 (N6814, N6805, N4411, N5383);
not NOT1 (N6815, N6813);
and AND4 (N6816, N6808, N5717, N6357, N1155);
not NOT1 (N6817, N6816);
and AND3 (N6818, N6814, N6272, N618);
and AND2 (N6819, N6802, N6160);
nand NAND4 (N6820, N6818, N1410, N518, N2612);
and AND4 (N6821, N6817, N4423, N5286, N6561);
and AND2 (N6822, N6815, N5352);
or OR2 (N6823, N6804, N6383);
buf BUF1 (N6824, N6782);
or OR3 (N6825, N6822, N897, N1080);
nor NOR4 (N6826, N6825, N5902, N2693, N3944);
and AND4 (N6827, N6812, N3780, N5333, N6094);
nor NOR2 (N6828, N6819, N705);
xor XOR2 (N6829, N6810, N919);
not NOT1 (N6830, N6826);
xor XOR2 (N6831, N6820, N1935);
buf BUF1 (N6832, N6829);
and AND4 (N6833, N6795, N906, N6097, N4200);
nand NAND2 (N6834, N6830, N2749);
or OR4 (N6835, N6833, N3368, N3957, N5675);
nand NAND4 (N6836, N6827, N5930, N2076, N2862);
nand NAND3 (N6837, N6832, N5030, N3534);
buf BUF1 (N6838, N6831);
and AND3 (N6839, N6828, N1455, N437);
xor XOR2 (N6840, N6834, N1948);
xor XOR2 (N6841, N6839, N6668);
nand NAND4 (N6842, N6811, N5619, N2576, N6454);
and AND3 (N6843, N6838, N2873, N1176);
buf BUF1 (N6844, N6837);
xor XOR2 (N6845, N6835, N6502);
nor NOR4 (N6846, N6841, N2467, N945, N1153);
nor NOR4 (N6847, N6844, N6722, N6109, N5627);
xor XOR2 (N6848, N6842, N1795);
nand NAND4 (N6849, N6823, N4023, N5853, N3959);
xor XOR2 (N6850, N6847, N2494);
nand NAND2 (N6851, N6846, N4926);
buf BUF1 (N6852, N6850);
not NOT1 (N6853, N6849);
or OR4 (N6854, N6845, N987, N3593, N1716);
nand NAND3 (N6855, N6821, N4158, N6809);
xor XOR2 (N6856, N6843, N2069);
buf BUF1 (N6857, N6852);
xor XOR2 (N6858, N6824, N1580);
buf BUF1 (N6859, N6836);
xor XOR2 (N6860, N6855, N4745);
nand NAND3 (N6861, N6857, N4287, N3530);
nor NOR3 (N6862, N6840, N822, N214);
not NOT1 (N6863, N6851);
nor NOR2 (N6864, N6858, N1111);
not NOT1 (N6865, N6853);
buf BUF1 (N6866, N6854);
or OR4 (N6867, N6859, N504, N2038, N1902);
buf BUF1 (N6868, N6864);
and AND2 (N6869, N6866, N4108);
nand NAND4 (N6870, N6869, N1786, N4507, N3095);
nand NAND4 (N6871, N6848, N1657, N5845, N6113);
not NOT1 (N6872, N6867);
or OR3 (N6873, N6868, N5822, N2123);
nand NAND2 (N6874, N6860, N4215);
xor XOR2 (N6875, N6870, N3872);
and AND2 (N6876, N6875, N2666);
and AND2 (N6877, N6871, N528);
xor XOR2 (N6878, N6856, N4336);
nor NOR2 (N6879, N6873, N5248);
nand NAND3 (N6880, N6879, N652, N6674);
and AND4 (N6881, N6874, N671, N903, N4297);
buf BUF1 (N6882, N6878);
xor XOR2 (N6883, N6876, N800);
xor XOR2 (N6884, N6882, N730);
or OR2 (N6885, N6861, N1749);
not NOT1 (N6886, N6872);
xor XOR2 (N6887, N6881, N3525);
or OR3 (N6888, N6877, N4494, N354);
and AND3 (N6889, N6862, N1345, N2098);
and AND2 (N6890, N6863, N6313);
buf BUF1 (N6891, N6885);
buf BUF1 (N6892, N6889);
nor NOR2 (N6893, N6891, N2610);
nand NAND2 (N6894, N6888, N5829);
nand NAND2 (N6895, N6894, N4620);
nand NAND2 (N6896, N6887, N4527);
nor NOR4 (N6897, N6896, N372, N395, N2807);
nor NOR4 (N6898, N6865, N2592, N6669, N3989);
nor NOR4 (N6899, N6890, N2192, N860, N5526);
buf BUF1 (N6900, N6899);
xor XOR2 (N6901, N6900, N553);
nand NAND2 (N6902, N6895, N3248);
or OR3 (N6903, N6902, N5462, N2819);
and AND4 (N6904, N6883, N88, N2371, N1861);
xor XOR2 (N6905, N6904, N3169);
and AND2 (N6906, N6880, N801);
nand NAND4 (N6907, N6884, N305, N3942, N5234);
nor NOR4 (N6908, N6907, N1642, N5323, N1800);
xor XOR2 (N6909, N6906, N5419);
or OR4 (N6910, N6909, N4210, N6465, N1344);
not NOT1 (N6911, N6910);
nor NOR3 (N6912, N6892, N5404, N2567);
xor XOR2 (N6913, N6897, N582);
nand NAND2 (N6914, N6901, N6786);
nand NAND2 (N6915, N6903, N359);
nor NOR4 (N6916, N6913, N884, N4813, N3348);
or OR3 (N6917, N6908, N4230, N2937);
not NOT1 (N6918, N6916);
not NOT1 (N6919, N6918);
not NOT1 (N6920, N6911);
and AND3 (N6921, N6886, N631, N1855);
and AND2 (N6922, N6921, N158);
nor NOR3 (N6923, N6914, N4778, N516);
and AND4 (N6924, N6919, N882, N3526, N5911);
buf BUF1 (N6925, N6915);
nor NOR4 (N6926, N6920, N6785, N1924, N5736);
and AND4 (N6927, N6925, N2776, N5879, N2534);
buf BUF1 (N6928, N6926);
or OR2 (N6929, N6917, N4583);
not NOT1 (N6930, N6905);
or OR2 (N6931, N6930, N3131);
or OR4 (N6932, N6898, N3772, N2066, N344);
and AND3 (N6933, N6923, N4568, N2995);
or OR2 (N6934, N6922, N5356);
or OR2 (N6935, N6927, N4214);
and AND3 (N6936, N6935, N5950, N1573);
or OR3 (N6937, N6929, N2355, N160);
and AND3 (N6938, N6932, N6827, N6224);
not NOT1 (N6939, N6933);
buf BUF1 (N6940, N6934);
nand NAND3 (N6941, N6893, N1895, N1210);
not NOT1 (N6942, N6936);
xor XOR2 (N6943, N6931, N2114);
nor NOR3 (N6944, N6940, N3377, N3820);
xor XOR2 (N6945, N6943, N3200);
xor XOR2 (N6946, N6945, N5953);
or OR3 (N6947, N6942, N4387, N3697);
nand NAND4 (N6948, N6938, N2092, N3018, N1872);
nand NAND3 (N6949, N6912, N2687, N659);
or OR4 (N6950, N6941, N651, N4148, N6793);
xor XOR2 (N6951, N6947, N5741);
and AND3 (N6952, N6939, N5811, N2099);
xor XOR2 (N6953, N6952, N2358);
or OR3 (N6954, N6953, N1765, N2647);
not NOT1 (N6955, N6946);
or OR3 (N6956, N6955, N6768, N513);
nor NOR2 (N6957, N6956, N2720);
not NOT1 (N6958, N6949);
nor NOR3 (N6959, N6944, N6630, N4576);
buf BUF1 (N6960, N6928);
or OR3 (N6961, N6957, N1361, N4493);
xor XOR2 (N6962, N6954, N3707);
nand NAND2 (N6963, N6924, N1427);
not NOT1 (N6964, N6958);
and AND3 (N6965, N6962, N4185, N2973);
xor XOR2 (N6966, N6965, N1815);
and AND2 (N6967, N6959, N1365);
xor XOR2 (N6968, N6948, N2834);
buf BUF1 (N6969, N6950);
nand NAND2 (N6970, N6961, N2766);
buf BUF1 (N6971, N6963);
nor NOR2 (N6972, N6969, N4104);
buf BUF1 (N6973, N6960);
or OR3 (N6974, N6966, N1353, N1419);
xor XOR2 (N6975, N6937, N1555);
buf BUF1 (N6976, N6973);
and AND2 (N6977, N6964, N551);
buf BUF1 (N6978, N6967);
not NOT1 (N6979, N6978);
buf BUF1 (N6980, N6974);
buf BUF1 (N6981, N6972);
not NOT1 (N6982, N6977);
and AND3 (N6983, N6975, N2639, N1522);
buf BUF1 (N6984, N6968);
or OR2 (N6985, N6976, N6242);
xor XOR2 (N6986, N6984, N3638);
or OR3 (N6987, N6986, N255, N4517);
nor NOR4 (N6988, N6979, N1852, N4775, N3213);
nand NAND4 (N6989, N6983, N283, N4453, N2444);
nor NOR4 (N6990, N6987, N2620, N3682, N2411);
buf BUF1 (N6991, N6982);
and AND3 (N6992, N6989, N6714, N3553);
nor NOR4 (N6993, N6981, N6279, N5788, N6480);
nand NAND3 (N6994, N6985, N4615, N1334);
buf BUF1 (N6995, N6951);
and AND3 (N6996, N6971, N6232, N437);
nor NOR3 (N6997, N6988, N6851, N912);
buf BUF1 (N6998, N6993);
xor XOR2 (N6999, N6996, N3588);
or OR2 (N7000, N6992, N6192);
not NOT1 (N7001, N6994);
and AND3 (N7002, N6991, N103, N3618);
nor NOR4 (N7003, N6990, N6132, N3101, N4865);
nand NAND3 (N7004, N6980, N6399, N4606);
nor NOR3 (N7005, N7002, N4232, N78);
nand NAND4 (N7006, N7005, N468, N5682, N6278);
not NOT1 (N7007, N7006);
nand NAND3 (N7008, N7003, N2825, N262);
nand NAND4 (N7009, N6998, N5814, N7008, N2230);
nor NOR2 (N7010, N3786, N1207);
or OR2 (N7011, N6997, N816);
nand NAND2 (N7012, N7011, N6871);
nor NOR2 (N7013, N6999, N1640);
xor XOR2 (N7014, N7007, N2133);
buf BUF1 (N7015, N6970);
buf BUF1 (N7016, N7001);
and AND4 (N7017, N7012, N6993, N5733, N2311);
buf BUF1 (N7018, N7013);
xor XOR2 (N7019, N7018, N930);
nor NOR4 (N7020, N7010, N6464, N5151, N2515);
or OR3 (N7021, N7009, N5254, N3526);
xor XOR2 (N7022, N7020, N1029);
or OR2 (N7023, N7004, N3371);
nor NOR3 (N7024, N7023, N3448, N5359);
nor NOR4 (N7025, N7000, N592, N530, N1958);
or OR4 (N7026, N7017, N137, N1827, N985);
nor NOR3 (N7027, N7025, N3769, N1562);
or OR3 (N7028, N6995, N1353, N5245);
xor XOR2 (N7029, N7027, N5810);
and AND3 (N7030, N7019, N4457, N3291);
buf BUF1 (N7031, N7021);
not NOT1 (N7032, N7028);
xor XOR2 (N7033, N7015, N1339);
not NOT1 (N7034, N7016);
buf BUF1 (N7035, N7024);
xor XOR2 (N7036, N7034, N5487);
not NOT1 (N7037, N7026);
nor NOR2 (N7038, N7036, N141);
not NOT1 (N7039, N7035);
nand NAND4 (N7040, N7029, N3048, N450, N4622);
nand NAND4 (N7041, N7038, N5774, N3807, N5336);
nand NAND2 (N7042, N7031, N2547);
or OR2 (N7043, N7030, N6321);
nand NAND4 (N7044, N7039, N5007, N4484, N4548);
or OR3 (N7045, N7037, N3133, N6298);
nor NOR3 (N7046, N7045, N1876, N6348);
nor NOR2 (N7047, N7044, N6680);
or OR3 (N7048, N7041, N5410, N1027);
nor NOR2 (N7049, N7047, N4747);
buf BUF1 (N7050, N7022);
buf BUF1 (N7051, N7042);
buf BUF1 (N7052, N7014);
and AND2 (N7053, N7033, N1170);
and AND4 (N7054, N7050, N2863, N4997, N1504);
nand NAND3 (N7055, N7043, N5318, N2298);
buf BUF1 (N7056, N7046);
nor NOR3 (N7057, N7049, N1854, N6288);
and AND3 (N7058, N7054, N1890, N1654);
buf BUF1 (N7059, N7058);
nor NOR4 (N7060, N7055, N5369, N5603, N6986);
buf BUF1 (N7061, N7040);
not NOT1 (N7062, N7060);
not NOT1 (N7063, N7059);
nand NAND4 (N7064, N7053, N5443, N3338, N4128);
and AND3 (N7065, N7032, N1721, N4332);
or OR4 (N7066, N7051, N353, N2228, N3762);
nand NAND3 (N7067, N7062, N1137, N5941);
nand NAND2 (N7068, N7064, N189);
and AND2 (N7069, N7066, N3813);
and AND3 (N7070, N7069, N711, N4298);
or OR3 (N7071, N7061, N4945, N6095);
xor XOR2 (N7072, N7065, N3089);
or OR2 (N7073, N7071, N1933);
and AND2 (N7074, N7073, N3974);
not NOT1 (N7075, N7052);
buf BUF1 (N7076, N7067);
or OR3 (N7077, N7075, N4851, N3606);
and AND4 (N7078, N7077, N3787, N5788, N1966);
xor XOR2 (N7079, N7076, N3071);
not NOT1 (N7080, N7072);
nor NOR4 (N7081, N7074, N4964, N4890, N1217);
buf BUF1 (N7082, N7079);
or OR2 (N7083, N7048, N3066);
xor XOR2 (N7084, N7080, N59);
buf BUF1 (N7085, N7081);
nand NAND2 (N7086, N7063, N2419);
buf BUF1 (N7087, N7056);
nor NOR2 (N7088, N7084, N1230);
and AND3 (N7089, N7068, N2314, N2487);
not NOT1 (N7090, N7083);
buf BUF1 (N7091, N7086);
and AND3 (N7092, N7082, N1304, N5796);
and AND3 (N7093, N7089, N252, N3620);
nand NAND3 (N7094, N7087, N2993, N1892);
nand NAND2 (N7095, N7092, N14);
buf BUF1 (N7096, N7070);
buf BUF1 (N7097, N7095);
and AND4 (N7098, N7091, N4356, N5686, N1397);
or OR2 (N7099, N7093, N6041);
and AND3 (N7100, N7099, N2618, N3995);
buf BUF1 (N7101, N7094);
xor XOR2 (N7102, N7101, N4970);
xor XOR2 (N7103, N7097, N2978);
buf BUF1 (N7104, N7090);
nor NOR2 (N7105, N7104, N5015);
nand NAND2 (N7106, N7100, N4101);
not NOT1 (N7107, N7096);
and AND2 (N7108, N7103, N4284);
xor XOR2 (N7109, N7105, N6542);
nor NOR4 (N7110, N7109, N1227, N4382, N2519);
xor XOR2 (N7111, N7108, N1620);
nor NOR2 (N7112, N7057, N5190);
and AND4 (N7113, N7088, N3489, N77, N5564);
or OR2 (N7114, N7113, N853);
nor NOR3 (N7115, N7098, N5099, N1674);
nor NOR3 (N7116, N7114, N6654, N5041);
and AND4 (N7117, N7106, N5847, N1130, N3906);
nor NOR2 (N7118, N7117, N6367);
not NOT1 (N7119, N7110);
or OR2 (N7120, N7111, N725);
and AND4 (N7121, N7116, N5917, N4096, N866);
and AND2 (N7122, N7120, N4517);
nor NOR2 (N7123, N7119, N2143);
and AND3 (N7124, N7122, N4776, N4234);
and AND2 (N7125, N7102, N5166);
nand NAND2 (N7126, N7115, N2929);
nor NOR4 (N7127, N7085, N2023, N4401, N4949);
nor NOR2 (N7128, N7121, N1070);
not NOT1 (N7129, N7125);
not NOT1 (N7130, N7107);
or OR4 (N7131, N7129, N5789, N988, N1244);
buf BUF1 (N7132, N7112);
or OR2 (N7133, N7130, N4061);
or OR3 (N7134, N7127, N708, N5792);
buf BUF1 (N7135, N7118);
or OR3 (N7136, N7126, N5697, N424);
buf BUF1 (N7137, N7134);
nor NOR3 (N7138, N7136, N6363, N5445);
xor XOR2 (N7139, N7123, N3170);
buf BUF1 (N7140, N7128);
buf BUF1 (N7141, N7132);
not NOT1 (N7142, N7124);
nor NOR2 (N7143, N7131, N4527);
and AND2 (N7144, N7137, N378);
and AND3 (N7145, N7138, N240, N5239);
buf BUF1 (N7146, N7139);
and AND3 (N7147, N7143, N4571, N3546);
buf BUF1 (N7148, N7140);
not NOT1 (N7149, N7146);
and AND3 (N7150, N7144, N6789, N4716);
nor NOR2 (N7151, N7149, N3194);
nand NAND2 (N7152, N7147, N6343);
not NOT1 (N7153, N7151);
and AND4 (N7154, N7133, N6087, N6638, N3629);
buf BUF1 (N7155, N7154);
and AND3 (N7156, N7155, N4485, N809);
and AND2 (N7157, N7148, N5029);
buf BUF1 (N7158, N7150);
and AND3 (N7159, N7153, N5574, N5777);
buf BUF1 (N7160, N7142);
not NOT1 (N7161, N7135);
nor NOR2 (N7162, N7158, N6089);
or OR4 (N7163, N7078, N2977, N2157, N6152);
not NOT1 (N7164, N7157);
or OR3 (N7165, N7159, N1679, N2374);
or OR4 (N7166, N7156, N3552, N843, N2636);
nand NAND2 (N7167, N7145, N6396);
nor NOR3 (N7168, N7162, N4821, N4312);
or OR2 (N7169, N7163, N5122);
or OR3 (N7170, N7152, N4743, N5609);
or OR2 (N7171, N7164, N6870);
xor XOR2 (N7172, N7165, N2956);
or OR3 (N7173, N7141, N6658, N5801);
not NOT1 (N7174, N7161);
nand NAND3 (N7175, N7168, N3690, N38);
xor XOR2 (N7176, N7170, N1677);
not NOT1 (N7177, N7171);
buf BUF1 (N7178, N7177);
xor XOR2 (N7179, N7172, N5275);
buf BUF1 (N7180, N7169);
nor NOR4 (N7181, N7178, N3309, N2003, N1952);
nor NOR3 (N7182, N7180, N4221, N7104);
nor NOR4 (N7183, N7181, N705, N6719, N5909);
and AND4 (N7184, N7183, N5850, N2128, N5546);
xor XOR2 (N7185, N7166, N2867);
buf BUF1 (N7186, N7184);
nor NOR4 (N7187, N7182, N3583, N268, N2787);
buf BUF1 (N7188, N7174);
buf BUF1 (N7189, N7173);
not NOT1 (N7190, N7179);
xor XOR2 (N7191, N7188, N357);
buf BUF1 (N7192, N7186);
not NOT1 (N7193, N7185);
and AND4 (N7194, N7190, N7170, N127, N3930);
or OR2 (N7195, N7191, N3471);
not NOT1 (N7196, N7189);
and AND4 (N7197, N7195, N6340, N2139, N4698);
nor NOR4 (N7198, N7192, N4443, N4834, N5265);
xor XOR2 (N7199, N7194, N750);
xor XOR2 (N7200, N7199, N5369);
nor NOR2 (N7201, N7197, N5859);
nand NAND2 (N7202, N7201, N6684);
nand NAND4 (N7203, N7200, N1240, N7132, N397);
nand NAND2 (N7204, N7160, N3982);
buf BUF1 (N7205, N7203);
buf BUF1 (N7206, N7198);
xor XOR2 (N7207, N7175, N5709);
and AND4 (N7208, N7196, N477, N3555, N3928);
not NOT1 (N7209, N7206);
xor XOR2 (N7210, N7202, N326);
or OR4 (N7211, N7205, N6300, N6345, N5554);
xor XOR2 (N7212, N7167, N6590);
nand NAND4 (N7213, N7187, N6529, N3354, N5739);
nor NOR2 (N7214, N7210, N205);
nand NAND3 (N7215, N7209, N3015, N5118);
and AND3 (N7216, N7193, N45, N2154);
or OR2 (N7217, N7214, N4205);
nand NAND3 (N7218, N7213, N4783, N1971);
or OR2 (N7219, N7218, N5207);
not NOT1 (N7220, N7204);
and AND4 (N7221, N7176, N2661, N4508, N2382);
not NOT1 (N7222, N7220);
not NOT1 (N7223, N7211);
and AND4 (N7224, N7219, N2212, N4356, N2739);
not NOT1 (N7225, N7208);
and AND3 (N7226, N7217, N6534, N3049);
nand NAND3 (N7227, N7224, N6368, N711);
and AND4 (N7228, N7223, N2816, N5958, N37);
nor NOR4 (N7229, N7226, N3670, N180, N5015);
or OR3 (N7230, N7215, N6649, N449);
or OR4 (N7231, N7225, N1797, N7197, N1290);
and AND3 (N7232, N7221, N5865, N2552);
xor XOR2 (N7233, N7222, N268);
buf BUF1 (N7234, N7233);
nand NAND2 (N7235, N7234, N3976);
xor XOR2 (N7236, N7207, N952);
and AND3 (N7237, N7230, N2692, N4678);
nor NOR3 (N7238, N7228, N4144, N973);
and AND3 (N7239, N7216, N1721, N3992);
nand NAND4 (N7240, N7231, N6521, N1626, N2131);
xor XOR2 (N7241, N7212, N1690);
nand NAND3 (N7242, N7232, N363, N4032);
buf BUF1 (N7243, N7235);
buf BUF1 (N7244, N7241);
not NOT1 (N7245, N7239);
not NOT1 (N7246, N7243);
nor NOR4 (N7247, N7240, N2596, N4457, N53);
and AND4 (N7248, N7237, N2204, N5627, N6103);
and AND3 (N7249, N7247, N6412, N2196);
not NOT1 (N7250, N7249);
not NOT1 (N7251, N7245);
xor XOR2 (N7252, N7242, N3556);
xor XOR2 (N7253, N7248, N2683);
nand NAND2 (N7254, N7238, N4943);
buf BUF1 (N7255, N7251);
nor NOR2 (N7256, N7227, N5425);
and AND4 (N7257, N7255, N6491, N1002, N257);
buf BUF1 (N7258, N7229);
xor XOR2 (N7259, N7256, N5012);
xor XOR2 (N7260, N7252, N7150);
not NOT1 (N7261, N7253);
not NOT1 (N7262, N7261);
nand NAND2 (N7263, N7260, N1475);
nor NOR3 (N7264, N7257, N6508, N5916);
buf BUF1 (N7265, N7259);
or OR4 (N7266, N7265, N669, N3014, N5032);
and AND2 (N7267, N7266, N816);
and AND2 (N7268, N7236, N2741);
nor NOR4 (N7269, N7268, N4295, N2632, N6109);
nor NOR2 (N7270, N7244, N2445);
buf BUF1 (N7271, N7258);
nor NOR4 (N7272, N7270, N5040, N3652, N6103);
buf BUF1 (N7273, N7264);
and AND2 (N7274, N7267, N5072);
buf BUF1 (N7275, N7271);
and AND2 (N7276, N7254, N1327);
xor XOR2 (N7277, N7246, N3314);
nor NOR2 (N7278, N7275, N6141);
buf BUF1 (N7279, N7250);
nor NOR4 (N7280, N7279, N4647, N6805, N2693);
xor XOR2 (N7281, N7262, N2769);
nor NOR3 (N7282, N7277, N3385, N6400);
nand NAND3 (N7283, N7278, N5789, N6914);
nor NOR3 (N7284, N7281, N6303, N3480);
nand NAND4 (N7285, N7274, N3795, N4723, N7101);
buf BUF1 (N7286, N7280);
nor NOR3 (N7287, N7285, N1224, N2779);
and AND2 (N7288, N7269, N6622);
nor NOR3 (N7289, N7287, N4902, N787);
buf BUF1 (N7290, N7283);
buf BUF1 (N7291, N7272);
or OR4 (N7292, N7286, N1640, N6086, N2408);
buf BUF1 (N7293, N7291);
or OR3 (N7294, N7263, N2645, N6859);
nor NOR4 (N7295, N7292, N2560, N6696, N4004);
buf BUF1 (N7296, N7288);
or OR3 (N7297, N7290, N6861, N6003);
and AND3 (N7298, N7276, N3054, N5785);
nand NAND2 (N7299, N7284, N5151);
buf BUF1 (N7300, N7295);
or OR2 (N7301, N7289, N2713);
not NOT1 (N7302, N7299);
nor NOR2 (N7303, N7302, N466);
buf BUF1 (N7304, N7296);
nor NOR2 (N7305, N7273, N2919);
nand NAND3 (N7306, N7293, N7184, N3682);
nand NAND4 (N7307, N7298, N1197, N6678, N2922);
or OR2 (N7308, N7282, N6899);
and AND2 (N7309, N7307, N1198);
and AND4 (N7310, N7308, N5557, N4366, N460);
xor XOR2 (N7311, N7297, N5095);
and AND2 (N7312, N7310, N1222);
buf BUF1 (N7313, N7304);
buf BUF1 (N7314, N7305);
and AND4 (N7315, N7311, N616, N488, N1439);
nor NOR3 (N7316, N7306, N5183, N712);
not NOT1 (N7317, N7314);
xor XOR2 (N7318, N7317, N7248);
and AND2 (N7319, N7312, N2431);
or OR3 (N7320, N7300, N4376, N3022);
nand NAND2 (N7321, N7303, N1968);
nor NOR3 (N7322, N7320, N598, N5285);
not NOT1 (N7323, N7321);
nand NAND2 (N7324, N7316, N3007);
buf BUF1 (N7325, N7322);
nor NOR4 (N7326, N7318, N1423, N2996, N5280);
nand NAND4 (N7327, N7326, N2572, N4941, N5255);
and AND4 (N7328, N7294, N5888, N2730, N3197);
not NOT1 (N7329, N7327);
buf BUF1 (N7330, N7313);
nor NOR2 (N7331, N7330, N6605);
and AND4 (N7332, N7309, N3786, N6558, N3874);
xor XOR2 (N7333, N7315, N1989);
nand NAND3 (N7334, N7332, N4905, N3250);
nand NAND2 (N7335, N7329, N1456);
or OR4 (N7336, N7334, N2624, N1487, N5431);
buf BUF1 (N7337, N7301);
not NOT1 (N7338, N7324);
buf BUF1 (N7339, N7333);
buf BUF1 (N7340, N7335);
and AND3 (N7341, N7336, N7270, N3040);
and AND3 (N7342, N7328, N1250, N3553);
buf BUF1 (N7343, N7323);
nor NOR3 (N7344, N7325, N6150, N1040);
and AND4 (N7345, N7344, N3881, N2354, N4160);
nor NOR4 (N7346, N7342, N223, N1522, N5016);
and AND3 (N7347, N7346, N4604, N5992);
nand NAND2 (N7348, N7338, N2723);
not NOT1 (N7349, N7319);
buf BUF1 (N7350, N7341);
nor NOR2 (N7351, N7348, N5181);
xor XOR2 (N7352, N7350, N4735);
not NOT1 (N7353, N7337);
nor NOR3 (N7354, N7351, N1485, N4821);
nor NOR3 (N7355, N7339, N1395, N3881);
xor XOR2 (N7356, N7343, N4789);
not NOT1 (N7357, N7352);
xor XOR2 (N7358, N7357, N582);
xor XOR2 (N7359, N7353, N6588);
and AND3 (N7360, N7345, N7342, N6664);
not NOT1 (N7361, N7331);
nand NAND4 (N7362, N7349, N2193, N470, N2356);
and AND4 (N7363, N7347, N2182, N826, N4470);
not NOT1 (N7364, N7361);
buf BUF1 (N7365, N7340);
nand NAND2 (N7366, N7356, N1210);
and AND4 (N7367, N7358, N346, N6393, N5183);
buf BUF1 (N7368, N7367);
nand NAND4 (N7369, N7363, N91, N1098, N3801);
nand NAND4 (N7370, N7366, N1232, N6890, N2891);
nor NOR4 (N7371, N7354, N1472, N6511, N3330);
or OR3 (N7372, N7355, N4615, N2710);
not NOT1 (N7373, N7368);
and AND4 (N7374, N7371, N7218, N2154, N6636);
and AND4 (N7375, N7369, N1334, N5766, N2080);
not NOT1 (N7376, N7364);
nor NOR2 (N7377, N7370, N4178);
or OR4 (N7378, N7375, N2337, N1712, N2114);
or OR2 (N7379, N7377, N364);
buf BUF1 (N7380, N7362);
nor NOR2 (N7381, N7380, N6402);
buf BUF1 (N7382, N7372);
xor XOR2 (N7383, N7382, N3753);
xor XOR2 (N7384, N7383, N6400);
xor XOR2 (N7385, N7360, N4389);
nand NAND2 (N7386, N7385, N3133);
buf BUF1 (N7387, N7376);
xor XOR2 (N7388, N7384, N609);
nor NOR4 (N7389, N7374, N6212, N6459, N6197);
and AND3 (N7390, N7359, N5002, N4231);
nand NAND2 (N7391, N7373, N261);
nor NOR3 (N7392, N7389, N1231, N5031);
and AND4 (N7393, N7392, N897, N6539, N3937);
not NOT1 (N7394, N7381);
nand NAND2 (N7395, N7393, N4738);
xor XOR2 (N7396, N7394, N3521);
nor NOR3 (N7397, N7378, N3349, N1168);
and AND3 (N7398, N7365, N3881, N626);
and AND4 (N7399, N7396, N94, N3016, N2069);
buf BUF1 (N7400, N7388);
not NOT1 (N7401, N7397);
buf BUF1 (N7402, N7386);
nand NAND2 (N7403, N7402, N4735);
or OR4 (N7404, N7400, N3374, N5251, N5658);
nand NAND2 (N7405, N7403, N7393);
nor NOR2 (N7406, N7405, N23);
or OR2 (N7407, N7391, N2653);
nand NAND4 (N7408, N7399, N2904, N754, N2298);
or OR4 (N7409, N7395, N2070, N1085, N5290);
not NOT1 (N7410, N7387);
nand NAND4 (N7411, N7401, N3036, N7391, N7296);
nor NOR4 (N7412, N7406, N241, N1509, N3405);
nand NAND2 (N7413, N7408, N3765);
nor NOR4 (N7414, N7398, N2516, N1013, N2015);
not NOT1 (N7415, N7390);
nand NAND2 (N7416, N7415, N7098);
not NOT1 (N7417, N7411);
nor NOR3 (N7418, N7414, N4770, N231);
xor XOR2 (N7419, N7409, N4247);
or OR4 (N7420, N7404, N5772, N5949, N4737);
nand NAND2 (N7421, N7413, N6044);
or OR3 (N7422, N7412, N7395, N3131);
not NOT1 (N7423, N7418);
buf BUF1 (N7424, N7422);
nand NAND2 (N7425, N7407, N6475);
buf BUF1 (N7426, N7423);
and AND3 (N7427, N7379, N1472, N6758);
not NOT1 (N7428, N7417);
xor XOR2 (N7429, N7427, N6020);
nor NOR3 (N7430, N7428, N2145, N1893);
not NOT1 (N7431, N7416);
nor NOR2 (N7432, N7420, N5804);
buf BUF1 (N7433, N7432);
buf BUF1 (N7434, N7424);
and AND3 (N7435, N7426, N3605, N2630);
or OR3 (N7436, N7419, N5614, N2661);
and AND4 (N7437, N7434, N3961, N6084, N2957);
xor XOR2 (N7438, N7425, N3155);
nor NOR2 (N7439, N7421, N5125);
xor XOR2 (N7440, N7433, N6489);
buf BUF1 (N7441, N7439);
xor XOR2 (N7442, N7410, N2543);
not NOT1 (N7443, N7429);
not NOT1 (N7444, N7437);
xor XOR2 (N7445, N7444, N3327);
and AND2 (N7446, N7440, N3692);
nor NOR3 (N7447, N7435, N3782, N430);
buf BUF1 (N7448, N7441);
xor XOR2 (N7449, N7448, N66);
not NOT1 (N7450, N7438);
not NOT1 (N7451, N7443);
nor NOR2 (N7452, N7447, N4454);
nand NAND3 (N7453, N7446, N773, N513);
nand NAND2 (N7454, N7449, N6625);
and AND3 (N7455, N7442, N1749, N3534);
nor NOR3 (N7456, N7445, N3267, N1697);
not NOT1 (N7457, N7453);
nand NAND4 (N7458, N7452, N210, N5015, N1629);
nand NAND2 (N7459, N7458, N4159);
xor XOR2 (N7460, N7456, N5470);
nor NOR4 (N7461, N7430, N2041, N1817, N5865);
not NOT1 (N7462, N7451);
not NOT1 (N7463, N7455);
nand NAND4 (N7464, N7462, N4406, N3013, N4380);
nor NOR3 (N7465, N7461, N696, N5833);
not NOT1 (N7466, N7464);
not NOT1 (N7467, N7463);
nand NAND4 (N7468, N7466, N2831, N6732, N5478);
nor NOR3 (N7469, N7468, N2178, N5254);
not NOT1 (N7470, N7467);
nor NOR4 (N7471, N7469, N4912, N5935, N6146);
nand NAND4 (N7472, N7450, N5970, N5756, N4724);
and AND3 (N7473, N7460, N342, N5613);
buf BUF1 (N7474, N7431);
and AND4 (N7475, N7459, N6549, N1743, N3215);
nor NOR2 (N7476, N7454, N1279);
not NOT1 (N7477, N7465);
nor NOR4 (N7478, N7476, N5986, N4555, N6504);
and AND4 (N7479, N7472, N4190, N7354, N7082);
buf BUF1 (N7480, N7477);
buf BUF1 (N7481, N7436);
nand NAND3 (N7482, N7473, N4191, N7424);
nand NAND2 (N7483, N7457, N2234);
nor NOR4 (N7484, N7471, N579, N6978, N3853);
nand NAND4 (N7485, N7479, N2765, N3624, N6347);
and AND3 (N7486, N7470, N7435, N6538);
or OR3 (N7487, N7484, N5544, N3971);
nand NAND4 (N7488, N7483, N3279, N675, N1296);
buf BUF1 (N7489, N7487);
nor NOR2 (N7490, N7485, N2738);
nand NAND2 (N7491, N7482, N4965);
or OR3 (N7492, N7488, N5574, N7228);
and AND3 (N7493, N7478, N4577, N5220);
or OR3 (N7494, N7474, N3072, N2607);
nor NOR2 (N7495, N7481, N6337);
xor XOR2 (N7496, N7490, N5344);
or OR2 (N7497, N7489, N1153);
xor XOR2 (N7498, N7492, N5051);
or OR3 (N7499, N7493, N444, N1235);
nor NOR4 (N7500, N7486, N1589, N6477, N4225);
not NOT1 (N7501, N7475);
nor NOR4 (N7502, N7491, N1516, N1276, N3610);
or OR2 (N7503, N7497, N3818);
xor XOR2 (N7504, N7499, N3182);
nor NOR3 (N7505, N7501, N6398, N5553);
not NOT1 (N7506, N7498);
or OR3 (N7507, N7506, N1426, N5426);
nand NAND4 (N7508, N7500, N3169, N3860, N2666);
or OR4 (N7509, N7507, N6485, N714, N6810);
buf BUF1 (N7510, N7480);
buf BUF1 (N7511, N7509);
and AND3 (N7512, N7505, N4478, N169);
not NOT1 (N7513, N7508);
nor NOR2 (N7514, N7512, N5413);
xor XOR2 (N7515, N7514, N3503);
not NOT1 (N7516, N7494);
not NOT1 (N7517, N7516);
and AND4 (N7518, N7517, N5032, N6015, N559);
not NOT1 (N7519, N7515);
nor NOR3 (N7520, N7511, N6091, N5227);
buf BUF1 (N7521, N7513);
not NOT1 (N7522, N7518);
or OR4 (N7523, N7504, N6321, N190, N2080);
not NOT1 (N7524, N7496);
or OR4 (N7525, N7503, N7500, N5566, N6278);
and AND3 (N7526, N7519, N6609, N1529);
or OR2 (N7527, N7521, N2802);
not NOT1 (N7528, N7502);
nand NAND3 (N7529, N7495, N2043, N3410);
not NOT1 (N7530, N7510);
not NOT1 (N7531, N7523);
and AND4 (N7532, N7525, N1539, N4540, N2674);
nand NAND3 (N7533, N7522, N6098, N5910);
and AND4 (N7534, N7520, N3318, N3360, N4107);
xor XOR2 (N7535, N7526, N6283);
nand NAND4 (N7536, N7532, N466, N7166, N2881);
and AND3 (N7537, N7527, N3524, N1552);
and AND4 (N7538, N7536, N5074, N1195, N3305);
or OR2 (N7539, N7535, N3519);
buf BUF1 (N7540, N7534);
xor XOR2 (N7541, N7533, N729);
nand NAND2 (N7542, N7537, N156);
nand NAND3 (N7543, N7529, N4493, N4744);
xor XOR2 (N7544, N7528, N4359);
nand NAND3 (N7545, N7541, N2796, N7391);
or OR3 (N7546, N7544, N1466, N910);
buf BUF1 (N7547, N7524);
nand NAND2 (N7548, N7547, N2100);
or OR3 (N7549, N7542, N7026, N4653);
nor NOR3 (N7550, N7549, N5331, N3720);
not NOT1 (N7551, N7545);
nor NOR4 (N7552, N7538, N4035, N5471, N6767);
xor XOR2 (N7553, N7539, N4959);
nor NOR3 (N7554, N7550, N5586, N535);
buf BUF1 (N7555, N7554);
buf BUF1 (N7556, N7551);
and AND4 (N7557, N7548, N5706, N6851, N2888);
nor NOR4 (N7558, N7546, N2038, N1315, N5100);
nand NAND2 (N7559, N7553, N2977);
nand NAND4 (N7560, N7552, N2103, N149, N4482);
and AND3 (N7561, N7557, N7453, N4759);
xor XOR2 (N7562, N7559, N3996);
nor NOR4 (N7563, N7531, N3517, N3115, N4982);
nor NOR2 (N7564, N7556, N1460);
or OR4 (N7565, N7561, N6773, N4548, N532);
and AND2 (N7566, N7558, N5610);
and AND3 (N7567, N7564, N2251, N2829);
nand NAND2 (N7568, N7563, N2677);
buf BUF1 (N7569, N7565);
or OR2 (N7570, N7567, N6360);
xor XOR2 (N7571, N7555, N6093);
buf BUF1 (N7572, N7530);
xor XOR2 (N7573, N7572, N5031);
nor NOR3 (N7574, N7568, N381, N3601);
or OR4 (N7575, N7570, N2158, N6283, N990);
nand NAND2 (N7576, N7569, N3077);
nor NOR4 (N7577, N7575, N2638, N2568, N4070);
nor NOR4 (N7578, N7566, N609, N3486, N271);
buf BUF1 (N7579, N7562);
and AND3 (N7580, N7577, N1924, N2329);
xor XOR2 (N7581, N7540, N5080);
buf BUF1 (N7582, N7579);
not NOT1 (N7583, N7576);
and AND4 (N7584, N7578, N192, N2820, N2696);
or OR4 (N7585, N7583, N2140, N2602, N2608);
xor XOR2 (N7586, N7571, N5127);
or OR4 (N7587, N7573, N2351, N6228, N5215);
nand NAND3 (N7588, N7574, N3002, N6547);
or OR3 (N7589, N7585, N7519, N5003);
xor XOR2 (N7590, N7586, N6933);
or OR3 (N7591, N7582, N6661, N703);
nand NAND3 (N7592, N7580, N2306, N2199);
and AND3 (N7593, N7589, N144, N3119);
not NOT1 (N7594, N7592);
nor NOR3 (N7595, N7588, N4602, N7307);
xor XOR2 (N7596, N7590, N2536);
not NOT1 (N7597, N7591);
or OR2 (N7598, N7597, N6062);
not NOT1 (N7599, N7581);
and AND2 (N7600, N7560, N108);
xor XOR2 (N7601, N7593, N3820);
not NOT1 (N7602, N7594);
xor XOR2 (N7603, N7600, N1335);
or OR3 (N7604, N7603, N3190, N110);
not NOT1 (N7605, N7587);
not NOT1 (N7606, N7604);
and AND2 (N7607, N7596, N1940);
xor XOR2 (N7608, N7606, N3384);
and AND4 (N7609, N7608, N4941, N5728, N1882);
not NOT1 (N7610, N7609);
and AND3 (N7611, N7543, N4958, N1828);
not NOT1 (N7612, N7598);
nor NOR3 (N7613, N7610, N6485, N1381);
nand NAND3 (N7614, N7611, N6080, N4022);
xor XOR2 (N7615, N7601, N6836);
or OR2 (N7616, N7612, N2467);
and AND4 (N7617, N7602, N4592, N1074, N2785);
buf BUF1 (N7618, N7599);
xor XOR2 (N7619, N7615, N799);
and AND3 (N7620, N7595, N3206, N6553);
xor XOR2 (N7621, N7619, N5146);
and AND2 (N7622, N7617, N1826);
nand NAND4 (N7623, N7618, N5861, N458, N483);
xor XOR2 (N7624, N7613, N3510);
not NOT1 (N7625, N7621);
xor XOR2 (N7626, N7624, N5952);
or OR4 (N7627, N7626, N4219, N433, N5362);
xor XOR2 (N7628, N7622, N5311);
xor XOR2 (N7629, N7614, N6070);
xor XOR2 (N7630, N7605, N5072);
and AND4 (N7631, N7584, N2220, N2747, N3805);
nor NOR2 (N7632, N7627, N7313);
or OR3 (N7633, N7616, N5583, N5011);
or OR3 (N7634, N7633, N7605, N2204);
or OR4 (N7635, N7631, N4245, N3017, N5446);
or OR2 (N7636, N7625, N4262);
and AND2 (N7637, N7630, N4018);
or OR3 (N7638, N7635, N2932, N2300);
nand NAND2 (N7639, N7636, N6741);
and AND2 (N7640, N7639, N6551);
or OR4 (N7641, N7634, N5916, N4296, N5342);
and AND4 (N7642, N7637, N2663, N2345, N4763);
nand NAND2 (N7643, N7628, N1790);
xor XOR2 (N7644, N7623, N4191);
nand NAND2 (N7645, N7644, N6285);
nor NOR2 (N7646, N7642, N4446);
xor XOR2 (N7647, N7629, N2738);
xor XOR2 (N7648, N7643, N7185);
nor NOR4 (N7649, N7648, N1082, N4547, N5668);
or OR4 (N7650, N7641, N5254, N1439, N6074);
nor NOR3 (N7651, N7647, N1571, N4943);
and AND4 (N7652, N7645, N466, N838, N3310);
not NOT1 (N7653, N7652);
nor NOR2 (N7654, N7632, N5378);
xor XOR2 (N7655, N7638, N5440);
buf BUF1 (N7656, N7620);
and AND4 (N7657, N7649, N4652, N2035, N5863);
buf BUF1 (N7658, N7655);
nor NOR4 (N7659, N7653, N932, N5845, N6576);
or OR2 (N7660, N7607, N3199);
nor NOR2 (N7661, N7660, N7510);
nor NOR2 (N7662, N7656, N1145);
not NOT1 (N7663, N7662);
xor XOR2 (N7664, N7658, N6113);
and AND3 (N7665, N7657, N5798, N5649);
nor NOR2 (N7666, N7661, N3718);
xor XOR2 (N7667, N7651, N2534);
or OR4 (N7668, N7666, N4489, N3553, N715);
buf BUF1 (N7669, N7640);
buf BUF1 (N7670, N7646);
not NOT1 (N7671, N7664);
and AND4 (N7672, N7654, N414, N367, N4600);
not NOT1 (N7673, N7650);
or OR3 (N7674, N7663, N6637, N4632);
nor NOR3 (N7675, N7667, N2713, N5580);
buf BUF1 (N7676, N7674);
not NOT1 (N7677, N7672);
xor XOR2 (N7678, N7675, N3073);
xor XOR2 (N7679, N7668, N4649);
buf BUF1 (N7680, N7669);
or OR2 (N7681, N7673, N6192);
and AND2 (N7682, N7670, N6487);
not NOT1 (N7683, N7682);
nor NOR4 (N7684, N7665, N3892, N5545, N2493);
and AND2 (N7685, N7659, N1311);
nor NOR4 (N7686, N7671, N7095, N5791, N2463);
nor NOR3 (N7687, N7678, N1255, N6073);
and AND3 (N7688, N7681, N453, N4767);
buf BUF1 (N7689, N7688);
and AND4 (N7690, N7679, N2478, N4789, N4771);
and AND4 (N7691, N7680, N4018, N766, N4175);
and AND4 (N7692, N7676, N2141, N2784, N946);
nor NOR2 (N7693, N7687, N2317);
nand NAND2 (N7694, N7683, N6184);
nor NOR4 (N7695, N7691, N1575, N4439, N6864);
nor NOR2 (N7696, N7695, N1378);
buf BUF1 (N7697, N7690);
xor XOR2 (N7698, N7692, N4349);
or OR4 (N7699, N7698, N5244, N3196, N2208);
or OR3 (N7700, N7699, N1455, N5872);
and AND4 (N7701, N7700, N2945, N6351, N3291);
nor NOR4 (N7702, N7685, N559, N7408, N4668);
and AND2 (N7703, N7684, N3009);
or OR2 (N7704, N7686, N2907);
nand NAND4 (N7705, N7703, N212, N2727, N5780);
not NOT1 (N7706, N7689);
nand NAND3 (N7707, N7693, N7396, N5845);
or OR4 (N7708, N7704, N2695, N5296, N2931);
and AND2 (N7709, N7707, N4840);
buf BUF1 (N7710, N7706);
not NOT1 (N7711, N7677);
or OR3 (N7712, N7710, N7604, N3298);
nand NAND3 (N7713, N7702, N5278, N3950);
not NOT1 (N7714, N7708);
nor NOR3 (N7715, N7713, N2447, N6556);
or OR4 (N7716, N7715, N2796, N4359, N3055);
buf BUF1 (N7717, N7716);
nor NOR3 (N7718, N7696, N2525, N359);
xor XOR2 (N7719, N7709, N5282);
not NOT1 (N7720, N7714);
not NOT1 (N7721, N7711);
nand NAND4 (N7722, N7712, N2163, N7495, N2637);
xor XOR2 (N7723, N7718, N7148);
or OR3 (N7724, N7723, N1956, N7397);
or OR3 (N7725, N7720, N4908, N376);
or OR4 (N7726, N7724, N5928, N2168, N537);
nand NAND4 (N7727, N7725, N500, N5269, N2916);
not NOT1 (N7728, N7717);
nor NOR2 (N7729, N7694, N5629);
xor XOR2 (N7730, N7726, N4147);
not NOT1 (N7731, N7727);
nor NOR3 (N7732, N7730, N6447, N7017);
nand NAND3 (N7733, N7728, N3133, N5966);
and AND4 (N7734, N7731, N4303, N4503, N777);
nand NAND3 (N7735, N7734, N1043, N5699);
not NOT1 (N7736, N7732);
and AND3 (N7737, N7705, N6871, N5813);
nor NOR3 (N7738, N7737, N1531, N1237);
nand NAND3 (N7739, N7721, N2260, N3665);
xor XOR2 (N7740, N7738, N6369);
or OR3 (N7741, N7733, N6388, N1612);
nand NAND2 (N7742, N7736, N3277);
xor XOR2 (N7743, N7739, N3134);
and AND3 (N7744, N7740, N487, N5932);
and AND4 (N7745, N7701, N6518, N5819, N3211);
nor NOR2 (N7746, N7719, N3747);
buf BUF1 (N7747, N7742);
and AND4 (N7748, N7741, N2504, N7154, N934);
buf BUF1 (N7749, N7748);
or OR4 (N7750, N7744, N3637, N628, N819);
xor XOR2 (N7751, N7729, N6494);
buf BUF1 (N7752, N7697);
and AND4 (N7753, N7749, N1892, N6904, N3216);
nor NOR2 (N7754, N7743, N3526);
nor NOR3 (N7755, N7746, N7317, N3753);
or OR4 (N7756, N7747, N1954, N6119, N7590);
buf BUF1 (N7757, N7752);
not NOT1 (N7758, N7751);
xor XOR2 (N7759, N7745, N5298);
not NOT1 (N7760, N7758);
and AND2 (N7761, N7755, N2283);
or OR4 (N7762, N7761, N4876, N6369, N111);
nor NOR4 (N7763, N7756, N7325, N7200, N7099);
nand NAND4 (N7764, N7722, N7468, N1936, N1961);
and AND2 (N7765, N7764, N4470);
or OR4 (N7766, N7754, N1519, N1023, N2964);
or OR2 (N7767, N7762, N2501);
buf BUF1 (N7768, N7766);
nor NOR3 (N7769, N7757, N4097, N5321);
or OR2 (N7770, N7760, N228);
and AND4 (N7771, N7750, N1456, N6478, N6513);
xor XOR2 (N7772, N7765, N2754);
or OR4 (N7773, N7753, N7401, N6797, N1990);
not NOT1 (N7774, N7763);
or OR3 (N7775, N7769, N5504, N3322);
nand NAND3 (N7776, N7770, N4933, N720);
buf BUF1 (N7777, N7768);
nor NOR3 (N7778, N7771, N7727, N6768);
or OR3 (N7779, N7773, N356, N5408);
nand NAND4 (N7780, N7767, N168, N5297, N1566);
nand NAND4 (N7781, N7776, N1592, N4539, N5643);
buf BUF1 (N7782, N7774);
buf BUF1 (N7783, N7772);
xor XOR2 (N7784, N7779, N5689);
and AND4 (N7785, N7778, N2606, N5444, N6880);
or OR4 (N7786, N7735, N539, N5628, N2865);
xor XOR2 (N7787, N7780, N1690);
or OR4 (N7788, N7782, N6088, N4311, N4494);
nor NOR2 (N7789, N7788, N2922);
buf BUF1 (N7790, N7783);
or OR2 (N7791, N7790, N2930);
nor NOR2 (N7792, N7785, N563);
nand NAND3 (N7793, N7786, N3749, N2081);
or OR2 (N7794, N7775, N6944);
buf BUF1 (N7795, N7777);
and AND3 (N7796, N7784, N6651, N3568);
nand NAND4 (N7797, N7796, N5660, N1884, N6015);
nand NAND4 (N7798, N7795, N358, N2647, N240);
or OR2 (N7799, N7781, N4277);
and AND4 (N7800, N7787, N826, N2054, N2573);
or OR4 (N7801, N7791, N9, N1210, N3083);
or OR4 (N7802, N7759, N2109, N294, N7028);
and AND4 (N7803, N7792, N3482, N7524, N443);
not NOT1 (N7804, N7793);
not NOT1 (N7805, N7797);
nand NAND4 (N7806, N7798, N3921, N5970, N5117);
not NOT1 (N7807, N7806);
buf BUF1 (N7808, N7789);
buf BUF1 (N7809, N7803);
nor NOR4 (N7810, N7799, N1065, N2965, N5634);
nand NAND3 (N7811, N7801, N5484, N2471);
buf BUF1 (N7812, N7804);
not NOT1 (N7813, N7812);
nand NAND4 (N7814, N7811, N4909, N3080, N424);
nand NAND3 (N7815, N7814, N1356, N2091);
xor XOR2 (N7816, N7808, N1375);
not NOT1 (N7817, N7800);
or OR2 (N7818, N7813, N6650);
nand NAND2 (N7819, N7807, N1158);
not NOT1 (N7820, N7805);
xor XOR2 (N7821, N7819, N1394);
not NOT1 (N7822, N7821);
and AND3 (N7823, N7802, N6157, N6179);
nand NAND3 (N7824, N7822, N2537, N3846);
buf BUF1 (N7825, N7810);
and AND3 (N7826, N7820, N1010, N7680);
nor NOR3 (N7827, N7815, N6326, N6006);
nor NOR4 (N7828, N7823, N2081, N495, N4078);
xor XOR2 (N7829, N7827, N2192);
buf BUF1 (N7830, N7826);
nand NAND4 (N7831, N7824, N7222, N5813, N2749);
nor NOR3 (N7832, N7825, N843, N5597);
and AND2 (N7833, N7794, N5671);
or OR4 (N7834, N7833, N4702, N4244, N1489);
nor NOR4 (N7835, N7831, N4581, N455, N6759);
nor NOR2 (N7836, N7835, N5621);
not NOT1 (N7837, N7816);
buf BUF1 (N7838, N7837);
nor NOR4 (N7839, N7834, N7794, N5292, N7702);
xor XOR2 (N7840, N7828, N1915);
or OR3 (N7841, N7832, N4351, N4412);
nand NAND2 (N7842, N7838, N2808);
not NOT1 (N7843, N7840);
nand NAND4 (N7844, N7842, N2315, N3541, N859);
nand NAND3 (N7845, N7817, N2862, N5574);
not NOT1 (N7846, N7839);
not NOT1 (N7847, N7818);
buf BUF1 (N7848, N7841);
or OR2 (N7849, N7847, N6117);
not NOT1 (N7850, N7829);
xor XOR2 (N7851, N7846, N4886);
buf BUF1 (N7852, N7851);
or OR2 (N7853, N7852, N5366);
or OR4 (N7854, N7830, N1771, N3898, N4631);
and AND3 (N7855, N7809, N1255, N5929);
buf BUF1 (N7856, N7855);
or OR3 (N7857, N7853, N1473, N2015);
xor XOR2 (N7858, N7848, N5886);
xor XOR2 (N7859, N7844, N4922);
nand NAND3 (N7860, N7849, N5875, N2886);
not NOT1 (N7861, N7858);
buf BUF1 (N7862, N7845);
or OR3 (N7863, N7857, N3434, N6042);
not NOT1 (N7864, N7850);
nor NOR3 (N7865, N7854, N2805, N3364);
not NOT1 (N7866, N7864);
and AND4 (N7867, N7866, N5593, N7455, N3490);
buf BUF1 (N7868, N7843);
or OR2 (N7869, N7836, N1794);
nor NOR4 (N7870, N7860, N4400, N3608, N6311);
and AND3 (N7871, N7868, N591, N1673);
nor NOR4 (N7872, N7871, N7236, N5580, N271);
or OR4 (N7873, N7869, N104, N5899, N2912);
or OR4 (N7874, N7867, N7247, N2284, N3578);
not NOT1 (N7875, N7865);
or OR4 (N7876, N7872, N2728, N816, N2119);
nand NAND3 (N7877, N7873, N1303, N1740);
nor NOR2 (N7878, N7861, N7841);
nor NOR3 (N7879, N7876, N5750, N2140);
and AND3 (N7880, N7870, N5679, N1043);
nand NAND3 (N7881, N7863, N4716, N2328);
and AND4 (N7882, N7874, N3095, N3672, N3915);
not NOT1 (N7883, N7877);
nor NOR4 (N7884, N7879, N3609, N4543, N3826);
nand NAND3 (N7885, N7859, N5180, N4941);
nor NOR2 (N7886, N7882, N5986);
buf BUF1 (N7887, N7884);
nor NOR4 (N7888, N7875, N1045, N1168, N2045);
nor NOR4 (N7889, N7888, N7770, N4499, N2208);
and AND3 (N7890, N7883, N6313, N2350);
nor NOR3 (N7891, N7856, N5512, N458);
and AND4 (N7892, N7862, N5192, N2666, N5456);
and AND4 (N7893, N7890, N3352, N6183, N2080);
or OR3 (N7894, N7891, N737, N2287);
and AND3 (N7895, N7881, N752, N2164);
nor NOR2 (N7896, N7887, N7744);
not NOT1 (N7897, N7896);
nor NOR2 (N7898, N7885, N1819);
buf BUF1 (N7899, N7889);
or OR3 (N7900, N7880, N6264, N3795);
or OR3 (N7901, N7899, N4709, N3207);
not NOT1 (N7902, N7894);
buf BUF1 (N7903, N7898);
buf BUF1 (N7904, N7892);
and AND2 (N7905, N7900, N4042);
xor XOR2 (N7906, N7903, N649);
not NOT1 (N7907, N7904);
buf BUF1 (N7908, N7886);
and AND3 (N7909, N7905, N6434, N7519);
or OR3 (N7910, N7895, N1245, N3704);
not NOT1 (N7911, N7907);
and AND4 (N7912, N7902, N5835, N5653, N3139);
and AND2 (N7913, N7908, N859);
xor XOR2 (N7914, N7910, N6631);
nor NOR3 (N7915, N7911, N2582, N5406);
not NOT1 (N7916, N7913);
not NOT1 (N7917, N7878);
not NOT1 (N7918, N7901);
xor XOR2 (N7919, N7917, N4146);
or OR2 (N7920, N7916, N4489);
not NOT1 (N7921, N7914);
nand NAND4 (N7922, N7921, N6988, N373, N7342);
or OR3 (N7923, N7920, N3184, N69);
nor NOR4 (N7924, N7906, N1527, N2980, N1697);
xor XOR2 (N7925, N7924, N3519);
and AND4 (N7926, N7919, N5330, N4975, N2339);
xor XOR2 (N7927, N7915, N5270);
or OR3 (N7928, N7923, N4700, N1298);
or OR2 (N7929, N7922, N7792);
not NOT1 (N7930, N7926);
and AND2 (N7931, N7930, N520);
buf BUF1 (N7932, N7918);
or OR3 (N7933, N7897, N2248, N559);
nand NAND4 (N7934, N7932, N2969, N5319, N1852);
nand NAND4 (N7935, N7912, N2395, N5455, N2046);
nor NOR3 (N7936, N7928, N6975, N6178);
or OR2 (N7937, N7909, N224);
buf BUF1 (N7938, N7929);
nand NAND3 (N7939, N7936, N7034, N5269);
and AND4 (N7940, N7931, N4504, N1513, N6002);
and AND4 (N7941, N7935, N2907, N3118, N4016);
not NOT1 (N7942, N7933);
and AND4 (N7943, N7925, N932, N4116, N1310);
and AND4 (N7944, N7927, N6173, N3165, N236);
not NOT1 (N7945, N7893);
or OR2 (N7946, N7940, N5498);
or OR3 (N7947, N7939, N6434, N352);
xor XOR2 (N7948, N7938, N6345);
nor NOR3 (N7949, N7943, N2072, N5261);
nor NOR2 (N7950, N7946, N1199);
buf BUF1 (N7951, N7950);
xor XOR2 (N7952, N7942, N1444);
not NOT1 (N7953, N7934);
nor NOR4 (N7954, N7948, N6845, N7023, N3027);
nand NAND4 (N7955, N7952, N3160, N3950, N6169);
or OR4 (N7956, N7951, N5653, N135, N7230);
nor NOR2 (N7957, N7944, N2935);
not NOT1 (N7958, N7947);
or OR4 (N7959, N7937, N3888, N2325, N3276);
nor NOR2 (N7960, N7954, N3182);
nor NOR4 (N7961, N7949, N258, N1127, N3220);
and AND2 (N7962, N7941, N241);
not NOT1 (N7963, N7960);
xor XOR2 (N7964, N7959, N3171);
buf BUF1 (N7965, N7953);
nand NAND4 (N7966, N7956, N1952, N3213, N5963);
and AND4 (N7967, N7964, N4794, N5169, N5274);
and AND2 (N7968, N7958, N4801);
not NOT1 (N7969, N7945);
nor NOR4 (N7970, N7969, N7111, N690, N7346);
or OR2 (N7971, N7961, N2126);
buf BUF1 (N7972, N7965);
and AND4 (N7973, N7962, N6193, N3562, N5185);
xor XOR2 (N7974, N7955, N5719);
buf BUF1 (N7975, N7974);
buf BUF1 (N7976, N7966);
nor NOR4 (N7977, N7972, N3547, N3744, N5457);
and AND4 (N7978, N7976, N5101, N7791, N7210);
and AND3 (N7979, N7967, N4876, N930);
and AND3 (N7980, N7975, N6280, N7072);
or OR3 (N7981, N7963, N1900, N5810);
or OR3 (N7982, N7973, N6714, N2059);
nand NAND3 (N7983, N7982, N380, N4171);
and AND3 (N7984, N7983, N5225, N1518);
nor NOR3 (N7985, N7971, N932, N211);
not NOT1 (N7986, N7980);
not NOT1 (N7987, N7984);
xor XOR2 (N7988, N7978, N5220);
or OR2 (N7989, N7979, N5528);
buf BUF1 (N7990, N7987);
nor NOR3 (N7991, N7988, N1210, N3947);
not NOT1 (N7992, N7986);
nand NAND3 (N7993, N7989, N4307, N4784);
xor XOR2 (N7994, N7970, N410);
and AND3 (N7995, N7985, N768, N5190);
nand NAND3 (N7996, N7995, N1726, N2185);
buf BUF1 (N7997, N7992);
not NOT1 (N7998, N7990);
nor NOR3 (N7999, N7994, N2139, N7856);
and AND4 (N8000, N7968, N1059, N7543, N5318);
not NOT1 (N8001, N7981);
or OR2 (N8002, N7977, N7345);
xor XOR2 (N8003, N8001, N2926);
nand NAND3 (N8004, N7997, N2130, N5208);
or OR3 (N8005, N7991, N4152, N2876);
not NOT1 (N8006, N7957);
nand NAND4 (N8007, N8000, N7998, N7917, N6010);
not NOT1 (N8008, N3129);
not NOT1 (N8009, N8007);
not NOT1 (N8010, N7999);
and AND3 (N8011, N8010, N3717, N2218);
nor NOR3 (N8012, N7996, N5243, N6454);
buf BUF1 (N8013, N8004);
nand NAND4 (N8014, N8013, N5369, N1619, N5398);
and AND2 (N8015, N8008, N424);
buf BUF1 (N8016, N8009);
nor NOR3 (N8017, N8015, N4105, N1477);
or OR3 (N8018, N8014, N5530, N2518);
nor NOR3 (N8019, N8017, N239, N2712);
buf BUF1 (N8020, N8002);
nor NOR4 (N8021, N8019, N7805, N7048, N5052);
not NOT1 (N8022, N8021);
nor NOR3 (N8023, N8022, N5987, N2408);
nand NAND2 (N8024, N8005, N5909);
nor NOR3 (N8025, N8016, N5527, N1249);
nor NOR4 (N8026, N8011, N2869, N6078, N3438);
not NOT1 (N8027, N8026);
nand NAND3 (N8028, N8003, N891, N2263);
not NOT1 (N8029, N8024);
and AND2 (N8030, N8027, N3689);
and AND2 (N8031, N8018, N2581);
and AND4 (N8032, N8006, N7686, N5557, N3564);
nand NAND3 (N8033, N8020, N4638, N8006);
nor NOR2 (N8034, N8029, N5969);
not NOT1 (N8035, N7993);
nor NOR3 (N8036, N8012, N5892, N850);
not NOT1 (N8037, N8028);
xor XOR2 (N8038, N8032, N5963);
xor XOR2 (N8039, N8034, N6354);
nor NOR2 (N8040, N8035, N1891);
xor XOR2 (N8041, N8036, N1274);
xor XOR2 (N8042, N8037, N3472);
buf BUF1 (N8043, N8040);
not NOT1 (N8044, N8043);
xor XOR2 (N8045, N8023, N513);
buf BUF1 (N8046, N8031);
nor NOR3 (N8047, N8039, N1009, N6673);
nand NAND3 (N8048, N8025, N2432, N7380);
nand NAND2 (N8049, N8044, N60);
nand NAND3 (N8050, N8030, N4, N7450);
xor XOR2 (N8051, N8046, N1465);
not NOT1 (N8052, N8042);
and AND2 (N8053, N8050, N137);
nand NAND3 (N8054, N8045, N6601, N5002);
nand NAND3 (N8055, N8033, N1721, N4767);
nand NAND2 (N8056, N8049, N7107);
nor NOR2 (N8057, N8052, N1153);
or OR4 (N8058, N8038, N6437, N6295, N6394);
buf BUF1 (N8059, N8048);
nand NAND4 (N8060, N8057, N4259, N4219, N1835);
nor NOR2 (N8061, N8059, N3733);
or OR4 (N8062, N8055, N5550, N1033, N6153);
nand NAND4 (N8063, N8047, N1935, N4734, N5263);
buf BUF1 (N8064, N8053);
not NOT1 (N8065, N8060);
and AND2 (N8066, N8061, N2138);
not NOT1 (N8067, N8065);
and AND4 (N8068, N8066, N1712, N1617, N6210);
nand NAND3 (N8069, N8058, N1829, N551);
nor NOR2 (N8070, N8062, N3951);
buf BUF1 (N8071, N8064);
buf BUF1 (N8072, N8071);
not NOT1 (N8073, N8054);
xor XOR2 (N8074, N8063, N3178);
not NOT1 (N8075, N8069);
and AND3 (N8076, N8068, N387, N4739);
nand NAND3 (N8077, N8056, N7822, N1920);
nor NOR4 (N8078, N8077, N1645, N3907, N783);
nand NAND2 (N8079, N8072, N295);
and AND2 (N8080, N8051, N2909);
not NOT1 (N8081, N8078);
not NOT1 (N8082, N8075);
buf BUF1 (N8083, N8076);
nand NAND2 (N8084, N8082, N1664);
nor NOR4 (N8085, N8041, N8071, N4211, N4279);
not NOT1 (N8086, N8084);
nand NAND4 (N8087, N8081, N2959, N7097, N4429);
nor NOR2 (N8088, N8087, N1305);
nor NOR2 (N8089, N8086, N3477);
nor NOR4 (N8090, N8085, N3074, N3284, N4071);
nand NAND2 (N8091, N8073, N5510);
nor NOR2 (N8092, N8088, N849);
or OR3 (N8093, N8089, N6472, N4656);
xor XOR2 (N8094, N8067, N3516);
not NOT1 (N8095, N8079);
or OR3 (N8096, N8095, N2302, N3071);
xor XOR2 (N8097, N8083, N858);
xor XOR2 (N8098, N8094, N3771);
nor NOR3 (N8099, N8098, N3971, N4269);
and AND3 (N8100, N8080, N70, N2389);
buf BUF1 (N8101, N8070);
not NOT1 (N8102, N8099);
or OR3 (N8103, N8100, N336, N627);
nor NOR2 (N8104, N8092, N5308);
not NOT1 (N8105, N8101);
buf BUF1 (N8106, N8096);
xor XOR2 (N8107, N8103, N4774);
not NOT1 (N8108, N8074);
not NOT1 (N8109, N8106);
or OR4 (N8110, N8093, N2294, N6793, N3101);
nor NOR2 (N8111, N8108, N5112);
xor XOR2 (N8112, N8097, N4104);
or OR2 (N8113, N8112, N617);
and AND4 (N8114, N8110, N7634, N2433, N6332);
and AND2 (N8115, N8102, N2216);
and AND3 (N8116, N8090, N3941, N1515);
nand NAND4 (N8117, N8114, N142, N2171, N6668);
not NOT1 (N8118, N8117);
not NOT1 (N8119, N8113);
xor XOR2 (N8120, N8104, N7659);
nor NOR2 (N8121, N8107, N2549);
nor NOR4 (N8122, N8109, N3002, N923, N1646);
and AND4 (N8123, N8091, N4668, N2765, N4427);
not NOT1 (N8124, N8116);
xor XOR2 (N8125, N8105, N7118);
xor XOR2 (N8126, N8119, N6756);
buf BUF1 (N8127, N8121);
not NOT1 (N8128, N8126);
nor NOR3 (N8129, N8125, N2780, N1965);
xor XOR2 (N8130, N8124, N5751);
xor XOR2 (N8131, N8120, N3714);
nor NOR4 (N8132, N8129, N620, N4619, N2239);
not NOT1 (N8133, N8131);
not NOT1 (N8134, N8118);
or OR4 (N8135, N8111, N5131, N4031, N6867);
nor NOR4 (N8136, N8128, N1816, N5031, N5740);
xor XOR2 (N8137, N8123, N8071);
nor NOR3 (N8138, N8135, N5649, N978);
nand NAND2 (N8139, N8130, N3493);
nor NOR3 (N8140, N8132, N6482, N6773);
and AND3 (N8141, N8138, N4647, N3326);
nor NOR2 (N8142, N8136, N6272);
or OR2 (N8143, N8134, N7455);
xor XOR2 (N8144, N8142, N2952);
and AND2 (N8145, N8137, N5761);
and AND3 (N8146, N8133, N6671, N226);
buf BUF1 (N8147, N8141);
not NOT1 (N8148, N8143);
buf BUF1 (N8149, N8139);
nor NOR3 (N8150, N8144, N7351, N5777);
xor XOR2 (N8151, N8146, N3100);
buf BUF1 (N8152, N8147);
nor NOR4 (N8153, N8122, N4479, N7131, N5935);
nand NAND4 (N8154, N8145, N3773, N4880, N5924);
or OR2 (N8155, N8149, N3829);
nor NOR2 (N8156, N8150, N6116);
nor NOR3 (N8157, N8148, N4936, N225);
nand NAND3 (N8158, N8153, N4840, N1977);
not NOT1 (N8159, N8115);
nand NAND3 (N8160, N8157, N5296, N3632);
not NOT1 (N8161, N8151);
and AND3 (N8162, N8152, N5881, N7617);
nor NOR4 (N8163, N8159, N4902, N4504, N3976);
nor NOR2 (N8164, N8155, N6696);
nand NAND3 (N8165, N8127, N6592, N6560);
xor XOR2 (N8166, N8160, N3037);
xor XOR2 (N8167, N8166, N1402);
nor NOR2 (N8168, N8165, N1399);
buf BUF1 (N8169, N8158);
nor NOR3 (N8170, N8167, N7310, N49);
not NOT1 (N8171, N8156);
buf BUF1 (N8172, N8169);
nand NAND2 (N8173, N8161, N719);
buf BUF1 (N8174, N8140);
xor XOR2 (N8175, N8162, N3131);
buf BUF1 (N8176, N8163);
buf BUF1 (N8177, N8171);
or OR4 (N8178, N8154, N5211, N5905, N1699);
nor NOR3 (N8179, N8175, N5023, N2621);
buf BUF1 (N8180, N8168);
buf BUF1 (N8181, N8173);
xor XOR2 (N8182, N8164, N982);
buf BUF1 (N8183, N8172);
not NOT1 (N8184, N8179);
nand NAND4 (N8185, N8174, N6792, N3515, N7500);
nor NOR3 (N8186, N8183, N2615, N176);
not NOT1 (N8187, N8182);
xor XOR2 (N8188, N8170, N3232);
nand NAND3 (N8189, N8185, N2849, N3980);
buf BUF1 (N8190, N8189);
not NOT1 (N8191, N8176);
or OR3 (N8192, N8184, N3837, N4670);
buf BUF1 (N8193, N8178);
buf BUF1 (N8194, N8190);
or OR3 (N8195, N8188, N5818, N5562);
buf BUF1 (N8196, N8192);
xor XOR2 (N8197, N8196, N1080);
and AND4 (N8198, N8187, N1161, N1619, N4295);
or OR2 (N8199, N8180, N4095);
nand NAND4 (N8200, N8193, N6813, N3517, N6422);
nand NAND4 (N8201, N8195, N2725, N3556, N7400);
and AND4 (N8202, N8186, N4558, N4509, N2653);
nor NOR2 (N8203, N8191, N5494);
buf BUF1 (N8204, N8198);
and AND4 (N8205, N8202, N4158, N4989, N681);
xor XOR2 (N8206, N8204, N2564);
xor XOR2 (N8207, N8197, N2219);
and AND4 (N8208, N8205, N2963, N414, N6139);
nor NOR2 (N8209, N8194, N1419);
nand NAND3 (N8210, N8203, N2930, N4141);
or OR4 (N8211, N8199, N4164, N88, N5231);
xor XOR2 (N8212, N8209, N4235);
buf BUF1 (N8213, N8181);
not NOT1 (N8214, N8200);
not NOT1 (N8215, N8207);
nor NOR4 (N8216, N8213, N7636, N5735, N4565);
or OR4 (N8217, N8210, N6229, N1486, N6390);
buf BUF1 (N8218, N8211);
nor NOR3 (N8219, N8217, N3021, N3715);
or OR3 (N8220, N8218, N7682, N4482);
or OR3 (N8221, N8201, N1832, N3493);
nand NAND2 (N8222, N8206, N3834);
buf BUF1 (N8223, N8216);
xor XOR2 (N8224, N8221, N1615);
xor XOR2 (N8225, N8215, N4561);
not NOT1 (N8226, N8225);
nor NOR2 (N8227, N8220, N7950);
not NOT1 (N8228, N8214);
nor NOR3 (N8229, N8212, N7405, N7949);
and AND3 (N8230, N8229, N4846, N8070);
xor XOR2 (N8231, N8177, N4631);
nand NAND2 (N8232, N8228, N5329);
buf BUF1 (N8233, N8227);
not NOT1 (N8234, N8223);
not NOT1 (N8235, N8208);
xor XOR2 (N8236, N8224, N6855);
xor XOR2 (N8237, N8234, N5500);
not NOT1 (N8238, N8232);
not NOT1 (N8239, N8219);
xor XOR2 (N8240, N8235, N7590);
nand NAND3 (N8241, N8236, N1167, N992);
nor NOR3 (N8242, N8240, N1606, N5773);
or OR4 (N8243, N8233, N6790, N6802, N8100);
xor XOR2 (N8244, N8239, N7508);
nor NOR3 (N8245, N8241, N6939, N5907);
and AND4 (N8246, N8226, N5185, N1658, N7304);
nand NAND4 (N8247, N8222, N637, N2652, N550);
and AND3 (N8248, N8230, N841, N4107);
or OR2 (N8249, N8242, N5996);
or OR2 (N8250, N8244, N6916);
buf BUF1 (N8251, N8249);
not NOT1 (N8252, N8251);
or OR4 (N8253, N8250, N1951, N2853, N5740);
nor NOR4 (N8254, N8247, N1513, N891, N2324);
and AND4 (N8255, N8245, N2933, N133, N6418);
nor NOR3 (N8256, N8254, N1252, N1382);
buf BUF1 (N8257, N8238);
xor XOR2 (N8258, N8231, N4202);
xor XOR2 (N8259, N8252, N2880);
and AND4 (N8260, N8243, N3498, N5447, N7429);
and AND3 (N8261, N8237, N3530, N3752);
xor XOR2 (N8262, N8255, N3013);
not NOT1 (N8263, N8257);
xor XOR2 (N8264, N8262, N1258);
buf BUF1 (N8265, N8264);
nand NAND3 (N8266, N8248, N5109, N4037);
xor XOR2 (N8267, N8258, N6983);
xor XOR2 (N8268, N8261, N7846);
buf BUF1 (N8269, N8265);
nor NOR2 (N8270, N8259, N4387);
not NOT1 (N8271, N8256);
or OR3 (N8272, N8268, N3400, N6001);
buf BUF1 (N8273, N8246);
not NOT1 (N8274, N8269);
xor XOR2 (N8275, N8266, N1813);
nand NAND4 (N8276, N8271, N1872, N2304, N1442);
and AND3 (N8277, N8272, N5059, N1184);
nand NAND3 (N8278, N8270, N7149, N906);
xor XOR2 (N8279, N8273, N7776);
nor NOR3 (N8280, N8263, N4329, N2822);
or OR2 (N8281, N8260, N6472);
nor NOR2 (N8282, N8281, N842);
or OR4 (N8283, N8267, N6205, N291, N4611);
nand NAND4 (N8284, N8276, N6851, N6693, N6519);
nand NAND3 (N8285, N8280, N4346, N4548);
xor XOR2 (N8286, N8279, N5348);
xor XOR2 (N8287, N8278, N4820);
not NOT1 (N8288, N8285);
buf BUF1 (N8289, N8283);
nand NAND4 (N8290, N8277, N7388, N7886, N7014);
not NOT1 (N8291, N8253);
not NOT1 (N8292, N8287);
and AND4 (N8293, N8292, N7151, N5678, N6966);
buf BUF1 (N8294, N8275);
buf BUF1 (N8295, N8291);
buf BUF1 (N8296, N8288);
not NOT1 (N8297, N8290);
nor NOR3 (N8298, N8284, N1048, N2739);
and AND4 (N8299, N8274, N5599, N7384, N1473);
buf BUF1 (N8300, N8286);
buf BUF1 (N8301, N8294);
nand NAND2 (N8302, N8299, N2566);
nor NOR4 (N8303, N8296, N7028, N3385, N2416);
not NOT1 (N8304, N8289);
or OR3 (N8305, N8282, N7574, N4398);
not NOT1 (N8306, N8300);
nor NOR4 (N8307, N8301, N3826, N7846, N5507);
nand NAND2 (N8308, N8307, N1212);
xor XOR2 (N8309, N8295, N2711);
nor NOR4 (N8310, N8303, N731, N6153, N5985);
buf BUF1 (N8311, N8309);
nand NAND3 (N8312, N8310, N4195, N1103);
nand NAND4 (N8313, N8311, N3020, N48, N6593);
nand NAND2 (N8314, N8305, N6581);
nor NOR3 (N8315, N8304, N419, N2622);
nor NOR4 (N8316, N8308, N991, N5605, N2751);
and AND4 (N8317, N8313, N1063, N4972, N1587);
and AND3 (N8318, N8302, N2171, N3960);
nor NOR3 (N8319, N8297, N4887, N8038);
and AND2 (N8320, N8314, N7918);
and AND4 (N8321, N8315, N2589, N3734, N1344);
buf BUF1 (N8322, N8312);
and AND4 (N8323, N8306, N7153, N2271, N5304);
and AND4 (N8324, N8318, N2238, N6665, N188);
xor XOR2 (N8325, N8323, N218);
or OR4 (N8326, N8293, N5977, N5554, N5490);
and AND3 (N8327, N8324, N1197, N663);
buf BUF1 (N8328, N8319);
not NOT1 (N8329, N8326);
not NOT1 (N8330, N8329);
or OR2 (N8331, N8330, N2708);
not NOT1 (N8332, N8331);
buf BUF1 (N8333, N8316);
and AND3 (N8334, N8333, N4968, N5987);
xor XOR2 (N8335, N8298, N7601);
not NOT1 (N8336, N8328);
xor XOR2 (N8337, N8332, N7265);
buf BUF1 (N8338, N8337);
or OR3 (N8339, N8327, N3965, N1061);
xor XOR2 (N8340, N8334, N3499);
not NOT1 (N8341, N8320);
or OR2 (N8342, N8339, N2733);
buf BUF1 (N8343, N8321);
buf BUF1 (N8344, N8325);
and AND3 (N8345, N8343, N6883, N5537);
nand NAND4 (N8346, N8336, N3028, N2370, N6044);
xor XOR2 (N8347, N8344, N3660);
not NOT1 (N8348, N8346);
buf BUF1 (N8349, N8322);
xor XOR2 (N8350, N8340, N5380);
nand NAND4 (N8351, N8335, N3574, N393, N3934);
nand NAND4 (N8352, N8349, N2516, N7616, N6520);
buf BUF1 (N8353, N8348);
and AND3 (N8354, N8350, N2967, N7797);
and AND3 (N8355, N8352, N901, N4635);
nor NOR3 (N8356, N8354, N2741, N291);
buf BUF1 (N8357, N8317);
nor NOR2 (N8358, N8341, N2282);
buf BUF1 (N8359, N8358);
nand NAND4 (N8360, N8351, N4433, N4349, N8335);
or OR2 (N8361, N8356, N3441);
nor NOR2 (N8362, N8361, N7957);
nand NAND2 (N8363, N8359, N1932);
and AND3 (N8364, N8342, N4907, N4045);
not NOT1 (N8365, N8345);
or OR4 (N8366, N8357, N1465, N3726, N7226);
nand NAND3 (N8367, N8347, N4936, N4105);
or OR4 (N8368, N8360, N422, N4184, N410);
nand NAND4 (N8369, N8363, N3989, N865, N4854);
or OR3 (N8370, N8365, N793, N2143);
or OR3 (N8371, N8366, N3487, N7748);
or OR2 (N8372, N8369, N5680);
xor XOR2 (N8373, N8370, N8037);
not NOT1 (N8374, N8367);
nor NOR3 (N8375, N8338, N466, N1572);
nor NOR4 (N8376, N8371, N544, N5882, N7831);
buf BUF1 (N8377, N8374);
or OR3 (N8378, N8375, N8308, N4106);
xor XOR2 (N8379, N8378, N2876);
not NOT1 (N8380, N8362);
nor NOR4 (N8381, N8377, N5469, N3451, N2970);
xor XOR2 (N8382, N8373, N6931);
not NOT1 (N8383, N8381);
and AND3 (N8384, N8364, N8164, N5181);
buf BUF1 (N8385, N8379);
nor NOR4 (N8386, N8368, N6194, N8181, N5371);
nor NOR4 (N8387, N8355, N6656, N2827, N7163);
not NOT1 (N8388, N8380);
and AND2 (N8389, N8383, N2171);
nor NOR4 (N8390, N8385, N718, N2694, N562);
nand NAND3 (N8391, N8353, N3528, N702);
not NOT1 (N8392, N8390);
and AND4 (N8393, N8389, N4845, N1064, N3106);
xor XOR2 (N8394, N8392, N2669);
not NOT1 (N8395, N8393);
and AND4 (N8396, N8384, N1812, N6101, N7170);
not NOT1 (N8397, N8387);
nand NAND2 (N8398, N8396, N8382);
not NOT1 (N8399, N4090);
buf BUF1 (N8400, N8372);
or OR4 (N8401, N8395, N6626, N3373, N3762);
nand NAND3 (N8402, N8399, N1768, N2381);
nor NOR4 (N8403, N8376, N2745, N7761, N6920);
or OR3 (N8404, N8403, N5622, N3877);
nand NAND3 (N8405, N8397, N3013, N7272);
buf BUF1 (N8406, N8388);
or OR2 (N8407, N8386, N3139);
buf BUF1 (N8408, N8391);
nand NAND2 (N8409, N8404, N8289);
nand NAND4 (N8410, N8402, N1641, N1987, N1088);
nor NOR3 (N8411, N8407, N5149, N4514);
and AND4 (N8412, N8408, N860, N4840, N2618);
or OR4 (N8413, N8412, N6217, N5737, N2983);
buf BUF1 (N8414, N8409);
xor XOR2 (N8415, N8401, N2891);
nand NAND2 (N8416, N8400, N3003);
nand NAND3 (N8417, N8414, N5867, N708);
not NOT1 (N8418, N8406);
or OR4 (N8419, N8415, N2647, N8370, N4372);
buf BUF1 (N8420, N8417);
xor XOR2 (N8421, N8398, N3249);
nor NOR3 (N8422, N8405, N7907, N3540);
and AND4 (N8423, N8421, N3010, N6443, N4349);
and AND4 (N8424, N8422, N7508, N6689, N939);
nand NAND2 (N8425, N8411, N5209);
and AND2 (N8426, N8419, N2256);
xor XOR2 (N8427, N8413, N1839);
and AND3 (N8428, N8425, N1615, N889);
not NOT1 (N8429, N8426);
nor NOR2 (N8430, N8420, N5489);
not NOT1 (N8431, N8423);
xor XOR2 (N8432, N8410, N1550);
or OR2 (N8433, N8432, N65);
buf BUF1 (N8434, N8433);
nor NOR4 (N8435, N8431, N6132, N5130, N1057);
or OR4 (N8436, N8430, N2022, N3082, N3468);
not NOT1 (N8437, N8418);
nor NOR4 (N8438, N8394, N1972, N3347, N4235);
xor XOR2 (N8439, N8436, N252);
and AND4 (N8440, N8416, N7134, N6902, N410);
nand NAND4 (N8441, N8427, N7408, N3425, N1810);
and AND4 (N8442, N8424, N6871, N3637, N8185);
or OR2 (N8443, N8428, N1140);
nor NOR3 (N8444, N8435, N3131, N6990);
xor XOR2 (N8445, N8442, N5573);
xor XOR2 (N8446, N8444, N3204);
not NOT1 (N8447, N8441);
xor XOR2 (N8448, N8446, N6714);
and AND3 (N8449, N8440, N5535, N6072);
nor NOR4 (N8450, N8437, N1723, N6491, N1916);
or OR2 (N8451, N8439, N5001);
xor XOR2 (N8452, N8445, N5095);
and AND2 (N8453, N8452, N132);
and AND2 (N8454, N8448, N4625);
and AND2 (N8455, N8429, N6820);
not NOT1 (N8456, N8453);
xor XOR2 (N8457, N8443, N3211);
nand NAND4 (N8458, N8456, N7698, N6488, N1861);
nand NAND4 (N8459, N8447, N4329, N1610, N8298);
nor NOR3 (N8460, N8459, N7546, N6459);
and AND4 (N8461, N8454, N4412, N3115, N6776);
not NOT1 (N8462, N8458);
or OR4 (N8463, N8462, N8374, N8037, N6772);
nor NOR4 (N8464, N8450, N5476, N3368, N5922);
not NOT1 (N8465, N8451);
nand NAND2 (N8466, N8460, N1195);
or OR2 (N8467, N8463, N4488);
and AND2 (N8468, N8455, N4947);
nand NAND4 (N8469, N8461, N8377, N6690, N4695);
xor XOR2 (N8470, N8465, N1256);
xor XOR2 (N8471, N8466, N1079);
xor XOR2 (N8472, N8457, N5345);
xor XOR2 (N8473, N8469, N3626);
or OR2 (N8474, N8473, N1822);
buf BUF1 (N8475, N8438);
or OR3 (N8476, N8449, N7602, N2933);
or OR3 (N8477, N8464, N5188, N7856);
not NOT1 (N8478, N8471);
and AND4 (N8479, N8470, N5608, N2650, N2868);
and AND3 (N8480, N8479, N6371, N7942);
or OR2 (N8481, N8467, N2646);
buf BUF1 (N8482, N8472);
and AND4 (N8483, N8482, N217, N1398, N7042);
or OR4 (N8484, N8468, N8068, N7978, N6824);
nand NAND3 (N8485, N8483, N8422, N5575);
nand NAND2 (N8486, N8480, N7793);
xor XOR2 (N8487, N8486, N2515);
and AND4 (N8488, N8477, N2769, N4234, N1336);
xor XOR2 (N8489, N8487, N445);
nand NAND2 (N8490, N8481, N613);
and AND3 (N8491, N8434, N7942, N7915);
buf BUF1 (N8492, N8488);
xor XOR2 (N8493, N8485, N4015);
nor NOR2 (N8494, N8478, N2773);
buf BUF1 (N8495, N8492);
nor NOR4 (N8496, N8489, N2350, N7733, N8337);
nor NOR3 (N8497, N8475, N3363, N5549);
or OR4 (N8498, N8491, N8279, N4665, N1542);
xor XOR2 (N8499, N8495, N2351);
and AND4 (N8500, N8499, N7241, N2951, N8025);
or OR2 (N8501, N8476, N7817);
buf BUF1 (N8502, N8484);
and AND4 (N8503, N8498, N6004, N8056, N3239);
xor XOR2 (N8504, N8503, N6716);
nand NAND4 (N8505, N8497, N6319, N2824, N4533);
and AND4 (N8506, N8500, N1856, N4245, N6128);
nor NOR4 (N8507, N8494, N4447, N6312, N4364);
or OR4 (N8508, N8506, N4442, N6335, N2781);
and AND4 (N8509, N8501, N558, N4577, N4037);
xor XOR2 (N8510, N8507, N8139);
nand NAND4 (N8511, N8504, N179, N5911, N3699);
xor XOR2 (N8512, N8490, N5821);
buf BUF1 (N8513, N8509);
or OR4 (N8514, N8496, N4443, N6122, N785);
nand NAND3 (N8515, N8505, N3994, N6322);
nand NAND4 (N8516, N8515, N5791, N90, N6430);
or OR4 (N8517, N8514, N571, N4575, N4455);
buf BUF1 (N8518, N8516);
and AND3 (N8519, N8518, N2032, N5409);
not NOT1 (N8520, N8512);
buf BUF1 (N8521, N8502);
buf BUF1 (N8522, N8493);
nor NOR2 (N8523, N8522, N3317);
buf BUF1 (N8524, N8474);
or OR2 (N8525, N8510, N3502);
not NOT1 (N8526, N8508);
and AND3 (N8527, N8520, N3538, N5793);
nor NOR2 (N8528, N8511, N1471);
or OR4 (N8529, N8525, N880, N8069, N6497);
buf BUF1 (N8530, N8517);
buf BUF1 (N8531, N8529);
not NOT1 (N8532, N8527);
nand NAND4 (N8533, N8513, N7767, N7527, N4396);
not NOT1 (N8534, N8519);
buf BUF1 (N8535, N8528);
not NOT1 (N8536, N8530);
or OR2 (N8537, N8526, N2715);
and AND4 (N8538, N8532, N542, N8141, N6814);
nor NOR3 (N8539, N8537, N3228, N3365);
xor XOR2 (N8540, N8533, N233);
or OR4 (N8541, N8538, N4152, N2979, N4465);
xor XOR2 (N8542, N8531, N790);
nand NAND4 (N8543, N8534, N1023, N6551, N2248);
buf BUF1 (N8544, N8521);
buf BUF1 (N8545, N8544);
nand NAND3 (N8546, N8524, N271, N6831);
nor NOR3 (N8547, N8539, N693, N3118);
and AND4 (N8548, N8535, N942, N3877, N7671);
and AND2 (N8549, N8545, N5930);
buf BUF1 (N8550, N8548);
not NOT1 (N8551, N8542);
nor NOR4 (N8552, N8549, N6284, N8056, N8008);
xor XOR2 (N8553, N8551, N6546);
or OR4 (N8554, N8541, N6870, N6397, N3259);
buf BUF1 (N8555, N8543);
and AND4 (N8556, N8555, N6429, N4636, N2198);
not NOT1 (N8557, N8547);
and AND4 (N8558, N8554, N6651, N1746, N8235);
and AND3 (N8559, N8552, N8064, N397);
or OR4 (N8560, N8559, N3936, N925, N7215);
buf BUF1 (N8561, N8540);
nand NAND2 (N8562, N8550, N769);
nand NAND2 (N8563, N8562, N6710);
nor NOR2 (N8564, N8563, N3296);
xor XOR2 (N8565, N8560, N7441);
not NOT1 (N8566, N8557);
not NOT1 (N8567, N8561);
nor NOR3 (N8568, N8558, N8300, N623);
nor NOR3 (N8569, N8536, N5861, N2344);
nand NAND3 (N8570, N8546, N4901, N3850);
and AND4 (N8571, N8565, N5354, N1465, N3355);
and AND3 (N8572, N8571, N5558, N4566);
and AND3 (N8573, N8556, N3875, N7006);
buf BUF1 (N8574, N8570);
xor XOR2 (N8575, N8568, N7286);
nor NOR2 (N8576, N8569, N5651);
and AND2 (N8577, N8566, N777);
buf BUF1 (N8578, N8523);
and AND2 (N8579, N8578, N2345);
xor XOR2 (N8580, N8579, N8239);
or OR3 (N8581, N8567, N957, N4681);
not NOT1 (N8582, N8573);
buf BUF1 (N8583, N8564);
nor NOR4 (N8584, N8580, N1958, N6203, N5036);
not NOT1 (N8585, N8577);
xor XOR2 (N8586, N8574, N860);
xor XOR2 (N8587, N8584, N7433);
or OR4 (N8588, N8581, N4664, N5063, N5018);
nor NOR4 (N8589, N8582, N434, N2747, N6283);
nor NOR2 (N8590, N8585, N4627);
or OR4 (N8591, N8589, N3820, N6134, N2478);
or OR3 (N8592, N8587, N8035, N2631);
buf BUF1 (N8593, N8576);
xor XOR2 (N8594, N8572, N23);
or OR3 (N8595, N8594, N2698, N5556);
nand NAND3 (N8596, N8591, N4846, N8375);
xor XOR2 (N8597, N8575, N2961);
xor XOR2 (N8598, N8595, N2488);
buf BUF1 (N8599, N8597);
nand NAND3 (N8600, N8553, N6852, N4815);
nand NAND2 (N8601, N8593, N1661);
nor NOR2 (N8602, N8600, N3553);
not NOT1 (N8603, N8586);
nor NOR3 (N8604, N8588, N8318, N3337);
not NOT1 (N8605, N8596);
and AND3 (N8606, N8605, N5073, N2803);
and AND2 (N8607, N8606, N7389);
or OR4 (N8608, N8604, N1401, N3259, N777);
nand NAND4 (N8609, N8590, N4088, N1183, N7728);
or OR2 (N8610, N8601, N3248);
buf BUF1 (N8611, N8609);
and AND3 (N8612, N8611, N5376, N4206);
xor XOR2 (N8613, N8599, N8311);
and AND3 (N8614, N8602, N1677, N1851);
not NOT1 (N8615, N8603);
nor NOR3 (N8616, N8607, N3341, N2718);
nor NOR4 (N8617, N8613, N5863, N5206, N2654);
and AND2 (N8618, N8617, N7509);
not NOT1 (N8619, N8598);
and AND3 (N8620, N8615, N1783, N5581);
or OR2 (N8621, N8608, N4233);
nor NOR2 (N8622, N8618, N6634);
nand NAND4 (N8623, N8614, N8455, N410, N5858);
nand NAND4 (N8624, N8592, N8103, N1181, N6728);
xor XOR2 (N8625, N8620, N965);
or OR3 (N8626, N8622, N4236, N1276);
nand NAND2 (N8627, N8616, N4504);
buf BUF1 (N8628, N8623);
or OR4 (N8629, N8627, N5220, N8157, N2950);
buf BUF1 (N8630, N8624);
not NOT1 (N8631, N8612);
buf BUF1 (N8632, N8625);
and AND4 (N8633, N8629, N8417, N6168, N2817);
buf BUF1 (N8634, N8619);
xor XOR2 (N8635, N8634, N2186);
nand NAND2 (N8636, N8628, N2039);
xor XOR2 (N8637, N8631, N1671);
or OR4 (N8638, N8636, N8157, N6135, N4100);
not NOT1 (N8639, N8635);
buf BUF1 (N8640, N8633);
not NOT1 (N8641, N8632);
or OR4 (N8642, N8621, N585, N6399, N2556);
buf BUF1 (N8643, N8638);
buf BUF1 (N8644, N8643);
and AND2 (N8645, N8644, N3216);
nor NOR3 (N8646, N8626, N1046, N2695);
or OR2 (N8647, N8637, N3409);
or OR2 (N8648, N8642, N450);
xor XOR2 (N8649, N8583, N7304);
not NOT1 (N8650, N8648);
or OR4 (N8651, N8641, N6660, N5354, N6150);
nor NOR2 (N8652, N8646, N6612);
and AND2 (N8653, N8610, N5238);
buf BUF1 (N8654, N8652);
not NOT1 (N8655, N8647);
or OR2 (N8656, N8651, N3493);
buf BUF1 (N8657, N8649);
or OR2 (N8658, N8630, N5906);
or OR4 (N8659, N8650, N5461, N8194, N2113);
and AND3 (N8660, N8658, N4099, N7262);
buf BUF1 (N8661, N8656);
not NOT1 (N8662, N8645);
or OR4 (N8663, N8655, N5272, N6022, N8400);
xor XOR2 (N8664, N8660, N4088);
nor NOR4 (N8665, N8640, N1945, N5974, N7420);
xor XOR2 (N8666, N8657, N6888);
or OR4 (N8667, N8659, N2904, N2137, N542);
nand NAND4 (N8668, N8664, N6201, N6265, N3364);
buf BUF1 (N8669, N8665);
buf BUF1 (N8670, N8639);
nand NAND4 (N8671, N8663, N244, N3923, N70);
nor NOR2 (N8672, N8654, N8028);
and AND2 (N8673, N8671, N2705);
or OR3 (N8674, N8666, N479, N1956);
nor NOR4 (N8675, N8674, N7363, N8243, N53);
nor NOR4 (N8676, N8668, N3252, N1107, N7634);
buf BUF1 (N8677, N8670);
and AND3 (N8678, N8661, N6462, N4674);
and AND3 (N8679, N8673, N7050, N7951);
or OR4 (N8680, N8662, N2978, N3605, N6642);
nand NAND3 (N8681, N8678, N8147, N3363);
nand NAND3 (N8682, N8681, N6195, N1828);
not NOT1 (N8683, N8680);
xor XOR2 (N8684, N8683, N7802);
xor XOR2 (N8685, N8684, N5705);
xor XOR2 (N8686, N8672, N3557);
buf BUF1 (N8687, N8669);
xor XOR2 (N8688, N8675, N4965);
buf BUF1 (N8689, N8679);
and AND4 (N8690, N8685, N5527, N988, N3642);
buf BUF1 (N8691, N8677);
nor NOR2 (N8692, N8688, N8199);
xor XOR2 (N8693, N8682, N4458);
not NOT1 (N8694, N8686);
nand NAND3 (N8695, N8667, N3317, N8618);
and AND3 (N8696, N8653, N8070, N7677);
and AND2 (N8697, N8691, N3208);
nand NAND4 (N8698, N8689, N5018, N6935, N943);
buf BUF1 (N8699, N8687);
nand NAND2 (N8700, N8696, N4414);
nor NOR3 (N8701, N8697, N6802, N905);
nand NAND4 (N8702, N8700, N8482, N7874, N1974);
buf BUF1 (N8703, N8690);
not NOT1 (N8704, N8703);
buf BUF1 (N8705, N8695);
nand NAND4 (N8706, N8692, N318, N3888, N6827);
and AND2 (N8707, N8694, N4134);
nor NOR3 (N8708, N8707, N4293, N4829);
and AND2 (N8709, N8706, N8620);
and AND3 (N8710, N8701, N4535, N1941);
buf BUF1 (N8711, N8709);
nor NOR3 (N8712, N8698, N5317, N5338);
nand NAND3 (N8713, N8711, N1893, N7502);
or OR2 (N8714, N8699, N7789);
buf BUF1 (N8715, N8676);
nand NAND2 (N8716, N8693, N4192);
or OR3 (N8717, N8716, N8126, N7815);
and AND2 (N8718, N8705, N7155);
nand NAND2 (N8719, N8712, N1861);
and AND2 (N8720, N8717, N4573);
nand NAND2 (N8721, N8714, N5006);
not NOT1 (N8722, N8702);
nand NAND3 (N8723, N8715, N2700, N4229);
or OR4 (N8724, N8723, N1412, N6762, N7718);
or OR3 (N8725, N8722, N2594, N1211);
xor XOR2 (N8726, N8710, N8656);
xor XOR2 (N8727, N8721, N3954);
not NOT1 (N8728, N8727);
xor XOR2 (N8729, N8704, N2167);
buf BUF1 (N8730, N8726);
not NOT1 (N8731, N8724);
xor XOR2 (N8732, N8728, N4495);
buf BUF1 (N8733, N8725);
nor NOR4 (N8734, N8719, N4024, N4835, N7318);
not NOT1 (N8735, N8730);
and AND3 (N8736, N8735, N2272, N7464);
nand NAND3 (N8737, N8729, N1507, N6773);
nor NOR3 (N8738, N8733, N2806, N5222);
and AND4 (N8739, N8720, N8276, N5608, N3215);
buf BUF1 (N8740, N8739);
and AND2 (N8741, N8708, N3704);
and AND3 (N8742, N8731, N8350, N8581);
not NOT1 (N8743, N8713);
buf BUF1 (N8744, N8740);
not NOT1 (N8745, N8732);
buf BUF1 (N8746, N8738);
nor NOR3 (N8747, N8718, N1564, N3224);
and AND2 (N8748, N8741, N3218);
not NOT1 (N8749, N8736);
nand NAND4 (N8750, N8746, N787, N5756, N3354);
nor NOR3 (N8751, N8737, N1009, N8371);
and AND3 (N8752, N8748, N5194, N1124);
buf BUF1 (N8753, N8750);
not NOT1 (N8754, N8753);
or OR2 (N8755, N8743, N7641);
and AND4 (N8756, N8734, N4528, N8296, N3421);
nand NAND3 (N8757, N8752, N7848, N865);
buf BUF1 (N8758, N8751);
not NOT1 (N8759, N8758);
buf BUF1 (N8760, N8744);
nand NAND4 (N8761, N8755, N7805, N7777, N1478);
xor XOR2 (N8762, N8749, N1485);
not NOT1 (N8763, N8756);
nor NOR4 (N8764, N8759, N1860, N6182, N6354);
nand NAND4 (N8765, N8760, N6110, N5894, N3128);
or OR2 (N8766, N8747, N6717);
xor XOR2 (N8767, N8742, N5142);
and AND3 (N8768, N8766, N2689, N431);
and AND3 (N8769, N8767, N8644, N4745);
nand NAND2 (N8770, N8763, N524);
and AND4 (N8771, N8764, N7580, N6080, N339);
xor XOR2 (N8772, N8754, N392);
not NOT1 (N8773, N8772);
and AND3 (N8774, N8769, N1939, N1189);
nor NOR3 (N8775, N8771, N4702, N294);
buf BUF1 (N8776, N8775);
nor NOR2 (N8777, N8745, N2719);
xor XOR2 (N8778, N8770, N4688);
nor NOR3 (N8779, N8774, N4182, N5690);
buf BUF1 (N8780, N8777);
xor XOR2 (N8781, N8776, N6389);
nor NOR3 (N8782, N8768, N4102, N1601);
nor NOR4 (N8783, N8780, N797, N6731, N6081);
nand NAND3 (N8784, N8778, N8240, N5989);
nor NOR3 (N8785, N8779, N7880, N6453);
or OR2 (N8786, N8785, N4580);
and AND3 (N8787, N8773, N7782, N8515);
buf BUF1 (N8788, N8761);
nand NAND2 (N8789, N8762, N276);
nor NOR2 (N8790, N8781, N5125);
xor XOR2 (N8791, N8783, N1691);
or OR2 (N8792, N8786, N1730);
buf BUF1 (N8793, N8789);
and AND4 (N8794, N8765, N37, N5888, N3230);
or OR3 (N8795, N8794, N1051, N8631);
nand NAND2 (N8796, N8793, N6642);
and AND3 (N8797, N8782, N711, N1892);
not NOT1 (N8798, N8796);
and AND4 (N8799, N8788, N1940, N724, N3898);
and AND2 (N8800, N8790, N3509);
and AND3 (N8801, N8784, N3364, N6741);
nand NAND4 (N8802, N8795, N4182, N196, N7937);
nand NAND4 (N8803, N8800, N195, N2457, N3096);
nor NOR3 (N8804, N8757, N8461, N5564);
nor NOR2 (N8805, N8803, N2596);
or OR2 (N8806, N8802, N7087);
nand NAND2 (N8807, N8797, N1560);
nor NOR4 (N8808, N8801, N7559, N7653, N8682);
xor XOR2 (N8809, N8799, N7025);
not NOT1 (N8810, N8805);
nor NOR2 (N8811, N8809, N4491);
not NOT1 (N8812, N8806);
or OR2 (N8813, N8808, N4627);
xor XOR2 (N8814, N8787, N1228);
xor XOR2 (N8815, N8792, N681);
or OR4 (N8816, N8812, N8295, N8323, N664);
buf BUF1 (N8817, N8811);
nor NOR4 (N8818, N8810, N5145, N506, N2515);
nand NAND3 (N8819, N8814, N321, N3792);
not NOT1 (N8820, N8807);
and AND4 (N8821, N8816, N7770, N4766, N21);
nand NAND3 (N8822, N8821, N2257, N8816);
not NOT1 (N8823, N8813);
xor XOR2 (N8824, N8815, N8401);
buf BUF1 (N8825, N8791);
xor XOR2 (N8826, N8798, N7292);
or OR3 (N8827, N8819, N1736, N7654);
or OR4 (N8828, N8804, N2861, N7737, N6164);
or OR2 (N8829, N8820, N2663);
xor XOR2 (N8830, N8817, N2642);
and AND4 (N8831, N8829, N6475, N1387, N8404);
nor NOR4 (N8832, N8826, N4409, N5230, N3471);
or OR4 (N8833, N8831, N7500, N323, N6252);
or OR3 (N8834, N8818, N687, N8828);
nand NAND2 (N8835, N7607, N1852);
nor NOR2 (N8836, N8827, N6461);
and AND4 (N8837, N8835, N2729, N8328, N747);
and AND3 (N8838, N8822, N7657, N4353);
not NOT1 (N8839, N8823);
nand NAND4 (N8840, N8824, N7144, N6566, N6634);
and AND2 (N8841, N8825, N3004);
and AND2 (N8842, N8840, N3096);
nor NOR4 (N8843, N8839, N5627, N1353, N146);
not NOT1 (N8844, N8837);
buf BUF1 (N8845, N8838);
or OR3 (N8846, N8832, N7283, N8568);
nor NOR2 (N8847, N8830, N3792);
or OR4 (N8848, N8847, N5357, N6435, N1555);
buf BUF1 (N8849, N8844);
not NOT1 (N8850, N8846);
nor NOR2 (N8851, N8841, N4934);
not NOT1 (N8852, N8849);
not NOT1 (N8853, N8848);
nor NOR3 (N8854, N8850, N7799, N7750);
nand NAND3 (N8855, N8853, N8756, N2298);
not NOT1 (N8856, N8834);
or OR2 (N8857, N8851, N7192);
nor NOR2 (N8858, N8857, N7389);
and AND2 (N8859, N8854, N7555);
buf BUF1 (N8860, N8845);
nand NAND3 (N8861, N8842, N7398, N2338);
xor XOR2 (N8862, N8855, N7759);
buf BUF1 (N8863, N8836);
and AND3 (N8864, N8858, N591, N6111);
buf BUF1 (N8865, N8852);
nand NAND3 (N8866, N8865, N268, N1139);
not NOT1 (N8867, N8862);
nand NAND3 (N8868, N8843, N761, N2188);
or OR4 (N8869, N8867, N1339, N736, N3472);
and AND4 (N8870, N8863, N1069, N2869, N6052);
not NOT1 (N8871, N8856);
nand NAND2 (N8872, N8859, N6932);
nor NOR3 (N8873, N8872, N3180, N7769);
xor XOR2 (N8874, N8871, N1173);
xor XOR2 (N8875, N8861, N6739);
or OR2 (N8876, N8860, N4853);
buf BUF1 (N8877, N8874);
buf BUF1 (N8878, N8873);
xor XOR2 (N8879, N8833, N554);
and AND3 (N8880, N8870, N3907, N2971);
nor NOR2 (N8881, N8869, N5134);
nand NAND4 (N8882, N8864, N3394, N8572, N4308);
or OR4 (N8883, N8880, N4216, N6626, N2033);
nand NAND4 (N8884, N8877, N6357, N4624, N8372);
xor XOR2 (N8885, N8876, N5174);
nor NOR2 (N8886, N8866, N2782);
and AND4 (N8887, N8879, N3323, N8594, N4973);
nand NAND4 (N8888, N8882, N8350, N914, N6836);
buf BUF1 (N8889, N8881);
buf BUF1 (N8890, N8888);
buf BUF1 (N8891, N8889);
and AND3 (N8892, N8875, N2623, N6545);
nor NOR4 (N8893, N8868, N6207, N7656, N66);
not NOT1 (N8894, N8892);
xor XOR2 (N8895, N8894, N991);
not NOT1 (N8896, N8895);
nand NAND3 (N8897, N8890, N8390, N7792);
xor XOR2 (N8898, N8883, N2530);
or OR3 (N8899, N8886, N8128, N547);
and AND2 (N8900, N8885, N3775);
not NOT1 (N8901, N8878);
and AND3 (N8902, N8898, N4632, N3801);
buf BUF1 (N8903, N8887);
and AND2 (N8904, N8884, N6742);
nor NOR3 (N8905, N8904, N7661, N8357);
xor XOR2 (N8906, N8899, N2137);
buf BUF1 (N8907, N8902);
or OR2 (N8908, N8906, N6170);
or OR4 (N8909, N8900, N852, N8697, N8183);
not NOT1 (N8910, N8903);
and AND3 (N8911, N8905, N4219, N1312);
nor NOR2 (N8912, N8907, N5134);
or OR2 (N8913, N8910, N7198);
nand NAND4 (N8914, N8897, N5755, N8455, N8636);
buf BUF1 (N8915, N8896);
not NOT1 (N8916, N8893);
buf BUF1 (N8917, N8915);
and AND4 (N8918, N8911, N5261, N7943, N8140);
or OR4 (N8919, N8912, N2268, N5781, N1528);
nor NOR2 (N8920, N8916, N1948);
buf BUF1 (N8921, N8920);
and AND3 (N8922, N8918, N617, N6705);
buf BUF1 (N8923, N8921);
not NOT1 (N8924, N8909);
or OR3 (N8925, N8922, N1514, N3602);
xor XOR2 (N8926, N8913, N3906);
or OR3 (N8927, N8908, N2363, N1513);
and AND4 (N8928, N8926, N4889, N6361, N7207);
nand NAND3 (N8929, N8927, N2785, N3756);
nor NOR3 (N8930, N8891, N5860, N7852);
buf BUF1 (N8931, N8929);
or OR3 (N8932, N8901, N4289, N4969);
nor NOR4 (N8933, N8923, N3254, N214, N7023);
xor XOR2 (N8934, N8925, N8723);
and AND4 (N8935, N8917, N1235, N1959, N8296);
and AND4 (N8936, N8924, N1656, N1451, N3974);
buf BUF1 (N8937, N8914);
not NOT1 (N8938, N8919);
nand NAND4 (N8939, N8932, N8807, N6481, N450);
not NOT1 (N8940, N8938);
xor XOR2 (N8941, N8937, N5493);
xor XOR2 (N8942, N8934, N2485);
xor XOR2 (N8943, N8942, N2028);
buf BUF1 (N8944, N8931);
nor NOR3 (N8945, N8940, N8187, N5198);
nand NAND4 (N8946, N8939, N7772, N3072, N8044);
nand NAND2 (N8947, N8945, N6489);
and AND2 (N8948, N8943, N4563);
not NOT1 (N8949, N8933);
nand NAND2 (N8950, N8935, N8943);
xor XOR2 (N8951, N8949, N4927);
buf BUF1 (N8952, N8936);
xor XOR2 (N8953, N8944, N5425);
buf BUF1 (N8954, N8952);
buf BUF1 (N8955, N8951);
not NOT1 (N8956, N8930);
xor XOR2 (N8957, N8941, N8427);
or OR4 (N8958, N8950, N2881, N8573, N8061);
xor XOR2 (N8959, N8957, N5587);
nand NAND3 (N8960, N8959, N7187, N2957);
and AND4 (N8961, N8958, N6455, N7780, N6072);
nor NOR3 (N8962, N8955, N8357, N5794);
nor NOR4 (N8963, N8956, N8705, N8399, N2822);
buf BUF1 (N8964, N8946);
buf BUF1 (N8965, N8960);
nor NOR3 (N8966, N8961, N8463, N7525);
buf BUF1 (N8967, N8954);
nand NAND2 (N8968, N8947, N1374);
and AND4 (N8969, N8963, N5523, N4222, N6827);
and AND2 (N8970, N8968, N1553);
nand NAND2 (N8971, N8953, N1887);
nor NOR3 (N8972, N8969, N3579, N964);
xor XOR2 (N8973, N8967, N283);
buf BUF1 (N8974, N8964);
buf BUF1 (N8975, N8928);
nand NAND3 (N8976, N8975, N8676, N5360);
nor NOR4 (N8977, N8966, N2753, N8421, N5317);
not NOT1 (N8978, N8972);
buf BUF1 (N8979, N8948);
or OR4 (N8980, N8979, N369, N8235, N1896);
nor NOR2 (N8981, N8976, N1560);
or OR3 (N8982, N8978, N8063, N5407);
and AND3 (N8983, N8974, N2537, N4994);
or OR3 (N8984, N8982, N8209, N5665);
xor XOR2 (N8985, N8981, N6797);
not NOT1 (N8986, N8971);
xor XOR2 (N8987, N8977, N5947);
nand NAND2 (N8988, N8986, N7848);
xor XOR2 (N8989, N8983, N5824);
xor XOR2 (N8990, N8980, N2562);
not NOT1 (N8991, N8990);
not NOT1 (N8992, N8962);
buf BUF1 (N8993, N8987);
xor XOR2 (N8994, N8985, N6505);
buf BUF1 (N8995, N8973);
nor NOR4 (N8996, N8970, N872, N1546, N928);
not NOT1 (N8997, N8991);
nand NAND2 (N8998, N8994, N658);
nor NOR4 (N8999, N8996, N987, N5759, N6268);
xor XOR2 (N9000, N8997, N7167);
xor XOR2 (N9001, N9000, N8894);
nor NOR2 (N9002, N8998, N8269);
not NOT1 (N9003, N9002);
or OR3 (N9004, N8995, N904, N4993);
xor XOR2 (N9005, N9001, N5649);
nor NOR4 (N9006, N8988, N3091, N4751, N406);
not NOT1 (N9007, N9004);
xor XOR2 (N9008, N8999, N3350);
and AND2 (N9009, N8993, N8948);
and AND2 (N9010, N8965, N2323);
nor NOR4 (N9011, N9007, N5535, N6955, N8580);
nand NAND4 (N9012, N9010, N8351, N5319, N7524);
buf BUF1 (N9013, N9005);
buf BUF1 (N9014, N9006);
not NOT1 (N9015, N8984);
xor XOR2 (N9016, N8989, N7420);
nand NAND2 (N9017, N9015, N2677);
nor NOR2 (N9018, N9009, N1401);
buf BUF1 (N9019, N9013);
not NOT1 (N9020, N9014);
xor XOR2 (N9021, N9019, N4985);
and AND4 (N9022, N9020, N7760, N1841, N7943);
not NOT1 (N9023, N9017);
xor XOR2 (N9024, N9011, N2055);
not NOT1 (N9025, N9003);
nand NAND2 (N9026, N9023, N7676);
buf BUF1 (N9027, N9026);
or OR2 (N9028, N9018, N1238);
xor XOR2 (N9029, N8992, N7002);
and AND2 (N9030, N9029, N5639);
not NOT1 (N9031, N9016);
nand NAND2 (N9032, N9024, N5792);
and AND3 (N9033, N9030, N535, N2320);
not NOT1 (N9034, N9032);
nor NOR4 (N9035, N9008, N1601, N7084, N2319);
nor NOR2 (N9036, N9022, N6419);
nand NAND2 (N9037, N9025, N2538);
and AND2 (N9038, N9031, N1523);
nor NOR3 (N9039, N9033, N3732, N8492);
or OR3 (N9040, N9021, N6691, N2795);
or OR2 (N9041, N9037, N213);
nor NOR3 (N9042, N9012, N1913, N5637);
xor XOR2 (N9043, N9035, N1752);
nor NOR3 (N9044, N9038, N1098, N2561);
xor XOR2 (N9045, N9036, N4139);
buf BUF1 (N9046, N9043);
and AND4 (N9047, N9027, N3459, N6957, N631);
or OR4 (N9048, N9047, N1040, N3358, N5608);
nand NAND4 (N9049, N9044, N1131, N633, N1547);
or OR2 (N9050, N9046, N6380);
and AND4 (N9051, N9050, N1483, N2445, N749);
nand NAND4 (N9052, N9042, N4005, N8466, N3306);
and AND4 (N9053, N9028, N6295, N6533, N5658);
not NOT1 (N9054, N9049);
nand NAND4 (N9055, N9041, N8815, N8764, N4165);
not NOT1 (N9056, N9039);
xor XOR2 (N9057, N9055, N5259);
xor XOR2 (N9058, N9040, N1125);
xor XOR2 (N9059, N9057, N7541);
xor XOR2 (N9060, N9052, N2442);
not NOT1 (N9061, N9045);
buf BUF1 (N9062, N9061);
and AND3 (N9063, N9053, N8954, N5541);
not NOT1 (N9064, N9051);
nor NOR4 (N9065, N9056, N7870, N97, N4693);
buf BUF1 (N9066, N9062);
buf BUF1 (N9067, N9058);
and AND3 (N9068, N9048, N3985, N5913);
nand NAND3 (N9069, N9064, N4595, N2548);
nor NOR4 (N9070, N9066, N7813, N6892, N7855);
nand NAND4 (N9071, N9068, N55, N5858, N2842);
nor NOR4 (N9072, N9054, N3107, N5641, N8316);
xor XOR2 (N9073, N9034, N6045);
xor XOR2 (N9074, N9073, N7479);
nor NOR4 (N9075, N9074, N8242, N4020, N3796);
nand NAND2 (N9076, N9065, N4303);
nand NAND3 (N9077, N9067, N1772, N1630);
nand NAND2 (N9078, N9059, N6598);
not NOT1 (N9079, N9075);
and AND3 (N9080, N9063, N7110, N1363);
and AND3 (N9081, N9079, N6344, N4100);
xor XOR2 (N9082, N9070, N3178);
not NOT1 (N9083, N9080);
and AND3 (N9084, N9081, N5461, N4456);
nand NAND2 (N9085, N9069, N771);
buf BUF1 (N9086, N9082);
and AND2 (N9087, N9083, N3727);
xor XOR2 (N9088, N9060, N3877);
and AND2 (N9089, N9086, N7699);
buf BUF1 (N9090, N9089);
and AND3 (N9091, N9084, N7594, N4685);
nand NAND2 (N9092, N9072, N6207);
and AND3 (N9093, N9090, N3438, N227);
nand NAND3 (N9094, N9087, N1288, N6070);
nand NAND3 (N9095, N9091, N1317, N8391);
and AND2 (N9096, N9092, N7432);
not NOT1 (N9097, N9094);
nor NOR4 (N9098, N9078, N822, N3736, N8215);
xor XOR2 (N9099, N9093, N2780);
nor NOR4 (N9100, N9095, N8528, N512, N3868);
xor XOR2 (N9101, N9099, N3130);
and AND2 (N9102, N9101, N8961);
xor XOR2 (N9103, N9088, N1248);
buf BUF1 (N9104, N9097);
not NOT1 (N9105, N9103);
nand NAND3 (N9106, N9104, N2172, N5253);
not NOT1 (N9107, N9106);
and AND2 (N9108, N9105, N4858);
or OR2 (N9109, N9098, N3831);
xor XOR2 (N9110, N9076, N2716);
buf BUF1 (N9111, N9107);
nor NOR2 (N9112, N9077, N8894);
buf BUF1 (N9113, N9071);
nand NAND2 (N9114, N9096, N7173);
nand NAND3 (N9115, N9100, N1343, N504);
nor NOR4 (N9116, N9112, N8200, N4198, N6104);
buf BUF1 (N9117, N9114);
or OR3 (N9118, N9109, N3317, N2597);
buf BUF1 (N9119, N9118);
xor XOR2 (N9120, N9110, N2626);
not NOT1 (N9121, N9116);
buf BUF1 (N9122, N9085);
or OR3 (N9123, N9122, N1157, N3536);
or OR3 (N9124, N9120, N7023, N8717);
not NOT1 (N9125, N9111);
xor XOR2 (N9126, N9124, N3584);
nand NAND4 (N9127, N9115, N1245, N3527, N7845);
or OR3 (N9128, N9126, N1790, N6229);
nand NAND2 (N9129, N9102, N3510);
not NOT1 (N9130, N9117);
or OR4 (N9131, N9128, N5555, N332, N1797);
not NOT1 (N9132, N9130);
not NOT1 (N9133, N9125);
nand NAND3 (N9134, N9121, N8689, N7186);
buf BUF1 (N9135, N9119);
nor NOR2 (N9136, N9132, N4293);
or OR4 (N9137, N9134, N4812, N4138, N6057);
or OR3 (N9138, N9135, N1791, N7956);
and AND2 (N9139, N9131, N8931);
not NOT1 (N9140, N9137);
xor XOR2 (N9141, N9129, N4665);
or OR4 (N9142, N9140, N1089, N1924, N49);
and AND3 (N9143, N9123, N3599, N2132);
not NOT1 (N9144, N9142);
xor XOR2 (N9145, N9139, N5499);
and AND3 (N9146, N9113, N3858, N5815);
buf BUF1 (N9147, N9145);
nor NOR2 (N9148, N9146, N5976);
nand NAND3 (N9149, N9148, N6046, N3972);
buf BUF1 (N9150, N9108);
or OR3 (N9151, N9149, N7249, N2704);
nor NOR2 (N9152, N9136, N4324);
xor XOR2 (N9153, N9151, N2894);
nand NAND4 (N9154, N9141, N4173, N6693, N4810);
xor XOR2 (N9155, N9154, N2363);
not NOT1 (N9156, N9153);
or OR2 (N9157, N9133, N7079);
and AND4 (N9158, N9127, N404, N6849, N7327);
or OR3 (N9159, N9158, N8757, N9105);
buf BUF1 (N9160, N9156);
nand NAND3 (N9161, N9143, N2741, N2500);
nand NAND2 (N9162, N9144, N8057);
nor NOR4 (N9163, N9161, N7622, N2734, N5360);
or OR4 (N9164, N9159, N2262, N4799, N5461);
and AND4 (N9165, N9162, N3000, N1238, N4452);
xor XOR2 (N9166, N9150, N5704);
buf BUF1 (N9167, N9160);
xor XOR2 (N9168, N9152, N8695);
xor XOR2 (N9169, N9138, N4532);
and AND4 (N9170, N9164, N7956, N5569, N6713);
not NOT1 (N9171, N9169);
nand NAND2 (N9172, N9147, N4770);
nand NAND2 (N9173, N9155, N6822);
not NOT1 (N9174, N9170);
not NOT1 (N9175, N9168);
nand NAND2 (N9176, N9174, N5205);
nand NAND3 (N9177, N9163, N4470, N5326);
nand NAND4 (N9178, N9173, N7811, N3823, N7500);
xor XOR2 (N9179, N9172, N5440);
or OR3 (N9180, N9171, N7250, N3799);
xor XOR2 (N9181, N9176, N3273);
nand NAND4 (N9182, N9180, N860, N372, N5657);
nand NAND4 (N9183, N9182, N2539, N6382, N4059);
and AND4 (N9184, N9166, N2154, N3083, N1819);
or OR3 (N9185, N9177, N7579, N6217);
xor XOR2 (N9186, N9183, N2729);
buf BUF1 (N9187, N9184);
and AND2 (N9188, N9165, N6390);
or OR2 (N9189, N9157, N9117);
nor NOR2 (N9190, N9167, N6684);
buf BUF1 (N9191, N9187);
not NOT1 (N9192, N9185);
or OR3 (N9193, N9190, N1620, N2616);
nor NOR4 (N9194, N9192, N4672, N8360, N7694);
nor NOR2 (N9195, N9193, N3608);
not NOT1 (N9196, N9181);
and AND2 (N9197, N9175, N6446);
nor NOR3 (N9198, N9196, N8338, N8963);
nand NAND2 (N9199, N9195, N6213);
nor NOR3 (N9200, N9188, N7733, N8776);
or OR4 (N9201, N9186, N5622, N8213, N3016);
nor NOR3 (N9202, N9198, N8917, N7716);
not NOT1 (N9203, N9200);
not NOT1 (N9204, N9178);
buf BUF1 (N9205, N9179);
nor NOR3 (N9206, N9201, N6706, N7593);
not NOT1 (N9207, N9203);
nor NOR3 (N9208, N9189, N3306, N7789);
and AND3 (N9209, N9205, N4808, N1144);
buf BUF1 (N9210, N9204);
buf BUF1 (N9211, N9197);
or OR3 (N9212, N9209, N1533, N4460);
nor NOR3 (N9213, N9210, N1235, N657);
xor XOR2 (N9214, N9207, N4077);
and AND2 (N9215, N9202, N4917);
buf BUF1 (N9216, N9215);
xor XOR2 (N9217, N9206, N1555);
buf BUF1 (N9218, N9199);
nor NOR3 (N9219, N9217, N4680, N8437);
xor XOR2 (N9220, N9212, N4133);
xor XOR2 (N9221, N9216, N6177);
nand NAND3 (N9222, N9218, N6656, N4626);
nor NOR3 (N9223, N9220, N1370, N8700);
nand NAND3 (N9224, N9219, N6021, N5843);
buf BUF1 (N9225, N9213);
or OR3 (N9226, N9221, N5339, N5409);
buf BUF1 (N9227, N9222);
nor NOR3 (N9228, N9223, N485, N266);
nor NOR4 (N9229, N9194, N2561, N6428, N1155);
or OR3 (N9230, N9191, N6213, N708);
nand NAND2 (N9231, N9224, N7548);
or OR2 (N9232, N9227, N4833);
nand NAND3 (N9233, N9211, N8327, N9186);
xor XOR2 (N9234, N9228, N7164);
or OR2 (N9235, N9230, N8032);
nor NOR2 (N9236, N9225, N6214);
nand NAND2 (N9237, N9229, N6607);
or OR3 (N9238, N9233, N7794, N4247);
buf BUF1 (N9239, N9236);
nand NAND2 (N9240, N9239, N2127);
nand NAND2 (N9241, N9237, N8732);
or OR2 (N9242, N9231, N8842);
xor XOR2 (N9243, N9238, N624);
or OR2 (N9244, N9241, N2394);
or OR4 (N9245, N9234, N9035, N6065, N5175);
or OR4 (N9246, N9243, N380, N4010, N8155);
nand NAND3 (N9247, N9244, N7530, N3078);
and AND2 (N9248, N9247, N6364);
nor NOR4 (N9249, N9214, N8249, N6104, N8811);
or OR2 (N9250, N9235, N1370);
or OR3 (N9251, N9226, N2292, N2447);
or OR3 (N9252, N9240, N5052, N912);
buf BUF1 (N9253, N9250);
or OR3 (N9254, N9248, N1724, N4660);
nand NAND4 (N9255, N9252, N993, N4978, N4410);
and AND3 (N9256, N9255, N936, N4875);
and AND2 (N9257, N9232, N6614);
not NOT1 (N9258, N9254);
buf BUF1 (N9259, N9249);
not NOT1 (N9260, N9208);
nor NOR4 (N9261, N9253, N7382, N5956, N1287);
xor XOR2 (N9262, N9259, N4391);
or OR3 (N9263, N9251, N999, N1489);
nor NOR2 (N9264, N9245, N2532);
buf BUF1 (N9265, N9258);
nor NOR2 (N9266, N9242, N9111);
nor NOR4 (N9267, N9246, N4672, N4395, N8479);
buf BUF1 (N9268, N9257);
nor NOR3 (N9269, N9267, N8607, N1730);
and AND2 (N9270, N9263, N3786);
nor NOR2 (N9271, N9268, N3474);
buf BUF1 (N9272, N9266);
and AND2 (N9273, N9272, N2192);
not NOT1 (N9274, N9261);
or OR4 (N9275, N9264, N5583, N4480, N1954);
buf BUF1 (N9276, N9271);
buf BUF1 (N9277, N9260);
not NOT1 (N9278, N9276);
nand NAND3 (N9279, N9269, N2389, N8992);
buf BUF1 (N9280, N9262);
nor NOR4 (N9281, N9265, N7765, N2252, N888);
and AND3 (N9282, N9281, N6731, N3772);
nor NOR4 (N9283, N9278, N3445, N4169, N3194);
or OR3 (N9284, N9270, N2957, N8106);
xor XOR2 (N9285, N9277, N7930);
xor XOR2 (N9286, N9275, N863);
xor XOR2 (N9287, N9273, N614);
buf BUF1 (N9288, N9256);
nand NAND4 (N9289, N9285, N647, N4823, N6713);
not NOT1 (N9290, N9288);
buf BUF1 (N9291, N9280);
xor XOR2 (N9292, N9274, N5738);
xor XOR2 (N9293, N9289, N3594);
buf BUF1 (N9294, N9293);
xor XOR2 (N9295, N9291, N3758);
buf BUF1 (N9296, N9287);
nor NOR4 (N9297, N9292, N4756, N6867, N9086);
buf BUF1 (N9298, N9279);
not NOT1 (N9299, N9296);
not NOT1 (N9300, N9298);
nand NAND3 (N9301, N9283, N817, N7376);
nand NAND4 (N9302, N9290, N7617, N1171, N4113);
buf BUF1 (N9303, N9297);
nand NAND4 (N9304, N9299, N2479, N7974, N7289);
buf BUF1 (N9305, N9284);
and AND2 (N9306, N9302, N7560);
xor XOR2 (N9307, N9286, N1890);
and AND3 (N9308, N9282, N6581, N128);
nand NAND4 (N9309, N9301, N4398, N7394, N2803);
and AND3 (N9310, N9303, N5532, N5504);
and AND2 (N9311, N9295, N2917);
not NOT1 (N9312, N9307);
nor NOR3 (N9313, N9305, N4273, N4272);
and AND2 (N9314, N9312, N8019);
nor NOR2 (N9315, N9304, N4441);
buf BUF1 (N9316, N9294);
and AND2 (N9317, N9311, N8374);
xor XOR2 (N9318, N9314, N7460);
xor XOR2 (N9319, N9310, N7181);
and AND2 (N9320, N9316, N1522);
buf BUF1 (N9321, N9308);
not NOT1 (N9322, N9317);
buf BUF1 (N9323, N9309);
buf BUF1 (N9324, N9306);
nor NOR3 (N9325, N9318, N6507, N2100);
and AND2 (N9326, N9315, N3181);
nor NOR4 (N9327, N9321, N6857, N188, N3835);
nand NAND3 (N9328, N9327, N1458, N3629);
nor NOR2 (N9329, N9319, N3843);
and AND2 (N9330, N9325, N4010);
or OR2 (N9331, N9329, N8234);
buf BUF1 (N9332, N9328);
not NOT1 (N9333, N9332);
buf BUF1 (N9334, N9322);
or OR4 (N9335, N9313, N1274, N6982, N2816);
xor XOR2 (N9336, N9324, N135);
nor NOR4 (N9337, N9320, N636, N9272, N6360);
nor NOR2 (N9338, N9330, N6188);
nor NOR2 (N9339, N9337, N1192);
or OR3 (N9340, N9300, N3282, N2466);
buf BUF1 (N9341, N9323);
and AND2 (N9342, N9336, N5185);
not NOT1 (N9343, N9335);
xor XOR2 (N9344, N9340, N1440);
or OR4 (N9345, N9344, N4384, N6333, N6317);
not NOT1 (N9346, N9342);
nor NOR2 (N9347, N9333, N835);
buf BUF1 (N9348, N9346);
not NOT1 (N9349, N9343);
nor NOR4 (N9350, N9348, N2635, N7352, N2867);
and AND2 (N9351, N9341, N175);
not NOT1 (N9352, N9349);
buf BUF1 (N9353, N9352);
buf BUF1 (N9354, N9345);
buf BUF1 (N9355, N9334);
and AND3 (N9356, N9331, N3771, N7296);
or OR2 (N9357, N9338, N4599);
and AND2 (N9358, N9355, N6027);
and AND4 (N9359, N9347, N3986, N4237, N198);
xor XOR2 (N9360, N9354, N6468);
xor XOR2 (N9361, N9339, N4922);
and AND2 (N9362, N9356, N6320);
or OR2 (N9363, N9351, N253);
or OR2 (N9364, N9361, N8752);
nand NAND3 (N9365, N9363, N3183, N5191);
xor XOR2 (N9366, N9365, N4018);
or OR4 (N9367, N9359, N7865, N5445, N1560);
and AND2 (N9368, N9360, N88);
or OR4 (N9369, N9366, N2184, N4868, N898);
xor XOR2 (N9370, N9353, N756);
not NOT1 (N9371, N9368);
or OR4 (N9372, N9358, N1838, N3785, N5730);
xor XOR2 (N9373, N9372, N6068);
not NOT1 (N9374, N9357);
buf BUF1 (N9375, N9362);
nand NAND3 (N9376, N9374, N7052, N4520);
or OR3 (N9377, N9364, N3679, N1966);
or OR3 (N9378, N9370, N7254, N5039);
nand NAND2 (N9379, N9367, N6399);
xor XOR2 (N9380, N9326, N3163);
xor XOR2 (N9381, N9373, N5059);
and AND4 (N9382, N9375, N3797, N5204, N9275);
xor XOR2 (N9383, N9371, N5087);
nor NOR2 (N9384, N9369, N1855);
or OR2 (N9385, N9384, N506);
nand NAND3 (N9386, N9379, N2479, N401);
nor NOR2 (N9387, N9350, N9247);
xor XOR2 (N9388, N9380, N2341);
buf BUF1 (N9389, N9385);
nand NAND4 (N9390, N9389, N7785, N3516, N8370);
nor NOR2 (N9391, N9387, N5517);
and AND4 (N9392, N9378, N1127, N3005, N8999);
and AND2 (N9393, N9376, N2434);
not NOT1 (N9394, N9388);
and AND4 (N9395, N9391, N6687, N5295, N3458);
nor NOR4 (N9396, N9394, N1268, N6329, N5010);
nand NAND3 (N9397, N9386, N3340, N6152);
nor NOR4 (N9398, N9382, N1048, N1704, N8756);
nor NOR4 (N9399, N9396, N3259, N8457, N5744);
or OR4 (N9400, N9398, N8042, N7064, N8765);
nor NOR4 (N9401, N9399, N3468, N1156, N6059);
or OR3 (N9402, N9395, N986, N8927);
nand NAND2 (N9403, N9383, N1094);
nand NAND3 (N9404, N9402, N3176, N1865);
and AND3 (N9405, N9393, N8921, N7585);
nor NOR2 (N9406, N9403, N7308);
buf BUF1 (N9407, N9392);
or OR2 (N9408, N9407, N8717);
xor XOR2 (N9409, N9408, N1223);
not NOT1 (N9410, N9401);
not NOT1 (N9411, N9390);
nand NAND2 (N9412, N9397, N4149);
xor XOR2 (N9413, N9411, N1548);
not NOT1 (N9414, N9410);
and AND2 (N9415, N9377, N2739);
not NOT1 (N9416, N9409);
and AND2 (N9417, N9412, N6095);
not NOT1 (N9418, N9381);
nor NOR2 (N9419, N9415, N9126);
nor NOR3 (N9420, N9400, N6681, N4491);
nand NAND2 (N9421, N9420, N4793);
and AND2 (N9422, N9416, N1032);
buf BUF1 (N9423, N9419);
nor NOR2 (N9424, N9421, N393);
xor XOR2 (N9425, N9424, N1003);
nand NAND3 (N9426, N9414, N1141, N1839);
or OR4 (N9427, N9418, N8385, N2298, N6692);
xor XOR2 (N9428, N9413, N8237);
or OR4 (N9429, N9425, N553, N9145, N9022);
nand NAND4 (N9430, N9428, N7348, N1178, N1880);
nand NAND2 (N9431, N9423, N789);
xor XOR2 (N9432, N9406, N5394);
nand NAND3 (N9433, N9405, N427, N7046);
xor XOR2 (N9434, N9432, N4835);
buf BUF1 (N9435, N9426);
or OR4 (N9436, N9431, N3763, N8238, N6794);
or OR2 (N9437, N9404, N4030);
not NOT1 (N9438, N9437);
and AND3 (N9439, N9422, N8399, N6640);
buf BUF1 (N9440, N9434);
and AND4 (N9441, N9430, N7119, N6283, N8674);
nor NOR2 (N9442, N9440, N6218);
not NOT1 (N9443, N9441);
or OR4 (N9444, N9442, N1143, N3283, N1120);
not NOT1 (N9445, N9429);
or OR3 (N9446, N9443, N2851, N3829);
xor XOR2 (N9447, N9439, N8295);
not NOT1 (N9448, N9438);
xor XOR2 (N9449, N9448, N8859);
not NOT1 (N9450, N9447);
and AND2 (N9451, N9449, N6755);
and AND3 (N9452, N9446, N3275, N727);
nor NOR4 (N9453, N9450, N7559, N288, N7934);
and AND4 (N9454, N9453, N5429, N8678, N1043);
and AND4 (N9455, N9435, N6415, N4685, N5005);
not NOT1 (N9456, N9454);
or OR4 (N9457, N9436, N6045, N8398, N7007);
or OR2 (N9458, N9457, N1909);
or OR3 (N9459, N9458, N8735, N1589);
nor NOR4 (N9460, N9459, N4221, N7064, N2507);
not NOT1 (N9461, N9456);
nor NOR4 (N9462, N9445, N5054, N5091, N8739);
xor XOR2 (N9463, N9451, N2214);
nor NOR4 (N9464, N9427, N3080, N2532, N4042);
nor NOR3 (N9465, N9417, N3802, N7338);
and AND4 (N9466, N9452, N446, N6505, N7882);
nand NAND2 (N9467, N9444, N5724);
and AND2 (N9468, N9467, N7394);
nor NOR4 (N9469, N9466, N8009, N4008, N4183);
xor XOR2 (N9470, N9469, N2942);
or OR2 (N9471, N9463, N2315);
nor NOR4 (N9472, N9460, N4525, N7294, N1017);
not NOT1 (N9473, N9471);
nand NAND3 (N9474, N9464, N8975, N1018);
xor XOR2 (N9475, N9472, N4161);
and AND2 (N9476, N9461, N3599);
buf BUF1 (N9477, N9433);
and AND3 (N9478, N9462, N1102, N8221);
nor NOR4 (N9479, N9475, N4958, N6505, N5667);
nor NOR3 (N9480, N9473, N1154, N4137);
nand NAND2 (N9481, N9455, N4684);
not NOT1 (N9482, N9465);
and AND4 (N9483, N9474, N900, N3803, N8104);
buf BUF1 (N9484, N9483);
not NOT1 (N9485, N9479);
or OR4 (N9486, N9468, N6848, N2539, N1011);
not NOT1 (N9487, N9470);
or OR3 (N9488, N9478, N577, N6159);
nand NAND4 (N9489, N9477, N4671, N7387, N3019);
nand NAND4 (N9490, N9489, N4641, N1237, N1438);
xor XOR2 (N9491, N9490, N3681);
or OR2 (N9492, N9484, N3272);
not NOT1 (N9493, N9485);
buf BUF1 (N9494, N9493);
and AND2 (N9495, N9482, N3564);
nand NAND3 (N9496, N9481, N4032, N1837);
nor NOR2 (N9497, N9487, N8167);
nor NOR3 (N9498, N9497, N630, N2418);
or OR2 (N9499, N9496, N288);
and AND3 (N9500, N9495, N7300, N4309);
nand NAND2 (N9501, N9486, N6896);
nand NAND2 (N9502, N9480, N8887);
buf BUF1 (N9503, N9494);
buf BUF1 (N9504, N9501);
nand NAND4 (N9505, N9498, N1245, N9182, N6781);
and AND4 (N9506, N9504, N5698, N4191, N4716);
and AND3 (N9507, N9499, N465, N1112);
and AND4 (N9508, N9503, N3451, N1239, N7586);
and AND3 (N9509, N9502, N4838, N1554);
buf BUF1 (N9510, N9506);
nor NOR3 (N9511, N9500, N4218, N8665);
xor XOR2 (N9512, N9508, N1731);
and AND3 (N9513, N9510, N6589, N3962);
or OR4 (N9514, N9507, N8258, N2724, N516);
not NOT1 (N9515, N9476);
xor XOR2 (N9516, N9492, N224);
or OR4 (N9517, N9515, N4701, N4739, N2581);
or OR3 (N9518, N9512, N2051, N8253);
nand NAND2 (N9519, N9514, N3444);
nor NOR4 (N9520, N9511, N1440, N4799, N6968);
nor NOR3 (N9521, N9509, N8373, N2664);
nand NAND3 (N9522, N9520, N7663, N5677);
buf BUF1 (N9523, N9513);
buf BUF1 (N9524, N9488);
buf BUF1 (N9525, N9519);
buf BUF1 (N9526, N9523);
nand NAND4 (N9527, N9525, N2354, N1112, N3210);
or OR4 (N9528, N9524, N2150, N6119, N7022);
not NOT1 (N9529, N9528);
not NOT1 (N9530, N9527);
xor XOR2 (N9531, N9516, N7806);
nand NAND4 (N9532, N9522, N819, N861, N1780);
nand NAND4 (N9533, N9505, N2832, N2306, N1776);
or OR3 (N9534, N9526, N2694, N344);
or OR3 (N9535, N9532, N7826, N8333);
or OR3 (N9536, N9535, N1472, N6992);
xor XOR2 (N9537, N9517, N6813);
nor NOR4 (N9538, N9533, N6663, N8819, N8814);
nand NAND4 (N9539, N9529, N8223, N6287, N5931);
xor XOR2 (N9540, N9538, N1371);
or OR4 (N9541, N9539, N8275, N1373, N629);
and AND2 (N9542, N9518, N6538);
buf BUF1 (N9543, N9542);
not NOT1 (N9544, N9541);
not NOT1 (N9545, N9537);
or OR3 (N9546, N9543, N7303, N723);
nand NAND4 (N9547, N9491, N4520, N5101, N2694);
or OR3 (N9548, N9545, N1036, N5223);
nor NOR4 (N9549, N9521, N1539, N4723, N8292);
nand NAND3 (N9550, N9546, N1989, N8280);
nand NAND4 (N9551, N9547, N4752, N3665, N540);
nand NAND3 (N9552, N9540, N614, N2216);
buf BUF1 (N9553, N9548);
nand NAND3 (N9554, N9549, N6603, N4169);
nand NAND4 (N9555, N9544, N9296, N7837, N7408);
nor NOR2 (N9556, N9551, N4473);
nand NAND4 (N9557, N9554, N2323, N3630, N7764);
nor NOR2 (N9558, N9555, N8039);
buf BUF1 (N9559, N9531);
nor NOR2 (N9560, N9558, N6239);
buf BUF1 (N9561, N9550);
buf BUF1 (N9562, N9559);
xor XOR2 (N9563, N9560, N8879);
not NOT1 (N9564, N9553);
or OR2 (N9565, N9552, N7574);
xor XOR2 (N9566, N9557, N5648);
nor NOR2 (N9567, N9563, N4439);
or OR3 (N9568, N9564, N6958, N1081);
or OR2 (N9569, N9567, N2947);
nor NOR4 (N9570, N9562, N1337, N8551, N6045);
xor XOR2 (N9571, N9556, N6917);
and AND3 (N9572, N9569, N6888, N2852);
nor NOR2 (N9573, N9570, N3514);
and AND2 (N9574, N9566, N3301);
not NOT1 (N9575, N9534);
xor XOR2 (N9576, N9572, N953);
and AND2 (N9577, N9530, N8796);
nor NOR3 (N9578, N9571, N9262, N2765);
xor XOR2 (N9579, N9573, N596);
or OR4 (N9580, N9565, N3496, N5400, N4978);
or OR3 (N9581, N9579, N8679, N448);
nor NOR2 (N9582, N9576, N5130);
not NOT1 (N9583, N9575);
nand NAND4 (N9584, N9581, N572, N5383, N8355);
or OR3 (N9585, N9577, N3675, N762);
and AND2 (N9586, N9582, N5234);
and AND3 (N9587, N9585, N1270, N146);
nand NAND3 (N9588, N9578, N4059, N3650);
buf BUF1 (N9589, N9568);
and AND4 (N9590, N9586, N5205, N9526, N355);
xor XOR2 (N9591, N9580, N2373);
and AND3 (N9592, N9589, N8624, N5208);
and AND2 (N9593, N9561, N1139);
buf BUF1 (N9594, N9583);
or OR4 (N9595, N9536, N196, N1375, N7482);
xor XOR2 (N9596, N9592, N633);
not NOT1 (N9597, N9587);
not NOT1 (N9598, N9591);
xor XOR2 (N9599, N9597, N5394);
or OR2 (N9600, N9594, N7433);
buf BUF1 (N9601, N9574);
xor XOR2 (N9602, N9595, N9309);
and AND3 (N9603, N9599, N2913, N6519);
and AND4 (N9604, N9603, N7281, N6404, N7171);
nor NOR2 (N9605, N9602, N7557);
buf BUF1 (N9606, N9593);
nor NOR3 (N9607, N9606, N663, N7139);
buf BUF1 (N9608, N9590);
or OR3 (N9609, N9600, N4171, N13);
nor NOR2 (N9610, N9601, N5312);
and AND2 (N9611, N9609, N5510);
buf BUF1 (N9612, N9611);
nand NAND4 (N9613, N9610, N4233, N4769, N9365);
xor XOR2 (N9614, N9613, N2809);
buf BUF1 (N9615, N9598);
nor NOR2 (N9616, N9607, N8019);
or OR4 (N9617, N9588, N5046, N5393, N2981);
not NOT1 (N9618, N9612);
and AND2 (N9619, N9618, N6275);
xor XOR2 (N9620, N9615, N5809);
not NOT1 (N9621, N9596);
xor XOR2 (N9622, N9584, N6799);
and AND3 (N9623, N9614, N9093, N8603);
or OR4 (N9624, N9604, N4439, N5295, N1888);
and AND2 (N9625, N9605, N3385);
and AND4 (N9626, N9608, N6798, N5810, N2975);
not NOT1 (N9627, N9625);
nor NOR3 (N9628, N9616, N4557, N4785);
not NOT1 (N9629, N9627);
nor NOR2 (N9630, N9622, N1424);
nor NOR4 (N9631, N9623, N5784, N6041, N3349);
not NOT1 (N9632, N9617);
buf BUF1 (N9633, N9629);
nor NOR4 (N9634, N9633, N8184, N5080, N3210);
nor NOR2 (N9635, N9630, N5170);
xor XOR2 (N9636, N9634, N9457);
xor XOR2 (N9637, N9636, N7259);
not NOT1 (N9638, N9621);
buf BUF1 (N9639, N9624);
nor NOR2 (N9640, N9639, N2092);
nand NAND2 (N9641, N9628, N7383);
and AND3 (N9642, N9631, N1060, N5507);
nor NOR3 (N9643, N9641, N7862, N5412);
or OR3 (N9644, N9642, N5549, N2917);
nor NOR4 (N9645, N9626, N3691, N7414, N5561);
xor XOR2 (N9646, N9640, N5963);
nand NAND4 (N9647, N9645, N1478, N7468, N837);
nand NAND2 (N9648, N9643, N4691);
and AND2 (N9649, N9635, N1607);
not NOT1 (N9650, N9638);
nand NAND4 (N9651, N9620, N5581, N5484, N5001);
buf BUF1 (N9652, N9651);
or OR3 (N9653, N9647, N6922, N8897);
and AND3 (N9654, N9637, N7703, N5579);
not NOT1 (N9655, N9648);
buf BUF1 (N9656, N9652);
xor XOR2 (N9657, N9644, N4949);
nand NAND3 (N9658, N9646, N319, N7048);
and AND4 (N9659, N9632, N8957, N1760, N9512);
nand NAND2 (N9660, N9659, N6388);
xor XOR2 (N9661, N9619, N9210);
xor XOR2 (N9662, N9655, N4119);
buf BUF1 (N9663, N9654);
buf BUF1 (N9664, N9653);
or OR2 (N9665, N9650, N5583);
nand NAND4 (N9666, N9656, N5185, N4752, N4564);
xor XOR2 (N9667, N9666, N2245);
nand NAND2 (N9668, N9661, N3389);
xor XOR2 (N9669, N9665, N3869);
and AND2 (N9670, N9662, N6013);
buf BUF1 (N9671, N9660);
buf BUF1 (N9672, N9671);
buf BUF1 (N9673, N9649);
buf BUF1 (N9674, N9667);
not NOT1 (N9675, N9663);
nand NAND3 (N9676, N9675, N8119, N9011);
xor XOR2 (N9677, N9674, N8589);
not NOT1 (N9678, N9668);
buf BUF1 (N9679, N9658);
buf BUF1 (N9680, N9677);
and AND2 (N9681, N9673, N398);
not NOT1 (N9682, N9657);
or OR3 (N9683, N9669, N1516, N4637);
buf BUF1 (N9684, N9681);
xor XOR2 (N9685, N9678, N756);
nor NOR2 (N9686, N9672, N5911);
not NOT1 (N9687, N9670);
xor XOR2 (N9688, N9685, N8497);
buf BUF1 (N9689, N9688);
xor XOR2 (N9690, N9683, N1496);
and AND4 (N9691, N9690, N7820, N9535, N4661);
nand NAND2 (N9692, N9664, N4767);
xor XOR2 (N9693, N9680, N406);
not NOT1 (N9694, N9693);
nand NAND4 (N9695, N9686, N8113, N4964, N6521);
not NOT1 (N9696, N9676);
nand NAND4 (N9697, N9691, N9392, N5301, N8653);
buf BUF1 (N9698, N9692);
nor NOR4 (N9699, N9689, N8666, N7971, N8087);
nand NAND4 (N9700, N9684, N261, N4669, N2349);
and AND4 (N9701, N9694, N1891, N3899, N8960);
xor XOR2 (N9702, N9696, N1018);
buf BUF1 (N9703, N9702);
nand NAND2 (N9704, N9682, N787);
nand NAND4 (N9705, N9699, N1708, N7786, N7707);
buf BUF1 (N9706, N9701);
nand NAND2 (N9707, N9698, N8796);
not NOT1 (N9708, N9687);
not NOT1 (N9709, N9706);
not NOT1 (N9710, N9708);
not NOT1 (N9711, N9679);
and AND4 (N9712, N9705, N609, N2363, N281);
nand NAND4 (N9713, N9695, N2797, N8189, N2293);
xor XOR2 (N9714, N9697, N244);
and AND3 (N9715, N9712, N2231, N7416);
xor XOR2 (N9716, N9715, N1118);
xor XOR2 (N9717, N9704, N7794);
buf BUF1 (N9718, N9707);
or OR2 (N9719, N9718, N4242);
and AND4 (N9720, N9711, N5290, N348, N4368);
or OR3 (N9721, N9716, N9331, N3400);
xor XOR2 (N9722, N9703, N1618);
or OR4 (N9723, N9720, N38, N8884, N8277);
or OR3 (N9724, N9713, N6464, N219);
or OR4 (N9725, N9719, N4776, N5009, N5726);
or OR4 (N9726, N9709, N4105, N2318, N1417);
nor NOR3 (N9727, N9721, N782, N5106);
or OR2 (N9728, N9700, N5498);
xor XOR2 (N9729, N9717, N9410);
xor XOR2 (N9730, N9725, N8285);
xor XOR2 (N9731, N9722, N62);
not NOT1 (N9732, N9710);
buf BUF1 (N9733, N9730);
nand NAND3 (N9734, N9727, N632, N2577);
and AND2 (N9735, N9732, N1172);
and AND2 (N9736, N9724, N9664);
buf BUF1 (N9737, N9723);
and AND3 (N9738, N9734, N8990, N4527);
and AND3 (N9739, N9738, N7970, N7999);
nor NOR3 (N9740, N9726, N9230, N3315);
buf BUF1 (N9741, N9729);
nand NAND4 (N9742, N9714, N2417, N6152, N1722);
nand NAND3 (N9743, N9740, N7832, N1901);
buf BUF1 (N9744, N9736);
nand NAND2 (N9745, N9735, N1012);
nand NAND4 (N9746, N9733, N3350, N1068, N2346);
not NOT1 (N9747, N9739);
and AND4 (N9748, N9746, N3118, N7205, N6048);
xor XOR2 (N9749, N9744, N6257);
not NOT1 (N9750, N9742);
xor XOR2 (N9751, N9731, N3756);
or OR3 (N9752, N9751, N5063, N4059);
not NOT1 (N9753, N9749);
xor XOR2 (N9754, N9752, N1953);
xor XOR2 (N9755, N9728, N4552);
buf BUF1 (N9756, N9755);
nand NAND3 (N9757, N9737, N8294, N8180);
or OR4 (N9758, N9747, N9398, N2626, N499);
nand NAND3 (N9759, N9743, N115, N5055);
or OR4 (N9760, N9759, N4258, N7438, N9111);
nor NOR4 (N9761, N9745, N8463, N3853, N9094);
not NOT1 (N9762, N9758);
not NOT1 (N9763, N9760);
nor NOR2 (N9764, N9741, N3191);
or OR3 (N9765, N9754, N1849, N6407);
nand NAND3 (N9766, N9748, N7654, N7171);
buf BUF1 (N9767, N9761);
xor XOR2 (N9768, N9753, N9372);
buf BUF1 (N9769, N9765);
nand NAND2 (N9770, N9764, N905);
xor XOR2 (N9771, N9768, N4018);
not NOT1 (N9772, N9769);
not NOT1 (N9773, N9772);
xor XOR2 (N9774, N9756, N5178);
nor NOR4 (N9775, N9762, N1937, N5874, N1871);
not NOT1 (N9776, N9771);
or OR2 (N9777, N9757, N5);
not NOT1 (N9778, N9776);
nand NAND3 (N9779, N9775, N7233, N6757);
nor NOR2 (N9780, N9773, N7100);
xor XOR2 (N9781, N9778, N2661);
nor NOR3 (N9782, N9774, N2223, N4657);
or OR2 (N9783, N9782, N5881);
nor NOR3 (N9784, N9763, N1043, N5997);
not NOT1 (N9785, N9779);
xor XOR2 (N9786, N9766, N7556);
or OR3 (N9787, N9783, N4697, N9325);
or OR3 (N9788, N9777, N6006, N6770);
not NOT1 (N9789, N9786);
xor XOR2 (N9790, N9767, N5076);
buf BUF1 (N9791, N9789);
nand NAND4 (N9792, N9784, N7297, N3932, N5827);
buf BUF1 (N9793, N9792);
nor NOR3 (N9794, N9770, N7507, N9633);
xor XOR2 (N9795, N9790, N4808);
xor XOR2 (N9796, N9794, N3773);
or OR2 (N9797, N9788, N620);
nor NOR3 (N9798, N9750, N3717, N8964);
nand NAND2 (N9799, N9787, N3103);
and AND2 (N9800, N9798, N4304);
not NOT1 (N9801, N9800);
or OR2 (N9802, N9797, N3736);
nand NAND2 (N9803, N9785, N1070);
nand NAND2 (N9804, N9803, N9221);
nor NOR4 (N9805, N9801, N7494, N774, N7596);
xor XOR2 (N9806, N9781, N7742);
and AND2 (N9807, N9805, N9506);
and AND2 (N9808, N9791, N1968);
buf BUF1 (N9809, N9780);
nand NAND2 (N9810, N9796, N328);
and AND4 (N9811, N9802, N4011, N9122, N4173);
nor NOR4 (N9812, N9799, N7534, N229, N4234);
and AND4 (N9813, N9806, N2338, N6451, N1388);
and AND4 (N9814, N9811, N4796, N1764, N4012);
and AND2 (N9815, N9793, N2686);
or OR4 (N9816, N9812, N8976, N3802, N5737);
or OR3 (N9817, N9795, N5092, N975);
or OR2 (N9818, N9810, N6240);
and AND2 (N9819, N9818, N4875);
and AND3 (N9820, N9808, N1551, N3917);
buf BUF1 (N9821, N9820);
and AND3 (N9822, N9804, N93, N9667);
nor NOR4 (N9823, N9817, N6515, N7497, N8871);
nand NAND4 (N9824, N9822, N5031, N2531, N5057);
nand NAND4 (N9825, N9819, N9375, N9043, N8135);
xor XOR2 (N9826, N9815, N6555);
buf BUF1 (N9827, N9814);
and AND2 (N9828, N9823, N2264);
xor XOR2 (N9829, N9824, N6793);
xor XOR2 (N9830, N9816, N7174);
xor XOR2 (N9831, N9828, N1171);
buf BUF1 (N9832, N9831);
and AND2 (N9833, N9825, N9284);
and AND2 (N9834, N9813, N7653);
or OR3 (N9835, N9827, N4952, N9194);
and AND2 (N9836, N9832, N849);
or OR2 (N9837, N9835, N6532);
xor XOR2 (N9838, N9821, N6075);
or OR2 (N9839, N9830, N7965);
buf BUF1 (N9840, N9807);
and AND4 (N9841, N9837, N1717, N2947, N6057);
buf BUF1 (N9842, N9829);
buf BUF1 (N9843, N9841);
or OR2 (N9844, N9809, N4422);
xor XOR2 (N9845, N9840, N1758);
nor NOR4 (N9846, N9843, N6611, N8946, N8252);
not NOT1 (N9847, N9839);
buf BUF1 (N9848, N9847);
xor XOR2 (N9849, N9845, N6781);
xor XOR2 (N9850, N9846, N2262);
not NOT1 (N9851, N9849);
xor XOR2 (N9852, N9833, N2675);
or OR2 (N9853, N9844, N7402);
nand NAND4 (N9854, N9852, N7049, N5298, N420);
or OR2 (N9855, N9854, N1548);
xor XOR2 (N9856, N9851, N7290);
or OR2 (N9857, N9856, N5374);
nor NOR4 (N9858, N9850, N5568, N9169, N2736);
or OR4 (N9859, N9853, N2248, N6044, N9008);
and AND2 (N9860, N9842, N5406);
nor NOR4 (N9861, N9834, N7620, N9370, N7598);
nor NOR4 (N9862, N9860, N9785, N27, N5734);
and AND2 (N9863, N9848, N5889);
nor NOR3 (N9864, N9861, N1024, N3505);
or OR3 (N9865, N9862, N7222, N7230);
nor NOR4 (N9866, N9826, N5602, N5275, N8396);
or OR4 (N9867, N9858, N2904, N5766, N3289);
and AND4 (N9868, N9866, N1473, N5440, N7371);
and AND3 (N9869, N9855, N9398, N8855);
buf BUF1 (N9870, N9859);
or OR4 (N9871, N9864, N307, N1660, N5217);
not NOT1 (N9872, N9838);
xor XOR2 (N9873, N9870, N9795);
and AND2 (N9874, N9863, N9050);
nor NOR4 (N9875, N9836, N4343, N2866, N1883);
or OR4 (N9876, N9867, N3771, N5246, N3989);
not NOT1 (N9877, N9876);
and AND3 (N9878, N9874, N3863, N9018);
buf BUF1 (N9879, N9871);
not NOT1 (N9880, N9877);
nand NAND2 (N9881, N9872, N6065);
nor NOR2 (N9882, N9873, N4198);
nand NAND3 (N9883, N9865, N2312, N1358);
nor NOR3 (N9884, N9881, N7145, N6044);
nor NOR3 (N9885, N9884, N1321, N5717);
nand NAND4 (N9886, N9875, N742, N8089, N8499);
nor NOR2 (N9887, N9869, N5464);
xor XOR2 (N9888, N9880, N6776);
and AND3 (N9889, N9878, N4485, N6460);
nor NOR4 (N9890, N9857, N2435, N3855, N2306);
xor XOR2 (N9891, N9885, N1847);
or OR3 (N9892, N9886, N7272, N8777);
xor XOR2 (N9893, N9887, N5508);
xor XOR2 (N9894, N9893, N3766);
not NOT1 (N9895, N9868);
or OR4 (N9896, N9894, N429, N3589, N6996);
and AND3 (N9897, N9896, N8503, N5620);
nor NOR2 (N9898, N9892, N6965);
nand NAND3 (N9899, N9890, N7143, N7971);
and AND3 (N9900, N9899, N4662, N1310);
not NOT1 (N9901, N9898);
xor XOR2 (N9902, N9883, N9180);
nand NAND4 (N9903, N9889, N6442, N5528, N6132);
not NOT1 (N9904, N9903);
and AND3 (N9905, N9895, N2402, N3581);
or OR3 (N9906, N9901, N6251, N3585);
or OR2 (N9907, N9879, N9850);
buf BUF1 (N9908, N9897);
nor NOR2 (N9909, N9906, N4594);
not NOT1 (N9910, N9904);
or OR2 (N9911, N9882, N46);
nor NOR3 (N9912, N9902, N1527, N5197);
not NOT1 (N9913, N9908);
and AND4 (N9914, N9907, N7625, N8881, N5235);
buf BUF1 (N9915, N9905);
buf BUF1 (N9916, N9910);
buf BUF1 (N9917, N9913);
nor NOR3 (N9918, N9914, N6442, N5326);
buf BUF1 (N9919, N9909);
or OR3 (N9920, N9891, N1672, N1383);
not NOT1 (N9921, N9917);
nand NAND2 (N9922, N9920, N9447);
xor XOR2 (N9923, N9918, N1184);
nand NAND2 (N9924, N9922, N3327);
or OR2 (N9925, N9912, N9311);
nand NAND2 (N9926, N9921, N1482);
not NOT1 (N9927, N9915);
and AND4 (N9928, N9925, N3862, N9429, N7978);
buf BUF1 (N9929, N9888);
nor NOR3 (N9930, N9927, N1504, N8244);
nand NAND2 (N9931, N9928, N7217);
and AND2 (N9932, N9919, N8153);
or OR2 (N9933, N9930, N933);
nor NOR2 (N9934, N9924, N1794);
not NOT1 (N9935, N9916);
nand NAND3 (N9936, N9929, N2967, N420);
buf BUF1 (N9937, N9932);
nand NAND2 (N9938, N9933, N7992);
buf BUF1 (N9939, N9935);
nor NOR3 (N9940, N9939, N4317, N6991);
and AND2 (N9941, N9938, N2350);
or OR4 (N9942, N9926, N510, N6565, N6833);
buf BUF1 (N9943, N9942);
nand NAND4 (N9944, N9941, N4676, N5486, N9246);
nor NOR2 (N9945, N9943, N4193);
or OR2 (N9946, N9911, N548);
nor NOR4 (N9947, N9940, N2700, N2070, N6144);
nand NAND4 (N9948, N9931, N4934, N6623, N7166);
nor NOR2 (N9949, N9945, N2329);
or OR2 (N9950, N9936, N8177);
or OR2 (N9951, N9937, N4201);
xor XOR2 (N9952, N9923, N2419);
or OR3 (N9953, N9900, N4175, N4367);
not NOT1 (N9954, N9949);
nor NOR2 (N9955, N9953, N7872);
and AND4 (N9956, N9946, N2838, N8058, N6653);
nand NAND2 (N9957, N9944, N6342);
xor XOR2 (N9958, N9954, N3999);
not NOT1 (N9959, N9956);
xor XOR2 (N9960, N9948, N3860);
buf BUF1 (N9961, N9957);
xor XOR2 (N9962, N9960, N6870);
buf BUF1 (N9963, N9950);
buf BUF1 (N9964, N9947);
not NOT1 (N9965, N9961);
and AND4 (N9966, N9934, N996, N5333, N6508);
or OR2 (N9967, N9959, N9669);
or OR3 (N9968, N9967, N3201, N669);
nor NOR4 (N9969, N9955, N4025, N3350, N6406);
not NOT1 (N9970, N9965);
and AND2 (N9971, N9969, N1075);
or OR2 (N9972, N9952, N8594);
nor NOR3 (N9973, N9966, N8625, N27);
buf BUF1 (N9974, N9958);
or OR4 (N9975, N9964, N5800, N6188, N7300);
and AND2 (N9976, N9963, N4866);
buf BUF1 (N9977, N9970);
or OR3 (N9978, N9976, N1421, N7048);
xor XOR2 (N9979, N9971, N1203);
nor NOR4 (N9980, N9979, N3766, N3670, N6887);
nand NAND2 (N9981, N9975, N2252);
xor XOR2 (N9982, N9977, N501);
nor NOR2 (N9983, N9982, N1487);
nand NAND2 (N9984, N9978, N2614);
or OR4 (N9985, N9951, N6553, N2430, N3680);
and AND2 (N9986, N9973, N9889);
buf BUF1 (N9987, N9968);
nand NAND2 (N9988, N9985, N8868);
not NOT1 (N9989, N9984);
nor NOR2 (N9990, N9987, N4313);
buf BUF1 (N9991, N9972);
xor XOR2 (N9992, N9990, N2835);
or OR3 (N9993, N9989, N7017, N1751);
buf BUF1 (N9994, N9988);
buf BUF1 (N9995, N9986);
or OR3 (N9996, N9962, N3118, N9266);
or OR3 (N9997, N9974, N3479, N3850);
or OR2 (N9998, N9993, N6258);
nand NAND2 (N9999, N9983, N3369);
nor NOR3 (N10000, N9980, N1558, N6879);
nand NAND3 (N10001, N9991, N8850, N7839);
or OR3 (N10002, N9999, N6129, N4021);
nand NAND2 (N10003, N9992, N5804);
or OR3 (N10004, N10001, N141, N4426);
xor XOR2 (N10005, N10003, N9583);
not NOT1 (N10006, N10000);
not NOT1 (N10007, N10002);
and AND2 (N10008, N10005, N8452);
or OR4 (N10009, N10004, N3717, N4792, N381);
xor XOR2 (N10010, N9995, N5655);
nand NAND2 (N10011, N9981, N5688);
nand NAND4 (N10012, N9997, N6947, N8473, N3982);
not NOT1 (N10013, N9998);
xor XOR2 (N10014, N10006, N255);
nor NOR2 (N10015, N10012, N801);
buf BUF1 (N10016, N10011);
nor NOR2 (N10017, N9996, N557);
nand NAND4 (N10018, N10013, N8855, N5293, N9235);
buf BUF1 (N10019, N10008);
xor XOR2 (N10020, N10017, N9318);
or OR2 (N10021, N10010, N6201);
not NOT1 (N10022, N10015);
and AND2 (N10023, N10018, N8200);
nand NAND4 (N10024, N10019, N6203, N7603, N2168);
buf BUF1 (N10025, N10014);
buf BUF1 (N10026, N10023);
nand NAND2 (N10027, N10020, N7819);
not NOT1 (N10028, N10025);
or OR2 (N10029, N10026, N258);
buf BUF1 (N10030, N10009);
xor XOR2 (N10031, N10007, N7913);
nand NAND3 (N10032, N10022, N3574, N5979);
or OR4 (N10033, N10031, N4873, N1382, N4677);
nand NAND4 (N10034, N10016, N6999, N16, N8851);
nor NOR4 (N10035, N10021, N379, N3507, N8426);
nor NOR4 (N10036, N10024, N4089, N8749, N3933);
or OR4 (N10037, N10030, N6326, N8676, N3670);
or OR2 (N10038, N10034, N6344);
buf BUF1 (N10039, N10027);
xor XOR2 (N10040, N10036, N9686);
and AND4 (N10041, N10033, N7673, N6731, N344);
nand NAND3 (N10042, N10038, N3159, N9582);
not NOT1 (N10043, N10037);
nor NOR4 (N10044, N10043, N781, N5678, N5912);
or OR2 (N10045, N10042, N8158);
not NOT1 (N10046, N9994);
not NOT1 (N10047, N10040);
nand NAND3 (N10048, N10047, N7062, N4687);
nand NAND3 (N10049, N10032, N4789, N6518);
and AND2 (N10050, N10048, N6994);
nor NOR4 (N10051, N10041, N2869, N8734, N284);
not NOT1 (N10052, N10044);
or OR2 (N10053, N10029, N2703);
nand NAND4 (N10054, N10053, N1865, N8301, N8047);
nor NOR4 (N10055, N10050, N8083, N7216, N4391);
or OR2 (N10056, N10049, N8417);
and AND4 (N10057, N10054, N8720, N5006, N6745);
xor XOR2 (N10058, N10057, N5929);
nand NAND4 (N10059, N10051, N2546, N5115, N7418);
or OR3 (N10060, N10058, N9616, N3783);
xor XOR2 (N10061, N10055, N3232);
not NOT1 (N10062, N10045);
and AND4 (N10063, N10056, N8132, N4437, N7439);
and AND2 (N10064, N10052, N247);
or OR2 (N10065, N10064, N2101);
not NOT1 (N10066, N10060);
nand NAND4 (N10067, N10039, N4168, N5118, N9955);
nor NOR3 (N10068, N10059, N5636, N1359);
and AND3 (N10069, N10035, N7884, N3466);
and AND3 (N10070, N10028, N3767, N146);
nor NOR4 (N10071, N10069, N5531, N7596, N5057);
nor NOR4 (N10072, N10066, N7965, N6032, N6631);
and AND2 (N10073, N10065, N8846);
not NOT1 (N10074, N10068);
and AND3 (N10075, N10072, N1049, N628);
nor NOR3 (N10076, N10071, N596, N635);
not NOT1 (N10077, N10070);
buf BUF1 (N10078, N10067);
buf BUF1 (N10079, N10075);
nor NOR3 (N10080, N10046, N3558, N7659);
not NOT1 (N10081, N10078);
xor XOR2 (N10082, N10081, N794);
nor NOR3 (N10083, N10080, N47, N9863);
and AND3 (N10084, N10074, N5959, N9780);
and AND3 (N10085, N10061, N1405, N8935);
and AND4 (N10086, N10076, N1337, N4918, N2719);
nor NOR3 (N10087, N10082, N7270, N9230);
and AND3 (N10088, N10077, N9000, N8311);
buf BUF1 (N10089, N10088);
nand NAND3 (N10090, N10063, N1840, N3355);
nand NAND4 (N10091, N10085, N3384, N644, N7209);
not NOT1 (N10092, N10083);
xor XOR2 (N10093, N10089, N4796);
nand NAND2 (N10094, N10086, N2917);
nor NOR4 (N10095, N10062, N6309, N4721, N305);
buf BUF1 (N10096, N10091);
xor XOR2 (N10097, N10096, N2265);
not NOT1 (N10098, N10094);
or OR2 (N10099, N10087, N57);
xor XOR2 (N10100, N10093, N7178);
xor XOR2 (N10101, N10079, N19);
or OR4 (N10102, N10084, N7195, N7260, N1744);
buf BUF1 (N10103, N10098);
and AND2 (N10104, N10097, N1450);
and AND2 (N10105, N10073, N7335);
nor NOR3 (N10106, N10090, N4700, N9428);
and AND3 (N10107, N10104, N6640, N9879);
not NOT1 (N10108, N10099);
or OR3 (N10109, N10108, N469, N4669);
and AND2 (N10110, N10106, N1091);
or OR3 (N10111, N10102, N8640, N6995);
or OR2 (N10112, N10100, N6481);
buf BUF1 (N10113, N10101);
nor NOR4 (N10114, N10105, N2745, N3713, N4540);
nor NOR4 (N10115, N10111, N5738, N942, N5862);
xor XOR2 (N10116, N10103, N10004);
xor XOR2 (N10117, N10095, N841);
or OR3 (N10118, N10115, N1691, N8084);
and AND2 (N10119, N10118, N1949);
buf BUF1 (N10120, N10114);
nand NAND2 (N10121, N10120, N1638);
nand NAND3 (N10122, N10109, N6601, N10000);
xor XOR2 (N10123, N10110, N8739);
nand NAND3 (N10124, N10092, N6055, N4500);
or OR2 (N10125, N10122, N9098);
nand NAND4 (N10126, N10117, N415, N4015, N5385);
not NOT1 (N10127, N10119);
buf BUF1 (N10128, N10125);
or OR4 (N10129, N10126, N6725, N2278, N3659);
not NOT1 (N10130, N10129);
xor XOR2 (N10131, N10127, N6995);
nor NOR2 (N10132, N10124, N309);
xor XOR2 (N10133, N10130, N7344);
or OR4 (N10134, N10123, N4981, N8894, N5205);
nand NAND2 (N10135, N10116, N9419);
buf BUF1 (N10136, N10134);
buf BUF1 (N10137, N10131);
nor NOR2 (N10138, N10107, N6616);
xor XOR2 (N10139, N10132, N6495);
and AND4 (N10140, N10133, N6739, N6612, N8019);
or OR4 (N10141, N10136, N9302, N583, N3583);
nor NOR4 (N10142, N10113, N4145, N667, N8169);
xor XOR2 (N10143, N10137, N2805);
or OR2 (N10144, N10140, N8807);
xor XOR2 (N10145, N10142, N3687);
nand NAND4 (N10146, N10112, N2159, N6344, N7105);
and AND4 (N10147, N10139, N4939, N6428, N5122);
buf BUF1 (N10148, N10128);
not NOT1 (N10149, N10138);
buf BUF1 (N10150, N10148);
and AND3 (N10151, N10135, N3288, N9756);
and AND3 (N10152, N10146, N7783, N582);
or OR2 (N10153, N10145, N6602);
not NOT1 (N10154, N10149);
nand NAND3 (N10155, N10147, N1606, N7304);
nand NAND2 (N10156, N10154, N4099);
not NOT1 (N10157, N10150);
or OR3 (N10158, N10157, N4302, N1369);
not NOT1 (N10159, N10158);
not NOT1 (N10160, N10141);
nand NAND3 (N10161, N10144, N2558, N7683);
buf BUF1 (N10162, N10143);
nand NAND2 (N10163, N10151, N9089);
xor XOR2 (N10164, N10121, N7113);
xor XOR2 (N10165, N10159, N8498);
and AND3 (N10166, N10152, N9368, N7929);
nor NOR2 (N10167, N10166, N175);
xor XOR2 (N10168, N10163, N4936);
buf BUF1 (N10169, N10164);
not NOT1 (N10170, N10156);
or OR2 (N10171, N10155, N2564);
or OR2 (N10172, N10168, N5409);
and AND3 (N10173, N10167, N9886, N3412);
nor NOR3 (N10174, N10171, N1508, N4728);
buf BUF1 (N10175, N10169);
or OR3 (N10176, N10165, N9551, N5203);
and AND3 (N10177, N10170, N8328, N4540);
and AND4 (N10178, N10175, N1329, N5909, N6473);
xor XOR2 (N10179, N10177, N9015);
not NOT1 (N10180, N10173);
xor XOR2 (N10181, N10162, N3761);
and AND2 (N10182, N10161, N7229);
not NOT1 (N10183, N10182);
nor NOR3 (N10184, N10181, N23, N5683);
nor NOR2 (N10185, N10178, N90);
nor NOR3 (N10186, N10179, N6598, N9487);
xor XOR2 (N10187, N10174, N133);
nor NOR3 (N10188, N10153, N5347, N9479);
nor NOR4 (N10189, N10186, N8788, N10081, N251);
not NOT1 (N10190, N10180);
buf BUF1 (N10191, N10188);
and AND4 (N10192, N10191, N3369, N4043, N353);
and AND2 (N10193, N10184, N5323);
or OR2 (N10194, N10189, N960);
not NOT1 (N10195, N10185);
xor XOR2 (N10196, N10193, N2329);
nand NAND4 (N10197, N10172, N9824, N3458, N7901);
nor NOR3 (N10198, N10196, N3842, N2366);
not NOT1 (N10199, N10197);
or OR2 (N10200, N10192, N9089);
buf BUF1 (N10201, N10187);
not NOT1 (N10202, N10190);
nand NAND3 (N10203, N10201, N9234, N6327);
nor NOR3 (N10204, N10176, N7772, N6318);
nand NAND3 (N10205, N10183, N8756, N5729);
xor XOR2 (N10206, N10194, N5312);
or OR2 (N10207, N10198, N9606);
nor NOR2 (N10208, N10199, N5498);
buf BUF1 (N10209, N10207);
not NOT1 (N10210, N10204);
not NOT1 (N10211, N10200);
and AND4 (N10212, N10210, N8078, N3974, N8541);
xor XOR2 (N10213, N10195, N7101);
nand NAND2 (N10214, N10208, N771);
buf BUF1 (N10215, N10205);
not NOT1 (N10216, N10215);
xor XOR2 (N10217, N10213, N6879);
nor NOR3 (N10218, N10202, N8714, N5500);
buf BUF1 (N10219, N10211);
buf BUF1 (N10220, N10217);
nor NOR4 (N10221, N10216, N2438, N9917, N9413);
nand NAND3 (N10222, N10206, N2118, N5862);
or OR3 (N10223, N10203, N3615, N4030);
or OR4 (N10224, N10222, N8164, N689, N8563);
or OR4 (N10225, N10223, N4402, N8686, N3085);
buf BUF1 (N10226, N10209);
nand NAND2 (N10227, N10218, N5270);
nor NOR3 (N10228, N10219, N4692, N1552);
and AND4 (N10229, N10224, N9332, N1965, N6130);
or OR2 (N10230, N10226, N7873);
nor NOR3 (N10231, N10221, N213, N2977);
xor XOR2 (N10232, N10212, N6159);
or OR2 (N10233, N10232, N9869);
xor XOR2 (N10234, N10160, N6113);
nand NAND3 (N10235, N10231, N9419, N6981);
xor XOR2 (N10236, N10220, N1477);
nor NOR3 (N10237, N10214, N279, N5609);
nor NOR3 (N10238, N10229, N9993, N9245);
buf BUF1 (N10239, N10225);
and AND4 (N10240, N10239, N277, N6840, N2453);
buf BUF1 (N10241, N10240);
or OR3 (N10242, N10227, N3755, N4954);
or OR3 (N10243, N10238, N7786, N8973);
not NOT1 (N10244, N10242);
and AND3 (N10245, N10244, N788, N1117);
nand NAND4 (N10246, N10237, N9027, N4579, N4403);
not NOT1 (N10247, N10236);
or OR3 (N10248, N10234, N6501, N4534);
or OR3 (N10249, N10235, N2879, N8377);
xor XOR2 (N10250, N10230, N4162);
or OR4 (N10251, N10228, N286, N4911, N1231);
xor XOR2 (N10252, N10249, N6498);
nand NAND4 (N10253, N10241, N2488, N3372, N5216);
xor XOR2 (N10254, N10245, N6237);
not NOT1 (N10255, N10250);
nand NAND3 (N10256, N10254, N4497, N793);
and AND4 (N10257, N10248, N3787, N5518, N8327);
nor NOR3 (N10258, N10252, N4073, N3797);
nand NAND4 (N10259, N10257, N3666, N7994, N7122);
not NOT1 (N10260, N10251);
or OR4 (N10261, N10253, N3332, N3842, N361);
nand NAND4 (N10262, N10256, N6820, N7406, N4003);
nand NAND2 (N10263, N10260, N4139);
and AND3 (N10264, N10262, N8194, N8074);
and AND2 (N10265, N10233, N4490);
nand NAND4 (N10266, N10243, N3544, N3478, N586);
not NOT1 (N10267, N10258);
xor XOR2 (N10268, N10263, N6674);
or OR4 (N10269, N10264, N10123, N7316, N2527);
or OR4 (N10270, N10247, N9870, N3560, N8937);
nor NOR2 (N10271, N10255, N2095);
buf BUF1 (N10272, N10246);
nand NAND3 (N10273, N10268, N2079, N6005);
buf BUF1 (N10274, N10267);
xor XOR2 (N10275, N10261, N7703);
and AND4 (N10276, N10270, N5884, N10148, N9967);
not NOT1 (N10277, N10265);
nor NOR3 (N10278, N10277, N4593, N193);
buf BUF1 (N10279, N10271);
not NOT1 (N10280, N10276);
or OR3 (N10281, N10259, N3561, N9775);
buf BUF1 (N10282, N10272);
and AND4 (N10283, N10279, N8603, N1324, N9832);
buf BUF1 (N10284, N10274);
or OR4 (N10285, N10284, N7472, N1705, N8017);
and AND3 (N10286, N10275, N4413, N6893);
or OR4 (N10287, N10283, N6774, N148, N7354);
nand NAND3 (N10288, N10269, N7007, N1933);
and AND4 (N10289, N10286, N6571, N3166, N2898);
or OR3 (N10290, N10273, N5686, N982);
buf BUF1 (N10291, N10281);
buf BUF1 (N10292, N10282);
not NOT1 (N10293, N10266);
nand NAND2 (N10294, N10289, N8399);
xor XOR2 (N10295, N10287, N3204);
and AND3 (N10296, N10285, N9626, N950);
or OR3 (N10297, N10288, N4787, N337);
buf BUF1 (N10298, N10280);
or OR3 (N10299, N10291, N8119, N4098);
not NOT1 (N10300, N10278);
nor NOR3 (N10301, N10295, N2284, N6672);
or OR3 (N10302, N10297, N5399, N3498);
buf BUF1 (N10303, N10302);
or OR3 (N10304, N10292, N6578, N6334);
buf BUF1 (N10305, N10290);
or OR2 (N10306, N10298, N4920);
nor NOR2 (N10307, N10300, N707);
and AND3 (N10308, N10296, N4575, N4421);
xor XOR2 (N10309, N10305, N6384);
and AND3 (N10310, N10307, N6727, N2553);
nor NOR2 (N10311, N10310, N7319);
not NOT1 (N10312, N10303);
buf BUF1 (N10313, N10301);
nor NOR2 (N10314, N10309, N8837);
and AND2 (N10315, N10299, N3277);
or OR4 (N10316, N10308, N6967, N7991, N1946);
or OR3 (N10317, N10306, N4725, N1372);
nor NOR3 (N10318, N10304, N201, N7550);
and AND2 (N10319, N10318, N6372);
or OR4 (N10320, N10312, N7994, N2921, N2945);
nand NAND4 (N10321, N10320, N7782, N1368, N8683);
not NOT1 (N10322, N10317);
nand NAND3 (N10323, N10311, N3300, N8195);
xor XOR2 (N10324, N10319, N2115);
xor XOR2 (N10325, N10313, N2891);
nor NOR2 (N10326, N10325, N5018);
xor XOR2 (N10327, N10314, N2570);
and AND2 (N10328, N10316, N493);
nor NOR4 (N10329, N10323, N8757, N8222, N5700);
xor XOR2 (N10330, N10315, N862);
xor XOR2 (N10331, N10293, N1453);
and AND3 (N10332, N10331, N135, N7866);
or OR2 (N10333, N10326, N8649);
xor XOR2 (N10334, N10324, N6136);
buf BUF1 (N10335, N10329);
or OR3 (N10336, N10332, N4965, N4128);
not NOT1 (N10337, N10330);
or OR2 (N10338, N10322, N2853);
nand NAND4 (N10339, N10321, N2519, N372, N3452);
nor NOR3 (N10340, N10335, N948, N3631);
not NOT1 (N10341, N10327);
xor XOR2 (N10342, N10340, N3346);
nand NAND4 (N10343, N10328, N8550, N1445, N8834);
nand NAND3 (N10344, N10333, N5683, N8936);
nor NOR3 (N10345, N10339, N6982, N419);
not NOT1 (N10346, N10341);
or OR3 (N10347, N10345, N4338, N3412);
not NOT1 (N10348, N10347);
nor NOR2 (N10349, N10337, N9675);
and AND3 (N10350, N10338, N2928, N456);
and AND2 (N10351, N10348, N95);
or OR3 (N10352, N10343, N6137, N3398);
nand NAND4 (N10353, N10294, N911, N52, N5275);
nand NAND4 (N10354, N10336, N8715, N10110, N247);
nand NAND2 (N10355, N10334, N545);
and AND2 (N10356, N10354, N6133);
or OR3 (N10357, N10351, N3835, N822);
nand NAND3 (N10358, N10342, N4334, N1999);
nor NOR2 (N10359, N10344, N9031);
xor XOR2 (N10360, N10346, N4103);
and AND2 (N10361, N10353, N4076);
xor XOR2 (N10362, N10359, N977);
not NOT1 (N10363, N10350);
nand NAND3 (N10364, N10360, N1628, N9638);
xor XOR2 (N10365, N10356, N8778);
not NOT1 (N10366, N10364);
and AND2 (N10367, N10355, N3952);
and AND4 (N10368, N10361, N3370, N1776, N6217);
or OR3 (N10369, N10366, N2091, N175);
xor XOR2 (N10370, N10357, N6650);
and AND3 (N10371, N10369, N5174, N6098);
nor NOR4 (N10372, N10370, N429, N6322, N7188);
buf BUF1 (N10373, N10349);
xor XOR2 (N10374, N10358, N10121);
xor XOR2 (N10375, N10367, N7603);
not NOT1 (N10376, N10373);
not NOT1 (N10377, N10376);
buf BUF1 (N10378, N10362);
xor XOR2 (N10379, N10352, N2413);
nor NOR2 (N10380, N10371, N5489);
nor NOR4 (N10381, N10379, N7661, N5290, N186);
not NOT1 (N10382, N10380);
nand NAND4 (N10383, N10381, N3115, N2881, N10364);
nand NAND4 (N10384, N10368, N3527, N6460, N6472);
xor XOR2 (N10385, N10363, N1669);
or OR4 (N10386, N10384, N4987, N6423, N8180);
xor XOR2 (N10387, N10365, N3466);
or OR4 (N10388, N10386, N2329, N5963, N1105);
and AND3 (N10389, N10385, N3688, N8860);
nor NOR3 (N10390, N10375, N9461, N4771);
or OR4 (N10391, N10390, N5717, N3302, N5400);
xor XOR2 (N10392, N10372, N4117);
not NOT1 (N10393, N10388);
nor NOR2 (N10394, N10392, N5780);
and AND4 (N10395, N10382, N3946, N6444, N9049);
buf BUF1 (N10396, N10394);
not NOT1 (N10397, N10378);
not NOT1 (N10398, N10395);
not NOT1 (N10399, N10377);
buf BUF1 (N10400, N10396);
and AND4 (N10401, N10398, N3530, N1232, N898);
nand NAND4 (N10402, N10399, N9981, N5191, N10291);
not NOT1 (N10403, N10389);
xor XOR2 (N10404, N10397, N2767);
not NOT1 (N10405, N10400);
not NOT1 (N10406, N10393);
or OR3 (N10407, N10402, N6563, N3057);
and AND4 (N10408, N10403, N3647, N6541, N3571);
and AND3 (N10409, N10383, N9197, N3813);
nand NAND2 (N10410, N10387, N8660);
and AND2 (N10411, N10409, N9027);
nand NAND4 (N10412, N10407, N3933, N1674, N2490);
or OR3 (N10413, N10391, N1720, N5330);
and AND2 (N10414, N10412, N3853);
and AND4 (N10415, N10410, N5273, N8903, N1960);
buf BUF1 (N10416, N10401);
nand NAND4 (N10417, N10406, N3944, N578, N7579);
not NOT1 (N10418, N10404);
and AND2 (N10419, N10411, N8767);
nand NAND4 (N10420, N10419, N8002, N1389, N1585);
nand NAND4 (N10421, N10408, N3396, N408, N9320);
nand NAND3 (N10422, N10413, N767, N5387);
nand NAND2 (N10423, N10418, N5918);
or OR3 (N10424, N10414, N3746, N4171);
nand NAND3 (N10425, N10416, N8300, N6450);
and AND3 (N10426, N10423, N4187, N2079);
or OR2 (N10427, N10422, N5227);
nor NOR4 (N10428, N10405, N8247, N1274, N9446);
xor XOR2 (N10429, N10421, N2341);
nor NOR2 (N10430, N10426, N8404);
buf BUF1 (N10431, N10417);
not NOT1 (N10432, N10420);
nor NOR2 (N10433, N10430, N9153);
not NOT1 (N10434, N10424);
and AND2 (N10435, N10415, N8567);
or OR3 (N10436, N10425, N3793, N6223);
or OR2 (N10437, N10427, N3705);
nor NOR2 (N10438, N10431, N4149);
and AND2 (N10439, N10374, N2842);
nor NOR3 (N10440, N10429, N9191, N1223);
nand NAND4 (N10441, N10433, N66, N1526, N758);
not NOT1 (N10442, N10440);
nand NAND3 (N10443, N10435, N1322, N7359);
and AND2 (N10444, N10432, N5984);
buf BUF1 (N10445, N10436);
buf BUF1 (N10446, N10441);
nand NAND3 (N10447, N10437, N7621, N4998);
buf BUF1 (N10448, N10434);
nor NOR3 (N10449, N10447, N4364, N4204);
not NOT1 (N10450, N10428);
not NOT1 (N10451, N10446);
nand NAND3 (N10452, N10448, N9313, N5507);
or OR2 (N10453, N10449, N1236);
xor XOR2 (N10454, N10444, N10366);
nand NAND4 (N10455, N10454, N9834, N8078, N8868);
xor XOR2 (N10456, N10452, N3258);
not NOT1 (N10457, N10439);
nand NAND4 (N10458, N10455, N5072, N6418, N10420);
or OR3 (N10459, N10450, N8610, N8163);
and AND2 (N10460, N10458, N3620);
xor XOR2 (N10461, N10451, N7125);
or OR4 (N10462, N10438, N5007, N8785, N3708);
xor XOR2 (N10463, N10457, N9324);
nor NOR3 (N10464, N10442, N4746, N6356);
nand NAND4 (N10465, N10443, N6345, N2705, N1474);
nand NAND3 (N10466, N10460, N7467, N2884);
xor XOR2 (N10467, N10456, N6367);
not NOT1 (N10468, N10466);
xor XOR2 (N10469, N10465, N7945);
not NOT1 (N10470, N10468);
xor XOR2 (N10471, N10463, N5224);
nor NOR2 (N10472, N10470, N6996);
nand NAND4 (N10473, N10461, N203, N1428, N2105);
nor NOR2 (N10474, N10464, N2559);
buf BUF1 (N10475, N10459);
not NOT1 (N10476, N10471);
or OR4 (N10477, N10472, N2587, N9134, N9097);
and AND2 (N10478, N10469, N5178);
nand NAND2 (N10479, N10462, N7934);
or OR4 (N10480, N10479, N2483, N4261, N622);
nor NOR2 (N10481, N10474, N88);
or OR4 (N10482, N10476, N7035, N83, N8710);
xor XOR2 (N10483, N10475, N10051);
or OR2 (N10484, N10467, N5490);
and AND2 (N10485, N10477, N8949);
xor XOR2 (N10486, N10480, N8955);
not NOT1 (N10487, N10445);
xor XOR2 (N10488, N10478, N9779);
not NOT1 (N10489, N10486);
and AND3 (N10490, N10485, N7204, N2583);
or OR2 (N10491, N10482, N8434);
or OR2 (N10492, N10453, N808);
buf BUF1 (N10493, N10491);
nor NOR3 (N10494, N10492, N6766, N152);
and AND2 (N10495, N10490, N9674);
buf BUF1 (N10496, N10489);
xor XOR2 (N10497, N10481, N5509);
nor NOR3 (N10498, N10496, N4591, N8307);
buf BUF1 (N10499, N10493);
xor XOR2 (N10500, N10497, N158);
xor XOR2 (N10501, N10499, N4413);
nor NOR3 (N10502, N10483, N2071, N4016);
not NOT1 (N10503, N10502);
not NOT1 (N10504, N10501);
xor XOR2 (N10505, N10484, N5792);
or OR2 (N10506, N10473, N4684);
or OR4 (N10507, N10498, N8474, N4290, N6484);
nand NAND4 (N10508, N10505, N5160, N1947, N5498);
and AND3 (N10509, N10487, N10204, N3715);
nor NOR4 (N10510, N10500, N6386, N2448, N4742);
nor NOR4 (N10511, N10507, N9443, N9181, N7189);
nor NOR4 (N10512, N10488, N2273, N4582, N1226);
not NOT1 (N10513, N10512);
or OR4 (N10514, N10508, N9556, N9868, N5162);
buf BUF1 (N10515, N10503);
not NOT1 (N10516, N10509);
nor NOR2 (N10517, N10514, N9357);
buf BUF1 (N10518, N10494);
xor XOR2 (N10519, N10518, N5704);
buf BUF1 (N10520, N10506);
and AND3 (N10521, N10516, N6650, N7951);
xor XOR2 (N10522, N10519, N10118);
and AND2 (N10523, N10511, N2036);
xor XOR2 (N10524, N10520, N5334);
xor XOR2 (N10525, N10515, N4862);
buf BUF1 (N10526, N10495);
not NOT1 (N10527, N10510);
xor XOR2 (N10528, N10527, N6186);
nor NOR2 (N10529, N10526, N5212);
buf BUF1 (N10530, N10523);
xor XOR2 (N10531, N10521, N6396);
nand NAND3 (N10532, N10522, N10386, N7777);
or OR2 (N10533, N10504, N2441);
not NOT1 (N10534, N10525);
or OR3 (N10535, N10517, N9644, N8489);
buf BUF1 (N10536, N10528);
or OR3 (N10537, N10536, N3861, N5527);
nand NAND2 (N10538, N10537, N3638);
nor NOR2 (N10539, N10513, N1316);
or OR3 (N10540, N10529, N10046, N2334);
nand NAND2 (N10541, N10524, N5199);
buf BUF1 (N10542, N10530);
not NOT1 (N10543, N10533);
not NOT1 (N10544, N10543);
not NOT1 (N10545, N10539);
nor NOR3 (N10546, N10541, N3851, N3424);
nand NAND4 (N10547, N10545, N4595, N8815, N5045);
and AND2 (N10548, N10534, N2354);
or OR3 (N10549, N10544, N5982, N23);
or OR4 (N10550, N10532, N7182, N9803, N1950);
not NOT1 (N10551, N10531);
xor XOR2 (N10552, N10551, N9356);
xor XOR2 (N10553, N10542, N2479);
buf BUF1 (N10554, N10549);
nand NAND2 (N10555, N10554, N2266);
buf BUF1 (N10556, N10540);
or OR4 (N10557, N10550, N2113, N2097, N6755);
or OR2 (N10558, N10555, N10005);
xor XOR2 (N10559, N10552, N601);
xor XOR2 (N10560, N10553, N7524);
buf BUF1 (N10561, N10546);
and AND2 (N10562, N10559, N7035);
nor NOR4 (N10563, N10548, N4098, N498, N2315);
not NOT1 (N10564, N10535);
not NOT1 (N10565, N10561);
and AND4 (N10566, N10557, N4090, N8158, N3527);
xor XOR2 (N10567, N10558, N8723);
and AND4 (N10568, N10556, N8381, N1704, N7150);
and AND2 (N10569, N10538, N7543);
or OR4 (N10570, N10547, N612, N6534, N2678);
buf BUF1 (N10571, N10568);
nand NAND3 (N10572, N10564, N4599, N3796);
not NOT1 (N10573, N10572);
nand NAND4 (N10574, N10573, N4543, N6676, N5223);
xor XOR2 (N10575, N10574, N7555);
buf BUF1 (N10576, N10569);
nand NAND3 (N10577, N10571, N230, N985);
nand NAND2 (N10578, N10563, N5416);
and AND4 (N10579, N10566, N8537, N3592, N3241);
nor NOR3 (N10580, N10560, N5996, N4922);
xor XOR2 (N10581, N10562, N934);
and AND3 (N10582, N10570, N4412, N943);
xor XOR2 (N10583, N10579, N9857);
nor NOR3 (N10584, N10581, N5090, N8849);
or OR4 (N10585, N10567, N5865, N4037, N7071);
or OR4 (N10586, N10565, N5104, N10441, N5888);
nand NAND2 (N10587, N10577, N8131);
xor XOR2 (N10588, N10586, N614);
not NOT1 (N10589, N10587);
and AND2 (N10590, N10588, N4298);
or OR3 (N10591, N10580, N2236, N2300);
nand NAND2 (N10592, N10584, N4046);
buf BUF1 (N10593, N10585);
nand NAND2 (N10594, N10575, N4720);
nor NOR4 (N10595, N10589, N9028, N5442, N5976);
xor XOR2 (N10596, N10578, N1220);
or OR4 (N10597, N10592, N3640, N8256, N7151);
not NOT1 (N10598, N10596);
nor NOR2 (N10599, N10593, N1360);
buf BUF1 (N10600, N10576);
nand NAND4 (N10601, N10598, N6150, N3747, N2488);
or OR4 (N10602, N10594, N3492, N9527, N3430);
nor NOR2 (N10603, N10600, N263);
or OR3 (N10604, N10603, N216, N6537);
and AND4 (N10605, N10597, N4608, N8626, N7253);
nor NOR4 (N10606, N10591, N4246, N9714, N159);
nand NAND3 (N10607, N10606, N7667, N10074);
xor XOR2 (N10608, N10590, N10000);
or OR3 (N10609, N10607, N3256, N2696);
nor NOR2 (N10610, N10601, N736);
or OR3 (N10611, N10602, N4738, N10167);
or OR2 (N10612, N10609, N1798);
nand NAND3 (N10613, N10610, N10209, N3248);
nor NOR2 (N10614, N10599, N3704);
buf BUF1 (N10615, N10605);
and AND2 (N10616, N10604, N3536);
or OR3 (N10617, N10615, N9299, N8538);
and AND2 (N10618, N10608, N8911);
or OR2 (N10619, N10616, N9678);
nor NOR3 (N10620, N10583, N9400, N6117);
not NOT1 (N10621, N10620);
buf BUF1 (N10622, N10619);
nand NAND2 (N10623, N10613, N1823);
nand NAND2 (N10624, N10618, N5815);
xor XOR2 (N10625, N10614, N10028);
nor NOR2 (N10626, N10582, N4062);
buf BUF1 (N10627, N10624);
or OR2 (N10628, N10626, N4373);
nand NAND2 (N10629, N10611, N5412);
or OR3 (N10630, N10627, N376, N9635);
and AND2 (N10631, N10595, N2246);
or OR4 (N10632, N10631, N2544, N7341, N801);
not NOT1 (N10633, N10625);
or OR2 (N10634, N10623, N2073);
nor NOR3 (N10635, N10634, N5738, N10518);
nand NAND4 (N10636, N10629, N1524, N8154, N10108);
nor NOR2 (N10637, N10636, N3960);
nor NOR2 (N10638, N10622, N8015);
buf BUF1 (N10639, N10632);
nor NOR3 (N10640, N10633, N1119, N3895);
xor XOR2 (N10641, N10621, N4339);
or OR2 (N10642, N10617, N3260);
and AND3 (N10643, N10642, N4865, N3482);
nand NAND3 (N10644, N10630, N5705, N805);
not NOT1 (N10645, N10640);
nand NAND3 (N10646, N10639, N6817, N6656);
or OR4 (N10647, N10641, N7274, N4428, N4474);
or OR3 (N10648, N10645, N9316, N7625);
xor XOR2 (N10649, N10638, N6415);
nand NAND2 (N10650, N10643, N3471);
xor XOR2 (N10651, N10646, N4525);
and AND3 (N10652, N10647, N296, N9933);
buf BUF1 (N10653, N10637);
nor NOR2 (N10654, N10653, N6914);
buf BUF1 (N10655, N10612);
xor XOR2 (N10656, N10635, N9480);
and AND2 (N10657, N10628, N243);
and AND4 (N10658, N10651, N6424, N669, N10349);
nor NOR2 (N10659, N10654, N9494);
not NOT1 (N10660, N10657);
nand NAND2 (N10661, N10655, N6359);
not NOT1 (N10662, N10650);
or OR3 (N10663, N10658, N2766, N7040);
buf BUF1 (N10664, N10649);
buf BUF1 (N10665, N10660);
nand NAND2 (N10666, N10659, N8610);
nand NAND2 (N10667, N10661, N9431);
nor NOR4 (N10668, N10666, N4780, N9627, N5832);
or OR2 (N10669, N10648, N1882);
nor NOR2 (N10670, N10663, N2585);
or OR2 (N10671, N10668, N5855);
nand NAND3 (N10672, N10656, N6560, N9690);
nand NAND2 (N10673, N10671, N9548);
not NOT1 (N10674, N10669);
nand NAND4 (N10675, N10665, N6579, N6607, N899);
not NOT1 (N10676, N10674);
not NOT1 (N10677, N10667);
and AND4 (N10678, N10652, N3050, N3379, N1855);
not NOT1 (N10679, N10644);
or OR4 (N10680, N10677, N7022, N1910, N7219);
buf BUF1 (N10681, N10679);
nand NAND4 (N10682, N10664, N7436, N9091, N2748);
or OR2 (N10683, N10673, N2085);
or OR3 (N10684, N10675, N4498, N7894);
and AND4 (N10685, N10682, N5429, N5882, N375);
buf BUF1 (N10686, N10683);
buf BUF1 (N10687, N10678);
not NOT1 (N10688, N10680);
buf BUF1 (N10689, N10685);
or OR3 (N10690, N10670, N3182, N282);
not NOT1 (N10691, N10688);
nor NOR4 (N10692, N10687, N1986, N5380, N8002);
and AND4 (N10693, N10681, N10230, N5045, N2131);
and AND2 (N10694, N10686, N1616);
and AND2 (N10695, N10691, N4902);
buf BUF1 (N10696, N10672);
or OR4 (N10697, N10694, N6705, N10315, N9211);
not NOT1 (N10698, N10697);
nand NAND3 (N10699, N10693, N2865, N5598);
xor XOR2 (N10700, N10676, N6635);
buf BUF1 (N10701, N10700);
nand NAND3 (N10702, N10695, N1981, N7497);
nand NAND2 (N10703, N10701, N3534);
nor NOR3 (N10704, N10698, N984, N6251);
not NOT1 (N10705, N10689);
not NOT1 (N10706, N10662);
and AND2 (N10707, N10684, N5239);
or OR2 (N10708, N10707, N4965);
xor XOR2 (N10709, N10699, N5420);
nand NAND3 (N10710, N10690, N9395, N2493);
buf BUF1 (N10711, N10710);
not NOT1 (N10712, N10711);
buf BUF1 (N10713, N10705);
not NOT1 (N10714, N10703);
buf BUF1 (N10715, N10712);
xor XOR2 (N10716, N10696, N8899);
nor NOR3 (N10717, N10715, N9773, N8508);
and AND4 (N10718, N10714, N8339, N4140, N7251);
and AND4 (N10719, N10709, N834, N8584, N9615);
not NOT1 (N10720, N10702);
nand NAND4 (N10721, N10708, N4498, N3412, N1266);
or OR4 (N10722, N10713, N6215, N2235, N781);
xor XOR2 (N10723, N10692, N3926);
buf BUF1 (N10724, N10716);
not NOT1 (N10725, N10723);
and AND2 (N10726, N10706, N4262);
xor XOR2 (N10727, N10724, N8448);
buf BUF1 (N10728, N10721);
nor NOR4 (N10729, N10722, N8427, N4323, N8486);
xor XOR2 (N10730, N10704, N1519);
nor NOR2 (N10731, N10719, N5340);
xor XOR2 (N10732, N10717, N4762);
and AND3 (N10733, N10729, N7091, N6323);
nor NOR2 (N10734, N10726, N9785);
not NOT1 (N10735, N10731);
or OR3 (N10736, N10735, N1877, N10073);
or OR3 (N10737, N10734, N3143, N7106);
and AND3 (N10738, N10736, N3348, N1403);
not NOT1 (N10739, N10718);
nor NOR2 (N10740, N10727, N3797);
and AND4 (N10741, N10738, N2665, N1315, N9144);
or OR4 (N10742, N10739, N7765, N2775, N7539);
nand NAND3 (N10743, N10732, N5195, N9820);
xor XOR2 (N10744, N10741, N320);
and AND4 (N10745, N10720, N9836, N4854, N6031);
buf BUF1 (N10746, N10730);
nor NOR3 (N10747, N10737, N3580, N4774);
or OR2 (N10748, N10740, N3069);
not NOT1 (N10749, N10747);
nor NOR2 (N10750, N10748, N8667);
or OR2 (N10751, N10743, N295);
nor NOR2 (N10752, N10750, N10631);
or OR4 (N10753, N10728, N7604, N10317, N6369);
nand NAND4 (N10754, N10742, N629, N6070, N888);
buf BUF1 (N10755, N10733);
not NOT1 (N10756, N10753);
xor XOR2 (N10757, N10752, N1635);
nor NOR2 (N10758, N10754, N4941);
or OR3 (N10759, N10756, N9370, N10453);
nor NOR3 (N10760, N10746, N87, N2448);
not NOT1 (N10761, N10755);
xor XOR2 (N10762, N10725, N10761);
or OR4 (N10763, N1961, N3960, N5453, N8836);
nand NAND3 (N10764, N10757, N2301, N4855);
or OR3 (N10765, N10744, N2057, N6029);
xor XOR2 (N10766, N10760, N7947);
nand NAND2 (N10767, N10745, N8596);
not NOT1 (N10768, N10766);
not NOT1 (N10769, N10751);
buf BUF1 (N10770, N10769);
nand NAND2 (N10771, N10765, N9476);
xor XOR2 (N10772, N10768, N9146);
nor NOR2 (N10773, N10771, N2456);
xor XOR2 (N10774, N10749, N9651);
nor NOR4 (N10775, N10773, N2066, N3312, N955);
buf BUF1 (N10776, N10775);
and AND3 (N10777, N10776, N7795, N5052);
and AND3 (N10778, N10763, N6327, N7341);
xor XOR2 (N10779, N10774, N29);
xor XOR2 (N10780, N10758, N8300);
buf BUF1 (N10781, N10779);
not NOT1 (N10782, N10781);
or OR4 (N10783, N10759, N1301, N5279, N8134);
or OR2 (N10784, N10767, N5056);
and AND3 (N10785, N10762, N7534, N5425);
nor NOR3 (N10786, N10770, N1955, N448);
or OR2 (N10787, N10783, N3131);
nand NAND3 (N10788, N10778, N8502, N5641);
not NOT1 (N10789, N10780);
nor NOR2 (N10790, N10788, N1295);
nand NAND4 (N10791, N10772, N7568, N8994, N4912);
not NOT1 (N10792, N10777);
nand NAND4 (N10793, N10787, N10219, N4833, N5947);
or OR2 (N10794, N10786, N2787);
buf BUF1 (N10795, N10792);
and AND3 (N10796, N10795, N660, N4381);
not NOT1 (N10797, N10790);
xor XOR2 (N10798, N10794, N6121);
xor XOR2 (N10799, N10796, N10768);
and AND4 (N10800, N10793, N4149, N5070, N5331);
nor NOR4 (N10801, N10782, N6255, N3606, N9595);
nand NAND4 (N10802, N10784, N6132, N10684, N5155);
xor XOR2 (N10803, N10785, N8455);
xor XOR2 (N10804, N10798, N2439);
or OR4 (N10805, N10789, N3603, N2208, N761);
and AND4 (N10806, N10803, N1262, N787, N10006);
and AND2 (N10807, N10806, N4336);
and AND2 (N10808, N10800, N10739);
and AND2 (N10809, N10808, N8269);
nand NAND3 (N10810, N10791, N1576, N6581);
or OR3 (N10811, N10809, N1989, N357);
nor NOR4 (N10812, N10811, N834, N1249, N9644);
buf BUF1 (N10813, N10807);
or OR2 (N10814, N10810, N8625);
nor NOR4 (N10815, N10813, N3392, N6408, N9036);
and AND2 (N10816, N10801, N1413);
or OR3 (N10817, N10764, N3811, N8660);
and AND4 (N10818, N10799, N7807, N4016, N4836);
nor NOR2 (N10819, N10805, N2733);
xor XOR2 (N10820, N10797, N9207);
or OR3 (N10821, N10817, N4273, N4354);
or OR2 (N10822, N10818, N2649);
buf BUF1 (N10823, N10819);
nand NAND2 (N10824, N10812, N6498);
nand NAND2 (N10825, N10804, N8251);
nand NAND4 (N10826, N10821, N9325, N10348, N3608);
nand NAND3 (N10827, N10816, N8227, N10787);
not NOT1 (N10828, N10822);
nand NAND4 (N10829, N10823, N2348, N967, N9711);
buf BUF1 (N10830, N10820);
nand NAND4 (N10831, N10826, N8097, N9320, N9981);
nor NOR2 (N10832, N10802, N1925);
buf BUF1 (N10833, N10828);
buf BUF1 (N10834, N10815);
or OR3 (N10835, N10831, N4457, N9797);
xor XOR2 (N10836, N10834, N8213);
and AND3 (N10837, N10835, N10681, N6696);
or OR4 (N10838, N10829, N3635, N5683, N1954);
buf BUF1 (N10839, N10832);
or OR4 (N10840, N10824, N5748, N7452, N3734);
nor NOR4 (N10841, N10840, N6520, N44, N3336);
buf BUF1 (N10842, N10825);
not NOT1 (N10843, N10827);
nor NOR4 (N10844, N10839, N9848, N9276, N6760);
or OR3 (N10845, N10836, N8987, N8232);
or OR4 (N10846, N10837, N10000, N7476, N645);
buf BUF1 (N10847, N10814);
xor XOR2 (N10848, N10830, N3403);
buf BUF1 (N10849, N10845);
xor XOR2 (N10850, N10849, N7363);
xor XOR2 (N10851, N10841, N7261);
nor NOR4 (N10852, N10846, N5593, N3324, N823);
and AND3 (N10853, N10844, N6974, N2022);
and AND4 (N10854, N10843, N9851, N9291, N1356);
and AND4 (N10855, N10851, N9592, N5855, N7044);
not NOT1 (N10856, N10854);
xor XOR2 (N10857, N10833, N976);
buf BUF1 (N10858, N10850);
nor NOR3 (N10859, N10858, N5645, N5466);
and AND4 (N10860, N10838, N4347, N2756, N6854);
not NOT1 (N10861, N10842);
nand NAND4 (N10862, N10853, N1562, N7758, N1251);
not NOT1 (N10863, N10855);
buf BUF1 (N10864, N10848);
and AND2 (N10865, N10856, N526);
and AND2 (N10866, N10861, N5317);
and AND4 (N10867, N10860, N1772, N5037, N1253);
and AND4 (N10868, N10852, N10060, N3981, N8286);
nand NAND3 (N10869, N10864, N7786, N1563);
xor XOR2 (N10870, N10865, N435);
not NOT1 (N10871, N10863);
and AND2 (N10872, N10867, N8853);
nand NAND3 (N10873, N10869, N5951, N1910);
or OR2 (N10874, N10872, N5968);
and AND4 (N10875, N10868, N9855, N3670, N4300);
not NOT1 (N10876, N10870);
buf BUF1 (N10877, N10847);
not NOT1 (N10878, N10857);
not NOT1 (N10879, N10871);
nand NAND4 (N10880, N10875, N10568, N1657, N4140);
buf BUF1 (N10881, N10880);
xor XOR2 (N10882, N10859, N2376);
nor NOR3 (N10883, N10874, N9980, N8544);
nand NAND4 (N10884, N10873, N6093, N3311, N5832);
buf BUF1 (N10885, N10882);
nand NAND4 (N10886, N10877, N7379, N3136, N4558);
not NOT1 (N10887, N10885);
and AND4 (N10888, N10887, N6772, N9784, N8775);
or OR4 (N10889, N10888, N1416, N8636, N6184);
xor XOR2 (N10890, N10881, N599);
buf BUF1 (N10891, N10883);
and AND4 (N10892, N10876, N5692, N410, N2734);
nor NOR2 (N10893, N10890, N4460);
not NOT1 (N10894, N10891);
nand NAND3 (N10895, N10862, N3238, N562);
nand NAND2 (N10896, N10886, N6656);
nand NAND4 (N10897, N10889, N2953, N930, N9662);
or OR3 (N10898, N10894, N770, N5841);
xor XOR2 (N10899, N10897, N7234);
not NOT1 (N10900, N10893);
buf BUF1 (N10901, N10899);
xor XOR2 (N10902, N10895, N4889);
or OR3 (N10903, N10902, N8469, N9243);
xor XOR2 (N10904, N10892, N8676);
or OR4 (N10905, N10878, N5044, N4644, N8099);
nand NAND4 (N10906, N10904, N10295, N8508, N4454);
nand NAND3 (N10907, N10906, N3123, N454);
xor XOR2 (N10908, N10866, N3525);
nand NAND3 (N10909, N10896, N415, N4284);
or OR4 (N10910, N10898, N397, N5504, N3816);
buf BUF1 (N10911, N10901);
nand NAND3 (N10912, N10884, N3461, N304);
xor XOR2 (N10913, N10900, N7408);
nor NOR4 (N10914, N10909, N6446, N3592, N4008);
not NOT1 (N10915, N10910);
and AND4 (N10916, N10913, N5084, N1692, N847);
nand NAND4 (N10917, N10908, N6270, N6404, N844);
not NOT1 (N10918, N10917);
buf BUF1 (N10919, N10903);
nand NAND2 (N10920, N10915, N10155);
and AND3 (N10921, N10907, N6491, N653);
or OR3 (N10922, N10918, N8023, N3316);
nand NAND4 (N10923, N10879, N5926, N5571, N7925);
nor NOR2 (N10924, N10920, N3574);
buf BUF1 (N10925, N10922);
not NOT1 (N10926, N10916);
xor XOR2 (N10927, N10925, N6108);
not NOT1 (N10928, N10914);
or OR3 (N10929, N10911, N6051, N876);
or OR2 (N10930, N10927, N907);
or OR4 (N10931, N10930, N10311, N769, N1407);
nand NAND3 (N10932, N10929, N7674, N1260);
or OR3 (N10933, N10912, N1828, N6009);
and AND2 (N10934, N10919, N6264);
not NOT1 (N10935, N10932);
and AND4 (N10936, N10921, N2497, N6628, N616);
or OR2 (N10937, N10905, N936);
and AND2 (N10938, N10934, N9493);
not NOT1 (N10939, N10938);
or OR3 (N10940, N10935, N2130, N2610);
nand NAND3 (N10941, N10926, N9383, N4215);
buf BUF1 (N10942, N10924);
and AND3 (N10943, N10933, N81, N2702);
buf BUF1 (N10944, N10943);
nand NAND2 (N10945, N10944, N3954);
or OR3 (N10946, N10931, N2469, N273);
nor NOR2 (N10947, N10939, N4041);
nor NOR3 (N10948, N10945, N8890, N1151);
and AND2 (N10949, N10947, N4835);
not NOT1 (N10950, N10936);
not NOT1 (N10951, N10946);
and AND2 (N10952, N10942, N2198);
and AND4 (N10953, N10928, N6657, N9595, N2292);
or OR3 (N10954, N10923, N419, N2253);
xor XOR2 (N10955, N10949, N6854);
buf BUF1 (N10956, N10952);
not NOT1 (N10957, N10953);
or OR4 (N10958, N10951, N6437, N4733, N3536);
nor NOR3 (N10959, N10958, N6293, N5360);
and AND4 (N10960, N10937, N8303, N8902, N9450);
buf BUF1 (N10961, N10940);
xor XOR2 (N10962, N10950, N1106);
and AND3 (N10963, N10957, N5072, N5448);
nor NOR2 (N10964, N10962, N5307);
nand NAND2 (N10965, N10956, N8282);
or OR3 (N10966, N10961, N6809, N2793);
nor NOR2 (N10967, N10963, N10476);
not NOT1 (N10968, N10941);
nor NOR3 (N10969, N10960, N882, N3704);
not NOT1 (N10970, N10948);
and AND4 (N10971, N10964, N10248, N9489, N7415);
and AND4 (N10972, N10967, N5977, N927, N9148);
nand NAND2 (N10973, N10971, N5548);
nand NAND2 (N10974, N10965, N869);
xor XOR2 (N10975, N10954, N10294);
buf BUF1 (N10976, N10955);
not NOT1 (N10977, N10973);
and AND4 (N10978, N10970, N5167, N8678, N2187);
nor NOR4 (N10979, N10966, N8695, N10313, N8435);
or OR4 (N10980, N10969, N5277, N10165, N5535);
and AND3 (N10981, N10974, N34, N10405);
xor XOR2 (N10982, N10972, N9894);
and AND3 (N10983, N10980, N9069, N6164);
buf BUF1 (N10984, N10976);
nor NOR4 (N10985, N10983, N10983, N8631, N10125);
buf BUF1 (N10986, N10985);
not NOT1 (N10987, N10982);
nor NOR4 (N10988, N10984, N9782, N4998, N3038);
buf BUF1 (N10989, N10977);
or OR4 (N10990, N10959, N4867, N2528, N5649);
not NOT1 (N10991, N10986);
nor NOR2 (N10992, N10981, N10712);
buf BUF1 (N10993, N10979);
buf BUF1 (N10994, N10968);
nor NOR3 (N10995, N10975, N9140, N4064);
nand NAND2 (N10996, N10992, N6493);
nor NOR4 (N10997, N10978, N8412, N7826, N7806);
nand NAND2 (N10998, N10993, N7517);
not NOT1 (N10999, N10989);
nor NOR3 (N11000, N10998, N7584, N1589);
or OR3 (N11001, N10987, N9460, N7845);
buf BUF1 (N11002, N10990);
nor NOR4 (N11003, N11000, N6149, N3775, N7988);
and AND2 (N11004, N10999, N9048);
xor XOR2 (N11005, N11001, N1405);
buf BUF1 (N11006, N11003);
and AND4 (N11007, N10991, N1612, N2636, N3187);
or OR4 (N11008, N10988, N8824, N1385, N5254);
buf BUF1 (N11009, N11006);
not NOT1 (N11010, N11005);
and AND4 (N11011, N11007, N4769, N2318, N4044);
nand NAND2 (N11012, N11008, N7845);
or OR4 (N11013, N11004, N10055, N6121, N8208);
xor XOR2 (N11014, N11009, N7860);
xor XOR2 (N11015, N11011, N5007);
nor NOR4 (N11016, N11010, N8293, N9123, N3304);
or OR2 (N11017, N11016, N5451);
nor NOR2 (N11018, N11015, N6991);
xor XOR2 (N11019, N10995, N6078);
buf BUF1 (N11020, N11012);
and AND2 (N11021, N11019, N1200);
xor XOR2 (N11022, N10994, N5409);
and AND2 (N11023, N11021, N7337);
xor XOR2 (N11024, N11020, N7894);
nor NOR4 (N11025, N11024, N9425, N8914, N7694);
or OR3 (N11026, N11025, N7954, N971);
or OR2 (N11027, N11002, N5820);
nor NOR4 (N11028, N11026, N199, N8090, N8053);
or OR2 (N11029, N10996, N3756);
nand NAND4 (N11030, N11027, N3394, N7064, N8687);
not NOT1 (N11031, N11022);
xor XOR2 (N11032, N11018, N1314);
nand NAND3 (N11033, N11014, N3041, N5146);
nor NOR4 (N11034, N11023, N1734, N7992, N654);
nor NOR3 (N11035, N11032, N10031, N10392);
or OR3 (N11036, N11013, N10264, N8002);
or OR3 (N11037, N11031, N10286, N6545);
and AND3 (N11038, N10997, N9811, N5375);
not NOT1 (N11039, N11034);
and AND4 (N11040, N11029, N5156, N10087, N10591);
not NOT1 (N11041, N11039);
not NOT1 (N11042, N11038);
nand NAND4 (N11043, N11035, N1298, N8522, N2404);
nor NOR2 (N11044, N11036, N3471);
and AND4 (N11045, N11041, N10892, N5565, N9478);
nor NOR2 (N11046, N11033, N9900);
nand NAND3 (N11047, N11028, N2696, N9713);
nand NAND4 (N11048, N11017, N6754, N7334, N10024);
nand NAND3 (N11049, N11043, N6351, N10585);
buf BUF1 (N11050, N11044);
buf BUF1 (N11051, N11049);
not NOT1 (N11052, N11042);
xor XOR2 (N11053, N11050, N5193);
and AND4 (N11054, N11047, N2581, N5220, N4270);
xor XOR2 (N11055, N11030, N2592);
nor NOR2 (N11056, N11040, N9930);
not NOT1 (N11057, N11048);
and AND2 (N11058, N11057, N138);
or OR2 (N11059, N11056, N5905);
nand NAND3 (N11060, N11058, N9298, N5451);
or OR3 (N11061, N11052, N3495, N2387);
not NOT1 (N11062, N11061);
and AND4 (N11063, N11060, N10009, N1976, N7632);
buf BUF1 (N11064, N11059);
or OR3 (N11065, N11055, N135, N1897);
nand NAND3 (N11066, N11063, N5293, N651);
nand NAND2 (N11067, N11037, N10135);
or OR3 (N11068, N11046, N1971, N9933);
buf BUF1 (N11069, N11062);
nand NAND2 (N11070, N11066, N7586);
nand NAND3 (N11071, N11053, N4663, N3479);
nor NOR3 (N11072, N11045, N7664, N8016);
nor NOR4 (N11073, N11070, N2276, N3550, N8548);
xor XOR2 (N11074, N11054, N3472);
or OR2 (N11075, N11069, N4638);
nor NOR3 (N11076, N11065, N6384, N6262);
or OR4 (N11077, N11071, N2728, N8331, N2990);
nand NAND3 (N11078, N11077, N2897, N9970);
or OR2 (N11079, N11078, N6621);
not NOT1 (N11080, N11067);
not NOT1 (N11081, N11072);
xor XOR2 (N11082, N11081, N5899);
xor XOR2 (N11083, N11051, N2367);
not NOT1 (N11084, N11080);
nor NOR2 (N11085, N11083, N6038);
not NOT1 (N11086, N11075);
buf BUF1 (N11087, N11086);
or OR4 (N11088, N11079, N1746, N1205, N2448);
nor NOR3 (N11089, N11076, N5905, N1157);
or OR2 (N11090, N11088, N3755);
nor NOR2 (N11091, N11068, N5049);
nor NOR4 (N11092, N11091, N1254, N2607, N6391);
buf BUF1 (N11093, N11084);
xor XOR2 (N11094, N11089, N1538);
xor XOR2 (N11095, N11087, N3083);
buf BUF1 (N11096, N11092);
or OR2 (N11097, N11096, N5056);
and AND4 (N11098, N11097, N108, N2773, N3596);
and AND3 (N11099, N11094, N6990, N9541);
not NOT1 (N11100, N11064);
and AND2 (N11101, N11098, N8497);
nor NOR4 (N11102, N11090, N3497, N3689, N8911);
not NOT1 (N11103, N11093);
nor NOR2 (N11104, N11095, N3031);
buf BUF1 (N11105, N11103);
not NOT1 (N11106, N11073);
or OR2 (N11107, N11106, N4976);
nand NAND2 (N11108, N11099, N9079);
nand NAND4 (N11109, N11101, N4686, N4593, N69);
and AND4 (N11110, N11107, N1524, N5188, N817);
nor NOR3 (N11111, N11102, N1084, N345);
xor XOR2 (N11112, N11082, N1883);
not NOT1 (N11113, N11104);
nand NAND4 (N11114, N11112, N8168, N1980, N10939);
not NOT1 (N11115, N11109);
nor NOR3 (N11116, N11100, N10285, N3360);
buf BUF1 (N11117, N11108);
and AND4 (N11118, N11113, N6486, N4148, N2086);
or OR3 (N11119, N11105, N9110, N10270);
buf BUF1 (N11120, N11118);
xor XOR2 (N11121, N11116, N2256);
or OR4 (N11122, N11117, N6725, N6014, N2752);
or OR4 (N11123, N11085, N8703, N2993, N4883);
buf BUF1 (N11124, N11115);
xor XOR2 (N11125, N11123, N2678);
buf BUF1 (N11126, N11124);
nor NOR3 (N11127, N11111, N3907, N2514);
buf BUF1 (N11128, N11120);
nand NAND3 (N11129, N11114, N8601, N170);
buf BUF1 (N11130, N11119);
nand NAND2 (N11131, N11122, N7695);
not NOT1 (N11132, N11110);
and AND2 (N11133, N11126, N1776);
nand NAND2 (N11134, N11133, N1448);
not NOT1 (N11135, N11130);
buf BUF1 (N11136, N11135);
buf BUF1 (N11137, N11129);
nand NAND4 (N11138, N11132, N11041, N4036, N8503);
xor XOR2 (N11139, N11138, N3374);
nand NAND2 (N11140, N11131, N5383);
not NOT1 (N11141, N11127);
nand NAND3 (N11142, N11136, N4043, N1683);
not NOT1 (N11143, N11074);
buf BUF1 (N11144, N11137);
xor XOR2 (N11145, N11142, N4773);
and AND4 (N11146, N11134, N7690, N3718, N3192);
buf BUF1 (N11147, N11128);
xor XOR2 (N11148, N11145, N6680);
xor XOR2 (N11149, N11146, N6113);
or OR3 (N11150, N11147, N7175, N5540);
xor XOR2 (N11151, N11148, N10618);
and AND3 (N11152, N11144, N2628, N4496);
nand NAND4 (N11153, N11150, N4188, N8821, N1396);
xor XOR2 (N11154, N11141, N5988);
not NOT1 (N11155, N11153);
or OR4 (N11156, N11121, N2577, N2733, N5146);
nand NAND4 (N11157, N11139, N2221, N9331, N5925);
nand NAND2 (N11158, N11157, N6259);
or OR4 (N11159, N11156, N112, N355, N9936);
xor XOR2 (N11160, N11149, N5743);
not NOT1 (N11161, N11160);
and AND3 (N11162, N11158, N5788, N1211);
xor XOR2 (N11163, N11155, N7729);
and AND2 (N11164, N11163, N731);
and AND3 (N11165, N11162, N7462, N6113);
xor XOR2 (N11166, N11151, N7058);
and AND2 (N11167, N11164, N505);
or OR2 (N11168, N11167, N7104);
nor NOR3 (N11169, N11166, N10011, N6064);
buf BUF1 (N11170, N11143);
nand NAND3 (N11171, N11170, N5858, N9234);
nand NAND4 (N11172, N11125, N723, N6922, N5090);
nand NAND2 (N11173, N11165, N10665);
nor NOR3 (N11174, N11172, N992, N5496);
and AND4 (N11175, N11152, N9175, N6154, N9419);
xor XOR2 (N11176, N11140, N10864);
and AND4 (N11177, N11171, N889, N7736, N9286);
not NOT1 (N11178, N11174);
not NOT1 (N11179, N11175);
xor XOR2 (N11180, N11177, N30);
buf BUF1 (N11181, N11168);
nand NAND2 (N11182, N11169, N5875);
or OR3 (N11183, N11178, N3382, N8587);
or OR3 (N11184, N11154, N1028, N1902);
xor XOR2 (N11185, N11184, N3460);
nor NOR2 (N11186, N11161, N4544);
nor NOR4 (N11187, N11186, N5185, N10332, N8918);
buf BUF1 (N11188, N11182);
nand NAND2 (N11189, N11159, N9293);
not NOT1 (N11190, N11181);
not NOT1 (N11191, N11173);
nor NOR2 (N11192, N11188, N11009);
nand NAND2 (N11193, N11176, N8011);
not NOT1 (N11194, N11185);
and AND3 (N11195, N11180, N8191, N6480);
or OR4 (N11196, N11187, N1904, N4010, N8409);
nand NAND4 (N11197, N11183, N10769, N5557, N8901);
not NOT1 (N11198, N11192);
xor XOR2 (N11199, N11198, N5674);
nor NOR2 (N11200, N11196, N193);
not NOT1 (N11201, N11200);
nand NAND3 (N11202, N11194, N5030, N4718);
or OR2 (N11203, N11190, N9009);
nor NOR4 (N11204, N11197, N5565, N3385, N5823);
nand NAND2 (N11205, N11199, N10345);
and AND2 (N11206, N11205, N3423);
nor NOR4 (N11207, N11193, N2050, N8441, N10766);
xor XOR2 (N11208, N11179, N5545);
xor XOR2 (N11209, N11208, N11180);
xor XOR2 (N11210, N11203, N6045);
not NOT1 (N11211, N11210);
nor NOR4 (N11212, N11207, N6064, N127, N7775);
or OR4 (N11213, N11206, N2979, N6784, N4849);
nand NAND3 (N11214, N11204, N4273, N9199);
not NOT1 (N11215, N11213);
nor NOR2 (N11216, N11212, N5122);
and AND4 (N11217, N11211, N5432, N71, N1957);
and AND3 (N11218, N11202, N10968, N11172);
and AND3 (N11219, N11209, N9025, N2316);
not NOT1 (N11220, N11219);
nor NOR4 (N11221, N11215, N6471, N2129, N8048);
nor NOR4 (N11222, N11214, N5164, N5470, N2800);
nor NOR3 (N11223, N11217, N8170, N8783);
not NOT1 (N11224, N11223);
nor NOR2 (N11225, N11191, N9907);
xor XOR2 (N11226, N11224, N10921);
nor NOR3 (N11227, N11222, N3267, N10793);
not NOT1 (N11228, N11225);
nand NAND4 (N11229, N11226, N8336, N5450, N7304);
and AND2 (N11230, N11216, N3434);
and AND2 (N11231, N11220, N4725);
buf BUF1 (N11232, N11227);
xor XOR2 (N11233, N11195, N2360);
nand NAND2 (N11234, N11218, N4184);
nand NAND4 (N11235, N11228, N11128, N7627, N2984);
nor NOR4 (N11236, N11231, N2029, N6028, N4131);
and AND2 (N11237, N11201, N5545);
nand NAND2 (N11238, N11189, N7321);
and AND2 (N11239, N11230, N9060);
nor NOR3 (N11240, N11237, N7799, N2307);
and AND4 (N11241, N11239, N10395, N9296, N4235);
nor NOR2 (N11242, N11240, N6455);
nor NOR2 (N11243, N11236, N8490);
buf BUF1 (N11244, N11238);
buf BUF1 (N11245, N11244);
buf BUF1 (N11246, N11229);
not NOT1 (N11247, N11245);
buf BUF1 (N11248, N11232);
xor XOR2 (N11249, N11233, N1253);
nand NAND4 (N11250, N11235, N7836, N346, N6562);
nor NOR4 (N11251, N11241, N5457, N795, N4928);
xor XOR2 (N11252, N11247, N1483);
xor XOR2 (N11253, N11249, N7977);
nand NAND2 (N11254, N11246, N2092);
nor NOR3 (N11255, N11250, N5716, N1684);
or OR2 (N11256, N11252, N8318);
or OR4 (N11257, N11242, N8744, N9102, N1678);
nand NAND4 (N11258, N11243, N3806, N41, N5923);
buf BUF1 (N11259, N11234);
or OR3 (N11260, N11253, N2837, N10290);
not NOT1 (N11261, N11251);
buf BUF1 (N11262, N11261);
or OR4 (N11263, N11221, N9596, N6613, N6806);
xor XOR2 (N11264, N11254, N11166);
or OR4 (N11265, N11264, N9593, N927, N10862);
nand NAND4 (N11266, N11258, N2800, N632, N3414);
buf BUF1 (N11267, N11263);
buf BUF1 (N11268, N11266);
not NOT1 (N11269, N11260);
nand NAND3 (N11270, N11268, N1981, N4798);
and AND3 (N11271, N11269, N10220, N7419);
buf BUF1 (N11272, N11248);
buf BUF1 (N11273, N11259);
nor NOR3 (N11274, N11257, N11253, N8330);
nand NAND4 (N11275, N11273, N10779, N4458, N3654);
and AND3 (N11276, N11270, N9364, N733);
buf BUF1 (N11277, N11265);
xor XOR2 (N11278, N11262, N6425);
buf BUF1 (N11279, N11275);
buf BUF1 (N11280, N11279);
nand NAND2 (N11281, N11256, N10187);
nor NOR3 (N11282, N11274, N6798, N1540);
xor XOR2 (N11283, N11278, N4185);
nor NOR2 (N11284, N11272, N10762);
and AND3 (N11285, N11281, N7998, N5985);
not NOT1 (N11286, N11267);
nor NOR4 (N11287, N11282, N7625, N10211, N10208);
or OR3 (N11288, N11287, N3367, N1962);
nand NAND2 (N11289, N11284, N28);
nand NAND4 (N11290, N11255, N8317, N1203, N10680);
nor NOR2 (N11291, N11280, N3241);
nor NOR2 (N11292, N11276, N10456);
buf BUF1 (N11293, N11291);
xor XOR2 (N11294, N11286, N2007);
not NOT1 (N11295, N11271);
xor XOR2 (N11296, N11290, N7634);
not NOT1 (N11297, N11293);
nand NAND2 (N11298, N11295, N6836);
or OR3 (N11299, N11277, N6275, N1733);
or OR4 (N11300, N11299, N5652, N2081, N9325);
nor NOR2 (N11301, N11289, N1485);
or OR4 (N11302, N11285, N3533, N3318, N3923);
not NOT1 (N11303, N11294);
or OR4 (N11304, N11283, N7209, N713, N2669);
nand NAND2 (N11305, N11303, N1515);
xor XOR2 (N11306, N11300, N2466);
buf BUF1 (N11307, N11292);
and AND2 (N11308, N11306, N1721);
nor NOR3 (N11309, N11297, N8741, N831);
not NOT1 (N11310, N11302);
and AND2 (N11311, N11305, N643);
or OR4 (N11312, N11301, N10966, N7342, N3339);
and AND4 (N11313, N11308, N763, N4553, N11279);
nor NOR3 (N11314, N11309, N275, N4850);
or OR4 (N11315, N11307, N2212, N8024, N1210);
nand NAND2 (N11316, N11288, N9010);
nor NOR4 (N11317, N11316, N9287, N10748, N4744);
and AND3 (N11318, N11313, N44, N6224);
and AND4 (N11319, N11317, N10721, N7654, N1618);
nor NOR4 (N11320, N11298, N4392, N6673, N10824);
not NOT1 (N11321, N11318);
buf BUF1 (N11322, N11304);
or OR3 (N11323, N11321, N5170, N8993);
nor NOR3 (N11324, N11320, N3169, N7527);
or OR4 (N11325, N11319, N4846, N5753, N1108);
buf BUF1 (N11326, N11325);
not NOT1 (N11327, N11322);
not NOT1 (N11328, N11315);
or OR3 (N11329, N11327, N9564, N11234);
not NOT1 (N11330, N11324);
xor XOR2 (N11331, N11323, N698);
nor NOR3 (N11332, N11328, N3967, N8179);
buf BUF1 (N11333, N11331);
or OR4 (N11334, N11326, N10005, N10711, N888);
not NOT1 (N11335, N11311);
nand NAND3 (N11336, N11333, N6781, N6149);
and AND2 (N11337, N11312, N4099);
or OR2 (N11338, N11332, N7534);
buf BUF1 (N11339, N11334);
xor XOR2 (N11340, N11310, N8607);
buf BUF1 (N11341, N11296);
not NOT1 (N11342, N11338);
nor NOR4 (N11343, N11330, N10043, N7259, N955);
not NOT1 (N11344, N11343);
xor XOR2 (N11345, N11342, N5083);
buf BUF1 (N11346, N11335);
or OR2 (N11347, N11344, N10925);
xor XOR2 (N11348, N11346, N6222);
and AND4 (N11349, N11347, N9994, N8259, N10380);
nor NOR3 (N11350, N11339, N3904, N7524);
or OR3 (N11351, N11341, N9586, N9049);
nand NAND3 (N11352, N11336, N5707, N5353);
xor XOR2 (N11353, N11352, N4632);
nor NOR3 (N11354, N11353, N4341, N2541);
or OR3 (N11355, N11349, N8790, N11058);
nor NOR4 (N11356, N11354, N3780, N8778, N5587);
buf BUF1 (N11357, N11345);
xor XOR2 (N11358, N11351, N10306);
nand NAND2 (N11359, N11329, N4608);
and AND2 (N11360, N11340, N3206);
not NOT1 (N11361, N11356);
xor XOR2 (N11362, N11355, N2409);
or OR2 (N11363, N11362, N1918);
or OR3 (N11364, N11360, N2692, N787);
buf BUF1 (N11365, N11363);
and AND4 (N11366, N11364, N1521, N7445, N162);
xor XOR2 (N11367, N11350, N8832);
nand NAND2 (N11368, N11348, N3858);
not NOT1 (N11369, N11358);
and AND3 (N11370, N11365, N47, N7513);
or OR4 (N11371, N11337, N769, N1214, N4511);
buf BUF1 (N11372, N11371);
or OR2 (N11373, N11372, N4235);
xor XOR2 (N11374, N11359, N2557);
not NOT1 (N11375, N11357);
nand NAND2 (N11376, N11367, N5265);
buf BUF1 (N11377, N11366);
xor XOR2 (N11378, N11368, N5162);
not NOT1 (N11379, N11314);
not NOT1 (N11380, N11378);
xor XOR2 (N11381, N11361, N4467);
nand NAND3 (N11382, N11379, N391, N2312);
buf BUF1 (N11383, N11369);
buf BUF1 (N11384, N11375);
nand NAND2 (N11385, N11383, N5666);
nor NOR3 (N11386, N11373, N9835, N6130);
and AND4 (N11387, N11370, N2624, N3724, N7175);
or OR2 (N11388, N11387, N6027);
buf BUF1 (N11389, N11384);
nor NOR3 (N11390, N11381, N3184, N2488);
buf BUF1 (N11391, N11385);
xor XOR2 (N11392, N11382, N9282);
nand NAND3 (N11393, N11390, N9514, N969);
nor NOR4 (N11394, N11391, N4210, N1264, N8589);
nand NAND3 (N11395, N11393, N10852, N31);
xor XOR2 (N11396, N11392, N3053);
nand NAND4 (N11397, N11389, N11000, N4269, N6959);
and AND3 (N11398, N11376, N7184, N27);
xor XOR2 (N11399, N11398, N1979);
xor XOR2 (N11400, N11396, N3821);
buf BUF1 (N11401, N11377);
buf BUF1 (N11402, N11395);
nor NOR3 (N11403, N11397, N8124, N5137);
or OR2 (N11404, N11374, N5337);
nand NAND2 (N11405, N11394, N7071);
not NOT1 (N11406, N11386);
xor XOR2 (N11407, N11400, N1312);
nand NAND3 (N11408, N11399, N4463, N10041);
or OR4 (N11409, N11402, N7982, N9880, N9057);
and AND2 (N11410, N11409, N10388);
not NOT1 (N11411, N11404);
nand NAND3 (N11412, N11410, N4079, N8929);
nor NOR3 (N11413, N11412, N9389, N4067);
or OR3 (N11414, N11406, N10109, N6598);
nand NAND3 (N11415, N11405, N2867, N10382);
nand NAND3 (N11416, N11403, N4259, N5127);
nand NAND2 (N11417, N11411, N5737);
xor XOR2 (N11418, N11407, N6362);
nor NOR2 (N11419, N11417, N10788);
and AND2 (N11420, N11401, N9626);
and AND2 (N11421, N11388, N2068);
and AND3 (N11422, N11408, N4814, N5802);
and AND3 (N11423, N11415, N4803, N6872);
buf BUF1 (N11424, N11421);
nand NAND3 (N11425, N11423, N9082, N10031);
and AND4 (N11426, N11416, N9277, N3203, N1043);
not NOT1 (N11427, N11413);
nand NAND4 (N11428, N11420, N3075, N6913, N6520);
buf BUF1 (N11429, N11427);
and AND2 (N11430, N11422, N220);
or OR3 (N11431, N11426, N3119, N9227);
not NOT1 (N11432, N11424);
nand NAND2 (N11433, N11414, N5275);
nor NOR3 (N11434, N11419, N10764, N8796);
not NOT1 (N11435, N11433);
and AND4 (N11436, N11425, N9807, N11276, N5833);
and AND3 (N11437, N11430, N4769, N9717);
xor XOR2 (N11438, N11380, N6378);
nand NAND4 (N11439, N11432, N10656, N11436, N2771);
buf BUF1 (N11440, N7811);
nand NAND2 (N11441, N11439, N8458);
buf BUF1 (N11442, N11435);
and AND3 (N11443, N11441, N2433, N437);
not NOT1 (N11444, N11442);
xor XOR2 (N11445, N11418, N912);
and AND4 (N11446, N11443, N216, N985, N3010);
nor NOR3 (N11447, N11445, N3938, N1271);
or OR3 (N11448, N11431, N10436, N4622);
or OR4 (N11449, N11437, N6701, N4642, N9521);
not NOT1 (N11450, N11449);
or OR3 (N11451, N11448, N6548, N2413);
or OR3 (N11452, N11438, N638, N5170);
nand NAND4 (N11453, N11444, N6921, N11132, N3942);
not NOT1 (N11454, N11428);
and AND3 (N11455, N11440, N8575, N9169);
buf BUF1 (N11456, N11450);
buf BUF1 (N11457, N11452);
buf BUF1 (N11458, N11429);
and AND4 (N11459, N11457, N162, N6687, N3046);
or OR3 (N11460, N11456, N1813, N4942);
not NOT1 (N11461, N11453);
nand NAND4 (N11462, N11454, N7310, N8940, N8028);
buf BUF1 (N11463, N11458);
xor XOR2 (N11464, N11462, N9371);
nor NOR2 (N11465, N11463, N2537);
or OR3 (N11466, N11459, N4777, N10672);
xor XOR2 (N11467, N11464, N655);
buf BUF1 (N11468, N11434);
xor XOR2 (N11469, N11455, N8427);
nor NOR4 (N11470, N11447, N8728, N119, N6677);
nor NOR3 (N11471, N11470, N3372, N3035);
and AND4 (N11472, N11465, N6172, N2115, N3398);
nand NAND4 (N11473, N11446, N4009, N11198, N8604);
xor XOR2 (N11474, N11467, N5920);
and AND3 (N11475, N11468, N7550, N5312);
buf BUF1 (N11476, N11461);
xor XOR2 (N11477, N11471, N10634);
nor NOR4 (N11478, N11469, N5169, N9039, N1574);
buf BUF1 (N11479, N11473);
and AND4 (N11480, N11478, N144, N4909, N516);
nor NOR2 (N11481, N11451, N7770);
not NOT1 (N11482, N11481);
nand NAND2 (N11483, N11475, N6498);
nor NOR2 (N11484, N11480, N7702);
buf BUF1 (N11485, N11482);
nand NAND4 (N11486, N11476, N8097, N400, N1307);
nand NAND2 (N11487, N11466, N8342);
nor NOR2 (N11488, N11487, N2774);
not NOT1 (N11489, N11479);
and AND2 (N11490, N11474, N10432);
not NOT1 (N11491, N11488);
or OR2 (N11492, N11483, N10333);
buf BUF1 (N11493, N11460);
nand NAND2 (N11494, N11486, N7106);
nor NOR4 (N11495, N11485, N7033, N5935, N9101);
xor XOR2 (N11496, N11494, N5318);
or OR4 (N11497, N11491, N7135, N9206, N6990);
nand NAND4 (N11498, N11492, N4139, N8267, N6590);
and AND3 (N11499, N11484, N1197, N5873);
or OR4 (N11500, N11496, N6146, N10407, N10294);
or OR4 (N11501, N11489, N2687, N8976, N10157);
nand NAND4 (N11502, N11495, N3980, N5212, N8214);
buf BUF1 (N11503, N11502);
buf BUF1 (N11504, N11501);
and AND3 (N11505, N11497, N7492, N8713);
nand NAND3 (N11506, N11477, N1061, N3792);
xor XOR2 (N11507, N11505, N10963);
nor NOR4 (N11508, N11472, N5022, N11433, N9546);
buf BUF1 (N11509, N11504);
buf BUF1 (N11510, N11509);
xor XOR2 (N11511, N11503, N3023);
xor XOR2 (N11512, N11498, N8598);
and AND3 (N11513, N11512, N6030, N10787);
and AND3 (N11514, N11500, N2384, N458);
buf BUF1 (N11515, N11510);
not NOT1 (N11516, N11507);
buf BUF1 (N11517, N11515);
buf BUF1 (N11518, N11517);
nand NAND3 (N11519, N11508, N7440, N5940);
and AND3 (N11520, N11513, N6745, N10290);
xor XOR2 (N11521, N11493, N1744);
not NOT1 (N11522, N11519);
nand NAND2 (N11523, N11514, N2349);
buf BUF1 (N11524, N11518);
or OR2 (N11525, N11506, N9345);
and AND2 (N11526, N11524, N11471);
buf BUF1 (N11527, N11516);
nand NAND2 (N11528, N11526, N2170);
buf BUF1 (N11529, N11490);
buf BUF1 (N11530, N11511);
xor XOR2 (N11531, N11525, N10919);
and AND2 (N11532, N11520, N6509);
xor XOR2 (N11533, N11523, N9136);
nand NAND4 (N11534, N11531, N4309, N9684, N7752);
and AND4 (N11535, N11533, N54, N9025, N2197);
and AND3 (N11536, N11532, N7183, N11470);
or OR2 (N11537, N11530, N6824);
not NOT1 (N11538, N11537);
nand NAND3 (N11539, N11521, N4181, N10738);
xor XOR2 (N11540, N11528, N6793);
nor NOR4 (N11541, N11535, N6504, N4987, N2838);
xor XOR2 (N11542, N11538, N7406);
nor NOR2 (N11543, N11529, N3316);
buf BUF1 (N11544, N11543);
not NOT1 (N11545, N11536);
not NOT1 (N11546, N11539);
and AND2 (N11547, N11499, N9284);
buf BUF1 (N11548, N11547);
and AND4 (N11549, N11542, N7061, N8337, N2907);
xor XOR2 (N11550, N11549, N3525);
nand NAND3 (N11551, N11541, N4121, N1941);
xor XOR2 (N11552, N11527, N2701);
or OR4 (N11553, N11551, N3743, N11256, N3737);
xor XOR2 (N11554, N11546, N4769);
and AND2 (N11555, N11534, N6397);
or OR4 (N11556, N11545, N2377, N2573, N10605);
nor NOR4 (N11557, N11522, N10572, N3348, N6153);
xor XOR2 (N11558, N11556, N8153);
nor NOR2 (N11559, N11548, N11520);
and AND2 (N11560, N11553, N3109);
buf BUF1 (N11561, N11540);
buf BUF1 (N11562, N11552);
not NOT1 (N11563, N11550);
xor XOR2 (N11564, N11554, N3714);
buf BUF1 (N11565, N11559);
and AND3 (N11566, N11564, N5535, N8685);
nor NOR2 (N11567, N11558, N11060);
not NOT1 (N11568, N11555);
buf BUF1 (N11569, N11565);
not NOT1 (N11570, N11560);
and AND2 (N11571, N11563, N5892);
buf BUF1 (N11572, N11544);
and AND4 (N11573, N11572, N9652, N10512, N9699);
not NOT1 (N11574, N11566);
not NOT1 (N11575, N11561);
nand NAND4 (N11576, N11575, N1414, N10656, N9860);
and AND4 (N11577, N11568, N5612, N6992, N2535);
or OR4 (N11578, N11576, N6879, N4584, N6187);
not NOT1 (N11579, N11578);
or OR2 (N11580, N11579, N2847);
not NOT1 (N11581, N11577);
xor XOR2 (N11582, N11562, N1831);
not NOT1 (N11583, N11569);
and AND2 (N11584, N11557, N5676);
buf BUF1 (N11585, N11574);
and AND2 (N11586, N11573, N3233);
nand NAND2 (N11587, N11583, N4570);
nor NOR3 (N11588, N11584, N11117, N1992);
xor XOR2 (N11589, N11567, N10878);
nor NOR4 (N11590, N11587, N125, N3621, N10343);
and AND2 (N11591, N11589, N533);
xor XOR2 (N11592, N11590, N10254);
not NOT1 (N11593, N11570);
nand NAND3 (N11594, N11588, N244, N7924);
and AND3 (N11595, N11571, N4125, N4706);
and AND3 (N11596, N11593, N1490, N9857);
buf BUF1 (N11597, N11591);
and AND2 (N11598, N11581, N741);
xor XOR2 (N11599, N11595, N8480);
buf BUF1 (N11600, N11592);
nand NAND2 (N11601, N11582, N6002);
or OR2 (N11602, N11599, N2851);
nor NOR4 (N11603, N11602, N3819, N2890, N4485);
buf BUF1 (N11604, N11600);
nor NOR3 (N11605, N11585, N10573, N1233);
buf BUF1 (N11606, N11597);
and AND4 (N11607, N11598, N849, N5626, N7427);
nor NOR2 (N11608, N11606, N2354);
nand NAND3 (N11609, N11586, N10634, N9477);
and AND3 (N11610, N11604, N6599, N7178);
nand NAND3 (N11611, N11580, N9104, N11542);
not NOT1 (N11612, N11603);
or OR3 (N11613, N11596, N2928, N10032);
and AND2 (N11614, N11608, N1257);
xor XOR2 (N11615, N11613, N4488);
or OR2 (N11616, N11605, N181);
buf BUF1 (N11617, N11614);
xor XOR2 (N11618, N11594, N5426);
nor NOR3 (N11619, N11601, N7634, N3270);
xor XOR2 (N11620, N11618, N6311);
or OR4 (N11621, N11615, N10616, N10136, N5264);
and AND2 (N11622, N11610, N6353);
xor XOR2 (N11623, N11612, N4471);
nand NAND3 (N11624, N11611, N7025, N2755);
xor XOR2 (N11625, N11621, N11043);
or OR3 (N11626, N11609, N9810, N3965);
not NOT1 (N11627, N11620);
xor XOR2 (N11628, N11622, N6732);
nor NOR3 (N11629, N11617, N141, N7625);
buf BUF1 (N11630, N11629);
and AND3 (N11631, N11624, N6813, N3965);
xor XOR2 (N11632, N11628, N1492);
nand NAND3 (N11633, N11623, N73, N10999);
nor NOR4 (N11634, N11632, N2636, N10103, N7610);
and AND4 (N11635, N11627, N3895, N5325, N6653);
nand NAND4 (N11636, N11607, N1921, N3242, N5454);
buf BUF1 (N11637, N11634);
nand NAND4 (N11638, N11636, N4788, N1273, N9878);
or OR4 (N11639, N11630, N6043, N7571, N10051);
xor XOR2 (N11640, N11633, N5116);
or OR4 (N11641, N11631, N9511, N704, N3260);
nor NOR4 (N11642, N11626, N1819, N4999, N7553);
not NOT1 (N11643, N11638);
buf BUF1 (N11644, N11616);
nor NOR2 (N11645, N11637, N5827);
not NOT1 (N11646, N11639);
xor XOR2 (N11647, N11642, N9060);
xor XOR2 (N11648, N11625, N2825);
nor NOR3 (N11649, N11640, N1334, N7266);
nor NOR3 (N11650, N11646, N5285, N9523);
or OR3 (N11651, N11644, N9517, N5178);
nor NOR2 (N11652, N11647, N9236);
buf BUF1 (N11653, N11643);
nand NAND3 (N11654, N11651, N8666, N10873);
or OR4 (N11655, N11648, N2858, N2041, N2933);
buf BUF1 (N11656, N11619);
xor XOR2 (N11657, N11645, N4065);
and AND3 (N11658, N11635, N1820, N6842);
nor NOR4 (N11659, N11653, N1303, N11082, N6615);
not NOT1 (N11660, N11655);
xor XOR2 (N11661, N11656, N470);
not NOT1 (N11662, N11659);
xor XOR2 (N11663, N11662, N9846);
buf BUF1 (N11664, N11657);
nor NOR2 (N11665, N11641, N3507);
not NOT1 (N11666, N11652);
not NOT1 (N11667, N11664);
nor NOR3 (N11668, N11654, N6993, N5166);
xor XOR2 (N11669, N11660, N4469);
nor NOR2 (N11670, N11663, N1268);
buf BUF1 (N11671, N11658);
xor XOR2 (N11672, N11671, N10211);
not NOT1 (N11673, N11667);
and AND2 (N11674, N11665, N854);
nor NOR4 (N11675, N11674, N5147, N9894, N7583);
not NOT1 (N11676, N11649);
buf BUF1 (N11677, N11673);
and AND4 (N11678, N11661, N10238, N10394, N5842);
buf BUF1 (N11679, N11678);
nor NOR3 (N11680, N11672, N8802, N10004);
buf BUF1 (N11681, N11668);
buf BUF1 (N11682, N11666);
and AND3 (N11683, N11676, N7879, N11498);
buf BUF1 (N11684, N11669);
or OR3 (N11685, N11675, N10645, N9150);
or OR3 (N11686, N11682, N4539, N6536);
and AND3 (N11687, N11677, N4765, N9414);
and AND3 (N11688, N11687, N10444, N3748);
and AND2 (N11689, N11688, N6107);
and AND4 (N11690, N11680, N5385, N2405, N9203);
nor NOR2 (N11691, N11650, N10039);
nor NOR2 (N11692, N11679, N1403);
not NOT1 (N11693, N11684);
or OR4 (N11694, N11686, N38, N8723, N2649);
nand NAND4 (N11695, N11683, N9492, N3933, N10760);
not NOT1 (N11696, N11670);
and AND3 (N11697, N11694, N3265, N3439);
xor XOR2 (N11698, N11685, N5072);
buf BUF1 (N11699, N11692);
nand NAND2 (N11700, N11693, N219);
xor XOR2 (N11701, N11681, N7434);
or OR2 (N11702, N11697, N9469);
nand NAND4 (N11703, N11699, N4016, N2049, N7254);
xor XOR2 (N11704, N11690, N4373);
and AND4 (N11705, N11696, N7041, N2713, N370);
xor XOR2 (N11706, N11703, N9952);
nor NOR2 (N11707, N11702, N2124);
and AND4 (N11708, N11700, N875, N11546, N4220);
nor NOR3 (N11709, N11707, N6227, N5447);
and AND4 (N11710, N11701, N9870, N8691, N9464);
and AND3 (N11711, N11710, N8096, N9135);
buf BUF1 (N11712, N11704);
nor NOR2 (N11713, N11709, N10426);
nor NOR3 (N11714, N11689, N8998, N10024);
buf BUF1 (N11715, N11711);
or OR3 (N11716, N11706, N6121, N6156);
nand NAND4 (N11717, N11698, N11465, N1519, N465);
xor XOR2 (N11718, N11708, N675);
or OR2 (N11719, N11695, N10712);
nand NAND3 (N11720, N11712, N9591, N8561);
nand NAND3 (N11721, N11720, N7819, N8168);
nand NAND2 (N11722, N11715, N4562);
nand NAND2 (N11723, N11716, N4118);
not NOT1 (N11724, N11714);
not NOT1 (N11725, N11691);
buf BUF1 (N11726, N11722);
buf BUF1 (N11727, N11726);
nor NOR2 (N11728, N11718, N4267);
nand NAND3 (N11729, N11728, N5880, N9541);
xor XOR2 (N11730, N11705, N1616);
not NOT1 (N11731, N11719);
not NOT1 (N11732, N11717);
not NOT1 (N11733, N11730);
buf BUF1 (N11734, N11731);
not NOT1 (N11735, N11724);
nand NAND3 (N11736, N11723, N1523, N7031);
nor NOR4 (N11737, N11735, N1554, N2513, N6176);
not NOT1 (N11738, N11727);
nand NAND2 (N11739, N11729, N2738);
xor XOR2 (N11740, N11713, N5241);
buf BUF1 (N11741, N11738);
and AND3 (N11742, N11741, N5933, N8588);
not NOT1 (N11743, N11733);
nor NOR2 (N11744, N11725, N10711);
nand NAND3 (N11745, N11740, N7482, N745);
nor NOR4 (N11746, N11736, N9161, N6127, N10644);
nor NOR2 (N11747, N11743, N7179);
nor NOR4 (N11748, N11742, N7718, N2408, N8000);
xor XOR2 (N11749, N11745, N6665);
and AND2 (N11750, N11744, N6989);
and AND3 (N11751, N11721, N968, N4317);
or OR3 (N11752, N11746, N340, N9662);
or OR4 (N11753, N11750, N3871, N4646, N6222);
xor XOR2 (N11754, N11734, N6690);
buf BUF1 (N11755, N11752);
not NOT1 (N11756, N11747);
or OR3 (N11757, N11749, N7946, N1950);
xor XOR2 (N11758, N11756, N893);
buf BUF1 (N11759, N11739);
nor NOR3 (N11760, N11754, N2938, N2007);
or OR4 (N11761, N11759, N4798, N4952, N6154);
nor NOR2 (N11762, N11751, N8213);
buf BUF1 (N11763, N11761);
or OR3 (N11764, N11763, N1479, N524);
nand NAND4 (N11765, N11764, N1854, N4821, N11250);
or OR4 (N11766, N11753, N6329, N3615, N10284);
nand NAND2 (N11767, N11766, N8074);
nor NOR4 (N11768, N11765, N6739, N11230, N8547);
and AND2 (N11769, N11760, N8348);
and AND4 (N11770, N11748, N10479, N9064, N8220);
and AND4 (N11771, N11732, N1992, N5222, N11310);
not NOT1 (N11772, N11768);
or OR3 (N11773, N11757, N2643, N5756);
nor NOR2 (N11774, N11755, N2689);
not NOT1 (N11775, N11767);
buf BUF1 (N11776, N11773);
nand NAND2 (N11777, N11758, N5435);
not NOT1 (N11778, N11774);
and AND2 (N11779, N11762, N7303);
nand NAND3 (N11780, N11775, N3353, N1383);
buf BUF1 (N11781, N11737);
xor XOR2 (N11782, N11770, N8227);
buf BUF1 (N11783, N11779);
nand NAND3 (N11784, N11780, N2192, N8919);
nor NOR3 (N11785, N11772, N7511, N8693);
not NOT1 (N11786, N11784);
and AND4 (N11787, N11785, N9902, N2053, N531);
nor NOR3 (N11788, N11781, N4664, N262);
or OR2 (N11789, N11787, N7252);
xor XOR2 (N11790, N11771, N10476);
nand NAND4 (N11791, N11776, N915, N7216, N314);
nand NAND2 (N11792, N11790, N1588);
and AND4 (N11793, N11789, N3961, N692, N7919);
xor XOR2 (N11794, N11786, N1111);
nor NOR2 (N11795, N11777, N6603);
or OR3 (N11796, N11778, N1756, N1758);
nor NOR4 (N11797, N11792, N3964, N3038, N6667);
buf BUF1 (N11798, N11791);
nand NAND2 (N11799, N11797, N5815);
nor NOR4 (N11800, N11782, N9260, N4606, N8161);
nand NAND2 (N11801, N11799, N6626);
or OR4 (N11802, N11783, N5699, N3684, N6961);
xor XOR2 (N11803, N11793, N4963);
and AND3 (N11804, N11795, N6963, N458);
or OR2 (N11805, N11800, N10148);
or OR4 (N11806, N11803, N353, N6250, N7591);
nand NAND3 (N11807, N11802, N9659, N949);
nand NAND2 (N11808, N11801, N8291);
nor NOR4 (N11809, N11806, N2303, N1748, N7061);
nand NAND2 (N11810, N11798, N4066);
or OR2 (N11811, N11804, N8640);
nand NAND2 (N11812, N11805, N10295);
xor XOR2 (N11813, N11796, N5522);
xor XOR2 (N11814, N11769, N7491);
nand NAND4 (N11815, N11788, N6243, N1916, N8847);
nand NAND4 (N11816, N11809, N6470, N20, N321);
nor NOR3 (N11817, N11815, N6591, N7658);
nor NOR2 (N11818, N11808, N11185);
not NOT1 (N11819, N11813);
not NOT1 (N11820, N11810);
nand NAND2 (N11821, N11817, N9108);
and AND2 (N11822, N11820, N7696);
nor NOR2 (N11823, N11812, N3549);
nand NAND2 (N11824, N11821, N3281);
buf BUF1 (N11825, N11824);
xor XOR2 (N11826, N11816, N7293);
nor NOR2 (N11827, N11814, N5949);
not NOT1 (N11828, N11826);
nand NAND2 (N11829, N11794, N3795);
not NOT1 (N11830, N11807);
or OR3 (N11831, N11818, N2724, N7345);
nand NAND2 (N11832, N11822, N5860);
buf BUF1 (N11833, N11823);
and AND4 (N11834, N11828, N4442, N4548, N9961);
not NOT1 (N11835, N11811);
nand NAND3 (N11836, N11825, N9353, N4994);
nor NOR4 (N11837, N11829, N1038, N8698, N5434);
or OR4 (N11838, N11830, N7413, N1292, N4724);
or OR4 (N11839, N11831, N7264, N3528, N2650);
buf BUF1 (N11840, N11839);
xor XOR2 (N11841, N11838, N2384);
and AND3 (N11842, N11840, N563, N5048);
not NOT1 (N11843, N11837);
nand NAND2 (N11844, N11841, N9607);
nor NOR4 (N11845, N11842, N6523, N9927, N8310);
nand NAND4 (N11846, N11835, N5760, N10892, N4794);
xor XOR2 (N11847, N11843, N9969);
nor NOR2 (N11848, N11844, N4231);
buf BUF1 (N11849, N11836);
nand NAND4 (N11850, N11834, N7461, N1087, N9357);
and AND3 (N11851, N11827, N4746, N4302);
and AND4 (N11852, N11832, N280, N10945, N709);
not NOT1 (N11853, N11846);
nor NOR3 (N11854, N11819, N9515, N7356);
or OR2 (N11855, N11847, N11244);
and AND2 (N11856, N11854, N8197);
nand NAND2 (N11857, N11853, N331);
and AND2 (N11858, N11848, N2516);
nor NOR3 (N11859, N11857, N7297, N11242);
not NOT1 (N11860, N11850);
not NOT1 (N11861, N11860);
not NOT1 (N11862, N11833);
not NOT1 (N11863, N11845);
or OR2 (N11864, N11859, N5705);
nor NOR4 (N11865, N11851, N6283, N11509, N8907);
buf BUF1 (N11866, N11863);
not NOT1 (N11867, N11852);
or OR3 (N11868, N11855, N8867, N120);
xor XOR2 (N11869, N11867, N2228);
xor XOR2 (N11870, N11864, N6810);
nand NAND4 (N11871, N11849, N7172, N1259, N10677);
not NOT1 (N11872, N11856);
nor NOR3 (N11873, N11861, N9171, N9976);
xor XOR2 (N11874, N11862, N11480);
buf BUF1 (N11875, N11866);
xor XOR2 (N11876, N11875, N9141);
buf BUF1 (N11877, N11865);
buf BUF1 (N11878, N11877);
buf BUF1 (N11879, N11873);
not NOT1 (N11880, N11874);
nor NOR4 (N11881, N11872, N1616, N6457, N6146);
not NOT1 (N11882, N11881);
or OR2 (N11883, N11879, N960);
nand NAND2 (N11884, N11883, N10239);
and AND3 (N11885, N11880, N7596, N11874);
not NOT1 (N11886, N11878);
xor XOR2 (N11887, N11871, N11381);
and AND2 (N11888, N11884, N9422);
xor XOR2 (N11889, N11858, N4327);
nor NOR4 (N11890, N11868, N7116, N11622, N7413);
buf BUF1 (N11891, N11890);
nand NAND3 (N11892, N11870, N8966, N5929);
or OR2 (N11893, N11876, N8993);
nand NAND3 (N11894, N11882, N1062, N9244);
and AND2 (N11895, N11869, N6965);
buf BUF1 (N11896, N11894);
not NOT1 (N11897, N11885);
nand NAND2 (N11898, N11887, N3746);
nand NAND4 (N11899, N11892, N7246, N7462, N3460);
nor NOR2 (N11900, N11898, N2370);
nor NOR3 (N11901, N11895, N228, N1716);
xor XOR2 (N11902, N11897, N9084);
xor XOR2 (N11903, N11888, N7929);
nor NOR3 (N11904, N11902, N473, N37);
nor NOR3 (N11905, N11893, N7326, N473);
nand NAND2 (N11906, N11900, N10946);
xor XOR2 (N11907, N11905, N6197);
buf BUF1 (N11908, N11886);
xor XOR2 (N11909, N11908, N1547);
nor NOR2 (N11910, N11889, N8741);
buf BUF1 (N11911, N11906);
xor XOR2 (N11912, N11891, N1444);
and AND3 (N11913, N11903, N5492, N11008);
or OR4 (N11914, N11899, N3292, N2387, N11892);
not NOT1 (N11915, N11910);
xor XOR2 (N11916, N11909, N3828);
or OR2 (N11917, N11916, N8366);
and AND4 (N11918, N11907, N3518, N1058, N6547);
buf BUF1 (N11919, N11911);
not NOT1 (N11920, N11915);
or OR4 (N11921, N11920, N7793, N8436, N7177);
not NOT1 (N11922, N11896);
and AND2 (N11923, N11901, N3559);
or OR3 (N11924, N11917, N8748, N49);
buf BUF1 (N11925, N11921);
nand NAND4 (N11926, N11904, N8914, N292, N8353);
buf BUF1 (N11927, N11926);
nor NOR4 (N11928, N11912, N6071, N370, N5661);
xor XOR2 (N11929, N11918, N11697);
and AND3 (N11930, N11925, N4999, N376);
nor NOR4 (N11931, N11927, N6866, N8809, N4739);
not NOT1 (N11932, N11919);
xor XOR2 (N11933, N11928, N2703);
buf BUF1 (N11934, N11930);
and AND2 (N11935, N11932, N1680);
and AND2 (N11936, N11934, N4013);
nand NAND4 (N11937, N11933, N5093, N5055, N11877);
buf BUF1 (N11938, N11913);
or OR3 (N11939, N11923, N6492, N665);
nor NOR4 (N11940, N11937, N11411, N3151, N11076);
and AND3 (N11941, N11940, N11202, N2834);
and AND2 (N11942, N11929, N583);
buf BUF1 (N11943, N11914);
buf BUF1 (N11944, N11939);
nand NAND2 (N11945, N11941, N7948);
xor XOR2 (N11946, N11944, N3200);
nor NOR4 (N11947, N11935, N3210, N5554, N3612);
buf BUF1 (N11948, N11938);
and AND4 (N11949, N11948, N11781, N11478, N11149);
xor XOR2 (N11950, N11924, N3614);
not NOT1 (N11951, N11947);
nor NOR3 (N11952, N11950, N3248, N8271);
buf BUF1 (N11953, N11945);
or OR2 (N11954, N11942, N9581);
buf BUF1 (N11955, N11952);
or OR4 (N11956, N11949, N2295, N9790, N9628);
xor XOR2 (N11957, N11943, N9504);
and AND4 (N11958, N11931, N3843, N8319, N3763);
nand NAND2 (N11959, N11955, N11465);
xor XOR2 (N11960, N11951, N11105);
xor XOR2 (N11961, N11953, N3871);
or OR3 (N11962, N11959, N11050, N6380);
or OR3 (N11963, N11957, N7427, N8573);
nor NOR2 (N11964, N11956, N11857);
and AND3 (N11965, N11960, N3254, N1995);
nand NAND2 (N11966, N11946, N9977);
and AND4 (N11967, N11954, N1620, N6217, N3226);
not NOT1 (N11968, N11961);
xor XOR2 (N11969, N11964, N11000);
nand NAND3 (N11970, N11936, N2430, N9820);
xor XOR2 (N11971, N11970, N7652);
nand NAND3 (N11972, N11962, N10728, N9386);
nand NAND3 (N11973, N11958, N10814, N4851);
nand NAND3 (N11974, N11966, N1991, N540);
and AND2 (N11975, N11922, N5341);
not NOT1 (N11976, N11971);
nand NAND2 (N11977, N11963, N19);
buf BUF1 (N11978, N11965);
or OR3 (N11979, N11975, N8453, N4457);
nor NOR2 (N11980, N11973, N10569);
not NOT1 (N11981, N11972);
and AND2 (N11982, N11976, N2672);
not NOT1 (N11983, N11967);
and AND3 (N11984, N11978, N7363, N2776);
not NOT1 (N11985, N11979);
xor XOR2 (N11986, N11984, N1929);
nand NAND3 (N11987, N11983, N1952, N10462);
buf BUF1 (N11988, N11974);
or OR3 (N11989, N11969, N504, N11371);
or OR3 (N11990, N11985, N2798, N11190);
nor NOR2 (N11991, N11988, N6904);
not NOT1 (N11992, N11981);
xor XOR2 (N11993, N11977, N305);
not NOT1 (N11994, N11987);
or OR3 (N11995, N11990, N6959, N10069);
nand NAND3 (N11996, N11994, N11418, N11027);
nand NAND3 (N11997, N11991, N11469, N4518);
not NOT1 (N11998, N11992);
nor NOR4 (N11999, N11980, N2880, N19, N5785);
not NOT1 (N12000, N11989);
nor NOR3 (N12001, N11995, N10944, N6116);
nor NOR3 (N12002, N11982, N11806, N10694);
not NOT1 (N12003, N11986);
nand NAND4 (N12004, N11996, N3623, N5427, N3959);
and AND4 (N12005, N11993, N11292, N11118, N3917);
xor XOR2 (N12006, N12005, N7612);
and AND4 (N12007, N11998, N8654, N3904, N10739);
not NOT1 (N12008, N12002);
buf BUF1 (N12009, N12000);
not NOT1 (N12010, N12003);
or OR3 (N12011, N11968, N7131, N3918);
xor XOR2 (N12012, N11997, N11371);
xor XOR2 (N12013, N11999, N1945);
not NOT1 (N12014, N12004);
and AND3 (N12015, N12013, N10781, N11457);
and AND2 (N12016, N12001, N3995);
not NOT1 (N12017, N12012);
xor XOR2 (N12018, N12011, N10444);
nand NAND4 (N12019, N12006, N8945, N5692, N3193);
or OR3 (N12020, N12010, N5846, N11732);
buf BUF1 (N12021, N12016);
or OR2 (N12022, N12007, N958);
not NOT1 (N12023, N12022);
or OR4 (N12024, N12021, N10538, N5922, N2698);
buf BUF1 (N12025, N12020);
buf BUF1 (N12026, N12017);
not NOT1 (N12027, N12026);
buf BUF1 (N12028, N12024);
or OR4 (N12029, N12028, N2665, N4426, N3473);
and AND4 (N12030, N12027, N7650, N294, N5151);
nor NOR2 (N12031, N12023, N2913);
buf BUF1 (N12032, N12009);
not NOT1 (N12033, N12025);
and AND3 (N12034, N12008, N4338, N4420);
or OR4 (N12035, N12029, N8569, N5948, N811);
not NOT1 (N12036, N12031);
xor XOR2 (N12037, N12014, N206);
and AND4 (N12038, N12019, N629, N10738, N3380);
not NOT1 (N12039, N12030);
not NOT1 (N12040, N12036);
not NOT1 (N12041, N12018);
or OR4 (N12042, N12038, N4552, N3432, N844);
buf BUF1 (N12043, N12042);
and AND4 (N12044, N12032, N6710, N10349, N49);
or OR4 (N12045, N12015, N1506, N8836, N11088);
or OR4 (N12046, N12039, N5659, N11827, N6984);
and AND2 (N12047, N12034, N7085);
nand NAND3 (N12048, N12035, N1394, N11057);
not NOT1 (N12049, N12037);
and AND4 (N12050, N12043, N5731, N3192, N4026);
nor NOR3 (N12051, N12040, N5875, N1333);
nand NAND3 (N12052, N12051, N11680, N7773);
nand NAND3 (N12053, N12048, N581, N9444);
nand NAND3 (N12054, N12047, N11116, N3542);
nor NOR3 (N12055, N12045, N4056, N9215);
and AND2 (N12056, N12049, N8876);
or OR2 (N12057, N12054, N10570);
or OR3 (N12058, N12056, N7131, N10080);
nor NOR3 (N12059, N12041, N10045, N9876);
xor XOR2 (N12060, N12052, N9418);
nor NOR2 (N12061, N12057, N321);
or OR2 (N12062, N12060, N7818);
nand NAND3 (N12063, N12055, N1680, N11599);
not NOT1 (N12064, N12061);
and AND2 (N12065, N12050, N3174);
nor NOR3 (N12066, N12065, N5130, N5534);
nand NAND4 (N12067, N12033, N7233, N4153, N101);
nand NAND3 (N12068, N12067, N3079, N6829);
not NOT1 (N12069, N12068);
nand NAND4 (N12070, N12069, N11087, N2242, N796);
and AND2 (N12071, N12046, N5068);
or OR3 (N12072, N12058, N3710, N661);
and AND4 (N12073, N12062, N5889, N2749, N3540);
nor NOR3 (N12074, N12072, N5239, N11587);
or OR4 (N12075, N12044, N2426, N4482, N4831);
nand NAND2 (N12076, N12070, N10220);
buf BUF1 (N12077, N12074);
and AND3 (N12078, N12066, N7905, N3057);
not NOT1 (N12079, N12064);
not NOT1 (N12080, N12071);
or OR4 (N12081, N12080, N2073, N7211, N1867);
xor XOR2 (N12082, N12079, N11456);
xor XOR2 (N12083, N12081, N4109);
nand NAND4 (N12084, N12083, N1861, N594, N9811);
nor NOR3 (N12085, N12077, N7387, N11787);
nor NOR2 (N12086, N12073, N11740);
xor XOR2 (N12087, N12059, N5821);
buf BUF1 (N12088, N12086);
not NOT1 (N12089, N12053);
nand NAND3 (N12090, N12088, N11084, N6012);
nor NOR3 (N12091, N12085, N7026, N11791);
and AND2 (N12092, N12075, N9084);
or OR3 (N12093, N12091, N4495, N10265);
and AND4 (N12094, N12078, N11110, N11841, N1510);
and AND3 (N12095, N12092, N5784, N5496);
and AND3 (N12096, N12090, N5854, N5130);
buf BUF1 (N12097, N12076);
nand NAND2 (N12098, N12082, N6448);
or OR4 (N12099, N12094, N8225, N1707, N520);
and AND4 (N12100, N12095, N9536, N1102, N10864);
nand NAND3 (N12101, N12099, N4681, N5726);
nor NOR2 (N12102, N12097, N683);
nor NOR2 (N12103, N12101, N9000);
buf BUF1 (N12104, N12084);
nor NOR4 (N12105, N12087, N5113, N7586, N2700);
and AND2 (N12106, N12096, N8211);
nand NAND4 (N12107, N12089, N3143, N3032, N3795);
nor NOR4 (N12108, N12063, N7723, N3023, N7415);
nor NOR2 (N12109, N12102, N995);
nand NAND4 (N12110, N12093, N5280, N3900, N11398);
not NOT1 (N12111, N12107);
nor NOR3 (N12112, N12108, N1351, N1676);
xor XOR2 (N12113, N12112, N5469);
xor XOR2 (N12114, N12104, N4496);
and AND3 (N12115, N12110, N724, N1373);
nand NAND4 (N12116, N12115, N6363, N10806, N3681);
xor XOR2 (N12117, N12103, N4094);
and AND3 (N12118, N12114, N4768, N2742);
nand NAND3 (N12119, N12109, N10627, N1337);
xor XOR2 (N12120, N12100, N11707);
xor XOR2 (N12121, N12116, N11942);
buf BUF1 (N12122, N12117);
xor XOR2 (N12123, N12118, N5974);
nor NOR4 (N12124, N12098, N9436, N2866, N3936);
buf BUF1 (N12125, N12113);
nor NOR4 (N12126, N12123, N6680, N3100, N2398);
buf BUF1 (N12127, N12106);
and AND4 (N12128, N12105, N531, N6326, N11262);
xor XOR2 (N12129, N12128, N10238);
xor XOR2 (N12130, N12125, N3643);
and AND2 (N12131, N12120, N8047);
nor NOR3 (N12132, N12126, N2981, N9296);
xor XOR2 (N12133, N12129, N1561);
buf BUF1 (N12134, N12127);
and AND4 (N12135, N12131, N8024, N7304, N2905);
or OR3 (N12136, N12111, N4015, N1141);
not NOT1 (N12137, N12119);
not NOT1 (N12138, N12133);
or OR4 (N12139, N12122, N5575, N5913, N7429);
not NOT1 (N12140, N12134);
nor NOR3 (N12141, N12130, N2857, N2104);
xor XOR2 (N12142, N12136, N12117);
not NOT1 (N12143, N12138);
nor NOR2 (N12144, N12143, N615);
buf BUF1 (N12145, N12124);
not NOT1 (N12146, N12137);
or OR4 (N12147, N12140, N10475, N7287, N8427);
nand NAND3 (N12148, N12142, N9551, N9965);
nor NOR4 (N12149, N12121, N2738, N10483, N5498);
buf BUF1 (N12150, N12144);
nor NOR4 (N12151, N12150, N6487, N6321, N6929);
xor XOR2 (N12152, N12145, N3841);
buf BUF1 (N12153, N12139);
or OR2 (N12154, N12146, N3306);
or OR2 (N12155, N12153, N10884);
xor XOR2 (N12156, N12148, N7981);
xor XOR2 (N12157, N12149, N8295);
buf BUF1 (N12158, N12141);
xor XOR2 (N12159, N12155, N4442);
nor NOR3 (N12160, N12157, N11566, N2166);
not NOT1 (N12161, N12154);
not NOT1 (N12162, N12151);
nor NOR4 (N12163, N12158, N11015, N734, N5156);
nand NAND3 (N12164, N12156, N145, N8261);
and AND4 (N12165, N12132, N7601, N9318, N2487);
not NOT1 (N12166, N12159);
not NOT1 (N12167, N12163);
nand NAND3 (N12168, N12164, N10387, N11379);
buf BUF1 (N12169, N12147);
and AND2 (N12170, N12152, N5721);
nor NOR2 (N12171, N12167, N12100);
nor NOR2 (N12172, N12171, N915);
buf BUF1 (N12173, N12162);
or OR2 (N12174, N12135, N5516);
and AND2 (N12175, N12161, N9925);
buf BUF1 (N12176, N12169);
xor XOR2 (N12177, N12172, N2274);
nor NOR3 (N12178, N12177, N3858, N10711);
nand NAND4 (N12179, N12175, N6063, N6336, N11594);
or OR4 (N12180, N12170, N2688, N5662, N8783);
or OR3 (N12181, N12166, N11598, N3484);
not NOT1 (N12182, N12180);
buf BUF1 (N12183, N12174);
xor XOR2 (N12184, N12176, N11497);
nand NAND2 (N12185, N12181, N8208);
or OR4 (N12186, N12165, N9586, N2717, N710);
xor XOR2 (N12187, N12178, N6502);
not NOT1 (N12188, N12187);
not NOT1 (N12189, N12188);
nor NOR2 (N12190, N12184, N2057);
xor XOR2 (N12191, N12186, N4671);
buf BUF1 (N12192, N12173);
buf BUF1 (N12193, N12185);
or OR3 (N12194, N12168, N506, N4246);
nand NAND3 (N12195, N12190, N6569, N4166);
buf BUF1 (N12196, N12193);
xor XOR2 (N12197, N12192, N4167);
nor NOR3 (N12198, N12194, N11720, N11081);
or OR2 (N12199, N12198, N7452);
not NOT1 (N12200, N12183);
or OR3 (N12201, N12191, N8843, N5756);
nor NOR3 (N12202, N12199, N11788, N2259);
not NOT1 (N12203, N12200);
nand NAND3 (N12204, N12195, N3211, N11889);
xor XOR2 (N12205, N12179, N8792);
and AND2 (N12206, N12182, N7315);
not NOT1 (N12207, N12160);
nand NAND2 (N12208, N12201, N5232);
not NOT1 (N12209, N12207);
nor NOR4 (N12210, N12206, N4013, N9937, N5496);
xor XOR2 (N12211, N12197, N3289);
nor NOR4 (N12212, N12205, N11644, N1828, N11283);
xor XOR2 (N12213, N12203, N791);
buf BUF1 (N12214, N12208);
and AND4 (N12215, N12202, N7180, N35, N7996);
nand NAND4 (N12216, N12209, N6157, N6437, N6335);
or OR2 (N12217, N12214, N10815);
nor NOR2 (N12218, N12196, N7187);
or OR4 (N12219, N12216, N1514, N1834, N10901);
or OR4 (N12220, N12218, N5437, N9317, N1776);
nor NOR2 (N12221, N12210, N2364);
not NOT1 (N12222, N12213);
buf BUF1 (N12223, N12212);
buf BUF1 (N12224, N12219);
and AND4 (N12225, N12224, N4394, N5740, N3276);
and AND2 (N12226, N12211, N9836);
nand NAND4 (N12227, N12221, N5199, N1084, N1472);
xor XOR2 (N12228, N12204, N10914);
and AND3 (N12229, N12228, N9193, N8051);
nand NAND3 (N12230, N12215, N7549, N4090);
or OR3 (N12231, N12189, N9130, N96);
and AND4 (N12232, N12231, N3060, N5017, N7966);
buf BUF1 (N12233, N12217);
not NOT1 (N12234, N12227);
buf BUF1 (N12235, N12232);
or OR2 (N12236, N12222, N10379);
nor NOR2 (N12237, N12234, N388);
nand NAND3 (N12238, N12226, N5091, N6932);
xor XOR2 (N12239, N12223, N5534);
and AND2 (N12240, N12235, N2209);
and AND3 (N12241, N12225, N179, N2042);
nand NAND3 (N12242, N12220, N8915, N9727);
or OR2 (N12243, N12242, N4897);
or OR3 (N12244, N12237, N3010, N2558);
nand NAND3 (N12245, N12239, N3178, N4115);
xor XOR2 (N12246, N12240, N3065);
buf BUF1 (N12247, N12245);
xor XOR2 (N12248, N12238, N8225);
nand NAND4 (N12249, N12236, N11287, N6057, N9959);
or OR4 (N12250, N12233, N8848, N7194, N12157);
not NOT1 (N12251, N12241);
nand NAND2 (N12252, N12246, N8244);
nand NAND3 (N12253, N12250, N3156, N8574);
xor XOR2 (N12254, N12230, N6641);
xor XOR2 (N12255, N12248, N12125);
nand NAND2 (N12256, N12253, N10604);
and AND3 (N12257, N12256, N10641, N11462);
not NOT1 (N12258, N12252);
not NOT1 (N12259, N12257);
buf BUF1 (N12260, N12249);
nor NOR2 (N12261, N12244, N2392);
xor XOR2 (N12262, N12258, N10867);
or OR2 (N12263, N12229, N8120);
buf BUF1 (N12264, N12251);
nand NAND2 (N12265, N12260, N681);
and AND4 (N12266, N12259, N613, N6074, N2171);
xor XOR2 (N12267, N12264, N387);
or OR2 (N12268, N12243, N10633);
buf BUF1 (N12269, N12266);
nand NAND3 (N12270, N12261, N5072, N2117);
or OR2 (N12271, N12270, N3673);
nor NOR3 (N12272, N12268, N4176, N7170);
or OR4 (N12273, N12267, N7378, N7076, N6963);
or OR2 (N12274, N12255, N1778);
or OR3 (N12275, N12273, N12101, N4077);
and AND3 (N12276, N12269, N3552, N2459);
and AND3 (N12277, N12271, N7857, N2363);
nand NAND3 (N12278, N12276, N4139, N8487);
nor NOR2 (N12279, N12265, N808);
not NOT1 (N12280, N12262);
xor XOR2 (N12281, N12277, N2180);
not NOT1 (N12282, N12263);
not NOT1 (N12283, N12247);
nand NAND4 (N12284, N12281, N5758, N7188, N8026);
and AND4 (N12285, N12279, N10396, N421, N5585);
xor XOR2 (N12286, N12272, N4423);
nand NAND3 (N12287, N12280, N3578, N10804);
and AND3 (N12288, N12274, N8695, N4351);
and AND4 (N12289, N12254, N7240, N8500, N7849);
buf BUF1 (N12290, N12278);
buf BUF1 (N12291, N12289);
nand NAND3 (N12292, N12287, N9431, N2392);
or OR3 (N12293, N12290, N1188, N3133);
buf BUF1 (N12294, N12275);
nand NAND4 (N12295, N12292, N1805, N9978, N11870);
or OR2 (N12296, N12293, N11928);
not NOT1 (N12297, N12294);
nor NOR4 (N12298, N12291, N11447, N12258, N11905);
or OR3 (N12299, N12286, N4541, N799);
nor NOR4 (N12300, N12288, N869, N5108, N11123);
and AND2 (N12301, N12282, N7114);
buf BUF1 (N12302, N12298);
buf BUF1 (N12303, N12302);
nand NAND4 (N12304, N12284, N4023, N11167, N6856);
nand NAND3 (N12305, N12285, N2009, N9166);
buf BUF1 (N12306, N12304);
and AND2 (N12307, N12299, N3786);
not NOT1 (N12308, N12305);
and AND2 (N12309, N12300, N9432);
buf BUF1 (N12310, N12283);
nand NAND2 (N12311, N12295, N1239);
not NOT1 (N12312, N12311);
and AND4 (N12313, N12310, N8410, N102, N10653);
nand NAND2 (N12314, N12306, N2953);
not NOT1 (N12315, N12309);
or OR3 (N12316, N12303, N3140, N1475);
xor XOR2 (N12317, N12316, N10840);
and AND3 (N12318, N12315, N11406, N11061);
nand NAND2 (N12319, N12301, N1693);
nor NOR4 (N12320, N12319, N6979, N4909, N3296);
buf BUF1 (N12321, N12314);
and AND2 (N12322, N12318, N6841);
and AND3 (N12323, N12297, N9432, N7200);
and AND4 (N12324, N12323, N9159, N4024, N9361);
nor NOR2 (N12325, N12307, N47);
buf BUF1 (N12326, N12321);
xor XOR2 (N12327, N12324, N388);
xor XOR2 (N12328, N12296, N9070);
xor XOR2 (N12329, N12313, N4949);
not NOT1 (N12330, N12325);
buf BUF1 (N12331, N12322);
and AND2 (N12332, N12329, N9910);
nor NOR3 (N12333, N12332, N4305, N10068);
not NOT1 (N12334, N12331);
nor NOR3 (N12335, N12320, N12286, N7358);
nand NAND2 (N12336, N12333, N5116);
nor NOR3 (N12337, N12327, N5921, N4815);
xor XOR2 (N12338, N12326, N362);
xor XOR2 (N12339, N12338, N8922);
nor NOR4 (N12340, N12308, N8476, N1041, N8751);
and AND4 (N12341, N12312, N4961, N424, N11317);
or OR3 (N12342, N12330, N3882, N4293);
nor NOR2 (N12343, N12335, N4003);
nand NAND3 (N12344, N12328, N1501, N4731);
not NOT1 (N12345, N12341);
nor NOR4 (N12346, N12344, N11447, N4635, N398);
xor XOR2 (N12347, N12336, N8317);
nand NAND2 (N12348, N12347, N5352);
xor XOR2 (N12349, N12340, N10114);
and AND4 (N12350, N12334, N1622, N1838, N3055);
not NOT1 (N12351, N12350);
nand NAND3 (N12352, N12345, N3998, N8356);
xor XOR2 (N12353, N12343, N2001);
or OR2 (N12354, N12342, N11125);
not NOT1 (N12355, N12349);
xor XOR2 (N12356, N12337, N9498);
xor XOR2 (N12357, N12317, N2183);
xor XOR2 (N12358, N12351, N5944);
nand NAND3 (N12359, N12353, N3484, N8919);
and AND3 (N12360, N12359, N5657, N11181);
buf BUF1 (N12361, N12348);
or OR4 (N12362, N12352, N2605, N1399, N9606);
not NOT1 (N12363, N12357);
xor XOR2 (N12364, N12355, N10962);
xor XOR2 (N12365, N12358, N5530);
not NOT1 (N12366, N12362);
or OR3 (N12367, N12364, N7646, N6210);
nand NAND4 (N12368, N12363, N3206, N464, N1932);
nor NOR3 (N12369, N12356, N2860, N9997);
nand NAND2 (N12370, N12346, N7526);
not NOT1 (N12371, N12365);
and AND2 (N12372, N12369, N1012);
and AND3 (N12373, N12370, N11996, N4763);
nand NAND3 (N12374, N12366, N10029, N8422);
nor NOR4 (N12375, N12373, N2514, N7339, N7363);
xor XOR2 (N12376, N12339, N5482);
xor XOR2 (N12377, N12367, N4435);
xor XOR2 (N12378, N12354, N5328);
not NOT1 (N12379, N12378);
buf BUF1 (N12380, N12375);
xor XOR2 (N12381, N12380, N5551);
or OR2 (N12382, N12374, N2044);
not NOT1 (N12383, N12377);
nor NOR2 (N12384, N12383, N9180);
not NOT1 (N12385, N12381);
and AND2 (N12386, N12376, N1813);
nand NAND2 (N12387, N12371, N7735);
not NOT1 (N12388, N12385);
xor XOR2 (N12389, N12368, N9630);
nor NOR2 (N12390, N12361, N2617);
and AND4 (N12391, N12390, N5231, N1576, N6024);
buf BUF1 (N12392, N12379);
nand NAND4 (N12393, N12388, N12356, N9822, N4407);
not NOT1 (N12394, N12386);
xor XOR2 (N12395, N12393, N2419);
buf BUF1 (N12396, N12382);
and AND2 (N12397, N12387, N1424);
or OR3 (N12398, N12360, N8151, N8890);
nand NAND2 (N12399, N12384, N7401);
nor NOR2 (N12400, N12394, N5323);
nor NOR3 (N12401, N12389, N9060, N3281);
xor XOR2 (N12402, N12391, N2860);
buf BUF1 (N12403, N12399);
xor XOR2 (N12404, N12403, N12011);
buf BUF1 (N12405, N12402);
and AND3 (N12406, N12398, N4045, N1911);
buf BUF1 (N12407, N12372);
xor XOR2 (N12408, N12404, N4263);
not NOT1 (N12409, N12396);
or OR4 (N12410, N12400, N3396, N2108, N8005);
or OR3 (N12411, N12392, N3391, N139);
and AND3 (N12412, N12397, N1009, N1481);
xor XOR2 (N12413, N12407, N11742);
not NOT1 (N12414, N12409);
not NOT1 (N12415, N12395);
not NOT1 (N12416, N12401);
buf BUF1 (N12417, N12413);
nor NOR3 (N12418, N12412, N1090, N1620);
or OR4 (N12419, N12405, N10699, N11984, N5791);
or OR4 (N12420, N12418, N3302, N12075, N8179);
xor XOR2 (N12421, N12419, N1453);
nand NAND2 (N12422, N12414, N10501);
or OR2 (N12423, N12422, N5073);
buf BUF1 (N12424, N12406);
or OR4 (N12425, N12415, N5557, N7530, N2591);
xor XOR2 (N12426, N12425, N3772);
nor NOR3 (N12427, N12408, N4542, N64);
and AND2 (N12428, N12410, N11623);
or OR3 (N12429, N12428, N5608, N3249);
nor NOR2 (N12430, N12416, N9965);
nor NOR2 (N12431, N12426, N4625);
xor XOR2 (N12432, N12427, N1882);
xor XOR2 (N12433, N12432, N2237);
or OR2 (N12434, N12423, N6926);
xor XOR2 (N12435, N12434, N3702);
or OR4 (N12436, N12417, N2408, N8215, N9609);
buf BUF1 (N12437, N12421);
and AND3 (N12438, N12431, N1694, N8089);
and AND2 (N12439, N12420, N8335);
and AND4 (N12440, N12439, N5384, N10771, N2558);
or OR4 (N12441, N12411, N8254, N1859, N8560);
not NOT1 (N12442, N12438);
and AND3 (N12443, N12435, N3329, N3047);
buf BUF1 (N12444, N12429);
nand NAND3 (N12445, N12444, N8946, N2079);
nand NAND3 (N12446, N12433, N3740, N9834);
nor NOR2 (N12447, N12441, N10406);
xor XOR2 (N12448, N12424, N5301);
buf BUF1 (N12449, N12440);
and AND3 (N12450, N12447, N9150, N5468);
xor XOR2 (N12451, N12448, N242);
or OR2 (N12452, N12442, N9661);
xor XOR2 (N12453, N12443, N2757);
buf BUF1 (N12454, N12452);
nand NAND4 (N12455, N12450, N1420, N5636, N6072);
and AND4 (N12456, N12453, N4642, N8140, N5904);
buf BUF1 (N12457, N12430);
and AND2 (N12458, N12437, N890);
or OR3 (N12459, N12446, N4525, N7270);
nand NAND3 (N12460, N12458, N4827, N2526);
not NOT1 (N12461, N12457);
xor XOR2 (N12462, N12436, N8194);
nand NAND3 (N12463, N12455, N4657, N4219);
xor XOR2 (N12464, N12462, N11785);
xor XOR2 (N12465, N12445, N11643);
and AND4 (N12466, N12463, N8735, N12258, N9055);
and AND2 (N12467, N12451, N5701);
buf BUF1 (N12468, N12465);
not NOT1 (N12469, N12456);
or OR3 (N12470, N12454, N10513, N2564);
buf BUF1 (N12471, N12467);
nor NOR3 (N12472, N12469, N8095, N11750);
nand NAND3 (N12473, N12466, N9279, N5864);
and AND4 (N12474, N12472, N4880, N12337, N320);
buf BUF1 (N12475, N12449);
nor NOR4 (N12476, N12460, N7750, N4084, N7495);
xor XOR2 (N12477, N12459, N11847);
not NOT1 (N12478, N12470);
buf BUF1 (N12479, N12464);
not NOT1 (N12480, N12476);
buf BUF1 (N12481, N12461);
buf BUF1 (N12482, N12478);
nor NOR2 (N12483, N12468, N1574);
xor XOR2 (N12484, N12477, N2053);
nor NOR3 (N12485, N12473, N6804, N11927);
nor NOR2 (N12486, N12475, N6213);
xor XOR2 (N12487, N12483, N7792);
or OR4 (N12488, N12479, N363, N4432, N7039);
buf BUF1 (N12489, N12474);
nand NAND4 (N12490, N12480, N3794, N5049, N3708);
and AND4 (N12491, N12487, N6047, N10702, N3811);
nand NAND3 (N12492, N12485, N8691, N8479);
not NOT1 (N12493, N12492);
and AND4 (N12494, N12488, N3814, N6590, N11167);
and AND4 (N12495, N12490, N8074, N2851, N8768);
and AND2 (N12496, N12471, N5960);
or OR4 (N12497, N12482, N8475, N1996, N293);
or OR2 (N12498, N12491, N7867);
nor NOR2 (N12499, N12496, N4803);
not NOT1 (N12500, N12497);
buf BUF1 (N12501, N12489);
or OR4 (N12502, N12498, N10277, N7723, N10261);
nor NOR4 (N12503, N12495, N4248, N11727, N3191);
nand NAND2 (N12504, N12484, N1347);
buf BUF1 (N12505, N12504);
not NOT1 (N12506, N12500);
nor NOR3 (N12507, N12501, N8651, N3825);
and AND3 (N12508, N12494, N2282, N473);
or OR2 (N12509, N12481, N969);
and AND2 (N12510, N12486, N8860);
nor NOR2 (N12511, N12502, N12253);
buf BUF1 (N12512, N12507);
and AND3 (N12513, N12512, N11161, N7064);
nand NAND4 (N12514, N12503, N2172, N6764, N8867);
buf BUF1 (N12515, N12493);
buf BUF1 (N12516, N12513);
xor XOR2 (N12517, N12508, N3500);
or OR4 (N12518, N12506, N11470, N3413, N12298);
or OR3 (N12519, N12499, N9492, N9710);
nand NAND2 (N12520, N12518, N10757);
not NOT1 (N12521, N12515);
and AND3 (N12522, N12511, N1196, N7353);
nand NAND4 (N12523, N12521, N7728, N3552, N8291);
or OR4 (N12524, N12505, N11369, N2987, N4008);
not NOT1 (N12525, N12524);
xor XOR2 (N12526, N12523, N3168);
or OR3 (N12527, N12519, N10811, N5865);
nand NAND3 (N12528, N12525, N7297, N12181);
not NOT1 (N12529, N12517);
or OR4 (N12530, N12516, N12129, N2777, N277);
nor NOR4 (N12531, N12522, N4343, N7688, N3481);
buf BUF1 (N12532, N12527);
or OR2 (N12533, N12531, N10649);
not NOT1 (N12534, N12532);
xor XOR2 (N12535, N12533, N10336);
nand NAND3 (N12536, N12528, N167, N872);
xor XOR2 (N12537, N12509, N9572);
not NOT1 (N12538, N12537);
and AND3 (N12539, N12530, N11529, N7725);
nand NAND3 (N12540, N12514, N7888, N5972);
nand NAND3 (N12541, N12540, N4960, N4719);
nor NOR3 (N12542, N12536, N11517, N9144);
and AND3 (N12543, N12520, N183, N5850);
buf BUF1 (N12544, N12534);
xor XOR2 (N12545, N12542, N9594);
or OR2 (N12546, N12529, N6074);
or OR4 (N12547, N12545, N12432, N8387, N7016);
or OR3 (N12548, N12510, N3189, N6960);
nand NAND4 (N12549, N12548, N8002, N4642, N6468);
or OR3 (N12550, N12526, N6913, N5363);
nand NAND3 (N12551, N12541, N10886, N1027);
nand NAND2 (N12552, N12550, N1773);
nand NAND2 (N12553, N12551, N11828);
and AND4 (N12554, N12553, N2423, N7116, N7978);
buf BUF1 (N12555, N12549);
xor XOR2 (N12556, N12546, N7186);
buf BUF1 (N12557, N12539);
buf BUF1 (N12558, N12557);
nand NAND3 (N12559, N12552, N386, N3999);
nor NOR2 (N12560, N12555, N11170);
or OR2 (N12561, N12543, N10209);
and AND3 (N12562, N12547, N6300, N4002);
and AND2 (N12563, N12535, N6946);
xor XOR2 (N12564, N12556, N10896);
nor NOR3 (N12565, N12560, N12485, N8346);
or OR2 (N12566, N12563, N1814);
nand NAND2 (N12567, N12558, N452);
buf BUF1 (N12568, N12561);
or OR3 (N12569, N12562, N4314, N2337);
and AND4 (N12570, N12569, N2962, N3884, N4143);
buf BUF1 (N12571, N12565);
or OR3 (N12572, N12538, N11699, N691);
xor XOR2 (N12573, N12567, N3188);
not NOT1 (N12574, N12544);
nand NAND4 (N12575, N12573, N2759, N10180, N1466);
xor XOR2 (N12576, N12571, N11631);
or OR2 (N12577, N12576, N2346);
nand NAND2 (N12578, N12566, N8838);
xor XOR2 (N12579, N12572, N5291);
and AND3 (N12580, N12564, N352, N7042);
nor NOR3 (N12581, N12559, N5774, N203);
nor NOR3 (N12582, N12580, N369, N7360);
not NOT1 (N12583, N12575);
and AND4 (N12584, N12578, N2658, N6458, N6062);
not NOT1 (N12585, N12574);
buf BUF1 (N12586, N12570);
or OR3 (N12587, N12584, N9424, N11516);
xor XOR2 (N12588, N12579, N375);
xor XOR2 (N12589, N12587, N2423);
nand NAND3 (N12590, N12586, N434, N12404);
nor NOR2 (N12591, N12589, N11280);
or OR2 (N12592, N12583, N2101);
xor XOR2 (N12593, N12581, N10213);
nor NOR4 (N12594, N12577, N480, N7625, N7889);
nand NAND4 (N12595, N12568, N9172, N5984, N10128);
xor XOR2 (N12596, N12595, N12009);
not NOT1 (N12597, N12585);
xor XOR2 (N12598, N12593, N3440);
nand NAND3 (N12599, N12597, N11547, N8644);
or OR4 (N12600, N12596, N6465, N2379, N12059);
nand NAND3 (N12601, N12594, N10354, N1060);
or OR2 (N12602, N12588, N4578);
nand NAND4 (N12603, N12582, N462, N4732, N8071);
nor NOR4 (N12604, N12591, N1204, N2474, N12059);
xor XOR2 (N12605, N12599, N3942);
nand NAND3 (N12606, N12603, N2907, N6124);
or OR3 (N12607, N12605, N4682, N7303);
nor NOR3 (N12608, N12598, N1296, N11310);
and AND2 (N12609, N12608, N7714);
buf BUF1 (N12610, N12607);
buf BUF1 (N12611, N12609);
nor NOR4 (N12612, N12602, N8822, N4578, N7466);
nor NOR3 (N12613, N12601, N913, N8644);
buf BUF1 (N12614, N12612);
nor NOR3 (N12615, N12604, N2036, N9184);
and AND3 (N12616, N12610, N5279, N2649);
and AND2 (N12617, N12590, N11518);
and AND2 (N12618, N12554, N10657);
buf BUF1 (N12619, N12606);
nand NAND2 (N12620, N12615, N12463);
and AND3 (N12621, N12611, N2513, N5790);
nor NOR2 (N12622, N12619, N10029);
nand NAND4 (N12623, N12613, N1107, N6313, N5574);
not NOT1 (N12624, N12617);
and AND2 (N12625, N12592, N1995);
and AND4 (N12626, N12625, N8868, N10845, N743);
or OR4 (N12627, N12626, N929, N790, N6108);
and AND4 (N12628, N12616, N2749, N4912, N491);
nand NAND3 (N12629, N12627, N4943, N7365);
nand NAND2 (N12630, N12629, N6240);
buf BUF1 (N12631, N12621);
nand NAND3 (N12632, N12618, N12625, N2166);
or OR3 (N12633, N12624, N9306, N1740);
buf BUF1 (N12634, N12600);
not NOT1 (N12635, N12628);
not NOT1 (N12636, N12633);
or OR3 (N12637, N12614, N2747, N9003);
and AND4 (N12638, N12637, N4295, N9287, N1325);
nand NAND4 (N12639, N12631, N373, N3993, N1183);
and AND4 (N12640, N12634, N11581, N1954, N9438);
nor NOR3 (N12641, N12630, N6234, N5100);
and AND4 (N12642, N12632, N2558, N5884, N6920);
not NOT1 (N12643, N12620);
nand NAND4 (N12644, N12638, N3750, N4598, N8026);
not NOT1 (N12645, N12639);
not NOT1 (N12646, N12622);
not NOT1 (N12647, N12623);
not NOT1 (N12648, N12641);
xor XOR2 (N12649, N12642, N4339);
buf BUF1 (N12650, N12636);
nand NAND2 (N12651, N12643, N11144);
buf BUF1 (N12652, N12648);
xor XOR2 (N12653, N12646, N11451);
and AND4 (N12654, N12649, N7448, N12555, N11178);
not NOT1 (N12655, N12644);
nand NAND4 (N12656, N12652, N2676, N9204, N11084);
nor NOR2 (N12657, N12656, N11128);
nand NAND2 (N12658, N12651, N9458);
not NOT1 (N12659, N12658);
nor NOR3 (N12660, N12654, N1495, N830);
not NOT1 (N12661, N12650);
not NOT1 (N12662, N12661);
nor NOR3 (N12663, N12640, N3614, N2638);
or OR3 (N12664, N12647, N8806, N8156);
or OR4 (N12665, N12653, N8858, N2663, N2583);
and AND4 (N12666, N12663, N6523, N3939, N11464);
and AND3 (N12667, N12655, N9217, N1398);
nor NOR3 (N12668, N12664, N334, N8919);
xor XOR2 (N12669, N12668, N2622);
nor NOR4 (N12670, N12669, N9839, N5362, N9918);
or OR4 (N12671, N12670, N8960, N12097, N6464);
buf BUF1 (N12672, N12666);
buf BUF1 (N12673, N12645);
nand NAND4 (N12674, N12667, N7315, N5960, N8073);
not NOT1 (N12675, N12665);
nor NOR2 (N12676, N12635, N4458);
buf BUF1 (N12677, N12657);
buf BUF1 (N12678, N12677);
xor XOR2 (N12679, N12671, N12135);
buf BUF1 (N12680, N12676);
xor XOR2 (N12681, N12673, N11652);
xor XOR2 (N12682, N12662, N12455);
or OR2 (N12683, N12678, N7077);
or OR2 (N12684, N12672, N3164);
and AND2 (N12685, N12683, N8588);
and AND4 (N12686, N12674, N4954, N8680, N877);
buf BUF1 (N12687, N12680);
and AND4 (N12688, N12679, N5096, N7948, N6399);
nand NAND4 (N12689, N12660, N2471, N12604, N1359);
not NOT1 (N12690, N12659);
buf BUF1 (N12691, N12688);
or OR2 (N12692, N12681, N9059);
nand NAND3 (N12693, N12686, N1416, N4446);
and AND4 (N12694, N12693, N9477, N5851, N4917);
nor NOR3 (N12695, N12685, N10414, N2705);
not NOT1 (N12696, N12694);
xor XOR2 (N12697, N12675, N8743);
nor NOR2 (N12698, N12697, N10617);
nand NAND2 (N12699, N12690, N11745);
or OR4 (N12700, N12687, N1749, N1499, N11222);
buf BUF1 (N12701, N12700);
nand NAND3 (N12702, N12701, N7184, N9059);
or OR4 (N12703, N12684, N855, N5839, N4607);
buf BUF1 (N12704, N12691);
buf BUF1 (N12705, N12696);
not NOT1 (N12706, N12695);
nand NAND3 (N12707, N12702, N4218, N9605);
and AND2 (N12708, N12707, N4193);
and AND4 (N12709, N12704, N2337, N8510, N10147);
and AND3 (N12710, N12689, N9057, N6527);
buf BUF1 (N12711, N12708);
nand NAND4 (N12712, N12705, N11375, N1783, N5342);
nor NOR3 (N12713, N12682, N8182, N450);
buf BUF1 (N12714, N12713);
nand NAND3 (N12715, N12714, N6846, N8169);
or OR2 (N12716, N12698, N9597);
not NOT1 (N12717, N12711);
or OR3 (N12718, N12712, N9169, N6754);
and AND2 (N12719, N12715, N11228);
buf BUF1 (N12720, N12703);
or OR2 (N12721, N12720, N441);
not NOT1 (N12722, N12709);
nor NOR4 (N12723, N12706, N10849, N4621, N11693);
not NOT1 (N12724, N12723);
xor XOR2 (N12725, N12717, N3878);
xor XOR2 (N12726, N12692, N12581);
nand NAND2 (N12727, N12724, N9901);
xor XOR2 (N12728, N12722, N2847);
and AND3 (N12729, N12725, N5209, N5948);
buf BUF1 (N12730, N12729);
nand NAND4 (N12731, N12699, N850, N8350, N9951);
nor NOR3 (N12732, N12728, N2086, N9055);
not NOT1 (N12733, N12721);
buf BUF1 (N12734, N12716);
buf BUF1 (N12735, N12734);
not NOT1 (N12736, N12719);
nor NOR4 (N12737, N12727, N961, N2651, N11868);
buf BUF1 (N12738, N12731);
xor XOR2 (N12739, N12710, N9897);
and AND2 (N12740, N12736, N9320);
nand NAND3 (N12741, N12739, N1773, N9042);
and AND4 (N12742, N12735, N11555, N6281, N7324);
buf BUF1 (N12743, N12741);
buf BUF1 (N12744, N12726);
or OR3 (N12745, N12718, N3820, N1117);
xor XOR2 (N12746, N12744, N4267);
and AND4 (N12747, N12733, N2185, N3947, N9300);
and AND3 (N12748, N12738, N6410, N10895);
and AND3 (N12749, N12748, N7172, N5664);
and AND2 (N12750, N12747, N5322);
nand NAND3 (N12751, N12732, N420, N6655);
xor XOR2 (N12752, N12745, N8974);
xor XOR2 (N12753, N12746, N2971);
or OR2 (N12754, N12750, N6505);
or OR4 (N12755, N12743, N9382, N2573, N10786);
xor XOR2 (N12756, N12730, N4191);
or OR3 (N12757, N12737, N9810, N6149);
or OR4 (N12758, N12751, N10570, N5522, N2753);
nor NOR4 (N12759, N12742, N4931, N2606, N7534);
buf BUF1 (N12760, N12753);
xor XOR2 (N12761, N12759, N7349);
or OR4 (N12762, N12740, N11162, N3009, N4744);
nand NAND3 (N12763, N12757, N12725, N4535);
buf BUF1 (N12764, N12762);
buf BUF1 (N12765, N12752);
not NOT1 (N12766, N12765);
nand NAND3 (N12767, N12756, N10804, N12264);
xor XOR2 (N12768, N12767, N4479);
xor XOR2 (N12769, N12768, N10885);
not NOT1 (N12770, N12761);
xor XOR2 (N12771, N12763, N572);
xor XOR2 (N12772, N12764, N1539);
or OR3 (N12773, N12754, N10566, N3269);
or OR4 (N12774, N12770, N11250, N4111, N6628);
nand NAND3 (N12775, N12766, N5260, N4249);
xor XOR2 (N12776, N12772, N980);
or OR3 (N12777, N12773, N11985, N11995);
buf BUF1 (N12778, N12774);
and AND4 (N12779, N12777, N3837, N8545, N6858);
xor XOR2 (N12780, N12776, N2617);
or OR2 (N12781, N12780, N11692);
buf BUF1 (N12782, N12779);
and AND2 (N12783, N12778, N6792);
and AND4 (N12784, N12782, N11633, N7587, N6679);
nor NOR4 (N12785, N12769, N3000, N7353, N5769);
not NOT1 (N12786, N12783);
xor XOR2 (N12787, N12781, N9680);
and AND3 (N12788, N12755, N2346, N2649);
nor NOR2 (N12789, N12775, N9340);
and AND3 (N12790, N12760, N5449, N10575);
nor NOR3 (N12791, N12758, N8149, N2746);
not NOT1 (N12792, N12785);
or OR2 (N12793, N12787, N12519);
and AND3 (N12794, N12749, N7812, N1396);
xor XOR2 (N12795, N12792, N12293);
buf BUF1 (N12796, N12771);
nor NOR3 (N12797, N12791, N4886, N8946);
buf BUF1 (N12798, N12786);
nor NOR3 (N12799, N12788, N9773, N1856);
and AND3 (N12800, N12797, N6087, N640);
buf BUF1 (N12801, N12794);
buf BUF1 (N12802, N12799);
buf BUF1 (N12803, N12798);
or OR4 (N12804, N12796, N11795, N10393, N876);
not NOT1 (N12805, N12802);
nand NAND3 (N12806, N12801, N6230, N5569);
buf BUF1 (N12807, N12784);
nand NAND2 (N12808, N12806, N229);
or OR2 (N12809, N12805, N11323);
nand NAND4 (N12810, N12789, N2183, N2836, N12523);
nand NAND3 (N12811, N12790, N3222, N3045);
nor NOR3 (N12812, N12803, N10770, N9312);
nand NAND3 (N12813, N12800, N8534, N7250);
xor XOR2 (N12814, N12810, N9792);
nand NAND3 (N12815, N12811, N824, N8156);
buf BUF1 (N12816, N12813);
xor XOR2 (N12817, N12809, N8904);
or OR3 (N12818, N12815, N12442, N2844);
or OR2 (N12819, N12807, N4989);
and AND2 (N12820, N12819, N1521);
nor NOR2 (N12821, N12804, N10086);
xor XOR2 (N12822, N12814, N6044);
nor NOR2 (N12823, N12812, N1282);
or OR4 (N12824, N12795, N1270, N6658, N4142);
nand NAND2 (N12825, N12816, N2182);
nand NAND3 (N12826, N12820, N6932, N1808);
and AND4 (N12827, N12817, N9253, N7281, N6656);
nand NAND2 (N12828, N12823, N2278);
xor XOR2 (N12829, N12821, N6231);
or OR2 (N12830, N12828, N4140);
xor XOR2 (N12831, N12829, N6763);
nand NAND3 (N12832, N12824, N9498, N9296);
buf BUF1 (N12833, N12830);
or OR2 (N12834, N12827, N12426);
and AND4 (N12835, N12818, N9949, N3999, N6143);
buf BUF1 (N12836, N12826);
buf BUF1 (N12837, N12834);
buf BUF1 (N12838, N12835);
buf BUF1 (N12839, N12832);
and AND4 (N12840, N12822, N968, N2169, N3993);
buf BUF1 (N12841, N12839);
nor NOR4 (N12842, N12837, N11424, N9141, N5749);
or OR4 (N12843, N12841, N11698, N11757, N1677);
or OR3 (N12844, N12843, N1094, N1807);
buf BUF1 (N12845, N12840);
xor XOR2 (N12846, N12845, N10687);
xor XOR2 (N12847, N12846, N11541);
xor XOR2 (N12848, N12831, N7985);
and AND4 (N12849, N12848, N12590, N11373, N11195);
xor XOR2 (N12850, N12849, N5083);
not NOT1 (N12851, N12825);
nor NOR4 (N12852, N12844, N8427, N9371, N1761);
nor NOR3 (N12853, N12793, N5307, N6683);
and AND3 (N12854, N12850, N1789, N10455);
nand NAND3 (N12855, N12852, N1593, N10760);
nor NOR2 (N12856, N12842, N1693);
not NOT1 (N12857, N12855);
nor NOR3 (N12858, N12851, N8913, N5992);
xor XOR2 (N12859, N12856, N6985);
and AND4 (N12860, N12853, N5155, N8794, N5598);
and AND4 (N12861, N12854, N719, N2607, N4798);
buf BUF1 (N12862, N12847);
or OR4 (N12863, N12859, N8000, N8700, N2161);
xor XOR2 (N12864, N12836, N5581);
nor NOR4 (N12865, N12858, N6809, N2043, N61);
not NOT1 (N12866, N12860);
nor NOR3 (N12867, N12862, N6947, N12340);
xor XOR2 (N12868, N12865, N10588);
or OR3 (N12869, N12867, N8748, N503);
buf BUF1 (N12870, N12857);
and AND4 (N12871, N12868, N5544, N2385, N4543);
nor NOR3 (N12872, N12866, N1831, N11447);
nand NAND3 (N12873, N12838, N882, N3767);
nand NAND4 (N12874, N12861, N8099, N10592, N10558);
buf BUF1 (N12875, N12872);
not NOT1 (N12876, N12863);
xor XOR2 (N12877, N12870, N8374);
or OR2 (N12878, N12808, N8687);
not NOT1 (N12879, N12833);
nand NAND3 (N12880, N12875, N150, N633);
nand NAND4 (N12881, N12873, N11765, N1111, N2962);
or OR3 (N12882, N12864, N1453, N1354);
and AND4 (N12883, N12879, N4318, N9941, N11552);
not NOT1 (N12884, N12880);
and AND2 (N12885, N12878, N5872);
not NOT1 (N12886, N12882);
or OR4 (N12887, N12883, N2738, N9455, N12314);
xor XOR2 (N12888, N12876, N3609);
and AND2 (N12889, N12885, N10552);
nor NOR3 (N12890, N12884, N1754, N5729);
and AND2 (N12891, N12889, N6703);
or OR3 (N12892, N12891, N11840, N4800);
buf BUF1 (N12893, N12877);
xor XOR2 (N12894, N12888, N9135);
nand NAND3 (N12895, N12869, N5549, N7280);
and AND3 (N12896, N12893, N6778, N8669);
xor XOR2 (N12897, N12896, N6009);
nand NAND4 (N12898, N12894, N2837, N7338, N3443);
nand NAND4 (N12899, N12881, N9952, N9725, N7880);
xor XOR2 (N12900, N12874, N6384);
xor XOR2 (N12901, N12897, N5998);
nand NAND4 (N12902, N12898, N3169, N11201, N2650);
or OR2 (N12903, N12871, N11868);
buf BUF1 (N12904, N12899);
and AND4 (N12905, N12900, N2418, N4481, N12206);
xor XOR2 (N12906, N12901, N3491);
or OR4 (N12907, N12905, N353, N12301, N1326);
and AND4 (N12908, N12890, N6549, N10742, N8078);
buf BUF1 (N12909, N12902);
xor XOR2 (N12910, N12909, N10661);
and AND3 (N12911, N12908, N9390, N998);
buf BUF1 (N12912, N12910);
nor NOR4 (N12913, N12911, N10311, N3983, N11607);
nand NAND4 (N12914, N12892, N1498, N544, N10286);
nor NOR3 (N12915, N12886, N4205, N5566);
xor XOR2 (N12916, N12895, N7399);
nand NAND4 (N12917, N12915, N10535, N6423, N5695);
buf BUF1 (N12918, N12903);
not NOT1 (N12919, N12912);
and AND2 (N12920, N12913, N5710);
not NOT1 (N12921, N12907);
and AND3 (N12922, N12920, N2507, N1898);
or OR2 (N12923, N12916, N3137);
nor NOR2 (N12924, N12906, N12274);
or OR3 (N12925, N12904, N6372, N6597);
nand NAND4 (N12926, N12887, N7988, N1479, N7675);
nor NOR4 (N12927, N12923, N2614, N9815, N7819);
buf BUF1 (N12928, N12918);
buf BUF1 (N12929, N12922);
buf BUF1 (N12930, N12914);
or OR4 (N12931, N12926, N117, N3365, N7701);
nand NAND2 (N12932, N12921, N5136);
not NOT1 (N12933, N12925);
nor NOR2 (N12934, N12932, N7690);
xor XOR2 (N12935, N12934, N12178);
or OR3 (N12936, N12931, N6472, N2730);
buf BUF1 (N12937, N12917);
xor XOR2 (N12938, N12937, N2116);
nor NOR2 (N12939, N12927, N11661);
xor XOR2 (N12940, N12930, N5548);
and AND4 (N12941, N12940, N4896, N8803, N7010);
and AND2 (N12942, N12933, N2549);
or OR4 (N12943, N12928, N5165, N11839, N8531);
not NOT1 (N12944, N12919);
nor NOR3 (N12945, N12942, N9872, N12238);
not NOT1 (N12946, N12936);
nand NAND2 (N12947, N12929, N2086);
not NOT1 (N12948, N12939);
nor NOR2 (N12949, N12941, N2988);
not NOT1 (N12950, N12924);
not NOT1 (N12951, N12945);
xor XOR2 (N12952, N12946, N10406);
nand NAND3 (N12953, N12947, N6822, N11531);
nor NOR4 (N12954, N12948, N2409, N10736, N2647);
buf BUF1 (N12955, N12952);
and AND2 (N12956, N12949, N8402);
buf BUF1 (N12957, N12944);
or OR3 (N12958, N12953, N10220, N6828);
not NOT1 (N12959, N12958);
nand NAND3 (N12960, N12956, N5539, N9208);
nand NAND4 (N12961, N12951, N10712, N9447, N11411);
or OR3 (N12962, N12954, N1626, N9694);
not NOT1 (N12963, N12961);
not NOT1 (N12964, N12950);
and AND3 (N12965, N12955, N9847, N6329);
xor XOR2 (N12966, N12938, N5004);
not NOT1 (N12967, N12960);
not NOT1 (N12968, N12959);
not NOT1 (N12969, N12963);
not NOT1 (N12970, N12968);
nor NOR2 (N12971, N12935, N8652);
xor XOR2 (N12972, N12966, N11250);
nor NOR4 (N12973, N12965, N8706, N9873, N1673);
or OR3 (N12974, N12967, N10923, N1759);
not NOT1 (N12975, N12943);
or OR3 (N12976, N12969, N4404, N484);
xor XOR2 (N12977, N12970, N277);
nand NAND4 (N12978, N12973, N9040, N4655, N6641);
not NOT1 (N12979, N12957);
and AND4 (N12980, N12972, N4429, N8887, N2593);
not NOT1 (N12981, N12975);
buf BUF1 (N12982, N12980);
nand NAND2 (N12983, N12976, N6550);
or OR3 (N12984, N12983, N3396, N6947);
buf BUF1 (N12985, N12962);
xor XOR2 (N12986, N12978, N3569);
nand NAND4 (N12987, N12986, N11809, N1262, N7625);
buf BUF1 (N12988, N12981);
and AND3 (N12989, N12988, N2194, N1477);
and AND4 (N12990, N12987, N5195, N12184, N6155);
or OR2 (N12991, N12984, N4817);
nor NOR4 (N12992, N12971, N12983, N12534, N8301);
xor XOR2 (N12993, N12985, N6416);
not NOT1 (N12994, N12991);
and AND3 (N12995, N12990, N6959, N6428);
not NOT1 (N12996, N12995);
not NOT1 (N12997, N12979);
nor NOR4 (N12998, N12997, N1664, N6643, N2751);
nand NAND2 (N12999, N12992, N4128);
not NOT1 (N13000, N12982);
xor XOR2 (N13001, N12993, N4725);
xor XOR2 (N13002, N13000, N521);
and AND2 (N13003, N12974, N3576);
buf BUF1 (N13004, N12964);
xor XOR2 (N13005, N12996, N12887);
xor XOR2 (N13006, N12994, N11065);
nor NOR3 (N13007, N13004, N11459, N8382);
or OR2 (N13008, N13005, N11124);
nor NOR2 (N13009, N12989, N4582);
nand NAND4 (N13010, N13009, N9389, N7710, N7631);
buf BUF1 (N13011, N12977);
nand NAND2 (N13012, N13003, N11256);
or OR3 (N13013, N13007, N1072, N6026);
and AND3 (N13014, N13001, N12660, N1849);
xor XOR2 (N13015, N13012, N12324);
buf BUF1 (N13016, N13013);
xor XOR2 (N13017, N13016, N5710);
nor NOR2 (N13018, N13006, N5976);
xor XOR2 (N13019, N13015, N4754);
and AND4 (N13020, N13014, N11771, N6147, N3485);
nor NOR3 (N13021, N13020, N12327, N11234);
nand NAND4 (N13022, N13002, N8414, N10500, N3974);
nor NOR2 (N13023, N13022, N3423);
or OR3 (N13024, N13019, N11780, N4411);
and AND3 (N13025, N13010, N7705, N1660);
nor NOR3 (N13026, N12998, N6005, N5644);
nand NAND4 (N13027, N13023, N9557, N7787, N2289);
not NOT1 (N13028, N13027);
and AND3 (N13029, N13024, N7148, N7174);
and AND3 (N13030, N13021, N2272, N2033);
and AND4 (N13031, N13028, N1560, N8347, N11367);
and AND2 (N13032, N13017, N7982);
xor XOR2 (N13033, N13031, N999);
nand NAND3 (N13034, N13032, N9980, N8149);
not NOT1 (N13035, N13030);
nor NOR2 (N13036, N13011, N4667);
or OR4 (N13037, N12999, N10061, N8577, N7587);
and AND2 (N13038, N13033, N3021);
buf BUF1 (N13039, N13008);
nor NOR3 (N13040, N13037, N9498, N85);
not NOT1 (N13041, N13018);
nor NOR3 (N13042, N13034, N2773, N1045);
nand NAND2 (N13043, N13041, N3854);
nand NAND3 (N13044, N13038, N9097, N4799);
and AND2 (N13045, N13044, N11932);
xor XOR2 (N13046, N13036, N9126);
xor XOR2 (N13047, N13025, N9456);
buf BUF1 (N13048, N13042);
and AND3 (N13049, N13035, N10479, N853);
buf BUF1 (N13050, N13039);
nand NAND2 (N13051, N13043, N5626);
nor NOR2 (N13052, N13047, N3364);
nor NOR4 (N13053, N13048, N12628, N3900, N10327);
xor XOR2 (N13054, N13045, N9122);
and AND3 (N13055, N13051, N4323, N8097);
xor XOR2 (N13056, N13029, N10180);
not NOT1 (N13057, N13053);
nand NAND2 (N13058, N13040, N2226);
and AND3 (N13059, N13026, N7861, N4407);
and AND4 (N13060, N13052, N4661, N95, N10876);
not NOT1 (N13061, N13055);
or OR2 (N13062, N13059, N9790);
or OR4 (N13063, N13054, N3396, N5894, N5413);
not NOT1 (N13064, N13057);
or OR3 (N13065, N13062, N643, N11301);
xor XOR2 (N13066, N13063, N3274);
not NOT1 (N13067, N13058);
buf BUF1 (N13068, N13064);
not NOT1 (N13069, N13050);
nand NAND4 (N13070, N13067, N8647, N7090, N11029);
nand NAND3 (N13071, N13069, N5808, N9775);
nand NAND3 (N13072, N13060, N8794, N12288);
buf BUF1 (N13073, N13049);
xor XOR2 (N13074, N13073, N12887);
nor NOR4 (N13075, N13046, N142, N5697, N6997);
nand NAND3 (N13076, N13056, N336, N2932);
xor XOR2 (N13077, N13071, N4689);
or OR2 (N13078, N13068, N7087);
buf BUF1 (N13079, N13065);
nor NOR2 (N13080, N13076, N333);
xor XOR2 (N13081, N13075, N8322);
xor XOR2 (N13082, N13074, N2837);
or OR3 (N13083, N13077, N8674, N6822);
not NOT1 (N13084, N13082);
not NOT1 (N13085, N13083);
buf BUF1 (N13086, N13084);
buf BUF1 (N13087, N13085);
xor XOR2 (N13088, N13078, N1683);
and AND4 (N13089, N13086, N10800, N10836, N12347);
and AND3 (N13090, N13080, N5770, N6491);
nor NOR4 (N13091, N13090, N7566, N13070, N5143);
not NOT1 (N13092, N6651);
xor XOR2 (N13093, N13081, N11488);
nand NAND2 (N13094, N13079, N10717);
and AND4 (N13095, N13061, N623, N8359, N6162);
buf BUF1 (N13096, N13094);
buf BUF1 (N13097, N13087);
not NOT1 (N13098, N13096);
not NOT1 (N13099, N13088);
buf BUF1 (N13100, N13091);
xor XOR2 (N13101, N13095, N8362);
nand NAND4 (N13102, N13066, N5034, N9459, N9121);
not NOT1 (N13103, N13099);
nor NOR3 (N13104, N13089, N5120, N2279);
nor NOR3 (N13105, N13103, N343, N840);
buf BUF1 (N13106, N13072);
or OR2 (N13107, N13106, N9827);
xor XOR2 (N13108, N13104, N4810);
nand NAND2 (N13109, N13092, N470);
and AND3 (N13110, N13100, N6683, N7377);
or OR2 (N13111, N13107, N8963);
nand NAND2 (N13112, N13105, N10788);
not NOT1 (N13113, N13102);
buf BUF1 (N13114, N13101);
not NOT1 (N13115, N13112);
and AND3 (N13116, N13111, N4210, N7437);
xor XOR2 (N13117, N13110, N6727);
and AND2 (N13118, N13117, N3388);
or OR2 (N13119, N13097, N6788);
nor NOR3 (N13120, N13109, N10920, N2503);
nand NAND2 (N13121, N13116, N9401);
and AND2 (N13122, N13098, N6575);
and AND3 (N13123, N13120, N1951, N9616);
nor NOR2 (N13124, N13113, N4459);
xor XOR2 (N13125, N13119, N1788);
buf BUF1 (N13126, N13108);
nor NOR2 (N13127, N13115, N7946);
nor NOR4 (N13128, N13126, N4623, N12211, N12550);
or OR2 (N13129, N13128, N7467);
nand NAND4 (N13130, N13127, N12759, N9896, N5007);
and AND2 (N13131, N13093, N4614);
or OR4 (N13132, N13129, N7919, N3781, N10488);
nor NOR3 (N13133, N13124, N11368, N9116);
nor NOR3 (N13134, N13130, N2986, N9294);
or OR2 (N13135, N13118, N184);
nor NOR4 (N13136, N13134, N3291, N5541, N6264);
or OR3 (N13137, N13123, N9934, N3753);
buf BUF1 (N13138, N13114);
or OR4 (N13139, N13125, N3808, N8831, N7909);
and AND2 (N13140, N13136, N10092);
xor XOR2 (N13141, N13122, N8740);
nor NOR3 (N13142, N13135, N8957, N5321);
buf BUF1 (N13143, N13133);
or OR2 (N13144, N13131, N12074);
xor XOR2 (N13145, N13138, N3093);
nor NOR2 (N13146, N13121, N10206);
nand NAND3 (N13147, N13140, N3696, N7445);
nand NAND2 (N13148, N13142, N11102);
nor NOR3 (N13149, N13141, N9348, N4372);
nand NAND3 (N13150, N13144, N6478, N1605);
nand NAND4 (N13151, N13150, N3913, N11478, N3325);
nor NOR2 (N13152, N13148, N3336);
nor NOR3 (N13153, N13139, N8684, N6343);
and AND2 (N13154, N13147, N3368);
not NOT1 (N13155, N13151);
nand NAND2 (N13156, N13153, N482);
not NOT1 (N13157, N13137);
or OR2 (N13158, N13143, N8465);
buf BUF1 (N13159, N13156);
or OR3 (N13160, N13154, N12714, N252);
nand NAND4 (N13161, N13160, N6299, N739, N8632);
xor XOR2 (N13162, N13132, N3994);
xor XOR2 (N13163, N13146, N4877);
buf BUF1 (N13164, N13159);
and AND3 (N13165, N13158, N11619, N2610);
and AND3 (N13166, N13162, N8478, N7388);
buf BUF1 (N13167, N13166);
nand NAND3 (N13168, N13157, N6036, N9240);
nor NOR3 (N13169, N13145, N2075, N2478);
nor NOR2 (N13170, N13167, N3407);
buf BUF1 (N13171, N13164);
not NOT1 (N13172, N13171);
nand NAND2 (N13173, N13170, N5822);
nor NOR2 (N13174, N13172, N2286);
nor NOR4 (N13175, N13161, N7160, N4629, N10635);
buf BUF1 (N13176, N13152);
not NOT1 (N13177, N13169);
nor NOR2 (N13178, N13173, N13102);
nor NOR4 (N13179, N13168, N9831, N4173, N5538);
xor XOR2 (N13180, N13178, N11838);
buf BUF1 (N13181, N13155);
xor XOR2 (N13182, N13176, N11290);
nor NOR2 (N13183, N13165, N12884);
not NOT1 (N13184, N13163);
nand NAND3 (N13185, N13181, N9045, N7457);
not NOT1 (N13186, N13183);
not NOT1 (N13187, N13182);
buf BUF1 (N13188, N13184);
and AND3 (N13189, N13179, N7564, N3737);
nand NAND4 (N13190, N13187, N12644, N12649, N6670);
and AND4 (N13191, N13177, N6160, N3694, N4287);
xor XOR2 (N13192, N13185, N7024);
nor NOR2 (N13193, N13192, N7127);
or OR4 (N13194, N13188, N7010, N12485, N2073);
buf BUF1 (N13195, N13191);
xor XOR2 (N13196, N13195, N11401);
and AND3 (N13197, N13149, N1718, N5295);
nand NAND3 (N13198, N13197, N13009, N2110);
nor NOR4 (N13199, N13189, N3073, N372, N2441);
xor XOR2 (N13200, N13175, N3960);
and AND4 (N13201, N13186, N1815, N4940, N6551);
or OR3 (N13202, N13174, N6155, N5970);
nand NAND2 (N13203, N13196, N12608);
or OR2 (N13204, N13180, N11471);
buf BUF1 (N13205, N13202);
and AND3 (N13206, N13204, N11292, N9054);
xor XOR2 (N13207, N13200, N6551);
not NOT1 (N13208, N13198);
nand NAND3 (N13209, N13199, N7452, N10917);
and AND2 (N13210, N13203, N9446);
xor XOR2 (N13211, N13194, N9754);
buf BUF1 (N13212, N13190);
buf BUF1 (N13213, N13212);
or OR3 (N13214, N13213, N2546, N2549);
and AND2 (N13215, N13210, N3280);
or OR4 (N13216, N13211, N9723, N7583, N1655);
nand NAND2 (N13217, N13205, N8526);
xor XOR2 (N13218, N13214, N12169);
and AND3 (N13219, N13209, N8721, N10195);
buf BUF1 (N13220, N13217);
xor XOR2 (N13221, N13218, N8757);
nand NAND3 (N13222, N13208, N1079, N12365);
nand NAND2 (N13223, N13220, N11964);
xor XOR2 (N13224, N13206, N7006);
xor XOR2 (N13225, N13223, N129);
or OR2 (N13226, N13225, N11065);
buf BUF1 (N13227, N13219);
not NOT1 (N13228, N13207);
or OR3 (N13229, N13224, N2376, N4173);
or OR2 (N13230, N13221, N8538);
xor XOR2 (N13231, N13227, N12788);
not NOT1 (N13232, N13201);
nor NOR4 (N13233, N13229, N10584, N12489, N10849);
nand NAND3 (N13234, N13233, N626, N2159);
nor NOR4 (N13235, N13232, N11203, N8284, N1441);
xor XOR2 (N13236, N13215, N1155);
not NOT1 (N13237, N13230);
nor NOR2 (N13238, N13236, N636);
xor XOR2 (N13239, N13237, N13214);
not NOT1 (N13240, N13228);
or OR4 (N13241, N13238, N11518, N9867, N3606);
buf BUF1 (N13242, N13216);
or OR3 (N13243, N13240, N12278, N3027);
nor NOR3 (N13244, N13231, N10079, N9029);
buf BUF1 (N13245, N13242);
xor XOR2 (N13246, N13193, N9030);
nor NOR4 (N13247, N13226, N6198, N12790, N8441);
buf BUF1 (N13248, N13234);
xor XOR2 (N13249, N13241, N6389);
or OR3 (N13250, N13243, N8317, N3564);
nand NAND4 (N13251, N13245, N3467, N10874, N2022);
buf BUF1 (N13252, N13246);
and AND3 (N13253, N13248, N4941, N12661);
and AND2 (N13254, N13250, N5209);
or OR2 (N13255, N13247, N7714);
buf BUF1 (N13256, N13252);
nand NAND2 (N13257, N13256, N11107);
or OR2 (N13258, N13254, N8186);
buf BUF1 (N13259, N13244);
and AND2 (N13260, N13257, N3141);
nand NAND2 (N13261, N13249, N399);
or OR3 (N13262, N13251, N11727, N3957);
or OR2 (N13263, N13239, N2786);
and AND3 (N13264, N13263, N9582, N135);
or OR3 (N13265, N13235, N11365, N6392);
nand NAND2 (N13266, N13265, N9027);
not NOT1 (N13267, N13262);
not NOT1 (N13268, N13266);
not NOT1 (N13269, N13268);
or OR4 (N13270, N13259, N12459, N11499, N1518);
and AND4 (N13271, N13258, N6811, N8593, N2097);
not NOT1 (N13272, N13253);
nor NOR2 (N13273, N13222, N8626);
xor XOR2 (N13274, N13264, N9985);
not NOT1 (N13275, N13273);
or OR4 (N13276, N13275, N1923, N2611, N7801);
xor XOR2 (N13277, N13271, N12011);
not NOT1 (N13278, N13267);
buf BUF1 (N13279, N13274);
and AND3 (N13280, N13260, N11360, N3902);
and AND3 (N13281, N13278, N6187, N9387);
nor NOR3 (N13282, N13281, N2327, N1990);
or OR4 (N13283, N13279, N7791, N11864, N2435);
not NOT1 (N13284, N13255);
xor XOR2 (N13285, N13270, N4438);
buf BUF1 (N13286, N13283);
nand NAND4 (N13287, N13280, N12526, N5863, N5130);
or OR3 (N13288, N13285, N2330, N137);
nor NOR2 (N13289, N13272, N431);
nand NAND2 (N13290, N13284, N9909);
nand NAND3 (N13291, N13290, N9530, N7122);
buf BUF1 (N13292, N13282);
and AND4 (N13293, N13286, N12850, N5337, N3241);
buf BUF1 (N13294, N13269);
or OR4 (N13295, N13288, N10770, N11953, N12054);
not NOT1 (N13296, N13276);
xor XOR2 (N13297, N13289, N6222);
nand NAND3 (N13298, N13293, N8254, N4618);
not NOT1 (N13299, N13277);
not NOT1 (N13300, N13294);
or OR3 (N13301, N13300, N10170, N10671);
buf BUF1 (N13302, N13299);
buf BUF1 (N13303, N13287);
xor XOR2 (N13304, N13261, N2262);
or OR2 (N13305, N13301, N6972);
nand NAND4 (N13306, N13292, N11634, N10763, N9196);
or OR3 (N13307, N13304, N9304, N8670);
nand NAND2 (N13308, N13303, N4980);
nand NAND3 (N13309, N13295, N12468, N3985);
xor XOR2 (N13310, N13305, N5427);
and AND4 (N13311, N13297, N12649, N8862, N6491);
xor XOR2 (N13312, N13311, N2955);
xor XOR2 (N13313, N13309, N8890);
xor XOR2 (N13314, N13306, N1110);
or OR3 (N13315, N13310, N10358, N9592);
or OR3 (N13316, N13313, N2001, N2375);
nand NAND4 (N13317, N13315, N1288, N3397, N4743);
nand NAND4 (N13318, N13307, N4024, N2633, N8264);
buf BUF1 (N13319, N13296);
xor XOR2 (N13320, N13298, N565);
xor XOR2 (N13321, N13308, N3058);
not NOT1 (N13322, N13320);
not NOT1 (N13323, N13291);
xor XOR2 (N13324, N13321, N9420);
xor XOR2 (N13325, N13323, N7912);
and AND2 (N13326, N13319, N97);
not NOT1 (N13327, N13314);
buf BUF1 (N13328, N13327);
xor XOR2 (N13329, N13326, N11229);
or OR2 (N13330, N13325, N653);
or OR2 (N13331, N13302, N265);
and AND4 (N13332, N13330, N4201, N7171, N10124);
nor NOR3 (N13333, N13312, N7657, N3559);
buf BUF1 (N13334, N13322);
not NOT1 (N13335, N13318);
buf BUF1 (N13336, N13331);
not NOT1 (N13337, N13334);
nor NOR4 (N13338, N13333, N12491, N4088, N3870);
buf BUF1 (N13339, N13337);
nand NAND2 (N13340, N13336, N8748);
nand NAND3 (N13341, N13339, N12560, N8203);
buf BUF1 (N13342, N13341);
not NOT1 (N13343, N13340);
not NOT1 (N13344, N13342);
or OR3 (N13345, N13335, N4733, N7757);
xor XOR2 (N13346, N13316, N552);
and AND4 (N13347, N13338, N10174, N9392, N7085);
not NOT1 (N13348, N13332);
buf BUF1 (N13349, N13344);
nand NAND4 (N13350, N13343, N219, N6038, N5100);
buf BUF1 (N13351, N13347);
nor NOR4 (N13352, N13348, N9559, N9110, N4261);
or OR3 (N13353, N13346, N4102, N4566);
nor NOR4 (N13354, N13349, N4173, N8550, N12806);
and AND4 (N13355, N13324, N2082, N7091, N9269);
nor NOR4 (N13356, N13329, N1016, N372, N6901);
and AND4 (N13357, N13351, N7197, N5813, N13353);
xor XOR2 (N13358, N643, N7915);
nand NAND3 (N13359, N13355, N7313, N12378);
and AND3 (N13360, N13352, N11628, N11820);
not NOT1 (N13361, N13354);
nand NAND3 (N13362, N13328, N3255, N2628);
not NOT1 (N13363, N13361);
nand NAND4 (N13364, N13362, N1562, N3022, N659);
or OR3 (N13365, N13359, N12121, N3206);
nand NAND3 (N13366, N13360, N996, N9159);
buf BUF1 (N13367, N13365);
or OR2 (N13368, N13367, N6982);
xor XOR2 (N13369, N13364, N6935);
and AND4 (N13370, N13350, N8857, N12437, N9309);
not NOT1 (N13371, N13358);
not NOT1 (N13372, N13366);
or OR2 (N13373, N13371, N4872);
or OR3 (N13374, N13317, N3215, N6876);
not NOT1 (N13375, N13370);
not NOT1 (N13376, N13368);
and AND2 (N13377, N13357, N12624);
buf BUF1 (N13378, N13377);
nand NAND4 (N13379, N13376, N1125, N3972, N11696);
and AND3 (N13380, N13378, N11169, N11564);
xor XOR2 (N13381, N13372, N2193);
or OR4 (N13382, N13375, N10332, N7399, N8650);
xor XOR2 (N13383, N13381, N12957);
or OR3 (N13384, N13356, N4432, N11982);
nor NOR4 (N13385, N13363, N10673, N12275, N2682);
buf BUF1 (N13386, N13374);
xor XOR2 (N13387, N13379, N1221);
not NOT1 (N13388, N13345);
xor XOR2 (N13389, N13385, N5727);
nand NAND2 (N13390, N13382, N10009);
nand NAND3 (N13391, N13384, N394, N11075);
nand NAND2 (N13392, N13380, N4392);
or OR3 (N13393, N13389, N7612, N8209);
and AND3 (N13394, N13383, N6681, N3051);
xor XOR2 (N13395, N13386, N8956);
nand NAND2 (N13396, N13391, N7490);
and AND4 (N13397, N13395, N3754, N5112, N12192);
and AND2 (N13398, N13387, N566);
nand NAND3 (N13399, N13396, N2426, N8135);
buf BUF1 (N13400, N13392);
nor NOR2 (N13401, N13398, N4460);
buf BUF1 (N13402, N13390);
and AND3 (N13403, N13388, N2262, N9754);
xor XOR2 (N13404, N13397, N9715);
nand NAND3 (N13405, N13399, N7775, N548);
not NOT1 (N13406, N13369);
buf BUF1 (N13407, N13402);
or OR3 (N13408, N13373, N6085, N1660);
or OR4 (N13409, N13405, N4342, N8363, N7449);
nand NAND3 (N13410, N13394, N94, N9849);
nor NOR2 (N13411, N13404, N4200);
and AND2 (N13412, N13411, N3407);
buf BUF1 (N13413, N13412);
or OR3 (N13414, N13409, N2402, N5868);
buf BUF1 (N13415, N13393);
or OR2 (N13416, N13414, N4242);
nand NAND2 (N13417, N13410, N8444);
or OR2 (N13418, N13401, N230);
buf BUF1 (N13419, N13408);
nand NAND3 (N13420, N13400, N333, N8435);
buf BUF1 (N13421, N13415);
or OR3 (N13422, N13413, N1172, N5371);
or OR4 (N13423, N13418, N4993, N3913, N1615);
not NOT1 (N13424, N13422);
xor XOR2 (N13425, N13419, N13043);
not NOT1 (N13426, N13420);
buf BUF1 (N13427, N13425);
nor NOR3 (N13428, N13416, N1108, N5219);
buf BUF1 (N13429, N13417);
xor XOR2 (N13430, N13406, N6851);
not NOT1 (N13431, N13428);
buf BUF1 (N13432, N13430);
xor XOR2 (N13433, N13431, N9296);
buf BUF1 (N13434, N13427);
nor NOR4 (N13435, N13424, N11111, N5097, N10226);
xor XOR2 (N13436, N13403, N9555);
buf BUF1 (N13437, N13434);
not NOT1 (N13438, N13407);
or OR4 (N13439, N13433, N4558, N7143, N5066);
nor NOR3 (N13440, N13423, N12397, N4317);
or OR4 (N13441, N13437, N1041, N3881, N5237);
not NOT1 (N13442, N13438);
nand NAND3 (N13443, N13432, N11608, N12241);
xor XOR2 (N13444, N13426, N10938);
buf BUF1 (N13445, N13435);
nand NAND3 (N13446, N13440, N2726, N10920);
and AND3 (N13447, N13446, N5991, N3922);
buf BUF1 (N13448, N13443);
nand NAND3 (N13449, N13441, N1994, N103);
xor XOR2 (N13450, N13429, N9752);
xor XOR2 (N13451, N13445, N9364);
and AND2 (N13452, N13421, N6979);
and AND3 (N13453, N13436, N9401, N9610);
xor XOR2 (N13454, N13444, N2744);
xor XOR2 (N13455, N13448, N7308);
buf BUF1 (N13456, N13453);
nand NAND4 (N13457, N13454, N6, N6872, N5029);
nor NOR4 (N13458, N13450, N7120, N3901, N142);
or OR3 (N13459, N13452, N1419, N12790);
buf BUF1 (N13460, N13447);
buf BUF1 (N13461, N13455);
nand NAND3 (N13462, N13457, N5390, N10013);
not NOT1 (N13463, N13449);
and AND4 (N13464, N13439, N8701, N10463, N3287);
nand NAND2 (N13465, N13456, N6514);
nor NOR2 (N13466, N13462, N11601);
or OR4 (N13467, N13459, N8812, N4207, N3718);
and AND4 (N13468, N13466, N10532, N2456, N12229);
buf BUF1 (N13469, N13458);
xor XOR2 (N13470, N13469, N7164);
xor XOR2 (N13471, N13468, N12055);
xor XOR2 (N13472, N13451, N5296);
xor XOR2 (N13473, N13442, N6137);
or OR4 (N13474, N13460, N2274, N4412, N7904);
xor XOR2 (N13475, N13463, N9255);
buf BUF1 (N13476, N13461);
buf BUF1 (N13477, N13470);
nand NAND2 (N13478, N13471, N1440);
buf BUF1 (N13479, N13478);
not NOT1 (N13480, N13475);
nor NOR3 (N13481, N13479, N7801, N7067);
and AND4 (N13482, N13465, N13326, N13450, N9294);
or OR2 (N13483, N13481, N7087);
buf BUF1 (N13484, N13482);
buf BUF1 (N13485, N13473);
not NOT1 (N13486, N13476);
or OR4 (N13487, N13483, N1465, N3763, N6140);
nand NAND3 (N13488, N13485, N1707, N5746);
not NOT1 (N13489, N13477);
buf BUF1 (N13490, N13467);
or OR4 (N13491, N13488, N8840, N10693, N8365);
or OR4 (N13492, N13489, N3058, N1030, N8988);
or OR3 (N13493, N13490, N11970, N1852);
nand NAND2 (N13494, N13493, N2885);
not NOT1 (N13495, N13491);
nand NAND4 (N13496, N13492, N5209, N3955, N700);
buf BUF1 (N13497, N13487);
xor XOR2 (N13498, N13474, N9481);
or OR2 (N13499, N13495, N11);
and AND3 (N13500, N13464, N12381, N2721);
and AND2 (N13501, N13500, N2245);
buf BUF1 (N13502, N13486);
or OR2 (N13503, N13498, N5353);
and AND2 (N13504, N13494, N8351);
not NOT1 (N13505, N13501);
xor XOR2 (N13506, N13472, N5194);
not NOT1 (N13507, N13499);
not NOT1 (N13508, N13505);
xor XOR2 (N13509, N13503, N11403);
not NOT1 (N13510, N13504);
buf BUF1 (N13511, N13502);
nor NOR3 (N13512, N13509, N9346, N7940);
xor XOR2 (N13513, N13484, N9265);
nor NOR3 (N13514, N13506, N8332, N3048);
nor NOR2 (N13515, N13511, N1716);
nand NAND4 (N13516, N13512, N6864, N1716, N8222);
not NOT1 (N13517, N13480);
buf BUF1 (N13518, N13513);
nand NAND3 (N13519, N13510, N4711, N13083);
xor XOR2 (N13520, N13515, N6262);
not NOT1 (N13521, N13520);
not NOT1 (N13522, N13508);
nand NAND2 (N13523, N13507, N7554);
and AND4 (N13524, N13523, N5255, N1798, N9660);
buf BUF1 (N13525, N13524);
not NOT1 (N13526, N13516);
not NOT1 (N13527, N13497);
or OR3 (N13528, N13521, N7883, N6525);
and AND2 (N13529, N13522, N5658);
not NOT1 (N13530, N13518);
and AND2 (N13531, N13496, N3601);
and AND4 (N13532, N13514, N7500, N9406, N4914);
buf BUF1 (N13533, N13530);
xor XOR2 (N13534, N13528, N8979);
xor XOR2 (N13535, N13533, N13091);
xor XOR2 (N13536, N13525, N4686);
not NOT1 (N13537, N13519);
not NOT1 (N13538, N13526);
xor XOR2 (N13539, N13517, N12747);
nor NOR4 (N13540, N13537, N9081, N2819, N6508);
not NOT1 (N13541, N13532);
nor NOR4 (N13542, N13531, N1315, N6032, N12865);
and AND4 (N13543, N13536, N3912, N2962, N7858);
not NOT1 (N13544, N13540);
nor NOR2 (N13545, N13538, N10473);
buf BUF1 (N13546, N13529);
buf BUF1 (N13547, N13541);
xor XOR2 (N13548, N13539, N7275);
not NOT1 (N13549, N13546);
nand NAND3 (N13550, N13535, N7918, N540);
buf BUF1 (N13551, N13548);
not NOT1 (N13552, N13549);
or OR3 (N13553, N13544, N11056, N10270);
xor XOR2 (N13554, N13551, N9145);
and AND2 (N13555, N13547, N8234);
nand NAND3 (N13556, N13553, N2104, N6190);
xor XOR2 (N13557, N13550, N11181);
nor NOR4 (N13558, N13534, N3602, N5387, N9197);
buf BUF1 (N13559, N13545);
buf BUF1 (N13560, N13559);
buf BUF1 (N13561, N13542);
nand NAND3 (N13562, N13561, N5479, N7747);
or OR2 (N13563, N13557, N1531);
and AND3 (N13564, N13527, N8233, N3188);
and AND3 (N13565, N13563, N1749, N9400);
nand NAND4 (N13566, N13564, N10795, N5389, N11839);
xor XOR2 (N13567, N13554, N4408);
and AND3 (N13568, N13558, N1581, N5431);
nand NAND3 (N13569, N13556, N12739, N4958);
not NOT1 (N13570, N13569);
buf BUF1 (N13571, N13562);
nor NOR4 (N13572, N13565, N9969, N1401, N6702);
xor XOR2 (N13573, N13543, N4659);
xor XOR2 (N13574, N13573, N5025);
or OR3 (N13575, N13570, N1414, N11569);
not NOT1 (N13576, N13552);
xor XOR2 (N13577, N13574, N4273);
buf BUF1 (N13578, N13572);
xor XOR2 (N13579, N13578, N9307);
and AND2 (N13580, N13560, N507);
nand NAND4 (N13581, N13575, N3257, N2027, N5942);
not NOT1 (N13582, N13580);
not NOT1 (N13583, N13571);
buf BUF1 (N13584, N13576);
not NOT1 (N13585, N13555);
buf BUF1 (N13586, N13582);
buf BUF1 (N13587, N13586);
nand NAND4 (N13588, N13587, N3633, N11581, N11972);
or OR3 (N13589, N13568, N6658, N2113);
and AND4 (N13590, N13581, N2109, N5446, N908);
xor XOR2 (N13591, N13566, N2744);
xor XOR2 (N13592, N13589, N10709);
xor XOR2 (N13593, N13591, N721);
buf BUF1 (N13594, N13583);
nand NAND4 (N13595, N13594, N2052, N1333, N11685);
or OR3 (N13596, N13590, N2653, N5372);
nand NAND4 (N13597, N13593, N12750, N6975, N12557);
nand NAND2 (N13598, N13585, N2853);
or OR2 (N13599, N13597, N7485);
xor XOR2 (N13600, N13599, N3154);
nand NAND2 (N13601, N13592, N1308);
or OR3 (N13602, N13579, N10863, N6980);
nand NAND4 (N13603, N13567, N192, N12824, N8246);
not NOT1 (N13604, N13577);
not NOT1 (N13605, N13600);
and AND4 (N13606, N13605, N11099, N4045, N10807);
nand NAND3 (N13607, N13602, N6447, N8187);
not NOT1 (N13608, N13606);
or OR3 (N13609, N13603, N9033, N5667);
or OR2 (N13610, N13609, N2972);
not NOT1 (N13611, N13598);
and AND4 (N13612, N13607, N11674, N13425, N2022);
or OR2 (N13613, N13610, N3416);
or OR2 (N13614, N13604, N10462);
or OR3 (N13615, N13608, N299, N12938);
not NOT1 (N13616, N13584);
not NOT1 (N13617, N13588);
buf BUF1 (N13618, N13601);
not NOT1 (N13619, N13612);
buf BUF1 (N13620, N13613);
or OR4 (N13621, N13616, N912, N2085, N12174);
or OR2 (N13622, N13611, N8815);
nor NOR2 (N13623, N13620, N9633);
buf BUF1 (N13624, N13614);
nor NOR2 (N13625, N13595, N5291);
and AND2 (N13626, N13624, N6142);
xor XOR2 (N13627, N13625, N11873);
and AND2 (N13628, N13615, N4719);
buf BUF1 (N13629, N13627);
and AND4 (N13630, N13619, N6772, N1132, N1800);
and AND3 (N13631, N13630, N10172, N468);
xor XOR2 (N13632, N13617, N11218);
xor XOR2 (N13633, N13631, N13081);
nand NAND3 (N13634, N13621, N1896, N10594);
or OR3 (N13635, N13626, N8049, N7013);
nor NOR3 (N13636, N13629, N10878, N3864);
or OR4 (N13637, N13633, N12101, N7238, N6186);
buf BUF1 (N13638, N13622);
or OR4 (N13639, N13596, N8708, N10846, N2631);
nor NOR4 (N13640, N13636, N7806, N6313, N4598);
xor XOR2 (N13641, N13637, N10488);
and AND4 (N13642, N13634, N833, N9437, N7031);
and AND2 (N13643, N13628, N10694);
xor XOR2 (N13644, N13643, N5857);
xor XOR2 (N13645, N13644, N4351);
or OR4 (N13646, N13618, N9277, N5607, N7897);
not NOT1 (N13647, N13635);
not NOT1 (N13648, N13632);
and AND3 (N13649, N13646, N332, N6690);
nor NOR4 (N13650, N13638, N1720, N8829, N12131);
nor NOR2 (N13651, N13641, N8886);
xor XOR2 (N13652, N13648, N727);
xor XOR2 (N13653, N13645, N1811);
nor NOR2 (N13654, N13639, N12427);
xor XOR2 (N13655, N13642, N6261);
not NOT1 (N13656, N13653);
or OR2 (N13657, N13651, N12667);
not NOT1 (N13658, N13656);
or OR3 (N13659, N13640, N5739, N4069);
buf BUF1 (N13660, N13654);
xor XOR2 (N13661, N13647, N9739);
nand NAND4 (N13662, N13660, N504, N13247, N13418);
and AND4 (N13663, N13657, N6110, N9167, N5493);
and AND2 (N13664, N13650, N2090);
nand NAND3 (N13665, N13649, N2869, N9135);
xor XOR2 (N13666, N13661, N10672);
not NOT1 (N13667, N13655);
and AND2 (N13668, N13658, N5302);
xor XOR2 (N13669, N13659, N2102);
xor XOR2 (N13670, N13623, N1062);
or OR3 (N13671, N13665, N9448, N4556);
buf BUF1 (N13672, N13662);
nand NAND4 (N13673, N13668, N11876, N6632, N1896);
nor NOR2 (N13674, N13673, N13535);
buf BUF1 (N13675, N13652);
or OR4 (N13676, N13669, N7074, N9811, N3113);
nand NAND4 (N13677, N13671, N2116, N3024, N1977);
nand NAND4 (N13678, N13666, N7991, N2612, N4408);
nor NOR3 (N13679, N13678, N2955, N2633);
nand NAND2 (N13680, N13663, N7375);
nor NOR4 (N13681, N13664, N5894, N4520, N4433);
nand NAND4 (N13682, N13672, N722, N5714, N4516);
nor NOR3 (N13683, N13667, N6230, N12804);
xor XOR2 (N13684, N13676, N5147);
and AND2 (N13685, N13675, N2895);
nor NOR2 (N13686, N13679, N12867);
nor NOR2 (N13687, N13670, N7818);
not NOT1 (N13688, N13686);
nand NAND4 (N13689, N13687, N3099, N12887, N12642);
not NOT1 (N13690, N13674);
nand NAND3 (N13691, N13682, N13490, N12879);
buf BUF1 (N13692, N13685);
not NOT1 (N13693, N13677);
buf BUF1 (N13694, N13688);
nor NOR3 (N13695, N13681, N4174, N9335);
or OR4 (N13696, N13680, N9155, N11139, N10782);
buf BUF1 (N13697, N13683);
and AND3 (N13698, N13692, N7476, N2147);
not NOT1 (N13699, N13697);
nand NAND4 (N13700, N13684, N9924, N5374, N10721);
nand NAND3 (N13701, N13693, N10793, N4072);
buf BUF1 (N13702, N13691);
xor XOR2 (N13703, N13700, N643);
and AND4 (N13704, N13694, N7468, N4291, N3472);
xor XOR2 (N13705, N13689, N4594);
buf BUF1 (N13706, N13702);
and AND4 (N13707, N13706, N6239, N4865, N6863);
and AND2 (N13708, N13704, N12115);
nor NOR4 (N13709, N13696, N6582, N9985, N3438);
nor NOR3 (N13710, N13705, N12108, N5947);
buf BUF1 (N13711, N13701);
nand NAND2 (N13712, N13708, N3885);
buf BUF1 (N13713, N13710);
or OR4 (N13714, N13707, N10441, N8824, N2934);
buf BUF1 (N13715, N13695);
nor NOR2 (N13716, N13711, N5564);
not NOT1 (N13717, N13715);
and AND3 (N13718, N13699, N12872, N12422);
or OR2 (N13719, N13690, N2563);
not NOT1 (N13720, N13718);
nand NAND2 (N13721, N13717, N2196);
or OR3 (N13722, N13712, N5579, N11778);
nor NOR2 (N13723, N13722, N8785);
nand NAND2 (N13724, N13716, N8318);
xor XOR2 (N13725, N13703, N10471);
or OR4 (N13726, N13709, N4830, N3383, N9054);
and AND4 (N13727, N13725, N12177, N12576, N1283);
or OR3 (N13728, N13724, N3044, N7530);
buf BUF1 (N13729, N13720);
nand NAND4 (N13730, N13719, N10673, N11633, N4784);
and AND4 (N13731, N13726, N10183, N8487, N10631);
or OR2 (N13732, N13730, N9643);
and AND2 (N13733, N13723, N1351);
nand NAND4 (N13734, N13733, N3900, N13250, N1799);
nor NOR4 (N13735, N13721, N6403, N8963, N4351);
buf BUF1 (N13736, N13713);
xor XOR2 (N13737, N13728, N8566);
nand NAND4 (N13738, N13729, N4470, N2552, N7497);
nor NOR2 (N13739, N13737, N1520);
buf BUF1 (N13740, N13734);
nand NAND4 (N13741, N13731, N6853, N2407, N2915);
and AND4 (N13742, N13736, N6021, N3193, N13366);
xor XOR2 (N13743, N13742, N4738);
xor XOR2 (N13744, N13732, N13738);
buf BUF1 (N13745, N9626);
not NOT1 (N13746, N13735);
or OR4 (N13747, N13744, N642, N12664, N8433);
not NOT1 (N13748, N13743);
or OR4 (N13749, N13745, N5261, N892, N6523);
buf BUF1 (N13750, N13698);
nor NOR3 (N13751, N13748, N4125, N885);
not NOT1 (N13752, N13747);
not NOT1 (N13753, N13727);
or OR2 (N13754, N13714, N7694);
or OR3 (N13755, N13741, N9645, N12896);
buf BUF1 (N13756, N13753);
xor XOR2 (N13757, N13751, N6413);
xor XOR2 (N13758, N13749, N9678);
nor NOR4 (N13759, N13739, N1932, N7001, N493);
buf BUF1 (N13760, N13754);
and AND4 (N13761, N13758, N11562, N5278, N10237);
nand NAND2 (N13762, N13760, N5392);
and AND3 (N13763, N13757, N9344, N11697);
nand NAND3 (N13764, N13740, N10756, N4303);
nand NAND3 (N13765, N13755, N4260, N4633);
or OR3 (N13766, N13763, N4741, N13111);
buf BUF1 (N13767, N13766);
xor XOR2 (N13768, N13762, N614);
nor NOR2 (N13769, N13764, N9398);
and AND4 (N13770, N13752, N10046, N10705, N5463);
and AND4 (N13771, N13765, N5542, N7881, N10843);
nor NOR4 (N13772, N13759, N12184, N521, N723);
and AND3 (N13773, N13769, N12616, N9474);
xor XOR2 (N13774, N13767, N677);
not NOT1 (N13775, N13756);
and AND4 (N13776, N13775, N11551, N10780, N10032);
buf BUF1 (N13777, N13776);
xor XOR2 (N13778, N13774, N8170);
not NOT1 (N13779, N13778);
nand NAND2 (N13780, N13779, N11679);
not NOT1 (N13781, N13777);
not NOT1 (N13782, N13750);
and AND2 (N13783, N13761, N5457);
nand NAND2 (N13784, N13772, N3604);
nand NAND3 (N13785, N13768, N1755, N12567);
buf BUF1 (N13786, N13781);
nor NOR3 (N13787, N13770, N13683, N12902);
not NOT1 (N13788, N13782);
buf BUF1 (N13789, N13746);
or OR2 (N13790, N13773, N9086);
not NOT1 (N13791, N13788);
nor NOR4 (N13792, N13787, N12895, N2282, N4752);
and AND4 (N13793, N13792, N8190, N3146, N12687);
nor NOR2 (N13794, N13783, N2752);
and AND2 (N13795, N13785, N7442);
and AND2 (N13796, N13795, N9251);
nor NOR4 (N13797, N13784, N3784, N9378, N2185);
buf BUF1 (N13798, N13791);
or OR3 (N13799, N13793, N1910, N7726);
xor XOR2 (N13800, N13797, N675);
not NOT1 (N13801, N13771);
not NOT1 (N13802, N13800);
nor NOR2 (N13803, N13798, N8991);
and AND2 (N13804, N13803, N13243);
nand NAND3 (N13805, N13786, N13456, N1733);
nor NOR3 (N13806, N13794, N11709, N12782);
and AND3 (N13807, N13802, N4029, N1985);
and AND4 (N13808, N13801, N6189, N3788, N5767);
nand NAND3 (N13809, N13806, N6844, N142);
xor XOR2 (N13810, N13809, N1026);
buf BUF1 (N13811, N13807);
xor XOR2 (N13812, N13810, N240);
buf BUF1 (N13813, N13808);
nor NOR4 (N13814, N13804, N9700, N12498, N3341);
nand NAND4 (N13815, N13799, N755, N5099, N9902);
nand NAND4 (N13816, N13811, N8516, N7697, N8463);
nor NOR4 (N13817, N13796, N1775, N1969, N5811);
nand NAND3 (N13818, N13817, N6305, N87);
nand NAND2 (N13819, N13815, N10400);
and AND3 (N13820, N13805, N4774, N8153);
and AND4 (N13821, N13790, N10329, N7244, N6072);
nor NOR2 (N13822, N13789, N8155);
and AND2 (N13823, N13780, N4529);
or OR4 (N13824, N13813, N2255, N2666, N2718);
nor NOR3 (N13825, N13820, N5805, N3439);
nand NAND4 (N13826, N13812, N10792, N13568, N12899);
nor NOR4 (N13827, N13824, N2850, N880, N7800);
nand NAND4 (N13828, N13814, N6015, N12727, N1859);
not NOT1 (N13829, N13826);
and AND4 (N13830, N13822, N4215, N5659, N10496);
nand NAND2 (N13831, N13825, N1507);
nand NAND3 (N13832, N13830, N5729, N1101);
buf BUF1 (N13833, N13816);
or OR3 (N13834, N13821, N11609, N12685);
xor XOR2 (N13835, N13818, N12794);
or OR3 (N13836, N13833, N7402, N3073);
nand NAND2 (N13837, N13827, N13392);
buf BUF1 (N13838, N13834);
not NOT1 (N13839, N13838);
or OR2 (N13840, N13836, N3706);
and AND2 (N13841, N13832, N9059);
not NOT1 (N13842, N13837);
and AND3 (N13843, N13831, N3051, N8462);
buf BUF1 (N13844, N13842);
buf BUF1 (N13845, N13843);
or OR4 (N13846, N13845, N13151, N10775, N12534);
xor XOR2 (N13847, N13823, N9792);
and AND3 (N13848, N13828, N7202, N6562);
buf BUF1 (N13849, N13835);
and AND2 (N13850, N13829, N996);
buf BUF1 (N13851, N13849);
buf BUF1 (N13852, N13839);
nand NAND3 (N13853, N13840, N10047, N7100);
nor NOR2 (N13854, N13841, N11894);
not NOT1 (N13855, N13852);
not NOT1 (N13856, N13853);
not NOT1 (N13857, N13846);
nor NOR2 (N13858, N13855, N2084);
buf BUF1 (N13859, N13851);
not NOT1 (N13860, N13850);
nand NAND2 (N13861, N13819, N13708);
nand NAND4 (N13862, N13861, N12740, N7956, N11153);
not NOT1 (N13863, N13854);
nor NOR2 (N13864, N13857, N13318);
nand NAND4 (N13865, N13864, N7846, N3354, N400);
buf BUF1 (N13866, N13856);
nor NOR2 (N13867, N13865, N5753);
and AND2 (N13868, N13847, N1581);
xor XOR2 (N13869, N13866, N8194);
xor XOR2 (N13870, N13859, N7876);
or OR3 (N13871, N13869, N3841, N3126);
xor XOR2 (N13872, N13863, N12435);
not NOT1 (N13873, N13870);
not NOT1 (N13874, N13868);
or OR2 (N13875, N13872, N10454);
nor NOR2 (N13876, N13873, N7133);
not NOT1 (N13877, N13871);
nor NOR3 (N13878, N13877, N9130, N3497);
nand NAND3 (N13879, N13875, N5374, N6528);
or OR3 (N13880, N13867, N7290, N5957);
buf BUF1 (N13881, N13844);
nand NAND4 (N13882, N13858, N1492, N13050, N9680);
not NOT1 (N13883, N13874);
or OR2 (N13884, N13882, N6699);
not NOT1 (N13885, N13883);
buf BUF1 (N13886, N13879);
not NOT1 (N13887, N13876);
buf BUF1 (N13888, N13862);
nand NAND2 (N13889, N13884, N13716);
nand NAND3 (N13890, N13878, N2528, N4769);
and AND4 (N13891, N13886, N1992, N5698, N11340);
or OR3 (N13892, N13888, N3186, N8994);
xor XOR2 (N13893, N13890, N4323);
or OR3 (N13894, N13893, N1495, N6498);
nand NAND3 (N13895, N13881, N8577, N10465);
not NOT1 (N13896, N13887);
and AND2 (N13897, N13880, N6095);
and AND4 (N13898, N13848, N8258, N13273, N9285);
and AND4 (N13899, N13885, N11783, N5108, N9169);
xor XOR2 (N13900, N13898, N4951);
buf BUF1 (N13901, N13896);
nand NAND3 (N13902, N13900, N67, N11968);
not NOT1 (N13903, N13897);
or OR2 (N13904, N13902, N5511);
not NOT1 (N13905, N13894);
or OR4 (N13906, N13889, N2936, N11265, N5961);
xor XOR2 (N13907, N13906, N1225);
and AND3 (N13908, N13907, N998, N11503);
buf BUF1 (N13909, N13892);
xor XOR2 (N13910, N13905, N13883);
nand NAND2 (N13911, N13910, N930);
buf BUF1 (N13912, N13909);
buf BUF1 (N13913, N13903);
nand NAND3 (N13914, N13891, N9909, N13497);
and AND3 (N13915, N13908, N13007, N5655);
nor NOR4 (N13916, N13901, N12555, N1241, N3453);
xor XOR2 (N13917, N13913, N8850);
nor NOR4 (N13918, N13916, N8854, N11422, N5732);
buf BUF1 (N13919, N13911);
or OR4 (N13920, N13912, N1409, N5658, N6119);
and AND2 (N13921, N13919, N2802);
nand NAND4 (N13922, N13921, N4030, N4433, N12356);
and AND4 (N13923, N13917, N11082, N10702, N9103);
not NOT1 (N13924, N13922);
xor XOR2 (N13925, N13899, N10921);
nand NAND2 (N13926, N13860, N5723);
or OR2 (N13927, N13923, N4836);
not NOT1 (N13928, N13915);
xor XOR2 (N13929, N13928, N1251);
or OR3 (N13930, N13926, N10565, N12596);
not NOT1 (N13931, N13929);
nand NAND3 (N13932, N13930, N8817, N938);
and AND4 (N13933, N13925, N5118, N8975, N12143);
buf BUF1 (N13934, N13904);
buf BUF1 (N13935, N13933);
not NOT1 (N13936, N13918);
nand NAND3 (N13937, N13927, N11401, N8897);
xor XOR2 (N13938, N13895, N8357);
not NOT1 (N13939, N13914);
buf BUF1 (N13940, N13934);
nor NOR2 (N13941, N13940, N9374);
not NOT1 (N13942, N13937);
xor XOR2 (N13943, N13931, N4308);
nor NOR3 (N13944, N13935, N9852, N11993);
buf BUF1 (N13945, N13938);
or OR2 (N13946, N13936, N7879);
or OR2 (N13947, N13946, N12682);
buf BUF1 (N13948, N13942);
buf BUF1 (N13949, N13944);
nor NOR4 (N13950, N13945, N7868, N9273, N3037);
and AND2 (N13951, N13939, N12999);
buf BUF1 (N13952, N13932);
and AND3 (N13953, N13943, N4289, N13589);
buf BUF1 (N13954, N13953);
not NOT1 (N13955, N13941);
or OR3 (N13956, N13955, N3901, N10082);
buf BUF1 (N13957, N13924);
buf BUF1 (N13958, N13949);
buf BUF1 (N13959, N13954);
or OR3 (N13960, N13947, N6717, N1536);
not NOT1 (N13961, N13951);
buf BUF1 (N13962, N13920);
xor XOR2 (N13963, N13952, N5111);
nand NAND4 (N13964, N13959, N5578, N102, N5920);
nand NAND3 (N13965, N13950, N6794, N3715);
nand NAND4 (N13966, N13958, N2220, N11020, N8484);
nand NAND3 (N13967, N13965, N2235, N5192);
nand NAND3 (N13968, N13963, N2989, N10063);
or OR3 (N13969, N13966, N5173, N6508);
buf BUF1 (N13970, N13964);
buf BUF1 (N13971, N13962);
not NOT1 (N13972, N13960);
or OR4 (N13973, N13956, N7003, N2696, N656);
xor XOR2 (N13974, N13973, N5951);
nor NOR2 (N13975, N13957, N5323);
and AND2 (N13976, N13967, N5830);
nor NOR2 (N13977, N13969, N5907);
xor XOR2 (N13978, N13948, N13683);
buf BUF1 (N13979, N13976);
buf BUF1 (N13980, N13971);
nand NAND3 (N13981, N13972, N818, N8520);
nor NOR4 (N13982, N13977, N10879, N306, N6860);
not NOT1 (N13983, N13980);
buf BUF1 (N13984, N13983);
buf BUF1 (N13985, N13981);
nand NAND3 (N13986, N13984, N12775, N10373);
xor XOR2 (N13987, N13982, N12337);
nand NAND2 (N13988, N13979, N4639);
not NOT1 (N13989, N13975);
or OR2 (N13990, N13985, N1799);
buf BUF1 (N13991, N13974);
nand NAND4 (N13992, N13987, N5843, N8489, N6233);
buf BUF1 (N13993, N13986);
or OR2 (N13994, N13961, N3150);
nor NOR2 (N13995, N13978, N10276);
buf BUF1 (N13996, N13990);
buf BUF1 (N13997, N13996);
or OR4 (N13998, N13997, N966, N613, N13111);
and AND2 (N13999, N13968, N6565);
buf BUF1 (N14000, N13999);
xor XOR2 (N14001, N13994, N332);
or OR4 (N14002, N13970, N3671, N12213, N2758);
xor XOR2 (N14003, N13989, N12981);
not NOT1 (N14004, N14000);
not NOT1 (N14005, N13988);
or OR2 (N14006, N13992, N4885);
nor NOR3 (N14007, N13998, N12900, N2524);
nand NAND3 (N14008, N14004, N265, N10183);
nand NAND3 (N14009, N14001, N1997, N8987);
xor XOR2 (N14010, N14009, N2122);
buf BUF1 (N14011, N14010);
nor NOR2 (N14012, N13991, N10136);
or OR3 (N14013, N14003, N3072, N13910);
and AND4 (N14014, N14012, N3766, N4665, N7454);
and AND2 (N14015, N13993, N10533);
nor NOR2 (N14016, N14002, N10984);
nor NOR2 (N14017, N14006, N8658);
nand NAND3 (N14018, N13995, N4956, N9817);
or OR2 (N14019, N14017, N2891);
nand NAND2 (N14020, N14007, N12432);
not NOT1 (N14021, N14008);
buf BUF1 (N14022, N14018);
nand NAND3 (N14023, N14013, N10655, N8731);
and AND4 (N14024, N14020, N10280, N3084, N177);
or OR2 (N14025, N14015, N9633);
nand NAND4 (N14026, N14016, N2575, N13741, N12245);
buf BUF1 (N14027, N14023);
or OR2 (N14028, N14026, N7392);
xor XOR2 (N14029, N14021, N12847);
and AND3 (N14030, N14014, N9625, N1446);
nor NOR3 (N14031, N14019, N11026, N6573);
and AND3 (N14032, N14025, N7124, N7090);
nor NOR4 (N14033, N14005, N7675, N11990, N5648);
nor NOR2 (N14034, N14024, N111);
buf BUF1 (N14035, N14022);
nand NAND3 (N14036, N14030, N4272, N7889);
buf BUF1 (N14037, N14032);
or OR4 (N14038, N14035, N6133, N5085, N4395);
or OR4 (N14039, N14028, N9623, N12091, N10926);
xor XOR2 (N14040, N14034, N5153);
nor NOR4 (N14041, N14038, N8695, N3449, N4005);
and AND3 (N14042, N14041, N9430, N1499);
xor XOR2 (N14043, N14031, N8988);
nand NAND3 (N14044, N14042, N4539, N5059);
and AND3 (N14045, N14027, N10965, N1992);
xor XOR2 (N14046, N14037, N9936);
nor NOR2 (N14047, N14045, N841);
xor XOR2 (N14048, N14011, N7645);
and AND3 (N14049, N14036, N12905, N7287);
buf BUF1 (N14050, N14039);
or OR4 (N14051, N14043, N8330, N10216, N13337);
and AND3 (N14052, N14046, N7701, N5703);
xor XOR2 (N14053, N14029, N11752);
and AND3 (N14054, N14050, N11985, N3740);
or OR3 (N14055, N14048, N13687, N11494);
and AND3 (N14056, N14049, N3774, N4569);
buf BUF1 (N14057, N14052);
xor XOR2 (N14058, N14051, N12571);
xor XOR2 (N14059, N14054, N1064);
and AND2 (N14060, N14057, N9886);
buf BUF1 (N14061, N14056);
nand NAND3 (N14062, N14044, N9393, N56);
buf BUF1 (N14063, N14033);
nand NAND2 (N14064, N14060, N3229);
xor XOR2 (N14065, N14055, N2255);
and AND2 (N14066, N14063, N4171);
nor NOR2 (N14067, N14064, N8559);
or OR3 (N14068, N14047, N13036, N5240);
xor XOR2 (N14069, N14062, N11626);
not NOT1 (N14070, N14067);
nor NOR2 (N14071, N14070, N843);
buf BUF1 (N14072, N14059);
xor XOR2 (N14073, N14061, N7366);
nor NOR3 (N14074, N14065, N5424, N13935);
or OR4 (N14075, N14040, N4265, N13649, N12285);
or OR3 (N14076, N14066, N3917, N4354);
nand NAND3 (N14077, N14069, N987, N8447);
nor NOR2 (N14078, N14073, N12328);
nand NAND4 (N14079, N14058, N5566, N8276, N13375);
buf BUF1 (N14080, N14071);
or OR2 (N14081, N14068, N13909);
or OR4 (N14082, N14053, N5400, N11869, N10213);
or OR4 (N14083, N14077, N6815, N5729, N2405);
xor XOR2 (N14084, N14076, N13710);
xor XOR2 (N14085, N14074, N4054);
not NOT1 (N14086, N14080);
and AND3 (N14087, N14082, N1253, N11203);
nor NOR3 (N14088, N14083, N474, N7938);
and AND3 (N14089, N14087, N12703, N13431);
not NOT1 (N14090, N14089);
not NOT1 (N14091, N14085);
not NOT1 (N14092, N14091);
and AND2 (N14093, N14086, N1474);
xor XOR2 (N14094, N14081, N13650);
nor NOR4 (N14095, N14072, N3892, N4372, N9383);
xor XOR2 (N14096, N14079, N5498);
xor XOR2 (N14097, N14092, N3396);
buf BUF1 (N14098, N14096);
or OR2 (N14099, N14088, N2151);
xor XOR2 (N14100, N14093, N11050);
or OR4 (N14101, N14097, N10755, N10064, N3125);
xor XOR2 (N14102, N14090, N5523);
and AND4 (N14103, N14095, N3961, N2851, N10573);
nor NOR2 (N14104, N14101, N1815);
and AND2 (N14105, N14100, N1998);
and AND4 (N14106, N14075, N10885, N1360, N12706);
or OR3 (N14107, N14105, N2093, N12358);
xor XOR2 (N14108, N14078, N2678);
nor NOR3 (N14109, N14099, N4270, N5617);
not NOT1 (N14110, N14104);
and AND3 (N14111, N14094, N6208, N8937);
not NOT1 (N14112, N14110);
and AND3 (N14113, N14108, N3146, N6441);
nor NOR4 (N14114, N14109, N11094, N13925, N13869);
or OR3 (N14115, N14106, N1543, N8263);
nand NAND3 (N14116, N14112, N6002, N690);
not NOT1 (N14117, N14103);
buf BUF1 (N14118, N14116);
buf BUF1 (N14119, N14098);
nand NAND2 (N14120, N14118, N11658);
nor NOR3 (N14121, N14114, N12094, N4015);
buf BUF1 (N14122, N14102);
not NOT1 (N14123, N14121);
xor XOR2 (N14124, N14120, N5284);
buf BUF1 (N14125, N14107);
and AND3 (N14126, N14115, N9493, N5628);
nor NOR3 (N14127, N14125, N6692, N3969);
or OR4 (N14128, N14123, N5839, N801, N5471);
not NOT1 (N14129, N14084);
nand NAND4 (N14130, N14128, N5676, N4550, N7505);
buf BUF1 (N14131, N14119);
buf BUF1 (N14132, N14117);
and AND3 (N14133, N14126, N4992, N4506);
or OR4 (N14134, N14129, N9193, N13562, N10147);
or OR3 (N14135, N14124, N4182, N8114);
not NOT1 (N14136, N14134);
or OR4 (N14137, N14131, N90, N10699, N1633);
not NOT1 (N14138, N14137);
xor XOR2 (N14139, N14111, N13572);
or OR4 (N14140, N14139, N3613, N720, N9820);
buf BUF1 (N14141, N14132);
and AND4 (N14142, N14113, N9910, N12246, N7614);
buf BUF1 (N14143, N14140);
not NOT1 (N14144, N14143);
xor XOR2 (N14145, N14144, N9108);
buf BUF1 (N14146, N14127);
and AND3 (N14147, N14133, N2079, N13805);
not NOT1 (N14148, N14135);
nor NOR4 (N14149, N14147, N5283, N842, N8528);
xor XOR2 (N14150, N14149, N9801);
not NOT1 (N14151, N14141);
and AND3 (N14152, N14122, N964, N9430);
and AND2 (N14153, N14151, N11019);
or OR3 (N14154, N14136, N6694, N4075);
nor NOR2 (N14155, N14130, N3922);
or OR4 (N14156, N14142, N7078, N6188, N10622);
buf BUF1 (N14157, N14155);
buf BUF1 (N14158, N14156);
nand NAND4 (N14159, N14154, N8232, N8343, N12831);
nand NAND4 (N14160, N14148, N10684, N5797, N1731);
xor XOR2 (N14161, N14153, N11417);
and AND4 (N14162, N14145, N7941, N1108, N9495);
not NOT1 (N14163, N14158);
xor XOR2 (N14164, N14160, N11270);
buf BUF1 (N14165, N14157);
or OR2 (N14166, N14150, N11732);
nand NAND2 (N14167, N14164, N14024);
xor XOR2 (N14168, N14138, N1252);
buf BUF1 (N14169, N14163);
nor NOR2 (N14170, N14169, N11114);
buf BUF1 (N14171, N14167);
not NOT1 (N14172, N14159);
nand NAND3 (N14173, N14165, N13269, N707);
not NOT1 (N14174, N14173);
nand NAND2 (N14175, N14174, N13015);
and AND3 (N14176, N14175, N14085, N944);
not NOT1 (N14177, N14168);
not NOT1 (N14178, N14171);
and AND2 (N14179, N14146, N9433);
xor XOR2 (N14180, N14179, N9223);
nand NAND2 (N14181, N14178, N10515);
xor XOR2 (N14182, N14170, N10948);
and AND3 (N14183, N14177, N8789, N11848);
nor NOR3 (N14184, N14152, N12895, N544);
and AND3 (N14185, N14180, N9734, N12353);
nor NOR4 (N14186, N14183, N13408, N14118, N154);
and AND2 (N14187, N14184, N9199);
and AND3 (N14188, N14176, N3998, N4574);
not NOT1 (N14189, N14182);
and AND2 (N14190, N14162, N3554);
nor NOR3 (N14191, N14181, N11947, N12092);
nand NAND3 (N14192, N14187, N2118, N808);
xor XOR2 (N14193, N14189, N6404);
not NOT1 (N14194, N14172);
not NOT1 (N14195, N14194);
nor NOR2 (N14196, N14192, N12166);
and AND4 (N14197, N14190, N10223, N12346, N13660);
or OR3 (N14198, N14186, N6397, N2990);
buf BUF1 (N14199, N14166);
buf BUF1 (N14200, N14198);
or OR3 (N14201, N14193, N11137, N8315);
buf BUF1 (N14202, N14191);
not NOT1 (N14203, N14161);
buf BUF1 (N14204, N14188);
xor XOR2 (N14205, N14199, N3162);
buf BUF1 (N14206, N14204);
and AND3 (N14207, N14200, N11775, N10256);
and AND2 (N14208, N14205, N9332);
or OR4 (N14209, N14197, N9519, N11460, N2693);
xor XOR2 (N14210, N14185, N8614);
nor NOR4 (N14211, N14196, N2567, N11284, N1137);
xor XOR2 (N14212, N14211, N4038);
nand NAND4 (N14213, N14201, N12752, N1844, N11326);
or OR2 (N14214, N14212, N8637);
nor NOR3 (N14215, N14207, N8099, N11064);
not NOT1 (N14216, N14210);
or OR2 (N14217, N14208, N12783);
or OR3 (N14218, N14195, N3219, N1570);
not NOT1 (N14219, N14213);
nand NAND3 (N14220, N14215, N12870, N8804);
buf BUF1 (N14221, N14218);
buf BUF1 (N14222, N14217);
and AND4 (N14223, N14222, N5277, N5797, N5734);
nand NAND2 (N14224, N14220, N4568);
not NOT1 (N14225, N14223);
xor XOR2 (N14226, N14202, N72);
xor XOR2 (N14227, N14209, N9418);
not NOT1 (N14228, N14206);
not NOT1 (N14229, N14221);
xor XOR2 (N14230, N14228, N3206);
buf BUF1 (N14231, N14226);
xor XOR2 (N14232, N14216, N2802);
nand NAND3 (N14233, N14232, N2935, N599);
and AND3 (N14234, N14233, N12508, N8766);
nand NAND4 (N14235, N14203, N6127, N5980, N662);
and AND2 (N14236, N14229, N2134);
not NOT1 (N14237, N14236);
not NOT1 (N14238, N14214);
not NOT1 (N14239, N14235);
and AND2 (N14240, N14231, N7079);
xor XOR2 (N14241, N14238, N8318);
or OR4 (N14242, N14224, N2771, N1537, N11925);
nor NOR4 (N14243, N14241, N9650, N3418, N416);
nand NAND2 (N14244, N14243, N13361);
nand NAND4 (N14245, N14244, N10666, N7569, N397);
xor XOR2 (N14246, N14234, N6379);
nand NAND3 (N14247, N14225, N7398, N4201);
nor NOR2 (N14248, N14219, N11919);
not NOT1 (N14249, N14247);
not NOT1 (N14250, N14245);
or OR2 (N14251, N14239, N7320);
nor NOR2 (N14252, N14230, N14069);
nor NOR3 (N14253, N14251, N85, N10293);
xor XOR2 (N14254, N14237, N13507);
buf BUF1 (N14255, N14240);
or OR2 (N14256, N14248, N10061);
nor NOR3 (N14257, N14250, N12430, N7824);
and AND2 (N14258, N14252, N8253);
buf BUF1 (N14259, N14258);
and AND3 (N14260, N14255, N7711, N11283);
nand NAND3 (N14261, N14260, N13628, N4381);
xor XOR2 (N14262, N14259, N12789);
not NOT1 (N14263, N14257);
buf BUF1 (N14264, N14262);
not NOT1 (N14265, N14246);
buf BUF1 (N14266, N14227);
or OR4 (N14267, N14253, N5754, N10417, N1713);
buf BUF1 (N14268, N14242);
not NOT1 (N14269, N14249);
and AND4 (N14270, N14266, N9211, N12718, N11712);
not NOT1 (N14271, N14264);
nand NAND4 (N14272, N14261, N12011, N3627, N6199);
or OR4 (N14273, N14263, N6847, N9918, N8230);
xor XOR2 (N14274, N14270, N4664);
not NOT1 (N14275, N14273);
or OR3 (N14276, N14256, N7982, N11671);
or OR4 (N14277, N14268, N4154, N6798, N6229);
or OR3 (N14278, N14269, N7929, N4117);
nand NAND2 (N14279, N14278, N3857);
not NOT1 (N14280, N14265);
and AND3 (N14281, N14272, N1903, N5498);
buf BUF1 (N14282, N14277);
nand NAND3 (N14283, N14274, N7289, N6919);
xor XOR2 (N14284, N14283, N9677);
not NOT1 (N14285, N14282);
and AND2 (N14286, N14254, N2137);
or OR3 (N14287, N14281, N6930, N4424);
buf BUF1 (N14288, N14271);
or OR2 (N14289, N14279, N13093);
and AND3 (N14290, N14288, N5119, N1982);
or OR2 (N14291, N14284, N12226);
xor XOR2 (N14292, N14289, N12529);
nor NOR4 (N14293, N14276, N10787, N13137, N1382);
xor XOR2 (N14294, N14287, N12816);
buf BUF1 (N14295, N14294);
or OR3 (N14296, N14275, N6849, N200);
and AND2 (N14297, N14296, N13903);
not NOT1 (N14298, N14295);
xor XOR2 (N14299, N14291, N5976);
not NOT1 (N14300, N14299);
and AND4 (N14301, N14285, N2037, N13445, N9178);
nor NOR2 (N14302, N14301, N1797);
buf BUF1 (N14303, N14300);
xor XOR2 (N14304, N14267, N483);
buf BUF1 (N14305, N14297);
or OR2 (N14306, N14302, N7737);
xor XOR2 (N14307, N14304, N4879);
nand NAND3 (N14308, N14290, N13575, N12343);
buf BUF1 (N14309, N14303);
and AND4 (N14310, N14293, N538, N5439, N1321);
not NOT1 (N14311, N14292);
nor NOR2 (N14312, N14309, N3662);
or OR2 (N14313, N14312, N11555);
and AND2 (N14314, N14307, N8675);
and AND3 (N14315, N14308, N7796, N7363);
nand NAND3 (N14316, N14286, N1643, N1672);
buf BUF1 (N14317, N14298);
and AND2 (N14318, N14313, N12346);
not NOT1 (N14319, N14311);
not NOT1 (N14320, N14310);
xor XOR2 (N14321, N14316, N11473);
xor XOR2 (N14322, N14314, N9667);
buf BUF1 (N14323, N14322);
and AND4 (N14324, N14305, N6572, N10630, N2943);
or OR4 (N14325, N14280, N12312, N5106, N4802);
and AND2 (N14326, N14321, N6865);
buf BUF1 (N14327, N14324);
xor XOR2 (N14328, N14306, N12102);
and AND4 (N14329, N14319, N2680, N2500, N7020);
not NOT1 (N14330, N14329);
nor NOR4 (N14331, N14320, N7454, N2534, N9831);
not NOT1 (N14332, N14318);
xor XOR2 (N14333, N14328, N5993);
nand NAND4 (N14334, N14333, N8310, N6604, N4292);
nor NOR3 (N14335, N14334, N3791, N6073);
not NOT1 (N14336, N14315);
nor NOR4 (N14337, N14327, N2528, N11912, N9077);
xor XOR2 (N14338, N14326, N11871);
nor NOR4 (N14339, N14331, N2016, N10570, N2025);
buf BUF1 (N14340, N14332);
xor XOR2 (N14341, N14323, N8924);
not NOT1 (N14342, N14330);
nor NOR2 (N14343, N14341, N1909);
nand NAND2 (N14344, N14338, N12574);
and AND3 (N14345, N14335, N4608, N6762);
nand NAND3 (N14346, N14339, N13255, N4408);
and AND2 (N14347, N14344, N8066);
or OR3 (N14348, N14343, N1898, N12075);
and AND3 (N14349, N14325, N4072, N13734);
buf BUF1 (N14350, N14345);
and AND3 (N14351, N14346, N1386, N8595);
buf BUF1 (N14352, N14317);
xor XOR2 (N14353, N14348, N11038);
nor NOR2 (N14354, N14347, N5781);
not NOT1 (N14355, N14340);
xor XOR2 (N14356, N14337, N4586);
or OR3 (N14357, N14356, N13158, N2432);
not NOT1 (N14358, N14349);
xor XOR2 (N14359, N14336, N3790);
nor NOR2 (N14360, N14352, N11700);
and AND4 (N14361, N14342, N10263, N12223, N6353);
xor XOR2 (N14362, N14359, N1280);
nand NAND4 (N14363, N14357, N2936, N10559, N6000);
not NOT1 (N14364, N14361);
buf BUF1 (N14365, N14350);
and AND4 (N14366, N14364, N2985, N9269, N2781);
nor NOR4 (N14367, N14366, N4870, N3797, N5586);
nor NOR4 (N14368, N14358, N11464, N1520, N8098);
or OR4 (N14369, N14355, N6993, N7511, N11030);
not NOT1 (N14370, N14353);
or OR4 (N14371, N14365, N2662, N5983, N8736);
nand NAND2 (N14372, N14367, N10784);
nor NOR4 (N14373, N14360, N6193, N7293, N8105);
xor XOR2 (N14374, N14371, N7080);
buf BUF1 (N14375, N14374);
nor NOR3 (N14376, N14372, N13168, N208);
or OR4 (N14377, N14368, N148, N7672, N2597);
nand NAND4 (N14378, N14377, N2412, N8746, N13678);
nor NOR3 (N14379, N14351, N11590, N11267);
not NOT1 (N14380, N14370);
not NOT1 (N14381, N14376);
nand NAND3 (N14382, N14363, N4832, N10471);
nand NAND2 (N14383, N14380, N3877);
xor XOR2 (N14384, N14378, N10262);
xor XOR2 (N14385, N14382, N2926);
nor NOR2 (N14386, N14369, N8797);
nor NOR2 (N14387, N14354, N3716);
and AND3 (N14388, N14373, N1462, N3655);
buf BUF1 (N14389, N14383);
nand NAND3 (N14390, N14389, N5328, N1687);
nand NAND3 (N14391, N14375, N7594, N3228);
and AND2 (N14392, N14390, N7378);
and AND4 (N14393, N14386, N5166, N6826, N4864);
not NOT1 (N14394, N14387);
xor XOR2 (N14395, N14392, N7613);
xor XOR2 (N14396, N14381, N4418);
nor NOR3 (N14397, N14362, N13330, N1704);
not NOT1 (N14398, N14388);
xor XOR2 (N14399, N14391, N672);
buf BUF1 (N14400, N14395);
nor NOR4 (N14401, N14399, N13549, N3415, N6966);
and AND4 (N14402, N14400, N6381, N8008, N1664);
xor XOR2 (N14403, N14379, N2181);
nor NOR4 (N14404, N14385, N8220, N123, N13649);
not NOT1 (N14405, N14393);
or OR2 (N14406, N14404, N10501);
and AND4 (N14407, N14396, N3237, N8179, N12803);
or OR3 (N14408, N14397, N5667, N362);
nor NOR3 (N14409, N14384, N12617, N13626);
not NOT1 (N14410, N14403);
or OR4 (N14411, N14410, N7070, N6561, N5919);
or OR3 (N14412, N14408, N2924, N3091);
nor NOR3 (N14413, N14409, N4391, N9096);
and AND3 (N14414, N14411, N7345, N3292);
nand NAND3 (N14415, N14406, N5890, N13394);
buf BUF1 (N14416, N14413);
nand NAND3 (N14417, N14414, N14391, N13246);
not NOT1 (N14418, N14407);
nor NOR4 (N14419, N14394, N4254, N10702, N9803);
buf BUF1 (N14420, N14415);
nor NOR4 (N14421, N14412, N10339, N14107, N866);
nand NAND2 (N14422, N14418, N12084);
xor XOR2 (N14423, N14401, N11439);
nand NAND4 (N14424, N14422, N13695, N6890, N10310);
and AND2 (N14425, N14402, N13049);
not NOT1 (N14426, N14421);
xor XOR2 (N14427, N14398, N10930);
buf BUF1 (N14428, N14416);
buf BUF1 (N14429, N14420);
xor XOR2 (N14430, N14405, N5144);
xor XOR2 (N14431, N14428, N12063);
or OR4 (N14432, N14423, N11989, N14301, N7282);
buf BUF1 (N14433, N14430);
nand NAND4 (N14434, N14427, N12743, N12871, N2230);
nand NAND3 (N14435, N14431, N7329, N13872);
not NOT1 (N14436, N14426);
nand NAND3 (N14437, N14424, N11820, N4477);
nand NAND4 (N14438, N14437, N4919, N8161, N3516);
nand NAND3 (N14439, N14432, N4967, N2500);
and AND4 (N14440, N14436, N11041, N5002, N3328);
buf BUF1 (N14441, N14429);
xor XOR2 (N14442, N14438, N184);
nand NAND4 (N14443, N14442, N4375, N1853, N1351);
nor NOR3 (N14444, N14440, N2433, N10656);
nand NAND4 (N14445, N14443, N11266, N5078, N9518);
or OR2 (N14446, N14435, N5842);
nand NAND4 (N14447, N14417, N5250, N2677, N5911);
not NOT1 (N14448, N14444);
buf BUF1 (N14449, N14433);
nor NOR2 (N14450, N14448, N7448);
buf BUF1 (N14451, N14450);
not NOT1 (N14452, N14447);
buf BUF1 (N14453, N14452);
not NOT1 (N14454, N14441);
and AND3 (N14455, N14439, N2307, N1067);
xor XOR2 (N14456, N14445, N3456);
or OR4 (N14457, N14425, N8461, N9644, N9232);
xor XOR2 (N14458, N14457, N797);
or OR4 (N14459, N14453, N4397, N13079, N5888);
and AND3 (N14460, N14459, N8975, N13005);
and AND3 (N14461, N14446, N6760, N10101);
nor NOR3 (N14462, N14449, N5593, N9891);
or OR3 (N14463, N14454, N6958, N5847);
and AND4 (N14464, N14462, N11400, N7647, N8023);
buf BUF1 (N14465, N14434);
and AND4 (N14466, N14461, N10871, N3504, N8733);
buf BUF1 (N14467, N14419);
nand NAND2 (N14468, N14458, N13803);
not NOT1 (N14469, N14463);
nand NAND2 (N14470, N14460, N14433);
not NOT1 (N14471, N14470);
xor XOR2 (N14472, N14455, N9054);
not NOT1 (N14473, N14469);
nand NAND4 (N14474, N14466, N12030, N6232, N5800);
buf BUF1 (N14475, N14473);
buf BUF1 (N14476, N14465);
nor NOR2 (N14477, N14474, N7397);
not NOT1 (N14478, N14467);
nand NAND3 (N14479, N14468, N6064, N8871);
nor NOR4 (N14480, N14479, N13045, N12687, N7338);
nand NAND4 (N14481, N14477, N12254, N5113, N2951);
and AND2 (N14482, N14464, N13115);
or OR2 (N14483, N14471, N993);
or OR2 (N14484, N14478, N6881);
and AND4 (N14485, N14456, N10139, N5922, N11455);
not NOT1 (N14486, N14451);
buf BUF1 (N14487, N14475);
buf BUF1 (N14488, N14486);
buf BUF1 (N14489, N14484);
or OR4 (N14490, N14476, N332, N12011, N3607);
xor XOR2 (N14491, N14488, N6079);
or OR4 (N14492, N14483, N7905, N9250, N7424);
not NOT1 (N14493, N14485);
buf BUF1 (N14494, N14493);
and AND2 (N14495, N14482, N7559);
or OR3 (N14496, N14490, N9407, N468);
not NOT1 (N14497, N14495);
buf BUF1 (N14498, N14480);
xor XOR2 (N14499, N14494, N3861);
nor NOR3 (N14500, N14491, N13943, N8781);
nor NOR4 (N14501, N14472, N8920, N4853, N13540);
nand NAND3 (N14502, N14492, N13791, N1797);
buf BUF1 (N14503, N14497);
or OR3 (N14504, N14503, N12490, N3789);
and AND3 (N14505, N14499, N8620, N1422);
nor NOR2 (N14506, N14505, N11140);
nor NOR4 (N14507, N14506, N3062, N8124, N8032);
buf BUF1 (N14508, N14487);
buf BUF1 (N14509, N14481);
buf BUF1 (N14510, N14502);
not NOT1 (N14511, N14496);
buf BUF1 (N14512, N14511);
buf BUF1 (N14513, N14508);
nand NAND2 (N14514, N14498, N5300);
nor NOR4 (N14515, N14512, N903, N1240, N8459);
and AND3 (N14516, N14507, N1780, N8475);
buf BUF1 (N14517, N14513);
buf BUF1 (N14518, N14516);
not NOT1 (N14519, N14517);
xor XOR2 (N14520, N14518, N4960);
not NOT1 (N14521, N14510);
nor NOR4 (N14522, N14515, N1970, N235, N7670);
nand NAND4 (N14523, N14509, N4009, N10568, N7872);
not NOT1 (N14524, N14519);
not NOT1 (N14525, N14524);
or OR4 (N14526, N14500, N587, N1994, N1934);
xor XOR2 (N14527, N14525, N14170);
not NOT1 (N14528, N14527);
nor NOR4 (N14529, N14520, N12096, N10141, N1159);
xor XOR2 (N14530, N14523, N11954);
nor NOR2 (N14531, N14522, N10048);
buf BUF1 (N14532, N14530);
not NOT1 (N14533, N14529);
nor NOR4 (N14534, N14514, N1537, N8178, N6301);
nand NAND3 (N14535, N14533, N12048, N6320);
or OR2 (N14536, N14504, N11289);
xor XOR2 (N14537, N14501, N2611);
or OR4 (N14538, N14521, N6041, N5317, N2743);
or OR3 (N14539, N14489, N8839, N7380);
xor XOR2 (N14540, N14537, N13189);
xor XOR2 (N14541, N14534, N2452);
xor XOR2 (N14542, N14535, N7893);
nand NAND2 (N14543, N14532, N12922);
and AND2 (N14544, N14526, N12651);
and AND3 (N14545, N14536, N4292, N11182);
or OR4 (N14546, N14540, N814, N11848, N3895);
xor XOR2 (N14547, N14539, N10076);
xor XOR2 (N14548, N14538, N6619);
nand NAND4 (N14549, N14542, N7052, N13474, N6810);
not NOT1 (N14550, N14548);
not NOT1 (N14551, N14549);
nand NAND3 (N14552, N14546, N8009, N8312);
or OR2 (N14553, N14531, N1076);
and AND2 (N14554, N14541, N4073);
xor XOR2 (N14555, N14545, N3153);
not NOT1 (N14556, N14543);
nand NAND2 (N14557, N14555, N7267);
xor XOR2 (N14558, N14528, N8707);
xor XOR2 (N14559, N14554, N4961);
buf BUF1 (N14560, N14558);
xor XOR2 (N14561, N14560, N5000);
buf BUF1 (N14562, N14547);
nand NAND3 (N14563, N14561, N14000, N14400);
buf BUF1 (N14564, N14562);
buf BUF1 (N14565, N14556);
nand NAND3 (N14566, N14563, N5978, N2684);
or OR3 (N14567, N14565, N10751, N11855);
or OR2 (N14568, N14567, N2665);
nand NAND2 (N14569, N14550, N3866);
and AND4 (N14570, N14557, N10940, N8305, N11234);
and AND3 (N14571, N14559, N10130, N6440);
nor NOR3 (N14572, N14566, N5808, N454);
nand NAND3 (N14573, N14570, N8367, N11165);
and AND4 (N14574, N14551, N3044, N804, N13372);
nor NOR3 (N14575, N14571, N10841, N691);
nor NOR2 (N14576, N14574, N410);
and AND2 (N14577, N14553, N5240);
and AND2 (N14578, N14569, N1433);
or OR2 (N14579, N14573, N13387);
or OR4 (N14580, N14544, N7441, N2537, N2449);
nor NOR2 (N14581, N14579, N13743);
nor NOR4 (N14582, N14575, N14274, N10719, N2166);
buf BUF1 (N14583, N14577);
nand NAND2 (N14584, N14552, N5343);
or OR2 (N14585, N14582, N5560);
nand NAND2 (N14586, N14581, N6462);
nand NAND2 (N14587, N14564, N10086);
buf BUF1 (N14588, N14583);
and AND4 (N14589, N14587, N3212, N7185, N13952);
not NOT1 (N14590, N14568);
buf BUF1 (N14591, N14572);
nor NOR3 (N14592, N14578, N3540, N7681);
nor NOR2 (N14593, N14585, N9508);
buf BUF1 (N14594, N14589);
and AND2 (N14595, N14586, N13020);
nor NOR3 (N14596, N14594, N1304, N4247);
xor XOR2 (N14597, N14592, N6413);
buf BUF1 (N14598, N14591);
nor NOR2 (N14599, N14590, N2895);
or OR4 (N14600, N14593, N4201, N4546, N1462);
and AND3 (N14601, N14580, N11823, N6056);
nor NOR3 (N14602, N14588, N434, N6118);
xor XOR2 (N14603, N14595, N4098);
not NOT1 (N14604, N14596);
xor XOR2 (N14605, N14601, N5076);
and AND2 (N14606, N14603, N12976);
not NOT1 (N14607, N14598);
or OR3 (N14608, N14604, N11230, N10276);
or OR2 (N14609, N14607, N12475);
xor XOR2 (N14610, N14584, N338);
and AND4 (N14611, N14605, N14168, N13010, N755);
and AND4 (N14612, N14576, N14221, N13485, N2296);
nand NAND2 (N14613, N14597, N171);
not NOT1 (N14614, N14600);
or OR3 (N14615, N14599, N6035, N14611);
and AND3 (N14616, N7886, N3145, N4246);
nand NAND4 (N14617, N14613, N12185, N3579, N12836);
and AND2 (N14618, N14616, N253);
nand NAND4 (N14619, N14614, N4010, N2444, N9740);
and AND3 (N14620, N14606, N14454, N2632);
not NOT1 (N14621, N14617);
nand NAND4 (N14622, N14619, N8613, N13257, N7939);
not NOT1 (N14623, N14620);
nand NAND4 (N14624, N14615, N2407, N4123, N8434);
and AND3 (N14625, N14618, N13403, N1165);
or OR2 (N14626, N14612, N12093);
buf BUF1 (N14627, N14626);
buf BUF1 (N14628, N14625);
buf BUF1 (N14629, N14602);
or OR4 (N14630, N14608, N8157, N1697, N12109);
or OR4 (N14631, N14609, N6665, N4386, N4175);
not NOT1 (N14632, N14610);
or OR4 (N14633, N14624, N638, N1482, N5236);
not NOT1 (N14634, N14623);
nand NAND2 (N14635, N14631, N9975);
nor NOR4 (N14636, N14627, N12603, N11179, N11786);
not NOT1 (N14637, N14636);
or OR3 (N14638, N14629, N13349, N5315);
buf BUF1 (N14639, N14633);
not NOT1 (N14640, N14622);
nor NOR2 (N14641, N14628, N11694);
xor XOR2 (N14642, N14641, N11823);
and AND4 (N14643, N14621, N10281, N195, N1213);
nand NAND2 (N14644, N14643, N8082);
nand NAND4 (N14645, N14637, N2681, N8193, N7664);
buf BUF1 (N14646, N14638);
nor NOR4 (N14647, N14645, N11484, N8293, N9993);
nor NOR3 (N14648, N14647, N14042, N11208);
nor NOR4 (N14649, N14632, N8924, N6510, N8763);
buf BUF1 (N14650, N14639);
and AND2 (N14651, N14640, N996);
xor XOR2 (N14652, N14646, N728);
nand NAND2 (N14653, N14642, N12241);
and AND4 (N14654, N14644, N5607, N4178, N10340);
and AND2 (N14655, N14650, N14572);
xor XOR2 (N14656, N14649, N10682);
nand NAND3 (N14657, N14655, N809, N2815);
xor XOR2 (N14658, N14635, N468);
nand NAND2 (N14659, N14654, N6556);
not NOT1 (N14660, N14648);
and AND2 (N14661, N14659, N8683);
and AND2 (N14662, N14657, N7499);
not NOT1 (N14663, N14630);
not NOT1 (N14664, N14634);
nor NOR3 (N14665, N14658, N9478, N6731);
buf BUF1 (N14666, N14663);
nand NAND3 (N14667, N14653, N13738, N12231);
not NOT1 (N14668, N14665);
or OR4 (N14669, N14664, N5107, N11870, N10830);
buf BUF1 (N14670, N14661);
buf BUF1 (N14671, N14669);
not NOT1 (N14672, N14656);
nor NOR3 (N14673, N14662, N13983, N13623);
and AND2 (N14674, N14673, N5118);
and AND4 (N14675, N14651, N10633, N4098, N3381);
and AND3 (N14676, N14670, N12013, N7684);
or OR2 (N14677, N14671, N14350);
nor NOR2 (N14678, N14660, N9918);
or OR3 (N14679, N14666, N7031, N9009);
and AND4 (N14680, N14678, N9485, N4282, N10841);
nand NAND2 (N14681, N14652, N14402);
not NOT1 (N14682, N14679);
not NOT1 (N14683, N14668);
nand NAND4 (N14684, N14681, N11682, N618, N6512);
not NOT1 (N14685, N14680);
or OR4 (N14686, N14667, N573, N10324, N1496);
xor XOR2 (N14687, N14684, N9026);
nor NOR2 (N14688, N14682, N14192);
or OR3 (N14689, N14674, N10535, N1959);
and AND2 (N14690, N14675, N7629);
or OR3 (N14691, N14688, N8953, N8605);
xor XOR2 (N14692, N14683, N1382);
xor XOR2 (N14693, N14691, N12532);
nand NAND2 (N14694, N14686, N4429);
buf BUF1 (N14695, N14690);
nand NAND2 (N14696, N14694, N10504);
nor NOR2 (N14697, N14676, N13431);
or OR2 (N14698, N14672, N7532);
not NOT1 (N14699, N14697);
not NOT1 (N14700, N14696);
not NOT1 (N14701, N14699);
nand NAND3 (N14702, N14698, N10043, N3072);
or OR4 (N14703, N14685, N8429, N13672, N12819);
nor NOR3 (N14704, N14689, N6097, N6117);
or OR3 (N14705, N14687, N9945, N1332);
buf BUF1 (N14706, N14704);
buf BUF1 (N14707, N14693);
not NOT1 (N14708, N14692);
xor XOR2 (N14709, N14707, N8090);
or OR4 (N14710, N14700, N1650, N5593, N12705);
or OR4 (N14711, N14710, N3441, N9250, N12313);
not NOT1 (N14712, N14677);
nor NOR4 (N14713, N14702, N38, N5979, N6841);
and AND2 (N14714, N14711, N4243);
nor NOR4 (N14715, N14712, N8138, N7947, N2267);
buf BUF1 (N14716, N14708);
nor NOR3 (N14717, N14713, N10749, N12118);
buf BUF1 (N14718, N14709);
nand NAND4 (N14719, N14715, N8163, N7109, N12826);
or OR3 (N14720, N14695, N8051, N7811);
buf BUF1 (N14721, N14719);
xor XOR2 (N14722, N14721, N4964);
nand NAND4 (N14723, N14703, N11392, N14627, N3205);
xor XOR2 (N14724, N14717, N9590);
or OR3 (N14725, N14723, N2599, N9144);
nor NOR2 (N14726, N14705, N8141);
or OR3 (N14727, N14716, N11063, N14644);
not NOT1 (N14728, N14725);
not NOT1 (N14729, N14720);
xor XOR2 (N14730, N14728, N25);
buf BUF1 (N14731, N14701);
not NOT1 (N14732, N14718);
or OR4 (N14733, N14706, N11919, N8221, N2735);
not NOT1 (N14734, N14732);
and AND3 (N14735, N14727, N8913, N12478);
and AND3 (N14736, N14730, N11868, N13714);
nand NAND4 (N14737, N14722, N3491, N3061, N6923);
or OR2 (N14738, N14724, N8526);
xor XOR2 (N14739, N14735, N4643);
xor XOR2 (N14740, N14726, N13331);
and AND3 (N14741, N14739, N11726, N5170);
nand NAND2 (N14742, N14737, N13755);
and AND2 (N14743, N14714, N14492);
buf BUF1 (N14744, N14740);
nor NOR4 (N14745, N14744, N5459, N9172, N14048);
xor XOR2 (N14746, N14741, N5258);
nand NAND3 (N14747, N14734, N9416, N10090);
nor NOR2 (N14748, N14733, N5082);
buf BUF1 (N14749, N14745);
nand NAND3 (N14750, N14729, N10836, N14723);
nor NOR4 (N14751, N14743, N2182, N6784, N12636);
buf BUF1 (N14752, N14749);
and AND2 (N14753, N14751, N12280);
xor XOR2 (N14754, N14738, N8422);
xor XOR2 (N14755, N14747, N9498);
or OR4 (N14756, N14753, N1575, N2250, N5570);
or OR3 (N14757, N14756, N9821, N11357);
buf BUF1 (N14758, N14742);
nand NAND2 (N14759, N14748, N3972);
nand NAND4 (N14760, N14750, N14688, N9387, N8371);
nand NAND3 (N14761, N14754, N12301, N1289);
not NOT1 (N14762, N14755);
or OR3 (N14763, N14731, N11949, N10278);
nand NAND4 (N14764, N14758, N2447, N10454, N3024);
nor NOR2 (N14765, N14752, N4443);
not NOT1 (N14766, N14762);
nor NOR4 (N14767, N14766, N12724, N11936, N3801);
buf BUF1 (N14768, N14761);
or OR3 (N14769, N14764, N2098, N9285);
and AND2 (N14770, N14757, N13742);
buf BUF1 (N14771, N14769);
xor XOR2 (N14772, N14767, N3382);
xor XOR2 (N14773, N14770, N6297);
and AND3 (N14774, N14765, N10418, N8864);
buf BUF1 (N14775, N14774);
buf BUF1 (N14776, N14771);
xor XOR2 (N14777, N14768, N11180);
buf BUF1 (N14778, N14776);
and AND2 (N14779, N14759, N9219);
buf BUF1 (N14780, N14772);
xor XOR2 (N14781, N14746, N6626);
nor NOR4 (N14782, N14780, N1032, N4807, N10368);
nand NAND2 (N14783, N14760, N7379);
buf BUF1 (N14784, N14778);
buf BUF1 (N14785, N14775);
nor NOR4 (N14786, N14784, N1284, N12213, N13452);
xor XOR2 (N14787, N14785, N13125);
nor NOR3 (N14788, N14783, N11813, N7934);
or OR4 (N14789, N14782, N7420, N2679, N286);
nand NAND3 (N14790, N14773, N2587, N10494);
or OR2 (N14791, N14777, N11174);
nand NAND3 (N14792, N14788, N12055, N12383);
or OR3 (N14793, N14787, N7570, N10262);
and AND2 (N14794, N14790, N9640);
nor NOR2 (N14795, N14789, N9593);
nor NOR3 (N14796, N14791, N12167, N8605);
xor XOR2 (N14797, N14795, N13989);
not NOT1 (N14798, N14796);
nand NAND4 (N14799, N14779, N12958, N6089, N13099);
xor XOR2 (N14800, N14781, N12551);
nand NAND3 (N14801, N14799, N10386, N9947);
nor NOR2 (N14802, N14763, N6975);
xor XOR2 (N14803, N14736, N13504);
nor NOR2 (N14804, N14786, N10521);
and AND3 (N14805, N14794, N10736, N2953);
and AND3 (N14806, N14802, N11231, N6190);
or OR2 (N14807, N14800, N4170);
or OR4 (N14808, N14804, N3431, N10013, N14749);
or OR2 (N14809, N14803, N7220);
and AND4 (N14810, N14806, N8516, N3257, N10603);
and AND4 (N14811, N14807, N852, N677, N14154);
or OR3 (N14812, N14810, N5328, N10948);
not NOT1 (N14813, N14811);
buf BUF1 (N14814, N14792);
and AND2 (N14815, N14809, N10064);
nor NOR4 (N14816, N14808, N1569, N894, N226);
not NOT1 (N14817, N14812);
nand NAND3 (N14818, N14797, N6699, N12543);
buf BUF1 (N14819, N14818);
nor NOR4 (N14820, N14801, N1727, N712, N11693);
buf BUF1 (N14821, N14819);
not NOT1 (N14822, N14793);
nand NAND4 (N14823, N14822, N4386, N13295, N13295);
and AND3 (N14824, N14813, N8613, N3537);
nand NAND3 (N14825, N14820, N1168, N5140);
xor XOR2 (N14826, N14821, N2237);
nand NAND2 (N14827, N14816, N8479);
not NOT1 (N14828, N14824);
xor XOR2 (N14829, N14815, N5319);
nor NOR4 (N14830, N14823, N14208, N11513, N9808);
or OR3 (N14831, N14805, N7133, N1457);
or OR3 (N14832, N14826, N10691, N11472);
or OR4 (N14833, N14825, N7914, N2352, N3585);
xor XOR2 (N14834, N14832, N918);
buf BUF1 (N14835, N14830);
buf BUF1 (N14836, N14833);
buf BUF1 (N14837, N14817);
and AND3 (N14838, N14814, N1492, N2761);
or OR3 (N14839, N14829, N10386, N123);
not NOT1 (N14840, N14828);
and AND3 (N14841, N14835, N12492, N10886);
not NOT1 (N14842, N14798);
or OR4 (N14843, N14837, N12470, N6899, N2176);
buf BUF1 (N14844, N14827);
xor XOR2 (N14845, N14834, N14789);
or OR2 (N14846, N14840, N5528);
and AND3 (N14847, N14845, N7368, N11564);
or OR4 (N14848, N14831, N613, N9224, N10626);
nand NAND2 (N14849, N14843, N12160);
or OR4 (N14850, N14847, N4800, N10605, N2616);
nor NOR3 (N14851, N14836, N12434, N8149);
nor NOR3 (N14852, N14839, N11643, N6894);
nand NAND4 (N14853, N14848, N10613, N9549, N1171);
xor XOR2 (N14854, N14838, N13907);
nand NAND4 (N14855, N14842, N7638, N9337, N10235);
nand NAND2 (N14856, N14853, N9169);
and AND2 (N14857, N14855, N4802);
not NOT1 (N14858, N14856);
or OR2 (N14859, N14841, N10585);
buf BUF1 (N14860, N14859);
not NOT1 (N14861, N14857);
or OR2 (N14862, N14860, N10043);
nor NOR2 (N14863, N14852, N4582);
nor NOR4 (N14864, N14863, N6830, N10824, N10027);
and AND3 (N14865, N14846, N6999, N2112);
and AND3 (N14866, N14844, N3389, N968);
nor NOR4 (N14867, N14864, N7959, N4076, N9695);
buf BUF1 (N14868, N14850);
xor XOR2 (N14869, N14866, N1377);
nor NOR2 (N14870, N14854, N476);
nand NAND2 (N14871, N14849, N7299);
not NOT1 (N14872, N14867);
xor XOR2 (N14873, N14861, N8389);
xor XOR2 (N14874, N14858, N13571);
or OR3 (N14875, N14871, N11595, N12108);
nor NOR4 (N14876, N14851, N5451, N11087, N13257);
or OR2 (N14877, N14875, N11408);
and AND3 (N14878, N14873, N6434, N9737);
not NOT1 (N14879, N14869);
or OR3 (N14880, N14879, N2051, N8921);
xor XOR2 (N14881, N14872, N13105);
nand NAND3 (N14882, N14881, N10822, N5112);
or OR3 (N14883, N14878, N5756, N7822);
not NOT1 (N14884, N14883);
and AND4 (N14885, N14874, N14253, N8160, N6597);
and AND4 (N14886, N14862, N10856, N10822, N7061);
not NOT1 (N14887, N14885);
not NOT1 (N14888, N14877);
nand NAND3 (N14889, N14870, N4803, N8653);
not NOT1 (N14890, N14882);
or OR2 (N14891, N14889, N11737);
buf BUF1 (N14892, N14880);
not NOT1 (N14893, N14887);
not NOT1 (N14894, N14888);
buf BUF1 (N14895, N14893);
not NOT1 (N14896, N14891);
nor NOR3 (N14897, N14884, N12339, N2751);
nand NAND2 (N14898, N14886, N2175);
buf BUF1 (N14899, N14868);
buf BUF1 (N14900, N14894);
not NOT1 (N14901, N14899);
and AND3 (N14902, N14890, N1298, N9979);
not NOT1 (N14903, N14900);
not NOT1 (N14904, N14898);
buf BUF1 (N14905, N14865);
buf BUF1 (N14906, N14905);
nand NAND4 (N14907, N14876, N3170, N7855, N2195);
nand NAND2 (N14908, N14903, N2383);
or OR2 (N14909, N14908, N12444);
and AND2 (N14910, N14901, N4385);
or OR4 (N14911, N14910, N12088, N14809, N2322);
or OR3 (N14912, N14895, N2933, N1305);
not NOT1 (N14913, N14912);
nand NAND2 (N14914, N14906, N10868);
buf BUF1 (N14915, N14909);
not NOT1 (N14916, N14892);
nand NAND2 (N14917, N14907, N10086);
xor XOR2 (N14918, N14904, N12285);
nand NAND3 (N14919, N14915, N8281, N9955);
xor XOR2 (N14920, N14911, N7955);
buf BUF1 (N14921, N14913);
and AND4 (N14922, N14897, N4205, N10871, N4943);
nor NOR3 (N14923, N14916, N4688, N1805);
nand NAND2 (N14924, N14922, N1611);
nor NOR2 (N14925, N14902, N8111);
nor NOR3 (N14926, N14923, N10308, N10903);
nor NOR3 (N14927, N14926, N14478, N12713);
nand NAND2 (N14928, N14925, N10104);
nor NOR4 (N14929, N14924, N10383, N13174, N11616);
not NOT1 (N14930, N14921);
xor XOR2 (N14931, N14928, N5120);
buf BUF1 (N14932, N14896);
buf BUF1 (N14933, N14914);
not NOT1 (N14934, N14927);
or OR2 (N14935, N14931, N11221);
buf BUF1 (N14936, N14933);
and AND2 (N14937, N14918, N4430);
or OR4 (N14938, N14917, N8882, N7780, N12274);
nand NAND4 (N14939, N14937, N6998, N6730, N11678);
nor NOR2 (N14940, N14932, N4765);
or OR2 (N14941, N14938, N8298);
and AND2 (N14942, N14920, N6370);
not NOT1 (N14943, N14934);
buf BUF1 (N14944, N14941);
and AND4 (N14945, N14940, N8842, N344, N14448);
not NOT1 (N14946, N14939);
or OR3 (N14947, N14945, N6852, N14460);
not NOT1 (N14948, N14919);
nand NAND2 (N14949, N14942, N7705);
nor NOR2 (N14950, N14935, N5623);
xor XOR2 (N14951, N14936, N2135);
nor NOR3 (N14952, N14948, N7725, N8900);
nand NAND3 (N14953, N14943, N6260, N4384);
buf BUF1 (N14954, N14953);
buf BUF1 (N14955, N14951);
nor NOR3 (N14956, N14949, N13652, N4365);
xor XOR2 (N14957, N14950, N7869);
and AND2 (N14958, N14955, N13689);
and AND4 (N14959, N14952, N8011, N11366, N1419);
buf BUF1 (N14960, N14956);
not NOT1 (N14961, N14946);
nor NOR4 (N14962, N14957, N7245, N12202, N12575);
or OR4 (N14963, N14947, N7353, N8914, N13661);
nand NAND4 (N14964, N14963, N1239, N14514, N3230);
nor NOR3 (N14965, N14964, N13340, N7343);
xor XOR2 (N14966, N14958, N11374);
and AND4 (N14967, N14944, N7722, N406, N2006);
nor NOR4 (N14968, N14930, N11034, N11025, N6890);
xor XOR2 (N14969, N14966, N4417);
nand NAND3 (N14970, N14962, N4220, N10900);
and AND4 (N14971, N14968, N11938, N7881, N2591);
not NOT1 (N14972, N14970);
not NOT1 (N14973, N14965);
xor XOR2 (N14974, N14967, N14946);
or OR2 (N14975, N14972, N6337);
xor XOR2 (N14976, N14969, N3977);
buf BUF1 (N14977, N14974);
nand NAND2 (N14978, N14975, N2764);
not NOT1 (N14979, N14978);
and AND2 (N14980, N14971, N322);
nand NAND4 (N14981, N14980, N2494, N12304, N14699);
nand NAND3 (N14982, N14973, N4650, N12731);
or OR4 (N14983, N14976, N8684, N2708, N167);
xor XOR2 (N14984, N14981, N11493);
or OR2 (N14985, N14954, N12781);
nor NOR3 (N14986, N14982, N2966, N8911);
xor XOR2 (N14987, N14985, N1865);
not NOT1 (N14988, N14979);
or OR2 (N14989, N14986, N2811);
buf BUF1 (N14990, N14977);
nor NOR2 (N14991, N14961, N10810);
not NOT1 (N14992, N14987);
and AND2 (N14993, N14960, N8622);
and AND3 (N14994, N14989, N13397, N656);
nor NOR4 (N14995, N14991, N8092, N7593, N10355);
not NOT1 (N14996, N14993);
nand NAND2 (N14997, N14994, N10018);
xor XOR2 (N14998, N14997, N10827);
xor XOR2 (N14999, N14984, N824);
nand NAND3 (N15000, N14983, N11331, N2085);
or OR2 (N15001, N14959, N14032);
nor NOR3 (N15002, N15001, N14573, N6509);
and AND2 (N15003, N14996, N7277);
nand NAND4 (N15004, N15003, N6568, N4221, N6097);
nor NOR2 (N15005, N15004, N7586);
or OR2 (N15006, N14998, N13634);
buf BUF1 (N15007, N15000);
or OR3 (N15008, N15002, N6470, N14470);
xor XOR2 (N15009, N14995, N13871);
or OR3 (N15010, N15008, N12831, N2373);
buf BUF1 (N15011, N15006);
not NOT1 (N15012, N14929);
xor XOR2 (N15013, N14988, N4417);
and AND3 (N15014, N15013, N7368, N14329);
nand NAND4 (N15015, N15011, N9439, N8572, N5154);
buf BUF1 (N15016, N15007);
xor XOR2 (N15017, N14992, N6166);
nand NAND4 (N15018, N14990, N5165, N709, N9688);
nand NAND2 (N15019, N15010, N1371);
buf BUF1 (N15020, N15018);
xor XOR2 (N15021, N15015, N6264);
not NOT1 (N15022, N15016);
buf BUF1 (N15023, N15017);
or OR4 (N15024, N14999, N13667, N7881, N8022);
xor XOR2 (N15025, N15020, N2713);
nand NAND4 (N15026, N15012, N9180, N12971, N7940);
nor NOR3 (N15027, N15023, N8127, N9573);
nand NAND3 (N15028, N15025, N12249, N1609);
or OR3 (N15029, N15019, N8171, N4364);
buf BUF1 (N15030, N15026);
or OR4 (N15031, N15028, N5004, N2113, N9556);
or OR4 (N15032, N15029, N8095, N734, N12042);
nor NOR2 (N15033, N15024, N7316);
or OR4 (N15034, N15005, N5926, N8577, N1719);
and AND3 (N15035, N15033, N7552, N6383);
xor XOR2 (N15036, N15034, N3057);
nor NOR3 (N15037, N15036, N6234, N9699);
nor NOR4 (N15038, N15035, N14753, N3383, N11055);
nor NOR4 (N15039, N15014, N4923, N3108, N10008);
nand NAND4 (N15040, N15039, N765, N7317, N2375);
buf BUF1 (N15041, N15032);
nand NAND3 (N15042, N15037, N5571, N4289);
nor NOR3 (N15043, N15030, N13354, N7873);
and AND2 (N15044, N15031, N12064);
not NOT1 (N15045, N15038);
not NOT1 (N15046, N15027);
xor XOR2 (N15047, N15046, N3993);
nor NOR2 (N15048, N15041, N8936);
and AND3 (N15049, N15022, N7668, N7500);
not NOT1 (N15050, N15021);
not NOT1 (N15051, N15043);
or OR4 (N15052, N15044, N11757, N13347, N8083);
not NOT1 (N15053, N15040);
nor NOR4 (N15054, N15049, N10503, N8715, N10949);
nor NOR2 (N15055, N15045, N14491);
and AND3 (N15056, N15054, N2665, N9850);
or OR3 (N15057, N15055, N12156, N9454);
buf BUF1 (N15058, N15048);
xor XOR2 (N15059, N15050, N8498);
buf BUF1 (N15060, N15059);
not NOT1 (N15061, N15057);
buf BUF1 (N15062, N15060);
nor NOR4 (N15063, N15058, N11281, N1431, N2038);
or OR2 (N15064, N15056, N4003);
nor NOR2 (N15065, N15053, N6678);
not NOT1 (N15066, N15051);
xor XOR2 (N15067, N15062, N812);
nand NAND2 (N15068, N15047, N3998);
or OR3 (N15069, N15066, N13273, N9539);
not NOT1 (N15070, N15064);
xor XOR2 (N15071, N15042, N13269);
nand NAND2 (N15072, N15052, N2206);
buf BUF1 (N15073, N15070);
nand NAND3 (N15074, N15073, N8147, N3571);
nor NOR2 (N15075, N15068, N5359);
buf BUF1 (N15076, N15061);
xor XOR2 (N15077, N15065, N5433);
buf BUF1 (N15078, N15072);
and AND2 (N15079, N15069, N1183);
or OR3 (N15080, N15078, N12120, N13119);
and AND4 (N15081, N15067, N3187, N8398, N59);
nand NAND3 (N15082, N15081, N5849, N14864);
xor XOR2 (N15083, N15075, N1853);
nand NAND3 (N15084, N15082, N11900, N14441);
nand NAND4 (N15085, N15071, N12171, N11997, N14266);
nor NOR4 (N15086, N15009, N15043, N3605, N7413);
buf BUF1 (N15087, N15076);
nand NAND3 (N15088, N15083, N2860, N8709);
nand NAND2 (N15089, N15080, N3416);
and AND2 (N15090, N15085, N8347);
and AND4 (N15091, N15089, N4932, N12014, N3430);
nand NAND4 (N15092, N15088, N3937, N654, N13560);
or OR4 (N15093, N15087, N11537, N1239, N4734);
and AND4 (N15094, N15077, N5205, N5193, N6406);
not NOT1 (N15095, N15084);
nand NAND4 (N15096, N15079, N1966, N3189, N6234);
xor XOR2 (N15097, N15096, N1678);
not NOT1 (N15098, N15095);
and AND4 (N15099, N15063, N12452, N10913, N5056);
nor NOR4 (N15100, N15091, N1716, N362, N8868);
xor XOR2 (N15101, N15086, N6677);
or OR2 (N15102, N15099, N5225);
and AND3 (N15103, N15100, N8487, N11726);
or OR4 (N15104, N15093, N7186, N9976, N587);
buf BUF1 (N15105, N15090);
not NOT1 (N15106, N15098);
xor XOR2 (N15107, N15074, N11334);
and AND2 (N15108, N15101, N14168);
or OR2 (N15109, N15102, N10463);
or OR3 (N15110, N15103, N4702, N12414);
not NOT1 (N15111, N15094);
nand NAND2 (N15112, N15107, N14631);
nand NAND3 (N15113, N15109, N4396, N13944);
nand NAND4 (N15114, N15097, N2971, N13726, N1784);
buf BUF1 (N15115, N15112);
xor XOR2 (N15116, N15105, N9153);
and AND3 (N15117, N15110, N2926, N13916);
or OR2 (N15118, N15113, N9714);
nor NOR3 (N15119, N15116, N8603, N11119);
xor XOR2 (N15120, N15119, N3744);
buf BUF1 (N15121, N15114);
buf BUF1 (N15122, N15121);
nand NAND3 (N15123, N15115, N7570, N13035);
buf BUF1 (N15124, N15118);
nand NAND4 (N15125, N15106, N9687, N4446, N14724);
xor XOR2 (N15126, N15125, N5178);
or OR4 (N15127, N15092, N7156, N1774, N2890);
and AND4 (N15128, N15117, N4736, N1342, N6775);
nand NAND2 (N15129, N15104, N4495);
or OR2 (N15130, N15126, N9465);
nand NAND4 (N15131, N15124, N9816, N1486, N3115);
nor NOR4 (N15132, N15120, N7624, N786, N5538);
nor NOR2 (N15133, N15130, N14965);
and AND4 (N15134, N15123, N7439, N11598, N9630);
nor NOR4 (N15135, N15108, N685, N4817, N12903);
nor NOR4 (N15136, N15128, N11023, N5010, N9090);
and AND4 (N15137, N15135, N10843, N7896, N14376);
xor XOR2 (N15138, N15134, N7127);
buf BUF1 (N15139, N15122);
xor XOR2 (N15140, N15136, N12519);
xor XOR2 (N15141, N15140, N10550);
and AND3 (N15142, N15127, N4626, N8895);
not NOT1 (N15143, N15142);
not NOT1 (N15144, N15132);
buf BUF1 (N15145, N15144);
or OR3 (N15146, N15133, N15144, N13212);
and AND2 (N15147, N15139, N9720);
nand NAND2 (N15148, N15111, N13436);
nor NOR4 (N15149, N15146, N11160, N13883, N6103);
and AND3 (N15150, N15145, N11267, N584);
or OR4 (N15151, N15150, N13888, N8331, N5875);
nor NOR4 (N15152, N15137, N131, N4232, N8194);
buf BUF1 (N15153, N15138);
xor XOR2 (N15154, N15141, N4049);
or OR4 (N15155, N15148, N4762, N10603, N1572);
nand NAND3 (N15156, N15153, N11852, N8083);
not NOT1 (N15157, N15151);
or OR3 (N15158, N15156, N2168, N10792);
not NOT1 (N15159, N15147);
or OR4 (N15160, N15158, N4812, N9146, N10813);
xor XOR2 (N15161, N15154, N401);
not NOT1 (N15162, N15143);
and AND4 (N15163, N15155, N7730, N8674, N5299);
nand NAND2 (N15164, N15129, N9311);
not NOT1 (N15165, N15159);
buf BUF1 (N15166, N15164);
or OR4 (N15167, N15163, N12814, N12645, N6909);
buf BUF1 (N15168, N15161);
buf BUF1 (N15169, N15152);
buf BUF1 (N15170, N15157);
or OR3 (N15171, N15170, N2748, N13465);
nor NOR4 (N15172, N15168, N13572, N2202, N7067);
buf BUF1 (N15173, N15131);
not NOT1 (N15174, N15162);
or OR3 (N15175, N15173, N13973, N10259);
or OR2 (N15176, N15149, N948);
buf BUF1 (N15177, N15175);
nand NAND2 (N15178, N15174, N12001);
nand NAND3 (N15179, N15172, N14457, N1164);
buf BUF1 (N15180, N15167);
and AND4 (N15181, N15171, N93, N2172, N816);
not NOT1 (N15182, N15178);
nor NOR4 (N15183, N15177, N5204, N9327, N10544);
xor XOR2 (N15184, N15165, N8856);
or OR2 (N15185, N15183, N5635);
buf BUF1 (N15186, N15182);
xor XOR2 (N15187, N15179, N5767);
nor NOR4 (N15188, N15176, N9083, N8437, N7201);
and AND3 (N15189, N15184, N11239, N652);
and AND2 (N15190, N15188, N14789);
buf BUF1 (N15191, N15166);
or OR3 (N15192, N15185, N3000, N12863);
nand NAND3 (N15193, N15181, N107, N3279);
or OR2 (N15194, N15190, N7160);
nand NAND3 (N15195, N15187, N8750, N4163);
not NOT1 (N15196, N15186);
and AND2 (N15197, N15192, N12356);
not NOT1 (N15198, N15195);
nor NOR4 (N15199, N15194, N13829, N5909, N3395);
nand NAND2 (N15200, N15199, N9119);
buf BUF1 (N15201, N15169);
nor NOR2 (N15202, N15197, N5847);
or OR4 (N15203, N15191, N11560, N14685, N393);
nor NOR2 (N15204, N15203, N11886);
and AND3 (N15205, N15160, N11928, N1935);
and AND4 (N15206, N15189, N8063, N8499, N3794);
nand NAND2 (N15207, N15206, N12611);
xor XOR2 (N15208, N15180, N11558);
nand NAND3 (N15209, N15205, N3718, N8605);
or OR2 (N15210, N15202, N15016);
xor XOR2 (N15211, N15204, N289);
buf BUF1 (N15212, N15210);
nor NOR4 (N15213, N15209, N1026, N8397, N7404);
and AND2 (N15214, N15193, N1748);
not NOT1 (N15215, N15208);
buf BUF1 (N15216, N15200);
and AND4 (N15217, N15198, N796, N7216, N5674);
nor NOR4 (N15218, N15211, N1106, N1255, N7842);
nor NOR4 (N15219, N15216, N12172, N1315, N13823);
xor XOR2 (N15220, N15217, N5526);
nand NAND2 (N15221, N15219, N2599);
buf BUF1 (N15222, N15212);
nor NOR3 (N15223, N15214, N7732, N13085);
nor NOR3 (N15224, N15220, N14590, N10803);
xor XOR2 (N15225, N15201, N8506);
and AND4 (N15226, N15221, N2740, N10165, N402);
and AND3 (N15227, N15218, N7196, N14793);
and AND4 (N15228, N15223, N14066, N3994, N5443);
nand NAND4 (N15229, N15224, N11056, N8531, N10615);
not NOT1 (N15230, N15196);
xor XOR2 (N15231, N15225, N2851);
nor NOR2 (N15232, N15231, N15104);
xor XOR2 (N15233, N15213, N39);
or OR4 (N15234, N15207, N12335, N2514, N9549);
nand NAND3 (N15235, N15229, N5536, N206);
not NOT1 (N15236, N15234);
buf BUF1 (N15237, N15227);
not NOT1 (N15238, N15228);
or OR4 (N15239, N15222, N4768, N4109, N14252);
nand NAND4 (N15240, N15215, N9668, N5280, N8844);
nand NAND4 (N15241, N15237, N8821, N338, N14056);
buf BUF1 (N15242, N15226);
buf BUF1 (N15243, N15230);
or OR3 (N15244, N15241, N8907, N6688);
buf BUF1 (N15245, N15233);
not NOT1 (N15246, N15240);
buf BUF1 (N15247, N15235);
xor XOR2 (N15248, N15247, N4770);
xor XOR2 (N15249, N15236, N14209);
not NOT1 (N15250, N15245);
nand NAND2 (N15251, N15238, N3179);
and AND2 (N15252, N15242, N2270);
buf BUF1 (N15253, N15246);
not NOT1 (N15254, N15248);
buf BUF1 (N15255, N15249);
nor NOR4 (N15256, N15253, N9572, N9683, N11962);
buf BUF1 (N15257, N15250);
xor XOR2 (N15258, N15256, N2239);
and AND4 (N15259, N15251, N5898, N12460, N9766);
xor XOR2 (N15260, N15257, N10672);
buf BUF1 (N15261, N15258);
nor NOR3 (N15262, N15255, N12274, N7675);
xor XOR2 (N15263, N15260, N14945);
and AND2 (N15264, N15244, N10093);
and AND4 (N15265, N15232, N13633, N7464, N13874);
xor XOR2 (N15266, N15261, N13112);
nor NOR4 (N15267, N15259, N5163, N4917, N2696);
not NOT1 (N15268, N15252);
and AND3 (N15269, N15268, N12833, N4249);
buf BUF1 (N15270, N15264);
xor XOR2 (N15271, N15266, N14018);
xor XOR2 (N15272, N15269, N14350);
buf BUF1 (N15273, N15270);
and AND2 (N15274, N15267, N6546);
or OR4 (N15275, N15263, N3724, N10612, N4510);
buf BUF1 (N15276, N15265);
nor NOR4 (N15277, N15272, N2966, N14237, N9324);
or OR3 (N15278, N15262, N14956, N563);
nand NAND2 (N15279, N15271, N5016);
buf BUF1 (N15280, N15239);
and AND3 (N15281, N15280, N5838, N7042);
or OR4 (N15282, N15243, N4021, N11035, N7916);
not NOT1 (N15283, N15277);
not NOT1 (N15284, N15276);
xor XOR2 (N15285, N15282, N8781);
xor XOR2 (N15286, N15254, N700);
not NOT1 (N15287, N15278);
nor NOR4 (N15288, N15285, N14944, N14259, N6684);
buf BUF1 (N15289, N15273);
and AND4 (N15290, N15275, N86, N2706, N10318);
nand NAND3 (N15291, N15281, N13391, N7856);
or OR2 (N15292, N15291, N7811);
nor NOR2 (N15293, N15288, N11130);
and AND3 (N15294, N15274, N2623, N3984);
nand NAND3 (N15295, N15286, N6708, N6016);
or OR3 (N15296, N15294, N6795, N13278);
buf BUF1 (N15297, N15290);
buf BUF1 (N15298, N15289);
not NOT1 (N15299, N15287);
not NOT1 (N15300, N15293);
or OR2 (N15301, N15283, N10467);
not NOT1 (N15302, N15298);
nand NAND2 (N15303, N15297, N4250);
and AND3 (N15304, N15292, N4352, N13663);
buf BUF1 (N15305, N15304);
nand NAND4 (N15306, N15302, N11479, N7276, N12598);
xor XOR2 (N15307, N15279, N9865);
nor NOR3 (N15308, N15299, N3111, N7470);
not NOT1 (N15309, N15301);
buf BUF1 (N15310, N15300);
nand NAND3 (N15311, N15308, N3143, N11564);
or OR3 (N15312, N15284, N2351, N14930);
or OR3 (N15313, N15303, N88, N8568);
not NOT1 (N15314, N15310);
nand NAND4 (N15315, N15307, N13398, N3684, N71);
xor XOR2 (N15316, N15311, N474);
buf BUF1 (N15317, N15296);
nor NOR2 (N15318, N15312, N6582);
not NOT1 (N15319, N15314);
not NOT1 (N15320, N15319);
nor NOR3 (N15321, N15315, N8098, N4320);
nor NOR4 (N15322, N15313, N3054, N4788, N8352);
nand NAND2 (N15323, N15305, N12455);
and AND4 (N15324, N15316, N6562, N3379, N12352);
nor NOR3 (N15325, N15318, N732, N1528);
nand NAND3 (N15326, N15309, N3110, N3247);
buf BUF1 (N15327, N15322);
not NOT1 (N15328, N15327);
nand NAND4 (N15329, N15321, N1276, N7433, N11030);
not NOT1 (N15330, N15317);
or OR2 (N15331, N15329, N12036);
buf BUF1 (N15332, N15330);
buf BUF1 (N15333, N15325);
buf BUF1 (N15334, N15320);
or OR2 (N15335, N15326, N13437);
not NOT1 (N15336, N15306);
nor NOR2 (N15337, N15333, N265);
nand NAND4 (N15338, N15335, N12458, N14421, N5367);
and AND3 (N15339, N15332, N15324, N9386);
nor NOR3 (N15340, N2923, N14959, N3223);
or OR2 (N15341, N15334, N3381);
and AND4 (N15342, N15336, N5242, N9090, N14665);
nand NAND3 (N15343, N15295, N5324, N1619);
xor XOR2 (N15344, N15328, N1499);
not NOT1 (N15345, N15341);
buf BUF1 (N15346, N15343);
xor XOR2 (N15347, N15345, N6848);
xor XOR2 (N15348, N15342, N14110);
not NOT1 (N15349, N15348);
or OR4 (N15350, N15340, N3595, N14378, N5498);
buf BUF1 (N15351, N15346);
or OR2 (N15352, N15349, N9706);
and AND2 (N15353, N15351, N14733);
xor XOR2 (N15354, N15323, N14385);
nor NOR3 (N15355, N15331, N1329, N10998);
nor NOR4 (N15356, N15350, N3091, N6528, N11956);
not NOT1 (N15357, N15344);
nand NAND3 (N15358, N15354, N3383, N1223);
nand NAND4 (N15359, N15347, N9894, N12871, N14976);
or OR3 (N15360, N15353, N12635, N8347);
and AND3 (N15361, N15359, N238, N10352);
nor NOR2 (N15362, N15355, N4424);
nand NAND4 (N15363, N15352, N5312, N14834, N2511);
not NOT1 (N15364, N15362);
and AND2 (N15365, N15360, N581);
buf BUF1 (N15366, N15363);
or OR3 (N15367, N15338, N6459, N15079);
not NOT1 (N15368, N15366);
nor NOR4 (N15369, N15361, N13947, N10966, N11980);
xor XOR2 (N15370, N15339, N4385);
buf BUF1 (N15371, N15364);
buf BUF1 (N15372, N15370);
buf BUF1 (N15373, N15372);
nor NOR4 (N15374, N15357, N2251, N4387, N10891);
and AND3 (N15375, N15337, N3524, N6860);
or OR3 (N15376, N15368, N8604, N2071);
nand NAND3 (N15377, N15375, N4791, N4163);
nor NOR4 (N15378, N15374, N2418, N4973, N10123);
nand NAND2 (N15379, N15365, N9738);
nor NOR2 (N15380, N15379, N135);
or OR4 (N15381, N15358, N7765, N9294, N1913);
xor XOR2 (N15382, N15371, N1437);
nand NAND3 (N15383, N15376, N3663, N12468);
or OR3 (N15384, N15369, N1930, N14259);
and AND3 (N15385, N15367, N11746, N5388);
xor XOR2 (N15386, N15377, N3371);
and AND3 (N15387, N15378, N747, N6087);
nand NAND2 (N15388, N15383, N5986);
and AND2 (N15389, N15388, N13025);
and AND4 (N15390, N15386, N5150, N1422, N10740);
xor XOR2 (N15391, N15385, N8289);
and AND4 (N15392, N15391, N15083, N2357, N13916);
nand NAND4 (N15393, N15356, N6222, N1536, N7077);
buf BUF1 (N15394, N15389);
not NOT1 (N15395, N15394);
not NOT1 (N15396, N15382);
nand NAND4 (N15397, N15390, N9944, N4010, N4429);
xor XOR2 (N15398, N15380, N5948);
not NOT1 (N15399, N15397);
nand NAND2 (N15400, N15387, N5689);
and AND2 (N15401, N15400, N14638);
xor XOR2 (N15402, N15381, N5078);
xor XOR2 (N15403, N15396, N12795);
nand NAND4 (N15404, N15395, N9206, N9958, N10806);
or OR3 (N15405, N15403, N5473, N10720);
xor XOR2 (N15406, N15392, N5676);
buf BUF1 (N15407, N15393);
nand NAND4 (N15408, N15404, N5706, N1244, N2525);
and AND2 (N15409, N15401, N12484);
buf BUF1 (N15410, N15373);
not NOT1 (N15411, N15408);
xor XOR2 (N15412, N15411, N10950);
nand NAND2 (N15413, N15410, N2983);
buf BUF1 (N15414, N15406);
xor XOR2 (N15415, N15402, N14593);
and AND3 (N15416, N15398, N13327, N9323);
xor XOR2 (N15417, N15416, N8996);
or OR2 (N15418, N15412, N1877);
xor XOR2 (N15419, N15415, N14874);
and AND2 (N15420, N15407, N6600);
buf BUF1 (N15421, N15418);
nor NOR2 (N15422, N15384, N3775);
not NOT1 (N15423, N15409);
buf BUF1 (N15424, N15421);
nor NOR4 (N15425, N15419, N14907, N3212, N6811);
nand NAND2 (N15426, N15413, N1731);
nand NAND4 (N15427, N15422, N13865, N12206, N10442);
buf BUF1 (N15428, N15414);
xor XOR2 (N15429, N15423, N4725);
xor XOR2 (N15430, N15399, N11990);
not NOT1 (N15431, N15427);
nor NOR4 (N15432, N15430, N5038, N4112, N13302);
nand NAND2 (N15433, N15432, N10282);
not NOT1 (N15434, N15417);
and AND3 (N15435, N15420, N922, N13496);
nor NOR2 (N15436, N15429, N15150);
nand NAND2 (N15437, N15436, N555);
and AND3 (N15438, N15428, N12893, N1651);
not NOT1 (N15439, N15405);
and AND2 (N15440, N15439, N3903);
and AND4 (N15441, N15437, N9303, N8060, N14782);
not NOT1 (N15442, N15434);
nor NOR4 (N15443, N15435, N6886, N8233, N6603);
nor NOR3 (N15444, N15424, N14657, N10980);
xor XOR2 (N15445, N15443, N8789);
and AND4 (N15446, N15441, N9763, N8045, N2307);
xor XOR2 (N15447, N15445, N7722);
not NOT1 (N15448, N15431);
xor XOR2 (N15449, N15440, N1979);
or OR4 (N15450, N15449, N13486, N9455, N12671);
nand NAND3 (N15451, N15438, N11675, N15195);
and AND4 (N15452, N15448, N7442, N14009, N14347);
xor XOR2 (N15453, N15446, N11329);
buf BUF1 (N15454, N15450);
and AND4 (N15455, N15433, N3274, N12067, N2118);
or OR2 (N15456, N15444, N9347);
xor XOR2 (N15457, N15426, N8150);
nand NAND2 (N15458, N15457, N11947);
xor XOR2 (N15459, N15425, N11870);
buf BUF1 (N15460, N15453);
or OR4 (N15461, N15454, N976, N7809, N5542);
not NOT1 (N15462, N15455);
xor XOR2 (N15463, N15456, N8129);
xor XOR2 (N15464, N15452, N3442);
not NOT1 (N15465, N15442);
and AND2 (N15466, N15463, N8138);
not NOT1 (N15467, N15460);
or OR2 (N15468, N15462, N7344);
or OR2 (N15469, N15467, N12565);
xor XOR2 (N15470, N15469, N1954);
nor NOR3 (N15471, N15470, N15096, N7516);
and AND3 (N15472, N15464, N9545, N7844);
not NOT1 (N15473, N15465);
not NOT1 (N15474, N15461);
buf BUF1 (N15475, N15473);
nand NAND2 (N15476, N15459, N14735);
nand NAND2 (N15477, N15472, N8416);
not NOT1 (N15478, N15476);
not NOT1 (N15479, N15478);
nor NOR2 (N15480, N15479, N4031);
or OR4 (N15481, N15477, N5076, N15107, N9704);
or OR4 (N15482, N15481, N13205, N2938, N9152);
nor NOR4 (N15483, N15468, N10737, N1900, N14018);
xor XOR2 (N15484, N15474, N13798);
buf BUF1 (N15485, N15482);
and AND3 (N15486, N15458, N6508, N11847);
nor NOR4 (N15487, N15475, N13705, N12161, N4345);
buf BUF1 (N15488, N15487);
and AND3 (N15489, N15471, N7534, N4507);
and AND3 (N15490, N15447, N11133, N14512);
xor XOR2 (N15491, N15488, N8361);
and AND2 (N15492, N15483, N3165);
buf BUF1 (N15493, N15451);
and AND4 (N15494, N15491, N11863, N10800, N773);
nor NOR2 (N15495, N15492, N7144);
not NOT1 (N15496, N15490);
not NOT1 (N15497, N15494);
buf BUF1 (N15498, N15493);
and AND4 (N15499, N15497, N2651, N14985, N831);
nor NOR4 (N15500, N15484, N1530, N13306, N12042);
nand NAND2 (N15501, N15495, N2924);
buf BUF1 (N15502, N15500);
not NOT1 (N15503, N15501);
buf BUF1 (N15504, N15496);
or OR3 (N15505, N15486, N6677, N10524);
nor NOR3 (N15506, N15505, N4623, N1480);
or OR2 (N15507, N15506, N11326);
xor XOR2 (N15508, N15504, N14895);
nor NOR3 (N15509, N15503, N2584, N6077);
nand NAND2 (N15510, N15502, N13142);
not NOT1 (N15511, N15509);
nand NAND4 (N15512, N15499, N1203, N6819, N10339);
not NOT1 (N15513, N15507);
buf BUF1 (N15514, N15512);
xor XOR2 (N15515, N15485, N294);
xor XOR2 (N15516, N15498, N10811);
not NOT1 (N15517, N15508);
and AND3 (N15518, N15511, N10615, N1131);
or OR3 (N15519, N15489, N11999, N3736);
buf BUF1 (N15520, N15466);
nor NOR4 (N15521, N15510, N4009, N3515, N10306);
nand NAND2 (N15522, N15520, N12490);
buf BUF1 (N15523, N15522);
or OR2 (N15524, N15480, N14794);
buf BUF1 (N15525, N15519);
xor XOR2 (N15526, N15521, N12898);
nand NAND2 (N15527, N15525, N3937);
and AND3 (N15528, N15516, N11150, N1538);
not NOT1 (N15529, N15518);
buf BUF1 (N15530, N15523);
and AND3 (N15531, N15517, N8838, N8106);
not NOT1 (N15532, N15530);
or OR3 (N15533, N15524, N6006, N10001);
buf BUF1 (N15534, N15513);
nor NOR3 (N15535, N15531, N14685, N7411);
nand NAND2 (N15536, N15532, N2206);
nor NOR3 (N15537, N15536, N5612, N1054);
xor XOR2 (N15538, N15527, N8272);
buf BUF1 (N15539, N15535);
nand NAND3 (N15540, N15515, N6850, N2851);
buf BUF1 (N15541, N15529);
xor XOR2 (N15542, N15537, N6031);
nor NOR3 (N15543, N15514, N13070, N1291);
xor XOR2 (N15544, N15539, N9029);
or OR3 (N15545, N15542, N6166, N5641);
xor XOR2 (N15546, N15541, N2431);
buf BUF1 (N15547, N15543);
nor NOR3 (N15548, N15540, N7653, N3532);
and AND2 (N15549, N15545, N6553);
or OR4 (N15550, N15547, N6927, N12613, N9967);
and AND2 (N15551, N15538, N1950);
nand NAND2 (N15552, N15544, N7897);
and AND2 (N15553, N15550, N1145);
buf BUF1 (N15554, N15533);
and AND4 (N15555, N15549, N11842, N2913, N6916);
nor NOR2 (N15556, N15548, N12342);
not NOT1 (N15557, N15552);
buf BUF1 (N15558, N15534);
not NOT1 (N15559, N15546);
or OR2 (N15560, N15554, N10636);
nor NOR4 (N15561, N15551, N9238, N4209, N13271);
and AND3 (N15562, N15553, N14207, N3999);
nand NAND3 (N15563, N15559, N12111, N14195);
nor NOR4 (N15564, N15528, N12948, N3073, N12317);
and AND2 (N15565, N15563, N7141);
xor XOR2 (N15566, N15557, N11336);
nand NAND2 (N15567, N15562, N5909);
nand NAND3 (N15568, N15555, N366, N11066);
or OR4 (N15569, N15564, N6116, N13514, N11965);
and AND4 (N15570, N15561, N15139, N7733, N13773);
and AND4 (N15571, N15569, N1911, N719, N8466);
nor NOR3 (N15572, N15570, N3408, N9953);
not NOT1 (N15573, N15560);
nand NAND3 (N15574, N15568, N7771, N13115);
nor NOR4 (N15575, N15566, N13939, N8343, N10285);
xor XOR2 (N15576, N15567, N5432);
or OR4 (N15577, N15526, N311, N10913, N9612);
buf BUF1 (N15578, N15574);
nand NAND2 (N15579, N15573, N14294);
nand NAND4 (N15580, N15558, N13308, N1220, N7784);
nand NAND4 (N15581, N15575, N2017, N9728, N5340);
buf BUF1 (N15582, N15580);
not NOT1 (N15583, N15578);
not NOT1 (N15584, N15571);
not NOT1 (N15585, N15572);
xor XOR2 (N15586, N15576, N10106);
or OR3 (N15587, N15581, N9723, N11261);
nor NOR3 (N15588, N15584, N1523, N11002);
buf BUF1 (N15589, N15579);
and AND4 (N15590, N15585, N4374, N7757, N13665);
nor NOR3 (N15591, N15582, N15501, N8178);
and AND2 (N15592, N15583, N6977);
xor XOR2 (N15593, N15587, N13443);
nor NOR3 (N15594, N15586, N1870, N5877);
buf BUF1 (N15595, N15565);
nand NAND3 (N15596, N15590, N8141, N3981);
buf BUF1 (N15597, N15593);
not NOT1 (N15598, N15592);
xor XOR2 (N15599, N15594, N15491);
or OR4 (N15600, N15599, N15020, N14774, N7143);
or OR2 (N15601, N15598, N7216);
xor XOR2 (N15602, N15600, N9329);
xor XOR2 (N15603, N15556, N2550);
xor XOR2 (N15604, N15589, N14804);
buf BUF1 (N15605, N15603);
xor XOR2 (N15606, N15588, N14072);
not NOT1 (N15607, N15577);
and AND4 (N15608, N15606, N15178, N14815, N9995);
xor XOR2 (N15609, N15601, N10085);
nor NOR2 (N15610, N15604, N14577);
buf BUF1 (N15611, N15591);
xor XOR2 (N15612, N15611, N5020);
buf BUF1 (N15613, N15597);
not NOT1 (N15614, N15595);
nand NAND4 (N15615, N15605, N13046, N602, N5114);
nor NOR3 (N15616, N15612, N11498, N6293);
or OR2 (N15617, N15613, N7065);
not NOT1 (N15618, N15607);
nor NOR3 (N15619, N15616, N10151, N3065);
nor NOR4 (N15620, N15615, N6371, N15507, N5199);
nand NAND3 (N15621, N15609, N13556, N11057);
and AND3 (N15622, N15620, N8862, N10724);
nor NOR2 (N15623, N15618, N11347);
nor NOR4 (N15624, N15621, N8312, N13601, N4073);
or OR3 (N15625, N15602, N15501, N11158);
nand NAND3 (N15626, N15619, N10578, N5731);
nand NAND2 (N15627, N15625, N11420);
buf BUF1 (N15628, N15614);
nor NOR2 (N15629, N15596, N5147);
not NOT1 (N15630, N15622);
nand NAND2 (N15631, N15610, N3699);
nor NOR2 (N15632, N15623, N11759);
buf BUF1 (N15633, N15631);
nand NAND3 (N15634, N15629, N14548, N9957);
or OR2 (N15635, N15632, N6336);
and AND3 (N15636, N15630, N1048, N10279);
not NOT1 (N15637, N15617);
nor NOR3 (N15638, N15635, N15464, N507);
not NOT1 (N15639, N15633);
nand NAND3 (N15640, N15634, N12942, N8130);
and AND3 (N15641, N15627, N1726, N14256);
xor XOR2 (N15642, N15637, N6798);
xor XOR2 (N15643, N15626, N1328);
buf BUF1 (N15644, N15640);
nor NOR3 (N15645, N15628, N5898, N14226);
or OR4 (N15646, N15645, N8578, N9692, N12652);
and AND3 (N15647, N15643, N9402, N13278);
and AND2 (N15648, N15639, N8125);
nand NAND3 (N15649, N15648, N9657, N10257);
nand NAND3 (N15650, N15636, N3146, N4747);
nand NAND3 (N15651, N15644, N3154, N321);
or OR2 (N15652, N15642, N1552);
nand NAND3 (N15653, N15608, N9981, N4349);
buf BUF1 (N15654, N15651);
or OR2 (N15655, N15653, N13133);
and AND3 (N15656, N15646, N4165, N12749);
xor XOR2 (N15657, N15624, N5082);
not NOT1 (N15658, N15652);
nand NAND2 (N15659, N15654, N5237);
nor NOR3 (N15660, N15657, N3845, N14592);
not NOT1 (N15661, N15641);
buf BUF1 (N15662, N15659);
nor NOR2 (N15663, N15650, N347);
and AND4 (N15664, N15656, N4134, N9198, N3361);
nand NAND4 (N15665, N15649, N3558, N5258, N5062);
not NOT1 (N15666, N15638);
nor NOR4 (N15667, N15660, N13667, N213, N3728);
buf BUF1 (N15668, N15664);
nor NOR3 (N15669, N15667, N6888, N9736);
xor XOR2 (N15670, N15668, N1608);
xor XOR2 (N15671, N15663, N4381);
nand NAND2 (N15672, N15647, N1827);
and AND3 (N15673, N15669, N14658, N5905);
buf BUF1 (N15674, N15671);
xor XOR2 (N15675, N15674, N2336);
not NOT1 (N15676, N15675);
nor NOR2 (N15677, N15673, N7590);
or OR4 (N15678, N15662, N5555, N2710, N9725);
nand NAND4 (N15679, N15678, N4811, N7286, N15441);
and AND2 (N15680, N15679, N9584);
not NOT1 (N15681, N15666);
xor XOR2 (N15682, N15677, N7296);
buf BUF1 (N15683, N15672);
and AND3 (N15684, N15680, N578, N9790);
and AND3 (N15685, N15655, N10386, N7317);
and AND4 (N15686, N15681, N9732, N810, N13189);
or OR3 (N15687, N15661, N14942, N12126);
xor XOR2 (N15688, N15684, N7965);
not NOT1 (N15689, N15682);
nand NAND3 (N15690, N15687, N12151, N6838);
nand NAND4 (N15691, N15670, N14246, N433, N13754);
nor NOR3 (N15692, N15691, N11069, N15389);
nor NOR4 (N15693, N15686, N11182, N11101, N1578);
nand NAND3 (N15694, N15658, N144, N12613);
nand NAND3 (N15695, N15689, N12643, N11172);
xor XOR2 (N15696, N15690, N4274);
and AND3 (N15697, N15693, N6971, N3699);
xor XOR2 (N15698, N15697, N9618);
nand NAND2 (N15699, N15683, N10715);
nor NOR4 (N15700, N15695, N13626, N6982, N15187);
xor XOR2 (N15701, N15694, N318);
and AND4 (N15702, N15699, N1126, N11656, N6651);
or OR2 (N15703, N15696, N12273);
not NOT1 (N15704, N15688);
and AND2 (N15705, N15665, N11120);
nand NAND3 (N15706, N15704, N4831, N11813);
not NOT1 (N15707, N15702);
and AND4 (N15708, N15705, N13192, N10590, N10342);
or OR3 (N15709, N15698, N13844, N8055);
buf BUF1 (N15710, N15707);
nand NAND4 (N15711, N15701, N283, N2811, N7858);
xor XOR2 (N15712, N15676, N10158);
xor XOR2 (N15713, N15709, N9081);
and AND2 (N15714, N15703, N12594);
nand NAND3 (N15715, N15713, N4943, N3008);
nand NAND4 (N15716, N15685, N6650, N9479, N8170);
xor XOR2 (N15717, N15692, N7250);
nor NOR4 (N15718, N15714, N695, N8131, N6544);
not NOT1 (N15719, N15715);
or OR3 (N15720, N15716, N8450, N3234);
nand NAND2 (N15721, N15710, N9820);
not NOT1 (N15722, N15706);
xor XOR2 (N15723, N15712, N10497);
nor NOR2 (N15724, N15711, N7734);
not NOT1 (N15725, N15708);
or OR4 (N15726, N15720, N10866, N3968, N3937);
nor NOR2 (N15727, N15723, N1732);
not NOT1 (N15728, N15717);
xor XOR2 (N15729, N15722, N11111);
nor NOR3 (N15730, N15700, N1457, N10830);
and AND2 (N15731, N15727, N10827);
or OR3 (N15732, N15718, N12202, N9728);
and AND4 (N15733, N15725, N943, N6168, N14387);
and AND3 (N15734, N15721, N4616, N1565);
buf BUF1 (N15735, N15719);
and AND3 (N15736, N15735, N1752, N9164);
nand NAND2 (N15737, N15726, N2668);
and AND2 (N15738, N15734, N11667);
not NOT1 (N15739, N15736);
xor XOR2 (N15740, N15729, N1910);
xor XOR2 (N15741, N15724, N9274);
xor XOR2 (N15742, N15738, N11486);
and AND2 (N15743, N15733, N3579);
and AND2 (N15744, N15731, N12958);
nor NOR4 (N15745, N15737, N3043, N12747, N10030);
nand NAND2 (N15746, N15743, N9357);
buf BUF1 (N15747, N15742);
and AND4 (N15748, N15744, N8057, N3958, N682);
xor XOR2 (N15749, N15748, N13719);
nand NAND2 (N15750, N15745, N6069);
buf BUF1 (N15751, N15741);
xor XOR2 (N15752, N15750, N1382);
not NOT1 (N15753, N15751);
nor NOR3 (N15754, N15749, N6509, N9012);
xor XOR2 (N15755, N15747, N13629);
nand NAND4 (N15756, N15728, N10159, N10799, N1778);
buf BUF1 (N15757, N15739);
and AND2 (N15758, N15756, N2110);
not NOT1 (N15759, N15757);
nand NAND2 (N15760, N15755, N5202);
buf BUF1 (N15761, N15730);
not NOT1 (N15762, N15746);
or OR4 (N15763, N15753, N4246, N5478, N14081);
xor XOR2 (N15764, N15752, N790);
nand NAND4 (N15765, N15754, N10515, N2466, N1201);
or OR3 (N15766, N15758, N12145, N12670);
or OR2 (N15767, N15766, N5675);
buf BUF1 (N15768, N15763);
nand NAND4 (N15769, N15761, N107, N12016, N2556);
and AND4 (N15770, N15760, N5701, N4027, N15752);
or OR2 (N15771, N15759, N15146);
nor NOR4 (N15772, N15762, N11860, N15396, N13398);
nand NAND3 (N15773, N15740, N7347, N14273);
nand NAND2 (N15774, N15770, N2738);
and AND2 (N15775, N15773, N12987);
xor XOR2 (N15776, N15771, N8872);
not NOT1 (N15777, N15765);
and AND4 (N15778, N15764, N12019, N2823, N10755);
nand NAND4 (N15779, N15732, N14859, N12841, N4092);
not NOT1 (N15780, N15776);
nor NOR3 (N15781, N15778, N7899, N1156);
or OR4 (N15782, N15781, N638, N7572, N1256);
nand NAND3 (N15783, N15777, N15669, N2363);
or OR2 (N15784, N15775, N9825);
xor XOR2 (N15785, N15783, N10405);
and AND2 (N15786, N15774, N15035);
and AND4 (N15787, N15767, N1191, N449, N9290);
nor NOR3 (N15788, N15785, N6242, N11930);
nand NAND4 (N15789, N15784, N3540, N10958, N10283);
buf BUF1 (N15790, N15788);
and AND3 (N15791, N15790, N5225, N12998);
xor XOR2 (N15792, N15772, N15278);
buf BUF1 (N15793, N15779);
buf BUF1 (N15794, N15768);
buf BUF1 (N15795, N15787);
buf BUF1 (N15796, N15782);
xor XOR2 (N15797, N15789, N9201);
xor XOR2 (N15798, N15796, N1975);
xor XOR2 (N15799, N15798, N3726);
not NOT1 (N15800, N15797);
or OR3 (N15801, N15793, N8106, N10387);
xor XOR2 (N15802, N15799, N3193);
nor NOR3 (N15803, N15769, N5797, N10124);
xor XOR2 (N15804, N15780, N14570);
and AND4 (N15805, N15786, N13975, N5455, N423);
nand NAND4 (N15806, N15794, N9391, N4667, N12314);
buf BUF1 (N15807, N15801);
buf BUF1 (N15808, N15804);
nand NAND3 (N15809, N15803, N2383, N7518);
not NOT1 (N15810, N15795);
or OR3 (N15811, N15810, N7604, N6473);
not NOT1 (N15812, N15809);
nand NAND3 (N15813, N15807, N9816, N12426);
nor NOR2 (N15814, N15791, N9001);
buf BUF1 (N15815, N15811);
xor XOR2 (N15816, N15800, N6044);
nor NOR3 (N15817, N15792, N2711, N11375);
and AND4 (N15818, N15815, N8610, N8592, N13923);
nor NOR3 (N15819, N15818, N5229, N4040);
or OR3 (N15820, N15813, N2121, N4899);
xor XOR2 (N15821, N15814, N3928);
or OR4 (N15822, N15821, N14499, N11306, N4750);
buf BUF1 (N15823, N15805);
xor XOR2 (N15824, N15817, N3218);
not NOT1 (N15825, N15806);
or OR3 (N15826, N15819, N12466, N2862);
buf BUF1 (N15827, N15802);
buf BUF1 (N15828, N15808);
or OR3 (N15829, N15812, N1309, N5526);
buf BUF1 (N15830, N15823);
xor XOR2 (N15831, N15826, N10339);
xor XOR2 (N15832, N15822, N15028);
and AND2 (N15833, N15830, N8931);
or OR2 (N15834, N15832, N8307);
not NOT1 (N15835, N15825);
buf BUF1 (N15836, N15824);
buf BUF1 (N15837, N15827);
nand NAND4 (N15838, N15837, N13310, N12700, N8114);
or OR2 (N15839, N15836, N8140);
nand NAND3 (N15840, N15834, N3701, N14767);
nand NAND2 (N15841, N15839, N8667);
or OR4 (N15842, N15833, N4134, N15564, N12037);
nand NAND3 (N15843, N15820, N2703, N1526);
or OR4 (N15844, N15829, N75, N1434, N1969);
not NOT1 (N15845, N15828);
nor NOR4 (N15846, N15816, N10440, N11201, N3650);
or OR4 (N15847, N15838, N10293, N5574, N9048);
not NOT1 (N15848, N15844);
not NOT1 (N15849, N15847);
xor XOR2 (N15850, N15849, N6389);
xor XOR2 (N15851, N15831, N5693);
not NOT1 (N15852, N15842);
buf BUF1 (N15853, N15843);
and AND3 (N15854, N15845, N4085, N534);
buf BUF1 (N15855, N15852);
buf BUF1 (N15856, N15850);
nor NOR3 (N15857, N15840, N3625, N13761);
nand NAND3 (N15858, N15851, N15292, N2819);
buf BUF1 (N15859, N15857);
xor XOR2 (N15860, N15855, N9742);
xor XOR2 (N15861, N15859, N7569);
or OR4 (N15862, N15848, N463, N3382, N15367);
or OR2 (N15863, N15862, N910);
xor XOR2 (N15864, N15853, N10351);
buf BUF1 (N15865, N15846);
and AND4 (N15866, N15864, N5335, N7915, N2205);
not NOT1 (N15867, N15854);
nand NAND2 (N15868, N15863, N15799);
xor XOR2 (N15869, N15868, N4080);
xor XOR2 (N15870, N15865, N296);
xor XOR2 (N15871, N15869, N8910);
nor NOR2 (N15872, N15858, N14688);
buf BUF1 (N15873, N15860);
xor XOR2 (N15874, N15841, N8955);
nand NAND2 (N15875, N15873, N15052);
nand NAND3 (N15876, N15874, N4889, N6085);
xor XOR2 (N15877, N15871, N6408);
nand NAND3 (N15878, N15861, N7257, N4682);
buf BUF1 (N15879, N15866);
not NOT1 (N15880, N15856);
nor NOR3 (N15881, N15835, N1492, N2732);
not NOT1 (N15882, N15881);
nor NOR4 (N15883, N15878, N8995, N12069, N11167);
and AND3 (N15884, N15867, N6514, N5880);
buf BUF1 (N15885, N15882);
or OR3 (N15886, N15876, N6477, N9826);
xor XOR2 (N15887, N15872, N13460);
xor XOR2 (N15888, N15886, N224);
or OR3 (N15889, N15875, N2959, N14417);
or OR4 (N15890, N15880, N9596, N1750, N9777);
and AND2 (N15891, N15879, N3451);
xor XOR2 (N15892, N15877, N14808);
nand NAND4 (N15893, N15890, N3253, N9824, N3652);
or OR3 (N15894, N15892, N5158, N10708);
xor XOR2 (N15895, N15894, N15855);
nor NOR4 (N15896, N15895, N12802, N9009, N7785);
xor XOR2 (N15897, N15870, N7887);
nor NOR2 (N15898, N15897, N10611);
nand NAND4 (N15899, N15883, N14143, N8475, N4752);
nand NAND3 (N15900, N15889, N1556, N15075);
and AND3 (N15901, N15885, N10692, N9490);
xor XOR2 (N15902, N15898, N2690);
or OR2 (N15903, N15887, N3491);
or OR2 (N15904, N15893, N12237);
nand NAND2 (N15905, N15896, N5522);
nor NOR3 (N15906, N15905, N2368, N15113);
buf BUF1 (N15907, N15884);
nor NOR3 (N15908, N15902, N4714, N15631);
xor XOR2 (N15909, N15908, N7079);
nor NOR2 (N15910, N15906, N3171);
xor XOR2 (N15911, N15900, N12822);
buf BUF1 (N15912, N15891);
and AND4 (N15913, N15899, N3760, N12802, N5479);
xor XOR2 (N15914, N15904, N12521);
nand NAND4 (N15915, N15910, N6658, N2208, N1538);
not NOT1 (N15916, N15907);
xor XOR2 (N15917, N15916, N683);
nand NAND3 (N15918, N15888, N6589, N7602);
or OR3 (N15919, N15914, N9486, N10411);
and AND3 (N15920, N15915, N15416, N2438);
nor NOR3 (N15921, N15920, N11803, N9554);
not NOT1 (N15922, N15903);
or OR3 (N15923, N15909, N2782, N2502);
nand NAND3 (N15924, N15919, N3456, N8520);
or OR4 (N15925, N15923, N1324, N4326, N6229);
nor NOR2 (N15926, N15924, N8821);
nor NOR2 (N15927, N15925, N3249);
not NOT1 (N15928, N15913);
xor XOR2 (N15929, N15928, N1192);
xor XOR2 (N15930, N15911, N2422);
not NOT1 (N15931, N15921);
xor XOR2 (N15932, N15930, N2914);
and AND2 (N15933, N15901, N1403);
or OR2 (N15934, N15931, N2632);
nor NOR2 (N15935, N15932, N6049);
not NOT1 (N15936, N15922);
and AND2 (N15937, N15933, N7217);
and AND4 (N15938, N15926, N3902, N5326, N10020);
xor XOR2 (N15939, N15929, N11639);
and AND3 (N15940, N15927, N15248, N2887);
nor NOR2 (N15941, N15934, N15254);
buf BUF1 (N15942, N15912);
nor NOR4 (N15943, N15936, N10908, N7519, N14168);
nand NAND3 (N15944, N15943, N1360, N2405);
buf BUF1 (N15945, N15939);
buf BUF1 (N15946, N15918);
nor NOR4 (N15947, N15940, N8922, N15262, N2961);
xor XOR2 (N15948, N15947, N5422);
xor XOR2 (N15949, N15938, N10879);
not NOT1 (N15950, N15937);
buf BUF1 (N15951, N15935);
nor NOR3 (N15952, N15917, N10201, N7509);
xor XOR2 (N15953, N15946, N7730);
nor NOR2 (N15954, N15949, N2594);
buf BUF1 (N15955, N15945);
xor XOR2 (N15956, N15954, N11689);
nand NAND4 (N15957, N15955, N12030, N14, N15503);
or OR4 (N15958, N15952, N6055, N11845, N11476);
or OR4 (N15959, N15941, N14145, N2517, N1500);
not NOT1 (N15960, N15953);
and AND4 (N15961, N15957, N15226, N9651, N486);
and AND3 (N15962, N15958, N7191, N12728);
nor NOR2 (N15963, N15951, N4686);
and AND4 (N15964, N15944, N6020, N11992, N3397);
not NOT1 (N15965, N15961);
and AND4 (N15966, N15962, N15611, N9472, N7021);
xor XOR2 (N15967, N15965, N3135);
buf BUF1 (N15968, N15963);
or OR3 (N15969, N15948, N15897, N10441);
and AND3 (N15970, N15969, N14833, N2002);
xor XOR2 (N15971, N15960, N3676);
nor NOR2 (N15972, N15956, N7714);
or OR4 (N15973, N15942, N4816, N1625, N4441);
nand NAND4 (N15974, N15964, N15946, N1689, N8202);
xor XOR2 (N15975, N15971, N11771);
and AND4 (N15976, N15975, N10281, N14036, N12046);
nor NOR2 (N15977, N15967, N433);
nand NAND2 (N15978, N15966, N274);
and AND4 (N15979, N15977, N10034, N3223, N5785);
nor NOR3 (N15980, N15970, N4365, N5806);
xor XOR2 (N15981, N15950, N12790);
or OR4 (N15982, N15973, N965, N1170, N15148);
buf BUF1 (N15983, N15982);
nand NAND3 (N15984, N15980, N15197, N3197);
buf BUF1 (N15985, N15976);
not NOT1 (N15986, N15979);
and AND4 (N15987, N15985, N12635, N13232, N13581);
or OR4 (N15988, N15968, N11758, N7444, N10262);
xor XOR2 (N15989, N15983, N12220);
xor XOR2 (N15990, N15972, N13980);
and AND4 (N15991, N15984, N8295, N8904, N1102);
or OR4 (N15992, N15981, N14703, N15147, N1854);
buf BUF1 (N15993, N15974);
buf BUF1 (N15994, N15959);
nor NOR3 (N15995, N15987, N13330, N6438);
xor XOR2 (N15996, N15990, N739);
buf BUF1 (N15997, N15992);
xor XOR2 (N15998, N15988, N11956);
nor NOR3 (N15999, N15998, N7379, N5640);
nor NOR2 (N16000, N15978, N12812);
buf BUF1 (N16001, N15999);
and AND3 (N16002, N15994, N12919, N12598);
not NOT1 (N16003, N15986);
and AND4 (N16004, N15993, N12120, N3710, N5013);
or OR3 (N16005, N15997, N15020, N6067);
or OR3 (N16006, N16005, N1184, N4270);
nand NAND3 (N16007, N16000, N3750, N3492);
nor NOR3 (N16008, N15989, N4239, N11175);
not NOT1 (N16009, N16007);
and AND3 (N16010, N16006, N9552, N5881);
nor NOR3 (N16011, N16008, N8068, N4550);
nand NAND4 (N16012, N16011, N14263, N5658, N9375);
buf BUF1 (N16013, N15995);
nor NOR2 (N16014, N16001, N2148);
nand NAND4 (N16015, N16012, N14044, N9356, N9870);
and AND2 (N16016, N16010, N7799);
and AND4 (N16017, N16002, N10226, N13359, N1559);
and AND4 (N16018, N16017, N8632, N6247, N14796);
nand NAND2 (N16019, N16016, N13893);
nand NAND4 (N16020, N16003, N7364, N5119, N8134);
or OR2 (N16021, N16013, N1596);
or OR4 (N16022, N16014, N7089, N5616, N6591);
nand NAND2 (N16023, N16009, N7640);
nor NOR3 (N16024, N16019, N10557, N3442);
nand NAND2 (N16025, N16021, N15233);
or OR3 (N16026, N16024, N4780, N8691);
and AND2 (N16027, N16025, N1300);
xor XOR2 (N16028, N16023, N13733);
and AND4 (N16029, N15996, N15804, N5765, N5347);
nor NOR3 (N16030, N16004, N6783, N737);
and AND3 (N16031, N16028, N3216, N10657);
not NOT1 (N16032, N16020);
nand NAND2 (N16033, N16027, N4595);
and AND2 (N16034, N16031, N6702);
nand NAND4 (N16035, N16026, N11338, N3726, N8746);
not NOT1 (N16036, N16029);
buf BUF1 (N16037, N16022);
or OR2 (N16038, N16030, N3814);
or OR4 (N16039, N16034, N6822, N14177, N14375);
nand NAND4 (N16040, N16035, N5346, N5214, N5639);
nor NOR4 (N16041, N16040, N1566, N1707, N2208);
or OR2 (N16042, N16038, N3401);
or OR3 (N16043, N16018, N5255, N9970);
buf BUF1 (N16044, N16032);
nor NOR3 (N16045, N16033, N1337, N5536);
nor NOR3 (N16046, N15991, N15164, N7636);
nor NOR2 (N16047, N16044, N15923);
buf BUF1 (N16048, N16015);
not NOT1 (N16049, N16036);
nor NOR4 (N16050, N16041, N4214, N10213, N4508);
or OR3 (N16051, N16050, N11803, N1542);
not NOT1 (N16052, N16051);
not NOT1 (N16053, N16043);
and AND2 (N16054, N16042, N2828);
or OR4 (N16055, N16052, N12940, N7970, N8996);
nor NOR2 (N16056, N16055, N7510);
or OR4 (N16057, N16049, N8619, N1733, N12665);
nand NAND3 (N16058, N16047, N4649, N5215);
nand NAND2 (N16059, N16054, N361);
and AND3 (N16060, N16048, N2755, N7840);
nand NAND2 (N16061, N16058, N314);
nor NOR3 (N16062, N16046, N8014, N12529);
nand NAND3 (N16063, N16037, N14674, N4166);
nor NOR2 (N16064, N16039, N7887);
buf BUF1 (N16065, N16061);
or OR4 (N16066, N16053, N11037, N12421, N2100);
xor XOR2 (N16067, N16060, N1364);
nor NOR2 (N16068, N16062, N12780);
not NOT1 (N16069, N16064);
nand NAND2 (N16070, N16065, N12298);
nor NOR4 (N16071, N16066, N7884, N12768, N1136);
and AND4 (N16072, N16071, N5194, N11144, N11775);
not NOT1 (N16073, N16063);
not NOT1 (N16074, N16068);
not NOT1 (N16075, N16072);
buf BUF1 (N16076, N16070);
nor NOR4 (N16077, N16057, N382, N4316, N14543);
nand NAND3 (N16078, N16056, N11239, N9878);
or OR3 (N16079, N16075, N15651, N14210);
or OR4 (N16080, N16076, N8157, N8554, N4085);
not NOT1 (N16081, N16080);
xor XOR2 (N16082, N16059, N12813);
or OR4 (N16083, N16079, N275, N4229, N10708);
nand NAND3 (N16084, N16073, N13196, N13927);
and AND4 (N16085, N16084, N4152, N5615, N13223);
not NOT1 (N16086, N16078);
nor NOR2 (N16087, N16069, N11394);
and AND4 (N16088, N16087, N1202, N15992, N6748);
buf BUF1 (N16089, N16082);
buf BUF1 (N16090, N16086);
buf BUF1 (N16091, N16074);
and AND2 (N16092, N16081, N7225);
buf BUF1 (N16093, N16089);
xor XOR2 (N16094, N16091, N8441);
buf BUF1 (N16095, N16077);
nor NOR4 (N16096, N16067, N8676, N1959, N6268);
or OR4 (N16097, N16092, N267, N15162, N9921);
nand NAND3 (N16098, N16097, N14874, N9340);
not NOT1 (N16099, N16045);
nand NAND3 (N16100, N16096, N12798, N15757);
or OR2 (N16101, N16093, N12369);
xor XOR2 (N16102, N16098, N8326);
not NOT1 (N16103, N16102);
nor NOR3 (N16104, N16103, N12911, N14832);
or OR3 (N16105, N16100, N11655, N7224);
and AND3 (N16106, N16101, N12333, N10795);
nand NAND2 (N16107, N16095, N12240);
nor NOR3 (N16108, N16094, N3062, N7444);
buf BUF1 (N16109, N16088);
and AND2 (N16110, N16106, N1666);
and AND4 (N16111, N16083, N8493, N13828, N7144);
nor NOR4 (N16112, N16085, N1918, N14026, N1177);
nand NAND4 (N16113, N16110, N1556, N1218, N4020);
not NOT1 (N16114, N16109);
xor XOR2 (N16115, N16090, N6852);
not NOT1 (N16116, N16112);
nand NAND4 (N16117, N16108, N10694, N3290, N5377);
not NOT1 (N16118, N16114);
or OR4 (N16119, N16105, N1006, N11508, N10156);
xor XOR2 (N16120, N16116, N3892);
nor NOR3 (N16121, N16117, N11086, N6053);
xor XOR2 (N16122, N16121, N15463);
or OR3 (N16123, N16118, N13043, N15919);
and AND3 (N16124, N16113, N5396, N15457);
nor NOR2 (N16125, N16104, N8258);
or OR4 (N16126, N16115, N4160, N1360, N14207);
buf BUF1 (N16127, N16122);
not NOT1 (N16128, N16127);
buf BUF1 (N16129, N16125);
not NOT1 (N16130, N16129);
buf BUF1 (N16131, N16128);
or OR2 (N16132, N16130, N16018);
not NOT1 (N16133, N16107);
or OR3 (N16134, N16099, N523, N8916);
nand NAND4 (N16135, N16123, N15108, N12310, N13190);
xor XOR2 (N16136, N16120, N4045);
not NOT1 (N16137, N16132);
xor XOR2 (N16138, N16124, N4217);
buf BUF1 (N16139, N16133);
or OR4 (N16140, N16138, N8619, N5498, N1634);
xor XOR2 (N16141, N16126, N11029);
nor NOR2 (N16142, N16141, N7911);
not NOT1 (N16143, N16131);
and AND3 (N16144, N16139, N8391, N6604);
or OR3 (N16145, N16136, N13839, N5362);
nor NOR4 (N16146, N16134, N14102, N8959, N5720);
nand NAND3 (N16147, N16144, N8678, N4958);
or OR4 (N16148, N16135, N12465, N15636, N8820);
buf BUF1 (N16149, N16140);
not NOT1 (N16150, N16147);
nor NOR3 (N16151, N16148, N4671, N5178);
xor XOR2 (N16152, N16119, N10892);
nand NAND2 (N16153, N16152, N2380);
not NOT1 (N16154, N16111);
xor XOR2 (N16155, N16146, N2257);
nand NAND3 (N16156, N16142, N1725, N610);
or OR4 (N16157, N16150, N8951, N5925, N7365);
nor NOR2 (N16158, N16153, N3579);
or OR2 (N16159, N16145, N221);
or OR3 (N16160, N16143, N1138, N13731);
nor NOR2 (N16161, N16156, N12361);
nor NOR2 (N16162, N16159, N14244);
not NOT1 (N16163, N16157);
nor NOR4 (N16164, N16162, N9548, N9145, N10241);
buf BUF1 (N16165, N16149);
nor NOR4 (N16166, N16158, N15420, N14406, N3787);
xor XOR2 (N16167, N16160, N489);
and AND3 (N16168, N16166, N13044, N2748);
nand NAND3 (N16169, N16165, N8462, N14619);
not NOT1 (N16170, N16161);
not NOT1 (N16171, N16154);
or OR4 (N16172, N16163, N12441, N1568, N15982);
buf BUF1 (N16173, N16155);
buf BUF1 (N16174, N16173);
xor XOR2 (N16175, N16168, N10752);
nand NAND4 (N16176, N16172, N3825, N2658, N8689);
xor XOR2 (N16177, N16176, N13820);
or OR4 (N16178, N16164, N3777, N493, N1656);
and AND3 (N16179, N16175, N8924, N13106);
nand NAND4 (N16180, N16171, N934, N5808, N12667);
and AND4 (N16181, N16169, N932, N11460, N9264);
nand NAND3 (N16182, N16137, N4732, N10028);
and AND4 (N16183, N16178, N14222, N7787, N15091);
or OR4 (N16184, N16183, N7109, N8097, N13280);
nand NAND2 (N16185, N16174, N8923);
nor NOR4 (N16186, N16181, N5039, N999, N8336);
xor XOR2 (N16187, N16185, N7688);
nand NAND4 (N16188, N16186, N8102, N9377, N9383);
not NOT1 (N16189, N16184);
nand NAND4 (N16190, N16189, N15420, N12572, N15009);
not NOT1 (N16191, N16179);
not NOT1 (N16192, N16151);
nor NOR2 (N16193, N16190, N15030);
xor XOR2 (N16194, N16180, N8670);
nor NOR4 (N16195, N16188, N4335, N8447, N1974);
xor XOR2 (N16196, N16187, N7745);
not NOT1 (N16197, N16182);
nor NOR2 (N16198, N16197, N7678);
xor XOR2 (N16199, N16195, N5887);
and AND2 (N16200, N16194, N15214);
buf BUF1 (N16201, N16191);
buf BUF1 (N16202, N16193);
buf BUF1 (N16203, N16200);
buf BUF1 (N16204, N16196);
not NOT1 (N16205, N16198);
nand NAND4 (N16206, N16170, N14957, N8327, N10667);
buf BUF1 (N16207, N16204);
xor XOR2 (N16208, N16167, N12575);
buf BUF1 (N16209, N16201);
buf BUF1 (N16210, N16199);
nand NAND3 (N16211, N16202, N4876, N296);
and AND3 (N16212, N16203, N4091, N648);
not NOT1 (N16213, N16208);
and AND4 (N16214, N16205, N14774, N6254, N10632);
nand NAND2 (N16215, N16213, N14628);
or OR4 (N16216, N16212, N5229, N8864, N832);
not NOT1 (N16217, N16216);
buf BUF1 (N16218, N16192);
and AND4 (N16219, N16218, N10203, N9188, N14373);
nand NAND3 (N16220, N16207, N8776, N2268);
nor NOR2 (N16221, N16215, N12815);
nand NAND4 (N16222, N16214, N3111, N15204, N2549);
xor XOR2 (N16223, N16177, N4666);
buf BUF1 (N16224, N16210);
buf BUF1 (N16225, N16221);
not NOT1 (N16226, N16217);
xor XOR2 (N16227, N16222, N8378);
or OR4 (N16228, N16220, N6356, N15992, N11602);
and AND3 (N16229, N16209, N7737, N10142);
nor NOR4 (N16230, N16228, N11966, N4289, N15673);
not NOT1 (N16231, N16211);
buf BUF1 (N16232, N16231);
nand NAND3 (N16233, N16224, N12029, N4973);
nand NAND2 (N16234, N16225, N9972);
xor XOR2 (N16235, N16233, N13217);
buf BUF1 (N16236, N16219);
and AND2 (N16237, N16232, N4376);
buf BUF1 (N16238, N16237);
nand NAND2 (N16239, N16235, N11782);
not NOT1 (N16240, N16206);
or OR3 (N16241, N16234, N4174, N6941);
nor NOR3 (N16242, N16226, N16153, N11380);
or OR3 (N16243, N16238, N9920, N13494);
or OR3 (N16244, N16227, N12642, N5193);
not NOT1 (N16245, N16242);
xor XOR2 (N16246, N16229, N4660);
xor XOR2 (N16247, N16241, N1145);
nor NOR4 (N16248, N16247, N4101, N15415, N9816);
buf BUF1 (N16249, N16246);
and AND4 (N16250, N16248, N12322, N1178, N4001);
nor NOR4 (N16251, N16236, N4975, N4078, N14223);
or OR3 (N16252, N16251, N4456, N9965);
nand NAND3 (N16253, N16249, N240, N7661);
or OR3 (N16254, N16253, N4504, N6907);
and AND4 (N16255, N16230, N8931, N15175, N14713);
and AND2 (N16256, N16240, N12175);
or OR2 (N16257, N16244, N7808);
buf BUF1 (N16258, N16257);
nor NOR2 (N16259, N16252, N8103);
or OR3 (N16260, N16223, N5008, N10535);
not NOT1 (N16261, N16245);
or OR4 (N16262, N16260, N14416, N6218, N12085);
buf BUF1 (N16263, N16243);
not NOT1 (N16264, N16263);
xor XOR2 (N16265, N16250, N529);
buf BUF1 (N16266, N16262);
buf BUF1 (N16267, N16261);
or OR2 (N16268, N16258, N4854);
nand NAND4 (N16269, N16265, N992, N218, N498);
nor NOR2 (N16270, N16264, N10634);
buf BUF1 (N16271, N16239);
and AND3 (N16272, N16268, N8145, N8428);
xor XOR2 (N16273, N16256, N9319);
nor NOR4 (N16274, N16266, N14850, N5178, N9409);
not NOT1 (N16275, N16259);
not NOT1 (N16276, N16272);
nor NOR2 (N16277, N16273, N10946);
and AND2 (N16278, N16276, N3999);
or OR2 (N16279, N16269, N8878);
xor XOR2 (N16280, N16279, N3741);
or OR4 (N16281, N16275, N3840, N10585, N2162);
buf BUF1 (N16282, N16281);
buf BUF1 (N16283, N16254);
nor NOR2 (N16284, N16277, N8506);
xor XOR2 (N16285, N16280, N1720);
and AND3 (N16286, N16270, N6856, N307);
nor NOR3 (N16287, N16267, N13642, N818);
nand NAND3 (N16288, N16283, N2926, N2634);
or OR2 (N16289, N16274, N8281);
not NOT1 (N16290, N16288);
not NOT1 (N16291, N16287);
xor XOR2 (N16292, N16278, N11064);
and AND2 (N16293, N16271, N13569);
not NOT1 (N16294, N16290);
buf BUF1 (N16295, N16255);
xor XOR2 (N16296, N16289, N11631);
xor XOR2 (N16297, N16282, N7867);
not NOT1 (N16298, N16285);
and AND4 (N16299, N16295, N7841, N13684, N9285);
buf BUF1 (N16300, N16296);
and AND4 (N16301, N16297, N1977, N4710, N8311);
nor NOR3 (N16302, N16301, N13201, N7320);
buf BUF1 (N16303, N16291);
nor NOR4 (N16304, N16293, N16219, N1634, N13613);
xor XOR2 (N16305, N16294, N15953);
xor XOR2 (N16306, N16302, N558);
buf BUF1 (N16307, N16292);
buf BUF1 (N16308, N16298);
xor XOR2 (N16309, N16284, N15982);
buf BUF1 (N16310, N16308);
xor XOR2 (N16311, N16309, N5878);
nand NAND3 (N16312, N16306, N7602, N12235);
xor XOR2 (N16313, N16312, N7245);
nor NOR3 (N16314, N16300, N15884, N11190);
buf BUF1 (N16315, N16303);
not NOT1 (N16316, N16311);
nand NAND3 (N16317, N16304, N15345, N7347);
nor NOR4 (N16318, N16317, N4372, N4946, N1439);
nand NAND2 (N16319, N16305, N3457);
or OR3 (N16320, N16299, N11437, N15487);
not NOT1 (N16321, N16314);
nor NOR4 (N16322, N16321, N1573, N13995, N9975);
and AND4 (N16323, N16310, N2804, N8973, N7664);
nand NAND3 (N16324, N16322, N3316, N541);
not NOT1 (N16325, N16307);
nor NOR2 (N16326, N16316, N13434);
or OR2 (N16327, N16286, N5343);
not NOT1 (N16328, N16313);
and AND2 (N16329, N16319, N12962);
or OR4 (N16330, N16328, N2478, N4232, N8532);
buf BUF1 (N16331, N16315);
not NOT1 (N16332, N16329);
or OR3 (N16333, N16323, N13671, N16154);
buf BUF1 (N16334, N16320);
and AND2 (N16335, N16318, N5794);
not NOT1 (N16336, N16324);
and AND4 (N16337, N16326, N15811, N9919, N3108);
xor XOR2 (N16338, N16332, N15512);
or OR3 (N16339, N16335, N8061, N6659);
or OR4 (N16340, N16336, N3699, N7222, N12875);
and AND2 (N16341, N16327, N8005);
buf BUF1 (N16342, N16341);
nor NOR3 (N16343, N16333, N12078, N15537);
xor XOR2 (N16344, N16337, N13290);
xor XOR2 (N16345, N16342, N4909);
and AND3 (N16346, N16340, N12554, N15370);
buf BUF1 (N16347, N16344);
and AND3 (N16348, N16334, N8794, N350);
nor NOR3 (N16349, N16338, N3037, N14834);
and AND3 (N16350, N16349, N12854, N4389);
not NOT1 (N16351, N16345);
buf BUF1 (N16352, N16347);
nor NOR3 (N16353, N16346, N6693, N5543);
nand NAND4 (N16354, N16343, N11693, N10872, N9991);
or OR3 (N16355, N16339, N2575, N3422);
not NOT1 (N16356, N16355);
nand NAND2 (N16357, N16350, N15416);
not NOT1 (N16358, N16330);
and AND2 (N16359, N16354, N12517);
nor NOR2 (N16360, N16352, N2796);
xor XOR2 (N16361, N16351, N2462);
nand NAND2 (N16362, N16353, N5051);
and AND2 (N16363, N16325, N14376);
xor XOR2 (N16364, N16361, N9821);
or OR4 (N16365, N16360, N14759, N7439, N10877);
nor NOR4 (N16366, N16348, N4578, N1275, N13141);
not NOT1 (N16367, N16364);
and AND3 (N16368, N16331, N6624, N8247);
buf BUF1 (N16369, N16366);
and AND3 (N16370, N16358, N2888, N5447);
nand NAND4 (N16371, N16370, N8510, N4911, N6164);
and AND4 (N16372, N16362, N15941, N12688, N6540);
nand NAND3 (N16373, N16359, N14520, N12253);
nand NAND2 (N16374, N16357, N9446);
not NOT1 (N16375, N16363);
nor NOR2 (N16376, N16369, N11492);
nand NAND3 (N16377, N16372, N6131, N9068);
nand NAND4 (N16378, N16368, N13756, N16128, N15524);
buf BUF1 (N16379, N16377);
not NOT1 (N16380, N16373);
nand NAND3 (N16381, N16376, N9570, N3469);
not NOT1 (N16382, N16356);
xor XOR2 (N16383, N16380, N16025);
xor XOR2 (N16384, N16381, N69);
not NOT1 (N16385, N16382);
not NOT1 (N16386, N16385);
xor XOR2 (N16387, N16375, N15385);
and AND2 (N16388, N16367, N11624);
not NOT1 (N16389, N16378);
xor XOR2 (N16390, N16388, N1330);
xor XOR2 (N16391, N16379, N26);
nand NAND4 (N16392, N16365, N14936, N6547, N3261);
nand NAND4 (N16393, N16391, N13099, N12734, N5071);
nor NOR3 (N16394, N16393, N10835, N9328);
xor XOR2 (N16395, N16394, N4223);
xor XOR2 (N16396, N16383, N15297);
nor NOR3 (N16397, N16395, N13951, N10385);
nor NOR3 (N16398, N16392, N4941, N13815);
nor NOR3 (N16399, N16398, N8170, N9312);
nor NOR3 (N16400, N16399, N4143, N11202);
nand NAND3 (N16401, N16384, N7856, N12029);
nor NOR2 (N16402, N16374, N10953);
xor XOR2 (N16403, N16402, N3657);
or OR3 (N16404, N16387, N16301, N8191);
or OR3 (N16405, N16403, N15464, N6421);
nor NOR2 (N16406, N16401, N14170);
and AND2 (N16407, N16371, N2508);
and AND4 (N16408, N16396, N7700, N2296, N9976);
and AND4 (N16409, N16389, N4241, N6901, N10864);
and AND2 (N16410, N16409, N3819);
or OR2 (N16411, N16407, N8843);
and AND2 (N16412, N16400, N337);
not NOT1 (N16413, N16404);
xor XOR2 (N16414, N16405, N6324);
nand NAND2 (N16415, N16408, N14598);
xor XOR2 (N16416, N16390, N11435);
buf BUF1 (N16417, N16406);
nor NOR3 (N16418, N16411, N8939, N13217);
and AND2 (N16419, N16397, N6322);
nand NAND3 (N16420, N16415, N4041, N6843);
nor NOR3 (N16421, N16413, N1860, N13171);
buf BUF1 (N16422, N16421);
buf BUF1 (N16423, N16416);
buf BUF1 (N16424, N16419);
and AND3 (N16425, N16410, N7394, N4036);
not NOT1 (N16426, N16422);
and AND4 (N16427, N16424, N11170, N8858, N2651);
nor NOR4 (N16428, N16423, N10312, N8433, N5149);
and AND3 (N16429, N16428, N12322, N8746);
xor XOR2 (N16430, N16426, N1447);
buf BUF1 (N16431, N16418);
and AND4 (N16432, N16414, N11361, N12671, N6367);
buf BUF1 (N16433, N16420);
not NOT1 (N16434, N16429);
buf BUF1 (N16435, N16427);
nand NAND4 (N16436, N16430, N11691, N13657, N16029);
or OR2 (N16437, N16431, N11360);
xor XOR2 (N16438, N16425, N5016);
xor XOR2 (N16439, N16436, N1894);
nor NOR4 (N16440, N16433, N14466, N9959, N6266);
not NOT1 (N16441, N16435);
not NOT1 (N16442, N16438);
xor XOR2 (N16443, N16412, N293);
not NOT1 (N16444, N16437);
xor XOR2 (N16445, N16432, N9242);
and AND4 (N16446, N16444, N5893, N4390, N6216);
and AND2 (N16447, N16446, N12267);
buf BUF1 (N16448, N16440);
not NOT1 (N16449, N16417);
xor XOR2 (N16450, N16447, N55);
xor XOR2 (N16451, N16443, N9557);
nand NAND4 (N16452, N16445, N456, N5095, N1125);
nand NAND4 (N16453, N16434, N7533, N11383, N508);
buf BUF1 (N16454, N16439);
not NOT1 (N16455, N16449);
and AND4 (N16456, N16441, N5948, N4061, N12248);
nor NOR3 (N16457, N16456, N1072, N11052);
not NOT1 (N16458, N16442);
buf BUF1 (N16459, N16455);
and AND2 (N16460, N16386, N6702);
and AND2 (N16461, N16457, N12822);
not NOT1 (N16462, N16448);
buf BUF1 (N16463, N16450);
buf BUF1 (N16464, N16451);
nand NAND2 (N16465, N16452, N5512);
and AND4 (N16466, N16459, N5551, N13485, N16154);
or OR4 (N16467, N16466, N14288, N14663, N10585);
xor XOR2 (N16468, N16453, N1851);
or OR2 (N16469, N16463, N16082);
not NOT1 (N16470, N16469);
or OR3 (N16471, N16465, N10568, N9749);
nor NOR4 (N16472, N16461, N1785, N5943, N7629);
or OR4 (N16473, N16464, N8522, N3691, N15667);
xor XOR2 (N16474, N16472, N759);
buf BUF1 (N16475, N16473);
nand NAND4 (N16476, N16474, N4062, N1511, N2961);
or OR3 (N16477, N16470, N16370, N3057);
nand NAND4 (N16478, N16468, N10688, N5466, N8755);
not NOT1 (N16479, N16478);
or OR3 (N16480, N16476, N4074, N9114);
or OR4 (N16481, N16458, N929, N5769, N10517);
nor NOR3 (N16482, N16471, N3304, N16307);
nand NAND3 (N16483, N16462, N6723, N6311);
nand NAND2 (N16484, N16482, N11497);
nor NOR2 (N16485, N16467, N3844);
nand NAND4 (N16486, N16485, N1914, N14067, N9776);
xor XOR2 (N16487, N16480, N3247);
and AND4 (N16488, N16475, N14513, N5763, N4938);
nand NAND2 (N16489, N16483, N16028);
nand NAND4 (N16490, N16479, N16479, N7072, N8224);
nor NOR4 (N16491, N16486, N16046, N1220, N11807);
not NOT1 (N16492, N16489);
buf BUF1 (N16493, N16490);
buf BUF1 (N16494, N16492);
and AND3 (N16495, N16487, N2592, N4830);
xor XOR2 (N16496, N16477, N7659);
nor NOR4 (N16497, N16495, N14620, N1463, N3019);
and AND3 (N16498, N16460, N13425, N12317);
xor XOR2 (N16499, N16494, N6195);
not NOT1 (N16500, N16481);
nand NAND3 (N16501, N16499, N13710, N1138);
buf BUF1 (N16502, N16498);
buf BUF1 (N16503, N16500);
xor XOR2 (N16504, N16502, N8874);
not NOT1 (N16505, N16503);
xor XOR2 (N16506, N16496, N7693);
nand NAND3 (N16507, N16491, N13845, N14093);
xor XOR2 (N16508, N16484, N14330);
or OR3 (N16509, N16501, N9450, N11600);
buf BUF1 (N16510, N16505);
nor NOR4 (N16511, N16504, N3769, N14120, N14832);
not NOT1 (N16512, N16507);
not NOT1 (N16513, N16509);
nand NAND4 (N16514, N16506, N9608, N3097, N3361);
and AND3 (N16515, N16511, N221, N9699);
nor NOR4 (N16516, N16493, N4041, N46, N4332);
nand NAND3 (N16517, N16497, N10161, N14836);
nor NOR3 (N16518, N16508, N3466, N11705);
not NOT1 (N16519, N16514);
xor XOR2 (N16520, N16518, N8930);
nor NOR3 (N16521, N16515, N13403, N15046);
and AND2 (N16522, N16521, N6132);
nand NAND2 (N16523, N16516, N11476);
buf BUF1 (N16524, N16510);
or OR4 (N16525, N16512, N8983, N13431, N5470);
xor XOR2 (N16526, N16524, N3531);
not NOT1 (N16527, N16520);
and AND4 (N16528, N16527, N10005, N15767, N16321);
and AND3 (N16529, N16523, N4401, N3657);
buf BUF1 (N16530, N16454);
xor XOR2 (N16531, N16525, N12273);
and AND3 (N16532, N16513, N4384, N9963);
nand NAND3 (N16533, N16519, N8155, N12948);
nor NOR3 (N16534, N16522, N514, N9303);
nand NAND3 (N16535, N16517, N15581, N14415);
not NOT1 (N16536, N16532);
not NOT1 (N16537, N16529);
or OR2 (N16538, N16531, N14389);
not NOT1 (N16539, N16528);
nor NOR4 (N16540, N16488, N5749, N15193, N2162);
nand NAND3 (N16541, N16535, N3147, N4177);
nor NOR2 (N16542, N16536, N7668);
nand NAND4 (N16543, N16542, N12942, N10409, N6246);
and AND4 (N16544, N16530, N14904, N14619, N693);
buf BUF1 (N16545, N16537);
nor NOR4 (N16546, N16545, N15087, N16517, N10863);
and AND3 (N16547, N16543, N6651, N10265);
and AND2 (N16548, N16538, N15236);
and AND4 (N16549, N16539, N11925, N12831, N7527);
or OR2 (N16550, N16526, N8316);
not NOT1 (N16551, N16546);
xor XOR2 (N16552, N16548, N6436);
buf BUF1 (N16553, N16540);
buf BUF1 (N16554, N16534);
and AND3 (N16555, N16547, N10765, N11788);
not NOT1 (N16556, N16550);
nor NOR2 (N16557, N16552, N12843);
buf BUF1 (N16558, N16553);
nor NOR2 (N16559, N16541, N1054);
buf BUF1 (N16560, N16557);
nor NOR2 (N16561, N16560, N1812);
buf BUF1 (N16562, N16549);
nand NAND3 (N16563, N16544, N5478, N11503);
nor NOR4 (N16564, N16556, N11259, N2977, N4915);
nor NOR3 (N16565, N16555, N15409, N6851);
or OR2 (N16566, N16561, N8221);
nor NOR3 (N16567, N16565, N8334, N11387);
xor XOR2 (N16568, N16566, N5106);
xor XOR2 (N16569, N16559, N11680);
and AND2 (N16570, N16551, N9564);
and AND2 (N16571, N16562, N13351);
buf BUF1 (N16572, N16568);
or OR2 (N16573, N16563, N9221);
xor XOR2 (N16574, N16571, N1616);
nand NAND2 (N16575, N16574, N13914);
and AND3 (N16576, N16533, N11315, N3394);
xor XOR2 (N16577, N16576, N13944);
nand NAND3 (N16578, N16570, N11506, N12975);
nor NOR4 (N16579, N16554, N15298, N9636, N2929);
nand NAND3 (N16580, N16577, N15184, N13948);
xor XOR2 (N16581, N16580, N13207);
nor NOR4 (N16582, N16579, N15765, N13419, N9703);
or OR4 (N16583, N16582, N7700, N1757, N6165);
nand NAND4 (N16584, N16569, N8310, N14134, N1882);
xor XOR2 (N16585, N16584, N8695);
xor XOR2 (N16586, N16575, N10678);
buf BUF1 (N16587, N16558);
nand NAND4 (N16588, N16573, N10353, N4160, N3551);
xor XOR2 (N16589, N16564, N16578);
and AND3 (N16590, N15031, N14071, N7259);
xor XOR2 (N16591, N16587, N3575);
xor XOR2 (N16592, N16588, N1200);
xor XOR2 (N16593, N16567, N10265);
and AND3 (N16594, N16591, N9345, N16583);
nor NOR4 (N16595, N10248, N11770, N5743, N1036);
xor XOR2 (N16596, N16594, N10440);
buf BUF1 (N16597, N16585);
not NOT1 (N16598, N16593);
buf BUF1 (N16599, N16581);
buf BUF1 (N16600, N16590);
nand NAND2 (N16601, N16596, N6099);
or OR2 (N16602, N16595, N10299);
nand NAND3 (N16603, N16601, N9397, N4514);
or OR4 (N16604, N16586, N15823, N4245, N5512);
nand NAND2 (N16605, N16572, N4251);
nor NOR4 (N16606, N16599, N15770, N11782, N7534);
nand NAND2 (N16607, N16602, N9796);
xor XOR2 (N16608, N16589, N13306);
buf BUF1 (N16609, N16592);
nand NAND2 (N16610, N16609, N8222);
and AND4 (N16611, N16598, N155, N14462, N8384);
nand NAND4 (N16612, N16606, N9968, N3490, N11627);
xor XOR2 (N16613, N16610, N1942);
buf BUF1 (N16614, N16608);
nand NAND2 (N16615, N16604, N6285);
and AND2 (N16616, N16605, N2627);
buf BUF1 (N16617, N16600);
nor NOR2 (N16618, N16597, N6403);
nor NOR4 (N16619, N16607, N1477, N10991, N15238);
xor XOR2 (N16620, N16611, N1936);
nor NOR3 (N16621, N16615, N536, N6772);
not NOT1 (N16622, N16619);
not NOT1 (N16623, N16603);
and AND2 (N16624, N16621, N4093);
buf BUF1 (N16625, N16622);
buf BUF1 (N16626, N16624);
not NOT1 (N16627, N16614);
or OR2 (N16628, N16617, N4429);
nand NAND4 (N16629, N16620, N14270, N1350, N14033);
not NOT1 (N16630, N16616);
nand NAND2 (N16631, N16630, N1093);
xor XOR2 (N16632, N16628, N12614);
nor NOR3 (N16633, N16631, N8351, N8907);
not NOT1 (N16634, N16626);
or OR2 (N16635, N16625, N5135);
nand NAND2 (N16636, N16618, N11407);
and AND2 (N16637, N16632, N14007);
nand NAND2 (N16638, N16627, N10399);
nand NAND3 (N16639, N16613, N13621, N14440);
xor XOR2 (N16640, N16623, N14805);
nand NAND3 (N16641, N16633, N11438, N14387);
xor XOR2 (N16642, N16634, N12385);
buf BUF1 (N16643, N16636);
and AND2 (N16644, N16642, N12747);
xor XOR2 (N16645, N16639, N10225);
not NOT1 (N16646, N16638);
and AND4 (N16647, N16641, N11005, N8927, N7194);
and AND3 (N16648, N16635, N2770, N5062);
nor NOR4 (N16649, N16637, N1554, N4371, N6117);
not NOT1 (N16650, N16648);
or OR2 (N16651, N16646, N11745);
buf BUF1 (N16652, N16644);
buf BUF1 (N16653, N16649);
nor NOR3 (N16654, N16651, N788, N4013);
buf BUF1 (N16655, N16652);
nor NOR2 (N16656, N16653, N14336);
or OR4 (N16657, N16655, N9822, N6092, N12859);
not NOT1 (N16658, N16643);
xor XOR2 (N16659, N16657, N11373);
or OR2 (N16660, N16612, N6026);
nand NAND2 (N16661, N16650, N12586);
buf BUF1 (N16662, N16647);
xor XOR2 (N16663, N16645, N15977);
and AND2 (N16664, N16629, N2745);
or OR2 (N16665, N16656, N5055);
nand NAND3 (N16666, N16661, N3866, N6584);
buf BUF1 (N16667, N16640);
nor NOR4 (N16668, N16662, N12351, N4699, N9108);
and AND3 (N16669, N16664, N15422, N14735);
nand NAND2 (N16670, N16669, N3890);
nand NAND3 (N16671, N16670, N14941, N7110);
buf BUF1 (N16672, N16666);
or OR4 (N16673, N16668, N7392, N15373, N6261);
buf BUF1 (N16674, N16654);
xor XOR2 (N16675, N16667, N15052);
not NOT1 (N16676, N16671);
and AND3 (N16677, N16659, N4234, N10100);
and AND2 (N16678, N16677, N7018);
nand NAND3 (N16679, N16658, N15852, N1191);
buf BUF1 (N16680, N16674);
buf BUF1 (N16681, N16678);
nor NOR4 (N16682, N16676, N12298, N6754, N14248);
nor NOR2 (N16683, N16673, N6864);
or OR3 (N16684, N16683, N15527, N3115);
and AND4 (N16685, N16682, N8823, N9863, N14397);
nand NAND3 (N16686, N16679, N12896, N16553);
and AND2 (N16687, N16675, N6675);
buf BUF1 (N16688, N16686);
xor XOR2 (N16689, N16684, N7588);
not NOT1 (N16690, N16663);
or OR2 (N16691, N16690, N15778);
nand NAND2 (N16692, N16665, N8762);
nor NOR3 (N16693, N16692, N12421, N14918);
or OR2 (N16694, N16681, N12439);
buf BUF1 (N16695, N16693);
buf BUF1 (N16696, N16695);
not NOT1 (N16697, N16689);
nor NOR3 (N16698, N16685, N15834, N10172);
nand NAND2 (N16699, N16691, N4301);
not NOT1 (N16700, N16687);
or OR2 (N16701, N16696, N5358);
and AND3 (N16702, N16680, N16160, N11284);
not NOT1 (N16703, N16672);
and AND4 (N16704, N16660, N3561, N67, N10579);
and AND3 (N16705, N16702, N3693, N14622);
nor NOR3 (N16706, N16688, N6393, N16478);
nor NOR3 (N16707, N16701, N991, N16008);
and AND4 (N16708, N16700, N16586, N3811, N15152);
and AND2 (N16709, N16708, N2920);
not NOT1 (N16710, N16694);
not NOT1 (N16711, N16704);
not NOT1 (N16712, N16710);
not NOT1 (N16713, N16707);
and AND4 (N16714, N16705, N9148, N633, N13229);
and AND3 (N16715, N16699, N6934, N5810);
or OR2 (N16716, N16712, N987);
nand NAND3 (N16717, N16703, N3735, N8196);
not NOT1 (N16718, N16715);
nand NAND3 (N16719, N16717, N5044, N11339);
and AND4 (N16720, N16697, N2699, N1677, N12309);
buf BUF1 (N16721, N16711);
xor XOR2 (N16722, N16713, N898);
not NOT1 (N16723, N16720);
xor XOR2 (N16724, N16723, N13653);
nand NAND3 (N16725, N16716, N3144, N12);
buf BUF1 (N16726, N16725);
or OR3 (N16727, N16718, N13139, N15474);
nor NOR3 (N16728, N16719, N15589, N4974);
or OR2 (N16729, N16724, N12084);
xor XOR2 (N16730, N16729, N3165);
buf BUF1 (N16731, N16706);
xor XOR2 (N16732, N16730, N2800);
nor NOR3 (N16733, N16709, N10455, N1196);
buf BUF1 (N16734, N16727);
xor XOR2 (N16735, N16698, N6715);
or OR4 (N16736, N16722, N8702, N1036, N10574);
nor NOR4 (N16737, N16731, N14563, N1626, N416);
buf BUF1 (N16738, N16728);
xor XOR2 (N16739, N16737, N422);
xor XOR2 (N16740, N16738, N5346);
and AND2 (N16741, N16726, N16519);
not NOT1 (N16742, N16721);
xor XOR2 (N16743, N16736, N15742);
or OR3 (N16744, N16741, N8502, N10084);
buf BUF1 (N16745, N16740);
buf BUF1 (N16746, N16742);
nor NOR4 (N16747, N16733, N12509, N4044, N8378);
nor NOR2 (N16748, N16714, N14513);
xor XOR2 (N16749, N16735, N16405);
nor NOR3 (N16750, N16749, N6196, N934);
nor NOR4 (N16751, N16746, N5381, N6162, N12076);
xor XOR2 (N16752, N16745, N15995);
and AND4 (N16753, N16748, N1322, N2162, N15003);
buf BUF1 (N16754, N16739);
or OR4 (N16755, N16753, N222, N9412, N8104);
nand NAND2 (N16756, N16755, N3484);
xor XOR2 (N16757, N16732, N16340);
xor XOR2 (N16758, N16757, N2457);
not NOT1 (N16759, N16747);
and AND2 (N16760, N16751, N9701);
buf BUF1 (N16761, N16758);
not NOT1 (N16762, N16756);
not NOT1 (N16763, N16743);
nand NAND2 (N16764, N16754, N6910);
and AND2 (N16765, N16752, N1985);
nor NOR3 (N16766, N16750, N14586, N992);
and AND4 (N16767, N16761, N3636, N7160, N12321);
nor NOR2 (N16768, N16763, N4479);
nor NOR4 (N16769, N16734, N731, N11488, N13840);
and AND4 (N16770, N16762, N13287, N677, N13304);
and AND3 (N16771, N16770, N13649, N3606);
not NOT1 (N16772, N16765);
buf BUF1 (N16773, N16764);
or OR3 (N16774, N16771, N10797, N15109);
xor XOR2 (N16775, N16772, N4637);
and AND2 (N16776, N16768, N14129);
nand NAND4 (N16777, N16759, N1957, N11600, N13403);
not NOT1 (N16778, N16744);
xor XOR2 (N16779, N16775, N10770);
xor XOR2 (N16780, N16773, N4939);
not NOT1 (N16781, N16774);
not NOT1 (N16782, N16760);
buf BUF1 (N16783, N16777);
or OR2 (N16784, N16780, N15631);
buf BUF1 (N16785, N16778);
or OR4 (N16786, N16779, N11232, N2530, N7891);
xor XOR2 (N16787, N16769, N4277);
not NOT1 (N16788, N16786);
and AND2 (N16789, N16782, N13952);
nor NOR3 (N16790, N16766, N2534, N7616);
not NOT1 (N16791, N16781);
buf BUF1 (N16792, N16784);
buf BUF1 (N16793, N16789);
not NOT1 (N16794, N16792);
or OR2 (N16795, N16793, N7473);
buf BUF1 (N16796, N16776);
not NOT1 (N16797, N16787);
or OR2 (N16798, N16783, N3228);
nand NAND2 (N16799, N16796, N3310);
xor XOR2 (N16800, N16767, N5993);
nor NOR2 (N16801, N16799, N1366);
or OR3 (N16802, N16794, N7181, N11761);
not NOT1 (N16803, N16788);
nor NOR3 (N16804, N16803, N5120, N2759);
and AND4 (N16805, N16797, N13409, N3963, N15798);
nand NAND4 (N16806, N16785, N9122, N2231, N2178);
xor XOR2 (N16807, N16805, N13467);
xor XOR2 (N16808, N16798, N2392);
and AND2 (N16809, N16790, N877);
buf BUF1 (N16810, N16791);
or OR4 (N16811, N16802, N2102, N1639, N3266);
xor XOR2 (N16812, N16807, N15204);
not NOT1 (N16813, N16809);
nor NOR4 (N16814, N16801, N9673, N5578, N13972);
xor XOR2 (N16815, N16813, N12654);
and AND2 (N16816, N16800, N894);
buf BUF1 (N16817, N16795);
xor XOR2 (N16818, N16816, N16065);
or OR3 (N16819, N16804, N849, N13636);
nor NOR4 (N16820, N16814, N9212, N2873, N12392);
buf BUF1 (N16821, N16819);
not NOT1 (N16822, N16820);
xor XOR2 (N16823, N16808, N8934);
nor NOR3 (N16824, N16810, N8754, N10172);
and AND3 (N16825, N16817, N1890, N12058);
buf BUF1 (N16826, N16818);
not NOT1 (N16827, N16806);
buf BUF1 (N16828, N16821);
nor NOR4 (N16829, N16828, N9098, N3489, N16344);
not NOT1 (N16830, N16824);
xor XOR2 (N16831, N16827, N2911);
or OR4 (N16832, N16823, N9912, N7546, N10503);
xor XOR2 (N16833, N16830, N6191);
or OR3 (N16834, N16811, N5042, N9176);
nor NOR3 (N16835, N16833, N2880, N9124);
nor NOR4 (N16836, N16825, N10658, N8459, N7209);
xor XOR2 (N16837, N16834, N13210);
not NOT1 (N16838, N16829);
buf BUF1 (N16839, N16815);
buf BUF1 (N16840, N16838);
or OR3 (N16841, N16832, N10304, N1633);
and AND3 (N16842, N16840, N217, N5585);
xor XOR2 (N16843, N16841, N13057);
or OR2 (N16844, N16837, N11608);
or OR3 (N16845, N16839, N12372, N11240);
not NOT1 (N16846, N16812);
nor NOR3 (N16847, N16826, N5943, N4401);
and AND2 (N16848, N16836, N479);
nor NOR4 (N16849, N16844, N1199, N14294, N1249);
xor XOR2 (N16850, N16847, N4008);
xor XOR2 (N16851, N16850, N12341);
xor XOR2 (N16852, N16846, N15255);
and AND3 (N16853, N16851, N12313, N7852);
nand NAND2 (N16854, N16852, N16710);
or OR3 (N16855, N16835, N15086, N9641);
nor NOR4 (N16856, N16854, N1409, N7036, N7801);
and AND4 (N16857, N16845, N9862, N15205, N9101);
buf BUF1 (N16858, N16857);
or OR2 (N16859, N16849, N8293);
xor XOR2 (N16860, N16858, N9890);
not NOT1 (N16861, N16860);
nor NOR4 (N16862, N16843, N13622, N3191, N5504);
or OR3 (N16863, N16855, N12740, N214);
nand NAND3 (N16864, N16861, N14682, N2288);
nand NAND2 (N16865, N16863, N14982);
and AND2 (N16866, N16853, N15158);
nand NAND2 (N16867, N16866, N3506);
or OR2 (N16868, N16867, N4846);
or OR3 (N16869, N16864, N5224, N7792);
not NOT1 (N16870, N16842);
not NOT1 (N16871, N16848);
nand NAND3 (N16872, N16865, N6563, N3402);
or OR4 (N16873, N16872, N14961, N4960, N1316);
nor NOR3 (N16874, N16868, N5751, N7093);
nand NAND3 (N16875, N16871, N3055, N13769);
or OR2 (N16876, N16859, N1740);
buf BUF1 (N16877, N16831);
nand NAND3 (N16878, N16822, N10802, N14323);
nor NOR2 (N16879, N16873, N14948);
buf BUF1 (N16880, N16877);
buf BUF1 (N16881, N16876);
xor XOR2 (N16882, N16880, N6514);
nor NOR4 (N16883, N16881, N8472, N12676, N6759);
and AND3 (N16884, N16874, N2824, N6706);
buf BUF1 (N16885, N16875);
nand NAND4 (N16886, N16869, N55, N3975, N11193);
not NOT1 (N16887, N16879);
nand NAND3 (N16888, N16884, N13984, N10809);
buf BUF1 (N16889, N16885);
nor NOR4 (N16890, N16889, N13215, N9524, N15729);
buf BUF1 (N16891, N16890);
xor XOR2 (N16892, N16882, N13784);
buf BUF1 (N16893, N16886);
nand NAND4 (N16894, N16892, N8948, N3965, N1469);
nand NAND2 (N16895, N16893, N4068);
nand NAND2 (N16896, N16856, N6997);
nand NAND4 (N16897, N16887, N13648, N13894, N6829);
xor XOR2 (N16898, N16894, N2670);
or OR4 (N16899, N16895, N7390, N4672, N2125);
xor XOR2 (N16900, N16870, N9772);
not NOT1 (N16901, N16891);
not NOT1 (N16902, N16901);
and AND3 (N16903, N16897, N6170, N16198);
xor XOR2 (N16904, N16883, N12064);
nor NOR3 (N16905, N16888, N15917, N1627);
nand NAND3 (N16906, N16905, N10995, N1327);
nand NAND4 (N16907, N16862, N15082, N7825, N11749);
nor NOR3 (N16908, N16907, N4919, N11395);
or OR3 (N16909, N16904, N7414, N1291);
and AND3 (N16910, N16896, N7070, N13965);
nor NOR4 (N16911, N16908, N4018, N9165, N8262);
buf BUF1 (N16912, N16900);
nor NOR2 (N16913, N16909, N5650);
buf BUF1 (N16914, N16912);
not NOT1 (N16915, N16913);
buf BUF1 (N16916, N16906);
nor NOR2 (N16917, N16898, N4114);
nand NAND4 (N16918, N16902, N14580, N4482, N9679);
not NOT1 (N16919, N16917);
or OR4 (N16920, N16915, N9102, N5755, N9335);
buf BUF1 (N16921, N16911);
buf BUF1 (N16922, N16921);
nor NOR2 (N16923, N16920, N9968);
buf BUF1 (N16924, N16916);
and AND3 (N16925, N16924, N15344, N6857);
not NOT1 (N16926, N16899);
nand NAND3 (N16927, N16878, N14581, N14107);
not NOT1 (N16928, N16918);
xor XOR2 (N16929, N16925, N5209);
xor XOR2 (N16930, N16903, N13575);
buf BUF1 (N16931, N16923);
or OR3 (N16932, N16914, N10078, N5545);
xor XOR2 (N16933, N16927, N712);
nor NOR2 (N16934, N16928, N2053);
buf BUF1 (N16935, N16931);
nor NOR2 (N16936, N16922, N13784);
or OR2 (N16937, N16929, N2409);
or OR4 (N16938, N16926, N10255, N9683, N6865);
and AND3 (N16939, N16919, N11158, N14739);
and AND2 (N16940, N16933, N15373);
nand NAND3 (N16941, N16910, N4565, N12459);
nand NAND2 (N16942, N16934, N5340);
nand NAND3 (N16943, N16937, N15996, N8892);
and AND4 (N16944, N16940, N15985, N1486, N4141);
nand NAND4 (N16945, N16943, N11847, N16422, N14112);
nor NOR2 (N16946, N16935, N8970);
not NOT1 (N16947, N16939);
nor NOR3 (N16948, N16938, N13845, N11031);
or OR4 (N16949, N16946, N14487, N3667, N15579);
nand NAND2 (N16950, N16942, N4968);
nand NAND2 (N16951, N16949, N2181);
and AND2 (N16952, N16944, N206);
nand NAND2 (N16953, N16950, N8681);
buf BUF1 (N16954, N16941);
nor NOR4 (N16955, N16952, N15510, N10757, N4568);
nor NOR4 (N16956, N16954, N14569, N8059, N680);
and AND3 (N16957, N16948, N15216, N1207);
and AND2 (N16958, N16945, N10765);
xor XOR2 (N16959, N16956, N11545);
nor NOR2 (N16960, N16930, N7789);
or OR3 (N16961, N16947, N3885, N5664);
buf BUF1 (N16962, N16957);
nand NAND2 (N16963, N16960, N4636);
xor XOR2 (N16964, N16955, N4392);
buf BUF1 (N16965, N16951);
xor XOR2 (N16966, N16961, N7306);
or OR2 (N16967, N16936, N16532);
nand NAND2 (N16968, N16953, N12051);
or OR3 (N16969, N16958, N13181, N16742);
or OR4 (N16970, N16969, N4950, N16701, N1935);
xor XOR2 (N16971, N16959, N11760);
nand NAND4 (N16972, N16963, N8269, N2456, N15465);
and AND3 (N16973, N16962, N1256, N8101);
buf BUF1 (N16974, N16970);
xor XOR2 (N16975, N16968, N13718);
xor XOR2 (N16976, N16975, N14404);
not NOT1 (N16977, N16976);
buf BUF1 (N16978, N16932);
and AND3 (N16979, N16964, N13357, N3317);
not NOT1 (N16980, N16971);
xor XOR2 (N16981, N16965, N4047);
buf BUF1 (N16982, N16979);
xor XOR2 (N16983, N16966, N2490);
and AND2 (N16984, N16983, N14411);
buf BUF1 (N16985, N16984);
xor XOR2 (N16986, N16985, N7039);
nand NAND4 (N16987, N16972, N16122, N6121, N13020);
buf BUF1 (N16988, N16978);
or OR3 (N16989, N16967, N5393, N4717);
or OR2 (N16990, N16989, N16901);
xor XOR2 (N16991, N16986, N4459);
and AND2 (N16992, N16977, N14946);
and AND2 (N16993, N16991, N1503);
or OR3 (N16994, N16973, N1149, N7527);
nor NOR4 (N16995, N16988, N4472, N10595, N2451);
and AND4 (N16996, N16995, N5166, N6687, N6278);
not NOT1 (N16997, N16993);
xor XOR2 (N16998, N16992, N2647);
nor NOR2 (N16999, N16982, N16884);
nand NAND2 (N17000, N16997, N11764);
xor XOR2 (N17001, N16981, N10998);
or OR4 (N17002, N16990, N15859, N16596, N9);
not NOT1 (N17003, N16996);
or OR4 (N17004, N16999, N7867, N5406, N833);
and AND2 (N17005, N16998, N5588);
and AND3 (N17006, N16980, N12215, N8936);
xor XOR2 (N17007, N17003, N269);
or OR2 (N17008, N17000, N13161);
xor XOR2 (N17009, N16974, N4765);
and AND4 (N17010, N17008, N2624, N12821, N10943);
nand NAND3 (N17011, N17009, N14596, N12067);
nand NAND4 (N17012, N16987, N12555, N1859, N10017);
nand NAND4 (N17013, N17002, N15757, N15627, N790);
or OR4 (N17014, N17010, N12513, N415, N10228);
nand NAND2 (N17015, N17007, N9187);
or OR4 (N17016, N17006, N184, N9606, N13763);
nand NAND3 (N17017, N17014, N337, N43);
and AND2 (N17018, N17016, N6890);
or OR2 (N17019, N17001, N14520);
and AND3 (N17020, N17005, N7861, N404);
nand NAND4 (N17021, N17019, N14885, N6077, N2491);
nand NAND4 (N17022, N17018, N8627, N14752, N16093);
not NOT1 (N17023, N17013);
xor XOR2 (N17024, N17022, N3376);
nor NOR4 (N17025, N17012, N15754, N8353, N3453);
xor XOR2 (N17026, N17025, N15813);
xor XOR2 (N17027, N17011, N1906);
nand NAND2 (N17028, N17021, N9031);
buf BUF1 (N17029, N17023);
and AND4 (N17030, N17020, N5490, N3571, N7677);
and AND3 (N17031, N17004, N5308, N7871);
xor XOR2 (N17032, N17028, N3545);
not NOT1 (N17033, N17024);
nand NAND4 (N17034, N17030, N6790, N3917, N14912);
or OR4 (N17035, N17029, N12313, N6205, N11552);
and AND2 (N17036, N17032, N14263);
buf BUF1 (N17037, N17035);
buf BUF1 (N17038, N17017);
and AND2 (N17039, N17015, N1606);
and AND2 (N17040, N17033, N13506);
nor NOR3 (N17041, N17037, N6775, N8350);
not NOT1 (N17042, N17026);
not NOT1 (N17043, N17036);
and AND2 (N17044, N17027, N14606);
buf BUF1 (N17045, N17040);
nand NAND4 (N17046, N17041, N6539, N15107, N13146);
or OR3 (N17047, N17046, N2195, N11154);
buf BUF1 (N17048, N17042);
buf BUF1 (N17049, N17038);
and AND2 (N17050, N17049, N13530);
buf BUF1 (N17051, N16994);
buf BUF1 (N17052, N17031);
xor XOR2 (N17053, N17044, N1078);
or OR3 (N17054, N17034, N453, N13716);
xor XOR2 (N17055, N17043, N2404);
nand NAND3 (N17056, N17054, N6142, N14080);
not NOT1 (N17057, N17051);
buf BUF1 (N17058, N17039);
xor XOR2 (N17059, N17048, N1072);
nand NAND2 (N17060, N17047, N13269);
nand NAND2 (N17061, N17053, N9217);
and AND4 (N17062, N17058, N14964, N11484, N3830);
or OR2 (N17063, N17056, N8857);
buf BUF1 (N17064, N17062);
or OR4 (N17065, N17059, N8046, N14843, N5243);
buf BUF1 (N17066, N17055);
or OR2 (N17067, N17045, N14278);
buf BUF1 (N17068, N17061);
xor XOR2 (N17069, N17057, N1333);
nor NOR4 (N17070, N17066, N15075, N9206, N15489);
xor XOR2 (N17071, N17060, N7057);
buf BUF1 (N17072, N17070);
xor XOR2 (N17073, N17052, N4800);
nor NOR2 (N17074, N17068, N14963);
and AND2 (N17075, N17067, N15075);
not NOT1 (N17076, N17050);
nor NOR4 (N17077, N17065, N6512, N3440, N9967);
xor XOR2 (N17078, N17071, N10552);
not NOT1 (N17079, N17069);
and AND2 (N17080, N17075, N15184);
xor XOR2 (N17081, N17080, N6700);
buf BUF1 (N17082, N17078);
not NOT1 (N17083, N17072);
not NOT1 (N17084, N17076);
nor NOR4 (N17085, N17083, N8634, N6692, N3942);
nor NOR2 (N17086, N17081, N14908);
and AND3 (N17087, N17073, N3184, N9754);
buf BUF1 (N17088, N17079);
nand NAND2 (N17089, N17084, N12666);
nand NAND2 (N17090, N17089, N5131);
not NOT1 (N17091, N17085);
or OR3 (N17092, N17091, N3386, N9993);
and AND4 (N17093, N17077, N2298, N9421, N15587);
nand NAND2 (N17094, N17074, N10885);
or OR4 (N17095, N17094, N11203, N12515, N8133);
buf BUF1 (N17096, N17088);
or OR4 (N17097, N17095, N16953, N10922, N12354);
or OR3 (N17098, N17086, N15959, N12749);
nand NAND3 (N17099, N17063, N9498, N869);
not NOT1 (N17100, N17099);
buf BUF1 (N17101, N17098);
not NOT1 (N17102, N17092);
buf BUF1 (N17103, N17082);
nor NOR2 (N17104, N17093, N16856);
not NOT1 (N17105, N17104);
or OR3 (N17106, N17105, N370, N16319);
not NOT1 (N17107, N17106);
or OR4 (N17108, N17064, N14997, N5619, N7378);
buf BUF1 (N17109, N17101);
nand NAND4 (N17110, N17100, N2638, N4648, N2948);
not NOT1 (N17111, N17110);
nand NAND3 (N17112, N17111, N10281, N640);
or OR4 (N17113, N17087, N14067, N3903, N5804);
xor XOR2 (N17114, N17090, N12218);
or OR3 (N17115, N17112, N9459, N4255);
not NOT1 (N17116, N17113);
nand NAND4 (N17117, N17102, N16577, N13540, N7253);
not NOT1 (N17118, N17096);
not NOT1 (N17119, N17108);
nand NAND3 (N17120, N17097, N3459, N855);
nand NAND2 (N17121, N17117, N12922);
and AND3 (N17122, N17119, N857, N9231);
nor NOR4 (N17123, N17109, N13440, N2981, N14185);
nand NAND4 (N17124, N17118, N14835, N12807, N8366);
nand NAND4 (N17125, N17123, N5691, N8353, N16657);
and AND3 (N17126, N17115, N9995, N9274);
and AND2 (N17127, N17126, N11671);
not NOT1 (N17128, N17116);
nand NAND4 (N17129, N17114, N5555, N1874, N6666);
nor NOR4 (N17130, N17124, N3587, N2706, N2448);
buf BUF1 (N17131, N17122);
nor NOR4 (N17132, N17128, N10051, N13986, N10329);
and AND4 (N17133, N17127, N12913, N6847, N16860);
xor XOR2 (N17134, N17120, N9896);
xor XOR2 (N17135, N17130, N1639);
and AND4 (N17136, N17103, N16052, N14, N7044);
xor XOR2 (N17137, N17129, N9418);
or OR4 (N17138, N17121, N4076, N15474, N2655);
nor NOR4 (N17139, N17125, N4603, N4401, N2678);
not NOT1 (N17140, N17137);
buf BUF1 (N17141, N17134);
nand NAND4 (N17142, N17141, N3597, N7264, N8691);
or OR2 (N17143, N17142, N14269);
buf BUF1 (N17144, N17131);
and AND2 (N17145, N17135, N3498);
xor XOR2 (N17146, N17133, N2061);
not NOT1 (N17147, N17146);
xor XOR2 (N17148, N17144, N413);
or OR4 (N17149, N17143, N6475, N10732, N11172);
buf BUF1 (N17150, N17136);
and AND4 (N17151, N17139, N7689, N14732, N10611);
nand NAND4 (N17152, N17150, N1871, N2413, N5884);
nor NOR2 (N17153, N17138, N14789);
or OR3 (N17154, N17148, N12428, N15911);
nor NOR4 (N17155, N17107, N14900, N8464, N7001);
buf BUF1 (N17156, N17155);
not NOT1 (N17157, N17152);
not NOT1 (N17158, N17156);
and AND3 (N17159, N17140, N13446, N1923);
or OR2 (N17160, N17153, N9655);
buf BUF1 (N17161, N17145);
or OR2 (N17162, N17147, N14681);
buf BUF1 (N17163, N17151);
nand NAND2 (N17164, N17162, N9061);
buf BUF1 (N17165, N17163);
not NOT1 (N17166, N17164);
nor NOR3 (N17167, N17159, N9855, N6840);
and AND3 (N17168, N17157, N1846, N4303);
and AND2 (N17169, N17165, N17067);
xor XOR2 (N17170, N17161, N5594);
and AND2 (N17171, N17132, N2922);
or OR2 (N17172, N17169, N2815);
and AND2 (N17173, N17168, N592);
xor XOR2 (N17174, N17170, N149);
nor NOR2 (N17175, N17174, N2866);
and AND3 (N17176, N17160, N3312, N11519);
xor XOR2 (N17177, N17166, N4581);
or OR2 (N17178, N17167, N7078);
xor XOR2 (N17179, N17171, N10895);
and AND3 (N17180, N17172, N11751, N6720);
or OR2 (N17181, N17176, N16651);
and AND2 (N17182, N17149, N15372);
nand NAND3 (N17183, N17158, N15172, N4911);
nand NAND4 (N17184, N17180, N10678, N3060, N7524);
not NOT1 (N17185, N17178);
nor NOR2 (N17186, N17177, N10133);
and AND2 (N17187, N17181, N2124);
not NOT1 (N17188, N17175);
or OR4 (N17189, N17183, N5423, N6959, N10046);
xor XOR2 (N17190, N17154, N790);
buf BUF1 (N17191, N17179);
and AND2 (N17192, N17182, N10764);
nor NOR2 (N17193, N17191, N5367);
nand NAND2 (N17194, N17173, N7825);
and AND2 (N17195, N17193, N2989);
nand NAND2 (N17196, N17184, N12467);
nand NAND2 (N17197, N17188, N1299);
not NOT1 (N17198, N17194);
and AND3 (N17199, N17185, N14534, N3892);
nor NOR2 (N17200, N17199, N5466);
or OR3 (N17201, N17189, N4456, N7029);
xor XOR2 (N17202, N17196, N2525);
not NOT1 (N17203, N17190);
xor XOR2 (N17204, N17201, N8805);
nand NAND4 (N17205, N17197, N7375, N16340, N5814);
nand NAND3 (N17206, N17195, N2005, N12870);
and AND3 (N17207, N17206, N3327, N13457);
or OR2 (N17208, N17202, N10707);
and AND3 (N17209, N17205, N9770, N1720);
xor XOR2 (N17210, N17204, N6794);
or OR3 (N17211, N17209, N9917, N15583);
and AND2 (N17212, N17187, N7528);
nor NOR2 (N17213, N17211, N7462);
buf BUF1 (N17214, N17198);
and AND3 (N17215, N17192, N15668, N2508);
nor NOR2 (N17216, N17214, N8443);
nor NOR3 (N17217, N17208, N13910, N7915);
and AND4 (N17218, N17186, N5650, N613, N8649);
not NOT1 (N17219, N17200);
and AND2 (N17220, N17203, N12499);
buf BUF1 (N17221, N17220);
nor NOR4 (N17222, N17216, N15243, N14957, N4830);
nand NAND2 (N17223, N17219, N7147);
buf BUF1 (N17224, N17215);
buf BUF1 (N17225, N17224);
buf BUF1 (N17226, N17210);
and AND3 (N17227, N17213, N12072, N15738);
and AND4 (N17228, N17207, N17045, N14056, N5813);
nand NAND4 (N17229, N17221, N9491, N10621, N2116);
nor NOR4 (N17230, N17212, N7523, N6146, N7749);
xor XOR2 (N17231, N17225, N308);
or OR4 (N17232, N17229, N13676, N1822, N6534);
or OR3 (N17233, N17230, N16074, N9718);
nor NOR2 (N17234, N17217, N2004);
and AND2 (N17235, N17223, N5311);
nor NOR3 (N17236, N17232, N14302, N5546);
buf BUF1 (N17237, N17228);
buf BUF1 (N17238, N17235);
not NOT1 (N17239, N17237);
or OR2 (N17240, N17233, N11460);
nand NAND2 (N17241, N17234, N13931);
buf BUF1 (N17242, N17239);
and AND3 (N17243, N17242, N15016, N11579);
or OR4 (N17244, N17222, N328, N14146, N16519);
and AND2 (N17245, N17218, N9720);
nor NOR2 (N17246, N17238, N3441);
and AND2 (N17247, N17227, N9312);
nor NOR2 (N17248, N17243, N12103);
nor NOR4 (N17249, N17248, N15897, N1707, N8723);
xor XOR2 (N17250, N17245, N6621);
nor NOR3 (N17251, N17226, N3907, N8072);
or OR2 (N17252, N17241, N5659);
buf BUF1 (N17253, N17231);
xor XOR2 (N17254, N17246, N10182);
and AND4 (N17255, N17249, N2123, N12743, N3390);
nor NOR2 (N17256, N17254, N9725);
nand NAND4 (N17257, N17256, N14012, N6923, N8228);
nor NOR3 (N17258, N17236, N13643, N14924);
buf BUF1 (N17259, N17244);
nor NOR2 (N17260, N17251, N2715);
or OR3 (N17261, N17247, N6958, N2522);
and AND3 (N17262, N17259, N7841, N6132);
or OR3 (N17263, N17261, N1046, N14161);
not NOT1 (N17264, N17257);
nand NAND3 (N17265, N17240, N1270, N1670);
nand NAND2 (N17266, N17263, N454);
or OR3 (N17267, N17262, N6365, N12800);
not NOT1 (N17268, N17266);
or OR4 (N17269, N17250, N13856, N5943, N2456);
or OR4 (N17270, N17255, N3382, N4182, N5494);
or OR3 (N17271, N17270, N12720, N9466);
not NOT1 (N17272, N17252);
nor NOR4 (N17273, N17264, N10584, N11224, N16559);
nor NOR2 (N17274, N17272, N12955);
xor XOR2 (N17275, N17269, N1589);
buf BUF1 (N17276, N17271);
buf BUF1 (N17277, N17268);
nand NAND4 (N17278, N17267, N10713, N13128, N13329);
or OR3 (N17279, N17278, N16026, N4503);
and AND2 (N17280, N17279, N10337);
nor NOR3 (N17281, N17276, N16451, N14421);
buf BUF1 (N17282, N17281);
nor NOR2 (N17283, N17253, N8311);
nand NAND4 (N17284, N17274, N7946, N12806, N5267);
not NOT1 (N17285, N17265);
buf BUF1 (N17286, N17258);
buf BUF1 (N17287, N17284);
nor NOR4 (N17288, N17280, N13104, N6732, N1515);
nor NOR3 (N17289, N17286, N4398, N11361);
nand NAND2 (N17290, N17273, N4488);
not NOT1 (N17291, N17285);
nand NAND3 (N17292, N17288, N14942, N15652);
buf BUF1 (N17293, N17291);
buf BUF1 (N17294, N17293);
not NOT1 (N17295, N17283);
buf BUF1 (N17296, N17282);
xor XOR2 (N17297, N17294, N3883);
buf BUF1 (N17298, N17295);
xor XOR2 (N17299, N17287, N6817);
xor XOR2 (N17300, N17260, N6942);
nor NOR3 (N17301, N17298, N7440, N5457);
buf BUF1 (N17302, N17300);
not NOT1 (N17303, N17297);
and AND3 (N17304, N17296, N7716, N2334);
or OR3 (N17305, N17302, N16944, N4879);
and AND4 (N17306, N17289, N16217, N9483, N7798);
xor XOR2 (N17307, N17277, N9783);
buf BUF1 (N17308, N17303);
nor NOR4 (N17309, N17299, N15924, N3819, N14837);
nand NAND3 (N17310, N17304, N14447, N8655);
or OR3 (N17311, N17275, N8742, N13912);
buf BUF1 (N17312, N17306);
nor NOR4 (N17313, N17308, N15988, N14533, N8712);
nor NOR3 (N17314, N17312, N1081, N1195);
or OR3 (N17315, N17313, N113, N16619);
or OR3 (N17316, N17307, N909, N107);
xor XOR2 (N17317, N17314, N14155);
buf BUF1 (N17318, N17290);
and AND4 (N17319, N17318, N4286, N4774, N1547);
nand NAND4 (N17320, N17311, N9608, N1025, N16587);
nor NOR3 (N17321, N17292, N14043, N16392);
buf BUF1 (N17322, N17315);
not NOT1 (N17323, N17301);
and AND2 (N17324, N17322, N2167);
not NOT1 (N17325, N17323);
and AND3 (N17326, N17310, N15461, N16614);
buf BUF1 (N17327, N17321);
and AND3 (N17328, N17317, N5281, N7745);
buf BUF1 (N17329, N17305);
and AND4 (N17330, N17326, N1322, N1704, N4926);
and AND4 (N17331, N17327, N3503, N7010, N11546);
not NOT1 (N17332, N17319);
not NOT1 (N17333, N17330);
nand NAND3 (N17334, N17333, N2227, N17030);
nand NAND3 (N17335, N17329, N2266, N16171);
nor NOR4 (N17336, N17309, N7882, N2898, N3114);
not NOT1 (N17337, N17335);
nor NOR2 (N17338, N17325, N6443);
nor NOR4 (N17339, N17337, N16919, N11809, N13561);
or OR2 (N17340, N17338, N2995);
not NOT1 (N17341, N17339);
and AND2 (N17342, N17332, N11695);
buf BUF1 (N17343, N17340);
nor NOR4 (N17344, N17331, N1058, N10614, N1707);
and AND2 (N17345, N17328, N7991);
or OR3 (N17346, N17336, N11707, N3579);
nor NOR3 (N17347, N17316, N1841, N13911);
nand NAND4 (N17348, N17344, N13839, N10905, N10122);
buf BUF1 (N17349, N17345);
and AND2 (N17350, N17348, N449);
nor NOR4 (N17351, N17320, N14548, N13504, N15170);
xor XOR2 (N17352, N17349, N14565);
xor XOR2 (N17353, N17352, N13666);
nand NAND3 (N17354, N17334, N10565, N1410);
nor NOR2 (N17355, N17343, N6695);
and AND2 (N17356, N17350, N14779);
buf BUF1 (N17357, N17346);
xor XOR2 (N17358, N17347, N8406);
nand NAND4 (N17359, N17356, N3830, N7035, N4427);
buf BUF1 (N17360, N17351);
and AND3 (N17361, N17342, N8282, N5991);
not NOT1 (N17362, N17361);
nor NOR4 (N17363, N17359, N4741, N8160, N15125);
nor NOR2 (N17364, N17341, N13600);
or OR2 (N17365, N17363, N11515);
not NOT1 (N17366, N17324);
xor XOR2 (N17367, N17357, N116);
nor NOR4 (N17368, N17367, N7308, N5487, N5078);
and AND4 (N17369, N17355, N15269, N6390, N6199);
nand NAND3 (N17370, N17354, N14576, N578);
not NOT1 (N17371, N17369);
not NOT1 (N17372, N17370);
not NOT1 (N17373, N17372);
nand NAND3 (N17374, N17371, N1711, N13599);
or OR2 (N17375, N17374, N12094);
and AND2 (N17376, N17358, N11813);
xor XOR2 (N17377, N17364, N519);
xor XOR2 (N17378, N17360, N15947);
not NOT1 (N17379, N17373);
not NOT1 (N17380, N17376);
buf BUF1 (N17381, N17379);
nor NOR4 (N17382, N17375, N15795, N16588, N12941);
nand NAND4 (N17383, N17382, N10724, N6578, N6913);
nor NOR3 (N17384, N17378, N8722, N5564);
not NOT1 (N17385, N17381);
or OR4 (N17386, N17362, N9345, N7957, N5410);
buf BUF1 (N17387, N17366);
nand NAND2 (N17388, N17377, N12198);
and AND4 (N17389, N17368, N6875, N8221, N6452);
or OR3 (N17390, N17384, N4424, N10731);
and AND4 (N17391, N17365, N5005, N3793, N14317);
and AND4 (N17392, N17391, N12815, N251, N16138);
buf BUF1 (N17393, N17380);
xor XOR2 (N17394, N17387, N9500);
buf BUF1 (N17395, N17390);
or OR3 (N17396, N17394, N16385, N13379);
not NOT1 (N17397, N17396);
or OR2 (N17398, N17353, N17320);
nand NAND4 (N17399, N17385, N11084, N823, N5629);
nor NOR4 (N17400, N17383, N9498, N6815, N11762);
xor XOR2 (N17401, N17388, N1346);
or OR2 (N17402, N17386, N2274);
nand NAND3 (N17403, N17392, N8060, N2060);
xor XOR2 (N17404, N17399, N7421);
not NOT1 (N17405, N17402);
not NOT1 (N17406, N17404);
buf BUF1 (N17407, N17401);
or OR4 (N17408, N17407, N10038, N5410, N11117);
xor XOR2 (N17409, N17405, N16226);
xor XOR2 (N17410, N17408, N1852);
not NOT1 (N17411, N17398);
nor NOR4 (N17412, N17395, N14564, N11886, N3611);
xor XOR2 (N17413, N17406, N10415);
xor XOR2 (N17414, N17411, N10859);
buf BUF1 (N17415, N17413);
and AND4 (N17416, N17415, N7600, N12109, N13965);
not NOT1 (N17417, N17400);
and AND2 (N17418, N17416, N3535);
xor XOR2 (N17419, N17412, N16004);
nor NOR4 (N17420, N17397, N9391, N315, N16785);
and AND4 (N17421, N17420, N10617, N9377, N15319);
buf BUF1 (N17422, N17419);
not NOT1 (N17423, N17418);
and AND2 (N17424, N17403, N17057);
or OR4 (N17425, N17417, N8733, N15845, N616);
not NOT1 (N17426, N17422);
nor NOR4 (N17427, N17426, N14901, N4609, N10421);
xor XOR2 (N17428, N17393, N15139);
xor XOR2 (N17429, N17424, N14572);
xor XOR2 (N17430, N17414, N15792);
nand NAND2 (N17431, N17430, N1208);
buf BUF1 (N17432, N17423);
xor XOR2 (N17433, N17429, N8333);
xor XOR2 (N17434, N17425, N4713);
nor NOR2 (N17435, N17427, N10420);
not NOT1 (N17436, N17434);
nand NAND2 (N17437, N17433, N13623);
and AND3 (N17438, N17435, N14483, N12224);
buf BUF1 (N17439, N17432);
and AND2 (N17440, N17439, N8853);
or OR3 (N17441, N17438, N11920, N14683);
or OR3 (N17442, N17440, N8833, N10531);
nor NOR3 (N17443, N17442, N13166, N6479);
xor XOR2 (N17444, N17436, N6424);
and AND4 (N17445, N17437, N4733, N16660, N5411);
buf BUF1 (N17446, N17445);
buf BUF1 (N17447, N17446);
and AND4 (N17448, N17443, N15441, N13624, N6578);
or OR2 (N17449, N17410, N8291);
and AND4 (N17450, N17428, N1060, N16716, N8922);
nand NAND3 (N17451, N17431, N16508, N11503);
buf BUF1 (N17452, N17389);
not NOT1 (N17453, N17449);
nor NOR4 (N17454, N17421, N6690, N4582, N10679);
nor NOR4 (N17455, N17453, N5242, N12297, N6138);
xor XOR2 (N17456, N17444, N16102);
or OR3 (N17457, N17448, N13163, N6920);
or OR2 (N17458, N17450, N3015);
or OR3 (N17459, N17409, N8605, N15258);
or OR4 (N17460, N17457, N17274, N10843, N9347);
not NOT1 (N17461, N17458);
or OR2 (N17462, N17459, N12068);
nor NOR4 (N17463, N17462, N7590, N14371, N3390);
or OR3 (N17464, N17455, N9968, N6489);
nand NAND3 (N17465, N17454, N14516, N8131);
or OR2 (N17466, N17456, N6275);
nor NOR3 (N17467, N17451, N5505, N5021);
or OR2 (N17468, N17452, N11814);
xor XOR2 (N17469, N17467, N12122);
buf BUF1 (N17470, N17465);
nand NAND4 (N17471, N17470, N11859, N2110, N7621);
nor NOR4 (N17472, N17447, N2981, N1835, N9817);
not NOT1 (N17473, N17460);
or OR2 (N17474, N17466, N12307);
or OR2 (N17475, N17474, N5173);
nand NAND2 (N17476, N17441, N6808);
or OR4 (N17477, N17464, N9439, N12447, N2159);
nor NOR2 (N17478, N17461, N1411);
not NOT1 (N17479, N17473);
and AND4 (N17480, N17463, N1124, N16342, N8123);
xor XOR2 (N17481, N17480, N2357);
xor XOR2 (N17482, N17468, N6556);
xor XOR2 (N17483, N17475, N13406);
or OR3 (N17484, N17483, N9660, N17207);
nor NOR2 (N17485, N17471, N4100);
nor NOR4 (N17486, N17472, N14296, N8485, N9933);
xor XOR2 (N17487, N17485, N11597);
not NOT1 (N17488, N17477);
xor XOR2 (N17489, N17488, N11101);
xor XOR2 (N17490, N17482, N8028);
buf BUF1 (N17491, N17469);
buf BUF1 (N17492, N17487);
nor NOR2 (N17493, N17481, N4206);
buf BUF1 (N17494, N17490);
and AND2 (N17495, N17489, N1054);
buf BUF1 (N17496, N17484);
not NOT1 (N17497, N17478);
or OR4 (N17498, N17496, N7119, N10815, N17066);
or OR3 (N17499, N17494, N14865, N13369);
not NOT1 (N17500, N17486);
nand NAND4 (N17501, N17476, N5492, N3253, N169);
xor XOR2 (N17502, N17498, N11300);
and AND3 (N17503, N17500, N3965, N9351);
xor XOR2 (N17504, N17495, N7926);
xor XOR2 (N17505, N17491, N10848);
not NOT1 (N17506, N17505);
xor XOR2 (N17507, N17501, N7004);
or OR3 (N17508, N17492, N5983, N675);
nor NOR2 (N17509, N17504, N6318);
buf BUF1 (N17510, N17507);
buf BUF1 (N17511, N17497);
xor XOR2 (N17512, N17493, N5800);
buf BUF1 (N17513, N17511);
not NOT1 (N17514, N17499);
not NOT1 (N17515, N17509);
and AND4 (N17516, N17508, N7410, N489, N4040);
not NOT1 (N17517, N17510);
or OR2 (N17518, N17513, N12911);
nand NAND4 (N17519, N17502, N2383, N11085, N6043);
buf BUF1 (N17520, N17506);
nor NOR2 (N17521, N17517, N7585);
not NOT1 (N17522, N17521);
nor NOR2 (N17523, N17522, N5607);
and AND3 (N17524, N17518, N12991, N10553);
and AND3 (N17525, N17512, N2465, N14220);
not NOT1 (N17526, N17515);
not NOT1 (N17527, N17524);
not NOT1 (N17528, N17514);
not NOT1 (N17529, N17528);
xor XOR2 (N17530, N17527, N12041);
and AND2 (N17531, N17503, N15685);
and AND2 (N17532, N17530, N13407);
not NOT1 (N17533, N17526);
xor XOR2 (N17534, N17531, N8214);
nor NOR3 (N17535, N17520, N13658, N14005);
xor XOR2 (N17536, N17535, N9627);
and AND2 (N17537, N17532, N10572);
or OR2 (N17538, N17533, N1615);
not NOT1 (N17539, N17534);
not NOT1 (N17540, N17536);
or OR4 (N17541, N17519, N16596, N669, N14712);
and AND3 (N17542, N17537, N14875, N11696);
buf BUF1 (N17543, N17529);
not NOT1 (N17544, N17525);
and AND4 (N17545, N17516, N9907, N5706, N8605);
nand NAND3 (N17546, N17540, N13684, N14623);
and AND3 (N17547, N17546, N3465, N7931);
and AND4 (N17548, N17523, N10642, N2235, N2947);
nand NAND2 (N17549, N17548, N10344);
and AND4 (N17550, N17541, N4687, N10858, N12295);
nor NOR2 (N17551, N17545, N7171);
not NOT1 (N17552, N17551);
not NOT1 (N17553, N17543);
xor XOR2 (N17554, N17547, N15768);
nand NAND3 (N17555, N17552, N7459, N8448);
nand NAND3 (N17556, N17549, N15730, N12027);
not NOT1 (N17557, N17553);
not NOT1 (N17558, N17539);
xor XOR2 (N17559, N17479, N5770);
nor NOR2 (N17560, N17559, N5239);
not NOT1 (N17561, N17556);
and AND3 (N17562, N17558, N4318, N3224);
nand NAND4 (N17563, N17562, N12151, N17039, N12923);
buf BUF1 (N17564, N17544);
nand NAND2 (N17565, N17563, N5382);
and AND3 (N17566, N17560, N1372, N5915);
not NOT1 (N17567, N17557);
buf BUF1 (N17568, N17538);
not NOT1 (N17569, N17564);
and AND2 (N17570, N17555, N14179);
buf BUF1 (N17571, N17568);
nand NAND2 (N17572, N17569, N12674);
buf BUF1 (N17573, N17566);
nand NAND4 (N17574, N17561, N2176, N14524, N16214);
not NOT1 (N17575, N17567);
and AND4 (N17576, N17574, N9012, N15475, N13077);
nand NAND2 (N17577, N17554, N8817);
nand NAND4 (N17578, N17550, N16386, N3786, N15805);
nor NOR2 (N17579, N17573, N12907);
not NOT1 (N17580, N17575);
or OR2 (N17581, N17580, N16266);
nor NOR3 (N17582, N17542, N3668, N11262);
and AND3 (N17583, N17581, N16581, N17519);
nor NOR2 (N17584, N17572, N8266);
nand NAND4 (N17585, N17578, N5425, N7912, N6283);
nand NAND4 (N17586, N17585, N6767, N13111, N6621);
and AND2 (N17587, N17579, N10306);
xor XOR2 (N17588, N17586, N4134);
and AND2 (N17589, N17582, N9930);
buf BUF1 (N17590, N17584);
nand NAND2 (N17591, N17587, N4303);
and AND4 (N17592, N17583, N7488, N12210, N14008);
or OR4 (N17593, N17570, N14298, N714, N11447);
and AND4 (N17594, N17591, N8848, N7639, N3488);
nor NOR4 (N17595, N17592, N7655, N3775, N5561);
and AND4 (N17596, N17577, N12725, N13457, N7739);
xor XOR2 (N17597, N17571, N9892);
buf BUF1 (N17598, N17565);
nor NOR4 (N17599, N17598, N6704, N8893, N4241);
or OR4 (N17600, N17599, N11834, N11539, N164);
nand NAND2 (N17601, N17588, N2526);
or OR2 (N17602, N17594, N12926);
buf BUF1 (N17603, N17600);
or OR2 (N17604, N17590, N15977);
nor NOR2 (N17605, N17601, N12965);
nor NOR4 (N17606, N17597, N12244, N13909, N3173);
buf BUF1 (N17607, N17605);
nand NAND3 (N17608, N17593, N10924, N2521);
or OR4 (N17609, N17606, N14770, N2647, N16461);
buf BUF1 (N17610, N17576);
or OR4 (N17611, N17602, N14079, N7657, N6458);
and AND4 (N17612, N17610, N8776, N290, N2578);
nor NOR4 (N17613, N17589, N17468, N13583, N9354);
or OR3 (N17614, N17613, N6490, N822);
or OR2 (N17615, N17595, N9676);
and AND3 (N17616, N17614, N2149, N7348);
buf BUF1 (N17617, N17609);
xor XOR2 (N17618, N17616, N12777);
or OR2 (N17619, N17618, N13685);
nor NOR4 (N17620, N17615, N3674, N2458, N3543);
buf BUF1 (N17621, N17620);
not NOT1 (N17622, N17603);
nor NOR2 (N17623, N17608, N9876);
not NOT1 (N17624, N17622);
buf BUF1 (N17625, N17617);
or OR3 (N17626, N17624, N12120, N2732);
nand NAND4 (N17627, N17626, N11974, N12209, N12531);
nand NAND2 (N17628, N17627, N103);
xor XOR2 (N17629, N17628, N5698);
not NOT1 (N17630, N17629);
buf BUF1 (N17631, N17607);
nor NOR3 (N17632, N17623, N12029, N9893);
buf BUF1 (N17633, N17596);
or OR3 (N17634, N17611, N10080, N9243);
or OR2 (N17635, N17634, N6418);
nand NAND3 (N17636, N17604, N9132, N6641);
nand NAND2 (N17637, N17619, N2998);
or OR3 (N17638, N17621, N12572, N2794);
nor NOR2 (N17639, N17630, N14159);
buf BUF1 (N17640, N17638);
not NOT1 (N17641, N17635);
not NOT1 (N17642, N17636);
or OR2 (N17643, N17612, N765);
nor NOR3 (N17644, N17642, N1714, N3970);
and AND3 (N17645, N17644, N152, N6715);
or OR2 (N17646, N17645, N14019);
and AND4 (N17647, N17646, N968, N12760, N12699);
and AND3 (N17648, N17641, N17379, N8344);
xor XOR2 (N17649, N17631, N9905);
buf BUF1 (N17650, N17648);
or OR2 (N17651, N17625, N2699);
or OR3 (N17652, N17647, N4033, N13860);
and AND2 (N17653, N17643, N4713);
xor XOR2 (N17654, N17640, N7586);
not NOT1 (N17655, N17637);
xor XOR2 (N17656, N17632, N1142);
or OR4 (N17657, N17656, N165, N16967, N15470);
buf BUF1 (N17658, N17652);
not NOT1 (N17659, N17639);
nand NAND3 (N17660, N17657, N9953, N16791);
or OR4 (N17661, N17660, N13380, N5519, N3885);
not NOT1 (N17662, N17653);
xor XOR2 (N17663, N17658, N7838);
and AND3 (N17664, N17663, N5002, N17416);
nor NOR4 (N17665, N17654, N12069, N16494, N15332);
xor XOR2 (N17666, N17661, N597);
buf BUF1 (N17667, N17664);
xor XOR2 (N17668, N17665, N11643);
nand NAND3 (N17669, N17659, N5613, N15243);
buf BUF1 (N17670, N17649);
or OR4 (N17671, N17655, N7785, N9479, N9466);
buf BUF1 (N17672, N17651);
nor NOR4 (N17673, N17667, N8643, N6903, N12472);
buf BUF1 (N17674, N17666);
nor NOR2 (N17675, N17673, N10420);
xor XOR2 (N17676, N17672, N10542);
and AND4 (N17677, N17633, N9025, N10905, N15528);
or OR2 (N17678, N17671, N9482);
buf BUF1 (N17679, N17677);
not NOT1 (N17680, N17679);
buf BUF1 (N17681, N17675);
nor NOR3 (N17682, N17669, N1766, N10667);
xor XOR2 (N17683, N17668, N9226);
buf BUF1 (N17684, N17674);
not NOT1 (N17685, N17650);
or OR2 (N17686, N17683, N9412);
nor NOR2 (N17687, N17685, N1635);
and AND4 (N17688, N17676, N375, N6956, N4781);
and AND2 (N17689, N17684, N3079);
buf BUF1 (N17690, N17681);
buf BUF1 (N17691, N17688);
or OR2 (N17692, N17686, N15553);
xor XOR2 (N17693, N17690, N7917);
nor NOR3 (N17694, N17692, N4526, N396);
not NOT1 (N17695, N17694);
and AND3 (N17696, N17691, N6864, N9410);
nand NAND4 (N17697, N17696, N14729, N12605, N12972);
or OR4 (N17698, N17687, N7724, N16550, N9502);
nor NOR2 (N17699, N17680, N14475);
nor NOR2 (N17700, N17678, N17606);
or OR4 (N17701, N17682, N1874, N5089, N10197);
xor XOR2 (N17702, N17699, N11248);
xor XOR2 (N17703, N17670, N6441);
or OR4 (N17704, N17700, N15748, N16335, N10052);
buf BUF1 (N17705, N17704);
nor NOR3 (N17706, N17693, N12346, N3876);
and AND3 (N17707, N17703, N15892, N10373);
buf BUF1 (N17708, N17707);
and AND4 (N17709, N17708, N7558, N8512, N8933);
and AND2 (N17710, N17662, N14002);
buf BUF1 (N17711, N17705);
nor NOR3 (N17712, N17689, N12763, N13463);
or OR3 (N17713, N17706, N11776, N16746);
xor XOR2 (N17714, N17711, N12070);
nor NOR4 (N17715, N17697, N7542, N12905, N15061);
xor XOR2 (N17716, N17702, N10518);
xor XOR2 (N17717, N17709, N6859);
xor XOR2 (N17718, N17716, N9759);
xor XOR2 (N17719, N17717, N11207);
buf BUF1 (N17720, N17695);
and AND2 (N17721, N17713, N17100);
and AND2 (N17722, N17712, N15277);
not NOT1 (N17723, N17722);
nor NOR2 (N17724, N17715, N11216);
nor NOR4 (N17725, N17710, N8464, N15557, N2368);
and AND2 (N17726, N17724, N16186);
and AND2 (N17727, N17701, N7299);
nor NOR3 (N17728, N17720, N560, N16372);
and AND3 (N17729, N17723, N11246, N9660);
xor XOR2 (N17730, N17714, N15030);
and AND3 (N17731, N17719, N9383, N8877);
nor NOR2 (N17732, N17698, N3605);
buf BUF1 (N17733, N17726);
and AND4 (N17734, N17730, N17696, N12046, N13564);
nand NAND3 (N17735, N17728, N4908, N1183);
buf BUF1 (N17736, N17725);
nor NOR4 (N17737, N17731, N5615, N17050, N4945);
buf BUF1 (N17738, N17721);
not NOT1 (N17739, N17718);
nand NAND4 (N17740, N17733, N12263, N896, N7844);
not NOT1 (N17741, N17740);
nand NAND2 (N17742, N17741, N13937);
buf BUF1 (N17743, N17739);
buf BUF1 (N17744, N17737);
xor XOR2 (N17745, N17736, N14353);
nor NOR4 (N17746, N17744, N9879, N10151, N17699);
nor NOR3 (N17747, N17742, N16955, N16255);
buf BUF1 (N17748, N17729);
not NOT1 (N17749, N17747);
and AND2 (N17750, N17727, N4477);
and AND3 (N17751, N17738, N3393, N13725);
xor XOR2 (N17752, N17745, N9411);
and AND2 (N17753, N17746, N3863);
xor XOR2 (N17754, N17732, N6665);
nor NOR4 (N17755, N17754, N13628, N5640, N16559);
nand NAND4 (N17756, N17753, N14498, N3216, N9269);
buf BUF1 (N17757, N17752);
or OR4 (N17758, N17756, N2499, N1816, N15833);
not NOT1 (N17759, N17750);
buf BUF1 (N17760, N17757);
xor XOR2 (N17761, N17760, N13788);
nor NOR4 (N17762, N17761, N6337, N5237, N13574);
buf BUF1 (N17763, N17743);
nand NAND3 (N17764, N17759, N9891, N3655);
nor NOR4 (N17765, N17764, N2186, N271, N4575);
or OR3 (N17766, N17763, N15597, N7992);
xor XOR2 (N17767, N17755, N527);
not NOT1 (N17768, N17762);
buf BUF1 (N17769, N17768);
and AND2 (N17770, N17766, N13649);
xor XOR2 (N17771, N17769, N2628);
buf BUF1 (N17772, N17748);
and AND2 (N17773, N17758, N5410);
nor NOR4 (N17774, N17765, N15510, N11482, N5537);
and AND4 (N17775, N17749, N4279, N13862, N7023);
buf BUF1 (N17776, N17767);
nand NAND3 (N17777, N17773, N9099, N7427);
and AND4 (N17778, N17776, N843, N10526, N12818);
buf BUF1 (N17779, N17771);
and AND4 (N17780, N17734, N10739, N6023, N1230);
xor XOR2 (N17781, N17751, N4419);
and AND4 (N17782, N17778, N16464, N4442, N4131);
buf BUF1 (N17783, N17777);
and AND3 (N17784, N17781, N13581, N12660);
nand NAND3 (N17785, N17779, N17343, N16345);
buf BUF1 (N17786, N17735);
not NOT1 (N17787, N17785);
xor XOR2 (N17788, N17783, N11114);
nor NOR4 (N17789, N17772, N11733, N4300, N4436);
not NOT1 (N17790, N17770);
and AND2 (N17791, N17786, N17302);
nand NAND3 (N17792, N17790, N14502, N8020);
not NOT1 (N17793, N17788);
buf BUF1 (N17794, N17793);
nor NOR2 (N17795, N17792, N12496);
xor XOR2 (N17796, N17782, N16298);
or OR4 (N17797, N17774, N5081, N1388, N10854);
nand NAND3 (N17798, N17791, N4195, N8665);
or OR2 (N17799, N17795, N13541);
or OR4 (N17800, N17799, N4921, N8424, N14002);
xor XOR2 (N17801, N17787, N17467);
and AND3 (N17802, N17794, N16724, N16567);
nor NOR3 (N17803, N17796, N12766, N1901);
xor XOR2 (N17804, N17798, N16670);
xor XOR2 (N17805, N17784, N5698);
buf BUF1 (N17806, N17802);
buf BUF1 (N17807, N17805);
nand NAND4 (N17808, N17800, N15296, N1073, N13725);
or OR3 (N17809, N17801, N13784, N156);
nand NAND3 (N17810, N17804, N11678, N8702);
not NOT1 (N17811, N17780);
buf BUF1 (N17812, N17806);
not NOT1 (N17813, N17789);
nor NOR3 (N17814, N17775, N17238, N6785);
nand NAND4 (N17815, N17807, N16371, N4985, N416);
xor XOR2 (N17816, N17811, N9744);
buf BUF1 (N17817, N17812);
and AND4 (N17818, N17809, N17582, N3909, N16336);
buf BUF1 (N17819, N17803);
or OR2 (N17820, N17819, N7381);
nand NAND4 (N17821, N17797, N5134, N10534, N10338);
buf BUF1 (N17822, N17813);
xor XOR2 (N17823, N17821, N4231);
buf BUF1 (N17824, N17822);
nand NAND4 (N17825, N17823, N8015, N15883, N15283);
not NOT1 (N17826, N17824);
and AND4 (N17827, N17814, N13725, N3143, N11710);
and AND3 (N17828, N17818, N10146, N14353);
not NOT1 (N17829, N17826);
not NOT1 (N17830, N17808);
nand NAND3 (N17831, N17828, N14736, N187);
or OR4 (N17832, N17817, N6291, N11489, N4607);
nand NAND2 (N17833, N17831, N5882);
not NOT1 (N17834, N17830);
buf BUF1 (N17835, N17829);
not NOT1 (N17836, N17816);
buf BUF1 (N17837, N17834);
and AND2 (N17838, N17833, N6030);
buf BUF1 (N17839, N17832);
buf BUF1 (N17840, N17815);
and AND3 (N17841, N17836, N11330, N13403);
and AND3 (N17842, N17841, N17557, N5655);
nor NOR4 (N17843, N17837, N5257, N9136, N282);
not NOT1 (N17844, N17835);
xor XOR2 (N17845, N17838, N5309);
or OR4 (N17846, N17827, N16238, N6913, N9784);
xor XOR2 (N17847, N17845, N15155);
buf BUF1 (N17848, N17820);
not NOT1 (N17849, N17843);
xor XOR2 (N17850, N17839, N13366);
and AND4 (N17851, N17850, N16099, N11693, N11830);
and AND4 (N17852, N17842, N13354, N10810, N3610);
and AND4 (N17853, N17852, N3411, N11832, N9831);
buf BUF1 (N17854, N17849);
xor XOR2 (N17855, N17840, N5866);
and AND2 (N17856, N17851, N80);
xor XOR2 (N17857, N17856, N11281);
not NOT1 (N17858, N17825);
buf BUF1 (N17859, N17853);
xor XOR2 (N17860, N17859, N8378);
xor XOR2 (N17861, N17847, N16918);
nor NOR4 (N17862, N17810, N384, N17584, N1735);
or OR4 (N17863, N17855, N4883, N12635, N5927);
or OR4 (N17864, N17861, N2974, N13367, N673);
not NOT1 (N17865, N17848);
nor NOR3 (N17866, N17854, N3978, N4556);
or OR3 (N17867, N17862, N14115, N14036);
xor XOR2 (N17868, N17858, N14009);
buf BUF1 (N17869, N17866);
or OR2 (N17870, N17864, N3007);
and AND2 (N17871, N17868, N16650);
or OR3 (N17872, N17844, N15264, N1689);
nor NOR3 (N17873, N17867, N14372, N12318);
not NOT1 (N17874, N17873);
and AND3 (N17875, N17860, N3217, N2447);
and AND4 (N17876, N17869, N5586, N17657, N10555);
buf BUF1 (N17877, N17865);
buf BUF1 (N17878, N17875);
nand NAND3 (N17879, N17863, N3370, N15104);
or OR2 (N17880, N17857, N159);
or OR4 (N17881, N17874, N8996, N168, N7632);
or OR4 (N17882, N17871, N6920, N10168, N6245);
and AND3 (N17883, N17877, N9227, N8592);
nand NAND4 (N17884, N17882, N7215, N11928, N8437);
buf BUF1 (N17885, N17870);
buf BUF1 (N17886, N17878);
xor XOR2 (N17887, N17885, N4607);
xor XOR2 (N17888, N17887, N17579);
and AND4 (N17889, N17880, N2003, N7502, N10223);
buf BUF1 (N17890, N17886);
not NOT1 (N17891, N17879);
buf BUF1 (N17892, N17876);
nand NAND3 (N17893, N17890, N5858, N5271);
nand NAND3 (N17894, N17846, N15904, N11997);
nand NAND3 (N17895, N17888, N2830, N15043);
buf BUF1 (N17896, N17891);
xor XOR2 (N17897, N17889, N9078);
not NOT1 (N17898, N17895);
or OR4 (N17899, N17894, N34, N5394, N17584);
and AND2 (N17900, N17881, N4701);
buf BUF1 (N17901, N17892);
nand NAND4 (N17902, N17897, N5356, N6556, N10770);
xor XOR2 (N17903, N17872, N3617);
xor XOR2 (N17904, N17900, N9597);
nor NOR3 (N17905, N17903, N5469, N4618);
nand NAND3 (N17906, N17896, N3887, N13330);
or OR4 (N17907, N17905, N9616, N11585, N1713);
and AND3 (N17908, N17904, N5826, N11138);
nor NOR2 (N17909, N17884, N10518);
xor XOR2 (N17910, N17908, N9474);
not NOT1 (N17911, N17899);
nand NAND4 (N17912, N17907, N1346, N10701, N11526);
or OR4 (N17913, N17909, N5942, N12820, N7558);
and AND2 (N17914, N17902, N15103);
not NOT1 (N17915, N17906);
nor NOR2 (N17916, N17901, N1159);
xor XOR2 (N17917, N17916, N2542);
or OR3 (N17918, N17883, N521, N1482);
xor XOR2 (N17919, N17917, N17414);
xor XOR2 (N17920, N17915, N15407);
or OR2 (N17921, N17911, N7504);
nand NAND2 (N17922, N17918, N2901);
not NOT1 (N17923, N17913);
or OR2 (N17924, N17893, N8561);
not NOT1 (N17925, N17921);
not NOT1 (N17926, N17920);
buf BUF1 (N17927, N17923);
not NOT1 (N17928, N17914);
buf BUF1 (N17929, N17924);
xor XOR2 (N17930, N17912, N8707);
or OR4 (N17931, N17919, N5473, N2743, N572);
nor NOR2 (N17932, N17926, N3567);
buf BUF1 (N17933, N17922);
and AND3 (N17934, N17930, N13590, N13974);
nor NOR2 (N17935, N17898, N7696);
and AND3 (N17936, N17925, N7418, N7890);
not NOT1 (N17937, N17935);
or OR2 (N17938, N17927, N3165);
buf BUF1 (N17939, N17931);
nor NOR2 (N17940, N17938, N13492);
or OR4 (N17941, N17940, N3850, N14080, N9574);
and AND4 (N17942, N17928, N7869, N9074, N17312);
and AND4 (N17943, N17942, N3621, N3597, N11344);
not NOT1 (N17944, N17933);
or OR2 (N17945, N17941, N7204);
xor XOR2 (N17946, N17939, N11803);
and AND4 (N17947, N17944, N15894, N3649, N8178);
nor NOR4 (N17948, N17937, N6927, N8875, N2507);
xor XOR2 (N17949, N17932, N9505);
and AND3 (N17950, N17936, N2471, N7474);
nand NAND4 (N17951, N17950, N19, N16607, N7741);
nand NAND2 (N17952, N17943, N3738);
nor NOR3 (N17953, N17934, N3382, N9200);
xor XOR2 (N17954, N17947, N5144);
or OR4 (N17955, N17954, N3983, N5446, N6013);
and AND2 (N17956, N17946, N17762);
and AND2 (N17957, N17951, N217);
buf BUF1 (N17958, N17955);
buf BUF1 (N17959, N17952);
nand NAND4 (N17960, N17959, N2092, N1870, N16604);
nor NOR4 (N17961, N17956, N123, N6069, N8719);
nor NOR3 (N17962, N17948, N3455, N13005);
not NOT1 (N17963, N17929);
buf BUF1 (N17964, N17958);
xor XOR2 (N17965, N17949, N8384);
and AND4 (N17966, N17945, N9489, N3933, N11679);
and AND3 (N17967, N17953, N13450, N4332);
nor NOR3 (N17968, N17960, N9017, N16484);
and AND3 (N17969, N17968, N12, N13770);
nand NAND3 (N17970, N17966, N7586, N84);
buf BUF1 (N17971, N17967);
and AND3 (N17972, N17964, N3884, N5448);
xor XOR2 (N17973, N17965, N10968);
or OR4 (N17974, N17971, N13824, N2389, N11752);
not NOT1 (N17975, N17972);
not NOT1 (N17976, N17962);
and AND3 (N17977, N17970, N17387, N810);
nand NAND2 (N17978, N17974, N1126);
buf BUF1 (N17979, N17978);
and AND2 (N17980, N17957, N6952);
xor XOR2 (N17981, N17910, N17964);
nand NAND4 (N17982, N17976, N3279, N13336, N16673);
nand NAND4 (N17983, N17979, N8454, N15085, N509);
not NOT1 (N17984, N17961);
xor XOR2 (N17985, N17973, N5733);
not NOT1 (N17986, N17985);
nand NAND2 (N17987, N17975, N13731);
buf BUF1 (N17988, N17982);
and AND2 (N17989, N17983, N14321);
xor XOR2 (N17990, N17984, N17348);
buf BUF1 (N17991, N17981);
or OR3 (N17992, N17990, N11499, N6244);
and AND4 (N17993, N17992, N3230, N5256, N2970);
nand NAND4 (N17994, N17989, N6706, N6336, N6934);
nand NAND2 (N17995, N17963, N7464);
buf BUF1 (N17996, N17988);
xor XOR2 (N17997, N17996, N14345);
nand NAND2 (N17998, N17995, N7498);
buf BUF1 (N17999, N17969);
and AND2 (N18000, N17997, N14466);
nor NOR3 (N18001, N17987, N17584, N5826);
not NOT1 (N18002, N17994);
nand NAND3 (N18003, N17986, N2238, N8777);
not NOT1 (N18004, N17993);
and AND2 (N18005, N18003, N1027);
xor XOR2 (N18006, N17991, N17296);
not NOT1 (N18007, N17999);
not NOT1 (N18008, N18007);
nor NOR4 (N18009, N18008, N2599, N5801, N14825);
or OR3 (N18010, N18005, N5910, N10527);
nor NOR2 (N18011, N17980, N6257);
nand NAND4 (N18012, N18004, N374, N14491, N13583);
or OR3 (N18013, N18011, N1901, N14456);
xor XOR2 (N18014, N18001, N3016);
nand NAND3 (N18015, N18012, N7999, N3444);
xor XOR2 (N18016, N18014, N5201);
or OR2 (N18017, N18006, N15385);
not NOT1 (N18018, N18002);
nand NAND3 (N18019, N18017, N15811, N9317);
xor XOR2 (N18020, N18015, N7765);
nand NAND2 (N18021, N17977, N6542);
or OR3 (N18022, N18018, N6520, N8140);
nor NOR4 (N18023, N18020, N9084, N4095, N17251);
xor XOR2 (N18024, N18009, N5542);
buf BUF1 (N18025, N18021);
and AND4 (N18026, N18000, N16773, N8227, N9031);
and AND2 (N18027, N18026, N3321);
xor XOR2 (N18028, N18023, N3979);
or OR4 (N18029, N17998, N15996, N13844, N16005);
xor XOR2 (N18030, N18028, N615);
or OR2 (N18031, N18022, N8682);
nor NOR2 (N18032, N18010, N14700);
and AND2 (N18033, N18013, N13257);
and AND4 (N18034, N18029, N10825, N8840, N13791);
or OR4 (N18035, N18027, N14595, N488, N15037);
and AND2 (N18036, N18033, N10599);
nand NAND4 (N18037, N18019, N6254, N7465, N15474);
and AND3 (N18038, N18030, N5537, N1071);
and AND2 (N18039, N18031, N10295);
not NOT1 (N18040, N18034);
or OR2 (N18041, N18036, N2331);
not NOT1 (N18042, N18032);
or OR2 (N18043, N18040, N7478);
or OR3 (N18044, N18016, N12784, N5782);
nand NAND3 (N18045, N18037, N3803, N12299);
buf BUF1 (N18046, N18041);
nand NAND3 (N18047, N18045, N4589, N3845);
or OR2 (N18048, N18044, N13208);
xor XOR2 (N18049, N18047, N9807);
nand NAND3 (N18050, N18049, N17569, N12545);
buf BUF1 (N18051, N18050);
nor NOR3 (N18052, N18043, N11821, N1081);
buf BUF1 (N18053, N18042);
nand NAND3 (N18054, N18024, N470, N1324);
xor XOR2 (N18055, N18038, N15545);
not NOT1 (N18056, N18054);
not NOT1 (N18057, N18053);
nand NAND4 (N18058, N18025, N7776, N5445, N5260);
buf BUF1 (N18059, N18048);
not NOT1 (N18060, N18058);
and AND2 (N18061, N18039, N3439);
nand NAND3 (N18062, N18055, N10398, N13449);
xor XOR2 (N18063, N18035, N17671);
nor NOR4 (N18064, N18056, N3043, N9783, N4707);
not NOT1 (N18065, N18063);
nor NOR2 (N18066, N18061, N4625);
xor XOR2 (N18067, N18062, N8736);
not NOT1 (N18068, N18052);
nand NAND4 (N18069, N18066, N10716, N12033, N6790);
or OR4 (N18070, N18064, N10297, N14633, N13604);
nor NOR2 (N18071, N18065, N14806);
or OR3 (N18072, N18057, N12308, N268);
and AND2 (N18073, N18060, N4152);
and AND2 (N18074, N18069, N8990);
nand NAND2 (N18075, N18046, N15103);
and AND3 (N18076, N18067, N9112, N9761);
nand NAND2 (N18077, N18073, N1662);
and AND2 (N18078, N18076, N6781);
and AND4 (N18079, N18059, N13571, N15663, N3917);
and AND4 (N18080, N18051, N4922, N11967, N634);
xor XOR2 (N18081, N18071, N10421);
nand NAND4 (N18082, N18079, N322, N6673, N12635);
or OR4 (N18083, N18068, N327, N8508, N1126);
and AND3 (N18084, N18074, N16815, N17643);
nand NAND3 (N18085, N18072, N13019, N5278);
and AND2 (N18086, N18077, N1053);
buf BUF1 (N18087, N18082);
not NOT1 (N18088, N18085);
buf BUF1 (N18089, N18080);
xor XOR2 (N18090, N18078, N11696);
buf BUF1 (N18091, N18081);
and AND3 (N18092, N18075, N14310, N14646);
buf BUF1 (N18093, N18087);
nand NAND4 (N18094, N18088, N8397, N12732, N4071);
nor NOR4 (N18095, N18090, N1814, N4308, N11140);
nor NOR2 (N18096, N18092, N12294);
and AND4 (N18097, N18095, N9628, N5222, N9142);
nand NAND4 (N18098, N18084, N6094, N5338, N3982);
nand NAND3 (N18099, N18089, N16534, N720);
not NOT1 (N18100, N18093);
xor XOR2 (N18101, N18091, N13387);
xor XOR2 (N18102, N18086, N12623);
buf BUF1 (N18103, N18094);
nand NAND4 (N18104, N18070, N12125, N8930, N768);
or OR3 (N18105, N18103, N2062, N13623);
not NOT1 (N18106, N18098);
xor XOR2 (N18107, N18105, N3795);
nand NAND3 (N18108, N18106, N17082, N3449);
not NOT1 (N18109, N18083);
buf BUF1 (N18110, N18102);
or OR4 (N18111, N18110, N5480, N9005, N12644);
or OR4 (N18112, N18109, N1957, N9389, N8852);
and AND4 (N18113, N18101, N7320, N16886, N10922);
nand NAND2 (N18114, N18111, N2135);
and AND4 (N18115, N18100, N11038, N6212, N1231);
buf BUF1 (N18116, N18099);
nor NOR4 (N18117, N18112, N14313, N15772, N2097);
buf BUF1 (N18118, N18113);
and AND4 (N18119, N18096, N1920, N8676, N3502);
xor XOR2 (N18120, N18104, N3936);
not NOT1 (N18121, N18120);
not NOT1 (N18122, N18107);
and AND4 (N18123, N18118, N2827, N16410, N2779);
nor NOR3 (N18124, N18115, N13386, N15329);
nor NOR3 (N18125, N18121, N6442, N4058);
xor XOR2 (N18126, N18125, N10418);
or OR3 (N18127, N18122, N5973, N2067);
nand NAND2 (N18128, N18097, N4009);
buf BUF1 (N18129, N18127);
xor XOR2 (N18130, N18116, N1749);
nor NOR4 (N18131, N18129, N12880, N16199, N11517);
xor XOR2 (N18132, N18123, N6784);
not NOT1 (N18133, N18131);
nand NAND2 (N18134, N18108, N8947);
and AND2 (N18135, N18119, N3416);
and AND4 (N18136, N18128, N10941, N2400, N16055);
or OR4 (N18137, N18117, N4491, N12250, N5401);
nor NOR2 (N18138, N18136, N4907);
xor XOR2 (N18139, N18132, N11408);
not NOT1 (N18140, N18114);
nor NOR3 (N18141, N18135, N387, N15218);
not NOT1 (N18142, N18137);
not NOT1 (N18143, N18142);
xor XOR2 (N18144, N18138, N13494);
or OR4 (N18145, N18124, N9066, N973, N13643);
nand NAND3 (N18146, N18145, N9862, N2870);
or OR2 (N18147, N18143, N7874);
not NOT1 (N18148, N18141);
xor XOR2 (N18149, N18139, N16526);
or OR2 (N18150, N18149, N15902);
buf BUF1 (N18151, N18133);
and AND4 (N18152, N18151, N16368, N17323, N11465);
nand NAND2 (N18153, N18130, N13385);
and AND2 (N18154, N18153, N13028);
not NOT1 (N18155, N18134);
or OR2 (N18156, N18155, N6456);
and AND3 (N18157, N18156, N16427, N1567);
or OR2 (N18158, N18144, N15465);
xor XOR2 (N18159, N18126, N12435);
not NOT1 (N18160, N18159);
and AND4 (N18161, N18146, N1772, N260, N9274);
buf BUF1 (N18162, N18147);
xor XOR2 (N18163, N18140, N17752);
not NOT1 (N18164, N18154);
buf BUF1 (N18165, N18163);
xor XOR2 (N18166, N18152, N8897);
nand NAND3 (N18167, N18157, N54, N11430);
xor XOR2 (N18168, N18150, N4779);
or OR3 (N18169, N18165, N12282, N15873);
or OR4 (N18170, N18169, N12517, N4985, N12687);
nand NAND2 (N18171, N18167, N10303);
and AND4 (N18172, N18162, N1303, N1941, N17601);
or OR4 (N18173, N18161, N8559, N6295, N14478);
and AND4 (N18174, N18168, N13693, N5607, N4074);
and AND2 (N18175, N18148, N17360);
not NOT1 (N18176, N18160);
nand NAND4 (N18177, N18176, N10452, N11622, N4299);
and AND3 (N18178, N18175, N2200, N11445);
xor XOR2 (N18179, N18172, N9322);
and AND4 (N18180, N18174, N9940, N3578, N16763);
not NOT1 (N18181, N18173);
and AND2 (N18182, N18181, N8604);
nor NOR2 (N18183, N18180, N2733);
buf BUF1 (N18184, N18170);
and AND4 (N18185, N18177, N6099, N10180, N8322);
xor XOR2 (N18186, N18183, N1641);
xor XOR2 (N18187, N18184, N7529);
xor XOR2 (N18188, N18166, N9109);
nand NAND2 (N18189, N18186, N10785);
or OR3 (N18190, N18187, N13149, N4499);
and AND4 (N18191, N18190, N17711, N7864, N7961);
nand NAND4 (N18192, N18164, N2523, N11408, N8875);
xor XOR2 (N18193, N18192, N15482);
nand NAND4 (N18194, N18178, N6765, N12274, N10348);
or OR4 (N18195, N18182, N9280, N4822, N10370);
or OR4 (N18196, N18179, N5607, N3926, N18186);
buf BUF1 (N18197, N18158);
nor NOR2 (N18198, N18191, N818);
not NOT1 (N18199, N18196);
nor NOR3 (N18200, N18171, N8471, N6791);
nor NOR3 (N18201, N18197, N1454, N11807);
xor XOR2 (N18202, N18185, N4733);
and AND4 (N18203, N18200, N15899, N15668, N2782);
xor XOR2 (N18204, N18194, N12545);
nor NOR4 (N18205, N18201, N16683, N814, N5255);
nand NAND2 (N18206, N18193, N5110);
not NOT1 (N18207, N18199);
nand NAND2 (N18208, N18195, N14145);
buf BUF1 (N18209, N18189);
xor XOR2 (N18210, N18205, N5232);
or OR3 (N18211, N18209, N17460, N8282);
or OR3 (N18212, N18206, N13541, N8422);
buf BUF1 (N18213, N18202);
not NOT1 (N18214, N18207);
or OR2 (N18215, N18198, N16824);
nand NAND3 (N18216, N18188, N3182, N6352);
nor NOR3 (N18217, N18211, N16189, N15727);
not NOT1 (N18218, N18217);
not NOT1 (N18219, N18203);
or OR4 (N18220, N18208, N3923, N10039, N3252);
nor NOR3 (N18221, N18220, N13537, N4169);
xor XOR2 (N18222, N18214, N2978);
xor XOR2 (N18223, N18219, N16312);
and AND3 (N18224, N18218, N9186, N7681);
xor XOR2 (N18225, N18224, N13743);
and AND2 (N18226, N18223, N1066);
and AND4 (N18227, N18204, N15426, N13932, N3986);
buf BUF1 (N18228, N18212);
not NOT1 (N18229, N18225);
or OR3 (N18230, N18226, N10838, N5430);
xor XOR2 (N18231, N18229, N4861);
and AND2 (N18232, N18221, N14038);
nor NOR4 (N18233, N18228, N17011, N10626, N14222);
buf BUF1 (N18234, N18216);
xor XOR2 (N18235, N18213, N17510);
or OR3 (N18236, N18222, N16919, N4374);
buf BUF1 (N18237, N18215);
nor NOR2 (N18238, N18230, N13054);
nand NAND2 (N18239, N18231, N2840);
not NOT1 (N18240, N18238);
not NOT1 (N18241, N18239);
buf BUF1 (N18242, N18241);
nand NAND4 (N18243, N18234, N12698, N13916, N4495);
and AND3 (N18244, N18237, N15781, N598);
not NOT1 (N18245, N18232);
buf BUF1 (N18246, N18242);
or OR2 (N18247, N18245, N10309);
and AND2 (N18248, N18236, N9865);
nand NAND3 (N18249, N18210, N17594, N10630);
nand NAND4 (N18250, N18249, N11978, N8029, N16008);
xor XOR2 (N18251, N18248, N1213);
buf BUF1 (N18252, N18251);
xor XOR2 (N18253, N18240, N5647);
xor XOR2 (N18254, N18250, N9988);
nor NOR2 (N18255, N18227, N12925);
not NOT1 (N18256, N18254);
nor NOR4 (N18257, N18247, N746, N10860, N12908);
xor XOR2 (N18258, N18233, N7159);
buf BUF1 (N18259, N18253);
and AND2 (N18260, N18235, N2629);
and AND2 (N18261, N18257, N5579);
nand NAND4 (N18262, N18258, N668, N3321, N15108);
nand NAND4 (N18263, N18259, N2971, N12962, N13939);
nand NAND3 (N18264, N18246, N4368, N12989);
buf BUF1 (N18265, N18256);
or OR3 (N18266, N18252, N14577, N6);
and AND4 (N18267, N18262, N4203, N11908, N15951);
nor NOR2 (N18268, N18260, N7126);
or OR3 (N18269, N18263, N2895, N11829);
nor NOR4 (N18270, N18261, N10707, N3531, N12251);
buf BUF1 (N18271, N18255);
and AND4 (N18272, N18268, N2079, N3052, N15129);
nor NOR2 (N18273, N18243, N10885);
or OR4 (N18274, N18266, N8023, N17877, N3662);
buf BUF1 (N18275, N18271);
nor NOR3 (N18276, N18265, N8103, N11738);
buf BUF1 (N18277, N18276);
nor NOR2 (N18278, N18272, N4659);
nor NOR4 (N18279, N18267, N7788, N4886, N3506);
and AND2 (N18280, N18279, N16904);
xor XOR2 (N18281, N18273, N2612);
and AND3 (N18282, N18281, N450, N12937);
not NOT1 (N18283, N18278);
nand NAND4 (N18284, N18277, N716, N13133, N16377);
xor XOR2 (N18285, N18275, N3160);
nor NOR2 (N18286, N18284, N1503);
not NOT1 (N18287, N18286);
and AND4 (N18288, N18280, N16526, N1967, N12416);
xor XOR2 (N18289, N18288, N6717);
buf BUF1 (N18290, N18289);
not NOT1 (N18291, N18285);
xor XOR2 (N18292, N18282, N18091);
not NOT1 (N18293, N18287);
xor XOR2 (N18294, N18291, N2501);
nand NAND2 (N18295, N18264, N3544);
xor XOR2 (N18296, N18244, N15397);
xor XOR2 (N18297, N18283, N12470);
buf BUF1 (N18298, N18297);
and AND3 (N18299, N18274, N12049, N3466);
and AND3 (N18300, N18296, N17173, N16001);
or OR4 (N18301, N18294, N7583, N2440, N9749);
not NOT1 (N18302, N18269);
nor NOR3 (N18303, N18302, N10102, N6310);
not NOT1 (N18304, N18290);
xor XOR2 (N18305, N18298, N18285);
and AND2 (N18306, N18299, N15219);
or OR2 (N18307, N18305, N17440);
and AND3 (N18308, N18292, N7418, N4523);
or OR2 (N18309, N18270, N11741);
buf BUF1 (N18310, N18301);
or OR4 (N18311, N18309, N8059, N4342, N17527);
xor XOR2 (N18312, N18307, N7463);
xor XOR2 (N18313, N18306, N5880);
and AND3 (N18314, N18295, N15801, N6613);
xor XOR2 (N18315, N18303, N14968);
and AND4 (N18316, N18313, N17953, N3986, N14851);
or OR4 (N18317, N18314, N6624, N14470, N2832);
not NOT1 (N18318, N18311);
not NOT1 (N18319, N18304);
nor NOR3 (N18320, N18319, N6739, N8350);
nor NOR4 (N18321, N18310, N9150, N17418, N2928);
or OR4 (N18322, N18300, N193, N12522, N16971);
xor XOR2 (N18323, N18317, N4138);
xor XOR2 (N18324, N18308, N9652);
buf BUF1 (N18325, N18293);
nand NAND3 (N18326, N18325, N15205, N17734);
nor NOR4 (N18327, N18320, N15537, N646, N2210);
nand NAND3 (N18328, N18312, N13058, N3006);
nand NAND4 (N18329, N18316, N8764, N7258, N8107);
and AND4 (N18330, N18329, N1341, N2351, N8081);
nand NAND3 (N18331, N18318, N2558, N17495);
and AND3 (N18332, N18323, N12049, N12445);
not NOT1 (N18333, N18331);
nor NOR4 (N18334, N18327, N15721, N5862, N15621);
or OR4 (N18335, N18324, N899, N11210, N13241);
nand NAND2 (N18336, N18332, N6561);
or OR2 (N18337, N18321, N542);
nand NAND2 (N18338, N18328, N2344);
nand NAND2 (N18339, N18336, N4513);
nand NAND2 (N18340, N18315, N17230);
xor XOR2 (N18341, N18338, N4884);
nor NOR2 (N18342, N18334, N13923);
buf BUF1 (N18343, N18330);
nor NOR4 (N18344, N18342, N12898, N11919, N1285);
buf BUF1 (N18345, N18344);
or OR2 (N18346, N18340, N6256);
not NOT1 (N18347, N18337);
nand NAND2 (N18348, N18345, N14687);
not NOT1 (N18349, N18343);
nor NOR3 (N18350, N18333, N4555, N82);
or OR3 (N18351, N18350, N353, N11237);
nand NAND4 (N18352, N18351, N14971, N7925, N9156);
nand NAND4 (N18353, N18346, N10722, N16195, N3626);
not NOT1 (N18354, N18335);
and AND2 (N18355, N18326, N12239);
xor XOR2 (N18356, N18347, N5059);
buf BUF1 (N18357, N18349);
nand NAND2 (N18358, N18357, N7244);
buf BUF1 (N18359, N18339);
buf BUF1 (N18360, N18322);
nand NAND4 (N18361, N18358, N5004, N11768, N7688);
nor NOR4 (N18362, N18341, N4616, N15421, N8326);
and AND3 (N18363, N18362, N7702, N15673);
not NOT1 (N18364, N18361);
nand NAND2 (N18365, N18355, N4857);
xor XOR2 (N18366, N18360, N1643);
nor NOR2 (N18367, N18364, N14504);
or OR2 (N18368, N18352, N4793);
or OR2 (N18369, N18353, N14254);
or OR2 (N18370, N18368, N15488);
and AND4 (N18371, N18370, N15207, N232, N890);
nor NOR3 (N18372, N18363, N8378, N1535);
nor NOR2 (N18373, N18348, N11601);
nor NOR4 (N18374, N18373, N9476, N10829, N10809);
and AND4 (N18375, N18369, N8034, N7976, N4197);
buf BUF1 (N18376, N18367);
nor NOR4 (N18377, N18374, N11852, N16137, N14276);
nor NOR2 (N18378, N18366, N9363);
or OR3 (N18379, N18371, N3840, N6110);
nor NOR4 (N18380, N18354, N5079, N14701, N12779);
or OR3 (N18381, N18376, N5485, N3020);
xor XOR2 (N18382, N18365, N12015);
and AND2 (N18383, N18375, N11181);
or OR3 (N18384, N18380, N7531, N17578);
or OR4 (N18385, N18377, N4187, N5153, N17617);
xor XOR2 (N18386, N18359, N5632);
nand NAND3 (N18387, N18379, N17907, N15906);
not NOT1 (N18388, N18385);
xor XOR2 (N18389, N18388, N15337);
buf BUF1 (N18390, N18383);
and AND2 (N18391, N18372, N8090);
nor NOR3 (N18392, N18378, N11995, N7189);
and AND3 (N18393, N18390, N7129, N15761);
buf BUF1 (N18394, N18384);
nand NAND4 (N18395, N18394, N895, N11139, N7755);
nand NAND4 (N18396, N18389, N4809, N4821, N7844);
nand NAND4 (N18397, N18396, N11804, N1386, N8483);
or OR4 (N18398, N18381, N12655, N16615, N18107);
buf BUF1 (N18399, N18393);
nand NAND3 (N18400, N18386, N6506, N3638);
nor NOR3 (N18401, N18398, N682, N8218);
xor XOR2 (N18402, N18401, N10712);
nor NOR3 (N18403, N18391, N5166, N87);
nor NOR2 (N18404, N18356, N5542);
and AND4 (N18405, N18399, N14328, N18272, N9243);
nand NAND4 (N18406, N18405, N17558, N577, N13270);
nor NOR4 (N18407, N18397, N9689, N11747, N16649);
not NOT1 (N18408, N18406);
or OR3 (N18409, N18382, N246, N7180);
and AND4 (N18410, N18402, N13483, N12368, N2693);
or OR2 (N18411, N18392, N4336);
xor XOR2 (N18412, N18395, N14998);
and AND2 (N18413, N18403, N3957);
nor NOR2 (N18414, N18412, N8898);
nor NOR3 (N18415, N18410, N2195, N15181);
not NOT1 (N18416, N18411);
or OR3 (N18417, N18404, N12674, N17487);
or OR4 (N18418, N18416, N4361, N468, N6681);
not NOT1 (N18419, N18414);
nor NOR3 (N18420, N18400, N15109, N9775);
or OR4 (N18421, N18415, N5505, N2852, N748);
buf BUF1 (N18422, N18419);
nor NOR2 (N18423, N18407, N15691);
buf BUF1 (N18424, N18418);
not NOT1 (N18425, N18422);
nand NAND2 (N18426, N18417, N828);
not NOT1 (N18427, N18426);
or OR4 (N18428, N18408, N8708, N8919, N14747);
buf BUF1 (N18429, N18421);
nor NOR3 (N18430, N18429, N16691, N13925);
and AND4 (N18431, N18387, N11641, N7761, N2928);
not NOT1 (N18432, N18413);
and AND2 (N18433, N18431, N3851);
xor XOR2 (N18434, N18428, N13966);
buf BUF1 (N18435, N18425);
buf BUF1 (N18436, N18427);
not NOT1 (N18437, N18409);
xor XOR2 (N18438, N18430, N2544);
not NOT1 (N18439, N18433);
nor NOR4 (N18440, N18436, N2011, N11739, N5441);
and AND2 (N18441, N18435, N15659);
or OR4 (N18442, N18420, N10079, N12526, N14071);
buf BUF1 (N18443, N18424);
or OR2 (N18444, N18440, N6550);
or OR2 (N18445, N18437, N13950);
nand NAND3 (N18446, N18423, N3977, N11603);
and AND2 (N18447, N18442, N7154);
nor NOR4 (N18448, N18447, N309, N6308, N13792);
buf BUF1 (N18449, N18443);
or OR2 (N18450, N18441, N10347);
nand NAND3 (N18451, N18450, N8775, N4938);
not NOT1 (N18452, N18434);
nand NAND3 (N18453, N18448, N4407, N3695);
or OR2 (N18454, N18446, N9593);
xor XOR2 (N18455, N18432, N1293);
xor XOR2 (N18456, N18445, N9063);
and AND4 (N18457, N18456, N15434, N11489, N13063);
or OR2 (N18458, N18451, N16371);
nand NAND3 (N18459, N18444, N9923, N4387);
or OR3 (N18460, N18458, N12999, N6518);
buf BUF1 (N18461, N18460);
buf BUF1 (N18462, N18438);
nor NOR3 (N18463, N18459, N16723, N11408);
and AND4 (N18464, N18455, N6519, N2675, N4510);
nand NAND2 (N18465, N18464, N280);
not NOT1 (N18466, N18457);
or OR2 (N18467, N18463, N2129);
or OR3 (N18468, N18465, N9685, N11127);
and AND3 (N18469, N18468, N15324, N11991);
nor NOR3 (N18470, N18462, N4607, N15897);
or OR2 (N18471, N18470, N10670);
buf BUF1 (N18472, N18449);
not NOT1 (N18473, N18439);
xor XOR2 (N18474, N18469, N17303);
xor XOR2 (N18475, N18453, N13063);
and AND2 (N18476, N18467, N8836);
nor NOR2 (N18477, N18454, N16214);
and AND2 (N18478, N18477, N5904);
nor NOR2 (N18479, N18478, N17408);
xor XOR2 (N18480, N18475, N3537);
xor XOR2 (N18481, N18473, N10079);
nor NOR2 (N18482, N18452, N9473);
buf BUF1 (N18483, N18479);
buf BUF1 (N18484, N18461);
buf BUF1 (N18485, N18484);
nor NOR3 (N18486, N18466, N8799, N16932);
not NOT1 (N18487, N18474);
not NOT1 (N18488, N18487);
xor XOR2 (N18489, N18485, N15369);
buf BUF1 (N18490, N18483);
not NOT1 (N18491, N18480);
and AND4 (N18492, N18482, N12180, N865, N14700);
and AND4 (N18493, N18490, N1727, N17070, N13865);
buf BUF1 (N18494, N18492);
nand NAND2 (N18495, N18476, N7831);
or OR4 (N18496, N18481, N18425, N6773, N15638);
xor XOR2 (N18497, N18493, N5979);
or OR2 (N18498, N18497, N5202);
or OR3 (N18499, N18489, N7904, N12686);
not NOT1 (N18500, N18472);
buf BUF1 (N18501, N18499);
nor NOR3 (N18502, N18491, N9596, N14890);
not NOT1 (N18503, N18495);
not NOT1 (N18504, N18501);
and AND4 (N18505, N18471, N11146, N13884, N5797);
nand NAND3 (N18506, N18486, N2046, N2761);
and AND2 (N18507, N18498, N14198);
nand NAND4 (N18508, N18494, N1140, N15737, N4200);
nor NOR2 (N18509, N18504, N527);
buf BUF1 (N18510, N18503);
xor XOR2 (N18511, N18507, N11728);
nand NAND4 (N18512, N18502, N10335, N13925, N16486);
nand NAND3 (N18513, N18509, N1803, N13332);
nor NOR4 (N18514, N18496, N13007, N17814, N13597);
buf BUF1 (N18515, N18505);
xor XOR2 (N18516, N18506, N12963);
or OR3 (N18517, N18500, N12053, N1588);
nand NAND3 (N18518, N18515, N5123, N15515);
xor XOR2 (N18519, N18508, N15098);
and AND3 (N18520, N18510, N13100, N11001);
nor NOR4 (N18521, N18516, N5003, N2850, N3125);
xor XOR2 (N18522, N18511, N7189);
xor XOR2 (N18523, N18513, N9773);
buf BUF1 (N18524, N18517);
nor NOR2 (N18525, N18519, N7550);
not NOT1 (N18526, N18524);
buf BUF1 (N18527, N18525);
not NOT1 (N18528, N18527);
or OR4 (N18529, N18521, N10359, N1907, N14164);
nor NOR3 (N18530, N18526, N6044, N4840);
nor NOR2 (N18531, N18522, N11611);
nand NAND4 (N18532, N18514, N9893, N3925, N16200);
xor XOR2 (N18533, N18528, N12275);
or OR2 (N18534, N18518, N15731);
buf BUF1 (N18535, N18532);
and AND2 (N18536, N18534, N253);
buf BUF1 (N18537, N18512);
or OR2 (N18538, N18536, N12913);
and AND4 (N18539, N18538, N12995, N17867, N968);
or OR2 (N18540, N18533, N7751);
nand NAND2 (N18541, N18537, N5186);
and AND4 (N18542, N18488, N13007, N4706, N6021);
nor NOR2 (N18543, N18542, N18471);
nand NAND4 (N18544, N18523, N4998, N3112, N6750);
buf BUF1 (N18545, N18535);
nor NOR2 (N18546, N18539, N7785);
nand NAND3 (N18547, N18544, N9244, N3050);
and AND2 (N18548, N18531, N16596);
buf BUF1 (N18549, N18548);
not NOT1 (N18550, N18549);
not NOT1 (N18551, N18540);
nand NAND4 (N18552, N18543, N12219, N17188, N7754);
nor NOR4 (N18553, N18545, N4573, N2973, N17405);
nand NAND4 (N18554, N18551, N14961, N6529, N2561);
or OR4 (N18555, N18550, N16399, N7004, N11021);
xor XOR2 (N18556, N18553, N8451);
and AND4 (N18557, N18520, N18496, N5323, N2631);
buf BUF1 (N18558, N18530);
or OR4 (N18559, N18552, N16554, N9116, N11745);
not NOT1 (N18560, N18559);
not NOT1 (N18561, N18557);
buf BUF1 (N18562, N18547);
and AND3 (N18563, N18560, N7872, N410);
nand NAND4 (N18564, N18556, N14321, N5611, N11552);
and AND3 (N18565, N18563, N5051, N16884);
xor XOR2 (N18566, N18541, N6437);
nor NOR3 (N18567, N18565, N8294, N16577);
buf BUF1 (N18568, N18561);
nor NOR2 (N18569, N18529, N13326);
nor NOR2 (N18570, N18568, N2985);
and AND2 (N18571, N18570, N14557);
or OR3 (N18572, N18564, N1514, N11238);
nand NAND2 (N18573, N18572, N9837);
or OR2 (N18574, N18573, N7281);
buf BUF1 (N18575, N18574);
xor XOR2 (N18576, N18555, N1878);
nand NAND3 (N18577, N18562, N10180, N12819);
nand NAND3 (N18578, N18575, N4366, N16146);
nand NAND4 (N18579, N18569, N17094, N7854, N534);
xor XOR2 (N18580, N18554, N7923);
or OR3 (N18581, N18577, N8826, N12348);
nor NOR4 (N18582, N18580, N8883, N11145, N1140);
nand NAND4 (N18583, N18578, N8614, N18128, N6528);
nand NAND2 (N18584, N18576, N11873);
buf BUF1 (N18585, N18583);
xor XOR2 (N18586, N18584, N5239);
buf BUF1 (N18587, N18567);
xor XOR2 (N18588, N18581, N10179);
and AND3 (N18589, N18582, N16844, N1288);
not NOT1 (N18590, N18587);
and AND2 (N18591, N18571, N7366);
xor XOR2 (N18592, N18589, N2770);
nor NOR4 (N18593, N18585, N17420, N12141, N11673);
nand NAND2 (N18594, N18546, N14473);
buf BUF1 (N18595, N18558);
nand NAND2 (N18596, N18591, N14698);
or OR4 (N18597, N18586, N14056, N6499, N7911);
nand NAND3 (N18598, N18593, N4430, N13776);
or OR2 (N18599, N18598, N16532);
nor NOR2 (N18600, N18595, N12074);
xor XOR2 (N18601, N18579, N18203);
buf BUF1 (N18602, N18601);
or OR2 (N18603, N18590, N1998);
nor NOR2 (N18604, N18592, N18134);
buf BUF1 (N18605, N18599);
xor XOR2 (N18606, N18603, N17909);
nor NOR4 (N18607, N18566, N9092, N12336, N3146);
xor XOR2 (N18608, N18594, N5853);
buf BUF1 (N18609, N18602);
nand NAND3 (N18610, N18607, N16949, N13919);
or OR3 (N18611, N18609, N13523, N15033);
nand NAND2 (N18612, N18605, N15028);
nand NAND3 (N18613, N18610, N1691, N760);
not NOT1 (N18614, N18596);
nand NAND4 (N18615, N18613, N14600, N12566, N16682);
and AND3 (N18616, N18604, N12999, N3582);
nor NOR3 (N18617, N18588, N13502, N5606);
not NOT1 (N18618, N18615);
nor NOR4 (N18619, N18597, N8276, N3886, N1474);
xor XOR2 (N18620, N18611, N8472);
nor NOR4 (N18621, N18614, N11100, N7035, N14286);
nand NAND4 (N18622, N18617, N10210, N11212, N516);
or OR3 (N18623, N18620, N11603, N7684);
nand NAND2 (N18624, N18600, N5491);
nand NAND4 (N18625, N18621, N3930, N7578, N2910);
or OR2 (N18626, N18612, N5308);
and AND3 (N18627, N18616, N16455, N17062);
buf BUF1 (N18628, N18626);
not NOT1 (N18629, N18627);
nor NOR3 (N18630, N18623, N1146, N3801);
buf BUF1 (N18631, N18608);
nand NAND2 (N18632, N18629, N1373);
not NOT1 (N18633, N18624);
not NOT1 (N18634, N18632);
or OR2 (N18635, N18625, N5356);
nand NAND3 (N18636, N18634, N5371, N16547);
nor NOR3 (N18637, N18628, N9582, N106);
or OR3 (N18638, N18631, N14322, N804);
nor NOR3 (N18639, N18633, N9781, N13522);
xor XOR2 (N18640, N18606, N7413);
or OR2 (N18641, N18619, N6470);
xor XOR2 (N18642, N18636, N8916);
buf BUF1 (N18643, N18638);
not NOT1 (N18644, N18640);
nand NAND3 (N18645, N18637, N18116, N9004);
not NOT1 (N18646, N18630);
xor XOR2 (N18647, N18645, N13788);
xor XOR2 (N18648, N18647, N4709);
nor NOR3 (N18649, N18618, N990, N8113);
nand NAND3 (N18650, N18648, N2908, N2262);
xor XOR2 (N18651, N18635, N4799);
or OR4 (N18652, N18651, N8745, N10135, N6348);
buf BUF1 (N18653, N18639);
nand NAND2 (N18654, N18650, N9547);
or OR2 (N18655, N18641, N13954);
not NOT1 (N18656, N18649);
nor NOR2 (N18657, N18656, N8098);
xor XOR2 (N18658, N18646, N17621);
xor XOR2 (N18659, N18655, N2660);
not NOT1 (N18660, N18643);
or OR2 (N18661, N18653, N24);
xor XOR2 (N18662, N18654, N5388);
and AND2 (N18663, N18661, N16876);
nand NAND4 (N18664, N18622, N6214, N14550, N6111);
not NOT1 (N18665, N18662);
nor NOR3 (N18666, N18658, N17861, N18048);
and AND4 (N18667, N18666, N18520, N3394, N14769);
buf BUF1 (N18668, N18665);
and AND2 (N18669, N18659, N6037);
nand NAND4 (N18670, N18644, N2122, N5591, N13781);
not NOT1 (N18671, N18660);
not NOT1 (N18672, N18652);
buf BUF1 (N18673, N18670);
not NOT1 (N18674, N18671);
buf BUF1 (N18675, N18674);
xor XOR2 (N18676, N18657, N7952);
nor NOR4 (N18677, N18673, N13993, N17161, N8335);
xor XOR2 (N18678, N18668, N11232);
nor NOR4 (N18679, N18675, N1270, N15155, N15737);
nor NOR2 (N18680, N18664, N13775);
or OR2 (N18681, N18669, N4150);
not NOT1 (N18682, N18642);
xor XOR2 (N18683, N18676, N17089);
nor NOR4 (N18684, N18678, N12699, N17467, N2728);
nand NAND3 (N18685, N18682, N4105, N11758);
nor NOR3 (N18686, N18684, N14038, N3901);
buf BUF1 (N18687, N18680);
not NOT1 (N18688, N18679);
or OR4 (N18689, N18672, N8066, N4059, N16317);
or OR2 (N18690, N18687, N520);
xor XOR2 (N18691, N18667, N4797);
xor XOR2 (N18692, N18691, N8541);
and AND3 (N18693, N18677, N5009, N4374);
buf BUF1 (N18694, N18685);
nor NOR3 (N18695, N18686, N15678, N6595);
nor NOR3 (N18696, N18689, N12558, N10599);
not NOT1 (N18697, N18690);
and AND4 (N18698, N18697, N14007, N1714, N2326);
or OR4 (N18699, N18693, N13537, N16624, N18636);
xor XOR2 (N18700, N18692, N5342);
and AND4 (N18701, N18683, N6914, N2818, N10288);
xor XOR2 (N18702, N18699, N3848);
nor NOR3 (N18703, N18681, N7246, N8512);
xor XOR2 (N18704, N18701, N11103);
and AND4 (N18705, N18694, N6927, N1014, N9549);
and AND2 (N18706, N18688, N4732);
buf BUF1 (N18707, N18700);
nand NAND2 (N18708, N18695, N13396);
not NOT1 (N18709, N18706);
and AND2 (N18710, N18704, N4206);
nor NOR4 (N18711, N18696, N9502, N9073, N9235);
nand NAND2 (N18712, N18707, N988);
buf BUF1 (N18713, N18709);
not NOT1 (N18714, N18703);
and AND3 (N18715, N18702, N6595, N11829);
xor XOR2 (N18716, N18713, N55);
or OR3 (N18717, N18712, N17555, N8078);
xor XOR2 (N18718, N18711, N10291);
xor XOR2 (N18719, N18708, N5697);
nor NOR2 (N18720, N18698, N3472);
buf BUF1 (N18721, N18715);
not NOT1 (N18722, N18718);
nor NOR2 (N18723, N18705, N7514);
and AND4 (N18724, N18723, N4726, N10783, N14534);
and AND3 (N18725, N18721, N16854, N17451);
and AND4 (N18726, N18714, N17747, N13390, N10848);
and AND2 (N18727, N18717, N7127);
nor NOR4 (N18728, N18726, N8929, N4701, N3953);
and AND2 (N18729, N18722, N10899);
nand NAND3 (N18730, N18720, N9727, N17951);
buf BUF1 (N18731, N18710);
xor XOR2 (N18732, N18731, N18566);
and AND2 (N18733, N18729, N5767);
nand NAND4 (N18734, N18716, N6991, N17628, N2978);
nand NAND3 (N18735, N18725, N7043, N2085);
not NOT1 (N18736, N18730);
or OR4 (N18737, N18732, N4013, N15343, N2544);
buf BUF1 (N18738, N18727);
nand NAND2 (N18739, N18737, N12890);
xor XOR2 (N18740, N18735, N7948);
not NOT1 (N18741, N18719);
not NOT1 (N18742, N18724);
not NOT1 (N18743, N18663);
buf BUF1 (N18744, N18743);
nor NOR2 (N18745, N18728, N7386);
nor NOR3 (N18746, N18742, N16477, N7712);
xor XOR2 (N18747, N18738, N17486);
buf BUF1 (N18748, N18747);
not NOT1 (N18749, N18736);
and AND2 (N18750, N18745, N15736);
nor NOR3 (N18751, N18733, N11351, N12654);
xor XOR2 (N18752, N18749, N3282);
nand NAND3 (N18753, N18740, N18333, N3826);
nand NAND3 (N18754, N18748, N18617, N15409);
xor XOR2 (N18755, N18752, N6767);
and AND4 (N18756, N18744, N9317, N747, N9467);
buf BUF1 (N18757, N18751);
and AND2 (N18758, N18741, N15991);
nand NAND4 (N18759, N18746, N3700, N5599, N18676);
nand NAND3 (N18760, N18756, N7804, N12449);
buf BUF1 (N18761, N18754);
nor NOR4 (N18762, N18734, N5335, N9495, N10207);
buf BUF1 (N18763, N18755);
not NOT1 (N18764, N18762);
or OR2 (N18765, N18764, N5553);
and AND4 (N18766, N18761, N14410, N13895, N13655);
and AND2 (N18767, N18739, N16091);
xor XOR2 (N18768, N18760, N5751);
not NOT1 (N18769, N18767);
buf BUF1 (N18770, N18759);
buf BUF1 (N18771, N18765);
and AND4 (N18772, N18753, N11053, N3966, N4870);
or OR4 (N18773, N18758, N7481, N14297, N13982);
and AND4 (N18774, N18750, N18374, N9957, N163);
nand NAND4 (N18775, N18763, N16346, N12121, N5351);
nand NAND2 (N18776, N18766, N14854);
nor NOR2 (N18777, N18770, N9015);
nand NAND2 (N18778, N18774, N10571);
xor XOR2 (N18779, N18775, N10034);
not NOT1 (N18780, N18779);
buf BUF1 (N18781, N18778);
and AND3 (N18782, N18768, N15443, N3958);
nand NAND3 (N18783, N18769, N4653, N10609);
buf BUF1 (N18784, N18783);
nand NAND4 (N18785, N18772, N8864, N17503, N15149);
not NOT1 (N18786, N18780);
nor NOR2 (N18787, N18784, N6931);
nor NOR3 (N18788, N18777, N10231, N1506);
buf BUF1 (N18789, N18788);
buf BUF1 (N18790, N18786);
not NOT1 (N18791, N18785);
nor NOR2 (N18792, N18757, N13103);
and AND4 (N18793, N18791, N8489, N17834, N14500);
or OR2 (N18794, N18771, N5283);
or OR4 (N18795, N18790, N16734, N18490, N1492);
not NOT1 (N18796, N18787);
not NOT1 (N18797, N18792);
nand NAND3 (N18798, N18773, N15180, N8752);
buf BUF1 (N18799, N18798);
and AND3 (N18800, N18799, N4344, N10967);
and AND2 (N18801, N18776, N17789);
not NOT1 (N18802, N18781);
not NOT1 (N18803, N18782);
nor NOR3 (N18804, N18794, N16807, N6783);
not NOT1 (N18805, N18802);
not NOT1 (N18806, N18805);
nand NAND4 (N18807, N18806, N37, N16314, N7546);
not NOT1 (N18808, N18801);
nor NOR4 (N18809, N18808, N1082, N8261, N9510);
buf BUF1 (N18810, N18803);
not NOT1 (N18811, N18809);
nor NOR2 (N18812, N18800, N15692);
nor NOR4 (N18813, N18807, N2151, N6620, N1679);
not NOT1 (N18814, N18811);
not NOT1 (N18815, N18797);
nand NAND4 (N18816, N18795, N1016, N6390, N4737);
and AND3 (N18817, N18814, N11774, N11309);
buf BUF1 (N18818, N18815);
nor NOR3 (N18819, N18789, N947, N6615);
and AND4 (N18820, N18819, N1871, N15121, N768);
nand NAND3 (N18821, N18817, N7428, N7389);
buf BUF1 (N18822, N18818);
or OR3 (N18823, N18813, N4775, N9240);
nand NAND4 (N18824, N18822, N12623, N1493, N8693);
nand NAND4 (N18825, N18793, N903, N796, N12538);
and AND2 (N18826, N18823, N9851);
or OR4 (N18827, N18810, N8789, N7869, N4133);
or OR2 (N18828, N18804, N9241);
nand NAND2 (N18829, N18826, N8714);
buf BUF1 (N18830, N18824);
nor NOR4 (N18831, N18812, N12476, N11244, N15786);
or OR4 (N18832, N18825, N3931, N15103, N14809);
nor NOR3 (N18833, N18830, N14075, N7910);
or OR3 (N18834, N18833, N337, N12606);
or OR4 (N18835, N18828, N18326, N4623, N7097);
not NOT1 (N18836, N18835);
or OR2 (N18837, N18796, N871);
nand NAND4 (N18838, N18836, N10589, N18361, N373);
nand NAND2 (N18839, N18829, N8691);
not NOT1 (N18840, N18820);
nor NOR4 (N18841, N18816, N9421, N12889, N14712);
nand NAND4 (N18842, N18841, N16353, N10798, N2894);
nor NOR2 (N18843, N18840, N1772);
nor NOR2 (N18844, N18838, N16922);
xor XOR2 (N18845, N18842, N2180);
or OR3 (N18846, N18843, N15919, N783);
buf BUF1 (N18847, N18844);
nand NAND3 (N18848, N18832, N14200, N15361);
or OR4 (N18849, N18834, N16892, N2832, N16525);
or OR2 (N18850, N18827, N7643);
not NOT1 (N18851, N18846);
buf BUF1 (N18852, N18850);
nor NOR2 (N18853, N18851, N5508);
nand NAND4 (N18854, N18845, N6255, N12923, N11304);
buf BUF1 (N18855, N18848);
buf BUF1 (N18856, N18852);
not NOT1 (N18857, N18853);
nor NOR2 (N18858, N18837, N8292);
nor NOR4 (N18859, N18849, N6158, N5919, N13293);
buf BUF1 (N18860, N18858);
nor NOR3 (N18861, N18855, N3522, N14087);
or OR3 (N18862, N18831, N4985, N6311);
nand NAND3 (N18863, N18821, N10086, N15505);
or OR3 (N18864, N18860, N2901, N459);
nand NAND4 (N18865, N18857, N4346, N3905, N11645);
or OR4 (N18866, N18847, N941, N4033, N7329);
or OR3 (N18867, N18859, N15481, N12298);
nor NOR2 (N18868, N18856, N180);
nand NAND2 (N18869, N18865, N10185);
or OR2 (N18870, N18839, N12515);
and AND3 (N18871, N18866, N15284, N12402);
and AND4 (N18872, N18868, N16797, N7888, N4362);
not NOT1 (N18873, N18871);
buf BUF1 (N18874, N18870);
buf BUF1 (N18875, N18862);
and AND2 (N18876, N18867, N1481);
and AND2 (N18877, N18872, N6155);
or OR3 (N18878, N18863, N7242, N15440);
or OR2 (N18879, N18874, N717);
nor NOR4 (N18880, N18879, N9451, N5036, N17047);
nor NOR2 (N18881, N18880, N9036);
buf BUF1 (N18882, N18877);
not NOT1 (N18883, N18861);
or OR4 (N18884, N18881, N2048, N3485, N17322);
nor NOR4 (N18885, N18873, N10059, N2265, N17971);
nand NAND4 (N18886, N18876, N6544, N2041, N7798);
buf BUF1 (N18887, N18882);
xor XOR2 (N18888, N18885, N3906);
nand NAND3 (N18889, N18883, N13700, N13040);
or OR2 (N18890, N18869, N7679);
xor XOR2 (N18891, N18886, N3333);
nor NOR2 (N18892, N18864, N4131);
nor NOR2 (N18893, N18884, N18236);
or OR2 (N18894, N18887, N6054);
nor NOR3 (N18895, N18875, N6406, N1288);
or OR4 (N18896, N18893, N2105, N5909, N8486);
nor NOR4 (N18897, N18890, N237, N9573, N11921);
not NOT1 (N18898, N18888);
nand NAND2 (N18899, N18894, N11173);
not NOT1 (N18900, N18898);
or OR2 (N18901, N18891, N14988);
or OR2 (N18902, N18897, N11700);
and AND2 (N18903, N18892, N13006);
not NOT1 (N18904, N18889);
buf BUF1 (N18905, N18904);
xor XOR2 (N18906, N18854, N12884);
or OR4 (N18907, N18901, N125, N9568, N4317);
or OR4 (N18908, N18895, N7093, N4611, N9087);
buf BUF1 (N18909, N18905);
nor NOR2 (N18910, N18878, N3709);
buf BUF1 (N18911, N18902);
and AND3 (N18912, N18906, N10566, N9048);
and AND2 (N18913, N18912, N12388);
not NOT1 (N18914, N18911);
xor XOR2 (N18915, N18913, N14695);
xor XOR2 (N18916, N18899, N2188);
not NOT1 (N18917, N18896);
nand NAND3 (N18918, N18907, N5881, N14633);
nand NAND4 (N18919, N18917, N16137, N15589, N16653);
and AND3 (N18920, N18910, N3163, N2320);
xor XOR2 (N18921, N18918, N16483);
not NOT1 (N18922, N18909);
nand NAND2 (N18923, N18920, N4540);
buf BUF1 (N18924, N18900);
not NOT1 (N18925, N18919);
buf BUF1 (N18926, N18922);
nand NAND2 (N18927, N18924, N4149);
or OR4 (N18928, N18921, N1169, N4106, N10725);
or OR2 (N18929, N18928, N10121);
not NOT1 (N18930, N18903);
not NOT1 (N18931, N18927);
xor XOR2 (N18932, N18925, N7292);
xor XOR2 (N18933, N18926, N11388);
nor NOR4 (N18934, N18914, N5175, N6574, N11912);
and AND2 (N18935, N18932, N4239);
or OR3 (N18936, N18934, N2811, N4444);
xor XOR2 (N18937, N18915, N10510);
nand NAND2 (N18938, N18908, N16744);
buf BUF1 (N18939, N18933);
buf BUF1 (N18940, N18939);
nand NAND2 (N18941, N18936, N4016);
and AND3 (N18942, N18935, N4512, N9870);
not NOT1 (N18943, N18930);
buf BUF1 (N18944, N18938);
not NOT1 (N18945, N18937);
nand NAND2 (N18946, N18931, N17133);
not NOT1 (N18947, N18943);
or OR4 (N18948, N18945, N12123, N9388, N12999);
xor XOR2 (N18949, N18947, N16280);
buf BUF1 (N18950, N18916);
not NOT1 (N18951, N18949);
and AND3 (N18952, N18944, N12385, N11400);
and AND3 (N18953, N18950, N11477, N10729);
not NOT1 (N18954, N18946);
and AND3 (N18955, N18940, N14677, N17695);
and AND4 (N18956, N18923, N9304, N153, N2717);
nor NOR4 (N18957, N18956, N14808, N16898, N2323);
nor NOR3 (N18958, N18954, N11830, N17442);
or OR2 (N18959, N18951, N17040);
nor NOR2 (N18960, N18955, N15760);
not NOT1 (N18961, N18941);
and AND3 (N18962, N18942, N10914, N16170);
and AND3 (N18963, N18960, N5178, N14701);
nor NOR2 (N18964, N18952, N14340);
buf BUF1 (N18965, N18957);
xor XOR2 (N18966, N18958, N2031);
buf BUF1 (N18967, N18961);
not NOT1 (N18968, N18967);
and AND4 (N18969, N18953, N5351, N8353, N11371);
and AND4 (N18970, N18959, N11517, N13179, N769);
and AND4 (N18971, N18968, N14093, N7000, N13550);
xor XOR2 (N18972, N18962, N16268);
buf BUF1 (N18973, N18948);
xor XOR2 (N18974, N18972, N4205);
or OR2 (N18975, N18965, N7220);
not NOT1 (N18976, N18963);
not NOT1 (N18977, N18964);
xor XOR2 (N18978, N18976, N15773);
and AND3 (N18979, N18929, N2373, N7598);
nor NOR2 (N18980, N18973, N10395);
nand NAND3 (N18981, N18979, N14836, N6953);
nor NOR4 (N18982, N18975, N18227, N9115, N124);
not NOT1 (N18983, N18966);
nor NOR4 (N18984, N18970, N6670, N9390, N16631);
and AND4 (N18985, N18980, N13435, N17567, N4170);
not NOT1 (N18986, N18983);
or OR4 (N18987, N18978, N3409, N9363, N4682);
nor NOR3 (N18988, N18974, N17000, N15709);
xor XOR2 (N18989, N18969, N18368);
nor NOR2 (N18990, N18981, N3970);
not NOT1 (N18991, N18988);
nand NAND2 (N18992, N18991, N9425);
not NOT1 (N18993, N18986);
xor XOR2 (N18994, N18990, N5879);
and AND4 (N18995, N18982, N14250, N5058, N9382);
buf BUF1 (N18996, N18992);
nor NOR4 (N18997, N18993, N8732, N3015, N13041);
or OR2 (N18998, N18989, N11275);
xor XOR2 (N18999, N18984, N10190);
or OR3 (N19000, N18995, N1073, N12004);
and AND3 (N19001, N18999, N3202, N10017);
not NOT1 (N19002, N18994);
or OR3 (N19003, N19002, N14352, N9776);
buf BUF1 (N19004, N19000);
or OR4 (N19005, N19001, N13003, N371, N7539);
xor XOR2 (N19006, N18985, N18521);
nand NAND2 (N19007, N18998, N2955);
and AND3 (N19008, N18971, N2694, N16001);
or OR2 (N19009, N18997, N6012);
xor XOR2 (N19010, N19003, N5278);
or OR4 (N19011, N18987, N7989, N7861, N5251);
nor NOR3 (N19012, N18996, N10199, N16226);
not NOT1 (N19013, N18977);
and AND2 (N19014, N19007, N12382);
and AND3 (N19015, N19014, N7629, N9309);
nor NOR2 (N19016, N19011, N15094);
not NOT1 (N19017, N19012);
xor XOR2 (N19018, N19005, N8652);
or OR2 (N19019, N19008, N14306);
and AND3 (N19020, N19010, N15983, N14616);
buf BUF1 (N19021, N19019);
not NOT1 (N19022, N19009);
xor XOR2 (N19023, N19018, N14882);
and AND3 (N19024, N19021, N2204, N7218);
nand NAND2 (N19025, N19015, N2337);
not NOT1 (N19026, N19006);
or OR3 (N19027, N19022, N1216, N15407);
nand NAND4 (N19028, N19020, N15078, N150, N17512);
nor NOR2 (N19029, N19025, N8861);
xor XOR2 (N19030, N19023, N16314);
nand NAND3 (N19031, N19017, N7696, N3013);
xor XOR2 (N19032, N19024, N11981);
and AND3 (N19033, N19030, N55, N1543);
or OR2 (N19034, N19026, N16181);
buf BUF1 (N19035, N19027);
buf BUF1 (N19036, N19035);
buf BUF1 (N19037, N19031);
nand NAND3 (N19038, N19029, N5349, N4778);
or OR4 (N19039, N19032, N5071, N11967, N7112);
xor XOR2 (N19040, N19028, N3973);
or OR4 (N19041, N19039, N4604, N7152, N5136);
nand NAND3 (N19042, N19037, N16144, N18234);
nor NOR2 (N19043, N19004, N13606);
not NOT1 (N19044, N19036);
not NOT1 (N19045, N19041);
and AND4 (N19046, N19016, N14881, N7107, N1733);
not NOT1 (N19047, N19034);
not NOT1 (N19048, N19038);
not NOT1 (N19049, N19044);
xor XOR2 (N19050, N19047, N18704);
nand NAND2 (N19051, N19046, N7730);
nor NOR3 (N19052, N19051, N7833, N14281);
nor NOR4 (N19053, N19043, N4090, N17821, N10128);
buf BUF1 (N19054, N19052);
and AND4 (N19055, N19050, N18365, N13083, N14010);
xor XOR2 (N19056, N19040, N5309);
buf BUF1 (N19057, N19053);
nor NOR2 (N19058, N19054, N16141);
buf BUF1 (N19059, N19048);
nor NOR3 (N19060, N19055, N7405, N5780);
not NOT1 (N19061, N19059);
not NOT1 (N19062, N19056);
nor NOR2 (N19063, N19045, N18194);
buf BUF1 (N19064, N19013);
buf BUF1 (N19065, N19057);
buf BUF1 (N19066, N19058);
not NOT1 (N19067, N19042);
xor XOR2 (N19068, N19067, N13600);
nand NAND4 (N19069, N19049, N9532, N15072, N1594);
nor NOR2 (N19070, N19066, N345);
or OR4 (N19071, N19061, N5045, N10464, N8668);
nand NAND4 (N19072, N19068, N5226, N9163, N721);
nand NAND3 (N19073, N19065, N7622, N5953);
or OR4 (N19074, N19064, N8504, N3472, N13664);
buf BUF1 (N19075, N19070);
not NOT1 (N19076, N19072);
buf BUF1 (N19077, N19074);
not NOT1 (N19078, N19071);
nand NAND4 (N19079, N19033, N9768, N18788, N5792);
nor NOR3 (N19080, N19062, N8081, N4002);
or OR3 (N19081, N19063, N10078, N12131);
not NOT1 (N19082, N19078);
and AND2 (N19083, N19060, N18179);
not NOT1 (N19084, N19069);
or OR4 (N19085, N19081, N11452, N13897, N10289);
xor XOR2 (N19086, N19077, N12997);
buf BUF1 (N19087, N19082);
not NOT1 (N19088, N19087);
nand NAND4 (N19089, N19076, N7148, N5132, N14139);
and AND4 (N19090, N19086, N12250, N11090, N7659);
buf BUF1 (N19091, N19079);
not NOT1 (N19092, N19085);
not NOT1 (N19093, N19092);
buf BUF1 (N19094, N19075);
and AND3 (N19095, N19073, N6557, N9526);
or OR2 (N19096, N19090, N11781);
buf BUF1 (N19097, N19096);
nand NAND3 (N19098, N19083, N18288, N17795);
not NOT1 (N19099, N19097);
not NOT1 (N19100, N19088);
nand NAND4 (N19101, N19095, N1649, N9582, N6728);
and AND3 (N19102, N19093, N12673, N11311);
not NOT1 (N19103, N19089);
nand NAND4 (N19104, N19103, N9360, N5417, N4780);
not NOT1 (N19105, N19091);
xor XOR2 (N19106, N19080, N17019);
xor XOR2 (N19107, N19101, N7121);
buf BUF1 (N19108, N19084);
and AND4 (N19109, N19107, N17162, N4448, N18731);
buf BUF1 (N19110, N19094);
or OR4 (N19111, N19109, N571, N12237, N17732);
not NOT1 (N19112, N19099);
not NOT1 (N19113, N19098);
and AND3 (N19114, N19112, N16550, N13605);
and AND2 (N19115, N19102, N4641);
nor NOR3 (N19116, N19114, N11914, N8222);
or OR2 (N19117, N19115, N17771);
nand NAND3 (N19118, N19105, N4563, N5658);
and AND4 (N19119, N19117, N1592, N18017, N15347);
buf BUF1 (N19120, N19113);
nand NAND3 (N19121, N19104, N10072, N17186);
not NOT1 (N19122, N19108);
xor XOR2 (N19123, N19100, N15369);
nor NOR2 (N19124, N19110, N13676);
nor NOR4 (N19125, N19106, N17957, N884, N5715);
not NOT1 (N19126, N19123);
xor XOR2 (N19127, N19125, N11620);
or OR4 (N19128, N19126, N17629, N1312, N4971);
xor XOR2 (N19129, N19111, N19040);
xor XOR2 (N19130, N19124, N7348);
buf BUF1 (N19131, N19119);
nand NAND2 (N19132, N19131, N14556);
nor NOR4 (N19133, N19120, N7135, N3213, N6988);
buf BUF1 (N19134, N19121);
or OR3 (N19135, N19132, N14229, N17020);
xor XOR2 (N19136, N19118, N140);
buf BUF1 (N19137, N19122);
not NOT1 (N19138, N19133);
nor NOR2 (N19139, N19127, N9146);
nor NOR4 (N19140, N19138, N14091, N9075, N14679);
nor NOR3 (N19141, N19116, N18320, N7744);
or OR4 (N19142, N19141, N3355, N3761, N7330);
and AND2 (N19143, N19136, N12321);
buf BUF1 (N19144, N19140);
and AND4 (N19145, N19134, N19064, N16643, N14722);
xor XOR2 (N19146, N19137, N4125);
and AND4 (N19147, N19144, N7772, N5098, N667);
or OR3 (N19148, N19128, N5424, N8705);
nand NAND4 (N19149, N19147, N12324, N6689, N2818);
nor NOR4 (N19150, N19149, N8010, N5975, N3746);
buf BUF1 (N19151, N19146);
nand NAND2 (N19152, N19129, N11606);
not NOT1 (N19153, N19151);
not NOT1 (N19154, N19139);
buf BUF1 (N19155, N19154);
or OR2 (N19156, N19153, N19140);
nand NAND4 (N19157, N19148, N8693, N7680, N766);
buf BUF1 (N19158, N19143);
xor XOR2 (N19159, N19130, N18954);
xor XOR2 (N19160, N19150, N18442);
and AND4 (N19161, N19156, N16046, N9948, N12584);
xor XOR2 (N19162, N19159, N7793);
and AND4 (N19163, N19142, N13081, N5675, N18183);
nand NAND4 (N19164, N19163, N9801, N9289, N12313);
nor NOR2 (N19165, N19161, N3389);
buf BUF1 (N19166, N19158);
xor XOR2 (N19167, N19155, N11406);
nand NAND2 (N19168, N19165, N9556);
buf BUF1 (N19169, N19167);
buf BUF1 (N19170, N19162);
xor XOR2 (N19171, N19145, N9715);
xor XOR2 (N19172, N19152, N12523);
buf BUF1 (N19173, N19160);
xor XOR2 (N19174, N19168, N6051);
nor NOR3 (N19175, N19170, N2485, N4586);
nor NOR2 (N19176, N19164, N7009);
and AND3 (N19177, N19171, N15924, N14984);
nor NOR4 (N19178, N19169, N19027, N16763, N17775);
xor XOR2 (N19179, N19174, N4940);
not NOT1 (N19180, N19178);
nand NAND2 (N19181, N19180, N18343);
xor XOR2 (N19182, N19135, N5375);
or OR2 (N19183, N19172, N4235);
and AND2 (N19184, N19181, N17877);
buf BUF1 (N19185, N19184);
not NOT1 (N19186, N19173);
xor XOR2 (N19187, N19185, N5668);
nor NOR2 (N19188, N19183, N10421);
and AND2 (N19189, N19157, N19056);
not NOT1 (N19190, N19166);
xor XOR2 (N19191, N19175, N296);
nand NAND2 (N19192, N19189, N9199);
buf BUF1 (N19193, N19190);
nand NAND2 (N19194, N19179, N13194);
or OR2 (N19195, N19187, N17907);
nand NAND3 (N19196, N19193, N5363, N11625);
and AND4 (N19197, N19191, N17439, N15291, N12128);
nand NAND3 (N19198, N19182, N16631, N17564);
and AND4 (N19199, N19188, N17291, N7338, N15389);
buf BUF1 (N19200, N19186);
xor XOR2 (N19201, N19194, N11756);
nor NOR2 (N19202, N19201, N9972);
nor NOR2 (N19203, N19176, N14549);
or OR2 (N19204, N19203, N11286);
and AND3 (N19205, N19196, N1811, N8658);
nor NOR2 (N19206, N19200, N8677);
and AND2 (N19207, N19204, N5020);
buf BUF1 (N19208, N19195);
buf BUF1 (N19209, N19208);
and AND3 (N19210, N19199, N8452, N18016);
not NOT1 (N19211, N19205);
and AND4 (N19212, N19207, N6625, N5481, N8057);
buf BUF1 (N19213, N19210);
or OR2 (N19214, N19212, N13351);
nor NOR2 (N19215, N19213, N15543);
or OR4 (N19216, N19214, N14164, N8756, N9069);
and AND3 (N19217, N19206, N11317, N15766);
xor XOR2 (N19218, N19217, N12447);
nand NAND2 (N19219, N19198, N4364);
buf BUF1 (N19220, N19218);
not NOT1 (N19221, N19216);
nand NAND2 (N19222, N19177, N15384);
xor XOR2 (N19223, N19211, N17184);
buf BUF1 (N19224, N19219);
xor XOR2 (N19225, N19220, N7658);
not NOT1 (N19226, N19202);
nand NAND4 (N19227, N19222, N15045, N16510, N3828);
or OR4 (N19228, N19227, N2610, N4043, N1828);
nor NOR3 (N19229, N19221, N4076, N9464);
nand NAND4 (N19230, N19225, N10978, N6948, N3147);
and AND4 (N19231, N19192, N6422, N1011, N17028);
not NOT1 (N19232, N19230);
buf BUF1 (N19233, N19215);
nor NOR3 (N19234, N19224, N9843, N9662);
nor NOR2 (N19235, N19232, N36);
xor XOR2 (N19236, N19228, N2130);
or OR4 (N19237, N19197, N17569, N11762, N8816);
and AND4 (N19238, N19235, N10236, N2886, N3209);
nor NOR3 (N19239, N19238, N10317, N7466);
nor NOR2 (N19240, N19233, N1849);
and AND3 (N19241, N19229, N5370, N15071);
not NOT1 (N19242, N19239);
not NOT1 (N19243, N19234);
buf BUF1 (N19244, N19209);
xor XOR2 (N19245, N19236, N11418);
and AND2 (N19246, N19244, N12600);
buf BUF1 (N19247, N19237);
xor XOR2 (N19248, N19242, N3272);
xor XOR2 (N19249, N19241, N5264);
nand NAND4 (N19250, N19231, N13762, N1697, N13365);
not NOT1 (N19251, N19226);
or OR4 (N19252, N19246, N16025, N10987, N1991);
nor NOR4 (N19253, N19243, N101, N6462, N13096);
nand NAND2 (N19254, N19247, N4643);
and AND4 (N19255, N19250, N18656, N2210, N17823);
nor NOR2 (N19256, N19249, N15950);
or OR2 (N19257, N19255, N4529);
xor XOR2 (N19258, N19248, N14487);
buf BUF1 (N19259, N19252);
nand NAND3 (N19260, N19259, N16049, N11160);
not NOT1 (N19261, N19223);
or OR4 (N19262, N19240, N8986, N6341, N8261);
xor XOR2 (N19263, N19254, N9009);
nand NAND4 (N19264, N19253, N17915, N11281, N15166);
xor XOR2 (N19265, N19263, N18024);
buf BUF1 (N19266, N19261);
nor NOR2 (N19267, N19264, N11013);
xor XOR2 (N19268, N19257, N2728);
xor XOR2 (N19269, N19265, N18821);
and AND2 (N19270, N19267, N1040);
buf BUF1 (N19271, N19269);
or OR2 (N19272, N19262, N5865);
nor NOR4 (N19273, N19256, N4039, N1089, N12890);
buf BUF1 (N19274, N19251);
nand NAND2 (N19275, N19245, N17073);
buf BUF1 (N19276, N19271);
xor XOR2 (N19277, N19275, N4002);
nor NOR2 (N19278, N19272, N19124);
nor NOR2 (N19279, N19277, N7054);
or OR2 (N19280, N19260, N18079);
nor NOR2 (N19281, N19258, N18824);
not NOT1 (N19282, N19276);
nor NOR3 (N19283, N19281, N8112, N3338);
nand NAND2 (N19284, N19282, N8721);
not NOT1 (N19285, N19274);
nand NAND4 (N19286, N19285, N8803, N7639, N10311);
xor XOR2 (N19287, N19283, N8177);
xor XOR2 (N19288, N19287, N19235);
buf BUF1 (N19289, N19279);
nor NOR2 (N19290, N19278, N3027);
buf BUF1 (N19291, N19288);
buf BUF1 (N19292, N19280);
not NOT1 (N19293, N19270);
buf BUF1 (N19294, N19268);
not NOT1 (N19295, N19290);
not NOT1 (N19296, N19286);
xor XOR2 (N19297, N19292, N11730);
buf BUF1 (N19298, N19291);
nor NOR3 (N19299, N19266, N11639, N16386);
buf BUF1 (N19300, N19273);
xor XOR2 (N19301, N19293, N7359);
buf BUF1 (N19302, N19289);
nor NOR4 (N19303, N19298, N11627, N1614, N11342);
nand NAND4 (N19304, N19300, N5316, N962, N17472);
nor NOR4 (N19305, N19284, N6419, N4751, N10089);
xor XOR2 (N19306, N19302, N9002);
buf BUF1 (N19307, N19294);
or OR4 (N19308, N19296, N11599, N10737, N16976);
or OR3 (N19309, N19304, N6268, N12564);
not NOT1 (N19310, N19308);
nand NAND3 (N19311, N19305, N11635, N17197);
buf BUF1 (N19312, N19307);
buf BUF1 (N19313, N19295);
xor XOR2 (N19314, N19310, N16721);
not NOT1 (N19315, N19312);
not NOT1 (N19316, N19309);
nor NOR2 (N19317, N19311, N17685);
not NOT1 (N19318, N19314);
buf BUF1 (N19319, N19313);
or OR3 (N19320, N19303, N2240, N12884);
nand NAND3 (N19321, N19297, N17379, N663);
nor NOR2 (N19322, N19318, N5249);
xor XOR2 (N19323, N19321, N12802);
nand NAND2 (N19324, N19323, N17000);
nand NAND2 (N19325, N19316, N6510);
and AND3 (N19326, N19317, N4726, N13353);
and AND3 (N19327, N19299, N17150, N16377);
not NOT1 (N19328, N19324);
buf BUF1 (N19329, N19327);
nand NAND3 (N19330, N19322, N15534, N6179);
not NOT1 (N19331, N19306);
and AND3 (N19332, N19328, N2713, N8450);
nand NAND4 (N19333, N19320, N318, N4887, N7492);
not NOT1 (N19334, N19325);
and AND2 (N19335, N19315, N13686);
and AND4 (N19336, N19326, N859, N11452, N8165);
xor XOR2 (N19337, N19336, N8595);
nor NOR2 (N19338, N19330, N2509);
nand NAND2 (N19339, N19331, N17900);
not NOT1 (N19340, N19332);
xor XOR2 (N19341, N19334, N16284);
nand NAND3 (N19342, N19333, N14073, N1605);
not NOT1 (N19343, N19339);
nor NOR4 (N19344, N19341, N9612, N3636, N9760);
nor NOR4 (N19345, N19319, N15928, N14166, N3648);
not NOT1 (N19346, N19343);
nor NOR2 (N19347, N19301, N14219);
nor NOR2 (N19348, N19346, N5491);
buf BUF1 (N19349, N19338);
not NOT1 (N19350, N19340);
nand NAND2 (N19351, N19335, N8276);
nand NAND3 (N19352, N19342, N9948, N3401);
not NOT1 (N19353, N19348);
not NOT1 (N19354, N19350);
or OR2 (N19355, N19347, N11774);
nor NOR4 (N19356, N19352, N11588, N7996, N11882);
or OR4 (N19357, N19356, N6071, N14532, N16220);
nor NOR3 (N19358, N19354, N5211, N10456);
nand NAND3 (N19359, N19355, N18653, N5162);
buf BUF1 (N19360, N19357);
buf BUF1 (N19361, N19349);
not NOT1 (N19362, N19360);
xor XOR2 (N19363, N19358, N13392);
not NOT1 (N19364, N19351);
or OR4 (N19365, N19345, N7731, N5115, N3918);
not NOT1 (N19366, N19364);
or OR4 (N19367, N19359, N5728, N13880, N13771);
nand NAND2 (N19368, N19361, N9266);
buf BUF1 (N19369, N19363);
not NOT1 (N19370, N19329);
or OR2 (N19371, N19367, N4600);
buf BUF1 (N19372, N19370);
or OR3 (N19373, N19369, N9679, N5037);
nor NOR3 (N19374, N19344, N9535, N15547);
nand NAND3 (N19375, N19372, N10949, N15998);
not NOT1 (N19376, N19337);
nor NOR4 (N19377, N19376, N10292, N17179, N17958);
nor NOR2 (N19378, N19353, N11267);
nor NOR3 (N19379, N19365, N15605, N5718);
xor XOR2 (N19380, N19371, N10235);
xor XOR2 (N19381, N19375, N6249);
nand NAND4 (N19382, N19362, N13525, N3064, N12004);
not NOT1 (N19383, N19381);
and AND3 (N19384, N19382, N3795, N10910);
or OR2 (N19385, N19383, N13508);
buf BUF1 (N19386, N19368);
nor NOR4 (N19387, N19366, N13399, N4395, N11837);
not NOT1 (N19388, N19374);
nand NAND4 (N19389, N19379, N3752, N328, N17682);
nor NOR3 (N19390, N19385, N10771, N10193);
or OR2 (N19391, N19373, N8079);
or OR4 (N19392, N19384, N12634, N10199, N7619);
nand NAND4 (N19393, N19389, N12468, N11351, N2533);
nor NOR4 (N19394, N19388, N4027, N14917, N11509);
and AND2 (N19395, N19380, N620);
buf BUF1 (N19396, N19387);
nand NAND2 (N19397, N19396, N13557);
and AND4 (N19398, N19397, N3276, N10276, N12786);
and AND2 (N19399, N19395, N11812);
nor NOR4 (N19400, N19391, N14814, N19203, N805);
not NOT1 (N19401, N19400);
or OR4 (N19402, N19378, N18410, N8307, N18654);
xor XOR2 (N19403, N19398, N1890);
nor NOR4 (N19404, N19401, N34, N10902, N8007);
and AND4 (N19405, N19393, N10759, N4456, N10576);
nor NOR3 (N19406, N19403, N13674, N8355);
or OR3 (N19407, N19405, N1877, N9010);
and AND3 (N19408, N19394, N5997, N19200);
buf BUF1 (N19409, N19404);
nand NAND3 (N19410, N19409, N14641, N3005);
xor XOR2 (N19411, N19402, N7017);
or OR4 (N19412, N19392, N16162, N14708, N12974);
not NOT1 (N19413, N19411);
or OR4 (N19414, N19408, N14864, N17308, N7634);
or OR3 (N19415, N19406, N3913, N9584);
nor NOR4 (N19416, N19386, N9977, N5970, N1655);
nand NAND3 (N19417, N19399, N16025, N7395);
buf BUF1 (N19418, N19412);
or OR2 (N19419, N19407, N2290);
not NOT1 (N19420, N19410);
and AND3 (N19421, N19390, N14616, N253);
buf BUF1 (N19422, N19414);
xor XOR2 (N19423, N19419, N4952);
nand NAND3 (N19424, N19413, N5424, N14217);
buf BUF1 (N19425, N19418);
and AND3 (N19426, N19420, N18029, N3359);
not NOT1 (N19427, N19417);
nor NOR2 (N19428, N19426, N11358);
or OR3 (N19429, N19423, N16969, N7251);
buf BUF1 (N19430, N19429);
nand NAND3 (N19431, N19424, N15488, N2479);
not NOT1 (N19432, N19421);
or OR2 (N19433, N19428, N12084);
or OR4 (N19434, N19415, N11789, N9563, N16867);
not NOT1 (N19435, N19377);
not NOT1 (N19436, N19433);
nand NAND3 (N19437, N19436, N13637, N16621);
not NOT1 (N19438, N19437);
not NOT1 (N19439, N19416);
xor XOR2 (N19440, N19425, N14383);
nand NAND2 (N19441, N19432, N1185);
buf BUF1 (N19442, N19430);
xor XOR2 (N19443, N19434, N13414);
or OR2 (N19444, N19440, N15707);
nand NAND4 (N19445, N19444, N5906, N18549, N6594);
xor XOR2 (N19446, N19441, N14381);
nor NOR3 (N19447, N19435, N12107, N3494);
or OR3 (N19448, N19442, N11627, N2244);
nand NAND4 (N19449, N19445, N7768, N8231, N8328);
not NOT1 (N19450, N19427);
not NOT1 (N19451, N19450);
and AND3 (N19452, N19443, N7983, N5615);
nand NAND4 (N19453, N19438, N6631, N17845, N15043);
xor XOR2 (N19454, N19453, N2809);
xor XOR2 (N19455, N19451, N17466);
or OR3 (N19456, N19455, N11833, N726);
not NOT1 (N19457, N19422);
not NOT1 (N19458, N19439);
not NOT1 (N19459, N19449);
or OR3 (N19460, N19446, N13884, N7884);
buf BUF1 (N19461, N19457);
nand NAND2 (N19462, N19431, N12275);
xor XOR2 (N19463, N19447, N4326);
xor XOR2 (N19464, N19461, N2425);
nand NAND3 (N19465, N19458, N13273, N3692);
and AND3 (N19466, N19448, N3972, N15635);
buf BUF1 (N19467, N19464);
and AND4 (N19468, N19459, N1110, N146, N13255);
and AND2 (N19469, N19468, N12741);
xor XOR2 (N19470, N19454, N4803);
xor XOR2 (N19471, N19466, N13828);
nand NAND4 (N19472, N19462, N19056, N19149, N6747);
not NOT1 (N19473, N19469);
not NOT1 (N19474, N19473);
not NOT1 (N19475, N19463);
xor XOR2 (N19476, N19460, N16074);
xor XOR2 (N19477, N19475, N3047);
nor NOR4 (N19478, N19470, N15223, N4704, N828);
xor XOR2 (N19479, N19456, N1244);
nand NAND3 (N19480, N19467, N7497, N10521);
nor NOR2 (N19481, N19471, N2210);
nand NAND4 (N19482, N19465, N17286, N4127, N8870);
nor NOR2 (N19483, N19474, N7326);
and AND3 (N19484, N19477, N14189, N16414);
xor XOR2 (N19485, N19484, N12025);
not NOT1 (N19486, N19485);
buf BUF1 (N19487, N19480);
and AND4 (N19488, N19487, N12551, N17451, N7133);
xor XOR2 (N19489, N19483, N4071);
or OR3 (N19490, N19452, N3935, N3893);
nand NAND2 (N19491, N19490, N2897);
nand NAND3 (N19492, N19481, N19122, N2859);
not NOT1 (N19493, N19479);
buf BUF1 (N19494, N19478);
and AND3 (N19495, N19472, N5832, N4436);
nand NAND4 (N19496, N19491, N93, N8139, N11764);
nand NAND4 (N19497, N19494, N13123, N18277, N16715);
or OR3 (N19498, N19489, N12004, N9998);
xor XOR2 (N19499, N19482, N16675);
or OR3 (N19500, N19498, N7130, N1127);
not NOT1 (N19501, N19492);
nor NOR4 (N19502, N19493, N7568, N7179, N2167);
or OR3 (N19503, N19499, N6174, N9177);
and AND2 (N19504, N19486, N10363);
nand NAND2 (N19505, N19497, N5673);
buf BUF1 (N19506, N19501);
buf BUF1 (N19507, N19495);
nand NAND2 (N19508, N19506, N9319);
nand NAND4 (N19509, N19508, N6560, N1750, N3212);
xor XOR2 (N19510, N19496, N2159);
and AND4 (N19511, N19504, N11671, N12355, N13513);
or OR3 (N19512, N19505, N18809, N17624);
nand NAND4 (N19513, N19500, N11773, N6546, N18091);
or OR4 (N19514, N19509, N14417, N10462, N18577);
xor XOR2 (N19515, N19512, N13000);
not NOT1 (N19516, N19502);
or OR4 (N19517, N19516, N18053, N747, N18696);
or OR3 (N19518, N19503, N17255, N14101);
buf BUF1 (N19519, N19488);
or OR3 (N19520, N19507, N18797, N17214);
buf BUF1 (N19521, N19514);
nor NOR2 (N19522, N19476, N5289);
not NOT1 (N19523, N19519);
nor NOR4 (N19524, N19518, N15322, N14372, N11626);
nand NAND3 (N19525, N19520, N8956, N1057);
buf BUF1 (N19526, N19511);
or OR4 (N19527, N19510, N13656, N14203, N11423);
and AND4 (N19528, N19527, N17754, N220, N12945);
or OR4 (N19529, N19524, N6722, N7951, N10573);
or OR4 (N19530, N19515, N14149, N14699, N287);
buf BUF1 (N19531, N19523);
not NOT1 (N19532, N19528);
buf BUF1 (N19533, N19525);
and AND2 (N19534, N19531, N4996);
or OR4 (N19535, N19517, N1722, N4571, N14850);
nand NAND3 (N19536, N19535, N7760, N7237);
buf BUF1 (N19537, N19536);
and AND2 (N19538, N19529, N18966);
buf BUF1 (N19539, N19521);
not NOT1 (N19540, N19532);
nor NOR3 (N19541, N19513, N18814, N14593);
xor XOR2 (N19542, N19538, N19058);
buf BUF1 (N19543, N19541);
buf BUF1 (N19544, N19542);
or OR2 (N19545, N19530, N13907);
nand NAND3 (N19546, N19522, N15594, N5341);
or OR2 (N19547, N19544, N3538);
nor NOR3 (N19548, N19539, N6620, N7848);
not NOT1 (N19549, N19547);
xor XOR2 (N19550, N19526, N4259);
and AND3 (N19551, N19550, N5352, N887);
not NOT1 (N19552, N19543);
and AND4 (N19553, N19552, N17057, N11320, N16610);
and AND2 (N19554, N19551, N8037);
nor NOR3 (N19555, N19533, N15180, N16601);
xor XOR2 (N19556, N19546, N16109);
nand NAND2 (N19557, N19537, N17249);
buf BUF1 (N19558, N19548);
or OR4 (N19559, N19540, N3098, N11219, N8016);
xor XOR2 (N19560, N19545, N12106);
and AND4 (N19561, N19553, N12195, N5604, N2408);
xor XOR2 (N19562, N19558, N4248);
not NOT1 (N19563, N19557);
nor NOR2 (N19564, N19556, N6651);
buf BUF1 (N19565, N19563);
nand NAND4 (N19566, N19565, N17816, N7290, N14935);
nand NAND2 (N19567, N19566, N1184);
nor NOR4 (N19568, N19559, N4330, N8062, N6043);
not NOT1 (N19569, N19555);
not NOT1 (N19570, N19561);
not NOT1 (N19571, N19567);
nand NAND4 (N19572, N19549, N17848, N18645, N18147);
nand NAND4 (N19573, N19564, N5628, N4381, N14684);
xor XOR2 (N19574, N19562, N16969);
or OR2 (N19575, N19560, N18677);
not NOT1 (N19576, N19568);
and AND3 (N19577, N19572, N13408, N8524);
nand NAND3 (N19578, N19577, N10688, N14590);
not NOT1 (N19579, N19573);
not NOT1 (N19580, N19569);
and AND4 (N19581, N19571, N12605, N18839, N14422);
nor NOR4 (N19582, N19580, N2212, N16962, N8483);
not NOT1 (N19583, N19579);
and AND2 (N19584, N19583, N14024);
xor XOR2 (N19585, N19582, N3905);
buf BUF1 (N19586, N19585);
xor XOR2 (N19587, N19584, N18669);
or OR3 (N19588, N19534, N10246, N1598);
nand NAND4 (N19589, N19578, N6933, N12641, N722);
not NOT1 (N19590, N19586);
not NOT1 (N19591, N19570);
nand NAND4 (N19592, N19589, N4926, N4565, N15546);
and AND2 (N19593, N19591, N9116);
buf BUF1 (N19594, N19587);
nor NOR3 (N19595, N19574, N15291, N12620);
or OR2 (N19596, N19581, N10658);
nand NAND3 (N19597, N19576, N18563, N10768);
or OR2 (N19598, N19554, N16262);
not NOT1 (N19599, N19575);
nand NAND3 (N19600, N19598, N19515, N11326);
buf BUF1 (N19601, N19599);
buf BUF1 (N19602, N19601);
and AND4 (N19603, N19600, N8490, N9710, N13666);
xor XOR2 (N19604, N19588, N14068);
buf BUF1 (N19605, N19593);
and AND3 (N19606, N19596, N5598, N18046);
and AND4 (N19607, N19592, N7000, N3972, N6743);
nor NOR4 (N19608, N19606, N4973, N11242, N7073);
and AND3 (N19609, N19607, N4983, N2809);
nor NOR4 (N19610, N19594, N15310, N18783, N11450);
xor XOR2 (N19611, N19605, N910);
nor NOR2 (N19612, N19604, N2673);
and AND3 (N19613, N19602, N1751, N10504);
or OR4 (N19614, N19595, N11028, N14629, N16293);
buf BUF1 (N19615, N19613);
buf BUF1 (N19616, N19610);
nand NAND4 (N19617, N19611, N5323, N14868, N14874);
not NOT1 (N19618, N19603);
not NOT1 (N19619, N19614);
nor NOR3 (N19620, N19608, N7507, N3111);
and AND3 (N19621, N19612, N3991, N11636);
nor NOR3 (N19622, N19615, N7211, N16272);
xor XOR2 (N19623, N19597, N3278);
buf BUF1 (N19624, N19621);
xor XOR2 (N19625, N19617, N3935);
xor XOR2 (N19626, N19622, N1729);
nand NAND2 (N19627, N19590, N3204);
or OR2 (N19628, N19620, N9164);
nand NAND2 (N19629, N19623, N1654);
buf BUF1 (N19630, N19626);
and AND3 (N19631, N19619, N2503, N18293);
buf BUF1 (N19632, N19631);
or OR2 (N19633, N19618, N16450);
xor XOR2 (N19634, N19616, N6942);
nor NOR3 (N19635, N19625, N4432, N16479);
xor XOR2 (N19636, N19627, N15592);
not NOT1 (N19637, N19632);
and AND3 (N19638, N19636, N18065, N9857);
or OR4 (N19639, N19624, N2438, N3039, N5867);
buf BUF1 (N19640, N19609);
not NOT1 (N19641, N19640);
or OR2 (N19642, N19634, N9059);
and AND2 (N19643, N19630, N4635);
nor NOR4 (N19644, N19641, N14636, N10060, N8602);
or OR2 (N19645, N19642, N12972);
xor XOR2 (N19646, N19645, N11315);
nand NAND2 (N19647, N19638, N793);
and AND3 (N19648, N19637, N3957, N17089);
nand NAND2 (N19649, N19635, N10819);
nor NOR4 (N19650, N19647, N5968, N16849, N1471);
and AND3 (N19651, N19639, N14336, N15657);
or OR2 (N19652, N19643, N2733);
not NOT1 (N19653, N19644);
buf BUF1 (N19654, N19646);
nand NAND4 (N19655, N19649, N11553, N11058, N12872);
and AND2 (N19656, N19653, N2709);
buf BUF1 (N19657, N19652);
buf BUF1 (N19658, N19633);
nand NAND2 (N19659, N19658, N17535);
not NOT1 (N19660, N19628);
xor XOR2 (N19661, N19629, N13301);
buf BUF1 (N19662, N19651);
buf BUF1 (N19663, N19657);
nand NAND3 (N19664, N19656, N8745, N14822);
and AND4 (N19665, N19664, N13628, N4798, N9022);
xor XOR2 (N19666, N19659, N13301);
or OR4 (N19667, N19662, N882, N4714, N16867);
nand NAND4 (N19668, N19666, N17281, N1120, N16682);
buf BUF1 (N19669, N19661);
xor XOR2 (N19670, N19668, N19189);
nor NOR3 (N19671, N19670, N2644, N19393);
nor NOR4 (N19672, N19654, N19485, N3380, N15767);
xor XOR2 (N19673, N19672, N13885);
or OR3 (N19674, N19671, N5741, N16854);
nand NAND3 (N19675, N19674, N9170, N8172);
not NOT1 (N19676, N19655);
and AND4 (N19677, N19650, N15792, N9865, N11942);
not NOT1 (N19678, N19667);
nor NOR2 (N19679, N19669, N508);
or OR2 (N19680, N19648, N17755);
and AND2 (N19681, N19665, N12008);
nand NAND4 (N19682, N19663, N10268, N5347, N10517);
nand NAND2 (N19683, N19677, N9154);
buf BUF1 (N19684, N19680);
xor XOR2 (N19685, N19673, N19335);
or OR4 (N19686, N19660, N714, N2843, N557);
and AND4 (N19687, N19682, N16002, N6937, N8407);
nand NAND3 (N19688, N19686, N8583, N14714);
and AND3 (N19689, N19688, N15297, N15786);
buf BUF1 (N19690, N19685);
and AND4 (N19691, N19684, N381, N8714, N15054);
or OR4 (N19692, N19675, N13913, N2489, N17358);
xor XOR2 (N19693, N19691, N19606);
and AND4 (N19694, N19689, N11242, N8685, N15721);
or OR3 (N19695, N19678, N12173, N13568);
nand NAND3 (N19696, N19695, N13613, N15871);
buf BUF1 (N19697, N19681);
nor NOR4 (N19698, N19690, N2798, N10926, N3504);
xor XOR2 (N19699, N19687, N19526);
or OR3 (N19700, N19697, N317, N18037);
or OR4 (N19701, N19692, N3432, N4187, N8316);
nor NOR2 (N19702, N19679, N13480);
xor XOR2 (N19703, N19700, N12243);
not NOT1 (N19704, N19699);
nand NAND4 (N19705, N19676, N6444, N1372, N960);
not NOT1 (N19706, N19701);
xor XOR2 (N19707, N19706, N8887);
or OR2 (N19708, N19683, N18535);
or OR4 (N19709, N19702, N6306, N10233, N3216);
xor XOR2 (N19710, N19693, N14495);
xor XOR2 (N19711, N19698, N130);
not NOT1 (N19712, N19696);
not NOT1 (N19713, N19704);
and AND2 (N19714, N19713, N6581);
xor XOR2 (N19715, N19709, N9810);
buf BUF1 (N19716, N19711);
not NOT1 (N19717, N19714);
or OR2 (N19718, N19710, N2910);
nand NAND3 (N19719, N19703, N898, N9845);
nand NAND4 (N19720, N19712, N1160, N5110, N4882);
not NOT1 (N19721, N19705);
xor XOR2 (N19722, N19717, N1383);
or OR4 (N19723, N19722, N12055, N151, N12688);
and AND2 (N19724, N19707, N10869);
buf BUF1 (N19725, N19724);
or OR2 (N19726, N19725, N6683);
xor XOR2 (N19727, N19708, N16202);
and AND2 (N19728, N19715, N2753);
and AND3 (N19729, N19716, N14502, N1954);
and AND3 (N19730, N19729, N6892, N16548);
not NOT1 (N19731, N19726);
nor NOR3 (N19732, N19731, N6380, N16528);
xor XOR2 (N19733, N19723, N19523);
or OR4 (N19734, N19694, N7831, N2789, N18464);
nor NOR3 (N19735, N19719, N19565, N277);
nor NOR4 (N19736, N19730, N17619, N19050, N15038);
and AND3 (N19737, N19734, N5748, N4470);
buf BUF1 (N19738, N19733);
not NOT1 (N19739, N19728);
or OR3 (N19740, N19727, N1633, N7947);
or OR3 (N19741, N19738, N13360, N10054);
nor NOR4 (N19742, N19718, N19628, N3139, N4087);
and AND2 (N19743, N19741, N19372);
or OR2 (N19744, N19739, N18785);
nand NAND3 (N19745, N19732, N17652, N12637);
not NOT1 (N19746, N19721);
nor NOR2 (N19747, N19742, N11675);
not NOT1 (N19748, N19737);
nor NOR4 (N19749, N19746, N10230, N4264, N496);
nand NAND4 (N19750, N19747, N17269, N19079, N2328);
not NOT1 (N19751, N19743);
buf BUF1 (N19752, N19736);
nand NAND4 (N19753, N19750, N16603, N19677, N11766);
nand NAND2 (N19754, N19735, N13958);
not NOT1 (N19755, N19749);
buf BUF1 (N19756, N19745);
buf BUF1 (N19757, N19748);
buf BUF1 (N19758, N19752);
nor NOR4 (N19759, N19758, N11218, N13954, N4050);
xor XOR2 (N19760, N19720, N13384);
or OR3 (N19761, N19760, N17207, N19397);
and AND3 (N19762, N19757, N3803, N16910);
nor NOR2 (N19763, N19762, N3885);
nor NOR4 (N19764, N19759, N15600, N14263, N9006);
buf BUF1 (N19765, N19751);
or OR3 (N19766, N19761, N15329, N14827);
or OR4 (N19767, N19744, N423, N157, N12760);
nand NAND3 (N19768, N19756, N4413, N8822);
and AND4 (N19769, N19766, N19503, N2559, N17171);
nand NAND3 (N19770, N19769, N8820, N5165);
and AND4 (N19771, N19763, N2380, N17599, N4723);
buf BUF1 (N19772, N19771);
xor XOR2 (N19773, N19770, N2161);
xor XOR2 (N19774, N19765, N10354);
nor NOR2 (N19775, N19754, N10164);
nand NAND3 (N19776, N19755, N15746, N10553);
buf BUF1 (N19777, N19776);
buf BUF1 (N19778, N19774);
nor NOR4 (N19779, N19767, N14006, N19569, N17132);
not NOT1 (N19780, N19779);
nand NAND3 (N19781, N19772, N4940, N10468);
nor NOR2 (N19782, N19768, N8456);
buf BUF1 (N19783, N19777);
nand NAND4 (N19784, N19753, N1484, N10506, N3901);
nor NOR2 (N19785, N19784, N10143);
or OR3 (N19786, N19785, N10721, N8136);
buf BUF1 (N19787, N19778);
xor XOR2 (N19788, N19781, N10640);
xor XOR2 (N19789, N19780, N19005);
or OR2 (N19790, N19783, N10595);
nand NAND4 (N19791, N19790, N19481, N8069, N9670);
not NOT1 (N19792, N19740);
nand NAND3 (N19793, N19791, N8240, N19746);
and AND2 (N19794, N19793, N16908);
xor XOR2 (N19795, N19789, N4360);
nand NAND3 (N19796, N19764, N11640, N59);
and AND2 (N19797, N19782, N9684);
not NOT1 (N19798, N19794);
nor NOR2 (N19799, N19797, N18491);
not NOT1 (N19800, N19773);
or OR2 (N19801, N19796, N14849);
xor XOR2 (N19802, N19787, N5053);
xor XOR2 (N19803, N19801, N575);
buf BUF1 (N19804, N19802);
not NOT1 (N19805, N19795);
xor XOR2 (N19806, N19775, N15349);
buf BUF1 (N19807, N19792);
nor NOR3 (N19808, N19804, N2157, N3598);
buf BUF1 (N19809, N19805);
nand NAND4 (N19810, N19788, N10187, N334, N907);
or OR3 (N19811, N19786, N128, N2732);
xor XOR2 (N19812, N19811, N8523);
and AND3 (N19813, N19810, N14682, N7895);
nor NOR2 (N19814, N19813, N14834);
not NOT1 (N19815, N19812);
nor NOR2 (N19816, N19808, N17455);
xor XOR2 (N19817, N19807, N9963);
not NOT1 (N19818, N19800);
and AND3 (N19819, N19799, N12583, N18714);
and AND4 (N19820, N19798, N19075, N18196, N1101);
and AND4 (N19821, N19816, N15187, N7743, N9071);
nand NAND4 (N19822, N19803, N7742, N10723, N8765);
nand NAND3 (N19823, N19814, N15926, N19335);
nand NAND3 (N19824, N19823, N151, N624);
and AND4 (N19825, N19819, N3690, N13421, N3340);
xor XOR2 (N19826, N19806, N6683);
and AND2 (N19827, N19817, N18784);
not NOT1 (N19828, N19822);
xor XOR2 (N19829, N19826, N18686);
nand NAND3 (N19830, N19809, N9094, N18587);
or OR4 (N19831, N19815, N6619, N7166, N10155);
buf BUF1 (N19832, N19830);
and AND3 (N19833, N19820, N15621, N6218);
and AND4 (N19834, N19827, N7986, N7466, N6926);
and AND2 (N19835, N19821, N11220);
nor NOR4 (N19836, N19824, N15242, N4721, N15899);
or OR3 (N19837, N19829, N17289, N10429);
buf BUF1 (N19838, N19818);
xor XOR2 (N19839, N19834, N422);
nor NOR2 (N19840, N19825, N19070);
or OR4 (N19841, N19828, N4624, N1585, N16918);
xor XOR2 (N19842, N19837, N13716);
or OR3 (N19843, N19836, N5381, N11209);
buf BUF1 (N19844, N19835);
or OR2 (N19845, N19840, N1635);
nor NOR3 (N19846, N19833, N16239, N10501);
xor XOR2 (N19847, N19839, N1003);
or OR2 (N19848, N19838, N18691);
buf BUF1 (N19849, N19841);
not NOT1 (N19850, N19848);
buf BUF1 (N19851, N19843);
xor XOR2 (N19852, N19846, N166);
buf BUF1 (N19853, N19850);
buf BUF1 (N19854, N19851);
xor XOR2 (N19855, N19842, N5168);
xor XOR2 (N19856, N19855, N7609);
nor NOR4 (N19857, N19832, N5000, N1926, N17113);
or OR4 (N19858, N19853, N8801, N19642, N3073);
nor NOR3 (N19859, N19847, N4165, N7676);
nor NOR3 (N19860, N19856, N19564, N3166);
nand NAND3 (N19861, N19859, N10095, N12301);
or OR4 (N19862, N19844, N18891, N7895, N18057);
nor NOR3 (N19863, N19831, N12019, N11438);
buf BUF1 (N19864, N19845);
not NOT1 (N19865, N19849);
and AND3 (N19866, N19861, N14404, N12723);
nor NOR2 (N19867, N19857, N5966);
or OR2 (N19868, N19858, N8395);
nor NOR3 (N19869, N19867, N7000, N1957);
not NOT1 (N19870, N19860);
not NOT1 (N19871, N19865);
nand NAND4 (N19872, N19870, N10534, N4599, N6361);
not NOT1 (N19873, N19871);
nor NOR4 (N19874, N19862, N7169, N14987, N9996);
or OR2 (N19875, N19852, N9674);
and AND4 (N19876, N19864, N4851, N12028, N7209);
nand NAND3 (N19877, N19873, N12163, N3070);
nor NOR3 (N19878, N19877, N9846, N19699);
not NOT1 (N19879, N19868);
not NOT1 (N19880, N19875);
xor XOR2 (N19881, N19866, N7472);
not NOT1 (N19882, N19881);
nor NOR4 (N19883, N19874, N1144, N5480, N10091);
not NOT1 (N19884, N19872);
buf BUF1 (N19885, N19883);
or OR2 (N19886, N19878, N1022);
nor NOR3 (N19887, N19885, N7494, N1615);
nor NOR3 (N19888, N19882, N1633, N8919);
xor XOR2 (N19889, N19886, N8919);
and AND2 (N19890, N19863, N65);
and AND4 (N19891, N19879, N15052, N19624, N574);
not NOT1 (N19892, N19887);
xor XOR2 (N19893, N19884, N2743);
nand NAND2 (N19894, N19893, N7790);
nor NOR2 (N19895, N19876, N2065);
and AND2 (N19896, N19880, N8883);
and AND4 (N19897, N19891, N18067, N19578, N12253);
or OR4 (N19898, N19892, N18849, N3123, N2541);
nand NAND2 (N19899, N19889, N10905);
buf BUF1 (N19900, N19897);
xor XOR2 (N19901, N19900, N10648);
xor XOR2 (N19902, N19854, N15071);
nand NAND2 (N19903, N19901, N11728);
or OR2 (N19904, N19903, N2843);
not NOT1 (N19905, N19894);
or OR3 (N19906, N19896, N14574, N9027);
xor XOR2 (N19907, N19906, N10609);
not NOT1 (N19908, N19888);
not NOT1 (N19909, N19869);
and AND2 (N19910, N19898, N12241);
buf BUF1 (N19911, N19907);
or OR4 (N19912, N19910, N7516, N3527, N16820);
nor NOR2 (N19913, N19899, N7769);
or OR3 (N19914, N19908, N18202, N6176);
nand NAND2 (N19915, N19905, N10494);
nand NAND3 (N19916, N19915, N1602, N8964);
or OR3 (N19917, N19916, N14826, N12989);
buf BUF1 (N19918, N19917);
not NOT1 (N19919, N19904);
nand NAND3 (N19920, N19911, N4330, N5124);
buf BUF1 (N19921, N19914);
nor NOR4 (N19922, N19890, N6726, N4947, N10856);
and AND2 (N19923, N19895, N16288);
nand NAND4 (N19924, N19909, N3563, N12253, N7284);
and AND3 (N19925, N19913, N13785, N2822);
nand NAND3 (N19926, N19918, N17774, N9755);
buf BUF1 (N19927, N19924);
nor NOR3 (N19928, N19926, N11485, N10042);
and AND4 (N19929, N19919, N1426, N11504, N19624);
nor NOR4 (N19930, N19929, N880, N48, N15157);
buf BUF1 (N19931, N19912);
nand NAND4 (N19932, N19921, N13988, N16168, N8700);
buf BUF1 (N19933, N19902);
nor NOR3 (N19934, N19927, N82, N10293);
buf BUF1 (N19935, N19934);
and AND2 (N19936, N19925, N2411);
and AND4 (N19937, N19923, N8770, N13249, N2141);
not NOT1 (N19938, N19931);
xor XOR2 (N19939, N19933, N13333);
nand NAND3 (N19940, N19932, N15875, N13745);
nor NOR2 (N19941, N19940, N3328);
nor NOR2 (N19942, N19930, N17193);
xor XOR2 (N19943, N19920, N11331);
nor NOR4 (N19944, N19941, N112, N14632, N19140);
nand NAND4 (N19945, N19943, N10097, N15644, N18109);
buf BUF1 (N19946, N19936);
nor NOR3 (N19947, N19945, N11630, N11513);
not NOT1 (N19948, N19928);
or OR3 (N19949, N19942, N6790, N19898);
nor NOR3 (N19950, N19947, N19144, N12151);
nor NOR3 (N19951, N19922, N11121, N19284);
nor NOR4 (N19952, N19950, N11359, N4361, N16442);
and AND2 (N19953, N19951, N7291);
nand NAND4 (N19954, N19935, N17797, N18872, N15098);
or OR3 (N19955, N19946, N13524, N7713);
and AND4 (N19956, N19954, N1935, N7798, N1795);
or OR3 (N19957, N19937, N12405, N8190);
buf BUF1 (N19958, N19949);
nand NAND4 (N19959, N19953, N5496, N16329, N19378);
and AND4 (N19960, N19958, N8468, N2319, N13790);
not NOT1 (N19961, N19948);
buf BUF1 (N19962, N19961);
nand NAND3 (N19963, N19939, N12970, N11315);
buf BUF1 (N19964, N19960);
nand NAND2 (N19965, N19962, N12250);
or OR4 (N19966, N19938, N12684, N16932, N16124);
xor XOR2 (N19967, N19966, N2618);
and AND3 (N19968, N19944, N13782, N2895);
and AND4 (N19969, N19968, N11244, N17504, N10654);
and AND4 (N19970, N19969, N4666, N13338, N13417);
and AND4 (N19971, N19964, N16453, N11256, N8747);
or OR4 (N19972, N19965, N806, N14800, N16373);
nor NOR4 (N19973, N19959, N13144, N15580, N6366);
nor NOR4 (N19974, N19973, N1160, N3542, N5422);
xor XOR2 (N19975, N19952, N18078);
buf BUF1 (N19976, N19974);
nor NOR3 (N19977, N19956, N12992, N15156);
nand NAND4 (N19978, N19967, N5383, N970, N5459);
and AND3 (N19979, N19972, N17090, N7151);
buf BUF1 (N19980, N19955);
nand NAND4 (N19981, N19970, N13428, N6532, N5461);
nor NOR2 (N19982, N19963, N3767);
xor XOR2 (N19983, N19979, N3339);
buf BUF1 (N19984, N19981);
nand NAND3 (N19985, N19980, N15797, N17613);
buf BUF1 (N19986, N19975);
not NOT1 (N19987, N19983);
xor XOR2 (N19988, N19985, N489);
or OR4 (N19989, N19987, N1676, N8959, N18300);
nand NAND2 (N19990, N19957, N4128);
buf BUF1 (N19991, N19976);
nor NOR3 (N19992, N19990, N4014, N169);
nand NAND2 (N19993, N19986, N10387);
xor XOR2 (N19994, N19991, N8209);
buf BUF1 (N19995, N19994);
not NOT1 (N19996, N19982);
xor XOR2 (N19997, N19993, N19007);
not NOT1 (N19998, N19989);
nor NOR2 (N19999, N19995, N10051);
and AND2 (N20000, N19996, N3202);
and AND3 (N20001, N19999, N12916, N6159);
buf BUF1 (N20002, N19998);
or OR2 (N20003, N20002, N11558);
nand NAND2 (N20004, N19978, N12348);
xor XOR2 (N20005, N19988, N16208);
nor NOR3 (N20006, N19977, N15596, N8482);
and AND4 (N20007, N20006, N7975, N2925, N5447);
xor XOR2 (N20008, N20004, N258);
not NOT1 (N20009, N20003);
or OR3 (N20010, N20001, N2901, N20005);
xor XOR2 (N20011, N6232, N6205);
nor NOR3 (N20012, N20010, N13458, N14337);
and AND2 (N20013, N20008, N3272);
buf BUF1 (N20014, N20000);
xor XOR2 (N20015, N19971, N1547);
not NOT1 (N20016, N19997);
not NOT1 (N20017, N20013);
xor XOR2 (N20018, N20007, N13354);
buf BUF1 (N20019, N20018);
or OR4 (N20020, N20011, N15533, N6730, N12024);
or OR3 (N20021, N20019, N3383, N16775);
or OR3 (N20022, N20016, N6345, N929);
nor NOR3 (N20023, N20012, N16509, N19992);
buf BUF1 (N20024, N5917);
nor NOR2 (N20025, N20023, N14853);
or OR4 (N20026, N20025, N11887, N5864, N5601);
nor NOR4 (N20027, N20009, N14670, N6448, N8423);
buf BUF1 (N20028, N20014);
nand NAND3 (N20029, N20017, N17125, N18619);
and AND2 (N20030, N20028, N9929);
nand NAND2 (N20031, N20026, N6680);
nand NAND4 (N20032, N20022, N5264, N2787, N15869);
xor XOR2 (N20033, N20027, N17536);
nand NAND3 (N20034, N20030, N8028, N12117);
not NOT1 (N20035, N20024);
or OR3 (N20036, N20033, N10171, N10630);
nand NAND2 (N20037, N20021, N17948);
buf BUF1 (N20038, N20037);
nor NOR3 (N20039, N20015, N9711, N6420);
xor XOR2 (N20040, N20036, N10925);
not NOT1 (N20041, N20039);
nor NOR3 (N20042, N20034, N3099, N11346);
xor XOR2 (N20043, N20042, N17324);
buf BUF1 (N20044, N20035);
buf BUF1 (N20045, N20043);
xor XOR2 (N20046, N20031, N13961);
nor NOR3 (N20047, N20020, N3516, N9967);
nand NAND3 (N20048, N20040, N10179, N11322);
buf BUF1 (N20049, N20046);
or OR3 (N20050, N20041, N14661, N116);
xor XOR2 (N20051, N20048, N5152);
buf BUF1 (N20052, N20044);
not NOT1 (N20053, N19984);
buf BUF1 (N20054, N20029);
nor NOR3 (N20055, N20051, N6417, N7672);
nand NAND2 (N20056, N20038, N4073);
nor NOR3 (N20057, N20052, N19634, N10914);
not NOT1 (N20058, N20050);
not NOT1 (N20059, N20049);
or OR2 (N20060, N20045, N1573);
or OR2 (N20061, N20032, N14558);
buf BUF1 (N20062, N20053);
not NOT1 (N20063, N20058);
or OR4 (N20064, N20057, N861, N18432, N2174);
or OR3 (N20065, N20054, N3905, N14810);
buf BUF1 (N20066, N20062);
xor XOR2 (N20067, N20047, N1063);
nand NAND2 (N20068, N20066, N2650);
nor NOR2 (N20069, N20056, N3469);
buf BUF1 (N20070, N20063);
nor NOR4 (N20071, N20069, N11259, N11715, N16897);
buf BUF1 (N20072, N20059);
nor NOR3 (N20073, N20071, N19024, N17460);
not NOT1 (N20074, N20064);
nor NOR4 (N20075, N20055, N17592, N14567, N11323);
and AND2 (N20076, N20060, N7927);
nand NAND4 (N20077, N20076, N3928, N2161, N11930);
or OR4 (N20078, N20075, N6378, N14078, N4309);
not NOT1 (N20079, N20074);
xor XOR2 (N20080, N20068, N1643);
not NOT1 (N20081, N20073);
xor XOR2 (N20082, N20081, N1969);
nand NAND2 (N20083, N20067, N5181);
or OR2 (N20084, N20070, N14618);
and AND4 (N20085, N20061, N16464, N13737, N4850);
not NOT1 (N20086, N20077);
nand NAND4 (N20087, N20079, N16948, N3592, N5861);
xor XOR2 (N20088, N20083, N9126);
nor NOR2 (N20089, N20086, N15655);
nand NAND3 (N20090, N20089, N10179, N10709);
nor NOR4 (N20091, N20087, N19566, N877, N19493);
and AND3 (N20092, N20082, N15682, N6265);
buf BUF1 (N20093, N20065);
not NOT1 (N20094, N20085);
nand NAND2 (N20095, N20092, N382);
buf BUF1 (N20096, N20078);
or OR4 (N20097, N20094, N13725, N15234, N2538);
or OR4 (N20098, N20097, N19009, N9130, N16967);
buf BUF1 (N20099, N20093);
nand NAND4 (N20100, N20080, N3417, N7800, N8657);
or OR3 (N20101, N20099, N8104, N19732);
and AND2 (N20102, N20084, N5701);
nor NOR4 (N20103, N20090, N9173, N4592, N4571);
not NOT1 (N20104, N20095);
buf BUF1 (N20105, N20091);
and AND4 (N20106, N20101, N18625, N11289, N20053);
nand NAND2 (N20107, N20072, N5183);
or OR4 (N20108, N20106, N10735, N3672, N7619);
not NOT1 (N20109, N20102);
buf BUF1 (N20110, N20105);
and AND4 (N20111, N20107, N11914, N7880, N10027);
or OR2 (N20112, N20100, N13981);
xor XOR2 (N20113, N20098, N15565);
not NOT1 (N20114, N20112);
nand NAND2 (N20115, N20111, N6256);
buf BUF1 (N20116, N20096);
nor NOR3 (N20117, N20088, N14425, N17465);
not NOT1 (N20118, N20103);
xor XOR2 (N20119, N20118, N1475);
nand NAND4 (N20120, N20119, N2852, N421, N13189);
xor XOR2 (N20121, N20115, N12414);
and AND3 (N20122, N20116, N13458, N3027);
nand NAND2 (N20123, N20121, N1155);
xor XOR2 (N20124, N20104, N18465);
not NOT1 (N20125, N20120);
nand NAND3 (N20126, N20114, N14880, N8258);
or OR3 (N20127, N20117, N11619, N11190);
buf BUF1 (N20128, N20109);
nor NOR2 (N20129, N20128, N16081);
not NOT1 (N20130, N20125);
nand NAND3 (N20131, N20127, N18292, N3605);
and AND3 (N20132, N20126, N19596, N14857);
nand NAND4 (N20133, N20123, N4186, N13678, N16175);
buf BUF1 (N20134, N20110);
or OR4 (N20135, N20132, N10077, N19055, N11578);
and AND4 (N20136, N20129, N7850, N427, N3029);
xor XOR2 (N20137, N20136, N14807);
buf BUF1 (N20138, N20133);
or OR4 (N20139, N20131, N17873, N350, N19415);
not NOT1 (N20140, N20139);
or OR4 (N20141, N20124, N433, N9859, N1674);
nor NOR3 (N20142, N20134, N11501, N5944);
nor NOR3 (N20143, N20140, N20049, N20009);
or OR2 (N20144, N20135, N7159);
or OR2 (N20145, N20144, N13625);
not NOT1 (N20146, N20130);
and AND4 (N20147, N20137, N6597, N5015, N13341);
xor XOR2 (N20148, N20143, N12996);
nor NOR4 (N20149, N20141, N18365, N3872, N9376);
xor XOR2 (N20150, N20122, N19032);
nand NAND3 (N20151, N20113, N12194, N13693);
and AND2 (N20152, N20151, N11181);
not NOT1 (N20153, N20148);
not NOT1 (N20154, N20108);
buf BUF1 (N20155, N20145);
nand NAND4 (N20156, N20138, N15377, N11025, N1904);
not NOT1 (N20157, N20146);
nand NAND3 (N20158, N20142, N11744, N2455);
and AND3 (N20159, N20152, N18095, N3656);
nand NAND3 (N20160, N20159, N3043, N2259);
or OR3 (N20161, N20153, N19120, N17162);
nand NAND2 (N20162, N20161, N4705);
buf BUF1 (N20163, N20150);
or OR2 (N20164, N20160, N6250);
nand NAND2 (N20165, N20154, N6854);
xor XOR2 (N20166, N20147, N10045);
not NOT1 (N20167, N20164);
not NOT1 (N20168, N20149);
xor XOR2 (N20169, N20158, N409);
not NOT1 (N20170, N20162);
or OR2 (N20171, N20169, N8519);
xor XOR2 (N20172, N20167, N13335);
or OR4 (N20173, N20166, N5553, N18529, N17263);
nand NAND3 (N20174, N20170, N10369, N3473);
and AND3 (N20175, N20174, N5105, N4491);
nand NAND3 (N20176, N20171, N10499, N7930);
or OR2 (N20177, N20176, N15807);
or OR4 (N20178, N20157, N3825, N17652, N2103);
nor NOR4 (N20179, N20175, N8742, N5215, N5484);
nor NOR4 (N20180, N20155, N14647, N6751, N2024);
buf BUF1 (N20181, N20165);
buf BUF1 (N20182, N20168);
nand NAND4 (N20183, N20178, N7523, N17200, N8144);
nand NAND4 (N20184, N20183, N15939, N1026, N8383);
xor XOR2 (N20185, N20184, N10162);
or OR2 (N20186, N20182, N9530);
nor NOR2 (N20187, N20173, N13320);
nor NOR2 (N20188, N20179, N4822);
buf BUF1 (N20189, N20186);
xor XOR2 (N20190, N20181, N2221);
xor XOR2 (N20191, N20189, N19347);
buf BUF1 (N20192, N20156);
nor NOR4 (N20193, N20188, N7501, N11800, N13125);
nand NAND3 (N20194, N20172, N17462, N16290);
nor NOR3 (N20195, N20193, N6794, N15591);
and AND3 (N20196, N20187, N9692, N13477);
and AND2 (N20197, N20194, N4488);
nand NAND3 (N20198, N20195, N12612, N6053);
nand NAND2 (N20199, N20196, N18540);
or OR4 (N20200, N20191, N12672, N13607, N3437);
nor NOR3 (N20201, N20185, N16920, N18616);
nand NAND3 (N20202, N20177, N15480, N10570);
and AND2 (N20203, N20192, N15250);
nor NOR3 (N20204, N20180, N8564, N19163);
buf BUF1 (N20205, N20190);
not NOT1 (N20206, N20202);
or OR2 (N20207, N20201, N3922);
nor NOR3 (N20208, N20204, N7480, N20131);
and AND3 (N20209, N20206, N6845, N10311);
or OR3 (N20210, N20208, N7701, N6811);
and AND2 (N20211, N20203, N13237);
or OR4 (N20212, N20207, N14928, N19824, N10281);
not NOT1 (N20213, N20210);
and AND2 (N20214, N20209, N10775);
or OR3 (N20215, N20205, N18715, N9913);
nand NAND2 (N20216, N20198, N19366);
and AND2 (N20217, N20215, N6355);
and AND4 (N20218, N20163, N3830, N18169, N3079);
xor XOR2 (N20219, N20213, N17899);
buf BUF1 (N20220, N20197);
or OR3 (N20221, N20211, N6878, N16035);
nand NAND2 (N20222, N20220, N17667);
and AND4 (N20223, N20221, N12878, N5766, N15278);
xor XOR2 (N20224, N20200, N16365);
nor NOR4 (N20225, N20214, N4345, N17329, N6779);
buf BUF1 (N20226, N20199);
xor XOR2 (N20227, N20218, N1265);
nand NAND2 (N20228, N20227, N11133);
nand NAND3 (N20229, N20225, N13094, N8095);
not NOT1 (N20230, N20216);
nor NOR2 (N20231, N20223, N13646);
buf BUF1 (N20232, N20222);
nand NAND2 (N20233, N20224, N2334);
or OR2 (N20234, N20226, N11814);
nand NAND2 (N20235, N20219, N3800);
and AND2 (N20236, N20229, N11700);
buf BUF1 (N20237, N20236);
xor XOR2 (N20238, N20231, N10507);
and AND3 (N20239, N20228, N11923, N8580);
buf BUF1 (N20240, N20233);
and AND2 (N20241, N20238, N17868);
buf BUF1 (N20242, N20235);
xor XOR2 (N20243, N20242, N16751);
buf BUF1 (N20244, N20241);
nand NAND4 (N20245, N20212, N19918, N18616, N16047);
buf BUF1 (N20246, N20237);
nand NAND4 (N20247, N20246, N15829, N6280, N624);
nor NOR2 (N20248, N20247, N11721);
or OR4 (N20249, N20232, N9646, N10442, N16036);
nand NAND4 (N20250, N20245, N12490, N3422, N10567);
buf BUF1 (N20251, N20250);
or OR4 (N20252, N20240, N13954, N8180, N6407);
not NOT1 (N20253, N20249);
nor NOR2 (N20254, N20252, N12249);
not NOT1 (N20255, N20251);
or OR2 (N20256, N20248, N10300);
nand NAND3 (N20257, N20243, N13383, N12438);
buf BUF1 (N20258, N20230);
buf BUF1 (N20259, N20234);
nor NOR2 (N20260, N20257, N665);
or OR2 (N20261, N20256, N167);
nand NAND4 (N20262, N20255, N5578, N2006, N4359);
xor XOR2 (N20263, N20258, N15405);
nand NAND2 (N20264, N20261, N12196);
nor NOR3 (N20265, N20239, N20109, N14443);
or OR2 (N20266, N20263, N4570);
or OR4 (N20267, N20254, N13649, N12330, N15190);
not NOT1 (N20268, N20267);
buf BUF1 (N20269, N20268);
xor XOR2 (N20270, N20262, N2067);
buf BUF1 (N20271, N20265);
or OR3 (N20272, N20253, N7830, N17907);
and AND3 (N20273, N20244, N10248, N15016);
buf BUF1 (N20274, N20271);
or OR3 (N20275, N20260, N17145, N9716);
nand NAND2 (N20276, N20274, N13097);
not NOT1 (N20277, N20275);
nand NAND4 (N20278, N20273, N5931, N3219, N14625);
nor NOR2 (N20279, N20217, N12675);
and AND3 (N20280, N20269, N8931, N10237);
not NOT1 (N20281, N20278);
or OR2 (N20282, N20266, N5481);
and AND4 (N20283, N20264, N18873, N18468, N12793);
or OR4 (N20284, N20259, N19488, N14101, N17429);
nand NAND4 (N20285, N20279, N2993, N6778, N12027);
nor NOR3 (N20286, N20285, N11462, N117);
buf BUF1 (N20287, N20282);
or OR4 (N20288, N20284, N7753, N12056, N4257);
or OR4 (N20289, N20272, N1137, N19028, N6840);
xor XOR2 (N20290, N20276, N7133);
or OR3 (N20291, N20277, N6195, N14621);
and AND3 (N20292, N20288, N11243, N3958);
or OR4 (N20293, N20291, N7520, N9301, N18872);
or OR3 (N20294, N20293, N7148, N8830);
buf BUF1 (N20295, N20294);
buf BUF1 (N20296, N20281);
nand NAND4 (N20297, N20270, N11793, N3693, N906);
not NOT1 (N20298, N20289);
xor XOR2 (N20299, N20286, N19052);
nor NOR4 (N20300, N20298, N5106, N8655, N1437);
buf BUF1 (N20301, N20300);
buf BUF1 (N20302, N20299);
and AND4 (N20303, N20302, N4218, N19948, N10472);
and AND3 (N20304, N20295, N3531, N6611);
and AND2 (N20305, N20280, N16819);
or OR3 (N20306, N20296, N18879, N14820);
or OR3 (N20307, N20290, N12296, N17130);
and AND2 (N20308, N20287, N5515);
and AND3 (N20309, N20304, N19383, N5322);
buf BUF1 (N20310, N20292);
or OR2 (N20311, N20307, N4766);
nor NOR2 (N20312, N20303, N10170);
buf BUF1 (N20313, N20308);
and AND4 (N20314, N20305, N7767, N969, N3938);
nor NOR2 (N20315, N20306, N1967);
not NOT1 (N20316, N20312);
xor XOR2 (N20317, N20310, N8816);
not NOT1 (N20318, N20314);
xor XOR2 (N20319, N20317, N5756);
and AND2 (N20320, N20319, N700);
or OR3 (N20321, N20318, N10470, N4726);
and AND2 (N20322, N20316, N19573);
nand NAND4 (N20323, N20309, N14349, N7212, N18181);
or OR4 (N20324, N20322, N8692, N5869, N6986);
nand NAND4 (N20325, N20324, N13851, N11193, N7320);
or OR2 (N20326, N20320, N18189);
xor XOR2 (N20327, N20326, N13844);
buf BUF1 (N20328, N20297);
buf BUF1 (N20329, N20313);
not NOT1 (N20330, N20325);
nand NAND4 (N20331, N20321, N8884, N3707, N5753);
buf BUF1 (N20332, N20315);
buf BUF1 (N20333, N20331);
and AND2 (N20334, N20330, N10428);
buf BUF1 (N20335, N20333);
nand NAND2 (N20336, N20334, N3301);
buf BUF1 (N20337, N20327);
xor XOR2 (N20338, N20336, N17172);
nor NOR3 (N20339, N20337, N11501, N9034);
not NOT1 (N20340, N20311);
not NOT1 (N20341, N20323);
nor NOR2 (N20342, N20341, N12874);
not NOT1 (N20343, N20328);
xor XOR2 (N20344, N20335, N9402);
nand NAND3 (N20345, N20340, N10189, N6385);
nor NOR3 (N20346, N20342, N17261, N5959);
or OR2 (N20347, N20329, N1461);
not NOT1 (N20348, N20338);
nand NAND3 (N20349, N20345, N6667, N10362);
and AND3 (N20350, N20332, N4856, N13931);
nor NOR3 (N20351, N20350, N19642, N12382);
not NOT1 (N20352, N20339);
and AND3 (N20353, N20344, N9898, N789);
nor NOR3 (N20354, N20352, N12013, N16820);
xor XOR2 (N20355, N20353, N3553);
and AND4 (N20356, N20351, N16984, N18376, N4173);
not NOT1 (N20357, N20346);
not NOT1 (N20358, N20347);
buf BUF1 (N20359, N20348);
buf BUF1 (N20360, N20349);
xor XOR2 (N20361, N20354, N647);
nor NOR4 (N20362, N20360, N5893, N2461, N5994);
nand NAND2 (N20363, N20357, N12136);
xor XOR2 (N20364, N20358, N14934);
buf BUF1 (N20365, N20355);
buf BUF1 (N20366, N20356);
not NOT1 (N20367, N20283);
or OR3 (N20368, N20359, N9507, N1584);
nor NOR3 (N20369, N20361, N17763, N18931);
nand NAND4 (N20370, N20364, N7158, N4853, N10342);
nor NOR2 (N20371, N20370, N6323);
nor NOR4 (N20372, N20367, N10952, N11641, N17637);
and AND3 (N20373, N20372, N10218, N13853);
not NOT1 (N20374, N20369);
buf BUF1 (N20375, N20365);
buf BUF1 (N20376, N20362);
or OR3 (N20377, N20301, N12786, N6685);
nand NAND4 (N20378, N20366, N18705, N1244, N14274);
and AND3 (N20379, N20368, N17574, N5868);
and AND2 (N20380, N20374, N2521);
nor NOR2 (N20381, N20377, N4462);
nor NOR4 (N20382, N20380, N10171, N5120, N1710);
or OR2 (N20383, N20371, N11694);
not NOT1 (N20384, N20378);
nor NOR4 (N20385, N20383, N11137, N4369, N2026);
and AND3 (N20386, N20379, N8944, N11667);
buf BUF1 (N20387, N20373);
xor XOR2 (N20388, N20386, N9944);
nand NAND4 (N20389, N20376, N13697, N1721, N20338);
nor NOR3 (N20390, N20375, N5574, N1305);
or OR3 (N20391, N20389, N13447, N19477);
and AND4 (N20392, N20382, N630, N15403, N3541);
buf BUF1 (N20393, N20343);
xor XOR2 (N20394, N20384, N6162);
not NOT1 (N20395, N20394);
not NOT1 (N20396, N20363);
nor NOR2 (N20397, N20387, N5264);
buf BUF1 (N20398, N20393);
not NOT1 (N20399, N20391);
xor XOR2 (N20400, N20399, N16677);
nand NAND2 (N20401, N20385, N6805);
buf BUF1 (N20402, N20397);
or OR2 (N20403, N20401, N3923);
not NOT1 (N20404, N20400);
and AND3 (N20405, N20390, N11308, N9360);
nand NAND3 (N20406, N20404, N4618, N4801);
buf BUF1 (N20407, N20405);
nor NOR4 (N20408, N20381, N4668, N7401, N8140);
nor NOR3 (N20409, N20407, N19505, N17424);
and AND3 (N20410, N20388, N1531, N6153);
not NOT1 (N20411, N20398);
nor NOR2 (N20412, N20409, N554);
or OR4 (N20413, N20412, N12644, N8745, N2191);
and AND4 (N20414, N20395, N1591, N18184, N11287);
buf BUF1 (N20415, N20413);
not NOT1 (N20416, N20392);
nor NOR4 (N20417, N20411, N6963, N14607, N2186);
not NOT1 (N20418, N20416);
nor NOR3 (N20419, N20418, N8813, N15524);
or OR4 (N20420, N20419, N1862, N12313, N20166);
nor NOR2 (N20421, N20406, N13744);
xor XOR2 (N20422, N20396, N17671);
or OR4 (N20423, N20402, N12329, N11834, N3010);
nand NAND2 (N20424, N20410, N2080);
and AND4 (N20425, N20424, N6910, N4598, N10178);
and AND4 (N20426, N20421, N13118, N9714, N12738);
nand NAND4 (N20427, N20423, N17414, N10690, N10743);
nor NOR2 (N20428, N20408, N17645);
buf BUF1 (N20429, N20414);
xor XOR2 (N20430, N20428, N3436);
buf BUF1 (N20431, N20426);
buf BUF1 (N20432, N20415);
xor XOR2 (N20433, N20403, N5117);
and AND3 (N20434, N20420, N16528, N11150);
and AND3 (N20435, N20425, N6069, N7587);
not NOT1 (N20436, N20433);
xor XOR2 (N20437, N20422, N15938);
nand NAND4 (N20438, N20435, N17062, N10926, N1193);
nor NOR2 (N20439, N20417, N12012);
not NOT1 (N20440, N20429);
not NOT1 (N20441, N20431);
nor NOR2 (N20442, N20434, N15327);
buf BUF1 (N20443, N20437);
nand NAND2 (N20444, N20432, N296);
nand NAND3 (N20445, N20442, N739, N17733);
and AND4 (N20446, N20444, N9554, N432, N10994);
nand NAND4 (N20447, N20439, N12844, N8283, N15298);
or OR4 (N20448, N20441, N4476, N19756, N7051);
not NOT1 (N20449, N20443);
or OR3 (N20450, N20427, N14759, N12313);
buf BUF1 (N20451, N20447);
nor NOR2 (N20452, N20451, N19004);
and AND2 (N20453, N20430, N16057);
or OR3 (N20454, N20438, N18779, N18411);
and AND4 (N20455, N20448, N1934, N15321, N13876);
nor NOR4 (N20456, N20446, N18878, N17968, N18426);
buf BUF1 (N20457, N20436);
or OR2 (N20458, N20450, N1799);
not NOT1 (N20459, N20449);
buf BUF1 (N20460, N20440);
buf BUF1 (N20461, N20445);
not NOT1 (N20462, N20454);
nor NOR4 (N20463, N20456, N9405, N1093, N15289);
or OR2 (N20464, N20457, N877);
nand NAND2 (N20465, N20464, N12226);
or OR3 (N20466, N20455, N665, N6060);
nand NAND4 (N20467, N20452, N3191, N11529, N3805);
xor XOR2 (N20468, N20460, N19998);
and AND3 (N20469, N20468, N8482, N19055);
nand NAND3 (N20470, N20458, N17413, N10732);
nand NAND2 (N20471, N20459, N19453);
and AND2 (N20472, N20463, N16173);
and AND3 (N20473, N20472, N14064, N10865);
nand NAND2 (N20474, N20470, N13138);
and AND3 (N20475, N20467, N9818, N19913);
and AND2 (N20476, N20473, N19076);
nor NOR4 (N20477, N20469, N15904, N10603, N8442);
nand NAND4 (N20478, N20465, N9768, N10371, N4752);
buf BUF1 (N20479, N20461);
or OR2 (N20480, N20476, N12412);
and AND2 (N20481, N20453, N9943);
buf BUF1 (N20482, N20481);
and AND3 (N20483, N20471, N9073, N14626);
buf BUF1 (N20484, N20479);
and AND3 (N20485, N20475, N7341, N18384);
and AND2 (N20486, N20480, N14936);
nand NAND3 (N20487, N20474, N3625, N16073);
not NOT1 (N20488, N20485);
buf BUF1 (N20489, N20483);
buf BUF1 (N20490, N20488);
not NOT1 (N20491, N20466);
xor XOR2 (N20492, N20489, N2774);
buf BUF1 (N20493, N20484);
nor NOR4 (N20494, N20477, N7532, N4933, N195);
or OR4 (N20495, N20486, N5696, N4872, N16532);
or OR3 (N20496, N20494, N18183, N3082);
or OR3 (N20497, N20487, N1783, N12032);
xor XOR2 (N20498, N20492, N12059);
buf BUF1 (N20499, N20462);
and AND3 (N20500, N20490, N18733, N1053);
or OR3 (N20501, N20496, N18561, N8063);
nand NAND4 (N20502, N20499, N1285, N4647, N6146);
xor XOR2 (N20503, N20495, N3366);
nor NOR4 (N20504, N20493, N17098, N12538, N15971);
xor XOR2 (N20505, N20500, N2535);
not NOT1 (N20506, N20505);
and AND3 (N20507, N20502, N15028, N10391);
xor XOR2 (N20508, N20497, N12338);
and AND4 (N20509, N20498, N8308, N3339, N2224);
nand NAND3 (N20510, N20507, N2647, N13640);
and AND4 (N20511, N20509, N10165, N14668, N10887);
nand NAND2 (N20512, N20511, N5534);
not NOT1 (N20513, N20501);
buf BUF1 (N20514, N20478);
and AND4 (N20515, N20482, N12826, N19882, N14065);
nand NAND3 (N20516, N20512, N9917, N7237);
nor NOR2 (N20517, N20515, N12481);
buf BUF1 (N20518, N20510);
nand NAND3 (N20519, N20517, N18155, N8217);
not NOT1 (N20520, N20516);
xor XOR2 (N20521, N20506, N18949);
or OR3 (N20522, N20519, N12174, N19102);
xor XOR2 (N20523, N20513, N19360);
xor XOR2 (N20524, N20523, N6132);
nand NAND2 (N20525, N20504, N2979);
buf BUF1 (N20526, N20491);
or OR2 (N20527, N20522, N11304);
xor XOR2 (N20528, N20520, N15907);
buf BUF1 (N20529, N20503);
nand NAND2 (N20530, N20521, N5551);
buf BUF1 (N20531, N20527);
or OR4 (N20532, N20525, N8214, N8072, N12433);
buf BUF1 (N20533, N20529);
xor XOR2 (N20534, N20531, N9860);
xor XOR2 (N20535, N20526, N20494);
not NOT1 (N20536, N20518);
xor XOR2 (N20537, N20508, N15431);
buf BUF1 (N20538, N20528);
xor XOR2 (N20539, N20533, N9532);
xor XOR2 (N20540, N20535, N2919);
nor NOR4 (N20541, N20540, N16846, N4302, N6562);
xor XOR2 (N20542, N20536, N15006);
nand NAND4 (N20543, N20539, N19031, N20187, N20128);
not NOT1 (N20544, N20541);
buf BUF1 (N20545, N20514);
buf BUF1 (N20546, N20544);
nand NAND3 (N20547, N20546, N4804, N16398);
xor XOR2 (N20548, N20530, N6838);
and AND3 (N20549, N20548, N3388, N11621);
not NOT1 (N20550, N20547);
xor XOR2 (N20551, N20534, N17465);
xor XOR2 (N20552, N20532, N3643);
xor XOR2 (N20553, N20542, N17016);
and AND4 (N20554, N20551, N7469, N9722, N12019);
buf BUF1 (N20555, N20538);
and AND4 (N20556, N20543, N13967, N11265, N12130);
nor NOR4 (N20557, N20556, N4650, N4885, N14763);
nor NOR3 (N20558, N20552, N6657, N1155);
not NOT1 (N20559, N20553);
not NOT1 (N20560, N20559);
not NOT1 (N20561, N20554);
xor XOR2 (N20562, N20545, N17606);
nand NAND3 (N20563, N20561, N1594, N6911);
and AND4 (N20564, N20558, N16442, N6673, N7692);
buf BUF1 (N20565, N20524);
buf BUF1 (N20566, N20562);
not NOT1 (N20567, N20555);
and AND3 (N20568, N20549, N14141, N4964);
buf BUF1 (N20569, N20563);
and AND3 (N20570, N20566, N10383, N3757);
buf BUF1 (N20571, N20570);
nand NAND4 (N20572, N20569, N2451, N13057, N12500);
nand NAND4 (N20573, N20571, N4371, N12483, N17375);
not NOT1 (N20574, N20537);
nand NAND4 (N20575, N20574, N20074, N20451, N18513);
nor NOR3 (N20576, N20565, N1560, N19712);
buf BUF1 (N20577, N20568);
nand NAND3 (N20578, N20567, N5691, N18277);
nor NOR4 (N20579, N20578, N18546, N13476, N13046);
nor NOR2 (N20580, N20575, N14991);
or OR2 (N20581, N20577, N2229);
xor XOR2 (N20582, N20557, N7859);
xor XOR2 (N20583, N20580, N15836);
xor XOR2 (N20584, N20579, N14896);
nand NAND4 (N20585, N20576, N14853, N5701, N12845);
nor NOR3 (N20586, N20572, N10400, N14181);
and AND4 (N20587, N20550, N3548, N15716, N17054);
or OR2 (N20588, N20581, N5574);
and AND3 (N20589, N20585, N9651, N20072);
nor NOR4 (N20590, N20582, N19337, N17741, N5115);
and AND4 (N20591, N20588, N8872, N11053, N3554);
xor XOR2 (N20592, N20584, N488);
not NOT1 (N20593, N20564);
nor NOR2 (N20594, N20586, N233);
or OR3 (N20595, N20594, N3885, N12324);
or OR4 (N20596, N20583, N13511, N16506, N3446);
nand NAND3 (N20597, N20596, N16605, N7264);
nor NOR2 (N20598, N20593, N12794);
or OR2 (N20599, N20587, N17977);
nor NOR2 (N20600, N20595, N4563);
buf BUF1 (N20601, N20590);
nor NOR2 (N20602, N20601, N12983);
xor XOR2 (N20603, N20589, N3931);
and AND3 (N20604, N20592, N13296, N8896);
or OR4 (N20605, N20600, N11070, N4728, N239);
buf BUF1 (N20606, N20603);
nand NAND4 (N20607, N20602, N7011, N12330, N20594);
or OR4 (N20608, N20597, N12158, N9510, N16986);
buf BUF1 (N20609, N20608);
or OR3 (N20610, N20598, N19040, N11449);
nor NOR4 (N20611, N20605, N19175, N4203, N5118);
xor XOR2 (N20612, N20611, N19092);
nand NAND4 (N20613, N20604, N8231, N11649, N1527);
nand NAND3 (N20614, N20612, N20146, N3821);
and AND2 (N20615, N20613, N8525);
nor NOR4 (N20616, N20591, N9544, N3490, N11024);
not NOT1 (N20617, N20573);
buf BUF1 (N20618, N20614);
and AND3 (N20619, N20615, N11851, N15472);
and AND2 (N20620, N20606, N17326);
xor XOR2 (N20621, N20599, N15767);
nor NOR4 (N20622, N20610, N16568, N6111, N16698);
or OR2 (N20623, N20620, N6085);
and AND4 (N20624, N20622, N15655, N689, N6768);
or OR3 (N20625, N20621, N302, N17244);
or OR4 (N20626, N20609, N354, N11922, N17780);
xor XOR2 (N20627, N20616, N2594);
xor XOR2 (N20628, N20607, N15942);
nor NOR2 (N20629, N20626, N14482);
or OR4 (N20630, N20624, N7913, N14939, N16599);
xor XOR2 (N20631, N20625, N11717);
buf BUF1 (N20632, N20617);
nand NAND2 (N20633, N20629, N1360);
or OR2 (N20634, N20627, N14905);
or OR4 (N20635, N20632, N4410, N15391, N9548);
buf BUF1 (N20636, N20560);
not NOT1 (N20637, N20628);
nor NOR4 (N20638, N20634, N4356, N2888, N18845);
nor NOR3 (N20639, N20619, N1301, N8291);
xor XOR2 (N20640, N20631, N19503);
or OR2 (N20641, N20618, N16600);
nor NOR3 (N20642, N20640, N12878, N16083);
nand NAND2 (N20643, N20633, N15907);
nor NOR2 (N20644, N20638, N9770);
buf BUF1 (N20645, N20644);
buf BUF1 (N20646, N20642);
nor NOR4 (N20647, N20643, N13596, N16857, N1745);
nand NAND4 (N20648, N20630, N15997, N12854, N11680);
nand NAND3 (N20649, N20641, N229, N14998);
nor NOR3 (N20650, N20647, N14004, N12489);
not NOT1 (N20651, N20646);
nand NAND3 (N20652, N20645, N5113, N14404);
nand NAND4 (N20653, N20652, N16042, N8846, N8028);
buf BUF1 (N20654, N20637);
and AND3 (N20655, N20636, N8213, N6198);
nand NAND4 (N20656, N20650, N1644, N11960, N18756);
xor XOR2 (N20657, N20654, N2347);
not NOT1 (N20658, N20649);
and AND4 (N20659, N20653, N6055, N16969, N16372);
not NOT1 (N20660, N20655);
nor NOR4 (N20661, N20658, N15040, N14021, N12524);
buf BUF1 (N20662, N20660);
nor NOR3 (N20663, N20661, N2295, N16872);
not NOT1 (N20664, N20663);
buf BUF1 (N20665, N20657);
xor XOR2 (N20666, N20648, N11237);
or OR3 (N20667, N20639, N6454, N14920);
nand NAND4 (N20668, N20651, N628, N14137, N6824);
buf BUF1 (N20669, N20667);
nor NOR2 (N20670, N20665, N1035);
nand NAND3 (N20671, N20635, N19201, N12783);
and AND4 (N20672, N20670, N6424, N20048, N522);
nor NOR4 (N20673, N20664, N16218, N4559, N6002);
and AND3 (N20674, N20668, N15143, N19856);
nor NOR2 (N20675, N20656, N13059);
nor NOR2 (N20676, N20659, N3974);
or OR4 (N20677, N20669, N10501, N16785, N16701);
nand NAND4 (N20678, N20671, N3859, N12930, N15122);
buf BUF1 (N20679, N20677);
nor NOR2 (N20680, N20662, N10460);
nor NOR4 (N20681, N20680, N19705, N12237, N4547);
and AND3 (N20682, N20672, N18387, N15909);
not NOT1 (N20683, N20682);
nand NAND3 (N20684, N20679, N12971, N1503);
buf BUF1 (N20685, N20673);
nor NOR3 (N20686, N20666, N16438, N1725);
buf BUF1 (N20687, N20681);
xor XOR2 (N20688, N20678, N19838);
xor XOR2 (N20689, N20686, N18827);
xor XOR2 (N20690, N20687, N1642);
nand NAND2 (N20691, N20683, N16450);
not NOT1 (N20692, N20688);
or OR2 (N20693, N20684, N14591);
nor NOR3 (N20694, N20693, N19786, N3552);
nor NOR4 (N20695, N20692, N1602, N12828, N14368);
or OR2 (N20696, N20690, N11224);
and AND4 (N20697, N20694, N3386, N16170, N10164);
nor NOR2 (N20698, N20623, N16938);
buf BUF1 (N20699, N20696);
or OR2 (N20700, N20697, N20443);
not NOT1 (N20701, N20691);
not NOT1 (N20702, N20695);
and AND2 (N20703, N20676, N19508);
nor NOR2 (N20704, N20702, N2506);
or OR4 (N20705, N20674, N17373, N18073, N14100);
xor XOR2 (N20706, N20701, N10265);
nand NAND4 (N20707, N20689, N5235, N13966, N436);
and AND3 (N20708, N20703, N10875, N2577);
not NOT1 (N20709, N20698);
and AND3 (N20710, N20704, N16060, N16446);
xor XOR2 (N20711, N20707, N15671);
nand NAND3 (N20712, N20708, N442, N9990);
nor NOR2 (N20713, N20712, N16381);
not NOT1 (N20714, N20713);
nor NOR2 (N20715, N20685, N1694);
nor NOR3 (N20716, N20706, N14542, N14989);
buf BUF1 (N20717, N20705);
buf BUF1 (N20718, N20711);
xor XOR2 (N20719, N20715, N20458);
nor NOR4 (N20720, N20710, N7322, N18264, N15881);
nor NOR2 (N20721, N20714, N19675);
and AND2 (N20722, N20700, N18074);
nand NAND2 (N20723, N20722, N3202);
not NOT1 (N20724, N20699);
buf BUF1 (N20725, N20721);
xor XOR2 (N20726, N20716, N13225);
or OR2 (N20727, N20720, N15422);
nand NAND2 (N20728, N20717, N18257);
and AND4 (N20729, N20725, N11738, N19805, N911);
nor NOR4 (N20730, N20718, N413, N6304, N18369);
not NOT1 (N20731, N20724);
nand NAND4 (N20732, N20719, N13626, N19036, N11369);
xor XOR2 (N20733, N20726, N1788);
and AND2 (N20734, N20728, N5112);
nor NOR4 (N20735, N20730, N10668, N3171, N3433);
or OR2 (N20736, N20732, N3753);
and AND3 (N20737, N20709, N14453, N11719);
nand NAND3 (N20738, N20733, N17735, N19758);
xor XOR2 (N20739, N20737, N2657);
buf BUF1 (N20740, N20729);
not NOT1 (N20741, N20735);
nand NAND3 (N20742, N20740, N18539, N660);
and AND2 (N20743, N20734, N10038);
not NOT1 (N20744, N20739);
xor XOR2 (N20745, N20741, N15800);
nor NOR2 (N20746, N20738, N7332);
and AND2 (N20747, N20744, N5048);
or OR3 (N20748, N20731, N16694, N1814);
xor XOR2 (N20749, N20736, N10530);
not NOT1 (N20750, N20727);
or OR4 (N20751, N20742, N14798, N10533, N19130);
or OR4 (N20752, N20750, N14396, N11069, N19714);
xor XOR2 (N20753, N20675, N6840);
nor NOR2 (N20754, N20753, N3355);
not NOT1 (N20755, N20745);
or OR2 (N20756, N20755, N18435);
nor NOR2 (N20757, N20743, N17838);
nand NAND3 (N20758, N20723, N18094, N8075);
nand NAND3 (N20759, N20746, N16174, N7703);
buf BUF1 (N20760, N20747);
buf BUF1 (N20761, N20758);
xor XOR2 (N20762, N20748, N14177);
xor XOR2 (N20763, N20756, N12682);
nor NOR3 (N20764, N20759, N13659, N4116);
not NOT1 (N20765, N20761);
and AND4 (N20766, N20760, N5006, N13466, N20537);
nand NAND3 (N20767, N20751, N8412, N14211);
or OR4 (N20768, N20762, N17948, N988, N15548);
and AND3 (N20769, N20749, N2717, N6258);
and AND3 (N20770, N20752, N13702, N8824);
buf BUF1 (N20771, N20769);
xor XOR2 (N20772, N20768, N16420);
nor NOR4 (N20773, N20771, N4052, N748, N14684);
or OR4 (N20774, N20764, N17203, N13947, N3747);
nor NOR3 (N20775, N20757, N11942, N1017);
nor NOR4 (N20776, N20772, N3158, N828, N7098);
not NOT1 (N20777, N20766);
nand NAND3 (N20778, N20763, N6398, N2185);
or OR3 (N20779, N20776, N18895, N11809);
not NOT1 (N20780, N20774);
or OR4 (N20781, N20773, N7315, N6586, N6159);
nand NAND4 (N20782, N20778, N790, N10480, N5369);
buf BUF1 (N20783, N20779);
nand NAND2 (N20784, N20775, N1319);
nor NOR2 (N20785, N20765, N20759);
nand NAND3 (N20786, N20781, N5651, N16024);
not NOT1 (N20787, N20777);
nor NOR4 (N20788, N20784, N14124, N20062, N763);
xor XOR2 (N20789, N20767, N11097);
nand NAND4 (N20790, N20787, N916, N15571, N17426);
or OR3 (N20791, N20782, N3900, N114);
or OR2 (N20792, N20791, N545);
nor NOR3 (N20793, N20770, N5366, N10825);
or OR2 (N20794, N20790, N11918);
nand NAND2 (N20795, N20789, N14848);
buf BUF1 (N20796, N20786);
or OR4 (N20797, N20794, N1850, N18289, N4757);
not NOT1 (N20798, N20792);
buf BUF1 (N20799, N20754);
or OR2 (N20800, N20796, N19023);
nor NOR4 (N20801, N20798, N733, N10552, N14463);
buf BUF1 (N20802, N20793);
nor NOR4 (N20803, N20799, N1745, N7014, N3352);
and AND3 (N20804, N20800, N7893, N17191);
xor XOR2 (N20805, N20795, N14456);
nor NOR3 (N20806, N20780, N6330, N19481);
buf BUF1 (N20807, N20802);
and AND3 (N20808, N20788, N11474, N19478);
nor NOR2 (N20809, N20807, N9832);
or OR3 (N20810, N20803, N6932, N12271);
and AND4 (N20811, N20804, N4884, N11513, N2359);
not NOT1 (N20812, N20810);
nand NAND3 (N20813, N20797, N13103, N15317);
or OR2 (N20814, N20805, N14228);
not NOT1 (N20815, N20814);
nand NAND4 (N20816, N20809, N7700, N11250, N13922);
and AND2 (N20817, N20811, N8296);
nand NAND2 (N20818, N20815, N12580);
xor XOR2 (N20819, N20812, N5032);
xor XOR2 (N20820, N20813, N10202);
nor NOR2 (N20821, N20783, N18699);
buf BUF1 (N20822, N20816);
buf BUF1 (N20823, N20822);
nor NOR2 (N20824, N20817, N6070);
nand NAND2 (N20825, N20824, N11776);
buf BUF1 (N20826, N20808);
buf BUF1 (N20827, N20785);
or OR3 (N20828, N20821, N14770, N6589);
nor NOR3 (N20829, N20826, N4271, N19462);
buf BUF1 (N20830, N20827);
nor NOR2 (N20831, N20818, N17301);
nor NOR4 (N20832, N20820, N7066, N12271, N6788);
nor NOR4 (N20833, N20832, N19164, N1917, N2877);
or OR2 (N20834, N20829, N16310);
xor XOR2 (N20835, N20806, N529);
and AND2 (N20836, N20801, N6819);
or OR2 (N20837, N20823, N4996);
not NOT1 (N20838, N20825);
nand NAND3 (N20839, N20838, N18070, N7123);
and AND2 (N20840, N20831, N5744);
and AND4 (N20841, N20819, N18508, N10912, N18434);
nor NOR4 (N20842, N20841, N14687, N7784, N11844);
or OR2 (N20843, N20837, N19981);
not NOT1 (N20844, N20835);
nor NOR3 (N20845, N20836, N7893, N13337);
nor NOR3 (N20846, N20834, N2446, N10725);
nor NOR3 (N20847, N20844, N3678, N16550);
nor NOR2 (N20848, N20843, N12041);
buf BUF1 (N20849, N20842);
buf BUF1 (N20850, N20839);
xor XOR2 (N20851, N20830, N3954);
or OR3 (N20852, N20828, N14062, N16151);
nand NAND2 (N20853, N20833, N7323);
or OR2 (N20854, N20849, N13659);
buf BUF1 (N20855, N20840);
xor XOR2 (N20856, N20845, N10505);
buf BUF1 (N20857, N20847);
buf BUF1 (N20858, N20855);
nor NOR3 (N20859, N20852, N2871, N9218);
nand NAND2 (N20860, N20857, N4106);
or OR3 (N20861, N20854, N17618, N2144);
nor NOR2 (N20862, N20848, N13305);
xor XOR2 (N20863, N20853, N13331);
nand NAND2 (N20864, N20858, N5369);
not NOT1 (N20865, N20851);
nand NAND3 (N20866, N20861, N4485, N15996);
not NOT1 (N20867, N20860);
or OR2 (N20868, N20862, N12006);
nor NOR4 (N20869, N20867, N11767, N6799, N17713);
nor NOR3 (N20870, N20863, N16048, N13886);
xor XOR2 (N20871, N20859, N5718);
and AND3 (N20872, N20866, N7710, N9563);
xor XOR2 (N20873, N20864, N6521);
nand NAND2 (N20874, N20873, N1482);
or OR4 (N20875, N20850, N13429, N4679, N7625);
and AND4 (N20876, N20872, N16715, N2890, N8748);
buf BUF1 (N20877, N20875);
xor XOR2 (N20878, N20869, N10739);
or OR2 (N20879, N20871, N19829);
xor XOR2 (N20880, N20870, N4920);
nor NOR3 (N20881, N20868, N19126, N2419);
buf BUF1 (N20882, N20881);
nor NOR3 (N20883, N20846, N20556, N15710);
and AND3 (N20884, N20856, N13826, N19366);
nand NAND3 (N20885, N20882, N16512, N11948);
not NOT1 (N20886, N20865);
xor XOR2 (N20887, N20886, N16067);
and AND3 (N20888, N20878, N15964, N3183);
or OR4 (N20889, N20883, N8625, N2226, N13608);
buf BUF1 (N20890, N20879);
and AND4 (N20891, N20889, N16870, N16273, N18583);
not NOT1 (N20892, N20877);
nand NAND3 (N20893, N20874, N8956, N17256);
nand NAND4 (N20894, N20891, N17956, N9887, N9606);
xor XOR2 (N20895, N20885, N10820);
nor NOR2 (N20896, N20888, N20757);
not NOT1 (N20897, N20884);
or OR4 (N20898, N20893, N15346, N715, N17949);
nand NAND3 (N20899, N20894, N11946, N2805);
nand NAND2 (N20900, N20897, N2253);
xor XOR2 (N20901, N20892, N3765);
and AND3 (N20902, N20896, N802, N11798);
not NOT1 (N20903, N20887);
buf BUF1 (N20904, N20898);
buf BUF1 (N20905, N20902);
and AND3 (N20906, N20905, N6942, N1568);
xor XOR2 (N20907, N20876, N19177);
xor XOR2 (N20908, N20904, N10151);
or OR3 (N20909, N20895, N6191, N15750);
nor NOR3 (N20910, N20906, N11910, N2504);
not NOT1 (N20911, N20908);
xor XOR2 (N20912, N20909, N20575);
not NOT1 (N20913, N20901);
and AND3 (N20914, N20890, N11584, N2513);
not NOT1 (N20915, N20911);
not NOT1 (N20916, N20900);
buf BUF1 (N20917, N20903);
nor NOR3 (N20918, N20914, N16656, N12783);
not NOT1 (N20919, N20917);
nand NAND4 (N20920, N20907, N13029, N17337, N5898);
not NOT1 (N20921, N20899);
or OR4 (N20922, N20912, N14670, N1197, N8371);
and AND2 (N20923, N20910, N14407);
nor NOR4 (N20924, N20913, N448, N14831, N6196);
nand NAND4 (N20925, N20924, N5527, N10719, N11228);
nor NOR2 (N20926, N20925, N9213);
not NOT1 (N20927, N20919);
nor NOR3 (N20928, N20927, N20908, N6554);
and AND3 (N20929, N20880, N11544, N4763);
or OR2 (N20930, N20918, N5368);
or OR4 (N20931, N20915, N12774, N19209, N338);
xor XOR2 (N20932, N20922, N17192);
or OR4 (N20933, N20916, N14322, N7942, N14247);
nand NAND2 (N20934, N20923, N15797);
nand NAND3 (N20935, N20931, N12335, N1722);
and AND3 (N20936, N20933, N16717, N16907);
nand NAND4 (N20937, N20928, N18951, N2213, N19896);
or OR3 (N20938, N20920, N20459, N11368);
or OR4 (N20939, N20929, N11549, N16081, N16443);
or OR3 (N20940, N20930, N3464, N7766);
nand NAND3 (N20941, N20938, N9095, N10434);
not NOT1 (N20942, N20935);
not NOT1 (N20943, N20939);
xor XOR2 (N20944, N20926, N1430);
not NOT1 (N20945, N20936);
xor XOR2 (N20946, N20944, N10689);
buf BUF1 (N20947, N20937);
not NOT1 (N20948, N20945);
nand NAND2 (N20949, N20948, N2836);
or OR2 (N20950, N20946, N7722);
and AND2 (N20951, N20921, N1409);
not NOT1 (N20952, N20949);
nor NOR4 (N20953, N20941, N14531, N10817, N1565);
not NOT1 (N20954, N20952);
nand NAND4 (N20955, N20943, N3849, N5674, N15394);
buf BUF1 (N20956, N20934);
or OR4 (N20957, N20932, N9668, N1247, N12964);
not NOT1 (N20958, N20940);
nor NOR2 (N20959, N20947, N12459);
not NOT1 (N20960, N20950);
xor XOR2 (N20961, N20953, N6747);
not NOT1 (N20962, N20955);
nand NAND3 (N20963, N20956, N7366, N3268);
nor NOR3 (N20964, N20963, N3769, N13222);
nor NOR3 (N20965, N20961, N11808, N20702);
and AND4 (N20966, N20962, N5548, N12902, N3178);
nor NOR2 (N20967, N20954, N6767);
nand NAND4 (N20968, N20958, N15524, N13788, N7131);
and AND3 (N20969, N20959, N18257, N2089);
nand NAND4 (N20970, N20951, N5299, N1452, N13286);
or OR3 (N20971, N20965, N7201, N2219);
and AND2 (N20972, N20966, N19192);
buf BUF1 (N20973, N20971);
nand NAND2 (N20974, N20967, N20424);
or OR3 (N20975, N20957, N6242, N15199);
and AND4 (N20976, N20973, N15040, N11334, N11669);
xor XOR2 (N20977, N20968, N4330);
not NOT1 (N20978, N20975);
and AND3 (N20979, N20976, N17699, N9833);
nand NAND4 (N20980, N20964, N4237, N20099, N8083);
nand NAND4 (N20981, N20978, N12789, N7943, N2746);
nand NAND3 (N20982, N20977, N2820, N14044);
xor XOR2 (N20983, N20970, N6049);
or OR2 (N20984, N20942, N17112);
or OR4 (N20985, N20974, N14894, N13861, N9788);
or OR4 (N20986, N20983, N11164, N13980, N10322);
and AND2 (N20987, N20984, N17432);
xor XOR2 (N20988, N20979, N12982);
nor NOR2 (N20989, N20969, N17084);
or OR4 (N20990, N20981, N20517, N15321, N20093);
and AND4 (N20991, N20990, N17021, N13416, N3370);
or OR4 (N20992, N20989, N14864, N421, N9673);
not NOT1 (N20993, N20992);
buf BUF1 (N20994, N20960);
nand NAND3 (N20995, N20980, N13191, N3520);
or OR2 (N20996, N20995, N3834);
or OR3 (N20997, N20991, N16200, N12861);
nand NAND3 (N20998, N20986, N20780, N19508);
xor XOR2 (N20999, N20982, N7302);
buf BUF1 (N21000, N20988);
and AND4 (N21001, N20996, N11997, N16049, N13562);
nor NOR3 (N21002, N20999, N4920, N14702);
or OR4 (N21003, N20998, N16132, N9513, N8607);
xor XOR2 (N21004, N21002, N20874);
or OR4 (N21005, N20997, N15896, N2955, N15647);
nor NOR2 (N21006, N21001, N11194);
and AND2 (N21007, N21004, N1111);
or OR2 (N21008, N21007, N10312);
xor XOR2 (N21009, N20994, N18231);
nand NAND3 (N21010, N21003, N263, N2462);
and AND2 (N21011, N21000, N47);
nand NAND3 (N21012, N20972, N15379, N4993);
buf BUF1 (N21013, N21009);
xor XOR2 (N21014, N21008, N1983);
or OR4 (N21015, N21011, N11505, N17874, N4917);
nand NAND2 (N21016, N21010, N8218);
xor XOR2 (N21017, N21015, N18846);
buf BUF1 (N21018, N21014);
buf BUF1 (N21019, N21005);
nor NOR2 (N21020, N21019, N1493);
and AND3 (N21021, N21020, N4835, N3116);
not NOT1 (N21022, N21006);
not NOT1 (N21023, N20985);
buf BUF1 (N21024, N21022);
buf BUF1 (N21025, N21024);
nor NOR4 (N21026, N21017, N14682, N8671, N13324);
not NOT1 (N21027, N21013);
xor XOR2 (N21028, N21021, N10047);
or OR2 (N21029, N21027, N13033);
buf BUF1 (N21030, N21025);
xor XOR2 (N21031, N21012, N3284);
or OR3 (N21032, N20993, N10634, N6276);
nor NOR3 (N21033, N21023, N15437, N1869);
nor NOR2 (N21034, N21018, N6396);
or OR2 (N21035, N21026, N19745);
and AND4 (N21036, N20987, N3794, N8284, N18601);
buf BUF1 (N21037, N21032);
nand NAND3 (N21038, N21016, N12042, N12094);
nand NAND3 (N21039, N21037, N387, N9462);
and AND3 (N21040, N21031, N14441, N8858);
xor XOR2 (N21041, N21034, N18547);
and AND3 (N21042, N21030, N17354, N15147);
or OR4 (N21043, N21042, N7050, N7139, N1196);
or OR4 (N21044, N21028, N16188, N10800, N9661);
and AND2 (N21045, N21029, N8933);
not NOT1 (N21046, N21044);
and AND2 (N21047, N21040, N12965);
nand NAND4 (N21048, N21043, N1296, N12996, N8843);
or OR2 (N21049, N21033, N16004);
and AND3 (N21050, N21045, N6306, N18533);
or OR3 (N21051, N21036, N17692, N2350);
nor NOR2 (N21052, N21041, N8515);
or OR2 (N21053, N21047, N587);
and AND4 (N21054, N21039, N4962, N12270, N20211);
and AND4 (N21055, N21046, N2476, N18459, N14380);
not NOT1 (N21056, N21048);
nor NOR2 (N21057, N21056, N9516);
nor NOR3 (N21058, N21055, N2277, N9816);
or OR3 (N21059, N21057, N4446, N1823);
not NOT1 (N21060, N21049);
not NOT1 (N21061, N21035);
buf BUF1 (N21062, N21059);
buf BUF1 (N21063, N21052);
and AND2 (N21064, N21038, N6488);
buf BUF1 (N21065, N21060);
nor NOR3 (N21066, N21065, N2320, N8873);
nand NAND3 (N21067, N21062, N11867, N10482);
xor XOR2 (N21068, N21066, N16858);
and AND2 (N21069, N21067, N18252);
xor XOR2 (N21070, N21051, N312);
buf BUF1 (N21071, N21061);
and AND3 (N21072, N21053, N7818, N20417);
and AND2 (N21073, N21069, N5694);
or OR3 (N21074, N21050, N11552, N9259);
not NOT1 (N21075, N21071);
and AND3 (N21076, N21058, N7170, N4077);
or OR2 (N21077, N21070, N19955);
or OR4 (N21078, N21054, N21034, N12325, N17344);
nand NAND4 (N21079, N21068, N526, N2589, N7295);
xor XOR2 (N21080, N21079, N20117);
nor NOR4 (N21081, N21063, N19938, N6523, N21037);
nand NAND2 (N21082, N21064, N11790);
buf BUF1 (N21083, N21082);
not NOT1 (N21084, N21077);
buf BUF1 (N21085, N21078);
buf BUF1 (N21086, N21075);
and AND2 (N21087, N21072, N6308);
nand NAND2 (N21088, N21083, N2624);
nor NOR4 (N21089, N21088, N2318, N14139, N11977);
or OR2 (N21090, N21076, N4404);
and AND2 (N21091, N21080, N20463);
nor NOR2 (N21092, N21073, N18236);
nor NOR4 (N21093, N21091, N12633, N14235, N4520);
and AND2 (N21094, N21093, N1443);
nor NOR2 (N21095, N21090, N5747);
or OR3 (N21096, N21089, N14084, N8412);
xor XOR2 (N21097, N21085, N13590);
xor XOR2 (N21098, N21092, N3808);
nor NOR3 (N21099, N21097, N18229, N4566);
not NOT1 (N21100, N21074);
and AND3 (N21101, N21087, N2329, N20039);
and AND3 (N21102, N21086, N14102, N11663);
nor NOR2 (N21103, N21081, N13639);
nand NAND3 (N21104, N21096, N12896, N1377);
nor NOR3 (N21105, N21099, N403, N17532);
or OR2 (N21106, N21101, N13590);
not NOT1 (N21107, N21095);
nor NOR3 (N21108, N21084, N919, N16707);
buf BUF1 (N21109, N21107);
nand NAND3 (N21110, N21106, N7446, N4790);
buf BUF1 (N21111, N21102);
and AND3 (N21112, N21109, N15005, N3395);
buf BUF1 (N21113, N21110);
nor NOR4 (N21114, N21094, N17769, N12864, N18150);
nor NOR4 (N21115, N21104, N1578, N4457, N7974);
and AND3 (N21116, N21105, N4615, N1485);
xor XOR2 (N21117, N21111, N8228);
nor NOR4 (N21118, N21103, N17715, N11028, N545);
and AND2 (N21119, N21118, N8053);
nand NAND4 (N21120, N21114, N6386, N5206, N7833);
and AND4 (N21121, N21120, N7579, N13850, N1844);
xor XOR2 (N21122, N21119, N9009);
not NOT1 (N21123, N21113);
nand NAND2 (N21124, N21123, N7602);
xor XOR2 (N21125, N21112, N11795);
and AND2 (N21126, N21108, N15618);
not NOT1 (N21127, N21121);
xor XOR2 (N21128, N21116, N17913);
or OR4 (N21129, N21127, N12670, N5238, N15127);
not NOT1 (N21130, N21125);
nor NOR2 (N21131, N21098, N10409);
and AND4 (N21132, N21128, N9766, N492, N20108);
buf BUF1 (N21133, N21129);
nand NAND4 (N21134, N21126, N10040, N9502, N5340);
and AND3 (N21135, N21124, N17958, N6285);
nor NOR4 (N21136, N21132, N19437, N15442, N14970);
and AND2 (N21137, N21135, N241);
and AND3 (N21138, N21130, N19314, N20194);
or OR2 (N21139, N21138, N20908);
not NOT1 (N21140, N21131);
and AND3 (N21141, N21137, N7459, N3034);
or OR3 (N21142, N21139, N8668, N3500);
and AND4 (N21143, N21122, N7125, N4424, N14443);
or OR2 (N21144, N21115, N2446);
or OR2 (N21145, N21117, N20519);
xor XOR2 (N21146, N21134, N9661);
buf BUF1 (N21147, N21146);
or OR2 (N21148, N21143, N3196);
or OR2 (N21149, N21100, N5320);
buf BUF1 (N21150, N21140);
nor NOR2 (N21151, N21136, N6553);
xor XOR2 (N21152, N21149, N3241);
nor NOR3 (N21153, N21147, N3677, N20410);
and AND2 (N21154, N21152, N20969);
xor XOR2 (N21155, N21142, N15447);
nand NAND3 (N21156, N21151, N15716, N9367);
or OR3 (N21157, N21156, N820, N14396);
nor NOR4 (N21158, N21155, N11215, N2400, N6376);
nand NAND3 (N21159, N21158, N10776, N1272);
xor XOR2 (N21160, N21159, N16263);
and AND3 (N21161, N21154, N4611, N10099);
buf BUF1 (N21162, N21133);
not NOT1 (N21163, N21161);
nor NOR3 (N21164, N21160, N647, N9618);
nor NOR2 (N21165, N21141, N20039);
nor NOR3 (N21166, N21162, N15216, N17179);
and AND2 (N21167, N21144, N13692);
nor NOR2 (N21168, N21164, N2413);
and AND4 (N21169, N21165, N18802, N5900, N10664);
not NOT1 (N21170, N21150);
buf BUF1 (N21171, N21148);
buf BUF1 (N21172, N21169);
nor NOR3 (N21173, N21166, N18053, N3795);
buf BUF1 (N21174, N21145);
nand NAND4 (N21175, N21163, N7264, N10847, N10513);
nand NAND3 (N21176, N21174, N2447, N10184);
or OR4 (N21177, N21157, N13472, N6070, N5376);
xor XOR2 (N21178, N21171, N12355);
and AND2 (N21179, N21170, N17617);
or OR3 (N21180, N21172, N968, N4355);
buf BUF1 (N21181, N21180);
xor XOR2 (N21182, N21179, N15338);
xor XOR2 (N21183, N21177, N3617);
nor NOR4 (N21184, N21168, N6176, N15401, N14714);
or OR4 (N21185, N21167, N1703, N6699, N6648);
buf BUF1 (N21186, N21184);
and AND2 (N21187, N21183, N15753);
or OR2 (N21188, N21186, N19625);
nand NAND3 (N21189, N21153, N20166, N6784);
or OR4 (N21190, N21173, N12273, N11537, N12959);
not NOT1 (N21191, N21175);
not NOT1 (N21192, N21185);
and AND3 (N21193, N21178, N5627, N7475);
buf BUF1 (N21194, N21192);
xor XOR2 (N21195, N21181, N12900);
not NOT1 (N21196, N21193);
nand NAND4 (N21197, N21182, N12741, N123, N10971);
nor NOR4 (N21198, N21197, N1427, N252, N18788);
xor XOR2 (N21199, N21176, N10822);
xor XOR2 (N21200, N21199, N4472);
nor NOR4 (N21201, N21188, N16381, N5751, N6397);
or OR4 (N21202, N21198, N10411, N1997, N3944);
nand NAND3 (N21203, N21196, N3504, N3860);
and AND2 (N21204, N21195, N14);
nand NAND4 (N21205, N21202, N11240, N13901, N2841);
nand NAND2 (N21206, N21187, N13977);
and AND3 (N21207, N21201, N2425, N7705);
nor NOR2 (N21208, N21189, N17640);
and AND3 (N21209, N21205, N15291, N18499);
xor XOR2 (N21210, N21204, N1104);
or OR3 (N21211, N21190, N14361, N11653);
or OR2 (N21212, N21200, N5461);
nand NAND4 (N21213, N21203, N8239, N18283, N5108);
buf BUF1 (N21214, N21209);
or OR3 (N21215, N21208, N6579, N10300);
not NOT1 (N21216, N21191);
nand NAND3 (N21217, N21211, N3154, N2593);
nand NAND3 (N21218, N21215, N19479, N12098);
not NOT1 (N21219, N21212);
not NOT1 (N21220, N21214);
and AND2 (N21221, N21207, N6067);
and AND4 (N21222, N21194, N14358, N343, N11262);
nand NAND4 (N21223, N21219, N4502, N12681, N12464);
buf BUF1 (N21224, N21221);
and AND4 (N21225, N21213, N4935, N17981, N13872);
buf BUF1 (N21226, N21223);
and AND2 (N21227, N21210, N20997);
not NOT1 (N21228, N21224);
xor XOR2 (N21229, N21217, N13152);
or OR4 (N21230, N21226, N14486, N6361, N19557);
nor NOR3 (N21231, N21206, N20057, N11689);
and AND4 (N21232, N21222, N7236, N191, N644);
and AND4 (N21233, N21216, N12884, N384, N5155);
or OR3 (N21234, N21229, N12291, N16621);
xor XOR2 (N21235, N21220, N20419);
or OR2 (N21236, N21235, N3281);
or OR2 (N21237, N21231, N3813);
not NOT1 (N21238, N21237);
not NOT1 (N21239, N21230);
xor XOR2 (N21240, N21236, N1080);
or OR3 (N21241, N21238, N6981, N3543);
or OR2 (N21242, N21241, N6636);
nor NOR3 (N21243, N21225, N10561, N10052);
and AND3 (N21244, N21239, N13407, N20586);
buf BUF1 (N21245, N21240);
xor XOR2 (N21246, N21242, N719);
nand NAND4 (N21247, N21244, N16965, N17036, N4433);
xor XOR2 (N21248, N21234, N31);
nand NAND2 (N21249, N21227, N11518);
or OR2 (N21250, N21245, N7962);
nand NAND3 (N21251, N21250, N14707, N4407);
xor XOR2 (N21252, N21243, N5294);
buf BUF1 (N21253, N21252);
and AND4 (N21254, N21228, N18792, N7049, N12828);
and AND4 (N21255, N21254, N2695, N7166, N5118);
not NOT1 (N21256, N21246);
and AND4 (N21257, N21247, N18331, N7320, N14185);
or OR2 (N21258, N21248, N11875);
xor XOR2 (N21259, N21257, N2767);
buf BUF1 (N21260, N21253);
nor NOR3 (N21261, N21218, N15858, N7965);
buf BUF1 (N21262, N21249);
xor XOR2 (N21263, N21256, N1648);
buf BUF1 (N21264, N21262);
buf BUF1 (N21265, N21251);
nor NOR4 (N21266, N21258, N15226, N6723, N14315);
nor NOR2 (N21267, N21255, N6581);
nor NOR3 (N21268, N21259, N7192, N13516);
not NOT1 (N21269, N21233);
buf BUF1 (N21270, N21261);
or OR4 (N21271, N21267, N18513, N8428, N15567);
xor XOR2 (N21272, N21260, N18742);
and AND4 (N21273, N21269, N16979, N3488, N240);
not NOT1 (N21274, N21270);
nor NOR3 (N21275, N21273, N1436, N11798);
nor NOR3 (N21276, N21264, N15143, N20288);
and AND3 (N21277, N21265, N18767, N3093);
not NOT1 (N21278, N21277);
not NOT1 (N21279, N21276);
not NOT1 (N21280, N21274);
buf BUF1 (N21281, N21280);
buf BUF1 (N21282, N21263);
and AND3 (N21283, N21279, N6325, N17061);
nand NAND2 (N21284, N21275, N15243);
and AND2 (N21285, N21281, N21001);
not NOT1 (N21286, N21232);
xor XOR2 (N21287, N21283, N10637);
buf BUF1 (N21288, N21271);
or OR3 (N21289, N21282, N8298, N16116);
xor XOR2 (N21290, N21284, N7629);
xor XOR2 (N21291, N21278, N2173);
not NOT1 (N21292, N21286);
and AND2 (N21293, N21291, N14101);
nor NOR2 (N21294, N21292, N5774);
not NOT1 (N21295, N21294);
buf BUF1 (N21296, N21295);
and AND2 (N21297, N21285, N18463);
nor NOR4 (N21298, N21287, N12049, N3552, N2463);
not NOT1 (N21299, N21293);
buf BUF1 (N21300, N21296);
or OR2 (N21301, N21268, N5667);
not NOT1 (N21302, N21298);
or OR3 (N21303, N21297, N18992, N15110);
buf BUF1 (N21304, N21272);
and AND2 (N21305, N21289, N18187);
nand NAND3 (N21306, N21305, N8546, N2665);
nor NOR3 (N21307, N21301, N6235, N16171);
nor NOR4 (N21308, N21290, N21061, N1914, N16539);
not NOT1 (N21309, N21302);
or OR3 (N21310, N21306, N11446, N2255);
nor NOR2 (N21311, N21303, N4190);
nor NOR3 (N21312, N21310, N10915, N9435);
not NOT1 (N21313, N21304);
or OR4 (N21314, N21288, N10779, N7463, N3022);
buf BUF1 (N21315, N21311);
not NOT1 (N21316, N21300);
nand NAND3 (N21317, N21307, N2728, N1394);
buf BUF1 (N21318, N21314);
xor XOR2 (N21319, N21266, N6830);
not NOT1 (N21320, N21316);
or OR4 (N21321, N21320, N1128, N3114, N17604);
buf BUF1 (N21322, N21319);
xor XOR2 (N21323, N21313, N8413);
and AND3 (N21324, N21299, N12993, N16);
buf BUF1 (N21325, N21318);
or OR2 (N21326, N21322, N13874);
and AND2 (N21327, N21323, N5358);
nor NOR4 (N21328, N21309, N18194, N8094, N9991);
buf BUF1 (N21329, N21321);
xor XOR2 (N21330, N21324, N1508);
not NOT1 (N21331, N21328);
buf BUF1 (N21332, N21326);
not NOT1 (N21333, N21330);
xor XOR2 (N21334, N21317, N9088);
not NOT1 (N21335, N21315);
or OR3 (N21336, N21312, N20940, N13848);
nor NOR3 (N21337, N21334, N5795, N2944);
and AND2 (N21338, N21333, N16114);
and AND2 (N21339, N21327, N4015);
or OR4 (N21340, N21329, N17408, N12707, N18146);
xor XOR2 (N21341, N21335, N12047);
not NOT1 (N21342, N21308);
nand NAND4 (N21343, N21325, N19096, N15348, N19349);
buf BUF1 (N21344, N21331);
not NOT1 (N21345, N21332);
or OR4 (N21346, N21344, N14358, N8061, N4087);
buf BUF1 (N21347, N21336);
and AND2 (N21348, N21340, N13261);
not NOT1 (N21349, N21345);
and AND2 (N21350, N21339, N20119);
nor NOR4 (N21351, N21350, N4475, N20447, N13825);
or OR4 (N21352, N21343, N7707, N4590, N2193);
xor XOR2 (N21353, N21341, N2878);
xor XOR2 (N21354, N21338, N9239);
and AND3 (N21355, N21346, N5495, N7348);
xor XOR2 (N21356, N21355, N8195);
nor NOR3 (N21357, N21348, N548, N3186);
and AND3 (N21358, N21357, N17293, N6830);
and AND3 (N21359, N21342, N8648, N7474);
nand NAND2 (N21360, N21337, N9938);
buf BUF1 (N21361, N21347);
xor XOR2 (N21362, N21353, N14653);
buf BUF1 (N21363, N21351);
not NOT1 (N21364, N21352);
xor XOR2 (N21365, N21354, N6606);
not NOT1 (N21366, N21358);
xor XOR2 (N21367, N21363, N10429);
nand NAND4 (N21368, N21361, N2047, N221, N18493);
not NOT1 (N21369, N21366);
not NOT1 (N21370, N21360);
or OR2 (N21371, N21356, N10414);
nand NAND3 (N21372, N21365, N215, N2137);
or OR2 (N21373, N21364, N496);
and AND2 (N21374, N21368, N13712);
nand NAND2 (N21375, N21367, N3421);
nand NAND2 (N21376, N21374, N4679);
nand NAND4 (N21377, N21372, N21245, N17936, N15781);
not NOT1 (N21378, N21362);
and AND2 (N21379, N21376, N13263);
nor NOR4 (N21380, N21371, N20007, N19064, N4006);
nor NOR3 (N21381, N21369, N14386, N8801);
not NOT1 (N21382, N21380);
nor NOR4 (N21383, N21378, N15718, N15166, N13997);
nand NAND3 (N21384, N21375, N19546, N7253);
buf BUF1 (N21385, N21382);
buf BUF1 (N21386, N21385);
not NOT1 (N21387, N21377);
nand NAND3 (N21388, N21386, N3483, N19899);
buf BUF1 (N21389, N21379);
nand NAND4 (N21390, N21384, N11212, N1420, N6559);
or OR2 (N21391, N21349, N12652);
and AND2 (N21392, N21383, N16977);
nand NAND4 (N21393, N21370, N7171, N20353, N4763);
nor NOR4 (N21394, N21389, N12412, N18612, N8682);
buf BUF1 (N21395, N21394);
nand NAND2 (N21396, N21373, N8566);
nor NOR2 (N21397, N21359, N18862);
not NOT1 (N21398, N21397);
or OR2 (N21399, N21395, N16485);
and AND4 (N21400, N21398, N17610, N10159, N16915);
not NOT1 (N21401, N21388);
or OR4 (N21402, N21396, N12574, N3140, N19729);
not NOT1 (N21403, N21393);
nand NAND3 (N21404, N21381, N1846, N10654);
nor NOR3 (N21405, N21391, N17387, N2413);
buf BUF1 (N21406, N21387);
and AND2 (N21407, N21400, N2192);
not NOT1 (N21408, N21403);
and AND3 (N21409, N21402, N7810, N9675);
nor NOR4 (N21410, N21408, N3746, N11446, N3442);
nor NOR3 (N21411, N21401, N7445, N4114);
not NOT1 (N21412, N21411);
not NOT1 (N21413, N21406);
or OR2 (N21414, N21412, N5553);
nor NOR3 (N21415, N21404, N13832, N17383);
or OR2 (N21416, N21405, N14703);
xor XOR2 (N21417, N21409, N19818);
or OR2 (N21418, N21416, N13179);
or OR4 (N21419, N21417, N11294, N2478, N17053);
buf BUF1 (N21420, N21407);
buf BUF1 (N21421, N21418);
not NOT1 (N21422, N21420);
buf BUF1 (N21423, N21414);
buf BUF1 (N21424, N21423);
nand NAND4 (N21425, N21415, N13285, N18696, N15669);
and AND4 (N21426, N21424, N18172, N590, N3738);
buf BUF1 (N21427, N21413);
buf BUF1 (N21428, N21390);
nand NAND2 (N21429, N21428, N10847);
and AND4 (N21430, N21410, N16684, N6573, N7022);
buf BUF1 (N21431, N21427);
nor NOR3 (N21432, N21392, N18784, N8229);
or OR4 (N21433, N21399, N19255, N11836, N12228);
not NOT1 (N21434, N21432);
xor XOR2 (N21435, N21419, N12257);
xor XOR2 (N21436, N21435, N18137);
nand NAND4 (N21437, N21430, N10807, N3625, N2862);
and AND2 (N21438, N21433, N14817);
xor XOR2 (N21439, N21429, N10676);
nor NOR3 (N21440, N21422, N1945, N20545);
or OR2 (N21441, N21421, N12273);
and AND2 (N21442, N21441, N8166);
or OR4 (N21443, N21438, N2067, N19886, N1353);
nand NAND2 (N21444, N21425, N11028);
or OR4 (N21445, N21442, N15298, N18561, N2249);
nor NOR2 (N21446, N21436, N10495);
and AND2 (N21447, N21426, N771);
nand NAND3 (N21448, N21440, N10671, N99);
and AND2 (N21449, N21434, N17420);
nand NAND3 (N21450, N21444, N10362, N12945);
nor NOR4 (N21451, N21445, N16385, N10706, N12145);
nor NOR2 (N21452, N21446, N1948);
xor XOR2 (N21453, N21448, N1223);
nand NAND4 (N21454, N21431, N14991, N19273, N12530);
nor NOR3 (N21455, N21447, N11860, N10106);
or OR3 (N21456, N21454, N15511, N15451);
or OR4 (N21457, N21450, N10125, N16057, N7795);
buf BUF1 (N21458, N21437);
or OR3 (N21459, N21449, N2725, N14695);
buf BUF1 (N21460, N21453);
xor XOR2 (N21461, N21456, N15109);
and AND2 (N21462, N21459, N2610);
nor NOR3 (N21463, N21460, N3967, N21237);
nand NAND3 (N21464, N21451, N12508, N19575);
or OR4 (N21465, N21439, N3172, N3242, N12968);
and AND4 (N21466, N21457, N21062, N12166, N1274);
xor XOR2 (N21467, N21464, N4225);
and AND2 (N21468, N21462, N6008);
nand NAND2 (N21469, N21463, N2370);
buf BUF1 (N21470, N21455);
xor XOR2 (N21471, N21465, N8711);
not NOT1 (N21472, N21458);
buf BUF1 (N21473, N21467);
buf BUF1 (N21474, N21470);
and AND2 (N21475, N21466, N8991);
not NOT1 (N21476, N21443);
xor XOR2 (N21477, N21472, N20718);
or OR3 (N21478, N21473, N16938, N8200);
nand NAND2 (N21479, N21468, N700);
or OR3 (N21480, N21474, N1985, N6763);
nand NAND4 (N21481, N21469, N5140, N7715, N17424);
and AND2 (N21482, N21480, N3855);
buf BUF1 (N21483, N21476);
nand NAND4 (N21484, N21479, N13304, N5342, N5894);
nor NOR2 (N21485, N21481, N18133);
or OR4 (N21486, N21485, N12023, N13250, N19361);
nand NAND4 (N21487, N21478, N2605, N13432, N3953);
nor NOR4 (N21488, N21482, N5913, N20972, N13056);
nand NAND3 (N21489, N21475, N289, N11641);
buf BUF1 (N21490, N21471);
buf BUF1 (N21491, N21489);
xor XOR2 (N21492, N21477, N17953);
nor NOR4 (N21493, N21492, N14268, N1779, N12432);
nand NAND4 (N21494, N21452, N6502, N20257, N4580);
nand NAND2 (N21495, N21486, N4456);
not NOT1 (N21496, N21491);
and AND4 (N21497, N21483, N8119, N10439, N18651);
xor XOR2 (N21498, N21494, N14937);
buf BUF1 (N21499, N21461);
not NOT1 (N21500, N21487);
nor NOR3 (N21501, N21496, N11513, N3919);
buf BUF1 (N21502, N21500);
or OR2 (N21503, N21495, N5383);
and AND3 (N21504, N21488, N7430, N11125);
and AND4 (N21505, N21499, N6568, N11606, N17730);
nor NOR2 (N21506, N21502, N20037);
and AND2 (N21507, N21505, N419);
nand NAND2 (N21508, N21490, N20106);
not NOT1 (N21509, N21504);
nand NAND3 (N21510, N21498, N4334, N3591);
or OR4 (N21511, N21507, N6515, N17011, N199);
nand NAND3 (N21512, N21501, N16358, N3240);
buf BUF1 (N21513, N21509);
nor NOR3 (N21514, N21503, N19629, N13547);
nand NAND3 (N21515, N21512, N14679, N5072);
or OR4 (N21516, N21508, N10807, N8534, N5219);
nand NAND3 (N21517, N21484, N11107, N198);
not NOT1 (N21518, N21510);
nand NAND3 (N21519, N21511, N9198, N7896);
nor NOR2 (N21520, N21519, N5984);
nor NOR2 (N21521, N21493, N8302);
not NOT1 (N21522, N21518);
buf BUF1 (N21523, N21515);
not NOT1 (N21524, N21497);
nand NAND2 (N21525, N21517, N378);
and AND3 (N21526, N21514, N19734, N4466);
xor XOR2 (N21527, N21523, N14805);
buf BUF1 (N21528, N21527);
not NOT1 (N21529, N21525);
buf BUF1 (N21530, N21526);
not NOT1 (N21531, N21513);
xor XOR2 (N21532, N21531, N7653);
nor NOR3 (N21533, N21516, N14160, N1151);
buf BUF1 (N21534, N21532);
nor NOR4 (N21535, N21521, N11851, N20976, N21360);
xor XOR2 (N21536, N21529, N635);
buf BUF1 (N21537, N21524);
buf BUF1 (N21538, N21530);
xor XOR2 (N21539, N21506, N6869);
or OR2 (N21540, N21538, N138);
nand NAND2 (N21541, N21534, N3183);
nand NAND3 (N21542, N21528, N20113, N1129);
and AND2 (N21543, N21539, N7195);
nor NOR3 (N21544, N21520, N7092, N13310);
and AND3 (N21545, N21540, N10254, N20589);
xor XOR2 (N21546, N21537, N7610);
and AND4 (N21547, N21536, N13476, N11074, N5356);
buf BUF1 (N21548, N21547);
xor XOR2 (N21549, N21543, N18780);
buf BUF1 (N21550, N21546);
not NOT1 (N21551, N21533);
nand NAND3 (N21552, N21522, N5611, N13694);
and AND2 (N21553, N21552, N5129);
nand NAND3 (N21554, N21544, N12006, N5517);
nor NOR4 (N21555, N21554, N13491, N20277, N8565);
nand NAND2 (N21556, N21555, N2969);
nand NAND4 (N21557, N21535, N18956, N2840, N17490);
not NOT1 (N21558, N21541);
xor XOR2 (N21559, N21542, N363);
or OR3 (N21560, N21551, N18310, N21288);
and AND3 (N21561, N21560, N12153, N12800);
not NOT1 (N21562, N21545);
buf BUF1 (N21563, N21561);
or OR2 (N21564, N21557, N13903);
nor NOR3 (N21565, N21553, N14423, N10974);
nor NOR3 (N21566, N21562, N17678, N13371);
nor NOR4 (N21567, N21566, N4812, N1508, N16178);
or OR4 (N21568, N21549, N16809, N4848, N335);
not NOT1 (N21569, N21567);
buf BUF1 (N21570, N21556);
not NOT1 (N21571, N21568);
not NOT1 (N21572, N21550);
xor XOR2 (N21573, N21570, N5889);
and AND3 (N21574, N21573, N16079, N14685);
or OR3 (N21575, N21571, N3941, N5288);
not NOT1 (N21576, N21564);
nand NAND2 (N21577, N21559, N10460);
and AND2 (N21578, N21558, N11444);
buf BUF1 (N21579, N21563);
xor XOR2 (N21580, N21548, N6496);
nor NOR3 (N21581, N21575, N5150, N7875);
or OR4 (N21582, N21565, N11025, N17433, N15057);
xor XOR2 (N21583, N21579, N5623);
xor XOR2 (N21584, N21576, N19568);
or OR2 (N21585, N21581, N16640);
buf BUF1 (N21586, N21574);
buf BUF1 (N21587, N21585);
xor XOR2 (N21588, N21586, N1522);
nor NOR2 (N21589, N21577, N2265);
nor NOR2 (N21590, N21584, N276);
buf BUF1 (N21591, N21589);
or OR2 (N21592, N21580, N2293);
not NOT1 (N21593, N21569);
buf BUF1 (N21594, N21593);
nor NOR2 (N21595, N21594, N15376);
buf BUF1 (N21596, N21572);
xor XOR2 (N21597, N21583, N7349);
buf BUF1 (N21598, N21588);
xor XOR2 (N21599, N21595, N19615);
or OR4 (N21600, N21592, N13895, N7024, N19438);
buf BUF1 (N21601, N21596);
or OR2 (N21602, N21599, N874);
nor NOR2 (N21603, N21591, N15726);
or OR4 (N21604, N21601, N1179, N10716, N17696);
and AND2 (N21605, N21602, N18980);
xor XOR2 (N21606, N21603, N15644);
and AND3 (N21607, N21598, N6673, N12262);
and AND2 (N21608, N21604, N19683);
buf BUF1 (N21609, N21597);
not NOT1 (N21610, N21600);
buf BUF1 (N21611, N21587);
nor NOR4 (N21612, N21609, N10477, N8006, N17465);
nor NOR4 (N21613, N21608, N748, N265, N376);
buf BUF1 (N21614, N21607);
nor NOR2 (N21615, N21610, N15267);
or OR2 (N21616, N21605, N20306);
buf BUF1 (N21617, N21616);
nor NOR4 (N21618, N21590, N8985, N17387, N7835);
nand NAND4 (N21619, N21615, N8110, N7573, N17384);
not NOT1 (N21620, N21614);
xor XOR2 (N21621, N21611, N6624);
nor NOR4 (N21622, N21612, N12626, N13929, N8568);
not NOT1 (N21623, N21578);
nor NOR2 (N21624, N21613, N481);
not NOT1 (N21625, N21623);
buf BUF1 (N21626, N21622);
nor NOR2 (N21627, N21626, N6696);
nor NOR2 (N21628, N21582, N7500);
buf BUF1 (N21629, N21624);
not NOT1 (N21630, N21621);
buf BUF1 (N21631, N21625);
or OR3 (N21632, N21629, N14748, N21119);
xor XOR2 (N21633, N21617, N6150);
xor XOR2 (N21634, N21628, N11766);
nor NOR4 (N21635, N21627, N7311, N20645, N16614);
nor NOR4 (N21636, N21633, N400, N15315, N16467);
or OR4 (N21637, N21619, N16519, N8149, N10490);
buf BUF1 (N21638, N21637);
xor XOR2 (N21639, N21634, N12053);
or OR3 (N21640, N21630, N13507, N17343);
nor NOR4 (N21641, N21640, N9526, N10108, N16755);
buf BUF1 (N21642, N21632);
nand NAND3 (N21643, N21635, N6310, N18150);
xor XOR2 (N21644, N21618, N2440);
not NOT1 (N21645, N21638);
and AND4 (N21646, N21645, N4385, N9240, N18158);
or OR4 (N21647, N21642, N4088, N15270, N9019);
nor NOR2 (N21648, N21606, N11344);
and AND3 (N21649, N21648, N2604, N15278);
nor NOR4 (N21650, N21631, N12103, N796, N7306);
buf BUF1 (N21651, N21636);
not NOT1 (N21652, N21643);
and AND2 (N21653, N21641, N4972);
or OR3 (N21654, N21646, N10212, N9650);
and AND3 (N21655, N21652, N2537, N7111);
nand NAND3 (N21656, N21639, N3271, N8791);
not NOT1 (N21657, N21656);
or OR4 (N21658, N21651, N1436, N18866, N16733);
or OR4 (N21659, N21655, N19833, N1049, N4130);
and AND3 (N21660, N21647, N3577, N5829);
nand NAND3 (N21661, N21653, N7837, N14101);
xor XOR2 (N21662, N21659, N11153);
buf BUF1 (N21663, N21657);
and AND2 (N21664, N21644, N4929);
buf BUF1 (N21665, N21649);
or OR2 (N21666, N21620, N13075);
buf BUF1 (N21667, N21661);
buf BUF1 (N21668, N21662);
not NOT1 (N21669, N21654);
xor XOR2 (N21670, N21668, N16390);
xor XOR2 (N21671, N21665, N18315);
or OR3 (N21672, N21663, N6847, N2959);
nand NAND4 (N21673, N21672, N20003, N14653, N11131);
not NOT1 (N21674, N21671);
and AND3 (N21675, N21673, N20975, N19118);
or OR4 (N21676, N21667, N16235, N6008, N5210);
nand NAND2 (N21677, N21674, N5154);
not NOT1 (N21678, N21676);
nor NOR2 (N21679, N21660, N8324);
or OR4 (N21680, N21658, N1267, N11411, N10750);
xor XOR2 (N21681, N21666, N9533);
xor XOR2 (N21682, N21664, N15832);
or OR3 (N21683, N21678, N7036, N5781);
buf BUF1 (N21684, N21679);
or OR2 (N21685, N21650, N457);
buf BUF1 (N21686, N21684);
nand NAND3 (N21687, N21683, N7465, N9043);
nand NAND4 (N21688, N21670, N9262, N5821, N4937);
or OR4 (N21689, N21681, N8691, N4903, N6676);
nor NOR4 (N21690, N21677, N5606, N9242, N7479);
and AND2 (N21691, N21689, N11518);
or OR2 (N21692, N21691, N12845);
or OR3 (N21693, N21675, N16037, N11258);
or OR2 (N21694, N21690, N15471);
or OR3 (N21695, N21686, N20976, N13889);
buf BUF1 (N21696, N21688);
nand NAND4 (N21697, N21682, N14920, N10648, N538);
or OR4 (N21698, N21685, N17295, N4738, N21002);
xor XOR2 (N21699, N21695, N3592);
xor XOR2 (N21700, N21698, N13993);
and AND4 (N21701, N21693, N11072, N9286, N17500);
and AND4 (N21702, N21687, N11481, N18172, N878);
xor XOR2 (N21703, N21699, N2114);
buf BUF1 (N21704, N21692);
not NOT1 (N21705, N21702);
xor XOR2 (N21706, N21696, N5620);
buf BUF1 (N21707, N21694);
xor XOR2 (N21708, N21700, N2788);
not NOT1 (N21709, N21697);
nand NAND4 (N21710, N21703, N5507, N16741, N21261);
and AND3 (N21711, N21709, N5029, N8304);
and AND4 (N21712, N21701, N395, N21291, N11727);
or OR3 (N21713, N21705, N2697, N12634);
nand NAND3 (N21714, N21712, N10778, N10635);
nor NOR4 (N21715, N21680, N5387, N2352, N2548);
nor NOR3 (N21716, N21708, N9578, N15203);
nand NAND4 (N21717, N21711, N20674, N5264, N4122);
not NOT1 (N21718, N21714);
xor XOR2 (N21719, N21717, N20604);
nor NOR4 (N21720, N21713, N21130, N15336, N10247);
not NOT1 (N21721, N21710);
nor NOR4 (N21722, N21707, N12414, N3398, N16944);
buf BUF1 (N21723, N21721);
nand NAND2 (N21724, N21715, N18864);
nor NOR3 (N21725, N21706, N9761, N5871);
not NOT1 (N21726, N21720);
nor NOR3 (N21727, N21725, N16308, N17622);
not NOT1 (N21728, N21718);
xor XOR2 (N21729, N21722, N3768);
nand NAND2 (N21730, N21716, N3102);
not NOT1 (N21731, N21728);
buf BUF1 (N21732, N21723);
buf BUF1 (N21733, N21729);
buf BUF1 (N21734, N21732);
not NOT1 (N21735, N21730);
or OR3 (N21736, N21726, N1850, N17369);
nor NOR2 (N21737, N21736, N16983);
nand NAND2 (N21738, N21669, N10819);
buf BUF1 (N21739, N21737);
not NOT1 (N21740, N21724);
and AND4 (N21741, N21733, N1796, N5992, N9827);
nor NOR4 (N21742, N21738, N5511, N10265, N4147);
buf BUF1 (N21743, N21719);
nor NOR3 (N21744, N21704, N13251, N11863);
nor NOR4 (N21745, N21741, N2289, N8366, N8670);
nand NAND2 (N21746, N21731, N2633);
nand NAND3 (N21747, N21746, N18450, N15975);
buf BUF1 (N21748, N21742);
buf BUF1 (N21749, N21743);
nand NAND3 (N21750, N21734, N21003, N2471);
and AND2 (N21751, N21740, N20769);
xor XOR2 (N21752, N21744, N5400);
nand NAND4 (N21753, N21748, N215, N10816, N3537);
or OR4 (N21754, N21753, N9967, N15787, N165);
or OR4 (N21755, N21749, N17364, N21624, N6487);
not NOT1 (N21756, N21752);
not NOT1 (N21757, N21727);
not NOT1 (N21758, N21755);
and AND2 (N21759, N21751, N2583);
nand NAND3 (N21760, N21754, N9427, N10187);
not NOT1 (N21761, N21735);
nor NOR3 (N21762, N21759, N7044, N8545);
nor NOR4 (N21763, N21745, N12806, N14820, N18076);
not NOT1 (N21764, N21756);
and AND2 (N21765, N21750, N1759);
xor XOR2 (N21766, N21764, N19062);
nand NAND3 (N21767, N21757, N18395, N1867);
xor XOR2 (N21768, N21761, N17274);
nor NOR3 (N21769, N21739, N18524, N12554);
buf BUF1 (N21770, N21760);
not NOT1 (N21771, N21766);
nor NOR2 (N21772, N21767, N12704);
nor NOR3 (N21773, N21768, N2500, N6697);
nor NOR2 (N21774, N21762, N10201);
nor NOR2 (N21775, N21774, N17946);
and AND4 (N21776, N21775, N3463, N1996, N2165);
not NOT1 (N21777, N21769);
nor NOR3 (N21778, N21771, N5933, N2801);
nor NOR4 (N21779, N21758, N8205, N3039, N7893);
xor XOR2 (N21780, N21773, N4999);
not NOT1 (N21781, N21763);
not NOT1 (N21782, N21780);
nor NOR3 (N21783, N21776, N4650, N3298);
xor XOR2 (N21784, N21765, N16344);
or OR4 (N21785, N21778, N1745, N5538, N17339);
xor XOR2 (N21786, N21781, N20229);
nor NOR2 (N21787, N21785, N7650);
or OR2 (N21788, N21779, N3785);
or OR2 (N21789, N21784, N12974);
buf BUF1 (N21790, N21770);
buf BUF1 (N21791, N21787);
not NOT1 (N21792, N21788);
nand NAND3 (N21793, N21747, N19034, N7364);
xor XOR2 (N21794, N21786, N6679);
not NOT1 (N21795, N21789);
nor NOR4 (N21796, N21790, N20482, N7914, N18278);
xor XOR2 (N21797, N21772, N149);
nor NOR2 (N21798, N21794, N5514);
xor XOR2 (N21799, N21798, N1311);
nand NAND3 (N21800, N21797, N5212, N3482);
or OR2 (N21801, N21796, N1141);
nand NAND3 (N21802, N21793, N12873, N19873);
or OR2 (N21803, N21802, N2710);
buf BUF1 (N21804, N21800);
nor NOR3 (N21805, N21803, N71, N14806);
not NOT1 (N21806, N21804);
and AND2 (N21807, N21777, N15293);
not NOT1 (N21808, N21795);
nand NAND3 (N21809, N21808, N3637, N1479);
nand NAND3 (N21810, N21792, N15466, N14292);
not NOT1 (N21811, N21807);
xor XOR2 (N21812, N21806, N10344);
and AND4 (N21813, N21799, N11686, N10237, N1113);
xor XOR2 (N21814, N21805, N4303);
buf BUF1 (N21815, N21791);
buf BUF1 (N21816, N21801);
or OR2 (N21817, N21815, N3965);
and AND2 (N21818, N21783, N18200);
xor XOR2 (N21819, N21812, N1818);
not NOT1 (N21820, N21809);
or OR2 (N21821, N21816, N343);
or OR3 (N21822, N21819, N8497, N10853);
and AND3 (N21823, N21813, N11632, N20219);
nor NOR4 (N21824, N21823, N19847, N1080, N9355);
buf BUF1 (N21825, N21782);
nand NAND4 (N21826, N21821, N17068, N20540, N1383);
nor NOR3 (N21827, N21817, N16250, N12791);
or OR2 (N21828, N21827, N3648);
and AND4 (N21829, N21811, N6644, N19043, N13263);
nand NAND3 (N21830, N21820, N2703, N15727);
and AND2 (N21831, N21824, N1491);
nand NAND3 (N21832, N21826, N12719, N15141);
nor NOR3 (N21833, N21814, N8320, N1739);
nand NAND2 (N21834, N21810, N7043);
xor XOR2 (N21835, N21831, N20641);
or OR4 (N21836, N21832, N3173, N3036, N11215);
or OR3 (N21837, N21834, N13070, N9852);
buf BUF1 (N21838, N21828);
not NOT1 (N21839, N21830);
and AND3 (N21840, N21836, N1767, N17929);
buf BUF1 (N21841, N21833);
xor XOR2 (N21842, N21835, N18658);
xor XOR2 (N21843, N21829, N5612);
not NOT1 (N21844, N21839);
nor NOR3 (N21845, N21841, N20839, N11279);
not NOT1 (N21846, N21822);
buf BUF1 (N21847, N21842);
buf BUF1 (N21848, N21837);
nand NAND3 (N21849, N21844, N9123, N6617);
or OR2 (N21850, N21838, N17316);
nand NAND4 (N21851, N21825, N16687, N8159, N9485);
nand NAND4 (N21852, N21847, N17839, N1622, N9402);
or OR3 (N21853, N21845, N16824, N15556);
xor XOR2 (N21854, N21853, N18409);
xor XOR2 (N21855, N21849, N5376);
and AND2 (N21856, N21852, N8561);
nor NOR3 (N21857, N21840, N4891, N8175);
nand NAND2 (N21858, N21850, N11378);
or OR3 (N21859, N21858, N15581, N4069);
buf BUF1 (N21860, N21818);
not NOT1 (N21861, N21846);
nor NOR3 (N21862, N21854, N5373, N6242);
xor XOR2 (N21863, N21843, N4522);
not NOT1 (N21864, N21855);
not NOT1 (N21865, N21860);
xor XOR2 (N21866, N21864, N1265);
xor XOR2 (N21867, N21851, N20356);
xor XOR2 (N21868, N21863, N16911);
nand NAND2 (N21869, N21859, N2579);
nor NOR3 (N21870, N21866, N2915, N8780);
and AND4 (N21871, N21848, N535, N4383, N12301);
buf BUF1 (N21872, N21867);
xor XOR2 (N21873, N21861, N17168);
xor XOR2 (N21874, N21868, N9686);
xor XOR2 (N21875, N21862, N4704);
xor XOR2 (N21876, N21869, N5364);
or OR4 (N21877, N21865, N21352, N11880, N14959);
not NOT1 (N21878, N21872);
nor NOR3 (N21879, N21857, N793, N19823);
nor NOR2 (N21880, N21871, N12675);
and AND2 (N21881, N21878, N2466);
nor NOR2 (N21882, N21880, N2908);
nor NOR3 (N21883, N21882, N20319, N17582);
xor XOR2 (N21884, N21870, N6287);
not NOT1 (N21885, N21884);
and AND2 (N21886, N21883, N19090);
and AND3 (N21887, N21876, N13025, N3810);
or OR3 (N21888, N21873, N13183, N9077);
nor NOR2 (N21889, N21881, N6049);
xor XOR2 (N21890, N21886, N4961);
nor NOR4 (N21891, N21877, N1664, N2436, N7106);
xor XOR2 (N21892, N21891, N12009);
nor NOR2 (N21893, N21885, N1583);
nor NOR2 (N21894, N21887, N15839);
and AND2 (N21895, N21892, N1083);
nand NAND4 (N21896, N21879, N973, N21893, N12124);
nor NOR2 (N21897, N4364, N5785);
not NOT1 (N21898, N21896);
and AND2 (N21899, N21890, N11726);
or OR3 (N21900, N21856, N7303, N3837);
not NOT1 (N21901, N21875);
nor NOR4 (N21902, N21894, N2984, N8054, N15438);
xor XOR2 (N21903, N21889, N9535);
xor XOR2 (N21904, N21895, N4131);
nand NAND2 (N21905, N21900, N16364);
xor XOR2 (N21906, N21901, N11247);
or OR4 (N21907, N21904, N2486, N16085, N10969);
nor NOR4 (N21908, N21907, N21006, N12784, N11290);
not NOT1 (N21909, N21906);
nand NAND3 (N21910, N21888, N5620, N13037);
nor NOR3 (N21911, N21897, N21355, N19770);
not NOT1 (N21912, N21909);
buf BUF1 (N21913, N21902);
xor XOR2 (N21914, N21898, N5173);
buf BUF1 (N21915, N21899);
not NOT1 (N21916, N21912);
and AND4 (N21917, N21874, N11033, N6396, N4471);
nor NOR4 (N21918, N21905, N7364, N2173, N19014);
buf BUF1 (N21919, N21913);
and AND2 (N21920, N21918, N19749);
nor NOR3 (N21921, N21916, N9101, N20043);
buf BUF1 (N21922, N21903);
nor NOR2 (N21923, N21922, N18663);
and AND4 (N21924, N21908, N7254, N7633, N2396);
not NOT1 (N21925, N21917);
buf BUF1 (N21926, N21920);
or OR2 (N21927, N21923, N17305);
nand NAND2 (N21928, N21915, N1075);
nor NOR3 (N21929, N21921, N12727, N2352);
and AND3 (N21930, N21910, N5981, N5559);
nand NAND2 (N21931, N21926, N8132);
or OR2 (N21932, N21930, N1908);
or OR4 (N21933, N21932, N17695, N12914, N7566);
buf BUF1 (N21934, N21925);
or OR4 (N21935, N21927, N15461, N20051, N12540);
nor NOR3 (N21936, N21935, N17911, N10710);
nor NOR3 (N21937, N21914, N3461, N775);
buf BUF1 (N21938, N21911);
xor XOR2 (N21939, N21919, N10446);
not NOT1 (N21940, N21924);
nor NOR3 (N21941, N21936, N8665, N2316);
not NOT1 (N21942, N21933);
nand NAND2 (N21943, N21938, N1080);
nor NOR4 (N21944, N21942, N3260, N5128, N3379);
nor NOR2 (N21945, N21939, N3313);
or OR2 (N21946, N21940, N6440);
and AND3 (N21947, N21944, N7996, N3335);
buf BUF1 (N21948, N21931);
and AND2 (N21949, N21941, N6784);
nand NAND3 (N21950, N21943, N7325, N18437);
nand NAND2 (N21951, N21929, N5710);
and AND2 (N21952, N21937, N11835);
not NOT1 (N21953, N21947);
xor XOR2 (N21954, N21951, N13349);
xor XOR2 (N21955, N21948, N3670);
and AND3 (N21956, N21952, N4478, N3687);
xor XOR2 (N21957, N21956, N825);
and AND4 (N21958, N21955, N21884, N4382, N17067);
nand NAND4 (N21959, N21928, N20335, N5538, N987);
buf BUF1 (N21960, N21949);
xor XOR2 (N21961, N21953, N979);
nand NAND3 (N21962, N21958, N16228, N5925);
nor NOR3 (N21963, N21954, N15245, N21211);
or OR3 (N21964, N21950, N13090, N20328);
nor NOR4 (N21965, N21960, N10658, N13295, N3501);
buf BUF1 (N21966, N21963);
not NOT1 (N21967, N21959);
xor XOR2 (N21968, N21962, N13873);
or OR2 (N21969, N21964, N20833);
xor XOR2 (N21970, N21961, N21879);
xor XOR2 (N21971, N21934, N2861);
xor XOR2 (N21972, N21970, N21244);
not NOT1 (N21973, N21969);
nand NAND3 (N21974, N21946, N5830, N21166);
nand NAND2 (N21975, N21957, N74);
nor NOR4 (N21976, N21974, N9356, N15337, N13152);
xor XOR2 (N21977, N21973, N16566);
or OR4 (N21978, N21966, N13413, N6821, N18876);
or OR2 (N21979, N21977, N13484);
or OR3 (N21980, N21967, N11302, N4553);
xor XOR2 (N21981, N21976, N16854);
nand NAND3 (N21982, N21978, N1140, N886);
and AND3 (N21983, N21979, N17046, N926);
or OR2 (N21984, N21983, N8091);
nor NOR2 (N21985, N21945, N16204);
nand NAND2 (N21986, N21975, N1757);
not NOT1 (N21987, N21972);
and AND3 (N21988, N21968, N20958, N8252);
or OR3 (N21989, N21965, N15412, N18755);
xor XOR2 (N21990, N21987, N13253);
nor NOR3 (N21991, N21984, N3931, N1820);
and AND4 (N21992, N21985, N15037, N14415, N4509);
nand NAND3 (N21993, N21992, N5243, N16433);
and AND2 (N21994, N21988, N8792);
and AND2 (N21995, N21981, N12802);
xor XOR2 (N21996, N21994, N6159);
not NOT1 (N21997, N21990);
nand NAND2 (N21998, N21989, N7410);
nor NOR4 (N21999, N21997, N17796, N2032, N9472);
not NOT1 (N22000, N21991);
nor NOR3 (N22001, N21999, N1512, N4395);
or OR2 (N22002, N21998, N21917);
and AND2 (N22003, N21996, N3567);
and AND3 (N22004, N22001, N7765, N7030);
and AND3 (N22005, N21971, N15907, N11314);
buf BUF1 (N22006, N21986);
nand NAND2 (N22007, N22000, N18591);
xor XOR2 (N22008, N22005, N8452);
xor XOR2 (N22009, N22006, N18332);
xor XOR2 (N22010, N22007, N21487);
xor XOR2 (N22011, N22009, N20173);
xor XOR2 (N22012, N22008, N16070);
buf BUF1 (N22013, N22010);
xor XOR2 (N22014, N22013, N5748);
and AND4 (N22015, N22003, N15568, N697, N1086);
or OR3 (N22016, N21982, N19978, N16169);
nand NAND3 (N22017, N21993, N966, N17306);
nor NOR2 (N22018, N22012, N21405);
nor NOR3 (N22019, N22018, N262, N16926);
or OR4 (N22020, N22014, N18804, N17257, N18372);
xor XOR2 (N22021, N22019, N5013);
nand NAND3 (N22022, N22002, N9993, N14143);
xor XOR2 (N22023, N22017, N14612);
nand NAND3 (N22024, N22023, N16930, N18041);
nand NAND3 (N22025, N21980, N19339, N3184);
buf BUF1 (N22026, N22022);
nand NAND3 (N22027, N22015, N14423, N15146);
xor XOR2 (N22028, N22004, N1686);
nor NOR4 (N22029, N22016, N19412, N5733, N13817);
xor XOR2 (N22030, N22021, N6259);
and AND3 (N22031, N22030, N675, N13616);
nand NAND4 (N22032, N22027, N195, N13311, N4113);
nor NOR4 (N22033, N22028, N21442, N1907, N1549);
or OR2 (N22034, N22033, N10179);
buf BUF1 (N22035, N22020);
or OR3 (N22036, N22025, N4425, N18444);
nor NOR4 (N22037, N22029, N17403, N20356, N3662);
not NOT1 (N22038, N22032);
not NOT1 (N22039, N22024);
nand NAND4 (N22040, N22035, N13987, N10079, N16454);
nand NAND2 (N22041, N22034, N15602);
nand NAND2 (N22042, N22031, N11617);
not NOT1 (N22043, N22038);
xor XOR2 (N22044, N22039, N21893);
buf BUF1 (N22045, N22026);
or OR3 (N22046, N21995, N4815, N4737);
or OR2 (N22047, N22041, N3140);
or OR4 (N22048, N22037, N2306, N21158, N21210);
nand NAND2 (N22049, N22047, N19669);
xor XOR2 (N22050, N22036, N16658);
not NOT1 (N22051, N22043);
or OR3 (N22052, N22044, N16253, N7772);
nor NOR3 (N22053, N22045, N150, N9399);
and AND4 (N22054, N22051, N967, N19129, N6);
xor XOR2 (N22055, N22054, N18933);
buf BUF1 (N22056, N22050);
buf BUF1 (N22057, N22056);
or OR4 (N22058, N22053, N17570, N20320, N11733);
and AND4 (N22059, N22046, N17614, N7426, N16372);
xor XOR2 (N22060, N22048, N13399);
or OR3 (N22061, N22058, N21449, N11999);
xor XOR2 (N22062, N22040, N10959);
buf BUF1 (N22063, N22052);
not NOT1 (N22064, N22062);
nand NAND4 (N22065, N22064, N8988, N13555, N5450);
nor NOR3 (N22066, N22061, N21220, N993);
or OR3 (N22067, N22057, N13193, N8575);
buf BUF1 (N22068, N22049);
and AND2 (N22069, N22060, N6294);
nand NAND3 (N22070, N22065, N14367, N227);
and AND3 (N22071, N22070, N14021, N14475);
buf BUF1 (N22072, N22066);
not NOT1 (N22073, N22011);
xor XOR2 (N22074, N22042, N4818);
buf BUF1 (N22075, N22072);
nor NOR3 (N22076, N22063, N4477, N21913);
xor XOR2 (N22077, N22073, N10210);
or OR3 (N22078, N22059, N9757, N6997);
nand NAND4 (N22079, N22055, N8559, N1894, N16601);
xor XOR2 (N22080, N22069, N3626);
or OR4 (N22081, N22074, N19804, N19760, N10270);
xor XOR2 (N22082, N22075, N3401);
and AND4 (N22083, N22076, N6478, N15806, N13928);
and AND4 (N22084, N22077, N15072, N15610, N8524);
xor XOR2 (N22085, N22071, N6628);
xor XOR2 (N22086, N22083, N3531);
or OR3 (N22087, N22085, N4993, N19767);
and AND4 (N22088, N22067, N10948, N17621, N17286);
nor NOR4 (N22089, N22081, N19991, N383, N19596);
and AND4 (N22090, N22086, N9277, N8728, N9979);
buf BUF1 (N22091, N22087);
or OR4 (N22092, N22088, N3868, N6942, N3535);
nand NAND2 (N22093, N22090, N8726);
nor NOR4 (N22094, N22092, N18523, N3720, N21209);
nor NOR4 (N22095, N22080, N7060, N14425, N8852);
xor XOR2 (N22096, N22078, N10448);
not NOT1 (N22097, N22096);
and AND4 (N22098, N22082, N5789, N1001, N4796);
not NOT1 (N22099, N22095);
and AND4 (N22100, N22068, N19194, N15306, N18888);
and AND4 (N22101, N22093, N18335, N17762, N14902);
nor NOR3 (N22102, N22094, N14570, N7331);
and AND3 (N22103, N22084, N11566, N19340);
or OR4 (N22104, N22098, N6144, N19143, N3876);
xor XOR2 (N22105, N22100, N1500);
and AND4 (N22106, N22091, N2151, N4693, N4007);
or OR4 (N22107, N22106, N6101, N21630, N8357);
or OR3 (N22108, N22101, N12345, N8731);
not NOT1 (N22109, N22104);
not NOT1 (N22110, N22105);
and AND4 (N22111, N22109, N4241, N3206, N9218);
nor NOR2 (N22112, N22107, N7556);
xor XOR2 (N22113, N22103, N6534);
or OR2 (N22114, N22097, N16138);
nand NAND4 (N22115, N22110, N13094, N21642, N20436);
nand NAND3 (N22116, N22115, N20859, N11255);
nand NAND4 (N22117, N22099, N15191, N5819, N5391);
and AND2 (N22118, N22112, N8487);
not NOT1 (N22119, N22108);
and AND4 (N22120, N22102, N7359, N16175, N18152);
and AND4 (N22121, N22119, N11078, N2199, N1313);
xor XOR2 (N22122, N22117, N10131);
or OR3 (N22123, N22116, N12207, N2776);
xor XOR2 (N22124, N22121, N5342);
nor NOR3 (N22125, N22079, N20224, N10628);
or OR3 (N22126, N22118, N19115, N6316);
not NOT1 (N22127, N22122);
xor XOR2 (N22128, N22123, N2827);
not NOT1 (N22129, N22120);
nand NAND4 (N22130, N22126, N6034, N3422, N19773);
or OR4 (N22131, N22129, N1157, N9856, N13321);
nor NOR4 (N22132, N22125, N3845, N11327, N4888);
and AND3 (N22133, N22127, N16870, N12960);
not NOT1 (N22134, N22111);
nor NOR2 (N22135, N22114, N6740);
nand NAND4 (N22136, N22130, N3702, N16179, N14938);
xor XOR2 (N22137, N22132, N2976);
and AND4 (N22138, N22134, N11503, N8249, N14436);
xor XOR2 (N22139, N22135, N9747);
not NOT1 (N22140, N22139);
nand NAND4 (N22141, N22140, N9271, N5795, N1);
xor XOR2 (N22142, N22089, N735);
nor NOR2 (N22143, N22113, N17990);
buf BUF1 (N22144, N22142);
not NOT1 (N22145, N22141);
xor XOR2 (N22146, N22124, N4075);
xor XOR2 (N22147, N22143, N12681);
nand NAND3 (N22148, N22137, N12682, N8899);
and AND2 (N22149, N22144, N4094);
not NOT1 (N22150, N22128);
and AND4 (N22151, N22146, N17984, N4476, N15535);
and AND3 (N22152, N22131, N17007, N14909);
nor NOR2 (N22153, N22151, N4457);
nor NOR3 (N22154, N22153, N5284, N13449);
nand NAND4 (N22155, N22152, N8839, N10924, N4964);
nor NOR4 (N22156, N22133, N4918, N14870, N12100);
xor XOR2 (N22157, N22154, N13243);
xor XOR2 (N22158, N22148, N4426);
nand NAND3 (N22159, N22150, N6316, N9452);
or OR4 (N22160, N22157, N10451, N8584, N21747);
xor XOR2 (N22161, N22147, N7258);
nor NOR4 (N22162, N22161, N16722, N19208, N9371);
nor NOR4 (N22163, N22149, N10062, N20354, N9844);
nor NOR3 (N22164, N22158, N9161, N19174);
and AND3 (N22165, N22155, N15154, N10036);
nor NOR2 (N22166, N22163, N16428);
xor XOR2 (N22167, N22138, N343);
nand NAND4 (N22168, N22162, N14950, N16029, N14958);
xor XOR2 (N22169, N22165, N14144);
buf BUF1 (N22170, N22167);
nand NAND2 (N22171, N22156, N9007);
not NOT1 (N22172, N22159);
nor NOR3 (N22173, N22136, N17851, N1672);
nor NOR2 (N22174, N22169, N4642);
and AND3 (N22175, N22173, N6684, N11438);
buf BUF1 (N22176, N22145);
or OR3 (N22177, N22170, N17214, N5498);
nor NOR2 (N22178, N22171, N12401);
nor NOR2 (N22179, N22174, N16414);
nor NOR4 (N22180, N22168, N7022, N4684, N7037);
buf BUF1 (N22181, N22175);
or OR2 (N22182, N22178, N20798);
not NOT1 (N22183, N22172);
xor XOR2 (N22184, N22179, N5742);
nor NOR4 (N22185, N22164, N6627, N11567, N13337);
and AND3 (N22186, N22181, N4762, N8041);
and AND4 (N22187, N22182, N3232, N10321, N17485);
nor NOR3 (N22188, N22186, N16731, N9194);
xor XOR2 (N22189, N22176, N9019);
not NOT1 (N22190, N22184);
not NOT1 (N22191, N22185);
and AND3 (N22192, N22187, N17835, N10539);
and AND4 (N22193, N22180, N19956, N14128, N15270);
and AND4 (N22194, N22193, N20859, N11607, N17265);
not NOT1 (N22195, N22183);
or OR2 (N22196, N22195, N1620);
buf BUF1 (N22197, N22189);
nand NAND4 (N22198, N22177, N6911, N1973, N20189);
buf BUF1 (N22199, N22196);
nor NOR2 (N22200, N22194, N3808);
nand NAND3 (N22201, N22198, N3, N11976);
xor XOR2 (N22202, N22201, N3063);
xor XOR2 (N22203, N22160, N1154);
xor XOR2 (N22204, N22191, N21584);
not NOT1 (N22205, N22203);
or OR3 (N22206, N22205, N14481, N18646);
xor XOR2 (N22207, N22166, N9360);
xor XOR2 (N22208, N22188, N4143);
buf BUF1 (N22209, N22204);
nand NAND4 (N22210, N22207, N31, N2081, N1714);
and AND3 (N22211, N22190, N19038, N15559);
nand NAND3 (N22212, N22206, N2056, N20712);
not NOT1 (N22213, N22200);
buf BUF1 (N22214, N22197);
nand NAND2 (N22215, N22212, N7569);
nor NOR3 (N22216, N22199, N11187, N20384);
buf BUF1 (N22217, N22202);
buf BUF1 (N22218, N22209);
and AND3 (N22219, N22211, N2900, N19678);
xor XOR2 (N22220, N22219, N21010);
not NOT1 (N22221, N22217);
buf BUF1 (N22222, N22218);
not NOT1 (N22223, N22221);
nor NOR3 (N22224, N22216, N8529, N13586);
nor NOR3 (N22225, N22210, N1383, N4984);
or OR2 (N22226, N22192, N17399);
xor XOR2 (N22227, N22213, N21626);
and AND2 (N22228, N22220, N4209);
not NOT1 (N22229, N22226);
nor NOR3 (N22230, N22227, N14179, N9216);
not NOT1 (N22231, N22214);
not NOT1 (N22232, N22229);
buf BUF1 (N22233, N22215);
xor XOR2 (N22234, N22233, N17728);
and AND3 (N22235, N22230, N6577, N7104);
buf BUF1 (N22236, N22223);
nor NOR2 (N22237, N22225, N4221);
or OR2 (N22238, N22237, N13005);
not NOT1 (N22239, N22232);
xor XOR2 (N22240, N22238, N4028);
and AND2 (N22241, N22236, N5538);
or OR2 (N22242, N22222, N15738);
nor NOR2 (N22243, N22239, N21917);
nor NOR2 (N22244, N22231, N397);
xor XOR2 (N22245, N22228, N20242);
and AND4 (N22246, N22245, N22113, N20240, N18765);
not NOT1 (N22247, N22234);
not NOT1 (N22248, N22247);
nand NAND4 (N22249, N22235, N941, N17505, N426);
buf BUF1 (N22250, N22242);
not NOT1 (N22251, N22244);
buf BUF1 (N22252, N22241);
nor NOR3 (N22253, N22248, N18996, N15949);
xor XOR2 (N22254, N22251, N8941);
nand NAND2 (N22255, N22252, N44);
buf BUF1 (N22256, N22254);
and AND4 (N22257, N22208, N8342, N4411, N14335);
xor XOR2 (N22258, N22257, N6006);
nor NOR4 (N22259, N22258, N11665, N3646, N3558);
and AND3 (N22260, N22259, N21533, N18089);
xor XOR2 (N22261, N22224, N10800);
buf BUF1 (N22262, N22243);
and AND2 (N22263, N22249, N21307);
or OR2 (N22264, N22256, N11535);
xor XOR2 (N22265, N22263, N21668);
xor XOR2 (N22266, N22250, N17074);
nand NAND4 (N22267, N22246, N12177, N15732, N2295);
and AND4 (N22268, N22266, N11215, N5335, N4190);
xor XOR2 (N22269, N22260, N14773);
or OR3 (N22270, N22261, N17039, N8371);
and AND2 (N22271, N22269, N6362);
buf BUF1 (N22272, N22240);
xor XOR2 (N22273, N22255, N19838);
xor XOR2 (N22274, N22262, N12076);
nand NAND4 (N22275, N22270, N10898, N19128, N1733);
and AND4 (N22276, N22275, N12695, N2307, N524);
not NOT1 (N22277, N22267);
xor XOR2 (N22278, N22271, N13467);
or OR3 (N22279, N22277, N18324, N18152);
xor XOR2 (N22280, N22268, N7462);
not NOT1 (N22281, N22253);
not NOT1 (N22282, N22273);
buf BUF1 (N22283, N22276);
nor NOR4 (N22284, N22280, N7087, N21726, N19464);
nand NAND4 (N22285, N22283, N13905, N11626, N16694);
not NOT1 (N22286, N22282);
nor NOR4 (N22287, N22285, N8181, N20169, N17385);
xor XOR2 (N22288, N22287, N20511);
nand NAND4 (N22289, N22278, N13302, N20066, N8743);
and AND4 (N22290, N22264, N1238, N2886, N8332);
and AND2 (N22291, N22281, N21348);
and AND3 (N22292, N22288, N7542, N1719);
or OR4 (N22293, N22292, N7276, N12266, N7060);
or OR4 (N22294, N22286, N7869, N8780, N15114);
nand NAND4 (N22295, N22293, N4032, N17888, N10731);
or OR2 (N22296, N22289, N4495);
buf BUF1 (N22297, N22279);
nand NAND4 (N22298, N22294, N14196, N3630, N14637);
nor NOR2 (N22299, N22295, N7517);
nand NAND3 (N22300, N22291, N2087, N10054);
not NOT1 (N22301, N22274);
xor XOR2 (N22302, N22298, N5317);
nor NOR3 (N22303, N22290, N21876, N14319);
buf BUF1 (N22304, N22265);
and AND2 (N22305, N22302, N6405);
and AND3 (N22306, N22299, N20346, N1525);
xor XOR2 (N22307, N22303, N19137);
and AND4 (N22308, N22307, N10481, N19262, N19867);
nor NOR3 (N22309, N22284, N10078, N5034);
or OR2 (N22310, N22272, N18006);
buf BUF1 (N22311, N22306);
or OR2 (N22312, N22310, N15973);
buf BUF1 (N22313, N22308);
nand NAND2 (N22314, N22301, N20276);
xor XOR2 (N22315, N22296, N17219);
or OR2 (N22316, N22304, N21871);
buf BUF1 (N22317, N22316);
and AND4 (N22318, N22317, N14121, N21132, N11117);
xor XOR2 (N22319, N22297, N11595);
or OR3 (N22320, N22318, N5590, N309);
xor XOR2 (N22321, N22315, N13576);
not NOT1 (N22322, N22319);
and AND2 (N22323, N22305, N9577);
and AND3 (N22324, N22300, N14412, N3352);
xor XOR2 (N22325, N22313, N19126);
nor NOR2 (N22326, N22323, N11538);
not NOT1 (N22327, N22320);
nand NAND3 (N22328, N22314, N13958, N2597);
nor NOR3 (N22329, N22326, N4924, N22185);
and AND3 (N22330, N22322, N11, N497);
nor NOR2 (N22331, N22309, N17399);
nand NAND3 (N22332, N22329, N7479, N20387);
xor XOR2 (N22333, N22331, N15275);
not NOT1 (N22334, N22311);
not NOT1 (N22335, N22332);
not NOT1 (N22336, N22325);
nor NOR3 (N22337, N22324, N7121, N4288);
and AND3 (N22338, N22312, N2760, N20635);
nand NAND3 (N22339, N22321, N5501, N9029);
nand NAND4 (N22340, N22328, N21507, N197, N17305);
nor NOR2 (N22341, N22334, N16609);
nand NAND2 (N22342, N22327, N14516);
or OR3 (N22343, N22340, N20844, N15414);
or OR2 (N22344, N22330, N15556);
not NOT1 (N22345, N22342);
or OR3 (N22346, N22341, N177, N9285);
nor NOR2 (N22347, N22336, N7066);
xor XOR2 (N22348, N22346, N4726);
nor NOR3 (N22349, N22347, N15758, N19546);
nor NOR3 (N22350, N22333, N2622, N11631);
or OR2 (N22351, N22345, N9412);
not NOT1 (N22352, N22350);
not NOT1 (N22353, N22337);
nor NOR2 (N22354, N22351, N8673);
or OR2 (N22355, N22339, N18421);
and AND2 (N22356, N22355, N8220);
nor NOR4 (N22357, N22344, N16722, N7280, N1060);
xor XOR2 (N22358, N22356, N14822);
not NOT1 (N22359, N22335);
and AND4 (N22360, N22354, N793, N17833, N13714);
nor NOR2 (N22361, N22358, N3388);
and AND3 (N22362, N22360, N8849, N2804);
and AND3 (N22363, N22357, N10241, N22280);
and AND2 (N22364, N22361, N730);
xor XOR2 (N22365, N22348, N6721);
nand NAND3 (N22366, N22363, N8633, N21997);
nor NOR4 (N22367, N22338, N1965, N20176, N14900);
nor NOR2 (N22368, N22364, N3136);
nor NOR3 (N22369, N22352, N7012, N8655);
buf BUF1 (N22370, N22368);
not NOT1 (N22371, N22366);
and AND3 (N22372, N22371, N21177, N571);
xor XOR2 (N22373, N22343, N14214);
and AND4 (N22374, N22349, N16766, N14936, N21118);
buf BUF1 (N22375, N22359);
or OR4 (N22376, N22375, N17228, N12940, N7161);
nand NAND4 (N22377, N22365, N10694, N20907, N2764);
and AND2 (N22378, N22369, N11336);
nand NAND4 (N22379, N22372, N18430, N15708, N21650);
buf BUF1 (N22380, N22373);
not NOT1 (N22381, N22374);
nor NOR4 (N22382, N22362, N8218, N1177, N2336);
not NOT1 (N22383, N22378);
buf BUF1 (N22384, N22377);
buf BUF1 (N22385, N22367);
or OR3 (N22386, N22379, N12465, N19871);
not NOT1 (N22387, N22384);
and AND3 (N22388, N22386, N4114, N16787);
and AND4 (N22389, N22385, N12344, N1529, N18600);
nor NOR3 (N22390, N22382, N15403, N1810);
xor XOR2 (N22391, N22370, N11018);
xor XOR2 (N22392, N22376, N708);
not NOT1 (N22393, N22387);
nor NOR3 (N22394, N22390, N12326, N7686);
buf BUF1 (N22395, N22388);
nand NAND4 (N22396, N22394, N818, N18692, N11996);
or OR3 (N22397, N22389, N6693, N11944);
or OR4 (N22398, N22380, N5159, N4587, N17698);
nand NAND3 (N22399, N22396, N6783, N14867);
and AND4 (N22400, N22395, N8475, N21472, N14800);
not NOT1 (N22401, N22399);
xor XOR2 (N22402, N22397, N5276);
xor XOR2 (N22403, N22401, N7700);
xor XOR2 (N22404, N22402, N21892);
nor NOR3 (N22405, N22404, N17790, N17723);
nand NAND3 (N22406, N22398, N16036, N4805);
nor NOR3 (N22407, N22381, N7596, N16532);
and AND3 (N22408, N22391, N17087, N20076);
xor XOR2 (N22409, N22407, N10424);
not NOT1 (N22410, N22383);
xor XOR2 (N22411, N22410, N8598);
nand NAND2 (N22412, N22405, N8568);
buf BUF1 (N22413, N22406);
xor XOR2 (N22414, N22393, N6431);
or OR4 (N22415, N22392, N3254, N7104, N12184);
and AND4 (N22416, N22408, N368, N5015, N8453);
nand NAND4 (N22417, N22415, N12297, N14232, N2573);
nor NOR4 (N22418, N22403, N14688, N6792, N19045);
xor XOR2 (N22419, N22409, N17143);
xor XOR2 (N22420, N22414, N13413);
or OR3 (N22421, N22416, N14478, N5537);
or OR4 (N22422, N22411, N21634, N60, N11531);
or OR4 (N22423, N22400, N11330, N5885, N8724);
xor XOR2 (N22424, N22423, N21678);
nor NOR2 (N22425, N22418, N13665);
or OR4 (N22426, N22422, N15835, N5688, N13700);
nor NOR2 (N22427, N22413, N20543);
xor XOR2 (N22428, N22425, N3444);
or OR2 (N22429, N22412, N166);
not NOT1 (N22430, N22426);
xor XOR2 (N22431, N22428, N6892);
and AND3 (N22432, N22421, N6694, N20786);
or OR4 (N22433, N22420, N6322, N15938, N589);
not NOT1 (N22434, N22432);
not NOT1 (N22435, N22434);
nand NAND4 (N22436, N22419, N4475, N9780, N14819);
nor NOR2 (N22437, N22429, N17682);
nand NAND4 (N22438, N22427, N14682, N9091, N6235);
not NOT1 (N22439, N22417);
buf BUF1 (N22440, N22439);
and AND4 (N22441, N22424, N2226, N12675, N8501);
nand NAND4 (N22442, N22436, N7465, N19465, N17191);
not NOT1 (N22443, N22438);
xor XOR2 (N22444, N22435, N243);
or OR3 (N22445, N22440, N14442, N13303);
xor XOR2 (N22446, N22437, N18559);
nand NAND3 (N22447, N22442, N8401, N7299);
buf BUF1 (N22448, N22353);
nor NOR4 (N22449, N22447, N12818, N14241, N17611);
nand NAND3 (N22450, N22430, N17961, N17085);
nand NAND4 (N22451, N22444, N14192, N15127, N1815);
and AND2 (N22452, N22448, N16625);
not NOT1 (N22453, N22441);
or OR3 (N22454, N22451, N8825, N18535);
and AND2 (N22455, N22449, N3157);
not NOT1 (N22456, N22453);
xor XOR2 (N22457, N22431, N6104);
xor XOR2 (N22458, N22446, N10295);
nor NOR3 (N22459, N22450, N17107, N15501);
buf BUF1 (N22460, N22456);
or OR2 (N22461, N22443, N10999);
and AND3 (N22462, N22433, N12562, N9200);
buf BUF1 (N22463, N22445);
not NOT1 (N22464, N22460);
not NOT1 (N22465, N22462);
not NOT1 (N22466, N22465);
or OR4 (N22467, N22464, N18934, N11311, N6238);
and AND2 (N22468, N22463, N3112);
buf BUF1 (N22469, N22467);
nor NOR2 (N22470, N22466, N18910);
not NOT1 (N22471, N22458);
and AND2 (N22472, N22468, N11368);
and AND4 (N22473, N22472, N5984, N12954, N16243);
xor XOR2 (N22474, N22473, N16416);
and AND4 (N22475, N22457, N19305, N18980, N20086);
not NOT1 (N22476, N22469);
xor XOR2 (N22477, N22455, N11957);
nand NAND2 (N22478, N22475, N15866);
buf BUF1 (N22479, N22454);
buf BUF1 (N22480, N22479);
xor XOR2 (N22481, N22461, N22448);
xor XOR2 (N22482, N22478, N19162);
nor NOR4 (N22483, N22452, N20222, N7124, N5820);
buf BUF1 (N22484, N22483);
nor NOR2 (N22485, N22480, N8028);
or OR2 (N22486, N22477, N2887);
nand NAND4 (N22487, N22482, N13698, N2770, N17861);
and AND2 (N22488, N22485, N11552);
nor NOR4 (N22489, N22488, N10003, N11525, N7375);
and AND2 (N22490, N22487, N15977);
or OR4 (N22491, N22474, N17237, N18240, N10619);
and AND2 (N22492, N22490, N4064);
and AND2 (N22493, N22484, N22382);
nand NAND2 (N22494, N22489, N20228);
buf BUF1 (N22495, N22491);
and AND4 (N22496, N22494, N3531, N16150, N480);
or OR4 (N22497, N22496, N1768, N13638, N7378);
or OR3 (N22498, N22493, N15120, N9390);
nor NOR4 (N22499, N22495, N17961, N13427, N18657);
or OR4 (N22500, N22499, N9251, N9547, N14032);
not NOT1 (N22501, N22486);
nand NAND2 (N22502, N22492, N11492);
not NOT1 (N22503, N22502);
xor XOR2 (N22504, N22498, N15478);
nand NAND4 (N22505, N22501, N9167, N6464, N16756);
nor NOR2 (N22506, N22471, N6550);
or OR4 (N22507, N22497, N22292, N8601, N4350);
nand NAND3 (N22508, N22459, N17006, N14183);
buf BUF1 (N22509, N22500);
or OR4 (N22510, N22470, N11939, N17427, N13650);
nand NAND4 (N22511, N22476, N16250, N3747, N2646);
buf BUF1 (N22512, N22481);
not NOT1 (N22513, N22510);
nor NOR2 (N22514, N22504, N2868);
not NOT1 (N22515, N22508);
nor NOR3 (N22516, N22507, N21104, N4512);
or OR2 (N22517, N22515, N22113);
xor XOR2 (N22518, N22505, N12186);
not NOT1 (N22519, N22512);
not NOT1 (N22520, N22509);
not NOT1 (N22521, N22506);
and AND2 (N22522, N22514, N1007);
nor NOR3 (N22523, N22522, N8338, N3344);
or OR4 (N22524, N22511, N15329, N21745, N365);
nand NAND3 (N22525, N22519, N22498, N19519);
not NOT1 (N22526, N22525);
xor XOR2 (N22527, N22518, N17879);
and AND3 (N22528, N22526, N6921, N8421);
buf BUF1 (N22529, N22520);
nand NAND2 (N22530, N22529, N1192);
or OR3 (N22531, N22516, N1936, N21222);
nor NOR3 (N22532, N22531, N16920, N2258);
nand NAND3 (N22533, N22532, N15754, N9331);
nor NOR4 (N22534, N22533, N19207, N13037, N22020);
and AND2 (N22535, N22513, N2129);
and AND4 (N22536, N22524, N16490, N7437, N14956);
nor NOR2 (N22537, N22536, N8474);
or OR2 (N22538, N22535, N22263);
and AND3 (N22539, N22538, N2073, N19048);
nor NOR3 (N22540, N22534, N15969, N5625);
nand NAND2 (N22541, N22530, N21973);
or OR3 (N22542, N22503, N20799, N11599);
xor XOR2 (N22543, N22521, N10732);
or OR2 (N22544, N22537, N22021);
buf BUF1 (N22545, N22528);
buf BUF1 (N22546, N22539);
buf BUF1 (N22547, N22541);
and AND4 (N22548, N22542, N7865, N6602, N17418);
xor XOR2 (N22549, N22527, N20498);
or OR2 (N22550, N22544, N14425);
nand NAND4 (N22551, N22546, N11859, N11522, N17715);
buf BUF1 (N22552, N22523);
buf BUF1 (N22553, N22548);
not NOT1 (N22554, N22543);
buf BUF1 (N22555, N22547);
buf BUF1 (N22556, N22555);
nor NOR2 (N22557, N22551, N9920);
and AND4 (N22558, N22553, N17190, N2798, N13430);
nand NAND3 (N22559, N22554, N3145, N12330);
and AND3 (N22560, N22559, N14376, N1235);
xor XOR2 (N22561, N22549, N7656);
xor XOR2 (N22562, N22558, N13102);
xor XOR2 (N22563, N22556, N5012);
not NOT1 (N22564, N22561);
buf BUF1 (N22565, N22517);
nor NOR2 (N22566, N22564, N20032);
nand NAND2 (N22567, N22552, N6014);
nor NOR4 (N22568, N22565, N20942, N22518, N15002);
buf BUF1 (N22569, N22563);
and AND3 (N22570, N22557, N2504, N19098);
buf BUF1 (N22571, N22570);
and AND2 (N22572, N22567, N4816);
not NOT1 (N22573, N22568);
buf BUF1 (N22574, N22571);
buf BUF1 (N22575, N22545);
and AND3 (N22576, N22550, N15540, N8211);
xor XOR2 (N22577, N22576, N11854);
or OR3 (N22578, N22560, N4551, N305);
and AND2 (N22579, N22578, N10930);
or OR3 (N22580, N22575, N19761, N5694);
xor XOR2 (N22581, N22540, N18474);
nand NAND3 (N22582, N22574, N569, N5210);
nor NOR4 (N22583, N22579, N1756, N6289, N8901);
and AND3 (N22584, N22569, N20237, N15740);
and AND3 (N22585, N22581, N9345, N9149);
nor NOR4 (N22586, N22572, N12452, N2833, N608);
and AND4 (N22587, N22585, N7286, N8927, N72);
and AND4 (N22588, N22586, N9810, N16842, N7716);
xor XOR2 (N22589, N22566, N11153);
or OR3 (N22590, N22584, N18130, N5619);
not NOT1 (N22591, N22589);
nor NOR3 (N22592, N22590, N16871, N839);
and AND4 (N22593, N22587, N2443, N3664, N15451);
not NOT1 (N22594, N22593);
not NOT1 (N22595, N22562);
nor NOR3 (N22596, N22592, N19177, N12373);
and AND4 (N22597, N22588, N11294, N10735, N3330);
nor NOR3 (N22598, N22594, N20417, N18237);
or OR4 (N22599, N22597, N8991, N14532, N15340);
buf BUF1 (N22600, N22573);
not NOT1 (N22601, N22591);
buf BUF1 (N22602, N22600);
not NOT1 (N22603, N22601);
xor XOR2 (N22604, N22602, N22236);
nor NOR2 (N22605, N22580, N193);
xor XOR2 (N22606, N22599, N3137);
nor NOR2 (N22607, N22604, N12314);
nand NAND2 (N22608, N22582, N11046);
not NOT1 (N22609, N22598);
nand NAND2 (N22610, N22583, N12028);
nor NOR4 (N22611, N22610, N8954, N4849, N8915);
buf BUF1 (N22612, N22603);
xor XOR2 (N22613, N22608, N10043);
or OR3 (N22614, N22577, N5759, N13192);
nand NAND4 (N22615, N22611, N20077, N15249, N21934);
and AND2 (N22616, N22613, N3113);
not NOT1 (N22617, N22616);
xor XOR2 (N22618, N22596, N13286);
or OR2 (N22619, N22607, N16777);
nor NOR3 (N22620, N22614, N4859, N19065);
buf BUF1 (N22621, N22605);
and AND4 (N22622, N22620, N22535, N18901, N6412);
not NOT1 (N22623, N22612);
and AND2 (N22624, N22618, N13850);
nor NOR4 (N22625, N22606, N10363, N15491, N7747);
nand NAND3 (N22626, N22624, N10474, N14394);
nor NOR4 (N22627, N22617, N10481, N18387, N17298);
and AND2 (N22628, N22595, N15565);
or OR2 (N22629, N22625, N22158);
xor XOR2 (N22630, N22619, N5919);
xor XOR2 (N22631, N22623, N15777);
buf BUF1 (N22632, N22621);
nor NOR2 (N22633, N22615, N4369);
xor XOR2 (N22634, N22632, N3841);
nand NAND3 (N22635, N22622, N14056, N9169);
nor NOR2 (N22636, N22626, N22584);
buf BUF1 (N22637, N22634);
xor XOR2 (N22638, N22631, N21333);
nand NAND3 (N22639, N22627, N16953, N14716);
nor NOR2 (N22640, N22630, N1585);
and AND2 (N22641, N22628, N13877);
nand NAND2 (N22642, N22629, N13249);
and AND4 (N22643, N22640, N6372, N8870, N2619);
not NOT1 (N22644, N22609);
or OR2 (N22645, N22636, N18705);
not NOT1 (N22646, N22633);
buf BUF1 (N22647, N22635);
nor NOR2 (N22648, N22639, N20885);
and AND3 (N22649, N22642, N19510, N21659);
nand NAND4 (N22650, N22641, N17534, N14454, N17204);
nor NOR3 (N22651, N22650, N18175, N1245);
buf BUF1 (N22652, N22645);
and AND2 (N22653, N22646, N9368);
not NOT1 (N22654, N22653);
xor XOR2 (N22655, N22652, N14848);
buf BUF1 (N22656, N22651);
buf BUF1 (N22657, N22655);
buf BUF1 (N22658, N22649);
nand NAND4 (N22659, N22647, N15259, N1896, N13849);
or OR3 (N22660, N22658, N14887, N1752);
and AND2 (N22661, N22637, N15198);
not NOT1 (N22662, N22648);
nor NOR4 (N22663, N22661, N13505, N15293, N11859);
and AND4 (N22664, N22638, N14031, N5086, N568);
and AND2 (N22665, N22643, N18014);
and AND2 (N22666, N22659, N18990);
xor XOR2 (N22667, N22665, N1928);
or OR2 (N22668, N22663, N4128);
nand NAND4 (N22669, N22662, N14571, N16627, N7561);
nand NAND4 (N22670, N22656, N16050, N9013, N1731);
nor NOR3 (N22671, N22670, N18287, N7491);
nor NOR2 (N22672, N22666, N21620);
buf BUF1 (N22673, N22660);
and AND3 (N22674, N22673, N1214, N12180);
buf BUF1 (N22675, N22674);
xor XOR2 (N22676, N22672, N21517);
nor NOR4 (N22677, N22664, N6905, N4271, N16418);
nand NAND2 (N22678, N22654, N19458);
and AND2 (N22679, N22668, N11734);
nor NOR4 (N22680, N22678, N950, N13729, N4607);
nand NAND2 (N22681, N22680, N2247);
xor XOR2 (N22682, N22667, N19342);
not NOT1 (N22683, N22682);
nand NAND4 (N22684, N22657, N17313, N15691, N8507);
xor XOR2 (N22685, N22677, N20614);
not NOT1 (N22686, N22684);
buf BUF1 (N22687, N22686);
nand NAND4 (N22688, N22669, N1373, N11794, N16412);
buf BUF1 (N22689, N22679);
nand NAND4 (N22690, N22683, N9577, N15109, N2833);
not NOT1 (N22691, N22671);
and AND4 (N22692, N22688, N20889, N2041, N2400);
or OR4 (N22693, N22675, N13289, N1323, N6271);
nor NOR4 (N22694, N22692, N6912, N6281, N7312);
buf BUF1 (N22695, N22687);
not NOT1 (N22696, N22695);
not NOT1 (N22697, N22644);
nand NAND4 (N22698, N22697, N8683, N4672, N15588);
nor NOR4 (N22699, N22696, N8704, N17638, N18630);
nand NAND3 (N22700, N22681, N13389, N18361);
or OR4 (N22701, N22676, N10503, N14726, N15740);
buf BUF1 (N22702, N22701);
buf BUF1 (N22703, N22690);
xor XOR2 (N22704, N22685, N8553);
or OR4 (N22705, N22689, N20193, N6567, N8413);
or OR4 (N22706, N22700, N5263, N16632, N7428);
buf BUF1 (N22707, N22691);
nand NAND3 (N22708, N22703, N6836, N17302);
nor NOR4 (N22709, N22704, N3820, N17886, N6400);
not NOT1 (N22710, N22694);
not NOT1 (N22711, N22693);
buf BUF1 (N22712, N22706);
not NOT1 (N22713, N22708);
xor XOR2 (N22714, N22711, N9853);
nor NOR3 (N22715, N22699, N12353, N4453);
xor XOR2 (N22716, N22714, N14008);
nor NOR2 (N22717, N22715, N21403);
and AND4 (N22718, N22702, N3433, N13185, N4975);
nor NOR2 (N22719, N22707, N20745);
or OR2 (N22720, N22718, N15953);
not NOT1 (N22721, N22719);
xor XOR2 (N22722, N22709, N10221);
buf BUF1 (N22723, N22716);
nor NOR3 (N22724, N22720, N12543, N11852);
nor NOR2 (N22725, N22723, N5493);
xor XOR2 (N22726, N22721, N21432);
and AND3 (N22727, N22726, N18846, N14494);
or OR2 (N22728, N22698, N5389);
nand NAND4 (N22729, N22717, N7797, N22479, N2083);
buf BUF1 (N22730, N22710);
xor XOR2 (N22731, N22713, N16753);
nand NAND3 (N22732, N22731, N2305, N22723);
not NOT1 (N22733, N22712);
and AND4 (N22734, N22727, N1116, N20828, N12344);
and AND3 (N22735, N22732, N17904, N6118);
or OR2 (N22736, N22725, N4463);
or OR2 (N22737, N22729, N14552);
nor NOR3 (N22738, N22733, N637, N5497);
nand NAND4 (N22739, N22734, N8217, N2761, N13421);
buf BUF1 (N22740, N22705);
or OR4 (N22741, N22722, N1650, N3437, N17147);
nor NOR2 (N22742, N22728, N5631);
xor XOR2 (N22743, N22742, N20130);
nor NOR2 (N22744, N22737, N16705);
and AND3 (N22745, N22744, N13954, N2010);
buf BUF1 (N22746, N22735);
buf BUF1 (N22747, N22730);
xor XOR2 (N22748, N22746, N21280);
nand NAND4 (N22749, N22738, N17533, N18540, N16299);
nand NAND2 (N22750, N22739, N7214);
nor NOR4 (N22751, N22743, N15409, N11509, N1050);
buf BUF1 (N22752, N22745);
or OR4 (N22753, N22724, N10766, N7169, N10326);
or OR2 (N22754, N22740, N1970);
or OR4 (N22755, N22752, N18046, N10925, N9230);
not NOT1 (N22756, N22747);
xor XOR2 (N22757, N22755, N10360);
nor NOR3 (N22758, N22741, N18186, N16370);
buf BUF1 (N22759, N22751);
xor XOR2 (N22760, N22749, N20554);
and AND3 (N22761, N22753, N12624, N5985);
xor XOR2 (N22762, N22756, N15639);
nand NAND4 (N22763, N22760, N7489, N203, N17928);
nand NAND2 (N22764, N22757, N1557);
nand NAND4 (N22765, N22764, N11716, N16981, N10926);
nand NAND3 (N22766, N22750, N17587, N13110);
xor XOR2 (N22767, N22762, N2207);
and AND4 (N22768, N22748, N5822, N16118, N14542);
xor XOR2 (N22769, N22767, N21403);
xor XOR2 (N22770, N22768, N18426);
buf BUF1 (N22771, N22758);
nor NOR4 (N22772, N22765, N3050, N10305, N3176);
nand NAND3 (N22773, N22770, N20262, N12902);
nor NOR4 (N22774, N22773, N7486, N1606, N14252);
xor XOR2 (N22775, N22772, N17100);
xor XOR2 (N22776, N22774, N10997);
nand NAND2 (N22777, N22766, N16108);
or OR4 (N22778, N22759, N4371, N5522, N2649);
not NOT1 (N22779, N22763);
xor XOR2 (N22780, N22775, N666);
and AND4 (N22781, N22778, N7981, N15849, N7557);
or OR2 (N22782, N22754, N357);
xor XOR2 (N22783, N22779, N7413);
nor NOR4 (N22784, N22777, N14185, N9257, N7766);
xor XOR2 (N22785, N22784, N21850);
buf BUF1 (N22786, N22782);
and AND4 (N22787, N22771, N1678, N14220, N15574);
or OR3 (N22788, N22787, N7393, N22401);
and AND2 (N22789, N22761, N9023);
xor XOR2 (N22790, N22783, N7003);
or OR2 (N22791, N22790, N16667);
and AND3 (N22792, N22788, N8580, N21586);
not NOT1 (N22793, N22769);
or OR2 (N22794, N22780, N14704);
not NOT1 (N22795, N22786);
and AND4 (N22796, N22776, N8998, N12674, N13538);
and AND3 (N22797, N22794, N12193, N9852);
buf BUF1 (N22798, N22736);
xor XOR2 (N22799, N22793, N9750);
not NOT1 (N22800, N22785);
nor NOR4 (N22801, N22781, N7295, N22762, N17986);
not NOT1 (N22802, N22801);
nor NOR3 (N22803, N22795, N18207, N5808);
nor NOR4 (N22804, N22798, N11871, N15474, N5306);
xor XOR2 (N22805, N22799, N6324);
nand NAND3 (N22806, N22805, N5062, N2114);
nor NOR3 (N22807, N22791, N15049, N19391);
xor XOR2 (N22808, N22806, N17174);
or OR2 (N22809, N22797, N2767);
not NOT1 (N22810, N22807);
buf BUF1 (N22811, N22789);
buf BUF1 (N22812, N22792);
xor XOR2 (N22813, N22810, N9581);
and AND4 (N22814, N22804, N10903, N5636, N8130);
nand NAND4 (N22815, N22802, N11238, N1486, N5105);
nor NOR3 (N22816, N22796, N16732, N7237);
xor XOR2 (N22817, N22813, N19450);
xor XOR2 (N22818, N22815, N18079);
or OR2 (N22819, N22809, N5876);
xor XOR2 (N22820, N22818, N4630);
nor NOR3 (N22821, N22800, N19246, N259);
and AND4 (N22822, N22816, N335, N17865, N18780);
and AND3 (N22823, N22819, N19371, N1467);
xor XOR2 (N22824, N22811, N5638);
buf BUF1 (N22825, N22824);
not NOT1 (N22826, N22803);
not NOT1 (N22827, N22821);
nand NAND4 (N22828, N22826, N6962, N1895, N18071);
or OR2 (N22829, N22822, N9019);
and AND3 (N22830, N22829, N18372, N10272);
not NOT1 (N22831, N22827);
xor XOR2 (N22832, N22830, N10582);
nand NAND3 (N22833, N22823, N5185, N9634);
xor XOR2 (N22834, N22812, N10700);
nand NAND2 (N22835, N22831, N22820);
not NOT1 (N22836, N21464);
nand NAND3 (N22837, N22836, N4226, N7046);
nor NOR2 (N22838, N22833, N17401);
buf BUF1 (N22839, N22835);
or OR4 (N22840, N22828, N18966, N13501, N4370);
buf BUF1 (N22841, N22834);
xor XOR2 (N22842, N22808, N10476);
and AND4 (N22843, N22839, N2306, N5432, N7371);
xor XOR2 (N22844, N22825, N5344);
not NOT1 (N22845, N22843);
nor NOR3 (N22846, N22840, N20289, N20517);
xor XOR2 (N22847, N22838, N13464);
nand NAND3 (N22848, N22837, N920, N10700);
not NOT1 (N22849, N22814);
nand NAND2 (N22850, N22841, N9418);
nor NOR4 (N22851, N22817, N13370, N2853, N13305);
or OR2 (N22852, N22851, N8629);
nor NOR2 (N22853, N22842, N22603);
nand NAND4 (N22854, N22846, N10865, N5320, N20729);
and AND2 (N22855, N22854, N10170);
or OR4 (N22856, N22850, N10113, N5013, N12198);
nand NAND2 (N22857, N22832, N13751);
not NOT1 (N22858, N22852);
nand NAND2 (N22859, N22856, N3621);
or OR4 (N22860, N22858, N16462, N9215, N21094);
or OR2 (N22861, N22855, N5629);
and AND4 (N22862, N22857, N12090, N12149, N11168);
nor NOR3 (N22863, N22849, N19310, N17267);
nand NAND4 (N22864, N22847, N4832, N9119, N19562);
xor XOR2 (N22865, N22860, N19026);
not NOT1 (N22866, N22864);
nand NAND4 (N22867, N22845, N9062, N13758, N10119);
and AND4 (N22868, N22867, N13718, N22721, N22740);
nand NAND2 (N22869, N22853, N14443);
or OR3 (N22870, N22862, N6272, N3169);
not NOT1 (N22871, N22868);
and AND3 (N22872, N22848, N2031, N7304);
and AND3 (N22873, N22872, N5126, N17517);
or OR4 (N22874, N22861, N13209, N9179, N8650);
not NOT1 (N22875, N22863);
buf BUF1 (N22876, N22866);
or OR4 (N22877, N22865, N8650, N8610, N17563);
not NOT1 (N22878, N22875);
nand NAND3 (N22879, N22869, N14159, N12243);
not NOT1 (N22880, N22877);
nand NAND3 (N22881, N22870, N8125, N19859);
buf BUF1 (N22882, N22874);
xor XOR2 (N22883, N22879, N18234);
buf BUF1 (N22884, N22844);
xor XOR2 (N22885, N22873, N9282);
not NOT1 (N22886, N22883);
not NOT1 (N22887, N22884);
buf BUF1 (N22888, N22882);
nand NAND2 (N22889, N22886, N618);
xor XOR2 (N22890, N22887, N12799);
nand NAND3 (N22891, N22880, N4751, N19380);
not NOT1 (N22892, N22885);
buf BUF1 (N22893, N22881);
xor XOR2 (N22894, N22878, N18751);
nand NAND2 (N22895, N22888, N21789);
xor XOR2 (N22896, N22859, N3424);
not NOT1 (N22897, N22891);
and AND2 (N22898, N22876, N6409);
xor XOR2 (N22899, N22890, N15754);
xor XOR2 (N22900, N22897, N17870);
and AND2 (N22901, N22889, N9038);
not NOT1 (N22902, N22899);
or OR3 (N22903, N22900, N10070, N3287);
not NOT1 (N22904, N22902);
xor XOR2 (N22905, N22895, N22528);
or OR3 (N22906, N22901, N13214, N18825);
nor NOR3 (N22907, N22903, N9123, N3069);
and AND3 (N22908, N22893, N1191, N19746);
xor XOR2 (N22909, N22896, N18647);
and AND3 (N22910, N22907, N18762, N4082);
xor XOR2 (N22911, N22871, N6143);
nand NAND2 (N22912, N22904, N6740);
xor XOR2 (N22913, N22909, N20653);
not NOT1 (N22914, N22898);
nor NOR3 (N22915, N22913, N11913, N5930);
not NOT1 (N22916, N22905);
or OR3 (N22917, N22910, N21368, N8344);
and AND2 (N22918, N22911, N3734);
and AND2 (N22919, N22894, N21301);
and AND2 (N22920, N22906, N3495);
buf BUF1 (N22921, N22918);
xor XOR2 (N22922, N22920, N11444);
xor XOR2 (N22923, N22922, N10239);
and AND2 (N22924, N22917, N9776);
xor XOR2 (N22925, N22923, N8148);
not NOT1 (N22926, N22915);
not NOT1 (N22927, N22925);
not NOT1 (N22928, N22919);
buf BUF1 (N22929, N22926);
xor XOR2 (N22930, N22916, N11439);
xor XOR2 (N22931, N22892, N7832);
buf BUF1 (N22932, N22928);
not NOT1 (N22933, N22932);
or OR2 (N22934, N22930, N18220);
xor XOR2 (N22935, N22934, N20555);
nand NAND3 (N22936, N22924, N9234, N14926);
not NOT1 (N22937, N22908);
not NOT1 (N22938, N22935);
nor NOR4 (N22939, N22936, N19113, N17453, N9205);
nor NOR4 (N22940, N22914, N12597, N773, N549);
nor NOR4 (N22941, N22940, N11448, N5386, N22323);
nor NOR4 (N22942, N22927, N21638, N8680, N7186);
nor NOR2 (N22943, N22912, N21604);
and AND2 (N22944, N22942, N13294);
xor XOR2 (N22945, N22933, N8682);
or OR3 (N22946, N22945, N9934, N2148);
xor XOR2 (N22947, N22944, N8992);
not NOT1 (N22948, N22938);
buf BUF1 (N22949, N22929);
and AND3 (N22950, N22941, N7205, N21426);
buf BUF1 (N22951, N22931);
nor NOR3 (N22952, N22946, N17086, N9557);
and AND3 (N22953, N22921, N10062, N15329);
not NOT1 (N22954, N22953);
and AND3 (N22955, N22950, N17883, N22107);
buf BUF1 (N22956, N22955);
nor NOR3 (N22957, N22952, N4604, N2092);
nand NAND3 (N22958, N22939, N10893, N22301);
and AND4 (N22959, N22943, N4872, N4122, N11277);
xor XOR2 (N22960, N22958, N12221);
not NOT1 (N22961, N22959);
buf BUF1 (N22962, N22949);
nor NOR3 (N22963, N22951, N16008, N7837);
buf BUF1 (N22964, N22963);
and AND4 (N22965, N22956, N22821, N4208, N5268);
buf BUF1 (N22966, N22962);
nand NAND4 (N22967, N22947, N8470, N14837, N22405);
not NOT1 (N22968, N22954);
or OR3 (N22969, N22948, N22121, N11006);
nor NOR2 (N22970, N22961, N10171);
nand NAND2 (N22971, N22969, N1105);
nand NAND3 (N22972, N22967, N15386, N2356);
not NOT1 (N22973, N22972);
nand NAND2 (N22974, N22973, N1966);
and AND4 (N22975, N22968, N10350, N16564, N19592);
not NOT1 (N22976, N22966);
xor XOR2 (N22977, N22974, N11532);
nand NAND4 (N22978, N22960, N15063, N21134, N17541);
nor NOR3 (N22979, N22964, N8336, N20156);
nor NOR2 (N22980, N22937, N10067);
nand NAND2 (N22981, N22971, N1329);
nor NOR2 (N22982, N22980, N4750);
nand NAND2 (N22983, N22965, N14821);
buf BUF1 (N22984, N22976);
buf BUF1 (N22985, N22977);
not NOT1 (N22986, N22984);
xor XOR2 (N22987, N22981, N11769);
nand NAND2 (N22988, N22957, N21580);
not NOT1 (N22989, N22970);
nor NOR4 (N22990, N22987, N5849, N2580, N6463);
xor XOR2 (N22991, N22988, N14057);
and AND2 (N22992, N22979, N4072);
xor XOR2 (N22993, N22992, N13802);
or OR4 (N22994, N22985, N13464, N20202, N1340);
and AND4 (N22995, N22983, N1661, N6536, N18288);
buf BUF1 (N22996, N22994);
not NOT1 (N22997, N22991);
nand NAND3 (N22998, N22996, N2706, N15154);
xor XOR2 (N22999, N22990, N8215);
or OR3 (N23000, N22982, N16964, N12109);
xor XOR2 (N23001, N22978, N16921);
buf BUF1 (N23002, N22999);
or OR3 (N23003, N22997, N1382, N18139);
nand NAND4 (N23004, N22975, N14782, N22182, N10209);
nor NOR4 (N23005, N23000, N3571, N18395, N14001);
nor NOR4 (N23006, N23004, N10400, N8084, N13883);
xor XOR2 (N23007, N22995, N18519);
and AND4 (N23008, N22989, N17781, N1769, N294);
nand NAND2 (N23009, N23003, N5115);
or OR2 (N23010, N23008, N7712);
or OR3 (N23011, N22998, N19364, N18053);
not NOT1 (N23012, N23006);
buf BUF1 (N23013, N23009);
nor NOR2 (N23014, N22986, N8586);
xor XOR2 (N23015, N23001, N2282);
nor NOR3 (N23016, N23014, N15884, N10273);
nand NAND2 (N23017, N23011, N15962);
xor XOR2 (N23018, N23010, N5109);
and AND2 (N23019, N23012, N547);
not NOT1 (N23020, N23018);
or OR2 (N23021, N23007, N17477);
buf BUF1 (N23022, N23002);
and AND4 (N23023, N23019, N9268, N10987, N8532);
buf BUF1 (N23024, N23021);
nor NOR3 (N23025, N23023, N20473, N22161);
nor NOR4 (N23026, N23020, N12901, N7530, N22712);
or OR2 (N23027, N23026, N9937);
or OR4 (N23028, N23027, N9937, N14514, N20742);
nand NAND2 (N23029, N23005, N10292);
not NOT1 (N23030, N23024);
xor XOR2 (N23031, N23017, N13824);
buf BUF1 (N23032, N23022);
or OR2 (N23033, N23029, N20890);
not NOT1 (N23034, N23016);
or OR2 (N23035, N23033, N14818);
nor NOR2 (N23036, N23035, N1423);
not NOT1 (N23037, N23030);
or OR4 (N23038, N23028, N10688, N4673, N5561);
buf BUF1 (N23039, N23038);
not NOT1 (N23040, N23036);
xor XOR2 (N23041, N23031, N218);
and AND2 (N23042, N23015, N4353);
xor XOR2 (N23043, N23040, N18411);
and AND4 (N23044, N23037, N2012, N13708, N8115);
not NOT1 (N23045, N23044);
or OR2 (N23046, N23032, N16389);
and AND2 (N23047, N23042, N15666);
nand NAND3 (N23048, N23039, N3450, N2678);
nor NOR4 (N23049, N23025, N20628, N19542, N2312);
nand NAND2 (N23050, N23013, N8350);
nand NAND4 (N23051, N23034, N19809, N6331, N13398);
or OR3 (N23052, N23046, N14582, N14583);
not NOT1 (N23053, N23048);
or OR4 (N23054, N23053, N4194, N5395, N1979);
nor NOR2 (N23055, N23050, N11816);
buf BUF1 (N23056, N23054);
xor XOR2 (N23057, N23041, N7230);
not NOT1 (N23058, N22993);
or OR2 (N23059, N23049, N12243);
buf BUF1 (N23060, N23058);
buf BUF1 (N23061, N23045);
buf BUF1 (N23062, N23055);
nor NOR3 (N23063, N23051, N21544, N2753);
xor XOR2 (N23064, N23062, N13253);
not NOT1 (N23065, N23052);
not NOT1 (N23066, N23063);
nand NAND4 (N23067, N23043, N21786, N21983, N22805);
nand NAND4 (N23068, N23064, N8962, N642, N3819);
not NOT1 (N23069, N23047);
buf BUF1 (N23070, N23069);
not NOT1 (N23071, N23061);
or OR2 (N23072, N23057, N11729);
nand NAND3 (N23073, N23067, N20710, N8514);
not NOT1 (N23074, N23073);
nor NOR4 (N23075, N23070, N3300, N15929, N3584);
buf BUF1 (N23076, N23071);
or OR2 (N23077, N23060, N2639);
or OR3 (N23078, N23059, N1418, N16386);
xor XOR2 (N23079, N23077, N18246);
buf BUF1 (N23080, N23065);
or OR2 (N23081, N23056, N811);
or OR3 (N23082, N23072, N15863, N3214);
nor NOR2 (N23083, N23080, N20375);
not NOT1 (N23084, N23068);
buf BUF1 (N23085, N23075);
not NOT1 (N23086, N23079);
not NOT1 (N23087, N23076);
nor NOR4 (N23088, N23084, N13827, N20645, N15974);
and AND4 (N23089, N23085, N12969, N1774, N16649);
buf BUF1 (N23090, N23083);
or OR2 (N23091, N23089, N8826);
nor NOR2 (N23092, N23081, N23041);
xor XOR2 (N23093, N23091, N3468);
xor XOR2 (N23094, N23078, N20309);
and AND3 (N23095, N23094, N4568, N22249);
xor XOR2 (N23096, N23074, N22386);
xor XOR2 (N23097, N23090, N8936);
and AND2 (N23098, N23092, N2242);
xor XOR2 (N23099, N23087, N8308);
buf BUF1 (N23100, N23097);
not NOT1 (N23101, N23099);
nor NOR2 (N23102, N23088, N4371);
nand NAND4 (N23103, N23082, N4848, N19278, N16909);
nor NOR3 (N23104, N23101, N7059, N4403);
or OR4 (N23105, N23100, N13277, N13571, N22732);
nor NOR2 (N23106, N23098, N2832);
nand NAND4 (N23107, N23102, N12385, N2387, N13999);
or OR3 (N23108, N23107, N6028, N16186);
nor NOR4 (N23109, N23096, N1999, N11771, N17452);
and AND3 (N23110, N23086, N23048, N6564);
not NOT1 (N23111, N23066);
not NOT1 (N23112, N23105);
or OR2 (N23113, N23095, N1530);
buf BUF1 (N23114, N23106);
or OR3 (N23115, N23104, N99, N4514);
buf BUF1 (N23116, N23109);
nor NOR3 (N23117, N23116, N11861, N14334);
nand NAND4 (N23118, N23093, N8648, N14897, N435);
xor XOR2 (N23119, N23112, N21316);
and AND2 (N23120, N23115, N11190);
xor XOR2 (N23121, N23114, N20050);
not NOT1 (N23122, N23111);
and AND3 (N23123, N23110, N633, N8029);
or OR3 (N23124, N23122, N21677, N3903);
nor NOR3 (N23125, N23120, N22621, N4322);
not NOT1 (N23126, N23103);
nor NOR4 (N23127, N23125, N9807, N7392, N3235);
or OR4 (N23128, N23127, N6126, N18744, N9272);
and AND3 (N23129, N23121, N3134, N4175);
nor NOR4 (N23130, N23129, N2291, N3385, N23080);
nand NAND4 (N23131, N23118, N12541, N2053, N21963);
and AND3 (N23132, N23124, N1066, N11542);
and AND4 (N23133, N23131, N22782, N953, N17282);
buf BUF1 (N23134, N23113);
xor XOR2 (N23135, N23134, N6926);
and AND3 (N23136, N23117, N9575, N18059);
nor NOR2 (N23137, N23126, N16989);
buf BUF1 (N23138, N23136);
xor XOR2 (N23139, N23128, N3888);
not NOT1 (N23140, N23133);
nand NAND2 (N23141, N23132, N18720);
buf BUF1 (N23142, N23140);
xor XOR2 (N23143, N23119, N2948);
and AND2 (N23144, N23138, N10849);
nor NOR4 (N23145, N23142, N14965, N16028, N16157);
not NOT1 (N23146, N23145);
nor NOR2 (N23147, N23141, N19165);
not NOT1 (N23148, N23108);
buf BUF1 (N23149, N23146);
not NOT1 (N23150, N23147);
nand NAND3 (N23151, N23137, N13182, N8683);
or OR2 (N23152, N23139, N13094);
not NOT1 (N23153, N23151);
nor NOR4 (N23154, N23143, N11032, N8963, N19550);
xor XOR2 (N23155, N23149, N16481);
and AND2 (N23156, N23155, N12386);
xor XOR2 (N23157, N23130, N2472);
and AND4 (N23158, N23123, N18726, N5639, N9778);
not NOT1 (N23159, N23157);
xor XOR2 (N23160, N23150, N6383);
nand NAND2 (N23161, N23135, N20799);
and AND4 (N23162, N23148, N20408, N17402, N15578);
and AND4 (N23163, N23159, N6479, N5254, N11785);
not NOT1 (N23164, N23144);
nor NOR3 (N23165, N23163, N4031, N10804);
or OR3 (N23166, N23161, N19646, N2868);
or OR4 (N23167, N23162, N19092, N2847, N16067);
nor NOR4 (N23168, N23166, N6669, N17903, N19640);
or OR3 (N23169, N23158, N6195, N18712);
buf BUF1 (N23170, N23167);
buf BUF1 (N23171, N23154);
xor XOR2 (N23172, N23171, N17098);
xor XOR2 (N23173, N23153, N20878);
and AND2 (N23174, N23173, N5841);
or OR2 (N23175, N23168, N7635);
or OR4 (N23176, N23165, N5774, N17397, N16529);
nand NAND2 (N23177, N23164, N7250);
nor NOR2 (N23178, N23177, N21496);
buf BUF1 (N23179, N23178);
or OR2 (N23180, N23175, N13831);
nand NAND4 (N23181, N23169, N15737, N6618, N22366);
and AND3 (N23182, N23160, N11804, N5554);
nor NOR3 (N23183, N23172, N13524, N8604);
or OR4 (N23184, N23183, N6276, N19291, N3575);
buf BUF1 (N23185, N23174);
or OR4 (N23186, N23176, N5013, N5000, N20742);
and AND4 (N23187, N23182, N4390, N5518, N3264);
nor NOR4 (N23188, N23181, N20372, N8316, N8717);
nand NAND4 (N23189, N23170, N14536, N9494, N155);
nor NOR2 (N23190, N23185, N6278);
or OR4 (N23191, N23180, N10266, N22169, N23025);
not NOT1 (N23192, N23188);
not NOT1 (N23193, N23191);
buf BUF1 (N23194, N23192);
nor NOR3 (N23195, N23190, N7217, N6073);
buf BUF1 (N23196, N23184);
or OR4 (N23197, N23189, N6531, N9975, N15389);
or OR2 (N23198, N23193, N1515);
nand NAND3 (N23199, N23186, N11109, N21692);
not NOT1 (N23200, N23187);
xor XOR2 (N23201, N23196, N1912);
not NOT1 (N23202, N23197);
buf BUF1 (N23203, N23194);
and AND4 (N23204, N23199, N11237, N2356, N16324);
buf BUF1 (N23205, N23179);
and AND4 (N23206, N23198, N4353, N6375, N16557);
or OR2 (N23207, N23206, N5131);
not NOT1 (N23208, N23205);
nand NAND2 (N23209, N23200, N14023);
nor NOR2 (N23210, N23204, N2175);
and AND3 (N23211, N23207, N3823, N21768);
not NOT1 (N23212, N23202);
or OR2 (N23213, N23201, N9179);
and AND2 (N23214, N23210, N15337);
or OR4 (N23215, N23152, N6748, N3490, N16103);
nor NOR2 (N23216, N23214, N17957);
nand NAND2 (N23217, N23216, N5955);
buf BUF1 (N23218, N23217);
and AND3 (N23219, N23203, N7972, N9242);
and AND2 (N23220, N23211, N5933);
not NOT1 (N23221, N23195);
buf BUF1 (N23222, N23215);
nand NAND2 (N23223, N23220, N6726);
and AND3 (N23224, N23221, N12830, N10511);
xor XOR2 (N23225, N23219, N8742);
not NOT1 (N23226, N23209);
nor NOR4 (N23227, N23223, N12971, N12948, N15410);
and AND3 (N23228, N23222, N2763, N1458);
xor XOR2 (N23229, N23225, N4753);
xor XOR2 (N23230, N23208, N15455);
nor NOR4 (N23231, N23212, N71, N14823, N6594);
nand NAND2 (N23232, N23231, N21150);
nand NAND2 (N23233, N23156, N7360);
not NOT1 (N23234, N23227);
buf BUF1 (N23235, N23228);
buf BUF1 (N23236, N23218);
buf BUF1 (N23237, N23229);
and AND2 (N23238, N23224, N19965);
or OR3 (N23239, N23226, N17628, N14107);
and AND4 (N23240, N23230, N7576, N21036, N7302);
xor XOR2 (N23241, N23236, N4595);
buf BUF1 (N23242, N23238);
nand NAND2 (N23243, N23241, N7532);
buf BUF1 (N23244, N23237);
nand NAND3 (N23245, N23234, N19282, N21761);
nor NOR4 (N23246, N23243, N3078, N10988, N8965);
and AND3 (N23247, N23235, N10975, N21927);
nand NAND3 (N23248, N23247, N21354, N15404);
nand NAND4 (N23249, N23240, N20221, N8608, N18987);
or OR4 (N23250, N23249, N19173, N5569, N15285);
or OR2 (N23251, N23239, N14056);
and AND4 (N23252, N23251, N1660, N17982, N9352);
nor NOR3 (N23253, N23250, N1516, N20827);
nand NAND4 (N23254, N23232, N21851, N17627, N5281);
or OR4 (N23255, N23252, N3876, N20146, N14401);
buf BUF1 (N23256, N23244);
and AND3 (N23257, N23242, N22970, N17294);
nor NOR2 (N23258, N23233, N19401);
xor XOR2 (N23259, N23256, N15631);
not NOT1 (N23260, N23245);
or OR3 (N23261, N23248, N5296, N596);
and AND4 (N23262, N23261, N22533, N14689, N1674);
not NOT1 (N23263, N23253);
and AND4 (N23264, N23257, N19271, N6870, N16059);
nor NOR3 (N23265, N23258, N1167, N18421);
xor XOR2 (N23266, N23255, N20638);
nand NAND2 (N23267, N23266, N15968);
nand NAND2 (N23268, N23213, N17047);
or OR2 (N23269, N23259, N5488);
or OR3 (N23270, N23263, N10038, N20095);
nand NAND2 (N23271, N23262, N22415);
and AND2 (N23272, N23264, N14139);
buf BUF1 (N23273, N23254);
not NOT1 (N23274, N23269);
nor NOR4 (N23275, N23268, N1653, N17741, N20826);
and AND3 (N23276, N23267, N5651, N19615);
xor XOR2 (N23277, N23270, N10305);
xor XOR2 (N23278, N23276, N15357);
nand NAND2 (N23279, N23278, N14551);
buf BUF1 (N23280, N23274);
not NOT1 (N23281, N23260);
and AND3 (N23282, N23265, N22787, N1034);
nand NAND2 (N23283, N23282, N10187);
or OR4 (N23284, N23275, N12649, N21344, N2689);
not NOT1 (N23285, N23281);
nand NAND4 (N23286, N23273, N13359, N9190, N12385);
or OR4 (N23287, N23280, N223, N6981, N12969);
xor XOR2 (N23288, N23284, N8806);
not NOT1 (N23289, N23279);
buf BUF1 (N23290, N23277);
nor NOR4 (N23291, N23246, N10604, N19704, N8368);
nor NOR4 (N23292, N23283, N16033, N4224, N11433);
nand NAND4 (N23293, N23286, N10105, N4598, N23056);
and AND2 (N23294, N23287, N22938);
not NOT1 (N23295, N23294);
nand NAND4 (N23296, N23295, N21740, N23167, N9900);
or OR2 (N23297, N23272, N18698);
or OR4 (N23298, N23291, N3119, N3056, N5285);
nand NAND4 (N23299, N23297, N4231, N14355, N7573);
nor NOR2 (N23300, N23296, N18745);
buf BUF1 (N23301, N23292);
xor XOR2 (N23302, N23285, N1951);
not NOT1 (N23303, N23300);
or OR2 (N23304, N23290, N11037);
and AND3 (N23305, N23299, N14537, N15449);
xor XOR2 (N23306, N23298, N1789);
nand NAND4 (N23307, N23303, N447, N6739, N22767);
nor NOR2 (N23308, N23293, N21544);
and AND4 (N23309, N23288, N20839, N6468, N2012);
nor NOR2 (N23310, N23301, N14823);
xor XOR2 (N23311, N23302, N3650);
xor XOR2 (N23312, N23289, N10039);
nand NAND2 (N23313, N23308, N3619);
and AND3 (N23314, N23307, N20719, N16224);
and AND4 (N23315, N23311, N1037, N7952, N7130);
buf BUF1 (N23316, N23310);
not NOT1 (N23317, N23316);
xor XOR2 (N23318, N23271, N9998);
not NOT1 (N23319, N23305);
or OR4 (N23320, N23304, N8403, N7987, N5983);
or OR3 (N23321, N23314, N6827, N17608);
buf BUF1 (N23322, N23312);
or OR3 (N23323, N23322, N20966, N632);
xor XOR2 (N23324, N23320, N14675);
and AND3 (N23325, N23306, N16827, N5351);
nand NAND4 (N23326, N23313, N5670, N7737, N16907);
not NOT1 (N23327, N23323);
or OR4 (N23328, N23317, N21502, N578, N21704);
and AND4 (N23329, N23326, N5032, N14437, N15799);
and AND2 (N23330, N23319, N9729);
not NOT1 (N23331, N23318);
nor NOR3 (N23332, N23328, N12093, N20775);
not NOT1 (N23333, N23329);
not NOT1 (N23334, N23324);
buf BUF1 (N23335, N23330);
buf BUF1 (N23336, N23327);
or OR4 (N23337, N23315, N13180, N6732, N10754);
buf BUF1 (N23338, N23334);
or OR4 (N23339, N23338, N13121, N12522, N16701);
or OR4 (N23340, N23336, N2021, N17460, N13102);
nor NOR3 (N23341, N23337, N10340, N21923);
buf BUF1 (N23342, N23333);
or OR3 (N23343, N23331, N9156, N13744);
nor NOR3 (N23344, N23339, N6366, N254);
buf BUF1 (N23345, N23341);
nand NAND4 (N23346, N23340, N1798, N7747, N17061);
and AND4 (N23347, N23345, N20600, N11901, N410);
nand NAND2 (N23348, N23335, N12805);
nand NAND4 (N23349, N23347, N7300, N17975, N9761);
xor XOR2 (N23350, N23309, N21117);
and AND2 (N23351, N23342, N15896);
or OR2 (N23352, N23348, N9354);
buf BUF1 (N23353, N23325);
or OR4 (N23354, N23343, N19290, N14674, N7417);
not NOT1 (N23355, N23346);
and AND2 (N23356, N23321, N19907);
nor NOR2 (N23357, N23355, N1);
or OR3 (N23358, N23356, N4787, N18926);
nor NOR3 (N23359, N23351, N12838, N13130);
and AND2 (N23360, N23349, N21686);
nor NOR3 (N23361, N23352, N17177, N945);
nor NOR2 (N23362, N23354, N13616);
and AND4 (N23363, N23344, N14251, N14164, N23221);
or OR4 (N23364, N23360, N4725, N22587, N2228);
or OR3 (N23365, N23362, N11356, N3765);
and AND4 (N23366, N23359, N7536, N13629, N4849);
or OR2 (N23367, N23363, N11328);
and AND2 (N23368, N23361, N18061);
and AND4 (N23369, N23365, N8720, N2601, N5367);
nor NOR2 (N23370, N23332, N17301);
nand NAND4 (N23371, N23370, N15476, N4981, N9735);
buf BUF1 (N23372, N23350);
or OR4 (N23373, N23366, N14752, N20500, N22379);
not NOT1 (N23374, N23358);
and AND2 (N23375, N23367, N9538);
xor XOR2 (N23376, N23373, N11343);
nand NAND2 (N23377, N23375, N11093);
xor XOR2 (N23378, N23369, N12399);
nand NAND4 (N23379, N23372, N10162, N5314, N21312);
buf BUF1 (N23380, N23379);
nand NAND4 (N23381, N23378, N1022, N634, N2523);
nand NAND4 (N23382, N23374, N17139, N22208, N10450);
and AND2 (N23383, N23376, N2725);
xor XOR2 (N23384, N23381, N1391);
nor NOR4 (N23385, N23357, N6802, N11821, N11505);
buf BUF1 (N23386, N23371);
and AND3 (N23387, N23386, N21849, N14101);
xor XOR2 (N23388, N23387, N2922);
buf BUF1 (N23389, N23380);
xor XOR2 (N23390, N23382, N12338);
nor NOR3 (N23391, N23368, N22233, N2629);
buf BUF1 (N23392, N23389);
nor NOR4 (N23393, N23391, N9686, N18633, N5885);
or OR3 (N23394, N23383, N6377, N10485);
and AND3 (N23395, N23364, N5375, N7078);
buf BUF1 (N23396, N23392);
xor XOR2 (N23397, N23395, N22591);
xor XOR2 (N23398, N23384, N15486);
nor NOR3 (N23399, N23353, N16603, N22364);
not NOT1 (N23400, N23398);
nor NOR3 (N23401, N23397, N20056, N13096);
or OR3 (N23402, N23394, N2194, N2668);
nor NOR3 (N23403, N23402, N20416, N23355);
not NOT1 (N23404, N23400);
nor NOR2 (N23405, N23403, N2826);
buf BUF1 (N23406, N23385);
nand NAND2 (N23407, N23405, N16925);
nand NAND2 (N23408, N23407, N11901);
nand NAND3 (N23409, N23388, N3196, N22676);
and AND2 (N23410, N23404, N13037);
not NOT1 (N23411, N23399);
nand NAND4 (N23412, N23410, N4714, N19778, N7813);
and AND3 (N23413, N23401, N6610, N16203);
nor NOR3 (N23414, N23377, N2288, N2217);
nand NAND4 (N23415, N23390, N6936, N15392, N5017);
xor XOR2 (N23416, N23412, N6597);
buf BUF1 (N23417, N23413);
or OR3 (N23418, N23409, N11112, N23188);
not NOT1 (N23419, N23396);
and AND4 (N23420, N23408, N2161, N2908, N7756);
and AND3 (N23421, N23419, N14, N8361);
xor XOR2 (N23422, N23414, N14276);
buf BUF1 (N23423, N23415);
buf BUF1 (N23424, N23411);
or OR3 (N23425, N23416, N12496, N7131);
and AND4 (N23426, N23424, N6586, N4758, N13771);
not NOT1 (N23427, N23418);
nor NOR2 (N23428, N23425, N20729);
xor XOR2 (N23429, N23423, N22496);
buf BUF1 (N23430, N23420);
nand NAND3 (N23431, N23422, N8879, N164);
nor NOR4 (N23432, N23431, N19623, N19659, N5650);
and AND2 (N23433, N23427, N20777);
buf BUF1 (N23434, N23426);
xor XOR2 (N23435, N23430, N9810);
or OR2 (N23436, N23417, N13590);
nand NAND3 (N23437, N23433, N13834, N3684);
not NOT1 (N23438, N23428);
nand NAND4 (N23439, N23434, N6147, N14512, N7695);
not NOT1 (N23440, N23429);
or OR2 (N23441, N23432, N14811);
not NOT1 (N23442, N23435);
nor NOR2 (N23443, N23393, N23427);
and AND4 (N23444, N23421, N14081, N12847, N19738);
or OR4 (N23445, N23406, N22836, N9545, N17553);
buf BUF1 (N23446, N23444);
nand NAND2 (N23447, N23441, N833);
xor XOR2 (N23448, N23442, N17182);
xor XOR2 (N23449, N23438, N2665);
nor NOR4 (N23450, N23448, N12531, N9122, N12396);
buf BUF1 (N23451, N23437);
nand NAND3 (N23452, N23447, N22293, N21510);
nand NAND3 (N23453, N23443, N21738, N1722);
xor XOR2 (N23454, N23449, N20472);
buf BUF1 (N23455, N23454);
nand NAND3 (N23456, N23439, N1022, N6737);
buf BUF1 (N23457, N23456);
or OR3 (N23458, N23436, N10980, N9799);
nand NAND3 (N23459, N23440, N15094, N19129);
xor XOR2 (N23460, N23450, N17228);
and AND3 (N23461, N23460, N13263, N16747);
or OR4 (N23462, N23446, N2694, N19865, N20940);
nor NOR2 (N23463, N23461, N6493);
not NOT1 (N23464, N23458);
or OR4 (N23465, N23462, N18328, N5139, N5559);
and AND4 (N23466, N23459, N3173, N2070, N20453);
not NOT1 (N23467, N23463);
xor XOR2 (N23468, N23451, N23068);
buf BUF1 (N23469, N23453);
or OR4 (N23470, N23455, N9049, N11193, N10131);
buf BUF1 (N23471, N23470);
and AND3 (N23472, N23465, N4991, N21743);
xor XOR2 (N23473, N23445, N19138);
or OR2 (N23474, N23464, N4365);
and AND2 (N23475, N23471, N5605);
nor NOR4 (N23476, N23468, N14754, N10439, N13573);
nand NAND2 (N23477, N23457, N17288);
or OR2 (N23478, N23469, N13590);
and AND4 (N23479, N23473, N23442, N13658, N11245);
not NOT1 (N23480, N23452);
buf BUF1 (N23481, N23475);
xor XOR2 (N23482, N23478, N1808);
buf BUF1 (N23483, N23472);
nand NAND4 (N23484, N23474, N2940, N709, N15484);
nor NOR2 (N23485, N23483, N10873);
or OR3 (N23486, N23484, N4396, N22039);
and AND4 (N23487, N23477, N244, N16953, N18451);
buf BUF1 (N23488, N23479);
not NOT1 (N23489, N23488);
or OR4 (N23490, N23489, N14750, N16622, N1837);
nand NAND3 (N23491, N23480, N3796, N11312);
and AND2 (N23492, N23491, N6419);
nand NAND2 (N23493, N23485, N6279);
nand NAND2 (N23494, N23466, N20245);
not NOT1 (N23495, N23494);
buf BUF1 (N23496, N23482);
buf BUF1 (N23497, N23476);
and AND3 (N23498, N23490, N904, N19544);
not NOT1 (N23499, N23467);
not NOT1 (N23500, N23497);
buf BUF1 (N23501, N23496);
xor XOR2 (N23502, N23487, N2031);
buf BUF1 (N23503, N23502);
buf BUF1 (N23504, N23498);
not NOT1 (N23505, N23486);
or OR3 (N23506, N23481, N14879, N18541);
xor XOR2 (N23507, N23504, N19309);
not NOT1 (N23508, N23507);
nor NOR2 (N23509, N23501, N16338);
buf BUF1 (N23510, N23503);
buf BUF1 (N23511, N23509);
not NOT1 (N23512, N23500);
or OR4 (N23513, N23492, N9539, N13459, N21195);
nor NOR4 (N23514, N23495, N23072, N21470, N10446);
not NOT1 (N23515, N23513);
nor NOR2 (N23516, N23514, N1138);
xor XOR2 (N23517, N23505, N23161);
buf BUF1 (N23518, N23506);
nor NOR4 (N23519, N23517, N10387, N13459, N22973);
and AND3 (N23520, N23518, N4382, N21297);
nand NAND2 (N23521, N23511, N16573);
nand NAND2 (N23522, N23519, N15199);
buf BUF1 (N23523, N23515);
and AND3 (N23524, N23522, N6145, N12866);
nor NOR3 (N23525, N23499, N17627, N20034);
xor XOR2 (N23526, N23508, N4867);
and AND3 (N23527, N23523, N18192, N2975);
nand NAND2 (N23528, N23493, N6723);
and AND3 (N23529, N23528, N11642, N21977);
and AND4 (N23530, N23512, N19466, N23131, N14936);
and AND2 (N23531, N23524, N9522);
xor XOR2 (N23532, N23531, N9819);
not NOT1 (N23533, N23510);
not NOT1 (N23534, N23526);
xor XOR2 (N23535, N23516, N8825);
nor NOR2 (N23536, N23532, N4856);
and AND2 (N23537, N23534, N7394);
nand NAND3 (N23538, N23530, N15778, N11088);
nand NAND4 (N23539, N23529, N17247, N16083, N15828);
or OR2 (N23540, N23527, N5891);
or OR3 (N23541, N23535, N15736, N14096);
not NOT1 (N23542, N23537);
nor NOR4 (N23543, N23540, N7994, N4116, N3713);
or OR3 (N23544, N23541, N13565, N12933);
buf BUF1 (N23545, N23533);
buf BUF1 (N23546, N23545);
nand NAND4 (N23547, N23539, N22445, N20713, N9481);
not NOT1 (N23548, N23525);
xor XOR2 (N23549, N23547, N14968);
nor NOR4 (N23550, N23536, N650, N23037, N8506);
and AND3 (N23551, N23538, N9304, N6368);
buf BUF1 (N23552, N23548);
not NOT1 (N23553, N23520);
and AND4 (N23554, N23550, N9081, N10090, N5420);
not NOT1 (N23555, N23544);
xor XOR2 (N23556, N23546, N22968);
nand NAND3 (N23557, N23556, N10862, N11683);
buf BUF1 (N23558, N23521);
or OR2 (N23559, N23542, N21620);
buf BUF1 (N23560, N23553);
or OR4 (N23561, N23560, N12033, N6047, N7278);
buf BUF1 (N23562, N23558);
or OR2 (N23563, N23554, N14437);
buf BUF1 (N23564, N23549);
nand NAND3 (N23565, N23551, N15485, N15836);
or OR2 (N23566, N23559, N793);
xor XOR2 (N23567, N23566, N5204);
and AND4 (N23568, N23543, N14732, N22561, N7210);
buf BUF1 (N23569, N23568);
or OR2 (N23570, N23567, N5967);
xor XOR2 (N23571, N23563, N15589);
xor XOR2 (N23572, N23552, N19898);
or OR3 (N23573, N23570, N10869, N23023);
and AND3 (N23574, N23557, N19001, N7977);
nand NAND3 (N23575, N23571, N6263, N151);
xor XOR2 (N23576, N23561, N18723);
xor XOR2 (N23577, N23574, N812);
and AND2 (N23578, N23572, N19405);
nand NAND4 (N23579, N23575, N18651, N21886, N459);
or OR3 (N23580, N23565, N5514, N21706);
not NOT1 (N23581, N23579);
buf BUF1 (N23582, N23581);
nor NOR3 (N23583, N23580, N7315, N2522);
and AND2 (N23584, N23569, N3062);
not NOT1 (N23585, N23564);
nor NOR3 (N23586, N23576, N15331, N4314);
nand NAND2 (N23587, N23584, N5300);
or OR3 (N23588, N23577, N14215, N14274);
nand NAND3 (N23589, N23582, N20294, N4694);
or OR3 (N23590, N23555, N21750, N22040);
and AND2 (N23591, N23573, N14967);
buf BUF1 (N23592, N23586);
not NOT1 (N23593, N23585);
buf BUF1 (N23594, N23593);
not NOT1 (N23595, N23591);
xor XOR2 (N23596, N23594, N20675);
nor NOR2 (N23597, N23592, N16810);
and AND3 (N23598, N23588, N227, N19183);
nand NAND3 (N23599, N23596, N13618, N1228);
and AND3 (N23600, N23595, N4221, N13916);
nand NAND2 (N23601, N23578, N6536);
xor XOR2 (N23602, N23583, N8678);
or OR2 (N23603, N23600, N16210);
or OR2 (N23604, N23601, N9302);
nor NOR3 (N23605, N23587, N3969, N6380);
and AND2 (N23606, N23604, N9443);
and AND4 (N23607, N23597, N4799, N9122, N21035);
xor XOR2 (N23608, N23589, N15990);
nor NOR4 (N23609, N23602, N19599, N16222, N3428);
or OR2 (N23610, N23606, N16650);
xor XOR2 (N23611, N23599, N8914);
and AND2 (N23612, N23605, N13169);
not NOT1 (N23613, N23598);
and AND2 (N23614, N23590, N15284);
nand NAND2 (N23615, N23608, N19812);
or OR2 (N23616, N23562, N12705);
nand NAND2 (N23617, N23603, N20397);
buf BUF1 (N23618, N23610);
not NOT1 (N23619, N23617);
not NOT1 (N23620, N23607);
and AND4 (N23621, N23620, N19643, N10645, N7102);
and AND3 (N23622, N23616, N21655, N19779);
not NOT1 (N23623, N23611);
or OR3 (N23624, N23622, N22700, N14043);
nand NAND3 (N23625, N23613, N14601, N22386);
and AND4 (N23626, N23621, N16202, N2649, N12902);
not NOT1 (N23627, N23623);
not NOT1 (N23628, N23614);
not NOT1 (N23629, N23626);
xor XOR2 (N23630, N23618, N21732);
xor XOR2 (N23631, N23615, N9154);
nand NAND2 (N23632, N23628, N16686);
not NOT1 (N23633, N23629);
xor XOR2 (N23634, N23612, N11304);
nor NOR2 (N23635, N23634, N11579);
and AND4 (N23636, N23625, N8873, N13974, N14271);
and AND3 (N23637, N23633, N11495, N12649);
nor NOR3 (N23638, N23609, N16431, N5243);
or OR4 (N23639, N23632, N1765, N2718, N354);
buf BUF1 (N23640, N23619);
or OR2 (N23641, N23627, N8344);
nand NAND4 (N23642, N23636, N9320, N10629, N22080);
xor XOR2 (N23643, N23639, N20066);
nand NAND2 (N23644, N23638, N6078);
xor XOR2 (N23645, N23640, N6230);
or OR2 (N23646, N23643, N11252);
buf BUF1 (N23647, N23642);
xor XOR2 (N23648, N23624, N6018);
nor NOR4 (N23649, N23646, N23175, N5764, N6674);
buf BUF1 (N23650, N23630);
and AND4 (N23651, N23637, N15686, N10384, N18479);
and AND3 (N23652, N23648, N9603, N776);
xor XOR2 (N23653, N23647, N16308);
nor NOR3 (N23654, N23645, N1440, N10177);
not NOT1 (N23655, N23653);
nand NAND4 (N23656, N23649, N13223, N3973, N219);
buf BUF1 (N23657, N23635);
and AND2 (N23658, N23654, N22109);
not NOT1 (N23659, N23652);
buf BUF1 (N23660, N23641);
buf BUF1 (N23661, N23655);
not NOT1 (N23662, N23644);
or OR4 (N23663, N23662, N16536, N19590, N2660);
buf BUF1 (N23664, N23651);
buf BUF1 (N23665, N23631);
nor NOR4 (N23666, N23657, N755, N22779, N1590);
and AND4 (N23667, N23666, N11580, N66, N16651);
nor NOR4 (N23668, N23659, N9564, N12640, N21629);
not NOT1 (N23669, N23665);
not NOT1 (N23670, N23667);
nand NAND2 (N23671, N23650, N20390);
nand NAND4 (N23672, N23658, N13176, N3061, N15414);
not NOT1 (N23673, N23663);
buf BUF1 (N23674, N23668);
buf BUF1 (N23675, N23656);
nand NAND3 (N23676, N23673, N12763, N5747);
and AND3 (N23677, N23671, N21940, N682);
nand NAND2 (N23678, N23661, N11346);
not NOT1 (N23679, N23677);
buf BUF1 (N23680, N23675);
nor NOR2 (N23681, N23669, N6433);
xor XOR2 (N23682, N23679, N4110);
nor NOR4 (N23683, N23660, N7989, N16318, N23654);
xor XOR2 (N23684, N23683, N5459);
buf BUF1 (N23685, N23674);
and AND4 (N23686, N23672, N14335, N634, N10628);
and AND2 (N23687, N23676, N7959);
buf BUF1 (N23688, N23686);
or OR3 (N23689, N23685, N14255, N3302);
and AND2 (N23690, N23689, N5467);
nand NAND2 (N23691, N23670, N4470);
nand NAND4 (N23692, N23680, N18402, N22691, N21807);
nor NOR4 (N23693, N23681, N9189, N16546, N7005);
or OR3 (N23694, N23691, N12970, N22356);
not NOT1 (N23695, N23688);
nand NAND4 (N23696, N23682, N2626, N19772, N2468);
xor XOR2 (N23697, N23696, N9356);
nand NAND3 (N23698, N23684, N15272, N9212);
xor XOR2 (N23699, N23693, N8813);
and AND4 (N23700, N23694, N19455, N5090, N11011);
buf BUF1 (N23701, N23678);
or OR4 (N23702, N23692, N20005, N5219, N4882);
xor XOR2 (N23703, N23701, N20678);
buf BUF1 (N23704, N23699);
and AND3 (N23705, N23703, N12240, N3481);
nor NOR3 (N23706, N23690, N2962, N13262);
and AND4 (N23707, N23695, N16021, N3801, N6571);
buf BUF1 (N23708, N23707);
nand NAND3 (N23709, N23664, N6415, N7032);
or OR3 (N23710, N23700, N22664, N21933);
or OR2 (N23711, N23698, N2585);
not NOT1 (N23712, N23705);
or OR4 (N23713, N23706, N3141, N23320, N10240);
nor NOR2 (N23714, N23704, N7592);
nand NAND4 (N23715, N23710, N16128, N23182, N1122);
buf BUF1 (N23716, N23687);
or OR2 (N23717, N23708, N5490);
not NOT1 (N23718, N23713);
and AND4 (N23719, N23709, N14917, N16562, N19517);
or OR3 (N23720, N23716, N20385, N4940);
nand NAND4 (N23721, N23702, N6644, N9519, N2556);
and AND3 (N23722, N23718, N12477, N16895);
nand NAND2 (N23723, N23721, N15680);
or OR3 (N23724, N23697, N22912, N18996);
nor NOR4 (N23725, N23712, N20759, N7526, N17517);
nand NAND2 (N23726, N23717, N14078);
nand NAND2 (N23727, N23725, N12216);
not NOT1 (N23728, N23727);
or OR4 (N23729, N23724, N11037, N2127, N13089);
nor NOR3 (N23730, N23720, N12956, N4590);
not NOT1 (N23731, N23728);
buf BUF1 (N23732, N23731);
not NOT1 (N23733, N23732);
and AND3 (N23734, N23719, N4556, N9206);
not NOT1 (N23735, N23711);
buf BUF1 (N23736, N23734);
nor NOR3 (N23737, N23736, N22464, N5887);
or OR4 (N23738, N23715, N22277, N3630, N22528);
not NOT1 (N23739, N23726);
xor XOR2 (N23740, N23729, N12280);
and AND4 (N23741, N23733, N13638, N4364, N7555);
not NOT1 (N23742, N23730);
xor XOR2 (N23743, N23740, N18603);
nor NOR2 (N23744, N23737, N14733);
nand NAND4 (N23745, N23743, N7794, N15056, N5822);
xor XOR2 (N23746, N23745, N12873);
buf BUF1 (N23747, N23735);
or OR3 (N23748, N23739, N20818, N13406);
nand NAND4 (N23749, N23722, N5561, N10133, N9341);
or OR2 (N23750, N23723, N9950);
not NOT1 (N23751, N23742);
not NOT1 (N23752, N23744);
not NOT1 (N23753, N23749);
not NOT1 (N23754, N23747);
and AND4 (N23755, N23753, N9652, N16900, N22377);
and AND4 (N23756, N23738, N12052, N10374, N11037);
buf BUF1 (N23757, N23748);
nand NAND2 (N23758, N23751, N23346);
buf BUF1 (N23759, N23757);
nand NAND2 (N23760, N23741, N16102);
or OR3 (N23761, N23754, N11643, N4823);
buf BUF1 (N23762, N23756);
buf BUF1 (N23763, N23758);
and AND3 (N23764, N23763, N1405, N21721);
or OR3 (N23765, N23755, N4321, N6132);
xor XOR2 (N23766, N23759, N21455);
nand NAND3 (N23767, N23714, N9567, N11625);
or OR2 (N23768, N23761, N15323);
and AND3 (N23769, N23766, N12895, N22135);
nor NOR2 (N23770, N23769, N22466);
xor XOR2 (N23771, N23765, N15642);
nor NOR3 (N23772, N23762, N15137, N5433);
and AND2 (N23773, N23752, N6179);
buf BUF1 (N23774, N23767);
and AND2 (N23775, N23773, N20480);
and AND3 (N23776, N23774, N9861, N13945);
nand NAND4 (N23777, N23776, N1411, N5270, N17156);
and AND2 (N23778, N23771, N22695);
and AND4 (N23779, N23768, N14187, N14193, N12672);
and AND3 (N23780, N23778, N22383, N16317);
not NOT1 (N23781, N23779);
buf BUF1 (N23782, N23746);
nand NAND2 (N23783, N23770, N8595);
nor NOR4 (N23784, N23750, N1026, N7721, N8040);
xor XOR2 (N23785, N23775, N18739);
xor XOR2 (N23786, N23781, N20685);
buf BUF1 (N23787, N23783);
xor XOR2 (N23788, N23786, N22294);
xor XOR2 (N23789, N23780, N10473);
and AND4 (N23790, N23782, N11944, N13861, N9487);
not NOT1 (N23791, N23789);
nor NOR2 (N23792, N23784, N10275);
buf BUF1 (N23793, N23772);
not NOT1 (N23794, N23760);
buf BUF1 (N23795, N23792);
or OR2 (N23796, N23764, N4519);
and AND4 (N23797, N23796, N12755, N1175, N12163);
nor NOR2 (N23798, N23788, N3170);
and AND2 (N23799, N23777, N12974);
nand NAND3 (N23800, N23790, N5673, N4559);
nor NOR2 (N23801, N23799, N5870);
and AND3 (N23802, N23794, N4522, N22563);
xor XOR2 (N23803, N23793, N23605);
nand NAND3 (N23804, N23797, N14203, N4095);
nand NAND2 (N23805, N23791, N21532);
nand NAND2 (N23806, N23802, N13562);
buf BUF1 (N23807, N23785);
not NOT1 (N23808, N23787);
nand NAND2 (N23809, N23800, N9224);
buf BUF1 (N23810, N23805);
xor XOR2 (N23811, N23803, N21827);
buf BUF1 (N23812, N23809);
nor NOR4 (N23813, N23806, N9836, N10322, N4605);
buf BUF1 (N23814, N23801);
nor NOR3 (N23815, N23810, N417, N18323);
xor XOR2 (N23816, N23815, N22495);
xor XOR2 (N23817, N23811, N12536);
not NOT1 (N23818, N23804);
xor XOR2 (N23819, N23817, N7540);
buf BUF1 (N23820, N23819);
nand NAND2 (N23821, N23795, N22987);
nor NOR2 (N23822, N23808, N2914);
and AND3 (N23823, N23798, N15632, N16433);
nand NAND2 (N23824, N23823, N17525);
not NOT1 (N23825, N23813);
buf BUF1 (N23826, N23820);
xor XOR2 (N23827, N23807, N2113);
nor NOR3 (N23828, N23824, N13119, N21060);
nor NOR2 (N23829, N23812, N23424);
or OR4 (N23830, N23822, N20866, N13455, N7028);
nor NOR4 (N23831, N23814, N2647, N2333, N13090);
and AND2 (N23832, N23828, N16611);
or OR3 (N23833, N23831, N1292, N12022);
and AND4 (N23834, N23827, N7908, N11451, N2335);
not NOT1 (N23835, N23818);
buf BUF1 (N23836, N23826);
nor NOR2 (N23837, N23830, N843);
nand NAND4 (N23838, N23834, N3, N13934, N8772);
or OR4 (N23839, N23833, N13659, N23436, N21235);
not NOT1 (N23840, N23825);
buf BUF1 (N23841, N23821);
buf BUF1 (N23842, N23832);
buf BUF1 (N23843, N23829);
nor NOR2 (N23844, N23842, N9827);
nand NAND2 (N23845, N23839, N3913);
buf BUF1 (N23846, N23838);
and AND4 (N23847, N23846, N9485, N13510, N14087);
and AND2 (N23848, N23843, N5995);
nor NOR3 (N23849, N23835, N18970, N187);
nand NAND4 (N23850, N23840, N14763, N18477, N9327);
or OR3 (N23851, N23847, N17482, N19545);
nand NAND4 (N23852, N23844, N6081, N7482, N13980);
not NOT1 (N23853, N23850);
xor XOR2 (N23854, N23848, N22147);
or OR4 (N23855, N23852, N5374, N15426, N18449);
xor XOR2 (N23856, N23837, N22276);
not NOT1 (N23857, N23853);
and AND3 (N23858, N23836, N23273, N11717);
not NOT1 (N23859, N23858);
buf BUF1 (N23860, N23851);
or OR4 (N23861, N23854, N20203, N4071, N6059);
and AND3 (N23862, N23849, N504, N4165);
not NOT1 (N23863, N23855);
and AND4 (N23864, N23861, N22018, N1568, N6973);
not NOT1 (N23865, N23860);
and AND2 (N23866, N23816, N6960);
buf BUF1 (N23867, N23841);
not NOT1 (N23868, N23862);
nand NAND3 (N23869, N23864, N2159, N9393);
nor NOR4 (N23870, N23863, N5802, N21777, N21989);
or OR3 (N23871, N23867, N12180, N13787);
nand NAND2 (N23872, N23868, N16721);
nor NOR3 (N23873, N23856, N18934, N22266);
buf BUF1 (N23874, N23871);
nor NOR4 (N23875, N23873, N15475, N17619, N17766);
or OR2 (N23876, N23874, N860);
nor NOR2 (N23877, N23875, N6747);
not NOT1 (N23878, N23869);
xor XOR2 (N23879, N23877, N21739);
nor NOR3 (N23880, N23857, N11960, N2799);
or OR2 (N23881, N23865, N4017);
and AND4 (N23882, N23878, N1378, N21794, N8969);
buf BUF1 (N23883, N23870);
not NOT1 (N23884, N23883);
or OR4 (N23885, N23884, N19933, N431, N23600);
xor XOR2 (N23886, N23872, N3440);
nor NOR4 (N23887, N23866, N18190, N19990, N19114);
nor NOR3 (N23888, N23885, N3116, N6756);
nand NAND4 (N23889, N23845, N14352, N7391, N1138);
buf BUF1 (N23890, N23879);
and AND4 (N23891, N23880, N23827, N19536, N7259);
buf BUF1 (N23892, N23890);
buf BUF1 (N23893, N23889);
and AND4 (N23894, N23893, N11532, N22935, N2166);
and AND2 (N23895, N23888, N397);
or OR4 (N23896, N23891, N11511, N15581, N20128);
nand NAND3 (N23897, N23887, N19168, N17964);
buf BUF1 (N23898, N23876);
buf BUF1 (N23899, N23896);
and AND2 (N23900, N23897, N13079);
and AND2 (N23901, N23886, N19304);
nor NOR4 (N23902, N23898, N10476, N16500, N2010);
buf BUF1 (N23903, N23894);
or OR2 (N23904, N23902, N18194);
buf BUF1 (N23905, N23904);
nor NOR4 (N23906, N23901, N21515, N19572, N10484);
not NOT1 (N23907, N23903);
and AND4 (N23908, N23882, N23192, N16937, N7725);
nand NAND2 (N23909, N23908, N17565);
nand NAND2 (N23910, N23899, N1614);
xor XOR2 (N23911, N23900, N19030);
not NOT1 (N23912, N23911);
and AND3 (N23913, N23905, N8128, N23663);
nand NAND4 (N23914, N23909, N12871, N23729, N3561);
or OR3 (N23915, N23859, N10535, N8331);
nand NAND3 (N23916, N23906, N21940, N17837);
nor NOR3 (N23917, N23913, N22767, N15025);
xor XOR2 (N23918, N23914, N21643);
not NOT1 (N23919, N23917);
nand NAND2 (N23920, N23915, N13671);
nor NOR3 (N23921, N23910, N9885, N20949);
xor XOR2 (N23922, N23916, N4075);
nor NOR4 (N23923, N23881, N9447, N3835, N11522);
nor NOR4 (N23924, N23892, N1658, N9256, N17104);
not NOT1 (N23925, N23919);
buf BUF1 (N23926, N23922);
buf BUF1 (N23927, N23912);
nand NAND2 (N23928, N23923, N3083);
nor NOR2 (N23929, N23907, N5342);
nor NOR4 (N23930, N23924, N2382, N14866, N16672);
nor NOR4 (N23931, N23927, N22187, N22498, N5273);
xor XOR2 (N23932, N23921, N4757);
or OR4 (N23933, N23930, N3250, N17021, N7836);
buf BUF1 (N23934, N23933);
not NOT1 (N23935, N23926);
xor XOR2 (N23936, N23932, N609);
xor XOR2 (N23937, N23936, N10653);
nand NAND2 (N23938, N23937, N7866);
or OR2 (N23939, N23935, N16765);
or OR3 (N23940, N23920, N3838, N19642);
xor XOR2 (N23941, N23938, N14751);
not NOT1 (N23942, N23928);
nor NOR2 (N23943, N23918, N14484);
not NOT1 (N23944, N23925);
or OR4 (N23945, N23941, N21531, N6946, N4256);
and AND3 (N23946, N23895, N12281, N22806);
not NOT1 (N23947, N23942);
xor XOR2 (N23948, N23946, N228);
buf BUF1 (N23949, N23948);
nor NOR4 (N23950, N23931, N7759, N4058, N5455);
nand NAND2 (N23951, N23939, N2350);
nor NOR3 (N23952, N23940, N2215, N838);
nand NAND2 (N23953, N23944, N10131);
nor NOR3 (N23954, N23951, N14315, N10545);
and AND3 (N23955, N23945, N9530, N2587);
xor XOR2 (N23956, N23952, N13545);
not NOT1 (N23957, N23950);
nand NAND4 (N23958, N23955, N211, N1749, N22778);
buf BUF1 (N23959, N23957);
or OR3 (N23960, N23954, N6148, N21154);
xor XOR2 (N23961, N23949, N2366);
xor XOR2 (N23962, N23953, N2143);
buf BUF1 (N23963, N23929);
nand NAND3 (N23964, N23960, N22804, N13872);
xor XOR2 (N23965, N23961, N5543);
or OR2 (N23966, N23959, N10374);
xor XOR2 (N23967, N23958, N19718);
nand NAND3 (N23968, N23947, N5637, N8039);
and AND2 (N23969, N23963, N14303);
and AND4 (N23970, N23956, N16995, N9421, N19842);
or OR4 (N23971, N23934, N19022, N4837, N9873);
nand NAND4 (N23972, N23969, N5111, N6735, N7243);
buf BUF1 (N23973, N23965);
buf BUF1 (N23974, N23967);
and AND4 (N23975, N23970, N3281, N11745, N14217);
xor XOR2 (N23976, N23966, N7424);
buf BUF1 (N23977, N23964);
and AND3 (N23978, N23971, N6104, N829);
and AND4 (N23979, N23962, N2714, N22212, N11347);
xor XOR2 (N23980, N23977, N15735);
xor XOR2 (N23981, N23978, N15150);
xor XOR2 (N23982, N23981, N21655);
not NOT1 (N23983, N23976);
nand NAND3 (N23984, N23943, N16884, N5531);
xor XOR2 (N23985, N23979, N17420);
or OR3 (N23986, N23974, N5079, N7317);
nand NAND2 (N23987, N23985, N20366);
nor NOR4 (N23988, N23987, N12753, N21132, N19331);
and AND3 (N23989, N23972, N3728, N18828);
and AND3 (N23990, N23973, N19452, N9558);
or OR2 (N23991, N23984, N8173);
buf BUF1 (N23992, N23989);
nand NAND3 (N23993, N23983, N7578, N19550);
not NOT1 (N23994, N23988);
not NOT1 (N23995, N23980);
not NOT1 (N23996, N23992);
or OR2 (N23997, N23968, N8213);
nor NOR2 (N23998, N23994, N15990);
buf BUF1 (N23999, N23991);
xor XOR2 (N24000, N23997, N16327);
buf BUF1 (N24001, N23996);
not NOT1 (N24002, N24001);
and AND2 (N24003, N23982, N23336);
and AND4 (N24004, N24003, N21956, N12010, N20844);
and AND3 (N24005, N23999, N4648, N21271);
nor NOR4 (N24006, N23990, N9171, N19625, N22551);
and AND2 (N24007, N24004, N11999);
not NOT1 (N24008, N24000);
and AND3 (N24009, N23995, N18654, N5612);
buf BUF1 (N24010, N23998);
or OR4 (N24011, N24002, N5147, N10899, N1071);
xor XOR2 (N24012, N24008, N6118);
buf BUF1 (N24013, N24012);
nor NOR4 (N24014, N23993, N19054, N12497, N16676);
or OR4 (N24015, N24013, N15315, N2667, N16339);
buf BUF1 (N24016, N23975);
not NOT1 (N24017, N24014);
nand NAND3 (N24018, N23986, N15936, N22694);
xor XOR2 (N24019, N24018, N22815);
xor XOR2 (N24020, N24019, N9559);
xor XOR2 (N24021, N24009, N11641);
buf BUF1 (N24022, N24020);
and AND4 (N24023, N24006, N10677, N23212, N22834);
buf BUF1 (N24024, N24007);
or OR3 (N24025, N24022, N2842, N23934);
nor NOR4 (N24026, N24010, N17116, N4142, N5417);
or OR2 (N24027, N24011, N5929);
nand NAND2 (N24028, N24024, N10356);
not NOT1 (N24029, N24005);
buf BUF1 (N24030, N24028);
xor XOR2 (N24031, N24021, N3932);
nand NAND4 (N24032, N24027, N17678, N21245, N13268);
and AND4 (N24033, N24029, N21918, N1796, N22333);
buf BUF1 (N24034, N24026);
nand NAND2 (N24035, N24034, N16857);
or OR4 (N24036, N24016, N24032, N17612, N19705);
and AND2 (N24037, N23781, N9364);
not NOT1 (N24038, N24023);
and AND3 (N24039, N24030, N3440, N15331);
not NOT1 (N24040, N24037);
and AND2 (N24041, N24031, N6749);
and AND3 (N24042, N24025, N3692, N21394);
nand NAND4 (N24043, N24040, N11892, N13004, N16611);
and AND3 (N24044, N24017, N3914, N23488);
xor XOR2 (N24045, N24044, N4129);
nand NAND3 (N24046, N24045, N8056, N1669);
nand NAND4 (N24047, N24039, N18271, N4032, N19975);
nand NAND2 (N24048, N24036, N21298);
nand NAND3 (N24049, N24046, N16979, N2848);
nand NAND2 (N24050, N24015, N21772);
or OR4 (N24051, N24050, N5447, N23744, N8623);
not NOT1 (N24052, N24035);
buf BUF1 (N24053, N24033);
nor NOR3 (N24054, N24043, N6134, N23707);
and AND3 (N24055, N24054, N16839, N5317);
buf BUF1 (N24056, N24055);
not NOT1 (N24057, N24047);
and AND2 (N24058, N24048, N7885);
and AND3 (N24059, N24042, N17812, N15331);
or OR2 (N24060, N24057, N13267);
xor XOR2 (N24061, N24049, N3425);
buf BUF1 (N24062, N24060);
buf BUF1 (N24063, N24058);
xor XOR2 (N24064, N24051, N3322);
nor NOR4 (N24065, N24056, N5621, N11414, N8783);
not NOT1 (N24066, N24065);
nor NOR4 (N24067, N24059, N1380, N22183, N6971);
or OR2 (N24068, N24061, N13675);
not NOT1 (N24069, N24063);
nor NOR4 (N24070, N24038, N23600, N3949, N2625);
nor NOR4 (N24071, N24052, N21414, N11550, N22910);
and AND4 (N24072, N24071, N254, N12887, N4781);
xor XOR2 (N24073, N24053, N19060);
nand NAND2 (N24074, N24062, N18076);
xor XOR2 (N24075, N24073, N21398);
or OR3 (N24076, N24067, N22019, N11296);
not NOT1 (N24077, N24076);
or OR2 (N24078, N24066, N21111);
and AND4 (N24079, N24068, N1924, N5988, N468);
nand NAND2 (N24080, N24064, N1123);
buf BUF1 (N24081, N24041);
or OR2 (N24082, N24078, N14303);
nand NAND3 (N24083, N24070, N1691, N19621);
and AND4 (N24084, N24074, N7360, N4439, N14590);
and AND2 (N24085, N24069, N446);
not NOT1 (N24086, N24079);
and AND4 (N24087, N24085, N18772, N6316, N23451);
xor XOR2 (N24088, N24084, N13469);
nand NAND3 (N24089, N24080, N1567, N7911);
buf BUF1 (N24090, N24072);
nand NAND3 (N24091, N24077, N15875, N12704);
nand NAND2 (N24092, N24082, N19763);
buf BUF1 (N24093, N24092);
buf BUF1 (N24094, N24083);
buf BUF1 (N24095, N24087);
not NOT1 (N24096, N24094);
and AND2 (N24097, N24096, N10375);
nand NAND2 (N24098, N24093, N14964);
or OR2 (N24099, N24089, N16113);
xor XOR2 (N24100, N24095, N17764);
and AND2 (N24101, N24099, N5383);
nand NAND2 (N24102, N24098, N7381);
or OR2 (N24103, N24091, N22817);
nand NAND4 (N24104, N24075, N16474, N7595, N1776);
not NOT1 (N24105, N24088);
and AND2 (N24106, N24101, N8088);
xor XOR2 (N24107, N24102, N1982);
and AND2 (N24108, N24105, N548);
or OR3 (N24109, N24106, N3684, N11509);
and AND2 (N24110, N24097, N12094);
not NOT1 (N24111, N24103);
xor XOR2 (N24112, N24111, N21900);
and AND2 (N24113, N24081, N15076);
xor XOR2 (N24114, N24100, N14807);
and AND3 (N24115, N24112, N6112, N4962);
not NOT1 (N24116, N24109);
xor XOR2 (N24117, N24108, N15209);
not NOT1 (N24118, N24090);
and AND4 (N24119, N24104, N13300, N7396, N14502);
buf BUF1 (N24120, N24107);
nand NAND2 (N24121, N24086, N6331);
nor NOR2 (N24122, N24120, N21460);
nand NAND3 (N24123, N24114, N5890, N8598);
and AND4 (N24124, N24121, N1101, N8222, N20309);
or OR3 (N24125, N24119, N21732, N18201);
not NOT1 (N24126, N24118);
nand NAND2 (N24127, N24115, N3667);
nor NOR3 (N24128, N24127, N5291, N12507);
or OR3 (N24129, N24122, N3271, N21152);
xor XOR2 (N24130, N24116, N6958);
buf BUF1 (N24131, N24130);
not NOT1 (N24132, N24131);
xor XOR2 (N24133, N24129, N16459);
nand NAND2 (N24134, N24117, N4182);
not NOT1 (N24135, N24110);
and AND4 (N24136, N24128, N1905, N11479, N23747);
nor NOR3 (N24137, N24135, N3405, N12409);
nand NAND3 (N24138, N24133, N22858, N17818);
buf BUF1 (N24139, N24136);
nor NOR4 (N24140, N24139, N10086, N4628, N5267);
xor XOR2 (N24141, N24138, N13863);
buf BUF1 (N24142, N24123);
not NOT1 (N24143, N24141);
nor NOR2 (N24144, N24134, N4005);
or OR2 (N24145, N24132, N23779);
and AND2 (N24146, N24113, N22416);
and AND4 (N24147, N24137, N21358, N23350, N8351);
and AND4 (N24148, N24126, N11846, N11495, N3405);
buf BUF1 (N24149, N24142);
buf BUF1 (N24150, N24149);
or OR4 (N24151, N24150, N4976, N2455, N10873);
xor XOR2 (N24152, N24148, N12418);
and AND3 (N24153, N24144, N21941, N3536);
xor XOR2 (N24154, N24124, N15508);
xor XOR2 (N24155, N24146, N21594);
nor NOR3 (N24156, N24155, N16330, N14139);
and AND4 (N24157, N24152, N20663, N20606, N3662);
nor NOR3 (N24158, N24153, N21347, N10555);
not NOT1 (N24159, N24154);
nor NOR2 (N24160, N24145, N17570);
buf BUF1 (N24161, N24125);
or OR3 (N24162, N24158, N13238, N14331);
or OR4 (N24163, N24157, N296, N20356, N14976);
buf BUF1 (N24164, N24162);
or OR2 (N24165, N24161, N23600);
not NOT1 (N24166, N24164);
xor XOR2 (N24167, N24156, N6036);
xor XOR2 (N24168, N24166, N8414);
buf BUF1 (N24169, N24167);
not NOT1 (N24170, N24168);
nor NOR3 (N24171, N24140, N19166, N6969);
or OR2 (N24172, N24169, N3967);
nand NAND3 (N24173, N24160, N79, N23830);
nand NAND3 (N24174, N24143, N22490, N5674);
nand NAND2 (N24175, N24170, N22824);
buf BUF1 (N24176, N24165);
and AND2 (N24177, N24147, N14924);
xor XOR2 (N24178, N24177, N11676);
nand NAND3 (N24179, N24163, N18419, N5851);
not NOT1 (N24180, N24171);
nor NOR4 (N24181, N24173, N8655, N5745, N17641);
nand NAND3 (N24182, N24159, N2905, N13453);
nor NOR2 (N24183, N24181, N19393);
or OR4 (N24184, N24180, N23383, N920, N22668);
xor XOR2 (N24185, N24151, N5913);
not NOT1 (N24186, N24175);
buf BUF1 (N24187, N24178);
not NOT1 (N24188, N24186);
not NOT1 (N24189, N24182);
xor XOR2 (N24190, N24172, N24041);
nor NOR2 (N24191, N24185, N3580);
not NOT1 (N24192, N24187);
nand NAND2 (N24193, N24191, N8118);
and AND2 (N24194, N24174, N18907);
nor NOR3 (N24195, N24188, N9734, N9026);
buf BUF1 (N24196, N24176);
nor NOR4 (N24197, N24194, N75, N482, N14226);
buf BUF1 (N24198, N24195);
not NOT1 (N24199, N24196);
nand NAND2 (N24200, N24198, N7143);
or OR4 (N24201, N24189, N12717, N16691, N12290);
xor XOR2 (N24202, N24183, N9356);
nor NOR4 (N24203, N24201, N852, N22706, N19403);
not NOT1 (N24204, N24193);
xor XOR2 (N24205, N24184, N17837);
and AND2 (N24206, N24204, N5);
nand NAND2 (N24207, N24197, N6190);
buf BUF1 (N24208, N24207);
and AND2 (N24209, N24190, N17393);
xor XOR2 (N24210, N24200, N20888);
nor NOR3 (N24211, N24205, N13842, N23310);
not NOT1 (N24212, N24208);
or OR4 (N24213, N24209, N3184, N15308, N12355);
or OR3 (N24214, N24192, N5187, N22759);
nor NOR2 (N24215, N24202, N6611);
or OR2 (N24216, N24213, N1974);
or OR4 (N24217, N24214, N20774, N8911, N17742);
or OR4 (N24218, N24216, N8532, N1583, N5126);
nand NAND4 (N24219, N24210, N20992, N4879, N5135);
or OR3 (N24220, N24203, N4419, N7445);
and AND4 (N24221, N24219, N7890, N19117, N22483);
or OR3 (N24222, N24218, N5716, N66);
xor XOR2 (N24223, N24217, N11085);
and AND3 (N24224, N24223, N11237, N12373);
or OR4 (N24225, N24220, N23437, N2973, N14267);
xor XOR2 (N24226, N24221, N22120);
or OR4 (N24227, N24212, N9140, N4974, N4230);
not NOT1 (N24228, N24215);
not NOT1 (N24229, N24199);
buf BUF1 (N24230, N24228);
and AND3 (N24231, N24179, N2441, N12512);
nand NAND4 (N24232, N24227, N13715, N23228, N11136);
not NOT1 (N24233, N24225);
and AND4 (N24234, N24224, N6262, N2686, N5302);
and AND2 (N24235, N24222, N23057);
nor NOR4 (N24236, N24234, N9817, N11240, N8544);
buf BUF1 (N24237, N24206);
nor NOR2 (N24238, N24211, N22566);
and AND2 (N24239, N24231, N4966);
or OR2 (N24240, N24229, N6496);
nand NAND2 (N24241, N24233, N1774);
nand NAND4 (N24242, N24236, N14395, N3574, N373);
xor XOR2 (N24243, N24242, N22950);
xor XOR2 (N24244, N24243, N11590);
buf BUF1 (N24245, N24232);
or OR2 (N24246, N24235, N18546);
nor NOR4 (N24247, N24240, N15679, N3574, N17056);
buf BUF1 (N24248, N24226);
and AND2 (N24249, N24241, N12645);
xor XOR2 (N24250, N24247, N5488);
xor XOR2 (N24251, N24239, N5501);
nand NAND4 (N24252, N24237, N12067, N195, N643);
and AND4 (N24253, N24248, N550, N16092, N3837);
not NOT1 (N24254, N24230);
buf BUF1 (N24255, N24250);
and AND2 (N24256, N24253, N12921);
buf BUF1 (N24257, N24249);
or OR4 (N24258, N24244, N985, N17822, N19244);
xor XOR2 (N24259, N24238, N19782);
and AND4 (N24260, N24257, N24018, N8316, N21616);
not NOT1 (N24261, N24251);
buf BUF1 (N24262, N24258);
and AND3 (N24263, N24261, N18096, N13414);
and AND3 (N24264, N24255, N12515, N17085);
and AND4 (N24265, N24246, N3572, N21875, N225);
nor NOR4 (N24266, N24260, N22567, N16431, N12936);
not NOT1 (N24267, N24254);
or OR4 (N24268, N24252, N9969, N17130, N6655);
nor NOR3 (N24269, N24259, N11894, N7834);
nand NAND3 (N24270, N24245, N3220, N11391);
not NOT1 (N24271, N24270);
xor XOR2 (N24272, N24269, N7054);
and AND3 (N24273, N24267, N6841, N19520);
not NOT1 (N24274, N24256);
or OR4 (N24275, N24262, N3887, N8897, N7568);
nand NAND2 (N24276, N24265, N12857);
nor NOR2 (N24277, N24271, N9550);
and AND2 (N24278, N24263, N3984);
and AND3 (N24279, N24274, N22739, N11171);
not NOT1 (N24280, N24272);
nor NOR3 (N24281, N24273, N10931, N11075);
or OR4 (N24282, N24275, N7864, N12510, N19393);
nor NOR4 (N24283, N24277, N20379, N913, N23439);
xor XOR2 (N24284, N24280, N21743);
not NOT1 (N24285, N24281);
buf BUF1 (N24286, N24283);
nand NAND2 (N24287, N24266, N9276);
nand NAND3 (N24288, N24278, N4423, N6742);
xor XOR2 (N24289, N24276, N1284);
buf BUF1 (N24290, N24264);
or OR3 (N24291, N24268, N12878, N12800);
and AND2 (N24292, N24290, N21031);
xor XOR2 (N24293, N24289, N513);
not NOT1 (N24294, N24284);
nand NAND2 (N24295, N24282, N19156);
nand NAND4 (N24296, N24293, N4278, N20173, N3534);
buf BUF1 (N24297, N24295);
buf BUF1 (N24298, N24286);
not NOT1 (N24299, N24285);
and AND3 (N24300, N24296, N11507, N10899);
or OR2 (N24301, N24291, N3603);
not NOT1 (N24302, N24299);
and AND4 (N24303, N24279, N21213, N1007, N17631);
nor NOR4 (N24304, N24300, N11494, N3760, N18241);
xor XOR2 (N24305, N24288, N21608);
xor XOR2 (N24306, N24303, N7854);
and AND4 (N24307, N24298, N16447, N11565, N6002);
or OR3 (N24308, N24292, N8646, N21723);
not NOT1 (N24309, N24304);
buf BUF1 (N24310, N24307);
nand NAND3 (N24311, N24306, N4562, N1466);
not NOT1 (N24312, N24301);
and AND3 (N24313, N24312, N19187, N21813);
not NOT1 (N24314, N24297);
and AND2 (N24315, N24305, N5385);
not NOT1 (N24316, N24302);
xor XOR2 (N24317, N24294, N3429);
nand NAND4 (N24318, N24310, N19024, N4082, N502);
or OR4 (N24319, N24315, N18920, N8320, N2123);
nor NOR2 (N24320, N24308, N6720);
nand NAND3 (N24321, N24311, N2309, N7934);
not NOT1 (N24322, N24318);
not NOT1 (N24323, N24316);
or OR4 (N24324, N24322, N1173, N21897, N21460);
and AND4 (N24325, N24287, N14857, N17345, N7886);
or OR4 (N24326, N24317, N2742, N22541, N285);
nand NAND4 (N24327, N24314, N15941, N1589, N4265);
or OR3 (N24328, N24325, N15851, N14143);
not NOT1 (N24329, N24327);
or OR2 (N24330, N24326, N14898);
nor NOR3 (N24331, N24324, N18348, N7511);
buf BUF1 (N24332, N24328);
not NOT1 (N24333, N24320);
or OR2 (N24334, N24331, N23568);
xor XOR2 (N24335, N24319, N24269);
nor NOR4 (N24336, N24321, N16210, N11990, N14605);
nor NOR4 (N24337, N24335, N20915, N18125, N20665);
and AND3 (N24338, N24334, N17604, N10738);
and AND3 (N24339, N24313, N11387, N23642);
or OR2 (N24340, N24337, N17329);
not NOT1 (N24341, N24336);
or OR2 (N24342, N24341, N19137);
buf BUF1 (N24343, N24338);
buf BUF1 (N24344, N24340);
and AND3 (N24345, N24342, N19630, N5715);
or OR4 (N24346, N24339, N17889, N2781, N19420);
buf BUF1 (N24347, N24309);
buf BUF1 (N24348, N24323);
xor XOR2 (N24349, N24330, N21459);
not NOT1 (N24350, N24348);
and AND4 (N24351, N24344, N8374, N6748, N23985);
and AND3 (N24352, N24332, N10562, N2515);
nor NOR4 (N24353, N24350, N5371, N22889, N17300);
and AND2 (N24354, N24347, N13738);
buf BUF1 (N24355, N24349);
nand NAND2 (N24356, N24345, N12498);
and AND2 (N24357, N24353, N2579);
nand NAND4 (N24358, N24329, N8509, N877, N9731);
buf BUF1 (N24359, N24333);
or OR3 (N24360, N24357, N7025, N23155);
buf BUF1 (N24361, N24354);
nand NAND3 (N24362, N24359, N9268, N2717);
nand NAND3 (N24363, N24361, N7317, N20509);
nor NOR4 (N24364, N24343, N11335, N17074, N15506);
or OR4 (N24365, N24356, N21261, N22779, N15406);
xor XOR2 (N24366, N24346, N7958);
buf BUF1 (N24367, N24365);
and AND2 (N24368, N24358, N12584);
xor XOR2 (N24369, N24366, N18429);
nand NAND3 (N24370, N24363, N24327, N11098);
nor NOR4 (N24371, N24360, N5689, N1471, N9339);
not NOT1 (N24372, N24351);
or OR2 (N24373, N24371, N12317);
not NOT1 (N24374, N24369);
nand NAND2 (N24375, N24367, N15772);
not NOT1 (N24376, N24362);
nor NOR2 (N24377, N24374, N305);
buf BUF1 (N24378, N24352);
not NOT1 (N24379, N24378);
nor NOR3 (N24380, N24368, N7239, N12962);
nor NOR4 (N24381, N24364, N11318, N3092, N19658);
not NOT1 (N24382, N24355);
or OR3 (N24383, N24381, N5719, N13563);
xor XOR2 (N24384, N24370, N7825);
not NOT1 (N24385, N24384);
buf BUF1 (N24386, N24375);
xor XOR2 (N24387, N24377, N10417);
buf BUF1 (N24388, N24373);
xor XOR2 (N24389, N24383, N24177);
not NOT1 (N24390, N24387);
nor NOR3 (N24391, N24382, N17717, N12666);
nand NAND2 (N24392, N24380, N18364);
not NOT1 (N24393, N24390);
nor NOR3 (N24394, N24376, N15192, N12526);
xor XOR2 (N24395, N24394, N21682);
xor XOR2 (N24396, N24395, N10876);
and AND2 (N24397, N24372, N21199);
not NOT1 (N24398, N24391);
xor XOR2 (N24399, N24389, N11343);
or OR3 (N24400, N24399, N20047, N23653);
buf BUF1 (N24401, N24379);
or OR4 (N24402, N24400, N9673, N18805, N13975);
and AND3 (N24403, N24393, N10622, N16776);
nand NAND3 (N24404, N24388, N6501, N3084);
buf BUF1 (N24405, N24402);
nor NOR3 (N24406, N24403, N7454, N6265);
buf BUF1 (N24407, N24385);
or OR4 (N24408, N24405, N7494, N8265, N19966);
buf BUF1 (N24409, N24407);
nand NAND3 (N24410, N24386, N14895, N3144);
and AND4 (N24411, N24406, N24174, N22824, N352);
nand NAND3 (N24412, N24404, N12542, N24195);
not NOT1 (N24413, N24410);
buf BUF1 (N24414, N24396);
nor NOR2 (N24415, N24411, N23489);
not NOT1 (N24416, N24414);
nand NAND4 (N24417, N24392, N15760, N9120, N2089);
buf BUF1 (N24418, N24408);
xor XOR2 (N24419, N24416, N3608);
and AND3 (N24420, N24397, N13616, N1954);
nand NAND4 (N24421, N24417, N21045, N20604, N13713);
and AND2 (N24422, N24421, N7843);
xor XOR2 (N24423, N24401, N14031);
buf BUF1 (N24424, N24415);
not NOT1 (N24425, N24419);
not NOT1 (N24426, N24413);
and AND3 (N24427, N24398, N2202, N9874);
nor NOR2 (N24428, N24420, N10359);
xor XOR2 (N24429, N24423, N22029);
and AND4 (N24430, N24429, N18911, N3560, N2143);
nor NOR4 (N24431, N24418, N21992, N9915, N5552);
nand NAND4 (N24432, N24426, N17273, N967, N16264);
nor NOR4 (N24433, N24430, N6697, N10753, N13255);
xor XOR2 (N24434, N24409, N6375);
xor XOR2 (N24435, N24432, N2207);
buf BUF1 (N24436, N24435);
nand NAND4 (N24437, N24428, N20131, N2428, N6194);
and AND2 (N24438, N24425, N8069);
nand NAND4 (N24439, N24431, N14484, N8279, N14374);
nand NAND3 (N24440, N24433, N22497, N24070);
nand NAND4 (N24441, N24412, N4197, N14337, N24209);
not NOT1 (N24442, N24424);
nand NAND4 (N24443, N24434, N4882, N6612, N22592);
nor NOR2 (N24444, N24443, N2172);
and AND2 (N24445, N24438, N9797);
xor XOR2 (N24446, N24441, N11979);
or OR2 (N24447, N24440, N13073);
and AND3 (N24448, N24427, N19876, N7924);
not NOT1 (N24449, N24437);
or OR3 (N24450, N24449, N17365, N4144);
nor NOR2 (N24451, N24450, N13070);
not NOT1 (N24452, N24448);
xor XOR2 (N24453, N24446, N14300);
not NOT1 (N24454, N24451);
or OR3 (N24455, N24454, N23596, N23581);
buf BUF1 (N24456, N24445);
or OR4 (N24457, N24436, N2796, N20950, N18811);
nand NAND4 (N24458, N24456, N1423, N1936, N21932);
not NOT1 (N24459, N24455);
or OR4 (N24460, N24442, N17210, N7057, N17438);
and AND2 (N24461, N24459, N13277);
nor NOR2 (N24462, N24460, N3157);
nor NOR3 (N24463, N24439, N20434, N4889);
nand NAND3 (N24464, N24422, N21036, N18712);
nand NAND3 (N24465, N24462, N20824, N7834);
or OR4 (N24466, N24458, N4667, N19967, N19583);
and AND4 (N24467, N24465, N3374, N19586, N5072);
nor NOR4 (N24468, N24452, N198, N18344, N19588);
nand NAND4 (N24469, N24453, N11443, N341, N12990);
not NOT1 (N24470, N24467);
nand NAND2 (N24471, N24470, N17477);
xor XOR2 (N24472, N24444, N17795);
buf BUF1 (N24473, N24471);
xor XOR2 (N24474, N24463, N15188);
nand NAND4 (N24475, N24464, N15838, N13169, N5851);
or OR2 (N24476, N24466, N20132);
nand NAND4 (N24477, N24447, N20776, N14366, N524);
or OR2 (N24478, N24476, N5010);
or OR4 (N24479, N24475, N22760, N8599, N13872);
nor NOR4 (N24480, N24477, N10996, N12464, N190);
nand NAND4 (N24481, N24479, N4684, N20366, N119);
or OR3 (N24482, N24474, N5176, N10562);
nor NOR4 (N24483, N24473, N5741, N10810, N17257);
not NOT1 (N24484, N24472);
nor NOR2 (N24485, N24478, N14124);
or OR2 (N24486, N24468, N501);
or OR4 (N24487, N24485, N7184, N12644, N7439);
nor NOR4 (N24488, N24457, N24426, N19692, N5959);
not NOT1 (N24489, N24486);
and AND4 (N24490, N24487, N5428, N16506, N9516);
or OR3 (N24491, N24480, N19714, N16949);
xor XOR2 (N24492, N24484, N21465);
nor NOR4 (N24493, N24490, N17751, N2007, N8222);
xor XOR2 (N24494, N24488, N21422);
buf BUF1 (N24495, N24489);
xor XOR2 (N24496, N24493, N1041);
nand NAND3 (N24497, N24495, N875, N14439);
xor XOR2 (N24498, N24481, N18247);
nor NOR4 (N24499, N24461, N22710, N7998, N19392);
buf BUF1 (N24500, N24491);
xor XOR2 (N24501, N24496, N17366);
not NOT1 (N24502, N24498);
or OR3 (N24503, N24492, N4969, N3644);
buf BUF1 (N24504, N24501);
nand NAND3 (N24505, N24482, N24423, N210);
not NOT1 (N24506, N24504);
buf BUF1 (N24507, N24505);
nor NOR3 (N24508, N24483, N10685, N17674);
and AND2 (N24509, N24497, N9520);
not NOT1 (N24510, N24509);
or OR3 (N24511, N24502, N19307, N20233);
nor NOR2 (N24512, N24503, N19207);
not NOT1 (N24513, N24510);
nor NOR2 (N24514, N24499, N314);
or OR3 (N24515, N24508, N7265, N1598);
nor NOR3 (N24516, N24513, N20880, N23710);
or OR4 (N24517, N24516, N214, N18797, N12011);
not NOT1 (N24518, N24514);
nand NAND4 (N24519, N24500, N20040, N8212, N12734);
not NOT1 (N24520, N24512);
not NOT1 (N24521, N24506);
not NOT1 (N24522, N24517);
and AND2 (N24523, N24520, N22499);
nor NOR2 (N24524, N24511, N12871);
not NOT1 (N24525, N24523);
xor XOR2 (N24526, N24522, N19645);
or OR3 (N24527, N24521, N20749, N4591);
nand NAND3 (N24528, N24524, N5618, N6627);
and AND2 (N24529, N24469, N5580);
xor XOR2 (N24530, N24529, N12691);
nor NOR4 (N24531, N24519, N4202, N17474, N11215);
not NOT1 (N24532, N24531);
and AND3 (N24533, N24527, N12871, N12261);
and AND4 (N24534, N24525, N15378, N10289, N11007);
or OR4 (N24535, N24507, N2024, N4654, N7122);
and AND3 (N24536, N24518, N11913, N8892);
nor NOR2 (N24537, N24532, N6958);
and AND4 (N24538, N24536, N11729, N5253, N18856);
nor NOR2 (N24539, N24526, N20670);
not NOT1 (N24540, N24535);
and AND3 (N24541, N24534, N4037, N11131);
not NOT1 (N24542, N24541);
nor NOR2 (N24543, N24530, N19692);
or OR2 (N24544, N24533, N21577);
and AND3 (N24545, N24542, N625, N6388);
nor NOR3 (N24546, N24540, N5136, N21906);
or OR2 (N24547, N24537, N8581);
nor NOR4 (N24548, N24515, N21947, N11405, N17277);
nand NAND4 (N24549, N24546, N13407, N17536, N21770);
not NOT1 (N24550, N24538);
xor XOR2 (N24551, N24543, N15026);
or OR4 (N24552, N24549, N16509, N2375, N5592);
and AND4 (N24553, N24545, N23467, N10605, N18387);
not NOT1 (N24554, N24539);
not NOT1 (N24555, N24553);
and AND2 (N24556, N24551, N7151);
nand NAND4 (N24557, N24556, N14768, N17676, N20213);
nor NOR2 (N24558, N24552, N12832);
nor NOR2 (N24559, N24494, N8292);
or OR4 (N24560, N24557, N17699, N5865, N15684);
and AND4 (N24561, N24560, N23207, N2062, N18018);
buf BUF1 (N24562, N24547);
and AND3 (N24563, N24562, N13405, N11524);
not NOT1 (N24564, N24554);
or OR4 (N24565, N24544, N11980, N6372, N7559);
nand NAND4 (N24566, N24563, N5101, N16988, N19465);
nand NAND3 (N24567, N24548, N290, N19290);
buf BUF1 (N24568, N24555);
buf BUF1 (N24569, N24550);
nand NAND4 (N24570, N24567, N19318, N21005, N2784);
or OR4 (N24571, N24566, N5877, N10146, N23719);
or OR4 (N24572, N24558, N8271, N1675, N3102);
nor NOR3 (N24573, N24561, N24185, N17018);
nor NOR2 (N24574, N24564, N19202);
buf BUF1 (N24575, N24528);
and AND3 (N24576, N24574, N22045, N24209);
not NOT1 (N24577, N24575);
nor NOR2 (N24578, N24568, N16044);
not NOT1 (N24579, N24576);
not NOT1 (N24580, N24571);
not NOT1 (N24581, N24570);
nand NAND2 (N24582, N24573, N3029);
nor NOR4 (N24583, N24565, N3675, N17704, N2993);
nor NOR2 (N24584, N24572, N18488);
nor NOR2 (N24585, N24569, N19650);
or OR4 (N24586, N24584, N17563, N18031, N16072);
nor NOR3 (N24587, N24579, N12669, N10566);
not NOT1 (N24588, N24577);
buf BUF1 (N24589, N24559);
nor NOR2 (N24590, N24580, N7373);
buf BUF1 (N24591, N24585);
or OR4 (N24592, N24591, N1189, N2576, N7812);
xor XOR2 (N24593, N24581, N9770);
xor XOR2 (N24594, N24583, N914);
buf BUF1 (N24595, N24588);
not NOT1 (N24596, N24586);
and AND2 (N24597, N24595, N23358);
buf BUF1 (N24598, N24590);
xor XOR2 (N24599, N24593, N12949);
and AND3 (N24600, N24599, N3438, N4835);
nand NAND4 (N24601, N24594, N6696, N3553, N14018);
buf BUF1 (N24602, N24587);
xor XOR2 (N24603, N24601, N785);
buf BUF1 (N24604, N24597);
not NOT1 (N24605, N24578);
and AND4 (N24606, N24596, N21237, N10284, N21904);
or OR4 (N24607, N24582, N14127, N12545, N19432);
buf BUF1 (N24608, N24600);
buf BUF1 (N24609, N24608);
or OR3 (N24610, N24606, N18919, N5985);
or OR3 (N24611, N24592, N14894, N9803);
xor XOR2 (N24612, N24589, N21933);
nand NAND2 (N24613, N24611, N23446);
nor NOR2 (N24614, N24612, N1325);
or OR3 (N24615, N24607, N3520, N16519);
and AND3 (N24616, N24602, N13928, N21233);
buf BUF1 (N24617, N24605);
not NOT1 (N24618, N24616);
and AND2 (N24619, N24617, N5236);
not NOT1 (N24620, N24615);
xor XOR2 (N24621, N24604, N19333);
and AND2 (N24622, N24619, N12790);
buf BUF1 (N24623, N24613);
nor NOR3 (N24624, N24618, N17340, N15070);
buf BUF1 (N24625, N24621);
xor XOR2 (N24626, N24622, N5968);
not NOT1 (N24627, N24609);
nor NOR3 (N24628, N24624, N13243, N8755);
or OR4 (N24629, N24627, N20604, N17343, N8668);
or OR3 (N24630, N24610, N9246, N12589);
xor XOR2 (N24631, N24623, N18714);
buf BUF1 (N24632, N24598);
buf BUF1 (N24633, N24603);
nor NOR2 (N24634, N24628, N7438);
not NOT1 (N24635, N24614);
nand NAND3 (N24636, N24620, N13503, N252);
and AND4 (N24637, N24636, N10238, N5178, N12066);
or OR4 (N24638, N24626, N9318, N23383, N7841);
xor XOR2 (N24639, N24637, N18085);
xor XOR2 (N24640, N24630, N13180);
buf BUF1 (N24641, N24631);
or OR2 (N24642, N24641, N11795);
nand NAND3 (N24643, N24638, N6164, N9102);
and AND3 (N24644, N24642, N21300, N4223);
nand NAND4 (N24645, N24640, N3901, N21014, N22126);
and AND3 (N24646, N24625, N20472, N1536);
buf BUF1 (N24647, N24645);
nand NAND2 (N24648, N24643, N13001);
and AND2 (N24649, N24635, N14535);
xor XOR2 (N24650, N24639, N13790);
or OR2 (N24651, N24647, N21551);
nand NAND4 (N24652, N24650, N15452, N11139, N821);
and AND4 (N24653, N24644, N17578, N14991, N11569);
and AND4 (N24654, N24629, N896, N14341, N20951);
buf BUF1 (N24655, N24646);
and AND3 (N24656, N24651, N16810, N8404);
not NOT1 (N24657, N24652);
nand NAND4 (N24658, N24655, N23331, N5539, N24489);
buf BUF1 (N24659, N24653);
or OR4 (N24660, N24649, N20925, N24190, N16869);
not NOT1 (N24661, N24656);
nand NAND2 (N24662, N24634, N16124);
buf BUF1 (N24663, N24662);
and AND3 (N24664, N24657, N16990, N19302);
nand NAND4 (N24665, N24658, N3867, N14866, N2233);
and AND2 (N24666, N24661, N11214);
nor NOR2 (N24667, N24633, N3678);
nand NAND4 (N24668, N24632, N17268, N9558, N8463);
not NOT1 (N24669, N24660);
buf BUF1 (N24670, N24654);
xor XOR2 (N24671, N24664, N4545);
and AND3 (N24672, N24671, N14394, N2315);
xor XOR2 (N24673, N24667, N21586);
or OR3 (N24674, N24648, N20932, N3819);
buf BUF1 (N24675, N24663);
not NOT1 (N24676, N24672);
buf BUF1 (N24677, N24675);
nand NAND2 (N24678, N24674, N1998);
nor NOR4 (N24679, N24666, N485, N15508, N3712);
and AND2 (N24680, N24679, N11796);
and AND4 (N24681, N24669, N10252, N2757, N2455);
nand NAND4 (N24682, N24678, N12250, N15556, N6488);
or OR3 (N24683, N24665, N835, N18161);
nand NAND3 (N24684, N24677, N6240, N16395);
or OR2 (N24685, N24659, N7987);
xor XOR2 (N24686, N24676, N8898);
or OR2 (N24687, N24682, N4808);
or OR4 (N24688, N24687, N23505, N4574, N22000);
or OR2 (N24689, N24681, N292);
or OR4 (N24690, N24685, N10306, N21137, N18992);
nand NAND4 (N24691, N24670, N24483, N21682, N14960);
nor NOR4 (N24692, N24673, N22655, N19717, N11669);
or OR3 (N24693, N24689, N22119, N15246);
or OR2 (N24694, N24668, N12590);
not NOT1 (N24695, N24690);
not NOT1 (N24696, N24686);
not NOT1 (N24697, N24693);
xor XOR2 (N24698, N24684, N506);
nor NOR2 (N24699, N24697, N17084);
nor NOR2 (N24700, N24696, N11305);
xor XOR2 (N24701, N24695, N13580);
and AND2 (N24702, N24691, N10765);
and AND3 (N24703, N24701, N4465, N8928);
nand NAND3 (N24704, N24700, N1825, N1873);
xor XOR2 (N24705, N24703, N9194);
buf BUF1 (N24706, N24705);
nand NAND4 (N24707, N24692, N12649, N17373, N15755);
xor XOR2 (N24708, N24683, N3300);
nand NAND3 (N24709, N24708, N19843, N23308);
nand NAND4 (N24710, N24707, N10752, N7475, N3447);
xor XOR2 (N24711, N24710, N8713);
nand NAND3 (N24712, N24704, N14789, N2626);
nor NOR4 (N24713, N24706, N9637, N11134, N5166);
and AND3 (N24714, N24680, N20956, N12372);
xor XOR2 (N24715, N24698, N23517);
nand NAND2 (N24716, N24694, N23179);
or OR2 (N24717, N24716, N1476);
not NOT1 (N24718, N24711);
nand NAND3 (N24719, N24699, N13219, N212);
nor NOR2 (N24720, N24709, N14472);
buf BUF1 (N24721, N24717);
nand NAND4 (N24722, N24688, N12857, N20388, N3288);
buf BUF1 (N24723, N24715);
not NOT1 (N24724, N24721);
nor NOR3 (N24725, N24714, N2366, N23994);
buf BUF1 (N24726, N24724);
not NOT1 (N24727, N24725);
not NOT1 (N24728, N24727);
not NOT1 (N24729, N24726);
buf BUF1 (N24730, N24702);
xor XOR2 (N24731, N24713, N11483);
and AND2 (N24732, N24722, N17391);
nand NAND4 (N24733, N24712, N4155, N7826, N16478);
nor NOR4 (N24734, N24729, N4721, N2223, N17854);
not NOT1 (N24735, N24728);
and AND4 (N24736, N24731, N14812, N23708, N16096);
nor NOR4 (N24737, N24720, N24695, N1311, N2430);
or OR2 (N24738, N24719, N7370);
nor NOR4 (N24739, N24737, N11983, N11300, N19730);
nor NOR2 (N24740, N24739, N1511);
not NOT1 (N24741, N24736);
or OR3 (N24742, N24740, N13330, N2335);
nor NOR2 (N24743, N24735, N9870);
nor NOR4 (N24744, N24732, N3773, N14431, N7583);
buf BUF1 (N24745, N24742);
not NOT1 (N24746, N24744);
or OR3 (N24747, N24743, N14660, N9585);
nand NAND4 (N24748, N24723, N16645, N10861, N13628);
not NOT1 (N24749, N24730);
and AND4 (N24750, N24733, N3696, N1091, N1853);
and AND3 (N24751, N24745, N10844, N4806);
and AND2 (N24752, N24749, N19162);
and AND4 (N24753, N24718, N17342, N15315, N13890);
nor NOR2 (N24754, N24748, N4197);
and AND4 (N24755, N24753, N11243, N17018, N14095);
xor XOR2 (N24756, N24750, N5420);
xor XOR2 (N24757, N24747, N4388);
not NOT1 (N24758, N24755);
nand NAND3 (N24759, N24741, N13773, N19614);
not NOT1 (N24760, N24734);
nand NAND2 (N24761, N24751, N166);
buf BUF1 (N24762, N24738);
buf BUF1 (N24763, N24762);
nand NAND4 (N24764, N24758, N11219, N20084, N24231);
and AND3 (N24765, N24761, N21531, N15718);
or OR4 (N24766, N24763, N5345, N12253, N12221);
xor XOR2 (N24767, N24760, N17159);
xor XOR2 (N24768, N24752, N11802);
xor XOR2 (N24769, N24765, N23385);
nor NOR3 (N24770, N24756, N8097, N17351);
nand NAND3 (N24771, N24767, N16258, N1577);
xor XOR2 (N24772, N24746, N23955);
xor XOR2 (N24773, N24754, N2376);
nor NOR4 (N24774, N24773, N18258, N18462, N16487);
not NOT1 (N24775, N24757);
buf BUF1 (N24776, N24759);
nand NAND4 (N24777, N24776, N3674, N7262, N23544);
or OR4 (N24778, N24764, N1018, N19321, N17763);
xor XOR2 (N24779, N24769, N16188);
buf BUF1 (N24780, N24778);
nor NOR3 (N24781, N24772, N5875, N21665);
or OR2 (N24782, N24771, N16719);
not NOT1 (N24783, N24766);
nand NAND3 (N24784, N24781, N15559, N7412);
and AND4 (N24785, N24780, N11455, N17531, N10482);
nand NAND4 (N24786, N24777, N19784, N4322, N8350);
nor NOR4 (N24787, N24783, N2067, N10624, N19877);
buf BUF1 (N24788, N24775);
buf BUF1 (N24789, N24785);
xor XOR2 (N24790, N24779, N20222);
not NOT1 (N24791, N24774);
nand NAND4 (N24792, N24770, N6340, N10827, N24412);
and AND3 (N24793, N24782, N1045, N6616);
nand NAND2 (N24794, N24787, N14911);
xor XOR2 (N24795, N24794, N9192);
not NOT1 (N24796, N24768);
nand NAND4 (N24797, N24788, N7553, N6270, N6109);
and AND2 (N24798, N24796, N943);
xor XOR2 (N24799, N24792, N2976);
or OR2 (N24800, N24793, N11943);
and AND2 (N24801, N24797, N13817);
and AND4 (N24802, N24798, N13248, N19375, N17172);
nand NAND3 (N24803, N24801, N19464, N16542);
or OR2 (N24804, N24784, N17486);
buf BUF1 (N24805, N24804);
nand NAND4 (N24806, N24789, N13549, N4305, N849);
nor NOR4 (N24807, N24791, N21597, N8430, N12003);
nand NAND4 (N24808, N24802, N13506, N13791, N20319);
not NOT1 (N24809, N24805);
and AND2 (N24810, N24808, N21592);
nor NOR3 (N24811, N24795, N5326, N18143);
nand NAND2 (N24812, N24807, N18288);
buf BUF1 (N24813, N24786);
xor XOR2 (N24814, N24803, N11839);
nand NAND3 (N24815, N24814, N12373, N8667);
and AND3 (N24816, N24812, N13925, N2883);
buf BUF1 (N24817, N24800);
not NOT1 (N24818, N24813);
or OR3 (N24819, N24809, N15391, N12049);
not NOT1 (N24820, N24816);
xor XOR2 (N24821, N24818, N18737);
nand NAND2 (N24822, N24821, N15993);
nand NAND4 (N24823, N24799, N12737, N14663, N8614);
xor XOR2 (N24824, N24823, N13353);
not NOT1 (N24825, N24790);
or OR2 (N24826, N24824, N8020);
nor NOR4 (N24827, N24819, N14247, N8224, N415);
or OR3 (N24828, N24825, N12104, N9651);
xor XOR2 (N24829, N24828, N23279);
nand NAND4 (N24830, N24811, N18776, N6582, N9259);
and AND3 (N24831, N24822, N23800, N14652);
nand NAND3 (N24832, N24831, N23870, N4195);
or OR4 (N24833, N24815, N4692, N15491, N20917);
not NOT1 (N24834, N24817);
xor XOR2 (N24835, N24829, N15905);
or OR2 (N24836, N24833, N17824);
xor XOR2 (N24837, N24830, N9956);
buf BUF1 (N24838, N24806);
not NOT1 (N24839, N24836);
xor XOR2 (N24840, N24820, N14778);
buf BUF1 (N24841, N24835);
xor XOR2 (N24842, N24827, N24080);
xor XOR2 (N24843, N24839, N12541);
buf BUF1 (N24844, N24826);
buf BUF1 (N24845, N24838);
not NOT1 (N24846, N24810);
or OR3 (N24847, N24846, N17676, N8727);
or OR4 (N24848, N24832, N5640, N4361, N6150);
nand NAND2 (N24849, N24841, N4708);
nand NAND3 (N24850, N24842, N3310, N8319);
buf BUF1 (N24851, N24849);
not NOT1 (N24852, N24840);
nor NOR3 (N24853, N24834, N819, N19126);
buf BUF1 (N24854, N24843);
and AND4 (N24855, N24845, N21326, N24121, N4685);
not NOT1 (N24856, N24852);
xor XOR2 (N24857, N24848, N16493);
xor XOR2 (N24858, N24847, N1424);
not NOT1 (N24859, N24858);
nor NOR4 (N24860, N24859, N1977, N1905, N22514);
xor XOR2 (N24861, N24844, N22418);
or OR2 (N24862, N24837, N9786);
xor XOR2 (N24863, N24850, N6338);
buf BUF1 (N24864, N24857);
and AND4 (N24865, N24853, N18157, N4679, N8548);
and AND4 (N24866, N24862, N23463, N16145, N17028);
nor NOR2 (N24867, N24860, N19677);
nand NAND3 (N24868, N24861, N22247, N24637);
xor XOR2 (N24869, N24864, N13291);
nor NOR4 (N24870, N24866, N5110, N19899, N14558);
or OR2 (N24871, N24854, N12060);
xor XOR2 (N24872, N24855, N17443);
or OR2 (N24873, N24870, N14682);
nor NOR4 (N24874, N24872, N8743, N23647, N4056);
and AND2 (N24875, N24873, N14688);
xor XOR2 (N24876, N24856, N17075);
xor XOR2 (N24877, N24865, N6274);
nor NOR3 (N24878, N24874, N8084, N11478);
nand NAND3 (N24879, N24869, N5694, N16321);
and AND4 (N24880, N24851, N19856, N15304, N18062);
nand NAND3 (N24881, N24876, N7061, N18782);
not NOT1 (N24882, N24878);
nand NAND2 (N24883, N24881, N22448);
and AND2 (N24884, N24871, N8612);
and AND4 (N24885, N24883, N17748, N3935, N11804);
nor NOR3 (N24886, N24879, N2669, N24654);
nand NAND3 (N24887, N24868, N18223, N17424);
nor NOR4 (N24888, N24863, N4178, N1286, N24379);
buf BUF1 (N24889, N24886);
not NOT1 (N24890, N24885);
and AND3 (N24891, N24882, N15920, N3628);
and AND2 (N24892, N24887, N4495);
xor XOR2 (N24893, N24877, N24205);
or OR4 (N24894, N24893, N3717, N13350, N5506);
xor XOR2 (N24895, N24891, N12129);
nor NOR3 (N24896, N24894, N20975, N17824);
and AND3 (N24897, N24875, N20151, N6535);
buf BUF1 (N24898, N24890);
buf BUF1 (N24899, N24892);
and AND3 (N24900, N24889, N12371, N17710);
nand NAND4 (N24901, N24884, N13507, N15984, N22182);
nor NOR3 (N24902, N24895, N8437, N9468);
xor XOR2 (N24903, N24880, N2079);
and AND2 (N24904, N24903, N18615);
nor NOR4 (N24905, N24900, N24275, N12165, N12173);
and AND3 (N24906, N24896, N24685, N12456);
nand NAND3 (N24907, N24905, N16707, N23321);
and AND4 (N24908, N24888, N12060, N15930, N8663);
and AND2 (N24909, N24908, N18009);
buf BUF1 (N24910, N24901);
or OR3 (N24911, N24910, N22763, N16892);
xor XOR2 (N24912, N24906, N16931);
nor NOR2 (N24913, N24902, N1973);
not NOT1 (N24914, N24899);
not NOT1 (N24915, N24911);
buf BUF1 (N24916, N24867);
buf BUF1 (N24917, N24909);
nor NOR4 (N24918, N24915, N18560, N2570, N23145);
nor NOR2 (N24919, N24916, N2923);
nor NOR2 (N24920, N24913, N6504);
buf BUF1 (N24921, N24898);
nand NAND2 (N24922, N24920, N12723);
nand NAND2 (N24923, N24907, N11352);
xor XOR2 (N24924, N24923, N15480);
and AND4 (N24925, N24914, N17171, N14173, N4631);
nor NOR3 (N24926, N24919, N8477, N8839);
nor NOR4 (N24927, N24912, N4467, N15964, N23509);
not NOT1 (N24928, N24927);
not NOT1 (N24929, N24922);
buf BUF1 (N24930, N24921);
nand NAND3 (N24931, N24926, N20746, N18942);
nand NAND2 (N24932, N24917, N19891);
nor NOR4 (N24933, N24924, N13412, N20091, N21309);
nand NAND2 (N24934, N24930, N15227);
nor NOR4 (N24935, N24931, N16241, N24742, N3630);
and AND4 (N24936, N24925, N19930, N21406, N12083);
nand NAND4 (N24937, N24935, N20845, N12031, N20523);
xor XOR2 (N24938, N24929, N12958);
xor XOR2 (N24939, N24928, N12988);
and AND3 (N24940, N24932, N9966, N11833);
buf BUF1 (N24941, N24936);
or OR2 (N24942, N24934, N14032);
nand NAND4 (N24943, N24940, N14730, N274, N9273);
not NOT1 (N24944, N24941);
nor NOR2 (N24945, N24944, N7698);
or OR4 (N24946, N24904, N13951, N18118, N11989);
and AND2 (N24947, N24897, N5847);
or OR2 (N24948, N24918, N5867);
or OR4 (N24949, N24946, N19715, N693, N18702);
xor XOR2 (N24950, N24949, N14514);
xor XOR2 (N24951, N24938, N18583);
nor NOR3 (N24952, N24948, N11956, N17209);
nor NOR2 (N24953, N24952, N4773);
nand NAND4 (N24954, N24953, N7633, N2006, N24458);
not NOT1 (N24955, N24947);
nand NAND3 (N24956, N24942, N6598, N3452);
nand NAND2 (N24957, N24933, N15260);
and AND4 (N24958, N24939, N12636, N21588, N9597);
or OR3 (N24959, N24954, N19802, N3194);
not NOT1 (N24960, N24943);
xor XOR2 (N24961, N24955, N3181);
buf BUF1 (N24962, N24960);
nor NOR2 (N24963, N24958, N10188);
or OR3 (N24964, N24962, N11037, N13182);
xor XOR2 (N24965, N24964, N15197);
or OR4 (N24966, N24961, N164, N13968, N15434);
nor NOR4 (N24967, N24945, N8974, N8583, N21776);
and AND2 (N24968, N24966, N4943);
and AND4 (N24969, N24937, N10731, N14347, N22004);
or OR3 (N24970, N24967, N14826, N2830);
nor NOR4 (N24971, N24963, N345, N9222, N7569);
buf BUF1 (N24972, N24950);
and AND3 (N24973, N24968, N5437, N21904);
nand NAND3 (N24974, N24969, N353, N17718);
or OR4 (N24975, N24959, N15283, N15580, N13639);
or OR2 (N24976, N24965, N11060);
and AND2 (N24977, N24971, N4752);
nor NOR3 (N24978, N24977, N3351, N23484);
or OR3 (N24979, N24956, N19112, N13986);
not NOT1 (N24980, N24978);
not NOT1 (N24981, N24980);
nor NOR4 (N24982, N24975, N19070, N7467, N15982);
or OR4 (N24983, N24951, N925, N19871, N20276);
nand NAND4 (N24984, N24957, N9218, N18245, N24914);
nor NOR4 (N24985, N24981, N18571, N19306, N14514);
or OR2 (N24986, N24982, N12270);
nor NOR2 (N24987, N24986, N796);
xor XOR2 (N24988, N24972, N221);
and AND2 (N24989, N24983, N24086);
xor XOR2 (N24990, N24974, N12240);
xor XOR2 (N24991, N24976, N1874);
or OR2 (N24992, N24991, N10553);
or OR3 (N24993, N24973, N14454, N7791);
or OR3 (N24994, N24984, N11794, N4123);
or OR2 (N24995, N24994, N15843);
nor NOR4 (N24996, N24970, N8414, N14827, N16701);
and AND4 (N24997, N24990, N9171, N19070, N16879);
and AND4 (N24998, N24993, N234, N13381, N24017);
xor XOR2 (N24999, N24992, N1720);
or OR4 (N25000, N24995, N1904, N11501, N1515);
buf BUF1 (N25001, N24999);
not NOT1 (N25002, N24997);
nor NOR3 (N25003, N24987, N20132, N6897);
or OR4 (N25004, N24998, N1188, N20876, N18457);
and AND3 (N25005, N25001, N5292, N16803);
nor NOR2 (N25006, N24979, N1425);
or OR3 (N25007, N24988, N6610, N16083);
nor NOR4 (N25008, N25006, N8317, N17162, N20129);
and AND3 (N25009, N24996, N19787, N14920);
or OR4 (N25010, N25000, N23381, N6332, N5271);
not NOT1 (N25011, N25004);
xor XOR2 (N25012, N25003, N6944);
nand NAND4 (N25013, N25002, N14464, N3995, N6049);
nand NAND2 (N25014, N25005, N10279);
or OR3 (N25015, N25014, N461, N22684);
not NOT1 (N25016, N25015);
or OR2 (N25017, N25008, N8245);
and AND4 (N25018, N25012, N8297, N22451, N17093);
and AND2 (N25019, N25011, N17804);
or OR2 (N25020, N25017, N17962);
or OR2 (N25021, N25019, N9034);
nor NOR4 (N25022, N25009, N14725, N14362, N24791);
xor XOR2 (N25023, N25007, N12795);
buf BUF1 (N25024, N24989);
nand NAND2 (N25025, N25018, N893);
nand NAND4 (N25026, N25021, N19151, N2313, N16982);
or OR3 (N25027, N24985, N12586, N23531);
xor XOR2 (N25028, N25026, N9930);
and AND4 (N25029, N25024, N6974, N21403, N11494);
not NOT1 (N25030, N25013);
and AND2 (N25031, N25022, N21106);
nor NOR4 (N25032, N25025, N14684, N24975, N17738);
nand NAND3 (N25033, N25030, N24798, N19288);
and AND2 (N25034, N25029, N6353);
xor XOR2 (N25035, N25031, N7704);
nor NOR4 (N25036, N25035, N9650, N14348, N21362);
buf BUF1 (N25037, N25032);
buf BUF1 (N25038, N25016);
not NOT1 (N25039, N25038);
buf BUF1 (N25040, N25039);
and AND3 (N25041, N25028, N12760, N3729);
buf BUF1 (N25042, N25033);
nor NOR4 (N25043, N25040, N21201, N342, N18819);
nor NOR2 (N25044, N25034, N18095);
buf BUF1 (N25045, N25037);
or OR3 (N25046, N25042, N6585, N8028);
nand NAND4 (N25047, N25045, N18736, N21270, N20787);
buf BUF1 (N25048, N25043);
xor XOR2 (N25049, N25010, N13772);
nand NAND3 (N25050, N25027, N18437, N12130);
xor XOR2 (N25051, N25023, N19568);
or OR2 (N25052, N25049, N15609);
not NOT1 (N25053, N25048);
buf BUF1 (N25054, N25020);
buf BUF1 (N25055, N25046);
and AND2 (N25056, N25044, N5120);
and AND3 (N25057, N25052, N16015, N22784);
nand NAND4 (N25058, N25047, N9908, N7904, N23204);
and AND4 (N25059, N25050, N16724, N22838, N6148);
nor NOR2 (N25060, N25054, N14536);
nor NOR2 (N25061, N25055, N19577);
buf BUF1 (N25062, N25053);
nor NOR4 (N25063, N25051, N13546, N19472, N12517);
buf BUF1 (N25064, N25058);
or OR4 (N25065, N25061, N15440, N17873, N12597);
and AND4 (N25066, N25041, N15808, N16212, N17860);
or OR4 (N25067, N25060, N23629, N11714, N13168);
buf BUF1 (N25068, N25059);
nand NAND2 (N25069, N25062, N10431);
nor NOR4 (N25070, N25066, N13172, N24996, N677);
xor XOR2 (N25071, N25063, N11985);
nor NOR4 (N25072, N25036, N1, N13033, N12774);
nand NAND3 (N25073, N25057, N21928, N17949);
or OR4 (N25074, N25073, N16063, N16493, N14847);
and AND4 (N25075, N25072, N13500, N4359, N3868);
nand NAND4 (N25076, N25069, N8416, N15902, N14543);
nand NAND3 (N25077, N25064, N18222, N6842);
buf BUF1 (N25078, N25070);
not NOT1 (N25079, N25075);
xor XOR2 (N25080, N25077, N12101);
nand NAND4 (N25081, N25074, N170, N16233, N23622);
and AND3 (N25082, N25067, N22062, N19746);
nor NOR3 (N25083, N25081, N19396, N11228);
buf BUF1 (N25084, N25078);
and AND2 (N25085, N25082, N2320);
or OR2 (N25086, N25068, N791);
nand NAND2 (N25087, N25071, N611);
or OR3 (N25088, N25086, N23199, N4910);
nand NAND3 (N25089, N25056, N21781, N477);
buf BUF1 (N25090, N25080);
nor NOR2 (N25091, N25076, N24748);
nand NAND2 (N25092, N25065, N5766);
or OR3 (N25093, N25091, N6280, N16305);
xor XOR2 (N25094, N25083, N14628);
nand NAND4 (N25095, N25093, N18141, N6076, N5206);
nand NAND4 (N25096, N25084, N13834, N16805, N18291);
or OR3 (N25097, N25088, N1903, N17719);
not NOT1 (N25098, N25087);
buf BUF1 (N25099, N25097);
and AND2 (N25100, N25098, N24882);
xor XOR2 (N25101, N25099, N1261);
and AND4 (N25102, N25079, N15995, N8980, N17577);
xor XOR2 (N25103, N25101, N22711);
nor NOR4 (N25104, N25085, N12659, N11324, N19135);
not NOT1 (N25105, N25103);
nor NOR4 (N25106, N25094, N1867, N11833, N2481);
nor NOR4 (N25107, N25102, N20548, N19270, N15530);
xor XOR2 (N25108, N25104, N19925);
and AND4 (N25109, N25100, N8285, N24871, N20741);
nand NAND3 (N25110, N25108, N20757, N4880);
nor NOR2 (N25111, N25105, N22190);
nand NAND2 (N25112, N25089, N10645);
and AND4 (N25113, N25111, N16918, N2988, N1899);
not NOT1 (N25114, N25090);
xor XOR2 (N25115, N25092, N13858);
xor XOR2 (N25116, N25106, N1355);
buf BUF1 (N25117, N25116);
and AND4 (N25118, N25113, N18998, N15143, N21688);
and AND4 (N25119, N25114, N17738, N13507, N16530);
nor NOR4 (N25120, N25119, N3617, N19155, N18547);
buf BUF1 (N25121, N25107);
nor NOR2 (N25122, N25096, N12769);
not NOT1 (N25123, N25118);
nor NOR3 (N25124, N25110, N11937, N14787);
nand NAND2 (N25125, N25115, N822);
xor XOR2 (N25126, N25112, N4839);
or OR4 (N25127, N25123, N19086, N23834, N14170);
nor NOR4 (N25128, N25109, N4081, N21436, N14944);
nand NAND4 (N25129, N25125, N9851, N16383, N20547);
xor XOR2 (N25130, N25124, N7265);
xor XOR2 (N25131, N25128, N6759);
and AND2 (N25132, N25127, N13625);
not NOT1 (N25133, N25126);
xor XOR2 (N25134, N25129, N23365);
xor XOR2 (N25135, N25130, N15659);
xor XOR2 (N25136, N25131, N13695);
not NOT1 (N25137, N25121);
nor NOR2 (N25138, N25134, N13744);
not NOT1 (N25139, N25117);
and AND4 (N25140, N25132, N15038, N9853, N1303);
or OR4 (N25141, N25120, N7979, N2827, N18781);
nor NOR2 (N25142, N25122, N14896);
xor XOR2 (N25143, N25139, N8304);
nand NAND4 (N25144, N25142, N3533, N13907, N1230);
nand NAND2 (N25145, N25135, N18193);
not NOT1 (N25146, N25143);
or OR2 (N25147, N25144, N24877);
not NOT1 (N25148, N25136);
xor XOR2 (N25149, N25147, N24643);
not NOT1 (N25150, N25149);
xor XOR2 (N25151, N25146, N23923);
not NOT1 (N25152, N25148);
nor NOR2 (N25153, N25133, N9982);
not NOT1 (N25154, N25153);
nand NAND2 (N25155, N25154, N21960);
xor XOR2 (N25156, N25145, N20687);
nor NOR4 (N25157, N25138, N10344, N9240, N7172);
xor XOR2 (N25158, N25150, N20143);
or OR2 (N25159, N25155, N20451);
nor NOR2 (N25160, N25140, N20994);
or OR2 (N25161, N25151, N6736);
not NOT1 (N25162, N25159);
nor NOR4 (N25163, N25162, N18538, N20481, N3711);
not NOT1 (N25164, N25163);
not NOT1 (N25165, N25137);
buf BUF1 (N25166, N25141);
buf BUF1 (N25167, N25161);
not NOT1 (N25168, N25167);
nand NAND2 (N25169, N25158, N21865);
buf BUF1 (N25170, N25157);
nand NAND3 (N25171, N25156, N3086, N22137);
and AND2 (N25172, N25152, N1547);
and AND4 (N25173, N25165, N14662, N14058, N2573);
not NOT1 (N25174, N25095);
and AND4 (N25175, N25166, N12, N7232, N16019);
or OR2 (N25176, N25174, N8430);
or OR3 (N25177, N25171, N19423, N628);
nor NOR3 (N25178, N25170, N11115, N22394);
nor NOR4 (N25179, N25176, N5979, N23368, N12536);
xor XOR2 (N25180, N25177, N14162);
not NOT1 (N25181, N25172);
buf BUF1 (N25182, N25168);
not NOT1 (N25183, N25178);
not NOT1 (N25184, N25182);
xor XOR2 (N25185, N25179, N12727);
and AND3 (N25186, N25185, N15451, N9626);
not NOT1 (N25187, N25175);
nor NOR3 (N25188, N25187, N1410, N10305);
buf BUF1 (N25189, N25181);
nand NAND3 (N25190, N25160, N4303, N22129);
not NOT1 (N25191, N25189);
xor XOR2 (N25192, N25183, N5560);
xor XOR2 (N25193, N25164, N20282);
and AND3 (N25194, N25192, N19995, N20302);
xor XOR2 (N25195, N25194, N4914);
buf BUF1 (N25196, N25184);
nand NAND4 (N25197, N25188, N17349, N1787, N10517);
or OR2 (N25198, N25180, N8781);
nand NAND4 (N25199, N25198, N11778, N12238, N20611);
buf BUF1 (N25200, N25173);
or OR4 (N25201, N25191, N11898, N10783, N21674);
buf BUF1 (N25202, N25186);
not NOT1 (N25203, N25197);
nor NOR4 (N25204, N25202, N6256, N24730, N16662);
xor XOR2 (N25205, N25201, N5434);
buf BUF1 (N25206, N25169);
and AND4 (N25207, N25200, N19315, N14543, N13998);
buf BUF1 (N25208, N25199);
nand NAND3 (N25209, N25205, N20417, N20449);
xor XOR2 (N25210, N25209, N3415);
or OR3 (N25211, N25210, N1324, N1214);
nand NAND4 (N25212, N25190, N6042, N18690, N22426);
buf BUF1 (N25213, N25211);
or OR3 (N25214, N25207, N18443, N2342);
xor XOR2 (N25215, N25208, N14145);
buf BUF1 (N25216, N25193);
or OR2 (N25217, N25203, N22245);
buf BUF1 (N25218, N25196);
and AND2 (N25219, N25195, N4585);
nor NOR4 (N25220, N25219, N12546, N24423, N23099);
nand NAND2 (N25221, N25206, N19033);
nand NAND3 (N25222, N25221, N24540, N13018);
or OR2 (N25223, N25204, N5277);
buf BUF1 (N25224, N25223);
nor NOR2 (N25225, N25224, N4268);
or OR2 (N25226, N25212, N2900);
nor NOR3 (N25227, N25225, N22608, N16010);
buf BUF1 (N25228, N25218);
or OR3 (N25229, N25213, N1166, N10160);
or OR4 (N25230, N25217, N1470, N6405, N21493);
or OR4 (N25231, N25222, N19779, N51, N12730);
nor NOR2 (N25232, N25228, N8746);
nand NAND3 (N25233, N25214, N8916, N21072);
and AND3 (N25234, N25226, N11866, N8870);
and AND2 (N25235, N25230, N8628);
or OR4 (N25236, N25220, N21966, N8353, N23459);
buf BUF1 (N25237, N25233);
nand NAND2 (N25238, N25227, N13858);
and AND4 (N25239, N25216, N21349, N7444, N24115);
nor NOR3 (N25240, N25239, N3283, N17645);
nand NAND2 (N25241, N25240, N4908);
buf BUF1 (N25242, N25236);
not NOT1 (N25243, N25234);
nand NAND2 (N25244, N25241, N8534);
not NOT1 (N25245, N25229);
and AND4 (N25246, N25235, N14064, N7838, N4861);
nor NOR4 (N25247, N25243, N4130, N21166, N3413);
nand NAND4 (N25248, N25244, N3055, N9089, N12982);
nor NOR4 (N25249, N25232, N17901, N13216, N22141);
xor XOR2 (N25250, N25238, N9688);
or OR2 (N25251, N25242, N5234);
or OR3 (N25252, N25245, N16443, N2508);
and AND3 (N25253, N25237, N2001, N3427);
not NOT1 (N25254, N25252);
nand NAND3 (N25255, N25251, N20297, N15749);
not NOT1 (N25256, N25250);
or OR4 (N25257, N25246, N17008, N9055, N4778);
nor NOR4 (N25258, N25248, N1573, N22361, N12241);
xor XOR2 (N25259, N25247, N18658);
xor XOR2 (N25260, N25256, N21730);
nand NAND3 (N25261, N25259, N15854, N9299);
xor XOR2 (N25262, N25231, N24310);
or OR2 (N25263, N25260, N12154);
buf BUF1 (N25264, N25257);
xor XOR2 (N25265, N25215, N15178);
nand NAND2 (N25266, N25262, N14549);
nor NOR2 (N25267, N25254, N9017);
or OR4 (N25268, N25264, N4309, N6589, N15815);
or OR2 (N25269, N25255, N22396);
and AND3 (N25270, N25269, N19971, N7232);
or OR3 (N25271, N25267, N4801, N1245);
xor XOR2 (N25272, N25270, N8395);
buf BUF1 (N25273, N25272);
not NOT1 (N25274, N25258);
nor NOR4 (N25275, N25253, N15029, N1675, N22372);
not NOT1 (N25276, N25261);
not NOT1 (N25277, N25276);
nand NAND2 (N25278, N25273, N15608);
xor XOR2 (N25279, N25274, N23168);
and AND2 (N25280, N25266, N22073);
not NOT1 (N25281, N25279);
and AND4 (N25282, N25275, N16934, N19054, N19177);
xor XOR2 (N25283, N25268, N22328);
not NOT1 (N25284, N25263);
or OR3 (N25285, N25277, N4559, N365);
nand NAND2 (N25286, N25278, N4938);
xor XOR2 (N25287, N25286, N21878);
and AND4 (N25288, N25285, N2514, N18523, N5692);
nand NAND4 (N25289, N25280, N22811, N18330, N6554);
or OR3 (N25290, N25287, N16183, N18223);
nand NAND4 (N25291, N25265, N1865, N1899, N24653);
not NOT1 (N25292, N25289);
xor XOR2 (N25293, N25249, N14332);
and AND2 (N25294, N25283, N14638);
not NOT1 (N25295, N25271);
not NOT1 (N25296, N25291);
nand NAND3 (N25297, N25281, N1942, N22115);
and AND3 (N25298, N25292, N9369, N13258);
buf BUF1 (N25299, N25284);
buf BUF1 (N25300, N25297);
or OR4 (N25301, N25299, N18070, N15626, N21251);
nand NAND4 (N25302, N25282, N22258, N16343, N8122);
and AND2 (N25303, N25288, N5027);
nor NOR2 (N25304, N25301, N2897);
buf BUF1 (N25305, N25304);
buf BUF1 (N25306, N25300);
not NOT1 (N25307, N25306);
xor XOR2 (N25308, N25294, N24609);
nand NAND2 (N25309, N25293, N20773);
xor XOR2 (N25310, N25308, N13601);
and AND3 (N25311, N25298, N6415, N15461);
nor NOR4 (N25312, N25296, N5519, N14807, N2286);
not NOT1 (N25313, N25290);
buf BUF1 (N25314, N25313);
xor XOR2 (N25315, N25309, N24739);
xor XOR2 (N25316, N25303, N16768);
xor XOR2 (N25317, N25316, N1246);
not NOT1 (N25318, N25315);
not NOT1 (N25319, N25295);
nor NOR2 (N25320, N25302, N25006);
buf BUF1 (N25321, N25317);
xor XOR2 (N25322, N25321, N4446);
xor XOR2 (N25323, N25319, N5036);
not NOT1 (N25324, N25312);
buf BUF1 (N25325, N25314);
xor XOR2 (N25326, N25318, N3598);
nor NOR2 (N25327, N25311, N22094);
and AND4 (N25328, N25327, N5424, N9941, N7910);
buf BUF1 (N25329, N25323);
buf BUF1 (N25330, N25328);
and AND2 (N25331, N25330, N14236);
buf BUF1 (N25332, N25329);
not NOT1 (N25333, N25325);
and AND3 (N25334, N25322, N17200, N24625);
buf BUF1 (N25335, N25324);
buf BUF1 (N25336, N25310);
buf BUF1 (N25337, N25333);
not NOT1 (N25338, N25335);
nand NAND3 (N25339, N25331, N13199, N6545);
or OR4 (N25340, N25307, N5454, N9197, N23041);
nand NAND4 (N25341, N25338, N18171, N10452, N20494);
nand NAND4 (N25342, N25340, N24041, N14459, N12332);
nand NAND2 (N25343, N25332, N9939);
and AND3 (N25344, N25326, N4840, N4661);
buf BUF1 (N25345, N25343);
not NOT1 (N25346, N25339);
and AND2 (N25347, N25337, N7744);
not NOT1 (N25348, N25341);
nand NAND2 (N25349, N25346, N17910);
nand NAND3 (N25350, N25305, N12695, N24387);
xor XOR2 (N25351, N25347, N23094);
and AND3 (N25352, N25345, N21239, N12707);
and AND4 (N25353, N25348, N25112, N8142, N20319);
nor NOR4 (N25354, N25334, N17313, N3044, N18816);
xor XOR2 (N25355, N25354, N23594);
and AND3 (N25356, N25336, N9352, N3025);
or OR3 (N25357, N25320, N21743, N20502);
and AND3 (N25358, N25349, N16904, N18731);
nand NAND4 (N25359, N25357, N9920, N21968, N20197);
and AND4 (N25360, N25344, N21474, N7232, N6149);
buf BUF1 (N25361, N25356);
and AND3 (N25362, N25360, N23636, N8876);
nor NOR2 (N25363, N25352, N10921);
xor XOR2 (N25364, N25361, N15644);
nor NOR3 (N25365, N25355, N12648, N356);
xor XOR2 (N25366, N25350, N18269);
buf BUF1 (N25367, N25362);
or OR4 (N25368, N25359, N21099, N9828, N15184);
nor NOR3 (N25369, N25358, N10308, N4570);
buf BUF1 (N25370, N25365);
and AND3 (N25371, N25367, N427, N11762);
and AND4 (N25372, N25369, N15062, N11635, N18491);
nand NAND4 (N25373, N25372, N5199, N12362, N14579);
or OR3 (N25374, N25368, N20485, N12755);
and AND4 (N25375, N25363, N17401, N10801, N9150);
nand NAND4 (N25376, N25375, N12651, N20278, N13450);
buf BUF1 (N25377, N25353);
or OR3 (N25378, N25373, N2700, N9427);
buf BUF1 (N25379, N25374);
buf BUF1 (N25380, N25342);
or OR2 (N25381, N25370, N91);
not NOT1 (N25382, N25371);
xor XOR2 (N25383, N25376, N15422);
nor NOR3 (N25384, N25351, N8533, N8126);
nand NAND2 (N25385, N25380, N25117);
nor NOR2 (N25386, N25383, N18482);
buf BUF1 (N25387, N25366);
xor XOR2 (N25388, N25384, N13569);
xor XOR2 (N25389, N25388, N3991);
or OR4 (N25390, N25386, N21083, N20947, N17472);
buf BUF1 (N25391, N25382);
and AND2 (N25392, N25381, N21547);
not NOT1 (N25393, N25391);
nand NAND2 (N25394, N25392, N3737);
not NOT1 (N25395, N25377);
nor NOR4 (N25396, N25394, N13107, N8794, N17338);
and AND2 (N25397, N25378, N2237);
not NOT1 (N25398, N25379);
not NOT1 (N25399, N25398);
nor NOR2 (N25400, N25364, N24777);
xor XOR2 (N25401, N25395, N6598);
buf BUF1 (N25402, N25399);
and AND4 (N25403, N25396, N7711, N19635, N21825);
or OR4 (N25404, N25385, N21523, N10918, N21006);
and AND2 (N25405, N25389, N2517);
nand NAND4 (N25406, N25387, N15317, N22899, N6025);
and AND3 (N25407, N25401, N6497, N9163);
buf BUF1 (N25408, N25397);
buf BUF1 (N25409, N25400);
xor XOR2 (N25410, N25409, N12926);
nand NAND3 (N25411, N25407, N12616, N198);
xor XOR2 (N25412, N25410, N22426);
and AND4 (N25413, N25406, N322, N17172, N8327);
xor XOR2 (N25414, N25408, N25009);
xor XOR2 (N25415, N25412, N20805);
not NOT1 (N25416, N25415);
or OR2 (N25417, N25414, N8394);
xor XOR2 (N25418, N25390, N8512);
or OR4 (N25419, N25393, N2255, N6600, N14722);
not NOT1 (N25420, N25403);
not NOT1 (N25421, N25417);
not NOT1 (N25422, N25402);
not NOT1 (N25423, N25422);
not NOT1 (N25424, N25419);
or OR2 (N25425, N25416, N1740);
or OR2 (N25426, N25404, N5292);
and AND2 (N25427, N25413, N6093);
not NOT1 (N25428, N25420);
and AND3 (N25429, N25427, N18081, N22316);
nand NAND3 (N25430, N25421, N23158, N3993);
or OR2 (N25431, N25428, N4087);
nand NAND3 (N25432, N25423, N16949, N11297);
xor XOR2 (N25433, N25418, N7697);
nor NOR4 (N25434, N25424, N19113, N8183, N14057);
xor XOR2 (N25435, N25432, N15612);
not NOT1 (N25436, N25433);
buf BUF1 (N25437, N25426);
and AND3 (N25438, N25405, N2997, N13843);
not NOT1 (N25439, N25430);
not NOT1 (N25440, N25438);
not NOT1 (N25441, N25411);
or OR2 (N25442, N25435, N23589);
xor XOR2 (N25443, N25437, N5990);
nand NAND2 (N25444, N25436, N10794);
or OR4 (N25445, N25425, N18281, N1497, N17284);
nor NOR2 (N25446, N25441, N25379);
nand NAND4 (N25447, N25444, N5044, N19981, N8797);
xor XOR2 (N25448, N25439, N2396);
xor XOR2 (N25449, N25447, N22597);
and AND3 (N25450, N25434, N16731, N15672);
nand NAND3 (N25451, N25450, N9560, N15460);
not NOT1 (N25452, N25446);
nand NAND3 (N25453, N25452, N5070, N20474);
nand NAND4 (N25454, N25431, N10694, N10604, N21722);
xor XOR2 (N25455, N25451, N2746);
or OR4 (N25456, N25448, N1179, N15964, N9077);
not NOT1 (N25457, N25449);
buf BUF1 (N25458, N25440);
nor NOR4 (N25459, N25458, N5799, N13244, N23008);
nor NOR4 (N25460, N25442, N7204, N22888, N4377);
nand NAND2 (N25461, N25443, N23251);
or OR2 (N25462, N25429, N19873);
xor XOR2 (N25463, N25454, N17609);
buf BUF1 (N25464, N25461);
not NOT1 (N25465, N25453);
nand NAND3 (N25466, N25462, N15414, N23903);
nand NAND2 (N25467, N25455, N191);
nand NAND3 (N25468, N25464, N12184, N78);
or OR3 (N25469, N25459, N17522, N5407);
nor NOR2 (N25470, N25468, N9760);
nor NOR4 (N25471, N25460, N7305, N19590, N8917);
or OR3 (N25472, N25456, N1816, N17199);
xor XOR2 (N25473, N25463, N18703);
xor XOR2 (N25474, N25465, N6777);
xor XOR2 (N25475, N25469, N21500);
nor NOR3 (N25476, N25445, N20026, N7686);
and AND4 (N25477, N25470, N16487, N8773, N13646);
nand NAND2 (N25478, N25475, N8284);
nor NOR4 (N25479, N25466, N9075, N22480, N25148);
xor XOR2 (N25480, N25472, N19311);
buf BUF1 (N25481, N25479);
nand NAND4 (N25482, N25476, N22869, N13019, N17166);
xor XOR2 (N25483, N25457, N25456);
xor XOR2 (N25484, N25482, N17551);
or OR3 (N25485, N25483, N8646, N25235);
and AND3 (N25486, N25474, N12381, N18170);
nor NOR4 (N25487, N25473, N24492, N19019, N11732);
not NOT1 (N25488, N25467);
nand NAND2 (N25489, N25487, N6960);
xor XOR2 (N25490, N25489, N16648);
xor XOR2 (N25491, N25488, N13296);
or OR2 (N25492, N25478, N23400);
buf BUF1 (N25493, N25485);
nor NOR2 (N25494, N25491, N14775);
or OR3 (N25495, N25480, N21460, N10979);
not NOT1 (N25496, N25486);
nand NAND2 (N25497, N25477, N22219);
xor XOR2 (N25498, N25496, N24008);
or OR3 (N25499, N25490, N22851, N18543);
nand NAND4 (N25500, N25495, N18198, N14159, N20842);
xor XOR2 (N25501, N25499, N16003);
or OR4 (N25502, N25494, N10134, N246, N19931);
or OR2 (N25503, N25492, N20207);
or OR3 (N25504, N25503, N12449, N15255);
nand NAND4 (N25505, N25484, N16763, N18536, N13022);
buf BUF1 (N25506, N25502);
nand NAND4 (N25507, N25506, N8728, N14217, N22805);
buf BUF1 (N25508, N25493);
buf BUF1 (N25509, N25508);
buf BUF1 (N25510, N25504);
buf BUF1 (N25511, N25498);
nor NOR3 (N25512, N25509, N22948, N13391);
nor NOR2 (N25513, N25507, N3781);
nor NOR3 (N25514, N25481, N19228, N2148);
nor NOR3 (N25515, N25505, N18428, N18067);
and AND3 (N25516, N25511, N12466, N21323);
nand NAND4 (N25517, N25500, N12528, N22197, N9980);
buf BUF1 (N25518, N25510);
nor NOR3 (N25519, N25513, N15083, N7074);
buf BUF1 (N25520, N25471);
nor NOR4 (N25521, N25501, N19006, N13609, N20454);
nor NOR3 (N25522, N25520, N3530, N8826);
or OR3 (N25523, N25517, N6227, N21558);
nand NAND2 (N25524, N25497, N451);
not NOT1 (N25525, N25522);
and AND4 (N25526, N25524, N10608, N721, N896);
nor NOR2 (N25527, N25518, N18168);
nor NOR2 (N25528, N25526, N11466);
xor XOR2 (N25529, N25521, N18232);
xor XOR2 (N25530, N25523, N1578);
nand NAND3 (N25531, N25525, N13045, N1126);
xor XOR2 (N25532, N25514, N4310);
nand NAND2 (N25533, N25531, N17020);
not NOT1 (N25534, N25512);
or OR4 (N25535, N25533, N11331, N10351, N13132);
not NOT1 (N25536, N25529);
nand NAND4 (N25537, N25515, N2478, N19978, N22180);
xor XOR2 (N25538, N25532, N19515);
nor NOR2 (N25539, N25538, N16532);
buf BUF1 (N25540, N25537);
nor NOR2 (N25541, N25534, N13371);
nor NOR3 (N25542, N25527, N5587, N6993);
nand NAND2 (N25543, N25535, N9048);
or OR2 (N25544, N25528, N21427);
xor XOR2 (N25545, N25530, N4577);
nor NOR3 (N25546, N25516, N16827, N22227);
nand NAND2 (N25547, N25546, N4449);
nand NAND3 (N25548, N25536, N535, N746);
not NOT1 (N25549, N25547);
not NOT1 (N25550, N25543);
xor XOR2 (N25551, N25519, N6169);
buf BUF1 (N25552, N25539);
not NOT1 (N25553, N25551);
not NOT1 (N25554, N25553);
and AND2 (N25555, N25542, N18011);
nor NOR2 (N25556, N25550, N21697);
or OR2 (N25557, N25549, N19850);
buf BUF1 (N25558, N25552);
nor NOR2 (N25559, N25554, N17554);
nand NAND4 (N25560, N25544, N6413, N23271, N25345);
or OR4 (N25561, N25540, N11178, N6247, N7177);
xor XOR2 (N25562, N25545, N10545);
and AND3 (N25563, N25562, N9842, N2442);
xor XOR2 (N25564, N25541, N746);
not NOT1 (N25565, N25555);
and AND2 (N25566, N25548, N5964);
nor NOR4 (N25567, N25557, N3076, N18176, N7933);
and AND4 (N25568, N25556, N24114, N8949, N18280);
or OR2 (N25569, N25568, N22676);
or OR3 (N25570, N25569, N25506, N10356);
or OR4 (N25571, N25564, N23369, N648, N22157);
buf BUF1 (N25572, N25567);
buf BUF1 (N25573, N25558);
or OR2 (N25574, N25572, N23361);
and AND4 (N25575, N25571, N14702, N4699, N6768);
xor XOR2 (N25576, N25575, N1954);
and AND3 (N25577, N25576, N24867, N14159);
buf BUF1 (N25578, N25566);
xor XOR2 (N25579, N25561, N14360);
buf BUF1 (N25580, N25565);
nor NOR2 (N25581, N25574, N5336);
nand NAND4 (N25582, N25559, N25157, N17653, N5589);
nor NOR3 (N25583, N25579, N17704, N5759);
and AND2 (N25584, N25573, N22179);
or OR2 (N25585, N25582, N20393);
nor NOR4 (N25586, N25577, N9204, N5286, N6245);
and AND4 (N25587, N25583, N14288, N14470, N21615);
and AND4 (N25588, N25580, N23601, N11848, N6152);
buf BUF1 (N25589, N25584);
nand NAND4 (N25590, N25588, N9869, N13385, N862);
not NOT1 (N25591, N25587);
or OR2 (N25592, N25591, N25039);
and AND4 (N25593, N25586, N907, N7352, N860);
xor XOR2 (N25594, N25570, N8647);
and AND4 (N25595, N25593, N423, N12271, N23017);
xor XOR2 (N25596, N25578, N16142);
and AND3 (N25597, N25590, N8535, N14355);
nand NAND4 (N25598, N25589, N8002, N19819, N12185);
not NOT1 (N25599, N25592);
not NOT1 (N25600, N25596);
or OR4 (N25601, N25563, N17456, N5077, N20971);
and AND3 (N25602, N25601, N1672, N13630);
or OR3 (N25603, N25594, N6986, N2759);
nor NOR3 (N25604, N25560, N7422, N6828);
and AND2 (N25605, N25598, N22622);
and AND2 (N25606, N25604, N3159);
or OR2 (N25607, N25605, N7913);
xor XOR2 (N25608, N25606, N10177);
nand NAND2 (N25609, N25595, N9161);
buf BUF1 (N25610, N25597);
xor XOR2 (N25611, N25599, N17306);
and AND3 (N25612, N25610, N21517, N23812);
and AND2 (N25613, N25581, N1115);
or OR2 (N25614, N25602, N25135);
buf BUF1 (N25615, N25607);
xor XOR2 (N25616, N25585, N3086);
not NOT1 (N25617, N25611);
xor XOR2 (N25618, N25612, N7913);
xor XOR2 (N25619, N25617, N127);
not NOT1 (N25620, N25603);
buf BUF1 (N25621, N25613);
nor NOR4 (N25622, N25608, N19162, N7681, N23374);
xor XOR2 (N25623, N25620, N19498);
not NOT1 (N25624, N25618);
endmodule