// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N2500,N2506,N2507,N2491,N2510,N2511,N2497,N2509,N2495,N2512;

not NOT1 (N13, N2);
not NOT1 (N14, N6);
nand NAND4 (N15, N10, N12, N9, N10);
nand NAND3 (N16, N5, N14, N2);
nor NOR4 (N17, N4, N1, N14, N4);
buf BUF1 (N18, N5);
not NOT1 (N19, N12);
or OR2 (N20, N17, N13);
xor XOR2 (N21, N14, N1);
nand NAND3 (N22, N13, N17, N19);
nand NAND4 (N23, N1, N12, N19, N19);
buf BUF1 (N24, N18);
or OR4 (N25, N22, N19, N7, N22);
buf BUF1 (N26, N25);
nor NOR3 (N27, N3, N6, N7);
not NOT1 (N28, N22);
not NOT1 (N29, N21);
xor XOR2 (N30, N26, N10);
and AND3 (N31, N11, N25, N14);
buf BUF1 (N32, N28);
and AND4 (N33, N27, N7, N25, N4);
or OR2 (N34, N24, N21);
nand NAND4 (N35, N23, N32, N28, N19);
nor NOR4 (N36, N18, N29, N11, N35);
or OR3 (N37, N12, N23, N31);
nand NAND4 (N38, N16, N9, N37, N33);
and AND4 (N39, N10, N23, N10, N24);
not NOT1 (N40, N15);
not NOT1 (N41, N13);
nand NAND3 (N42, N28, N8, N18);
not NOT1 (N43, N29);
nor NOR2 (N44, N20, N42);
or OR4 (N45, N19, N10, N44, N8);
and AND4 (N46, N5, N25, N22, N32);
not NOT1 (N47, N41);
nor NOR2 (N48, N36, N42);
buf BUF1 (N49, N34);
nor NOR3 (N50, N46, N37, N39);
nand NAND2 (N51, N9, N47);
or OR4 (N52, N51, N22, N8, N13);
xor XOR2 (N53, N42, N17);
or OR2 (N54, N45, N35);
nand NAND2 (N55, N52, N3);
xor XOR2 (N56, N54, N30);
nor NOR3 (N57, N7, N12, N38);
or OR3 (N58, N36, N24, N49);
nor NOR3 (N59, N50, N51, N46);
and AND4 (N60, N37, N30, N54, N20);
not NOT1 (N61, N58);
nand NAND3 (N62, N43, N27, N16);
nand NAND3 (N63, N48, N3, N5);
or OR2 (N64, N55, N30);
xor XOR2 (N65, N60, N43);
or OR2 (N66, N61, N48);
nand NAND3 (N67, N64, N4, N48);
and AND2 (N68, N65, N37);
xor XOR2 (N69, N59, N11);
not NOT1 (N70, N57);
xor XOR2 (N71, N63, N70);
xor XOR2 (N72, N71, N38);
and AND4 (N73, N7, N36, N27, N24);
and AND2 (N74, N53, N58);
nor NOR3 (N75, N66, N9, N56);
nand NAND2 (N76, N15, N38);
nand NAND3 (N77, N72, N30, N2);
and AND2 (N78, N40, N59);
buf BUF1 (N79, N68);
nand NAND4 (N80, N62, N30, N38, N20);
not NOT1 (N81, N76);
or OR4 (N82, N75, N22, N34, N70);
nor NOR3 (N83, N78, N29, N23);
and AND3 (N84, N69, N52, N30);
xor XOR2 (N85, N77, N24);
and AND3 (N86, N79, N28, N41);
nand NAND3 (N87, N84, N77, N35);
nor NOR2 (N88, N67, N78);
or OR3 (N89, N80, N82, N35);
xor XOR2 (N90, N77, N88);
buf BUF1 (N91, N40);
and AND2 (N92, N85, N5);
buf BUF1 (N93, N87);
nand NAND4 (N94, N90, N62, N87, N30);
xor XOR2 (N95, N91, N84);
buf BUF1 (N96, N74);
or OR2 (N97, N93, N74);
and AND3 (N98, N81, N42, N21);
or OR2 (N99, N83, N1);
or OR3 (N100, N95, N92, N31);
xor XOR2 (N101, N65, N23);
nand NAND3 (N102, N73, N59, N72);
nand NAND4 (N103, N99, N1, N73, N10);
buf BUF1 (N104, N97);
buf BUF1 (N105, N86);
buf BUF1 (N106, N104);
or OR2 (N107, N94, N96);
or OR2 (N108, N55, N38);
xor XOR2 (N109, N105, N26);
xor XOR2 (N110, N108, N32);
not NOT1 (N111, N100);
xor XOR2 (N112, N102, N71);
nand NAND3 (N113, N89, N79, N67);
or OR3 (N114, N98, N24, N14);
buf BUF1 (N115, N103);
not NOT1 (N116, N112);
or OR4 (N117, N107, N89, N48, N89);
buf BUF1 (N118, N109);
nor NOR3 (N119, N116, N69, N67);
buf BUF1 (N120, N113);
or OR2 (N121, N118, N41);
buf BUF1 (N122, N115);
buf BUF1 (N123, N117);
not NOT1 (N124, N119);
nor NOR4 (N125, N111, N18, N111, N104);
buf BUF1 (N126, N120);
nor NOR3 (N127, N106, N87, N68);
and AND3 (N128, N124, N109, N119);
buf BUF1 (N129, N121);
buf BUF1 (N130, N122);
nor NOR2 (N131, N123, N112);
nand NAND2 (N132, N101, N2);
buf BUF1 (N133, N128);
or OR4 (N134, N130, N60, N126, N125);
xor XOR2 (N135, N92, N63);
nor NOR2 (N136, N47, N8);
not NOT1 (N137, N114);
and AND3 (N138, N135, N80, N121);
buf BUF1 (N139, N133);
not NOT1 (N140, N110);
nand NAND4 (N141, N139, N69, N74, N23);
or OR3 (N142, N136, N3, N102);
and AND4 (N143, N137, N52, N141, N22);
nand NAND4 (N144, N133, N25, N107, N105);
or OR3 (N145, N127, N122, N101);
nand NAND4 (N146, N131, N59, N140, N88);
nor NOR3 (N147, N116, N119, N139);
buf BUF1 (N148, N134);
nor NOR4 (N149, N147, N89, N3, N126);
xor XOR2 (N150, N145, N72);
xor XOR2 (N151, N138, N17);
not NOT1 (N152, N148);
buf BUF1 (N153, N146);
xor XOR2 (N154, N142, N32);
or OR3 (N155, N129, N62, N147);
or OR2 (N156, N150, N6);
not NOT1 (N157, N153);
not NOT1 (N158, N156);
nand NAND3 (N159, N144, N17, N141);
buf BUF1 (N160, N155);
nand NAND4 (N161, N154, N91, N71, N38);
nor NOR2 (N162, N160, N72);
buf BUF1 (N163, N157);
or OR4 (N164, N161, N34, N157, N141);
and AND4 (N165, N162, N80, N57, N24);
or OR3 (N166, N151, N105, N89);
xor XOR2 (N167, N149, N133);
nand NAND4 (N168, N158, N149, N141, N18);
xor XOR2 (N169, N164, N35);
buf BUF1 (N170, N166);
nor NOR2 (N171, N143, N108);
nand NAND3 (N172, N167, N49, N167);
xor XOR2 (N173, N169, N119);
and AND3 (N174, N152, N88, N25);
or OR3 (N175, N173, N148, N96);
and AND2 (N176, N170, N121);
or OR3 (N177, N175, N43, N120);
not NOT1 (N178, N177);
nor NOR3 (N179, N174, N62, N32);
nand NAND2 (N180, N176, N132);
xor XOR2 (N181, N110, N152);
xor XOR2 (N182, N180, N89);
not NOT1 (N183, N171);
and AND4 (N184, N179, N99, N78, N1);
not NOT1 (N185, N159);
nand NAND3 (N186, N182, N54, N29);
or OR3 (N187, N178, N110, N33);
nor NOR4 (N188, N183, N21, N108, N62);
xor XOR2 (N189, N163, N114);
nand NAND4 (N190, N185, N40, N144, N41);
not NOT1 (N191, N165);
xor XOR2 (N192, N190, N174);
xor XOR2 (N193, N186, N123);
buf BUF1 (N194, N191);
not NOT1 (N195, N188);
or OR3 (N196, N172, N70, N57);
not NOT1 (N197, N195);
xor XOR2 (N198, N194, N67);
not NOT1 (N199, N198);
not NOT1 (N200, N168);
or OR4 (N201, N197, N136, N190, N186);
and AND3 (N202, N181, N141, N146);
or OR2 (N203, N202, N19);
not NOT1 (N204, N192);
or OR2 (N205, N189, N92);
xor XOR2 (N206, N204, N162);
not NOT1 (N207, N200);
nand NAND2 (N208, N196, N201);
xor XOR2 (N209, N34, N135);
nand NAND3 (N210, N205, N76, N174);
and AND3 (N211, N187, N88, N209);
not NOT1 (N212, N34);
or OR2 (N213, N212, N172);
and AND3 (N214, N206, N122, N51);
or OR4 (N215, N210, N14, N33, N206);
and AND3 (N216, N207, N37, N66);
nand NAND4 (N217, N193, N201, N44, N47);
not NOT1 (N218, N215);
or OR3 (N219, N203, N186, N14);
xor XOR2 (N220, N219, N218);
buf BUF1 (N221, N42);
and AND3 (N222, N211, N158, N120);
and AND4 (N223, N217, N137, N153, N18);
and AND3 (N224, N184, N222, N222);
not NOT1 (N225, N184);
not NOT1 (N226, N220);
nand NAND2 (N227, N221, N39);
xor XOR2 (N228, N225, N31);
nor NOR2 (N229, N228, N124);
nand NAND2 (N230, N223, N174);
buf BUF1 (N231, N227);
nor NOR3 (N232, N208, N222, N204);
buf BUF1 (N233, N216);
nand NAND4 (N234, N226, N100, N47, N108);
nand NAND3 (N235, N234, N228, N216);
buf BUF1 (N236, N230);
and AND4 (N237, N231, N169, N226, N22);
nand NAND4 (N238, N235, N166, N160, N128);
and AND2 (N239, N199, N206);
not NOT1 (N240, N237);
and AND2 (N241, N233, N144);
nand NAND4 (N242, N241, N165, N231, N191);
or OR4 (N243, N224, N64, N169, N11);
nand NAND4 (N244, N236, N98, N114, N228);
xor XOR2 (N245, N229, N117);
nor NOR4 (N246, N242, N203, N41, N98);
nor NOR3 (N247, N213, N167, N84);
xor XOR2 (N248, N214, N74);
and AND3 (N249, N232, N6, N32);
and AND4 (N250, N244, N184, N91, N120);
xor XOR2 (N251, N248, N137);
xor XOR2 (N252, N250, N69);
not NOT1 (N253, N251);
or OR2 (N254, N253, N93);
and AND3 (N255, N243, N5, N76);
xor XOR2 (N256, N254, N233);
buf BUF1 (N257, N252);
nor NOR2 (N258, N255, N99);
nand NAND4 (N259, N246, N253, N125, N5);
nor NOR3 (N260, N247, N247, N216);
and AND4 (N261, N249, N11, N260, N211);
nand NAND3 (N262, N219, N254, N219);
not NOT1 (N263, N240);
nand NAND4 (N264, N263, N166, N158, N89);
not NOT1 (N265, N257);
nor NOR2 (N266, N261, N73);
and AND3 (N267, N238, N48, N201);
nor NOR2 (N268, N267, N126);
not NOT1 (N269, N265);
xor XOR2 (N270, N264, N63);
xor XOR2 (N271, N259, N198);
buf BUF1 (N272, N268);
xor XOR2 (N273, N272, N59);
nand NAND2 (N274, N262, N16);
not NOT1 (N275, N256);
and AND2 (N276, N266, N5);
and AND4 (N277, N276, N75, N184, N71);
and AND3 (N278, N273, N40, N94);
not NOT1 (N279, N269);
xor XOR2 (N280, N274, N40);
and AND3 (N281, N239, N154, N134);
and AND4 (N282, N271, N41, N70, N50);
buf BUF1 (N283, N277);
xor XOR2 (N284, N282, N276);
xor XOR2 (N285, N283, N134);
and AND4 (N286, N279, N103, N202, N13);
or OR3 (N287, N258, N72, N211);
and AND3 (N288, N286, N146, N148);
xor XOR2 (N289, N275, N93);
nor NOR3 (N290, N280, N250, N36);
not NOT1 (N291, N284);
and AND2 (N292, N281, N291);
buf BUF1 (N293, N49);
nand NAND3 (N294, N292, N74, N37);
or OR2 (N295, N285, N231);
and AND2 (N296, N294, N95);
nand NAND4 (N297, N296, N4, N259, N65);
or OR4 (N298, N287, N185, N40, N191);
or OR2 (N299, N278, N184);
xor XOR2 (N300, N290, N26);
and AND3 (N301, N300, N145, N266);
not NOT1 (N302, N270);
not NOT1 (N303, N293);
or OR2 (N304, N302, N218);
buf BUF1 (N305, N245);
and AND2 (N306, N304, N166);
not NOT1 (N307, N298);
xor XOR2 (N308, N295, N278);
nand NAND4 (N309, N306, N71, N232, N114);
nand NAND4 (N310, N288, N268, N286, N285);
buf BUF1 (N311, N297);
not NOT1 (N312, N303);
nor NOR2 (N313, N311, N269);
nor NOR3 (N314, N305, N29, N268);
nor NOR4 (N315, N301, N63, N267, N213);
or OR3 (N316, N313, N19, N266);
and AND2 (N317, N307, N313);
buf BUF1 (N318, N317);
buf BUF1 (N319, N289);
buf BUF1 (N320, N310);
xor XOR2 (N321, N315, N15);
and AND4 (N322, N314, N20, N237, N311);
and AND4 (N323, N320, N63, N107, N270);
buf BUF1 (N324, N319);
and AND3 (N325, N309, N103, N169);
nor NOR3 (N326, N321, N246, N143);
nor NOR2 (N327, N316, N254);
nand NAND3 (N328, N327, N145, N317);
or OR4 (N329, N325, N137, N172, N114);
not NOT1 (N330, N308);
buf BUF1 (N331, N312);
or OR2 (N332, N330, N26);
or OR4 (N333, N318, N268, N91, N1);
and AND4 (N334, N299, N280, N250, N14);
not NOT1 (N335, N334);
or OR2 (N336, N322, N252);
xor XOR2 (N337, N333, N318);
not NOT1 (N338, N335);
nor NOR4 (N339, N337, N300, N198, N149);
xor XOR2 (N340, N339, N128);
nand NAND3 (N341, N324, N107, N13);
buf BUF1 (N342, N331);
nand NAND3 (N343, N341, N320, N184);
xor XOR2 (N344, N323, N323);
xor XOR2 (N345, N338, N194);
xor XOR2 (N346, N336, N85);
buf BUF1 (N347, N326);
nor NOR3 (N348, N347, N26, N92);
nand NAND2 (N349, N344, N305);
nand NAND2 (N350, N348, N280);
buf BUF1 (N351, N340);
nor NOR3 (N352, N343, N270, N247);
nor NOR3 (N353, N332, N103, N289);
xor XOR2 (N354, N349, N344);
or OR4 (N355, N329, N258, N343, N62);
and AND3 (N356, N353, N312, N333);
not NOT1 (N357, N342);
buf BUF1 (N358, N328);
and AND2 (N359, N346, N99);
or OR4 (N360, N359, N138, N12, N194);
and AND2 (N361, N358, N19);
buf BUF1 (N362, N345);
buf BUF1 (N363, N357);
buf BUF1 (N364, N355);
xor XOR2 (N365, N363, N42);
or OR2 (N366, N361, N126);
or OR3 (N367, N350, N135, N54);
or OR3 (N368, N351, N325, N283);
not NOT1 (N369, N364);
not NOT1 (N370, N367);
nor NOR3 (N371, N362, N234, N310);
and AND2 (N372, N369, N357);
xor XOR2 (N373, N360, N208);
and AND4 (N374, N366, N316, N125, N341);
xor XOR2 (N375, N370, N12);
and AND3 (N376, N368, N40, N337);
buf BUF1 (N377, N352);
and AND3 (N378, N372, N19, N46);
not NOT1 (N379, N374);
or OR2 (N380, N375, N362);
or OR3 (N381, N379, N116, N161);
buf BUF1 (N382, N376);
nor NOR3 (N383, N377, N372, N84);
xor XOR2 (N384, N381, N222);
xor XOR2 (N385, N378, N218);
or OR4 (N386, N380, N351, N123, N240);
xor XOR2 (N387, N385, N300);
nor NOR4 (N388, N356, N220, N295, N295);
nand NAND4 (N389, N386, N16, N331, N294);
xor XOR2 (N390, N383, N237);
buf BUF1 (N391, N387);
xor XOR2 (N392, N382, N191);
or OR2 (N393, N371, N306);
buf BUF1 (N394, N354);
buf BUF1 (N395, N365);
buf BUF1 (N396, N373);
buf BUF1 (N397, N384);
and AND3 (N398, N390, N68, N25);
buf BUF1 (N399, N392);
nand NAND2 (N400, N398, N138);
nand NAND4 (N401, N397, N373, N100, N370);
nor NOR2 (N402, N395, N30);
xor XOR2 (N403, N389, N372);
xor XOR2 (N404, N388, N106);
nand NAND3 (N405, N403, N243, N51);
or OR3 (N406, N405, N165, N173);
and AND2 (N407, N394, N32);
nor NOR2 (N408, N404, N239);
xor XOR2 (N409, N406, N237);
not NOT1 (N410, N408);
or OR4 (N411, N399, N74, N230, N71);
xor XOR2 (N412, N411, N200);
or OR4 (N413, N391, N103, N154, N314);
and AND2 (N414, N412, N392);
and AND4 (N415, N407, N63, N371, N318);
nor NOR3 (N416, N396, N104, N3);
not NOT1 (N417, N414);
buf BUF1 (N418, N393);
and AND2 (N419, N418, N13);
not NOT1 (N420, N402);
not NOT1 (N421, N419);
nand NAND3 (N422, N415, N51, N379);
nor NOR4 (N423, N413, N88, N415, N116);
nor NOR3 (N424, N409, N334, N157);
not NOT1 (N425, N420);
and AND4 (N426, N425, N387, N249, N160);
not NOT1 (N427, N401);
and AND2 (N428, N427, N92);
nand NAND3 (N429, N424, N191, N192);
and AND3 (N430, N421, N149, N54);
nor NOR4 (N431, N416, N281, N179, N117);
xor XOR2 (N432, N417, N146);
nor NOR3 (N433, N430, N116, N223);
nor NOR2 (N434, N432, N143);
nand NAND3 (N435, N434, N355, N37);
not NOT1 (N436, N423);
and AND3 (N437, N426, N289, N184);
nor NOR2 (N438, N435, N327);
and AND2 (N439, N400, N434);
nand NAND3 (N440, N437, N399, N356);
xor XOR2 (N441, N439, N260);
not NOT1 (N442, N431);
not NOT1 (N443, N440);
nor NOR2 (N444, N441, N274);
and AND2 (N445, N444, N95);
nand NAND3 (N446, N438, N115, N434);
buf BUF1 (N447, N429);
nor NOR2 (N448, N446, N384);
nand NAND3 (N449, N448, N287, N313);
nor NOR4 (N450, N422, N331, N407, N131);
or OR3 (N451, N449, N337, N297);
not NOT1 (N452, N445);
nor NOR2 (N453, N410, N242);
xor XOR2 (N454, N436, N314);
and AND4 (N455, N442, N449, N402, N412);
nand NAND2 (N456, N443, N177);
buf BUF1 (N457, N428);
nand NAND4 (N458, N450, N91, N252, N382);
buf BUF1 (N459, N447);
nor NOR2 (N460, N458, N133);
and AND3 (N461, N455, N146, N209);
nand NAND2 (N462, N459, N379);
xor XOR2 (N463, N457, N373);
nand NAND3 (N464, N460, N107, N133);
nand NAND3 (N465, N453, N152, N348);
nor NOR3 (N466, N463, N444, N239);
or OR4 (N467, N452, N253, N75, N376);
buf BUF1 (N468, N456);
not NOT1 (N469, N433);
and AND4 (N470, N465, N53, N381, N276);
or OR3 (N471, N461, N392, N155);
xor XOR2 (N472, N468, N148);
nand NAND3 (N473, N466, N408, N268);
and AND4 (N474, N473, N311, N353, N457);
xor XOR2 (N475, N462, N72);
buf BUF1 (N476, N471);
nor NOR2 (N477, N454, N449);
nor NOR4 (N478, N469, N425, N282, N140);
not NOT1 (N479, N451);
and AND2 (N480, N478, N410);
xor XOR2 (N481, N467, N387);
nand NAND2 (N482, N476, N350);
nor NOR4 (N483, N480, N341, N56, N108);
not NOT1 (N484, N474);
or OR3 (N485, N481, N16, N398);
xor XOR2 (N486, N483, N375);
nand NAND4 (N487, N477, N334, N286, N291);
and AND3 (N488, N485, N406, N195);
nand NAND2 (N489, N488, N10);
or OR3 (N490, N482, N150, N17);
and AND2 (N491, N484, N192);
not NOT1 (N492, N490);
nand NAND2 (N493, N472, N421);
not NOT1 (N494, N475);
not NOT1 (N495, N487);
and AND4 (N496, N479, N22, N353, N462);
nand NAND2 (N497, N496, N356);
nor NOR2 (N498, N494, N443);
xor XOR2 (N499, N470, N94);
buf BUF1 (N500, N492);
nor NOR4 (N501, N486, N181, N450, N457);
or OR4 (N502, N489, N257, N101, N404);
nor NOR2 (N503, N495, N158);
and AND4 (N504, N491, N22, N212, N310);
and AND3 (N505, N500, N266, N75);
xor XOR2 (N506, N464, N11);
and AND3 (N507, N502, N353, N397);
buf BUF1 (N508, N501);
nor NOR2 (N509, N503, N109);
buf BUF1 (N510, N507);
and AND4 (N511, N508, N264, N263, N205);
or OR4 (N512, N511, N34, N362, N57);
or OR4 (N513, N499, N234, N347, N460);
and AND4 (N514, N505, N465, N36, N368);
not NOT1 (N515, N497);
xor XOR2 (N516, N506, N411);
buf BUF1 (N517, N509);
nand NAND3 (N518, N514, N480, N212);
and AND3 (N519, N517, N348, N498);
nand NAND2 (N520, N98, N172);
or OR3 (N521, N493, N255, N218);
or OR4 (N522, N520, N517, N240, N308);
nand NAND4 (N523, N522, N370, N345, N236);
buf BUF1 (N524, N519);
and AND2 (N525, N521, N200);
buf BUF1 (N526, N504);
not NOT1 (N527, N513);
and AND4 (N528, N515, N17, N281, N456);
buf BUF1 (N529, N526);
xor XOR2 (N530, N510, N236);
not NOT1 (N531, N516);
nor NOR3 (N532, N523, N395, N23);
or OR3 (N533, N524, N332, N59);
and AND2 (N534, N530, N418);
xor XOR2 (N535, N532, N163);
buf BUF1 (N536, N533);
xor XOR2 (N537, N527, N152);
and AND4 (N538, N531, N317, N409, N378);
nand NAND3 (N539, N512, N201, N504);
not NOT1 (N540, N518);
nor NOR4 (N541, N525, N369, N483, N184);
xor XOR2 (N542, N535, N173);
xor XOR2 (N543, N528, N214);
buf BUF1 (N544, N537);
and AND2 (N545, N540, N359);
nor NOR2 (N546, N543, N67);
and AND2 (N547, N538, N353);
and AND4 (N548, N541, N158, N176, N30);
nand NAND3 (N549, N539, N136, N211);
xor XOR2 (N550, N549, N173);
not NOT1 (N551, N536);
nor NOR3 (N552, N534, N510, N148);
buf BUF1 (N553, N546);
or OR4 (N554, N550, N116, N289, N330);
nand NAND2 (N555, N551, N515);
not NOT1 (N556, N552);
and AND4 (N557, N555, N30, N73, N39);
buf BUF1 (N558, N547);
and AND4 (N559, N542, N557, N533, N443);
buf BUF1 (N560, N101);
xor XOR2 (N561, N556, N297);
xor XOR2 (N562, N560, N234);
xor XOR2 (N563, N545, N448);
nand NAND2 (N564, N548, N393);
nand NAND4 (N565, N561, N191, N563, N184);
buf BUF1 (N566, N399);
and AND4 (N567, N565, N216, N464, N36);
xor XOR2 (N568, N562, N244);
nand NAND4 (N569, N553, N219, N404, N23);
not NOT1 (N570, N544);
or OR4 (N571, N529, N384, N34, N80);
buf BUF1 (N572, N558);
xor XOR2 (N573, N569, N334);
xor XOR2 (N574, N567, N458);
nor NOR4 (N575, N572, N534, N381, N379);
xor XOR2 (N576, N570, N328);
xor XOR2 (N577, N576, N27);
xor XOR2 (N578, N575, N214);
not NOT1 (N579, N554);
buf BUF1 (N580, N566);
or OR2 (N581, N577, N249);
nor NOR4 (N582, N568, N222, N267, N47);
not NOT1 (N583, N581);
xor XOR2 (N584, N579, N134);
not NOT1 (N585, N578);
xor XOR2 (N586, N580, N401);
or OR4 (N587, N574, N227, N178, N155);
buf BUF1 (N588, N564);
and AND3 (N589, N559, N474, N86);
buf BUF1 (N590, N584);
or OR3 (N591, N590, N258, N122);
and AND2 (N592, N585, N141);
xor XOR2 (N593, N573, N226);
and AND4 (N594, N586, N447, N201, N280);
xor XOR2 (N595, N594, N80);
buf BUF1 (N596, N588);
xor XOR2 (N597, N582, N138);
not NOT1 (N598, N589);
or OR3 (N599, N596, N122, N363);
not NOT1 (N600, N599);
nor NOR4 (N601, N591, N236, N274, N463);
nand NAND4 (N602, N593, N293, N499, N452);
nor NOR2 (N603, N601, N564);
or OR4 (N604, N603, N343, N180, N466);
or OR4 (N605, N602, N487, N154, N23);
xor XOR2 (N606, N587, N59);
and AND4 (N607, N600, N458, N159, N5);
and AND2 (N608, N583, N191);
nor NOR2 (N609, N571, N206);
or OR3 (N610, N597, N506, N520);
and AND3 (N611, N605, N137, N195);
buf BUF1 (N612, N609);
nor NOR3 (N613, N607, N184, N103);
buf BUF1 (N614, N611);
and AND2 (N615, N612, N286);
not NOT1 (N616, N614);
not NOT1 (N617, N616);
nand NAND4 (N618, N598, N69, N84, N393);
xor XOR2 (N619, N604, N97);
nand NAND3 (N620, N610, N18, N94);
xor XOR2 (N621, N595, N114);
not NOT1 (N622, N619);
nand NAND2 (N623, N608, N217);
xor XOR2 (N624, N592, N256);
not NOT1 (N625, N623);
nor NOR3 (N626, N625, N193, N174);
xor XOR2 (N627, N621, N546);
buf BUF1 (N628, N618);
xor XOR2 (N629, N620, N507);
and AND2 (N630, N627, N608);
or OR4 (N631, N628, N89, N251, N238);
nand NAND4 (N632, N613, N530, N622, N275);
or OR3 (N633, N295, N208, N264);
nor NOR2 (N634, N631, N378);
and AND4 (N635, N626, N124, N383, N119);
nand NAND4 (N636, N632, N173, N175, N35);
or OR4 (N637, N615, N301, N174, N411);
or OR3 (N638, N617, N29, N337);
and AND3 (N639, N634, N361, N500);
xor XOR2 (N640, N606, N235);
and AND4 (N641, N630, N55, N391, N613);
not NOT1 (N642, N624);
not NOT1 (N643, N636);
not NOT1 (N644, N635);
not NOT1 (N645, N640);
nor NOR4 (N646, N643, N527, N513, N577);
or OR4 (N647, N629, N304, N274, N620);
nor NOR2 (N648, N633, N220);
not NOT1 (N649, N639);
nor NOR3 (N650, N645, N186, N298);
xor XOR2 (N651, N638, N638);
nor NOR2 (N652, N641, N118);
not NOT1 (N653, N644);
or OR4 (N654, N637, N297, N431, N90);
or OR4 (N655, N642, N567, N142, N369);
xor XOR2 (N656, N652, N8);
not NOT1 (N657, N653);
not NOT1 (N658, N647);
and AND2 (N659, N654, N187);
nor NOR2 (N660, N646, N611);
or OR4 (N661, N658, N344, N101, N585);
nor NOR4 (N662, N650, N431, N625, N577);
buf BUF1 (N663, N661);
buf BUF1 (N664, N656);
xor XOR2 (N665, N659, N473);
and AND4 (N666, N648, N119, N308, N60);
or OR4 (N667, N665, N582, N233, N539);
nand NAND2 (N668, N664, N502);
nor NOR4 (N669, N663, N655, N288, N43);
nand NAND2 (N670, N463, N425);
and AND2 (N671, N649, N449);
not NOT1 (N672, N669);
or OR2 (N673, N671, N631);
and AND2 (N674, N662, N88);
and AND3 (N675, N651, N615, N146);
not NOT1 (N676, N657);
nand NAND3 (N677, N675, N289, N222);
and AND4 (N678, N666, N459, N323, N276);
buf BUF1 (N679, N670);
xor XOR2 (N680, N673, N423);
nor NOR2 (N681, N677, N370);
xor XOR2 (N682, N672, N201);
nor NOR2 (N683, N679, N356);
xor XOR2 (N684, N674, N652);
not NOT1 (N685, N678);
xor XOR2 (N686, N681, N537);
nand NAND2 (N687, N682, N289);
nor NOR4 (N688, N686, N10, N404, N437);
or OR4 (N689, N660, N478, N514, N452);
buf BUF1 (N690, N676);
or OR2 (N691, N668, N477);
buf BUF1 (N692, N689);
or OR4 (N693, N690, N449, N649, N527);
not NOT1 (N694, N692);
or OR2 (N695, N694, N159);
not NOT1 (N696, N695);
nor NOR4 (N697, N696, N654, N135, N420);
nand NAND4 (N698, N680, N623, N313, N251);
xor XOR2 (N699, N684, N171);
not NOT1 (N700, N697);
and AND2 (N701, N685, N586);
nand NAND2 (N702, N667, N263);
nand NAND3 (N703, N699, N138, N682);
xor XOR2 (N704, N687, N179);
nand NAND2 (N705, N698, N289);
nand NAND4 (N706, N704, N403, N406, N15);
nand NAND3 (N707, N700, N10, N666);
nand NAND4 (N708, N706, N170, N62, N49);
and AND3 (N709, N702, N216, N467);
nor NOR4 (N710, N693, N520, N521, N648);
nand NAND3 (N711, N707, N155, N374);
nor NOR3 (N712, N708, N86, N49);
not NOT1 (N713, N712);
nor NOR2 (N714, N709, N152);
buf BUF1 (N715, N710);
nor NOR4 (N716, N683, N281, N294, N474);
nor NOR2 (N717, N701, N9);
not NOT1 (N718, N711);
nand NAND2 (N719, N691, N119);
not NOT1 (N720, N719);
nand NAND4 (N721, N715, N594, N362, N279);
xor XOR2 (N722, N703, N385);
nor NOR3 (N723, N716, N43, N86);
nor NOR2 (N724, N720, N526);
nor NOR2 (N725, N718, N152);
or OR4 (N726, N722, N126, N676, N650);
xor XOR2 (N727, N726, N5);
nor NOR3 (N728, N721, N101, N291);
nor NOR2 (N729, N713, N424);
and AND4 (N730, N725, N140, N118, N288);
buf BUF1 (N731, N717);
not NOT1 (N732, N727);
buf BUF1 (N733, N688);
nor NOR4 (N734, N724, N119, N282, N340);
and AND4 (N735, N734, N255, N299, N730);
xor XOR2 (N736, N710, N583);
nor NOR3 (N737, N723, N34, N678);
buf BUF1 (N738, N731);
or OR3 (N739, N732, N653, N44);
nor NOR2 (N740, N737, N309);
nor NOR3 (N741, N736, N551, N669);
nand NAND3 (N742, N738, N182, N413);
and AND2 (N743, N714, N194);
buf BUF1 (N744, N729);
nand NAND4 (N745, N741, N714, N462, N404);
xor XOR2 (N746, N743, N463);
nand NAND3 (N747, N744, N110, N71);
xor XOR2 (N748, N740, N518);
not NOT1 (N749, N745);
nand NAND2 (N750, N749, N623);
not NOT1 (N751, N742);
nor NOR2 (N752, N728, N612);
nand NAND2 (N753, N746, N341);
nand NAND3 (N754, N735, N258, N192);
xor XOR2 (N755, N705, N552);
not NOT1 (N756, N733);
nor NOR2 (N757, N756, N688);
xor XOR2 (N758, N750, N721);
nor NOR4 (N759, N754, N525, N62, N89);
nor NOR4 (N760, N752, N511, N708, N510);
nor NOR3 (N761, N753, N450, N254);
not NOT1 (N762, N757);
or OR3 (N763, N739, N220, N385);
buf BUF1 (N764, N761);
or OR4 (N765, N760, N490, N622, N389);
nor NOR3 (N766, N751, N11, N559);
xor XOR2 (N767, N755, N679);
or OR2 (N768, N767, N254);
buf BUF1 (N769, N765);
buf BUF1 (N770, N759);
or OR4 (N771, N766, N383, N18, N523);
nand NAND2 (N772, N770, N478);
xor XOR2 (N773, N769, N137);
nand NAND4 (N774, N762, N197, N228, N198);
nor NOR4 (N775, N771, N534, N436, N388);
nor NOR2 (N776, N775, N27);
xor XOR2 (N777, N763, N373);
not NOT1 (N778, N768);
or OR3 (N779, N774, N379, N393);
or OR4 (N780, N758, N129, N323, N330);
xor XOR2 (N781, N748, N725);
and AND4 (N782, N776, N497, N628, N321);
or OR4 (N783, N777, N428, N226, N26);
buf BUF1 (N784, N779);
xor XOR2 (N785, N747, N528);
buf BUF1 (N786, N773);
xor XOR2 (N787, N781, N422);
and AND2 (N788, N787, N432);
buf BUF1 (N789, N772);
xor XOR2 (N790, N764, N100);
nor NOR3 (N791, N790, N195, N147);
and AND3 (N792, N782, N710, N587);
buf BUF1 (N793, N791);
nand NAND2 (N794, N784, N412);
nand NAND2 (N795, N785, N20);
xor XOR2 (N796, N789, N737);
or OR2 (N797, N780, N294);
not NOT1 (N798, N793);
nor NOR3 (N799, N786, N570, N734);
buf BUF1 (N800, N799);
nand NAND2 (N801, N795, N212);
or OR3 (N802, N796, N311, N798);
nand NAND2 (N803, N66, N639);
nand NAND2 (N804, N778, N56);
buf BUF1 (N805, N797);
xor XOR2 (N806, N800, N756);
nand NAND2 (N807, N801, N313);
nor NOR3 (N808, N805, N346, N30);
xor XOR2 (N809, N808, N599);
buf BUF1 (N810, N809);
nand NAND3 (N811, N806, N408, N213);
xor XOR2 (N812, N807, N145);
nor NOR2 (N813, N810, N694);
or OR4 (N814, N803, N238, N731, N593);
xor XOR2 (N815, N792, N194);
xor XOR2 (N816, N794, N507);
nand NAND3 (N817, N816, N123, N174);
nand NAND2 (N818, N812, N59);
or OR2 (N819, N811, N434);
nor NOR2 (N820, N783, N791);
xor XOR2 (N821, N814, N270);
buf BUF1 (N822, N820);
buf BUF1 (N823, N813);
nor NOR3 (N824, N822, N3, N229);
xor XOR2 (N825, N802, N569);
xor XOR2 (N826, N788, N150);
or OR2 (N827, N817, N361);
nand NAND2 (N828, N819, N509);
xor XOR2 (N829, N815, N282);
buf BUF1 (N830, N826);
buf BUF1 (N831, N829);
nand NAND2 (N832, N824, N336);
nor NOR2 (N833, N804, N470);
not NOT1 (N834, N821);
or OR4 (N835, N825, N809, N358, N770);
and AND4 (N836, N830, N326, N654, N302);
or OR4 (N837, N828, N41, N485, N621);
xor XOR2 (N838, N837, N620);
buf BUF1 (N839, N838);
or OR4 (N840, N818, N702, N449, N611);
nand NAND3 (N841, N834, N257, N808);
not NOT1 (N842, N827);
xor XOR2 (N843, N831, N751);
or OR3 (N844, N839, N26, N379);
xor XOR2 (N845, N841, N376);
and AND4 (N846, N833, N659, N70, N619);
nand NAND4 (N847, N843, N100, N781, N490);
not NOT1 (N848, N835);
not NOT1 (N849, N848);
buf BUF1 (N850, N845);
not NOT1 (N851, N844);
nand NAND4 (N852, N850, N481, N16, N39);
or OR2 (N853, N852, N274);
nand NAND2 (N854, N823, N579);
nor NOR4 (N855, N832, N478, N544, N58);
nand NAND2 (N856, N847, N580);
not NOT1 (N857, N856);
not NOT1 (N858, N851);
xor XOR2 (N859, N854, N482);
or OR3 (N860, N855, N48, N538);
not NOT1 (N861, N840);
nand NAND2 (N862, N846, N482);
nand NAND3 (N863, N860, N330, N793);
nand NAND3 (N864, N857, N488, N259);
xor XOR2 (N865, N858, N140);
xor XOR2 (N866, N861, N79);
nand NAND3 (N867, N842, N780, N688);
xor XOR2 (N868, N853, N369);
nand NAND2 (N869, N864, N269);
nor NOR3 (N870, N868, N862, N197);
xor XOR2 (N871, N409, N332);
nand NAND4 (N872, N870, N227, N661, N648);
or OR2 (N873, N872, N783);
xor XOR2 (N874, N871, N861);
not NOT1 (N875, N869);
nand NAND4 (N876, N867, N285, N695, N742);
or OR4 (N877, N873, N42, N786, N461);
and AND2 (N878, N863, N669);
or OR2 (N879, N836, N65);
buf BUF1 (N880, N865);
not NOT1 (N881, N877);
not NOT1 (N882, N866);
xor XOR2 (N883, N876, N147);
nand NAND4 (N884, N874, N526, N758, N733);
xor XOR2 (N885, N879, N755);
and AND4 (N886, N882, N804, N415, N498);
or OR3 (N887, N878, N336, N374);
nand NAND2 (N888, N883, N88);
nand NAND2 (N889, N885, N182);
not NOT1 (N890, N889);
nor NOR4 (N891, N881, N94, N302, N662);
nor NOR4 (N892, N887, N758, N558, N394);
or OR3 (N893, N880, N219, N61);
buf BUF1 (N894, N888);
xor XOR2 (N895, N859, N131);
and AND3 (N896, N875, N42, N546);
and AND2 (N897, N895, N480);
xor XOR2 (N898, N896, N509);
buf BUF1 (N899, N891);
nand NAND3 (N900, N892, N587, N257);
or OR4 (N901, N893, N510, N304, N127);
xor XOR2 (N902, N884, N487);
xor XOR2 (N903, N849, N315);
buf BUF1 (N904, N894);
or OR3 (N905, N898, N151, N256);
not NOT1 (N906, N905);
and AND3 (N907, N899, N606, N15);
and AND4 (N908, N886, N366, N631, N57);
or OR2 (N909, N901, N503);
nand NAND4 (N910, N906, N351, N436, N389);
and AND3 (N911, N909, N387, N7);
not NOT1 (N912, N890);
xor XOR2 (N913, N902, N240);
and AND4 (N914, N900, N543, N523, N406);
nand NAND4 (N915, N904, N228, N257, N628);
or OR4 (N916, N908, N475, N762, N808);
nor NOR2 (N917, N916, N913);
or OR4 (N918, N175, N152, N187, N12);
buf BUF1 (N919, N914);
nor NOR2 (N920, N903, N802);
nand NAND3 (N921, N911, N335, N546);
nor NOR4 (N922, N907, N140, N796, N720);
xor XOR2 (N923, N915, N592);
or OR3 (N924, N921, N46, N167);
xor XOR2 (N925, N924, N10);
buf BUF1 (N926, N922);
or OR3 (N927, N923, N106, N857);
not NOT1 (N928, N920);
xor XOR2 (N929, N928, N790);
xor XOR2 (N930, N919, N70);
or OR3 (N931, N927, N869, N31);
buf BUF1 (N932, N918);
buf BUF1 (N933, N897);
and AND4 (N934, N912, N727, N317, N460);
nor NOR3 (N935, N930, N914, N750);
buf BUF1 (N936, N931);
nand NAND3 (N937, N936, N134, N849);
or OR4 (N938, N929, N321, N451, N366);
buf BUF1 (N939, N910);
not NOT1 (N940, N933);
or OR3 (N941, N935, N500, N368);
not NOT1 (N942, N940);
xor XOR2 (N943, N925, N22);
not NOT1 (N944, N943);
nor NOR4 (N945, N938, N562, N795, N419);
buf BUF1 (N946, N941);
nor NOR3 (N947, N944, N672, N475);
or OR4 (N948, N932, N944, N710, N920);
nand NAND4 (N949, N939, N551, N215, N71);
buf BUF1 (N950, N937);
buf BUF1 (N951, N948);
and AND2 (N952, N926, N883);
not NOT1 (N953, N934);
xor XOR2 (N954, N949, N892);
nand NAND3 (N955, N954, N243, N192);
xor XOR2 (N956, N917, N335);
or OR4 (N957, N951, N565, N564, N586);
buf BUF1 (N958, N956);
buf BUF1 (N959, N947);
or OR2 (N960, N942, N513);
and AND2 (N961, N950, N485);
nand NAND4 (N962, N945, N382, N564, N947);
and AND4 (N963, N955, N249, N813, N400);
and AND4 (N964, N953, N179, N664, N187);
or OR4 (N965, N964, N639, N307, N513);
nor NOR2 (N966, N952, N949);
nor NOR3 (N967, N957, N352, N834);
not NOT1 (N968, N959);
buf BUF1 (N969, N968);
nand NAND3 (N970, N966, N60, N944);
not NOT1 (N971, N946);
nor NOR3 (N972, N971, N768, N939);
and AND3 (N973, N965, N200, N721);
or OR3 (N974, N969, N116, N926);
or OR4 (N975, N972, N869, N901, N348);
nand NAND3 (N976, N974, N896, N893);
xor XOR2 (N977, N973, N502);
buf BUF1 (N978, N967);
xor XOR2 (N979, N975, N128);
nand NAND2 (N980, N978, N608);
nand NAND3 (N981, N958, N412, N329);
buf BUF1 (N982, N963);
nand NAND3 (N983, N962, N201, N135);
xor XOR2 (N984, N981, N300);
buf BUF1 (N985, N983);
not NOT1 (N986, N976);
or OR2 (N987, N986, N289);
not NOT1 (N988, N982);
or OR3 (N989, N984, N661, N752);
not NOT1 (N990, N980);
not NOT1 (N991, N960);
or OR4 (N992, N990, N97, N363, N956);
and AND3 (N993, N979, N854, N421);
not NOT1 (N994, N993);
xor XOR2 (N995, N992, N2);
not NOT1 (N996, N988);
nor NOR4 (N997, N996, N612, N532, N932);
xor XOR2 (N998, N991, N997);
xor XOR2 (N999, N322, N122);
nand NAND4 (N1000, N970, N227, N180, N859);
not NOT1 (N1001, N995);
and AND3 (N1002, N961, N385, N269);
not NOT1 (N1003, N987);
not NOT1 (N1004, N994);
nand NAND3 (N1005, N999, N591, N937);
buf BUF1 (N1006, N1005);
or OR2 (N1007, N989, N251);
not NOT1 (N1008, N1007);
buf BUF1 (N1009, N998);
not NOT1 (N1010, N1006);
nor NOR3 (N1011, N1009, N410, N346);
xor XOR2 (N1012, N977, N420);
or OR4 (N1013, N1003, N556, N686, N622);
nor NOR3 (N1014, N1008, N2, N914);
xor XOR2 (N1015, N1013, N247);
nand NAND2 (N1016, N1000, N348);
nand NAND2 (N1017, N1016, N58);
not NOT1 (N1018, N985);
or OR3 (N1019, N1011, N618, N304);
xor XOR2 (N1020, N1017, N533);
not NOT1 (N1021, N1018);
buf BUF1 (N1022, N1019);
buf BUF1 (N1023, N1002);
not NOT1 (N1024, N1022);
nor NOR4 (N1025, N1020, N719, N313, N941);
buf BUF1 (N1026, N1023);
not NOT1 (N1027, N1001);
nor NOR4 (N1028, N1012, N516, N276, N929);
nand NAND3 (N1029, N1024, N479, N946);
and AND2 (N1030, N1026, N990);
and AND2 (N1031, N1029, N135);
buf BUF1 (N1032, N1027);
not NOT1 (N1033, N1032);
nand NAND4 (N1034, N1031, N537, N142, N729);
nor NOR2 (N1035, N1025, N652);
xor XOR2 (N1036, N1014, N61);
nand NAND2 (N1037, N1036, N23);
xor XOR2 (N1038, N1033, N464);
and AND3 (N1039, N1038, N817, N877);
or OR2 (N1040, N1004, N761);
and AND4 (N1041, N1010, N54, N720, N937);
buf BUF1 (N1042, N1037);
buf BUF1 (N1043, N1041);
xor XOR2 (N1044, N1042, N418);
buf BUF1 (N1045, N1044);
buf BUF1 (N1046, N1039);
or OR2 (N1047, N1043, N563);
and AND3 (N1048, N1028, N33, N953);
not NOT1 (N1049, N1040);
and AND2 (N1050, N1045, N506);
nand NAND2 (N1051, N1048, N139);
not NOT1 (N1052, N1051);
xor XOR2 (N1053, N1021, N863);
and AND4 (N1054, N1049, N698, N899, N609);
nand NAND3 (N1055, N1046, N449, N207);
nand NAND2 (N1056, N1015, N541);
nand NAND4 (N1057, N1054, N744, N320, N434);
xor XOR2 (N1058, N1055, N970);
not NOT1 (N1059, N1053);
and AND4 (N1060, N1047, N500, N564, N97);
buf BUF1 (N1061, N1030);
and AND3 (N1062, N1061, N366, N428);
not NOT1 (N1063, N1057);
xor XOR2 (N1064, N1056, N315);
or OR3 (N1065, N1034, N275, N517);
nand NAND2 (N1066, N1065, N1053);
nor NOR2 (N1067, N1058, N868);
nor NOR4 (N1068, N1050, N257, N43, N640);
and AND2 (N1069, N1052, N1042);
nand NAND3 (N1070, N1064, N1055, N821);
and AND3 (N1071, N1068, N296, N20);
nand NAND2 (N1072, N1062, N763);
nand NAND4 (N1073, N1063, N386, N332, N32);
xor XOR2 (N1074, N1071, N209);
and AND2 (N1075, N1070, N587);
or OR4 (N1076, N1060, N554, N38, N45);
xor XOR2 (N1077, N1073, N148);
nand NAND3 (N1078, N1035, N315, N414);
not NOT1 (N1079, N1076);
or OR3 (N1080, N1059, N695, N354);
xor XOR2 (N1081, N1066, N477);
not NOT1 (N1082, N1069);
xor XOR2 (N1083, N1067, N485);
not NOT1 (N1084, N1077);
xor XOR2 (N1085, N1082, N1033);
not NOT1 (N1086, N1079);
nor NOR2 (N1087, N1072, N264);
and AND2 (N1088, N1084, N629);
and AND3 (N1089, N1080, N620, N207);
and AND3 (N1090, N1081, N706, N297);
or OR3 (N1091, N1090, N603, N1034);
buf BUF1 (N1092, N1088);
buf BUF1 (N1093, N1086);
not NOT1 (N1094, N1093);
buf BUF1 (N1095, N1085);
nand NAND4 (N1096, N1078, N967, N964, N706);
not NOT1 (N1097, N1087);
and AND3 (N1098, N1089, N272, N974);
xor XOR2 (N1099, N1074, N463);
or OR2 (N1100, N1075, N585);
xor XOR2 (N1101, N1083, N512);
xor XOR2 (N1102, N1100, N505);
buf BUF1 (N1103, N1097);
nand NAND4 (N1104, N1092, N949, N38, N937);
nor NOR3 (N1105, N1104, N1059, N969);
nor NOR2 (N1106, N1096, N577);
nor NOR3 (N1107, N1094, N331, N121);
or OR4 (N1108, N1103, N400, N72, N212);
and AND2 (N1109, N1095, N382);
or OR4 (N1110, N1102, N485, N483, N256);
nor NOR3 (N1111, N1106, N603, N750);
nor NOR2 (N1112, N1109, N154);
or OR4 (N1113, N1108, N664, N694, N1088);
not NOT1 (N1114, N1101);
xor XOR2 (N1115, N1110, N281);
nand NAND4 (N1116, N1107, N166, N892, N312);
buf BUF1 (N1117, N1091);
buf BUF1 (N1118, N1113);
not NOT1 (N1119, N1114);
nand NAND4 (N1120, N1115, N719, N593, N379);
and AND2 (N1121, N1112, N816);
not NOT1 (N1122, N1121);
and AND4 (N1123, N1119, N264, N1003, N247);
xor XOR2 (N1124, N1120, N1064);
nor NOR2 (N1125, N1124, N401);
or OR4 (N1126, N1117, N521, N1040, N836);
or OR4 (N1127, N1098, N576, N49, N1041);
not NOT1 (N1128, N1125);
buf BUF1 (N1129, N1105);
buf BUF1 (N1130, N1111);
nand NAND4 (N1131, N1116, N127, N849, N153);
and AND2 (N1132, N1127, N234);
nor NOR4 (N1133, N1131, N112, N1110, N721);
nor NOR2 (N1134, N1122, N40);
nand NAND2 (N1135, N1126, N831);
nor NOR3 (N1136, N1123, N336, N10);
or OR2 (N1137, N1128, N740);
nand NAND3 (N1138, N1099, N964, N334);
buf BUF1 (N1139, N1129);
nor NOR4 (N1140, N1139, N74, N436, N195);
nand NAND2 (N1141, N1134, N11);
or OR2 (N1142, N1136, N574);
nor NOR4 (N1143, N1140, N999, N417, N1045);
nor NOR4 (N1144, N1141, N540, N1032, N700);
nand NAND4 (N1145, N1135, N220, N1016, N179);
xor XOR2 (N1146, N1143, N299);
nor NOR3 (N1147, N1144, N1112, N93);
nor NOR2 (N1148, N1130, N759);
or OR2 (N1149, N1146, N676);
and AND2 (N1150, N1148, N1035);
nor NOR4 (N1151, N1133, N761, N214, N288);
or OR3 (N1152, N1142, N79, N1090);
xor XOR2 (N1153, N1152, N382);
nor NOR4 (N1154, N1147, N810, N751, N439);
and AND3 (N1155, N1149, N635, N537);
and AND2 (N1156, N1150, N380);
nand NAND3 (N1157, N1132, N949, N1141);
and AND3 (N1158, N1138, N416, N1003);
and AND4 (N1159, N1151, N827, N1141, N574);
not NOT1 (N1160, N1145);
and AND2 (N1161, N1137, N1090);
buf BUF1 (N1162, N1156);
and AND4 (N1163, N1161, N972, N1048, N843);
xor XOR2 (N1164, N1118, N494);
xor XOR2 (N1165, N1162, N761);
or OR3 (N1166, N1155, N124, N1128);
not NOT1 (N1167, N1159);
buf BUF1 (N1168, N1167);
and AND3 (N1169, N1160, N496, N130);
xor XOR2 (N1170, N1169, N1149);
nor NOR2 (N1171, N1165, N940);
nor NOR2 (N1172, N1164, N911);
not NOT1 (N1173, N1163);
nor NOR2 (N1174, N1168, N332);
nand NAND2 (N1175, N1174, N787);
and AND3 (N1176, N1158, N725, N565);
buf BUF1 (N1177, N1172);
or OR2 (N1178, N1170, N826);
buf BUF1 (N1179, N1177);
xor XOR2 (N1180, N1179, N361);
or OR2 (N1181, N1153, N392);
nor NOR3 (N1182, N1181, N1161, N334);
or OR4 (N1183, N1173, N1092, N1164, N219);
xor XOR2 (N1184, N1175, N154);
nor NOR2 (N1185, N1157, N778);
nor NOR4 (N1186, N1182, N1075, N1153, N760);
nand NAND4 (N1187, N1184, N232, N1091, N380);
nand NAND4 (N1188, N1185, N1118, N703, N1185);
xor XOR2 (N1189, N1176, N1013);
buf BUF1 (N1190, N1171);
or OR3 (N1191, N1183, N441, N941);
and AND2 (N1192, N1154, N583);
not NOT1 (N1193, N1180);
and AND2 (N1194, N1192, N441);
or OR3 (N1195, N1187, N299, N710);
buf BUF1 (N1196, N1186);
and AND2 (N1197, N1191, N250);
and AND4 (N1198, N1193, N281, N385, N832);
or OR2 (N1199, N1195, N1127);
not NOT1 (N1200, N1196);
nand NAND3 (N1201, N1200, N815, N1168);
xor XOR2 (N1202, N1194, N213);
and AND2 (N1203, N1197, N1055);
xor XOR2 (N1204, N1198, N606);
and AND2 (N1205, N1204, N156);
not NOT1 (N1206, N1201);
xor XOR2 (N1207, N1206, N637);
not NOT1 (N1208, N1190);
and AND3 (N1209, N1203, N520, N739);
buf BUF1 (N1210, N1205);
not NOT1 (N1211, N1208);
not NOT1 (N1212, N1209);
nand NAND4 (N1213, N1189, N1095, N969, N1010);
not NOT1 (N1214, N1213);
or OR2 (N1215, N1212, N384);
or OR2 (N1216, N1188, N1051);
not NOT1 (N1217, N1178);
and AND3 (N1218, N1217, N802, N15);
nor NOR4 (N1219, N1211, N987, N662, N814);
buf BUF1 (N1220, N1199);
and AND2 (N1221, N1166, N626);
or OR4 (N1222, N1220, N283, N187, N146);
buf BUF1 (N1223, N1214);
nor NOR4 (N1224, N1207, N528, N1169, N207);
buf BUF1 (N1225, N1210);
nor NOR4 (N1226, N1216, N727, N1125, N207);
buf BUF1 (N1227, N1202);
and AND3 (N1228, N1218, N577, N67);
nor NOR2 (N1229, N1222, N1098);
not NOT1 (N1230, N1228);
buf BUF1 (N1231, N1219);
nor NOR3 (N1232, N1223, N1002, N1051);
nand NAND4 (N1233, N1227, N288, N719, N13);
nand NAND3 (N1234, N1225, N252, N681);
nor NOR4 (N1235, N1233, N1207, N246, N975);
and AND3 (N1236, N1232, N523, N735);
and AND4 (N1237, N1230, N419, N455, N363);
nor NOR4 (N1238, N1231, N379, N462, N864);
not NOT1 (N1239, N1215);
or OR3 (N1240, N1234, N923, N1223);
or OR4 (N1241, N1240, N252, N1116, N457);
nand NAND3 (N1242, N1235, N301, N19);
not NOT1 (N1243, N1237);
and AND3 (N1244, N1241, N177, N1198);
not NOT1 (N1245, N1226);
buf BUF1 (N1246, N1229);
nor NOR2 (N1247, N1242, N861);
nand NAND3 (N1248, N1236, N544, N498);
not NOT1 (N1249, N1246);
xor XOR2 (N1250, N1238, N894);
xor XOR2 (N1251, N1239, N414);
nor NOR2 (N1252, N1251, N918);
buf BUF1 (N1253, N1252);
xor XOR2 (N1254, N1250, N2);
and AND2 (N1255, N1249, N730);
or OR3 (N1256, N1221, N988, N939);
or OR2 (N1257, N1253, N962);
buf BUF1 (N1258, N1243);
or OR2 (N1259, N1256, N1093);
nand NAND4 (N1260, N1244, N83, N920, N937);
or OR3 (N1261, N1254, N1188, N870);
xor XOR2 (N1262, N1255, N732);
or OR4 (N1263, N1261, N1070, N616, N133);
not NOT1 (N1264, N1257);
buf BUF1 (N1265, N1264);
xor XOR2 (N1266, N1260, N318);
and AND2 (N1267, N1248, N457);
nand NAND4 (N1268, N1247, N621, N493, N1079);
and AND2 (N1269, N1263, N577);
buf BUF1 (N1270, N1265);
not NOT1 (N1271, N1267);
and AND2 (N1272, N1259, N500);
nand NAND4 (N1273, N1266, N123, N1063, N151);
or OR2 (N1274, N1271, N394);
xor XOR2 (N1275, N1274, N458);
and AND4 (N1276, N1224, N373, N124, N65);
nor NOR3 (N1277, N1245, N119, N647);
nor NOR4 (N1278, N1275, N329, N213, N593);
nand NAND4 (N1279, N1273, N1220, N197, N1066);
nand NAND2 (N1280, N1258, N1040);
buf BUF1 (N1281, N1269);
nor NOR2 (N1282, N1280, N232);
not NOT1 (N1283, N1281);
and AND2 (N1284, N1283, N1204);
nand NAND4 (N1285, N1278, N971, N517, N631);
nand NAND4 (N1286, N1276, N498, N618, N595);
and AND2 (N1287, N1277, N546);
nor NOR2 (N1288, N1272, N391);
or OR2 (N1289, N1282, N299);
xor XOR2 (N1290, N1270, N15);
or OR2 (N1291, N1290, N955);
nor NOR4 (N1292, N1268, N890, N186, N548);
nand NAND2 (N1293, N1285, N404);
and AND3 (N1294, N1286, N691, N602);
xor XOR2 (N1295, N1288, N259);
nand NAND3 (N1296, N1291, N905, N1232);
nand NAND3 (N1297, N1296, N701, N1129);
and AND2 (N1298, N1294, N913);
nor NOR3 (N1299, N1289, N601, N897);
not NOT1 (N1300, N1292);
nor NOR3 (N1301, N1298, N567, N32);
xor XOR2 (N1302, N1301, N643);
xor XOR2 (N1303, N1279, N654);
nor NOR2 (N1304, N1295, N58);
xor XOR2 (N1305, N1304, N67);
and AND4 (N1306, N1299, N1161, N191, N78);
buf BUF1 (N1307, N1297);
not NOT1 (N1308, N1306);
or OR2 (N1309, N1284, N966);
buf BUF1 (N1310, N1303);
or OR3 (N1311, N1309, N692, N30);
nor NOR3 (N1312, N1307, N161, N1296);
or OR2 (N1313, N1312, N893);
not NOT1 (N1314, N1311);
nand NAND4 (N1315, N1308, N1031, N1159, N254);
xor XOR2 (N1316, N1315, N77);
nand NAND4 (N1317, N1310, N1092, N127, N990);
nor NOR4 (N1318, N1316, N944, N1317, N163);
and AND2 (N1319, N375, N1129);
nor NOR2 (N1320, N1302, N191);
buf BUF1 (N1321, N1318);
nand NAND4 (N1322, N1321, N701, N707, N1041);
not NOT1 (N1323, N1314);
not NOT1 (N1324, N1262);
and AND4 (N1325, N1324, N836, N280, N957);
or OR3 (N1326, N1322, N93, N562);
nor NOR4 (N1327, N1326, N21, N1121, N84);
nand NAND4 (N1328, N1327, N899, N608, N1293);
and AND2 (N1329, N948, N781);
nand NAND3 (N1330, N1323, N1310, N12);
or OR2 (N1331, N1330, N417);
or OR4 (N1332, N1320, N655, N626, N907);
buf BUF1 (N1333, N1305);
xor XOR2 (N1334, N1319, N319);
and AND3 (N1335, N1333, N686, N1227);
and AND2 (N1336, N1325, N829);
nand NAND4 (N1337, N1335, N911, N1027, N628);
nor NOR2 (N1338, N1329, N649);
not NOT1 (N1339, N1336);
and AND2 (N1340, N1334, N635);
not NOT1 (N1341, N1313);
buf BUF1 (N1342, N1331);
not NOT1 (N1343, N1332);
nand NAND2 (N1344, N1340, N215);
xor XOR2 (N1345, N1344, N781);
nor NOR3 (N1346, N1342, N1255, N607);
not NOT1 (N1347, N1345);
nor NOR4 (N1348, N1337, N1212, N313, N1302);
or OR4 (N1349, N1338, N692, N633, N726);
or OR4 (N1350, N1349, N436, N463, N806);
not NOT1 (N1351, N1350);
buf BUF1 (N1352, N1348);
buf BUF1 (N1353, N1287);
nor NOR3 (N1354, N1341, N896, N1160);
and AND4 (N1355, N1328, N240, N1090, N611);
buf BUF1 (N1356, N1352);
buf BUF1 (N1357, N1355);
nand NAND2 (N1358, N1346, N406);
and AND2 (N1359, N1351, N383);
or OR3 (N1360, N1358, N901, N1005);
xor XOR2 (N1361, N1356, N549);
not NOT1 (N1362, N1354);
nand NAND2 (N1363, N1339, N272);
nor NOR2 (N1364, N1363, N950);
nor NOR4 (N1365, N1360, N1068, N976, N1105);
and AND3 (N1366, N1359, N353, N703);
nor NOR4 (N1367, N1362, N409, N1294, N173);
nand NAND2 (N1368, N1367, N572);
and AND3 (N1369, N1343, N797, N700);
xor XOR2 (N1370, N1300, N497);
not NOT1 (N1371, N1368);
buf BUF1 (N1372, N1371);
or OR2 (N1373, N1372, N857);
nand NAND4 (N1374, N1366, N151, N1046, N79);
xor XOR2 (N1375, N1357, N1106);
buf BUF1 (N1376, N1347);
and AND2 (N1377, N1353, N373);
or OR3 (N1378, N1369, N441, N406);
nor NOR3 (N1379, N1361, N724, N1331);
nand NAND2 (N1380, N1365, N297);
or OR4 (N1381, N1374, N157, N525, N643);
and AND4 (N1382, N1376, N311, N869, N943);
nand NAND4 (N1383, N1364, N717, N74, N847);
buf BUF1 (N1384, N1380);
xor XOR2 (N1385, N1373, N1190);
xor XOR2 (N1386, N1370, N808);
xor XOR2 (N1387, N1381, N1134);
nor NOR4 (N1388, N1383, N377, N943, N211);
nor NOR4 (N1389, N1379, N449, N1100, N740);
xor XOR2 (N1390, N1385, N911);
not NOT1 (N1391, N1386);
not NOT1 (N1392, N1389);
nor NOR4 (N1393, N1387, N673, N11, N1151);
or OR2 (N1394, N1378, N235);
or OR2 (N1395, N1382, N599);
and AND3 (N1396, N1384, N832, N55);
xor XOR2 (N1397, N1391, N199);
not NOT1 (N1398, N1397);
nor NOR3 (N1399, N1375, N1387, N1163);
or OR2 (N1400, N1396, N322);
nor NOR3 (N1401, N1398, N1117, N231);
nand NAND2 (N1402, N1392, N1042);
xor XOR2 (N1403, N1399, N50);
or OR3 (N1404, N1400, N1380, N36);
buf BUF1 (N1405, N1404);
and AND2 (N1406, N1405, N671);
nor NOR4 (N1407, N1403, N216, N1050, N652);
or OR3 (N1408, N1390, N12, N1077);
not NOT1 (N1409, N1377);
nand NAND4 (N1410, N1401, N663, N1132, N1186);
and AND4 (N1411, N1388, N1086, N1278, N818);
nand NAND2 (N1412, N1394, N872);
and AND2 (N1413, N1408, N197);
xor XOR2 (N1414, N1407, N687);
not NOT1 (N1415, N1402);
and AND4 (N1416, N1413, N995, N1352, N144);
nand NAND3 (N1417, N1393, N886, N465);
and AND3 (N1418, N1417, N911, N1215);
and AND3 (N1419, N1410, N1094, N236);
or OR2 (N1420, N1418, N244);
nand NAND3 (N1421, N1420, N305, N1301);
nor NOR2 (N1422, N1411, N778);
nand NAND2 (N1423, N1412, N591);
not NOT1 (N1424, N1419);
not NOT1 (N1425, N1414);
and AND4 (N1426, N1415, N306, N614, N1202);
xor XOR2 (N1427, N1416, N121);
buf BUF1 (N1428, N1425);
xor XOR2 (N1429, N1426, N467);
xor XOR2 (N1430, N1423, N869);
and AND4 (N1431, N1424, N449, N629, N929);
and AND3 (N1432, N1428, N564, N461);
not NOT1 (N1433, N1421);
xor XOR2 (N1434, N1395, N663);
buf BUF1 (N1435, N1431);
not NOT1 (N1436, N1433);
nand NAND4 (N1437, N1436, N966, N1063, N1176);
xor XOR2 (N1438, N1409, N204);
nand NAND2 (N1439, N1437, N240);
or OR4 (N1440, N1422, N186, N917, N1149);
nand NAND2 (N1441, N1440, N495);
nor NOR2 (N1442, N1430, N684);
not NOT1 (N1443, N1441);
and AND2 (N1444, N1434, N59);
nand NAND2 (N1445, N1432, N1294);
xor XOR2 (N1446, N1438, N690);
not NOT1 (N1447, N1446);
or OR2 (N1448, N1442, N1021);
and AND2 (N1449, N1445, N232);
xor XOR2 (N1450, N1427, N733);
nor NOR4 (N1451, N1429, N431, N112, N317);
buf BUF1 (N1452, N1447);
and AND4 (N1453, N1443, N92, N538, N346);
buf BUF1 (N1454, N1451);
xor XOR2 (N1455, N1452, N1306);
nand NAND2 (N1456, N1448, N915);
xor XOR2 (N1457, N1444, N1414);
xor XOR2 (N1458, N1453, N653);
nor NOR4 (N1459, N1435, N100, N379, N530);
nand NAND2 (N1460, N1457, N1037);
nand NAND3 (N1461, N1450, N881, N231);
or OR4 (N1462, N1406, N659, N1272, N683);
nand NAND3 (N1463, N1462, N24, N1366);
buf BUF1 (N1464, N1461);
nand NAND3 (N1465, N1460, N1415, N973);
and AND3 (N1466, N1463, N674, N96);
buf BUF1 (N1467, N1454);
buf BUF1 (N1468, N1467);
not NOT1 (N1469, N1466);
xor XOR2 (N1470, N1464, N1338);
or OR4 (N1471, N1455, N938, N869, N102);
nand NAND4 (N1472, N1471, N318, N357, N611);
not NOT1 (N1473, N1465);
xor XOR2 (N1474, N1472, N429);
nand NAND4 (N1475, N1473, N1057, N789, N1019);
xor XOR2 (N1476, N1468, N1161);
nand NAND3 (N1477, N1456, N176, N416);
or OR2 (N1478, N1458, N1300);
xor XOR2 (N1479, N1478, N76);
nor NOR2 (N1480, N1476, N817);
or OR2 (N1481, N1477, N1134);
xor XOR2 (N1482, N1469, N1425);
xor XOR2 (N1483, N1482, N618);
or OR2 (N1484, N1449, N129);
and AND4 (N1485, N1439, N1035, N1338, N1106);
buf BUF1 (N1486, N1459);
nand NAND4 (N1487, N1470, N939, N530, N1107);
or OR4 (N1488, N1487, N1156, N662, N1203);
or OR2 (N1489, N1480, N1226);
not NOT1 (N1490, N1489);
buf BUF1 (N1491, N1483);
or OR3 (N1492, N1479, N150, N1061);
not NOT1 (N1493, N1481);
and AND2 (N1494, N1475, N642);
not NOT1 (N1495, N1491);
xor XOR2 (N1496, N1474, N30);
xor XOR2 (N1497, N1490, N1222);
xor XOR2 (N1498, N1493, N988);
and AND2 (N1499, N1492, N258);
xor XOR2 (N1500, N1499, N550);
or OR2 (N1501, N1495, N366);
nor NOR4 (N1502, N1497, N890, N886, N1417);
or OR3 (N1503, N1502, N1496, N1459);
or OR2 (N1504, N1441, N511);
not NOT1 (N1505, N1485);
nand NAND3 (N1506, N1486, N596, N1195);
and AND2 (N1507, N1501, N782);
or OR4 (N1508, N1503, N1019, N135, N509);
buf BUF1 (N1509, N1494);
nand NAND4 (N1510, N1507, N607, N104, N371);
buf BUF1 (N1511, N1484);
buf BUF1 (N1512, N1511);
xor XOR2 (N1513, N1498, N733);
and AND4 (N1514, N1506, N631, N360, N683);
buf BUF1 (N1515, N1514);
not NOT1 (N1516, N1512);
nor NOR2 (N1517, N1504, N894);
nor NOR2 (N1518, N1500, N918);
not NOT1 (N1519, N1488);
not NOT1 (N1520, N1510);
nand NAND3 (N1521, N1520, N1106, N1120);
xor XOR2 (N1522, N1508, N216);
nand NAND4 (N1523, N1516, N566, N1182, N21);
nor NOR3 (N1524, N1523, N1432, N1474);
xor XOR2 (N1525, N1519, N1137);
xor XOR2 (N1526, N1518, N290);
xor XOR2 (N1527, N1525, N623);
xor XOR2 (N1528, N1505, N1483);
xor XOR2 (N1529, N1522, N193);
nor NOR3 (N1530, N1509, N92, N416);
nor NOR2 (N1531, N1521, N1266);
buf BUF1 (N1532, N1529);
and AND4 (N1533, N1517, N446, N931, N1341);
and AND4 (N1534, N1527, N339, N1067, N1212);
and AND2 (N1535, N1530, N639);
xor XOR2 (N1536, N1535, N85);
nand NAND2 (N1537, N1531, N1253);
and AND2 (N1538, N1513, N1085);
or OR2 (N1539, N1536, N190);
xor XOR2 (N1540, N1528, N1405);
not NOT1 (N1541, N1515);
or OR2 (N1542, N1537, N259);
nand NAND4 (N1543, N1533, N1399, N665, N1162);
not NOT1 (N1544, N1539);
buf BUF1 (N1545, N1534);
not NOT1 (N1546, N1542);
or OR3 (N1547, N1541, N577, N1257);
buf BUF1 (N1548, N1526);
xor XOR2 (N1549, N1538, N462);
not NOT1 (N1550, N1546);
or OR2 (N1551, N1545, N190);
nand NAND4 (N1552, N1550, N1260, N218, N434);
nand NAND2 (N1553, N1549, N410);
nand NAND3 (N1554, N1524, N631, N179);
and AND2 (N1555, N1544, N1215);
nand NAND4 (N1556, N1551, N1007, N1145, N793);
buf BUF1 (N1557, N1552);
not NOT1 (N1558, N1555);
or OR3 (N1559, N1540, N207, N1263);
and AND2 (N1560, N1547, N11);
or OR4 (N1561, N1532, N1289, N238, N596);
xor XOR2 (N1562, N1558, N776);
xor XOR2 (N1563, N1554, N668);
not NOT1 (N1564, N1557);
buf BUF1 (N1565, N1563);
and AND4 (N1566, N1543, N1353, N136, N1565);
nor NOR3 (N1567, N434, N116, N1168);
nand NAND3 (N1568, N1567, N927, N1408);
xor XOR2 (N1569, N1561, N394);
or OR4 (N1570, N1566, N1045, N461, N643);
and AND3 (N1571, N1560, N1414, N995);
or OR4 (N1572, N1564, N967, N1528, N1481);
nor NOR3 (N1573, N1556, N1091, N639);
not NOT1 (N1574, N1571);
buf BUF1 (N1575, N1562);
or OR4 (N1576, N1548, N402, N937, N165);
nor NOR3 (N1577, N1572, N1114, N1424);
not NOT1 (N1578, N1569);
not NOT1 (N1579, N1568);
nand NAND3 (N1580, N1559, N1009, N533);
nand NAND3 (N1581, N1574, N463, N193);
buf BUF1 (N1582, N1581);
nor NOR2 (N1583, N1575, N331);
or OR4 (N1584, N1582, N426, N758, N1343);
xor XOR2 (N1585, N1577, N1163);
not NOT1 (N1586, N1553);
not NOT1 (N1587, N1578);
buf BUF1 (N1588, N1585);
nand NAND2 (N1589, N1579, N1352);
xor XOR2 (N1590, N1583, N1140);
xor XOR2 (N1591, N1576, N711);
not NOT1 (N1592, N1589);
or OR4 (N1593, N1588, N707, N611, N739);
or OR2 (N1594, N1573, N1478);
xor XOR2 (N1595, N1593, N561);
nand NAND2 (N1596, N1584, N873);
not NOT1 (N1597, N1595);
not NOT1 (N1598, N1587);
xor XOR2 (N1599, N1586, N809);
buf BUF1 (N1600, N1591);
and AND4 (N1601, N1594, N325, N1323, N221);
buf BUF1 (N1602, N1597);
xor XOR2 (N1603, N1598, N773);
nand NAND3 (N1604, N1580, N715, N911);
nor NOR3 (N1605, N1602, N1211, N635);
or OR4 (N1606, N1570, N258, N347, N25);
nand NAND2 (N1607, N1590, N598);
not NOT1 (N1608, N1601);
nand NAND4 (N1609, N1592, N348, N611, N401);
or OR2 (N1610, N1608, N1025);
nand NAND3 (N1611, N1596, N1181, N152);
and AND4 (N1612, N1605, N105, N1400, N1579);
or OR3 (N1613, N1599, N771, N1136);
nand NAND4 (N1614, N1604, N887, N1357, N663);
or OR2 (N1615, N1612, N1524);
nor NOR2 (N1616, N1606, N945);
buf BUF1 (N1617, N1610);
and AND4 (N1618, N1607, N1341, N574, N101);
nand NAND4 (N1619, N1615, N998, N123, N988);
buf BUF1 (N1620, N1611);
nor NOR2 (N1621, N1600, N845);
nand NAND2 (N1622, N1609, N792);
buf BUF1 (N1623, N1621);
xor XOR2 (N1624, N1622, N1552);
xor XOR2 (N1625, N1613, N1491);
buf BUF1 (N1626, N1619);
not NOT1 (N1627, N1618);
nand NAND3 (N1628, N1603, N608, N547);
and AND2 (N1629, N1623, N1586);
and AND2 (N1630, N1624, N858);
or OR4 (N1631, N1627, N405, N454, N412);
buf BUF1 (N1632, N1631);
buf BUF1 (N1633, N1632);
xor XOR2 (N1634, N1630, N1477);
xor XOR2 (N1635, N1625, N710);
or OR4 (N1636, N1620, N1563, N1215, N1173);
xor XOR2 (N1637, N1617, N814);
or OR4 (N1638, N1634, N147, N1551, N1016);
nand NAND3 (N1639, N1638, N804, N1112);
buf BUF1 (N1640, N1628);
nor NOR4 (N1641, N1637, N472, N414, N1425);
nor NOR2 (N1642, N1636, N823);
nor NOR3 (N1643, N1642, N1077, N1043);
or OR3 (N1644, N1641, N216, N1544);
buf BUF1 (N1645, N1626);
nor NOR3 (N1646, N1643, N932, N1012);
not NOT1 (N1647, N1645);
buf BUF1 (N1648, N1629);
not NOT1 (N1649, N1616);
xor XOR2 (N1650, N1649, N1563);
and AND3 (N1651, N1640, N1356, N1449);
or OR3 (N1652, N1648, N1512, N1338);
nor NOR4 (N1653, N1651, N418, N525, N491);
or OR3 (N1654, N1644, N1111, N1116);
and AND2 (N1655, N1654, N527);
or OR4 (N1656, N1614, N138, N1562, N36);
xor XOR2 (N1657, N1650, N1635);
buf BUF1 (N1658, N885);
not NOT1 (N1659, N1658);
xor XOR2 (N1660, N1655, N1266);
nor NOR2 (N1661, N1660, N651);
not NOT1 (N1662, N1633);
not NOT1 (N1663, N1656);
nor NOR3 (N1664, N1653, N170, N1198);
nand NAND4 (N1665, N1663, N1544, N960, N150);
nand NAND3 (N1666, N1665, N1369, N1588);
or OR2 (N1667, N1657, N1622);
or OR4 (N1668, N1652, N67, N108, N429);
not NOT1 (N1669, N1661);
not NOT1 (N1670, N1659);
and AND3 (N1671, N1669, N1558, N281);
nor NOR4 (N1672, N1639, N476, N459, N975);
nor NOR2 (N1673, N1670, N625);
xor XOR2 (N1674, N1673, N713);
nor NOR3 (N1675, N1664, N1186, N1616);
or OR4 (N1676, N1647, N1041, N1465, N418);
nor NOR4 (N1677, N1676, N1101, N1193, N157);
xor XOR2 (N1678, N1677, N1158);
and AND4 (N1679, N1667, N897, N190, N1426);
and AND4 (N1680, N1678, N1674, N34, N845);
buf BUF1 (N1681, N698);
nor NOR3 (N1682, N1646, N1110, N1641);
buf BUF1 (N1683, N1668);
and AND2 (N1684, N1679, N736);
nor NOR2 (N1685, N1684, N894);
buf BUF1 (N1686, N1682);
not NOT1 (N1687, N1671);
or OR4 (N1688, N1680, N628, N144, N267);
nand NAND4 (N1689, N1675, N1453, N66, N1042);
and AND3 (N1690, N1686, N318, N1078);
xor XOR2 (N1691, N1690, N221);
xor XOR2 (N1692, N1687, N1366);
nand NAND4 (N1693, N1672, N1684, N485, N1449);
nor NOR2 (N1694, N1688, N1025);
or OR2 (N1695, N1694, N457);
xor XOR2 (N1696, N1691, N594);
and AND3 (N1697, N1666, N1675, N787);
nand NAND3 (N1698, N1696, N551, N854);
nor NOR3 (N1699, N1697, N921, N730);
not NOT1 (N1700, N1685);
nand NAND4 (N1701, N1681, N199, N519, N388);
xor XOR2 (N1702, N1662, N1076);
nand NAND4 (N1703, N1692, N689, N1088, N1374);
nor NOR4 (N1704, N1703, N1237, N891, N415);
nor NOR2 (N1705, N1695, N955);
xor XOR2 (N1706, N1700, N760);
xor XOR2 (N1707, N1699, N1031);
xor XOR2 (N1708, N1706, N1415);
nor NOR2 (N1709, N1707, N137);
not NOT1 (N1710, N1704);
or OR2 (N1711, N1708, N1424);
or OR4 (N1712, N1693, N679, N1241, N970);
and AND2 (N1713, N1698, N1173);
buf BUF1 (N1714, N1713);
and AND2 (N1715, N1702, N770);
xor XOR2 (N1716, N1701, N92);
xor XOR2 (N1717, N1689, N1410);
xor XOR2 (N1718, N1683, N562);
nor NOR2 (N1719, N1715, N1646);
nor NOR2 (N1720, N1716, N564);
buf BUF1 (N1721, N1705);
nor NOR3 (N1722, N1712, N1647, N1376);
nand NAND2 (N1723, N1714, N262);
and AND4 (N1724, N1710, N902, N848, N1426);
xor XOR2 (N1725, N1722, N892);
nand NAND4 (N1726, N1709, N940, N376, N1029);
not NOT1 (N1727, N1725);
not NOT1 (N1728, N1723);
buf BUF1 (N1729, N1717);
or OR3 (N1730, N1711, N1257, N291);
nand NAND4 (N1731, N1727, N21, N447, N32);
nor NOR4 (N1732, N1718, N76, N1050, N171);
nand NAND3 (N1733, N1732, N1719, N798);
not NOT1 (N1734, N1503);
xor XOR2 (N1735, N1728, N823);
buf BUF1 (N1736, N1735);
nand NAND4 (N1737, N1721, N882, N646, N18);
buf BUF1 (N1738, N1731);
xor XOR2 (N1739, N1733, N589);
nor NOR3 (N1740, N1724, N488, N1524);
nor NOR2 (N1741, N1740, N689);
nor NOR2 (N1742, N1738, N1463);
and AND4 (N1743, N1729, N320, N1333, N934);
nand NAND4 (N1744, N1736, N1436, N319, N152);
or OR3 (N1745, N1743, N1496, N262);
or OR3 (N1746, N1720, N464, N102);
or OR2 (N1747, N1739, N700);
not NOT1 (N1748, N1726);
not NOT1 (N1749, N1737);
nand NAND2 (N1750, N1734, N1565);
or OR2 (N1751, N1745, N1398);
or OR3 (N1752, N1741, N371, N857);
nand NAND3 (N1753, N1748, N270, N641);
and AND4 (N1754, N1746, N97, N1001, N1374);
xor XOR2 (N1755, N1730, N383);
nand NAND4 (N1756, N1752, N1258, N1549, N1576);
nor NOR3 (N1757, N1749, N1582, N439);
and AND3 (N1758, N1747, N1287, N156);
xor XOR2 (N1759, N1750, N1745);
buf BUF1 (N1760, N1755);
nand NAND2 (N1761, N1759, N1604);
and AND3 (N1762, N1753, N1141, N484);
nor NOR4 (N1763, N1744, N386, N73, N1550);
or OR4 (N1764, N1762, N912, N1037, N1105);
xor XOR2 (N1765, N1763, N1727);
nor NOR3 (N1766, N1751, N1650, N649);
buf BUF1 (N1767, N1766);
and AND2 (N1768, N1761, N970);
not NOT1 (N1769, N1757);
nor NOR4 (N1770, N1742, N1243, N1279, N1735);
buf BUF1 (N1771, N1769);
buf BUF1 (N1772, N1754);
and AND4 (N1773, N1756, N1233, N634, N1587);
and AND4 (N1774, N1772, N98, N1603, N243);
and AND4 (N1775, N1768, N680, N283, N574);
buf BUF1 (N1776, N1774);
or OR4 (N1777, N1765, N216, N1257, N1320);
not NOT1 (N1778, N1764);
buf BUF1 (N1779, N1760);
nand NAND4 (N1780, N1779, N304, N485, N247);
buf BUF1 (N1781, N1780);
or OR3 (N1782, N1771, N1313, N1465);
nor NOR2 (N1783, N1782, N1093);
xor XOR2 (N1784, N1783, N1768);
xor XOR2 (N1785, N1767, N699);
not NOT1 (N1786, N1781);
and AND3 (N1787, N1776, N1646, N947);
nand NAND4 (N1788, N1786, N129, N207, N371);
or OR3 (N1789, N1758, N1116, N756);
not NOT1 (N1790, N1778);
nand NAND3 (N1791, N1789, N583, N254);
buf BUF1 (N1792, N1791);
buf BUF1 (N1793, N1790);
not NOT1 (N1794, N1773);
or OR3 (N1795, N1785, N1315, N1054);
and AND2 (N1796, N1777, N111);
nor NOR4 (N1797, N1796, N971, N292, N1530);
nand NAND2 (N1798, N1788, N1503);
buf BUF1 (N1799, N1795);
nor NOR2 (N1800, N1793, N1106);
and AND4 (N1801, N1787, N746, N1233, N1115);
and AND2 (N1802, N1799, N1140);
and AND2 (N1803, N1797, N244);
nor NOR4 (N1804, N1802, N1590, N1393, N930);
or OR3 (N1805, N1803, N1510, N525);
and AND3 (N1806, N1801, N1532, N992);
or OR4 (N1807, N1800, N1777, N621, N1685);
not NOT1 (N1808, N1784);
not NOT1 (N1809, N1806);
nand NAND3 (N1810, N1770, N258, N1039);
nand NAND2 (N1811, N1805, N1789);
nor NOR4 (N1812, N1811, N903, N1029, N1410);
or OR4 (N1813, N1798, N912, N27, N1306);
and AND4 (N1814, N1807, N1213, N20, N536);
xor XOR2 (N1815, N1809, N540);
and AND2 (N1816, N1815, N1802);
buf BUF1 (N1817, N1804);
nand NAND3 (N1818, N1792, N1343, N985);
or OR2 (N1819, N1812, N925);
nand NAND2 (N1820, N1817, N225);
nand NAND2 (N1821, N1819, N1610);
nor NOR3 (N1822, N1808, N912, N241);
or OR4 (N1823, N1822, N1257, N755, N1301);
nand NAND2 (N1824, N1821, N1751);
nand NAND2 (N1825, N1820, N900);
xor XOR2 (N1826, N1816, N405);
buf BUF1 (N1827, N1818);
nor NOR2 (N1828, N1810, N1213);
nor NOR3 (N1829, N1823, N26, N660);
nand NAND4 (N1830, N1828, N271, N350, N1061);
not NOT1 (N1831, N1826);
not NOT1 (N1832, N1829);
or OR4 (N1833, N1775, N48, N582, N254);
xor XOR2 (N1834, N1827, N1485);
nand NAND3 (N1835, N1833, N1697, N835);
not NOT1 (N1836, N1794);
or OR4 (N1837, N1831, N229, N718, N1397);
and AND3 (N1838, N1830, N748, N1761);
or OR3 (N1839, N1824, N1451, N1690);
nand NAND3 (N1840, N1813, N306, N766);
nand NAND4 (N1841, N1835, N332, N964, N1281);
nor NOR2 (N1842, N1841, N1674);
nand NAND2 (N1843, N1838, N105);
not NOT1 (N1844, N1843);
and AND3 (N1845, N1844, N1459, N70);
and AND3 (N1846, N1837, N484, N1384);
not NOT1 (N1847, N1836);
and AND3 (N1848, N1842, N216, N71);
buf BUF1 (N1849, N1845);
buf BUF1 (N1850, N1846);
nor NOR4 (N1851, N1839, N1653, N1493, N1748);
nor NOR2 (N1852, N1834, N874);
buf BUF1 (N1853, N1814);
and AND3 (N1854, N1852, N1099, N1055);
not NOT1 (N1855, N1832);
nor NOR2 (N1856, N1847, N1347);
nand NAND3 (N1857, N1855, N238, N571);
xor XOR2 (N1858, N1848, N1777);
buf BUF1 (N1859, N1857);
and AND3 (N1860, N1854, N381, N1103);
nand NAND4 (N1861, N1853, N1300, N1160, N161);
xor XOR2 (N1862, N1840, N51);
and AND2 (N1863, N1851, N238);
not NOT1 (N1864, N1850);
nor NOR2 (N1865, N1861, N289);
nand NAND3 (N1866, N1863, N109, N1663);
buf BUF1 (N1867, N1866);
and AND3 (N1868, N1862, N653, N1726);
nand NAND3 (N1869, N1856, N933, N56);
buf BUF1 (N1870, N1868);
buf BUF1 (N1871, N1864);
and AND2 (N1872, N1871, N1427);
xor XOR2 (N1873, N1859, N38);
or OR3 (N1874, N1825, N1240, N589);
not NOT1 (N1875, N1873);
nand NAND3 (N1876, N1849, N977, N3);
nand NAND4 (N1877, N1870, N619, N205, N143);
nor NOR2 (N1878, N1858, N886);
xor XOR2 (N1879, N1872, N1373);
not NOT1 (N1880, N1879);
xor XOR2 (N1881, N1877, N1412);
not NOT1 (N1882, N1880);
not NOT1 (N1883, N1874);
nand NAND2 (N1884, N1875, N570);
nor NOR3 (N1885, N1865, N841, N1756);
buf BUF1 (N1886, N1876);
buf BUF1 (N1887, N1860);
nand NAND2 (N1888, N1883, N1222);
or OR3 (N1889, N1887, N964, N466);
nand NAND4 (N1890, N1867, N1019, N67, N1888);
nor NOR3 (N1891, N101, N1722, N1748);
or OR3 (N1892, N1889, N1624, N154);
and AND4 (N1893, N1892, N507, N134, N1827);
nor NOR3 (N1894, N1886, N587, N887);
xor XOR2 (N1895, N1894, N590);
or OR3 (N1896, N1882, N1338, N1469);
nand NAND4 (N1897, N1881, N1082, N468, N279);
nand NAND3 (N1898, N1885, N1158, N225);
nand NAND4 (N1899, N1898, N1331, N1786, N928);
nor NOR3 (N1900, N1895, N52, N1040);
or OR4 (N1901, N1878, N186, N1818, N492);
xor XOR2 (N1902, N1884, N853);
and AND4 (N1903, N1869, N10, N930, N500);
nor NOR4 (N1904, N1897, N762, N1724, N1739);
xor XOR2 (N1905, N1899, N1766);
buf BUF1 (N1906, N1893);
nor NOR2 (N1907, N1904, N1578);
xor XOR2 (N1908, N1903, N1235);
not NOT1 (N1909, N1905);
not NOT1 (N1910, N1902);
nand NAND2 (N1911, N1896, N1465);
xor XOR2 (N1912, N1891, N396);
and AND3 (N1913, N1908, N1830, N1393);
buf BUF1 (N1914, N1906);
nand NAND2 (N1915, N1890, N341);
and AND4 (N1916, N1910, N305, N288, N1033);
xor XOR2 (N1917, N1912, N701);
buf BUF1 (N1918, N1911);
nand NAND4 (N1919, N1909, N847, N1880, N1911);
nor NOR3 (N1920, N1900, N1721, N140);
nor NOR4 (N1921, N1920, N343, N1909, N1597);
xor XOR2 (N1922, N1901, N545);
and AND2 (N1923, N1919, N1360);
nand NAND3 (N1924, N1918, N1255, N1134);
buf BUF1 (N1925, N1916);
nand NAND3 (N1926, N1922, N1084, N1739);
nor NOR4 (N1927, N1915, N842, N1716, N655);
and AND4 (N1928, N1926, N1113, N234, N615);
not NOT1 (N1929, N1928);
buf BUF1 (N1930, N1914);
nand NAND3 (N1931, N1930, N1465, N1517);
not NOT1 (N1932, N1921);
and AND2 (N1933, N1932, N397);
xor XOR2 (N1934, N1931, N940);
buf BUF1 (N1935, N1927);
not NOT1 (N1936, N1913);
nor NOR2 (N1937, N1907, N1406);
xor XOR2 (N1938, N1923, N723);
nand NAND3 (N1939, N1938, N1670, N889);
buf BUF1 (N1940, N1937);
nor NOR4 (N1941, N1934, N150, N796, N1798);
and AND2 (N1942, N1917, N987);
not NOT1 (N1943, N1935);
buf BUF1 (N1944, N1941);
or OR3 (N1945, N1936, N1904, N1499);
buf BUF1 (N1946, N1945);
or OR2 (N1947, N1943, N398);
nand NAND2 (N1948, N1939, N750);
nand NAND2 (N1949, N1944, N1254);
not NOT1 (N1950, N1942);
not NOT1 (N1951, N1929);
or OR4 (N1952, N1951, N408, N1552, N1101);
buf BUF1 (N1953, N1949);
not NOT1 (N1954, N1948);
not NOT1 (N1955, N1953);
not NOT1 (N1956, N1954);
not NOT1 (N1957, N1924);
nor NOR2 (N1958, N1933, N141);
nand NAND2 (N1959, N1958, N1296);
nand NAND2 (N1960, N1950, N694);
xor XOR2 (N1961, N1940, N1669);
xor XOR2 (N1962, N1946, N1864);
and AND3 (N1963, N1925, N1368, N1538);
nand NAND2 (N1964, N1955, N79);
xor XOR2 (N1965, N1960, N1170);
nand NAND3 (N1966, N1964, N1322, N633);
not NOT1 (N1967, N1956);
not NOT1 (N1968, N1966);
nand NAND3 (N1969, N1963, N1323, N590);
buf BUF1 (N1970, N1952);
not NOT1 (N1971, N1959);
not NOT1 (N1972, N1969);
buf BUF1 (N1973, N1957);
or OR2 (N1974, N1967, N1465);
buf BUF1 (N1975, N1973);
not NOT1 (N1976, N1972);
nand NAND4 (N1977, N1961, N1918, N449, N1475);
buf BUF1 (N1978, N1970);
or OR3 (N1979, N1976, N142, N777);
or OR3 (N1980, N1971, N505, N977);
and AND2 (N1981, N1979, N1675);
or OR3 (N1982, N1947, N1531, N1001);
or OR4 (N1983, N1982, N1071, N739, N753);
nand NAND3 (N1984, N1981, N105, N1099);
or OR2 (N1985, N1965, N349);
and AND2 (N1986, N1977, N585);
buf BUF1 (N1987, N1984);
nor NOR4 (N1988, N1985, N1431, N1742, N426);
nand NAND2 (N1989, N1988, N34);
or OR4 (N1990, N1974, N1732, N209, N1396);
nor NOR4 (N1991, N1962, N790, N713, N212);
not NOT1 (N1992, N1978);
and AND2 (N1993, N1983, N665);
and AND2 (N1994, N1990, N981);
xor XOR2 (N1995, N1992, N740);
nand NAND3 (N1996, N1980, N794, N1076);
not NOT1 (N1997, N1994);
nand NAND4 (N1998, N1995, N1134, N1853, N1483);
xor XOR2 (N1999, N1986, N1476);
not NOT1 (N2000, N1999);
or OR3 (N2001, N1998, N832, N1228);
and AND3 (N2002, N2001, N1024, N583);
buf BUF1 (N2003, N2002);
buf BUF1 (N2004, N1996);
not NOT1 (N2005, N1987);
nand NAND4 (N2006, N1968, N1819, N659, N927);
not NOT1 (N2007, N2006);
or OR3 (N2008, N1997, N993, N67);
nand NAND3 (N2009, N2004, N1150, N683);
buf BUF1 (N2010, N2007);
or OR2 (N2011, N2005, N1055);
nand NAND2 (N2012, N1993, N1095);
and AND2 (N2013, N2012, N1922);
and AND2 (N2014, N2000, N719);
nand NAND3 (N2015, N2008, N1648, N48);
or OR3 (N2016, N2014, N1878, N666);
nand NAND4 (N2017, N1975, N1405, N1288, N606);
and AND4 (N2018, N2013, N710, N412, N887);
and AND2 (N2019, N2017, N1802);
nor NOR2 (N2020, N2018, N1370);
nor NOR2 (N2021, N2019, N1305);
and AND4 (N2022, N2016, N851, N1683, N628);
xor XOR2 (N2023, N1989, N2017);
nand NAND3 (N2024, N2020, N773, N164);
nand NAND2 (N2025, N2022, N223);
xor XOR2 (N2026, N2015, N922);
and AND3 (N2027, N2011, N1833, N1074);
buf BUF1 (N2028, N1991);
and AND4 (N2029, N2028, N1205, N814, N1935);
buf BUF1 (N2030, N2009);
or OR3 (N2031, N2025, N1068, N1802);
nor NOR2 (N2032, N2023, N665);
nand NAND2 (N2033, N2003, N1144);
or OR3 (N2034, N2029, N963, N1704);
nand NAND3 (N2035, N2033, N428, N181);
not NOT1 (N2036, N2027);
and AND4 (N2037, N2034, N1799, N691, N1832);
or OR4 (N2038, N2021, N1770, N831, N104);
nand NAND4 (N2039, N2030, N1626, N242, N1812);
buf BUF1 (N2040, N2038);
nand NAND3 (N2041, N2026, N1019, N326);
or OR3 (N2042, N2041, N1041, N1243);
xor XOR2 (N2043, N2037, N432);
not NOT1 (N2044, N2032);
nand NAND2 (N2045, N2031, N1367);
xor XOR2 (N2046, N2043, N1284);
not NOT1 (N2047, N2045);
buf BUF1 (N2048, N2046);
nor NOR4 (N2049, N2024, N1019, N785, N556);
and AND3 (N2050, N2049, N526, N73);
and AND3 (N2051, N2050, N522, N981);
not NOT1 (N2052, N2048);
or OR3 (N2053, N2042, N1456, N1829);
nor NOR3 (N2054, N2035, N1445, N134);
not NOT1 (N2055, N2051);
not NOT1 (N2056, N2055);
buf BUF1 (N2057, N2044);
xor XOR2 (N2058, N2057, N369);
or OR4 (N2059, N2036, N1878, N1707, N283);
not NOT1 (N2060, N2039);
and AND3 (N2061, N2047, N294, N1766);
not NOT1 (N2062, N2060);
xor XOR2 (N2063, N2010, N1513);
nand NAND4 (N2064, N2059, N1884, N1391, N1272);
not NOT1 (N2065, N2058);
not NOT1 (N2066, N2061);
nand NAND3 (N2067, N2056, N448, N1126);
buf BUF1 (N2068, N2064);
buf BUF1 (N2069, N2063);
buf BUF1 (N2070, N2066);
and AND2 (N2071, N2053, N541);
xor XOR2 (N2072, N2054, N262);
buf BUF1 (N2073, N2068);
not NOT1 (N2074, N2072);
not NOT1 (N2075, N2069);
nor NOR4 (N2076, N2075, N1463, N310, N1676);
buf BUF1 (N2077, N2073);
xor XOR2 (N2078, N2074, N366);
nand NAND3 (N2079, N2077, N294, N1120);
nor NOR3 (N2080, N2052, N792, N940);
and AND2 (N2081, N2070, N1791);
not NOT1 (N2082, N2076);
and AND3 (N2083, N2082, N226, N2000);
and AND2 (N2084, N2081, N19);
and AND4 (N2085, N2083, N898, N1045, N157);
or OR2 (N2086, N2085, N301);
or OR4 (N2087, N2086, N599, N659, N1391);
or OR2 (N2088, N2078, N229);
nand NAND4 (N2089, N2080, N23, N1499, N1755);
xor XOR2 (N2090, N2079, N210);
nand NAND2 (N2091, N2040, N1300);
xor XOR2 (N2092, N2091, N1982);
nor NOR4 (N2093, N2071, N328, N130, N520);
not NOT1 (N2094, N2089);
xor XOR2 (N2095, N2062, N1361);
xor XOR2 (N2096, N2065, N1405);
or OR3 (N2097, N2088, N864, N1732);
xor XOR2 (N2098, N2084, N522);
or OR4 (N2099, N2087, N602, N395, N980);
and AND2 (N2100, N2092, N1707);
nand NAND4 (N2101, N2098, N323, N2036, N144);
nor NOR2 (N2102, N2093, N551);
and AND4 (N2103, N2095, N1675, N1410, N1022);
or OR4 (N2104, N2096, N1735, N507, N226);
nand NAND3 (N2105, N2094, N491, N163);
not NOT1 (N2106, N2067);
xor XOR2 (N2107, N2106, N629);
nor NOR4 (N2108, N2090, N341, N1335, N1541);
and AND3 (N2109, N2108, N736, N746);
not NOT1 (N2110, N2104);
nor NOR2 (N2111, N2110, N1568);
buf BUF1 (N2112, N2097);
buf BUF1 (N2113, N2105);
xor XOR2 (N2114, N2101, N826);
or OR3 (N2115, N2111, N1172, N996);
nand NAND4 (N2116, N2114, N1736, N1840, N1944);
xor XOR2 (N2117, N2109, N1126);
or OR4 (N2118, N2116, N790, N1159, N1940);
xor XOR2 (N2119, N2115, N265);
buf BUF1 (N2120, N2113);
xor XOR2 (N2121, N2118, N1482);
buf BUF1 (N2122, N2102);
or OR3 (N2123, N2121, N746, N1820);
not NOT1 (N2124, N2107);
nor NOR2 (N2125, N2119, N467);
not NOT1 (N2126, N2124);
xor XOR2 (N2127, N2123, N2025);
or OR3 (N2128, N2103, N1986, N1655);
and AND4 (N2129, N2100, N1011, N542, N425);
xor XOR2 (N2130, N2099, N1582);
nand NAND4 (N2131, N2112, N4, N1768, N1486);
nand NAND3 (N2132, N2122, N1717, N159);
xor XOR2 (N2133, N2120, N1809);
nand NAND4 (N2134, N2126, N1454, N1557, N1085);
buf BUF1 (N2135, N2134);
xor XOR2 (N2136, N2133, N634);
or OR3 (N2137, N2132, N1516, N1295);
and AND4 (N2138, N2117, N2048, N223, N1806);
nand NAND4 (N2139, N2135, N932, N517, N326);
nand NAND2 (N2140, N2125, N648);
not NOT1 (N2141, N2128);
buf BUF1 (N2142, N2130);
nor NOR3 (N2143, N2141, N845, N390);
nand NAND2 (N2144, N2131, N943);
buf BUF1 (N2145, N2140);
buf BUF1 (N2146, N2136);
nor NOR3 (N2147, N2138, N219, N410);
or OR3 (N2148, N2144, N1745, N93);
not NOT1 (N2149, N2147);
xor XOR2 (N2150, N2129, N249);
xor XOR2 (N2151, N2148, N1664);
nor NOR2 (N2152, N2137, N1835);
nand NAND4 (N2153, N2142, N1535, N561, N2067);
or OR4 (N2154, N2145, N951, N140, N1962);
buf BUF1 (N2155, N2149);
not NOT1 (N2156, N2154);
nand NAND2 (N2157, N2153, N295);
nand NAND4 (N2158, N2143, N2008, N247, N97);
and AND3 (N2159, N2146, N1772, N1598);
buf BUF1 (N2160, N2139);
and AND3 (N2161, N2158, N607, N70);
nor NOR4 (N2162, N2157, N1646, N887, N727);
and AND2 (N2163, N2127, N178);
or OR4 (N2164, N2151, N1891, N396, N1696);
xor XOR2 (N2165, N2152, N1933);
or OR4 (N2166, N2162, N2009, N1279, N1840);
nand NAND3 (N2167, N2161, N732, N1151);
or OR2 (N2168, N2167, N170);
and AND2 (N2169, N2160, N2072);
not NOT1 (N2170, N2166);
and AND2 (N2171, N2156, N821);
nand NAND2 (N2172, N2163, N1815);
and AND4 (N2173, N2169, N602, N2060, N105);
nand NAND2 (N2174, N2168, N1778);
xor XOR2 (N2175, N2150, N1985);
buf BUF1 (N2176, N2159);
xor XOR2 (N2177, N2165, N139);
or OR2 (N2178, N2175, N318);
or OR3 (N2179, N2177, N1251, N2012);
or OR4 (N2180, N2170, N1667, N1091, N899);
buf BUF1 (N2181, N2155);
not NOT1 (N2182, N2171);
xor XOR2 (N2183, N2164, N526);
nand NAND3 (N2184, N2176, N1617, N886);
xor XOR2 (N2185, N2182, N226);
nor NOR2 (N2186, N2185, N237);
xor XOR2 (N2187, N2180, N486);
and AND2 (N2188, N2184, N1255);
buf BUF1 (N2189, N2172);
or OR3 (N2190, N2188, N637, N45);
and AND4 (N2191, N2183, N987, N545, N517);
and AND4 (N2192, N2189, N1769, N738, N310);
and AND3 (N2193, N2178, N1758, N506);
xor XOR2 (N2194, N2191, N491);
or OR3 (N2195, N2186, N1509, N1153);
or OR3 (N2196, N2179, N1104, N273);
nor NOR2 (N2197, N2190, N325);
nand NAND4 (N2198, N2187, N1758, N286, N1406);
nor NOR3 (N2199, N2174, N788, N1505);
or OR3 (N2200, N2199, N205, N1106);
nand NAND4 (N2201, N2173, N1430, N1152, N1714);
buf BUF1 (N2202, N2196);
xor XOR2 (N2203, N2181, N680);
or OR2 (N2204, N2202, N1578);
not NOT1 (N2205, N2193);
nor NOR2 (N2206, N2198, N2068);
buf BUF1 (N2207, N2206);
nor NOR2 (N2208, N2197, N669);
and AND4 (N2209, N2200, N1098, N991, N1727);
nand NAND4 (N2210, N2208, N1347, N1448, N689);
nor NOR3 (N2211, N2201, N1529, N2030);
not NOT1 (N2212, N2204);
and AND2 (N2213, N2203, N1158);
nor NOR2 (N2214, N2205, N1376);
xor XOR2 (N2215, N2195, N467);
or OR3 (N2216, N2209, N1230, N1348);
not NOT1 (N2217, N2194);
xor XOR2 (N2218, N2210, N924);
not NOT1 (N2219, N2216);
buf BUF1 (N2220, N2207);
xor XOR2 (N2221, N2218, N402);
nand NAND3 (N2222, N2221, N1970, N1937);
nor NOR2 (N2223, N2215, N1615);
xor XOR2 (N2224, N2192, N365);
not NOT1 (N2225, N2214);
xor XOR2 (N2226, N2225, N923);
nor NOR4 (N2227, N2219, N1886, N2001, N1314);
buf BUF1 (N2228, N2227);
nor NOR4 (N2229, N2226, N589, N1603, N1049);
nor NOR2 (N2230, N2217, N186);
or OR3 (N2231, N2220, N2060, N1245);
and AND3 (N2232, N2224, N177, N226);
and AND3 (N2233, N2213, N1595, N447);
nor NOR3 (N2234, N2223, N419, N1133);
buf BUF1 (N2235, N2229);
nand NAND3 (N2236, N2230, N1102, N1116);
and AND3 (N2237, N2222, N1484, N1377);
and AND2 (N2238, N2236, N567);
or OR4 (N2239, N2237, N2080, N1712, N1780);
xor XOR2 (N2240, N2238, N1875);
nand NAND4 (N2241, N2231, N1757, N1059, N1453);
xor XOR2 (N2242, N2233, N852);
nor NOR2 (N2243, N2234, N1915);
not NOT1 (N2244, N2211);
or OR4 (N2245, N2242, N1379, N909, N232);
xor XOR2 (N2246, N2228, N1941);
buf BUF1 (N2247, N2240);
nor NOR2 (N2248, N2245, N602);
not NOT1 (N2249, N2243);
xor XOR2 (N2250, N2248, N256);
nor NOR4 (N2251, N2212, N1001, N2049, N2174);
not NOT1 (N2252, N2241);
nor NOR3 (N2253, N2246, N835, N311);
xor XOR2 (N2254, N2239, N584);
or OR4 (N2255, N2235, N351, N1117, N1292);
nor NOR3 (N2256, N2253, N1276, N297);
not NOT1 (N2257, N2247);
and AND3 (N2258, N2254, N466, N1647);
or OR2 (N2259, N2249, N479);
nor NOR3 (N2260, N2258, N13, N860);
nor NOR4 (N2261, N2232, N1468, N730, N778);
nor NOR3 (N2262, N2256, N2081, N2214);
nand NAND3 (N2263, N2262, N2007, N321);
xor XOR2 (N2264, N2261, N1684);
or OR2 (N2265, N2260, N264);
and AND2 (N2266, N2264, N1499);
or OR4 (N2267, N2251, N756, N1942, N1189);
and AND2 (N2268, N2255, N1406);
or OR4 (N2269, N2259, N595, N749, N1613);
nand NAND2 (N2270, N2244, N834);
nor NOR3 (N2271, N2270, N661, N1956);
nand NAND2 (N2272, N2250, N413);
and AND2 (N2273, N2263, N478);
nor NOR4 (N2274, N2267, N1820, N924, N1618);
not NOT1 (N2275, N2271);
or OR3 (N2276, N2252, N175, N746);
xor XOR2 (N2277, N2274, N1198);
and AND2 (N2278, N2275, N639);
or OR4 (N2279, N2278, N2108, N969, N1637);
xor XOR2 (N2280, N2273, N1329);
nor NOR3 (N2281, N2280, N1201, N329);
xor XOR2 (N2282, N2257, N1217);
nand NAND4 (N2283, N2266, N2064, N1598, N1959);
or OR4 (N2284, N2269, N1587, N1844, N2187);
nor NOR3 (N2285, N2277, N2069, N378);
not NOT1 (N2286, N2268);
nand NAND3 (N2287, N2283, N1634, N2211);
buf BUF1 (N2288, N2276);
nand NAND4 (N2289, N2286, N621, N1676, N2066);
and AND2 (N2290, N2285, N424);
nand NAND4 (N2291, N2288, N114, N887, N356);
xor XOR2 (N2292, N2265, N1707);
nor NOR4 (N2293, N2287, N1076, N2227, N1788);
not NOT1 (N2294, N2290);
and AND2 (N2295, N2291, N1140);
nor NOR3 (N2296, N2281, N2162, N651);
xor XOR2 (N2297, N2296, N1491);
buf BUF1 (N2298, N2282);
not NOT1 (N2299, N2284);
nand NAND4 (N2300, N2297, N1926, N1772, N791);
and AND4 (N2301, N2289, N198, N2264, N611);
nand NAND4 (N2302, N2299, N11, N398, N1470);
not NOT1 (N2303, N2301);
or OR4 (N2304, N2292, N811, N423, N1264);
not NOT1 (N2305, N2302);
not NOT1 (N2306, N2294);
and AND3 (N2307, N2304, N2039, N106);
nand NAND3 (N2308, N2279, N511, N2027);
nand NAND4 (N2309, N2298, N1765, N1584, N1195);
not NOT1 (N2310, N2272);
xor XOR2 (N2311, N2307, N44);
buf BUF1 (N2312, N2303);
not NOT1 (N2313, N2312);
and AND2 (N2314, N2308, N2089);
xor XOR2 (N2315, N2293, N834);
and AND3 (N2316, N2305, N912, N776);
nor NOR2 (N2317, N2313, N898);
not NOT1 (N2318, N2314);
and AND4 (N2319, N2317, N196, N902, N1009);
nand NAND3 (N2320, N2318, N1880, N1137);
nand NAND2 (N2321, N2300, N2125);
buf BUF1 (N2322, N2310);
xor XOR2 (N2323, N2295, N1954);
buf BUF1 (N2324, N2321);
nor NOR2 (N2325, N2322, N1115);
buf BUF1 (N2326, N2311);
xor XOR2 (N2327, N2326, N1602);
nand NAND3 (N2328, N2320, N1654, N627);
xor XOR2 (N2329, N2315, N2218);
xor XOR2 (N2330, N2309, N1202);
or OR2 (N2331, N2328, N1658);
nor NOR3 (N2332, N2306, N1203, N259);
nand NAND4 (N2333, N2323, N1225, N1134, N2127);
xor XOR2 (N2334, N2332, N1124);
buf BUF1 (N2335, N2324);
nor NOR2 (N2336, N2330, N986);
nor NOR3 (N2337, N2329, N1999, N1103);
xor XOR2 (N2338, N2316, N236);
xor XOR2 (N2339, N2319, N2003);
and AND2 (N2340, N2334, N594);
nor NOR3 (N2341, N2338, N1895, N1481);
not NOT1 (N2342, N2340);
nor NOR3 (N2343, N2331, N1472, N1997);
xor XOR2 (N2344, N2342, N597);
or OR2 (N2345, N2344, N1419);
buf BUF1 (N2346, N2337);
nand NAND2 (N2347, N2343, N1154);
not NOT1 (N2348, N2327);
and AND2 (N2349, N2339, N1206);
xor XOR2 (N2350, N2341, N1638);
buf BUF1 (N2351, N2336);
not NOT1 (N2352, N2350);
buf BUF1 (N2353, N2346);
nor NOR2 (N2354, N2351, N1389);
nand NAND2 (N2355, N2353, N742);
xor XOR2 (N2356, N2335, N2026);
nand NAND2 (N2357, N2333, N629);
not NOT1 (N2358, N2348);
nor NOR4 (N2359, N2325, N317, N2004, N288);
buf BUF1 (N2360, N2355);
buf BUF1 (N2361, N2358);
and AND3 (N2362, N2347, N1637, N789);
nor NOR3 (N2363, N2362, N1445, N952);
not NOT1 (N2364, N2359);
nor NOR4 (N2365, N2352, N649, N1500, N390);
buf BUF1 (N2366, N2364);
nor NOR4 (N2367, N2363, N1273, N54, N1307);
nand NAND3 (N2368, N2354, N2025, N2243);
nor NOR2 (N2369, N2345, N1289);
xor XOR2 (N2370, N2367, N948);
buf BUF1 (N2371, N2369);
buf BUF1 (N2372, N2366);
not NOT1 (N2373, N2360);
xor XOR2 (N2374, N2357, N1452);
and AND2 (N2375, N2365, N58);
buf BUF1 (N2376, N2375);
or OR4 (N2377, N2372, N1347, N344, N902);
xor XOR2 (N2378, N2370, N910);
xor XOR2 (N2379, N2361, N1625);
nor NOR2 (N2380, N2377, N2271);
or OR4 (N2381, N2376, N145, N689, N1667);
nor NOR3 (N2382, N2381, N142, N717);
or OR4 (N2383, N2380, N56, N386, N334);
nand NAND3 (N2384, N2379, N181, N161);
not NOT1 (N2385, N2378);
and AND4 (N2386, N2349, N396, N1190, N391);
nand NAND3 (N2387, N2385, N831, N302);
buf BUF1 (N2388, N2383);
buf BUF1 (N2389, N2386);
nor NOR3 (N2390, N2374, N1722, N1563);
nor NOR4 (N2391, N2384, N1963, N1529, N1008);
nand NAND4 (N2392, N2389, N553, N1068, N1966);
not NOT1 (N2393, N2387);
nand NAND4 (N2394, N2388, N1544, N970, N2022);
not NOT1 (N2395, N2371);
and AND2 (N2396, N2368, N827);
nand NAND2 (N2397, N2393, N1286);
not NOT1 (N2398, N2390);
xor XOR2 (N2399, N2392, N279);
and AND3 (N2400, N2398, N1534, N317);
not NOT1 (N2401, N2356);
buf BUF1 (N2402, N2396);
nor NOR3 (N2403, N2391, N2067, N2077);
nor NOR2 (N2404, N2382, N1463);
nor NOR4 (N2405, N2394, N1292, N334, N1187);
not NOT1 (N2406, N2403);
not NOT1 (N2407, N2395);
not NOT1 (N2408, N2405);
not NOT1 (N2409, N2402);
buf BUF1 (N2410, N2399);
nand NAND3 (N2411, N2407, N94, N1139);
xor XOR2 (N2412, N2411, N605);
xor XOR2 (N2413, N2401, N1135);
nor NOR2 (N2414, N2412, N1336);
nand NAND3 (N2415, N2409, N1706, N1993);
not NOT1 (N2416, N2397);
nor NOR4 (N2417, N2373, N139, N1248, N2020);
xor XOR2 (N2418, N2414, N1955);
xor XOR2 (N2419, N2400, N196);
nor NOR2 (N2420, N2419, N1227);
nand NAND3 (N2421, N2410, N1189, N1789);
or OR4 (N2422, N2404, N2028, N1639, N1434);
nor NOR4 (N2423, N2406, N406, N430, N2296);
or OR4 (N2424, N2415, N929, N2259, N1093);
buf BUF1 (N2425, N2413);
nor NOR2 (N2426, N2423, N63);
nand NAND3 (N2427, N2422, N1668, N1589);
nand NAND3 (N2428, N2426, N1731, N603);
and AND4 (N2429, N2417, N194, N19, N1879);
buf BUF1 (N2430, N2416);
and AND4 (N2431, N2418, N220, N1309, N84);
and AND2 (N2432, N2427, N1240);
or OR4 (N2433, N2420, N998, N1926, N2287);
or OR2 (N2434, N2430, N38);
nor NOR4 (N2435, N2408, N707, N1053, N1963);
nand NAND4 (N2436, N2433, N2192, N100, N1582);
not NOT1 (N2437, N2421);
buf BUF1 (N2438, N2428);
xor XOR2 (N2439, N2436, N131);
or OR2 (N2440, N2425, N508);
nor NOR3 (N2441, N2440, N982, N679);
or OR4 (N2442, N2432, N565, N2324, N179);
or OR3 (N2443, N2434, N2007, N1374);
buf BUF1 (N2444, N2429);
nor NOR4 (N2445, N2437, N523, N1507, N2230);
or OR3 (N2446, N2424, N1738, N800);
nor NOR3 (N2447, N2439, N1359, N35);
and AND3 (N2448, N2444, N1324, N418);
xor XOR2 (N2449, N2447, N1266);
nand NAND2 (N2450, N2435, N899);
nor NOR3 (N2451, N2445, N715, N1264);
xor XOR2 (N2452, N2443, N696);
nand NAND4 (N2453, N2449, N1966, N1325, N2148);
nand NAND2 (N2454, N2438, N2254);
or OR4 (N2455, N2453, N334, N2204, N2025);
buf BUF1 (N2456, N2448);
nand NAND3 (N2457, N2441, N1588, N2176);
buf BUF1 (N2458, N2457);
buf BUF1 (N2459, N2442);
not NOT1 (N2460, N2451);
and AND2 (N2461, N2459, N1764);
buf BUF1 (N2462, N2452);
nand NAND4 (N2463, N2450, N49, N1686, N1566);
and AND4 (N2464, N2461, N2130, N313, N1129);
or OR4 (N2465, N2458, N1716, N1778, N2119);
not NOT1 (N2466, N2455);
buf BUF1 (N2467, N2464);
and AND4 (N2468, N2465, N1423, N1110, N1884);
nor NOR2 (N2469, N2463, N1374);
not NOT1 (N2470, N2456);
nor NOR2 (N2471, N2462, N761);
xor XOR2 (N2472, N2470, N387);
or OR3 (N2473, N2460, N295, N500);
xor XOR2 (N2474, N2467, N2012);
not NOT1 (N2475, N2454);
nand NAND4 (N2476, N2471, N2206, N497, N1320);
nor NOR3 (N2477, N2469, N351, N1205);
not NOT1 (N2478, N2474);
and AND3 (N2479, N2466, N1766, N407);
nor NOR3 (N2480, N2479, N1337, N176);
nor NOR3 (N2481, N2478, N920, N62);
or OR4 (N2482, N2475, N785, N1361, N2292);
buf BUF1 (N2483, N2473);
not NOT1 (N2484, N2483);
nand NAND3 (N2485, N2431, N351, N729);
nor NOR4 (N2486, N2485, N1457, N2102, N1950);
nand NAND2 (N2487, N2484, N1684);
buf BUF1 (N2488, N2446);
nand NAND2 (N2489, N2480, N42);
buf BUF1 (N2490, N2477);
or OR2 (N2491, N2486, N2403);
and AND4 (N2492, N2487, N1095, N438, N635);
not NOT1 (N2493, N2492);
or OR2 (N2494, N2489, N182);
or OR4 (N2495, N2468, N1213, N410, N2279);
or OR2 (N2496, N2494, N548);
xor XOR2 (N2497, N2496, N2315);
nand NAND2 (N2498, N2493, N294);
xor XOR2 (N2499, N2482, N2085);
xor XOR2 (N2500, N2499, N573);
nand NAND3 (N2501, N2498, N1657, N1378);
not NOT1 (N2502, N2472);
or OR3 (N2503, N2501, N1074, N1673);
nand NAND3 (N2504, N2481, N279, N773);
nand NAND4 (N2505, N2504, N1568, N2191, N538);
nand NAND2 (N2506, N2488, N934);
xor XOR2 (N2507, N2503, N1490);
or OR4 (N2508, N2490, N2023, N496, N696);
nor NOR3 (N2509, N2508, N2089, N2380);
not NOT1 (N2510, N2505);
or OR3 (N2511, N2476, N725, N847);
and AND3 (N2512, N2502, N199, N1344);
endmodule