// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N8016,N8019,N8020,N8012,N8014,N8021,N8009,N7992,N8017,N8022;

nor NOR3 (N23, N21, N3, N4);
and AND3 (N24, N20, N2, N8);
or OR3 (N25, N23, N17, N21);
nor NOR3 (N26, N21, N18, N11);
or OR2 (N27, N21, N12);
not NOT1 (N28, N15);
not NOT1 (N29, N13);
xor XOR2 (N30, N25, N17);
nand NAND2 (N31, N3, N2);
xor XOR2 (N32, N17, N5);
and AND4 (N33, N11, N25, N19, N5);
or OR2 (N34, N2, N10);
nor NOR4 (N35, N34, N24, N7, N32);
xor XOR2 (N36, N33, N27);
nor NOR3 (N37, N20, N33, N30);
and AND2 (N38, N10, N29);
or OR4 (N39, N1, N2, N32, N9);
nand NAND3 (N40, N13, N36, N23);
nand NAND4 (N41, N14, N32, N40, N29);
and AND2 (N42, N31, N38);
nand NAND2 (N43, N33, N34);
nand NAND4 (N44, N10, N14, N19, N27);
nand NAND4 (N45, N26, N29, N12, N12);
nor NOR2 (N46, N2, N28);
not NOT1 (N47, N38);
and AND2 (N48, N41, N24);
not NOT1 (N49, N39);
not NOT1 (N50, N48);
or OR4 (N51, N37, N39, N28, N44);
buf BUF1 (N52, N3);
xor XOR2 (N53, N42, N16);
not NOT1 (N54, N46);
and AND3 (N55, N49, N8, N49);
buf BUF1 (N56, N55);
not NOT1 (N57, N45);
nor NOR4 (N58, N47, N48, N32, N2);
nor NOR4 (N59, N57, N20, N12, N11);
or OR2 (N60, N51, N3);
xor XOR2 (N61, N53, N13);
not NOT1 (N62, N59);
or OR2 (N63, N60, N45);
or OR3 (N64, N56, N54, N43);
xor XOR2 (N65, N37, N33);
nand NAND4 (N66, N26, N12, N2, N56);
xor XOR2 (N67, N63, N27);
and AND3 (N68, N58, N27, N19);
nor NOR3 (N69, N52, N44, N68);
nor NOR3 (N70, N42, N2, N69);
nor NOR4 (N71, N8, N70, N15, N30);
and AND2 (N72, N47, N2);
and AND2 (N73, N67, N64);
buf BUF1 (N74, N44);
nor NOR4 (N75, N65, N12, N62, N41);
not NOT1 (N76, N36);
or OR4 (N77, N61, N67, N45, N27);
or OR4 (N78, N50, N31, N15, N13);
and AND2 (N79, N74, N63);
buf BUF1 (N80, N77);
and AND3 (N81, N73, N59, N24);
nand NAND4 (N82, N76, N41, N36, N31);
not NOT1 (N83, N72);
and AND3 (N84, N79, N35, N59);
not NOT1 (N85, N42);
xor XOR2 (N86, N80, N70);
xor XOR2 (N87, N84, N61);
xor XOR2 (N88, N86, N8);
xor XOR2 (N89, N81, N28);
buf BUF1 (N90, N71);
nand NAND2 (N91, N90, N46);
nand NAND4 (N92, N66, N34, N24, N57);
nor NOR4 (N93, N91, N58, N47, N41);
nand NAND4 (N94, N83, N11, N58, N31);
xor XOR2 (N95, N87, N2);
buf BUF1 (N96, N95);
or OR2 (N97, N88, N91);
nor NOR2 (N98, N78, N87);
buf BUF1 (N99, N82);
and AND3 (N100, N85, N2, N69);
and AND4 (N101, N97, N61, N16, N29);
and AND4 (N102, N99, N67, N50, N37);
not NOT1 (N103, N75);
not NOT1 (N104, N96);
and AND3 (N105, N98, N58, N51);
xor XOR2 (N106, N92, N89);
buf BUF1 (N107, N28);
not NOT1 (N108, N105);
xor XOR2 (N109, N93, N1);
or OR4 (N110, N109, N1, N105, N100);
nor NOR3 (N111, N35, N82, N29);
nor NOR4 (N112, N108, N104, N80, N59);
or OR4 (N113, N44, N98, N34, N65);
or OR3 (N114, N111, N46, N87);
and AND4 (N115, N102, N102, N51, N92);
buf BUF1 (N116, N113);
nor NOR2 (N117, N106, N59);
or OR4 (N118, N117, N37, N66, N41);
not NOT1 (N119, N101);
nand NAND3 (N120, N114, N23, N83);
not NOT1 (N121, N120);
or OR3 (N122, N112, N69, N24);
buf BUF1 (N123, N115);
buf BUF1 (N124, N94);
and AND2 (N125, N103, N28);
buf BUF1 (N126, N119);
and AND3 (N127, N116, N72, N57);
nor NOR2 (N128, N107, N80);
nor NOR4 (N129, N123, N52, N59, N109);
and AND2 (N130, N118, N110);
or OR2 (N131, N12, N67);
xor XOR2 (N132, N130, N65);
not NOT1 (N133, N132);
xor XOR2 (N134, N131, N34);
xor XOR2 (N135, N121, N45);
xor XOR2 (N136, N134, N50);
buf BUF1 (N137, N136);
nand NAND2 (N138, N126, N42);
or OR3 (N139, N133, N79, N116);
not NOT1 (N140, N135);
xor XOR2 (N141, N122, N39);
nor NOR3 (N142, N124, N12, N127);
and AND3 (N143, N31, N96, N120);
nor NOR3 (N144, N125, N127, N86);
nor NOR3 (N145, N129, N61, N107);
not NOT1 (N146, N141);
or OR3 (N147, N145, N34, N128);
or OR2 (N148, N96, N69);
nand NAND2 (N149, N140, N127);
or OR4 (N150, N138, N36, N58, N109);
nand NAND3 (N151, N139, N68, N57);
xor XOR2 (N152, N143, N12);
and AND4 (N153, N144, N148, N132, N73);
buf BUF1 (N154, N131);
nor NOR4 (N155, N153, N107, N123, N71);
or OR4 (N156, N149, N1, N22, N110);
not NOT1 (N157, N155);
not NOT1 (N158, N146);
and AND4 (N159, N151, N87, N131, N12);
nor NOR3 (N160, N159, N81, N45);
nand NAND3 (N161, N152, N72, N142);
not NOT1 (N162, N40);
xor XOR2 (N163, N158, N144);
not NOT1 (N164, N154);
buf BUF1 (N165, N156);
not NOT1 (N166, N157);
and AND4 (N167, N150, N154, N145, N2);
buf BUF1 (N168, N164);
or OR4 (N169, N165, N28, N51, N65);
xor XOR2 (N170, N167, N96);
buf BUF1 (N171, N137);
nand NAND3 (N172, N168, N93, N54);
xor XOR2 (N173, N160, N48);
nand NAND3 (N174, N162, N171, N74);
and AND4 (N175, N42, N70, N12, N80);
nor NOR4 (N176, N173, N144, N71, N118);
not NOT1 (N177, N170);
or OR4 (N178, N177, N170, N149, N113);
xor XOR2 (N179, N163, N69);
buf BUF1 (N180, N169);
or OR3 (N181, N161, N149, N98);
and AND3 (N182, N178, N8, N141);
buf BUF1 (N183, N166);
or OR4 (N184, N182, N52, N126, N183);
xor XOR2 (N185, N23, N28);
nand NAND4 (N186, N176, N139, N49, N113);
not NOT1 (N187, N186);
xor XOR2 (N188, N172, N96);
nand NAND2 (N189, N188, N44);
xor XOR2 (N190, N180, N144);
and AND4 (N191, N147, N40, N57, N139);
and AND4 (N192, N190, N132, N137, N182);
nand NAND4 (N193, N184, N178, N118, N127);
not NOT1 (N194, N191);
buf BUF1 (N195, N179);
or OR2 (N196, N192, N45);
nand NAND3 (N197, N194, N182, N165);
nor NOR4 (N198, N187, N190, N143, N146);
xor XOR2 (N199, N198, N132);
xor XOR2 (N200, N195, N27);
buf BUF1 (N201, N199);
nor NOR3 (N202, N193, N154, N171);
or OR2 (N203, N197, N176);
nor NOR4 (N204, N201, N101, N126, N57);
or OR2 (N205, N204, N152);
or OR3 (N206, N205, N15, N167);
or OR4 (N207, N203, N48, N167, N10);
buf BUF1 (N208, N202);
nand NAND4 (N209, N196, N38, N36, N127);
or OR2 (N210, N174, N78);
nand NAND2 (N211, N210, N66);
nor NOR3 (N212, N211, N184, N147);
and AND4 (N213, N185, N106, N177, N172);
nand NAND4 (N214, N189, N62, N101, N160);
nand NAND4 (N215, N209, N210, N64, N40);
not NOT1 (N216, N200);
xor XOR2 (N217, N213, N194);
or OR3 (N218, N212, N171, N48);
or OR2 (N219, N216, N163);
nor NOR2 (N220, N175, N154);
nand NAND4 (N221, N218, N3, N36, N220);
or OR3 (N222, N134, N176, N67);
nand NAND3 (N223, N206, N42, N113);
and AND3 (N224, N214, N137, N126);
not NOT1 (N225, N181);
nand NAND2 (N226, N207, N143);
or OR2 (N227, N222, N33);
or OR3 (N228, N223, N197, N79);
or OR2 (N229, N228, N175);
and AND3 (N230, N224, N143, N33);
or OR4 (N231, N217, N36, N212, N119);
and AND3 (N232, N226, N154, N49);
and AND3 (N233, N219, N62, N159);
buf BUF1 (N234, N227);
not NOT1 (N235, N229);
xor XOR2 (N236, N234, N111);
buf BUF1 (N237, N215);
or OR2 (N238, N221, N117);
or OR4 (N239, N236, N138, N236, N30);
not NOT1 (N240, N232);
not NOT1 (N241, N230);
or OR4 (N242, N235, N42, N235, N130);
nor NOR4 (N243, N225, N65, N65, N214);
nand NAND3 (N244, N239, N10, N81);
nor NOR2 (N245, N244, N33);
nand NAND2 (N246, N245, N133);
and AND2 (N247, N238, N51);
xor XOR2 (N248, N247, N211);
not NOT1 (N249, N233);
or OR4 (N250, N241, N211, N62, N106);
or OR2 (N251, N248, N235);
xor XOR2 (N252, N240, N223);
nor NOR3 (N253, N208, N87, N29);
nor NOR3 (N254, N246, N69, N99);
not NOT1 (N255, N231);
buf BUF1 (N256, N253);
or OR4 (N257, N249, N164, N207, N61);
nor NOR4 (N258, N243, N29, N82, N184);
nand NAND3 (N259, N256, N161, N106);
not NOT1 (N260, N237);
or OR4 (N261, N252, N174, N78, N242);
and AND2 (N262, N78, N211);
nor NOR4 (N263, N258, N68, N131, N46);
nor NOR2 (N264, N262, N169);
buf BUF1 (N265, N264);
not NOT1 (N266, N259);
not NOT1 (N267, N257);
xor XOR2 (N268, N251, N207);
not NOT1 (N269, N267);
and AND3 (N270, N261, N187, N174);
xor XOR2 (N271, N269, N258);
buf BUF1 (N272, N271);
xor XOR2 (N273, N250, N258);
buf BUF1 (N274, N263);
or OR2 (N275, N255, N53);
nand NAND3 (N276, N270, N83, N43);
nor NOR3 (N277, N268, N248, N53);
or OR3 (N278, N272, N166, N203);
and AND3 (N279, N266, N82, N248);
xor XOR2 (N280, N273, N176);
not NOT1 (N281, N278);
not NOT1 (N282, N260);
or OR2 (N283, N281, N28);
and AND4 (N284, N277, N11, N41, N250);
or OR3 (N285, N283, N92, N86);
nor NOR2 (N286, N254, N243);
or OR2 (N287, N282, N265);
and AND3 (N288, N7, N141, N190);
xor XOR2 (N289, N284, N181);
or OR2 (N290, N280, N239);
xor XOR2 (N291, N287, N230);
buf BUF1 (N292, N285);
xor XOR2 (N293, N279, N101);
or OR4 (N294, N291, N53, N201, N80);
xor XOR2 (N295, N294, N114);
buf BUF1 (N296, N293);
not NOT1 (N297, N275);
xor XOR2 (N298, N274, N182);
nand NAND3 (N299, N286, N193, N22);
xor XOR2 (N300, N290, N33);
nand NAND4 (N301, N292, N5, N118, N237);
xor XOR2 (N302, N296, N171);
nor NOR4 (N303, N289, N104, N193, N268);
nand NAND4 (N304, N299, N251, N301, N31);
or OR2 (N305, N242, N149);
xor XOR2 (N306, N297, N63);
nand NAND4 (N307, N300, N118, N4, N46);
buf BUF1 (N308, N298);
xor XOR2 (N309, N306, N279);
or OR4 (N310, N308, N307, N221, N216);
or OR4 (N311, N115, N267, N172, N190);
not NOT1 (N312, N276);
and AND2 (N313, N310, N52);
buf BUF1 (N314, N313);
and AND2 (N315, N314, N131);
xor XOR2 (N316, N312, N112);
and AND4 (N317, N315, N284, N57, N154);
or OR2 (N318, N302, N49);
xor XOR2 (N319, N305, N314);
nor NOR2 (N320, N303, N140);
buf BUF1 (N321, N317);
not NOT1 (N322, N319);
or OR3 (N323, N304, N106, N107);
not NOT1 (N324, N316);
or OR4 (N325, N318, N21, N279, N192);
nor NOR3 (N326, N321, N260, N206);
nand NAND4 (N327, N324, N295, N236, N158);
buf BUF1 (N328, N49);
buf BUF1 (N329, N311);
not NOT1 (N330, N288);
nand NAND2 (N331, N328, N153);
or OR3 (N332, N327, N283, N73);
not NOT1 (N333, N309);
buf BUF1 (N334, N325);
buf BUF1 (N335, N332);
or OR2 (N336, N330, N272);
not NOT1 (N337, N320);
or OR2 (N338, N323, N66);
or OR2 (N339, N338, N219);
nand NAND2 (N340, N337, N178);
buf BUF1 (N341, N336);
nand NAND3 (N342, N341, N246, N71);
or OR2 (N343, N329, N280);
nand NAND4 (N344, N335, N282, N57, N318);
nand NAND3 (N345, N333, N327, N30);
buf BUF1 (N346, N331);
xor XOR2 (N347, N334, N143);
nand NAND4 (N348, N345, N326, N104, N285);
nor NOR3 (N349, N136, N176, N119);
nor NOR3 (N350, N340, N172, N249);
nor NOR3 (N351, N339, N344, N109);
and AND2 (N352, N294, N5);
nor NOR3 (N353, N343, N177, N206);
or OR2 (N354, N347, N305);
nor NOR4 (N355, N346, N35, N22, N151);
nand NAND4 (N356, N353, N140, N351, N346);
buf BUF1 (N357, N257);
nor NOR2 (N358, N322, N28);
not NOT1 (N359, N356);
not NOT1 (N360, N357);
not NOT1 (N361, N342);
nand NAND2 (N362, N360, N189);
nor NOR2 (N363, N362, N181);
or OR3 (N364, N359, N6, N183);
not NOT1 (N365, N348);
not NOT1 (N366, N361);
or OR4 (N367, N366, N168, N70, N351);
nor NOR4 (N368, N365, N306, N199, N138);
and AND2 (N369, N367, N311);
and AND3 (N370, N364, N261, N160);
not NOT1 (N371, N352);
nor NOR3 (N372, N358, N307, N3);
or OR4 (N373, N372, N108, N76, N252);
and AND3 (N374, N370, N59, N127);
or OR4 (N375, N369, N308, N78, N98);
not NOT1 (N376, N350);
or OR3 (N377, N355, N93, N25);
or OR3 (N378, N371, N253, N271);
xor XOR2 (N379, N373, N348);
xor XOR2 (N380, N363, N76);
nor NOR4 (N381, N376, N92, N105, N138);
buf BUF1 (N382, N379);
and AND4 (N383, N377, N220, N302, N373);
buf BUF1 (N384, N374);
not NOT1 (N385, N349);
or OR3 (N386, N375, N384, N99);
buf BUF1 (N387, N43);
not NOT1 (N388, N386);
or OR3 (N389, N382, N224, N301);
nor NOR2 (N390, N387, N289);
and AND3 (N391, N354, N138, N173);
xor XOR2 (N392, N391, N361);
or OR4 (N393, N390, N85, N246, N256);
or OR4 (N394, N381, N225, N356, N272);
nor NOR3 (N395, N383, N192, N3);
xor XOR2 (N396, N380, N173);
not NOT1 (N397, N395);
buf BUF1 (N398, N385);
and AND4 (N399, N389, N42, N331, N248);
buf BUF1 (N400, N393);
and AND4 (N401, N368, N274, N306, N224);
xor XOR2 (N402, N400, N183);
not NOT1 (N403, N397);
buf BUF1 (N404, N398);
nand NAND3 (N405, N388, N53, N302);
nand NAND3 (N406, N392, N207, N120);
nor NOR2 (N407, N404, N351);
nor NOR4 (N408, N407, N280, N135, N15);
nor NOR4 (N409, N406, N373, N275, N100);
nand NAND2 (N410, N409, N183);
buf BUF1 (N411, N402);
and AND2 (N412, N394, N104);
nor NOR2 (N413, N399, N25);
nor NOR3 (N414, N401, N36, N168);
or OR2 (N415, N403, N67);
nand NAND3 (N416, N405, N398, N176);
or OR4 (N417, N413, N167, N35, N401);
nor NOR2 (N418, N412, N3);
xor XOR2 (N419, N417, N319);
nand NAND3 (N420, N410, N56, N80);
and AND3 (N421, N378, N28, N347);
and AND2 (N422, N420, N152);
nor NOR4 (N423, N415, N83, N162, N81);
nor NOR3 (N424, N408, N340, N12);
and AND4 (N425, N396, N307, N234, N105);
nor NOR4 (N426, N422, N185, N343, N382);
or OR3 (N427, N426, N389, N320);
nand NAND3 (N428, N418, N236, N288);
or OR4 (N429, N423, N20, N119, N166);
or OR3 (N430, N428, N318, N167);
or OR3 (N431, N429, N347, N148);
and AND4 (N432, N411, N234, N76, N82);
xor XOR2 (N433, N419, N361);
buf BUF1 (N434, N424);
not NOT1 (N435, N427);
xor XOR2 (N436, N431, N384);
xor XOR2 (N437, N435, N295);
or OR4 (N438, N421, N157, N53, N46);
nor NOR3 (N439, N438, N219, N181);
nand NAND4 (N440, N439, N78, N292, N72);
nand NAND2 (N441, N416, N164);
or OR3 (N442, N433, N246, N431);
buf BUF1 (N443, N434);
buf BUF1 (N444, N442);
not NOT1 (N445, N441);
not NOT1 (N446, N443);
not NOT1 (N447, N430);
xor XOR2 (N448, N444, N129);
nand NAND2 (N449, N432, N214);
and AND3 (N450, N445, N231, N305);
or OR4 (N451, N448, N142, N398, N19);
and AND4 (N452, N414, N146, N256, N126);
nor NOR3 (N453, N436, N101, N3);
and AND3 (N454, N453, N386, N18);
xor XOR2 (N455, N440, N38);
nor NOR2 (N456, N451, N83);
nand NAND4 (N457, N454, N55, N301, N378);
not NOT1 (N458, N437);
xor XOR2 (N459, N446, N45);
or OR2 (N460, N425, N333);
buf BUF1 (N461, N456);
or OR4 (N462, N447, N444, N67, N189);
nor NOR2 (N463, N449, N456);
nand NAND3 (N464, N459, N19, N217);
buf BUF1 (N465, N461);
nand NAND2 (N466, N463, N399);
nand NAND3 (N467, N465, N232, N399);
xor XOR2 (N468, N460, N214);
nor NOR2 (N469, N466, N7);
nand NAND3 (N470, N457, N448, N46);
not NOT1 (N471, N469);
nand NAND2 (N472, N452, N437);
buf BUF1 (N473, N471);
or OR4 (N474, N468, N244, N34, N406);
nor NOR2 (N475, N450, N450);
nand NAND3 (N476, N464, N178, N168);
nand NAND4 (N477, N462, N347, N386, N220);
nor NOR2 (N478, N458, N247);
buf BUF1 (N479, N475);
xor XOR2 (N480, N470, N417);
buf BUF1 (N481, N472);
xor XOR2 (N482, N476, N89);
buf BUF1 (N483, N455);
not NOT1 (N484, N474);
not NOT1 (N485, N467);
not NOT1 (N486, N478);
nand NAND2 (N487, N486, N420);
nor NOR3 (N488, N482, N247, N392);
xor XOR2 (N489, N477, N49);
and AND3 (N490, N484, N208, N393);
xor XOR2 (N491, N485, N325);
or OR2 (N492, N473, N241);
nand NAND4 (N493, N488, N376, N40, N449);
nor NOR4 (N494, N489, N2, N430, N192);
nor NOR2 (N495, N481, N354);
xor XOR2 (N496, N490, N91);
nand NAND4 (N497, N491, N108, N133, N459);
and AND2 (N498, N494, N280);
nor NOR4 (N499, N496, N235, N423, N376);
nor NOR4 (N500, N498, N434, N375, N480);
buf BUF1 (N501, N101);
xor XOR2 (N502, N483, N56);
nand NAND2 (N503, N497, N493);
xor XOR2 (N504, N97, N371);
nand NAND3 (N505, N500, N50, N499);
or OR4 (N506, N44, N97, N472, N398);
xor XOR2 (N507, N487, N331);
nor NOR3 (N508, N495, N37, N34);
nand NAND4 (N509, N508, N434, N44, N84);
nor NOR3 (N510, N507, N152, N254);
nor NOR3 (N511, N506, N125, N183);
buf BUF1 (N512, N510);
and AND2 (N513, N505, N464);
buf BUF1 (N514, N503);
or OR2 (N515, N512, N265);
nor NOR2 (N516, N515, N78);
and AND2 (N517, N504, N486);
nand NAND2 (N518, N514, N161);
nor NOR4 (N519, N513, N38, N132, N367);
not NOT1 (N520, N501);
not NOT1 (N521, N519);
xor XOR2 (N522, N521, N245);
nor NOR2 (N523, N511, N338);
not NOT1 (N524, N523);
nand NAND2 (N525, N517, N5);
xor XOR2 (N526, N479, N149);
or OR4 (N527, N492, N285, N496, N114);
nor NOR3 (N528, N525, N270, N458);
nor NOR3 (N529, N509, N12, N141);
xor XOR2 (N530, N527, N12);
buf BUF1 (N531, N516);
xor XOR2 (N532, N524, N63);
not NOT1 (N533, N532);
nand NAND2 (N534, N502, N359);
nand NAND4 (N535, N533, N238, N90, N304);
buf BUF1 (N536, N530);
and AND3 (N537, N522, N465, N451);
buf BUF1 (N538, N535);
xor XOR2 (N539, N528, N264);
nand NAND4 (N540, N537, N65, N352, N475);
not NOT1 (N541, N518);
xor XOR2 (N542, N531, N146);
buf BUF1 (N543, N540);
and AND3 (N544, N534, N450, N156);
not NOT1 (N545, N526);
nor NOR3 (N546, N536, N144, N464);
nor NOR2 (N547, N546, N282);
or OR4 (N548, N543, N22, N336, N8);
and AND4 (N549, N539, N380, N101, N230);
not NOT1 (N550, N538);
nand NAND4 (N551, N544, N154, N366, N82);
nand NAND3 (N552, N548, N70, N322);
nand NAND4 (N553, N529, N73, N187, N297);
buf BUF1 (N554, N520);
xor XOR2 (N555, N545, N58);
nand NAND4 (N556, N542, N455, N236, N46);
or OR3 (N557, N547, N74, N303);
not NOT1 (N558, N541);
and AND3 (N559, N558, N43, N481);
not NOT1 (N560, N556);
not NOT1 (N561, N557);
nand NAND2 (N562, N551, N280);
nand NAND2 (N563, N562, N364);
buf BUF1 (N564, N561);
buf BUF1 (N565, N550);
nand NAND4 (N566, N559, N552, N392, N178);
xor XOR2 (N567, N63, N555);
nor NOR2 (N568, N297, N105);
and AND2 (N569, N549, N235);
or OR2 (N570, N568, N287);
nor NOR3 (N571, N564, N537, N418);
not NOT1 (N572, N554);
and AND4 (N573, N570, N264, N422, N487);
or OR3 (N574, N560, N251, N429);
or OR2 (N575, N553, N16);
xor XOR2 (N576, N563, N327);
and AND2 (N577, N576, N175);
nor NOR2 (N578, N572, N184);
and AND2 (N579, N569, N9);
buf BUF1 (N580, N578);
nor NOR3 (N581, N579, N305, N25);
or OR3 (N582, N574, N249, N378);
or OR2 (N583, N577, N293);
nand NAND3 (N584, N565, N434, N195);
xor XOR2 (N585, N566, N537);
not NOT1 (N586, N582);
xor XOR2 (N587, N584, N350);
buf BUF1 (N588, N573);
not NOT1 (N589, N583);
buf BUF1 (N590, N587);
buf BUF1 (N591, N571);
nand NAND2 (N592, N589, N472);
xor XOR2 (N593, N592, N572);
and AND2 (N594, N591, N283);
not NOT1 (N595, N575);
buf BUF1 (N596, N586);
not NOT1 (N597, N588);
nor NOR3 (N598, N581, N55, N391);
and AND3 (N599, N593, N112, N360);
or OR2 (N600, N585, N429);
nor NOR4 (N601, N580, N343, N417, N409);
or OR4 (N602, N597, N478, N58, N539);
xor XOR2 (N603, N602, N310);
not NOT1 (N604, N600);
or OR4 (N605, N590, N206, N265, N38);
nand NAND3 (N606, N595, N580, N141);
xor XOR2 (N607, N598, N551);
nor NOR2 (N608, N594, N120);
xor XOR2 (N609, N567, N513);
nor NOR4 (N610, N604, N385, N179, N387);
xor XOR2 (N611, N610, N415);
or OR2 (N612, N599, N205);
nor NOR4 (N613, N608, N386, N591, N95);
buf BUF1 (N614, N606);
xor XOR2 (N615, N613, N33);
buf BUF1 (N616, N615);
buf BUF1 (N617, N603);
xor XOR2 (N618, N605, N196);
not NOT1 (N619, N601);
nor NOR2 (N620, N611, N425);
nand NAND4 (N621, N596, N403, N44, N500);
not NOT1 (N622, N607);
buf BUF1 (N623, N617);
not NOT1 (N624, N619);
buf BUF1 (N625, N618);
xor XOR2 (N626, N623, N262);
xor XOR2 (N627, N625, N493);
buf BUF1 (N628, N627);
not NOT1 (N629, N614);
xor XOR2 (N630, N620, N395);
xor XOR2 (N631, N626, N341);
nor NOR4 (N632, N628, N251, N575, N223);
not NOT1 (N633, N632);
nor NOR4 (N634, N630, N537, N205, N250);
nor NOR4 (N635, N616, N622, N14, N355);
not NOT1 (N636, N22);
buf BUF1 (N637, N635);
not NOT1 (N638, N631);
and AND4 (N639, N638, N519, N124, N327);
nor NOR2 (N640, N609, N565);
buf BUF1 (N641, N633);
not NOT1 (N642, N637);
not NOT1 (N643, N624);
nor NOR4 (N644, N640, N390, N3, N246);
not NOT1 (N645, N636);
buf BUF1 (N646, N612);
or OR4 (N647, N634, N535, N645, N240);
xor XOR2 (N648, N324, N557);
xor XOR2 (N649, N647, N149);
buf BUF1 (N650, N644);
or OR4 (N651, N650, N427, N111, N289);
and AND3 (N652, N641, N565, N607);
nand NAND2 (N653, N629, N256);
nor NOR4 (N654, N646, N374, N190, N31);
nand NAND4 (N655, N651, N354, N448, N647);
and AND3 (N656, N639, N543, N39);
nand NAND2 (N657, N652, N539);
or OR2 (N658, N642, N279);
or OR4 (N659, N655, N302, N524, N492);
nor NOR3 (N660, N654, N44, N18);
and AND3 (N661, N658, N284, N513);
nor NOR3 (N662, N657, N450, N471);
and AND3 (N663, N649, N535, N331);
buf BUF1 (N664, N663);
xor XOR2 (N665, N656, N178);
nand NAND4 (N666, N664, N25, N549, N333);
nand NAND2 (N667, N666, N39);
and AND2 (N668, N643, N171);
nand NAND2 (N669, N659, N343);
not NOT1 (N670, N621);
not NOT1 (N671, N669);
or OR3 (N672, N648, N640, N166);
not NOT1 (N673, N660);
and AND4 (N674, N671, N431, N463, N536);
nand NAND4 (N675, N674, N467, N656, N571);
xor XOR2 (N676, N662, N391);
nand NAND2 (N677, N670, N73);
nand NAND3 (N678, N653, N108, N242);
nand NAND4 (N679, N675, N347, N111, N125);
buf BUF1 (N680, N679);
and AND3 (N681, N677, N153, N50);
and AND4 (N682, N667, N443, N664, N458);
nand NAND3 (N683, N681, N46, N336);
nor NOR4 (N684, N682, N26, N405, N570);
nand NAND2 (N685, N684, N71);
nand NAND2 (N686, N680, N106);
not NOT1 (N687, N678);
nand NAND4 (N688, N665, N273, N371, N590);
and AND2 (N689, N686, N460);
xor XOR2 (N690, N661, N649);
nor NOR4 (N691, N672, N76, N339, N217);
not NOT1 (N692, N685);
and AND3 (N693, N668, N646, N84);
nand NAND3 (N694, N688, N419, N332);
nor NOR2 (N695, N690, N493);
buf BUF1 (N696, N693);
nor NOR3 (N697, N673, N44, N373);
or OR4 (N698, N697, N282, N264, N537);
nand NAND4 (N699, N698, N45, N253, N258);
nor NOR2 (N700, N689, N563);
buf BUF1 (N701, N694);
xor XOR2 (N702, N683, N211);
nand NAND3 (N703, N691, N55, N631);
or OR4 (N704, N701, N699, N258, N641);
xor XOR2 (N705, N542, N429);
or OR3 (N706, N692, N444, N200);
and AND2 (N707, N705, N426);
xor XOR2 (N708, N703, N228);
nor NOR2 (N709, N706, N418);
xor XOR2 (N710, N687, N655);
xor XOR2 (N711, N696, N401);
nand NAND2 (N712, N707, N541);
not NOT1 (N713, N700);
nand NAND2 (N714, N708, N17);
not NOT1 (N715, N714);
buf BUF1 (N716, N711);
not NOT1 (N717, N702);
buf BUF1 (N718, N695);
not NOT1 (N719, N717);
nand NAND2 (N720, N704, N130);
nand NAND2 (N721, N676, N489);
nor NOR3 (N722, N709, N595, N477);
or OR4 (N723, N719, N604, N601, N510);
nand NAND4 (N724, N722, N300, N93, N723);
and AND3 (N725, N300, N433, N17);
or OR3 (N726, N713, N567, N555);
xor XOR2 (N727, N716, N298);
and AND3 (N728, N725, N638, N669);
nand NAND4 (N729, N712, N533, N567, N567);
or OR3 (N730, N710, N239, N278);
xor XOR2 (N731, N721, N623);
not NOT1 (N732, N729);
not NOT1 (N733, N718);
nor NOR3 (N734, N730, N543, N516);
xor XOR2 (N735, N732, N134);
not NOT1 (N736, N715);
not NOT1 (N737, N724);
nand NAND4 (N738, N737, N457, N107, N578);
and AND3 (N739, N734, N594, N207);
nand NAND3 (N740, N726, N411, N39);
xor XOR2 (N741, N740, N525);
and AND2 (N742, N731, N501);
xor XOR2 (N743, N739, N321);
not NOT1 (N744, N742);
nor NOR2 (N745, N743, N203);
nand NAND4 (N746, N738, N502, N409, N332);
xor XOR2 (N747, N735, N102);
and AND4 (N748, N747, N533, N430, N18);
and AND2 (N749, N744, N98);
or OR3 (N750, N733, N581, N58);
and AND2 (N751, N748, N297);
xor XOR2 (N752, N720, N373);
buf BUF1 (N753, N750);
not NOT1 (N754, N727);
buf BUF1 (N755, N745);
xor XOR2 (N756, N751, N106);
not NOT1 (N757, N746);
and AND4 (N758, N752, N263, N29, N129);
nor NOR3 (N759, N741, N513, N708);
nand NAND2 (N760, N755, N334);
nand NAND2 (N761, N753, N509);
xor XOR2 (N762, N758, N484);
nor NOR2 (N763, N728, N504);
nor NOR2 (N764, N763, N423);
not NOT1 (N765, N764);
xor XOR2 (N766, N754, N253);
or OR4 (N767, N766, N744, N54, N573);
buf BUF1 (N768, N757);
nor NOR3 (N769, N749, N619, N460);
not NOT1 (N770, N765);
or OR3 (N771, N759, N233, N3);
buf BUF1 (N772, N767);
nor NOR3 (N773, N768, N495, N127);
and AND2 (N774, N773, N595);
nand NAND4 (N775, N771, N383, N14, N463);
nand NAND2 (N776, N760, N222);
not NOT1 (N777, N772);
not NOT1 (N778, N761);
nand NAND4 (N779, N775, N56, N418, N58);
not NOT1 (N780, N777);
buf BUF1 (N781, N736);
xor XOR2 (N782, N781, N526);
or OR2 (N783, N778, N466);
nor NOR4 (N784, N774, N712, N77, N712);
not NOT1 (N785, N762);
xor XOR2 (N786, N785, N288);
buf BUF1 (N787, N783);
xor XOR2 (N788, N776, N335);
and AND3 (N789, N786, N354, N151);
not NOT1 (N790, N770);
or OR3 (N791, N779, N280, N445);
and AND2 (N792, N787, N686);
nand NAND4 (N793, N788, N179, N633, N709);
nand NAND3 (N794, N782, N762, N500);
nand NAND2 (N795, N789, N80);
xor XOR2 (N796, N792, N414);
or OR2 (N797, N793, N729);
xor XOR2 (N798, N794, N27);
and AND4 (N799, N769, N744, N477, N419);
nor NOR4 (N800, N796, N755, N750, N51);
nor NOR2 (N801, N790, N442);
buf BUF1 (N802, N797);
buf BUF1 (N803, N795);
buf BUF1 (N804, N803);
not NOT1 (N805, N799);
or OR4 (N806, N791, N444, N409, N363);
and AND4 (N807, N802, N38, N587, N675);
not NOT1 (N808, N780);
buf BUF1 (N809, N800);
xor XOR2 (N810, N798, N484);
and AND3 (N811, N804, N479, N753);
and AND2 (N812, N810, N694);
and AND2 (N813, N805, N236);
or OR3 (N814, N807, N442, N367);
nor NOR4 (N815, N813, N775, N471, N308);
not NOT1 (N816, N814);
xor XOR2 (N817, N816, N804);
nor NOR3 (N818, N811, N624, N709);
nor NOR4 (N819, N784, N813, N589, N244);
nand NAND3 (N820, N817, N506, N555);
and AND3 (N821, N806, N537, N195);
xor XOR2 (N822, N815, N685);
xor XOR2 (N823, N756, N245);
nor NOR4 (N824, N809, N807, N188, N310);
or OR3 (N825, N808, N95, N590);
not NOT1 (N826, N825);
nor NOR4 (N827, N812, N215, N145, N353);
and AND4 (N828, N822, N255, N282, N457);
and AND3 (N829, N827, N279, N59);
buf BUF1 (N830, N819);
buf BUF1 (N831, N830);
not NOT1 (N832, N831);
and AND3 (N833, N832, N153, N207);
not NOT1 (N834, N818);
not NOT1 (N835, N821);
and AND4 (N836, N834, N262, N195, N660);
buf BUF1 (N837, N828);
nand NAND2 (N838, N820, N158);
buf BUF1 (N839, N835);
nor NOR4 (N840, N837, N394, N434, N278);
not NOT1 (N841, N823);
nand NAND2 (N842, N836, N557);
and AND3 (N843, N841, N75, N823);
nor NOR2 (N844, N839, N270);
not NOT1 (N845, N840);
not NOT1 (N846, N842);
nor NOR3 (N847, N844, N651, N349);
buf BUF1 (N848, N833);
nor NOR3 (N849, N848, N227, N93);
buf BUF1 (N850, N838);
xor XOR2 (N851, N826, N801);
nand NAND2 (N852, N375, N418);
nand NAND3 (N853, N843, N440, N522);
nand NAND4 (N854, N851, N248, N523, N672);
nand NAND2 (N855, N849, N104);
nand NAND2 (N856, N850, N421);
xor XOR2 (N857, N846, N237);
nand NAND2 (N858, N829, N517);
and AND4 (N859, N845, N384, N8, N369);
and AND3 (N860, N853, N550, N290);
or OR3 (N861, N852, N410, N118);
nor NOR2 (N862, N824, N510);
nor NOR2 (N863, N847, N80);
or OR4 (N864, N862, N139, N827, N71);
nand NAND3 (N865, N858, N227, N6);
xor XOR2 (N866, N855, N250);
not NOT1 (N867, N861);
and AND4 (N868, N864, N632, N224, N635);
nand NAND3 (N869, N859, N450, N173);
or OR4 (N870, N865, N442, N751, N360);
nand NAND2 (N871, N868, N724);
not NOT1 (N872, N857);
nor NOR2 (N873, N872, N676);
nor NOR4 (N874, N854, N53, N268, N505);
xor XOR2 (N875, N856, N717);
not NOT1 (N876, N869);
buf BUF1 (N877, N871);
not NOT1 (N878, N873);
buf BUF1 (N879, N874);
or OR2 (N880, N863, N484);
xor XOR2 (N881, N877, N89);
or OR2 (N882, N870, N529);
nor NOR2 (N883, N878, N769);
buf BUF1 (N884, N867);
or OR3 (N885, N881, N460, N739);
and AND2 (N886, N879, N800);
nor NOR4 (N887, N860, N135, N417, N774);
and AND2 (N888, N880, N803);
nand NAND2 (N889, N885, N423);
or OR2 (N890, N875, N432);
buf BUF1 (N891, N886);
buf BUF1 (N892, N889);
or OR3 (N893, N883, N347, N437);
or OR3 (N894, N890, N683, N474);
not NOT1 (N895, N882);
nand NAND2 (N896, N876, N765);
not NOT1 (N897, N884);
and AND3 (N898, N896, N705, N248);
nand NAND2 (N899, N891, N796);
not NOT1 (N900, N892);
and AND3 (N901, N887, N483, N634);
not NOT1 (N902, N901);
and AND2 (N903, N894, N218);
not NOT1 (N904, N893);
buf BUF1 (N905, N866);
xor XOR2 (N906, N902, N607);
nor NOR4 (N907, N906, N483, N61, N390);
nand NAND3 (N908, N898, N130, N23);
nand NAND2 (N909, N895, N491);
xor XOR2 (N910, N904, N739);
not NOT1 (N911, N888);
not NOT1 (N912, N899);
and AND4 (N913, N909, N394, N463, N331);
and AND2 (N914, N911, N373);
nand NAND4 (N915, N912, N640, N870, N820);
or OR2 (N916, N914, N771);
nand NAND2 (N917, N910, N473);
buf BUF1 (N918, N905);
buf BUF1 (N919, N913);
and AND4 (N920, N897, N193, N539, N103);
nand NAND2 (N921, N900, N278);
buf BUF1 (N922, N920);
xor XOR2 (N923, N922, N308);
nand NAND4 (N924, N903, N389, N627, N862);
and AND4 (N925, N908, N889, N139, N716);
buf BUF1 (N926, N907);
buf BUF1 (N927, N917);
nor NOR4 (N928, N927, N719, N398, N896);
buf BUF1 (N929, N919);
nand NAND4 (N930, N926, N909, N658, N276);
or OR2 (N931, N921, N115);
xor XOR2 (N932, N915, N76);
and AND4 (N933, N923, N112, N35, N364);
nor NOR3 (N934, N924, N96, N283);
nand NAND3 (N935, N932, N122, N727);
nor NOR4 (N936, N935, N753, N357, N206);
nand NAND4 (N937, N934, N910, N694, N147);
nor NOR2 (N938, N925, N854);
nor NOR3 (N939, N937, N784, N664);
buf BUF1 (N940, N939);
not NOT1 (N941, N938);
nor NOR4 (N942, N930, N51, N498, N932);
nor NOR4 (N943, N941, N299, N81, N102);
nor NOR4 (N944, N931, N739, N799, N817);
buf BUF1 (N945, N916);
nor NOR2 (N946, N943, N69);
buf BUF1 (N947, N918);
not NOT1 (N948, N946);
not NOT1 (N949, N947);
not NOT1 (N950, N928);
or OR4 (N951, N949, N562, N203, N499);
xor XOR2 (N952, N942, N304);
buf BUF1 (N953, N933);
and AND2 (N954, N936, N676);
nand NAND4 (N955, N944, N865, N550, N339);
nand NAND2 (N956, N929, N670);
and AND2 (N957, N952, N866);
or OR2 (N958, N953, N189);
not NOT1 (N959, N958);
not NOT1 (N960, N948);
or OR2 (N961, N945, N494);
xor XOR2 (N962, N957, N437);
not NOT1 (N963, N962);
not NOT1 (N964, N963);
buf BUF1 (N965, N955);
buf BUF1 (N966, N960);
buf BUF1 (N967, N966);
xor XOR2 (N968, N967, N463);
nor NOR4 (N969, N950, N711, N819, N566);
xor XOR2 (N970, N965, N966);
not NOT1 (N971, N951);
and AND2 (N972, N969, N498);
xor XOR2 (N973, N961, N448);
or OR3 (N974, N954, N589, N780);
buf BUF1 (N975, N959);
xor XOR2 (N976, N974, N90);
or OR4 (N977, N973, N63, N720, N335);
nand NAND2 (N978, N976, N96);
nand NAND4 (N979, N964, N113, N866, N200);
xor XOR2 (N980, N977, N257);
or OR3 (N981, N940, N412, N286);
or OR4 (N982, N968, N450, N474, N864);
xor XOR2 (N983, N975, N131);
buf BUF1 (N984, N981);
nand NAND2 (N985, N956, N951);
buf BUF1 (N986, N982);
not NOT1 (N987, N970);
or OR4 (N988, N971, N766, N47, N521);
or OR3 (N989, N986, N634, N772);
nand NAND3 (N990, N980, N946, N390);
buf BUF1 (N991, N984);
or OR4 (N992, N987, N392, N300, N448);
buf BUF1 (N993, N979);
nand NAND3 (N994, N972, N924, N160);
and AND2 (N995, N994, N230);
not NOT1 (N996, N992);
and AND2 (N997, N995, N480);
and AND2 (N998, N990, N391);
and AND4 (N999, N991, N894, N930, N144);
or OR2 (N1000, N988, N718);
buf BUF1 (N1001, N997);
nor NOR3 (N1002, N1000, N954, N78);
not NOT1 (N1003, N1001);
and AND4 (N1004, N989, N272, N306, N736);
not NOT1 (N1005, N998);
not NOT1 (N1006, N985);
nor NOR2 (N1007, N996, N251);
nor NOR2 (N1008, N1005, N513);
buf BUF1 (N1009, N1006);
nor NOR2 (N1010, N1008, N731);
nand NAND3 (N1011, N1009, N131, N724);
or OR3 (N1012, N993, N98, N547);
xor XOR2 (N1013, N999, N78);
not NOT1 (N1014, N978);
nand NAND3 (N1015, N1002, N678, N873);
and AND4 (N1016, N1013, N406, N427, N157);
or OR4 (N1017, N983, N690, N577, N451);
xor XOR2 (N1018, N1011, N465);
and AND4 (N1019, N1016, N608, N481, N125);
or OR3 (N1020, N1010, N955, N499);
buf BUF1 (N1021, N1007);
or OR4 (N1022, N1015, N21, N98, N272);
or OR3 (N1023, N1003, N656, N616);
and AND4 (N1024, N1014, N276, N156, N16);
nand NAND4 (N1025, N1017, N813, N357, N681);
or OR3 (N1026, N1022, N674, N643);
nand NAND3 (N1027, N1020, N377, N261);
nand NAND4 (N1028, N1012, N722, N436, N108);
or OR2 (N1029, N1025, N60);
nand NAND3 (N1030, N1023, N307, N442);
not NOT1 (N1031, N1029);
nor NOR2 (N1032, N1021, N899);
and AND2 (N1033, N1030, N298);
nor NOR2 (N1034, N1033, N215);
and AND4 (N1035, N1026, N985, N111, N30);
xor XOR2 (N1036, N1027, N477);
and AND2 (N1037, N1034, N833);
xor XOR2 (N1038, N1036, N199);
or OR4 (N1039, N1018, N966, N865, N30);
or OR2 (N1040, N1028, N17);
not NOT1 (N1041, N1024);
buf BUF1 (N1042, N1037);
and AND3 (N1043, N1041, N156, N438);
and AND4 (N1044, N1038, N467, N226, N721);
nand NAND2 (N1045, N1040, N209);
buf BUF1 (N1046, N1035);
buf BUF1 (N1047, N1004);
nand NAND4 (N1048, N1043, N653, N651, N926);
not NOT1 (N1049, N1045);
nand NAND2 (N1050, N1044, N963);
xor XOR2 (N1051, N1042, N973);
xor XOR2 (N1052, N1051, N726);
nor NOR2 (N1053, N1050, N592);
nor NOR4 (N1054, N1048, N265, N968, N193);
nand NAND2 (N1055, N1031, N738);
or OR2 (N1056, N1053, N497);
or OR2 (N1057, N1039, N271);
and AND4 (N1058, N1032, N192, N607, N300);
nand NAND3 (N1059, N1052, N145, N435);
buf BUF1 (N1060, N1049);
not NOT1 (N1061, N1060);
and AND4 (N1062, N1047, N457, N898, N684);
nand NAND2 (N1063, N1061, N535);
not NOT1 (N1064, N1054);
not NOT1 (N1065, N1056);
xor XOR2 (N1066, N1064, N325);
nand NAND4 (N1067, N1046, N438, N143, N496);
xor XOR2 (N1068, N1062, N268);
nor NOR2 (N1069, N1066, N369);
nor NOR2 (N1070, N1019, N849);
nor NOR3 (N1071, N1058, N827, N896);
or OR2 (N1072, N1071, N1010);
nor NOR4 (N1073, N1072, N296, N977, N94);
nor NOR4 (N1074, N1055, N371, N223, N808);
nor NOR4 (N1075, N1063, N1022, N405, N875);
buf BUF1 (N1076, N1073);
nand NAND2 (N1077, N1069, N106);
buf BUF1 (N1078, N1075);
nand NAND4 (N1079, N1078, N886, N316, N151);
or OR3 (N1080, N1076, N994, N445);
nor NOR2 (N1081, N1059, N785);
buf BUF1 (N1082, N1077);
and AND4 (N1083, N1074, N576, N930, N371);
not NOT1 (N1084, N1067);
nand NAND2 (N1085, N1068, N94);
nor NOR4 (N1086, N1081, N430, N599, N449);
and AND4 (N1087, N1070, N604, N579, N113);
not NOT1 (N1088, N1080);
and AND2 (N1089, N1079, N393);
nor NOR3 (N1090, N1085, N525, N1068);
xor XOR2 (N1091, N1057, N235);
buf BUF1 (N1092, N1089);
or OR4 (N1093, N1087, N109, N422, N852);
and AND2 (N1094, N1083, N1054);
and AND3 (N1095, N1092, N1075, N14);
or OR4 (N1096, N1086, N393, N817, N1077);
nor NOR2 (N1097, N1096, N634);
or OR3 (N1098, N1097, N302, N767);
xor XOR2 (N1099, N1065, N1006);
nand NAND4 (N1100, N1091, N110, N88, N684);
xor XOR2 (N1101, N1088, N1079);
nand NAND4 (N1102, N1100, N625, N702, N793);
or OR2 (N1103, N1090, N497);
and AND3 (N1104, N1082, N39, N791);
buf BUF1 (N1105, N1101);
xor XOR2 (N1106, N1095, N1040);
not NOT1 (N1107, N1099);
and AND2 (N1108, N1106, N584);
buf BUF1 (N1109, N1107);
nand NAND4 (N1110, N1093, N199, N714, N249);
and AND3 (N1111, N1103, N1073, N671);
xor XOR2 (N1112, N1084, N639);
not NOT1 (N1113, N1094);
not NOT1 (N1114, N1104);
not NOT1 (N1115, N1108);
buf BUF1 (N1116, N1098);
not NOT1 (N1117, N1113);
and AND3 (N1118, N1115, N1060, N130);
nand NAND3 (N1119, N1117, N873, N704);
nor NOR2 (N1120, N1110, N966);
or OR2 (N1121, N1109, N79);
nand NAND4 (N1122, N1112, N185, N348, N35);
nand NAND4 (N1123, N1121, N262, N267, N1011);
not NOT1 (N1124, N1120);
not NOT1 (N1125, N1119);
buf BUF1 (N1126, N1125);
nand NAND2 (N1127, N1116, N562);
buf BUF1 (N1128, N1111);
nor NOR3 (N1129, N1128, N909, N806);
not NOT1 (N1130, N1126);
not NOT1 (N1131, N1122);
nand NAND4 (N1132, N1114, N554, N259, N137);
and AND4 (N1133, N1124, N440, N191, N911);
not NOT1 (N1134, N1129);
xor XOR2 (N1135, N1105, N483);
xor XOR2 (N1136, N1123, N141);
or OR3 (N1137, N1130, N1043, N806);
buf BUF1 (N1138, N1118);
not NOT1 (N1139, N1136);
not NOT1 (N1140, N1137);
and AND2 (N1141, N1133, N568);
or OR3 (N1142, N1127, N552, N333);
and AND2 (N1143, N1134, N24);
nand NAND4 (N1144, N1140, N410, N1055, N767);
and AND3 (N1145, N1144, N131, N813);
and AND4 (N1146, N1102, N18, N609, N3);
not NOT1 (N1147, N1146);
or OR3 (N1148, N1132, N901, N630);
nand NAND3 (N1149, N1139, N375, N430);
xor XOR2 (N1150, N1131, N1097);
nor NOR2 (N1151, N1142, N982);
nand NAND3 (N1152, N1143, N744, N507);
nand NAND2 (N1153, N1141, N432);
nand NAND4 (N1154, N1135, N748, N840, N136);
buf BUF1 (N1155, N1149);
not NOT1 (N1156, N1148);
or OR3 (N1157, N1145, N987, N175);
not NOT1 (N1158, N1155);
buf BUF1 (N1159, N1157);
not NOT1 (N1160, N1147);
nand NAND3 (N1161, N1154, N17, N248);
or OR2 (N1162, N1159, N727);
or OR4 (N1163, N1153, N111, N548, N912);
nand NAND4 (N1164, N1150, N869, N427, N818);
nand NAND3 (N1165, N1162, N541, N12);
nor NOR4 (N1166, N1160, N502, N1027, N931);
and AND4 (N1167, N1163, N193, N1074, N316);
xor XOR2 (N1168, N1167, N872);
xor XOR2 (N1169, N1156, N997);
xor XOR2 (N1170, N1151, N36);
nor NOR2 (N1171, N1158, N766);
buf BUF1 (N1172, N1170);
nand NAND4 (N1173, N1152, N374, N639, N481);
nand NAND3 (N1174, N1168, N309, N254);
nand NAND2 (N1175, N1166, N493);
xor XOR2 (N1176, N1161, N721);
not NOT1 (N1177, N1174);
and AND4 (N1178, N1138, N700, N531, N822);
not NOT1 (N1179, N1176);
nand NAND2 (N1180, N1178, N717);
or OR3 (N1181, N1179, N184, N1066);
and AND3 (N1182, N1181, N1138, N436);
nand NAND4 (N1183, N1182, N16, N591, N578);
xor XOR2 (N1184, N1171, N702);
buf BUF1 (N1185, N1164);
and AND3 (N1186, N1169, N500, N866);
xor XOR2 (N1187, N1165, N214);
and AND4 (N1188, N1183, N404, N825, N405);
buf BUF1 (N1189, N1177);
nor NOR3 (N1190, N1172, N409, N410);
nor NOR2 (N1191, N1190, N379);
not NOT1 (N1192, N1173);
xor XOR2 (N1193, N1184, N299);
xor XOR2 (N1194, N1185, N452);
or OR4 (N1195, N1186, N944, N720, N539);
nor NOR3 (N1196, N1194, N1029, N607);
buf BUF1 (N1197, N1191);
nand NAND4 (N1198, N1188, N1175, N1175, N472);
or OR3 (N1199, N354, N1182, N945);
and AND3 (N1200, N1193, N729, N529);
not NOT1 (N1201, N1200);
xor XOR2 (N1202, N1199, N1149);
xor XOR2 (N1203, N1192, N190);
nor NOR2 (N1204, N1198, N336);
buf BUF1 (N1205, N1189);
nor NOR3 (N1206, N1196, N737, N885);
and AND3 (N1207, N1197, N892, N392);
nor NOR4 (N1208, N1202, N821, N300, N909);
nand NAND4 (N1209, N1204, N277, N842, N30);
nor NOR4 (N1210, N1180, N104, N136, N1095);
nand NAND3 (N1211, N1208, N48, N1029);
not NOT1 (N1212, N1187);
nor NOR2 (N1213, N1205, N749);
buf BUF1 (N1214, N1203);
nor NOR4 (N1215, N1210, N116, N619, N1117);
nor NOR2 (N1216, N1211, N172);
not NOT1 (N1217, N1207);
nand NAND2 (N1218, N1209, N894);
or OR4 (N1219, N1217, N193, N382, N839);
or OR3 (N1220, N1201, N329, N581);
nand NAND3 (N1221, N1220, N574, N573);
xor XOR2 (N1222, N1214, N411);
nor NOR4 (N1223, N1195, N155, N535, N1077);
or OR2 (N1224, N1219, N972);
not NOT1 (N1225, N1218);
nand NAND3 (N1226, N1206, N497, N1005);
buf BUF1 (N1227, N1213);
and AND4 (N1228, N1226, N1208, N1126, N440);
buf BUF1 (N1229, N1221);
nor NOR4 (N1230, N1223, N166, N703, N581);
xor XOR2 (N1231, N1228, N155);
or OR4 (N1232, N1225, N98, N426, N485);
xor XOR2 (N1233, N1222, N823);
nand NAND3 (N1234, N1230, N175, N497);
nand NAND4 (N1235, N1227, N596, N147, N741);
xor XOR2 (N1236, N1235, N344);
xor XOR2 (N1237, N1215, N584);
not NOT1 (N1238, N1234);
or OR3 (N1239, N1229, N536, N637);
nand NAND3 (N1240, N1212, N1226, N1025);
or OR3 (N1241, N1237, N915, N435);
and AND2 (N1242, N1241, N762);
nor NOR4 (N1243, N1236, N692, N387, N620);
nor NOR3 (N1244, N1233, N1016, N315);
xor XOR2 (N1245, N1244, N653);
nor NOR2 (N1246, N1242, N337);
buf BUF1 (N1247, N1243);
and AND2 (N1248, N1238, N32);
nand NAND2 (N1249, N1247, N247);
buf BUF1 (N1250, N1248);
or OR3 (N1251, N1232, N1102, N798);
xor XOR2 (N1252, N1224, N631);
nor NOR4 (N1253, N1251, N608, N1026, N333);
not NOT1 (N1254, N1252);
or OR4 (N1255, N1249, N148, N1188, N24);
not NOT1 (N1256, N1246);
not NOT1 (N1257, N1255);
or OR4 (N1258, N1254, N806, N557, N153);
nand NAND2 (N1259, N1245, N244);
and AND3 (N1260, N1257, N324, N249);
nor NOR2 (N1261, N1253, N1255);
or OR3 (N1262, N1250, N70, N184);
or OR3 (N1263, N1231, N1178, N86);
nand NAND2 (N1264, N1259, N60);
buf BUF1 (N1265, N1260);
nor NOR2 (N1266, N1216, N809);
buf BUF1 (N1267, N1263);
or OR4 (N1268, N1258, N1175, N485, N537);
and AND2 (N1269, N1239, N805);
nand NAND2 (N1270, N1264, N375);
or OR2 (N1271, N1270, N791);
buf BUF1 (N1272, N1269);
or OR3 (N1273, N1272, N966, N1139);
nor NOR4 (N1274, N1268, N904, N148, N747);
not NOT1 (N1275, N1256);
not NOT1 (N1276, N1271);
not NOT1 (N1277, N1240);
nor NOR3 (N1278, N1276, N728, N509);
or OR4 (N1279, N1274, N1058, N913, N698);
nor NOR2 (N1280, N1273, N65);
not NOT1 (N1281, N1266);
buf BUF1 (N1282, N1280);
buf BUF1 (N1283, N1265);
or OR2 (N1284, N1267, N246);
nor NOR3 (N1285, N1284, N74, N1128);
not NOT1 (N1286, N1278);
and AND3 (N1287, N1285, N75, N21);
nor NOR2 (N1288, N1277, N502);
xor XOR2 (N1289, N1288, N457);
buf BUF1 (N1290, N1287);
xor XOR2 (N1291, N1281, N625);
and AND4 (N1292, N1262, N58, N45, N256);
or OR2 (N1293, N1289, N1229);
nand NAND4 (N1294, N1290, N613, N1290, N1066);
or OR4 (N1295, N1291, N5, N171, N301);
buf BUF1 (N1296, N1261);
xor XOR2 (N1297, N1294, N782);
not NOT1 (N1298, N1293);
buf BUF1 (N1299, N1297);
or OR4 (N1300, N1295, N1284, N210, N135);
not NOT1 (N1301, N1296);
and AND2 (N1302, N1279, N452);
xor XOR2 (N1303, N1300, N888);
and AND4 (N1304, N1282, N230, N1122, N656);
not NOT1 (N1305, N1303);
nand NAND2 (N1306, N1298, N912);
buf BUF1 (N1307, N1305);
nand NAND2 (N1308, N1302, N249);
not NOT1 (N1309, N1299);
buf BUF1 (N1310, N1306);
nand NAND3 (N1311, N1292, N789, N512);
and AND4 (N1312, N1307, N61, N339, N567);
not NOT1 (N1313, N1310);
nand NAND3 (N1314, N1309, N38, N1279);
nand NAND4 (N1315, N1301, N797, N515, N819);
not NOT1 (N1316, N1308);
nor NOR3 (N1317, N1316, N977, N28);
buf BUF1 (N1318, N1286);
nand NAND3 (N1319, N1315, N1238, N1243);
nor NOR4 (N1320, N1319, N605, N205, N631);
buf BUF1 (N1321, N1317);
and AND3 (N1322, N1314, N1033, N410);
and AND4 (N1323, N1311, N1243, N1244, N266);
or OR3 (N1324, N1318, N1037, N873);
not NOT1 (N1325, N1322);
or OR2 (N1326, N1320, N541);
buf BUF1 (N1327, N1283);
nand NAND2 (N1328, N1327, N883);
not NOT1 (N1329, N1304);
nor NOR2 (N1330, N1313, N896);
and AND2 (N1331, N1325, N953);
or OR2 (N1332, N1326, N405);
or OR4 (N1333, N1328, N62, N830, N985);
nand NAND3 (N1334, N1323, N757, N452);
nand NAND2 (N1335, N1275, N1189);
or OR3 (N1336, N1331, N507, N1247);
not NOT1 (N1337, N1336);
xor XOR2 (N1338, N1324, N1193);
and AND3 (N1339, N1312, N802, N90);
and AND3 (N1340, N1337, N915, N341);
not NOT1 (N1341, N1330);
nor NOR4 (N1342, N1340, N1043, N449, N953);
nor NOR4 (N1343, N1333, N459, N206, N686);
and AND2 (N1344, N1332, N269);
buf BUF1 (N1345, N1335);
nand NAND2 (N1346, N1345, N376);
or OR2 (N1347, N1339, N80);
nor NOR3 (N1348, N1344, N238, N709);
and AND2 (N1349, N1338, N1028);
not NOT1 (N1350, N1347);
buf BUF1 (N1351, N1334);
or OR2 (N1352, N1350, N1237);
and AND2 (N1353, N1351, N338);
xor XOR2 (N1354, N1343, N970);
buf BUF1 (N1355, N1346);
buf BUF1 (N1356, N1348);
not NOT1 (N1357, N1356);
xor XOR2 (N1358, N1355, N186);
nor NOR4 (N1359, N1354, N728, N242, N793);
nor NOR2 (N1360, N1321, N762);
not NOT1 (N1361, N1341);
nand NAND2 (N1362, N1342, N1086);
or OR3 (N1363, N1360, N197, N1260);
or OR4 (N1364, N1349, N720, N1150, N438);
xor XOR2 (N1365, N1363, N129);
not NOT1 (N1366, N1352);
not NOT1 (N1367, N1361);
xor XOR2 (N1368, N1365, N979);
buf BUF1 (N1369, N1364);
nor NOR2 (N1370, N1368, N534);
and AND3 (N1371, N1367, N862, N266);
or OR4 (N1372, N1357, N568, N591, N928);
nor NOR2 (N1373, N1366, N763);
and AND2 (N1374, N1373, N1087);
or OR2 (N1375, N1353, N385);
buf BUF1 (N1376, N1375);
nand NAND2 (N1377, N1362, N211);
or OR3 (N1378, N1376, N802, N1082);
buf BUF1 (N1379, N1359);
nor NOR4 (N1380, N1358, N644, N902, N618);
nand NAND3 (N1381, N1370, N909, N233);
nor NOR2 (N1382, N1369, N1269);
nor NOR3 (N1383, N1371, N43, N548);
xor XOR2 (N1384, N1374, N945);
xor XOR2 (N1385, N1329, N529);
buf BUF1 (N1386, N1383);
and AND4 (N1387, N1385, N786, N899, N308);
xor XOR2 (N1388, N1384, N998);
xor XOR2 (N1389, N1382, N828);
nor NOR4 (N1390, N1387, N864, N230, N235);
nand NAND2 (N1391, N1378, N940);
nor NOR3 (N1392, N1391, N823, N425);
not NOT1 (N1393, N1390);
nor NOR3 (N1394, N1392, N127, N741);
and AND3 (N1395, N1388, N428, N302);
not NOT1 (N1396, N1381);
nand NAND4 (N1397, N1380, N710, N405, N734);
nor NOR2 (N1398, N1397, N778);
nor NOR4 (N1399, N1398, N1241, N391, N353);
not NOT1 (N1400, N1386);
not NOT1 (N1401, N1372);
xor XOR2 (N1402, N1394, N1387);
buf BUF1 (N1403, N1395);
buf BUF1 (N1404, N1379);
nand NAND2 (N1405, N1401, N609);
or OR4 (N1406, N1400, N804, N1327, N728);
not NOT1 (N1407, N1406);
xor XOR2 (N1408, N1377, N1128);
not NOT1 (N1409, N1393);
and AND4 (N1410, N1399, N613, N242, N585);
not NOT1 (N1411, N1404);
or OR2 (N1412, N1409, N143);
xor XOR2 (N1413, N1410, N1005);
xor XOR2 (N1414, N1413, N999);
buf BUF1 (N1415, N1402);
xor XOR2 (N1416, N1407, N105);
buf BUF1 (N1417, N1415);
or OR4 (N1418, N1389, N957, N818, N830);
or OR4 (N1419, N1416, N813, N1373, N923);
not NOT1 (N1420, N1403);
buf BUF1 (N1421, N1414);
or OR4 (N1422, N1419, N354, N523, N617);
not NOT1 (N1423, N1422);
nor NOR2 (N1424, N1408, N594);
or OR2 (N1425, N1423, N1080);
nor NOR2 (N1426, N1418, N770);
or OR4 (N1427, N1426, N213, N1103, N1050);
and AND4 (N1428, N1411, N1137, N1099, N275);
not NOT1 (N1429, N1427);
nor NOR4 (N1430, N1429, N1098, N1053, N1209);
and AND4 (N1431, N1396, N699, N802, N765);
and AND4 (N1432, N1420, N1428, N1244, N163);
and AND4 (N1433, N1268, N843, N842, N450);
buf BUF1 (N1434, N1430);
xor XOR2 (N1435, N1421, N599);
not NOT1 (N1436, N1424);
xor XOR2 (N1437, N1431, N1069);
nand NAND3 (N1438, N1436, N339, N1434);
nor NOR2 (N1439, N946, N1124);
or OR2 (N1440, N1437, N332);
or OR2 (N1441, N1439, N537);
and AND3 (N1442, N1405, N1392, N376);
nor NOR3 (N1443, N1412, N698, N782);
xor XOR2 (N1444, N1443, N181);
and AND3 (N1445, N1432, N193, N1078);
not NOT1 (N1446, N1425);
nand NAND4 (N1447, N1417, N151, N461, N590);
nand NAND2 (N1448, N1442, N1420);
xor XOR2 (N1449, N1446, N582);
and AND2 (N1450, N1447, N897);
and AND4 (N1451, N1441, N733, N779, N512);
buf BUF1 (N1452, N1444);
nor NOR4 (N1453, N1438, N395, N753, N529);
buf BUF1 (N1454, N1452);
xor XOR2 (N1455, N1445, N1317);
and AND4 (N1456, N1451, N935, N97, N455);
or OR2 (N1457, N1454, N398);
nand NAND4 (N1458, N1440, N1088, N1385, N1065);
xor XOR2 (N1459, N1455, N1146);
and AND3 (N1460, N1435, N1058, N130);
or OR4 (N1461, N1449, N667, N573, N328);
xor XOR2 (N1462, N1459, N864);
buf BUF1 (N1463, N1462);
nand NAND3 (N1464, N1458, N674, N640);
nand NAND4 (N1465, N1464, N1153, N155, N1205);
nand NAND4 (N1466, N1463, N1393, N839, N1462);
nor NOR4 (N1467, N1466, N954, N558, N77);
and AND4 (N1468, N1456, N28, N224, N22);
nand NAND4 (N1469, N1450, N108, N548, N1079);
nor NOR2 (N1470, N1460, N1101);
buf BUF1 (N1471, N1433);
xor XOR2 (N1472, N1457, N706);
xor XOR2 (N1473, N1448, N1470);
nand NAND3 (N1474, N947, N29, N970);
and AND4 (N1475, N1471, N1404, N414, N255);
or OR3 (N1476, N1461, N493, N746);
xor XOR2 (N1477, N1473, N1282);
not NOT1 (N1478, N1467);
and AND3 (N1479, N1474, N626, N819);
buf BUF1 (N1480, N1478);
nor NOR4 (N1481, N1469, N1380, N573, N338);
nor NOR4 (N1482, N1472, N89, N267, N598);
xor XOR2 (N1483, N1481, N47);
nor NOR3 (N1484, N1479, N597, N581);
xor XOR2 (N1485, N1482, N1236);
xor XOR2 (N1486, N1480, N100);
not NOT1 (N1487, N1483);
or OR4 (N1488, N1477, N196, N1129, N530);
nor NOR3 (N1489, N1465, N52, N557);
not NOT1 (N1490, N1468);
not NOT1 (N1491, N1484);
nand NAND4 (N1492, N1487, N1306, N30, N466);
nand NAND3 (N1493, N1488, N715, N258);
nand NAND4 (N1494, N1486, N33, N907, N1396);
or OR3 (N1495, N1453, N605, N1091);
and AND2 (N1496, N1475, N454);
buf BUF1 (N1497, N1485);
nand NAND2 (N1498, N1493, N310);
nor NOR3 (N1499, N1494, N1252, N866);
not NOT1 (N1500, N1495);
nand NAND4 (N1501, N1491, N1423, N1425, N1430);
xor XOR2 (N1502, N1501, N602);
buf BUF1 (N1503, N1498);
or OR4 (N1504, N1499, N393, N572, N934);
and AND4 (N1505, N1504, N710, N1345, N966);
nand NAND4 (N1506, N1497, N480, N122, N1107);
or OR2 (N1507, N1492, N1222);
nor NOR2 (N1508, N1505, N460);
nand NAND3 (N1509, N1503, N80, N784);
nor NOR3 (N1510, N1502, N1447, N917);
nand NAND2 (N1511, N1508, N443);
nand NAND3 (N1512, N1489, N393, N1405);
or OR2 (N1513, N1507, N900);
not NOT1 (N1514, N1512);
not NOT1 (N1515, N1513);
not NOT1 (N1516, N1476);
xor XOR2 (N1517, N1506, N327);
and AND4 (N1518, N1496, N353, N353, N1188);
buf BUF1 (N1519, N1515);
nor NOR2 (N1520, N1500, N694);
not NOT1 (N1521, N1519);
and AND3 (N1522, N1517, N788, N1243);
not NOT1 (N1523, N1518);
xor XOR2 (N1524, N1510, N917);
nor NOR2 (N1525, N1509, N1084);
buf BUF1 (N1526, N1514);
or OR3 (N1527, N1490, N1118, N500);
and AND2 (N1528, N1516, N412);
and AND3 (N1529, N1524, N497, N443);
and AND2 (N1530, N1528, N1193);
nor NOR2 (N1531, N1529, N173);
buf BUF1 (N1532, N1527);
or OR4 (N1533, N1531, N1153, N598, N891);
not NOT1 (N1534, N1523);
not NOT1 (N1535, N1526);
nand NAND2 (N1536, N1534, N1288);
and AND2 (N1537, N1522, N1352);
and AND4 (N1538, N1511, N844, N890, N1208);
and AND4 (N1539, N1536, N297, N1145, N162);
xor XOR2 (N1540, N1538, N951);
nand NAND2 (N1541, N1535, N996);
xor XOR2 (N1542, N1530, N1432);
buf BUF1 (N1543, N1540);
buf BUF1 (N1544, N1525);
xor XOR2 (N1545, N1542, N838);
and AND2 (N1546, N1543, N247);
or OR3 (N1547, N1544, N337, N394);
nor NOR4 (N1548, N1537, N1490, N1353, N127);
nand NAND4 (N1549, N1521, N312, N351, N868);
not NOT1 (N1550, N1539);
or OR3 (N1551, N1533, N863, N729);
nand NAND2 (N1552, N1532, N1218);
buf BUF1 (N1553, N1541);
xor XOR2 (N1554, N1551, N810);
buf BUF1 (N1555, N1548);
xor XOR2 (N1556, N1546, N159);
not NOT1 (N1557, N1545);
not NOT1 (N1558, N1557);
buf BUF1 (N1559, N1553);
nor NOR4 (N1560, N1552, N1315, N132, N232);
or OR3 (N1561, N1547, N495, N945);
or OR2 (N1562, N1561, N347);
nand NAND4 (N1563, N1558, N1144, N446, N1200);
xor XOR2 (N1564, N1559, N136);
nor NOR2 (N1565, N1563, N1518);
xor XOR2 (N1566, N1565, N67);
not NOT1 (N1567, N1556);
buf BUF1 (N1568, N1550);
or OR3 (N1569, N1560, N895, N942);
buf BUF1 (N1570, N1564);
xor XOR2 (N1571, N1520, N210);
nor NOR2 (N1572, N1549, N1423);
nand NAND4 (N1573, N1555, N246, N342, N121);
buf BUF1 (N1574, N1566);
and AND4 (N1575, N1570, N763, N1407, N661);
and AND3 (N1576, N1571, N876, N1536);
nor NOR4 (N1577, N1576, N154, N1484, N734);
buf BUF1 (N1578, N1562);
not NOT1 (N1579, N1578);
xor XOR2 (N1580, N1574, N541);
xor XOR2 (N1581, N1567, N248);
xor XOR2 (N1582, N1568, N522);
not NOT1 (N1583, N1575);
nor NOR4 (N1584, N1579, N461, N1477, N744);
xor XOR2 (N1585, N1580, N198);
xor XOR2 (N1586, N1582, N164);
or OR2 (N1587, N1573, N1226);
not NOT1 (N1588, N1577);
and AND4 (N1589, N1572, N192, N1487, N83);
xor XOR2 (N1590, N1554, N265);
or OR3 (N1591, N1588, N114, N497);
not NOT1 (N1592, N1569);
nand NAND3 (N1593, N1589, N303, N986);
nor NOR4 (N1594, N1590, N489, N117, N1412);
xor XOR2 (N1595, N1581, N193);
or OR2 (N1596, N1592, N920);
or OR2 (N1597, N1584, N682);
xor XOR2 (N1598, N1587, N681);
xor XOR2 (N1599, N1593, N1062);
buf BUF1 (N1600, N1596);
not NOT1 (N1601, N1583);
xor XOR2 (N1602, N1600, N1027);
or OR2 (N1603, N1597, N212);
xor XOR2 (N1604, N1585, N784);
xor XOR2 (N1605, N1591, N757);
buf BUF1 (N1606, N1601);
xor XOR2 (N1607, N1604, N868);
not NOT1 (N1608, N1607);
or OR3 (N1609, N1594, N747, N449);
nor NOR2 (N1610, N1606, N183);
nand NAND2 (N1611, N1595, N425);
nor NOR3 (N1612, N1605, N597, N1592);
not NOT1 (N1613, N1611);
not NOT1 (N1614, N1612);
nor NOR4 (N1615, N1613, N372, N838, N512);
not NOT1 (N1616, N1598);
not NOT1 (N1617, N1610);
buf BUF1 (N1618, N1599);
xor XOR2 (N1619, N1586, N664);
xor XOR2 (N1620, N1617, N1578);
nor NOR4 (N1621, N1609, N1334, N1449, N172);
or OR4 (N1622, N1603, N547, N877, N341);
not NOT1 (N1623, N1621);
or OR4 (N1624, N1614, N176, N78, N436);
nand NAND2 (N1625, N1618, N1485);
or OR3 (N1626, N1623, N1372, N1170);
xor XOR2 (N1627, N1615, N1091);
not NOT1 (N1628, N1619);
and AND3 (N1629, N1620, N689, N1292);
not NOT1 (N1630, N1608);
buf BUF1 (N1631, N1616);
nor NOR2 (N1632, N1625, N437);
and AND2 (N1633, N1629, N1094);
and AND2 (N1634, N1630, N52);
nor NOR3 (N1635, N1634, N192, N104);
or OR4 (N1636, N1626, N1019, N316, N84);
or OR3 (N1637, N1636, N629, N677);
and AND2 (N1638, N1627, N1572);
xor XOR2 (N1639, N1628, N807);
or OR2 (N1640, N1635, N26);
or OR2 (N1641, N1638, N1457);
nand NAND3 (N1642, N1637, N1216, N735);
or OR2 (N1643, N1624, N1472);
and AND4 (N1644, N1639, N1101, N1215, N759);
nor NOR2 (N1645, N1642, N267);
buf BUF1 (N1646, N1640);
xor XOR2 (N1647, N1602, N1315);
buf BUF1 (N1648, N1641);
xor XOR2 (N1649, N1644, N235);
xor XOR2 (N1650, N1643, N345);
xor XOR2 (N1651, N1633, N1285);
xor XOR2 (N1652, N1648, N993);
or OR3 (N1653, N1651, N719, N830);
or OR3 (N1654, N1645, N155, N1459);
not NOT1 (N1655, N1647);
or OR4 (N1656, N1650, N130, N885, N1159);
xor XOR2 (N1657, N1646, N648);
not NOT1 (N1658, N1654);
xor XOR2 (N1659, N1653, N698);
buf BUF1 (N1660, N1649);
or OR2 (N1661, N1631, N1075);
not NOT1 (N1662, N1632);
not NOT1 (N1663, N1658);
buf BUF1 (N1664, N1622);
buf BUF1 (N1665, N1657);
xor XOR2 (N1666, N1652, N708);
nand NAND3 (N1667, N1659, N162, N422);
or OR2 (N1668, N1662, N1102);
nor NOR2 (N1669, N1664, N13);
xor XOR2 (N1670, N1669, N1383);
nand NAND3 (N1671, N1666, N472, N1499);
buf BUF1 (N1672, N1670);
nand NAND3 (N1673, N1667, N402, N15);
nor NOR3 (N1674, N1655, N1485, N1442);
nand NAND4 (N1675, N1674, N25, N1442, N251);
nand NAND2 (N1676, N1668, N250);
buf BUF1 (N1677, N1665);
nand NAND2 (N1678, N1661, N939);
nor NOR4 (N1679, N1676, N749, N215, N832);
xor XOR2 (N1680, N1656, N167);
nand NAND2 (N1681, N1660, N1567);
buf BUF1 (N1682, N1677);
nand NAND4 (N1683, N1663, N1222, N190, N946);
xor XOR2 (N1684, N1675, N422);
nand NAND2 (N1685, N1683, N1258);
not NOT1 (N1686, N1679);
not NOT1 (N1687, N1680);
not NOT1 (N1688, N1686);
or OR4 (N1689, N1671, N726, N1235, N1572);
and AND2 (N1690, N1682, N754);
not NOT1 (N1691, N1689);
nand NAND2 (N1692, N1690, N1661);
xor XOR2 (N1693, N1672, N367);
not NOT1 (N1694, N1673);
nor NOR3 (N1695, N1681, N564, N632);
buf BUF1 (N1696, N1695);
xor XOR2 (N1697, N1691, N1666);
not NOT1 (N1698, N1687);
nor NOR2 (N1699, N1696, N1101);
nor NOR4 (N1700, N1678, N491, N190, N487);
buf BUF1 (N1701, N1700);
xor XOR2 (N1702, N1699, N641);
nor NOR3 (N1703, N1693, N1318, N931);
or OR4 (N1704, N1692, N367, N290, N1291);
nand NAND4 (N1705, N1703, N1415, N638, N50);
not NOT1 (N1706, N1704);
or OR3 (N1707, N1706, N625, N1189);
not NOT1 (N1708, N1694);
not NOT1 (N1709, N1707);
or OR3 (N1710, N1698, N440, N541);
or OR4 (N1711, N1701, N1297, N759, N1088);
not NOT1 (N1712, N1697);
not NOT1 (N1713, N1708);
or OR4 (N1714, N1709, N44, N508, N976);
xor XOR2 (N1715, N1714, N832);
or OR3 (N1716, N1684, N1192, N1472);
and AND2 (N1717, N1710, N402);
nor NOR2 (N1718, N1716, N778);
and AND4 (N1719, N1711, N1341, N37, N591);
buf BUF1 (N1720, N1685);
nand NAND3 (N1721, N1720, N189, N1413);
nor NOR3 (N1722, N1719, N710, N340);
xor XOR2 (N1723, N1721, N1434);
buf BUF1 (N1724, N1713);
xor XOR2 (N1725, N1712, N948);
nand NAND3 (N1726, N1688, N983, N842);
nand NAND3 (N1727, N1724, N1625, N936);
nand NAND4 (N1728, N1725, N899, N1377, N40);
or OR4 (N1729, N1715, N36, N1452, N435);
nand NAND4 (N1730, N1718, N1247, N249, N484);
buf BUF1 (N1731, N1729);
nand NAND3 (N1732, N1730, N1159, N75);
nor NOR3 (N1733, N1731, N253, N945);
nand NAND3 (N1734, N1717, N1472, N66);
not NOT1 (N1735, N1726);
or OR2 (N1736, N1735, N153);
nor NOR4 (N1737, N1723, N1012, N383, N1577);
and AND3 (N1738, N1728, N983, N1691);
and AND3 (N1739, N1736, N1641, N1403);
or OR2 (N1740, N1733, N969);
nor NOR4 (N1741, N1734, N1131, N1469, N969);
not NOT1 (N1742, N1738);
or OR4 (N1743, N1742, N1227, N558, N607);
nor NOR2 (N1744, N1741, N1232);
buf BUF1 (N1745, N1739);
xor XOR2 (N1746, N1745, N600);
nor NOR3 (N1747, N1702, N1352, N17);
xor XOR2 (N1748, N1747, N795);
or OR3 (N1749, N1744, N1524, N1630);
xor XOR2 (N1750, N1722, N492);
and AND2 (N1751, N1732, N1432);
buf BUF1 (N1752, N1750);
nor NOR2 (N1753, N1727, N125);
xor XOR2 (N1754, N1748, N1160);
and AND2 (N1755, N1751, N165);
xor XOR2 (N1756, N1754, N1066);
or OR2 (N1757, N1705, N1653);
xor XOR2 (N1758, N1746, N1217);
buf BUF1 (N1759, N1757);
and AND3 (N1760, N1753, N1725, N1448);
nand NAND4 (N1761, N1749, N1593, N194, N669);
xor XOR2 (N1762, N1758, N671);
buf BUF1 (N1763, N1756);
and AND4 (N1764, N1763, N855, N194, N985);
xor XOR2 (N1765, N1743, N742);
not NOT1 (N1766, N1762);
and AND3 (N1767, N1760, N1685, N1436);
and AND3 (N1768, N1767, N1586, N334);
and AND2 (N1769, N1764, N400);
nand NAND4 (N1770, N1737, N575, N1761, N1009);
nor NOR2 (N1771, N854, N1470);
xor XOR2 (N1772, N1768, N62);
not NOT1 (N1773, N1771);
not NOT1 (N1774, N1770);
xor XOR2 (N1775, N1773, N1177);
and AND2 (N1776, N1775, N666);
xor XOR2 (N1777, N1766, N683);
buf BUF1 (N1778, N1752);
not NOT1 (N1779, N1769);
and AND4 (N1780, N1759, N224, N1426, N1529);
nand NAND2 (N1781, N1755, N69);
or OR3 (N1782, N1765, N1468, N1073);
nor NOR4 (N1783, N1776, N759, N1451, N974);
nand NAND4 (N1784, N1781, N49, N1468, N1180);
nor NOR3 (N1785, N1784, N496, N597);
buf BUF1 (N1786, N1783);
xor XOR2 (N1787, N1740, N1123);
or OR4 (N1788, N1782, N105, N1516, N1208);
xor XOR2 (N1789, N1772, N725);
nor NOR3 (N1790, N1788, N1425, N441);
not NOT1 (N1791, N1789);
not NOT1 (N1792, N1787);
nor NOR2 (N1793, N1779, N1758);
not NOT1 (N1794, N1780);
buf BUF1 (N1795, N1793);
nand NAND4 (N1796, N1795, N180, N979, N1615);
not NOT1 (N1797, N1790);
nor NOR2 (N1798, N1792, N282);
buf BUF1 (N1799, N1774);
and AND2 (N1800, N1799, N1683);
xor XOR2 (N1801, N1798, N1551);
and AND2 (N1802, N1797, N192);
or OR2 (N1803, N1800, N1776);
nand NAND3 (N1804, N1801, N744, N439);
nand NAND3 (N1805, N1791, N143, N1097);
buf BUF1 (N1806, N1778);
buf BUF1 (N1807, N1796);
xor XOR2 (N1808, N1785, N1022);
and AND2 (N1809, N1807, N582);
or OR2 (N1810, N1805, N323);
xor XOR2 (N1811, N1803, N694);
buf BUF1 (N1812, N1786);
nand NAND2 (N1813, N1806, N1209);
nand NAND4 (N1814, N1808, N1409, N1351, N155);
buf BUF1 (N1815, N1810);
xor XOR2 (N1816, N1814, N1470);
nor NOR4 (N1817, N1816, N1781, N1159, N623);
nor NOR4 (N1818, N1809, N15, N278, N1273);
or OR4 (N1819, N1812, N250, N1684, N609);
not NOT1 (N1820, N1804);
or OR4 (N1821, N1794, N925, N822, N420);
xor XOR2 (N1822, N1811, N1055);
not NOT1 (N1823, N1821);
or OR3 (N1824, N1777, N1362, N1510);
or OR2 (N1825, N1802, N948);
or OR3 (N1826, N1819, N658, N822);
not NOT1 (N1827, N1823);
and AND3 (N1828, N1827, N1476, N1136);
nand NAND4 (N1829, N1820, N208, N725, N1512);
buf BUF1 (N1830, N1822);
nand NAND3 (N1831, N1825, N79, N333);
or OR4 (N1832, N1831, N1046, N85, N691);
nor NOR4 (N1833, N1829, N1621, N1501, N816);
or OR2 (N1834, N1815, N1396);
nand NAND2 (N1835, N1813, N438);
or OR2 (N1836, N1818, N1467);
and AND3 (N1837, N1817, N311, N692);
and AND4 (N1838, N1833, N1537, N11, N1484);
xor XOR2 (N1839, N1828, N473);
nor NOR4 (N1840, N1832, N1826, N1227, N172);
buf BUF1 (N1841, N1042);
nand NAND4 (N1842, N1837, N1818, N43, N825);
not NOT1 (N1843, N1835);
xor XOR2 (N1844, N1824, N466);
buf BUF1 (N1845, N1839);
buf BUF1 (N1846, N1844);
and AND2 (N1847, N1841, N899);
buf BUF1 (N1848, N1842);
or OR2 (N1849, N1840, N134);
not NOT1 (N1850, N1834);
nor NOR2 (N1851, N1838, N1456);
nor NOR3 (N1852, N1846, N1520, N1512);
buf BUF1 (N1853, N1849);
and AND3 (N1854, N1836, N1237, N156);
or OR2 (N1855, N1851, N651);
nor NOR4 (N1856, N1855, N1602, N169, N1463);
buf BUF1 (N1857, N1847);
not NOT1 (N1858, N1830);
or OR3 (N1859, N1856, N1449, N779);
nor NOR3 (N1860, N1858, N135, N1081);
nor NOR3 (N1861, N1859, N497, N1343);
nand NAND3 (N1862, N1845, N342, N1249);
or OR2 (N1863, N1850, N533);
nand NAND2 (N1864, N1852, N447);
nor NOR2 (N1865, N1860, N1155);
not NOT1 (N1866, N1848);
buf BUF1 (N1867, N1843);
xor XOR2 (N1868, N1853, N1319);
and AND4 (N1869, N1862, N746, N22, N1135);
nand NAND2 (N1870, N1869, N1044);
buf BUF1 (N1871, N1865);
and AND2 (N1872, N1864, N1142);
nand NAND3 (N1873, N1857, N699, N199);
or OR2 (N1874, N1873, N569);
or OR3 (N1875, N1874, N1110, N1708);
nor NOR4 (N1876, N1867, N1159, N1261, N673);
and AND2 (N1877, N1854, N1236);
buf BUF1 (N1878, N1863);
xor XOR2 (N1879, N1868, N1209);
xor XOR2 (N1880, N1876, N1074);
nor NOR3 (N1881, N1871, N924, N846);
not NOT1 (N1882, N1879);
or OR4 (N1883, N1880, N600, N1717, N1108);
buf BUF1 (N1884, N1861);
buf BUF1 (N1885, N1875);
nand NAND2 (N1886, N1883, N1674);
or OR3 (N1887, N1885, N1496, N375);
and AND3 (N1888, N1872, N1872, N409);
and AND2 (N1889, N1882, N817);
nor NOR3 (N1890, N1877, N646, N1779);
xor XOR2 (N1891, N1870, N634);
xor XOR2 (N1892, N1888, N1007);
nor NOR3 (N1893, N1884, N1024, N719);
not NOT1 (N1894, N1893);
not NOT1 (N1895, N1886);
nand NAND2 (N1896, N1878, N845);
nand NAND2 (N1897, N1887, N1775);
nand NAND4 (N1898, N1891, N471, N1010, N1154);
and AND3 (N1899, N1894, N93, N590);
not NOT1 (N1900, N1898);
or OR2 (N1901, N1900, N243);
nor NOR3 (N1902, N1890, N1662, N372);
and AND3 (N1903, N1866, N1852, N1319);
not NOT1 (N1904, N1889);
not NOT1 (N1905, N1897);
xor XOR2 (N1906, N1899, N888);
nand NAND2 (N1907, N1904, N1543);
buf BUF1 (N1908, N1902);
not NOT1 (N1909, N1901);
buf BUF1 (N1910, N1905);
and AND2 (N1911, N1892, N1528);
nor NOR3 (N1912, N1911, N1516, N561);
not NOT1 (N1913, N1909);
xor XOR2 (N1914, N1906, N858);
and AND4 (N1915, N1910, N922, N1737, N1785);
and AND2 (N1916, N1903, N1671);
not NOT1 (N1917, N1914);
not NOT1 (N1918, N1881);
xor XOR2 (N1919, N1907, N303);
or OR2 (N1920, N1913, N948);
or OR3 (N1921, N1908, N37, N1162);
nor NOR2 (N1922, N1917, N546);
not NOT1 (N1923, N1919);
not NOT1 (N1924, N1915);
buf BUF1 (N1925, N1924);
not NOT1 (N1926, N1925);
or OR2 (N1927, N1912, N771);
xor XOR2 (N1928, N1895, N737);
xor XOR2 (N1929, N1922, N1458);
nor NOR2 (N1930, N1923, N1593);
xor XOR2 (N1931, N1928, N1481);
and AND4 (N1932, N1931, N689, N1761, N1036);
not NOT1 (N1933, N1932);
or OR2 (N1934, N1920, N689);
not NOT1 (N1935, N1896);
not NOT1 (N1936, N1930);
xor XOR2 (N1937, N1927, N1887);
not NOT1 (N1938, N1934);
xor XOR2 (N1939, N1929, N315);
or OR3 (N1940, N1937, N1756, N911);
not NOT1 (N1941, N1938);
not NOT1 (N1942, N1940);
xor XOR2 (N1943, N1926, N226);
not NOT1 (N1944, N1921);
and AND3 (N1945, N1933, N1245, N764);
and AND3 (N1946, N1939, N1416, N242);
buf BUF1 (N1947, N1941);
or OR2 (N1948, N1918, N555);
xor XOR2 (N1949, N1935, N970);
or OR2 (N1950, N1916, N1102);
nor NOR2 (N1951, N1936, N1281);
buf BUF1 (N1952, N1942);
nand NAND4 (N1953, N1946, N504, N606, N1053);
and AND4 (N1954, N1943, N439, N74, N653);
nor NOR4 (N1955, N1951, N1107, N966, N349);
or OR2 (N1956, N1954, N1091);
not NOT1 (N1957, N1956);
not NOT1 (N1958, N1950);
nand NAND4 (N1959, N1958, N535, N679, N383);
not NOT1 (N1960, N1947);
nor NOR2 (N1961, N1945, N707);
xor XOR2 (N1962, N1961, N1716);
and AND3 (N1963, N1962, N1089, N1437);
not NOT1 (N1964, N1960);
or OR2 (N1965, N1953, N29);
not NOT1 (N1966, N1955);
nor NOR2 (N1967, N1965, N668);
nand NAND3 (N1968, N1966, N1626, N1148);
nand NAND3 (N1969, N1968, N1201, N797);
xor XOR2 (N1970, N1944, N1958);
and AND4 (N1971, N1949, N246, N1256, N802);
not NOT1 (N1972, N1952);
or OR3 (N1973, N1969, N1404, N1049);
xor XOR2 (N1974, N1957, N411);
nand NAND2 (N1975, N1948, N228);
buf BUF1 (N1976, N1972);
buf BUF1 (N1977, N1967);
buf BUF1 (N1978, N1959);
nor NOR2 (N1979, N1978, N591);
nand NAND3 (N1980, N1979, N285, N509);
and AND3 (N1981, N1977, N1178, N1517);
buf BUF1 (N1982, N1976);
not NOT1 (N1983, N1975);
not NOT1 (N1984, N1964);
buf BUF1 (N1985, N1983);
nand NAND3 (N1986, N1974, N1366, N564);
not NOT1 (N1987, N1963);
xor XOR2 (N1988, N1987, N1984);
nand NAND3 (N1989, N482, N33, N105);
nand NAND4 (N1990, N1989, N756, N470, N1957);
nand NAND4 (N1991, N1981, N1511, N1439, N227);
and AND4 (N1992, N1971, N476, N1241, N1563);
or OR3 (N1993, N1992, N14, N916);
nand NAND3 (N1994, N1988, N1328, N1878);
or OR3 (N1995, N1994, N302, N122);
and AND3 (N1996, N1982, N199, N686);
not NOT1 (N1997, N1986);
not NOT1 (N1998, N1996);
buf BUF1 (N1999, N1985);
buf BUF1 (N2000, N1970);
and AND3 (N2001, N1997, N925, N1723);
and AND2 (N2002, N1990, N501);
not NOT1 (N2003, N2000);
and AND2 (N2004, N1993, N1540);
nand NAND2 (N2005, N2002, N1344);
not NOT1 (N2006, N1991);
and AND3 (N2007, N1998, N1315, N1543);
and AND4 (N2008, N2001, N1669, N884, N243);
not NOT1 (N2009, N2008);
or OR2 (N2010, N2006, N555);
buf BUF1 (N2011, N1973);
xor XOR2 (N2012, N2005, N1064);
buf BUF1 (N2013, N2009);
xor XOR2 (N2014, N2012, N245);
nor NOR3 (N2015, N2003, N1421, N1418);
nand NAND2 (N2016, N2015, N1349);
and AND3 (N2017, N2010, N1880, N317);
nand NAND4 (N2018, N1980, N571, N224, N826);
not NOT1 (N2019, N2004);
xor XOR2 (N2020, N2017, N611);
nor NOR4 (N2021, N2011, N171, N450, N1778);
and AND4 (N2022, N2019, N1476, N1484, N1365);
nor NOR4 (N2023, N1999, N851, N1233, N1567);
nor NOR3 (N2024, N2007, N573, N1450);
or OR2 (N2025, N2016, N635);
xor XOR2 (N2026, N2013, N440);
not NOT1 (N2027, N2026);
xor XOR2 (N2028, N1995, N1202);
or OR2 (N2029, N2028, N1706);
xor XOR2 (N2030, N2021, N1069);
nor NOR4 (N2031, N2023, N248, N25, N728);
buf BUF1 (N2032, N2024);
nor NOR3 (N2033, N2032, N474, N749);
buf BUF1 (N2034, N2030);
not NOT1 (N2035, N2031);
nor NOR4 (N2036, N2034, N1225, N136, N584);
buf BUF1 (N2037, N2035);
not NOT1 (N2038, N2037);
and AND2 (N2039, N2018, N86);
nor NOR4 (N2040, N2039, N1344, N188, N4);
or OR3 (N2041, N2029, N874, N408);
buf BUF1 (N2042, N2020);
not NOT1 (N2043, N2040);
or OR4 (N2044, N2042, N68, N1325, N1180);
not NOT1 (N2045, N2043);
not NOT1 (N2046, N2025);
and AND2 (N2047, N2041, N875);
nand NAND4 (N2048, N2027, N2032, N91, N1361);
not NOT1 (N2049, N2014);
and AND3 (N2050, N2033, N1812, N35);
not NOT1 (N2051, N2038);
and AND2 (N2052, N2049, N1991);
or OR2 (N2053, N2052, N631);
nor NOR3 (N2054, N2053, N12, N199);
buf BUF1 (N2055, N2048);
not NOT1 (N2056, N2054);
buf BUF1 (N2057, N2047);
nand NAND2 (N2058, N2022, N1921);
nand NAND4 (N2059, N2044, N862, N865, N1193);
nor NOR4 (N2060, N2055, N1126, N52, N1469);
buf BUF1 (N2061, N2056);
nand NAND4 (N2062, N2045, N1037, N236, N1877);
and AND3 (N2063, N2057, N1462, N853);
or OR4 (N2064, N2061, N960, N1668, N1595);
not NOT1 (N2065, N2063);
and AND2 (N2066, N2062, N2064);
or OR2 (N2067, N1609, N1989);
or OR3 (N2068, N2058, N1708, N152);
nor NOR2 (N2069, N2036, N476);
or OR2 (N2070, N2067, N1383);
nor NOR3 (N2071, N2060, N1976, N1823);
nand NAND2 (N2072, N2046, N442);
not NOT1 (N2073, N2068);
xor XOR2 (N2074, N2072, N367);
xor XOR2 (N2075, N2059, N834);
xor XOR2 (N2076, N2075, N335);
and AND2 (N2077, N2076, N24);
not NOT1 (N2078, N2051);
and AND2 (N2079, N2073, N481);
nand NAND4 (N2080, N2077, N320, N500, N1709);
or OR4 (N2081, N2070, N1750, N325, N761);
not NOT1 (N2082, N2066);
xor XOR2 (N2083, N2082, N1550);
or OR3 (N2084, N2079, N867, N1612);
buf BUF1 (N2085, N2078);
nand NAND3 (N2086, N2069, N833, N782);
and AND4 (N2087, N2085, N328, N1893, N1526);
nor NOR4 (N2088, N2080, N380, N491, N1341);
or OR3 (N2089, N2083, N56, N22);
and AND3 (N2090, N2081, N1881, N1567);
nor NOR3 (N2091, N2087, N827, N1589);
not NOT1 (N2092, N2090);
not NOT1 (N2093, N2050);
not NOT1 (N2094, N2093);
nand NAND2 (N2095, N2088, N1796);
xor XOR2 (N2096, N2084, N1137);
nand NAND3 (N2097, N2091, N14, N357);
xor XOR2 (N2098, N2092, N478);
nor NOR2 (N2099, N2097, N1080);
nor NOR2 (N2100, N2065, N1344);
nand NAND4 (N2101, N2096, N570, N1693, N1608);
not NOT1 (N2102, N2101);
nand NAND2 (N2103, N2094, N1727);
and AND4 (N2104, N2086, N1069, N223, N885);
and AND4 (N2105, N2071, N151, N1593, N236);
not NOT1 (N2106, N2095);
or OR2 (N2107, N2102, N1936);
xor XOR2 (N2108, N2100, N1416);
nor NOR2 (N2109, N2107, N1105);
nand NAND4 (N2110, N2105, N1429, N597, N666);
and AND4 (N2111, N2099, N781, N1289, N1846);
not NOT1 (N2112, N2106);
nand NAND2 (N2113, N2074, N1550);
not NOT1 (N2114, N2112);
xor XOR2 (N2115, N2109, N1334);
nand NAND3 (N2116, N2104, N2016, N87);
or OR2 (N2117, N2113, N224);
xor XOR2 (N2118, N2115, N764);
xor XOR2 (N2119, N2103, N865);
and AND2 (N2120, N2119, N805);
buf BUF1 (N2121, N2111);
buf BUF1 (N2122, N2120);
nor NOR3 (N2123, N2116, N936, N179);
nand NAND2 (N2124, N2110, N1662);
or OR4 (N2125, N2118, N860, N1586, N453);
nor NOR3 (N2126, N2122, N417, N1210);
nand NAND4 (N2127, N2121, N1562, N293, N1546);
xor XOR2 (N2128, N2098, N1495);
not NOT1 (N2129, N2127);
buf BUF1 (N2130, N2089);
and AND4 (N2131, N2124, N1442, N312, N929);
nor NOR4 (N2132, N2123, N1660, N467, N2087);
and AND2 (N2133, N2129, N877);
and AND4 (N2134, N2131, N1473, N173, N736);
nor NOR2 (N2135, N2128, N1799);
nand NAND4 (N2136, N2134, N1766, N1648, N1814);
buf BUF1 (N2137, N2135);
nand NAND4 (N2138, N2117, N158, N345, N1000);
or OR2 (N2139, N2132, N1706);
xor XOR2 (N2140, N2136, N680);
xor XOR2 (N2141, N2126, N1901);
and AND4 (N2142, N2138, N1623, N746, N1476);
or OR2 (N2143, N2108, N1526);
buf BUF1 (N2144, N2133);
nor NOR4 (N2145, N2141, N231, N220, N1493);
or OR4 (N2146, N2145, N1331, N1942, N1786);
nand NAND4 (N2147, N2143, N259, N1317, N1571);
xor XOR2 (N2148, N2142, N780);
xor XOR2 (N2149, N2146, N1009);
and AND2 (N2150, N2137, N1272);
nand NAND2 (N2151, N2149, N109);
xor XOR2 (N2152, N2144, N1621);
nand NAND3 (N2153, N2125, N884, N702);
buf BUF1 (N2154, N2153);
nor NOR4 (N2155, N2140, N1100, N712, N1109);
and AND4 (N2156, N2130, N1019, N216, N1847);
not NOT1 (N2157, N2150);
not NOT1 (N2158, N2152);
nor NOR3 (N2159, N2154, N436, N514);
nand NAND2 (N2160, N2159, N291);
not NOT1 (N2161, N2139);
and AND2 (N2162, N2155, N1466);
not NOT1 (N2163, N2148);
not NOT1 (N2164, N2162);
or OR4 (N2165, N2156, N758, N48, N278);
xor XOR2 (N2166, N2165, N304);
nand NAND2 (N2167, N2151, N1550);
or OR3 (N2168, N2164, N135, N253);
and AND3 (N2169, N2114, N1827, N253);
not NOT1 (N2170, N2167);
buf BUF1 (N2171, N2170);
nor NOR2 (N2172, N2169, N1719);
buf BUF1 (N2173, N2157);
and AND4 (N2174, N2166, N129, N1840, N392);
not NOT1 (N2175, N2174);
nor NOR3 (N2176, N2168, N487, N1174);
buf BUF1 (N2177, N2176);
xor XOR2 (N2178, N2158, N910);
nor NOR3 (N2179, N2175, N2064, N924);
nand NAND2 (N2180, N2177, N1622);
and AND3 (N2181, N2179, N1254, N935);
nand NAND4 (N2182, N2173, N1531, N1262, N1939);
and AND4 (N2183, N2182, N386, N1754, N1735);
xor XOR2 (N2184, N2172, N1430);
and AND4 (N2185, N2147, N603, N1035, N1740);
or OR3 (N2186, N2181, N1067, N1072);
nand NAND4 (N2187, N2171, N720, N1192, N435);
and AND3 (N2188, N2163, N1477, N1198);
or OR2 (N2189, N2184, N715);
nor NOR4 (N2190, N2178, N1009, N1564, N2081);
not NOT1 (N2191, N2160);
buf BUF1 (N2192, N2185);
and AND2 (N2193, N2161, N470);
buf BUF1 (N2194, N2180);
or OR2 (N2195, N2192, N1039);
and AND2 (N2196, N2183, N1612);
or OR3 (N2197, N2194, N1844, N1266);
nand NAND2 (N2198, N2195, N85);
and AND3 (N2199, N2187, N2086, N1865);
buf BUF1 (N2200, N2190);
nand NAND2 (N2201, N2191, N1101);
and AND4 (N2202, N2188, N800, N220, N634);
nand NAND2 (N2203, N2186, N2053);
xor XOR2 (N2204, N2199, N1428);
nor NOR2 (N2205, N2204, N1918);
not NOT1 (N2206, N2205);
nand NAND4 (N2207, N2202, N2167, N1620, N832);
nor NOR2 (N2208, N2207, N660);
not NOT1 (N2209, N2193);
buf BUF1 (N2210, N2196);
nand NAND3 (N2211, N2201, N1235, N459);
nand NAND4 (N2212, N2211, N156, N1958, N888);
not NOT1 (N2213, N2200);
or OR2 (N2214, N2209, N169);
buf BUF1 (N2215, N2197);
xor XOR2 (N2216, N2189, N1269);
xor XOR2 (N2217, N2206, N1297);
and AND4 (N2218, N2215, N1438, N647, N2205);
and AND4 (N2219, N2217, N1016, N412, N330);
xor XOR2 (N2220, N2219, N1299);
buf BUF1 (N2221, N2218);
nand NAND2 (N2222, N2220, N880);
nand NAND4 (N2223, N2208, N345, N2015, N331);
or OR4 (N2224, N2221, N1790, N892, N1638);
not NOT1 (N2225, N2224);
buf BUF1 (N2226, N2216);
and AND3 (N2227, N2210, N792, N948);
xor XOR2 (N2228, N2222, N476);
nand NAND3 (N2229, N2223, N923, N731);
xor XOR2 (N2230, N2214, N145);
or OR4 (N2231, N2228, N1117, N1899, N2059);
nor NOR2 (N2232, N2231, N1671);
or OR4 (N2233, N2227, N1382, N1828, N781);
nand NAND4 (N2234, N2233, N1809, N510, N523);
nand NAND3 (N2235, N2226, N305, N302);
nand NAND2 (N2236, N2229, N406);
xor XOR2 (N2237, N2225, N1347);
not NOT1 (N2238, N2237);
or OR3 (N2239, N2198, N1565, N1325);
xor XOR2 (N2240, N2232, N1772);
nor NOR4 (N2241, N2235, N2052, N352, N1725);
xor XOR2 (N2242, N2234, N178);
buf BUF1 (N2243, N2238);
or OR2 (N2244, N2203, N1547);
buf BUF1 (N2245, N2240);
or OR4 (N2246, N2239, N483, N207, N1110);
buf BUF1 (N2247, N2212);
not NOT1 (N2248, N2246);
nor NOR2 (N2249, N2236, N516);
xor XOR2 (N2250, N2244, N1560);
nor NOR2 (N2251, N2248, N1789);
and AND4 (N2252, N2250, N1512, N482, N200);
xor XOR2 (N2253, N2251, N984);
or OR4 (N2254, N2252, N542, N1610, N517);
not NOT1 (N2255, N2213);
buf BUF1 (N2256, N2247);
and AND3 (N2257, N2242, N551, N944);
or OR4 (N2258, N2230, N469, N575, N1173);
or OR4 (N2259, N2245, N820, N1941, N133);
buf BUF1 (N2260, N2243);
and AND4 (N2261, N2249, N995, N1742, N2249);
xor XOR2 (N2262, N2261, N840);
or OR3 (N2263, N2258, N2198, N787);
or OR3 (N2264, N2256, N1757, N1420);
buf BUF1 (N2265, N2260);
or OR4 (N2266, N2265, N1834, N696, N1399);
xor XOR2 (N2267, N2266, N66);
buf BUF1 (N2268, N2267);
buf BUF1 (N2269, N2263);
not NOT1 (N2270, N2254);
nor NOR4 (N2271, N2264, N1309, N1852, N2122);
nor NOR4 (N2272, N2259, N1107, N1824, N647);
not NOT1 (N2273, N2268);
buf BUF1 (N2274, N2269);
not NOT1 (N2275, N2271);
buf BUF1 (N2276, N2273);
not NOT1 (N2277, N2253);
not NOT1 (N2278, N2255);
nand NAND2 (N2279, N2262, N1142);
nand NAND3 (N2280, N2275, N340, N1973);
buf BUF1 (N2281, N2279);
xor XOR2 (N2282, N2257, N664);
and AND4 (N2283, N2278, N2154, N507, N1363);
xor XOR2 (N2284, N2272, N937);
not NOT1 (N2285, N2280);
and AND4 (N2286, N2270, N1874, N891, N74);
buf BUF1 (N2287, N2277);
and AND3 (N2288, N2282, N294, N1945);
xor XOR2 (N2289, N2283, N2121);
buf BUF1 (N2290, N2288);
buf BUF1 (N2291, N2289);
or OR2 (N2292, N2276, N211);
xor XOR2 (N2293, N2292, N807);
nand NAND3 (N2294, N2274, N729, N2290);
or OR2 (N2295, N503, N1044);
or OR4 (N2296, N2295, N1399, N200, N1408);
buf BUF1 (N2297, N2294);
nand NAND4 (N2298, N2241, N986, N152, N2193);
xor XOR2 (N2299, N2291, N1610);
not NOT1 (N2300, N2287);
and AND2 (N2301, N2300, N1715);
xor XOR2 (N2302, N2299, N1953);
xor XOR2 (N2303, N2296, N1065);
or OR3 (N2304, N2285, N1498, N1881);
nand NAND2 (N2305, N2297, N869);
xor XOR2 (N2306, N2281, N2199);
buf BUF1 (N2307, N2284);
nand NAND3 (N2308, N2302, N56, N172);
and AND4 (N2309, N2286, N903, N672, N1622);
nor NOR4 (N2310, N2293, N964, N1013, N666);
and AND4 (N2311, N2298, N282, N681, N713);
buf BUF1 (N2312, N2310);
or OR4 (N2313, N2304, N721, N1904, N378);
buf BUF1 (N2314, N2307);
nand NAND2 (N2315, N2313, N1612);
and AND4 (N2316, N2306, N141, N1889, N216);
and AND2 (N2317, N2303, N728);
nor NOR4 (N2318, N2316, N631, N1847, N1192);
nand NAND4 (N2319, N2301, N1588, N216, N203);
and AND3 (N2320, N2308, N451, N559);
nor NOR3 (N2321, N2305, N631, N448);
nor NOR3 (N2322, N2311, N1587, N2299);
xor XOR2 (N2323, N2317, N1688);
buf BUF1 (N2324, N2315);
and AND2 (N2325, N2324, N288);
or OR3 (N2326, N2321, N464, N1848);
not NOT1 (N2327, N2320);
nand NAND2 (N2328, N2327, N1147);
not NOT1 (N2329, N2328);
nor NOR4 (N2330, N2309, N2000, N843, N418);
or OR3 (N2331, N2329, N1368, N1176);
buf BUF1 (N2332, N2330);
xor XOR2 (N2333, N2326, N348);
not NOT1 (N2334, N2325);
or OR4 (N2335, N2322, N1172, N1232, N1423);
or OR2 (N2336, N2335, N260);
buf BUF1 (N2337, N2333);
nor NOR4 (N2338, N2336, N489, N523, N293);
nand NAND4 (N2339, N2332, N591, N2072, N1367);
buf BUF1 (N2340, N2334);
nor NOR4 (N2341, N2338, N2325, N2074, N1565);
xor XOR2 (N2342, N2341, N1843);
buf BUF1 (N2343, N2314);
nor NOR2 (N2344, N2342, N2261);
buf BUF1 (N2345, N2323);
xor XOR2 (N2346, N2319, N2043);
nor NOR2 (N2347, N2343, N147);
nor NOR3 (N2348, N2331, N1360, N623);
nor NOR3 (N2349, N2347, N509, N2001);
nor NOR3 (N2350, N2346, N663, N1583);
or OR3 (N2351, N2348, N270, N2015);
xor XOR2 (N2352, N2350, N1773);
nor NOR4 (N2353, N2337, N1563, N878, N1922);
buf BUF1 (N2354, N2349);
buf BUF1 (N2355, N2353);
not NOT1 (N2356, N2340);
not NOT1 (N2357, N2339);
nor NOR4 (N2358, N2352, N1031, N648, N719);
not NOT1 (N2359, N2356);
nor NOR4 (N2360, N2318, N1010, N1754, N1077);
nor NOR2 (N2361, N2358, N528);
nand NAND3 (N2362, N2357, N1976, N1897);
not NOT1 (N2363, N2345);
and AND4 (N2364, N2360, N592, N2051, N1982);
or OR4 (N2365, N2361, N2323, N719, N1429);
nand NAND3 (N2366, N2363, N1290, N641);
nor NOR3 (N2367, N2354, N595, N143);
nand NAND3 (N2368, N2366, N1845, N2291);
or OR3 (N2369, N2355, N1607, N832);
buf BUF1 (N2370, N2368);
and AND4 (N2371, N2369, N2116, N1801, N1885);
nor NOR2 (N2372, N2351, N197);
xor XOR2 (N2373, N2364, N1778);
xor XOR2 (N2374, N2359, N60);
buf BUF1 (N2375, N2362);
not NOT1 (N2376, N2373);
xor XOR2 (N2377, N2374, N248);
nand NAND4 (N2378, N2372, N2307, N1938, N1042);
nand NAND2 (N2379, N2376, N1290);
buf BUF1 (N2380, N2370);
not NOT1 (N2381, N2312);
xor XOR2 (N2382, N2367, N1509);
and AND2 (N2383, N2382, N989);
nor NOR4 (N2384, N2378, N698, N2190, N329);
and AND2 (N2385, N2380, N1073);
nor NOR3 (N2386, N2371, N1293, N903);
and AND3 (N2387, N2365, N1505, N1186);
and AND2 (N2388, N2386, N1860);
buf BUF1 (N2389, N2388);
nor NOR4 (N2390, N2385, N695, N1707, N1397);
not NOT1 (N2391, N2390);
xor XOR2 (N2392, N2379, N880);
not NOT1 (N2393, N2392);
and AND4 (N2394, N2393, N1571, N1397, N1829);
nand NAND4 (N2395, N2391, N2368, N606, N1247);
buf BUF1 (N2396, N2389);
nand NAND4 (N2397, N2394, N1930, N911, N994);
buf BUF1 (N2398, N2383);
xor XOR2 (N2399, N2384, N645);
not NOT1 (N2400, N2395);
not NOT1 (N2401, N2396);
and AND4 (N2402, N2377, N937, N467, N828);
xor XOR2 (N2403, N2399, N167);
nand NAND4 (N2404, N2381, N608, N346, N2057);
nand NAND4 (N2405, N2397, N923, N1451, N166);
not NOT1 (N2406, N2344);
xor XOR2 (N2407, N2403, N1107);
nor NOR2 (N2408, N2406, N2085);
nand NAND3 (N2409, N2404, N1081, N1991);
and AND3 (N2410, N2407, N148, N564);
not NOT1 (N2411, N2398);
not NOT1 (N2412, N2402);
nand NAND2 (N2413, N2410, N1244);
nand NAND4 (N2414, N2401, N2044, N1521, N254);
nor NOR4 (N2415, N2409, N172, N564, N77);
buf BUF1 (N2416, N2414);
and AND2 (N2417, N2412, N2192);
or OR4 (N2418, N2415, N1243, N1698, N2050);
or OR3 (N2419, N2416, N1516, N2364);
not NOT1 (N2420, N2405);
buf BUF1 (N2421, N2411);
or OR3 (N2422, N2413, N1381, N2007);
nand NAND3 (N2423, N2418, N1159, N2379);
nand NAND2 (N2424, N2421, N457);
nand NAND3 (N2425, N2420, N2420, N2060);
buf BUF1 (N2426, N2400);
nand NAND3 (N2427, N2425, N1753, N826);
nor NOR4 (N2428, N2375, N2309, N683, N239);
or OR2 (N2429, N2387, N1763);
xor XOR2 (N2430, N2422, N441);
nor NOR3 (N2431, N2429, N1006, N790);
not NOT1 (N2432, N2424);
nor NOR2 (N2433, N2408, N1643);
or OR2 (N2434, N2427, N1);
not NOT1 (N2435, N2428);
and AND3 (N2436, N2423, N1743, N1648);
nor NOR2 (N2437, N2432, N285);
or OR3 (N2438, N2430, N1828, N556);
buf BUF1 (N2439, N2435);
or OR4 (N2440, N2417, N315, N957, N598);
nor NOR2 (N2441, N2439, N564);
or OR4 (N2442, N2434, N187, N1791, N1095);
xor XOR2 (N2443, N2419, N1064);
buf BUF1 (N2444, N2426);
nor NOR4 (N2445, N2441, N1004, N1458, N2034);
not NOT1 (N2446, N2438);
not NOT1 (N2447, N2433);
not NOT1 (N2448, N2447);
nand NAND2 (N2449, N2440, N1891);
or OR4 (N2450, N2442, N2053, N94, N2191);
nor NOR4 (N2451, N2448, N367, N185, N1445);
nand NAND2 (N2452, N2431, N1592);
nor NOR4 (N2453, N2449, N1538, N106, N2070);
and AND3 (N2454, N2444, N963, N793);
nor NOR3 (N2455, N2445, N982, N1239);
xor XOR2 (N2456, N2436, N2070);
not NOT1 (N2457, N2455);
not NOT1 (N2458, N2443);
xor XOR2 (N2459, N2457, N2414);
and AND3 (N2460, N2452, N1943, N294);
buf BUF1 (N2461, N2460);
xor XOR2 (N2462, N2446, N1641);
xor XOR2 (N2463, N2456, N1643);
not NOT1 (N2464, N2461);
nor NOR4 (N2465, N2453, N1258, N1202, N2235);
nor NOR4 (N2466, N2454, N858, N1605, N2105);
not NOT1 (N2467, N2458);
nand NAND3 (N2468, N2466, N2138, N1524);
not NOT1 (N2469, N2463);
not NOT1 (N2470, N2469);
and AND2 (N2471, N2462, N473);
not NOT1 (N2472, N2465);
xor XOR2 (N2473, N2467, N1256);
not NOT1 (N2474, N2437);
or OR2 (N2475, N2450, N899);
xor XOR2 (N2476, N2474, N238);
nand NAND4 (N2477, N2471, N653, N780, N438);
nand NAND4 (N2478, N2475, N1716, N386, N1833);
nor NOR3 (N2479, N2451, N2159, N1950);
xor XOR2 (N2480, N2476, N1145);
xor XOR2 (N2481, N2479, N1675);
xor XOR2 (N2482, N2464, N315);
and AND2 (N2483, N2470, N721);
or OR2 (N2484, N2480, N2080);
nand NAND2 (N2485, N2472, N1913);
not NOT1 (N2486, N2484);
or OR2 (N2487, N2483, N1002);
buf BUF1 (N2488, N2485);
buf BUF1 (N2489, N2478);
xor XOR2 (N2490, N2468, N657);
nor NOR2 (N2491, N2486, N634);
not NOT1 (N2492, N2482);
buf BUF1 (N2493, N2487);
buf BUF1 (N2494, N2459);
nor NOR3 (N2495, N2494, N2353, N934);
or OR2 (N2496, N2495, N1212);
xor XOR2 (N2497, N2490, N2039);
nand NAND3 (N2498, N2496, N89, N1717);
and AND2 (N2499, N2492, N2044);
and AND4 (N2500, N2493, N1721, N26, N379);
nor NOR3 (N2501, N2473, N141, N2229);
buf BUF1 (N2502, N2497);
or OR2 (N2503, N2499, N886);
nor NOR4 (N2504, N2498, N2027, N1324, N1);
nor NOR3 (N2505, N2500, N584, N902);
or OR4 (N2506, N2488, N370, N222, N1279);
buf BUF1 (N2507, N2503);
nand NAND2 (N2508, N2481, N234);
nand NAND4 (N2509, N2506, N1124, N1168, N2485);
not NOT1 (N2510, N2489);
nand NAND3 (N2511, N2502, N1436, N1172);
and AND4 (N2512, N2507, N1343, N1077, N1973);
buf BUF1 (N2513, N2505);
nand NAND3 (N2514, N2508, N1488, N1123);
and AND3 (N2515, N2477, N28, N1786);
not NOT1 (N2516, N2504);
xor XOR2 (N2517, N2514, N2179);
nand NAND3 (N2518, N2513, N1162, N1218);
buf BUF1 (N2519, N2491);
not NOT1 (N2520, N2510);
nor NOR2 (N2521, N2511, N459);
and AND3 (N2522, N2509, N107, N2508);
buf BUF1 (N2523, N2515);
buf BUF1 (N2524, N2516);
and AND2 (N2525, N2521, N2099);
buf BUF1 (N2526, N2520);
nand NAND2 (N2527, N2525, N714);
and AND4 (N2528, N2501, N1326, N429, N721);
nand NAND4 (N2529, N2517, N482, N231, N11);
nand NAND4 (N2530, N2526, N1843, N998, N671);
or OR3 (N2531, N2524, N31, N323);
nor NOR3 (N2532, N2529, N2146, N2201);
xor XOR2 (N2533, N2527, N42);
or OR4 (N2534, N2512, N285, N1005, N2344);
xor XOR2 (N2535, N2519, N50);
or OR4 (N2536, N2534, N1659, N1579, N1064);
nand NAND2 (N2537, N2533, N1912);
nand NAND2 (N2538, N2522, N1509);
xor XOR2 (N2539, N2538, N1640);
not NOT1 (N2540, N2537);
nand NAND2 (N2541, N2528, N2072);
not NOT1 (N2542, N2536);
nand NAND4 (N2543, N2539, N1063, N1553, N1168);
buf BUF1 (N2544, N2531);
or OR2 (N2545, N2535, N546);
nand NAND2 (N2546, N2532, N2438);
and AND2 (N2547, N2541, N2021);
xor XOR2 (N2548, N2542, N168);
nor NOR4 (N2549, N2544, N11, N719, N1918);
nor NOR2 (N2550, N2549, N281);
xor XOR2 (N2551, N2545, N856);
and AND3 (N2552, N2547, N1753, N2348);
or OR4 (N2553, N2551, N805, N2424, N2108);
or OR2 (N2554, N2550, N1617);
and AND2 (N2555, N2518, N239);
not NOT1 (N2556, N2555);
xor XOR2 (N2557, N2530, N1072);
nor NOR4 (N2558, N2523, N881, N1158, N393);
xor XOR2 (N2559, N2548, N1938);
xor XOR2 (N2560, N2552, N1343);
not NOT1 (N2561, N2540);
and AND4 (N2562, N2546, N348, N342, N429);
nand NAND3 (N2563, N2560, N929, N591);
or OR3 (N2564, N2543, N2492, N825);
nand NAND2 (N2565, N2556, N1448);
buf BUF1 (N2566, N2562);
nor NOR3 (N2567, N2554, N908, N904);
or OR4 (N2568, N2564, N1736, N183, N2170);
nor NOR3 (N2569, N2553, N2056, N427);
xor XOR2 (N2570, N2569, N399);
buf BUF1 (N2571, N2566);
and AND2 (N2572, N2561, N2518);
xor XOR2 (N2573, N2568, N763);
not NOT1 (N2574, N2563);
nand NAND4 (N2575, N2557, N1736, N953, N1270);
or OR3 (N2576, N2572, N1140, N2098);
nand NAND2 (N2577, N2571, N1522);
xor XOR2 (N2578, N2574, N2255);
and AND3 (N2579, N2573, N1836, N541);
buf BUF1 (N2580, N2558);
not NOT1 (N2581, N2578);
buf BUF1 (N2582, N2567);
or OR3 (N2583, N2580, N67, N2493);
and AND4 (N2584, N2582, N1988, N893, N68);
and AND3 (N2585, N2575, N2554, N1957);
nand NAND4 (N2586, N2565, N445, N2564, N995);
xor XOR2 (N2587, N2559, N2471);
or OR2 (N2588, N2586, N2095);
or OR2 (N2589, N2588, N85);
and AND3 (N2590, N2577, N2042, N2130);
nand NAND2 (N2591, N2583, N1723);
nand NAND2 (N2592, N2579, N63);
xor XOR2 (N2593, N2591, N489);
nor NOR2 (N2594, N2576, N417);
buf BUF1 (N2595, N2587);
not NOT1 (N2596, N2595);
xor XOR2 (N2597, N2584, N1821);
xor XOR2 (N2598, N2594, N2141);
buf BUF1 (N2599, N2589);
buf BUF1 (N2600, N2596);
not NOT1 (N2601, N2581);
nor NOR3 (N2602, N2570, N833, N1872);
xor XOR2 (N2603, N2590, N1294);
and AND2 (N2604, N2601, N241);
xor XOR2 (N2605, N2602, N1749);
not NOT1 (N2606, N2598);
xor XOR2 (N2607, N2600, N1912);
nor NOR4 (N2608, N2592, N857, N740, N299);
xor XOR2 (N2609, N2608, N1699);
or OR4 (N2610, N2585, N1582, N1857, N807);
not NOT1 (N2611, N2597);
nand NAND3 (N2612, N2607, N2080, N1045);
not NOT1 (N2613, N2610);
nor NOR3 (N2614, N2609, N1079, N1701);
nor NOR3 (N2615, N2603, N1605, N1888);
buf BUF1 (N2616, N2615);
nor NOR4 (N2617, N2605, N674, N332, N2336);
not NOT1 (N2618, N2612);
and AND3 (N2619, N2617, N1820, N2035);
xor XOR2 (N2620, N2616, N470);
nand NAND3 (N2621, N2611, N279, N244);
buf BUF1 (N2622, N2618);
and AND2 (N2623, N2593, N2362);
nand NAND3 (N2624, N2599, N1226, N2249);
nor NOR2 (N2625, N2606, N472);
and AND3 (N2626, N2614, N2501, N1390);
buf BUF1 (N2627, N2625);
or OR3 (N2628, N2613, N1112, N1837);
or OR2 (N2629, N2628, N700);
nor NOR4 (N2630, N2622, N1610, N1748, N270);
buf BUF1 (N2631, N2624);
nand NAND4 (N2632, N2621, N445, N1431, N802);
nor NOR4 (N2633, N2629, N1684, N281, N1564);
not NOT1 (N2634, N2604);
nor NOR3 (N2635, N2631, N816, N1004);
nand NAND4 (N2636, N2619, N2290, N727, N2434);
xor XOR2 (N2637, N2626, N91);
buf BUF1 (N2638, N2633);
xor XOR2 (N2639, N2620, N2549);
and AND4 (N2640, N2632, N2028, N1089, N507);
nand NAND3 (N2641, N2634, N354, N2078);
buf BUF1 (N2642, N2630);
and AND4 (N2643, N2635, N2486, N2403, N315);
not NOT1 (N2644, N2627);
nor NOR4 (N2645, N2637, N1766, N2327, N167);
nor NOR4 (N2646, N2636, N1432, N2498, N1778);
or OR2 (N2647, N2641, N1826);
nand NAND3 (N2648, N2638, N1270, N876);
and AND2 (N2649, N2647, N1873);
not NOT1 (N2650, N2639);
not NOT1 (N2651, N2623);
or OR4 (N2652, N2646, N2429, N1953, N669);
xor XOR2 (N2653, N2651, N909);
nand NAND4 (N2654, N2645, N2180, N1029, N1679);
and AND3 (N2655, N2653, N1880, N2034);
not NOT1 (N2656, N2643);
or OR3 (N2657, N2642, N1376, N1124);
or OR2 (N2658, N2657, N1005);
nand NAND3 (N2659, N2658, N493, N768);
xor XOR2 (N2660, N2649, N1784);
xor XOR2 (N2661, N2650, N390);
nor NOR2 (N2662, N2659, N1144);
not NOT1 (N2663, N2660);
nand NAND2 (N2664, N2656, N1963);
nor NOR3 (N2665, N2663, N1642, N583);
nor NOR4 (N2666, N2652, N1001, N56, N2044);
nand NAND3 (N2667, N2665, N1096, N633);
buf BUF1 (N2668, N2662);
nor NOR3 (N2669, N2640, N705, N2011);
nand NAND3 (N2670, N2661, N377, N1352);
not NOT1 (N2671, N2648);
nand NAND2 (N2672, N2664, N218);
nor NOR2 (N2673, N2667, N968);
and AND4 (N2674, N2644, N131, N294, N2503);
nand NAND2 (N2675, N2668, N577);
and AND2 (N2676, N2673, N477);
or OR2 (N2677, N2672, N169);
buf BUF1 (N2678, N2671);
not NOT1 (N2679, N2670);
or OR4 (N2680, N2669, N68, N330, N1428);
buf BUF1 (N2681, N2654);
or OR4 (N2682, N2675, N592, N2175, N1054);
xor XOR2 (N2683, N2681, N2068);
nor NOR4 (N2684, N2677, N317, N1518, N1206);
or OR3 (N2685, N2679, N1700, N956);
xor XOR2 (N2686, N2666, N904);
not NOT1 (N2687, N2686);
nand NAND3 (N2688, N2676, N2371, N2018);
nand NAND3 (N2689, N2684, N234, N2364);
xor XOR2 (N2690, N2687, N2418);
not NOT1 (N2691, N2680);
buf BUF1 (N2692, N2689);
not NOT1 (N2693, N2678);
xor XOR2 (N2694, N2692, N354);
nor NOR3 (N2695, N2688, N1186, N2590);
nor NOR4 (N2696, N2690, N777, N2071, N1887);
nand NAND2 (N2697, N2696, N1134);
or OR3 (N2698, N2695, N1193, N1973);
and AND4 (N2699, N2693, N79, N841, N1273);
nor NOR3 (N2700, N2655, N1744, N1025);
and AND3 (N2701, N2682, N1441, N1059);
nand NAND4 (N2702, N2698, N680, N1469, N995);
xor XOR2 (N2703, N2697, N1571);
nand NAND4 (N2704, N2694, N558, N1829, N1650);
nand NAND2 (N2705, N2702, N411);
xor XOR2 (N2706, N2701, N1215);
nor NOR2 (N2707, N2703, N885);
xor XOR2 (N2708, N2705, N2293);
nor NOR2 (N2709, N2700, N2201);
nand NAND2 (N2710, N2691, N140);
not NOT1 (N2711, N2704);
and AND4 (N2712, N2709, N2054, N2095, N2212);
nand NAND2 (N2713, N2674, N402);
nand NAND3 (N2714, N2710, N1550, N506);
nor NOR3 (N2715, N2699, N2681, N14);
xor XOR2 (N2716, N2715, N1165);
or OR2 (N2717, N2706, N276);
nand NAND3 (N2718, N2712, N1417, N1605);
buf BUF1 (N2719, N2718);
nor NOR3 (N2720, N2719, N521, N514);
buf BUF1 (N2721, N2707);
buf BUF1 (N2722, N2713);
buf BUF1 (N2723, N2721);
not NOT1 (N2724, N2722);
nor NOR3 (N2725, N2685, N1439, N2257);
not NOT1 (N2726, N2714);
nand NAND2 (N2727, N2708, N1963);
nand NAND4 (N2728, N2725, N2037, N1315, N2409);
nand NAND2 (N2729, N2717, N450);
xor XOR2 (N2730, N2729, N234);
and AND3 (N2731, N2683, N2469, N442);
nor NOR2 (N2732, N2724, N2210);
not NOT1 (N2733, N2727);
or OR4 (N2734, N2711, N886, N969, N1133);
or OR3 (N2735, N2734, N707, N2526);
nor NOR4 (N2736, N2720, N1970, N1691, N36);
buf BUF1 (N2737, N2731);
nor NOR2 (N2738, N2726, N786);
buf BUF1 (N2739, N2732);
not NOT1 (N2740, N2723);
or OR2 (N2741, N2737, N2590);
and AND4 (N2742, N2735, N2345, N1304, N1799);
nor NOR2 (N2743, N2716, N1257);
xor XOR2 (N2744, N2736, N435);
or OR2 (N2745, N2743, N540);
buf BUF1 (N2746, N2733);
or OR3 (N2747, N2730, N74, N602);
xor XOR2 (N2748, N2742, N386);
or OR4 (N2749, N2748, N325, N848, N2495);
buf BUF1 (N2750, N2739);
xor XOR2 (N2751, N2750, N833);
not NOT1 (N2752, N2746);
or OR3 (N2753, N2741, N2669, N2315);
or OR3 (N2754, N2751, N1395, N1693);
and AND2 (N2755, N2745, N1014);
nand NAND2 (N2756, N2749, N2486);
nor NOR4 (N2757, N2754, N650, N1984, N579);
buf BUF1 (N2758, N2738);
and AND4 (N2759, N2753, N845, N623, N2477);
xor XOR2 (N2760, N2759, N801);
nand NAND4 (N2761, N2747, N103, N2188, N1269);
buf BUF1 (N2762, N2760);
xor XOR2 (N2763, N2728, N83);
not NOT1 (N2764, N2762);
nor NOR2 (N2765, N2755, N359);
nand NAND2 (N2766, N2756, N110);
nand NAND3 (N2767, N2744, N400, N2380);
nor NOR4 (N2768, N2761, N792, N49, N2174);
buf BUF1 (N2769, N2766);
and AND3 (N2770, N2758, N1840, N1155);
nand NAND3 (N2771, N2767, N1884, N1255);
nand NAND4 (N2772, N2764, N308, N1658, N620);
xor XOR2 (N2773, N2752, N2023);
or OR2 (N2774, N2768, N394);
nand NAND2 (N2775, N2770, N419);
buf BUF1 (N2776, N2773);
buf BUF1 (N2777, N2771);
buf BUF1 (N2778, N2775);
xor XOR2 (N2779, N2777, N1234);
not NOT1 (N2780, N2740);
xor XOR2 (N2781, N2763, N2054);
and AND3 (N2782, N2774, N766, N542);
and AND4 (N2783, N2769, N70, N797, N1839);
buf BUF1 (N2784, N2779);
nor NOR2 (N2785, N2780, N2292);
nand NAND4 (N2786, N2778, N601, N875, N985);
nand NAND3 (N2787, N2757, N644, N736);
nor NOR4 (N2788, N2787, N2173, N2069, N2702);
nand NAND2 (N2789, N2785, N1916);
not NOT1 (N2790, N2781);
not NOT1 (N2791, N2786);
or OR2 (N2792, N2783, N818);
nand NAND4 (N2793, N2772, N1369, N1167, N805);
nand NAND2 (N2794, N2792, N1398);
xor XOR2 (N2795, N2789, N243);
nor NOR2 (N2796, N2795, N982);
buf BUF1 (N2797, N2793);
buf BUF1 (N2798, N2797);
xor XOR2 (N2799, N2788, N1899);
buf BUF1 (N2800, N2784);
buf BUF1 (N2801, N2776);
xor XOR2 (N2802, N2794, N2379);
and AND4 (N2803, N2782, N1265, N1737, N1349);
or OR2 (N2804, N2802, N2119);
or OR3 (N2805, N2800, N558, N773);
not NOT1 (N2806, N2803);
and AND2 (N2807, N2799, N371);
not NOT1 (N2808, N2807);
nor NOR2 (N2809, N2806, N1258);
nand NAND2 (N2810, N2805, N493);
nand NAND4 (N2811, N2804, N1982, N719, N2601);
buf BUF1 (N2812, N2809);
xor XOR2 (N2813, N2765, N2333);
not NOT1 (N2814, N2801);
nand NAND4 (N2815, N2813, N669, N2648, N1411);
nor NOR3 (N2816, N2791, N726, N1870);
xor XOR2 (N2817, N2790, N2711);
xor XOR2 (N2818, N2814, N1049);
nand NAND3 (N2819, N2811, N2324, N378);
nor NOR2 (N2820, N2819, N433);
nor NOR3 (N2821, N2818, N709, N1508);
xor XOR2 (N2822, N2821, N1274);
and AND2 (N2823, N2815, N2337);
xor XOR2 (N2824, N2822, N1463);
not NOT1 (N2825, N2812);
not NOT1 (N2826, N2796);
buf BUF1 (N2827, N2820);
or OR2 (N2828, N2816, N2243);
or OR4 (N2829, N2824, N5, N792, N413);
nand NAND4 (N2830, N2808, N395, N2606, N1471);
and AND3 (N2831, N2829, N1516, N2242);
nand NAND3 (N2832, N2798, N1065, N1454);
nand NAND3 (N2833, N2826, N83, N133);
buf BUF1 (N2834, N2830);
or OR4 (N2835, N2831, N1882, N2545, N2192);
xor XOR2 (N2836, N2823, N738);
or OR4 (N2837, N2835, N1284, N1067, N1611);
not NOT1 (N2838, N2810);
nor NOR3 (N2839, N2837, N430, N834);
and AND2 (N2840, N2836, N916);
or OR2 (N2841, N2825, N2059);
and AND4 (N2842, N2827, N1596, N2689, N915);
nor NOR3 (N2843, N2817, N2791, N2113);
and AND2 (N2844, N2833, N2055);
nand NAND2 (N2845, N2842, N575);
nor NOR2 (N2846, N2834, N1358);
or OR2 (N2847, N2846, N2264);
xor XOR2 (N2848, N2841, N1550);
and AND4 (N2849, N2844, N989, N2530, N1086);
xor XOR2 (N2850, N2845, N2166);
buf BUF1 (N2851, N2832);
buf BUF1 (N2852, N2828);
nor NOR2 (N2853, N2852, N44);
buf BUF1 (N2854, N2840);
nand NAND3 (N2855, N2851, N2097, N815);
and AND3 (N2856, N2838, N825, N1353);
nor NOR4 (N2857, N2853, N1919, N1518, N2441);
nor NOR2 (N2858, N2856, N68);
buf BUF1 (N2859, N2839);
xor XOR2 (N2860, N2848, N1008);
and AND4 (N2861, N2847, N552, N2178, N2400);
and AND3 (N2862, N2850, N1197, N2858);
xor XOR2 (N2863, N1075, N2519);
not NOT1 (N2864, N2862);
nand NAND2 (N2865, N2864, N2457);
xor XOR2 (N2866, N2860, N108);
buf BUF1 (N2867, N2859);
nand NAND2 (N2868, N2861, N353);
xor XOR2 (N2869, N2868, N110);
and AND4 (N2870, N2866, N1644, N2390, N2596);
or OR3 (N2871, N2857, N464, N1637);
or OR4 (N2872, N2855, N1737, N1012, N1919);
and AND3 (N2873, N2849, N446, N329);
nand NAND2 (N2874, N2872, N1661);
and AND3 (N2875, N2870, N1437, N1544);
not NOT1 (N2876, N2843);
xor XOR2 (N2877, N2869, N2204);
not NOT1 (N2878, N2865);
nand NAND4 (N2879, N2878, N1380, N2867, N2589);
and AND3 (N2880, N2353, N895, N291);
or OR4 (N2881, N2879, N2856, N456, N1369);
xor XOR2 (N2882, N2875, N805);
nand NAND4 (N2883, N2871, N1927, N785, N1659);
or OR3 (N2884, N2863, N364, N228);
and AND2 (N2885, N2873, N2093);
xor XOR2 (N2886, N2876, N1556);
and AND2 (N2887, N2884, N609);
not NOT1 (N2888, N2883);
or OR2 (N2889, N2887, N848);
nor NOR3 (N2890, N2854, N1017, N2691);
or OR3 (N2891, N2874, N2718, N1840);
or OR3 (N2892, N2891, N762, N2382);
and AND3 (N2893, N2877, N2782, N455);
not NOT1 (N2894, N2885);
xor XOR2 (N2895, N2882, N1430);
xor XOR2 (N2896, N2881, N599);
and AND3 (N2897, N2893, N2083, N1125);
xor XOR2 (N2898, N2895, N765);
nor NOR4 (N2899, N2886, N929, N2483, N362);
not NOT1 (N2900, N2897);
not NOT1 (N2901, N2880);
not NOT1 (N2902, N2888);
nor NOR4 (N2903, N2898, N2542, N1253, N1663);
buf BUF1 (N2904, N2890);
buf BUF1 (N2905, N2900);
not NOT1 (N2906, N2905);
nor NOR4 (N2907, N2901, N890, N1496, N1942);
or OR4 (N2908, N2894, N26, N763, N1813);
and AND3 (N2909, N2903, N2689, N1189);
nand NAND2 (N2910, N2902, N1381);
not NOT1 (N2911, N2899);
nand NAND2 (N2912, N2907, N643);
xor XOR2 (N2913, N2910, N663);
nor NOR3 (N2914, N2909, N1855, N2635);
or OR3 (N2915, N2911, N50, N12);
xor XOR2 (N2916, N2906, N2057);
nand NAND4 (N2917, N2912, N871, N1273, N388);
not NOT1 (N2918, N2908);
not NOT1 (N2919, N2918);
not NOT1 (N2920, N2916);
and AND3 (N2921, N2913, N2422, N1878);
nor NOR2 (N2922, N2917, N618);
buf BUF1 (N2923, N2914);
nand NAND4 (N2924, N2896, N1519, N449, N858);
nor NOR4 (N2925, N2904, N1475, N1753, N1534);
nand NAND4 (N2926, N2920, N1984, N1621, N335);
nand NAND2 (N2927, N2919, N475);
nand NAND2 (N2928, N2922, N1529);
or OR4 (N2929, N2915, N649, N522, N2889);
xor XOR2 (N2930, N2379, N2281);
or OR3 (N2931, N2930, N108, N2328);
and AND2 (N2932, N2921, N1657);
and AND4 (N2933, N2928, N2014, N1211, N1355);
and AND4 (N2934, N2933, N2189, N2346, N2125);
nor NOR3 (N2935, N2926, N1670, N2094);
buf BUF1 (N2936, N2929);
or OR2 (N2937, N2923, N793);
buf BUF1 (N2938, N2927);
or OR4 (N2939, N2934, N1998, N2560, N1436);
nand NAND3 (N2940, N2936, N1302, N1698);
nor NOR3 (N2941, N2931, N2351, N1029);
and AND2 (N2942, N2925, N27);
nor NOR4 (N2943, N2937, N1511, N173, N2520);
xor XOR2 (N2944, N2941, N2204);
nor NOR3 (N2945, N2944, N519, N2112);
or OR2 (N2946, N2935, N2888);
nand NAND3 (N2947, N2924, N1256, N2120);
nand NAND2 (N2948, N2892, N1271);
or OR2 (N2949, N2938, N2248);
xor XOR2 (N2950, N2947, N2241);
nor NOR2 (N2951, N2945, N1052);
nand NAND2 (N2952, N2943, N1326);
nand NAND2 (N2953, N2948, N1302);
xor XOR2 (N2954, N2932, N1302);
buf BUF1 (N2955, N2939);
nor NOR4 (N2956, N2953, N1497, N2902, N1155);
and AND3 (N2957, N2952, N1542, N2314);
or OR2 (N2958, N2942, N2332);
xor XOR2 (N2959, N2946, N2018);
not NOT1 (N2960, N2956);
nor NOR2 (N2961, N2949, N2280);
nor NOR3 (N2962, N2958, N1716, N1732);
buf BUF1 (N2963, N2957);
buf BUF1 (N2964, N2951);
nor NOR4 (N2965, N2961, N1928, N817, N2539);
nand NAND2 (N2966, N2950, N983);
xor XOR2 (N2967, N2959, N2582);
nor NOR2 (N2968, N2965, N1119);
and AND3 (N2969, N2966, N2449, N1037);
or OR4 (N2970, N2955, N188, N1459, N1427);
xor XOR2 (N2971, N2968, N1193);
not NOT1 (N2972, N2969);
not NOT1 (N2973, N2967);
and AND3 (N2974, N2964, N1421, N288);
nor NOR3 (N2975, N2971, N2524, N337);
buf BUF1 (N2976, N2960);
or OR2 (N2977, N2954, N2495);
buf BUF1 (N2978, N2972);
nor NOR2 (N2979, N2978, N2073);
buf BUF1 (N2980, N2973);
and AND2 (N2981, N2977, N565);
nor NOR2 (N2982, N2940, N1405);
nand NAND3 (N2983, N2980, N578, N1270);
nand NAND3 (N2984, N2983, N1871, N1028);
or OR4 (N2985, N2982, N1189, N2609, N2175);
buf BUF1 (N2986, N2976);
and AND4 (N2987, N2963, N1745, N452, N1021);
or OR3 (N2988, N2974, N246, N161);
xor XOR2 (N2989, N2981, N2692);
nor NOR3 (N2990, N2986, N588, N2196);
nor NOR2 (N2991, N2975, N2437);
nor NOR3 (N2992, N2991, N2303, N2404);
nand NAND3 (N2993, N2985, N2815, N2597);
or OR3 (N2994, N2970, N2633, N385);
nor NOR3 (N2995, N2990, N2943, N1290);
nand NAND3 (N2996, N2984, N2331, N618);
and AND2 (N2997, N2992, N1995);
nor NOR2 (N2998, N2989, N1690);
or OR3 (N2999, N2995, N73, N1802);
nor NOR3 (N3000, N2997, N84, N714);
buf BUF1 (N3001, N3000);
buf BUF1 (N3002, N2962);
not NOT1 (N3003, N2998);
nand NAND4 (N3004, N2996, N133, N96, N2730);
and AND3 (N3005, N3003, N115, N877);
not NOT1 (N3006, N2987);
and AND2 (N3007, N2994, N2001);
or OR2 (N3008, N2979, N562);
buf BUF1 (N3009, N3007);
nor NOR3 (N3010, N3002, N1731, N2848);
not NOT1 (N3011, N3005);
nand NAND4 (N3012, N2999, N1415, N615, N608);
nand NAND2 (N3013, N3001, N149);
xor XOR2 (N3014, N3004, N2941);
nor NOR4 (N3015, N2993, N1444, N474, N259);
xor XOR2 (N3016, N3013, N1453);
xor XOR2 (N3017, N3016, N2270);
nor NOR2 (N3018, N3008, N1498);
nand NAND2 (N3019, N3006, N145);
xor XOR2 (N3020, N3019, N2074);
xor XOR2 (N3021, N3017, N172);
not NOT1 (N3022, N3015);
and AND2 (N3023, N3009, N152);
nand NAND2 (N3024, N3010, N1900);
not NOT1 (N3025, N2988);
or OR2 (N3026, N3011, N2702);
not NOT1 (N3027, N3018);
xor XOR2 (N3028, N3022, N2298);
buf BUF1 (N3029, N3014);
buf BUF1 (N3030, N3026);
or OR2 (N3031, N3030, N91);
nand NAND2 (N3032, N3027, N2563);
and AND3 (N3033, N3031, N2645, N1071);
nand NAND4 (N3034, N3023, N1616, N1626, N247);
buf BUF1 (N3035, N3024);
xor XOR2 (N3036, N3012, N2642);
nor NOR2 (N3037, N3025, N2032);
nand NAND2 (N3038, N3029, N2808);
or OR4 (N3039, N3036, N2772, N1711, N258);
not NOT1 (N3040, N3033);
buf BUF1 (N3041, N3028);
nor NOR3 (N3042, N3039, N2331, N644);
buf BUF1 (N3043, N3037);
buf BUF1 (N3044, N3020);
nand NAND3 (N3045, N3035, N505, N1892);
buf BUF1 (N3046, N3021);
xor XOR2 (N3047, N3038, N1439);
nor NOR2 (N3048, N3040, N2255);
nand NAND3 (N3049, N3048, N2682, N2111);
and AND4 (N3050, N3034, N2165, N1632, N1000);
and AND2 (N3051, N3044, N620);
nand NAND2 (N3052, N3042, N832);
buf BUF1 (N3053, N3050);
nor NOR3 (N3054, N3053, N1781, N2321);
not NOT1 (N3055, N3043);
nor NOR4 (N3056, N3041, N1187, N901, N642);
or OR4 (N3057, N3045, N1846, N628, N2054);
nand NAND3 (N3058, N3057, N2844, N3028);
xor XOR2 (N3059, N3051, N1465);
buf BUF1 (N3060, N3059);
or OR4 (N3061, N3055, N70, N1829, N850);
and AND3 (N3062, N3052, N1505, N903);
nand NAND3 (N3063, N3047, N1996, N49);
nor NOR2 (N3064, N3060, N388);
not NOT1 (N3065, N3049);
or OR4 (N3066, N3065, N1637, N1072, N2975);
nor NOR4 (N3067, N3054, N221, N2285, N549);
not NOT1 (N3068, N3067);
and AND2 (N3069, N3068, N430);
nand NAND3 (N3070, N3058, N327, N2966);
and AND2 (N3071, N3070, N446);
nand NAND3 (N3072, N3066, N1616, N198);
nand NAND4 (N3073, N3072, N884, N2769, N677);
nor NOR3 (N3074, N3046, N1277, N698);
and AND2 (N3075, N3056, N2000);
nand NAND4 (N3076, N3073, N2618, N1158, N2696);
xor XOR2 (N3077, N3069, N1520);
and AND2 (N3078, N3074, N733);
xor XOR2 (N3079, N3078, N249);
buf BUF1 (N3080, N3076);
nor NOR3 (N3081, N3079, N1579, N2481);
xor XOR2 (N3082, N3063, N94);
or OR3 (N3083, N3082, N2690, N2645);
nand NAND2 (N3084, N3080, N2603);
not NOT1 (N3085, N3032);
not NOT1 (N3086, N3075);
or OR4 (N3087, N3077, N2599, N2832, N357);
nor NOR4 (N3088, N3062, N2799, N2578, N1571);
or OR4 (N3089, N3071, N3046, N2815, N2903);
nor NOR4 (N3090, N3085, N2274, N497, N1949);
buf BUF1 (N3091, N3089);
xor XOR2 (N3092, N3090, N56);
or OR3 (N3093, N3083, N734, N1382);
nand NAND3 (N3094, N3081, N1005, N212);
and AND4 (N3095, N3086, N329, N2205, N2022);
or OR2 (N3096, N3088, N1461);
buf BUF1 (N3097, N3096);
buf BUF1 (N3098, N3095);
buf BUF1 (N3099, N3061);
not NOT1 (N3100, N3099);
not NOT1 (N3101, N3097);
and AND4 (N3102, N3091, N1231, N2328, N431);
or OR3 (N3103, N3101, N1328, N1516);
and AND2 (N3104, N3087, N1318);
not NOT1 (N3105, N3102);
xor XOR2 (N3106, N3103, N1699);
and AND2 (N3107, N3084, N1432);
nor NOR3 (N3108, N3064, N331, N1449);
nor NOR4 (N3109, N3092, N661, N2459, N200);
and AND3 (N3110, N3105, N2700, N2842);
nor NOR3 (N3111, N3108, N1002, N2173);
nand NAND3 (N3112, N3093, N1451, N2821);
xor XOR2 (N3113, N3109, N2825);
nor NOR3 (N3114, N3107, N2115, N1644);
buf BUF1 (N3115, N3106);
nand NAND3 (N3116, N3094, N1986, N2559);
nor NOR2 (N3117, N3100, N2370);
not NOT1 (N3118, N3117);
nand NAND3 (N3119, N3110, N80, N1834);
nor NOR4 (N3120, N3115, N1960, N735, N1236);
or OR4 (N3121, N3112, N1543, N1198, N1500);
xor XOR2 (N3122, N3119, N1230);
xor XOR2 (N3123, N3121, N437);
not NOT1 (N3124, N3104);
not NOT1 (N3125, N3122);
and AND2 (N3126, N3098, N1477);
xor XOR2 (N3127, N3120, N2580);
not NOT1 (N3128, N3127);
nand NAND4 (N3129, N3114, N2062, N2548, N2120);
not NOT1 (N3130, N3111);
not NOT1 (N3131, N3113);
or OR4 (N3132, N3125, N2479, N1277, N118);
nand NAND4 (N3133, N3129, N2004, N1166, N189);
not NOT1 (N3134, N3123);
or OR2 (N3135, N3116, N2828);
and AND2 (N3136, N3124, N1653);
nand NAND3 (N3137, N3134, N964, N932);
buf BUF1 (N3138, N3118);
and AND4 (N3139, N3130, N287, N1152, N842);
xor XOR2 (N3140, N3136, N1020);
nor NOR3 (N3141, N3128, N1757, N11);
or OR2 (N3142, N3138, N39);
and AND2 (N3143, N3135, N2077);
or OR4 (N3144, N3142, N94, N548, N1163);
buf BUF1 (N3145, N3140);
nand NAND4 (N3146, N3144, N1487, N493, N1185);
and AND3 (N3147, N3132, N61, N361);
nor NOR2 (N3148, N3141, N1116);
or OR2 (N3149, N3133, N1217);
nor NOR3 (N3150, N3143, N916, N128);
nand NAND3 (N3151, N3146, N653, N1718);
or OR4 (N3152, N3147, N3061, N876, N814);
not NOT1 (N3153, N3152);
or OR3 (N3154, N3137, N1477, N1973);
nor NOR4 (N3155, N3139, N2085, N1617, N1650);
and AND3 (N3156, N3145, N2371, N524);
xor XOR2 (N3157, N3151, N1353);
and AND4 (N3158, N3149, N404, N2341, N1146);
not NOT1 (N3159, N3131);
not NOT1 (N3160, N3158);
nor NOR2 (N3161, N3159, N1628);
nand NAND4 (N3162, N3161, N1367, N1011, N2673);
nor NOR2 (N3163, N3154, N2477);
or OR3 (N3164, N3163, N2928, N1214);
buf BUF1 (N3165, N3126);
not NOT1 (N3166, N3162);
xor XOR2 (N3167, N3165, N2740);
nand NAND3 (N3168, N3150, N2106, N1738);
buf BUF1 (N3169, N3156);
not NOT1 (N3170, N3168);
xor XOR2 (N3171, N3160, N3132);
and AND2 (N3172, N3171, N3113);
buf BUF1 (N3173, N3148);
and AND2 (N3174, N3172, N1397);
nand NAND3 (N3175, N3173, N2452, N2517);
nor NOR3 (N3176, N3169, N2300, N2937);
and AND2 (N3177, N3157, N2167);
or OR4 (N3178, N3153, N1385, N3056, N2925);
nor NOR2 (N3179, N3175, N236);
or OR2 (N3180, N3179, N1397);
xor XOR2 (N3181, N3166, N2022);
buf BUF1 (N3182, N3178);
not NOT1 (N3183, N3177);
not NOT1 (N3184, N3167);
and AND2 (N3185, N3180, N1352);
xor XOR2 (N3186, N3181, N395);
or OR2 (N3187, N3174, N9);
nor NOR4 (N3188, N3186, N1896, N1470, N123);
not NOT1 (N3189, N3182);
or OR4 (N3190, N3155, N2749, N265, N2837);
or OR2 (N3191, N3187, N3032);
buf BUF1 (N3192, N3164);
not NOT1 (N3193, N3190);
not NOT1 (N3194, N3191);
not NOT1 (N3195, N3183);
or OR4 (N3196, N3188, N808, N1858, N1491);
or OR2 (N3197, N3184, N1127);
or OR4 (N3198, N3196, N1514, N144, N1098);
not NOT1 (N3199, N3198);
or OR3 (N3200, N3195, N1905, N1480);
or OR3 (N3201, N3194, N533, N1110);
nor NOR3 (N3202, N3199, N473, N673);
or OR4 (N3203, N3202, N2780, N1631, N1904);
not NOT1 (N3204, N3203);
xor XOR2 (N3205, N3176, N2961);
or OR3 (N3206, N3193, N2985, N2015);
nand NAND2 (N3207, N3206, N2637);
not NOT1 (N3208, N3201);
xor XOR2 (N3209, N3192, N2414);
xor XOR2 (N3210, N3205, N1497);
xor XOR2 (N3211, N3207, N930);
nand NAND2 (N3212, N3185, N815);
not NOT1 (N3213, N3212);
nor NOR4 (N3214, N3200, N117, N1079, N2259);
and AND4 (N3215, N3210, N1229, N2436, N2316);
buf BUF1 (N3216, N3211);
or OR2 (N3217, N3216, N1056);
or OR3 (N3218, N3208, N2333, N2252);
or OR4 (N3219, N3218, N72, N1527, N1969);
or OR3 (N3220, N3213, N1803, N1240);
buf BUF1 (N3221, N3170);
not NOT1 (N3222, N3217);
nor NOR2 (N3223, N3197, N2590);
nor NOR4 (N3224, N3223, N1779, N1332, N2102);
nor NOR4 (N3225, N3189, N2830, N705, N209);
buf BUF1 (N3226, N3221);
nor NOR2 (N3227, N3222, N908);
or OR3 (N3228, N3204, N1644, N1539);
nand NAND4 (N3229, N3225, N108, N2925, N1178);
and AND4 (N3230, N3227, N3149, N999, N1155);
nor NOR4 (N3231, N3229, N1135, N1223, N1544);
nor NOR3 (N3232, N3214, N999, N1170);
buf BUF1 (N3233, N3231);
or OR3 (N3234, N3230, N2550, N936);
nand NAND3 (N3235, N3219, N3165, N2131);
not NOT1 (N3236, N3234);
and AND3 (N3237, N3228, N987, N1762);
or OR2 (N3238, N3215, N1860);
or OR2 (N3239, N3236, N1983);
nand NAND2 (N3240, N3232, N3188);
buf BUF1 (N3241, N3237);
not NOT1 (N3242, N3239);
nor NOR3 (N3243, N3226, N708, N468);
nand NAND4 (N3244, N3209, N1423, N1434, N2199);
and AND3 (N3245, N3242, N1323, N2743);
nor NOR4 (N3246, N3233, N969, N579, N1850);
not NOT1 (N3247, N3245);
nor NOR4 (N3248, N3240, N2518, N1501, N1641);
xor XOR2 (N3249, N3244, N164);
not NOT1 (N3250, N3241);
buf BUF1 (N3251, N3243);
nand NAND4 (N3252, N3220, N1273, N757, N852);
nand NAND4 (N3253, N3238, N844, N3154, N1366);
nor NOR3 (N3254, N3252, N3174, N1177);
xor XOR2 (N3255, N3254, N733);
buf BUF1 (N3256, N3251);
buf BUF1 (N3257, N3235);
and AND4 (N3258, N3257, N1213, N2481, N1519);
nand NAND2 (N3259, N3250, N939);
and AND4 (N3260, N3258, N2514, N201, N2184);
buf BUF1 (N3261, N3253);
buf BUF1 (N3262, N3246);
buf BUF1 (N3263, N3249);
buf BUF1 (N3264, N3224);
nand NAND3 (N3265, N3263, N2405, N2024);
not NOT1 (N3266, N3247);
or OR4 (N3267, N3259, N1954, N219, N186);
nor NOR2 (N3268, N3256, N2954);
and AND3 (N3269, N3265, N981, N3012);
nor NOR3 (N3270, N3266, N715, N2586);
nor NOR3 (N3271, N3255, N1678, N2203);
and AND4 (N3272, N3268, N1806, N292, N2155);
nand NAND4 (N3273, N3261, N547, N3260, N3239);
not NOT1 (N3274, N354);
not NOT1 (N3275, N3270);
and AND2 (N3276, N3248, N168);
nor NOR2 (N3277, N3276, N2481);
xor XOR2 (N3278, N3267, N198);
and AND2 (N3279, N3264, N1041);
or OR3 (N3280, N3262, N1426, N1878);
not NOT1 (N3281, N3273);
buf BUF1 (N3282, N3271);
buf BUF1 (N3283, N3272);
xor XOR2 (N3284, N3280, N2290);
or OR4 (N3285, N3275, N2298, N1678, N1412);
not NOT1 (N3286, N3274);
or OR4 (N3287, N3269, N1715, N546, N2032);
nor NOR2 (N3288, N3281, N2264);
buf BUF1 (N3289, N3284);
xor XOR2 (N3290, N3278, N595);
not NOT1 (N3291, N3288);
xor XOR2 (N3292, N3291, N352);
and AND3 (N3293, N3282, N1971, N117);
nor NOR4 (N3294, N3292, N1666, N1995, N2264);
nor NOR3 (N3295, N3293, N2326, N484);
and AND2 (N3296, N3283, N1564);
nor NOR3 (N3297, N3277, N179, N311);
and AND3 (N3298, N3279, N3207, N2886);
and AND3 (N3299, N3295, N1324, N619);
or OR4 (N3300, N3294, N1701, N2308, N213);
xor XOR2 (N3301, N3286, N1444);
not NOT1 (N3302, N3301);
buf BUF1 (N3303, N3297);
or OR3 (N3304, N3289, N1533, N1023);
nor NOR2 (N3305, N3304, N2236);
and AND3 (N3306, N3287, N3, N1091);
not NOT1 (N3307, N3296);
and AND4 (N3308, N3300, N100, N825, N270);
nor NOR3 (N3309, N3290, N481, N2991);
nand NAND2 (N3310, N3305, N1786);
and AND4 (N3311, N3303, N1931, N1201, N2573);
nand NAND2 (N3312, N3302, N2456);
xor XOR2 (N3313, N3310, N903);
and AND3 (N3314, N3309, N1864, N1122);
nor NOR3 (N3315, N3312, N1794, N3007);
buf BUF1 (N3316, N3311);
nand NAND2 (N3317, N3285, N530);
not NOT1 (N3318, N3298);
buf BUF1 (N3319, N3315);
not NOT1 (N3320, N3318);
nor NOR3 (N3321, N3308, N519, N197);
nand NAND3 (N3322, N3299, N2792, N1269);
xor XOR2 (N3323, N3307, N2124);
or OR3 (N3324, N3317, N1846, N114);
not NOT1 (N3325, N3321);
xor XOR2 (N3326, N3320, N2877);
nor NOR4 (N3327, N3314, N1115, N2529, N2559);
or OR3 (N3328, N3325, N1876, N893);
and AND2 (N3329, N3323, N486);
xor XOR2 (N3330, N3329, N3253);
not NOT1 (N3331, N3327);
nor NOR4 (N3332, N3306, N2278, N86, N2939);
not NOT1 (N3333, N3331);
or OR4 (N3334, N3328, N2712, N1770, N3053);
buf BUF1 (N3335, N3330);
or OR2 (N3336, N3319, N1981);
nor NOR2 (N3337, N3316, N2671);
not NOT1 (N3338, N3324);
nor NOR4 (N3339, N3338, N1105, N892, N3004);
not NOT1 (N3340, N3326);
and AND3 (N3341, N3332, N2586, N3098);
and AND3 (N3342, N3337, N3138, N444);
and AND4 (N3343, N3341, N2748, N3115, N742);
xor XOR2 (N3344, N3339, N1448);
not NOT1 (N3345, N3322);
xor XOR2 (N3346, N3345, N1612);
nor NOR3 (N3347, N3342, N698, N939);
and AND2 (N3348, N3343, N1050);
xor XOR2 (N3349, N3335, N177);
and AND4 (N3350, N3344, N2076, N2243, N2557);
xor XOR2 (N3351, N3349, N183);
nand NAND2 (N3352, N3347, N3217);
buf BUF1 (N3353, N3340);
nand NAND4 (N3354, N3334, N228, N2909, N2049);
and AND4 (N3355, N3313, N1544, N1982, N393);
not NOT1 (N3356, N3348);
xor XOR2 (N3357, N3356, N2529);
or OR4 (N3358, N3355, N1536, N2805, N2077);
xor XOR2 (N3359, N3358, N2039);
and AND4 (N3360, N3336, N786, N521, N31);
not NOT1 (N3361, N3360);
and AND3 (N3362, N3353, N771, N2633);
or OR4 (N3363, N3346, N3240, N518, N2446);
or OR4 (N3364, N3362, N2726, N2573, N3066);
nand NAND2 (N3365, N3364, N2465);
and AND3 (N3366, N3363, N1296, N2526);
nand NAND2 (N3367, N3333, N2967);
or OR4 (N3368, N3361, N2040, N2195, N2232);
nand NAND2 (N3369, N3368, N2400);
xor XOR2 (N3370, N3367, N1660);
and AND2 (N3371, N3370, N1901);
nand NAND3 (N3372, N3359, N1484, N2203);
buf BUF1 (N3373, N3354);
nand NAND3 (N3374, N3369, N117, N1004);
nand NAND3 (N3375, N3350, N113, N978);
nand NAND2 (N3376, N3374, N3103);
xor XOR2 (N3377, N3357, N643);
nand NAND3 (N3378, N3351, N1661, N497);
or OR2 (N3379, N3371, N2524);
buf BUF1 (N3380, N3352);
not NOT1 (N3381, N3366);
or OR2 (N3382, N3372, N2559);
not NOT1 (N3383, N3377);
and AND2 (N3384, N3381, N2352);
xor XOR2 (N3385, N3373, N810);
not NOT1 (N3386, N3375);
and AND3 (N3387, N3376, N2394, N1776);
and AND3 (N3388, N3384, N410, N3078);
buf BUF1 (N3389, N3382);
and AND3 (N3390, N3383, N418, N2814);
xor XOR2 (N3391, N3379, N1458);
nand NAND2 (N3392, N3387, N502);
nor NOR2 (N3393, N3386, N131);
not NOT1 (N3394, N3391);
not NOT1 (N3395, N3390);
not NOT1 (N3396, N3385);
or OR4 (N3397, N3394, N437, N340, N1450);
xor XOR2 (N3398, N3396, N1195);
and AND4 (N3399, N3380, N3132, N2027, N970);
buf BUF1 (N3400, N3392);
or OR4 (N3401, N3395, N2042, N1634, N2496);
xor XOR2 (N3402, N3378, N283);
not NOT1 (N3403, N3397);
not NOT1 (N3404, N3401);
and AND3 (N3405, N3393, N707, N3356);
xor XOR2 (N3406, N3405, N3075);
nor NOR4 (N3407, N3388, N2449, N810, N3003);
buf BUF1 (N3408, N3402);
buf BUF1 (N3409, N3365);
buf BUF1 (N3410, N3403);
or OR4 (N3411, N3398, N3347, N2826, N686);
buf BUF1 (N3412, N3404);
and AND4 (N3413, N3409, N1400, N2786, N357);
not NOT1 (N3414, N3410);
not NOT1 (N3415, N3407);
xor XOR2 (N3416, N3399, N3008);
nand NAND2 (N3417, N3415, N3051);
xor XOR2 (N3418, N3411, N935);
and AND4 (N3419, N3408, N434, N826, N3391);
and AND3 (N3420, N3414, N2399, N1766);
nand NAND2 (N3421, N3406, N383);
xor XOR2 (N3422, N3389, N1620);
and AND3 (N3423, N3400, N2390, N2110);
xor XOR2 (N3424, N3419, N2616);
or OR2 (N3425, N3413, N979);
not NOT1 (N3426, N3421);
nand NAND3 (N3427, N3420, N2433, N1014);
buf BUF1 (N3428, N3422);
xor XOR2 (N3429, N3425, N2778);
and AND2 (N3430, N3427, N1264);
nand NAND4 (N3431, N3424, N2134, N2413, N1796);
not NOT1 (N3432, N3428);
xor XOR2 (N3433, N3431, N2366);
buf BUF1 (N3434, N3430);
nand NAND2 (N3435, N3434, N2781);
or OR3 (N3436, N3426, N1197, N1285);
nor NOR3 (N3437, N3423, N2644, N1686);
buf BUF1 (N3438, N3432);
buf BUF1 (N3439, N3429);
not NOT1 (N3440, N3436);
and AND4 (N3441, N3416, N2643, N3038, N513);
nor NOR3 (N3442, N3417, N921, N3298);
not NOT1 (N3443, N3442);
or OR2 (N3444, N3438, N95);
not NOT1 (N3445, N3441);
nor NOR4 (N3446, N3418, N1289, N2468, N862);
xor XOR2 (N3447, N3445, N1003);
nand NAND3 (N3448, N3412, N2945, N3116);
nand NAND4 (N3449, N3448, N431, N1194, N2001);
and AND3 (N3450, N3446, N960, N696);
and AND2 (N3451, N3437, N2091);
or OR3 (N3452, N3443, N1543, N530);
xor XOR2 (N3453, N3447, N2507);
nand NAND2 (N3454, N3433, N2501);
or OR3 (N3455, N3440, N2595, N222);
and AND4 (N3456, N3449, N1671, N3004, N2275);
and AND2 (N3457, N3439, N3198);
nor NOR4 (N3458, N3435, N1687, N3337, N311);
buf BUF1 (N3459, N3444);
xor XOR2 (N3460, N3454, N743);
or OR4 (N3461, N3450, N1816, N1897, N1836);
or OR3 (N3462, N3457, N2069, N389);
or OR4 (N3463, N3462, N3075, N1623, N2431);
and AND2 (N3464, N3461, N2539);
buf BUF1 (N3465, N3463);
nor NOR3 (N3466, N3460, N2705, N411);
buf BUF1 (N3467, N3453);
nand NAND4 (N3468, N3465, N631, N3090, N2756);
nor NOR3 (N3469, N3456, N996, N1961);
or OR2 (N3470, N3451, N1727);
or OR2 (N3471, N3466, N1765);
nor NOR4 (N3472, N3455, N1052, N16, N3286);
not NOT1 (N3473, N3472);
not NOT1 (N3474, N3458);
xor XOR2 (N3475, N3470, N2667);
buf BUF1 (N3476, N3452);
and AND2 (N3477, N3467, N422);
not NOT1 (N3478, N3475);
and AND3 (N3479, N3471, N1517, N2445);
buf BUF1 (N3480, N3473);
not NOT1 (N3481, N3478);
or OR4 (N3482, N3469, N553, N334, N468);
buf BUF1 (N3483, N3476);
and AND3 (N3484, N3482, N6, N1618);
xor XOR2 (N3485, N3459, N2341);
nand NAND3 (N3486, N3480, N670, N689);
or OR4 (N3487, N3483, N3422, N3335, N3121);
or OR2 (N3488, N3486, N2376);
or OR3 (N3489, N3481, N719, N154);
nand NAND4 (N3490, N3489, N951, N1473, N3012);
xor XOR2 (N3491, N3479, N1569);
not NOT1 (N3492, N3474);
nand NAND4 (N3493, N3491, N2972, N1604, N86);
xor XOR2 (N3494, N3488, N1471);
and AND3 (N3495, N3485, N3033, N2324);
xor XOR2 (N3496, N3484, N2084);
and AND4 (N3497, N3492, N1680, N403, N926);
not NOT1 (N3498, N3494);
buf BUF1 (N3499, N3496);
nand NAND2 (N3500, N3498, N2724);
nand NAND4 (N3501, N3493, N495, N1828, N2654);
nand NAND3 (N3502, N3500, N2, N540);
or OR3 (N3503, N3501, N1404, N883);
nand NAND2 (N3504, N3490, N709);
xor XOR2 (N3505, N3495, N998);
buf BUF1 (N3506, N3487);
xor XOR2 (N3507, N3477, N3108);
and AND4 (N3508, N3505, N377, N1640, N764);
nor NOR3 (N3509, N3499, N1392, N3405);
and AND4 (N3510, N3504, N2813, N1755, N3278);
nand NAND4 (N3511, N3507, N735, N1184, N182);
nand NAND2 (N3512, N3468, N1122);
nor NOR2 (N3513, N3503, N1603);
or OR3 (N3514, N3502, N2072, N3072);
buf BUF1 (N3515, N3511);
nand NAND2 (N3516, N3512, N2598);
xor XOR2 (N3517, N3506, N673);
nor NOR3 (N3518, N3508, N656, N790);
or OR2 (N3519, N3515, N1414);
or OR2 (N3520, N3517, N2520);
buf BUF1 (N3521, N3516);
buf BUF1 (N3522, N3510);
and AND4 (N3523, N3513, N887, N2546, N1947);
buf BUF1 (N3524, N3514);
and AND2 (N3525, N3464, N1967);
and AND2 (N3526, N3518, N1932);
xor XOR2 (N3527, N3526, N1761);
nand NAND4 (N3528, N3524, N2819, N2468, N1822);
xor XOR2 (N3529, N3497, N126);
and AND3 (N3530, N3523, N388, N2854);
or OR2 (N3531, N3525, N699);
not NOT1 (N3532, N3522);
xor XOR2 (N3533, N3529, N2414);
or OR3 (N3534, N3531, N2405, N1675);
not NOT1 (N3535, N3521);
or OR2 (N3536, N3509, N665);
buf BUF1 (N3537, N3528);
or OR2 (N3538, N3534, N1198);
xor XOR2 (N3539, N3533, N3358);
xor XOR2 (N3540, N3532, N1599);
xor XOR2 (N3541, N3535, N159);
not NOT1 (N3542, N3519);
not NOT1 (N3543, N3530);
xor XOR2 (N3544, N3541, N1911);
or OR3 (N3545, N3520, N2468, N87);
xor XOR2 (N3546, N3540, N187);
xor XOR2 (N3547, N3545, N1295);
not NOT1 (N3548, N3546);
nor NOR2 (N3549, N3536, N1265);
nor NOR4 (N3550, N3549, N1340, N1139, N3529);
nand NAND2 (N3551, N3538, N183);
and AND3 (N3552, N3542, N1040, N19);
xor XOR2 (N3553, N3548, N3412);
nand NAND4 (N3554, N3547, N2633, N1075, N2639);
not NOT1 (N3555, N3543);
and AND4 (N3556, N3527, N589, N3525, N1266);
nand NAND4 (N3557, N3553, N2761, N2627, N2303);
or OR4 (N3558, N3556, N514, N1264, N2642);
buf BUF1 (N3559, N3544);
nand NAND2 (N3560, N3557, N2199);
and AND2 (N3561, N3537, N3546);
nor NOR4 (N3562, N3558, N1551, N2074, N593);
xor XOR2 (N3563, N3554, N3014);
and AND2 (N3564, N3562, N144);
and AND3 (N3565, N3550, N1695, N1719);
nor NOR3 (N3566, N3539, N2344, N222);
not NOT1 (N3567, N3551);
and AND2 (N3568, N3560, N3166);
nand NAND4 (N3569, N3568, N2149, N2355, N2713);
nand NAND3 (N3570, N3555, N2640, N962);
not NOT1 (N3571, N3559);
not NOT1 (N3572, N3563);
and AND2 (N3573, N3552, N3375);
buf BUF1 (N3574, N3571);
xor XOR2 (N3575, N3569, N557);
and AND2 (N3576, N3566, N343);
nand NAND2 (N3577, N3574, N2328);
buf BUF1 (N3578, N3573);
buf BUF1 (N3579, N3578);
nand NAND3 (N3580, N3577, N1844, N3533);
nor NOR2 (N3581, N3580, N2335);
nand NAND4 (N3582, N3575, N1559, N629, N3030);
nor NOR4 (N3583, N3582, N1307, N1785, N609);
not NOT1 (N3584, N3564);
nor NOR3 (N3585, N3565, N359, N574);
xor XOR2 (N3586, N3579, N500);
or OR2 (N3587, N3583, N1593);
xor XOR2 (N3588, N3585, N283);
buf BUF1 (N3589, N3586);
nor NOR4 (N3590, N3561, N1731, N1696, N1783);
buf BUF1 (N3591, N3590);
not NOT1 (N3592, N3567);
xor XOR2 (N3593, N3588, N705);
nor NOR2 (N3594, N3591, N2673);
not NOT1 (N3595, N3570);
nand NAND3 (N3596, N3576, N1556, N1443);
nor NOR2 (N3597, N3584, N306);
nor NOR4 (N3598, N3587, N2438, N1664, N71);
xor XOR2 (N3599, N3598, N2470);
or OR2 (N3600, N3581, N142);
nand NAND4 (N3601, N3596, N1636, N3546, N1214);
buf BUF1 (N3602, N3589);
xor XOR2 (N3603, N3572, N1874);
nor NOR4 (N3604, N3602, N338, N893, N2171);
xor XOR2 (N3605, N3597, N1260);
or OR2 (N3606, N3594, N1850);
nand NAND4 (N3607, N3603, N559, N1104, N556);
nor NOR3 (N3608, N3599, N3340, N2437);
nand NAND2 (N3609, N3605, N381);
xor XOR2 (N3610, N3595, N2436);
nand NAND3 (N3611, N3607, N1618, N2055);
nand NAND4 (N3612, N3604, N513, N1764, N1022);
not NOT1 (N3613, N3609);
nor NOR4 (N3614, N3610, N2926, N1111, N2522);
nor NOR3 (N3615, N3614, N2692, N3369);
xor XOR2 (N3616, N3593, N2493);
nand NAND3 (N3617, N3608, N3401, N1648);
nand NAND3 (N3618, N3611, N2107, N2490);
or OR3 (N3619, N3616, N2972, N2569);
nand NAND3 (N3620, N3612, N1697, N3228);
buf BUF1 (N3621, N3619);
nand NAND2 (N3622, N3592, N2736);
and AND2 (N3623, N3617, N3476);
and AND3 (N3624, N3615, N2589, N957);
nand NAND3 (N3625, N3621, N2718, N1628);
nor NOR4 (N3626, N3620, N520, N1308, N2944);
nor NOR2 (N3627, N3601, N498);
xor XOR2 (N3628, N3627, N1762);
buf BUF1 (N3629, N3600);
nand NAND3 (N3630, N3623, N2551, N2205);
buf BUF1 (N3631, N3618);
nand NAND4 (N3632, N3629, N2548, N238, N1999);
or OR4 (N3633, N3613, N2771, N2804, N3130);
buf BUF1 (N3634, N3631);
xor XOR2 (N3635, N3630, N805);
xor XOR2 (N3636, N3632, N803);
and AND2 (N3637, N3622, N3029);
buf BUF1 (N3638, N3624);
nor NOR4 (N3639, N3637, N2896, N2497, N2616);
or OR4 (N3640, N3639, N2095, N3374, N3217);
nor NOR3 (N3641, N3638, N2992, N2764);
nor NOR3 (N3642, N3606, N2950, N1811);
xor XOR2 (N3643, N3635, N116);
buf BUF1 (N3644, N3626);
not NOT1 (N3645, N3634);
not NOT1 (N3646, N3628);
not NOT1 (N3647, N3645);
buf BUF1 (N3648, N3643);
buf BUF1 (N3649, N3648);
buf BUF1 (N3650, N3625);
not NOT1 (N3651, N3649);
nand NAND2 (N3652, N3641, N2308);
nor NOR2 (N3653, N3646, N2481);
nand NAND4 (N3654, N3650, N947, N3161, N267);
and AND2 (N3655, N3654, N742);
or OR3 (N3656, N3644, N933, N2907);
or OR3 (N3657, N3655, N3398, N710);
not NOT1 (N3658, N3657);
nor NOR4 (N3659, N3656, N488, N304, N112);
buf BUF1 (N3660, N3647);
nand NAND2 (N3661, N3659, N2605);
not NOT1 (N3662, N3651);
or OR4 (N3663, N3652, N1992, N1822, N1542);
not NOT1 (N3664, N3653);
nand NAND2 (N3665, N3636, N1951);
and AND3 (N3666, N3662, N377, N421);
nor NOR4 (N3667, N3660, N1420, N1313, N3370);
nor NOR4 (N3668, N3665, N1217, N2862, N3619);
xor XOR2 (N3669, N3668, N1666);
buf BUF1 (N3670, N3667);
nand NAND4 (N3671, N3670, N2296, N1746, N744);
not NOT1 (N3672, N3642);
and AND2 (N3673, N3669, N1286);
nor NOR2 (N3674, N3666, N117);
nand NAND4 (N3675, N3658, N535, N1730, N3277);
and AND2 (N3676, N3661, N335);
xor XOR2 (N3677, N3633, N2565);
nand NAND2 (N3678, N3676, N3189);
nand NAND4 (N3679, N3664, N599, N442, N3599);
xor XOR2 (N3680, N3663, N3298);
nand NAND4 (N3681, N3678, N2913, N1871, N969);
not NOT1 (N3682, N3640);
nand NAND4 (N3683, N3674, N61, N2120, N489);
not NOT1 (N3684, N3671);
or OR2 (N3685, N3675, N1923);
or OR2 (N3686, N3682, N1199);
or OR3 (N3687, N3681, N2042, N781);
or OR3 (N3688, N3677, N904, N3178);
and AND2 (N3689, N3684, N1896);
not NOT1 (N3690, N3672);
or OR2 (N3691, N3679, N2269);
and AND4 (N3692, N3691, N2901, N3169, N3053);
or OR3 (N3693, N3688, N2436, N1658);
nand NAND3 (N3694, N3686, N2438, N2492);
buf BUF1 (N3695, N3689);
or OR4 (N3696, N3694, N84, N349, N3578);
and AND3 (N3697, N3680, N563, N2724);
xor XOR2 (N3698, N3693, N2637);
xor XOR2 (N3699, N3698, N1629);
or OR3 (N3700, N3683, N2843, N2642);
buf BUF1 (N3701, N3696);
nor NOR3 (N3702, N3699, N793, N2178);
buf BUF1 (N3703, N3687);
not NOT1 (N3704, N3673);
nand NAND3 (N3705, N3695, N670, N2566);
nand NAND4 (N3706, N3697, N2431, N372, N3232);
nand NAND3 (N3707, N3692, N32, N1743);
or OR3 (N3708, N3700, N2587, N1935);
or OR2 (N3709, N3704, N877);
buf BUF1 (N3710, N3708);
xor XOR2 (N3711, N3701, N2479);
and AND2 (N3712, N3709, N2981);
nor NOR4 (N3713, N3711, N1587, N3182, N1113);
xor XOR2 (N3714, N3712, N923);
nor NOR4 (N3715, N3690, N1612, N2292, N1799);
xor XOR2 (N3716, N3685, N2428);
or OR3 (N3717, N3713, N1735, N2987);
xor XOR2 (N3718, N3707, N2389);
buf BUF1 (N3719, N3706);
nand NAND4 (N3720, N3703, N877, N3130, N25);
and AND2 (N3721, N3702, N232);
not NOT1 (N3722, N3719);
or OR2 (N3723, N3716, N1066);
nand NAND3 (N3724, N3715, N1397, N1800);
not NOT1 (N3725, N3723);
or OR2 (N3726, N3705, N1160);
or OR2 (N3727, N3726, N3111);
buf BUF1 (N3728, N3717);
buf BUF1 (N3729, N3721);
and AND3 (N3730, N3724, N2251, N2723);
xor XOR2 (N3731, N3727, N2753);
nor NOR4 (N3732, N3714, N611, N1699, N2843);
not NOT1 (N3733, N3720);
not NOT1 (N3734, N3730);
or OR4 (N3735, N3733, N2328, N3095, N2940);
or OR2 (N3736, N3735, N1997);
nand NAND4 (N3737, N3731, N941, N1510, N950);
xor XOR2 (N3738, N3725, N1066);
nor NOR4 (N3739, N3737, N3074, N3350, N3009);
and AND3 (N3740, N3729, N730, N3347);
and AND2 (N3741, N3732, N3623);
buf BUF1 (N3742, N3740);
nand NAND3 (N3743, N3739, N824, N1222);
nand NAND2 (N3744, N3741, N2445);
buf BUF1 (N3745, N3742);
nand NAND3 (N3746, N3745, N505, N3185);
xor XOR2 (N3747, N3722, N15);
buf BUF1 (N3748, N3747);
or OR2 (N3749, N3734, N742);
nor NOR4 (N3750, N3749, N3335, N2301, N2621);
or OR4 (N3751, N3718, N3381, N443, N2841);
xor XOR2 (N3752, N3728, N3241);
nand NAND3 (N3753, N3738, N3655, N671);
and AND3 (N3754, N3751, N2987, N1616);
nand NAND4 (N3755, N3743, N2897, N2922, N1682);
xor XOR2 (N3756, N3748, N168);
buf BUF1 (N3757, N3746);
not NOT1 (N3758, N3736);
or OR2 (N3759, N3750, N2192);
nor NOR4 (N3760, N3759, N2779, N1339, N3661);
not NOT1 (N3761, N3760);
not NOT1 (N3762, N3756);
nand NAND2 (N3763, N3755, N3707);
nor NOR4 (N3764, N3763, N1732, N1521, N602);
and AND4 (N3765, N3762, N2894, N2002, N2795);
or OR4 (N3766, N3757, N52, N2410, N2821);
not NOT1 (N3767, N3765);
not NOT1 (N3768, N3754);
or OR4 (N3769, N3761, N3047, N886, N724);
and AND2 (N3770, N3766, N3469);
xor XOR2 (N3771, N3764, N3035);
not NOT1 (N3772, N3768);
xor XOR2 (N3773, N3770, N3480);
and AND2 (N3774, N3752, N1877);
or OR4 (N3775, N3769, N610, N3555, N167);
not NOT1 (N3776, N3774);
not NOT1 (N3777, N3772);
and AND3 (N3778, N3744, N2206, N3267);
and AND4 (N3779, N3773, N1335, N3420, N1396);
and AND2 (N3780, N3767, N738);
xor XOR2 (N3781, N3776, N1642);
xor XOR2 (N3782, N3753, N1036);
nand NAND2 (N3783, N3710, N3758);
xor XOR2 (N3784, N974, N3065);
and AND4 (N3785, N3771, N2577, N2979, N1310);
or OR2 (N3786, N3782, N302);
xor XOR2 (N3787, N3781, N1655);
nor NOR2 (N3788, N3783, N2196);
xor XOR2 (N3789, N3780, N507);
xor XOR2 (N3790, N3789, N740);
buf BUF1 (N3791, N3786);
nand NAND4 (N3792, N3784, N903, N1104, N2341);
and AND4 (N3793, N3785, N3491, N3134, N288);
or OR4 (N3794, N3775, N117, N2142, N2503);
xor XOR2 (N3795, N3794, N1192);
not NOT1 (N3796, N3778);
nand NAND2 (N3797, N3777, N263);
nand NAND2 (N3798, N3788, N2230);
not NOT1 (N3799, N3792);
buf BUF1 (N3800, N3791);
xor XOR2 (N3801, N3796, N2005);
nor NOR4 (N3802, N3795, N2521, N3480, N340);
nand NAND3 (N3803, N3801, N1671, N2155);
or OR2 (N3804, N3800, N2645);
not NOT1 (N3805, N3797);
and AND2 (N3806, N3805, N1887);
not NOT1 (N3807, N3779);
nand NAND3 (N3808, N3798, N146, N2200);
not NOT1 (N3809, N3803);
nor NOR3 (N3810, N3809, N2967, N2575);
not NOT1 (N3811, N3807);
nand NAND3 (N3812, N3799, N533, N2324);
not NOT1 (N3813, N3802);
xor XOR2 (N3814, N3808, N2268);
nor NOR4 (N3815, N3814, N135, N3143, N24);
nand NAND2 (N3816, N3811, N1179);
xor XOR2 (N3817, N3806, N1475);
not NOT1 (N3818, N3790);
nand NAND2 (N3819, N3810, N861);
not NOT1 (N3820, N3816);
buf BUF1 (N3821, N3818);
or OR2 (N3822, N3820, N589);
and AND2 (N3823, N3787, N763);
not NOT1 (N3824, N3815);
buf BUF1 (N3825, N3822);
nor NOR2 (N3826, N3804, N2508);
xor XOR2 (N3827, N3819, N3425);
nor NOR3 (N3828, N3824, N1238, N1709);
not NOT1 (N3829, N3823);
nor NOR4 (N3830, N3827, N2801, N337, N2447);
nand NAND4 (N3831, N3821, N1330, N2856, N1377);
not NOT1 (N3832, N3825);
and AND2 (N3833, N3829, N2204);
or OR2 (N3834, N3832, N2768);
nand NAND4 (N3835, N3813, N2919, N3647, N2136);
or OR3 (N3836, N3817, N2672, N1465);
and AND3 (N3837, N3834, N809, N3800);
buf BUF1 (N3838, N3828);
not NOT1 (N3839, N3793);
or OR4 (N3840, N3830, N3670, N980, N391);
or OR3 (N3841, N3839, N1847, N1540);
and AND3 (N3842, N3838, N3711, N2110);
buf BUF1 (N3843, N3831);
xor XOR2 (N3844, N3837, N368);
nor NOR4 (N3845, N3844, N1064, N1922, N2336);
nand NAND2 (N3846, N3843, N2662);
nand NAND2 (N3847, N3845, N2884);
and AND4 (N3848, N3840, N3546, N1979, N2877);
and AND3 (N3849, N3842, N1364, N1743);
and AND3 (N3850, N3826, N3660, N3366);
or OR4 (N3851, N3846, N205, N1944, N3593);
nor NOR2 (N3852, N3849, N338);
and AND2 (N3853, N3851, N1556);
nand NAND2 (N3854, N3850, N1067);
nand NAND3 (N3855, N3847, N3495, N45);
and AND4 (N3856, N3835, N1319, N2390, N701);
or OR4 (N3857, N3841, N3756, N3548, N1948);
nor NOR4 (N3858, N3853, N1302, N1898, N1442);
nand NAND4 (N3859, N3812, N397, N1009, N3839);
nor NOR3 (N3860, N3848, N1825, N1106);
not NOT1 (N3861, N3858);
nor NOR4 (N3862, N3859, N2210, N1992, N3734);
nor NOR2 (N3863, N3854, N262);
nor NOR4 (N3864, N3836, N3717, N851, N221);
nor NOR4 (N3865, N3860, N3514, N1047, N2841);
nor NOR3 (N3866, N3863, N2988, N2891);
not NOT1 (N3867, N3864);
xor XOR2 (N3868, N3833, N2229);
or OR3 (N3869, N3856, N2627, N2448);
buf BUF1 (N3870, N3852);
xor XOR2 (N3871, N3867, N904);
or OR2 (N3872, N3866, N3002);
and AND2 (N3873, N3855, N1262);
nand NAND2 (N3874, N3869, N556);
or OR2 (N3875, N3870, N3036);
nand NAND2 (N3876, N3857, N2062);
not NOT1 (N3877, N3876);
buf BUF1 (N3878, N3861);
or OR2 (N3879, N3868, N2293);
not NOT1 (N3880, N3865);
nand NAND2 (N3881, N3880, N984);
buf BUF1 (N3882, N3875);
and AND3 (N3883, N3879, N1329, N1539);
nand NAND2 (N3884, N3871, N2728);
buf BUF1 (N3885, N3862);
nor NOR3 (N3886, N3878, N3597, N3547);
not NOT1 (N3887, N3885);
not NOT1 (N3888, N3883);
or OR4 (N3889, N3884, N410, N2527, N3448);
not NOT1 (N3890, N3877);
or OR3 (N3891, N3874, N363, N2429);
nand NAND3 (N3892, N3889, N2416, N2075);
not NOT1 (N3893, N3890);
nand NAND4 (N3894, N3881, N2662, N2789, N515);
buf BUF1 (N3895, N3893);
and AND2 (N3896, N3886, N3395);
and AND2 (N3897, N3887, N1941);
not NOT1 (N3898, N3897);
or OR2 (N3899, N3898, N3163);
xor XOR2 (N3900, N3888, N868);
nor NOR4 (N3901, N3872, N2705, N2448, N967);
not NOT1 (N3902, N3900);
buf BUF1 (N3903, N3902);
nand NAND2 (N3904, N3899, N1186);
and AND2 (N3905, N3895, N3662);
buf BUF1 (N3906, N3896);
xor XOR2 (N3907, N3882, N1037);
nor NOR4 (N3908, N3906, N2647, N2734, N2836);
nand NAND4 (N3909, N3873, N1952, N2177, N326);
buf BUF1 (N3910, N3905);
nor NOR4 (N3911, N3903, N2674, N2846, N372);
xor XOR2 (N3912, N3908, N1626);
nand NAND4 (N3913, N3912, N2580, N2961, N1774);
xor XOR2 (N3914, N3909, N3763);
and AND3 (N3915, N3914, N2491, N2672);
buf BUF1 (N3916, N3913);
and AND3 (N3917, N3907, N2965, N989);
xor XOR2 (N3918, N3910, N3690);
buf BUF1 (N3919, N3904);
buf BUF1 (N3920, N3915);
buf BUF1 (N3921, N3920);
xor XOR2 (N3922, N3891, N1958);
not NOT1 (N3923, N3922);
xor XOR2 (N3924, N3892, N2194);
xor XOR2 (N3925, N3916, N1915);
nand NAND4 (N3926, N3925, N728, N2688, N2661);
xor XOR2 (N3927, N3919, N2087);
not NOT1 (N3928, N3927);
and AND3 (N3929, N3926, N2976, N2835);
or OR4 (N3930, N3929, N2451, N1886, N83);
not NOT1 (N3931, N3924);
and AND2 (N3932, N3931, N586);
not NOT1 (N3933, N3932);
or OR3 (N3934, N3923, N523, N1431);
buf BUF1 (N3935, N3933);
xor XOR2 (N3936, N3934, N3457);
or OR2 (N3937, N3928, N1487);
not NOT1 (N3938, N3901);
or OR4 (N3939, N3911, N1455, N1301, N3496);
buf BUF1 (N3940, N3894);
or OR3 (N3941, N3918, N2941, N3725);
or OR4 (N3942, N3938, N2393, N3363, N1051);
buf BUF1 (N3943, N3939);
or OR3 (N3944, N3921, N2399, N2554);
xor XOR2 (N3945, N3944, N3593);
not NOT1 (N3946, N3917);
nor NOR2 (N3947, N3941, N623);
not NOT1 (N3948, N3945);
buf BUF1 (N3949, N3946);
nor NOR4 (N3950, N3942, N726, N2223, N3638);
nor NOR4 (N3951, N3947, N2328, N1564, N3090);
nor NOR4 (N3952, N3940, N627, N512, N2430);
buf BUF1 (N3953, N3937);
nand NAND4 (N3954, N3949, N1889, N2158, N1487);
buf BUF1 (N3955, N3954);
nor NOR4 (N3956, N3955, N2691, N3316, N2093);
nand NAND4 (N3957, N3943, N3449, N991, N2586);
not NOT1 (N3958, N3950);
xor XOR2 (N3959, N3952, N677);
nand NAND2 (N3960, N3953, N3148);
or OR2 (N3961, N3957, N2958);
and AND2 (N3962, N3948, N1170);
and AND4 (N3963, N3930, N1875, N2485, N2324);
or OR3 (N3964, N3956, N403, N2115);
nand NAND2 (N3965, N3963, N2804);
buf BUF1 (N3966, N3965);
and AND3 (N3967, N3962, N3114, N36);
not NOT1 (N3968, N3951);
or OR4 (N3969, N3966, N396, N105, N2663);
and AND4 (N3970, N3958, N1106, N1125, N1007);
not NOT1 (N3971, N3935);
buf BUF1 (N3972, N3969);
nor NOR2 (N3973, N3961, N47);
or OR3 (N3974, N3973, N3123, N3858);
not NOT1 (N3975, N3960);
xor XOR2 (N3976, N3971, N1287);
not NOT1 (N3977, N3972);
nor NOR2 (N3978, N3975, N191);
or OR3 (N3979, N3967, N2575, N2233);
xor XOR2 (N3980, N3974, N1415);
xor XOR2 (N3981, N3968, N1807);
nand NAND2 (N3982, N3964, N1598);
not NOT1 (N3983, N3979);
not NOT1 (N3984, N3983);
nand NAND4 (N3985, N3977, N2064, N3069, N2555);
not NOT1 (N3986, N3978);
not NOT1 (N3987, N3970);
and AND3 (N3988, N3984, N3308, N1950);
nor NOR2 (N3989, N3980, N2757);
and AND4 (N3990, N3976, N2429, N3388, N1926);
nor NOR4 (N3991, N3982, N3932, N2846, N2738);
xor XOR2 (N3992, N3989, N2879);
xor XOR2 (N3993, N3990, N2144);
nand NAND3 (N3994, N3988, N2827, N2779);
nor NOR3 (N3995, N3985, N2086, N898);
xor XOR2 (N3996, N3936, N609);
not NOT1 (N3997, N3992);
buf BUF1 (N3998, N3959);
buf BUF1 (N3999, N3998);
not NOT1 (N4000, N3993);
buf BUF1 (N4001, N3994);
nand NAND3 (N4002, N3999, N1173, N2830);
not NOT1 (N4003, N4000);
buf BUF1 (N4004, N3986);
nor NOR4 (N4005, N3987, N56, N766, N707);
buf BUF1 (N4006, N4005);
nand NAND4 (N4007, N3981, N1458, N975, N1758);
nor NOR4 (N4008, N4007, N708, N713, N3023);
buf BUF1 (N4009, N4004);
xor XOR2 (N4010, N3997, N1030);
not NOT1 (N4011, N3991);
buf BUF1 (N4012, N3996);
and AND4 (N4013, N4006, N2435, N1600, N3837);
or OR4 (N4014, N4003, N2235, N99, N860);
not NOT1 (N4015, N4009);
buf BUF1 (N4016, N3995);
and AND2 (N4017, N4002, N2451);
or OR2 (N4018, N4001, N2273);
buf BUF1 (N4019, N4016);
nor NOR4 (N4020, N4015, N1667, N56, N1848);
nor NOR4 (N4021, N4012, N1342, N811, N1552);
nor NOR2 (N4022, N4018, N3976);
xor XOR2 (N4023, N4019, N778);
not NOT1 (N4024, N4017);
xor XOR2 (N4025, N4021, N3317);
and AND3 (N4026, N4022, N1003, N2285);
buf BUF1 (N4027, N4014);
nor NOR2 (N4028, N4026, N3317);
buf BUF1 (N4029, N4008);
and AND3 (N4030, N4025, N3115, N1684);
xor XOR2 (N4031, N4013, N3976);
xor XOR2 (N4032, N4020, N578);
and AND4 (N4033, N4032, N3668, N1259, N1444);
and AND3 (N4034, N4027, N861, N2641);
or OR2 (N4035, N4024, N1119);
or OR2 (N4036, N4034, N711);
and AND2 (N4037, N4029, N2009);
nand NAND4 (N4038, N4023, N3174, N34, N653);
and AND3 (N4039, N4036, N3434, N1698);
and AND3 (N4040, N4037, N1624, N3239);
xor XOR2 (N4041, N4030, N731);
not NOT1 (N4042, N4041);
not NOT1 (N4043, N4039);
nand NAND4 (N4044, N4038, N3062, N3947, N1376);
nand NAND2 (N4045, N4011, N3419);
nor NOR4 (N4046, N4035, N3326, N3046, N810);
not NOT1 (N4047, N4010);
xor XOR2 (N4048, N4040, N490);
or OR2 (N4049, N4042, N939);
buf BUF1 (N4050, N4031);
nand NAND3 (N4051, N4050, N389, N1900);
xor XOR2 (N4052, N4033, N2355);
not NOT1 (N4053, N4045);
or OR2 (N4054, N4044, N1301);
buf BUF1 (N4055, N4052);
xor XOR2 (N4056, N4055, N86);
buf BUF1 (N4057, N4049);
buf BUF1 (N4058, N4057);
nand NAND2 (N4059, N4053, N2678);
buf BUF1 (N4060, N4051);
nor NOR3 (N4061, N4048, N2636, N2791);
and AND3 (N4062, N4058, N2614, N2576);
buf BUF1 (N4063, N4054);
not NOT1 (N4064, N4063);
and AND4 (N4065, N4061, N1570, N59, N1053);
nor NOR4 (N4066, N4065, N3954, N689, N3180);
not NOT1 (N4067, N4046);
nor NOR3 (N4068, N4062, N1634, N1316);
nor NOR4 (N4069, N4064, N652, N1308, N2762);
not NOT1 (N4070, N4060);
and AND3 (N4071, N4028, N3347, N3851);
buf BUF1 (N4072, N4067);
not NOT1 (N4073, N4047);
nand NAND3 (N4074, N4069, N3150, N1758);
not NOT1 (N4075, N4056);
xor XOR2 (N4076, N4043, N2550);
xor XOR2 (N4077, N4075, N2838);
or OR3 (N4078, N4070, N114, N1232);
not NOT1 (N4079, N4068);
and AND3 (N4080, N4071, N412, N2803);
xor XOR2 (N4081, N4066, N284);
or OR2 (N4082, N4080, N3196);
xor XOR2 (N4083, N4079, N1659);
nand NAND2 (N4084, N4072, N2124);
xor XOR2 (N4085, N4073, N2331);
not NOT1 (N4086, N4082);
buf BUF1 (N4087, N4083);
and AND3 (N4088, N4059, N3726, N52);
or OR4 (N4089, N4085, N220, N1926, N1481);
and AND4 (N4090, N4088, N2392, N3154, N2048);
nand NAND3 (N4091, N4077, N1765, N1798);
and AND4 (N4092, N4086, N3531, N3241, N2246);
or OR3 (N4093, N4091, N901, N2738);
buf BUF1 (N4094, N4090);
not NOT1 (N4095, N4076);
and AND2 (N4096, N4094, N1082);
nor NOR2 (N4097, N4095, N4009);
nor NOR4 (N4098, N4092, N2834, N1031, N2169);
buf BUF1 (N4099, N4093);
buf BUF1 (N4100, N4084);
xor XOR2 (N4101, N4098, N4036);
and AND2 (N4102, N4074, N1249);
nand NAND2 (N4103, N4097, N3790);
xor XOR2 (N4104, N4081, N2902);
xor XOR2 (N4105, N4102, N1485);
or OR3 (N4106, N4104, N1371, N3900);
xor XOR2 (N4107, N4105, N338);
and AND3 (N4108, N4103, N3754, N3521);
not NOT1 (N4109, N4078);
or OR4 (N4110, N4109, N2722, N2441, N3830);
buf BUF1 (N4111, N4100);
buf BUF1 (N4112, N4108);
buf BUF1 (N4113, N4107);
or OR2 (N4114, N4087, N2081);
xor XOR2 (N4115, N4089, N1549);
nand NAND3 (N4116, N4112, N2322, N913);
nand NAND3 (N4117, N4116, N3480, N2406);
and AND4 (N4118, N4114, N2634, N3187, N953);
xor XOR2 (N4119, N4106, N2508);
buf BUF1 (N4120, N4115);
or OR2 (N4121, N4096, N3234);
buf BUF1 (N4122, N4113);
or OR3 (N4123, N4110, N3392, N2716);
nor NOR3 (N4124, N4119, N168, N2393);
or OR2 (N4125, N4099, N3601);
nand NAND3 (N4126, N4101, N4, N410);
nor NOR4 (N4127, N4118, N2717, N3642, N1974);
nand NAND3 (N4128, N4117, N3283, N1252);
not NOT1 (N4129, N4122);
nand NAND3 (N4130, N4129, N1154, N3551);
xor XOR2 (N4131, N4126, N1607);
buf BUF1 (N4132, N4111);
xor XOR2 (N4133, N4128, N2488);
or OR3 (N4134, N4121, N2381, N923);
xor XOR2 (N4135, N4130, N2277);
xor XOR2 (N4136, N4134, N3349);
not NOT1 (N4137, N4131);
or OR3 (N4138, N4135, N2711, N2166);
nor NOR3 (N4139, N4136, N1505, N1231);
xor XOR2 (N4140, N4123, N3242);
or OR3 (N4141, N4140, N1503, N1441);
xor XOR2 (N4142, N4124, N1776);
not NOT1 (N4143, N4120);
buf BUF1 (N4144, N4141);
nor NOR4 (N4145, N4127, N3868, N3445, N2337);
nor NOR2 (N4146, N4143, N2209);
and AND2 (N4147, N4145, N444);
nor NOR2 (N4148, N4142, N2268);
buf BUF1 (N4149, N4148);
nor NOR4 (N4150, N4125, N248, N1156, N1840);
buf BUF1 (N4151, N4149);
buf BUF1 (N4152, N4137);
or OR2 (N4153, N4151, N3934);
buf BUF1 (N4154, N4138);
nor NOR4 (N4155, N4132, N2587, N2029, N2455);
buf BUF1 (N4156, N4139);
nor NOR2 (N4157, N4154, N4021);
nand NAND4 (N4158, N4133, N2982, N264, N2413);
not NOT1 (N4159, N4158);
not NOT1 (N4160, N4147);
and AND3 (N4161, N4159, N1181, N3847);
nor NOR2 (N4162, N4157, N3860);
nand NAND4 (N4163, N4144, N3793, N1164, N428);
or OR3 (N4164, N4153, N2623, N307);
buf BUF1 (N4165, N4146);
and AND4 (N4166, N4156, N3438, N2598, N1968);
xor XOR2 (N4167, N4161, N2626);
not NOT1 (N4168, N4162);
not NOT1 (N4169, N4167);
nand NAND3 (N4170, N4150, N299, N2369);
and AND4 (N4171, N4155, N3342, N2122, N2084);
nor NOR3 (N4172, N4163, N2919, N2983);
not NOT1 (N4173, N4164);
and AND4 (N4174, N4171, N2253, N2384, N3415);
and AND2 (N4175, N4174, N1535);
nor NOR4 (N4176, N4152, N139, N1955, N3088);
not NOT1 (N4177, N4175);
and AND2 (N4178, N4160, N1184);
or OR2 (N4179, N4165, N636);
buf BUF1 (N4180, N4173);
not NOT1 (N4181, N4169);
not NOT1 (N4182, N4178);
nor NOR3 (N4183, N4166, N1838, N1890);
nor NOR4 (N4184, N4181, N2326, N2374, N1202);
and AND4 (N4185, N4182, N3909, N3843, N2980);
and AND3 (N4186, N4179, N1522, N1571);
and AND2 (N4187, N4177, N1848);
nand NAND3 (N4188, N4176, N585, N3315);
not NOT1 (N4189, N4180);
or OR3 (N4190, N4187, N1202, N1890);
buf BUF1 (N4191, N4170);
and AND3 (N4192, N4188, N2511, N3662);
and AND4 (N4193, N4172, N4023, N3055, N3693);
nand NAND3 (N4194, N4186, N2169, N251);
buf BUF1 (N4195, N4168);
or OR2 (N4196, N4191, N1238);
and AND2 (N4197, N4194, N3175);
and AND3 (N4198, N4195, N3962, N49);
or OR4 (N4199, N4190, N294, N2205, N2095);
not NOT1 (N4200, N4183);
xor XOR2 (N4201, N4196, N2130);
xor XOR2 (N4202, N4192, N827);
and AND2 (N4203, N4184, N3609);
nor NOR2 (N4204, N4202, N535);
nand NAND2 (N4205, N4189, N1282);
and AND4 (N4206, N4197, N928, N930, N3397);
xor XOR2 (N4207, N4198, N3775);
buf BUF1 (N4208, N4199);
buf BUF1 (N4209, N4205);
nand NAND2 (N4210, N4208, N608);
buf BUF1 (N4211, N4209);
buf BUF1 (N4212, N4207);
nand NAND2 (N4213, N4206, N634);
and AND3 (N4214, N4203, N3926, N1664);
buf BUF1 (N4215, N4185);
buf BUF1 (N4216, N4211);
and AND2 (N4217, N4214, N2966);
or OR3 (N4218, N4216, N1857, N2057);
buf BUF1 (N4219, N4217);
or OR3 (N4220, N4212, N2740, N41);
xor XOR2 (N4221, N4213, N2966);
xor XOR2 (N4222, N4221, N2505);
nor NOR2 (N4223, N4215, N3512);
not NOT1 (N4224, N4218);
xor XOR2 (N4225, N4210, N3800);
nand NAND3 (N4226, N4193, N2449, N137);
nand NAND4 (N4227, N4201, N2722, N889, N2880);
and AND2 (N4228, N4223, N602);
or OR2 (N4229, N4227, N3222);
nand NAND3 (N4230, N4204, N1675, N4129);
nor NOR2 (N4231, N4222, N2939);
not NOT1 (N4232, N4224);
buf BUF1 (N4233, N4220);
buf BUF1 (N4234, N4225);
not NOT1 (N4235, N4232);
or OR4 (N4236, N4229, N2009, N1131, N2034);
buf BUF1 (N4237, N4219);
not NOT1 (N4238, N4231);
nand NAND4 (N4239, N4233, N689, N3854, N1305);
or OR4 (N4240, N4237, N2192, N212, N3208);
not NOT1 (N4241, N4235);
nor NOR2 (N4242, N4226, N2020);
and AND4 (N4243, N4242, N2354, N4210, N4177);
or OR3 (N4244, N4241, N1366, N1474);
buf BUF1 (N4245, N4239);
buf BUF1 (N4246, N4236);
nor NOR4 (N4247, N4228, N706, N28, N1376);
xor XOR2 (N4248, N4240, N3649);
buf BUF1 (N4249, N4234);
nor NOR4 (N4250, N4243, N4139, N897, N3254);
nor NOR4 (N4251, N4244, N2292, N2604, N877);
nand NAND3 (N4252, N4238, N2039, N3500);
nand NAND3 (N4253, N4245, N344, N4117);
nand NAND2 (N4254, N4246, N865);
xor XOR2 (N4255, N4249, N625);
and AND3 (N4256, N4230, N1572, N2464);
not NOT1 (N4257, N4247);
or OR3 (N4258, N4257, N1780, N3107);
and AND2 (N4259, N4255, N510);
nor NOR2 (N4260, N4254, N3409);
nor NOR2 (N4261, N4251, N1743);
not NOT1 (N4262, N4200);
not NOT1 (N4263, N4259);
xor XOR2 (N4264, N4263, N133);
or OR2 (N4265, N4250, N3274);
not NOT1 (N4266, N4253);
nor NOR4 (N4267, N4260, N199, N1, N321);
not NOT1 (N4268, N4264);
or OR2 (N4269, N4258, N1596);
and AND4 (N4270, N4265, N788, N1409, N3106);
not NOT1 (N4271, N4270);
not NOT1 (N4272, N4252);
buf BUF1 (N4273, N4266);
and AND4 (N4274, N4267, N552, N32, N1967);
and AND3 (N4275, N4273, N2500, N3459);
not NOT1 (N4276, N4271);
nand NAND2 (N4277, N4261, N395);
nor NOR4 (N4278, N4272, N1205, N355, N314);
buf BUF1 (N4279, N4269);
xor XOR2 (N4280, N4275, N3862);
or OR3 (N4281, N4248, N3574, N918);
nand NAND3 (N4282, N4268, N3199, N268);
xor XOR2 (N4283, N4274, N3472);
or OR2 (N4284, N4256, N3942);
or OR3 (N4285, N4276, N927, N1236);
xor XOR2 (N4286, N4277, N1398);
buf BUF1 (N4287, N4262);
nor NOR3 (N4288, N4280, N3226, N965);
buf BUF1 (N4289, N4279);
nor NOR3 (N4290, N4281, N3253, N3507);
or OR3 (N4291, N4286, N3731, N3274);
not NOT1 (N4292, N4284);
xor XOR2 (N4293, N4278, N451);
and AND2 (N4294, N4292, N4114);
nor NOR4 (N4295, N4282, N2438, N3359, N3177);
or OR4 (N4296, N4289, N4228, N3186, N3310);
nand NAND3 (N4297, N4293, N1082, N933);
nand NAND2 (N4298, N4288, N2607);
xor XOR2 (N4299, N4290, N584);
not NOT1 (N4300, N4291);
or OR2 (N4301, N4296, N2878);
xor XOR2 (N4302, N4287, N3794);
xor XOR2 (N4303, N4283, N4054);
nand NAND2 (N4304, N4301, N1106);
xor XOR2 (N4305, N4304, N2880);
nand NAND4 (N4306, N4294, N2313, N892, N2436);
nor NOR3 (N4307, N4300, N1424, N3136);
nor NOR4 (N4308, N4307, N2191, N877, N154);
nand NAND2 (N4309, N4297, N3252);
nor NOR3 (N4310, N4303, N1675, N446);
xor XOR2 (N4311, N4299, N919);
and AND4 (N4312, N4309, N3535, N2149, N1830);
or OR2 (N4313, N4302, N374);
buf BUF1 (N4314, N4306);
nand NAND4 (N4315, N4310, N403, N567, N243);
or OR4 (N4316, N4298, N1301, N101, N1324);
not NOT1 (N4317, N4314);
and AND4 (N4318, N4311, N635, N1220, N814);
nand NAND3 (N4319, N4285, N1601, N582);
xor XOR2 (N4320, N4295, N101);
nor NOR4 (N4321, N4319, N4162, N2542, N3746);
buf BUF1 (N4322, N4312);
buf BUF1 (N4323, N4315);
buf BUF1 (N4324, N4318);
xor XOR2 (N4325, N4313, N2740);
not NOT1 (N4326, N4308);
nand NAND2 (N4327, N4317, N592);
nor NOR3 (N4328, N4322, N3627, N3579);
not NOT1 (N4329, N4325);
nand NAND4 (N4330, N4328, N2449, N4196, N2879);
not NOT1 (N4331, N4326);
and AND2 (N4332, N4305, N3810);
buf BUF1 (N4333, N4329);
and AND2 (N4334, N4316, N2097);
nor NOR4 (N4335, N4334, N3715, N120, N1258);
nor NOR2 (N4336, N4324, N629);
buf BUF1 (N4337, N4335);
not NOT1 (N4338, N4332);
nand NAND3 (N4339, N4327, N3448, N86);
buf BUF1 (N4340, N4323);
and AND3 (N4341, N4320, N3422, N2329);
not NOT1 (N4342, N4330);
buf BUF1 (N4343, N4336);
nand NAND4 (N4344, N4343, N497, N2827, N3776);
nor NOR4 (N4345, N4341, N4207, N2497, N995);
not NOT1 (N4346, N4339);
nand NAND2 (N4347, N4331, N1607);
buf BUF1 (N4348, N4340);
or OR3 (N4349, N4321, N3381, N521);
nand NAND4 (N4350, N4337, N418, N1367, N552);
or OR3 (N4351, N4349, N1694, N3503);
or OR3 (N4352, N4338, N3188, N1721);
xor XOR2 (N4353, N4342, N2750);
nand NAND2 (N4354, N4348, N645);
buf BUF1 (N4355, N4352);
nor NOR4 (N4356, N4354, N592, N443, N3500);
xor XOR2 (N4357, N4333, N1458);
nor NOR4 (N4358, N4356, N3260, N1503, N3013);
and AND4 (N4359, N4353, N3466, N1213, N49);
buf BUF1 (N4360, N4344);
xor XOR2 (N4361, N4359, N3938);
and AND2 (N4362, N4351, N3916);
nand NAND3 (N4363, N4362, N2957, N371);
or OR2 (N4364, N4345, N4239);
nand NAND3 (N4365, N4347, N416, N3124);
or OR3 (N4366, N4364, N2035, N511);
xor XOR2 (N4367, N4346, N486);
and AND3 (N4368, N4365, N21, N216);
nor NOR4 (N4369, N4350, N4191, N567, N727);
nand NAND3 (N4370, N4367, N928, N3051);
buf BUF1 (N4371, N4355);
buf BUF1 (N4372, N4357);
and AND3 (N4373, N4360, N4002, N3640);
or OR3 (N4374, N4369, N252, N3984);
xor XOR2 (N4375, N4368, N1364);
nor NOR4 (N4376, N4366, N2395, N606, N2168);
or OR4 (N4377, N4373, N4016, N2894, N1356);
or OR4 (N4378, N4377, N1551, N825, N3585);
not NOT1 (N4379, N4363);
buf BUF1 (N4380, N4361);
xor XOR2 (N4381, N4371, N2483);
xor XOR2 (N4382, N4370, N3121);
nor NOR3 (N4383, N4374, N1928, N2188);
and AND2 (N4384, N4358, N3066);
not NOT1 (N4385, N4378);
xor XOR2 (N4386, N4383, N333);
or OR4 (N4387, N4382, N2771, N1015, N3916);
nor NOR3 (N4388, N4386, N1214, N1570);
xor XOR2 (N4389, N4379, N1883);
nor NOR4 (N4390, N4381, N2418, N83, N1625);
not NOT1 (N4391, N4390);
and AND3 (N4392, N4380, N2763, N4081);
not NOT1 (N4393, N4387);
buf BUF1 (N4394, N4391);
not NOT1 (N4395, N4394);
nand NAND2 (N4396, N4393, N3219);
buf BUF1 (N4397, N4389);
and AND3 (N4398, N4372, N3998, N778);
nor NOR4 (N4399, N4397, N2719, N2674, N48);
not NOT1 (N4400, N4392);
not NOT1 (N4401, N4388);
not NOT1 (N4402, N4399);
xor XOR2 (N4403, N4385, N4335);
nand NAND4 (N4404, N4395, N1273, N606, N4217);
or OR4 (N4405, N4384, N4227, N3774, N3301);
buf BUF1 (N4406, N4405);
buf BUF1 (N4407, N4406);
and AND2 (N4408, N4400, N2610);
or OR3 (N4409, N4404, N1645, N1572);
and AND2 (N4410, N4396, N3408);
xor XOR2 (N4411, N4407, N916);
xor XOR2 (N4412, N4398, N2718);
nor NOR4 (N4413, N4376, N347, N26, N3689);
and AND3 (N4414, N4375, N2350, N414);
or OR4 (N4415, N4413, N2981, N4079, N1569);
and AND4 (N4416, N4412, N2065, N4018, N250);
xor XOR2 (N4417, N4415, N3740);
buf BUF1 (N4418, N4403);
nand NAND2 (N4419, N4416, N2833);
or OR4 (N4420, N4401, N1160, N2607, N2829);
or OR3 (N4421, N4402, N1707, N3987);
and AND2 (N4422, N4408, N1681);
or OR3 (N4423, N4417, N3601, N149);
nand NAND3 (N4424, N4419, N31, N3244);
xor XOR2 (N4425, N4423, N2508);
buf BUF1 (N4426, N4425);
or OR4 (N4427, N4410, N4295, N921, N4124);
and AND3 (N4428, N4418, N4076, N3682);
xor XOR2 (N4429, N4414, N1013);
not NOT1 (N4430, N4429);
nand NAND2 (N4431, N4420, N1403);
nand NAND2 (N4432, N4409, N1891);
and AND2 (N4433, N4421, N629);
or OR3 (N4434, N4411, N4098, N151);
not NOT1 (N4435, N4432);
nand NAND4 (N4436, N4434, N1046, N1786, N1839);
nand NAND4 (N4437, N4436, N3099, N149, N3495);
not NOT1 (N4438, N4428);
nand NAND3 (N4439, N4438, N4418, N63);
xor XOR2 (N4440, N4435, N2680);
nand NAND4 (N4441, N4440, N3459, N726, N837);
nor NOR3 (N4442, N4437, N2580, N3282);
buf BUF1 (N4443, N4441);
nor NOR3 (N4444, N4422, N4425, N2416);
not NOT1 (N4445, N4443);
and AND3 (N4446, N4442, N1896, N1192);
nand NAND3 (N4447, N4431, N4231, N92);
nand NAND4 (N4448, N4426, N1697, N1848, N2584);
nand NAND4 (N4449, N4448, N2840, N4012, N2730);
nand NAND3 (N4450, N4433, N3082, N2468);
not NOT1 (N4451, N4427);
or OR4 (N4452, N4447, N1023, N2893, N3296);
not NOT1 (N4453, N4444);
and AND2 (N4454, N4445, N808);
nand NAND3 (N4455, N4424, N4199, N4230);
xor XOR2 (N4456, N4439, N3187);
buf BUF1 (N4457, N4450);
xor XOR2 (N4458, N4457, N2098);
not NOT1 (N4459, N4453);
or OR2 (N4460, N4456, N1837);
or OR2 (N4461, N4454, N4236);
nand NAND3 (N4462, N4449, N2676, N3086);
nand NAND3 (N4463, N4459, N3127, N4090);
xor XOR2 (N4464, N4446, N1616);
and AND2 (N4465, N4455, N146);
or OR3 (N4466, N4451, N4411, N4187);
buf BUF1 (N4467, N4463);
nand NAND4 (N4468, N4466, N814, N1484, N3386);
or OR3 (N4469, N4461, N781, N1167);
xor XOR2 (N4470, N4460, N1365);
nor NOR2 (N4471, N4469, N1126);
buf BUF1 (N4472, N4430);
xor XOR2 (N4473, N4470, N1065);
nor NOR3 (N4474, N4471, N1936, N1753);
xor XOR2 (N4475, N4458, N4336);
nand NAND3 (N4476, N4465, N2323, N694);
or OR3 (N4477, N4464, N362, N3755);
buf BUF1 (N4478, N4473);
nand NAND3 (N4479, N4478, N2929, N4305);
nand NAND2 (N4480, N4472, N2021);
buf BUF1 (N4481, N4477);
not NOT1 (N4482, N4480);
xor XOR2 (N4483, N4462, N80);
nand NAND4 (N4484, N4467, N926, N2075, N3416);
or OR3 (N4485, N4484, N4227, N2252);
buf BUF1 (N4486, N4452);
nor NOR3 (N4487, N4485, N2845, N3449);
buf BUF1 (N4488, N4483);
xor XOR2 (N4489, N4482, N3477);
and AND2 (N4490, N4488, N1214);
not NOT1 (N4491, N4487);
nand NAND4 (N4492, N4481, N3390, N3605, N3857);
not NOT1 (N4493, N4476);
xor XOR2 (N4494, N4486, N2493);
nor NOR4 (N4495, N4468, N4289, N1181, N2462);
nor NOR4 (N4496, N4490, N554, N589, N3798);
nor NOR4 (N4497, N4475, N4476, N3835, N459);
buf BUF1 (N4498, N4497);
nor NOR3 (N4499, N4494, N4302, N3106);
and AND4 (N4500, N4493, N4048, N1586, N1098);
nand NAND4 (N4501, N4496, N2454, N249, N3423);
and AND3 (N4502, N4474, N3643, N3133);
xor XOR2 (N4503, N4492, N1304);
not NOT1 (N4504, N4495);
xor XOR2 (N4505, N4502, N1561);
or OR4 (N4506, N4499, N146, N414, N3873);
and AND4 (N4507, N4501, N2959, N1873, N3268);
and AND4 (N4508, N4500, N2920, N4473, N4344);
xor XOR2 (N4509, N4508, N2822);
or OR3 (N4510, N4491, N3380, N1527);
not NOT1 (N4511, N4503);
or OR4 (N4512, N4507, N1898, N1589, N1783);
xor XOR2 (N4513, N4510, N4486);
buf BUF1 (N4514, N4505);
nor NOR3 (N4515, N4504, N2973, N2696);
or OR2 (N4516, N4512, N290);
or OR4 (N4517, N4509, N3112, N3939, N1317);
and AND4 (N4518, N4515, N3543, N3227, N1635);
not NOT1 (N4519, N4506);
nand NAND4 (N4520, N4489, N4514, N744, N263);
buf BUF1 (N4521, N1498);
or OR3 (N4522, N4517, N2897, N2124);
nand NAND4 (N4523, N4511, N2190, N3959, N1583);
not NOT1 (N4524, N4519);
nor NOR2 (N4525, N4479, N2638);
buf BUF1 (N4526, N4513);
nand NAND4 (N4527, N4526, N145, N1297, N355);
nand NAND2 (N4528, N4521, N11);
buf BUF1 (N4529, N4523);
or OR3 (N4530, N4522, N866, N1584);
or OR2 (N4531, N4528, N2857);
nor NOR4 (N4532, N4520, N1211, N301, N4076);
not NOT1 (N4533, N4529);
buf BUF1 (N4534, N4527);
nor NOR2 (N4535, N4532, N916);
nor NOR3 (N4536, N4518, N2873, N3971);
buf BUF1 (N4537, N4530);
xor XOR2 (N4538, N4531, N575);
not NOT1 (N4539, N4538);
or OR4 (N4540, N4537, N3453, N2440, N3085);
or OR3 (N4541, N4534, N3440, N2877);
buf BUF1 (N4542, N4536);
xor XOR2 (N4543, N4541, N4394);
not NOT1 (N4544, N4535);
nand NAND2 (N4545, N4539, N4157);
and AND2 (N4546, N4525, N1031);
not NOT1 (N4547, N4524);
nor NOR3 (N4548, N4546, N3975, N3613);
or OR4 (N4549, N4548, N2709, N3056, N1097);
not NOT1 (N4550, N4547);
nor NOR4 (N4551, N4533, N3429, N1133, N1263);
or OR2 (N4552, N4544, N1819);
xor XOR2 (N4553, N4551, N1375);
nor NOR2 (N4554, N4540, N2268);
nor NOR2 (N4555, N4542, N1942);
buf BUF1 (N4556, N4549);
xor XOR2 (N4557, N4554, N3127);
nand NAND3 (N4558, N4545, N4036, N1550);
or OR3 (N4559, N4555, N1566, N1183);
nand NAND3 (N4560, N4557, N4529, N3724);
or OR3 (N4561, N4543, N2860, N3702);
buf BUF1 (N4562, N4560);
or OR2 (N4563, N4559, N2818);
nand NAND3 (N4564, N4498, N1991, N682);
nand NAND3 (N4565, N4561, N3630, N1062);
nand NAND4 (N4566, N4516, N2597, N4471, N2201);
or OR3 (N4567, N4558, N1897, N4331);
buf BUF1 (N4568, N4566);
or OR4 (N4569, N4556, N1558, N1380, N4047);
and AND4 (N4570, N4569, N1330, N3832, N4529);
buf BUF1 (N4571, N4550);
xor XOR2 (N4572, N4565, N4483);
not NOT1 (N4573, N4568);
buf BUF1 (N4574, N4571);
nand NAND4 (N4575, N4552, N1924, N1467, N1224);
and AND3 (N4576, N4567, N483, N3847);
nor NOR2 (N4577, N4563, N3383);
and AND2 (N4578, N4576, N2404);
xor XOR2 (N4579, N4562, N1797);
not NOT1 (N4580, N4578);
not NOT1 (N4581, N4579);
xor XOR2 (N4582, N4572, N4571);
or OR2 (N4583, N4580, N1825);
not NOT1 (N4584, N4577);
and AND3 (N4585, N4583, N4082, N3235);
not NOT1 (N4586, N4582);
nand NAND3 (N4587, N4574, N969, N3204);
and AND4 (N4588, N4553, N4056, N4347, N4184);
nand NAND2 (N4589, N4588, N2617);
and AND3 (N4590, N4564, N959, N3052);
nor NOR3 (N4591, N4585, N2084, N4224);
nor NOR4 (N4592, N4584, N1484, N2430, N356);
nor NOR2 (N4593, N4590, N580);
or OR4 (N4594, N4581, N2917, N2974, N2768);
nor NOR4 (N4595, N4591, N3079, N2611, N1565);
not NOT1 (N4596, N4570);
nand NAND3 (N4597, N4593, N3520, N1859);
and AND3 (N4598, N4573, N401, N352);
buf BUF1 (N4599, N4598);
or OR2 (N4600, N4599, N1344);
buf BUF1 (N4601, N4587);
buf BUF1 (N4602, N4575);
nand NAND2 (N4603, N4597, N558);
buf BUF1 (N4604, N4596);
not NOT1 (N4605, N4601);
nor NOR3 (N4606, N4586, N3107, N3270);
nor NOR3 (N4607, N4594, N2105, N1005);
nand NAND3 (N4608, N4604, N3828, N405);
and AND4 (N4609, N4608, N1926, N987, N2842);
or OR3 (N4610, N4603, N2507, N4447);
nor NOR2 (N4611, N4609, N1238);
xor XOR2 (N4612, N4611, N3924);
buf BUF1 (N4613, N4600);
buf BUF1 (N4614, N4592);
or OR4 (N4615, N4610, N11, N3522, N1211);
xor XOR2 (N4616, N4605, N4425);
or OR4 (N4617, N4606, N3565, N2290, N3563);
and AND4 (N4618, N4614, N3054, N1520, N3820);
xor XOR2 (N4619, N4612, N4442);
buf BUF1 (N4620, N4619);
buf BUF1 (N4621, N4617);
xor XOR2 (N4622, N4589, N3346);
or OR4 (N4623, N4615, N1430, N4301, N2824);
nand NAND2 (N4624, N4621, N4447);
and AND3 (N4625, N4624, N1939, N901);
not NOT1 (N4626, N4602);
xor XOR2 (N4627, N4620, N3801);
or OR3 (N4628, N4622, N3190, N1499);
xor XOR2 (N4629, N4595, N217);
and AND2 (N4630, N4626, N555);
nor NOR2 (N4631, N4629, N3758);
buf BUF1 (N4632, N4613);
nand NAND4 (N4633, N4607, N3481, N4126, N2435);
nand NAND2 (N4634, N4618, N2882);
and AND2 (N4635, N4632, N928);
not NOT1 (N4636, N4634);
not NOT1 (N4637, N4625);
buf BUF1 (N4638, N4623);
or OR2 (N4639, N4635, N2989);
buf BUF1 (N4640, N4636);
or OR4 (N4641, N4640, N1002, N3838, N2531);
nor NOR3 (N4642, N4639, N4541, N4382);
or OR2 (N4643, N4637, N2208);
nand NAND3 (N4644, N4631, N4374, N4209);
buf BUF1 (N4645, N4616);
or OR4 (N4646, N4633, N1076, N2813, N2100);
nand NAND2 (N4647, N4646, N2514);
and AND2 (N4648, N4644, N1645);
or OR4 (N4649, N4648, N1710, N1218, N981);
nor NOR2 (N4650, N4627, N1521);
nor NOR3 (N4651, N4643, N1871, N748);
nor NOR3 (N4652, N4642, N1600, N4112);
buf BUF1 (N4653, N4652);
nor NOR4 (N4654, N4649, N4437, N483, N4146);
nor NOR4 (N4655, N4645, N4650, N3468, N502);
or OR4 (N4656, N4049, N1445, N3039, N2507);
nand NAND4 (N4657, N4656, N4104, N4513, N120);
or OR3 (N4658, N4628, N1327, N2342);
nor NOR3 (N4659, N4654, N2975, N3630);
nor NOR2 (N4660, N4638, N2846);
or OR4 (N4661, N4630, N4246, N1561, N3620);
nor NOR4 (N4662, N4655, N4412, N1785, N3533);
nand NAND3 (N4663, N4662, N4017, N1931);
nand NAND3 (N4664, N4653, N277, N1504);
nor NOR4 (N4665, N4657, N3143, N4132, N470);
nand NAND3 (N4666, N4663, N2175, N1571);
not NOT1 (N4667, N4665);
xor XOR2 (N4668, N4659, N283);
nor NOR4 (N4669, N4667, N3399, N321, N3494);
buf BUF1 (N4670, N4669);
not NOT1 (N4671, N4666);
buf BUF1 (N4672, N4668);
nor NOR2 (N4673, N4664, N834);
buf BUF1 (N4674, N4673);
or OR3 (N4675, N4647, N2295, N837);
xor XOR2 (N4676, N4672, N4009);
buf BUF1 (N4677, N4676);
nand NAND3 (N4678, N4658, N2514, N3770);
nor NOR3 (N4679, N4677, N649, N1775);
nand NAND2 (N4680, N4651, N271);
not NOT1 (N4681, N4670);
nand NAND4 (N4682, N4674, N2370, N392, N2157);
or OR3 (N4683, N4682, N4114, N2993);
nor NOR2 (N4684, N4671, N2926);
or OR2 (N4685, N4681, N1781);
not NOT1 (N4686, N4683);
buf BUF1 (N4687, N4661);
or OR4 (N4688, N4685, N1589, N3889, N3509);
nor NOR4 (N4689, N4678, N606, N4381, N3042);
xor XOR2 (N4690, N4689, N3139);
not NOT1 (N4691, N4680);
and AND3 (N4692, N4641, N4637, N3106);
buf BUF1 (N4693, N4660);
or OR2 (N4694, N4686, N3210);
not NOT1 (N4695, N4694);
xor XOR2 (N4696, N4690, N4140);
nor NOR3 (N4697, N4684, N3018, N2510);
or OR3 (N4698, N4693, N2289, N3041);
nor NOR3 (N4699, N4688, N4682, N2104);
xor XOR2 (N4700, N4695, N2572);
and AND4 (N4701, N4696, N3257, N3266, N701);
xor XOR2 (N4702, N4698, N3657);
not NOT1 (N4703, N4697);
or OR4 (N4704, N4691, N1509, N2002, N2545);
nand NAND3 (N4705, N4702, N252, N745);
not NOT1 (N4706, N4703);
xor XOR2 (N4707, N4706, N3722);
buf BUF1 (N4708, N4679);
nand NAND2 (N4709, N4700, N2163);
buf BUF1 (N4710, N4692);
not NOT1 (N4711, N4709);
or OR4 (N4712, N4699, N3530, N2255, N4178);
nand NAND2 (N4713, N4675, N3965);
nor NOR2 (N4714, N4701, N2173);
nand NAND4 (N4715, N4714, N1414, N1852, N1574);
nor NOR3 (N4716, N4708, N4371, N698);
not NOT1 (N4717, N4711);
or OR3 (N4718, N4713, N2967, N3480);
buf BUF1 (N4719, N4715);
buf BUF1 (N4720, N4716);
xor XOR2 (N4721, N4704, N4094);
xor XOR2 (N4722, N4687, N417);
nor NOR3 (N4723, N4719, N2635, N1011);
not NOT1 (N4724, N4710);
not NOT1 (N4725, N4721);
buf BUF1 (N4726, N4718);
and AND4 (N4727, N4725, N2771, N1407, N1268);
buf BUF1 (N4728, N4707);
nand NAND2 (N4729, N4726, N819);
not NOT1 (N4730, N4717);
and AND3 (N4731, N4724, N322, N3105);
nand NAND2 (N4732, N4730, N2469);
not NOT1 (N4733, N4705);
nand NAND4 (N4734, N4723, N1557, N2939, N2284);
or OR2 (N4735, N4731, N1174);
or OR3 (N4736, N4720, N801, N2886);
not NOT1 (N4737, N4728);
and AND3 (N4738, N4712, N1283, N3006);
and AND4 (N4739, N4733, N2133, N3003, N1841);
buf BUF1 (N4740, N4722);
nand NAND2 (N4741, N4737, N3342);
xor XOR2 (N4742, N4738, N4536);
xor XOR2 (N4743, N4735, N734);
nand NAND3 (N4744, N4742, N4526, N3903);
or OR2 (N4745, N4736, N2155);
and AND4 (N4746, N4744, N302, N3144, N3157);
xor XOR2 (N4747, N4727, N383);
buf BUF1 (N4748, N4743);
buf BUF1 (N4749, N4729);
buf BUF1 (N4750, N4741);
not NOT1 (N4751, N4746);
nand NAND2 (N4752, N4751, N1775);
buf BUF1 (N4753, N4734);
or OR3 (N4754, N4750, N832, N4190);
nor NOR2 (N4755, N4748, N9);
buf BUF1 (N4756, N4740);
or OR2 (N4757, N4755, N2216);
not NOT1 (N4758, N4739);
xor XOR2 (N4759, N4758, N2032);
nand NAND3 (N4760, N4753, N2818, N666);
nor NOR3 (N4761, N4752, N2869, N174);
or OR2 (N4762, N4759, N4683);
buf BUF1 (N4763, N4762);
not NOT1 (N4764, N4749);
or OR3 (N4765, N4732, N494, N4729);
nor NOR2 (N4766, N4747, N3779);
xor XOR2 (N4767, N4745, N4599);
xor XOR2 (N4768, N4754, N1980);
xor XOR2 (N4769, N4765, N289);
and AND4 (N4770, N4764, N2834, N1814, N4437);
or OR2 (N4771, N4770, N2567);
nor NOR3 (N4772, N4771, N2087, N3883);
buf BUF1 (N4773, N4760);
not NOT1 (N4774, N4772);
and AND2 (N4775, N4773, N1488);
not NOT1 (N4776, N4763);
and AND3 (N4777, N4761, N235, N2037);
or OR4 (N4778, N4776, N665, N358, N3552);
not NOT1 (N4779, N4766);
or OR2 (N4780, N4757, N742);
not NOT1 (N4781, N4767);
xor XOR2 (N4782, N4775, N1364);
nor NOR4 (N4783, N4779, N4436, N4443, N2636);
nand NAND2 (N4784, N4768, N413);
and AND3 (N4785, N4769, N1924, N4554);
nor NOR2 (N4786, N4756, N4569);
or OR3 (N4787, N4782, N2565, N4478);
nand NAND2 (N4788, N4774, N4561);
not NOT1 (N4789, N4781);
nor NOR3 (N4790, N4784, N766, N850);
buf BUF1 (N4791, N4778);
not NOT1 (N4792, N4789);
or OR2 (N4793, N4780, N1058);
nand NAND3 (N4794, N4786, N3097, N722);
xor XOR2 (N4795, N4787, N3056);
or OR4 (N4796, N4785, N3243, N726, N54);
not NOT1 (N4797, N4788);
buf BUF1 (N4798, N4794);
not NOT1 (N4799, N4797);
and AND2 (N4800, N4796, N1454);
xor XOR2 (N4801, N4791, N3085);
or OR2 (N4802, N4798, N1223);
nor NOR3 (N4803, N4793, N3028, N3003);
nand NAND3 (N4804, N4801, N3386, N1952);
or OR2 (N4805, N4792, N4031);
and AND2 (N4806, N4800, N138);
nor NOR2 (N4807, N4795, N3369);
or OR3 (N4808, N4803, N3440, N3705);
nor NOR3 (N4809, N4802, N3548, N311);
buf BUF1 (N4810, N4807);
and AND4 (N4811, N4783, N787, N3506, N129);
not NOT1 (N4812, N4790);
not NOT1 (N4813, N4812);
or OR2 (N4814, N4804, N1933);
nor NOR2 (N4815, N4806, N911);
and AND2 (N4816, N4811, N1251);
and AND4 (N4817, N4813, N3178, N3665, N1282);
nand NAND4 (N4818, N4809, N4304, N3178, N412);
buf BUF1 (N4819, N4808);
and AND4 (N4820, N4818, N4815, N3506, N2486);
nor NOR2 (N4821, N4780, N4037);
nor NOR2 (N4822, N4799, N2132);
or OR4 (N4823, N4821, N2800, N3182, N1592);
buf BUF1 (N4824, N4810);
xor XOR2 (N4825, N4823, N1801);
nand NAND3 (N4826, N4824, N1340, N251);
xor XOR2 (N4827, N4819, N3603);
or OR2 (N4828, N4817, N1686);
nand NAND3 (N4829, N4825, N2331, N3617);
or OR3 (N4830, N4829, N1890, N3316);
or OR3 (N4831, N4828, N3367, N4098);
not NOT1 (N4832, N4814);
buf BUF1 (N4833, N4827);
or OR4 (N4834, N4832, N3472, N2754, N2094);
xor XOR2 (N4835, N4822, N1743);
not NOT1 (N4836, N4820);
not NOT1 (N4837, N4816);
and AND2 (N4838, N4805, N2844);
nand NAND4 (N4839, N4830, N2617, N1337, N3089);
buf BUF1 (N4840, N4837);
not NOT1 (N4841, N4838);
and AND3 (N4842, N4836, N3061, N48);
xor XOR2 (N4843, N4839, N4364);
and AND2 (N4844, N4842, N2271);
nor NOR3 (N4845, N4777, N2445, N3869);
xor XOR2 (N4846, N4834, N4165);
or OR3 (N4847, N4840, N427, N4015);
not NOT1 (N4848, N4847);
nor NOR4 (N4849, N4846, N1067, N618, N2769);
xor XOR2 (N4850, N4843, N4312);
nor NOR4 (N4851, N4831, N1833, N2863, N2991);
xor XOR2 (N4852, N4833, N2020);
nor NOR2 (N4853, N4844, N3037);
xor XOR2 (N4854, N4826, N1446);
and AND2 (N4855, N4845, N1336);
nand NAND4 (N4856, N4854, N2772, N176, N1644);
buf BUF1 (N4857, N4835);
xor XOR2 (N4858, N4855, N2205);
nor NOR4 (N4859, N4853, N1336, N1645, N1921);
nand NAND2 (N4860, N4858, N4573);
or OR2 (N4861, N4859, N4567);
nor NOR2 (N4862, N4860, N518);
xor XOR2 (N4863, N4856, N3027);
and AND4 (N4864, N4863, N2384, N1635, N4113);
xor XOR2 (N4865, N4850, N3062);
not NOT1 (N4866, N4849);
or OR2 (N4867, N4861, N4775);
nand NAND2 (N4868, N4857, N1761);
nor NOR4 (N4869, N4867, N2570, N2081, N1902);
not NOT1 (N4870, N4848);
and AND2 (N4871, N4841, N2301);
nand NAND3 (N4872, N4851, N3987, N2830);
or OR2 (N4873, N4865, N4026);
and AND3 (N4874, N4862, N118, N2183);
xor XOR2 (N4875, N4852, N1612);
and AND3 (N4876, N4869, N1244, N2727);
xor XOR2 (N4877, N4873, N1895);
nor NOR4 (N4878, N4871, N2140, N3910, N428);
xor XOR2 (N4879, N4874, N3623);
nand NAND3 (N4880, N4876, N763, N2030);
and AND4 (N4881, N4864, N2521, N2975, N4358);
buf BUF1 (N4882, N4881);
nand NAND4 (N4883, N4870, N3738, N3126, N1737);
xor XOR2 (N4884, N4866, N2860);
buf BUF1 (N4885, N4872);
and AND4 (N4886, N4868, N483, N1471, N2753);
and AND2 (N4887, N4885, N3590);
not NOT1 (N4888, N4879);
buf BUF1 (N4889, N4882);
buf BUF1 (N4890, N4883);
xor XOR2 (N4891, N4877, N2455);
xor XOR2 (N4892, N4887, N2647);
or OR2 (N4893, N4884, N3447);
not NOT1 (N4894, N4892);
or OR3 (N4895, N4891, N3606, N1870);
buf BUF1 (N4896, N4875);
nor NOR2 (N4897, N4888, N4847);
not NOT1 (N4898, N4878);
not NOT1 (N4899, N4898);
and AND2 (N4900, N4897, N2691);
nand NAND3 (N4901, N4894, N3135, N3587);
nand NAND2 (N4902, N4890, N4269);
and AND3 (N4903, N4896, N4142, N1484);
xor XOR2 (N4904, N4903, N513);
xor XOR2 (N4905, N4902, N1430);
not NOT1 (N4906, N4901);
nor NOR4 (N4907, N4893, N1782, N95, N119);
or OR2 (N4908, N4886, N3413);
nand NAND3 (N4909, N4906, N1627, N3935);
or OR2 (N4910, N4904, N4059);
buf BUF1 (N4911, N4899);
nor NOR2 (N4912, N4895, N2477);
nor NOR2 (N4913, N4889, N3117);
nand NAND4 (N4914, N4905, N4160, N3834, N2837);
nand NAND3 (N4915, N4900, N174, N2965);
nand NAND4 (N4916, N4912, N1438, N3135, N831);
and AND4 (N4917, N4913, N1548, N2281, N551);
nand NAND2 (N4918, N4910, N1823);
xor XOR2 (N4919, N4915, N4130);
or OR4 (N4920, N4909, N4672, N3013, N2681);
not NOT1 (N4921, N4916);
xor XOR2 (N4922, N4921, N3785);
and AND3 (N4923, N4911, N1020, N3003);
nor NOR4 (N4924, N4914, N1718, N4425, N4579);
and AND3 (N4925, N4907, N866, N3329);
and AND2 (N4926, N4923, N1200);
or OR3 (N4927, N4925, N109, N4191);
buf BUF1 (N4928, N4922);
nand NAND3 (N4929, N4926, N820, N991);
nand NAND3 (N4930, N4880, N1740, N2353);
or OR2 (N4931, N4929, N982);
nand NAND2 (N4932, N4918, N2327);
nand NAND3 (N4933, N4928, N3614, N3572);
not NOT1 (N4934, N4930);
and AND3 (N4935, N4920, N2011, N34);
nor NOR3 (N4936, N4931, N2556, N4727);
and AND3 (N4937, N4934, N662, N4537);
not NOT1 (N4938, N4932);
xor XOR2 (N4939, N4933, N1707);
nand NAND3 (N4940, N4938, N4322, N1528);
and AND4 (N4941, N4917, N1863, N2802, N4466);
nor NOR2 (N4942, N4936, N4348);
not NOT1 (N4943, N4924);
and AND3 (N4944, N4919, N3906, N2649);
xor XOR2 (N4945, N4935, N3372);
not NOT1 (N4946, N4937);
and AND4 (N4947, N4927, N1255, N171, N4467);
xor XOR2 (N4948, N4908, N904);
or OR2 (N4949, N4943, N639);
buf BUF1 (N4950, N4942);
buf BUF1 (N4951, N4950);
not NOT1 (N4952, N4946);
not NOT1 (N4953, N4944);
and AND3 (N4954, N4945, N94, N1387);
not NOT1 (N4955, N4939);
xor XOR2 (N4956, N4951, N3657);
not NOT1 (N4957, N4956);
nand NAND2 (N4958, N4955, N2247);
nor NOR3 (N4959, N4954, N1077, N637);
or OR3 (N4960, N4940, N437, N609);
buf BUF1 (N4961, N4953);
buf BUF1 (N4962, N4947);
and AND2 (N4963, N4962, N3756);
or OR3 (N4964, N4941, N712, N4432);
not NOT1 (N4965, N4961);
xor XOR2 (N4966, N4963, N3274);
or OR3 (N4967, N4966, N2835, N4360);
xor XOR2 (N4968, N4949, N73);
or OR4 (N4969, N4968, N4602, N3279, N355);
nor NOR3 (N4970, N4952, N445, N3368);
or OR4 (N4971, N4970, N2279, N2867, N1146);
or OR2 (N4972, N4964, N2067);
nor NOR3 (N4973, N4958, N879, N441);
and AND4 (N4974, N4965, N469, N1636, N465);
not NOT1 (N4975, N4959);
nand NAND4 (N4976, N4972, N4028, N4578, N1601);
or OR4 (N4977, N4967, N329, N4901, N2140);
not NOT1 (N4978, N4957);
nand NAND2 (N4979, N4978, N3979);
or OR4 (N4980, N4960, N3508, N717, N1263);
or OR4 (N4981, N4948, N2835, N2601, N2475);
not NOT1 (N4982, N4971);
not NOT1 (N4983, N4982);
not NOT1 (N4984, N4980);
or OR4 (N4985, N4975, N2278, N2529, N81);
nor NOR3 (N4986, N4981, N3213, N601);
xor XOR2 (N4987, N4983, N2527);
not NOT1 (N4988, N4976);
xor XOR2 (N4989, N4987, N3428);
nor NOR4 (N4990, N4985, N4146, N4828, N815);
not NOT1 (N4991, N4979);
nand NAND2 (N4992, N4986, N4654);
or OR3 (N4993, N4974, N962, N1524);
not NOT1 (N4994, N4977);
nor NOR2 (N4995, N4993, N1230);
xor XOR2 (N4996, N4988, N2147);
nor NOR3 (N4997, N4996, N1222, N4425);
and AND2 (N4998, N4995, N407);
nand NAND3 (N4999, N4989, N106, N4450);
buf BUF1 (N5000, N4998);
nor NOR2 (N5001, N4992, N4795);
buf BUF1 (N5002, N4969);
buf BUF1 (N5003, N4997);
nand NAND3 (N5004, N5002, N3819, N2866);
not NOT1 (N5005, N4984);
xor XOR2 (N5006, N5005, N2823);
nor NOR2 (N5007, N5001, N4190);
and AND2 (N5008, N5004, N2185);
nor NOR3 (N5009, N5008, N1049, N4991);
nand NAND4 (N5010, N2110, N497, N1524, N1128);
nand NAND4 (N5011, N4994, N1610, N1598, N4939);
and AND2 (N5012, N5000, N2033);
not NOT1 (N5013, N4999);
nor NOR3 (N5014, N5009, N2879, N2426);
and AND3 (N5015, N5014, N4431, N4293);
or OR2 (N5016, N4990, N2664);
buf BUF1 (N5017, N5012);
or OR2 (N5018, N5016, N779);
buf BUF1 (N5019, N4973);
and AND4 (N5020, N5006, N814, N2781, N1792);
xor XOR2 (N5021, N5015, N3153);
or OR3 (N5022, N5013, N673, N3887);
nand NAND3 (N5023, N5020, N4836, N3981);
xor XOR2 (N5024, N5007, N3939);
xor XOR2 (N5025, N5011, N4572);
not NOT1 (N5026, N5025);
and AND4 (N5027, N5017, N4995, N1294, N4472);
xor XOR2 (N5028, N5019, N2920);
not NOT1 (N5029, N5003);
or OR3 (N5030, N5023, N1474, N3480);
nand NAND3 (N5031, N5028, N3917, N2997);
or OR2 (N5032, N5027, N1832);
not NOT1 (N5033, N5018);
xor XOR2 (N5034, N5022, N3732);
xor XOR2 (N5035, N5021, N3684);
nand NAND4 (N5036, N5033, N1418, N2867, N1766);
not NOT1 (N5037, N5034);
and AND3 (N5038, N5024, N4037, N2029);
or OR2 (N5039, N5031, N523);
xor XOR2 (N5040, N5036, N2487);
nor NOR3 (N5041, N5029, N2730, N3954);
buf BUF1 (N5042, N5039);
xor XOR2 (N5043, N5030, N3498);
buf BUF1 (N5044, N5041);
nand NAND4 (N5045, N5038, N1597, N5021, N3428);
nand NAND3 (N5046, N5035, N4672, N3316);
and AND4 (N5047, N5037, N4048, N2454, N996);
xor XOR2 (N5048, N5040, N4675);
not NOT1 (N5049, N5042);
and AND3 (N5050, N5044, N4937, N2068);
and AND3 (N5051, N5026, N2506, N3899);
nand NAND2 (N5052, N5051, N1827);
buf BUF1 (N5053, N5045);
and AND3 (N5054, N5048, N2926, N2263);
xor XOR2 (N5055, N5032, N4035);
buf BUF1 (N5056, N5043);
xor XOR2 (N5057, N5046, N4633);
nand NAND2 (N5058, N5056, N3275);
nand NAND4 (N5059, N5055, N1631, N3482, N3683);
or OR2 (N5060, N5053, N2171);
and AND2 (N5061, N5047, N4165);
buf BUF1 (N5062, N5050);
nor NOR4 (N5063, N5062, N2225, N4354, N2956);
nand NAND3 (N5064, N5054, N1058, N3085);
not NOT1 (N5065, N5064);
nor NOR4 (N5066, N5058, N3974, N1134, N4217);
nor NOR2 (N5067, N5061, N2727);
buf BUF1 (N5068, N5066);
buf BUF1 (N5069, N5052);
buf BUF1 (N5070, N5060);
not NOT1 (N5071, N5068);
not NOT1 (N5072, N5067);
nor NOR3 (N5073, N5049, N2748, N1277);
or OR2 (N5074, N5071, N2412);
nor NOR3 (N5075, N5070, N4270, N3999);
buf BUF1 (N5076, N5065);
nor NOR2 (N5077, N5063, N2648);
nand NAND3 (N5078, N5073, N1113, N5056);
nand NAND4 (N5079, N5076, N5050, N681, N1709);
nor NOR4 (N5080, N5057, N2748, N4507, N1676);
or OR2 (N5081, N5079, N3642);
and AND4 (N5082, N5077, N1109, N4357, N1363);
not NOT1 (N5083, N5059);
xor XOR2 (N5084, N5069, N197);
xor XOR2 (N5085, N5084, N41);
not NOT1 (N5086, N5082);
not NOT1 (N5087, N5080);
and AND4 (N5088, N5074, N624, N2983, N1874);
buf BUF1 (N5089, N5083);
xor XOR2 (N5090, N5078, N3468);
and AND4 (N5091, N5075, N4686, N1038, N4809);
nor NOR4 (N5092, N5085, N5058, N3994, N3020);
nor NOR4 (N5093, N5010, N2947, N4352, N3432);
and AND4 (N5094, N5088, N103, N2141, N3752);
or OR3 (N5095, N5087, N3777, N1247);
not NOT1 (N5096, N5095);
and AND4 (N5097, N5093, N2694, N3878, N3877);
not NOT1 (N5098, N5097);
buf BUF1 (N5099, N5086);
nor NOR3 (N5100, N5091, N4174, N1513);
nor NOR3 (N5101, N5092, N2836, N3934);
nand NAND3 (N5102, N5096, N1313, N3949);
buf BUF1 (N5103, N5098);
buf BUF1 (N5104, N5100);
or OR2 (N5105, N5099, N1520);
nor NOR3 (N5106, N5105, N2658, N338);
buf BUF1 (N5107, N5081);
nand NAND4 (N5108, N5089, N3937, N3971, N885);
not NOT1 (N5109, N5101);
buf BUF1 (N5110, N5104);
buf BUF1 (N5111, N5110);
nand NAND4 (N5112, N5102, N4680, N2269, N359);
nor NOR3 (N5113, N5109, N767, N4695);
not NOT1 (N5114, N5094);
not NOT1 (N5115, N5112);
nor NOR2 (N5116, N5111, N3117);
and AND3 (N5117, N5106, N712, N811);
nor NOR3 (N5118, N5090, N494, N3392);
xor XOR2 (N5119, N5113, N1699);
not NOT1 (N5120, N5072);
buf BUF1 (N5121, N5108);
or OR3 (N5122, N5107, N3440, N2425);
xor XOR2 (N5123, N5118, N3509);
or OR3 (N5124, N5121, N5084, N842);
buf BUF1 (N5125, N5119);
nand NAND2 (N5126, N5117, N3048);
not NOT1 (N5127, N5115);
nand NAND2 (N5128, N5116, N4878);
buf BUF1 (N5129, N5128);
nand NAND3 (N5130, N5125, N2951, N1463);
nor NOR2 (N5131, N5120, N4045);
buf BUF1 (N5132, N5114);
xor XOR2 (N5133, N5129, N2411);
nand NAND2 (N5134, N5133, N2397);
xor XOR2 (N5135, N5134, N628);
or OR4 (N5136, N5122, N866, N4476, N390);
xor XOR2 (N5137, N5130, N114);
or OR3 (N5138, N5135, N2275, N1859);
or OR4 (N5139, N5137, N808, N80, N199);
nor NOR3 (N5140, N5139, N2509, N4622);
buf BUF1 (N5141, N5140);
nor NOR2 (N5142, N5138, N1785);
not NOT1 (N5143, N5126);
nor NOR3 (N5144, N5124, N4595, N2173);
or OR2 (N5145, N5136, N3914);
nor NOR2 (N5146, N5131, N2526);
buf BUF1 (N5147, N5141);
or OR4 (N5148, N5123, N240, N572, N1770);
nand NAND2 (N5149, N5132, N168);
nand NAND3 (N5150, N5127, N1048, N1441);
buf BUF1 (N5151, N5146);
xor XOR2 (N5152, N5147, N3626);
and AND2 (N5153, N5149, N2949);
and AND3 (N5154, N5145, N738, N3034);
and AND2 (N5155, N5142, N1300);
buf BUF1 (N5156, N5155);
xor XOR2 (N5157, N5151, N2844);
nor NOR3 (N5158, N5152, N3443, N2511);
buf BUF1 (N5159, N5103);
buf BUF1 (N5160, N5159);
or OR2 (N5161, N5156, N2923);
or OR2 (N5162, N5158, N1993);
nor NOR2 (N5163, N5153, N3900);
and AND3 (N5164, N5150, N945, N30);
or OR2 (N5165, N5157, N3526);
not NOT1 (N5166, N5164);
nand NAND2 (N5167, N5154, N1023);
nor NOR4 (N5168, N5144, N150, N416, N2873);
nor NOR4 (N5169, N5160, N135, N4968, N698);
nor NOR3 (N5170, N5161, N1009, N526);
nand NAND3 (N5171, N5163, N1355, N4254);
and AND4 (N5172, N5165, N3667, N2679, N4843);
not NOT1 (N5173, N5171);
nor NOR2 (N5174, N5167, N4160);
and AND4 (N5175, N5173, N2867, N1643, N4569);
nor NOR4 (N5176, N5170, N4193, N2365, N2146);
or OR2 (N5177, N5143, N1348);
xor XOR2 (N5178, N5169, N3277);
not NOT1 (N5179, N5177);
and AND3 (N5180, N5172, N999, N3614);
nand NAND3 (N5181, N5176, N2379, N4125);
nand NAND2 (N5182, N5178, N1421);
nor NOR3 (N5183, N5166, N3524, N556);
not NOT1 (N5184, N5175);
and AND4 (N5185, N5174, N2529, N4964, N474);
or OR3 (N5186, N5148, N591, N2890);
xor XOR2 (N5187, N5186, N4675);
not NOT1 (N5188, N5181);
xor XOR2 (N5189, N5180, N4887);
xor XOR2 (N5190, N5183, N3009);
or OR2 (N5191, N5187, N2563);
and AND4 (N5192, N5182, N607, N1932, N3979);
or OR3 (N5193, N5192, N2526, N3971);
or OR4 (N5194, N5191, N4223, N1600, N2849);
buf BUF1 (N5195, N5168);
and AND4 (N5196, N5190, N3627, N1466, N1843);
nor NOR3 (N5197, N5179, N2499, N3118);
buf BUF1 (N5198, N5193);
not NOT1 (N5199, N5195);
xor XOR2 (N5200, N5199, N169);
and AND3 (N5201, N5198, N2041, N1126);
and AND3 (N5202, N5200, N3659, N1799);
not NOT1 (N5203, N5188);
xor XOR2 (N5204, N5203, N1601);
xor XOR2 (N5205, N5189, N1681);
buf BUF1 (N5206, N5202);
buf BUF1 (N5207, N5184);
xor XOR2 (N5208, N5194, N1935);
and AND4 (N5209, N5197, N3765, N1778, N1976);
buf BUF1 (N5210, N5207);
nor NOR2 (N5211, N5162, N4726);
and AND4 (N5212, N5196, N694, N277, N1608);
or OR2 (N5213, N5209, N3311);
and AND3 (N5214, N5208, N1615, N5015);
not NOT1 (N5215, N5213);
and AND2 (N5216, N5185, N1873);
nor NOR2 (N5217, N5214, N2971);
and AND3 (N5218, N5211, N3175, N1695);
and AND3 (N5219, N5218, N5007, N1398);
nand NAND2 (N5220, N5204, N3137);
not NOT1 (N5221, N5201);
nor NOR2 (N5222, N5221, N4272);
or OR3 (N5223, N5206, N3527, N3315);
buf BUF1 (N5224, N5220);
and AND4 (N5225, N5219, N5207, N134, N2862);
nand NAND3 (N5226, N5216, N4994, N4995);
buf BUF1 (N5227, N5225);
nand NAND4 (N5228, N5223, N4868, N1521, N5040);
nand NAND4 (N5229, N5210, N875, N1703, N669);
and AND4 (N5230, N5212, N354, N5032, N2482);
nor NOR2 (N5231, N5224, N279);
nand NAND3 (N5232, N5229, N3411, N188);
and AND4 (N5233, N5226, N2570, N2985, N328);
not NOT1 (N5234, N5215);
nand NAND2 (N5235, N5222, N3718);
nor NOR2 (N5236, N5217, N3979);
nor NOR2 (N5237, N5228, N4793);
buf BUF1 (N5238, N5205);
and AND2 (N5239, N5233, N4501);
nor NOR4 (N5240, N5235, N847, N3665, N4207);
not NOT1 (N5241, N5232);
nor NOR4 (N5242, N5241, N4800, N3016, N1223);
and AND2 (N5243, N5240, N3123);
or OR4 (N5244, N5237, N2328, N3460, N2159);
nor NOR2 (N5245, N5230, N3270);
not NOT1 (N5246, N5242);
nor NOR2 (N5247, N5245, N2256);
and AND3 (N5248, N5239, N297, N2819);
nor NOR3 (N5249, N5236, N923, N667);
and AND4 (N5250, N5234, N3474, N351, N2563);
xor XOR2 (N5251, N5249, N4934);
nand NAND3 (N5252, N5250, N3905, N3565);
not NOT1 (N5253, N5244);
not NOT1 (N5254, N5231);
or OR2 (N5255, N5247, N2521);
nor NOR4 (N5256, N5254, N452, N1879, N1025);
nor NOR2 (N5257, N5227, N361);
nand NAND4 (N5258, N5246, N3038, N1562, N1230);
buf BUF1 (N5259, N5255);
and AND3 (N5260, N5243, N2145, N1862);
and AND4 (N5261, N5252, N347, N2764, N910);
or OR2 (N5262, N5259, N835);
nor NOR3 (N5263, N5256, N1919, N2131);
xor XOR2 (N5264, N5260, N1822);
buf BUF1 (N5265, N5248);
or OR4 (N5266, N5251, N95, N589, N871);
and AND2 (N5267, N5265, N1179);
xor XOR2 (N5268, N5253, N4551);
buf BUF1 (N5269, N5263);
xor XOR2 (N5270, N5269, N1846);
nand NAND2 (N5271, N5261, N2920);
and AND2 (N5272, N5238, N3205);
xor XOR2 (N5273, N5264, N4745);
not NOT1 (N5274, N5270);
and AND4 (N5275, N5257, N4277, N4118, N2138);
nand NAND2 (N5276, N5274, N3020);
nor NOR2 (N5277, N5272, N1730);
buf BUF1 (N5278, N5275);
not NOT1 (N5279, N5262);
or OR3 (N5280, N5279, N1743, N275);
or OR3 (N5281, N5268, N3901, N614);
buf BUF1 (N5282, N5258);
buf BUF1 (N5283, N5277);
or OR2 (N5284, N5280, N1372);
and AND4 (N5285, N5276, N3662, N489, N370);
buf BUF1 (N5286, N5273);
or OR2 (N5287, N5283, N863);
or OR4 (N5288, N5267, N3179, N622, N1066);
and AND2 (N5289, N5286, N76);
buf BUF1 (N5290, N5287);
or OR3 (N5291, N5278, N10, N218);
nor NOR4 (N5292, N5289, N582, N3551, N2944);
not NOT1 (N5293, N5288);
and AND3 (N5294, N5285, N3274, N4761);
and AND2 (N5295, N5281, N2894);
buf BUF1 (N5296, N5290);
and AND2 (N5297, N5292, N1148);
nand NAND2 (N5298, N5296, N2944);
or OR2 (N5299, N5266, N1416);
xor XOR2 (N5300, N5294, N1709);
and AND3 (N5301, N5295, N3915, N4004);
or OR2 (N5302, N5301, N3851);
or OR4 (N5303, N5298, N4529, N4322, N1623);
buf BUF1 (N5304, N5282);
nand NAND2 (N5305, N5299, N4434);
xor XOR2 (N5306, N5284, N38);
nor NOR2 (N5307, N5300, N1346);
xor XOR2 (N5308, N5297, N331);
nand NAND2 (N5309, N5304, N2496);
buf BUF1 (N5310, N5307);
nand NAND2 (N5311, N5305, N3898);
not NOT1 (N5312, N5302);
and AND2 (N5313, N5311, N498);
nor NOR3 (N5314, N5271, N4318, N5026);
nand NAND4 (N5315, N5309, N3369, N1153, N3382);
nor NOR2 (N5316, N5306, N852);
xor XOR2 (N5317, N5308, N4114);
or OR2 (N5318, N5293, N631);
or OR4 (N5319, N5314, N4128, N3046, N1942);
buf BUF1 (N5320, N5316);
not NOT1 (N5321, N5317);
buf BUF1 (N5322, N5315);
not NOT1 (N5323, N5310);
xor XOR2 (N5324, N5291, N3443);
xor XOR2 (N5325, N5321, N3208);
nor NOR2 (N5326, N5325, N2627);
nand NAND3 (N5327, N5324, N1056, N280);
nor NOR2 (N5328, N5323, N4530);
buf BUF1 (N5329, N5320);
nor NOR2 (N5330, N5322, N3517);
nor NOR4 (N5331, N5327, N3666, N3427, N3978);
not NOT1 (N5332, N5326);
or OR4 (N5333, N5312, N2904, N4029, N4044);
nand NAND3 (N5334, N5329, N3269, N2553);
xor XOR2 (N5335, N5333, N4956);
nand NAND4 (N5336, N5319, N3129, N4539, N5178);
buf BUF1 (N5337, N5313);
not NOT1 (N5338, N5328);
xor XOR2 (N5339, N5331, N4543);
not NOT1 (N5340, N5336);
xor XOR2 (N5341, N5335, N1991);
buf BUF1 (N5342, N5330);
and AND4 (N5343, N5332, N2622, N890, N2985);
buf BUF1 (N5344, N5338);
nand NAND4 (N5345, N5339, N1979, N679, N3791);
buf BUF1 (N5346, N5343);
xor XOR2 (N5347, N5342, N2192);
xor XOR2 (N5348, N5340, N2643);
or OR2 (N5349, N5344, N4778);
buf BUF1 (N5350, N5348);
xor XOR2 (N5351, N5350, N4909);
xor XOR2 (N5352, N5347, N3702);
nand NAND4 (N5353, N5345, N2797, N1645, N310);
and AND2 (N5354, N5341, N3935);
and AND2 (N5355, N5354, N1260);
xor XOR2 (N5356, N5352, N2426);
nor NOR2 (N5357, N5318, N1972);
and AND3 (N5358, N5334, N4541, N2474);
and AND2 (N5359, N5351, N3435);
xor XOR2 (N5360, N5346, N3151);
and AND2 (N5361, N5359, N2961);
not NOT1 (N5362, N5361);
nand NAND3 (N5363, N5355, N3047, N2105);
xor XOR2 (N5364, N5356, N4661);
xor XOR2 (N5365, N5349, N5170);
not NOT1 (N5366, N5337);
nor NOR4 (N5367, N5357, N50, N3650, N337);
nor NOR4 (N5368, N5353, N5060, N2177, N3229);
nand NAND3 (N5369, N5362, N1383, N2695);
not NOT1 (N5370, N5363);
xor XOR2 (N5371, N5366, N3098);
and AND2 (N5372, N5360, N3739);
or OR3 (N5373, N5370, N4156, N1218);
not NOT1 (N5374, N5358);
or OR3 (N5375, N5365, N698, N3878);
not NOT1 (N5376, N5372);
or OR3 (N5377, N5374, N3147, N3907);
nand NAND2 (N5378, N5368, N3334);
or OR3 (N5379, N5377, N4222, N1442);
buf BUF1 (N5380, N5375);
nand NAND4 (N5381, N5379, N3104, N5048, N5204);
not NOT1 (N5382, N5371);
or OR2 (N5383, N5378, N624);
nor NOR2 (N5384, N5373, N1204);
and AND3 (N5385, N5382, N1541, N1455);
and AND3 (N5386, N5369, N514, N5366);
buf BUF1 (N5387, N5381);
not NOT1 (N5388, N5385);
not NOT1 (N5389, N5386);
xor XOR2 (N5390, N5376, N2005);
and AND4 (N5391, N5389, N5165, N3232, N981);
or OR4 (N5392, N5303, N3586, N4541, N462);
xor XOR2 (N5393, N5384, N1528);
not NOT1 (N5394, N5393);
nor NOR3 (N5395, N5367, N1207, N2590);
nand NAND2 (N5396, N5394, N3469);
and AND3 (N5397, N5388, N2601, N342);
xor XOR2 (N5398, N5390, N227);
and AND4 (N5399, N5396, N5312, N4984, N4986);
nor NOR3 (N5400, N5399, N105, N208);
not NOT1 (N5401, N5392);
nand NAND4 (N5402, N5401, N1799, N3662, N656);
nand NAND3 (N5403, N5383, N3311, N4074);
nor NOR4 (N5404, N5395, N1553, N4332, N399);
xor XOR2 (N5405, N5404, N3406);
xor XOR2 (N5406, N5400, N5351);
and AND3 (N5407, N5387, N3087, N4228);
xor XOR2 (N5408, N5391, N4637);
xor XOR2 (N5409, N5402, N4052);
nor NOR4 (N5410, N5397, N164, N2331, N2177);
and AND3 (N5411, N5410, N2783, N1383);
not NOT1 (N5412, N5408);
nand NAND4 (N5413, N5364, N1121, N4819, N132);
nor NOR2 (N5414, N5409, N3060);
xor XOR2 (N5415, N5407, N2124);
xor XOR2 (N5416, N5398, N579);
or OR3 (N5417, N5411, N3326, N2129);
and AND3 (N5418, N5406, N954, N4358);
not NOT1 (N5419, N5415);
or OR4 (N5420, N5405, N4193, N5039, N3809);
or OR3 (N5421, N5413, N3013, N1511);
buf BUF1 (N5422, N5403);
buf BUF1 (N5423, N5416);
nor NOR3 (N5424, N5380, N2061, N4975);
nor NOR2 (N5425, N5420, N4458);
xor XOR2 (N5426, N5421, N1415);
buf BUF1 (N5427, N5423);
or OR2 (N5428, N5412, N4734);
nand NAND2 (N5429, N5428, N1012);
or OR2 (N5430, N5426, N222);
nor NOR4 (N5431, N5424, N5266, N3652, N3449);
nand NAND4 (N5432, N5429, N2537, N1432, N1910);
or OR2 (N5433, N5418, N3440);
nand NAND2 (N5434, N5422, N667);
nand NAND4 (N5435, N5434, N3183, N3300, N3816);
or OR4 (N5436, N5435, N1737, N3069, N2148);
nor NOR4 (N5437, N5433, N1491, N4961, N4478);
buf BUF1 (N5438, N5436);
nor NOR2 (N5439, N5425, N2020);
not NOT1 (N5440, N5419);
buf BUF1 (N5441, N5427);
or OR2 (N5442, N5432, N481);
nor NOR3 (N5443, N5437, N4582, N2646);
or OR2 (N5444, N5442, N795);
or OR4 (N5445, N5417, N2248, N1645, N1285);
xor XOR2 (N5446, N5438, N259);
or OR2 (N5447, N5446, N1157);
buf BUF1 (N5448, N5445);
buf BUF1 (N5449, N5430);
or OR3 (N5450, N5444, N4735, N445);
and AND2 (N5451, N5447, N4714);
xor XOR2 (N5452, N5431, N4737);
not NOT1 (N5453, N5449);
buf BUF1 (N5454, N5448);
and AND2 (N5455, N5443, N2376);
and AND3 (N5456, N5455, N891, N3239);
xor XOR2 (N5457, N5440, N69);
buf BUF1 (N5458, N5441);
or OR2 (N5459, N5458, N4435);
not NOT1 (N5460, N5457);
xor XOR2 (N5461, N5451, N1544);
and AND2 (N5462, N5461, N1856);
nand NAND3 (N5463, N5462, N2542, N2280);
nand NAND3 (N5464, N5463, N1958, N837);
xor XOR2 (N5465, N5464, N3494);
or OR4 (N5466, N5456, N1824, N1534, N4569);
xor XOR2 (N5467, N5452, N4395);
and AND4 (N5468, N5460, N3350, N3447, N2809);
or OR3 (N5469, N5414, N1644, N23);
nand NAND4 (N5470, N5454, N408, N1875, N1893);
xor XOR2 (N5471, N5469, N2395);
and AND2 (N5472, N5471, N1271);
buf BUF1 (N5473, N5467);
and AND2 (N5474, N5472, N4822);
not NOT1 (N5475, N5459);
and AND3 (N5476, N5439, N3121, N958);
xor XOR2 (N5477, N5450, N4254);
not NOT1 (N5478, N5453);
and AND3 (N5479, N5466, N981, N2537);
and AND3 (N5480, N5477, N3736, N4185);
buf BUF1 (N5481, N5479);
nor NOR3 (N5482, N5474, N597, N1792);
nand NAND2 (N5483, N5476, N742);
or OR2 (N5484, N5470, N210);
nand NAND4 (N5485, N5482, N2774, N1327, N4457);
xor XOR2 (N5486, N5478, N4748);
not NOT1 (N5487, N5483);
or OR4 (N5488, N5468, N5394, N3275, N839);
buf BUF1 (N5489, N5465);
and AND4 (N5490, N5473, N876, N4586, N3776);
xor XOR2 (N5491, N5487, N4679);
xor XOR2 (N5492, N5480, N4027);
not NOT1 (N5493, N5488);
not NOT1 (N5494, N5492);
nor NOR3 (N5495, N5490, N5215, N3268);
not NOT1 (N5496, N5481);
buf BUF1 (N5497, N5496);
nor NOR4 (N5498, N5493, N2436, N4995, N2781);
not NOT1 (N5499, N5475);
not NOT1 (N5500, N5494);
or OR2 (N5501, N5491, N3960);
and AND4 (N5502, N5486, N4684, N3749, N1625);
not NOT1 (N5503, N5498);
not NOT1 (N5504, N5485);
and AND3 (N5505, N5484, N5351, N4192);
buf BUF1 (N5506, N5500);
nor NOR4 (N5507, N5501, N4367, N1225, N3383);
and AND2 (N5508, N5489, N1629);
not NOT1 (N5509, N5497);
or OR4 (N5510, N5504, N2512, N4689, N3688);
buf BUF1 (N5511, N5503);
nor NOR3 (N5512, N5502, N2713, N2177);
nand NAND4 (N5513, N5505, N4706, N5261, N3539);
and AND2 (N5514, N5506, N4030);
buf BUF1 (N5515, N5508);
buf BUF1 (N5516, N5510);
or OR2 (N5517, N5509, N1959);
nor NOR3 (N5518, N5514, N1641, N5399);
and AND4 (N5519, N5507, N1760, N274, N5325);
nand NAND3 (N5520, N5513, N1261, N3501);
not NOT1 (N5521, N5519);
xor XOR2 (N5522, N5511, N3527);
xor XOR2 (N5523, N5495, N2576);
nor NOR3 (N5524, N5516, N2204, N377);
nand NAND4 (N5525, N5517, N3860, N689, N770);
and AND4 (N5526, N5518, N4146, N4966, N553);
xor XOR2 (N5527, N5521, N572);
or OR4 (N5528, N5499, N5177, N1415, N5359);
and AND3 (N5529, N5528, N2243, N1239);
xor XOR2 (N5530, N5526, N133);
and AND3 (N5531, N5527, N1274, N5456);
nand NAND2 (N5532, N5515, N2731);
or OR2 (N5533, N5524, N1350);
and AND2 (N5534, N5522, N1079);
buf BUF1 (N5535, N5529);
nand NAND4 (N5536, N5531, N3756, N4563, N324);
or OR3 (N5537, N5520, N2228, N4068);
xor XOR2 (N5538, N5533, N5325);
xor XOR2 (N5539, N5538, N3548);
not NOT1 (N5540, N5525);
or OR4 (N5541, N5512, N3932, N4493, N683);
buf BUF1 (N5542, N5537);
xor XOR2 (N5543, N5539, N4690);
nand NAND2 (N5544, N5543, N3523);
buf BUF1 (N5545, N5532);
not NOT1 (N5546, N5541);
nand NAND4 (N5547, N5523, N527, N2763, N1352);
or OR3 (N5548, N5547, N3953, N3921);
nor NOR2 (N5549, N5544, N5238);
not NOT1 (N5550, N5545);
buf BUF1 (N5551, N5535);
nor NOR3 (N5552, N5551, N5209, N547);
buf BUF1 (N5553, N5542);
and AND3 (N5554, N5546, N3931, N3762);
buf BUF1 (N5555, N5549);
nor NOR2 (N5556, N5554, N2144);
nor NOR3 (N5557, N5556, N470, N3676);
nand NAND2 (N5558, N5540, N196);
not NOT1 (N5559, N5555);
nor NOR3 (N5560, N5536, N2123, N3117);
not NOT1 (N5561, N5530);
not NOT1 (N5562, N5550);
not NOT1 (N5563, N5548);
buf BUF1 (N5564, N5553);
or OR4 (N5565, N5534, N2368, N329, N4321);
or OR2 (N5566, N5562, N2);
and AND4 (N5567, N5566, N954, N4351, N1975);
nand NAND2 (N5568, N5563, N4391);
buf BUF1 (N5569, N5564);
or OR3 (N5570, N5552, N1967, N3674);
xor XOR2 (N5571, N5559, N5401);
or OR3 (N5572, N5561, N296, N1199);
nor NOR2 (N5573, N5567, N5044);
buf BUF1 (N5574, N5569);
nand NAND4 (N5575, N5573, N5404, N3781, N1193);
buf BUF1 (N5576, N5558);
nor NOR2 (N5577, N5560, N3638);
and AND4 (N5578, N5577, N557, N5540, N3712);
nor NOR2 (N5579, N5557, N2550);
xor XOR2 (N5580, N5578, N2095);
and AND2 (N5581, N5568, N5516);
not NOT1 (N5582, N5576);
buf BUF1 (N5583, N5575);
xor XOR2 (N5584, N5571, N343);
not NOT1 (N5585, N5579);
buf BUF1 (N5586, N5582);
and AND4 (N5587, N5586, N3139, N69, N2387);
buf BUF1 (N5588, N5572);
nand NAND3 (N5589, N5580, N3079, N4997);
buf BUF1 (N5590, N5589);
xor XOR2 (N5591, N5574, N4048);
or OR2 (N5592, N5587, N2112);
nor NOR2 (N5593, N5592, N266);
xor XOR2 (N5594, N5583, N3571);
nor NOR4 (N5595, N5593, N1422, N4412, N3157);
and AND2 (N5596, N5570, N5212);
xor XOR2 (N5597, N5584, N4886);
not NOT1 (N5598, N5591);
nand NAND3 (N5599, N5594, N3837, N4566);
not NOT1 (N5600, N5598);
nor NOR3 (N5601, N5585, N4706, N2095);
nor NOR3 (N5602, N5597, N4203, N1734);
buf BUF1 (N5603, N5602);
buf BUF1 (N5604, N5595);
not NOT1 (N5605, N5596);
or OR2 (N5606, N5581, N3167);
xor XOR2 (N5607, N5604, N1224);
nor NOR3 (N5608, N5601, N2979, N5151);
xor XOR2 (N5609, N5565, N4431);
nand NAND3 (N5610, N5590, N103, N5211);
nand NAND3 (N5611, N5608, N3146, N3532);
nor NOR2 (N5612, N5607, N5031);
not NOT1 (N5613, N5600);
or OR3 (N5614, N5611, N691, N1739);
buf BUF1 (N5615, N5610);
not NOT1 (N5616, N5609);
and AND2 (N5617, N5614, N1508);
buf BUF1 (N5618, N5603);
or OR3 (N5619, N5617, N2238, N4615);
xor XOR2 (N5620, N5615, N1409);
xor XOR2 (N5621, N5619, N2160);
xor XOR2 (N5622, N5613, N4930);
nor NOR3 (N5623, N5621, N1395, N4870);
buf BUF1 (N5624, N5599);
and AND3 (N5625, N5612, N3907, N250);
and AND4 (N5626, N5605, N4647, N723, N2214);
buf BUF1 (N5627, N5625);
and AND2 (N5628, N5623, N2271);
nand NAND2 (N5629, N5606, N3962);
nand NAND2 (N5630, N5626, N1875);
xor XOR2 (N5631, N5620, N791);
and AND2 (N5632, N5616, N2878);
or OR2 (N5633, N5627, N3625);
nand NAND2 (N5634, N5628, N3831);
and AND4 (N5635, N5634, N2591, N341, N1543);
and AND4 (N5636, N5630, N3328, N4126, N3211);
xor XOR2 (N5637, N5635, N2847);
xor XOR2 (N5638, N5637, N3838);
nand NAND2 (N5639, N5632, N1640);
and AND3 (N5640, N5631, N3906, N1472);
and AND2 (N5641, N5622, N1193);
and AND2 (N5642, N5636, N5182);
buf BUF1 (N5643, N5629);
or OR2 (N5644, N5638, N2225);
nor NOR4 (N5645, N5624, N5156, N2752, N2033);
not NOT1 (N5646, N5641);
or OR4 (N5647, N5633, N1523, N4743, N965);
or OR3 (N5648, N5644, N573, N3360);
buf BUF1 (N5649, N5643);
buf BUF1 (N5650, N5648);
nand NAND3 (N5651, N5588, N2156, N4564);
xor XOR2 (N5652, N5639, N4923);
not NOT1 (N5653, N5640);
nor NOR4 (N5654, N5650, N5242, N1349, N5069);
buf BUF1 (N5655, N5651);
and AND2 (N5656, N5647, N4770);
or OR2 (N5657, N5656, N4382);
nor NOR3 (N5658, N5653, N5537, N1192);
buf BUF1 (N5659, N5657);
buf BUF1 (N5660, N5655);
nand NAND4 (N5661, N5652, N5258, N4411, N5054);
nor NOR2 (N5662, N5658, N2263);
buf BUF1 (N5663, N5645);
not NOT1 (N5664, N5661);
buf BUF1 (N5665, N5654);
or OR2 (N5666, N5662, N721);
xor XOR2 (N5667, N5642, N4518);
or OR2 (N5668, N5659, N40);
and AND4 (N5669, N5666, N5412, N4870, N3967);
buf BUF1 (N5670, N5646);
nand NAND2 (N5671, N5670, N5151);
or OR2 (N5672, N5618, N5086);
buf BUF1 (N5673, N5663);
nand NAND3 (N5674, N5665, N5204, N4618);
xor XOR2 (N5675, N5660, N2314);
xor XOR2 (N5676, N5671, N1385);
not NOT1 (N5677, N5675);
buf BUF1 (N5678, N5649);
nor NOR4 (N5679, N5677, N1318, N4654, N434);
nand NAND4 (N5680, N5672, N1782, N3094, N3747);
nand NAND3 (N5681, N5676, N3612, N2433);
buf BUF1 (N5682, N5669);
xor XOR2 (N5683, N5680, N5012);
nand NAND2 (N5684, N5682, N116);
nor NOR2 (N5685, N5684, N1688);
xor XOR2 (N5686, N5679, N1661);
buf BUF1 (N5687, N5664);
xor XOR2 (N5688, N5683, N2219);
nand NAND4 (N5689, N5686, N1520, N4343, N4745);
nand NAND4 (N5690, N5687, N4821, N868, N3437);
buf BUF1 (N5691, N5668);
or OR3 (N5692, N5673, N2250, N1445);
xor XOR2 (N5693, N5691, N4285);
buf BUF1 (N5694, N5678);
or OR3 (N5695, N5694, N3042, N1303);
or OR2 (N5696, N5667, N1436);
or OR3 (N5697, N5695, N781, N4308);
not NOT1 (N5698, N5690);
not NOT1 (N5699, N5681);
xor XOR2 (N5700, N5697, N5424);
and AND3 (N5701, N5689, N4139, N5305);
or OR4 (N5702, N5674, N5405, N1132, N4451);
nor NOR2 (N5703, N5699, N1861);
buf BUF1 (N5704, N5700);
or OR3 (N5705, N5685, N3659, N3816);
not NOT1 (N5706, N5696);
and AND4 (N5707, N5701, N1715, N1831, N3213);
not NOT1 (N5708, N5688);
nor NOR2 (N5709, N5705, N4517);
nand NAND2 (N5710, N5702, N4248);
or OR4 (N5711, N5704, N4374, N4257, N2579);
nor NOR4 (N5712, N5707, N2235, N4458, N1517);
nand NAND4 (N5713, N5698, N2799, N4682, N548);
nand NAND4 (N5714, N5709, N5363, N3388, N2391);
or OR2 (N5715, N5692, N879);
and AND4 (N5716, N5714, N1223, N695, N1864);
xor XOR2 (N5717, N5715, N1009);
buf BUF1 (N5718, N5717);
and AND4 (N5719, N5710, N4143, N4518, N2691);
not NOT1 (N5720, N5703);
not NOT1 (N5721, N5712);
buf BUF1 (N5722, N5716);
and AND4 (N5723, N5720, N91, N5104, N1941);
not NOT1 (N5724, N5719);
nand NAND3 (N5725, N5693, N896, N3710);
nor NOR2 (N5726, N5723, N1170);
not NOT1 (N5727, N5724);
nor NOR2 (N5728, N5713, N3037);
or OR4 (N5729, N5725, N2227, N768, N2881);
buf BUF1 (N5730, N5727);
nor NOR2 (N5731, N5726, N3494);
buf BUF1 (N5732, N5711);
nand NAND2 (N5733, N5721, N1850);
nand NAND3 (N5734, N5718, N767, N3767);
and AND2 (N5735, N5733, N5232);
buf BUF1 (N5736, N5735);
and AND4 (N5737, N5708, N5250, N2097, N5387);
nor NOR4 (N5738, N5734, N1175, N4281, N3053);
nor NOR3 (N5739, N5728, N109, N3148);
nand NAND3 (N5740, N5738, N5001, N2667);
not NOT1 (N5741, N5730);
not NOT1 (N5742, N5706);
buf BUF1 (N5743, N5741);
buf BUF1 (N5744, N5732);
and AND2 (N5745, N5731, N1254);
xor XOR2 (N5746, N5739, N2568);
buf BUF1 (N5747, N5742);
nor NOR3 (N5748, N5740, N444, N5390);
buf BUF1 (N5749, N5747);
nand NAND4 (N5750, N5749, N3831, N5390, N3103);
buf BUF1 (N5751, N5745);
and AND4 (N5752, N5744, N2573, N989, N4519);
nor NOR4 (N5753, N5722, N394, N1740, N4663);
xor XOR2 (N5754, N5737, N3021);
or OR4 (N5755, N5748, N537, N5169, N1646);
xor XOR2 (N5756, N5746, N2929);
buf BUF1 (N5757, N5751);
or OR3 (N5758, N5756, N3670, N3336);
and AND4 (N5759, N5752, N3014, N5318, N826);
not NOT1 (N5760, N5736);
xor XOR2 (N5761, N5755, N4246);
and AND2 (N5762, N5757, N2217);
xor XOR2 (N5763, N5762, N540);
nand NAND4 (N5764, N5750, N2697, N962, N2338);
not NOT1 (N5765, N5758);
xor XOR2 (N5766, N5753, N2680);
nor NOR4 (N5767, N5761, N3143, N1844, N250);
xor XOR2 (N5768, N5766, N4412);
or OR3 (N5769, N5760, N4674, N2872);
buf BUF1 (N5770, N5767);
xor XOR2 (N5771, N5759, N3753);
nand NAND3 (N5772, N5765, N5519, N3844);
not NOT1 (N5773, N5754);
nor NOR3 (N5774, N5729, N1026, N4282);
and AND2 (N5775, N5772, N3773);
or OR3 (N5776, N5773, N2664, N2709);
nor NOR3 (N5777, N5764, N2171, N4960);
or OR2 (N5778, N5763, N2474);
buf BUF1 (N5779, N5777);
buf BUF1 (N5780, N5743);
nand NAND4 (N5781, N5776, N4675, N4212, N3223);
xor XOR2 (N5782, N5770, N4058);
nand NAND3 (N5783, N5775, N451, N2640);
not NOT1 (N5784, N5774);
nor NOR2 (N5785, N5769, N1477);
buf BUF1 (N5786, N5771);
nand NAND2 (N5787, N5768, N4200);
not NOT1 (N5788, N5779);
buf BUF1 (N5789, N5788);
nor NOR4 (N5790, N5785, N2459, N4607, N902);
not NOT1 (N5791, N5783);
nand NAND2 (N5792, N5790, N5305);
nand NAND3 (N5793, N5784, N3553, N4186);
nand NAND4 (N5794, N5789, N2896, N367, N2643);
nand NAND2 (N5795, N5781, N4649);
not NOT1 (N5796, N5787);
or OR2 (N5797, N5792, N1928);
xor XOR2 (N5798, N5786, N2839);
and AND3 (N5799, N5796, N5244, N2587);
not NOT1 (N5800, N5797);
buf BUF1 (N5801, N5782);
nor NOR4 (N5802, N5800, N1850, N5127, N2743);
xor XOR2 (N5803, N5801, N765);
and AND3 (N5804, N5791, N1636, N833);
nor NOR4 (N5805, N5802, N1641, N3839, N290);
xor XOR2 (N5806, N5794, N968);
and AND3 (N5807, N5804, N2590, N68);
buf BUF1 (N5808, N5799);
nor NOR2 (N5809, N5798, N98);
nand NAND2 (N5810, N5793, N2700);
and AND2 (N5811, N5778, N3870);
and AND4 (N5812, N5780, N3352, N352, N1883);
or OR3 (N5813, N5811, N3947, N5710);
and AND3 (N5814, N5795, N3745, N1299);
nand NAND2 (N5815, N5809, N844);
xor XOR2 (N5816, N5806, N2977);
or OR3 (N5817, N5813, N3377, N1417);
or OR2 (N5818, N5815, N4519);
not NOT1 (N5819, N5812);
nor NOR2 (N5820, N5819, N2127);
and AND2 (N5821, N5807, N3630);
not NOT1 (N5822, N5817);
nor NOR4 (N5823, N5805, N1844, N3088, N2951);
xor XOR2 (N5824, N5822, N1090);
buf BUF1 (N5825, N5820);
not NOT1 (N5826, N5816);
nor NOR3 (N5827, N5803, N3111, N1848);
nor NOR4 (N5828, N5823, N60, N2262, N3518);
xor XOR2 (N5829, N5824, N748);
nor NOR4 (N5830, N5828, N4250, N4397, N5392);
or OR2 (N5831, N5827, N2616);
or OR2 (N5832, N5814, N2569);
xor XOR2 (N5833, N5832, N720);
nand NAND4 (N5834, N5821, N5695, N2706, N3214);
xor XOR2 (N5835, N5810, N1778);
xor XOR2 (N5836, N5818, N4574);
or OR2 (N5837, N5830, N3609);
not NOT1 (N5838, N5837);
or OR4 (N5839, N5835, N4591, N1423, N1959);
nand NAND3 (N5840, N5838, N1301, N2405);
nor NOR4 (N5841, N5825, N1985, N3312, N3408);
xor XOR2 (N5842, N5840, N4349);
and AND3 (N5843, N5836, N3969, N3934);
nand NAND2 (N5844, N5843, N4195);
and AND3 (N5845, N5842, N5626, N1050);
xor XOR2 (N5846, N5834, N4557);
nor NOR4 (N5847, N5831, N5435, N5091, N365);
and AND2 (N5848, N5844, N154);
not NOT1 (N5849, N5846);
nor NOR4 (N5850, N5826, N2123, N2043, N2866);
not NOT1 (N5851, N5841);
xor XOR2 (N5852, N5850, N2832);
buf BUF1 (N5853, N5849);
or OR2 (N5854, N5851, N2816);
not NOT1 (N5855, N5852);
nand NAND4 (N5856, N5847, N697, N3348, N5651);
and AND2 (N5857, N5854, N6);
nor NOR2 (N5858, N5808, N1766);
xor XOR2 (N5859, N5839, N2306);
and AND2 (N5860, N5853, N2134);
nand NAND4 (N5861, N5833, N3980, N2100, N3340);
nor NOR4 (N5862, N5856, N2427, N1603, N1013);
nand NAND4 (N5863, N5862, N5154, N1474, N2566);
not NOT1 (N5864, N5845);
nor NOR2 (N5865, N5860, N4684);
xor XOR2 (N5866, N5829, N5059);
not NOT1 (N5867, N5864);
nor NOR2 (N5868, N5855, N2220);
or OR2 (N5869, N5868, N4178);
nand NAND4 (N5870, N5865, N2749, N2059, N5119);
xor XOR2 (N5871, N5861, N4605);
xor XOR2 (N5872, N5870, N3044);
buf BUF1 (N5873, N5871);
nand NAND4 (N5874, N5859, N4022, N1876, N3796);
buf BUF1 (N5875, N5857);
or OR4 (N5876, N5866, N468, N5182, N2053);
or OR4 (N5877, N5848, N2842, N4277, N794);
and AND2 (N5878, N5858, N3194);
not NOT1 (N5879, N5876);
and AND3 (N5880, N5873, N3099, N140);
nor NOR3 (N5881, N5875, N1260, N1617);
not NOT1 (N5882, N5863);
nand NAND3 (N5883, N5877, N1558, N2545);
xor XOR2 (N5884, N5881, N392);
and AND4 (N5885, N5874, N1114, N1189, N5811);
or OR3 (N5886, N5884, N3863, N4377);
xor XOR2 (N5887, N5869, N3892);
buf BUF1 (N5888, N5880);
buf BUF1 (N5889, N5885);
and AND2 (N5890, N5887, N4343);
not NOT1 (N5891, N5879);
not NOT1 (N5892, N5882);
or OR2 (N5893, N5890, N2698);
buf BUF1 (N5894, N5893);
or OR2 (N5895, N5878, N5839);
buf BUF1 (N5896, N5895);
and AND3 (N5897, N5883, N1106, N1248);
and AND4 (N5898, N5897, N3963, N3075, N1825);
xor XOR2 (N5899, N5886, N1140);
buf BUF1 (N5900, N5896);
or OR2 (N5901, N5892, N4157);
xor XOR2 (N5902, N5901, N5113);
nor NOR4 (N5903, N5898, N5434, N1795, N143);
buf BUF1 (N5904, N5894);
nand NAND3 (N5905, N5903, N3057, N3034);
buf BUF1 (N5906, N5902);
not NOT1 (N5907, N5906);
or OR4 (N5908, N5904, N4587, N1349, N4666);
nor NOR4 (N5909, N5900, N179, N1089, N301);
nor NOR3 (N5910, N5908, N4898, N3960);
xor XOR2 (N5911, N5872, N1920);
nor NOR2 (N5912, N5911, N5180);
and AND3 (N5913, N5899, N2775, N4137);
xor XOR2 (N5914, N5912, N2255);
nand NAND3 (N5915, N5867, N435, N3748);
or OR2 (N5916, N5914, N2976);
buf BUF1 (N5917, N5916);
nor NOR4 (N5918, N5915, N5286, N4791, N136);
nand NAND3 (N5919, N5917, N5604, N3594);
or OR2 (N5920, N5910, N3104);
xor XOR2 (N5921, N5909, N906);
nor NOR3 (N5922, N5888, N2735, N3807);
and AND4 (N5923, N5889, N5439, N1810, N5470);
nand NAND3 (N5924, N5891, N4424, N559);
nand NAND3 (N5925, N5918, N995, N4459);
xor XOR2 (N5926, N5922, N218);
xor XOR2 (N5927, N5920, N3849);
nor NOR3 (N5928, N5926, N384, N4620);
nand NAND3 (N5929, N5925, N2527, N4352);
not NOT1 (N5930, N5907);
and AND2 (N5931, N5913, N4241);
nor NOR4 (N5932, N5927, N2435, N5098, N888);
or OR4 (N5933, N5923, N2132, N5386, N486);
nor NOR3 (N5934, N5905, N2376, N150);
or OR3 (N5935, N5930, N5844, N5190);
nand NAND2 (N5936, N5919, N5510);
xor XOR2 (N5937, N5928, N2892);
buf BUF1 (N5938, N5937);
and AND2 (N5939, N5921, N1776);
buf BUF1 (N5940, N5938);
not NOT1 (N5941, N5932);
or OR4 (N5942, N5935, N660, N5104, N1340);
xor XOR2 (N5943, N5933, N2449);
or OR3 (N5944, N5931, N1902, N4429);
nand NAND2 (N5945, N5939, N521);
or OR3 (N5946, N5943, N1550, N3029);
or OR3 (N5947, N5946, N3176, N3405);
nor NOR3 (N5948, N5941, N5395, N1853);
buf BUF1 (N5949, N5947);
nand NAND4 (N5950, N5936, N431, N4809, N1181);
nor NOR4 (N5951, N5945, N4641, N2679, N832);
not NOT1 (N5952, N5929);
nand NAND2 (N5953, N5952, N4347);
and AND2 (N5954, N5950, N2197);
buf BUF1 (N5955, N5949);
xor XOR2 (N5956, N5940, N4834);
or OR3 (N5957, N5954, N1974, N267);
and AND2 (N5958, N5957, N1733);
and AND4 (N5959, N5951, N5909, N255, N4758);
buf BUF1 (N5960, N5948);
or OR3 (N5961, N5960, N378, N5145);
not NOT1 (N5962, N5955);
nor NOR4 (N5963, N5942, N1677, N766, N4620);
or OR2 (N5964, N5962, N2574);
xor XOR2 (N5965, N5924, N1842);
buf BUF1 (N5966, N5953);
and AND3 (N5967, N5963, N2091, N2507);
or OR3 (N5968, N5934, N2889, N2115);
buf BUF1 (N5969, N5965);
not NOT1 (N5970, N5961);
and AND2 (N5971, N5966, N5210);
buf BUF1 (N5972, N5969);
not NOT1 (N5973, N5968);
and AND4 (N5974, N5972, N131, N4474, N4444);
nor NOR4 (N5975, N5970, N4664, N4727, N4232);
buf BUF1 (N5976, N5964);
and AND2 (N5977, N5971, N2798);
and AND3 (N5978, N5959, N2310, N2489);
xor XOR2 (N5979, N5977, N3902);
not NOT1 (N5980, N5976);
and AND4 (N5981, N5967, N1297, N4365, N4247);
nand NAND4 (N5982, N5975, N5012, N2812, N2818);
nand NAND4 (N5983, N5978, N470, N2273, N2138);
nor NOR3 (N5984, N5956, N2443, N1642);
and AND3 (N5985, N5983, N3349, N3646);
buf BUF1 (N5986, N5944);
and AND4 (N5987, N5980, N2291, N333, N5804);
not NOT1 (N5988, N5985);
not NOT1 (N5989, N5987);
buf BUF1 (N5990, N5984);
xor XOR2 (N5991, N5989, N3993);
not NOT1 (N5992, N5986);
buf BUF1 (N5993, N5982);
xor XOR2 (N5994, N5958, N3243);
xor XOR2 (N5995, N5993, N2153);
nand NAND3 (N5996, N5973, N777, N4137);
nand NAND3 (N5997, N5994, N997, N2250);
buf BUF1 (N5998, N5974);
and AND3 (N5999, N5990, N2144, N5590);
not NOT1 (N6000, N5998);
or OR3 (N6001, N5988, N5621, N336);
or OR2 (N6002, N6001, N250);
and AND2 (N6003, N5981, N5442);
nand NAND3 (N6004, N5999, N5108, N3623);
not NOT1 (N6005, N5992);
nand NAND3 (N6006, N5991, N4406, N5186);
nand NAND3 (N6007, N5979, N1748, N1695);
nor NOR2 (N6008, N6004, N2721);
not NOT1 (N6009, N6006);
and AND3 (N6010, N6009, N1509, N3482);
buf BUF1 (N6011, N5997);
not NOT1 (N6012, N6005);
not NOT1 (N6013, N6012);
xor XOR2 (N6014, N6011, N5481);
not NOT1 (N6015, N6003);
buf BUF1 (N6016, N6014);
xor XOR2 (N6017, N6002, N525);
buf BUF1 (N6018, N5996);
and AND2 (N6019, N6008, N135);
and AND3 (N6020, N6017, N5611, N1307);
or OR4 (N6021, N6000, N3872, N5801, N2556);
nand NAND4 (N6022, N6013, N5259, N1732, N4349);
nor NOR3 (N6023, N6020, N4682, N910);
not NOT1 (N6024, N6019);
nand NAND4 (N6025, N6010, N5866, N4930, N225);
or OR4 (N6026, N6025, N1723, N5118, N5729);
and AND4 (N6027, N6018, N333, N5376, N2825);
or OR4 (N6028, N6024, N2308, N2411, N3350);
or OR2 (N6029, N6016, N1558);
nor NOR4 (N6030, N6023, N4781, N3324, N3501);
buf BUF1 (N6031, N5995);
or OR3 (N6032, N6026, N5137, N3107);
nor NOR4 (N6033, N6031, N4898, N5442, N5859);
and AND3 (N6034, N6028, N1260, N4860);
xor XOR2 (N6035, N6034, N5329);
xor XOR2 (N6036, N6015, N410);
nand NAND4 (N6037, N6033, N4972, N4371, N4781);
xor XOR2 (N6038, N6030, N465);
nor NOR4 (N6039, N6037, N3178, N2821, N5845);
and AND2 (N6040, N6027, N908);
xor XOR2 (N6041, N6036, N2075);
nor NOR2 (N6042, N6035, N4994);
buf BUF1 (N6043, N6021);
and AND2 (N6044, N6043, N4549);
buf BUF1 (N6045, N6042);
nor NOR4 (N6046, N6039, N223, N1223, N1760);
nor NOR3 (N6047, N6007, N3871, N3055);
xor XOR2 (N6048, N6032, N2735);
not NOT1 (N6049, N6022);
buf BUF1 (N6050, N6040);
nand NAND4 (N6051, N6041, N2863, N2349, N1485);
and AND4 (N6052, N6046, N5413, N5494, N4087);
xor XOR2 (N6053, N6052, N2049);
buf BUF1 (N6054, N6038);
buf BUF1 (N6055, N6049);
nand NAND2 (N6056, N6054, N1797);
xor XOR2 (N6057, N6055, N2269);
or OR4 (N6058, N6047, N4532, N787, N827);
nor NOR4 (N6059, N6057, N3837, N4528, N5770);
nor NOR2 (N6060, N6056, N1033);
and AND2 (N6061, N6058, N286);
buf BUF1 (N6062, N6053);
buf BUF1 (N6063, N6051);
and AND2 (N6064, N6060, N4137);
not NOT1 (N6065, N6044);
xor XOR2 (N6066, N6050, N4910);
nor NOR4 (N6067, N6065, N5845, N3840, N190);
buf BUF1 (N6068, N6045);
and AND3 (N6069, N6064, N544, N6019);
and AND4 (N6070, N6062, N1308, N2655, N5580);
not NOT1 (N6071, N6048);
buf BUF1 (N6072, N6059);
nor NOR3 (N6073, N6066, N18, N3513);
nor NOR4 (N6074, N6067, N2478, N2720, N4689);
and AND3 (N6075, N6061, N3010, N2206);
xor XOR2 (N6076, N6071, N1777);
buf BUF1 (N6077, N6072);
and AND4 (N6078, N6073, N5374, N4159, N1878);
or OR2 (N6079, N6063, N5023);
xor XOR2 (N6080, N6068, N1482);
xor XOR2 (N6081, N6077, N2108);
buf BUF1 (N6082, N6075);
xor XOR2 (N6083, N6079, N1588);
buf BUF1 (N6084, N6029);
not NOT1 (N6085, N6083);
or OR3 (N6086, N6076, N234, N5002);
xor XOR2 (N6087, N6080, N3114);
not NOT1 (N6088, N6070);
not NOT1 (N6089, N6085);
and AND4 (N6090, N6074, N154, N968, N321);
xor XOR2 (N6091, N6090, N2931);
and AND3 (N6092, N6082, N2428, N2265);
buf BUF1 (N6093, N6089);
nor NOR4 (N6094, N6086, N4, N5351, N406);
xor XOR2 (N6095, N6094, N2583);
or OR3 (N6096, N6084, N5990, N1115);
nor NOR3 (N6097, N6096, N1276, N5910);
xor XOR2 (N6098, N6091, N5278);
nand NAND4 (N6099, N6081, N5823, N1557, N5535);
and AND4 (N6100, N6078, N3648, N4845, N4361);
and AND2 (N6101, N6092, N3190);
nor NOR4 (N6102, N6099, N2697, N5909, N2839);
nor NOR3 (N6103, N6095, N4360, N5335);
or OR4 (N6104, N6101, N3091, N1861, N2311);
or OR2 (N6105, N6098, N848);
not NOT1 (N6106, N6105);
nor NOR4 (N6107, N6093, N1319, N6080, N2720);
nand NAND4 (N6108, N6087, N2221, N2931, N5468);
xor XOR2 (N6109, N6107, N5272);
buf BUF1 (N6110, N6106);
or OR3 (N6111, N6104, N3397, N664);
xor XOR2 (N6112, N6102, N4664);
not NOT1 (N6113, N6100);
and AND3 (N6114, N6113, N2212, N4864);
nor NOR2 (N6115, N6108, N4518);
nand NAND2 (N6116, N6103, N3473);
buf BUF1 (N6117, N6109);
nand NAND4 (N6118, N6114, N4887, N4594, N365);
or OR2 (N6119, N6112, N6066);
nor NOR3 (N6120, N6097, N5391, N1426);
buf BUF1 (N6121, N6110);
nand NAND2 (N6122, N6111, N1399);
nor NOR3 (N6123, N6121, N1871, N2517);
and AND2 (N6124, N6118, N1866);
nor NOR4 (N6125, N6069, N1508, N1751, N1991);
nor NOR3 (N6126, N6122, N5484, N265);
nor NOR4 (N6127, N6123, N2455, N598, N3770);
not NOT1 (N6128, N6088);
xor XOR2 (N6129, N6115, N2344);
xor XOR2 (N6130, N6117, N5545);
not NOT1 (N6131, N6124);
xor XOR2 (N6132, N6131, N3325);
xor XOR2 (N6133, N6132, N4696);
nor NOR4 (N6134, N6116, N5101, N5714, N1295);
or OR3 (N6135, N6125, N3972, N264);
or OR4 (N6136, N6130, N696, N1543, N4625);
xor XOR2 (N6137, N6120, N5410);
nand NAND4 (N6138, N6135, N5870, N1548, N4551);
nand NAND4 (N6139, N6138, N2268, N2641, N120);
or OR2 (N6140, N6134, N2262);
nor NOR4 (N6141, N6128, N2720, N5241, N2410);
not NOT1 (N6142, N6129);
and AND4 (N6143, N6141, N1399, N3546, N54);
buf BUF1 (N6144, N6133);
and AND2 (N6145, N6142, N1947);
buf BUF1 (N6146, N6137);
and AND2 (N6147, N6139, N1573);
or OR3 (N6148, N6145, N3454, N1004);
buf BUF1 (N6149, N6127);
nand NAND4 (N6150, N6126, N4663, N4770, N3830);
xor XOR2 (N6151, N6149, N2756);
xor XOR2 (N6152, N6151, N5704);
nor NOR4 (N6153, N6119, N73, N858, N4399);
not NOT1 (N6154, N6152);
xor XOR2 (N6155, N6140, N1983);
nand NAND2 (N6156, N6155, N1887);
nor NOR4 (N6157, N6144, N2620, N2565, N4369);
nor NOR3 (N6158, N6153, N5719, N3164);
and AND2 (N6159, N6156, N1893);
not NOT1 (N6160, N6148);
nor NOR4 (N6161, N6147, N1868, N1293, N348);
nand NAND4 (N6162, N6150, N2063, N5237, N5468);
nand NAND3 (N6163, N6146, N4047, N453);
or OR3 (N6164, N6154, N1073, N2992);
nand NAND4 (N6165, N6143, N2148, N451, N3843);
nand NAND2 (N6166, N6165, N3970);
nor NOR3 (N6167, N6164, N910, N3870);
xor XOR2 (N6168, N6163, N3922);
nor NOR2 (N6169, N6167, N5863);
nand NAND3 (N6170, N6159, N3942, N2985);
buf BUF1 (N6171, N6166);
or OR4 (N6172, N6170, N139, N4498, N688);
nor NOR3 (N6173, N6171, N489, N4123);
nand NAND2 (N6174, N6160, N1026);
xor XOR2 (N6175, N6172, N2700);
nor NOR3 (N6176, N6173, N2696, N866);
not NOT1 (N6177, N6174);
or OR2 (N6178, N6158, N2389);
nor NOR4 (N6179, N6176, N226, N4473, N926);
or OR4 (N6180, N6162, N1349, N2236, N5326);
not NOT1 (N6181, N6178);
not NOT1 (N6182, N6157);
xor XOR2 (N6183, N6179, N1269);
nand NAND3 (N6184, N6183, N288, N508);
buf BUF1 (N6185, N6177);
xor XOR2 (N6186, N6175, N1928);
nand NAND3 (N6187, N6168, N3849, N1545);
nor NOR3 (N6188, N6136, N5584, N3377);
not NOT1 (N6189, N6186);
not NOT1 (N6190, N6169);
and AND4 (N6191, N6187, N1363, N5639, N5335);
or OR3 (N6192, N6181, N2600, N6083);
and AND3 (N6193, N6188, N3096, N3294);
not NOT1 (N6194, N6192);
or OR4 (N6195, N6193, N3330, N3565, N5078);
not NOT1 (N6196, N6190);
nor NOR3 (N6197, N6184, N4785, N5499);
buf BUF1 (N6198, N6196);
xor XOR2 (N6199, N6194, N4686);
xor XOR2 (N6200, N6191, N1115);
buf BUF1 (N6201, N6185);
buf BUF1 (N6202, N6200);
buf BUF1 (N6203, N6180);
nand NAND2 (N6204, N6201, N5451);
buf BUF1 (N6205, N6204);
xor XOR2 (N6206, N6205, N331);
buf BUF1 (N6207, N6203);
nand NAND2 (N6208, N6199, N5846);
or OR2 (N6209, N6206, N5397);
nand NAND2 (N6210, N6182, N3764);
and AND4 (N6211, N6207, N1501, N3965, N102);
or OR4 (N6212, N6211, N4246, N5036, N3673);
or OR3 (N6213, N6198, N5671, N1077);
buf BUF1 (N6214, N6208);
buf BUF1 (N6215, N6213);
and AND4 (N6216, N6209, N2393, N1203, N5184);
and AND4 (N6217, N6212, N6146, N998, N94);
nor NOR4 (N6218, N6195, N2150, N2473, N3877);
or OR3 (N6219, N6216, N6174, N5903);
or OR3 (N6220, N6189, N1866, N4503);
buf BUF1 (N6221, N6219);
and AND2 (N6222, N6220, N2533);
xor XOR2 (N6223, N6215, N888);
or OR3 (N6224, N6214, N6175, N5547);
nand NAND3 (N6225, N6197, N1805, N233);
buf BUF1 (N6226, N6218);
nor NOR3 (N6227, N6161, N4648, N665);
not NOT1 (N6228, N6225);
nand NAND3 (N6229, N6210, N5857, N3178);
or OR4 (N6230, N6222, N4116, N1584, N2503);
and AND4 (N6231, N6227, N2395, N294, N3613);
xor XOR2 (N6232, N6224, N1496);
xor XOR2 (N6233, N6202, N3298);
xor XOR2 (N6234, N6221, N2977);
or OR2 (N6235, N6234, N3052);
buf BUF1 (N6236, N6217);
xor XOR2 (N6237, N6236, N3465);
and AND2 (N6238, N6231, N2819);
nand NAND2 (N6239, N6232, N2904);
xor XOR2 (N6240, N6239, N5747);
and AND4 (N6241, N6223, N1450, N1454, N3719);
buf BUF1 (N6242, N6233);
or OR4 (N6243, N6241, N5162, N4549, N3162);
nor NOR4 (N6244, N6242, N2479, N1787, N539);
buf BUF1 (N6245, N6228);
or OR3 (N6246, N6238, N2582, N3717);
nor NOR2 (N6247, N6230, N5161);
not NOT1 (N6248, N6235);
and AND2 (N6249, N6243, N2817);
xor XOR2 (N6250, N6248, N2181);
not NOT1 (N6251, N6247);
nand NAND3 (N6252, N6237, N1473, N3495);
buf BUF1 (N6253, N6250);
and AND3 (N6254, N6252, N5919, N6173);
buf BUF1 (N6255, N6254);
nand NAND2 (N6256, N6255, N607);
buf BUF1 (N6257, N6240);
nand NAND3 (N6258, N6244, N2766, N3595);
or OR3 (N6259, N6249, N4532, N2010);
buf BUF1 (N6260, N6256);
not NOT1 (N6261, N6226);
and AND4 (N6262, N6246, N5642, N1461, N1027);
nor NOR3 (N6263, N6258, N4255, N4670);
not NOT1 (N6264, N6262);
not NOT1 (N6265, N6261);
nor NOR2 (N6266, N6259, N5787);
nor NOR2 (N6267, N6263, N1126);
nand NAND4 (N6268, N6267, N2452, N940, N3522);
xor XOR2 (N6269, N6268, N5503);
nor NOR3 (N6270, N6253, N3436, N2675);
and AND4 (N6271, N6260, N186, N4658, N3910);
and AND4 (N6272, N6265, N4723, N557, N434);
or OR2 (N6273, N6266, N4991);
not NOT1 (N6274, N6251);
nor NOR3 (N6275, N6274, N3327, N4658);
buf BUF1 (N6276, N6264);
not NOT1 (N6277, N6275);
or OR3 (N6278, N6270, N4452, N1310);
buf BUF1 (N6279, N6276);
not NOT1 (N6280, N6277);
buf BUF1 (N6281, N6280);
xor XOR2 (N6282, N6272, N1180);
nor NOR2 (N6283, N6281, N4515);
or OR2 (N6284, N6282, N6002);
nor NOR3 (N6285, N6245, N686, N59);
or OR4 (N6286, N6279, N2431, N132, N6185);
nand NAND2 (N6287, N6278, N3326);
and AND2 (N6288, N6269, N869);
nor NOR4 (N6289, N6229, N5895, N3565, N4168);
buf BUF1 (N6290, N6289);
nand NAND4 (N6291, N6273, N1911, N564, N2138);
buf BUF1 (N6292, N6271);
nand NAND3 (N6293, N6285, N338, N1342);
buf BUF1 (N6294, N6286);
nand NAND3 (N6295, N6293, N85, N4384);
and AND2 (N6296, N6291, N656);
not NOT1 (N6297, N6292);
and AND2 (N6298, N6284, N6208);
or OR3 (N6299, N6296, N5027, N2656);
or OR3 (N6300, N6297, N533, N2896);
xor XOR2 (N6301, N6290, N4710);
or OR4 (N6302, N6300, N3192, N1710, N3620);
buf BUF1 (N6303, N6295);
xor XOR2 (N6304, N6303, N5968);
xor XOR2 (N6305, N6294, N517);
nand NAND2 (N6306, N6299, N5545);
or OR2 (N6307, N6301, N5355);
nand NAND2 (N6308, N6298, N5683);
and AND4 (N6309, N6307, N2348, N2755, N58);
not NOT1 (N6310, N6306);
not NOT1 (N6311, N6287);
and AND3 (N6312, N6309, N5914, N628);
or OR2 (N6313, N6310, N5394);
nand NAND2 (N6314, N6283, N1552);
nand NAND2 (N6315, N6302, N1298);
nor NOR3 (N6316, N6288, N2406, N5909);
nand NAND3 (N6317, N6315, N3010, N2364);
nand NAND2 (N6318, N6313, N5657);
buf BUF1 (N6319, N6312);
and AND4 (N6320, N6305, N1030, N640, N4209);
nand NAND2 (N6321, N6304, N6202);
buf BUF1 (N6322, N6320);
buf BUF1 (N6323, N6308);
and AND2 (N6324, N6321, N1855);
nand NAND2 (N6325, N6324, N2649);
xor XOR2 (N6326, N6311, N1812);
nand NAND4 (N6327, N6318, N5926, N1190, N5491);
or OR3 (N6328, N6326, N1736, N6091);
or OR2 (N6329, N6316, N4254);
not NOT1 (N6330, N6329);
not NOT1 (N6331, N6330);
and AND4 (N6332, N6314, N2762, N2022, N4243);
nor NOR2 (N6333, N6319, N1908);
not NOT1 (N6334, N6327);
and AND3 (N6335, N6323, N4839, N4734);
nor NOR2 (N6336, N6325, N4678);
or OR4 (N6337, N6317, N3921, N1312, N4005);
or OR4 (N6338, N6337, N4244, N4096, N6261);
and AND4 (N6339, N6257, N919, N5924, N3615);
and AND4 (N6340, N6331, N3349, N4242, N3895);
nor NOR3 (N6341, N6338, N1865, N2433);
not NOT1 (N6342, N6339);
and AND4 (N6343, N6333, N4611, N5692, N3974);
buf BUF1 (N6344, N6340);
or OR3 (N6345, N6342, N1090, N1140);
nor NOR4 (N6346, N6341, N5598, N487, N6298);
xor XOR2 (N6347, N6344, N2331);
and AND4 (N6348, N6332, N1681, N3389, N453);
or OR3 (N6349, N6328, N1780, N5496);
and AND4 (N6350, N6346, N881, N3192, N4853);
or OR4 (N6351, N6343, N4536, N4801, N2535);
nand NAND3 (N6352, N6336, N1921, N3256);
buf BUF1 (N6353, N6348);
and AND3 (N6354, N6322, N4443, N1386);
xor XOR2 (N6355, N6334, N4192);
and AND2 (N6356, N6351, N5872);
or OR4 (N6357, N6345, N2037, N3656, N2140);
not NOT1 (N6358, N6349);
nor NOR4 (N6359, N6357, N6352, N3442, N3500);
buf BUF1 (N6360, N6312);
and AND4 (N6361, N6354, N5916, N2531, N957);
and AND4 (N6362, N6350, N4834, N3388, N4882);
or OR2 (N6363, N6335, N4763);
nor NOR2 (N6364, N6353, N2966);
nor NOR4 (N6365, N6360, N4756, N1136, N180);
not NOT1 (N6366, N6365);
or OR2 (N6367, N6361, N5665);
nor NOR4 (N6368, N6366, N1235, N216, N4274);
buf BUF1 (N6369, N6355);
nor NOR4 (N6370, N6362, N2911, N4536, N355);
or OR3 (N6371, N6369, N4747, N2895);
and AND3 (N6372, N6356, N2433, N658);
buf BUF1 (N6373, N6372);
nand NAND2 (N6374, N6368, N3015);
not NOT1 (N6375, N6364);
xor XOR2 (N6376, N6359, N4005);
nand NAND4 (N6377, N6370, N1269, N2423, N1909);
nor NOR4 (N6378, N6373, N2883, N3778, N380);
or OR3 (N6379, N6358, N2235, N1472);
nor NOR4 (N6380, N6378, N1961, N3420, N146);
or OR3 (N6381, N6347, N4330, N5705);
buf BUF1 (N6382, N6381);
buf BUF1 (N6383, N6382);
xor XOR2 (N6384, N6367, N1121);
and AND2 (N6385, N6384, N1833);
nor NOR4 (N6386, N6363, N4608, N6286, N306);
buf BUF1 (N6387, N6374);
not NOT1 (N6388, N6376);
and AND4 (N6389, N6383, N6265, N915, N3875);
or OR4 (N6390, N6377, N2416, N145, N4942);
xor XOR2 (N6391, N6375, N5896);
not NOT1 (N6392, N6391);
xor XOR2 (N6393, N6389, N6130);
or OR2 (N6394, N6388, N246);
buf BUF1 (N6395, N6393);
buf BUF1 (N6396, N6386);
and AND2 (N6397, N6394, N1058);
nand NAND3 (N6398, N6392, N4302, N182);
not NOT1 (N6399, N6379);
or OR2 (N6400, N6398, N1725);
and AND4 (N6401, N6397, N4882, N4627, N5975);
or OR4 (N6402, N6401, N5430, N4143, N4715);
and AND4 (N6403, N6380, N2640, N694, N3135);
buf BUF1 (N6404, N6403);
or OR4 (N6405, N6395, N2529, N5856, N2663);
not NOT1 (N6406, N6404);
buf BUF1 (N6407, N6405);
or OR4 (N6408, N6385, N1101, N1089, N4597);
buf BUF1 (N6409, N6399);
nor NOR2 (N6410, N6396, N1981);
or OR3 (N6411, N6387, N1449, N1495);
not NOT1 (N6412, N6402);
xor XOR2 (N6413, N6400, N708);
or OR4 (N6414, N6406, N374, N5939, N3080);
nand NAND4 (N6415, N6390, N4998, N4901, N4554);
nand NAND4 (N6416, N6407, N5911, N2229, N6390);
buf BUF1 (N6417, N6411);
or OR4 (N6418, N6416, N3613, N53, N2115);
not NOT1 (N6419, N6415);
nand NAND3 (N6420, N6410, N953, N2005);
nand NAND4 (N6421, N6417, N2417, N2036, N4736);
and AND3 (N6422, N6414, N4784, N4319);
xor XOR2 (N6423, N6420, N1402);
or OR2 (N6424, N6408, N850);
not NOT1 (N6425, N6409);
nand NAND2 (N6426, N6371, N4778);
buf BUF1 (N6427, N6421);
or OR4 (N6428, N6425, N2291, N4883, N3182);
or OR2 (N6429, N6426, N4436);
or OR4 (N6430, N6422, N1382, N3924, N1160);
nand NAND3 (N6431, N6418, N298, N6324);
buf BUF1 (N6432, N6429);
buf BUF1 (N6433, N6430);
nor NOR2 (N6434, N6433, N634);
and AND4 (N6435, N6419, N2818, N3705, N140);
nor NOR3 (N6436, N6413, N4501, N3616);
and AND3 (N6437, N6432, N1409, N3717);
and AND3 (N6438, N6423, N5563, N545);
buf BUF1 (N6439, N6436);
and AND2 (N6440, N6412, N5942);
and AND3 (N6441, N6427, N490, N560);
and AND3 (N6442, N6439, N1216, N1919);
buf BUF1 (N6443, N6424);
nor NOR2 (N6444, N6428, N6354);
and AND4 (N6445, N6435, N1823, N1487, N79);
not NOT1 (N6446, N6442);
buf BUF1 (N6447, N6441);
not NOT1 (N6448, N6445);
nand NAND2 (N6449, N6431, N541);
buf BUF1 (N6450, N6449);
buf BUF1 (N6451, N6434);
nor NOR4 (N6452, N6440, N6375, N5774, N6271);
or OR2 (N6453, N6437, N3712);
nor NOR4 (N6454, N6452, N4254, N374, N1798);
nor NOR2 (N6455, N6447, N4634);
buf BUF1 (N6456, N6450);
or OR2 (N6457, N6448, N5691);
buf BUF1 (N6458, N6451);
not NOT1 (N6459, N6453);
buf BUF1 (N6460, N6443);
xor XOR2 (N6461, N6459, N106);
not NOT1 (N6462, N6458);
xor XOR2 (N6463, N6461, N3829);
not NOT1 (N6464, N6455);
buf BUF1 (N6465, N6454);
not NOT1 (N6466, N6446);
and AND2 (N6467, N6444, N6186);
nor NOR2 (N6468, N6463, N326);
nor NOR3 (N6469, N6457, N4643, N2506);
nor NOR3 (N6470, N6456, N2445, N1902);
not NOT1 (N6471, N6470);
nand NAND4 (N6472, N6466, N4153, N1258, N1752);
nand NAND3 (N6473, N6462, N672, N1738);
xor XOR2 (N6474, N6471, N1777);
not NOT1 (N6475, N6473);
and AND3 (N6476, N6472, N5237, N4086);
and AND4 (N6477, N6474, N4962, N5327, N5883);
and AND3 (N6478, N6476, N2984, N2301);
or OR4 (N6479, N6438, N3279, N672, N1885);
nor NOR3 (N6480, N6460, N2740, N2864);
or OR3 (N6481, N6475, N5560, N958);
nand NAND4 (N6482, N6467, N1185, N4152, N1862);
nor NOR4 (N6483, N6468, N999, N2349, N4945);
buf BUF1 (N6484, N6477);
or OR4 (N6485, N6465, N3623, N660, N1594);
and AND3 (N6486, N6479, N2683, N5457);
and AND3 (N6487, N6469, N3276, N3280);
buf BUF1 (N6488, N6484);
and AND4 (N6489, N6485, N4898, N4072, N1061);
buf BUF1 (N6490, N6488);
buf BUF1 (N6491, N6482);
nor NOR3 (N6492, N6489, N3044, N4796);
buf BUF1 (N6493, N6492);
buf BUF1 (N6494, N6493);
buf BUF1 (N6495, N6480);
and AND4 (N6496, N6487, N1442, N792, N2022);
buf BUF1 (N6497, N6464);
or OR2 (N6498, N6497, N754);
not NOT1 (N6499, N6478);
buf BUF1 (N6500, N6491);
nor NOR2 (N6501, N6496, N5649);
nand NAND2 (N6502, N6499, N3835);
not NOT1 (N6503, N6490);
nand NAND4 (N6504, N6494, N6389, N1623, N5760);
and AND2 (N6505, N6483, N3764);
not NOT1 (N6506, N6505);
nand NAND4 (N6507, N6504, N1036, N644, N824);
and AND3 (N6508, N6502, N5268, N3201);
buf BUF1 (N6509, N6501);
or OR3 (N6510, N6481, N684, N5373);
and AND2 (N6511, N6495, N4098);
nand NAND4 (N6512, N6510, N5135, N120, N2252);
nor NOR3 (N6513, N6500, N4323, N4787);
and AND3 (N6514, N6507, N5870, N1142);
not NOT1 (N6515, N6513);
nor NOR4 (N6516, N6486, N4540, N1681, N6047);
buf BUF1 (N6517, N6515);
or OR4 (N6518, N6511, N5223, N4678, N1747);
not NOT1 (N6519, N6517);
nor NOR4 (N6520, N6498, N3463, N2656, N1494);
buf BUF1 (N6521, N6518);
not NOT1 (N6522, N6521);
xor XOR2 (N6523, N6522, N5587);
not NOT1 (N6524, N6506);
nor NOR4 (N6525, N6520, N1167, N529, N2979);
not NOT1 (N6526, N6524);
nor NOR4 (N6527, N6509, N1534, N4965, N2444);
and AND2 (N6528, N6523, N3301);
or OR4 (N6529, N6528, N2627, N1645, N2068);
buf BUF1 (N6530, N6514);
and AND4 (N6531, N6516, N3427, N6324, N4441);
nand NAND4 (N6532, N6530, N1261, N852, N2956);
buf BUF1 (N6533, N6525);
buf BUF1 (N6534, N6533);
xor XOR2 (N6535, N6512, N5769);
not NOT1 (N6536, N6535);
xor XOR2 (N6537, N6519, N4861);
xor XOR2 (N6538, N6529, N5829);
nand NAND3 (N6539, N6503, N5931, N1598);
not NOT1 (N6540, N6538);
or OR2 (N6541, N6536, N1786);
nor NOR2 (N6542, N6531, N3789);
nor NOR4 (N6543, N6542, N1844, N2640, N6512);
and AND2 (N6544, N6534, N376);
nor NOR2 (N6545, N6537, N1168);
or OR3 (N6546, N6545, N1437, N594);
nor NOR2 (N6547, N6546, N4192);
xor XOR2 (N6548, N6526, N680);
or OR3 (N6549, N6527, N2112, N1740);
not NOT1 (N6550, N6543);
xor XOR2 (N6551, N6540, N557);
not NOT1 (N6552, N6508);
buf BUF1 (N6553, N6552);
xor XOR2 (N6554, N6539, N668);
nand NAND3 (N6555, N6532, N5440, N392);
nor NOR3 (N6556, N6554, N5210, N4815);
nor NOR2 (N6557, N6548, N4450);
nand NAND2 (N6558, N6550, N6305);
xor XOR2 (N6559, N6551, N4714);
xor XOR2 (N6560, N6547, N4477);
buf BUF1 (N6561, N6553);
buf BUF1 (N6562, N6544);
xor XOR2 (N6563, N6562, N6142);
nand NAND2 (N6564, N6559, N1572);
nand NAND3 (N6565, N6555, N2090, N4612);
not NOT1 (N6566, N6556);
xor XOR2 (N6567, N6557, N690);
nor NOR4 (N6568, N6564, N2505, N6541, N6155);
xor XOR2 (N6569, N4749, N258);
not NOT1 (N6570, N6563);
xor XOR2 (N6571, N6567, N501);
nand NAND3 (N6572, N6549, N1614, N5737);
xor XOR2 (N6573, N6568, N6233);
and AND4 (N6574, N6566, N6217, N1114, N6065);
xor XOR2 (N6575, N6569, N4776);
nor NOR4 (N6576, N6571, N4484, N1568, N2115);
buf BUF1 (N6577, N6575);
buf BUF1 (N6578, N6561);
buf BUF1 (N6579, N6573);
buf BUF1 (N6580, N6558);
nand NAND3 (N6581, N6576, N437, N1605);
xor XOR2 (N6582, N6578, N920);
and AND3 (N6583, N6565, N5018, N4654);
buf BUF1 (N6584, N6574);
and AND3 (N6585, N6582, N6521, N658);
and AND4 (N6586, N6579, N2493, N6009, N2755);
xor XOR2 (N6587, N6586, N6136);
and AND3 (N6588, N6572, N4079, N3005);
or OR2 (N6589, N6583, N2007);
not NOT1 (N6590, N6581);
nor NOR2 (N6591, N6590, N6148);
buf BUF1 (N6592, N6589);
buf BUF1 (N6593, N6592);
nand NAND2 (N6594, N6593, N4576);
and AND2 (N6595, N6580, N2859);
and AND4 (N6596, N6560, N4386, N2823, N3974);
nor NOR4 (N6597, N6595, N1991, N1023, N2520);
not NOT1 (N6598, N6577);
nor NOR4 (N6599, N6587, N1891, N378, N853);
nor NOR3 (N6600, N6591, N2313, N3728);
nand NAND3 (N6601, N6598, N2026, N2138);
nor NOR2 (N6602, N6585, N888);
nand NAND2 (N6603, N6600, N2185);
or OR4 (N6604, N6603, N2559, N2707, N5733);
not NOT1 (N6605, N6570);
xor XOR2 (N6606, N6597, N2598);
xor XOR2 (N6607, N6588, N2671);
nor NOR3 (N6608, N6596, N3365, N5419);
and AND3 (N6609, N6604, N4576, N103);
nand NAND2 (N6610, N6609, N146);
or OR4 (N6611, N6608, N1468, N727, N814);
or OR2 (N6612, N6599, N2904);
nor NOR3 (N6613, N6605, N1224, N1246);
nor NOR4 (N6614, N6607, N3409, N4131, N4517);
nor NOR2 (N6615, N6606, N5589);
xor XOR2 (N6616, N6614, N4048);
not NOT1 (N6617, N6610);
xor XOR2 (N6618, N6601, N3154);
not NOT1 (N6619, N6617);
nor NOR3 (N6620, N6616, N3625, N6141);
nor NOR2 (N6621, N6612, N5042);
xor XOR2 (N6622, N6594, N1154);
buf BUF1 (N6623, N6618);
not NOT1 (N6624, N6611);
xor XOR2 (N6625, N6584, N6442);
nand NAND2 (N6626, N6619, N181);
buf BUF1 (N6627, N6620);
and AND2 (N6628, N6621, N1565);
not NOT1 (N6629, N6602);
buf BUF1 (N6630, N6628);
nor NOR4 (N6631, N6630, N3512, N4821, N368);
buf BUF1 (N6632, N6615);
or OR3 (N6633, N6629, N6145, N465);
buf BUF1 (N6634, N6633);
not NOT1 (N6635, N6622);
and AND2 (N6636, N6626, N2949);
nor NOR2 (N6637, N6624, N3555);
nand NAND2 (N6638, N6636, N5479);
and AND4 (N6639, N6634, N1373, N6055, N2763);
or OR3 (N6640, N6638, N3554, N1833);
buf BUF1 (N6641, N6635);
and AND3 (N6642, N6641, N6598, N1574);
buf BUF1 (N6643, N6631);
and AND2 (N6644, N6642, N4185);
or OR4 (N6645, N6644, N1314, N4582, N227);
nand NAND3 (N6646, N6640, N4154, N2870);
nand NAND3 (N6647, N6646, N4457, N2524);
nor NOR2 (N6648, N6627, N6458);
xor XOR2 (N6649, N6637, N6326);
or OR2 (N6650, N6639, N5132);
nand NAND4 (N6651, N6632, N3013, N3126, N4494);
xor XOR2 (N6652, N6625, N1815);
buf BUF1 (N6653, N6647);
xor XOR2 (N6654, N6651, N4029);
and AND2 (N6655, N6654, N355);
and AND2 (N6656, N6648, N3671);
xor XOR2 (N6657, N6650, N4319);
nor NOR4 (N6658, N6645, N5335, N2049, N5290);
nor NOR2 (N6659, N6656, N217);
nand NAND3 (N6660, N6613, N5665, N169);
not NOT1 (N6661, N6623);
or OR4 (N6662, N6653, N6438, N5585, N184);
and AND2 (N6663, N6649, N4490);
or OR3 (N6664, N6657, N4137, N1052);
buf BUF1 (N6665, N6655);
xor XOR2 (N6666, N6658, N3033);
nand NAND3 (N6667, N6643, N1315, N980);
buf BUF1 (N6668, N6666);
and AND3 (N6669, N6661, N5847, N5665);
and AND2 (N6670, N6665, N3502);
not NOT1 (N6671, N6667);
not NOT1 (N6672, N6662);
nor NOR2 (N6673, N6660, N459);
and AND4 (N6674, N6659, N3010, N200, N1873);
nand NAND2 (N6675, N6673, N3985);
nand NAND2 (N6676, N6668, N5665);
buf BUF1 (N6677, N6674);
and AND2 (N6678, N6669, N4667);
xor XOR2 (N6679, N6663, N5075);
and AND3 (N6680, N6664, N6664, N5158);
not NOT1 (N6681, N6680);
or OR2 (N6682, N6679, N281);
xor XOR2 (N6683, N6682, N1162);
nor NOR2 (N6684, N6681, N350);
and AND2 (N6685, N6676, N2111);
buf BUF1 (N6686, N6652);
or OR3 (N6687, N6671, N2724, N3163);
or OR4 (N6688, N6677, N1609, N3808, N672);
nor NOR2 (N6689, N6685, N700);
buf BUF1 (N6690, N6678);
nor NOR2 (N6691, N6689, N5638);
nor NOR3 (N6692, N6687, N4133, N3127);
nand NAND2 (N6693, N6675, N4524);
xor XOR2 (N6694, N6672, N4375);
and AND4 (N6695, N6693, N1423, N3347, N109);
xor XOR2 (N6696, N6670, N4354);
nor NOR2 (N6697, N6686, N4073);
nand NAND4 (N6698, N6691, N2263, N4000, N3856);
or OR3 (N6699, N6692, N694, N4008);
not NOT1 (N6700, N6694);
xor XOR2 (N6701, N6698, N1032);
nor NOR2 (N6702, N6688, N1924);
nor NOR4 (N6703, N6696, N2344, N3694, N2022);
or OR2 (N6704, N6701, N2367);
not NOT1 (N6705, N6703);
nor NOR2 (N6706, N6705, N4504);
or OR4 (N6707, N6702, N5680, N3233, N580);
or OR4 (N6708, N6700, N4167, N6088, N6222);
nand NAND4 (N6709, N6699, N3011, N2577, N86);
buf BUF1 (N6710, N6704);
nand NAND3 (N6711, N6706, N5568, N5617);
or OR2 (N6712, N6711, N2074);
nand NAND2 (N6713, N6709, N6457);
xor XOR2 (N6714, N6684, N3333);
or OR3 (N6715, N6708, N4610, N2172);
buf BUF1 (N6716, N6710);
nor NOR3 (N6717, N6712, N2370, N944);
nand NAND3 (N6718, N6714, N291, N592);
and AND2 (N6719, N6717, N6703);
buf BUF1 (N6720, N6697);
buf BUF1 (N6721, N6695);
xor XOR2 (N6722, N6713, N6486);
nand NAND3 (N6723, N6722, N5604, N4242);
buf BUF1 (N6724, N6723);
and AND4 (N6725, N6716, N6045, N895, N329);
not NOT1 (N6726, N6718);
nand NAND4 (N6727, N6683, N122, N6101, N4446);
nand NAND4 (N6728, N6720, N2387, N2340, N3212);
nand NAND4 (N6729, N6707, N6276, N849, N1397);
buf BUF1 (N6730, N6690);
and AND3 (N6731, N6715, N5807, N2606);
nor NOR2 (N6732, N6721, N1657);
xor XOR2 (N6733, N6726, N1277);
not NOT1 (N6734, N6727);
nand NAND4 (N6735, N6733, N4347, N848, N1428);
nand NAND3 (N6736, N6734, N3230, N127);
nor NOR2 (N6737, N6725, N691);
or OR2 (N6738, N6728, N874);
and AND3 (N6739, N6730, N3948, N3310);
nor NOR4 (N6740, N6737, N4263, N722, N6131);
buf BUF1 (N6741, N6732);
not NOT1 (N6742, N6735);
and AND4 (N6743, N6740, N1784, N5952, N4247);
xor XOR2 (N6744, N6739, N781);
buf BUF1 (N6745, N6729);
nand NAND2 (N6746, N6741, N1442);
and AND3 (N6747, N6738, N6309, N62);
and AND4 (N6748, N6736, N2374, N4841, N5030);
nand NAND2 (N6749, N6742, N3798);
not NOT1 (N6750, N6743);
xor XOR2 (N6751, N6747, N3521);
not NOT1 (N6752, N6751);
not NOT1 (N6753, N6750);
nor NOR3 (N6754, N6749, N2252, N1029);
nand NAND4 (N6755, N6731, N1959, N4989, N4016);
and AND2 (N6756, N6754, N3439);
not NOT1 (N6757, N6745);
nand NAND2 (N6758, N6748, N2710);
and AND4 (N6759, N6757, N726, N3714, N3530);
buf BUF1 (N6760, N6755);
buf BUF1 (N6761, N6756);
nand NAND4 (N6762, N6746, N5530, N1823, N3724);
and AND3 (N6763, N6762, N5482, N667);
xor XOR2 (N6764, N6763, N3691);
not NOT1 (N6765, N6724);
and AND3 (N6766, N6744, N5442, N1737);
or OR3 (N6767, N6766, N3198, N92);
not NOT1 (N6768, N6759);
or OR4 (N6769, N6752, N4833, N2480, N2482);
nor NOR4 (N6770, N6768, N779, N6062, N4552);
and AND2 (N6771, N6769, N1416);
or OR3 (N6772, N6770, N4130, N2361);
or OR2 (N6773, N6758, N4321);
xor XOR2 (N6774, N6753, N1095);
not NOT1 (N6775, N6764);
nor NOR4 (N6776, N6719, N3872, N1886, N6416);
not NOT1 (N6777, N6773);
or OR4 (N6778, N6777, N5896, N3199, N6265);
xor XOR2 (N6779, N6767, N56);
xor XOR2 (N6780, N6776, N573);
not NOT1 (N6781, N6772);
or OR3 (N6782, N6775, N1903, N6489);
or OR3 (N6783, N6760, N2224, N908);
not NOT1 (N6784, N6778);
or OR2 (N6785, N6761, N1577);
or OR2 (N6786, N6774, N1443);
nor NOR2 (N6787, N6783, N5576);
buf BUF1 (N6788, N6771);
not NOT1 (N6789, N6787);
or OR4 (N6790, N6785, N5756, N5054, N4281);
nor NOR2 (N6791, N6788, N2074);
xor XOR2 (N6792, N6786, N4397);
xor XOR2 (N6793, N6784, N3827);
nand NAND3 (N6794, N6790, N536, N4327);
xor XOR2 (N6795, N6782, N1643);
or OR2 (N6796, N6794, N5879);
and AND2 (N6797, N6789, N6175);
and AND3 (N6798, N6781, N1412, N4953);
nand NAND3 (N6799, N6779, N2801, N3302);
nor NOR4 (N6800, N6797, N422, N3595, N5241);
buf BUF1 (N6801, N6796);
and AND4 (N6802, N6793, N398, N6640, N5451);
or OR4 (N6803, N6800, N3335, N4312, N5929);
buf BUF1 (N6804, N6765);
nand NAND3 (N6805, N6804, N4507, N4114);
nand NAND3 (N6806, N6798, N2852, N3434);
buf BUF1 (N6807, N6803);
nand NAND2 (N6808, N6791, N4779);
nand NAND3 (N6809, N6802, N6064, N4521);
and AND2 (N6810, N6805, N1099);
not NOT1 (N6811, N6808);
nand NAND4 (N6812, N6810, N2704, N1897, N1408);
nor NOR2 (N6813, N6809, N824);
and AND4 (N6814, N6795, N6420, N2929, N681);
and AND2 (N6815, N6813, N2412);
and AND2 (N6816, N6792, N4467);
buf BUF1 (N6817, N6816);
nand NAND2 (N6818, N6801, N6291);
buf BUF1 (N6819, N6818);
nor NOR4 (N6820, N6807, N2553, N639, N6746);
nor NOR3 (N6821, N6812, N216, N829);
nand NAND3 (N6822, N6820, N4347, N3439);
not NOT1 (N6823, N6815);
buf BUF1 (N6824, N6806);
or OR3 (N6825, N6814, N6302, N5564);
buf BUF1 (N6826, N6811);
not NOT1 (N6827, N6817);
nand NAND3 (N6828, N6826, N1852, N3591);
xor XOR2 (N6829, N6827, N4864);
or OR3 (N6830, N6828, N2678, N307);
or OR2 (N6831, N6823, N3859);
and AND3 (N6832, N6819, N6120, N2863);
nor NOR4 (N6833, N6780, N364, N518, N3805);
not NOT1 (N6834, N6832);
xor XOR2 (N6835, N6821, N148);
xor XOR2 (N6836, N6831, N133);
nand NAND2 (N6837, N6836, N5359);
not NOT1 (N6838, N6825);
and AND4 (N6839, N6834, N5912, N5921, N3144);
xor XOR2 (N6840, N6799, N4028);
and AND4 (N6841, N6837, N1931, N3336, N5268);
xor XOR2 (N6842, N6833, N6349);
xor XOR2 (N6843, N6822, N6052);
buf BUF1 (N6844, N6838);
nand NAND2 (N6845, N6842, N3679);
xor XOR2 (N6846, N6835, N4458);
buf BUF1 (N6847, N6829);
and AND2 (N6848, N6843, N6005);
not NOT1 (N6849, N6839);
not NOT1 (N6850, N6841);
and AND4 (N6851, N6824, N2715, N3936, N4414);
nor NOR2 (N6852, N6830, N118);
or OR2 (N6853, N6852, N3412);
nor NOR4 (N6854, N6845, N75, N1866, N3225);
not NOT1 (N6855, N6848);
and AND4 (N6856, N6853, N2859, N887, N3052);
nor NOR2 (N6857, N6851, N1778);
and AND4 (N6858, N6854, N372, N4975, N5378);
nor NOR4 (N6859, N6847, N2653, N4948, N2706);
or OR4 (N6860, N6858, N3566, N6719, N3205);
nand NAND2 (N6861, N6855, N5102);
and AND3 (N6862, N6850, N4817, N1486);
and AND3 (N6863, N6860, N3006, N4043);
and AND2 (N6864, N6859, N5719);
not NOT1 (N6865, N6864);
not NOT1 (N6866, N6846);
nor NOR4 (N6867, N6844, N3072, N1330, N5234);
xor XOR2 (N6868, N6840, N1022);
xor XOR2 (N6869, N6865, N5425);
xor XOR2 (N6870, N6849, N6136);
and AND4 (N6871, N6856, N5382, N674, N416);
nand NAND2 (N6872, N6868, N6137);
buf BUF1 (N6873, N6869);
buf BUF1 (N6874, N6863);
xor XOR2 (N6875, N6866, N843);
not NOT1 (N6876, N6872);
xor XOR2 (N6877, N6870, N3016);
or OR4 (N6878, N6867, N1436, N5274, N6382);
or OR4 (N6879, N6873, N3832, N6124, N276);
buf BUF1 (N6880, N6862);
xor XOR2 (N6881, N6879, N3131);
or OR3 (N6882, N6881, N953, N1173);
and AND2 (N6883, N6880, N6407);
nand NAND3 (N6884, N6861, N5249, N2099);
xor XOR2 (N6885, N6877, N2998);
not NOT1 (N6886, N6878);
nor NOR2 (N6887, N6886, N5535);
not NOT1 (N6888, N6882);
or OR2 (N6889, N6871, N1207);
or OR2 (N6890, N6887, N5016);
or OR4 (N6891, N6874, N6220, N2828, N477);
or OR2 (N6892, N6876, N1621);
nor NOR4 (N6893, N6884, N2644, N125, N3900);
xor XOR2 (N6894, N6891, N2970);
nand NAND4 (N6895, N6885, N6451, N810, N162);
and AND3 (N6896, N6895, N217, N3768);
buf BUF1 (N6897, N6857);
not NOT1 (N6898, N6888);
nor NOR4 (N6899, N6898, N5134, N2583, N4356);
not NOT1 (N6900, N6897);
not NOT1 (N6901, N6896);
nor NOR3 (N6902, N6900, N5058, N6149);
buf BUF1 (N6903, N6875);
buf BUF1 (N6904, N6901);
buf BUF1 (N6905, N6902);
not NOT1 (N6906, N6903);
and AND4 (N6907, N6894, N6385, N6276, N398);
buf BUF1 (N6908, N6906);
or OR3 (N6909, N6889, N5981, N3789);
buf BUF1 (N6910, N6905);
or OR3 (N6911, N6908, N6331, N5498);
xor XOR2 (N6912, N6911, N2525);
and AND3 (N6913, N6892, N5503, N5007);
and AND2 (N6914, N6907, N6046);
buf BUF1 (N6915, N6910);
not NOT1 (N6916, N6912);
or OR2 (N6917, N6890, N48);
nand NAND4 (N6918, N6914, N4458, N1579, N5856);
not NOT1 (N6919, N6883);
and AND2 (N6920, N6913, N3545);
not NOT1 (N6921, N6920);
and AND2 (N6922, N6915, N5248);
not NOT1 (N6923, N6921);
and AND4 (N6924, N6899, N2224, N4501, N856);
xor XOR2 (N6925, N6924, N5364);
buf BUF1 (N6926, N6909);
xor XOR2 (N6927, N6925, N4930);
and AND2 (N6928, N6917, N3924);
buf BUF1 (N6929, N6919);
and AND3 (N6930, N6918, N4562, N3382);
and AND2 (N6931, N6893, N5554);
or OR3 (N6932, N6930, N2284, N3251);
not NOT1 (N6933, N6904);
or OR4 (N6934, N6916, N2128, N1305, N712);
nand NAND4 (N6935, N6928, N2818, N6298, N6710);
buf BUF1 (N6936, N6922);
and AND2 (N6937, N6932, N899);
buf BUF1 (N6938, N6933);
nand NAND4 (N6939, N6926, N3385, N5772, N4587);
buf BUF1 (N6940, N6927);
xor XOR2 (N6941, N6938, N5569);
nand NAND3 (N6942, N6935, N3455, N5066);
nor NOR4 (N6943, N6929, N6826, N3858, N5489);
not NOT1 (N6944, N6939);
or OR3 (N6945, N6936, N4669, N5100);
not NOT1 (N6946, N6941);
not NOT1 (N6947, N6945);
not NOT1 (N6948, N6943);
nand NAND4 (N6949, N6931, N703, N4308, N2495);
nor NOR2 (N6950, N6947, N2764);
not NOT1 (N6951, N6934);
not NOT1 (N6952, N6937);
and AND2 (N6953, N6923, N2418);
nor NOR3 (N6954, N6940, N5585, N2730);
and AND3 (N6955, N6954, N6743, N1164);
not NOT1 (N6956, N6942);
nand NAND3 (N6957, N6953, N6184, N5480);
or OR3 (N6958, N6946, N4804, N5191);
not NOT1 (N6959, N6951);
not NOT1 (N6960, N6958);
nand NAND4 (N6961, N6944, N5431, N1822, N455);
xor XOR2 (N6962, N6959, N2713);
or OR3 (N6963, N6957, N6073, N462);
buf BUF1 (N6964, N6952);
or OR4 (N6965, N6962, N1785, N671, N2828);
nor NOR3 (N6966, N6956, N2446, N4690);
xor XOR2 (N6967, N6961, N4139);
or OR3 (N6968, N6960, N3256, N2251);
or OR3 (N6969, N6963, N6299, N5341);
buf BUF1 (N6970, N6967);
and AND4 (N6971, N6966, N3011, N1938, N6455);
nand NAND4 (N6972, N6971, N2413, N54, N1191);
xor XOR2 (N6973, N6972, N5547);
not NOT1 (N6974, N6950);
nor NOR3 (N6975, N6949, N3406, N5565);
nor NOR3 (N6976, N6969, N3409, N648);
and AND3 (N6977, N6973, N3206, N1811);
nand NAND4 (N6978, N6965, N5883, N1971, N4362);
xor XOR2 (N6979, N6975, N565);
or OR2 (N6980, N6968, N2790);
or OR3 (N6981, N6955, N6635, N2841);
nor NOR2 (N6982, N6964, N5256);
and AND2 (N6983, N6982, N1472);
not NOT1 (N6984, N6977);
xor XOR2 (N6985, N6970, N6107);
or OR3 (N6986, N6979, N252, N414);
and AND3 (N6987, N6980, N357, N755);
and AND3 (N6988, N6984, N1227, N6625);
and AND3 (N6989, N6986, N3078, N2042);
and AND3 (N6990, N6987, N2320, N2364);
buf BUF1 (N6991, N6974);
or OR4 (N6992, N6988, N2096, N3065, N4264);
nor NOR3 (N6993, N6978, N4885, N6722);
and AND3 (N6994, N6985, N5512, N6648);
buf BUF1 (N6995, N6948);
xor XOR2 (N6996, N6995, N6058);
buf BUF1 (N6997, N6981);
not NOT1 (N6998, N6997);
buf BUF1 (N6999, N6976);
or OR3 (N7000, N6996, N1894, N867);
and AND2 (N7001, N7000, N3564);
or OR2 (N7002, N6990, N4550);
buf BUF1 (N7003, N6989);
not NOT1 (N7004, N6991);
nor NOR2 (N7005, N6999, N2854);
nand NAND2 (N7006, N6998, N5177);
buf BUF1 (N7007, N6994);
nor NOR4 (N7008, N7001, N2523, N2874, N1496);
buf BUF1 (N7009, N7002);
xor XOR2 (N7010, N7008, N3116);
buf BUF1 (N7011, N7004);
nor NOR3 (N7012, N6993, N860, N536);
nor NOR2 (N7013, N6992, N5297);
xor XOR2 (N7014, N6983, N227);
nor NOR2 (N7015, N7003, N5748);
nand NAND3 (N7016, N7015, N6444, N197);
or OR3 (N7017, N7006, N2110, N4294);
and AND3 (N7018, N7010, N1375, N785);
and AND4 (N7019, N7012, N241, N5840, N1993);
or OR4 (N7020, N7009, N3778, N4852, N6874);
nand NAND3 (N7021, N7011, N6766, N2817);
xor XOR2 (N7022, N7005, N238);
or OR2 (N7023, N7022, N2798);
nand NAND4 (N7024, N7016, N3196, N705, N6853);
xor XOR2 (N7025, N7023, N1997);
nor NOR4 (N7026, N7014, N404, N3515, N3477);
nand NAND2 (N7027, N7019, N3094);
or OR4 (N7028, N7021, N3245, N5843, N5611);
xor XOR2 (N7029, N7026, N3531);
or OR3 (N7030, N7028, N397, N2282);
nor NOR2 (N7031, N7030, N4791);
buf BUF1 (N7032, N7024);
not NOT1 (N7033, N7018);
nand NAND4 (N7034, N7020, N5009, N4996, N5021);
xor XOR2 (N7035, N7027, N2141);
and AND2 (N7036, N7017, N2521);
or OR2 (N7037, N7025, N4963);
nand NAND2 (N7038, N7035, N6793);
or OR3 (N7039, N7007, N3290, N5918);
and AND3 (N7040, N7031, N597, N4049);
or OR4 (N7041, N7013, N6326, N4568, N2517);
nand NAND2 (N7042, N7037, N2416);
nand NAND3 (N7043, N7042, N490, N4457);
nand NAND4 (N7044, N7033, N3573, N2659, N4047);
not NOT1 (N7045, N7032);
not NOT1 (N7046, N7038);
or OR2 (N7047, N7036, N1153);
xor XOR2 (N7048, N7034, N4766);
not NOT1 (N7049, N7047);
nand NAND2 (N7050, N7043, N2136);
xor XOR2 (N7051, N7039, N3946);
or OR2 (N7052, N7049, N484);
nor NOR4 (N7053, N7040, N6101, N2519, N685);
or OR3 (N7054, N7052, N4383, N3333);
xor XOR2 (N7055, N7044, N1170);
not NOT1 (N7056, N7054);
not NOT1 (N7057, N7046);
nor NOR4 (N7058, N7041, N2811, N2271, N3172);
and AND4 (N7059, N7048, N6154, N3817, N340);
nor NOR2 (N7060, N7055, N3566);
not NOT1 (N7061, N7029);
nor NOR4 (N7062, N7059, N2993, N3536, N987);
and AND2 (N7063, N7061, N1489);
buf BUF1 (N7064, N7063);
not NOT1 (N7065, N7060);
xor XOR2 (N7066, N7062, N2726);
and AND4 (N7067, N7056, N1925, N6967, N3718);
nor NOR3 (N7068, N7053, N2306, N3244);
buf BUF1 (N7069, N7050);
and AND3 (N7070, N7067, N1683, N5221);
nor NOR4 (N7071, N7051, N3706, N6411, N2320);
and AND4 (N7072, N7066, N206, N2164, N3283);
or OR4 (N7073, N7064, N2725, N4484, N6659);
nand NAND2 (N7074, N7068, N5342);
xor XOR2 (N7075, N7072, N6433);
xor XOR2 (N7076, N7065, N936);
and AND3 (N7077, N7075, N33, N5529);
or OR3 (N7078, N7073, N298, N438);
nor NOR3 (N7079, N7070, N5449, N3155);
xor XOR2 (N7080, N7074, N2532);
and AND3 (N7081, N7069, N4902, N3714);
buf BUF1 (N7082, N7081);
nand NAND2 (N7083, N7080, N685);
nor NOR4 (N7084, N7082, N729, N2552, N4469);
and AND2 (N7085, N7057, N4023);
xor XOR2 (N7086, N7083, N5973);
nand NAND3 (N7087, N7079, N3118, N6369);
not NOT1 (N7088, N7087);
not NOT1 (N7089, N7078);
or OR3 (N7090, N7077, N4094, N2746);
buf BUF1 (N7091, N7071);
xor XOR2 (N7092, N7085, N698);
buf BUF1 (N7093, N7090);
and AND4 (N7094, N7076, N5213, N1703, N6432);
nor NOR4 (N7095, N7058, N4376, N5252, N6052);
nor NOR4 (N7096, N7084, N355, N915, N6278);
buf BUF1 (N7097, N7091);
not NOT1 (N7098, N7095);
nand NAND2 (N7099, N7089, N750);
buf BUF1 (N7100, N7099);
nor NOR2 (N7101, N7088, N4815);
xor XOR2 (N7102, N7093, N1785);
not NOT1 (N7103, N7102);
buf BUF1 (N7104, N7086);
nand NAND4 (N7105, N7097, N577, N3267, N3809);
nor NOR2 (N7106, N7045, N4717);
not NOT1 (N7107, N7101);
nand NAND4 (N7108, N7103, N2257, N1032, N3602);
nor NOR3 (N7109, N7092, N639, N6077);
nor NOR2 (N7110, N7108, N3640);
nand NAND2 (N7111, N7098, N6876);
nand NAND2 (N7112, N7109, N4364);
or OR4 (N7113, N7106, N3628, N787, N6933);
nor NOR2 (N7114, N7113, N450);
buf BUF1 (N7115, N7104);
xor XOR2 (N7116, N7100, N156);
not NOT1 (N7117, N7107);
xor XOR2 (N7118, N7110, N6407);
buf BUF1 (N7119, N7116);
nor NOR3 (N7120, N7118, N631, N5529);
not NOT1 (N7121, N7094);
xor XOR2 (N7122, N7114, N6092);
buf BUF1 (N7123, N7105);
nand NAND2 (N7124, N7115, N2140);
nand NAND3 (N7125, N7120, N157, N1244);
nor NOR4 (N7126, N7122, N609, N2405, N2577);
and AND3 (N7127, N7096, N6713, N4852);
buf BUF1 (N7128, N7124);
xor XOR2 (N7129, N7123, N4084);
not NOT1 (N7130, N7125);
xor XOR2 (N7131, N7119, N6222);
and AND2 (N7132, N7111, N83);
nor NOR4 (N7133, N7129, N5095, N6257, N5508);
and AND2 (N7134, N7117, N305);
not NOT1 (N7135, N7121);
nand NAND4 (N7136, N7126, N1726, N679, N1129);
buf BUF1 (N7137, N7131);
buf BUF1 (N7138, N7130);
nand NAND4 (N7139, N7127, N6815, N4379, N5699);
nor NOR3 (N7140, N7139, N5209, N4687);
nor NOR3 (N7141, N7138, N341, N3146);
nand NAND4 (N7142, N7137, N628, N4536, N3315);
nor NOR3 (N7143, N7134, N6286, N2286);
not NOT1 (N7144, N7132);
nand NAND2 (N7145, N7112, N2224);
nor NOR4 (N7146, N7135, N2818, N5687, N5060);
xor XOR2 (N7147, N7128, N4039);
xor XOR2 (N7148, N7143, N2167);
nor NOR3 (N7149, N7142, N5163, N6135);
nor NOR3 (N7150, N7133, N4740, N5469);
nor NOR3 (N7151, N7147, N2147, N2046);
or OR4 (N7152, N7148, N6376, N5467, N1406);
xor XOR2 (N7153, N7150, N6046);
buf BUF1 (N7154, N7146);
xor XOR2 (N7155, N7151, N6005);
or OR2 (N7156, N7141, N5728);
nand NAND4 (N7157, N7155, N3116, N1963, N5902);
nor NOR3 (N7158, N7156, N3299, N5615);
and AND4 (N7159, N7157, N3295, N3846, N2986);
and AND4 (N7160, N7145, N3813, N3957, N1096);
not NOT1 (N7161, N7144);
not NOT1 (N7162, N7159);
nor NOR4 (N7163, N7161, N6588, N966, N5686);
nand NAND4 (N7164, N7163, N7030, N5103, N4477);
nor NOR2 (N7165, N7158, N186);
or OR2 (N7166, N7162, N2614);
not NOT1 (N7167, N7154);
not NOT1 (N7168, N7149);
and AND2 (N7169, N7164, N72);
xor XOR2 (N7170, N7160, N2017);
xor XOR2 (N7171, N7153, N1094);
not NOT1 (N7172, N7136);
nand NAND4 (N7173, N7170, N3192, N4433, N4637);
and AND3 (N7174, N7171, N2243, N4202);
xor XOR2 (N7175, N7172, N677);
and AND2 (N7176, N7167, N2246);
nor NOR3 (N7177, N7152, N59, N1522);
nor NOR3 (N7178, N7165, N3703, N2291);
nand NAND3 (N7179, N7166, N169, N5055);
xor XOR2 (N7180, N7168, N5267);
xor XOR2 (N7181, N7173, N789);
nor NOR2 (N7182, N7177, N341);
xor XOR2 (N7183, N7176, N11);
nand NAND2 (N7184, N7181, N4213);
and AND3 (N7185, N7175, N1885, N2398);
nor NOR3 (N7186, N7169, N7028, N404);
nand NAND2 (N7187, N7174, N2074);
xor XOR2 (N7188, N7178, N1158);
xor XOR2 (N7189, N7183, N5513);
nand NAND4 (N7190, N7140, N6995, N3684, N124);
nor NOR2 (N7191, N7182, N6851);
or OR2 (N7192, N7180, N5578);
xor XOR2 (N7193, N7186, N2996);
nor NOR3 (N7194, N7192, N364, N6874);
xor XOR2 (N7195, N7179, N190);
xor XOR2 (N7196, N7185, N3280);
nand NAND4 (N7197, N7188, N6205, N4045, N2425);
nand NAND3 (N7198, N7193, N152, N2066);
nand NAND3 (N7199, N7198, N2561, N6705);
nor NOR3 (N7200, N7194, N4982, N6695);
buf BUF1 (N7201, N7184);
xor XOR2 (N7202, N7196, N4840);
not NOT1 (N7203, N7191);
or OR3 (N7204, N7200, N905, N6641);
nand NAND3 (N7205, N7201, N6041, N6686);
and AND4 (N7206, N7189, N773, N1099, N5183);
nand NAND4 (N7207, N7199, N1994, N4357, N1212);
nand NAND2 (N7208, N7197, N4387);
and AND4 (N7209, N7190, N3428, N2357, N5498);
nand NAND3 (N7210, N7205, N2604, N5162);
nand NAND2 (N7211, N7208, N1448);
buf BUF1 (N7212, N7202);
nor NOR3 (N7213, N7207, N1500, N5870);
xor XOR2 (N7214, N7195, N263);
not NOT1 (N7215, N7187);
xor XOR2 (N7216, N7204, N778);
not NOT1 (N7217, N7203);
buf BUF1 (N7218, N7217);
nand NAND2 (N7219, N7214, N3200);
and AND4 (N7220, N7210, N7161, N2904, N2991);
nand NAND3 (N7221, N7209, N6763, N3833);
not NOT1 (N7222, N7206);
xor XOR2 (N7223, N7212, N3956);
buf BUF1 (N7224, N7220);
buf BUF1 (N7225, N7221);
not NOT1 (N7226, N7224);
or OR3 (N7227, N7223, N6282, N425);
xor XOR2 (N7228, N7213, N3208);
or OR3 (N7229, N7218, N7, N1100);
nor NOR2 (N7230, N7227, N236);
nor NOR4 (N7231, N7226, N5019, N1669, N4295);
xor XOR2 (N7232, N7222, N4847);
xor XOR2 (N7233, N7230, N2276);
buf BUF1 (N7234, N7233);
buf BUF1 (N7235, N7215);
xor XOR2 (N7236, N7228, N3574);
xor XOR2 (N7237, N7236, N1369);
not NOT1 (N7238, N7231);
buf BUF1 (N7239, N7211);
not NOT1 (N7240, N7219);
or OR3 (N7241, N7239, N825, N7085);
nand NAND2 (N7242, N7234, N6972);
or OR3 (N7243, N7235, N2490, N5317);
buf BUF1 (N7244, N7242);
and AND4 (N7245, N7241, N5489, N6330, N6398);
not NOT1 (N7246, N7243);
not NOT1 (N7247, N7244);
xor XOR2 (N7248, N7246, N3844);
not NOT1 (N7249, N7238);
or OR4 (N7250, N7248, N4372, N3600, N2304);
or OR2 (N7251, N7247, N168);
nand NAND3 (N7252, N7237, N171, N2672);
nor NOR3 (N7253, N7216, N4251, N3101);
or OR4 (N7254, N7253, N1956, N4691, N4382);
not NOT1 (N7255, N7254);
not NOT1 (N7256, N7232);
and AND4 (N7257, N7249, N5842, N1299, N2031);
or OR4 (N7258, N7255, N1267, N1380, N6427);
and AND4 (N7259, N7229, N1732, N2802, N5029);
or OR2 (N7260, N7250, N3365);
buf BUF1 (N7261, N7225);
nor NOR3 (N7262, N7251, N1401, N1922);
and AND2 (N7263, N7261, N3682);
and AND4 (N7264, N7257, N6684, N6033, N1866);
and AND4 (N7265, N7245, N5590, N7107, N1319);
nor NOR4 (N7266, N7262, N4071, N1244, N3034);
nand NAND4 (N7267, N7258, N5229, N1833, N4295);
or OR3 (N7268, N7252, N2288, N5951);
or OR4 (N7269, N7267, N3663, N775, N1698);
xor XOR2 (N7270, N7240, N1008);
buf BUF1 (N7271, N7269);
nor NOR3 (N7272, N7263, N2158, N4206);
or OR4 (N7273, N7270, N3556, N6732, N5116);
nor NOR2 (N7274, N7265, N5297);
and AND2 (N7275, N7268, N3888);
nand NAND4 (N7276, N7256, N3857, N6956, N2426);
xor XOR2 (N7277, N7266, N1846);
and AND2 (N7278, N7272, N6922);
not NOT1 (N7279, N7275);
buf BUF1 (N7280, N7279);
buf BUF1 (N7281, N7273);
and AND3 (N7282, N7274, N4915, N4104);
nand NAND3 (N7283, N7260, N4037, N150);
buf BUF1 (N7284, N7278);
xor XOR2 (N7285, N7284, N6112);
and AND3 (N7286, N7280, N1641, N6076);
nor NOR4 (N7287, N7277, N562, N5580, N5559);
not NOT1 (N7288, N7282);
not NOT1 (N7289, N7281);
nor NOR3 (N7290, N7283, N6460, N2026);
nor NOR4 (N7291, N7287, N1573, N2402, N3433);
buf BUF1 (N7292, N7285);
and AND3 (N7293, N7292, N1685, N2697);
xor XOR2 (N7294, N7289, N7143);
xor XOR2 (N7295, N7276, N2156);
nand NAND2 (N7296, N7295, N4347);
nor NOR2 (N7297, N7290, N1509);
not NOT1 (N7298, N7286);
nand NAND4 (N7299, N7291, N1339, N3131, N6922);
nor NOR2 (N7300, N7299, N4211);
nand NAND2 (N7301, N7297, N5661);
not NOT1 (N7302, N7300);
and AND3 (N7303, N7296, N3783, N6780);
and AND3 (N7304, N7264, N1404, N46);
nor NOR2 (N7305, N7302, N912);
nand NAND2 (N7306, N7304, N7227);
xor XOR2 (N7307, N7306, N3164);
nor NOR2 (N7308, N7293, N4409);
and AND2 (N7309, N7308, N2739);
nor NOR3 (N7310, N7259, N399, N838);
xor XOR2 (N7311, N7310, N4471);
nand NAND4 (N7312, N7301, N4566, N5864, N887);
or OR2 (N7313, N7298, N3939);
not NOT1 (N7314, N7288);
or OR2 (N7315, N7314, N1506);
nand NAND4 (N7316, N7271, N3605, N7313, N1097);
and AND3 (N7317, N3063, N5173, N97);
xor XOR2 (N7318, N7303, N1822);
not NOT1 (N7319, N7294);
nor NOR4 (N7320, N7305, N1395, N1977, N3145);
and AND3 (N7321, N7316, N3080, N6502);
nand NAND3 (N7322, N7318, N589, N3322);
nand NAND4 (N7323, N7315, N4800, N4390, N4161);
not NOT1 (N7324, N7319);
and AND4 (N7325, N7322, N759, N959, N991);
and AND4 (N7326, N7323, N2749, N6393, N4652);
buf BUF1 (N7327, N7326);
xor XOR2 (N7328, N7325, N68);
nand NAND3 (N7329, N7327, N4123, N1204);
buf BUF1 (N7330, N7329);
buf BUF1 (N7331, N7321);
nor NOR3 (N7332, N7317, N179, N2064);
nand NAND3 (N7333, N7328, N1679, N1580);
nor NOR2 (N7334, N7311, N4065);
nand NAND4 (N7335, N7324, N3277, N6564, N6263);
buf BUF1 (N7336, N7309);
nand NAND2 (N7337, N7333, N2528);
not NOT1 (N7338, N7330);
or OR2 (N7339, N7338, N845);
and AND2 (N7340, N7320, N2221);
buf BUF1 (N7341, N7331);
or OR3 (N7342, N7339, N5571, N6894);
nand NAND4 (N7343, N7334, N998, N6754, N3107);
nor NOR4 (N7344, N7307, N7338, N1123, N577);
xor XOR2 (N7345, N7342, N5772);
nand NAND3 (N7346, N7345, N638, N2601);
and AND3 (N7347, N7346, N3423, N3157);
xor XOR2 (N7348, N7343, N3481);
and AND4 (N7349, N7312, N5627, N2816, N1021);
buf BUF1 (N7350, N7348);
xor XOR2 (N7351, N7349, N7227);
xor XOR2 (N7352, N7344, N1756);
and AND3 (N7353, N7336, N6467, N2972);
not NOT1 (N7354, N7335);
nor NOR2 (N7355, N7352, N1955);
and AND3 (N7356, N7355, N4674, N5312);
not NOT1 (N7357, N7340);
xor XOR2 (N7358, N7356, N2265);
nor NOR2 (N7359, N7353, N6553);
nor NOR4 (N7360, N7341, N2819, N316, N158);
and AND2 (N7361, N7351, N1782);
nor NOR2 (N7362, N7347, N2744);
or OR3 (N7363, N7362, N1774, N379);
or OR4 (N7364, N7350, N6214, N1155, N821);
nand NAND3 (N7365, N7361, N1106, N753);
or OR3 (N7366, N7365, N6352, N3532);
not NOT1 (N7367, N7364);
buf BUF1 (N7368, N7363);
nand NAND3 (N7369, N7360, N3842, N337);
or OR2 (N7370, N7354, N846);
buf BUF1 (N7371, N7369);
xor XOR2 (N7372, N7359, N1678);
and AND4 (N7373, N7371, N468, N6518, N4700);
nor NOR2 (N7374, N7368, N6492);
buf BUF1 (N7375, N7370);
nand NAND3 (N7376, N7366, N782, N6853);
or OR2 (N7377, N7332, N6625);
buf BUF1 (N7378, N7367);
xor XOR2 (N7379, N7376, N3307);
or OR2 (N7380, N7372, N1444);
xor XOR2 (N7381, N7358, N5402);
buf BUF1 (N7382, N7378);
and AND2 (N7383, N7377, N3649);
not NOT1 (N7384, N7373);
buf BUF1 (N7385, N7379);
buf BUF1 (N7386, N7385);
nand NAND2 (N7387, N7383, N2285);
and AND4 (N7388, N7382, N5334, N6994, N4812);
or OR2 (N7389, N7388, N2250);
or OR3 (N7390, N7386, N5386, N3876);
buf BUF1 (N7391, N7374);
and AND4 (N7392, N7381, N13, N201, N206);
xor XOR2 (N7393, N7389, N6186);
and AND2 (N7394, N7390, N5078);
or OR3 (N7395, N7357, N3078, N1843);
buf BUF1 (N7396, N7391);
xor XOR2 (N7397, N7392, N4737);
not NOT1 (N7398, N7397);
nor NOR4 (N7399, N7393, N1355, N1155, N1429);
buf BUF1 (N7400, N7380);
nand NAND2 (N7401, N7400, N775);
xor XOR2 (N7402, N7396, N4433);
nor NOR4 (N7403, N7401, N5799, N6754, N4806);
and AND4 (N7404, N7399, N5194, N4807, N6001);
nand NAND2 (N7405, N7398, N7298);
or OR2 (N7406, N7403, N2387);
not NOT1 (N7407, N7337);
buf BUF1 (N7408, N7387);
and AND3 (N7409, N7394, N2133, N933);
or OR4 (N7410, N7375, N1956, N2431, N1417);
not NOT1 (N7411, N7409);
buf BUF1 (N7412, N7410);
nand NAND2 (N7413, N7405, N4919);
or OR4 (N7414, N7395, N1912, N4668, N631);
xor XOR2 (N7415, N7413, N6417);
nand NAND3 (N7416, N7406, N40, N221);
nand NAND4 (N7417, N7407, N6336, N1349, N5984);
nand NAND2 (N7418, N7402, N3769);
and AND3 (N7419, N7411, N3506, N969);
or OR2 (N7420, N7384, N3982);
and AND3 (N7421, N7412, N1051, N3828);
and AND2 (N7422, N7418, N4852);
not NOT1 (N7423, N7422);
nor NOR3 (N7424, N7419, N2873, N6263);
buf BUF1 (N7425, N7414);
xor XOR2 (N7426, N7421, N1419);
not NOT1 (N7427, N7420);
xor XOR2 (N7428, N7425, N7049);
not NOT1 (N7429, N7415);
not NOT1 (N7430, N7427);
not NOT1 (N7431, N7416);
xor XOR2 (N7432, N7417, N5904);
nor NOR2 (N7433, N7429, N6497);
nor NOR2 (N7434, N7423, N751);
nand NAND3 (N7435, N7432, N2889, N7235);
or OR3 (N7436, N7428, N347, N1440);
buf BUF1 (N7437, N7404);
nand NAND2 (N7438, N7430, N2802);
nor NOR4 (N7439, N7436, N2354, N3911, N33);
xor XOR2 (N7440, N7435, N3366);
buf BUF1 (N7441, N7437);
and AND4 (N7442, N7431, N4244, N1570, N3820);
not NOT1 (N7443, N7424);
or OR2 (N7444, N7408, N2499);
and AND4 (N7445, N7438, N6545, N5476, N2955);
nor NOR3 (N7446, N7433, N3717, N5572);
nand NAND4 (N7447, N7442, N830, N6568, N2253);
xor XOR2 (N7448, N7446, N5723);
xor XOR2 (N7449, N7444, N2205);
or OR2 (N7450, N7426, N5251);
nor NOR2 (N7451, N7447, N5166);
xor XOR2 (N7452, N7440, N489);
and AND4 (N7453, N7449, N5859, N5952, N4059);
nor NOR2 (N7454, N7443, N6437);
not NOT1 (N7455, N7434);
and AND4 (N7456, N7453, N614, N6284, N7163);
xor XOR2 (N7457, N7452, N2597);
not NOT1 (N7458, N7448);
buf BUF1 (N7459, N7457);
xor XOR2 (N7460, N7445, N666);
or OR3 (N7461, N7441, N3083, N5760);
buf BUF1 (N7462, N7451);
nand NAND4 (N7463, N7439, N4509, N5259, N2554);
and AND3 (N7464, N7462, N4423, N6820);
and AND3 (N7465, N7461, N84, N1482);
and AND3 (N7466, N7456, N1663, N7445);
buf BUF1 (N7467, N7464);
nor NOR2 (N7468, N7454, N125);
or OR3 (N7469, N7463, N7441, N7282);
xor XOR2 (N7470, N7468, N5904);
not NOT1 (N7471, N7460);
xor XOR2 (N7472, N7469, N6052);
buf BUF1 (N7473, N7450);
or OR2 (N7474, N7473, N2244);
nand NAND3 (N7475, N7471, N1892, N4521);
nand NAND2 (N7476, N7472, N347);
xor XOR2 (N7477, N7467, N513);
not NOT1 (N7478, N7475);
buf BUF1 (N7479, N7465);
buf BUF1 (N7480, N7479);
or OR4 (N7481, N7466, N5551, N5458, N7386);
buf BUF1 (N7482, N7480);
and AND2 (N7483, N7470, N639);
xor XOR2 (N7484, N7483, N1926);
xor XOR2 (N7485, N7482, N3206);
or OR4 (N7486, N7459, N3367, N4962, N3293);
and AND2 (N7487, N7476, N1121);
xor XOR2 (N7488, N7455, N2276);
not NOT1 (N7489, N7488);
not NOT1 (N7490, N7474);
xor XOR2 (N7491, N7481, N1016);
not NOT1 (N7492, N7484);
and AND4 (N7493, N7485, N1474, N406, N6244);
and AND3 (N7494, N7493, N7109, N2401);
or OR2 (N7495, N7477, N1639);
xor XOR2 (N7496, N7478, N4301);
nand NAND3 (N7497, N7494, N1261, N2019);
not NOT1 (N7498, N7491);
or OR3 (N7499, N7496, N3822, N7242);
buf BUF1 (N7500, N7487);
or OR3 (N7501, N7489, N542, N1371);
xor XOR2 (N7502, N7495, N2630);
and AND4 (N7503, N7486, N5440, N1346, N5816);
buf BUF1 (N7504, N7497);
nor NOR3 (N7505, N7492, N2335, N3521);
buf BUF1 (N7506, N7502);
and AND4 (N7507, N7499, N2412, N5949, N7224);
buf BUF1 (N7508, N7498);
buf BUF1 (N7509, N7505);
nand NAND4 (N7510, N7507, N5042, N6984, N7302);
or OR4 (N7511, N7501, N4430, N3176, N3774);
and AND3 (N7512, N7490, N4100, N4660);
xor XOR2 (N7513, N7500, N3797);
xor XOR2 (N7514, N7510, N3773);
or OR4 (N7515, N7503, N5616, N4620, N3656);
nor NOR4 (N7516, N7508, N5607, N1262, N704);
nand NAND4 (N7517, N7515, N1771, N5797, N2216);
and AND2 (N7518, N7509, N3189);
or OR4 (N7519, N7514, N4109, N4752, N72);
xor XOR2 (N7520, N7518, N5239);
buf BUF1 (N7521, N7517);
buf BUF1 (N7522, N7504);
or OR2 (N7523, N7506, N2531);
nor NOR3 (N7524, N7519, N5727, N166);
not NOT1 (N7525, N7512);
or OR4 (N7526, N7516, N5399, N5494, N4257);
nor NOR3 (N7527, N7521, N4153, N5904);
and AND4 (N7528, N7522, N4133, N2668, N343);
and AND3 (N7529, N7527, N1552, N6878);
buf BUF1 (N7530, N7524);
and AND3 (N7531, N7529, N1078, N4525);
buf BUF1 (N7532, N7531);
nor NOR2 (N7533, N7523, N1532);
nand NAND2 (N7534, N7525, N4113);
buf BUF1 (N7535, N7520);
xor XOR2 (N7536, N7528, N4996);
nand NAND3 (N7537, N7526, N3952, N7128);
and AND4 (N7538, N7534, N5444, N1288, N3158);
or OR4 (N7539, N7530, N7028, N1160, N5859);
not NOT1 (N7540, N7537);
xor XOR2 (N7541, N7540, N6156);
nor NOR4 (N7542, N7458, N1599, N2966, N4032);
buf BUF1 (N7543, N7536);
nor NOR2 (N7544, N7532, N5906);
or OR4 (N7545, N7511, N407, N3208, N4387);
nand NAND3 (N7546, N7541, N2156, N1493);
nand NAND4 (N7547, N7533, N6876, N2188, N6989);
buf BUF1 (N7548, N7535);
nand NAND3 (N7549, N7543, N5174, N1507);
xor XOR2 (N7550, N7538, N1368);
or OR3 (N7551, N7546, N4345, N3646);
or OR4 (N7552, N7547, N1232, N7225, N6650);
nor NOR2 (N7553, N7544, N6884);
xor XOR2 (N7554, N7513, N4032);
nand NAND3 (N7555, N7550, N987, N4417);
xor XOR2 (N7556, N7539, N5166);
not NOT1 (N7557, N7542);
buf BUF1 (N7558, N7553);
or OR3 (N7559, N7555, N6965, N2185);
nor NOR2 (N7560, N7549, N688);
nor NOR4 (N7561, N7559, N6795, N3751, N5053);
xor XOR2 (N7562, N7561, N5150);
or OR3 (N7563, N7557, N266, N5341);
xor XOR2 (N7564, N7558, N2051);
and AND4 (N7565, N7551, N7513, N5489, N2509);
or OR2 (N7566, N7563, N6872);
nor NOR3 (N7567, N7554, N4701, N4236);
xor XOR2 (N7568, N7566, N1257);
buf BUF1 (N7569, N7565);
and AND2 (N7570, N7569, N451);
not NOT1 (N7571, N7568);
xor XOR2 (N7572, N7545, N6719);
and AND3 (N7573, N7570, N6825, N2795);
not NOT1 (N7574, N7572);
buf BUF1 (N7575, N7564);
nand NAND3 (N7576, N7552, N1177, N1788);
xor XOR2 (N7577, N7573, N1597);
not NOT1 (N7578, N7562);
not NOT1 (N7579, N7576);
nor NOR4 (N7580, N7575, N6121, N2229, N4491);
or OR4 (N7581, N7571, N4233, N568, N682);
or OR4 (N7582, N7548, N1383, N3708, N1960);
or OR4 (N7583, N7580, N5874, N6758, N1906);
and AND3 (N7584, N7583, N2381, N3804);
buf BUF1 (N7585, N7582);
buf BUF1 (N7586, N7577);
nor NOR2 (N7587, N7560, N7070);
or OR3 (N7588, N7574, N1325, N6165);
and AND4 (N7589, N7584, N484, N400, N263);
nand NAND4 (N7590, N7589, N3491, N1814, N1562);
buf BUF1 (N7591, N7587);
and AND3 (N7592, N7588, N6727, N1491);
not NOT1 (N7593, N7567);
not NOT1 (N7594, N7581);
not NOT1 (N7595, N7590);
nor NOR3 (N7596, N7585, N2610, N6265);
nand NAND3 (N7597, N7594, N6074, N4165);
nand NAND3 (N7598, N7593, N7569, N6081);
nand NAND2 (N7599, N7592, N4352);
buf BUF1 (N7600, N7591);
nand NAND3 (N7601, N7595, N5399, N5430);
or OR3 (N7602, N7601, N4930, N4653);
nor NOR3 (N7603, N7578, N3835, N2884);
xor XOR2 (N7604, N7603, N7182);
and AND4 (N7605, N7597, N126, N1813, N1462);
nor NOR4 (N7606, N7579, N6025, N4841, N2584);
xor XOR2 (N7607, N7596, N2370);
buf BUF1 (N7608, N7606);
nor NOR2 (N7609, N7602, N6320);
nor NOR4 (N7610, N7598, N1108, N5216, N3495);
not NOT1 (N7611, N7599);
xor XOR2 (N7612, N7605, N1317);
or OR3 (N7613, N7610, N4969, N5218);
xor XOR2 (N7614, N7586, N2718);
and AND3 (N7615, N7607, N5709, N5485);
xor XOR2 (N7616, N7612, N4639);
and AND2 (N7617, N7611, N5483);
xor XOR2 (N7618, N7604, N4127);
nor NOR2 (N7619, N7600, N2640);
or OR4 (N7620, N7614, N5372, N643, N6891);
or OR2 (N7621, N7609, N423);
or OR2 (N7622, N7617, N3545);
nand NAND4 (N7623, N7618, N4715, N7453, N1534);
not NOT1 (N7624, N7608);
xor XOR2 (N7625, N7615, N4506);
and AND4 (N7626, N7556, N691, N2926, N4542);
not NOT1 (N7627, N7616);
not NOT1 (N7628, N7622);
nor NOR2 (N7629, N7627, N2134);
buf BUF1 (N7630, N7628);
nor NOR2 (N7631, N7625, N4439);
xor XOR2 (N7632, N7623, N1223);
xor XOR2 (N7633, N7624, N3383);
or OR3 (N7634, N7631, N2588, N3568);
nor NOR3 (N7635, N7633, N5718, N5536);
buf BUF1 (N7636, N7613);
and AND4 (N7637, N7621, N2908, N5639, N1595);
nor NOR4 (N7638, N7620, N2249, N1838, N6369);
or OR3 (N7639, N7626, N2258, N6681);
not NOT1 (N7640, N7632);
buf BUF1 (N7641, N7637);
nor NOR2 (N7642, N7629, N942);
xor XOR2 (N7643, N7642, N5509);
and AND4 (N7644, N7639, N7359, N539, N5507);
buf BUF1 (N7645, N7641);
or OR3 (N7646, N7638, N1421, N6911);
nor NOR3 (N7647, N7643, N4601, N6375);
nor NOR3 (N7648, N7645, N279, N6817);
and AND4 (N7649, N7648, N7160, N7522, N3030);
xor XOR2 (N7650, N7644, N2467);
xor XOR2 (N7651, N7649, N7177);
and AND4 (N7652, N7634, N5255, N5948, N3901);
not NOT1 (N7653, N7650);
nand NAND2 (N7654, N7653, N6876);
and AND4 (N7655, N7652, N7316, N5746, N516);
and AND3 (N7656, N7655, N7489, N545);
and AND3 (N7657, N7654, N1807, N5995);
nand NAND3 (N7658, N7651, N6292, N4607);
nand NAND4 (N7659, N7635, N2097, N5921, N5829);
or OR4 (N7660, N7640, N2120, N4819, N3444);
buf BUF1 (N7661, N7660);
not NOT1 (N7662, N7619);
buf BUF1 (N7663, N7646);
xor XOR2 (N7664, N7656, N217);
buf BUF1 (N7665, N7664);
xor XOR2 (N7666, N7659, N6947);
buf BUF1 (N7667, N7630);
xor XOR2 (N7668, N7662, N363);
not NOT1 (N7669, N7663);
or OR2 (N7670, N7658, N2159);
not NOT1 (N7671, N7668);
nand NAND2 (N7672, N7666, N7460);
not NOT1 (N7673, N7661);
nor NOR4 (N7674, N7636, N6284, N4400, N6570);
nand NAND4 (N7675, N7671, N324, N910, N4420);
nor NOR2 (N7676, N7672, N6096);
nor NOR4 (N7677, N7647, N6842, N1939, N5284);
or OR2 (N7678, N7677, N6814);
or OR2 (N7679, N7674, N3781);
or OR2 (N7680, N7678, N5026);
nand NAND2 (N7681, N7669, N4647);
nand NAND2 (N7682, N7673, N5763);
xor XOR2 (N7683, N7679, N3095);
not NOT1 (N7684, N7667);
nand NAND2 (N7685, N7680, N6197);
xor XOR2 (N7686, N7665, N2311);
and AND3 (N7687, N7686, N2220, N6984);
buf BUF1 (N7688, N7657);
or OR2 (N7689, N7681, N4792);
nand NAND4 (N7690, N7676, N7082, N4060, N5791);
or OR4 (N7691, N7690, N996, N6106, N624);
not NOT1 (N7692, N7684);
xor XOR2 (N7693, N7689, N2470);
and AND3 (N7694, N7693, N2427, N4185);
xor XOR2 (N7695, N7685, N5176);
buf BUF1 (N7696, N7675);
nand NAND3 (N7697, N7687, N313, N6733);
or OR4 (N7698, N7697, N6316, N412, N3510);
nor NOR2 (N7699, N7682, N5839);
not NOT1 (N7700, N7692);
and AND2 (N7701, N7700, N2705);
and AND2 (N7702, N7688, N6180);
or OR2 (N7703, N7696, N1835);
not NOT1 (N7704, N7698);
nand NAND3 (N7705, N7695, N3608, N3231);
or OR3 (N7706, N7702, N4575, N1101);
not NOT1 (N7707, N7701);
or OR4 (N7708, N7694, N23, N1700, N1368);
nand NAND4 (N7709, N7670, N765, N2518, N7091);
and AND4 (N7710, N7706, N1204, N1329, N5947);
or OR2 (N7711, N7704, N6483);
or OR4 (N7712, N7709, N4759, N4532, N4433);
nand NAND4 (N7713, N7691, N2363, N5153, N5444);
and AND3 (N7714, N7699, N6395, N1904);
nor NOR2 (N7715, N7714, N4903);
and AND2 (N7716, N7705, N7204);
nand NAND4 (N7717, N7713, N4386, N3531, N7154);
nor NOR4 (N7718, N7707, N56, N386, N332);
xor XOR2 (N7719, N7715, N5251);
nor NOR3 (N7720, N7711, N1992, N3177);
nor NOR3 (N7721, N7717, N6619, N2329);
nand NAND3 (N7722, N7720, N4328, N3735);
and AND4 (N7723, N7708, N4481, N3655, N1076);
nand NAND2 (N7724, N7712, N2818);
or OR3 (N7725, N7724, N950, N2177);
xor XOR2 (N7726, N7683, N6780);
and AND4 (N7727, N7703, N5808, N6474, N5232);
or OR2 (N7728, N7727, N3010);
buf BUF1 (N7729, N7718);
buf BUF1 (N7730, N7729);
or OR3 (N7731, N7726, N2098, N3972);
or OR3 (N7732, N7719, N423, N560);
xor XOR2 (N7733, N7731, N7626);
buf BUF1 (N7734, N7722);
or OR4 (N7735, N7734, N3025, N2527, N6829);
and AND4 (N7736, N7728, N6933, N491, N5230);
or OR3 (N7737, N7725, N5080, N3278);
nor NOR3 (N7738, N7733, N1301, N6307);
buf BUF1 (N7739, N7732);
nor NOR4 (N7740, N7736, N5071, N2542, N4999);
not NOT1 (N7741, N7740);
nand NAND3 (N7742, N7739, N7333, N7242);
buf BUF1 (N7743, N7737);
not NOT1 (N7744, N7742);
and AND3 (N7745, N7744, N4751, N4311);
buf BUF1 (N7746, N7741);
not NOT1 (N7747, N7721);
nor NOR2 (N7748, N7746, N6513);
nand NAND4 (N7749, N7747, N5366, N4407, N3099);
nand NAND3 (N7750, N7743, N5980, N2016);
not NOT1 (N7751, N7749);
nor NOR3 (N7752, N7745, N3946, N1566);
nor NOR3 (N7753, N7730, N6751, N4845);
buf BUF1 (N7754, N7735);
buf BUF1 (N7755, N7753);
buf BUF1 (N7756, N7755);
nor NOR4 (N7757, N7716, N5940, N248, N1437);
not NOT1 (N7758, N7750);
or OR4 (N7759, N7754, N1532, N3939, N4794);
xor XOR2 (N7760, N7758, N3205);
nand NAND3 (N7761, N7760, N1856, N4701);
nor NOR3 (N7762, N7759, N5003, N2465);
nor NOR2 (N7763, N7762, N6635);
xor XOR2 (N7764, N7723, N4216);
nor NOR3 (N7765, N7761, N5626, N1023);
nor NOR4 (N7766, N7756, N3151, N6058, N1129);
or OR3 (N7767, N7757, N719, N5884);
nor NOR2 (N7768, N7710, N1233);
xor XOR2 (N7769, N7751, N4925);
buf BUF1 (N7770, N7768);
nor NOR3 (N7771, N7765, N970, N6958);
nand NAND4 (N7772, N7770, N2475, N6174, N244);
and AND2 (N7773, N7752, N2194);
and AND2 (N7774, N7771, N1605);
nand NAND4 (N7775, N7769, N5701, N6389, N987);
buf BUF1 (N7776, N7773);
not NOT1 (N7777, N7766);
or OR3 (N7778, N7776, N4708, N7740);
not NOT1 (N7779, N7748);
nor NOR2 (N7780, N7775, N2259);
or OR3 (N7781, N7779, N6842, N84);
and AND2 (N7782, N7781, N7196);
nor NOR2 (N7783, N7780, N7755);
buf BUF1 (N7784, N7783);
not NOT1 (N7785, N7763);
xor XOR2 (N7786, N7764, N2553);
nand NAND2 (N7787, N7785, N927);
and AND4 (N7788, N7774, N1906, N505, N1039);
nor NOR2 (N7789, N7777, N1862);
nor NOR2 (N7790, N7789, N2509);
buf BUF1 (N7791, N7738);
nand NAND3 (N7792, N7778, N6467, N1823);
and AND4 (N7793, N7782, N4259, N5212, N5641);
xor XOR2 (N7794, N7772, N6236);
xor XOR2 (N7795, N7794, N6988);
buf BUF1 (N7796, N7795);
and AND4 (N7797, N7790, N2541, N6277, N307);
buf BUF1 (N7798, N7797);
xor XOR2 (N7799, N7798, N3147);
xor XOR2 (N7800, N7799, N1712);
nand NAND2 (N7801, N7788, N934);
nor NOR3 (N7802, N7787, N3501, N7315);
xor XOR2 (N7803, N7791, N2483);
nor NOR4 (N7804, N7793, N6068, N6672, N3776);
and AND4 (N7805, N7802, N2786, N3621, N6627);
nand NAND2 (N7806, N7804, N6296);
not NOT1 (N7807, N7784);
and AND3 (N7808, N7792, N1417, N1943);
nand NAND2 (N7809, N7800, N97);
nand NAND2 (N7810, N7796, N4920);
or OR4 (N7811, N7807, N3867, N343, N6739);
and AND2 (N7812, N7808, N5770);
nor NOR4 (N7813, N7810, N4355, N6064, N7001);
nand NAND4 (N7814, N7801, N4816, N1236, N1586);
not NOT1 (N7815, N7811);
nor NOR3 (N7816, N7809, N554, N3561);
and AND4 (N7817, N7816, N266, N1653, N1552);
or OR3 (N7818, N7786, N535, N5655);
xor XOR2 (N7819, N7806, N5374);
not NOT1 (N7820, N7817);
buf BUF1 (N7821, N7767);
nand NAND4 (N7822, N7819, N2273, N2257, N1796);
nor NOR2 (N7823, N7813, N6596);
nor NOR3 (N7824, N7814, N1570, N3107);
nand NAND2 (N7825, N7818, N7136);
or OR2 (N7826, N7824, N37);
xor XOR2 (N7827, N7823, N5498);
nor NOR4 (N7828, N7822, N5173, N6154, N4409);
nor NOR3 (N7829, N7828, N1212, N875);
xor XOR2 (N7830, N7826, N5156);
nand NAND4 (N7831, N7812, N3374, N7249, N1376);
not NOT1 (N7832, N7829);
xor XOR2 (N7833, N7830, N730);
buf BUF1 (N7834, N7832);
and AND3 (N7835, N7805, N4206, N7814);
buf BUF1 (N7836, N7803);
buf BUF1 (N7837, N7831);
nor NOR4 (N7838, N7820, N557, N194, N5464);
nand NAND2 (N7839, N7834, N3544);
nor NOR3 (N7840, N7839, N542, N3710);
nor NOR2 (N7841, N7837, N332);
and AND2 (N7842, N7835, N2797);
buf BUF1 (N7843, N7825);
not NOT1 (N7844, N7836);
xor XOR2 (N7845, N7840, N465);
nor NOR2 (N7846, N7842, N3975);
or OR2 (N7847, N7843, N996);
nor NOR2 (N7848, N7844, N6091);
nor NOR3 (N7849, N7821, N4321, N1891);
or OR4 (N7850, N7848, N5589, N5502, N6236);
nor NOR3 (N7851, N7849, N4277, N3821);
xor XOR2 (N7852, N7847, N25);
buf BUF1 (N7853, N7845);
or OR3 (N7854, N7833, N242, N6773);
nor NOR2 (N7855, N7841, N3060);
or OR4 (N7856, N7846, N2073, N4630, N6550);
nand NAND2 (N7857, N7851, N1905);
buf BUF1 (N7858, N7857);
xor XOR2 (N7859, N7858, N5738);
nand NAND4 (N7860, N7815, N6946, N6116, N4626);
nor NOR2 (N7861, N7859, N1257);
nand NAND2 (N7862, N7856, N2183);
not NOT1 (N7863, N7860);
nand NAND4 (N7864, N7863, N7261, N1502, N7590);
buf BUF1 (N7865, N7838);
xor XOR2 (N7866, N7827, N6277);
and AND4 (N7867, N7864, N7396, N7342, N1949);
nor NOR2 (N7868, N7853, N3411);
buf BUF1 (N7869, N7854);
and AND2 (N7870, N7855, N4035);
nand NAND4 (N7871, N7867, N1185, N4959, N4963);
not NOT1 (N7872, N7865);
not NOT1 (N7873, N7870);
nor NOR2 (N7874, N7872, N7395);
buf BUF1 (N7875, N7852);
nand NAND2 (N7876, N7875, N2361);
nor NOR3 (N7877, N7873, N3592, N5076);
buf BUF1 (N7878, N7876);
xor XOR2 (N7879, N7861, N2740);
xor XOR2 (N7880, N7868, N7118);
or OR4 (N7881, N7869, N7089, N6208, N6574);
xor XOR2 (N7882, N7874, N2109);
nand NAND3 (N7883, N7882, N1240, N6161);
nand NAND2 (N7884, N7879, N4176);
buf BUF1 (N7885, N7884);
nand NAND4 (N7886, N7871, N7371, N3218, N1824);
not NOT1 (N7887, N7850);
nor NOR3 (N7888, N7877, N4054, N4357);
nor NOR4 (N7889, N7885, N1291, N2881, N4003);
and AND3 (N7890, N7878, N6041, N3158);
xor XOR2 (N7891, N7862, N1250);
xor XOR2 (N7892, N7881, N800);
nor NOR3 (N7893, N7889, N2154, N133);
xor XOR2 (N7894, N7891, N1929);
nor NOR3 (N7895, N7894, N3883, N6556);
not NOT1 (N7896, N7888);
nand NAND2 (N7897, N7890, N6824);
not NOT1 (N7898, N7893);
and AND3 (N7899, N7887, N2731, N2882);
buf BUF1 (N7900, N7898);
xor XOR2 (N7901, N7896, N3397);
xor XOR2 (N7902, N7900, N939);
xor XOR2 (N7903, N7899, N2702);
nand NAND4 (N7904, N7880, N4191, N4948, N3605);
or OR3 (N7905, N7903, N5092, N5620);
buf BUF1 (N7906, N7897);
nand NAND4 (N7907, N7904, N5043, N1221, N3057);
nand NAND3 (N7908, N7901, N7093, N7114);
and AND3 (N7909, N7907, N696, N4899);
nor NOR3 (N7910, N7883, N1181, N7405);
xor XOR2 (N7911, N7866, N1248);
or OR3 (N7912, N7895, N5009, N3781);
not NOT1 (N7913, N7892);
and AND2 (N7914, N7913, N4667);
buf BUF1 (N7915, N7908);
xor XOR2 (N7916, N7905, N3214);
nand NAND4 (N7917, N7911, N798, N2023, N3955);
and AND3 (N7918, N7914, N6926, N6238);
xor XOR2 (N7919, N7909, N5013);
xor XOR2 (N7920, N7906, N986);
not NOT1 (N7921, N7916);
and AND3 (N7922, N7910, N717, N4314);
nand NAND2 (N7923, N7902, N2106);
nand NAND4 (N7924, N7886, N1944, N924, N3885);
nand NAND3 (N7925, N7923, N5015, N877);
nand NAND2 (N7926, N7918, N1792);
nand NAND4 (N7927, N7925, N3058, N4610, N2060);
xor XOR2 (N7928, N7915, N684);
not NOT1 (N7929, N7920);
buf BUF1 (N7930, N7922);
nor NOR3 (N7931, N7917, N5653, N204);
xor XOR2 (N7932, N7927, N2660);
and AND2 (N7933, N7926, N2190);
and AND3 (N7934, N7932, N5457, N2438);
nand NAND2 (N7935, N7931, N4744);
nor NOR2 (N7936, N7928, N6780);
xor XOR2 (N7937, N7919, N6615);
buf BUF1 (N7938, N7929);
or OR4 (N7939, N7934, N3073, N5446, N7404);
and AND2 (N7940, N7930, N5296);
nand NAND3 (N7941, N7921, N2583, N3373);
and AND3 (N7942, N7933, N4019, N2584);
xor XOR2 (N7943, N7939, N6770);
xor XOR2 (N7944, N7942, N196);
nor NOR4 (N7945, N7941, N2719, N3224, N4192);
buf BUF1 (N7946, N7935);
nand NAND3 (N7947, N7940, N2171, N232);
not NOT1 (N7948, N7944);
xor XOR2 (N7949, N7947, N1800);
xor XOR2 (N7950, N7946, N6747);
xor XOR2 (N7951, N7937, N2339);
nand NAND2 (N7952, N7948, N5771);
nand NAND4 (N7953, N7938, N5005, N7917, N3805);
buf BUF1 (N7954, N7945);
buf BUF1 (N7955, N7952);
and AND2 (N7956, N7949, N2022);
not NOT1 (N7957, N7953);
xor XOR2 (N7958, N7912, N3778);
and AND2 (N7959, N7954, N4798);
and AND2 (N7960, N7951, N3333);
xor XOR2 (N7961, N7950, N5715);
not NOT1 (N7962, N7960);
buf BUF1 (N7963, N7962);
or OR4 (N7964, N7957, N6680, N2805, N3817);
xor XOR2 (N7965, N7963, N1380);
buf BUF1 (N7966, N7959);
nor NOR2 (N7967, N7965, N3163);
xor XOR2 (N7968, N7955, N864);
buf BUF1 (N7969, N7964);
or OR3 (N7970, N7969, N6605, N310);
xor XOR2 (N7971, N7966, N2274);
xor XOR2 (N7972, N7958, N7883);
nand NAND4 (N7973, N7961, N4541, N330, N5541);
not NOT1 (N7974, N7968);
and AND4 (N7975, N7924, N228, N4675, N6090);
not NOT1 (N7976, N7936);
nor NOR2 (N7977, N7975, N2200);
xor XOR2 (N7978, N7973, N3564);
nor NOR2 (N7979, N7970, N4939);
buf BUF1 (N7980, N7974);
not NOT1 (N7981, N7979);
xor XOR2 (N7982, N7956, N5875);
nor NOR3 (N7983, N7977, N6627, N3276);
and AND3 (N7984, N7943, N3621, N6878);
xor XOR2 (N7985, N7980, N7016);
nand NAND4 (N7986, N7971, N7890, N5902, N4270);
nand NAND3 (N7987, N7983, N1447, N1058);
not NOT1 (N7988, N7986);
or OR3 (N7989, N7987, N2245, N2933);
xor XOR2 (N7990, N7972, N5468);
not NOT1 (N7991, N7976);
nor NOR2 (N7992, N7988, N3910);
buf BUF1 (N7993, N7982);
not NOT1 (N7994, N7989);
xor XOR2 (N7995, N7981, N2836);
and AND3 (N7996, N7994, N1467, N7185);
buf BUF1 (N7997, N7990);
nand NAND3 (N7998, N7985, N7210, N1324);
nand NAND3 (N7999, N7998, N3498, N1294);
nand NAND4 (N8000, N7978, N6493, N2925, N1366);
xor XOR2 (N8001, N7999, N6388);
xor XOR2 (N8002, N7984, N4692);
buf BUF1 (N8003, N8002);
or OR4 (N8004, N7993, N1871, N1077, N5401);
or OR4 (N8005, N7991, N4070, N5170, N7249);
nor NOR4 (N8006, N8004, N3424, N1634, N7195);
buf BUF1 (N8007, N8005);
nor NOR2 (N8008, N8001, N5681);
or OR4 (N8009, N8003, N6448, N6066, N7259);
nand NAND2 (N8010, N8007, N897);
xor XOR2 (N8011, N7997, N2679);
or OR2 (N8012, N8011, N3509);
and AND4 (N8013, N8000, N3820, N7701, N7262);
nand NAND2 (N8014, N7995, N3891);
nor NOR3 (N8015, N8008, N3865, N4225);
not NOT1 (N8016, N8010);
nand NAND4 (N8017, N8006, N6504, N6816, N3732);
not NOT1 (N8018, N8015);
nand NAND2 (N8019, N8013, N7320);
xor XOR2 (N8020, N7996, N222);
and AND4 (N8021, N7967, N7716, N1500, N7135);
nand NAND4 (N8022, N8018, N1515, N7690, N6390);
endmodule