// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N784,N803,N804,N811,N794,N782,N809,N800,N806,N812;

and AND2 (N13, N8, N6);
xor XOR2 (N14, N6, N6);
nor NOR3 (N15, N6, N10, N14);
and AND2 (N16, N9, N12);
not NOT1 (N17, N5);
nor NOR3 (N18, N16, N11, N6);
buf BUF1 (N19, N17);
nand NAND4 (N20, N2, N16, N12, N6);
xor XOR2 (N21, N19, N5);
and AND2 (N22, N19, N1);
not NOT1 (N23, N2);
xor XOR2 (N24, N12, N17);
nor NOR4 (N25, N12, N22, N21, N3);
nor NOR3 (N26, N19, N12, N1);
nand NAND2 (N27, N14, N24);
or OR2 (N28, N19, N12);
nand NAND3 (N29, N11, N14, N4);
nand NAND3 (N30, N26, N4, N6);
buf BUF1 (N31, N25);
and AND2 (N32, N28, N15);
xor XOR2 (N33, N32, N7);
or OR3 (N34, N3, N27, N21);
and AND3 (N35, N20, N16, N7);
xor XOR2 (N36, N24, N10);
nor NOR3 (N37, N36, N10, N28);
and AND4 (N38, N18, N34, N34, N13);
or OR2 (N39, N33, N7);
buf BUF1 (N40, N25);
or OR3 (N41, N23, N6, N32);
nor NOR2 (N42, N21, N34);
nor NOR2 (N43, N31, N33);
nor NOR4 (N44, N29, N18, N5, N40);
not NOT1 (N45, N44);
not NOT1 (N46, N34);
and AND2 (N47, N46, N4);
not NOT1 (N48, N38);
and AND2 (N49, N48, N28);
or OR4 (N50, N39, N22, N29, N41);
nor NOR3 (N51, N20, N7, N26);
or OR2 (N52, N51, N25);
xor XOR2 (N53, N42, N27);
or OR3 (N54, N47, N27, N52);
and AND3 (N55, N16, N6, N1);
not NOT1 (N56, N35);
nand NAND3 (N57, N55, N33, N31);
xor XOR2 (N58, N57, N51);
not NOT1 (N59, N53);
or OR3 (N60, N50, N4, N44);
nor NOR3 (N61, N54, N60, N35);
buf BUF1 (N62, N43);
and AND3 (N63, N60, N55, N47);
buf BUF1 (N64, N30);
nor NOR3 (N65, N64, N64, N14);
nand NAND3 (N66, N63, N51, N64);
nor NOR3 (N67, N61, N44, N31);
or OR2 (N68, N67, N18);
or OR4 (N69, N65, N13, N25, N33);
nand NAND4 (N70, N49, N51, N67, N40);
xor XOR2 (N71, N66, N36);
and AND3 (N72, N62, N1, N28);
or OR3 (N73, N59, N51, N47);
and AND2 (N74, N37, N54);
not NOT1 (N75, N68);
or OR2 (N76, N56, N69);
buf BUF1 (N77, N10);
buf BUF1 (N78, N71);
nand NAND4 (N79, N73, N70, N69, N14);
xor XOR2 (N80, N22, N9);
and AND3 (N81, N75, N12, N37);
not NOT1 (N82, N81);
nand NAND2 (N83, N80, N36);
buf BUF1 (N84, N58);
and AND3 (N85, N77, N14, N74);
not NOT1 (N86, N68);
not NOT1 (N87, N84);
nand NAND4 (N88, N76, N19, N54, N31);
nor NOR4 (N89, N85, N41, N24, N53);
and AND4 (N90, N45, N82, N56, N15);
and AND2 (N91, N66, N62);
buf BUF1 (N92, N91);
buf BUF1 (N93, N87);
xor XOR2 (N94, N86, N44);
and AND4 (N95, N93, N39, N92, N49);
nand NAND2 (N96, N92, N70);
xor XOR2 (N97, N90, N68);
or OR4 (N98, N72, N33, N62, N36);
buf BUF1 (N99, N94);
nand NAND2 (N100, N98, N25);
and AND3 (N101, N79, N5, N20);
nor NOR4 (N102, N100, N47, N96, N29);
not NOT1 (N103, N98);
and AND4 (N104, N101, N43, N37, N65);
buf BUF1 (N105, N104);
and AND2 (N106, N89, N29);
nor NOR2 (N107, N97, N85);
buf BUF1 (N108, N78);
buf BUF1 (N109, N88);
nor NOR3 (N110, N109, N2, N5);
and AND2 (N111, N103, N7);
nor NOR4 (N112, N83, N7, N78, N77);
not NOT1 (N113, N95);
xor XOR2 (N114, N110, N73);
nor NOR3 (N115, N111, N94, N43);
nand NAND2 (N116, N105, N99);
buf BUF1 (N117, N68);
not NOT1 (N118, N117);
and AND2 (N119, N115, N57);
or OR2 (N120, N112, N85);
xor XOR2 (N121, N116, N116);
or OR4 (N122, N114, N91, N3, N116);
or OR4 (N123, N108, N103, N116, N6);
not NOT1 (N124, N102);
xor XOR2 (N125, N113, N79);
not NOT1 (N126, N120);
or OR2 (N127, N106, N109);
or OR2 (N128, N119, N44);
xor XOR2 (N129, N122, N93);
xor XOR2 (N130, N126, N81);
and AND3 (N131, N130, N61, N119);
not NOT1 (N132, N131);
buf BUF1 (N133, N125);
xor XOR2 (N134, N129, N92);
nand NAND3 (N135, N127, N124, N9);
nor NOR2 (N136, N44, N127);
xor XOR2 (N137, N134, N20);
and AND3 (N138, N107, N110, N106);
or OR2 (N139, N136, N112);
buf BUF1 (N140, N128);
nor NOR2 (N141, N133, N130);
nand NAND2 (N142, N118, N136);
xor XOR2 (N143, N138, N44);
and AND2 (N144, N137, N75);
buf BUF1 (N145, N139);
and AND2 (N146, N135, N125);
and AND4 (N147, N140, N95, N106, N132);
not NOT1 (N148, N53);
or OR3 (N149, N148, N19, N68);
and AND2 (N150, N149, N40);
and AND4 (N151, N142, N115, N105, N82);
nand NAND4 (N152, N143, N115, N74, N22);
nand NAND2 (N153, N145, N116);
nand NAND4 (N154, N123, N74, N12, N63);
nand NAND2 (N155, N153, N90);
buf BUF1 (N156, N155);
and AND3 (N157, N141, N69, N121);
nand NAND2 (N158, N72, N34);
nand NAND3 (N159, N157, N144, N22);
nor NOR3 (N160, N158, N114, N74);
buf BUF1 (N161, N159);
and AND2 (N162, N54, N129);
nor NOR4 (N163, N152, N124, N15, N66);
nand NAND4 (N164, N154, N162, N1, N117);
and AND4 (N165, N64, N14, N6, N35);
nand NAND4 (N166, N160, N10, N158, N74);
not NOT1 (N167, N164);
not NOT1 (N168, N163);
not NOT1 (N169, N165);
nand NAND3 (N170, N166, N29, N38);
buf BUF1 (N171, N161);
and AND4 (N172, N147, N106, N38, N57);
nand NAND2 (N173, N170, N33);
buf BUF1 (N174, N150);
nand NAND3 (N175, N173, N4, N80);
buf BUF1 (N176, N167);
nor NOR2 (N177, N172, N157);
not NOT1 (N178, N169);
or OR4 (N179, N171, N37, N153, N81);
and AND4 (N180, N178, N147, N123, N97);
buf BUF1 (N181, N179);
nor NOR2 (N182, N181, N74);
nand NAND3 (N183, N168, N171, N55);
buf BUF1 (N184, N175);
xor XOR2 (N185, N174, N71);
or OR2 (N186, N185, N61);
or OR4 (N187, N183, N63, N13, N165);
or OR3 (N188, N146, N183, N67);
xor XOR2 (N189, N186, N101);
nor NOR3 (N190, N187, N41, N56);
nand NAND2 (N191, N182, N60);
buf BUF1 (N192, N191);
buf BUF1 (N193, N180);
buf BUF1 (N194, N151);
buf BUF1 (N195, N192);
nand NAND4 (N196, N177, N69, N119, N49);
xor XOR2 (N197, N195, N144);
buf BUF1 (N198, N196);
nor NOR2 (N199, N197, N18);
buf BUF1 (N200, N199);
nor NOR4 (N201, N189, N99, N33, N12);
xor XOR2 (N202, N198, N144);
nand NAND3 (N203, N190, N59, N162);
nand NAND3 (N204, N203, N92, N43);
xor XOR2 (N205, N194, N132);
not NOT1 (N206, N176);
buf BUF1 (N207, N201);
nand NAND2 (N208, N207, N95);
xor XOR2 (N209, N202, N6);
xor XOR2 (N210, N188, N4);
buf BUF1 (N211, N156);
buf BUF1 (N212, N211);
buf BUF1 (N213, N212);
not NOT1 (N214, N210);
nor NOR2 (N215, N184, N182);
nand NAND3 (N216, N206, N147, N73);
xor XOR2 (N217, N204, N150);
and AND4 (N218, N209, N198, N118, N61);
nand NAND4 (N219, N215, N68, N207, N116);
not NOT1 (N220, N217);
and AND4 (N221, N193, N163, N176, N62);
nand NAND3 (N222, N205, N48, N80);
buf BUF1 (N223, N208);
and AND3 (N224, N213, N143, N146);
nand NAND2 (N225, N200, N22);
nand NAND3 (N226, N214, N171, N138);
and AND4 (N227, N216, N173, N149, N102);
buf BUF1 (N228, N220);
nor NOR2 (N229, N218, N73);
and AND4 (N230, N225, N61, N56, N109);
nand NAND4 (N231, N224, N35, N138, N42);
or OR4 (N232, N227, N175, N121, N19);
nand NAND4 (N233, N223, N102, N223, N20);
buf BUF1 (N234, N230);
xor XOR2 (N235, N226, N224);
or OR4 (N236, N229, N100, N134, N201);
xor XOR2 (N237, N219, N48);
and AND4 (N238, N232, N204, N194, N92);
xor XOR2 (N239, N233, N6);
and AND3 (N240, N238, N138, N105);
or OR3 (N241, N235, N23, N13);
nor NOR3 (N242, N240, N192, N232);
xor XOR2 (N243, N236, N237);
xor XOR2 (N244, N35, N30);
and AND4 (N245, N228, N132, N141, N10);
and AND4 (N246, N245, N20, N226, N69);
nand NAND4 (N247, N221, N228, N234, N139);
or OR2 (N248, N85, N169);
xor XOR2 (N249, N242, N247);
nand NAND3 (N250, N155, N31, N79);
not NOT1 (N251, N246);
xor XOR2 (N252, N250, N178);
buf BUF1 (N253, N241);
buf BUF1 (N254, N249);
xor XOR2 (N255, N222, N221);
or OR2 (N256, N239, N49);
nor NOR3 (N257, N248, N235, N221);
nand NAND3 (N258, N243, N40, N64);
nor NOR3 (N259, N244, N202, N112);
not NOT1 (N260, N255);
or OR2 (N261, N256, N150);
nand NAND2 (N262, N252, N162);
nor NOR3 (N263, N262, N120, N112);
buf BUF1 (N264, N261);
xor XOR2 (N265, N263, N124);
xor XOR2 (N266, N231, N66);
or OR2 (N267, N264, N19);
xor XOR2 (N268, N266, N179);
nor NOR2 (N269, N251, N73);
nand NAND4 (N270, N269, N60, N123, N149);
nor NOR3 (N271, N254, N169, N240);
not NOT1 (N272, N271);
buf BUF1 (N273, N267);
not NOT1 (N274, N259);
buf BUF1 (N275, N258);
not NOT1 (N276, N257);
xor XOR2 (N277, N270, N8);
not NOT1 (N278, N277);
and AND3 (N279, N260, N256, N261);
xor XOR2 (N280, N253, N101);
buf BUF1 (N281, N278);
and AND4 (N282, N268, N242, N53, N132);
nand NAND2 (N283, N282, N145);
nor NOR2 (N284, N281, N45);
buf BUF1 (N285, N284);
xor XOR2 (N286, N274, N276);
or OR4 (N287, N241, N111, N110, N2);
buf BUF1 (N288, N287);
and AND2 (N289, N286, N225);
buf BUF1 (N290, N288);
and AND4 (N291, N290, N119, N208, N162);
nand NAND3 (N292, N289, N17, N248);
nand NAND4 (N293, N291, N37, N84, N137);
xor XOR2 (N294, N292, N47);
or OR2 (N295, N294, N206);
and AND2 (N296, N283, N106);
xor XOR2 (N297, N293, N281);
buf BUF1 (N298, N273);
or OR4 (N299, N295, N108, N33, N138);
or OR4 (N300, N275, N113, N41, N136);
xor XOR2 (N301, N298, N263);
nor NOR2 (N302, N297, N252);
nor NOR2 (N303, N301, N197);
and AND4 (N304, N299, N205, N81, N105);
not NOT1 (N305, N272);
and AND3 (N306, N305, N195, N257);
xor XOR2 (N307, N304, N220);
buf BUF1 (N308, N279);
not NOT1 (N309, N303);
xor XOR2 (N310, N300, N236);
buf BUF1 (N311, N308);
xor XOR2 (N312, N310, N176);
not NOT1 (N313, N307);
nor NOR3 (N314, N285, N28, N60);
nand NAND4 (N315, N265, N119, N177, N232);
not NOT1 (N316, N306);
nand NAND4 (N317, N280, N284, N134, N119);
nor NOR2 (N318, N316, N136);
and AND4 (N319, N314, N282, N260, N206);
xor XOR2 (N320, N315, N79);
xor XOR2 (N321, N318, N162);
buf BUF1 (N322, N312);
and AND3 (N323, N302, N257, N7);
nand NAND4 (N324, N296, N63, N18, N116);
nand NAND3 (N325, N324, N194, N80);
and AND4 (N326, N309, N115, N114, N91);
xor XOR2 (N327, N323, N120);
nand NAND2 (N328, N321, N318);
xor XOR2 (N329, N317, N1);
nor NOR2 (N330, N319, N296);
not NOT1 (N331, N311);
buf BUF1 (N332, N322);
or OR3 (N333, N328, N86, N68);
or OR3 (N334, N333, N220, N71);
or OR2 (N335, N326, N291);
nand NAND4 (N336, N327, N72, N25, N119);
and AND4 (N337, N332, N263, N194, N332);
nor NOR3 (N338, N330, N288, N181);
or OR4 (N339, N313, N24, N302, N16);
and AND2 (N340, N329, N5);
not NOT1 (N341, N334);
and AND4 (N342, N338, N77, N65, N117);
nand NAND4 (N343, N331, N87, N259, N109);
nand NAND3 (N344, N325, N51, N267);
nor NOR3 (N345, N337, N160, N131);
or OR3 (N346, N345, N134, N108);
nor NOR4 (N347, N335, N344, N252, N37);
xor XOR2 (N348, N48, N53);
buf BUF1 (N349, N320);
buf BUF1 (N350, N336);
or OR2 (N351, N343, N130);
buf BUF1 (N352, N348);
nor NOR2 (N353, N350, N328);
buf BUF1 (N354, N347);
nand NAND4 (N355, N353, N116, N163, N115);
xor XOR2 (N356, N342, N89);
or OR4 (N357, N339, N9, N25, N189);
buf BUF1 (N358, N352);
xor XOR2 (N359, N341, N210);
xor XOR2 (N360, N358, N342);
xor XOR2 (N361, N346, N263);
and AND2 (N362, N349, N127);
nor NOR4 (N363, N340, N36, N55, N59);
xor XOR2 (N364, N360, N17);
buf BUF1 (N365, N364);
nand NAND2 (N366, N354, N49);
not NOT1 (N367, N363);
xor XOR2 (N368, N355, N182);
not NOT1 (N369, N365);
nand NAND4 (N370, N351, N60, N138, N260);
buf BUF1 (N371, N362);
nand NAND4 (N372, N371, N202, N341, N237);
or OR2 (N373, N366, N137);
or OR4 (N374, N372, N21, N311, N50);
nor NOR3 (N375, N367, N22, N267);
nand NAND2 (N376, N359, N315);
nand NAND2 (N377, N376, N97);
nand NAND3 (N378, N356, N176, N209);
xor XOR2 (N379, N370, N350);
nor NOR2 (N380, N374, N102);
or OR3 (N381, N373, N291, N232);
nor NOR3 (N382, N381, N56, N109);
or OR3 (N383, N380, N130, N96);
or OR3 (N384, N382, N79, N102);
nand NAND2 (N385, N383, N59);
or OR2 (N386, N384, N61);
xor XOR2 (N387, N386, N214);
or OR3 (N388, N377, N272, N214);
nand NAND2 (N389, N368, N351);
nor NOR3 (N390, N389, N346, N362);
not NOT1 (N391, N388);
buf BUF1 (N392, N361);
nand NAND2 (N393, N379, N93);
not NOT1 (N394, N390);
nand NAND3 (N395, N385, N213, N289);
and AND2 (N396, N391, N130);
xor XOR2 (N397, N394, N107);
nor NOR4 (N398, N369, N23, N316, N362);
nor NOR3 (N399, N396, N319, N346);
and AND4 (N400, N399, N45, N186, N284);
xor XOR2 (N401, N398, N359);
nor NOR2 (N402, N378, N83);
buf BUF1 (N403, N397);
nor NOR4 (N404, N392, N307, N95, N277);
buf BUF1 (N405, N395);
and AND2 (N406, N402, N20);
nor NOR4 (N407, N406, N51, N297, N76);
or OR2 (N408, N375, N112);
nand NAND4 (N409, N403, N90, N271, N143);
not NOT1 (N410, N401);
nand NAND4 (N411, N357, N285, N65, N363);
buf BUF1 (N412, N387);
and AND3 (N413, N412, N396, N340);
nand NAND2 (N414, N404, N349);
xor XOR2 (N415, N413, N308);
and AND2 (N416, N415, N240);
nor NOR2 (N417, N400, N106);
not NOT1 (N418, N407);
or OR2 (N419, N405, N142);
or OR2 (N420, N409, N43);
buf BUF1 (N421, N416);
nor NOR2 (N422, N411, N287);
nor NOR4 (N423, N417, N48, N320, N72);
or OR3 (N424, N421, N15, N163);
nand NAND3 (N425, N423, N233, N134);
or OR3 (N426, N408, N43, N359);
and AND4 (N427, N393, N107, N241, N165);
or OR3 (N428, N419, N50, N151);
not NOT1 (N429, N420);
or OR3 (N430, N426, N359, N365);
nor NOR4 (N431, N430, N301, N344, N55);
nor NOR4 (N432, N428, N266, N215, N97);
not NOT1 (N433, N414);
or OR2 (N434, N433, N165);
buf BUF1 (N435, N424);
or OR4 (N436, N425, N408, N217, N120);
or OR2 (N437, N436, N180);
and AND3 (N438, N418, N412, N315);
xor XOR2 (N439, N429, N397);
xor XOR2 (N440, N439, N315);
and AND2 (N441, N422, N306);
not NOT1 (N442, N410);
nor NOR4 (N443, N427, N354, N132, N44);
nand NAND4 (N444, N442, N16, N395, N20);
and AND2 (N445, N444, N378);
or OR4 (N446, N440, N189, N386, N420);
and AND3 (N447, N431, N50, N79);
or OR4 (N448, N446, N95, N436, N420);
and AND2 (N449, N432, N238);
xor XOR2 (N450, N441, N362);
and AND2 (N451, N447, N68);
nor NOR3 (N452, N443, N224, N201);
nand NAND2 (N453, N450, N271);
and AND4 (N454, N452, N135, N231, N239);
nand NAND3 (N455, N453, N37, N264);
buf BUF1 (N456, N438);
not NOT1 (N457, N454);
nand NAND2 (N458, N449, N327);
not NOT1 (N459, N434);
nor NOR2 (N460, N456, N433);
xor XOR2 (N461, N458, N232);
xor XOR2 (N462, N459, N36);
nand NAND3 (N463, N455, N215, N192);
and AND4 (N464, N463, N221, N418, N355);
xor XOR2 (N465, N437, N334);
xor XOR2 (N466, N435, N82);
nor NOR4 (N467, N460, N244, N129, N180);
or OR2 (N468, N465, N279);
nor NOR2 (N469, N445, N65);
buf BUF1 (N470, N468);
or OR4 (N471, N462, N145, N401, N452);
xor XOR2 (N472, N448, N379);
not NOT1 (N473, N461);
xor XOR2 (N474, N471, N395);
nor NOR4 (N475, N466, N195, N318, N199);
xor XOR2 (N476, N470, N177);
or OR2 (N477, N475, N336);
nand NAND3 (N478, N457, N336, N262);
nor NOR2 (N479, N477, N9);
and AND4 (N480, N451, N392, N373, N18);
not NOT1 (N481, N480);
nor NOR3 (N482, N478, N127, N157);
nor NOR3 (N483, N474, N477, N233);
nor NOR2 (N484, N469, N236);
and AND4 (N485, N467, N386, N460, N265);
or OR3 (N486, N479, N438, N377);
not NOT1 (N487, N476);
not NOT1 (N488, N485);
not NOT1 (N489, N484);
nand NAND4 (N490, N483, N482, N346, N130);
buf BUF1 (N491, N444);
or OR3 (N492, N486, N30, N455);
xor XOR2 (N493, N492, N98);
nor NOR4 (N494, N481, N286, N234, N484);
or OR4 (N495, N473, N458, N362, N350);
xor XOR2 (N496, N488, N94);
buf BUF1 (N497, N472);
buf BUF1 (N498, N495);
nor NOR2 (N499, N497, N42);
not NOT1 (N500, N491);
nor NOR2 (N501, N493, N271);
nor NOR4 (N502, N487, N463, N181, N86);
nand NAND4 (N503, N464, N337, N210, N385);
not NOT1 (N504, N496);
xor XOR2 (N505, N500, N4);
xor XOR2 (N506, N499, N131);
or OR2 (N507, N489, N340);
not NOT1 (N508, N507);
buf BUF1 (N509, N505);
nand NAND4 (N510, N494, N69, N65, N202);
xor XOR2 (N511, N501, N75);
and AND2 (N512, N509, N258);
buf BUF1 (N513, N503);
and AND2 (N514, N512, N423);
xor XOR2 (N515, N502, N273);
buf BUF1 (N516, N515);
or OR2 (N517, N513, N64);
xor XOR2 (N518, N498, N42);
buf BUF1 (N519, N514);
nand NAND2 (N520, N511, N423);
and AND2 (N521, N506, N421);
nand NAND2 (N522, N510, N471);
or OR3 (N523, N516, N449, N333);
not NOT1 (N524, N517);
or OR4 (N525, N508, N207, N8, N289);
or OR4 (N526, N520, N143, N199, N240);
xor XOR2 (N527, N521, N38);
nor NOR4 (N528, N504, N441, N414, N359);
nor NOR4 (N529, N519, N247, N176, N149);
buf BUF1 (N530, N528);
not NOT1 (N531, N526);
buf BUF1 (N532, N524);
nand NAND4 (N533, N523, N164, N122, N360);
nor NOR2 (N534, N527, N27);
buf BUF1 (N535, N530);
not NOT1 (N536, N532);
xor XOR2 (N537, N525, N96);
nand NAND3 (N538, N537, N376, N39);
xor XOR2 (N539, N490, N335);
nand NAND4 (N540, N531, N422, N404, N145);
or OR3 (N541, N538, N11, N306);
nor NOR4 (N542, N518, N302, N484, N254);
or OR3 (N543, N539, N173, N532);
nor NOR3 (N544, N540, N243, N411);
nor NOR4 (N545, N534, N312, N320, N535);
nor NOR3 (N546, N104, N330, N353);
nor NOR2 (N547, N533, N10);
buf BUF1 (N548, N544);
buf BUF1 (N549, N545);
xor XOR2 (N550, N536, N252);
or OR3 (N551, N522, N54, N197);
nand NAND2 (N552, N546, N499);
nor NOR3 (N553, N550, N374, N200);
nor NOR3 (N554, N548, N538, N384);
nand NAND4 (N555, N549, N549, N251, N431);
xor XOR2 (N556, N554, N42);
buf BUF1 (N557, N542);
buf BUF1 (N558, N557);
nand NAND4 (N559, N555, N388, N299, N317);
and AND4 (N560, N529, N443, N21, N195);
xor XOR2 (N561, N543, N295);
xor XOR2 (N562, N556, N241);
nand NAND4 (N563, N562, N139, N430, N137);
nand NAND2 (N564, N552, N521);
buf BUF1 (N565, N541);
xor XOR2 (N566, N559, N432);
and AND4 (N567, N564, N9, N243, N540);
xor XOR2 (N568, N567, N441);
and AND2 (N569, N563, N419);
not NOT1 (N570, N569);
xor XOR2 (N571, N558, N292);
buf BUF1 (N572, N570);
not NOT1 (N573, N551);
nand NAND2 (N574, N573, N530);
nand NAND3 (N575, N566, N400, N329);
nand NAND3 (N576, N560, N241, N144);
buf BUF1 (N577, N561);
xor XOR2 (N578, N577, N462);
nor NOR4 (N579, N572, N286, N319, N550);
xor XOR2 (N580, N568, N185);
or OR2 (N581, N553, N450);
or OR3 (N582, N574, N434, N361);
or OR4 (N583, N582, N382, N381, N113);
or OR2 (N584, N575, N294);
not NOT1 (N585, N571);
xor XOR2 (N586, N576, N545);
or OR4 (N587, N583, N152, N342, N483);
xor XOR2 (N588, N587, N528);
nand NAND2 (N589, N588, N452);
not NOT1 (N590, N589);
nor NOR3 (N591, N585, N99, N190);
not NOT1 (N592, N590);
buf BUF1 (N593, N579);
nand NAND3 (N594, N593, N289, N15);
nand NAND4 (N595, N584, N115, N496, N446);
xor XOR2 (N596, N547, N316);
or OR4 (N597, N596, N228, N102, N48);
nand NAND4 (N598, N591, N264, N254, N23);
not NOT1 (N599, N565);
or OR2 (N600, N581, N593);
buf BUF1 (N601, N595);
buf BUF1 (N602, N599);
xor XOR2 (N603, N601, N23);
and AND4 (N604, N594, N82, N326, N91);
and AND2 (N605, N586, N487);
or OR3 (N606, N578, N446, N539);
nand NAND2 (N607, N605, N48);
nor NOR2 (N608, N602, N210);
nor NOR4 (N609, N597, N572, N475, N133);
nand NAND4 (N610, N607, N534, N128, N120);
nor NOR3 (N611, N608, N57, N323);
nor NOR2 (N612, N604, N220);
or OR2 (N613, N600, N391);
buf BUF1 (N614, N580);
xor XOR2 (N615, N598, N419);
nor NOR4 (N616, N611, N580, N174, N347);
nor NOR4 (N617, N610, N175, N42, N419);
nor NOR3 (N618, N614, N476, N365);
or OR4 (N619, N603, N488, N600, N309);
nor NOR3 (N620, N613, N557, N224);
nor NOR4 (N621, N617, N564, N311, N143);
nand NAND2 (N622, N619, N307);
not NOT1 (N623, N621);
nor NOR4 (N624, N618, N569, N417, N452);
not NOT1 (N625, N609);
and AND3 (N626, N606, N224, N210);
nand NAND3 (N627, N625, N495, N153);
nor NOR4 (N628, N592, N48, N335, N451);
buf BUF1 (N629, N626);
or OR3 (N630, N629, N12, N549);
buf BUF1 (N631, N628);
not NOT1 (N632, N631);
or OR4 (N633, N630, N395, N224, N515);
nand NAND4 (N634, N620, N180, N482, N601);
buf BUF1 (N635, N627);
buf BUF1 (N636, N623);
nor NOR3 (N637, N636, N300, N517);
not NOT1 (N638, N616);
xor XOR2 (N639, N622, N397);
or OR2 (N640, N624, N58);
nand NAND2 (N641, N637, N218);
buf BUF1 (N642, N638);
buf BUF1 (N643, N641);
buf BUF1 (N644, N642);
or OR4 (N645, N612, N233, N322, N279);
or OR3 (N646, N643, N180, N7);
buf BUF1 (N647, N640);
buf BUF1 (N648, N647);
and AND4 (N649, N639, N56, N530, N201);
not NOT1 (N650, N615);
buf BUF1 (N651, N650);
and AND3 (N652, N632, N435, N15);
or OR2 (N653, N646, N166);
xor XOR2 (N654, N652, N314);
xor XOR2 (N655, N653, N466);
nand NAND2 (N656, N655, N96);
xor XOR2 (N657, N648, N411);
or OR4 (N658, N633, N227, N510, N22);
xor XOR2 (N659, N635, N66);
buf BUF1 (N660, N651);
nor NOR2 (N661, N634, N394);
xor XOR2 (N662, N649, N37);
not NOT1 (N663, N658);
nand NAND4 (N664, N662, N302, N496, N549);
buf BUF1 (N665, N656);
or OR4 (N666, N654, N176, N523, N655);
buf BUF1 (N667, N665);
nor NOR2 (N668, N660, N637);
xor XOR2 (N669, N645, N97);
or OR3 (N670, N657, N65, N360);
nand NAND4 (N671, N668, N583, N144, N326);
buf BUF1 (N672, N671);
and AND4 (N673, N644, N624, N108, N407);
nor NOR3 (N674, N661, N566, N31);
or OR4 (N675, N674, N332, N24, N100);
xor XOR2 (N676, N675, N105);
buf BUF1 (N677, N669);
nor NOR3 (N678, N666, N316, N370);
nor NOR3 (N679, N670, N67, N100);
not NOT1 (N680, N663);
xor XOR2 (N681, N680, N343);
and AND4 (N682, N659, N48, N146, N519);
xor XOR2 (N683, N667, N524);
buf BUF1 (N684, N672);
nand NAND2 (N685, N682, N65);
not NOT1 (N686, N684);
not NOT1 (N687, N679);
buf BUF1 (N688, N683);
or OR4 (N689, N676, N549, N306, N42);
xor XOR2 (N690, N673, N90);
buf BUF1 (N691, N687);
nor NOR2 (N692, N691, N428);
or OR2 (N693, N677, N435);
xor XOR2 (N694, N686, N232);
or OR2 (N695, N681, N234);
and AND2 (N696, N690, N236);
xor XOR2 (N697, N695, N632);
xor XOR2 (N698, N678, N118);
nand NAND2 (N699, N696, N520);
buf BUF1 (N700, N664);
nor NOR3 (N701, N689, N523, N336);
and AND2 (N702, N685, N177);
nor NOR2 (N703, N688, N574);
or OR4 (N704, N698, N523, N668, N266);
not NOT1 (N705, N697);
nand NAND4 (N706, N705, N105, N24, N230);
nor NOR2 (N707, N693, N397);
nand NAND3 (N708, N692, N527, N598);
nand NAND2 (N709, N707, N664);
xor XOR2 (N710, N699, N681);
nor NOR2 (N711, N701, N167);
or OR3 (N712, N711, N540, N195);
and AND4 (N713, N694, N97, N101, N3);
buf BUF1 (N714, N709);
xor XOR2 (N715, N713, N347);
buf BUF1 (N716, N703);
not NOT1 (N717, N712);
nand NAND3 (N718, N716, N558, N25);
and AND3 (N719, N702, N77, N681);
and AND3 (N720, N710, N204, N314);
and AND4 (N721, N717, N626, N313, N35);
nand NAND4 (N722, N706, N583, N380, N602);
or OR2 (N723, N720, N273);
nor NOR3 (N724, N723, N402, N289);
nor NOR4 (N725, N704, N381, N573, N658);
nor NOR4 (N726, N715, N246, N92, N103);
nor NOR3 (N727, N724, N436, N242);
xor XOR2 (N728, N708, N348);
nor NOR3 (N729, N718, N13, N257);
buf BUF1 (N730, N721);
not NOT1 (N731, N722);
xor XOR2 (N732, N719, N707);
and AND2 (N733, N732, N343);
and AND2 (N734, N725, N203);
nor NOR2 (N735, N733, N561);
xor XOR2 (N736, N734, N574);
not NOT1 (N737, N728);
not NOT1 (N738, N700);
nor NOR2 (N739, N714, N378);
not NOT1 (N740, N737);
nand NAND4 (N741, N736, N437, N711, N68);
xor XOR2 (N742, N730, N574);
not NOT1 (N743, N742);
and AND4 (N744, N740, N70, N302, N519);
xor XOR2 (N745, N739, N565);
or OR2 (N746, N731, N123);
xor XOR2 (N747, N746, N505);
and AND4 (N748, N745, N453, N667, N670);
nor NOR3 (N749, N747, N148, N748);
xor XOR2 (N750, N656, N455);
xor XOR2 (N751, N743, N291);
not NOT1 (N752, N750);
and AND4 (N753, N752, N572, N408, N323);
buf BUF1 (N754, N744);
not NOT1 (N755, N738);
and AND2 (N756, N729, N381);
not NOT1 (N757, N754);
buf BUF1 (N758, N741);
xor XOR2 (N759, N758, N719);
or OR4 (N760, N757, N24, N494, N119);
xor XOR2 (N761, N756, N674);
not NOT1 (N762, N759);
nand NAND4 (N763, N755, N227, N492, N348);
nor NOR3 (N764, N727, N204, N156);
not NOT1 (N765, N760);
buf BUF1 (N766, N765);
xor XOR2 (N767, N726, N288);
not NOT1 (N768, N749);
and AND3 (N769, N761, N44, N48);
nor NOR2 (N770, N753, N266);
not NOT1 (N771, N735);
nor NOR2 (N772, N768, N707);
buf BUF1 (N773, N771);
or OR2 (N774, N770, N480);
nand NAND2 (N775, N772, N30);
buf BUF1 (N776, N775);
buf BUF1 (N777, N773);
or OR2 (N778, N763, N314);
or OR2 (N779, N777, N746);
buf BUF1 (N780, N779);
or OR3 (N781, N769, N526, N687);
buf BUF1 (N782, N778);
buf BUF1 (N783, N767);
nor NOR2 (N784, N762, N104);
nand NAND2 (N785, N783, N720);
and AND4 (N786, N780, N189, N202, N261);
nand NAND4 (N787, N766, N721, N581, N551);
buf BUF1 (N788, N751);
xor XOR2 (N789, N776, N715);
or OR3 (N790, N786, N45, N319);
nand NAND4 (N791, N788, N687, N233, N723);
not NOT1 (N792, N791);
buf BUF1 (N793, N764);
not NOT1 (N794, N785);
or OR3 (N795, N774, N560, N724);
xor XOR2 (N796, N795, N301);
xor XOR2 (N797, N790, N149);
not NOT1 (N798, N793);
nand NAND2 (N799, N796, N21);
or OR2 (N800, N799, N391);
nand NAND3 (N801, N792, N139, N372);
or OR4 (N802, N797, N613, N273, N598);
not NOT1 (N803, N802);
nor NOR3 (N804, N798, N438, N365);
not NOT1 (N805, N781);
and AND2 (N806, N787, N723);
or OR2 (N807, N801, N757);
or OR4 (N808, N789, N631, N305, N442);
nand NAND4 (N809, N807, N709, N697, N225);
xor XOR2 (N810, N808, N571);
and AND2 (N811, N805, N71);
nand NAND4 (N812, N810, N337, N332, N587);
endmodule