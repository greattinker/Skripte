// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N323,N318,N312,N321,N305,N320,N310,N322,N315,N324;

not NOT1 (N25, N17);
buf BUF1 (N26, N25);
or OR2 (N27, N12, N22);
xor XOR2 (N28, N22, N1);
and AND2 (N29, N11, N25);
or OR4 (N30, N10, N3, N5, N29);
buf BUF1 (N31, N10);
not NOT1 (N32, N10);
nor NOR4 (N33, N12, N19, N13, N31);
nor NOR4 (N34, N3, N8, N17, N32);
or OR3 (N35, N33, N21, N4);
buf BUF1 (N36, N12);
and AND4 (N37, N23, N11, N17, N34);
nand NAND3 (N38, N31, N13, N20);
buf BUF1 (N39, N23);
not NOT1 (N40, N3);
nand NAND3 (N41, N39, N31, N28);
and AND4 (N42, N21, N19, N6, N12);
nand NAND2 (N43, N38, N1);
nand NAND2 (N44, N27, N4);
nand NAND3 (N45, N30, N17, N29);
not NOT1 (N46, N40);
nor NOR4 (N47, N37, N15, N22, N8);
and AND4 (N48, N26, N5, N47, N30);
or OR2 (N49, N8, N35);
buf BUF1 (N50, N28);
xor XOR2 (N51, N41, N46);
buf BUF1 (N52, N51);
xor XOR2 (N53, N50, N15);
not NOT1 (N54, N15);
not NOT1 (N55, N43);
buf BUF1 (N56, N45);
and AND2 (N57, N53, N24);
xor XOR2 (N58, N48, N35);
nor NOR4 (N59, N58, N3, N31, N19);
or OR4 (N60, N52, N22, N58, N32);
not NOT1 (N61, N44);
and AND4 (N62, N61, N50, N38, N55);
and AND2 (N63, N10, N52);
buf BUF1 (N64, N57);
and AND2 (N65, N59, N41);
not NOT1 (N66, N62);
nor NOR4 (N67, N42, N12, N1, N12);
nor NOR2 (N68, N60, N49);
not NOT1 (N69, N32);
xor XOR2 (N70, N36, N5);
xor XOR2 (N71, N68, N63);
xor XOR2 (N72, N51, N61);
buf BUF1 (N73, N72);
buf BUF1 (N74, N69);
or OR4 (N75, N66, N10, N65, N5);
nor NOR4 (N76, N22, N47, N72, N38);
not NOT1 (N77, N74);
buf BUF1 (N78, N77);
or OR3 (N79, N73, N65, N51);
and AND3 (N80, N64, N72, N55);
not NOT1 (N81, N67);
not NOT1 (N82, N56);
xor XOR2 (N83, N75, N82);
xor XOR2 (N84, N10, N82);
nor NOR3 (N85, N78, N46, N55);
or OR3 (N86, N80, N77, N65);
or OR4 (N87, N86, N53, N17, N33);
and AND4 (N88, N83, N51, N72, N28);
xor XOR2 (N89, N70, N53);
buf BUF1 (N90, N71);
nand NAND4 (N91, N81, N40, N71, N4);
or OR4 (N92, N76, N11, N33, N50);
or OR4 (N93, N84, N33, N8, N31);
nor NOR2 (N94, N93, N34);
nand NAND2 (N95, N90, N69);
xor XOR2 (N96, N91, N40);
xor XOR2 (N97, N94, N38);
and AND3 (N98, N89, N89, N79);
xor XOR2 (N99, N98, N30);
and AND2 (N100, N86, N46);
xor XOR2 (N101, N85, N85);
xor XOR2 (N102, N96, N64);
xor XOR2 (N103, N97, N55);
buf BUF1 (N104, N102);
xor XOR2 (N105, N101, N71);
xor XOR2 (N106, N87, N76);
nand NAND2 (N107, N103, N54);
nor NOR3 (N108, N95, N75, N25);
not NOT1 (N109, N78);
buf BUF1 (N110, N92);
and AND3 (N111, N106, N75, N86);
nand NAND3 (N112, N109, N51, N83);
xor XOR2 (N113, N112, N13);
nor NOR2 (N114, N104, N18);
buf BUF1 (N115, N88);
nand NAND4 (N116, N111, N83, N67, N23);
not NOT1 (N117, N110);
xor XOR2 (N118, N113, N17);
and AND4 (N119, N99, N57, N21, N30);
nand NAND2 (N120, N117, N59);
and AND2 (N121, N120, N59);
and AND4 (N122, N114, N120, N58, N15);
or OR2 (N123, N118, N57);
nand NAND3 (N124, N122, N26, N58);
nor NOR4 (N125, N107, N40, N28, N114);
and AND4 (N126, N123, N89, N34, N95);
nor NOR3 (N127, N125, N16, N64);
and AND2 (N128, N119, N116);
nor NOR3 (N129, N87, N87, N51);
buf BUF1 (N130, N121);
not NOT1 (N131, N108);
or OR4 (N132, N131, N79, N88, N59);
buf BUF1 (N133, N132);
nand NAND2 (N134, N129, N57);
nand NAND4 (N135, N133, N77, N23, N15);
and AND2 (N136, N126, N13);
and AND4 (N137, N134, N104, N46, N28);
buf BUF1 (N138, N115);
xor XOR2 (N139, N135, N90);
not NOT1 (N140, N127);
or OR3 (N141, N105, N8, N26);
nand NAND4 (N142, N100, N1, N82, N99);
xor XOR2 (N143, N140, N57);
nor NOR2 (N144, N130, N104);
xor XOR2 (N145, N139, N4);
nand NAND2 (N146, N143, N52);
xor XOR2 (N147, N124, N126);
not NOT1 (N148, N138);
or OR3 (N149, N144, N41, N135);
nor NOR4 (N150, N141, N118, N61, N83);
nor NOR4 (N151, N128, N103, N90, N53);
nand NAND3 (N152, N146, N87, N60);
xor XOR2 (N153, N145, N135);
nor NOR3 (N154, N150, N81, N94);
buf BUF1 (N155, N142);
xor XOR2 (N156, N137, N28);
and AND3 (N157, N156, N143, N53);
nor NOR3 (N158, N149, N154, N107);
or OR4 (N159, N105, N120, N48, N21);
or OR4 (N160, N153, N110, N44, N148);
nand NAND3 (N161, N103, N154, N20);
not NOT1 (N162, N151);
not NOT1 (N163, N136);
and AND3 (N164, N161, N143, N136);
nand NAND2 (N165, N163, N154);
or OR3 (N166, N147, N50, N92);
buf BUF1 (N167, N162);
not NOT1 (N168, N159);
not NOT1 (N169, N160);
nor NOR3 (N170, N168, N127, N51);
buf BUF1 (N171, N170);
nand NAND3 (N172, N169, N106, N119);
buf BUF1 (N173, N166);
xor XOR2 (N174, N172, N41);
or OR3 (N175, N164, N110, N136);
nor NOR2 (N176, N174, N12);
and AND3 (N177, N158, N111, N175);
or OR4 (N178, N14, N136, N94, N149);
not NOT1 (N179, N167);
buf BUF1 (N180, N177);
buf BUF1 (N181, N173);
buf BUF1 (N182, N178);
nor NOR4 (N183, N165, N44, N66, N39);
nor NOR2 (N184, N152, N165);
or OR2 (N185, N182, N116);
nor NOR3 (N186, N155, N2, N105);
and AND4 (N187, N176, N38, N181, N24);
or OR2 (N188, N8, N73);
nand NAND4 (N189, N157, N145, N118, N2);
nor NOR4 (N190, N179, N38, N124, N182);
or OR4 (N191, N186, N105, N148, N4);
nor NOR2 (N192, N184, N159);
or OR3 (N193, N183, N126, N52);
or OR2 (N194, N185, N65);
buf BUF1 (N195, N171);
and AND4 (N196, N188, N39, N2, N21);
xor XOR2 (N197, N180, N144);
nor NOR4 (N198, N193, N57, N118, N120);
nor NOR2 (N199, N198, N11);
buf BUF1 (N200, N190);
or OR3 (N201, N199, N53, N62);
nor NOR3 (N202, N195, N17, N15);
or OR3 (N203, N201, N99, N187);
and AND2 (N204, N20, N44);
and AND2 (N205, N196, N165);
or OR2 (N206, N197, N16);
xor XOR2 (N207, N194, N178);
or OR2 (N208, N204, N64);
xor XOR2 (N209, N202, N40);
nor NOR2 (N210, N189, N82);
nor NOR2 (N211, N192, N23);
or OR4 (N212, N207, N105, N155, N72);
nor NOR4 (N213, N211, N159, N125, N207);
or OR3 (N214, N200, N17, N43);
or OR4 (N215, N205, N185, N194, N125);
nand NAND4 (N216, N191, N70, N155, N13);
and AND2 (N217, N213, N147);
buf BUF1 (N218, N206);
and AND2 (N219, N210, N214);
not NOT1 (N220, N196);
and AND4 (N221, N219, N136, N33, N162);
nor NOR2 (N222, N209, N16);
not NOT1 (N223, N216);
xor XOR2 (N224, N223, N183);
nand NAND4 (N225, N208, N72, N99, N60);
nor NOR3 (N226, N220, N73, N161);
buf BUF1 (N227, N226);
buf BUF1 (N228, N224);
buf BUF1 (N229, N203);
nand NAND2 (N230, N222, N74);
nand NAND3 (N231, N228, N114, N205);
nand NAND2 (N232, N215, N66);
nand NAND3 (N233, N218, N223, N102);
buf BUF1 (N234, N217);
nor NOR3 (N235, N230, N22, N13);
xor XOR2 (N236, N234, N144);
nor NOR2 (N237, N231, N224);
not NOT1 (N238, N229);
not NOT1 (N239, N212);
not NOT1 (N240, N227);
nand NAND4 (N241, N235, N113, N5, N202);
not NOT1 (N242, N221);
nor NOR4 (N243, N240, N232, N1, N78);
buf BUF1 (N244, N203);
buf BUF1 (N245, N242);
nor NOR2 (N246, N236, N206);
buf BUF1 (N247, N237);
and AND3 (N248, N233, N224, N29);
not NOT1 (N249, N246);
buf BUF1 (N250, N239);
xor XOR2 (N251, N241, N160);
or OR3 (N252, N247, N160, N208);
xor XOR2 (N253, N243, N132);
nor NOR2 (N254, N249, N175);
not NOT1 (N255, N248);
nand NAND2 (N256, N252, N107);
nor NOR2 (N257, N245, N131);
nor NOR4 (N258, N255, N247, N237, N256);
not NOT1 (N259, N106);
buf BUF1 (N260, N257);
nor NOR2 (N261, N253, N10);
nand NAND2 (N262, N259, N142);
buf BUF1 (N263, N260);
nand NAND4 (N264, N254, N73, N200, N58);
and AND2 (N265, N238, N132);
buf BUF1 (N266, N265);
or OR3 (N267, N258, N155, N7);
nor NOR2 (N268, N267, N109);
and AND2 (N269, N264, N65);
not NOT1 (N270, N250);
buf BUF1 (N271, N251);
nand NAND3 (N272, N244, N68, N71);
buf BUF1 (N273, N272);
nor NOR3 (N274, N269, N60, N36);
or OR3 (N275, N266, N99, N79);
not NOT1 (N276, N271);
not NOT1 (N277, N274);
and AND2 (N278, N273, N86);
not NOT1 (N279, N262);
xor XOR2 (N280, N276, N48);
nor NOR3 (N281, N263, N58, N144);
nor NOR2 (N282, N277, N62);
xor XOR2 (N283, N278, N155);
or OR3 (N284, N283, N259, N173);
or OR2 (N285, N268, N149);
xor XOR2 (N286, N270, N158);
not NOT1 (N287, N225);
buf BUF1 (N288, N279);
or OR2 (N289, N275, N166);
or OR4 (N290, N282, N181, N258, N284);
nand NAND2 (N291, N130, N278);
and AND3 (N292, N281, N281, N180);
not NOT1 (N293, N289);
buf BUF1 (N294, N285);
nor NOR3 (N295, N286, N144, N28);
or OR4 (N296, N291, N166, N206, N51);
buf BUF1 (N297, N295);
xor XOR2 (N298, N294, N71);
or OR4 (N299, N297, N126, N290, N49);
nor NOR2 (N300, N60, N82);
not NOT1 (N301, N299);
nand NAND4 (N302, N292, N172, N170, N219);
and AND3 (N303, N293, N170, N109);
xor XOR2 (N304, N298, N166);
not NOT1 (N305, N296);
not NOT1 (N306, N302);
nor NOR2 (N307, N261, N161);
xor XOR2 (N308, N304, N6);
and AND3 (N309, N301, N131, N106);
or OR3 (N310, N308, N195, N88);
buf BUF1 (N311, N306);
nor NOR3 (N312, N280, N266, N16);
xor XOR2 (N313, N300, N158);
buf BUF1 (N314, N303);
or OR3 (N315, N313, N314, N63);
nand NAND3 (N316, N192, N182, N89);
nor NOR3 (N317, N307, N216, N39);
not NOT1 (N318, N288);
or OR4 (N319, N311, N131, N25, N63);
not NOT1 (N320, N316);
or OR2 (N321, N317, N117);
or OR2 (N322, N287, N51);
or OR4 (N323, N319, N21, N146, N249);
xor XOR2 (N324, N309, N210);
endmodule