// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N313,N319,N311,N321,N302,N318,N316,N286,N317,N322;

and AND3 (N23, N18, N15, N3);
buf BUF1 (N24, N1);
or OR4 (N25, N6, N15, N22, N16);
nor NOR3 (N26, N12, N4, N11);
buf BUF1 (N27, N12);
and AND4 (N28, N9, N19, N6, N5);
and AND4 (N29, N25, N20, N1, N10);
nor NOR4 (N30, N23, N24, N17, N24);
buf BUF1 (N31, N5);
buf BUF1 (N32, N26);
buf BUF1 (N33, N8);
xor XOR2 (N34, N7, N9);
nand NAND4 (N35, N22, N18, N18, N9);
nand NAND3 (N36, N35, N2, N12);
not NOT1 (N37, N23);
xor XOR2 (N38, N33, N18);
not NOT1 (N39, N37);
and AND3 (N40, N34, N33, N17);
xor XOR2 (N41, N27, N8);
or OR4 (N42, N40, N29, N34, N7);
nand NAND3 (N43, N33, N17, N19);
and AND3 (N44, N36, N29, N22);
nand NAND2 (N45, N41, N5);
nand NAND2 (N46, N28, N16);
and AND2 (N47, N30, N36);
or OR3 (N48, N47, N46, N6);
xor XOR2 (N49, N35, N30);
and AND2 (N50, N48, N37);
nor NOR3 (N51, N42, N26, N41);
nor NOR2 (N52, N31, N15);
buf BUF1 (N53, N45);
not NOT1 (N54, N44);
xor XOR2 (N55, N50, N16);
buf BUF1 (N56, N54);
or OR4 (N57, N38, N6, N24, N1);
not NOT1 (N58, N55);
or OR4 (N59, N58, N57, N29, N19);
not NOT1 (N60, N34);
xor XOR2 (N61, N59, N57);
and AND3 (N62, N32, N43, N16);
and AND4 (N63, N3, N17, N14, N50);
not NOT1 (N64, N60);
and AND4 (N65, N63, N35, N20, N50);
buf BUF1 (N66, N51);
not NOT1 (N67, N49);
nand NAND2 (N68, N53, N56);
nor NOR3 (N69, N54, N53, N32);
nand NAND2 (N70, N64, N5);
buf BUF1 (N71, N65);
buf BUF1 (N72, N62);
buf BUF1 (N73, N39);
or OR2 (N74, N52, N7);
buf BUF1 (N75, N74);
not NOT1 (N76, N69);
and AND3 (N77, N73, N18, N39);
nor NOR4 (N78, N77, N11, N59, N12);
nor NOR3 (N79, N67, N52, N69);
and AND4 (N80, N72, N78, N68, N5);
not NOT1 (N81, N1);
or OR4 (N82, N20, N26, N40, N42);
xor XOR2 (N83, N81, N77);
nand NAND3 (N84, N61, N9, N26);
nand NAND3 (N85, N75, N6, N79);
nand NAND3 (N86, N10, N10, N76);
and AND4 (N87, N65, N62, N46, N33);
not NOT1 (N88, N85);
buf BUF1 (N89, N80);
not NOT1 (N90, N88);
xor XOR2 (N91, N90, N42);
nor NOR2 (N92, N82, N58);
buf BUF1 (N93, N70);
buf BUF1 (N94, N86);
not NOT1 (N95, N92);
or OR3 (N96, N83, N2, N26);
nand NAND2 (N97, N66, N12);
nor NOR3 (N98, N94, N81, N35);
nor NOR3 (N99, N71, N50, N74);
buf BUF1 (N100, N97);
and AND3 (N101, N91, N12, N25);
xor XOR2 (N102, N99, N45);
and AND2 (N103, N89, N57);
buf BUF1 (N104, N98);
buf BUF1 (N105, N95);
nor NOR4 (N106, N96, N85, N59, N7);
and AND2 (N107, N100, N75);
and AND3 (N108, N84, N42, N24);
nand NAND3 (N109, N107, N22, N14);
or OR3 (N110, N109, N1, N82);
and AND3 (N111, N108, N1, N57);
and AND4 (N112, N87, N60, N93, N83);
nor NOR2 (N113, N80, N46);
xor XOR2 (N114, N111, N9);
nand NAND2 (N115, N106, N9);
nand NAND3 (N116, N114, N56, N105);
not NOT1 (N117, N26);
nand NAND2 (N118, N115, N74);
xor XOR2 (N119, N117, N3);
nor NOR4 (N120, N110, N67, N103, N81);
nand NAND3 (N121, N31, N5, N36);
and AND2 (N122, N102, N3);
not NOT1 (N123, N116);
nand NAND2 (N124, N122, N22);
not NOT1 (N125, N113);
nor NOR3 (N126, N120, N70, N70);
not NOT1 (N127, N112);
nor NOR3 (N128, N123, N60, N2);
and AND3 (N129, N104, N126, N122);
xor XOR2 (N130, N42, N71);
and AND2 (N131, N101, N62);
and AND2 (N132, N129, N44);
nand NAND2 (N133, N132, N88);
or OR4 (N134, N119, N107, N11, N57);
and AND3 (N135, N130, N107, N7);
or OR4 (N136, N127, N49, N22, N132);
and AND3 (N137, N121, N38, N107);
and AND3 (N138, N128, N27, N130);
or OR3 (N139, N133, N125, N134);
nand NAND4 (N140, N104, N27, N84, N137);
not NOT1 (N141, N110);
nor NOR4 (N142, N4, N108, N53, N37);
nor NOR3 (N143, N141, N10, N24);
xor XOR2 (N144, N140, N43);
nor NOR4 (N145, N143, N7, N71, N136);
buf BUF1 (N146, N109);
nor NOR4 (N147, N124, N117, N17, N95);
not NOT1 (N148, N146);
nand NAND2 (N149, N148, N109);
and AND3 (N150, N144, N141, N30);
and AND3 (N151, N145, N43, N11);
xor XOR2 (N152, N150, N34);
nand NAND3 (N153, N142, N131, N8);
nor NOR2 (N154, N64, N144);
xor XOR2 (N155, N154, N99);
nor NOR2 (N156, N139, N113);
and AND2 (N157, N147, N78);
not NOT1 (N158, N156);
not NOT1 (N159, N118);
nor NOR3 (N160, N153, N2, N11);
xor XOR2 (N161, N151, N139);
xor XOR2 (N162, N161, N142);
nor NOR2 (N163, N149, N108);
nand NAND4 (N164, N159, N66, N68, N40);
nor NOR2 (N165, N162, N13);
and AND2 (N166, N157, N115);
and AND4 (N167, N138, N38, N74, N76);
buf BUF1 (N168, N155);
buf BUF1 (N169, N164);
or OR2 (N170, N167, N131);
or OR3 (N171, N165, N146, N53);
or OR4 (N172, N135, N26, N160, N163);
nand NAND3 (N173, N125, N129, N120);
nand NAND4 (N174, N144, N164, N118, N92);
not NOT1 (N175, N173);
xor XOR2 (N176, N170, N22);
and AND2 (N177, N166, N4);
nor NOR3 (N178, N169, N142, N115);
xor XOR2 (N179, N177, N16);
and AND3 (N180, N168, N68, N139);
nand NAND2 (N181, N175, N3);
buf BUF1 (N182, N178);
nor NOR2 (N183, N181, N76);
buf BUF1 (N184, N176);
or OR4 (N185, N152, N49, N92, N39);
buf BUF1 (N186, N184);
nor NOR3 (N187, N172, N12, N171);
nor NOR2 (N188, N102, N92);
nor NOR4 (N189, N180, N31, N36, N55);
buf BUF1 (N190, N187);
xor XOR2 (N191, N174, N11);
nor NOR4 (N192, N179, N181, N159, N172);
nand NAND2 (N193, N188, N101);
nand NAND3 (N194, N193, N61, N102);
or OR4 (N195, N189, N128, N192, N41);
or OR2 (N196, N36, N18);
and AND3 (N197, N191, N134, N103);
or OR4 (N198, N185, N126, N187, N49);
and AND2 (N199, N198, N95);
buf BUF1 (N200, N182);
nand NAND4 (N201, N200, N27, N177, N136);
not NOT1 (N202, N183);
nor NOR3 (N203, N186, N148, N58);
and AND2 (N204, N199, N47);
nor NOR4 (N205, N203, N35, N120, N131);
nor NOR2 (N206, N194, N134);
or OR2 (N207, N206, N74);
or OR4 (N208, N207, N78, N35, N95);
xor XOR2 (N209, N197, N43);
buf BUF1 (N210, N201);
or OR3 (N211, N158, N39, N100);
nand NAND4 (N212, N208, N143, N92, N63);
xor XOR2 (N213, N210, N207);
nand NAND3 (N214, N212, N59, N204);
nor NOR4 (N215, N213, N128, N71, N67);
not NOT1 (N216, N95);
and AND2 (N217, N214, N87);
and AND4 (N218, N217, N53, N159, N28);
buf BUF1 (N219, N209);
and AND4 (N220, N202, N132, N79, N190);
nor NOR3 (N221, N40, N57, N205);
nor NOR3 (N222, N132, N72, N1);
and AND2 (N223, N218, N8);
nor NOR2 (N224, N219, N193);
not NOT1 (N225, N216);
buf BUF1 (N226, N222);
or OR3 (N227, N226, N94, N159);
buf BUF1 (N228, N211);
nor NOR3 (N229, N224, N129, N7);
and AND3 (N230, N223, N95, N23);
buf BUF1 (N231, N225);
or OR3 (N232, N196, N209, N193);
not NOT1 (N233, N220);
buf BUF1 (N234, N230);
and AND3 (N235, N228, N34, N92);
and AND2 (N236, N233, N232);
nand NAND4 (N237, N235, N196, N55, N63);
or OR3 (N238, N183, N91, N182);
buf BUF1 (N239, N234);
and AND2 (N240, N238, N48);
not NOT1 (N241, N237);
xor XOR2 (N242, N236, N27);
xor XOR2 (N243, N231, N139);
nor NOR3 (N244, N242, N207, N40);
nor NOR4 (N245, N241, N13, N62, N97);
xor XOR2 (N246, N245, N64);
nor NOR4 (N247, N239, N161, N241, N164);
and AND3 (N248, N240, N209, N104);
not NOT1 (N249, N215);
nor NOR3 (N250, N243, N195, N20);
and AND3 (N251, N71, N37, N145);
nand NAND3 (N252, N229, N121, N4);
xor XOR2 (N253, N252, N232);
xor XOR2 (N254, N227, N203);
buf BUF1 (N255, N247);
xor XOR2 (N256, N221, N194);
not NOT1 (N257, N251);
buf BUF1 (N258, N256);
nand NAND3 (N259, N248, N7, N26);
not NOT1 (N260, N257);
or OR4 (N261, N259, N187, N27, N187);
xor XOR2 (N262, N244, N39);
xor XOR2 (N263, N246, N253);
buf BUF1 (N264, N243);
not NOT1 (N265, N258);
or OR2 (N266, N250, N96);
nor NOR4 (N267, N254, N196, N119, N232);
xor XOR2 (N268, N266, N55);
nand NAND2 (N269, N263, N266);
buf BUF1 (N270, N264);
or OR4 (N271, N262, N253, N16, N239);
nor NOR3 (N272, N249, N98, N83);
not NOT1 (N273, N261);
or OR3 (N274, N260, N1, N253);
nand NAND2 (N275, N274, N243);
buf BUF1 (N276, N268);
xor XOR2 (N277, N270, N215);
buf BUF1 (N278, N265);
not NOT1 (N279, N278);
nor NOR2 (N280, N273, N263);
xor XOR2 (N281, N277, N84);
not NOT1 (N282, N255);
xor XOR2 (N283, N272, N197);
or OR3 (N284, N280, N279, N154);
or OR4 (N285, N162, N244, N100, N282);
nand NAND4 (N286, N82, N76, N281, N186);
xor XOR2 (N287, N187, N283);
not NOT1 (N288, N241);
not NOT1 (N289, N267);
nand NAND4 (N290, N288, N138, N58, N183);
nor NOR3 (N291, N285, N265, N79);
not NOT1 (N292, N287);
buf BUF1 (N293, N290);
and AND2 (N294, N289, N126);
and AND3 (N295, N275, N284, N175);
and AND2 (N296, N221, N5);
nand NAND4 (N297, N269, N228, N90, N211);
buf BUF1 (N298, N296);
not NOT1 (N299, N293);
nor NOR3 (N300, N292, N277, N168);
nor NOR2 (N301, N276, N99);
nand NAND2 (N302, N271, N145);
buf BUF1 (N303, N301);
not NOT1 (N304, N300);
nor NOR4 (N305, N297, N226, N39, N229);
and AND4 (N306, N304, N130, N147, N277);
and AND2 (N307, N303, N178);
and AND3 (N308, N307, N238, N94);
nor NOR2 (N309, N291, N84);
nor NOR3 (N310, N295, N225, N245);
nand NAND2 (N311, N294, N208);
not NOT1 (N312, N309);
nor NOR3 (N313, N298, N296, N201);
not NOT1 (N314, N299);
not NOT1 (N315, N308);
and AND3 (N316, N310, N143, N5);
xor XOR2 (N317, N314, N96);
and AND2 (N318, N305, N177);
nor NOR2 (N319, N306, N207);
or OR4 (N320, N315, N52, N312, N56);
nand NAND4 (N321, N172, N1, N30, N266);
or OR2 (N322, N320, N200);
endmodule