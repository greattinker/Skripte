// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N604,N605,N613,N590,N612,N607,N602,N603,N608,N614;

nand NAND2 (N15, N7, N11);
or OR4 (N16, N7, N8, N12, N2);
nor NOR3 (N17, N8, N4, N14);
and AND4 (N18, N9, N1, N12, N17);
xor XOR2 (N19, N10, N2);
or OR4 (N20, N15, N4, N16, N17);
and AND2 (N21, N1, N17);
or OR2 (N22, N7, N10);
buf BUF1 (N23, N21);
not NOT1 (N24, N8);
not NOT1 (N25, N19);
nor NOR4 (N26, N20, N12, N25, N15);
nand NAND4 (N27, N21, N11, N10, N17);
buf BUF1 (N28, N3);
xor XOR2 (N29, N11, N9);
and AND4 (N30, N21, N23, N27, N19);
nor NOR2 (N31, N4, N5);
nor NOR3 (N32, N2, N30, N24);
not NOT1 (N33, N12);
and AND3 (N34, N3, N22, N22);
or OR2 (N35, N19, N2);
not NOT1 (N36, N6);
nor NOR4 (N37, N18, N26, N12, N1);
and AND3 (N38, N21, N31, N7);
or OR4 (N39, N28, N38, N17, N31);
buf BUF1 (N40, N10);
and AND4 (N41, N33, N12, N21, N37);
xor XOR2 (N42, N2, N36);
nor NOR4 (N43, N31, N17, N28, N21);
buf BUF1 (N44, N35);
or OR3 (N45, N39, N9, N3);
nand NAND3 (N46, N11, N18, N23);
buf BUF1 (N47, N45);
not NOT1 (N48, N46);
nand NAND3 (N49, N29, N10, N35);
xor XOR2 (N50, N32, N32);
not NOT1 (N51, N44);
or OR4 (N52, N42, N32, N43, N26);
not NOT1 (N53, N22);
xor XOR2 (N54, N47, N2);
nor NOR2 (N55, N49, N46);
buf BUF1 (N56, N48);
or OR4 (N57, N55, N31, N13, N8);
not NOT1 (N58, N57);
nand NAND4 (N59, N41, N57, N50, N4);
nor NOR2 (N60, N40, N48);
or OR4 (N61, N15, N51, N2, N39);
buf BUF1 (N62, N53);
nand NAND3 (N63, N30, N33, N23);
nor NOR2 (N64, N54, N22);
and AND2 (N65, N61, N7);
and AND3 (N66, N58, N42, N41);
nor NOR3 (N67, N52, N51, N18);
and AND2 (N68, N64, N10);
or OR2 (N69, N60, N7);
not NOT1 (N70, N34);
buf BUF1 (N71, N59);
xor XOR2 (N72, N67, N71);
not NOT1 (N73, N70);
buf BUF1 (N74, N49);
nand NAND2 (N75, N72, N39);
xor XOR2 (N76, N69, N5);
buf BUF1 (N77, N75);
buf BUF1 (N78, N76);
xor XOR2 (N79, N68, N20);
or OR4 (N80, N78, N52, N52, N49);
or OR4 (N81, N80, N1, N52, N73);
and AND3 (N82, N61, N27, N8);
and AND2 (N83, N65, N71);
not NOT1 (N84, N66);
or OR3 (N85, N62, N73, N8);
not NOT1 (N86, N84);
not NOT1 (N87, N82);
nor NOR2 (N88, N87, N46);
and AND3 (N89, N56, N23, N30);
nor NOR4 (N90, N83, N30, N2, N83);
not NOT1 (N91, N81);
nand NAND3 (N92, N88, N66, N34);
buf BUF1 (N93, N92);
not NOT1 (N94, N89);
xor XOR2 (N95, N86, N37);
and AND2 (N96, N77, N46);
not NOT1 (N97, N90);
not NOT1 (N98, N63);
buf BUF1 (N99, N96);
buf BUF1 (N100, N94);
and AND4 (N101, N97, N4, N44, N34);
or OR4 (N102, N99, N31, N31, N45);
xor XOR2 (N103, N102, N43);
and AND3 (N104, N101, N95, N20);
or OR2 (N105, N29, N18);
and AND3 (N106, N74, N93, N18);
buf BUF1 (N107, N3);
not NOT1 (N108, N100);
nand NAND2 (N109, N103, N37);
nor NOR4 (N110, N98, N106, N50, N35);
and AND2 (N111, N63, N47);
or OR4 (N112, N109, N86, N39, N28);
nor NOR4 (N113, N85, N55, N69, N106);
and AND2 (N114, N105, N78);
nand NAND3 (N115, N114, N64, N92);
or OR2 (N116, N91, N11);
buf BUF1 (N117, N79);
nor NOR3 (N118, N111, N44, N98);
nand NAND4 (N119, N116, N57, N86, N86);
nand NAND2 (N120, N115, N43);
xor XOR2 (N121, N104, N56);
nor NOR2 (N122, N117, N63);
xor XOR2 (N123, N119, N101);
nand NAND2 (N124, N123, N83);
nand NAND3 (N125, N124, N29, N50);
and AND3 (N126, N112, N28, N29);
buf BUF1 (N127, N118);
xor XOR2 (N128, N108, N16);
nand NAND2 (N129, N121, N38);
xor XOR2 (N130, N125, N53);
xor XOR2 (N131, N127, N2);
not NOT1 (N132, N129);
nand NAND4 (N133, N113, N52, N42, N60);
not NOT1 (N134, N120);
not NOT1 (N135, N133);
xor XOR2 (N136, N132, N58);
nor NOR2 (N137, N135, N4);
nand NAND3 (N138, N136, N102, N65);
nand NAND3 (N139, N122, N17, N128);
not NOT1 (N140, N129);
and AND2 (N141, N107, N82);
nand NAND4 (N142, N131, N58, N66, N73);
not NOT1 (N143, N110);
not NOT1 (N144, N130);
buf BUF1 (N145, N137);
or OR4 (N146, N142, N79, N9, N85);
nor NOR3 (N147, N134, N126, N97);
nand NAND3 (N148, N144, N67, N68);
and AND3 (N149, N101, N71, N106);
or OR3 (N150, N145, N54, N122);
and AND4 (N151, N148, N123, N104, N91);
not NOT1 (N152, N140);
not NOT1 (N153, N141);
or OR3 (N154, N149, N120, N100);
not NOT1 (N155, N150);
nor NOR4 (N156, N146, N108, N89, N85);
xor XOR2 (N157, N139, N151);
xor XOR2 (N158, N68, N142);
and AND4 (N159, N158, N101, N140, N122);
buf BUF1 (N160, N157);
xor XOR2 (N161, N138, N6);
or OR4 (N162, N143, N94, N101, N141);
xor XOR2 (N163, N152, N109);
nor NOR3 (N164, N156, N162, N155);
xor XOR2 (N165, N9, N23);
or OR2 (N166, N44, N120);
xor XOR2 (N167, N159, N163);
buf BUF1 (N168, N8);
or OR2 (N169, N167, N45);
nor NOR2 (N170, N160, N89);
xor XOR2 (N171, N161, N102);
xor XOR2 (N172, N164, N95);
or OR2 (N173, N165, N41);
or OR2 (N174, N168, N24);
and AND4 (N175, N172, N79, N14, N124);
xor XOR2 (N176, N175, N32);
xor XOR2 (N177, N166, N170);
xor XOR2 (N178, N135, N139);
nand NAND2 (N179, N154, N79);
xor XOR2 (N180, N179, N36);
not NOT1 (N181, N169);
buf BUF1 (N182, N171);
nor NOR3 (N183, N177, N181, N10);
and AND2 (N184, N183, N64);
not NOT1 (N185, N133);
and AND4 (N186, N180, N133, N38, N156);
nor NOR2 (N187, N178, N76);
not NOT1 (N188, N153);
and AND3 (N189, N187, N107, N167);
and AND4 (N190, N174, N131, N172, N25);
and AND3 (N191, N189, N77, N52);
and AND3 (N192, N185, N144, N54);
buf BUF1 (N193, N182);
not NOT1 (N194, N191);
or OR4 (N195, N194, N131, N94, N36);
nor NOR4 (N196, N192, N136, N7, N37);
xor XOR2 (N197, N196, N48);
buf BUF1 (N198, N195);
nand NAND2 (N199, N188, N174);
and AND3 (N200, N198, N111, N132);
nand NAND2 (N201, N193, N62);
not NOT1 (N202, N176);
or OR3 (N203, N147, N126, N32);
and AND2 (N204, N203, N123);
nor NOR2 (N205, N197, N84);
and AND2 (N206, N202, N34);
buf BUF1 (N207, N206);
or OR4 (N208, N200, N194, N95, N59);
not NOT1 (N209, N186);
and AND2 (N210, N208, N200);
not NOT1 (N211, N207);
nand NAND2 (N212, N199, N104);
not NOT1 (N213, N184);
or OR3 (N214, N205, N104, N70);
or OR2 (N215, N213, N181);
nor NOR3 (N216, N212, N214, N35);
nand NAND4 (N217, N207, N73, N210, N100);
and AND4 (N218, N123, N64, N114, N43);
xor XOR2 (N219, N173, N7);
and AND3 (N220, N216, N167, N38);
or OR4 (N221, N211, N61, N110, N172);
not NOT1 (N222, N204);
buf BUF1 (N223, N220);
xor XOR2 (N224, N201, N178);
not NOT1 (N225, N222);
xor XOR2 (N226, N225, N95);
not NOT1 (N227, N221);
or OR3 (N228, N218, N160, N108);
nor NOR3 (N229, N190, N126, N120);
or OR3 (N230, N228, N122, N68);
or OR4 (N231, N209, N14, N230, N93);
nor NOR3 (N232, N223, N67, N22);
buf BUF1 (N233, N148);
xor XOR2 (N234, N227, N39);
not NOT1 (N235, N231);
not NOT1 (N236, N232);
or OR2 (N237, N224, N95);
nand NAND2 (N238, N215, N203);
xor XOR2 (N239, N237, N68);
nand NAND3 (N240, N226, N83, N31);
nand NAND2 (N241, N238, N147);
nand NAND2 (N242, N236, N21);
nand NAND3 (N243, N242, N179, N207);
and AND2 (N244, N243, N93);
nand NAND4 (N245, N234, N92, N186, N51);
and AND4 (N246, N229, N48, N81, N199);
nand NAND4 (N247, N245, N200, N185, N85);
nor NOR2 (N248, N246, N151);
not NOT1 (N249, N235);
xor XOR2 (N250, N217, N239);
nand NAND3 (N251, N129, N41, N8);
xor XOR2 (N252, N247, N163);
not NOT1 (N253, N219);
not NOT1 (N254, N244);
nand NAND3 (N255, N248, N35, N116);
and AND4 (N256, N250, N12, N245, N32);
nor NOR2 (N257, N233, N59);
nand NAND2 (N258, N251, N153);
nand NAND2 (N259, N249, N202);
and AND2 (N260, N256, N247);
xor XOR2 (N261, N258, N131);
nand NAND3 (N262, N240, N55, N16);
buf BUF1 (N263, N262);
nor NOR4 (N264, N263, N96, N45, N174);
nor NOR3 (N265, N254, N86, N107);
buf BUF1 (N266, N241);
buf BUF1 (N267, N252);
not NOT1 (N268, N261);
buf BUF1 (N269, N259);
or OR4 (N270, N268, N198, N70, N106);
and AND3 (N271, N267, N221, N96);
nor NOR2 (N272, N257, N63);
not NOT1 (N273, N253);
and AND4 (N274, N265, N247, N230, N90);
or OR3 (N275, N260, N28, N242);
nor NOR4 (N276, N264, N103, N60, N103);
not NOT1 (N277, N274);
or OR4 (N278, N272, N245, N6, N7);
nor NOR3 (N279, N255, N259, N134);
not NOT1 (N280, N269);
and AND3 (N281, N277, N209, N151);
nor NOR2 (N282, N280, N169);
buf BUF1 (N283, N279);
buf BUF1 (N284, N276);
and AND2 (N285, N266, N225);
nor NOR2 (N286, N282, N136);
and AND2 (N287, N285, N143);
and AND2 (N288, N287, N147);
not NOT1 (N289, N273);
nand NAND3 (N290, N288, N272, N70);
not NOT1 (N291, N278);
or OR4 (N292, N290, N5, N194, N165);
or OR2 (N293, N283, N130);
nand NAND4 (N294, N286, N121, N75, N196);
buf BUF1 (N295, N275);
xor XOR2 (N296, N291, N20);
buf BUF1 (N297, N293);
nand NAND2 (N298, N284, N17);
nand NAND2 (N299, N296, N66);
buf BUF1 (N300, N281);
and AND4 (N301, N299, N1, N172, N19);
nor NOR2 (N302, N297, N263);
buf BUF1 (N303, N270);
nor NOR3 (N304, N295, N239, N60);
xor XOR2 (N305, N294, N17);
not NOT1 (N306, N301);
or OR4 (N307, N303, N1, N155, N194);
not NOT1 (N308, N302);
nand NAND3 (N309, N304, N135, N79);
nor NOR4 (N310, N307, N217, N110, N225);
not NOT1 (N311, N308);
nand NAND3 (N312, N306, N66, N311);
or OR3 (N313, N123, N180, N196);
nor NOR4 (N314, N271, N273, N128, N298);
xor XOR2 (N315, N115, N236);
xor XOR2 (N316, N313, N25);
and AND3 (N317, N310, N41, N174);
buf BUF1 (N318, N305);
xor XOR2 (N319, N312, N186);
and AND3 (N320, N292, N177, N44);
nand NAND2 (N321, N289, N205);
nand NAND4 (N322, N318, N277, N54, N85);
nor NOR2 (N323, N314, N232);
nor NOR3 (N324, N309, N113, N285);
nand NAND2 (N325, N320, N153);
xor XOR2 (N326, N322, N133);
not NOT1 (N327, N321);
and AND2 (N328, N317, N71);
not NOT1 (N329, N315);
nor NOR4 (N330, N325, N166, N98, N267);
xor XOR2 (N331, N326, N202);
xor XOR2 (N332, N329, N123);
nand NAND2 (N333, N324, N122);
nand NAND2 (N334, N331, N244);
not NOT1 (N335, N327);
or OR4 (N336, N316, N306, N180, N226);
nor NOR3 (N337, N334, N188, N148);
and AND4 (N338, N328, N2, N113, N112);
not NOT1 (N339, N336);
nand NAND2 (N340, N333, N246);
nand NAND4 (N341, N319, N166, N151, N195);
buf BUF1 (N342, N341);
buf BUF1 (N343, N339);
nand NAND4 (N344, N332, N160, N50, N155);
and AND4 (N345, N337, N10, N108, N12);
buf BUF1 (N346, N300);
buf BUF1 (N347, N346);
not NOT1 (N348, N340);
buf BUF1 (N349, N347);
nand NAND4 (N350, N335, N82, N335, N153);
nor NOR2 (N351, N348, N137);
or OR2 (N352, N338, N316);
and AND3 (N353, N351, N276, N110);
not NOT1 (N354, N349);
xor XOR2 (N355, N342, N340);
xor XOR2 (N356, N344, N127);
and AND4 (N357, N356, N242, N178, N252);
not NOT1 (N358, N353);
buf BUF1 (N359, N345);
nand NAND2 (N360, N330, N81);
xor XOR2 (N361, N354, N202);
nand NAND4 (N362, N352, N2, N1, N59);
buf BUF1 (N363, N343);
nor NOR2 (N364, N358, N13);
not NOT1 (N365, N361);
not NOT1 (N366, N357);
not NOT1 (N367, N350);
buf BUF1 (N368, N364);
xor XOR2 (N369, N365, N209);
buf BUF1 (N370, N368);
xor XOR2 (N371, N362, N316);
or OR3 (N372, N370, N12, N23);
buf BUF1 (N373, N369);
nor NOR2 (N374, N360, N301);
nand NAND2 (N375, N374, N128);
and AND4 (N376, N367, N260, N63, N42);
nand NAND2 (N377, N373, N367);
not NOT1 (N378, N363);
not NOT1 (N379, N355);
or OR2 (N380, N379, N18);
nor NOR2 (N381, N377, N42);
nand NAND2 (N382, N366, N70);
and AND4 (N383, N375, N69, N187, N238);
nor NOR4 (N384, N371, N277, N317, N97);
and AND4 (N385, N378, N185, N312, N210);
buf BUF1 (N386, N372);
nor NOR2 (N387, N359, N108);
or OR3 (N388, N387, N273, N276);
not NOT1 (N389, N382);
not NOT1 (N390, N381);
nand NAND4 (N391, N384, N362, N35, N208);
or OR4 (N392, N389, N235, N13, N321);
and AND4 (N393, N385, N143, N49, N141);
nand NAND4 (N394, N383, N244, N47, N93);
and AND4 (N395, N388, N364, N186, N136);
xor XOR2 (N396, N376, N278);
xor XOR2 (N397, N390, N72);
and AND2 (N398, N393, N49);
xor XOR2 (N399, N397, N291);
xor XOR2 (N400, N391, N4);
buf BUF1 (N401, N323);
nand NAND2 (N402, N396, N246);
and AND3 (N403, N398, N200, N326);
nand NAND2 (N404, N399, N303);
or OR3 (N405, N404, N191, N54);
and AND2 (N406, N401, N343);
and AND4 (N407, N403, N226, N131, N209);
not NOT1 (N408, N405);
xor XOR2 (N409, N392, N351);
buf BUF1 (N410, N380);
xor XOR2 (N411, N408, N254);
xor XOR2 (N412, N394, N202);
nor NOR3 (N413, N407, N214, N393);
nand NAND3 (N414, N386, N108, N200);
not NOT1 (N415, N395);
xor XOR2 (N416, N409, N202);
nand NAND3 (N417, N416, N87, N133);
nor NOR2 (N418, N410, N389);
and AND4 (N419, N411, N13, N104, N410);
nand NAND2 (N420, N402, N206);
or OR4 (N421, N418, N189, N377, N28);
nand NAND2 (N422, N414, N62);
xor XOR2 (N423, N417, N317);
nor NOR3 (N424, N419, N241, N310);
not NOT1 (N425, N415);
xor XOR2 (N426, N423, N323);
or OR3 (N427, N413, N426, N353);
and AND2 (N428, N398, N233);
and AND4 (N429, N412, N96, N45, N186);
nand NAND3 (N430, N400, N395, N324);
or OR3 (N431, N428, N43, N157);
and AND2 (N432, N431, N46);
nand NAND3 (N433, N432, N2, N224);
and AND2 (N434, N430, N156);
nor NOR2 (N435, N406, N135);
xor XOR2 (N436, N422, N135);
nor NOR3 (N437, N420, N407, N252);
not NOT1 (N438, N434);
nor NOR2 (N439, N429, N149);
nand NAND2 (N440, N435, N439);
nand NAND4 (N441, N311, N405, N396, N116);
or OR3 (N442, N440, N98, N179);
not NOT1 (N443, N424);
and AND2 (N444, N443, N419);
nand NAND4 (N445, N438, N304, N202, N376);
and AND3 (N446, N441, N52, N250);
buf BUF1 (N447, N433);
not NOT1 (N448, N436);
or OR3 (N449, N421, N68, N239);
buf BUF1 (N450, N447);
xor XOR2 (N451, N437, N116);
and AND2 (N452, N442, N274);
nor NOR3 (N453, N448, N227, N40);
buf BUF1 (N454, N449);
and AND2 (N455, N427, N440);
buf BUF1 (N456, N444);
or OR4 (N457, N452, N282, N74, N7);
or OR3 (N458, N445, N175, N298);
not NOT1 (N459, N458);
nand NAND2 (N460, N455, N413);
nand NAND2 (N461, N451, N210);
not NOT1 (N462, N460);
buf BUF1 (N463, N453);
buf BUF1 (N464, N457);
buf BUF1 (N465, N446);
and AND2 (N466, N454, N280);
nand NAND3 (N467, N464, N391, N354);
buf BUF1 (N468, N461);
nand NAND4 (N469, N468, N96, N274, N13);
not NOT1 (N470, N450);
and AND4 (N471, N459, N21, N451, N38);
nor NOR3 (N472, N471, N263, N199);
nor NOR2 (N473, N466, N457);
or OR3 (N474, N472, N332, N43);
xor XOR2 (N475, N462, N425);
nor NOR3 (N476, N144, N23, N56);
or OR2 (N477, N475, N165);
and AND4 (N478, N474, N396, N363, N251);
nand NAND2 (N479, N476, N113);
and AND4 (N480, N456, N280, N408, N182);
and AND3 (N481, N480, N125, N136);
buf BUF1 (N482, N473);
or OR4 (N483, N479, N381, N463, N387);
and AND4 (N484, N303, N168, N130, N480);
and AND4 (N485, N478, N15, N271, N298);
nand NAND4 (N486, N483, N406, N451, N203);
not NOT1 (N487, N477);
or OR2 (N488, N484, N206);
not NOT1 (N489, N485);
buf BUF1 (N490, N489);
and AND2 (N491, N490, N71);
xor XOR2 (N492, N467, N330);
nor NOR2 (N493, N470, N123);
and AND2 (N494, N469, N77);
nor NOR2 (N495, N494, N457);
and AND4 (N496, N493, N478, N138, N177);
not NOT1 (N497, N486);
nand NAND3 (N498, N488, N29, N216);
or OR3 (N499, N497, N320, N199);
or OR2 (N500, N492, N394);
nand NAND2 (N501, N482, N471);
xor XOR2 (N502, N499, N25);
xor XOR2 (N503, N495, N414);
nand NAND4 (N504, N496, N231, N97, N140);
nand NAND2 (N505, N487, N495);
not NOT1 (N506, N501);
not NOT1 (N507, N498);
not NOT1 (N508, N502);
buf BUF1 (N509, N500);
or OR4 (N510, N505, N254, N231, N438);
nand NAND2 (N511, N481, N28);
or OR2 (N512, N509, N328);
nor NOR2 (N513, N511, N455);
xor XOR2 (N514, N504, N462);
not NOT1 (N515, N513);
and AND4 (N516, N514, N131, N388, N459);
or OR2 (N517, N508, N392);
nand NAND2 (N518, N510, N253);
and AND2 (N519, N516, N27);
buf BUF1 (N520, N518);
buf BUF1 (N521, N491);
buf BUF1 (N522, N465);
buf BUF1 (N523, N522);
not NOT1 (N524, N521);
nand NAND4 (N525, N520, N186, N411, N486);
buf BUF1 (N526, N524);
nor NOR4 (N527, N512, N115, N53, N502);
not NOT1 (N528, N525);
and AND2 (N529, N503, N95);
or OR4 (N530, N527, N326, N305, N133);
or OR3 (N531, N529, N420, N390);
or OR3 (N532, N526, N8, N146);
xor XOR2 (N533, N528, N106);
or OR3 (N534, N517, N475, N221);
nor NOR4 (N535, N507, N54, N361, N60);
nand NAND2 (N536, N515, N520);
nand NAND4 (N537, N506, N466, N123, N320);
nand NAND2 (N538, N535, N363);
and AND4 (N539, N519, N17, N391, N282);
or OR3 (N540, N538, N439, N395);
buf BUF1 (N541, N532);
xor XOR2 (N542, N531, N384);
and AND3 (N543, N533, N283, N307);
and AND3 (N544, N542, N23, N311);
nand NAND2 (N545, N544, N484);
xor XOR2 (N546, N537, N409);
nor NOR3 (N547, N530, N477, N429);
or OR2 (N548, N541, N294);
or OR3 (N549, N547, N422, N310);
buf BUF1 (N550, N545);
not NOT1 (N551, N550);
and AND3 (N552, N549, N82, N460);
and AND4 (N553, N539, N290, N413, N163);
or OR3 (N554, N551, N233, N445);
not NOT1 (N555, N534);
and AND3 (N556, N552, N532, N467);
or OR4 (N557, N546, N353, N540, N381);
nand NAND3 (N558, N464, N210, N112);
nor NOR4 (N559, N548, N211, N425, N157);
nor NOR4 (N560, N554, N514, N37, N371);
buf BUF1 (N561, N553);
nor NOR4 (N562, N560, N151, N305, N310);
and AND2 (N563, N543, N284);
and AND3 (N564, N558, N116, N178);
nor NOR2 (N565, N564, N536);
nand NAND4 (N566, N53, N236, N447, N206);
buf BUF1 (N567, N555);
not NOT1 (N568, N562);
buf BUF1 (N569, N559);
buf BUF1 (N570, N563);
or OR2 (N571, N569, N272);
or OR2 (N572, N570, N483);
xor XOR2 (N573, N572, N38);
nand NAND2 (N574, N568, N270);
nand NAND3 (N575, N557, N485, N57);
not NOT1 (N576, N523);
nand NAND4 (N577, N567, N460, N230, N228);
buf BUF1 (N578, N576);
or OR2 (N579, N575, N238);
nand NAND2 (N580, N577, N287);
nand NAND4 (N581, N566, N14, N87, N401);
or OR3 (N582, N571, N86, N12);
nor NOR2 (N583, N582, N478);
buf BUF1 (N584, N579);
and AND4 (N585, N561, N309, N7, N421);
and AND3 (N586, N556, N525, N91);
nor NOR3 (N587, N578, N418, N447);
or OR4 (N588, N581, N564, N538, N514);
nand NAND3 (N589, N573, N507, N457);
not NOT1 (N590, N587);
not NOT1 (N591, N583);
or OR4 (N592, N589, N147, N536, N414);
not NOT1 (N593, N591);
buf BUF1 (N594, N592);
buf BUF1 (N595, N584);
or OR4 (N596, N574, N509, N144, N574);
and AND3 (N597, N586, N555, N40);
buf BUF1 (N598, N595);
nor NOR3 (N599, N598, N261, N200);
not NOT1 (N600, N596);
xor XOR2 (N601, N565, N168);
and AND4 (N602, N585, N443, N115, N580);
nand NAND2 (N603, N209, N260);
nor NOR2 (N604, N588, N554);
nand NAND2 (N605, N593, N144);
not NOT1 (N606, N599);
xor XOR2 (N607, N600, N532);
and AND3 (N608, N606, N374, N414);
and AND2 (N609, N594, N472);
buf BUF1 (N610, N601);
buf BUF1 (N611, N597);
nor NOR3 (N612, N610, N261, N491);
and AND3 (N613, N609, N558, N203);
xor XOR2 (N614, N611, N234);
endmodule