// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N3514,N3512,N3515,N3518,N3517,N3510,N3513,N3516,N3507,N3519;

and AND2 (N20, N4, N16);
nor NOR2 (N21, N17, N2);
not NOT1 (N22, N6);
nand NAND3 (N23, N15, N13, N21);
buf BUF1 (N24, N12);
nor NOR2 (N25, N7, N11);
xor XOR2 (N26, N18, N25);
and AND2 (N27, N18, N10);
xor XOR2 (N28, N3, N2);
xor XOR2 (N29, N16, N18);
not NOT1 (N30, N16);
and AND2 (N31, N8, N25);
nor NOR4 (N32, N27, N10, N7, N9);
xor XOR2 (N33, N24, N24);
not NOT1 (N34, N22);
or OR3 (N35, N23, N21, N1);
buf BUF1 (N36, N31);
nand NAND4 (N37, N20, N26, N34, N19);
buf BUF1 (N38, N14);
or OR4 (N39, N24, N25, N9, N12);
buf BUF1 (N40, N28);
xor XOR2 (N41, N40, N32);
nand NAND3 (N42, N13, N28, N38);
buf BUF1 (N43, N31);
buf BUF1 (N44, N42);
nor NOR4 (N45, N44, N34, N29, N17);
buf BUF1 (N46, N28);
nand NAND3 (N47, N39, N25, N32);
buf BUF1 (N48, N43);
nor NOR3 (N49, N36, N23, N17);
nand NAND3 (N50, N48, N16, N38);
buf BUF1 (N51, N49);
or OR3 (N52, N51, N23, N39);
buf BUF1 (N53, N45);
and AND4 (N54, N46, N42, N22, N9);
not NOT1 (N55, N37);
not NOT1 (N56, N54);
nand NAND2 (N57, N47, N10);
and AND3 (N58, N53, N32, N40);
and AND4 (N59, N50, N40, N32, N15);
or OR3 (N60, N59, N16, N34);
not NOT1 (N61, N52);
nor NOR4 (N62, N30, N29, N56, N22);
nor NOR2 (N63, N58, N6);
nor NOR2 (N64, N3, N42);
buf BUF1 (N65, N57);
not NOT1 (N66, N61);
buf BUF1 (N67, N65);
or OR2 (N68, N33, N17);
xor XOR2 (N69, N66, N51);
or OR4 (N70, N67, N29, N46, N65);
nor NOR4 (N71, N70, N55, N48, N48);
or OR4 (N72, N58, N33, N71, N3);
nand NAND4 (N73, N37, N13, N5, N17);
not NOT1 (N74, N41);
or OR3 (N75, N63, N6, N2);
xor XOR2 (N76, N75, N24);
xor XOR2 (N77, N73, N50);
and AND4 (N78, N68, N21, N20, N73);
and AND3 (N79, N60, N38, N54);
not NOT1 (N80, N77);
and AND4 (N81, N74, N64, N40, N76);
nand NAND4 (N82, N76, N40, N65, N73);
nor NOR4 (N83, N67, N44, N1, N29);
not NOT1 (N84, N80);
buf BUF1 (N85, N81);
and AND4 (N86, N83, N24, N82, N16);
not NOT1 (N87, N11);
nand NAND4 (N88, N78, N30, N36, N11);
and AND2 (N89, N85, N19);
nor NOR4 (N90, N35, N61, N30, N53);
or OR4 (N91, N84, N19, N46, N74);
or OR2 (N92, N72, N60);
nand NAND2 (N93, N86, N56);
xor XOR2 (N94, N92, N85);
xor XOR2 (N95, N88, N24);
xor XOR2 (N96, N79, N70);
buf BUF1 (N97, N95);
nor NOR2 (N98, N93, N70);
buf BUF1 (N99, N62);
xor XOR2 (N100, N94, N16);
not NOT1 (N101, N99);
and AND3 (N102, N97, N49, N68);
buf BUF1 (N103, N102);
nor NOR2 (N104, N69, N62);
buf BUF1 (N105, N89);
not NOT1 (N106, N103);
not NOT1 (N107, N101);
not NOT1 (N108, N87);
nor NOR2 (N109, N98, N20);
nor NOR4 (N110, N100, N57, N96, N102);
or OR4 (N111, N60, N39, N104, N34);
and AND3 (N112, N78, N20, N41);
nor NOR2 (N113, N112, N103);
not NOT1 (N114, N111);
or OR4 (N115, N108, N79, N27, N51);
nor NOR4 (N116, N115, N22, N86, N94);
xor XOR2 (N117, N105, N92);
xor XOR2 (N118, N107, N46);
nand NAND2 (N119, N118, N86);
nand NAND4 (N120, N116, N16, N39, N69);
nor NOR3 (N121, N91, N43, N55);
not NOT1 (N122, N110);
buf BUF1 (N123, N117);
nand NAND4 (N124, N114, N77, N44, N52);
nor NOR4 (N125, N109, N118, N21, N71);
not NOT1 (N126, N120);
not NOT1 (N127, N113);
xor XOR2 (N128, N90, N113);
nand NAND3 (N129, N122, N2, N77);
and AND4 (N130, N128, N55, N53, N74);
xor XOR2 (N131, N106, N95);
nor NOR3 (N132, N129, N43, N44);
not NOT1 (N133, N123);
and AND2 (N134, N124, N4);
buf BUF1 (N135, N121);
buf BUF1 (N136, N127);
not NOT1 (N137, N134);
not NOT1 (N138, N136);
xor XOR2 (N139, N135, N101);
xor XOR2 (N140, N126, N21);
and AND4 (N141, N139, N78, N2, N80);
nor NOR2 (N142, N132, N128);
xor XOR2 (N143, N137, N11);
nor NOR2 (N144, N142, N87);
nor NOR3 (N145, N133, N15, N89);
or OR3 (N146, N125, N9, N28);
nor NOR4 (N147, N119, N103, N97, N110);
not NOT1 (N148, N146);
or OR3 (N149, N131, N113, N87);
nand NAND3 (N150, N145, N102, N22);
and AND4 (N151, N130, N5, N116, N79);
nand NAND2 (N152, N151, N91);
xor XOR2 (N153, N152, N99);
xor XOR2 (N154, N153, N133);
nand NAND2 (N155, N150, N149);
or OR4 (N156, N9, N150, N75, N20);
nor NOR3 (N157, N147, N91, N50);
buf BUF1 (N158, N141);
nor NOR2 (N159, N158, N146);
nor NOR4 (N160, N144, N154, N95, N11);
and AND2 (N161, N136, N109);
buf BUF1 (N162, N138);
buf BUF1 (N163, N162);
xor XOR2 (N164, N148, N107);
nand NAND4 (N165, N157, N113, N88, N157);
not NOT1 (N166, N164);
and AND4 (N167, N143, N43, N56, N3);
or OR2 (N168, N166, N138);
xor XOR2 (N169, N140, N162);
buf BUF1 (N170, N161);
nand NAND3 (N171, N170, N19, N113);
buf BUF1 (N172, N169);
nor NOR2 (N173, N156, N30);
xor XOR2 (N174, N159, N160);
buf BUF1 (N175, N25);
xor XOR2 (N176, N155, N6);
buf BUF1 (N177, N172);
and AND3 (N178, N168, N170, N169);
and AND3 (N179, N167, N133, N167);
buf BUF1 (N180, N163);
and AND2 (N181, N178, N49);
and AND3 (N182, N171, N123, N85);
nand NAND3 (N183, N180, N77, N72);
nand NAND4 (N184, N182, N47, N59, N149);
nand NAND3 (N185, N165, N125, N132);
or OR4 (N186, N173, N25, N176, N134);
and AND3 (N187, N77, N22, N122);
nand NAND3 (N188, N186, N63, N87);
or OR2 (N189, N184, N79);
or OR2 (N190, N187, N141);
xor XOR2 (N191, N183, N185);
xor XOR2 (N192, N40, N41);
xor XOR2 (N193, N181, N103);
nor NOR2 (N194, N179, N119);
and AND2 (N195, N190, N176);
buf BUF1 (N196, N192);
nand NAND4 (N197, N174, N51, N157, N167);
and AND3 (N198, N193, N150, N93);
nor NOR3 (N199, N197, N130, N34);
xor XOR2 (N200, N194, N187);
not NOT1 (N201, N188);
nor NOR3 (N202, N177, N59, N147);
not NOT1 (N203, N200);
nor NOR2 (N204, N196, N86);
or OR4 (N205, N195, N24, N186, N101);
or OR3 (N206, N205, N189, N171);
and AND2 (N207, N64, N104);
and AND3 (N208, N206, N150, N88);
not NOT1 (N209, N201);
buf BUF1 (N210, N203);
or OR4 (N211, N209, N17, N160, N177);
xor XOR2 (N212, N204, N93);
nor NOR2 (N213, N212, N111);
and AND2 (N214, N175, N177);
and AND3 (N215, N207, N57, N200);
and AND3 (N216, N215, N16, N27);
or OR4 (N217, N199, N107, N62, N61);
not NOT1 (N218, N191);
and AND3 (N219, N218, N93, N109);
and AND4 (N220, N210, N205, N203, N216);
buf BUF1 (N221, N72);
buf BUF1 (N222, N220);
or OR2 (N223, N219, N151);
nand NAND4 (N224, N208, N222, N129, N156);
nor NOR4 (N225, N185, N156, N42, N34);
and AND2 (N226, N217, N196);
nor NOR3 (N227, N224, N1, N142);
buf BUF1 (N228, N223);
nor NOR2 (N229, N202, N122);
xor XOR2 (N230, N228, N63);
xor XOR2 (N231, N225, N69);
nand NAND2 (N232, N227, N198);
xor XOR2 (N233, N36, N125);
and AND3 (N234, N214, N142, N232);
xor XOR2 (N235, N175, N191);
and AND4 (N236, N211, N27, N210, N140);
xor XOR2 (N237, N233, N54);
and AND4 (N238, N221, N177, N199, N124);
and AND3 (N239, N238, N199, N97);
xor XOR2 (N240, N231, N32);
nor NOR3 (N241, N235, N87, N2);
xor XOR2 (N242, N240, N98);
nand NAND2 (N243, N213, N178);
buf BUF1 (N244, N236);
buf BUF1 (N245, N230);
nand NAND2 (N246, N239, N222);
not NOT1 (N247, N245);
nor NOR2 (N248, N243, N208);
not NOT1 (N249, N242);
xor XOR2 (N250, N229, N57);
and AND3 (N251, N237, N237, N134);
not NOT1 (N252, N244);
and AND3 (N253, N248, N227, N93);
xor XOR2 (N254, N234, N81);
and AND2 (N255, N241, N232);
nor NOR3 (N256, N250, N97, N250);
not NOT1 (N257, N226);
xor XOR2 (N258, N246, N175);
xor XOR2 (N259, N249, N77);
buf BUF1 (N260, N251);
or OR2 (N261, N247, N222);
nand NAND2 (N262, N253, N106);
buf BUF1 (N263, N257);
or OR2 (N264, N261, N49);
and AND4 (N265, N255, N103, N192, N46);
nand NAND4 (N266, N259, N114, N196, N129);
and AND3 (N267, N264, N30, N184);
xor XOR2 (N268, N262, N192);
and AND4 (N269, N258, N127, N142, N180);
xor XOR2 (N270, N265, N209);
or OR3 (N271, N260, N252, N155);
not NOT1 (N272, N258);
buf BUF1 (N273, N267);
or OR4 (N274, N270, N161, N201, N167);
nand NAND4 (N275, N269, N177, N133, N118);
and AND2 (N276, N275, N220);
nand NAND4 (N277, N263, N168, N42, N129);
xor XOR2 (N278, N272, N50);
nor NOR4 (N279, N254, N173, N187, N249);
nand NAND3 (N280, N278, N208, N222);
xor XOR2 (N281, N277, N98);
nand NAND3 (N282, N271, N71, N4);
and AND2 (N283, N276, N68);
or OR2 (N284, N282, N154);
not NOT1 (N285, N274);
and AND4 (N286, N285, N202, N264, N28);
xor XOR2 (N287, N268, N238);
nand NAND2 (N288, N281, N155);
nand NAND4 (N289, N288, N6, N73, N104);
and AND3 (N290, N279, N234, N25);
nand NAND4 (N291, N283, N49, N269, N145);
xor XOR2 (N292, N289, N181);
xor XOR2 (N293, N266, N180);
nor NOR2 (N294, N291, N17);
buf BUF1 (N295, N280);
buf BUF1 (N296, N295);
or OR4 (N297, N286, N231, N13, N84);
and AND4 (N298, N273, N23, N281, N131);
nand NAND2 (N299, N293, N129);
xor XOR2 (N300, N298, N159);
not NOT1 (N301, N297);
xor XOR2 (N302, N294, N9);
and AND2 (N303, N284, N302);
buf BUF1 (N304, N36);
or OR3 (N305, N303, N74, N266);
nand NAND4 (N306, N292, N249, N217, N202);
xor XOR2 (N307, N256, N251);
nor NOR2 (N308, N306, N274);
or OR3 (N309, N300, N213, N255);
nand NAND2 (N310, N296, N208);
nand NAND4 (N311, N301, N100, N249, N281);
or OR2 (N312, N310, N189);
nand NAND2 (N313, N312, N186);
and AND3 (N314, N290, N143, N87);
buf BUF1 (N315, N305);
not NOT1 (N316, N313);
buf BUF1 (N317, N287);
and AND4 (N318, N304, N15, N304, N49);
xor XOR2 (N319, N299, N299);
or OR4 (N320, N311, N111, N116, N66);
nand NAND3 (N321, N307, N143, N257);
and AND4 (N322, N317, N102, N241, N284);
or OR3 (N323, N319, N249, N222);
nand NAND2 (N324, N323, N189);
and AND4 (N325, N320, N89, N66, N87);
buf BUF1 (N326, N318);
and AND2 (N327, N322, N122);
or OR4 (N328, N327, N253, N105, N147);
not NOT1 (N329, N308);
not NOT1 (N330, N326);
not NOT1 (N331, N330);
not NOT1 (N332, N314);
nor NOR3 (N333, N332, N94, N290);
or OR4 (N334, N333, N10, N158, N63);
nand NAND3 (N335, N331, N9, N242);
not NOT1 (N336, N325);
and AND3 (N337, N309, N177, N43);
nor NOR2 (N338, N335, N137);
nor NOR4 (N339, N321, N207, N260, N113);
or OR3 (N340, N338, N28, N156);
xor XOR2 (N341, N316, N81);
and AND4 (N342, N329, N129, N175, N320);
nor NOR2 (N343, N339, N256);
or OR4 (N344, N341, N181, N324, N234);
buf BUF1 (N345, N93);
buf BUF1 (N346, N342);
or OR2 (N347, N345, N47);
nor NOR4 (N348, N343, N175, N166, N336);
nand NAND4 (N349, N31, N181, N324, N99);
and AND2 (N350, N349, N333);
not NOT1 (N351, N315);
xor XOR2 (N352, N337, N238);
nor NOR2 (N353, N351, N251);
or OR3 (N354, N348, N15, N256);
xor XOR2 (N355, N334, N277);
buf BUF1 (N356, N352);
buf BUF1 (N357, N356);
or OR2 (N358, N344, N235);
nor NOR3 (N359, N340, N119, N155);
or OR2 (N360, N358, N315);
nand NAND3 (N361, N360, N43, N180);
or OR2 (N362, N361, N229);
xor XOR2 (N363, N350, N226);
buf BUF1 (N364, N357);
buf BUF1 (N365, N353);
or OR4 (N366, N363, N218, N104, N31);
not NOT1 (N367, N362);
nand NAND3 (N368, N364, N222, N341);
nor NOR3 (N369, N355, N73, N285);
not NOT1 (N370, N365);
not NOT1 (N371, N347);
nand NAND4 (N372, N370, N288, N228, N102);
buf BUF1 (N373, N354);
not NOT1 (N374, N372);
nand NAND4 (N375, N367, N112, N52, N222);
nor NOR2 (N376, N328, N47);
nand NAND2 (N377, N373, N99);
or OR2 (N378, N374, N153);
and AND3 (N379, N378, N194, N178);
nor NOR4 (N380, N371, N114, N368, N264);
xor XOR2 (N381, N161, N101);
buf BUF1 (N382, N359);
not NOT1 (N383, N377);
not NOT1 (N384, N383);
not NOT1 (N385, N369);
buf BUF1 (N386, N384);
and AND2 (N387, N346, N276);
or OR4 (N388, N382, N366, N96, N295);
buf BUF1 (N389, N209);
not NOT1 (N390, N386);
and AND2 (N391, N380, N40);
and AND2 (N392, N375, N262);
not NOT1 (N393, N391);
buf BUF1 (N394, N388);
and AND2 (N395, N381, N315);
buf BUF1 (N396, N385);
and AND2 (N397, N396, N77);
not NOT1 (N398, N392);
and AND2 (N399, N379, N297);
nand NAND3 (N400, N398, N21, N56);
nor NOR3 (N401, N389, N140, N313);
xor XOR2 (N402, N395, N163);
nand NAND4 (N403, N402, N118, N155, N36);
and AND4 (N404, N401, N52, N106, N17);
not NOT1 (N405, N393);
nor NOR4 (N406, N403, N265, N22, N76);
nor NOR4 (N407, N404, N196, N211, N264);
xor XOR2 (N408, N397, N25);
not NOT1 (N409, N406);
or OR4 (N410, N376, N375, N30, N190);
buf BUF1 (N411, N407);
or OR3 (N412, N394, N384, N66);
xor XOR2 (N413, N408, N173);
nor NOR3 (N414, N413, N283, N320);
nand NAND2 (N415, N399, N18);
nand NAND3 (N416, N409, N187, N54);
and AND3 (N417, N412, N88, N347);
or OR3 (N418, N417, N139, N157);
buf BUF1 (N419, N390);
and AND3 (N420, N410, N145, N121);
nor NOR4 (N421, N416, N366, N389, N85);
or OR2 (N422, N415, N317);
or OR4 (N423, N411, N414, N162, N267);
or OR4 (N424, N282, N320, N311, N277);
nor NOR3 (N425, N421, N77, N198);
nand NAND3 (N426, N422, N175, N355);
not NOT1 (N427, N405);
buf BUF1 (N428, N400);
nand NAND4 (N429, N420, N81, N110, N168);
nand NAND3 (N430, N429, N276, N55);
or OR3 (N431, N423, N407, N387);
nand NAND2 (N432, N272, N185);
xor XOR2 (N433, N431, N266);
and AND3 (N434, N433, N116, N54);
buf BUF1 (N435, N427);
nand NAND2 (N436, N419, N392);
nor NOR3 (N437, N426, N310, N80);
buf BUF1 (N438, N434);
or OR3 (N439, N436, N386, N229);
or OR2 (N440, N418, N34);
or OR3 (N441, N430, N98, N264);
nor NOR2 (N442, N438, N245);
xor XOR2 (N443, N428, N200);
or OR2 (N444, N424, N191);
xor XOR2 (N445, N425, N214);
buf BUF1 (N446, N437);
and AND4 (N447, N441, N193, N155, N390);
not NOT1 (N448, N445);
nand NAND3 (N449, N442, N114, N321);
or OR3 (N450, N440, N71, N33);
nand NAND3 (N451, N446, N180, N29);
buf BUF1 (N452, N448);
nor NOR4 (N453, N451, N72, N172, N61);
or OR3 (N454, N453, N187, N403);
or OR4 (N455, N452, N161, N73, N375);
nand NAND3 (N456, N435, N121, N358);
nand NAND2 (N457, N450, N195);
or OR4 (N458, N447, N376, N26, N362);
buf BUF1 (N459, N439);
or OR3 (N460, N457, N74, N177);
nor NOR3 (N461, N454, N275, N92);
xor XOR2 (N462, N443, N294);
xor XOR2 (N463, N455, N17);
and AND3 (N464, N444, N296, N348);
nor NOR3 (N465, N459, N72, N460);
buf BUF1 (N466, N208);
not NOT1 (N467, N449);
nor NOR2 (N468, N462, N112);
not NOT1 (N469, N466);
nand NAND4 (N470, N461, N21, N254, N359);
and AND2 (N471, N464, N283);
nand NAND2 (N472, N432, N195);
buf BUF1 (N473, N465);
and AND2 (N474, N463, N255);
buf BUF1 (N475, N456);
not NOT1 (N476, N458);
or OR3 (N477, N475, N335, N419);
xor XOR2 (N478, N477, N442);
nand NAND2 (N479, N467, N163);
buf BUF1 (N480, N478);
or OR2 (N481, N471, N343);
or OR4 (N482, N473, N98, N164, N196);
not NOT1 (N483, N469);
or OR2 (N484, N468, N398);
nand NAND3 (N485, N483, N259, N446);
buf BUF1 (N486, N476);
nand NAND4 (N487, N472, N117, N110, N175);
nor NOR2 (N488, N480, N458);
nor NOR4 (N489, N485, N128, N246, N50);
xor XOR2 (N490, N486, N31);
not NOT1 (N491, N474);
not NOT1 (N492, N481);
buf BUF1 (N493, N490);
or OR2 (N494, N493, N35);
or OR4 (N495, N484, N13, N202, N351);
not NOT1 (N496, N495);
not NOT1 (N497, N488);
xor XOR2 (N498, N487, N121);
and AND2 (N499, N479, N145);
and AND2 (N500, N497, N360);
buf BUF1 (N501, N491);
and AND3 (N502, N494, N339, N102);
not NOT1 (N503, N500);
nor NOR2 (N504, N489, N397);
or OR4 (N505, N503, N258, N120, N105);
nand NAND3 (N506, N499, N405, N131);
not NOT1 (N507, N496);
and AND2 (N508, N501, N33);
buf BUF1 (N509, N502);
buf BUF1 (N510, N504);
not NOT1 (N511, N498);
buf BUF1 (N512, N470);
nand NAND3 (N513, N507, N275, N210);
nor NOR2 (N514, N509, N27);
or OR2 (N515, N482, N399);
or OR3 (N516, N511, N226, N412);
nor NOR4 (N517, N512, N367, N327, N342);
or OR4 (N518, N515, N328, N139, N220);
buf BUF1 (N519, N513);
nor NOR2 (N520, N514, N256);
or OR2 (N521, N517, N116);
nand NAND4 (N522, N520, N252, N482, N376);
buf BUF1 (N523, N518);
buf BUF1 (N524, N506);
or OR4 (N525, N524, N204, N179, N13);
not NOT1 (N526, N525);
and AND3 (N527, N516, N264, N12);
or OR2 (N528, N521, N384);
buf BUF1 (N529, N492);
or OR3 (N530, N505, N368, N111);
and AND4 (N531, N519, N508, N27, N146);
and AND4 (N532, N208, N164, N361, N440);
buf BUF1 (N533, N530);
or OR4 (N534, N532, N141, N450, N532);
and AND3 (N535, N533, N104, N30);
xor XOR2 (N536, N535, N483);
xor XOR2 (N537, N536, N57);
nor NOR3 (N538, N531, N405, N162);
and AND2 (N539, N537, N399);
xor XOR2 (N540, N523, N390);
buf BUF1 (N541, N540);
or OR2 (N542, N534, N515);
xor XOR2 (N543, N542, N360);
or OR4 (N544, N539, N159, N496, N236);
or OR3 (N545, N529, N212, N520);
nor NOR3 (N546, N541, N267, N449);
buf BUF1 (N547, N538);
xor XOR2 (N548, N545, N33);
and AND2 (N549, N544, N290);
xor XOR2 (N550, N547, N517);
nand NAND3 (N551, N522, N268, N172);
or OR3 (N552, N526, N273, N401);
buf BUF1 (N553, N543);
nand NAND3 (N554, N553, N96, N88);
or OR4 (N555, N554, N307, N204, N364);
buf BUF1 (N556, N548);
buf BUF1 (N557, N527);
not NOT1 (N558, N551);
buf BUF1 (N559, N546);
nor NOR4 (N560, N558, N255, N268, N122);
nor NOR2 (N561, N560, N351);
xor XOR2 (N562, N561, N337);
nand NAND2 (N563, N549, N267);
xor XOR2 (N564, N552, N338);
or OR4 (N565, N550, N321, N184, N236);
not NOT1 (N566, N562);
and AND2 (N567, N556, N344);
buf BUF1 (N568, N557);
nor NOR4 (N569, N565, N27, N95, N194);
nor NOR3 (N570, N528, N348, N157);
buf BUF1 (N571, N564);
buf BUF1 (N572, N569);
xor XOR2 (N573, N566, N170);
and AND2 (N574, N568, N352);
xor XOR2 (N575, N574, N307);
nor NOR2 (N576, N575, N450);
xor XOR2 (N577, N567, N134);
not NOT1 (N578, N559);
and AND4 (N579, N572, N97, N549, N498);
buf BUF1 (N580, N570);
buf BUF1 (N581, N578);
xor XOR2 (N582, N510, N154);
and AND2 (N583, N582, N438);
nand NAND3 (N584, N555, N490, N329);
nand NAND4 (N585, N573, N473, N554, N247);
or OR2 (N586, N576, N333);
xor XOR2 (N587, N579, N459);
buf BUF1 (N588, N585);
and AND4 (N589, N581, N372, N205, N58);
nand NAND3 (N590, N580, N171, N168);
and AND2 (N591, N586, N315);
nor NOR2 (N592, N589, N332);
or OR2 (N593, N583, N187);
nand NAND2 (N594, N577, N259);
nand NAND3 (N595, N587, N327, N25);
xor XOR2 (N596, N595, N388);
buf BUF1 (N597, N596);
buf BUF1 (N598, N588);
nand NAND3 (N599, N598, N408, N345);
nand NAND4 (N600, N590, N200, N505, N214);
nor NOR4 (N601, N592, N77, N93, N333);
nor NOR2 (N602, N571, N413);
nand NAND4 (N603, N597, N413, N357, N277);
not NOT1 (N604, N603);
nor NOR3 (N605, N599, N207, N590);
xor XOR2 (N606, N601, N99);
and AND3 (N607, N602, N516, N376);
and AND2 (N608, N563, N126);
nor NOR3 (N609, N606, N295, N272);
xor XOR2 (N610, N600, N352);
or OR3 (N611, N605, N175, N340);
not NOT1 (N612, N593);
xor XOR2 (N613, N611, N82);
or OR4 (N614, N594, N604, N442, N220);
xor XOR2 (N615, N90, N69);
nand NAND4 (N616, N591, N108, N304, N79);
buf BUF1 (N617, N616);
and AND2 (N618, N613, N565);
xor XOR2 (N619, N612, N135);
and AND2 (N620, N608, N266);
nor NOR3 (N621, N610, N609, N42);
nand NAND3 (N622, N502, N549, N135);
and AND2 (N623, N621, N373);
buf BUF1 (N624, N618);
nor NOR3 (N625, N619, N44, N543);
xor XOR2 (N626, N614, N415);
or OR3 (N627, N584, N391, N114);
nand NAND4 (N628, N625, N588, N28, N101);
buf BUF1 (N629, N623);
xor XOR2 (N630, N607, N46);
buf BUF1 (N631, N629);
or OR4 (N632, N624, N295, N267, N82);
xor XOR2 (N633, N626, N348);
nand NAND4 (N634, N620, N539, N534, N392);
nor NOR4 (N635, N632, N9, N435, N364);
and AND4 (N636, N633, N616, N450, N466);
buf BUF1 (N637, N617);
and AND3 (N638, N628, N298, N56);
buf BUF1 (N639, N636);
xor XOR2 (N640, N615, N37);
buf BUF1 (N641, N639);
nor NOR2 (N642, N627, N18);
nor NOR2 (N643, N634, N10);
xor XOR2 (N644, N643, N270);
or OR4 (N645, N641, N17, N522, N526);
xor XOR2 (N646, N635, N185);
xor XOR2 (N647, N640, N445);
and AND4 (N648, N622, N420, N362, N248);
buf BUF1 (N649, N646);
buf BUF1 (N650, N647);
buf BUF1 (N651, N650);
buf BUF1 (N652, N642);
buf BUF1 (N653, N630);
nor NOR2 (N654, N631, N136);
and AND3 (N655, N645, N92, N131);
nor NOR4 (N656, N638, N283, N490, N32);
buf BUF1 (N657, N654);
nand NAND2 (N658, N651, N568);
not NOT1 (N659, N648);
or OR4 (N660, N659, N490, N267, N501);
buf BUF1 (N661, N655);
nand NAND3 (N662, N653, N110, N31);
buf BUF1 (N663, N649);
buf BUF1 (N664, N637);
and AND2 (N665, N656, N91);
xor XOR2 (N666, N660, N508);
and AND3 (N667, N666, N372, N228);
and AND2 (N668, N667, N499);
buf BUF1 (N669, N652);
nor NOR2 (N670, N665, N393);
not NOT1 (N671, N662);
buf BUF1 (N672, N671);
nand NAND3 (N673, N669, N290, N606);
xor XOR2 (N674, N668, N304);
buf BUF1 (N675, N673);
nor NOR4 (N676, N657, N616, N283, N495);
xor XOR2 (N677, N644, N168);
or OR4 (N678, N677, N577, N250, N166);
nand NAND4 (N679, N678, N519, N2, N225);
nor NOR2 (N680, N664, N679);
nand NAND3 (N681, N223, N181, N619);
xor XOR2 (N682, N670, N419);
xor XOR2 (N683, N682, N327);
nor NOR4 (N684, N683, N31, N497, N197);
nor NOR4 (N685, N661, N578, N422, N108);
buf BUF1 (N686, N672);
and AND2 (N687, N663, N74);
and AND2 (N688, N658, N603);
or OR4 (N689, N685, N639, N624, N206);
xor XOR2 (N690, N686, N669);
not NOT1 (N691, N687);
nand NAND4 (N692, N681, N651, N463, N114);
or OR3 (N693, N684, N356, N437);
nor NOR3 (N694, N688, N518, N318);
and AND2 (N695, N690, N333);
nand NAND3 (N696, N692, N552, N457);
nand NAND2 (N697, N680, N527);
xor XOR2 (N698, N689, N350);
xor XOR2 (N699, N696, N481);
xor XOR2 (N700, N691, N196);
or OR2 (N701, N674, N267);
nand NAND2 (N702, N676, N671);
not NOT1 (N703, N702);
not NOT1 (N704, N694);
and AND3 (N705, N698, N416, N98);
nor NOR3 (N706, N700, N337, N14);
nand NAND3 (N707, N699, N23, N38);
not NOT1 (N708, N675);
and AND4 (N709, N693, N230, N62, N395);
buf BUF1 (N710, N709);
nor NOR2 (N711, N704, N124);
nor NOR2 (N712, N701, N281);
not NOT1 (N713, N707);
not NOT1 (N714, N705);
xor XOR2 (N715, N695, N40);
buf BUF1 (N716, N708);
or OR3 (N717, N710, N302, N637);
nor NOR2 (N718, N706, N649);
and AND4 (N719, N716, N651, N80, N356);
nand NAND4 (N720, N711, N117, N368, N170);
nor NOR4 (N721, N713, N438, N407, N363);
xor XOR2 (N722, N720, N615);
not NOT1 (N723, N697);
and AND3 (N724, N721, N678, N410);
xor XOR2 (N725, N717, N315);
not NOT1 (N726, N714);
nand NAND2 (N727, N715, N28);
not NOT1 (N728, N723);
or OR3 (N729, N724, N640, N333);
nand NAND2 (N730, N703, N282);
nor NOR4 (N731, N726, N29, N387, N630);
buf BUF1 (N732, N731);
not NOT1 (N733, N725);
nand NAND4 (N734, N712, N727, N30, N328);
not NOT1 (N735, N214);
nand NAND2 (N736, N728, N30);
nand NAND2 (N737, N718, N235);
and AND2 (N738, N722, N472);
nand NAND3 (N739, N729, N74, N507);
buf BUF1 (N740, N736);
xor XOR2 (N741, N735, N85);
xor XOR2 (N742, N737, N541);
or OR2 (N743, N740, N99);
nand NAND3 (N744, N719, N726, N242);
nor NOR3 (N745, N734, N287, N645);
nor NOR4 (N746, N730, N223, N468, N299);
or OR2 (N747, N733, N5);
and AND2 (N748, N747, N67);
or OR3 (N749, N745, N244, N690);
buf BUF1 (N750, N746);
xor XOR2 (N751, N738, N446);
nor NOR4 (N752, N748, N126, N401, N505);
xor XOR2 (N753, N750, N640);
not NOT1 (N754, N749);
xor XOR2 (N755, N742, N94);
and AND2 (N756, N753, N678);
nand NAND4 (N757, N743, N621, N16, N655);
not NOT1 (N758, N751);
nand NAND4 (N759, N757, N613, N430, N418);
nor NOR2 (N760, N744, N401);
xor XOR2 (N761, N752, N536);
buf BUF1 (N762, N756);
nand NAND4 (N763, N739, N130, N229, N577);
nand NAND4 (N764, N763, N238, N621, N107);
and AND3 (N765, N759, N630, N240);
nor NOR3 (N766, N741, N634, N764);
and AND3 (N767, N302, N731, N328);
nand NAND3 (N768, N755, N351, N392);
nand NAND2 (N769, N761, N205);
or OR4 (N770, N769, N312, N261, N117);
buf BUF1 (N771, N732);
nor NOR4 (N772, N762, N630, N327, N10);
xor XOR2 (N773, N771, N213);
and AND2 (N774, N767, N482);
nor NOR3 (N775, N774, N368, N332);
xor XOR2 (N776, N772, N413);
buf BUF1 (N777, N754);
nand NAND3 (N778, N776, N601, N396);
xor XOR2 (N779, N777, N632);
nor NOR4 (N780, N758, N62, N485, N715);
not NOT1 (N781, N770);
xor XOR2 (N782, N781, N102);
nand NAND3 (N783, N775, N427, N420);
nand NAND2 (N784, N783, N653);
and AND3 (N785, N773, N408, N400);
and AND4 (N786, N760, N613, N496, N74);
buf BUF1 (N787, N779);
buf BUF1 (N788, N787);
xor XOR2 (N789, N768, N695);
or OR2 (N790, N778, N180);
and AND3 (N791, N789, N639, N150);
nor NOR4 (N792, N765, N456, N142, N505);
and AND3 (N793, N784, N346, N696);
not NOT1 (N794, N791);
nand NAND4 (N795, N782, N52, N84, N611);
xor XOR2 (N796, N788, N675);
not NOT1 (N797, N785);
and AND3 (N798, N793, N428, N184);
nand NAND4 (N799, N795, N435, N454, N268);
or OR4 (N800, N799, N193, N88, N459);
or OR2 (N801, N798, N471);
not NOT1 (N802, N780);
xor XOR2 (N803, N786, N129);
or OR3 (N804, N797, N267, N509);
not NOT1 (N805, N794);
or OR3 (N806, N805, N12, N557);
not NOT1 (N807, N803);
not NOT1 (N808, N807);
and AND2 (N809, N796, N28);
nor NOR4 (N810, N808, N168, N544, N401);
buf BUF1 (N811, N806);
nand NAND4 (N812, N766, N209, N141, N373);
nand NAND2 (N813, N810, N495);
nand NAND2 (N814, N813, N621);
not NOT1 (N815, N792);
and AND4 (N816, N814, N483, N456, N676);
nor NOR4 (N817, N802, N626, N199, N756);
nor NOR3 (N818, N817, N298, N583);
and AND4 (N819, N790, N198, N103, N83);
nand NAND2 (N820, N811, N41);
xor XOR2 (N821, N815, N16);
buf BUF1 (N822, N800);
not NOT1 (N823, N816);
or OR3 (N824, N812, N478, N107);
nor NOR3 (N825, N819, N82, N606);
or OR3 (N826, N824, N133, N704);
nor NOR4 (N827, N801, N645, N179, N279);
nor NOR2 (N828, N804, N131);
xor XOR2 (N829, N822, N596);
or OR3 (N830, N825, N437, N563);
nand NAND3 (N831, N809, N723, N465);
not NOT1 (N832, N821);
not NOT1 (N833, N831);
xor XOR2 (N834, N826, N47);
xor XOR2 (N835, N820, N787);
and AND3 (N836, N830, N577, N563);
and AND4 (N837, N835, N178, N149, N88);
buf BUF1 (N838, N829);
buf BUF1 (N839, N818);
nor NOR2 (N840, N838, N417);
and AND3 (N841, N837, N554, N365);
xor XOR2 (N842, N828, N47);
not NOT1 (N843, N841);
buf BUF1 (N844, N834);
xor XOR2 (N845, N823, N276);
xor XOR2 (N846, N842, N256);
not NOT1 (N847, N845);
nor NOR2 (N848, N847, N561);
or OR2 (N849, N827, N522);
not NOT1 (N850, N840);
not NOT1 (N851, N832);
or OR4 (N852, N844, N685, N63, N90);
nor NOR2 (N853, N839, N230);
or OR3 (N854, N833, N177, N129);
nand NAND2 (N855, N850, N846);
xor XOR2 (N856, N435, N710);
or OR3 (N857, N855, N766, N301);
nand NAND3 (N858, N857, N124, N458);
nand NAND3 (N859, N848, N545, N438);
and AND4 (N860, N843, N206, N125, N146);
and AND2 (N861, N856, N63);
not NOT1 (N862, N853);
xor XOR2 (N863, N862, N426);
and AND2 (N864, N836, N696);
nand NAND3 (N865, N854, N748, N524);
not NOT1 (N866, N861);
not NOT1 (N867, N851);
nand NAND4 (N868, N852, N195, N834, N224);
nor NOR4 (N869, N849, N622, N821, N807);
or OR2 (N870, N858, N804);
nand NAND2 (N871, N870, N775);
and AND3 (N872, N869, N78, N863);
nor NOR4 (N873, N675, N74, N604, N73);
and AND3 (N874, N865, N593, N497);
and AND4 (N875, N864, N516, N383, N109);
or OR4 (N876, N866, N65, N356, N794);
buf BUF1 (N877, N859);
nand NAND2 (N878, N874, N679);
nor NOR2 (N879, N875, N744);
not NOT1 (N880, N872);
xor XOR2 (N881, N877, N606);
xor XOR2 (N882, N871, N423);
or OR4 (N883, N873, N606, N245, N43);
and AND3 (N884, N881, N183, N292);
or OR2 (N885, N867, N821);
nand NAND4 (N886, N868, N286, N71, N466);
buf BUF1 (N887, N860);
and AND3 (N888, N887, N532, N5);
and AND4 (N889, N885, N170, N495, N824);
buf BUF1 (N890, N882);
not NOT1 (N891, N878);
not NOT1 (N892, N886);
and AND3 (N893, N880, N701, N54);
nand NAND2 (N894, N876, N66);
xor XOR2 (N895, N888, N325);
nor NOR4 (N896, N884, N377, N168, N460);
not NOT1 (N897, N883);
nand NAND4 (N898, N879, N250, N266, N628);
nor NOR4 (N899, N897, N426, N23, N312);
xor XOR2 (N900, N891, N580);
nand NAND3 (N901, N895, N769, N179);
or OR2 (N902, N894, N610);
xor XOR2 (N903, N902, N593);
buf BUF1 (N904, N893);
xor XOR2 (N905, N900, N26);
or OR4 (N906, N903, N848, N902, N634);
nand NAND3 (N907, N896, N690, N296);
nand NAND4 (N908, N905, N484, N873, N314);
or OR2 (N909, N904, N155);
nor NOR2 (N910, N889, N480);
not NOT1 (N911, N909);
or OR4 (N912, N908, N830, N91, N29);
xor XOR2 (N913, N906, N94);
not NOT1 (N914, N898);
or OR2 (N915, N910, N126);
xor XOR2 (N916, N912, N250);
nand NAND3 (N917, N901, N781, N16);
nor NOR4 (N918, N911, N776, N817, N588);
not NOT1 (N919, N913);
xor XOR2 (N920, N917, N264);
buf BUF1 (N921, N920);
buf BUF1 (N922, N915);
nor NOR3 (N923, N921, N590, N122);
nor NOR3 (N924, N907, N399, N917);
xor XOR2 (N925, N890, N592);
xor XOR2 (N926, N924, N50);
nor NOR2 (N927, N916, N407);
not NOT1 (N928, N923);
or OR2 (N929, N925, N785);
nor NOR2 (N930, N892, N81);
nor NOR2 (N931, N928, N597);
buf BUF1 (N932, N918);
buf BUF1 (N933, N922);
not NOT1 (N934, N930);
buf BUF1 (N935, N926);
buf BUF1 (N936, N899);
and AND3 (N937, N927, N844, N547);
nor NOR2 (N938, N932, N371);
and AND2 (N939, N914, N887);
buf BUF1 (N940, N935);
not NOT1 (N941, N933);
buf BUF1 (N942, N937);
nand NAND2 (N943, N934, N499);
and AND2 (N944, N943, N23);
xor XOR2 (N945, N929, N629);
xor XOR2 (N946, N919, N392);
or OR4 (N947, N944, N447, N941, N834);
not NOT1 (N948, N735);
not NOT1 (N949, N940);
nor NOR4 (N950, N931, N167, N662, N128);
nor NOR3 (N951, N947, N432, N226);
xor XOR2 (N952, N951, N413);
not NOT1 (N953, N939);
nand NAND4 (N954, N936, N190, N233, N861);
nor NOR2 (N955, N953, N287);
nor NOR4 (N956, N949, N285, N337, N173);
not NOT1 (N957, N945);
not NOT1 (N958, N955);
not NOT1 (N959, N946);
xor XOR2 (N960, N956, N733);
not NOT1 (N961, N938);
xor XOR2 (N962, N959, N427);
nand NAND2 (N963, N962, N425);
xor XOR2 (N964, N950, N37);
nand NAND4 (N965, N942, N381, N933, N874);
nor NOR4 (N966, N948, N269, N157, N217);
not NOT1 (N967, N954);
xor XOR2 (N968, N958, N451);
and AND2 (N969, N965, N150);
buf BUF1 (N970, N966);
nor NOR2 (N971, N967, N312);
nor NOR3 (N972, N970, N880, N970);
and AND2 (N973, N960, N338);
nand NAND2 (N974, N971, N389);
nor NOR4 (N975, N972, N348, N861, N972);
nor NOR4 (N976, N964, N862, N107, N248);
not NOT1 (N977, N961);
not NOT1 (N978, N975);
and AND3 (N979, N978, N291, N669);
xor XOR2 (N980, N976, N633);
and AND2 (N981, N968, N171);
xor XOR2 (N982, N973, N130);
buf BUF1 (N983, N977);
not NOT1 (N984, N974);
and AND2 (N985, N979, N819);
xor XOR2 (N986, N985, N208);
buf BUF1 (N987, N981);
or OR4 (N988, N983, N827, N798, N930);
not NOT1 (N989, N952);
nand NAND2 (N990, N969, N858);
and AND4 (N991, N990, N166, N740, N514);
nor NOR2 (N992, N984, N801);
and AND3 (N993, N989, N194, N685);
buf BUF1 (N994, N957);
nand NAND2 (N995, N991, N712);
nor NOR2 (N996, N963, N579);
not NOT1 (N997, N987);
buf BUF1 (N998, N995);
xor XOR2 (N999, N988, N850);
nor NOR3 (N1000, N980, N666, N758);
not NOT1 (N1001, N999);
buf BUF1 (N1002, N996);
nand NAND3 (N1003, N993, N883, N359);
and AND2 (N1004, N994, N907);
xor XOR2 (N1005, N998, N346);
buf BUF1 (N1006, N986);
xor XOR2 (N1007, N1005, N29);
xor XOR2 (N1008, N1000, N974);
or OR4 (N1009, N992, N990, N357, N468);
nor NOR4 (N1010, N1002, N12, N505, N293);
not NOT1 (N1011, N1001);
and AND3 (N1012, N997, N857, N890);
not NOT1 (N1013, N1003);
and AND3 (N1014, N1009, N141, N748);
or OR2 (N1015, N1010, N101);
xor XOR2 (N1016, N1004, N921);
or OR2 (N1017, N1008, N794);
and AND2 (N1018, N1007, N106);
nor NOR3 (N1019, N1006, N176, N984);
xor XOR2 (N1020, N1015, N976);
and AND3 (N1021, N982, N285, N905);
or OR2 (N1022, N1017, N372);
nand NAND3 (N1023, N1016, N165, N981);
buf BUF1 (N1024, N1014);
buf BUF1 (N1025, N1022);
nor NOR4 (N1026, N1024, N617, N346, N349);
and AND3 (N1027, N1018, N54, N23);
buf BUF1 (N1028, N1011);
and AND4 (N1029, N1012, N621, N506, N777);
buf BUF1 (N1030, N1029);
buf BUF1 (N1031, N1023);
or OR2 (N1032, N1028, N597);
or OR4 (N1033, N1026, N217, N530, N558);
not NOT1 (N1034, N1030);
buf BUF1 (N1035, N1019);
buf BUF1 (N1036, N1034);
and AND2 (N1037, N1032, N13);
buf BUF1 (N1038, N1027);
or OR3 (N1039, N1038, N230, N288);
or OR2 (N1040, N1021, N490);
buf BUF1 (N1041, N1037);
nor NOR2 (N1042, N1013, N8);
or OR4 (N1043, N1031, N292, N982, N603);
nor NOR3 (N1044, N1040, N481, N158);
buf BUF1 (N1045, N1041);
not NOT1 (N1046, N1045);
and AND3 (N1047, N1043, N553, N133);
not NOT1 (N1048, N1020);
nor NOR3 (N1049, N1046, N228, N901);
xor XOR2 (N1050, N1049, N1030);
nor NOR3 (N1051, N1025, N49, N624);
buf BUF1 (N1052, N1042);
nand NAND4 (N1053, N1035, N345, N836, N551);
nor NOR2 (N1054, N1053, N941);
not NOT1 (N1055, N1052);
and AND3 (N1056, N1054, N831, N568);
not NOT1 (N1057, N1051);
or OR2 (N1058, N1044, N364);
nand NAND4 (N1059, N1055, N361, N714, N767);
buf BUF1 (N1060, N1047);
nand NAND3 (N1061, N1039, N378, N242);
and AND3 (N1062, N1059, N142, N592);
buf BUF1 (N1063, N1056);
buf BUF1 (N1064, N1060);
nand NAND4 (N1065, N1062, N899, N421, N177);
and AND3 (N1066, N1058, N1039, N126);
xor XOR2 (N1067, N1061, N447);
nor NOR3 (N1068, N1063, N839, N825);
and AND2 (N1069, N1033, N696);
xor XOR2 (N1070, N1057, N165);
xor XOR2 (N1071, N1070, N380);
or OR2 (N1072, N1071, N409);
nand NAND4 (N1073, N1066, N720, N109, N606);
not NOT1 (N1074, N1067);
and AND2 (N1075, N1074, N113);
or OR4 (N1076, N1050, N483, N105, N540);
xor XOR2 (N1077, N1065, N327);
and AND2 (N1078, N1077, N1076);
xor XOR2 (N1079, N805, N691);
nor NOR2 (N1080, N1075, N304);
nand NAND2 (N1081, N1078, N611);
nand NAND4 (N1082, N1064, N258, N613, N486);
nand NAND3 (N1083, N1082, N229, N665);
buf BUF1 (N1084, N1068);
not NOT1 (N1085, N1072);
nor NOR3 (N1086, N1081, N483, N852);
xor XOR2 (N1087, N1083, N427);
not NOT1 (N1088, N1080);
not NOT1 (N1089, N1087);
nand NAND3 (N1090, N1073, N73, N428);
or OR4 (N1091, N1090, N760, N624, N299);
buf BUF1 (N1092, N1085);
and AND2 (N1093, N1036, N266);
xor XOR2 (N1094, N1086, N1009);
and AND2 (N1095, N1092, N349);
xor XOR2 (N1096, N1093, N825);
or OR3 (N1097, N1084, N327, N537);
nand NAND4 (N1098, N1069, N99, N692, N717);
or OR2 (N1099, N1091, N164);
xor XOR2 (N1100, N1048, N368);
nand NAND4 (N1101, N1088, N232, N611, N962);
xor XOR2 (N1102, N1094, N149);
nor NOR4 (N1103, N1100, N1028, N410, N657);
nor NOR4 (N1104, N1096, N150, N330, N524);
nand NAND2 (N1105, N1101, N114);
or OR4 (N1106, N1095, N804, N1035, N1082);
or OR2 (N1107, N1104, N760);
buf BUF1 (N1108, N1099);
xor XOR2 (N1109, N1098, N526);
or OR3 (N1110, N1106, N887, N923);
buf BUF1 (N1111, N1103);
not NOT1 (N1112, N1110);
nor NOR3 (N1113, N1105, N892, N322);
xor XOR2 (N1114, N1107, N1035);
and AND2 (N1115, N1102, N6);
nand NAND2 (N1116, N1089, N417);
and AND3 (N1117, N1114, N765, N749);
nand NAND2 (N1118, N1108, N1021);
not NOT1 (N1119, N1118);
nor NOR2 (N1120, N1116, N907);
buf BUF1 (N1121, N1113);
not NOT1 (N1122, N1097);
nor NOR3 (N1123, N1119, N797, N79);
nand NAND2 (N1124, N1121, N894);
not NOT1 (N1125, N1111);
buf BUF1 (N1126, N1109);
not NOT1 (N1127, N1124);
and AND4 (N1128, N1123, N1111, N363, N131);
nor NOR4 (N1129, N1128, N1114, N933, N370);
and AND3 (N1130, N1125, N84, N569);
and AND2 (N1131, N1112, N1011);
and AND4 (N1132, N1115, N554, N181, N403);
xor XOR2 (N1133, N1129, N514);
buf BUF1 (N1134, N1133);
nand NAND2 (N1135, N1117, N1134);
not NOT1 (N1136, N712);
not NOT1 (N1137, N1132);
not NOT1 (N1138, N1130);
nand NAND4 (N1139, N1137, N969, N896, N1016);
xor XOR2 (N1140, N1135, N208);
buf BUF1 (N1141, N1139);
and AND3 (N1142, N1131, N473, N729);
buf BUF1 (N1143, N1127);
or OR4 (N1144, N1122, N929, N1099, N563);
and AND3 (N1145, N1140, N287, N733);
nand NAND4 (N1146, N1138, N680, N383, N756);
nor NOR2 (N1147, N1144, N785);
not NOT1 (N1148, N1079);
nor NOR3 (N1149, N1147, N589, N237);
and AND2 (N1150, N1146, N507);
nor NOR3 (N1151, N1149, N938, N923);
or OR3 (N1152, N1150, N597, N183);
nor NOR4 (N1153, N1152, N94, N464, N863);
nor NOR3 (N1154, N1136, N261, N77);
or OR4 (N1155, N1151, N767, N442, N1035);
or OR4 (N1156, N1142, N116, N312, N1015);
xor XOR2 (N1157, N1143, N306);
buf BUF1 (N1158, N1145);
buf BUF1 (N1159, N1120);
and AND2 (N1160, N1154, N204);
xor XOR2 (N1161, N1160, N167);
and AND4 (N1162, N1157, N806, N909, N306);
not NOT1 (N1163, N1161);
or OR3 (N1164, N1156, N1080, N702);
and AND3 (N1165, N1126, N303, N127);
or OR2 (N1166, N1159, N80);
or OR2 (N1167, N1141, N380);
buf BUF1 (N1168, N1153);
xor XOR2 (N1169, N1164, N264);
not NOT1 (N1170, N1166);
nor NOR4 (N1171, N1168, N916, N66, N1069);
xor XOR2 (N1172, N1171, N175);
nand NAND4 (N1173, N1163, N543, N125, N1080);
not NOT1 (N1174, N1170);
nor NOR3 (N1175, N1174, N246, N796);
xor XOR2 (N1176, N1155, N542);
nor NOR3 (N1177, N1172, N139, N360);
nor NOR2 (N1178, N1167, N933);
buf BUF1 (N1179, N1175);
not NOT1 (N1180, N1162);
nor NOR4 (N1181, N1180, N196, N751, N672);
buf BUF1 (N1182, N1176);
nor NOR4 (N1183, N1179, N389, N433, N49);
nand NAND3 (N1184, N1148, N494, N513);
nand NAND4 (N1185, N1169, N628, N451, N62);
not NOT1 (N1186, N1182);
and AND4 (N1187, N1184, N1154, N730, N875);
nand NAND3 (N1188, N1158, N1101, N184);
and AND3 (N1189, N1185, N959, N877);
and AND3 (N1190, N1188, N844, N1155);
nand NAND3 (N1191, N1187, N466, N446);
xor XOR2 (N1192, N1189, N232);
not NOT1 (N1193, N1177);
not NOT1 (N1194, N1165);
buf BUF1 (N1195, N1181);
nand NAND2 (N1196, N1173, N974);
buf BUF1 (N1197, N1192);
or OR2 (N1198, N1190, N500);
nor NOR3 (N1199, N1191, N45, N1024);
nand NAND3 (N1200, N1194, N558, N114);
xor XOR2 (N1201, N1198, N305);
xor XOR2 (N1202, N1196, N1057);
or OR3 (N1203, N1199, N605, N1187);
and AND2 (N1204, N1201, N319);
nor NOR2 (N1205, N1204, N717);
xor XOR2 (N1206, N1193, N254);
xor XOR2 (N1207, N1205, N226);
nand NAND4 (N1208, N1206, N190, N425, N682);
and AND4 (N1209, N1195, N1136, N298, N428);
nor NOR2 (N1210, N1200, N336);
nand NAND3 (N1211, N1203, N450, N405);
nor NOR3 (N1212, N1209, N157, N733);
nor NOR4 (N1213, N1202, N536, N836, N476);
nand NAND3 (N1214, N1210, N50, N85);
and AND2 (N1215, N1207, N776);
and AND4 (N1216, N1215, N666, N736, N193);
nor NOR2 (N1217, N1213, N414);
xor XOR2 (N1218, N1208, N575);
nand NAND3 (N1219, N1214, N379, N891);
not NOT1 (N1220, N1178);
nand NAND2 (N1221, N1217, N1053);
and AND4 (N1222, N1219, N966, N982, N558);
nand NAND3 (N1223, N1222, N427, N1142);
nor NOR2 (N1224, N1197, N593);
xor XOR2 (N1225, N1221, N403);
and AND2 (N1226, N1186, N614);
xor XOR2 (N1227, N1224, N250);
nor NOR2 (N1228, N1225, N887);
not NOT1 (N1229, N1211);
and AND4 (N1230, N1229, N528, N1016, N626);
nand NAND3 (N1231, N1230, N428, N527);
or OR4 (N1232, N1218, N795, N906, N1224);
nand NAND3 (N1233, N1220, N1189, N74);
nor NOR3 (N1234, N1226, N476, N1105);
buf BUF1 (N1235, N1231);
or OR3 (N1236, N1233, N170, N388);
not NOT1 (N1237, N1216);
or OR2 (N1238, N1227, N913);
or OR3 (N1239, N1232, N86, N782);
xor XOR2 (N1240, N1236, N478);
nand NAND3 (N1241, N1237, N378, N215);
or OR4 (N1242, N1234, N969, N76, N120);
not NOT1 (N1243, N1238);
and AND2 (N1244, N1223, N652);
not NOT1 (N1245, N1243);
nor NOR2 (N1246, N1245, N124);
or OR4 (N1247, N1228, N437, N422, N101);
not NOT1 (N1248, N1212);
xor XOR2 (N1249, N1241, N1065);
xor XOR2 (N1250, N1183, N634);
nor NOR2 (N1251, N1248, N1045);
nor NOR2 (N1252, N1244, N954);
xor XOR2 (N1253, N1247, N639);
not NOT1 (N1254, N1250);
not NOT1 (N1255, N1254);
buf BUF1 (N1256, N1242);
and AND3 (N1257, N1253, N911, N89);
nand NAND2 (N1258, N1251, N909);
or OR2 (N1259, N1252, N93);
not NOT1 (N1260, N1240);
not NOT1 (N1261, N1255);
xor XOR2 (N1262, N1261, N1258);
xor XOR2 (N1263, N672, N53);
buf BUF1 (N1264, N1263);
or OR2 (N1265, N1264, N673);
nand NAND3 (N1266, N1235, N1160, N517);
or OR4 (N1267, N1246, N1037, N163, N786);
xor XOR2 (N1268, N1265, N800);
xor XOR2 (N1269, N1267, N414);
or OR2 (N1270, N1249, N238);
not NOT1 (N1271, N1270);
and AND2 (N1272, N1260, N1151);
xor XOR2 (N1273, N1271, N721);
not NOT1 (N1274, N1269);
nor NOR4 (N1275, N1274, N137, N446, N575);
and AND2 (N1276, N1262, N1160);
nand NAND3 (N1277, N1272, N522, N47);
nor NOR3 (N1278, N1273, N159, N639);
not NOT1 (N1279, N1259);
nand NAND3 (N1280, N1257, N303, N1160);
and AND2 (N1281, N1275, N667);
not NOT1 (N1282, N1279);
nand NAND3 (N1283, N1266, N584, N705);
nand NAND4 (N1284, N1278, N1208, N239, N1162);
buf BUF1 (N1285, N1276);
nand NAND2 (N1286, N1283, N172);
buf BUF1 (N1287, N1281);
not NOT1 (N1288, N1277);
nand NAND2 (N1289, N1287, N1222);
nand NAND3 (N1290, N1289, N563, N856);
nand NAND3 (N1291, N1288, N392, N557);
not NOT1 (N1292, N1286);
xor XOR2 (N1293, N1291, N958);
buf BUF1 (N1294, N1256);
xor XOR2 (N1295, N1239, N568);
not NOT1 (N1296, N1295);
buf BUF1 (N1297, N1285);
and AND3 (N1298, N1293, N927, N342);
and AND4 (N1299, N1296, N101, N877, N449);
nor NOR4 (N1300, N1290, N886, N502, N988);
nor NOR4 (N1301, N1298, N1058, N653, N328);
not NOT1 (N1302, N1268);
not NOT1 (N1303, N1297);
nand NAND3 (N1304, N1294, N467, N553);
not NOT1 (N1305, N1304);
and AND4 (N1306, N1280, N1147, N356, N576);
buf BUF1 (N1307, N1301);
xor XOR2 (N1308, N1292, N1167);
nand NAND3 (N1309, N1305, N155, N214);
not NOT1 (N1310, N1308);
and AND3 (N1311, N1303, N875, N998);
not NOT1 (N1312, N1310);
nor NOR3 (N1313, N1306, N538, N258);
nand NAND2 (N1314, N1299, N1048);
or OR2 (N1315, N1307, N776);
not NOT1 (N1316, N1302);
xor XOR2 (N1317, N1282, N1123);
and AND4 (N1318, N1317, N957, N379, N126);
buf BUF1 (N1319, N1318);
xor XOR2 (N1320, N1319, N238);
or OR2 (N1321, N1316, N1199);
or OR4 (N1322, N1313, N478, N919, N622);
and AND2 (N1323, N1315, N621);
not NOT1 (N1324, N1314);
nand NAND4 (N1325, N1309, N28, N737, N649);
xor XOR2 (N1326, N1312, N1061);
xor XOR2 (N1327, N1324, N1288);
not NOT1 (N1328, N1325);
nand NAND4 (N1329, N1322, N938, N709, N1228);
nor NOR2 (N1330, N1311, N1141);
and AND4 (N1331, N1284, N22, N461, N207);
xor XOR2 (N1332, N1331, N200);
or OR4 (N1333, N1332, N1190, N6, N1169);
or OR4 (N1334, N1333, N906, N1182, N711);
or OR4 (N1335, N1328, N116, N1287, N1049);
nor NOR2 (N1336, N1334, N930);
nand NAND2 (N1337, N1335, N514);
or OR3 (N1338, N1321, N1268, N445);
nor NOR4 (N1339, N1327, N379, N1257, N1124);
nor NOR3 (N1340, N1329, N439, N358);
nand NAND2 (N1341, N1337, N1327);
nor NOR3 (N1342, N1323, N242, N1066);
xor XOR2 (N1343, N1340, N625);
nand NAND3 (N1344, N1343, N1140, N1170);
xor XOR2 (N1345, N1330, N343);
nor NOR4 (N1346, N1345, N303, N824, N592);
or OR4 (N1347, N1339, N599, N1216, N1248);
and AND3 (N1348, N1346, N326, N218);
xor XOR2 (N1349, N1348, N1237);
and AND3 (N1350, N1338, N1145, N634);
or OR4 (N1351, N1320, N980, N1216, N156);
nor NOR2 (N1352, N1351, N471);
nand NAND2 (N1353, N1336, N572);
not NOT1 (N1354, N1326);
xor XOR2 (N1355, N1352, N1311);
or OR2 (N1356, N1354, N352);
nor NOR3 (N1357, N1300, N105, N310);
buf BUF1 (N1358, N1342);
nand NAND2 (N1359, N1356, N1183);
and AND3 (N1360, N1341, N52, N288);
and AND4 (N1361, N1349, N1083, N824, N376);
buf BUF1 (N1362, N1357);
not NOT1 (N1363, N1355);
or OR3 (N1364, N1362, N609, N851);
not NOT1 (N1365, N1361);
and AND3 (N1366, N1358, N1223, N79);
and AND2 (N1367, N1363, N1106);
not NOT1 (N1368, N1350);
and AND4 (N1369, N1364, N332, N652, N1042);
or OR3 (N1370, N1366, N176, N956);
xor XOR2 (N1371, N1370, N743);
xor XOR2 (N1372, N1347, N1112);
buf BUF1 (N1373, N1371);
or OR4 (N1374, N1360, N234, N685, N1126);
and AND2 (N1375, N1344, N69);
xor XOR2 (N1376, N1374, N850);
not NOT1 (N1377, N1368);
buf BUF1 (N1378, N1365);
nand NAND3 (N1379, N1375, N1251, N652);
xor XOR2 (N1380, N1353, N421);
xor XOR2 (N1381, N1373, N847);
nand NAND4 (N1382, N1367, N254, N471, N148);
and AND2 (N1383, N1379, N291);
not NOT1 (N1384, N1377);
xor XOR2 (N1385, N1376, N911);
or OR2 (N1386, N1359, N487);
not NOT1 (N1387, N1385);
xor XOR2 (N1388, N1382, N896);
and AND2 (N1389, N1380, N784);
and AND4 (N1390, N1388, N182, N1340, N399);
buf BUF1 (N1391, N1372);
and AND2 (N1392, N1384, N25);
nand NAND2 (N1393, N1369, N1312);
nand NAND4 (N1394, N1391, N633, N720, N1166);
and AND3 (N1395, N1393, N1164, N1195);
xor XOR2 (N1396, N1390, N953);
xor XOR2 (N1397, N1394, N272);
nor NOR3 (N1398, N1383, N892, N1238);
nand NAND4 (N1399, N1398, N622, N932, N500);
buf BUF1 (N1400, N1386);
buf BUF1 (N1401, N1392);
or OR2 (N1402, N1378, N283);
xor XOR2 (N1403, N1387, N677);
nand NAND4 (N1404, N1395, N1222, N1318, N959);
nor NOR4 (N1405, N1403, N564, N997, N644);
buf BUF1 (N1406, N1389);
nand NAND4 (N1407, N1402, N673, N1041, N642);
xor XOR2 (N1408, N1396, N924);
xor XOR2 (N1409, N1397, N660);
nand NAND2 (N1410, N1405, N1128);
nand NAND3 (N1411, N1381, N1397, N122);
nor NOR4 (N1412, N1399, N1350, N668, N257);
nor NOR4 (N1413, N1410, N433, N1239, N994);
xor XOR2 (N1414, N1408, N221);
buf BUF1 (N1415, N1411);
nand NAND4 (N1416, N1414, N115, N16, N397);
or OR2 (N1417, N1406, N547);
not NOT1 (N1418, N1412);
buf BUF1 (N1419, N1418);
or OR3 (N1420, N1400, N521, N958);
and AND4 (N1421, N1404, N554, N1117, N221);
nand NAND3 (N1422, N1421, N557, N522);
nand NAND3 (N1423, N1409, N377, N375);
nand NAND2 (N1424, N1420, N1017);
and AND2 (N1425, N1407, N68);
or OR3 (N1426, N1415, N408, N1007);
xor XOR2 (N1427, N1423, N726);
nor NOR4 (N1428, N1422, N1025, N1070, N1239);
not NOT1 (N1429, N1428);
or OR2 (N1430, N1416, N400);
nand NAND3 (N1431, N1401, N1031, N790);
xor XOR2 (N1432, N1424, N345);
buf BUF1 (N1433, N1429);
or OR2 (N1434, N1427, N335);
nand NAND2 (N1435, N1413, N593);
or OR4 (N1436, N1419, N58, N876, N166);
and AND3 (N1437, N1432, N326, N965);
not NOT1 (N1438, N1425);
or OR4 (N1439, N1435, N1186, N753, N128);
xor XOR2 (N1440, N1426, N480);
nor NOR4 (N1441, N1438, N1434, N1188, N62);
nor NOR4 (N1442, N1361, N1425, N1349, N839);
xor XOR2 (N1443, N1417, N1333);
nand NAND4 (N1444, N1431, N615, N1070, N389);
nand NAND2 (N1445, N1437, N651);
nand NAND3 (N1446, N1440, N370, N1196);
and AND4 (N1447, N1443, N636, N700, N49);
buf BUF1 (N1448, N1445);
or OR2 (N1449, N1448, N498);
nand NAND2 (N1450, N1449, N534);
and AND4 (N1451, N1444, N1131, N1441, N1244);
or OR3 (N1452, N466, N1087, N828);
or OR2 (N1453, N1442, N1202);
nand NAND4 (N1454, N1452, N1084, N232, N1261);
nand NAND3 (N1455, N1446, N872, N284);
nand NAND4 (N1456, N1436, N561, N241, N1035);
xor XOR2 (N1457, N1430, N723);
and AND2 (N1458, N1455, N1409);
not NOT1 (N1459, N1458);
xor XOR2 (N1460, N1457, N11);
buf BUF1 (N1461, N1450);
and AND2 (N1462, N1456, N545);
and AND2 (N1463, N1459, N687);
nor NOR3 (N1464, N1447, N1312, N485);
xor XOR2 (N1465, N1451, N462);
or OR2 (N1466, N1439, N770);
nor NOR4 (N1467, N1466, N232, N653, N598);
xor XOR2 (N1468, N1462, N181);
xor XOR2 (N1469, N1454, N714);
or OR3 (N1470, N1467, N337, N631);
buf BUF1 (N1471, N1464);
and AND4 (N1472, N1465, N363, N860, N31);
and AND3 (N1473, N1433, N1338, N1227);
xor XOR2 (N1474, N1471, N330);
and AND2 (N1475, N1470, N630);
nand NAND2 (N1476, N1461, N409);
xor XOR2 (N1477, N1476, N954);
buf BUF1 (N1478, N1472);
nor NOR4 (N1479, N1453, N1369, N1429, N62);
nand NAND4 (N1480, N1460, N1001, N1048, N856);
nand NAND2 (N1481, N1477, N831);
nand NAND3 (N1482, N1469, N101, N1412);
xor XOR2 (N1483, N1478, N960);
nand NAND2 (N1484, N1473, N1482);
and AND3 (N1485, N433, N1364, N1353);
or OR4 (N1486, N1475, N674, N1371, N960);
nor NOR2 (N1487, N1483, N101);
nor NOR3 (N1488, N1468, N143, N355);
xor XOR2 (N1489, N1474, N1034);
buf BUF1 (N1490, N1480);
buf BUF1 (N1491, N1485);
or OR4 (N1492, N1487, N189, N147, N266);
and AND4 (N1493, N1488, N1149, N104, N330);
buf BUF1 (N1494, N1492);
not NOT1 (N1495, N1490);
nand NAND3 (N1496, N1481, N1083, N840);
and AND4 (N1497, N1494, N758, N1052, N1152);
and AND3 (N1498, N1463, N92, N1196);
or OR3 (N1499, N1497, N327, N662);
or OR2 (N1500, N1484, N481);
buf BUF1 (N1501, N1499);
or OR3 (N1502, N1491, N752, N1355);
nor NOR4 (N1503, N1502, N85, N1253, N906);
not NOT1 (N1504, N1479);
buf BUF1 (N1505, N1504);
buf BUF1 (N1506, N1501);
and AND4 (N1507, N1493, N133, N178, N361);
or OR2 (N1508, N1489, N199);
and AND2 (N1509, N1486, N224);
and AND2 (N1510, N1506, N1050);
nand NAND4 (N1511, N1510, N1131, N1223, N1161);
xor XOR2 (N1512, N1511, N363);
nor NOR4 (N1513, N1495, N291, N594, N1207);
not NOT1 (N1514, N1512);
xor XOR2 (N1515, N1513, N1136);
nand NAND3 (N1516, N1498, N1397, N679);
or OR2 (N1517, N1515, N1026);
nor NOR3 (N1518, N1516, N75, N780);
not NOT1 (N1519, N1514);
nand NAND2 (N1520, N1505, N1271);
xor XOR2 (N1521, N1519, N845);
nor NOR4 (N1522, N1508, N1226, N1097, N1283);
xor XOR2 (N1523, N1518, N1082);
and AND2 (N1524, N1503, N284);
buf BUF1 (N1525, N1521);
nand NAND4 (N1526, N1496, N1380, N364, N612);
nand NAND3 (N1527, N1517, N1123, N133);
buf BUF1 (N1528, N1520);
nor NOR4 (N1529, N1525, N218, N545, N685);
and AND2 (N1530, N1523, N1426);
nor NOR3 (N1531, N1527, N716, N590);
not NOT1 (N1532, N1524);
and AND3 (N1533, N1500, N1138, N298);
or OR3 (N1534, N1507, N1280, N75);
nor NOR3 (N1535, N1522, N765, N799);
or OR2 (N1536, N1529, N651);
buf BUF1 (N1537, N1509);
not NOT1 (N1538, N1535);
buf BUF1 (N1539, N1526);
and AND2 (N1540, N1531, N330);
not NOT1 (N1541, N1537);
buf BUF1 (N1542, N1532);
nor NOR4 (N1543, N1536, N1510, N839, N47);
not NOT1 (N1544, N1538);
nand NAND2 (N1545, N1544, N168);
xor XOR2 (N1546, N1543, N12);
nand NAND2 (N1547, N1539, N779);
nor NOR3 (N1548, N1542, N378, N7);
not NOT1 (N1549, N1545);
or OR3 (N1550, N1540, N1510, N312);
or OR2 (N1551, N1546, N1513);
nand NAND3 (N1552, N1551, N68, N1442);
nand NAND4 (N1553, N1530, N1088, N264, N659);
nand NAND3 (N1554, N1550, N963, N593);
or OR3 (N1555, N1541, N1440, N184);
and AND3 (N1556, N1528, N499, N1427);
nand NAND4 (N1557, N1555, N1048, N220, N342);
nand NAND3 (N1558, N1557, N1034, N75);
and AND4 (N1559, N1534, N1503, N523, N55);
nand NAND2 (N1560, N1554, N720);
and AND4 (N1561, N1549, N481, N73, N531);
nor NOR4 (N1562, N1561, N1339, N116, N756);
nor NOR4 (N1563, N1547, N151, N595, N308);
nand NAND3 (N1564, N1563, N465, N196);
not NOT1 (N1565, N1548);
nand NAND2 (N1566, N1565, N1534);
buf BUF1 (N1567, N1566);
nor NOR3 (N1568, N1564, N974, N955);
buf BUF1 (N1569, N1552);
nand NAND3 (N1570, N1568, N734, N869);
or OR4 (N1571, N1533, N354, N1283, N1221);
buf BUF1 (N1572, N1556);
not NOT1 (N1573, N1562);
nand NAND4 (N1574, N1560, N1279, N1360, N968);
not NOT1 (N1575, N1567);
and AND2 (N1576, N1553, N925);
and AND4 (N1577, N1569, N571, N1394, N676);
and AND4 (N1578, N1574, N453, N187, N240);
xor XOR2 (N1579, N1575, N333);
nand NAND3 (N1580, N1573, N1549, N668);
or OR3 (N1581, N1570, N1079, N1164);
nor NOR4 (N1582, N1559, N1348, N647, N811);
not NOT1 (N1583, N1576);
nor NOR2 (N1584, N1581, N179);
nor NOR4 (N1585, N1584, N716, N227, N165);
nand NAND2 (N1586, N1571, N1301);
nor NOR3 (N1587, N1583, N978, N1230);
buf BUF1 (N1588, N1587);
nor NOR2 (N1589, N1577, N967);
xor XOR2 (N1590, N1585, N1058);
or OR3 (N1591, N1589, N717, N158);
nand NAND3 (N1592, N1579, N33, N593);
buf BUF1 (N1593, N1578);
nor NOR4 (N1594, N1580, N556, N100, N1021);
buf BUF1 (N1595, N1558);
nand NAND4 (N1596, N1572, N1530, N237, N1153);
and AND2 (N1597, N1590, N1046);
nor NOR4 (N1598, N1597, N322, N1260, N143);
not NOT1 (N1599, N1596);
and AND2 (N1600, N1592, N744);
nor NOR2 (N1601, N1586, N439);
xor XOR2 (N1602, N1599, N828);
or OR2 (N1603, N1582, N1170);
nor NOR2 (N1604, N1588, N853);
or OR3 (N1605, N1593, N238, N1539);
nand NAND4 (N1606, N1603, N687, N500, N375);
or OR3 (N1607, N1600, N576, N1558);
nor NOR4 (N1608, N1605, N1099, N1318, N1510);
nor NOR2 (N1609, N1602, N1045);
xor XOR2 (N1610, N1609, N1266);
or OR4 (N1611, N1591, N866, N1239, N416);
or OR2 (N1612, N1607, N718);
not NOT1 (N1613, N1610);
and AND2 (N1614, N1604, N577);
or OR4 (N1615, N1613, N5, N1163, N156);
or OR2 (N1616, N1615, N1096);
nor NOR4 (N1617, N1606, N993, N797, N440);
not NOT1 (N1618, N1611);
nand NAND4 (N1619, N1614, N1040, N897, N106);
nand NAND3 (N1620, N1601, N1483, N501);
nand NAND2 (N1621, N1620, N1234);
buf BUF1 (N1622, N1617);
nor NOR3 (N1623, N1594, N1531, N1517);
not NOT1 (N1624, N1622);
nand NAND3 (N1625, N1621, N1275, N446);
buf BUF1 (N1626, N1608);
xor XOR2 (N1627, N1616, N1007);
or OR4 (N1628, N1624, N1515, N759, N1467);
not NOT1 (N1629, N1627);
nand NAND4 (N1630, N1629, N1574, N1227, N261);
or OR4 (N1631, N1598, N517, N1041, N730);
or OR2 (N1632, N1625, N1340);
buf BUF1 (N1633, N1631);
nor NOR4 (N1634, N1612, N195, N812, N1264);
not NOT1 (N1635, N1618);
xor XOR2 (N1636, N1623, N990);
and AND4 (N1637, N1595, N1077, N668, N149);
buf BUF1 (N1638, N1637);
or OR3 (N1639, N1635, N1112, N1014);
nand NAND4 (N1640, N1628, N1034, N1407, N473);
nor NOR2 (N1641, N1636, N713);
not NOT1 (N1642, N1634);
xor XOR2 (N1643, N1632, N442);
and AND3 (N1644, N1643, N471, N1186);
or OR4 (N1645, N1630, N1611, N581, N327);
or OR3 (N1646, N1641, N42, N1338);
or OR3 (N1647, N1642, N962, N1412);
nand NAND4 (N1648, N1645, N1564, N1497, N566);
buf BUF1 (N1649, N1640);
buf BUF1 (N1650, N1619);
nand NAND3 (N1651, N1638, N333, N14);
or OR3 (N1652, N1626, N1531, N1417);
nor NOR4 (N1653, N1644, N768, N63, N289);
and AND3 (N1654, N1649, N41, N1125);
not NOT1 (N1655, N1651);
not NOT1 (N1656, N1652);
or OR3 (N1657, N1655, N1072, N683);
not NOT1 (N1658, N1657);
or OR2 (N1659, N1647, N734);
buf BUF1 (N1660, N1650);
buf BUF1 (N1661, N1658);
xor XOR2 (N1662, N1660, N750);
nor NOR3 (N1663, N1653, N1548, N785);
xor XOR2 (N1664, N1659, N1139);
and AND2 (N1665, N1654, N1617);
not NOT1 (N1666, N1648);
xor XOR2 (N1667, N1664, N169);
or OR2 (N1668, N1667, N954);
nand NAND4 (N1669, N1666, N945, N922, N1375);
xor XOR2 (N1670, N1662, N160);
xor XOR2 (N1671, N1633, N41);
and AND4 (N1672, N1646, N1082, N1252, N1503);
nand NAND3 (N1673, N1670, N311, N511);
or OR3 (N1674, N1668, N305, N1353);
buf BUF1 (N1675, N1656);
xor XOR2 (N1676, N1661, N1368);
xor XOR2 (N1677, N1671, N949);
buf BUF1 (N1678, N1669);
nand NAND4 (N1679, N1678, N356, N1332, N1129);
buf BUF1 (N1680, N1672);
nand NAND3 (N1681, N1677, N1533, N710);
buf BUF1 (N1682, N1639);
nand NAND3 (N1683, N1682, N182, N87);
buf BUF1 (N1684, N1665);
xor XOR2 (N1685, N1675, N384);
not NOT1 (N1686, N1663);
nand NAND2 (N1687, N1679, N336);
or OR2 (N1688, N1673, N519);
or OR2 (N1689, N1676, N879);
nor NOR4 (N1690, N1689, N1513, N449, N1222);
or OR3 (N1691, N1683, N335, N1168);
nor NOR3 (N1692, N1690, N494, N1128);
xor XOR2 (N1693, N1674, N855);
nand NAND2 (N1694, N1692, N901);
not NOT1 (N1695, N1688);
nand NAND4 (N1696, N1686, N1159, N703, N880);
and AND3 (N1697, N1680, N93, N76);
buf BUF1 (N1698, N1695);
nand NAND3 (N1699, N1693, N1500, N1155);
not NOT1 (N1700, N1698);
nand NAND4 (N1701, N1696, N320, N1402, N428);
or OR4 (N1702, N1700, N1375, N1266, N1618);
or OR4 (N1703, N1681, N978, N1088, N339);
not NOT1 (N1704, N1702);
or OR2 (N1705, N1694, N656);
or OR3 (N1706, N1691, N1229, N101);
or OR2 (N1707, N1706, N1696);
or OR2 (N1708, N1699, N1193);
nand NAND2 (N1709, N1708, N491);
buf BUF1 (N1710, N1684);
buf BUF1 (N1711, N1709);
buf BUF1 (N1712, N1697);
not NOT1 (N1713, N1710);
and AND4 (N1714, N1685, N1191, N532, N1511);
xor XOR2 (N1715, N1713, N311);
buf BUF1 (N1716, N1711);
xor XOR2 (N1717, N1687, N228);
xor XOR2 (N1718, N1703, N1583);
nor NOR4 (N1719, N1707, N266, N839, N345);
not NOT1 (N1720, N1719);
and AND4 (N1721, N1718, N1508, N585, N1088);
xor XOR2 (N1722, N1705, N1364);
xor XOR2 (N1723, N1715, N834);
xor XOR2 (N1724, N1704, N599);
nor NOR4 (N1725, N1723, N1723, N250, N1059);
xor XOR2 (N1726, N1716, N1552);
nand NAND4 (N1727, N1721, N1243, N875, N81);
xor XOR2 (N1728, N1722, N212);
buf BUF1 (N1729, N1726);
not NOT1 (N1730, N1714);
nand NAND2 (N1731, N1717, N422);
nand NAND2 (N1732, N1729, N1602);
buf BUF1 (N1733, N1731);
nor NOR3 (N1734, N1712, N1594, N1702);
not NOT1 (N1735, N1728);
or OR4 (N1736, N1720, N760, N782, N1663);
nor NOR4 (N1737, N1734, N1107, N1105, N871);
not NOT1 (N1738, N1730);
nor NOR4 (N1739, N1725, N1013, N938, N1522);
or OR4 (N1740, N1737, N1671, N536, N1319);
and AND3 (N1741, N1739, N1415, N542);
xor XOR2 (N1742, N1738, N1541);
nor NOR2 (N1743, N1735, N1249);
buf BUF1 (N1744, N1743);
nor NOR2 (N1745, N1741, N986);
or OR4 (N1746, N1744, N1279, N621, N1558);
buf BUF1 (N1747, N1746);
nor NOR4 (N1748, N1724, N1327, N308, N1736);
nand NAND3 (N1749, N1018, N1607, N1024);
and AND3 (N1750, N1742, N1114, N1358);
and AND2 (N1751, N1747, N21);
not NOT1 (N1752, N1701);
nand NAND2 (N1753, N1748, N265);
nor NOR2 (N1754, N1740, N1588);
nor NOR4 (N1755, N1727, N1444, N573, N1675);
or OR4 (N1756, N1749, N246, N458, N282);
and AND4 (N1757, N1752, N1510, N208, N804);
not NOT1 (N1758, N1745);
nand NAND4 (N1759, N1758, N1278, N705, N890);
nand NAND3 (N1760, N1732, N463, N1707);
nor NOR2 (N1761, N1760, N1200);
or OR4 (N1762, N1754, N155, N173, N922);
buf BUF1 (N1763, N1762);
not NOT1 (N1764, N1753);
nand NAND4 (N1765, N1733, N1339, N868, N491);
or OR3 (N1766, N1764, N570, N1018);
buf BUF1 (N1767, N1750);
xor XOR2 (N1768, N1765, N282);
buf BUF1 (N1769, N1763);
nand NAND4 (N1770, N1759, N727, N1174, N1734);
not NOT1 (N1771, N1767);
buf BUF1 (N1772, N1770);
buf BUF1 (N1773, N1768);
buf BUF1 (N1774, N1761);
and AND3 (N1775, N1756, N1109, N1377);
and AND3 (N1776, N1771, N908, N1447);
buf BUF1 (N1777, N1766);
not NOT1 (N1778, N1777);
xor XOR2 (N1779, N1778, N162);
and AND4 (N1780, N1772, N1457, N1631, N1696);
or OR2 (N1781, N1774, N46);
buf BUF1 (N1782, N1769);
and AND3 (N1783, N1751, N708, N1299);
not NOT1 (N1784, N1780);
or OR3 (N1785, N1783, N527, N632);
or OR4 (N1786, N1785, N454, N913, N793);
nor NOR3 (N1787, N1776, N1456, N77);
nand NAND3 (N1788, N1786, N44, N244);
and AND3 (N1789, N1755, N254, N616);
nand NAND4 (N1790, N1779, N256, N1077, N724);
xor XOR2 (N1791, N1790, N1148);
xor XOR2 (N1792, N1787, N1044);
not NOT1 (N1793, N1784);
nand NAND2 (N1794, N1789, N1190);
buf BUF1 (N1795, N1757);
or OR2 (N1796, N1782, N1735);
not NOT1 (N1797, N1793);
xor XOR2 (N1798, N1791, N1001);
xor XOR2 (N1799, N1798, N731);
not NOT1 (N1800, N1788);
nand NAND3 (N1801, N1775, N1462, N1093);
nor NOR4 (N1802, N1792, N501, N630, N421);
nand NAND4 (N1803, N1795, N415, N569, N1103);
not NOT1 (N1804, N1802);
nor NOR2 (N1805, N1794, N1184);
or OR3 (N1806, N1800, N323, N1601);
and AND3 (N1807, N1797, N1066, N1440);
not NOT1 (N1808, N1803);
or OR3 (N1809, N1773, N169, N832);
xor XOR2 (N1810, N1781, N303);
or OR3 (N1811, N1805, N58, N106);
and AND3 (N1812, N1808, N334, N440);
not NOT1 (N1813, N1801);
not NOT1 (N1814, N1812);
nand NAND3 (N1815, N1810, N1641, N941);
nand NAND3 (N1816, N1815, N32, N355);
nor NOR2 (N1817, N1806, N242);
xor XOR2 (N1818, N1809, N1734);
nor NOR4 (N1819, N1816, N177, N1616, N1233);
or OR2 (N1820, N1796, N437);
not NOT1 (N1821, N1819);
or OR4 (N1822, N1818, N1794, N1585, N669);
or OR4 (N1823, N1820, N1786, N1570, N1449);
nor NOR3 (N1824, N1821, N1421, N455);
or OR4 (N1825, N1823, N1522, N1818, N414);
or OR2 (N1826, N1807, N755);
not NOT1 (N1827, N1824);
nand NAND3 (N1828, N1811, N1078, N1421);
and AND4 (N1829, N1799, N1494, N1254, N1188);
nor NOR2 (N1830, N1829, N1365);
and AND4 (N1831, N1828, N483, N1245, N928);
or OR3 (N1832, N1814, N660, N67);
or OR4 (N1833, N1827, N943, N206, N793);
xor XOR2 (N1834, N1831, N981);
buf BUF1 (N1835, N1830);
nand NAND2 (N1836, N1833, N1656);
or OR3 (N1837, N1835, N891, N1272);
and AND3 (N1838, N1836, N1827, N1462);
or OR4 (N1839, N1832, N515, N44, N666);
xor XOR2 (N1840, N1813, N1805);
and AND2 (N1841, N1839, N786);
buf BUF1 (N1842, N1826);
nor NOR2 (N1843, N1817, N913);
not NOT1 (N1844, N1838);
xor XOR2 (N1845, N1844, N1226);
not NOT1 (N1846, N1841);
xor XOR2 (N1847, N1822, N385);
xor XOR2 (N1848, N1840, N286);
nor NOR2 (N1849, N1804, N99);
nand NAND2 (N1850, N1837, N534);
nor NOR3 (N1851, N1834, N1140, N138);
not NOT1 (N1852, N1845);
buf BUF1 (N1853, N1851);
xor XOR2 (N1854, N1853, N376);
buf BUF1 (N1855, N1854);
or OR4 (N1856, N1850, N150, N1402, N680);
not NOT1 (N1857, N1847);
nor NOR4 (N1858, N1852, N1717, N1673, N396);
or OR3 (N1859, N1842, N1115, N1153);
xor XOR2 (N1860, N1848, N1549);
not NOT1 (N1861, N1849);
and AND3 (N1862, N1825, N19, N1546);
and AND2 (N1863, N1861, N1394);
and AND3 (N1864, N1858, N1619, N777);
and AND3 (N1865, N1856, N1252, N736);
not NOT1 (N1866, N1864);
xor XOR2 (N1867, N1843, N1473);
nand NAND3 (N1868, N1866, N760, N527);
not NOT1 (N1869, N1857);
nor NOR2 (N1870, N1869, N1080);
nand NAND4 (N1871, N1868, N461, N822, N1204);
nand NAND2 (N1872, N1867, N1325);
nor NOR2 (N1873, N1855, N312);
buf BUF1 (N1874, N1859);
not NOT1 (N1875, N1865);
xor XOR2 (N1876, N1860, N1711);
nand NAND4 (N1877, N1863, N1768, N1817, N453);
buf BUF1 (N1878, N1873);
or OR2 (N1879, N1878, N1873);
or OR2 (N1880, N1862, N1535);
or OR4 (N1881, N1875, N570, N1604, N1653);
buf BUF1 (N1882, N1846);
or OR3 (N1883, N1876, N1088, N439);
and AND3 (N1884, N1870, N429, N1329);
or OR3 (N1885, N1883, N542, N398);
and AND3 (N1886, N1877, N1463, N125);
xor XOR2 (N1887, N1884, N1079);
buf BUF1 (N1888, N1874);
not NOT1 (N1889, N1887);
buf BUF1 (N1890, N1885);
xor XOR2 (N1891, N1881, N938);
not NOT1 (N1892, N1890);
nand NAND3 (N1893, N1892, N1617, N335);
or OR3 (N1894, N1886, N117, N1479);
not NOT1 (N1895, N1872);
nor NOR2 (N1896, N1882, N1299);
not NOT1 (N1897, N1880);
buf BUF1 (N1898, N1896);
or OR2 (N1899, N1871, N196);
nor NOR3 (N1900, N1893, N293, N1480);
not NOT1 (N1901, N1900);
not NOT1 (N1902, N1889);
and AND4 (N1903, N1888, N535, N447, N838);
nor NOR2 (N1904, N1891, N1304);
buf BUF1 (N1905, N1879);
nand NAND3 (N1906, N1902, N954, N740);
nand NAND4 (N1907, N1903, N700, N1771, N672);
nor NOR2 (N1908, N1895, N1010);
buf BUF1 (N1909, N1894);
nand NAND3 (N1910, N1908, N1393, N174);
nand NAND2 (N1911, N1904, N1347);
and AND2 (N1912, N1899, N1647);
or OR2 (N1913, N1905, N1113);
nand NAND2 (N1914, N1909, N1724);
and AND4 (N1915, N1911, N671, N1116, N844);
not NOT1 (N1916, N1913);
and AND2 (N1917, N1916, N115);
and AND4 (N1918, N1917, N800, N986, N1163);
nor NOR2 (N1919, N1914, N101);
xor XOR2 (N1920, N1901, N708);
nor NOR4 (N1921, N1912, N432, N1499, N830);
buf BUF1 (N1922, N1907);
or OR2 (N1923, N1906, N522);
nor NOR3 (N1924, N1918, N737, N979);
nor NOR3 (N1925, N1919, N1854, N277);
or OR3 (N1926, N1922, N1553, N1418);
nand NAND2 (N1927, N1898, N683);
and AND2 (N1928, N1925, N1515);
or OR2 (N1929, N1915, N1768);
and AND4 (N1930, N1927, N655, N739, N1783);
nand NAND2 (N1931, N1929, N1735);
not NOT1 (N1932, N1910);
and AND4 (N1933, N1923, N957, N507, N71);
nand NAND2 (N1934, N1932, N1566);
and AND4 (N1935, N1934, N427, N487, N785);
or OR2 (N1936, N1920, N417);
nor NOR2 (N1937, N1935, N932);
and AND4 (N1938, N1937, N1014, N1420, N1361);
nand NAND3 (N1939, N1897, N807, N1134);
or OR3 (N1940, N1938, N399, N354);
or OR3 (N1941, N1926, N979, N1682);
not NOT1 (N1942, N1933);
xor XOR2 (N1943, N1924, N1867);
or OR3 (N1944, N1942, N305, N329);
xor XOR2 (N1945, N1943, N1797);
or OR2 (N1946, N1921, N1240);
and AND4 (N1947, N1944, N932, N1266, N80);
and AND3 (N1948, N1939, N424, N1914);
nand NAND2 (N1949, N1945, N962);
nor NOR2 (N1950, N1936, N1574);
or OR2 (N1951, N1930, N1433);
xor XOR2 (N1952, N1947, N1058);
not NOT1 (N1953, N1928);
buf BUF1 (N1954, N1948);
xor XOR2 (N1955, N1931, N594);
buf BUF1 (N1956, N1953);
not NOT1 (N1957, N1949);
not NOT1 (N1958, N1954);
xor XOR2 (N1959, N1955, N1766);
and AND4 (N1960, N1957, N1946, N323, N777);
and AND3 (N1961, N813, N493, N937);
buf BUF1 (N1962, N1958);
not NOT1 (N1963, N1959);
not NOT1 (N1964, N1940);
nor NOR4 (N1965, N1941, N1675, N644, N27);
not NOT1 (N1966, N1956);
not NOT1 (N1967, N1950);
and AND4 (N1968, N1951, N977, N821, N815);
buf BUF1 (N1969, N1964);
and AND2 (N1970, N1966, N1139);
not NOT1 (N1971, N1962);
nand NAND3 (N1972, N1971, N861, N1257);
buf BUF1 (N1973, N1972);
nor NOR4 (N1974, N1960, N403, N1053, N380);
and AND3 (N1975, N1973, N248, N135);
or OR2 (N1976, N1967, N1195);
xor XOR2 (N1977, N1963, N1190);
buf BUF1 (N1978, N1965);
not NOT1 (N1979, N1975);
and AND2 (N1980, N1977, N1310);
buf BUF1 (N1981, N1970);
nor NOR3 (N1982, N1980, N211, N1150);
not NOT1 (N1983, N1969);
xor XOR2 (N1984, N1952, N1324);
nor NOR3 (N1985, N1982, N1516, N1172);
not NOT1 (N1986, N1978);
buf BUF1 (N1987, N1968);
not NOT1 (N1988, N1984);
nand NAND3 (N1989, N1987, N1499, N55);
and AND2 (N1990, N1974, N470);
xor XOR2 (N1991, N1961, N1764);
not NOT1 (N1992, N1983);
nor NOR3 (N1993, N1985, N890, N365);
buf BUF1 (N1994, N1992);
and AND3 (N1995, N1986, N1700, N865);
xor XOR2 (N1996, N1994, N1271);
buf BUF1 (N1997, N1996);
xor XOR2 (N1998, N1993, N1490);
buf BUF1 (N1999, N1998);
nand NAND2 (N2000, N1989, N283);
buf BUF1 (N2001, N1981);
not NOT1 (N2002, N1999);
nor NOR2 (N2003, N1990, N400);
xor XOR2 (N2004, N1979, N148);
and AND4 (N2005, N2004, N1991, N93, N1417);
and AND2 (N2006, N68, N798);
and AND3 (N2007, N2000, N1760, N1507);
buf BUF1 (N2008, N2002);
buf BUF1 (N2009, N1988);
nor NOR2 (N2010, N1976, N803);
nand NAND3 (N2011, N2001, N344, N288);
and AND3 (N2012, N2008, N1488, N1810);
and AND2 (N2013, N2009, N358);
nor NOR3 (N2014, N2010, N459, N918);
xor XOR2 (N2015, N2011, N458);
not NOT1 (N2016, N2014);
and AND3 (N2017, N2015, N318, N267);
or OR4 (N2018, N2016, N406, N1121, N1335);
and AND4 (N2019, N2013, N1847, N1673, N1064);
not NOT1 (N2020, N2005);
and AND4 (N2021, N1995, N2017, N670, N525);
nor NOR4 (N2022, N329, N623, N1122, N1532);
buf BUF1 (N2023, N2019);
buf BUF1 (N2024, N2021);
not NOT1 (N2025, N1997);
buf BUF1 (N2026, N2006);
nand NAND2 (N2027, N2018, N1300);
xor XOR2 (N2028, N2023, N595);
xor XOR2 (N2029, N2026, N1683);
buf BUF1 (N2030, N2028);
nor NOR4 (N2031, N2029, N1556, N193, N1071);
buf BUF1 (N2032, N2027);
buf BUF1 (N2033, N2031);
not NOT1 (N2034, N2030);
nor NOR4 (N2035, N2034, N594, N1053, N1342);
nor NOR2 (N2036, N2020, N605);
and AND2 (N2037, N2003, N118);
and AND2 (N2038, N2033, N1481);
and AND2 (N2039, N2037, N707);
nor NOR4 (N2040, N2038, N2006, N1174, N1649);
or OR4 (N2041, N2025, N1818, N1440, N1048);
and AND2 (N2042, N2032, N1059);
buf BUF1 (N2043, N2024);
nand NAND2 (N2044, N2039, N1288);
buf BUF1 (N2045, N2040);
or OR4 (N2046, N2044, N667, N1588, N1510);
xor XOR2 (N2047, N2042, N49);
or OR3 (N2048, N2007, N350, N890);
buf BUF1 (N2049, N2046);
not NOT1 (N2050, N2047);
and AND2 (N2051, N2035, N45);
not NOT1 (N2052, N2045);
buf BUF1 (N2053, N2041);
buf BUF1 (N2054, N2052);
nor NOR3 (N2055, N2012, N1115, N1067);
nand NAND3 (N2056, N2055, N1051, N460);
buf BUF1 (N2057, N2048);
xor XOR2 (N2058, N2022, N411);
nand NAND2 (N2059, N2053, N972);
not NOT1 (N2060, N2058);
xor XOR2 (N2061, N2050, N181);
buf BUF1 (N2062, N2059);
buf BUF1 (N2063, N2061);
or OR2 (N2064, N2060, N603);
or OR3 (N2065, N2051, N589, N451);
nor NOR2 (N2066, N2057, N940);
nand NAND4 (N2067, N2065, N489, N371, N1192);
xor XOR2 (N2068, N2066, N235);
xor XOR2 (N2069, N2068, N1837);
nor NOR3 (N2070, N2054, N1228, N477);
or OR4 (N2071, N2062, N664, N809, N412);
nor NOR2 (N2072, N2063, N497);
and AND4 (N2073, N2072, N49, N1996, N1167);
nand NAND3 (N2074, N2064, N600, N1068);
buf BUF1 (N2075, N2070);
xor XOR2 (N2076, N2071, N1943);
and AND2 (N2077, N2049, N762);
nor NOR2 (N2078, N2073, N1859);
xor XOR2 (N2079, N2056, N1645);
buf BUF1 (N2080, N2069);
and AND2 (N2081, N2077, N715);
or OR4 (N2082, N2081, N1267, N641, N565);
not NOT1 (N2083, N2078);
nor NOR4 (N2084, N2075, N1306, N214, N595);
buf BUF1 (N2085, N2082);
nor NOR4 (N2086, N2043, N1354, N1091, N1094);
and AND2 (N2087, N2076, N425);
or OR4 (N2088, N2067, N1494, N289, N1947);
or OR2 (N2089, N2083, N984);
and AND4 (N2090, N2086, N1409, N1187, N1851);
and AND4 (N2091, N2090, N1531, N724, N666);
nand NAND3 (N2092, N2085, N101, N19);
or OR4 (N2093, N2036, N526, N707, N1379);
not NOT1 (N2094, N2080);
not NOT1 (N2095, N2094);
xor XOR2 (N2096, N2087, N334);
nor NOR4 (N2097, N2095, N1343, N667, N1135);
nor NOR3 (N2098, N2097, N483, N115);
xor XOR2 (N2099, N2079, N1292);
buf BUF1 (N2100, N2099);
not NOT1 (N2101, N2074);
nor NOR4 (N2102, N2101, N1918, N1079, N56);
nand NAND3 (N2103, N2092, N606, N1710);
buf BUF1 (N2104, N2093);
nor NOR3 (N2105, N2091, N1781, N1562);
buf BUF1 (N2106, N2103);
buf BUF1 (N2107, N2105);
nor NOR3 (N2108, N2107, N1, N1906);
nand NAND2 (N2109, N2106, N1406);
nand NAND3 (N2110, N2108, N473, N1004);
and AND2 (N2111, N2104, N1787);
nor NOR3 (N2112, N2089, N1458, N96);
nor NOR2 (N2113, N2088, N1426);
not NOT1 (N2114, N2113);
nand NAND2 (N2115, N2084, N128);
nand NAND4 (N2116, N2115, N381, N1763, N682);
and AND3 (N2117, N2110, N441, N836);
not NOT1 (N2118, N2111);
not NOT1 (N2119, N2109);
nor NOR3 (N2120, N2117, N1760, N1132);
nand NAND4 (N2121, N2100, N2105, N596, N1418);
nor NOR2 (N2122, N2112, N1102);
nor NOR3 (N2123, N2102, N1710, N1366);
not NOT1 (N2124, N2120);
nand NAND2 (N2125, N2123, N864);
nand NAND4 (N2126, N2114, N1723, N1650, N938);
xor XOR2 (N2127, N2096, N1644);
not NOT1 (N2128, N2119);
and AND4 (N2129, N2122, N1721, N1248, N49);
nor NOR3 (N2130, N2116, N607, N1575);
and AND4 (N2131, N2126, N1449, N1907, N77);
nor NOR2 (N2132, N2121, N1472);
not NOT1 (N2133, N2131);
xor XOR2 (N2134, N2124, N168);
not NOT1 (N2135, N2118);
not NOT1 (N2136, N2127);
buf BUF1 (N2137, N2125);
or OR4 (N2138, N2129, N544, N817, N547);
nand NAND4 (N2139, N2137, N1881, N1804, N1315);
not NOT1 (N2140, N2139);
not NOT1 (N2141, N2136);
and AND2 (N2142, N2133, N1369);
not NOT1 (N2143, N2128);
or OR4 (N2144, N2135, N505, N1885, N66);
xor XOR2 (N2145, N2140, N380);
xor XOR2 (N2146, N2143, N2023);
not NOT1 (N2147, N2142);
xor XOR2 (N2148, N2130, N911);
or OR2 (N2149, N2134, N1560);
nor NOR4 (N2150, N2132, N524, N1330, N662);
not NOT1 (N2151, N2145);
xor XOR2 (N2152, N2151, N723);
nand NAND4 (N2153, N2152, N473, N1390, N1585);
nor NOR2 (N2154, N2150, N1818);
nand NAND4 (N2155, N2154, N936, N2069, N1730);
and AND2 (N2156, N2155, N788);
or OR2 (N2157, N2148, N409);
xor XOR2 (N2158, N2157, N404);
xor XOR2 (N2159, N2146, N1756);
buf BUF1 (N2160, N2147);
nor NOR3 (N2161, N2141, N1596, N1330);
or OR2 (N2162, N2098, N2008);
nor NOR4 (N2163, N2160, N1886, N1451, N1912);
or OR2 (N2164, N2153, N2020);
not NOT1 (N2165, N2156);
nor NOR4 (N2166, N2159, N388, N1394, N412);
buf BUF1 (N2167, N2165);
or OR3 (N2168, N2161, N1431, N381);
not NOT1 (N2169, N2163);
buf BUF1 (N2170, N2164);
not NOT1 (N2171, N2149);
nand NAND2 (N2172, N2138, N1021);
and AND2 (N2173, N2171, N1601);
not NOT1 (N2174, N2168);
buf BUF1 (N2175, N2166);
buf BUF1 (N2176, N2162);
buf BUF1 (N2177, N2172);
nor NOR3 (N2178, N2174, N766, N2099);
nor NOR3 (N2179, N2175, N230, N1346);
or OR4 (N2180, N2179, N514, N431, N1256);
buf BUF1 (N2181, N2180);
nor NOR4 (N2182, N2177, N964, N1382, N2109);
xor XOR2 (N2183, N2182, N1788);
and AND4 (N2184, N2183, N64, N115, N288);
nor NOR3 (N2185, N2170, N1075, N545);
or OR3 (N2186, N2184, N1755, N759);
not NOT1 (N2187, N2169);
or OR2 (N2188, N2185, N1243);
xor XOR2 (N2189, N2173, N2029);
not NOT1 (N2190, N2188);
not NOT1 (N2191, N2144);
buf BUF1 (N2192, N2178);
nor NOR3 (N2193, N2158, N205, N2188);
nand NAND2 (N2194, N2186, N445);
or OR2 (N2195, N2187, N2024);
not NOT1 (N2196, N2176);
xor XOR2 (N2197, N2192, N801);
xor XOR2 (N2198, N2195, N1325);
xor XOR2 (N2199, N2191, N645);
not NOT1 (N2200, N2196);
buf BUF1 (N2201, N2193);
not NOT1 (N2202, N2167);
and AND3 (N2203, N2198, N1912, N1571);
not NOT1 (N2204, N2199);
nand NAND2 (N2205, N2197, N283);
nand NAND4 (N2206, N2202, N1066, N883, N1323);
not NOT1 (N2207, N2189);
xor XOR2 (N2208, N2206, N381);
or OR2 (N2209, N2207, N484);
buf BUF1 (N2210, N2181);
nand NAND4 (N2211, N2210, N321, N530, N958);
or OR4 (N2212, N2194, N2000, N922, N948);
nand NAND3 (N2213, N2212, N743, N70);
nor NOR3 (N2214, N2205, N1715, N1123);
xor XOR2 (N2215, N2190, N1213);
buf BUF1 (N2216, N2213);
buf BUF1 (N2217, N2201);
xor XOR2 (N2218, N2203, N985);
buf BUF1 (N2219, N2215);
not NOT1 (N2220, N2218);
xor XOR2 (N2221, N2220, N662);
nand NAND3 (N2222, N2200, N1819, N1481);
and AND4 (N2223, N2211, N298, N1430, N1904);
nor NOR2 (N2224, N2223, N1719);
buf BUF1 (N2225, N2208);
nor NOR3 (N2226, N2214, N1464, N1348);
buf BUF1 (N2227, N2209);
or OR3 (N2228, N2217, N956, N1811);
xor XOR2 (N2229, N2227, N1452);
nand NAND2 (N2230, N2216, N278);
buf BUF1 (N2231, N2224);
and AND4 (N2232, N2231, N90, N1102, N1107);
and AND4 (N2233, N2232, N527, N988, N1787);
and AND3 (N2234, N2229, N515, N707);
and AND3 (N2235, N2233, N1990, N528);
and AND3 (N2236, N2221, N239, N1653);
buf BUF1 (N2237, N2235);
xor XOR2 (N2238, N2236, N2198);
xor XOR2 (N2239, N2238, N1646);
or OR4 (N2240, N2239, N2118, N975, N382);
or OR4 (N2241, N2237, N1822, N271, N883);
not NOT1 (N2242, N2225);
not NOT1 (N2243, N2234);
not NOT1 (N2244, N2228);
not NOT1 (N2245, N2241);
nand NAND2 (N2246, N2240, N247);
buf BUF1 (N2247, N2204);
not NOT1 (N2248, N2243);
nor NOR2 (N2249, N2242, N650);
and AND4 (N2250, N2226, N1165, N2062, N1704);
and AND4 (N2251, N2250, N1662, N373, N1437);
buf BUF1 (N2252, N2219);
nor NOR4 (N2253, N2247, N367, N1193, N790);
buf BUF1 (N2254, N2252);
or OR2 (N2255, N2245, N656);
not NOT1 (N2256, N2253);
buf BUF1 (N2257, N2251);
not NOT1 (N2258, N2248);
and AND4 (N2259, N2254, N1515, N1159, N302);
nand NAND4 (N2260, N2258, N213, N1957, N2011);
xor XOR2 (N2261, N2260, N1544);
not NOT1 (N2262, N2249);
nand NAND4 (N2263, N2257, N1795, N2190, N1482);
xor XOR2 (N2264, N2230, N1383);
not NOT1 (N2265, N2246);
and AND2 (N2266, N2244, N51);
and AND2 (N2267, N2266, N279);
nor NOR2 (N2268, N2263, N1747);
xor XOR2 (N2269, N2259, N416);
buf BUF1 (N2270, N2262);
or OR2 (N2271, N2256, N348);
buf BUF1 (N2272, N2222);
nand NAND2 (N2273, N2269, N914);
buf BUF1 (N2274, N2264);
or OR2 (N2275, N2274, N1197);
buf BUF1 (N2276, N2273);
or OR3 (N2277, N2276, N1673, N1302);
not NOT1 (N2278, N2272);
buf BUF1 (N2279, N2265);
xor XOR2 (N2280, N2255, N323);
nand NAND2 (N2281, N2271, N478);
and AND3 (N2282, N2281, N1676, N1460);
nand NAND2 (N2283, N2278, N1097);
and AND3 (N2284, N2282, N1089, N504);
buf BUF1 (N2285, N2275);
nand NAND3 (N2286, N2284, N1688, N1234);
or OR4 (N2287, N2267, N754, N1446, N986);
or OR4 (N2288, N2261, N275, N2011, N57);
nand NAND4 (N2289, N2270, N1352, N1678, N1130);
not NOT1 (N2290, N2283);
and AND4 (N2291, N2288, N138, N2086, N2142);
nand NAND3 (N2292, N2291, N197, N2249);
not NOT1 (N2293, N2268);
xor XOR2 (N2294, N2290, N1634);
nor NOR2 (N2295, N2289, N1237);
and AND4 (N2296, N2293, N1037, N102, N1760);
and AND2 (N2297, N2279, N17);
xor XOR2 (N2298, N2285, N1620);
not NOT1 (N2299, N2295);
or OR2 (N2300, N2299, N1973);
xor XOR2 (N2301, N2292, N409);
and AND3 (N2302, N2287, N1754, N945);
or OR4 (N2303, N2296, N925, N1997, N885);
nand NAND4 (N2304, N2286, N1425, N829, N2003);
xor XOR2 (N2305, N2300, N2276);
and AND4 (N2306, N2297, N1343, N212, N1896);
xor XOR2 (N2307, N2301, N648);
nand NAND4 (N2308, N2305, N1214, N619, N2288);
not NOT1 (N2309, N2280);
xor XOR2 (N2310, N2307, N2087);
nand NAND2 (N2311, N2306, N2053);
or OR3 (N2312, N2294, N1263, N277);
and AND4 (N2313, N2304, N1377, N1641, N641);
nand NAND4 (N2314, N2303, N1612, N1007, N814);
nor NOR4 (N2315, N2302, N2062, N940, N1958);
nor NOR2 (N2316, N2312, N1400);
nor NOR4 (N2317, N2315, N357, N1710, N2210);
or OR2 (N2318, N2277, N714);
not NOT1 (N2319, N2318);
not NOT1 (N2320, N2317);
nor NOR3 (N2321, N2311, N928, N1869);
nand NAND4 (N2322, N2321, N2295, N1341, N45);
buf BUF1 (N2323, N2316);
nand NAND4 (N2324, N2310, N1443, N1423, N36);
nand NAND4 (N2325, N2322, N544, N2131, N960);
buf BUF1 (N2326, N2323);
not NOT1 (N2327, N2308);
nand NAND4 (N2328, N2319, N487, N889, N1571);
nand NAND3 (N2329, N2313, N139, N708);
buf BUF1 (N2330, N2325);
nand NAND3 (N2331, N2320, N2251, N1514);
or OR4 (N2332, N2324, N1736, N1025, N1414);
nand NAND2 (N2333, N2330, N624);
not NOT1 (N2334, N2332);
or OR3 (N2335, N2327, N25, N641);
and AND2 (N2336, N2333, N1043);
and AND3 (N2337, N2328, N775, N1785);
nand NAND2 (N2338, N2335, N661);
xor XOR2 (N2339, N2338, N1792);
nand NAND2 (N2340, N2298, N919);
not NOT1 (N2341, N2314);
buf BUF1 (N2342, N2326);
buf BUF1 (N2343, N2339);
not NOT1 (N2344, N2329);
nor NOR3 (N2345, N2331, N1270, N150);
xor XOR2 (N2346, N2343, N1518);
not NOT1 (N2347, N2341);
nand NAND3 (N2348, N2309, N284, N830);
and AND2 (N2349, N2340, N1431);
buf BUF1 (N2350, N2337);
or OR3 (N2351, N2334, N2279, N341);
and AND4 (N2352, N2347, N130, N2157, N1627);
buf BUF1 (N2353, N2350);
buf BUF1 (N2354, N2351);
not NOT1 (N2355, N2348);
buf BUF1 (N2356, N2349);
nand NAND3 (N2357, N2344, N1076, N1131);
buf BUF1 (N2358, N2352);
buf BUF1 (N2359, N2353);
not NOT1 (N2360, N2354);
nand NAND2 (N2361, N2346, N1993);
buf BUF1 (N2362, N2336);
nor NOR2 (N2363, N2342, N943);
xor XOR2 (N2364, N2345, N1682);
xor XOR2 (N2365, N2358, N333);
xor XOR2 (N2366, N2357, N148);
nand NAND2 (N2367, N2356, N2037);
not NOT1 (N2368, N2361);
xor XOR2 (N2369, N2360, N2010);
nand NAND4 (N2370, N2359, N1187, N755, N148);
or OR2 (N2371, N2364, N133);
xor XOR2 (N2372, N2369, N1887);
or OR2 (N2373, N2363, N997);
xor XOR2 (N2374, N2365, N1421);
or OR3 (N2375, N2366, N2213, N2227);
or OR4 (N2376, N2375, N1321, N3, N692);
or OR2 (N2377, N2362, N1522);
or OR3 (N2378, N2377, N1621, N924);
nor NOR2 (N2379, N2371, N1525);
not NOT1 (N2380, N2368);
not NOT1 (N2381, N2376);
xor XOR2 (N2382, N2373, N1617);
nand NAND4 (N2383, N2372, N686, N898, N57);
nand NAND2 (N2384, N2378, N2028);
or OR3 (N2385, N2370, N705, N1744);
xor XOR2 (N2386, N2385, N493);
or OR4 (N2387, N2355, N1339, N1209, N1502);
nand NAND3 (N2388, N2374, N974, N1836);
buf BUF1 (N2389, N2386);
buf BUF1 (N2390, N2387);
buf BUF1 (N2391, N2384);
xor XOR2 (N2392, N2388, N688);
and AND3 (N2393, N2390, N292, N581);
and AND2 (N2394, N2379, N665);
nand NAND2 (N2395, N2382, N2148);
and AND2 (N2396, N2393, N204);
not NOT1 (N2397, N2394);
nand NAND3 (N2398, N2380, N2394, N1441);
or OR2 (N2399, N2389, N260);
not NOT1 (N2400, N2392);
nand NAND4 (N2401, N2367, N1418, N1962, N741);
xor XOR2 (N2402, N2383, N1227);
nand NAND3 (N2403, N2402, N510, N1482);
nor NOR2 (N2404, N2395, N895);
buf BUF1 (N2405, N2404);
xor XOR2 (N2406, N2397, N605);
xor XOR2 (N2407, N2403, N305);
not NOT1 (N2408, N2401);
or OR4 (N2409, N2400, N187, N1620, N1811);
not NOT1 (N2410, N2391);
nor NOR2 (N2411, N2408, N618);
not NOT1 (N2412, N2396);
nor NOR3 (N2413, N2399, N425, N1269);
buf BUF1 (N2414, N2405);
buf BUF1 (N2415, N2410);
nand NAND2 (N2416, N2398, N2120);
xor XOR2 (N2417, N2409, N1911);
or OR2 (N2418, N2412, N307);
nor NOR3 (N2419, N2381, N1085, N575);
or OR2 (N2420, N2417, N259);
buf BUF1 (N2421, N2419);
not NOT1 (N2422, N2406);
or OR3 (N2423, N2420, N1444, N921);
and AND3 (N2424, N2421, N1600, N979);
not NOT1 (N2425, N2411);
nand NAND2 (N2426, N2414, N1762);
nor NOR4 (N2427, N2416, N2207, N1159, N2103);
or OR2 (N2428, N2427, N2253);
buf BUF1 (N2429, N2426);
or OR2 (N2430, N2424, N1319);
not NOT1 (N2431, N2425);
and AND3 (N2432, N2428, N922, N1522);
and AND2 (N2433, N2431, N1449);
buf BUF1 (N2434, N2429);
or OR2 (N2435, N2423, N742);
nand NAND2 (N2436, N2432, N1623);
nor NOR2 (N2437, N2413, N1430);
buf BUF1 (N2438, N2422);
xor XOR2 (N2439, N2430, N1992);
not NOT1 (N2440, N2438);
not NOT1 (N2441, N2415);
buf BUF1 (N2442, N2441);
or OR4 (N2443, N2407, N651, N686, N1955);
xor XOR2 (N2444, N2433, N542);
and AND3 (N2445, N2443, N2064, N830);
xor XOR2 (N2446, N2435, N905);
nand NAND2 (N2447, N2418, N1957);
nand NAND4 (N2448, N2447, N99, N694, N829);
buf BUF1 (N2449, N2439);
buf BUF1 (N2450, N2434);
xor XOR2 (N2451, N2436, N861);
not NOT1 (N2452, N2442);
nand NAND2 (N2453, N2452, N621);
nand NAND3 (N2454, N2448, N977, N728);
or OR3 (N2455, N2445, N1913, N2449);
or OR4 (N2456, N335, N1568, N2323, N239);
and AND4 (N2457, N2444, N177, N265, N1229);
and AND2 (N2458, N2455, N308);
not NOT1 (N2459, N2440);
nor NOR4 (N2460, N2437, N1563, N2365, N2029);
not NOT1 (N2461, N2457);
xor XOR2 (N2462, N2451, N1688);
xor XOR2 (N2463, N2462, N1168);
not NOT1 (N2464, N2459);
xor XOR2 (N2465, N2446, N726);
nand NAND3 (N2466, N2461, N2081, N525);
buf BUF1 (N2467, N2466);
or OR3 (N2468, N2450, N207, N443);
and AND3 (N2469, N2464, N1876, N466);
xor XOR2 (N2470, N2463, N2334);
not NOT1 (N2471, N2453);
or OR3 (N2472, N2470, N2032, N2075);
and AND2 (N2473, N2469, N1770);
not NOT1 (N2474, N2467);
or OR4 (N2475, N2460, N957, N2300, N1753);
buf BUF1 (N2476, N2471);
xor XOR2 (N2477, N2454, N1092);
or OR2 (N2478, N2473, N1320);
nand NAND4 (N2479, N2474, N757, N1731, N73);
nor NOR3 (N2480, N2479, N947, N1291);
nand NAND4 (N2481, N2458, N2386, N1645, N410);
or OR3 (N2482, N2480, N853, N1924);
nand NAND4 (N2483, N2456, N880, N232, N594);
buf BUF1 (N2484, N2475);
or OR4 (N2485, N2483, N870, N719, N937);
not NOT1 (N2486, N2485);
or OR4 (N2487, N2468, N54, N1244, N2392);
nand NAND2 (N2488, N2465, N854);
xor XOR2 (N2489, N2484, N2114);
or OR2 (N2490, N2478, N1065);
and AND4 (N2491, N2486, N1571, N1380, N1385);
nand NAND3 (N2492, N2477, N1718, N1873);
buf BUF1 (N2493, N2491);
or OR4 (N2494, N2481, N2265, N778, N1626);
not NOT1 (N2495, N2490);
not NOT1 (N2496, N2472);
nand NAND2 (N2497, N2496, N1068);
not NOT1 (N2498, N2493);
or OR2 (N2499, N2498, N1250);
and AND2 (N2500, N2488, N1685);
or OR3 (N2501, N2495, N1343, N763);
and AND4 (N2502, N2492, N819, N2054, N325);
or OR3 (N2503, N2497, N1245, N1560);
xor XOR2 (N2504, N2503, N1846);
xor XOR2 (N2505, N2502, N2419);
nor NOR4 (N2506, N2489, N842, N1599, N645);
nand NAND2 (N2507, N2501, N620);
not NOT1 (N2508, N2494);
nand NAND2 (N2509, N2500, N926);
not NOT1 (N2510, N2506);
xor XOR2 (N2511, N2504, N211);
or OR3 (N2512, N2487, N2244, N901);
and AND3 (N2513, N2499, N2220, N2226);
or OR3 (N2514, N2507, N268, N1765);
xor XOR2 (N2515, N2505, N1020);
nand NAND2 (N2516, N2512, N503);
and AND2 (N2517, N2510, N2090);
nor NOR4 (N2518, N2514, N784, N2373, N2465);
and AND4 (N2519, N2518, N1205, N2072, N231);
not NOT1 (N2520, N2511);
nor NOR4 (N2521, N2517, N38, N1461, N335);
and AND2 (N2522, N2519, N806);
nand NAND4 (N2523, N2513, N2021, N27, N684);
xor XOR2 (N2524, N2508, N330);
not NOT1 (N2525, N2521);
or OR4 (N2526, N2523, N2164, N2284, N682);
xor XOR2 (N2527, N2476, N694);
nand NAND4 (N2528, N2522, N2370, N1103, N1037);
xor XOR2 (N2529, N2509, N887);
nor NOR4 (N2530, N2528, N1712, N941, N2480);
not NOT1 (N2531, N2524);
buf BUF1 (N2532, N2526);
or OR4 (N2533, N2529, N2039, N1058, N2266);
nor NOR3 (N2534, N2533, N1073, N171);
xor XOR2 (N2535, N2532, N1328);
nor NOR3 (N2536, N2525, N933, N2054);
and AND3 (N2537, N2536, N42, N2169);
xor XOR2 (N2538, N2527, N1767);
not NOT1 (N2539, N2537);
xor XOR2 (N2540, N2535, N1522);
nand NAND3 (N2541, N2531, N89, N1728);
not NOT1 (N2542, N2534);
buf BUF1 (N2543, N2538);
not NOT1 (N2544, N2515);
nand NAND3 (N2545, N2544, N2209, N2087);
not NOT1 (N2546, N2540);
xor XOR2 (N2547, N2516, N2306);
xor XOR2 (N2548, N2547, N481);
not NOT1 (N2549, N2545);
nor NOR3 (N2550, N2539, N2527, N1952);
not NOT1 (N2551, N2546);
and AND4 (N2552, N2551, N669, N1479, N1218);
nand NAND3 (N2553, N2482, N806, N1099);
nor NOR3 (N2554, N2541, N2329, N1999);
nand NAND2 (N2555, N2550, N142);
nand NAND4 (N2556, N2520, N1564, N809, N1034);
nor NOR3 (N2557, N2556, N1734, N159);
and AND3 (N2558, N2557, N1163, N2428);
nand NAND2 (N2559, N2554, N498);
nor NOR3 (N2560, N2558, N861, N1421);
nand NAND3 (N2561, N2559, N2338, N458);
not NOT1 (N2562, N2543);
nor NOR3 (N2563, N2561, N516, N770);
or OR4 (N2564, N2555, N1571, N2016, N148);
not NOT1 (N2565, N2549);
or OR3 (N2566, N2530, N1090, N1909);
or OR4 (N2567, N2565, N122, N722, N500);
not NOT1 (N2568, N2542);
and AND3 (N2569, N2553, N2417, N966);
and AND2 (N2570, N2560, N49);
or OR2 (N2571, N2563, N691);
xor XOR2 (N2572, N2566, N627);
buf BUF1 (N2573, N2548);
and AND3 (N2574, N2572, N1986, N13);
or OR2 (N2575, N2562, N831);
or OR4 (N2576, N2567, N2092, N137, N187);
nor NOR4 (N2577, N2568, N154, N1235, N148);
or OR2 (N2578, N2573, N33);
or OR2 (N2579, N2578, N1356);
buf BUF1 (N2580, N2552);
xor XOR2 (N2581, N2571, N2051);
buf BUF1 (N2582, N2576);
nor NOR2 (N2583, N2579, N552);
and AND3 (N2584, N2580, N2532, N1116);
or OR4 (N2585, N2575, N1083, N2302, N2023);
not NOT1 (N2586, N2583);
buf BUF1 (N2587, N2584);
xor XOR2 (N2588, N2585, N1298);
nand NAND2 (N2589, N2564, N11);
xor XOR2 (N2590, N2587, N229);
xor XOR2 (N2591, N2570, N371);
buf BUF1 (N2592, N2577);
buf BUF1 (N2593, N2586);
and AND4 (N2594, N2588, N194, N2297, N2413);
or OR4 (N2595, N2594, N1154, N1853, N2592);
nand NAND4 (N2596, N2393, N128, N235, N1819);
and AND2 (N2597, N2596, N2044);
nand NAND4 (N2598, N2595, N237, N2474, N1426);
xor XOR2 (N2599, N2591, N1920);
buf BUF1 (N2600, N2593);
and AND2 (N2601, N2581, N2391);
or OR4 (N2602, N2589, N2121, N132, N1893);
and AND4 (N2603, N2574, N34, N1019, N1955);
xor XOR2 (N2604, N2603, N2229);
not NOT1 (N2605, N2604);
or OR4 (N2606, N2582, N916, N285, N749);
or OR4 (N2607, N2598, N2419, N1605, N901);
xor XOR2 (N2608, N2606, N102);
and AND3 (N2609, N2590, N1332, N1406);
nor NOR2 (N2610, N2608, N2460);
and AND3 (N2611, N2597, N2460, N147);
nand NAND3 (N2612, N2600, N188, N1733);
xor XOR2 (N2613, N2599, N2175);
or OR3 (N2614, N2613, N1514, N2384);
and AND4 (N2615, N2605, N1868, N1890, N2171);
xor XOR2 (N2616, N2610, N124);
or OR4 (N2617, N2614, N1792, N1203, N1353);
and AND2 (N2618, N2602, N1815);
nand NAND4 (N2619, N2617, N2557, N1156, N1931);
or OR3 (N2620, N2612, N1241, N1516);
nand NAND2 (N2621, N2607, N1857);
or OR4 (N2622, N2615, N414, N1312, N1218);
or OR4 (N2623, N2609, N49, N876, N567);
not NOT1 (N2624, N2618);
or OR3 (N2625, N2623, N1352, N2397);
not NOT1 (N2626, N2622);
nor NOR3 (N2627, N2624, N122, N290);
and AND2 (N2628, N2601, N862);
not NOT1 (N2629, N2621);
buf BUF1 (N2630, N2625);
not NOT1 (N2631, N2628);
or OR3 (N2632, N2627, N654, N2434);
nor NOR3 (N2633, N2630, N2004, N1587);
buf BUF1 (N2634, N2633);
and AND4 (N2635, N2632, N2033, N2452, N1383);
xor XOR2 (N2636, N2629, N287);
nor NOR2 (N2637, N2616, N1598);
nand NAND3 (N2638, N2611, N2594, N2440);
nand NAND4 (N2639, N2626, N2494, N1247, N638);
nand NAND4 (N2640, N2634, N929, N2414, N2148);
nand NAND4 (N2641, N2637, N1993, N1733, N916);
nor NOR2 (N2642, N2619, N2102);
buf BUF1 (N2643, N2640);
or OR3 (N2644, N2631, N1059, N337);
nor NOR4 (N2645, N2635, N771, N2136, N2031);
nor NOR2 (N2646, N2643, N882);
buf BUF1 (N2647, N2645);
xor XOR2 (N2648, N2620, N662);
or OR3 (N2649, N2638, N750, N238);
buf BUF1 (N2650, N2649);
nand NAND2 (N2651, N2646, N305);
xor XOR2 (N2652, N2648, N2142);
or OR3 (N2653, N2639, N771, N1168);
or OR4 (N2654, N2651, N2476, N2589, N491);
not NOT1 (N2655, N2654);
and AND2 (N2656, N2655, N1951);
buf BUF1 (N2657, N2653);
nand NAND2 (N2658, N2657, N1817);
nor NOR2 (N2659, N2656, N932);
and AND2 (N2660, N2647, N1923);
nor NOR3 (N2661, N2660, N727, N1931);
nand NAND4 (N2662, N2642, N2257, N83, N90);
not NOT1 (N2663, N2652);
nand NAND2 (N2664, N2661, N195);
not NOT1 (N2665, N2658);
xor XOR2 (N2666, N2636, N1912);
buf BUF1 (N2667, N2666);
not NOT1 (N2668, N2663);
nand NAND4 (N2669, N2641, N1443, N2422, N383);
and AND2 (N2670, N2665, N1174);
xor XOR2 (N2671, N2644, N1856);
nand NAND4 (N2672, N2667, N2352, N137, N685);
or OR3 (N2673, N2662, N391, N1977);
nor NOR4 (N2674, N2671, N2651, N898, N1452);
and AND4 (N2675, N2569, N1743, N97, N212);
and AND4 (N2676, N2672, N1251, N188, N2661);
and AND2 (N2677, N2650, N782);
not NOT1 (N2678, N2670);
nor NOR4 (N2679, N2664, N2027, N1075, N1128);
nor NOR3 (N2680, N2675, N1712, N2236);
not NOT1 (N2681, N2677);
xor XOR2 (N2682, N2668, N623);
buf BUF1 (N2683, N2678);
nand NAND2 (N2684, N2669, N1324);
not NOT1 (N2685, N2684);
buf BUF1 (N2686, N2673);
buf BUF1 (N2687, N2682);
buf BUF1 (N2688, N2687);
not NOT1 (N2689, N2674);
nor NOR3 (N2690, N2681, N1489, N565);
nand NAND2 (N2691, N2679, N2500);
nor NOR3 (N2692, N2691, N2612, N756);
and AND3 (N2693, N2685, N1604, N2075);
nor NOR2 (N2694, N2676, N878);
buf BUF1 (N2695, N2688);
buf BUF1 (N2696, N2659);
buf BUF1 (N2697, N2686);
nor NOR3 (N2698, N2692, N259, N1207);
and AND3 (N2699, N2689, N925, N1433);
and AND4 (N2700, N2699, N2254, N182, N754);
xor XOR2 (N2701, N2695, N2318);
xor XOR2 (N2702, N2700, N82);
or OR3 (N2703, N2683, N2593, N1562);
buf BUF1 (N2704, N2696);
xor XOR2 (N2705, N2680, N1483);
nand NAND2 (N2706, N2702, N1105);
and AND4 (N2707, N2701, N1799, N1944, N60);
not NOT1 (N2708, N2690);
not NOT1 (N2709, N2708);
or OR2 (N2710, N2704, N2675);
xor XOR2 (N2711, N2707, N2144);
xor XOR2 (N2712, N2706, N1214);
nand NAND3 (N2713, N2703, N1567, N2228);
not NOT1 (N2714, N2711);
buf BUF1 (N2715, N2698);
and AND3 (N2716, N2712, N833, N1882);
xor XOR2 (N2717, N2714, N2696);
nor NOR4 (N2718, N2715, N1973, N1120, N829);
or OR3 (N2719, N2694, N921, N2546);
not NOT1 (N2720, N2716);
not NOT1 (N2721, N2719);
nand NAND3 (N2722, N2697, N968, N201);
not NOT1 (N2723, N2705);
or OR4 (N2724, N2709, N329, N2667, N1954);
xor XOR2 (N2725, N2723, N1982);
or OR2 (N2726, N2720, N2494);
nand NAND3 (N2727, N2721, N1210, N2726);
buf BUF1 (N2728, N487);
buf BUF1 (N2729, N2710);
and AND3 (N2730, N2713, N1694, N2419);
buf BUF1 (N2731, N2729);
or OR4 (N2732, N2724, N1147, N46, N1382);
xor XOR2 (N2733, N2730, N499);
nor NOR4 (N2734, N2725, N2595, N442, N1401);
xor XOR2 (N2735, N2717, N457);
xor XOR2 (N2736, N2727, N1191);
not NOT1 (N2737, N2722);
nand NAND2 (N2738, N2733, N1171);
nor NOR4 (N2739, N2732, N181, N998, N743);
nor NOR2 (N2740, N2735, N2685);
buf BUF1 (N2741, N2734);
and AND4 (N2742, N2740, N2263, N2517, N263);
nand NAND4 (N2743, N2739, N149, N1067, N2287);
nand NAND3 (N2744, N2731, N2475, N1794);
nor NOR4 (N2745, N2736, N2441, N1542, N931);
buf BUF1 (N2746, N2728);
xor XOR2 (N2747, N2741, N2228);
and AND2 (N2748, N2718, N779);
not NOT1 (N2749, N2744);
or OR2 (N2750, N2747, N2219);
not NOT1 (N2751, N2738);
or OR3 (N2752, N2693, N2040, N2552);
buf BUF1 (N2753, N2737);
xor XOR2 (N2754, N2748, N2024);
or OR3 (N2755, N2751, N522, N1057);
not NOT1 (N2756, N2754);
or OR2 (N2757, N2755, N450);
nand NAND2 (N2758, N2743, N2339);
not NOT1 (N2759, N2752);
xor XOR2 (N2760, N2757, N366);
and AND2 (N2761, N2749, N1165);
nand NAND2 (N2762, N2750, N1772);
not NOT1 (N2763, N2756);
or OR4 (N2764, N2753, N774, N1950, N2602);
and AND2 (N2765, N2764, N646);
nor NOR4 (N2766, N2745, N2052, N695, N900);
not NOT1 (N2767, N2759);
xor XOR2 (N2768, N2760, N947);
xor XOR2 (N2769, N2758, N2001);
and AND2 (N2770, N2766, N2507);
buf BUF1 (N2771, N2767);
xor XOR2 (N2772, N2761, N960);
buf BUF1 (N2773, N2742);
buf BUF1 (N2774, N2773);
xor XOR2 (N2775, N2774, N518);
xor XOR2 (N2776, N2769, N263);
and AND4 (N2777, N2765, N1846, N1479, N1853);
or OR3 (N2778, N2775, N1333, N434);
nand NAND4 (N2779, N2777, N1768, N1439, N202);
nand NAND3 (N2780, N2778, N1367, N625);
or OR2 (N2781, N2776, N1780);
nor NOR3 (N2782, N2781, N1125, N479);
buf BUF1 (N2783, N2772);
and AND3 (N2784, N2770, N1541, N1130);
not NOT1 (N2785, N2782);
xor XOR2 (N2786, N2771, N2551);
nand NAND3 (N2787, N2785, N1874, N435);
not NOT1 (N2788, N2786);
nor NOR3 (N2789, N2780, N276, N602);
nand NAND3 (N2790, N2763, N617, N2451);
or OR4 (N2791, N2788, N2762, N33, N1452);
and AND2 (N2792, N1657, N1678);
nor NOR2 (N2793, N2768, N907);
nand NAND2 (N2794, N2793, N2197);
buf BUF1 (N2795, N2789);
xor XOR2 (N2796, N2791, N2021);
buf BUF1 (N2797, N2795);
not NOT1 (N2798, N2794);
xor XOR2 (N2799, N2790, N199);
not NOT1 (N2800, N2799);
nor NOR3 (N2801, N2779, N48, N1611);
and AND3 (N2802, N2783, N2663, N540);
nor NOR4 (N2803, N2797, N959, N1561, N246);
and AND2 (N2804, N2801, N2152);
buf BUF1 (N2805, N2804);
or OR3 (N2806, N2798, N648, N458);
and AND3 (N2807, N2746, N1391, N2303);
or OR2 (N2808, N2792, N7);
nor NOR3 (N2809, N2806, N2412, N2646);
xor XOR2 (N2810, N2803, N908);
or OR3 (N2811, N2809, N1391, N1987);
and AND4 (N2812, N2802, N924, N609, N2544);
xor XOR2 (N2813, N2808, N676);
or OR4 (N2814, N2784, N1080, N1496, N46);
or OR3 (N2815, N2814, N529, N956);
not NOT1 (N2816, N2815);
buf BUF1 (N2817, N2812);
buf BUF1 (N2818, N2813);
nand NAND2 (N2819, N2810, N40);
or OR4 (N2820, N2805, N1461, N1761, N1713);
buf BUF1 (N2821, N2796);
or OR2 (N2822, N2807, N2367);
buf BUF1 (N2823, N2820);
and AND2 (N2824, N2817, N1005);
and AND3 (N2825, N2800, N372, N1323);
nor NOR3 (N2826, N2821, N1351, N1544);
xor XOR2 (N2827, N2819, N2371);
not NOT1 (N2828, N2825);
buf BUF1 (N2829, N2826);
xor XOR2 (N2830, N2787, N695);
xor XOR2 (N2831, N2830, N1391);
nor NOR2 (N2832, N2823, N859);
not NOT1 (N2833, N2824);
and AND4 (N2834, N2829, N1566, N39, N202);
buf BUF1 (N2835, N2822);
xor XOR2 (N2836, N2828, N39);
xor XOR2 (N2837, N2832, N1995);
not NOT1 (N2838, N2837);
nor NOR3 (N2839, N2834, N2195, N362);
buf BUF1 (N2840, N2816);
not NOT1 (N2841, N2831);
xor XOR2 (N2842, N2840, N519);
xor XOR2 (N2843, N2833, N1625);
buf BUF1 (N2844, N2842);
nor NOR2 (N2845, N2811, N1459);
nor NOR3 (N2846, N2838, N75, N2209);
not NOT1 (N2847, N2836);
nor NOR2 (N2848, N2847, N2089);
buf BUF1 (N2849, N2844);
buf BUF1 (N2850, N2835);
and AND2 (N2851, N2849, N1578);
and AND3 (N2852, N2839, N1303, N2008);
nor NOR2 (N2853, N2841, N2655);
nor NOR4 (N2854, N2846, N1, N980, N1559);
or OR3 (N2855, N2854, N2385, N685);
not NOT1 (N2856, N2848);
buf BUF1 (N2857, N2845);
or OR2 (N2858, N2850, N520);
or OR2 (N2859, N2843, N836);
xor XOR2 (N2860, N2827, N729);
not NOT1 (N2861, N2858);
or OR2 (N2862, N2859, N2845);
nor NOR2 (N2863, N2862, N1724);
nand NAND4 (N2864, N2861, N1256, N2850, N596);
buf BUF1 (N2865, N2855);
nor NOR3 (N2866, N2865, N835, N673);
or OR2 (N2867, N2857, N70);
not NOT1 (N2868, N2851);
or OR4 (N2869, N2818, N2567, N1258, N2012);
not NOT1 (N2870, N2856);
buf BUF1 (N2871, N2864);
and AND4 (N2872, N2869, N1701, N2733, N1571);
xor XOR2 (N2873, N2871, N1505);
nand NAND3 (N2874, N2872, N229, N772);
not NOT1 (N2875, N2853);
nand NAND3 (N2876, N2860, N964, N132);
or OR2 (N2877, N2874, N1703);
and AND3 (N2878, N2876, N2533, N773);
buf BUF1 (N2879, N2870);
not NOT1 (N2880, N2852);
xor XOR2 (N2881, N2875, N1887);
buf BUF1 (N2882, N2868);
buf BUF1 (N2883, N2873);
xor XOR2 (N2884, N2883, N1327);
nor NOR3 (N2885, N2863, N2250, N664);
or OR4 (N2886, N2878, N359, N1814, N795);
buf BUF1 (N2887, N2882);
not NOT1 (N2888, N2885);
nor NOR4 (N2889, N2866, N187, N1710, N952);
nor NOR2 (N2890, N2879, N1425);
xor XOR2 (N2891, N2884, N1598);
buf BUF1 (N2892, N2867);
nand NAND4 (N2893, N2887, N1002, N1251, N2038);
or OR3 (N2894, N2890, N884, N2758);
nand NAND3 (N2895, N2889, N1083, N1996);
and AND4 (N2896, N2893, N2109, N177, N1292);
buf BUF1 (N2897, N2881);
and AND2 (N2898, N2877, N2101);
xor XOR2 (N2899, N2886, N2177);
or OR3 (N2900, N2898, N1744, N195);
buf BUF1 (N2901, N2888);
xor XOR2 (N2902, N2892, N2266);
xor XOR2 (N2903, N2896, N1003);
nand NAND4 (N2904, N2903, N2580, N2344, N2684);
and AND4 (N2905, N2895, N976, N1933, N319);
or OR4 (N2906, N2902, N1194, N1972, N618);
xor XOR2 (N2907, N2900, N2267);
nand NAND4 (N2908, N2894, N2306, N318, N87);
xor XOR2 (N2909, N2901, N2565);
buf BUF1 (N2910, N2908);
or OR2 (N2911, N2906, N2799);
not NOT1 (N2912, N2904);
xor XOR2 (N2913, N2912, N636);
buf BUF1 (N2914, N2910);
and AND2 (N2915, N2907, N2376);
or OR3 (N2916, N2897, N86, N1174);
and AND2 (N2917, N2905, N706);
xor XOR2 (N2918, N2899, N641);
and AND4 (N2919, N2891, N745, N2745, N2440);
and AND3 (N2920, N2909, N2394, N2756);
xor XOR2 (N2921, N2920, N398);
not NOT1 (N2922, N2913);
or OR2 (N2923, N2917, N2756);
buf BUF1 (N2924, N2923);
buf BUF1 (N2925, N2918);
nor NOR4 (N2926, N2880, N2500, N554, N1645);
nand NAND4 (N2927, N2914, N379, N2022, N1518);
buf BUF1 (N2928, N2924);
or OR2 (N2929, N2925, N2271);
buf BUF1 (N2930, N2919);
nand NAND2 (N2931, N2911, N808);
and AND4 (N2932, N2921, N2557, N2861, N710);
nor NOR2 (N2933, N2929, N177);
and AND2 (N2934, N2916, N1102);
nor NOR3 (N2935, N2932, N1153, N1656);
nor NOR4 (N2936, N2928, N1555, N1711, N2912);
xor XOR2 (N2937, N2933, N2614);
and AND3 (N2938, N2937, N9, N1839);
and AND2 (N2939, N2934, N2546);
buf BUF1 (N2940, N2915);
xor XOR2 (N2941, N2927, N155);
or OR2 (N2942, N2931, N750);
not NOT1 (N2943, N2930);
xor XOR2 (N2944, N2941, N1803);
or OR4 (N2945, N2922, N2433, N971, N2670);
xor XOR2 (N2946, N2939, N2472);
and AND2 (N2947, N2935, N1175);
nor NOR3 (N2948, N2942, N210, N127);
nand NAND2 (N2949, N2948, N1317);
and AND4 (N2950, N2936, N234, N2000, N819);
xor XOR2 (N2951, N2943, N880);
buf BUF1 (N2952, N2944);
or OR3 (N2953, N2946, N1234, N1860);
and AND3 (N2954, N2926, N2327, N31);
xor XOR2 (N2955, N2938, N504);
or OR2 (N2956, N2947, N600);
xor XOR2 (N2957, N2953, N771);
not NOT1 (N2958, N2956);
nor NOR3 (N2959, N2951, N1524, N2028);
buf BUF1 (N2960, N2955);
nor NOR4 (N2961, N2949, N2207, N2262, N2657);
buf BUF1 (N2962, N2959);
nor NOR3 (N2963, N2952, N799, N271);
or OR3 (N2964, N2945, N2502, N2602);
not NOT1 (N2965, N2964);
nand NAND2 (N2966, N2962, N448);
buf BUF1 (N2967, N2950);
and AND4 (N2968, N2961, N2723, N2594, N2029);
not NOT1 (N2969, N2968);
xor XOR2 (N2970, N2967, N2639);
buf BUF1 (N2971, N2963);
or OR3 (N2972, N2970, N56, N1634);
nor NOR2 (N2973, N2971, N2535);
or OR3 (N2974, N2966, N2063, N141);
nor NOR3 (N2975, N2973, N820, N78);
not NOT1 (N2976, N2940);
nor NOR2 (N2977, N2960, N53);
or OR2 (N2978, N2976, N2279);
and AND3 (N2979, N2958, N1368, N2734);
and AND3 (N2980, N2972, N772, N1754);
and AND2 (N2981, N2957, N2264);
nor NOR4 (N2982, N2969, N313, N2662, N1909);
and AND4 (N2983, N2981, N1119, N288, N1166);
xor XOR2 (N2984, N2977, N1819);
not NOT1 (N2985, N2980);
nand NAND2 (N2986, N2975, N2604);
xor XOR2 (N2987, N2979, N426);
and AND3 (N2988, N2986, N2661, N322);
and AND4 (N2989, N2974, N666, N438, N2010);
or OR2 (N2990, N2978, N427);
not NOT1 (N2991, N2990);
not NOT1 (N2992, N2954);
nor NOR4 (N2993, N2992, N2791, N1299, N1622);
not NOT1 (N2994, N2982);
buf BUF1 (N2995, N2991);
buf BUF1 (N2996, N2983);
nand NAND4 (N2997, N2965, N1288, N2798, N1231);
nor NOR3 (N2998, N2987, N963, N1634);
and AND2 (N2999, N2997, N603);
nor NOR4 (N3000, N2993, N2505, N56, N1098);
buf BUF1 (N3001, N2984);
xor XOR2 (N3002, N2998, N2811);
nor NOR4 (N3003, N2995, N2660, N2584, N320);
or OR2 (N3004, N2994, N403);
nand NAND4 (N3005, N2989, N569, N2471, N2986);
nand NAND4 (N3006, N3003, N394, N2340, N289);
nor NOR3 (N3007, N2988, N1825, N1362);
xor XOR2 (N3008, N3001, N1296);
xor XOR2 (N3009, N3000, N1548);
nand NAND3 (N3010, N3006, N253, N1110);
nand NAND3 (N3011, N3008, N2251, N1706);
xor XOR2 (N3012, N2999, N1375);
buf BUF1 (N3013, N3002);
not NOT1 (N3014, N3013);
or OR3 (N3015, N3009, N517, N403);
xor XOR2 (N3016, N3015, N652);
buf BUF1 (N3017, N3010);
nand NAND2 (N3018, N3017, N1465);
nor NOR3 (N3019, N3007, N884, N754);
not NOT1 (N3020, N2996);
buf BUF1 (N3021, N3012);
or OR4 (N3022, N3018, N2754, N1294, N2120);
nor NOR4 (N3023, N3011, N137, N2651, N1682);
xor XOR2 (N3024, N3021, N1308);
nand NAND4 (N3025, N3019, N518, N87, N2029);
buf BUF1 (N3026, N3005);
nand NAND3 (N3027, N3014, N2444, N2539);
buf BUF1 (N3028, N3027);
or OR2 (N3029, N3004, N1134);
xor XOR2 (N3030, N3029, N1403);
and AND2 (N3031, N3022, N287);
xor XOR2 (N3032, N2985, N2517);
nor NOR4 (N3033, N3020, N2265, N1998, N2616);
xor XOR2 (N3034, N3030, N2336);
buf BUF1 (N3035, N3025);
not NOT1 (N3036, N3033);
nor NOR4 (N3037, N3016, N758, N2476, N2855);
xor XOR2 (N3038, N3036, N851);
or OR3 (N3039, N3031, N914, N503);
xor XOR2 (N3040, N3026, N806);
and AND4 (N3041, N3028, N1366, N1050, N1275);
buf BUF1 (N3042, N3023);
xor XOR2 (N3043, N3041, N2854);
nor NOR3 (N3044, N3042, N377, N872);
or OR3 (N3045, N3043, N635, N1831);
nand NAND2 (N3046, N3034, N1545);
and AND3 (N3047, N3024, N962, N2287);
or OR3 (N3048, N3047, N1084, N2486);
not NOT1 (N3049, N3038);
and AND4 (N3050, N3037, N818, N613, N307);
not NOT1 (N3051, N3045);
xor XOR2 (N3052, N3032, N1771);
nor NOR4 (N3053, N3051, N722, N1631, N1255);
buf BUF1 (N3054, N3052);
or OR2 (N3055, N3048, N2707);
nand NAND3 (N3056, N3050, N1243, N2254);
not NOT1 (N3057, N3054);
not NOT1 (N3058, N3046);
not NOT1 (N3059, N3055);
and AND4 (N3060, N3049, N1908, N2737, N967);
xor XOR2 (N3061, N3044, N868);
buf BUF1 (N3062, N3039);
nand NAND3 (N3063, N3062, N2452, N2509);
nand NAND2 (N3064, N3035, N564);
nand NAND3 (N3065, N3060, N1209, N1947);
xor XOR2 (N3066, N3040, N26);
or OR3 (N3067, N3061, N2361, N2412);
nand NAND3 (N3068, N3053, N1997, N535);
and AND3 (N3069, N3064, N2992, N1389);
nand NAND4 (N3070, N3068, N691, N1275, N694);
not NOT1 (N3071, N3069);
or OR4 (N3072, N3059, N866, N2956, N2110);
xor XOR2 (N3073, N3071, N2559);
buf BUF1 (N3074, N3070);
or OR2 (N3075, N3056, N2169);
and AND4 (N3076, N3074, N167, N1843, N2025);
or OR2 (N3077, N3058, N1958);
nand NAND2 (N3078, N3057, N239);
buf BUF1 (N3079, N3075);
not NOT1 (N3080, N3077);
buf BUF1 (N3081, N3078);
nand NAND2 (N3082, N3081, N1673);
or OR2 (N3083, N3082, N2573);
nor NOR2 (N3084, N3063, N1796);
not NOT1 (N3085, N3084);
nor NOR3 (N3086, N3076, N142, N403);
not NOT1 (N3087, N3086);
not NOT1 (N3088, N3072);
not NOT1 (N3089, N3083);
not NOT1 (N3090, N3085);
nand NAND3 (N3091, N3067, N584, N1504);
nor NOR3 (N3092, N3091, N1379, N836);
nand NAND2 (N3093, N3088, N2551);
nor NOR4 (N3094, N3065, N757, N2027, N2915);
xor XOR2 (N3095, N3066, N2708);
nand NAND2 (N3096, N3087, N217);
and AND2 (N3097, N3092, N2395);
nand NAND3 (N3098, N3090, N1065, N204);
buf BUF1 (N3099, N3073);
not NOT1 (N3100, N3079);
nand NAND4 (N3101, N3095, N2019, N2147, N506);
nand NAND4 (N3102, N3093, N428, N745, N2075);
or OR3 (N3103, N3080, N1553, N3097);
buf BUF1 (N3104, N493);
nand NAND2 (N3105, N3098, N45);
xor XOR2 (N3106, N3089, N765);
xor XOR2 (N3107, N3094, N1251);
nor NOR2 (N3108, N3106, N353);
or OR4 (N3109, N3096, N2999, N2663, N655);
nor NOR2 (N3110, N3109, N2505);
or OR2 (N3111, N3110, N904);
buf BUF1 (N3112, N3107);
buf BUF1 (N3113, N3103);
xor XOR2 (N3114, N3100, N2920);
nand NAND3 (N3115, N3104, N1596, N648);
or OR3 (N3116, N3101, N2636, N1803);
nand NAND3 (N3117, N3108, N2402, N2085);
nor NOR3 (N3118, N3111, N2340, N2935);
nand NAND3 (N3119, N3115, N79, N302);
and AND4 (N3120, N3114, N1464, N1465, N1329);
nor NOR4 (N3121, N3102, N23, N2344, N443);
and AND3 (N3122, N3121, N824, N1020);
or OR2 (N3123, N3122, N1409);
not NOT1 (N3124, N3105);
not NOT1 (N3125, N3124);
not NOT1 (N3126, N3120);
or OR2 (N3127, N3118, N1806);
or OR4 (N3128, N3123, N680, N689, N1575);
and AND2 (N3129, N3116, N1596);
nand NAND2 (N3130, N3099, N2184);
not NOT1 (N3131, N3125);
xor XOR2 (N3132, N3129, N2335);
buf BUF1 (N3133, N3127);
not NOT1 (N3134, N3117);
and AND2 (N3135, N3131, N2526);
xor XOR2 (N3136, N3128, N1802);
or OR4 (N3137, N3132, N1693, N111, N1123);
and AND4 (N3138, N3133, N1452, N822, N1959);
not NOT1 (N3139, N3130);
xor XOR2 (N3140, N3119, N205);
nand NAND2 (N3141, N3134, N2428);
xor XOR2 (N3142, N3136, N1699);
nor NOR3 (N3143, N3142, N1717, N836);
xor XOR2 (N3144, N3113, N520);
buf BUF1 (N3145, N3135);
nand NAND3 (N3146, N3138, N1059, N20);
or OR4 (N3147, N3144, N888, N1353, N2558);
xor XOR2 (N3148, N3141, N1672);
not NOT1 (N3149, N3139);
nand NAND4 (N3150, N3146, N2465, N2951, N1130);
xor XOR2 (N3151, N3143, N2901);
or OR2 (N3152, N3149, N3047);
buf BUF1 (N3153, N3148);
nand NAND4 (N3154, N3145, N2248, N1575, N616);
and AND4 (N3155, N3153, N1110, N2248, N373);
and AND2 (N3156, N3137, N1173);
nor NOR2 (N3157, N3150, N163);
and AND3 (N3158, N3126, N989, N1261);
buf BUF1 (N3159, N3147);
or OR3 (N3160, N3140, N2311, N2505);
buf BUF1 (N3161, N3156);
buf BUF1 (N3162, N3158);
buf BUF1 (N3163, N3112);
buf BUF1 (N3164, N3160);
and AND2 (N3165, N3157, N1500);
nor NOR4 (N3166, N3161, N204, N2381, N2176);
xor XOR2 (N3167, N3159, N1544);
xor XOR2 (N3168, N3154, N1261);
nand NAND3 (N3169, N3166, N619, N1851);
not NOT1 (N3170, N3169);
or OR2 (N3171, N3163, N789);
not NOT1 (N3172, N3165);
not NOT1 (N3173, N3171);
or OR3 (N3174, N3172, N1183, N1921);
nor NOR2 (N3175, N3173, N2753);
xor XOR2 (N3176, N3170, N258);
nand NAND3 (N3177, N3164, N2361, N2436);
or OR4 (N3178, N3176, N2357, N2851, N2102);
or OR3 (N3179, N3174, N1713, N939);
or OR4 (N3180, N3167, N1248, N847, N1247);
nor NOR2 (N3181, N3178, N72);
or OR4 (N3182, N3155, N1986, N37, N699);
nand NAND2 (N3183, N3182, N1080);
or OR2 (N3184, N3180, N2338);
nand NAND3 (N3185, N3179, N2663, N272);
and AND2 (N3186, N3184, N2533);
buf BUF1 (N3187, N3168);
not NOT1 (N3188, N3151);
nand NAND4 (N3189, N3152, N2532, N1762, N2583);
nor NOR3 (N3190, N3175, N1712, N1558);
buf BUF1 (N3191, N3186);
and AND2 (N3192, N3188, N2727);
and AND3 (N3193, N3162, N569, N270);
or OR4 (N3194, N3190, N415, N1054, N178);
and AND2 (N3195, N3185, N696);
nor NOR2 (N3196, N3189, N2614);
not NOT1 (N3197, N3196);
buf BUF1 (N3198, N3197);
and AND2 (N3199, N3192, N3151);
or OR3 (N3200, N3187, N2664, N1709);
and AND2 (N3201, N3199, N2879);
nor NOR4 (N3202, N3183, N1368, N151, N272);
xor XOR2 (N3203, N3200, N400);
or OR4 (N3204, N3194, N3075, N2374, N2416);
buf BUF1 (N3205, N3203);
and AND2 (N3206, N3181, N138);
not NOT1 (N3207, N3201);
nand NAND4 (N3208, N3177, N2913, N2801, N628);
buf BUF1 (N3209, N3204);
xor XOR2 (N3210, N3195, N2292);
nor NOR4 (N3211, N3208, N1339, N2401, N2700);
buf BUF1 (N3212, N3198);
or OR3 (N3213, N3212, N1405, N3004);
buf BUF1 (N3214, N3207);
nor NOR4 (N3215, N3205, N2395, N404, N40);
nor NOR2 (N3216, N3211, N3089);
nor NOR3 (N3217, N3210, N293, N2476);
not NOT1 (N3218, N3213);
or OR3 (N3219, N3206, N128, N2435);
not NOT1 (N3220, N3202);
xor XOR2 (N3221, N3191, N2474);
not NOT1 (N3222, N3193);
nor NOR4 (N3223, N3217, N1266, N3051, N870);
or OR3 (N3224, N3220, N2005, N1047);
nor NOR4 (N3225, N3223, N1486, N2879, N2413);
xor XOR2 (N3226, N3225, N1270);
nand NAND4 (N3227, N3214, N1710, N2348, N1479);
nor NOR3 (N3228, N3218, N3221, N2095);
or OR2 (N3229, N1336, N2907);
xor XOR2 (N3230, N3229, N199);
buf BUF1 (N3231, N3224);
nand NAND2 (N3232, N3228, N315);
nor NOR2 (N3233, N3209, N2679);
and AND3 (N3234, N3216, N575, N2644);
and AND3 (N3235, N3215, N528, N2423);
not NOT1 (N3236, N3231);
or OR2 (N3237, N3235, N2110);
and AND2 (N3238, N3237, N1399);
not NOT1 (N3239, N3219);
and AND3 (N3240, N3238, N2586, N299);
not NOT1 (N3241, N3240);
not NOT1 (N3242, N3239);
buf BUF1 (N3243, N3226);
xor XOR2 (N3244, N3230, N3164);
buf BUF1 (N3245, N3234);
nand NAND3 (N3246, N3236, N679, N1761);
not NOT1 (N3247, N3245);
and AND2 (N3248, N3222, N2059);
xor XOR2 (N3249, N3248, N2367);
nor NOR2 (N3250, N3227, N1215);
not NOT1 (N3251, N3232);
and AND2 (N3252, N3243, N2985);
not NOT1 (N3253, N3247);
or OR4 (N3254, N3233, N435, N2403, N2458);
and AND4 (N3255, N3253, N1326, N1235, N2012);
buf BUF1 (N3256, N3241);
nor NOR3 (N3257, N3250, N911, N2987);
and AND4 (N3258, N3251, N1415, N3232, N1129);
nor NOR3 (N3259, N3252, N1278, N1322);
and AND2 (N3260, N3258, N2375);
not NOT1 (N3261, N3259);
buf BUF1 (N3262, N3261);
buf BUF1 (N3263, N3254);
and AND2 (N3264, N3244, N855);
nor NOR2 (N3265, N3242, N1305);
not NOT1 (N3266, N3263);
and AND3 (N3267, N3264, N767, N1765);
not NOT1 (N3268, N3249);
not NOT1 (N3269, N3266);
buf BUF1 (N3270, N3267);
and AND3 (N3271, N3269, N1510, N2367);
and AND4 (N3272, N3270, N2111, N1295, N3229);
or OR2 (N3273, N3271, N335);
xor XOR2 (N3274, N3268, N1811);
or OR2 (N3275, N3246, N501);
or OR3 (N3276, N3274, N2470, N1543);
buf BUF1 (N3277, N3255);
or OR2 (N3278, N3276, N660);
xor XOR2 (N3279, N3265, N2558);
not NOT1 (N3280, N3275);
or OR4 (N3281, N3257, N2591, N2988, N148);
nand NAND3 (N3282, N3260, N2824, N2482);
xor XOR2 (N3283, N3278, N902);
or OR3 (N3284, N3283, N1913, N2987);
buf BUF1 (N3285, N3277);
or OR4 (N3286, N3256, N2704, N330, N575);
not NOT1 (N3287, N3281);
and AND4 (N3288, N3280, N1194, N1570, N143);
or OR3 (N3289, N3287, N3219, N227);
nand NAND4 (N3290, N3286, N2543, N1371, N366);
buf BUF1 (N3291, N3289);
nor NOR2 (N3292, N3273, N283);
nor NOR3 (N3293, N3279, N1117, N1590);
and AND4 (N3294, N3282, N1821, N2562, N2368);
nor NOR4 (N3295, N3288, N1513, N2707, N58);
not NOT1 (N3296, N3272);
or OR4 (N3297, N3293, N253, N348, N3065);
not NOT1 (N3298, N3291);
not NOT1 (N3299, N3298);
buf BUF1 (N3300, N3296);
nor NOR3 (N3301, N3299, N543, N136);
buf BUF1 (N3302, N3284);
xor XOR2 (N3303, N3262, N2390);
or OR4 (N3304, N3295, N2879, N288, N1074);
nor NOR2 (N3305, N3294, N2228);
not NOT1 (N3306, N3302);
buf BUF1 (N3307, N3303);
and AND4 (N3308, N3290, N2615, N1967, N2265);
and AND2 (N3309, N3306, N2586);
nand NAND2 (N3310, N3307, N385);
xor XOR2 (N3311, N3310, N2885);
nor NOR4 (N3312, N3308, N2282, N1656, N1033);
and AND3 (N3313, N3297, N601, N2012);
or OR4 (N3314, N3292, N3093, N3265, N794);
xor XOR2 (N3315, N3300, N1924);
nand NAND4 (N3316, N3314, N2988, N2144, N2365);
nand NAND2 (N3317, N3301, N1682);
and AND2 (N3318, N3317, N867);
buf BUF1 (N3319, N3315);
nand NAND4 (N3320, N3311, N2596, N1125, N1980);
xor XOR2 (N3321, N3313, N1897);
or OR2 (N3322, N3305, N1290);
or OR4 (N3323, N3285, N135, N490, N1954);
or OR2 (N3324, N3312, N595);
and AND4 (N3325, N3304, N1423, N1959, N2485);
nor NOR4 (N3326, N3320, N1937, N1387, N1564);
buf BUF1 (N3327, N3316);
and AND2 (N3328, N3327, N2312);
xor XOR2 (N3329, N3324, N1365);
xor XOR2 (N3330, N3322, N2076);
and AND2 (N3331, N3326, N2778);
not NOT1 (N3332, N3323);
not NOT1 (N3333, N3318);
or OR3 (N3334, N3332, N364, N519);
nand NAND2 (N3335, N3331, N881);
xor XOR2 (N3336, N3325, N973);
buf BUF1 (N3337, N3309);
xor XOR2 (N3338, N3334, N2801);
not NOT1 (N3339, N3336);
not NOT1 (N3340, N3321);
nand NAND4 (N3341, N3339, N1039, N2430, N1594);
buf BUF1 (N3342, N3338);
not NOT1 (N3343, N3328);
not NOT1 (N3344, N3329);
not NOT1 (N3345, N3340);
buf BUF1 (N3346, N3345);
not NOT1 (N3347, N3343);
buf BUF1 (N3348, N3341);
nor NOR4 (N3349, N3319, N664, N3192, N545);
nor NOR3 (N3350, N3347, N503, N340);
nand NAND4 (N3351, N3350, N2656, N1594, N1167);
xor XOR2 (N3352, N3348, N2193);
buf BUF1 (N3353, N3342);
nor NOR2 (N3354, N3352, N939);
or OR4 (N3355, N3344, N1155, N93, N3260);
nand NAND4 (N3356, N3346, N1071, N1527, N1297);
nor NOR4 (N3357, N3349, N2322, N1621, N292);
or OR3 (N3358, N3354, N2503, N2135);
and AND4 (N3359, N3357, N527, N1475, N2811);
or OR4 (N3360, N3335, N3270, N193, N195);
or OR3 (N3361, N3353, N439, N588);
or OR2 (N3362, N3333, N1275);
nor NOR3 (N3363, N3359, N599, N1960);
nor NOR3 (N3364, N3355, N650, N255);
and AND4 (N3365, N3360, N2162, N1824, N1916);
and AND3 (N3366, N3337, N2492, N2139);
buf BUF1 (N3367, N3356);
nor NOR2 (N3368, N3366, N3309);
nor NOR2 (N3369, N3358, N2695);
nor NOR2 (N3370, N3367, N347);
nand NAND2 (N3371, N3363, N3040);
and AND4 (N3372, N3369, N482, N1515, N2575);
nand NAND2 (N3373, N3361, N1736);
or OR4 (N3374, N3372, N595, N359, N2831);
and AND2 (N3375, N3351, N2455);
nor NOR2 (N3376, N3364, N246);
xor XOR2 (N3377, N3375, N2103);
or OR3 (N3378, N3371, N2791, N541);
or OR3 (N3379, N3376, N702, N3111);
and AND4 (N3380, N3365, N2709, N790, N2061);
and AND4 (N3381, N3380, N1735, N1645, N252);
nor NOR3 (N3382, N3379, N919, N1366);
and AND2 (N3383, N3378, N1269);
xor XOR2 (N3384, N3382, N1993);
and AND2 (N3385, N3377, N1776);
nand NAND3 (N3386, N3381, N1511, N1300);
xor XOR2 (N3387, N3373, N968);
xor XOR2 (N3388, N3330, N2807);
xor XOR2 (N3389, N3368, N569);
xor XOR2 (N3390, N3384, N307);
and AND2 (N3391, N3388, N1639);
nor NOR4 (N3392, N3389, N1191, N2044, N3152);
or OR4 (N3393, N3374, N1411, N1943, N2494);
xor XOR2 (N3394, N3391, N1827);
xor XOR2 (N3395, N3385, N1379);
or OR2 (N3396, N3387, N1174);
or OR4 (N3397, N3395, N2017, N1558, N2807);
or OR3 (N3398, N3362, N1602, N3292);
nand NAND3 (N3399, N3397, N1822, N1780);
not NOT1 (N3400, N3399);
nand NAND3 (N3401, N3400, N1823, N2338);
or OR3 (N3402, N3394, N2626, N3302);
and AND4 (N3403, N3386, N1611, N3319, N2686);
and AND3 (N3404, N3390, N143, N595);
not NOT1 (N3405, N3393);
xor XOR2 (N3406, N3404, N1049);
not NOT1 (N3407, N3406);
and AND3 (N3408, N3396, N1869, N1044);
and AND2 (N3409, N3401, N2405);
and AND3 (N3410, N3383, N2515, N1928);
nor NOR2 (N3411, N3408, N77);
xor XOR2 (N3412, N3403, N1900);
not NOT1 (N3413, N3410);
buf BUF1 (N3414, N3413);
nor NOR4 (N3415, N3407, N2406, N1342, N589);
not NOT1 (N3416, N3412);
buf BUF1 (N3417, N3414);
xor XOR2 (N3418, N3405, N129);
nor NOR3 (N3419, N3411, N3362, N57);
nor NOR2 (N3420, N3392, N1647);
buf BUF1 (N3421, N3402);
nor NOR2 (N3422, N3415, N1835);
nand NAND3 (N3423, N3419, N693, N375);
not NOT1 (N3424, N3417);
nor NOR2 (N3425, N3409, N586);
nor NOR3 (N3426, N3421, N1453, N3368);
nor NOR3 (N3427, N3422, N520, N66);
not NOT1 (N3428, N3416);
or OR4 (N3429, N3428, N1811, N1206, N296);
buf BUF1 (N3430, N3398);
and AND2 (N3431, N3420, N97);
xor XOR2 (N3432, N3425, N3291);
nor NOR3 (N3433, N3430, N1161, N794);
and AND3 (N3434, N3426, N1762, N1566);
nor NOR3 (N3435, N3423, N1244, N2809);
or OR2 (N3436, N3433, N1917);
or OR2 (N3437, N3432, N2742);
nand NAND4 (N3438, N3435, N630, N2190, N1681);
nand NAND4 (N3439, N3424, N2627, N700, N1444);
nand NAND3 (N3440, N3438, N99, N2240);
or OR3 (N3441, N3439, N568, N3136);
not NOT1 (N3442, N3436);
xor XOR2 (N3443, N3427, N2689);
buf BUF1 (N3444, N3442);
nor NOR2 (N3445, N3437, N345);
nor NOR4 (N3446, N3431, N1808, N33, N2986);
not NOT1 (N3447, N3445);
nand NAND3 (N3448, N3434, N494, N1146);
buf BUF1 (N3449, N3441);
or OR4 (N3450, N3448, N87, N2867, N629);
nand NAND3 (N3451, N3449, N2921, N681);
xor XOR2 (N3452, N3440, N2338);
not NOT1 (N3453, N3450);
not NOT1 (N3454, N3418);
or OR3 (N3455, N3447, N787, N2744);
not NOT1 (N3456, N3453);
nor NOR3 (N3457, N3446, N1255, N3125);
or OR4 (N3458, N3454, N1647, N1568, N1990);
buf BUF1 (N3459, N3452);
and AND3 (N3460, N3455, N2149, N683);
nand NAND2 (N3461, N3460, N3147);
not NOT1 (N3462, N3429);
nor NOR3 (N3463, N3456, N2694, N357);
xor XOR2 (N3464, N3370, N56);
and AND2 (N3465, N3458, N767);
buf BUF1 (N3466, N3443);
or OR4 (N3467, N3457, N2979, N1651, N2096);
or OR2 (N3468, N3464, N2864);
nand NAND4 (N3469, N3459, N2084, N3412, N254);
xor XOR2 (N3470, N3461, N1797);
nand NAND2 (N3471, N3465, N2085);
buf BUF1 (N3472, N3462);
or OR2 (N3473, N3451, N171);
nor NOR3 (N3474, N3472, N474, N2474);
xor XOR2 (N3475, N3469, N2884);
not NOT1 (N3476, N3468);
buf BUF1 (N3477, N3470);
not NOT1 (N3478, N3475);
and AND3 (N3479, N3444, N1331, N368);
nor NOR2 (N3480, N3467, N2086);
and AND4 (N3481, N3463, N576, N966, N1804);
and AND2 (N3482, N3471, N933);
buf BUF1 (N3483, N3480);
buf BUF1 (N3484, N3482);
nand NAND3 (N3485, N3477, N3241, N3257);
nand NAND2 (N3486, N3466, N1518);
xor XOR2 (N3487, N3485, N72);
nand NAND4 (N3488, N3483, N787, N1896, N650);
or OR4 (N3489, N3488, N1899, N1389, N2465);
nor NOR2 (N3490, N3489, N2588);
nor NOR3 (N3491, N3487, N2414, N832);
nor NOR4 (N3492, N3481, N2088, N2977, N2670);
and AND3 (N3493, N3491, N2110, N1992);
nor NOR2 (N3494, N3484, N2128);
or OR4 (N3495, N3479, N1362, N127, N1192);
not NOT1 (N3496, N3490);
not NOT1 (N3497, N3486);
nand NAND4 (N3498, N3492, N752, N451, N1533);
nand NAND4 (N3499, N3498, N2520, N3350, N1970);
nor NOR2 (N3500, N3497, N277);
buf BUF1 (N3501, N3500);
not NOT1 (N3502, N3478);
or OR3 (N3503, N3494, N1457, N1857);
xor XOR2 (N3504, N3501, N2233);
not NOT1 (N3505, N3496);
or OR3 (N3506, N3476, N2850, N1060);
or OR4 (N3507, N3495, N362, N1087, N1781);
buf BUF1 (N3508, N3503);
not NOT1 (N3509, N3505);
buf BUF1 (N3510, N3504);
nor NOR3 (N3511, N3499, N3447, N2056);
nand NAND2 (N3512, N3493, N2476);
nand NAND4 (N3513, N3509, N1994, N555, N2278);
nand NAND4 (N3514, N3508, N803, N80, N557);
nor NOR2 (N3515, N3474, N3454);
buf BUF1 (N3516, N3473);
and AND3 (N3517, N3511, N1391, N1807);
or OR4 (N3518, N3506, N2997, N1476, N1918);
or OR3 (N3519, N3502, N2407, N2493);
endmodule