// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N1013,N989,N995,N1014,N1018,N1016,N1017,N1000,N1012,N1019;

not NOT1 (N20, N13);
not NOT1 (N21, N13);
nand NAND4 (N22, N17, N21, N9, N11);
or OR2 (N23, N9, N8);
and AND2 (N24, N4, N10);
buf BUF1 (N25, N17);
buf BUF1 (N26, N20);
not NOT1 (N27, N15);
or OR4 (N28, N26, N25, N11, N8);
or OR4 (N29, N25, N17, N25, N23);
or OR3 (N30, N10, N28, N16);
nor NOR3 (N31, N8, N21, N12);
nand NAND3 (N32, N13, N1, N1);
xor XOR2 (N33, N1, N21);
and AND3 (N34, N18, N29, N31);
and AND2 (N35, N29, N23);
nor NOR2 (N36, N9, N25);
nor NOR3 (N37, N36, N11, N5);
buf BUF1 (N38, N29);
buf BUF1 (N39, N35);
not NOT1 (N40, N38);
buf BUF1 (N41, N24);
nand NAND4 (N42, N40, N40, N21, N9);
or OR3 (N43, N22, N11, N39);
xor XOR2 (N44, N16, N18);
not NOT1 (N45, N33);
nand NAND3 (N46, N30, N36, N16);
xor XOR2 (N47, N34, N6);
or OR4 (N48, N47, N26, N24, N3);
nor NOR4 (N49, N44, N3, N45, N20);
nor NOR3 (N50, N47, N43, N6);
buf BUF1 (N51, N28);
xor XOR2 (N52, N37, N33);
and AND4 (N53, N27, N27, N1, N4);
nand NAND3 (N54, N41, N22, N38);
nor NOR2 (N55, N50, N36);
and AND3 (N56, N49, N16, N43);
and AND2 (N57, N56, N46);
or OR4 (N58, N22, N38, N45, N23);
nor NOR4 (N59, N55, N20, N46, N1);
nand NAND4 (N60, N58, N55, N33, N42);
nor NOR4 (N61, N50, N9, N47, N16);
nand NAND3 (N62, N57, N50, N21);
nand NAND3 (N63, N62, N49, N25);
nor NOR3 (N64, N59, N53, N19);
nor NOR2 (N65, N41, N24);
not NOT1 (N66, N51);
nand NAND2 (N67, N60, N56);
not NOT1 (N68, N67);
xor XOR2 (N69, N64, N53);
nor NOR2 (N70, N61, N33);
nor NOR3 (N71, N52, N44, N39);
nor NOR3 (N72, N32, N17, N23);
and AND4 (N73, N71, N16, N31, N68);
buf BUF1 (N74, N34);
xor XOR2 (N75, N66, N37);
buf BUF1 (N76, N65);
nand NAND2 (N77, N74, N11);
nor NOR4 (N78, N75, N7, N66, N67);
xor XOR2 (N79, N70, N61);
nor NOR2 (N80, N72, N75);
xor XOR2 (N81, N54, N76);
nor NOR3 (N82, N74, N48, N13);
not NOT1 (N83, N56);
nor NOR3 (N84, N77, N77, N44);
buf BUF1 (N85, N78);
xor XOR2 (N86, N80, N15);
not NOT1 (N87, N69);
not NOT1 (N88, N87);
xor XOR2 (N89, N84, N24);
nor NOR3 (N90, N83, N58, N34);
nor NOR2 (N91, N85, N49);
xor XOR2 (N92, N82, N56);
not NOT1 (N93, N89);
not NOT1 (N94, N86);
nand NAND3 (N95, N81, N45, N30);
buf BUF1 (N96, N94);
buf BUF1 (N97, N88);
buf BUF1 (N98, N90);
buf BUF1 (N99, N95);
or OR3 (N100, N91, N46, N70);
and AND4 (N101, N93, N63, N43, N56);
buf BUF1 (N102, N89);
and AND4 (N103, N79, N21, N69, N48);
xor XOR2 (N104, N73, N54);
not NOT1 (N105, N96);
buf BUF1 (N106, N102);
nor NOR2 (N107, N105, N87);
or OR4 (N108, N99, N77, N81, N101);
buf BUF1 (N109, N60);
or OR4 (N110, N98, N77, N67, N44);
nand NAND4 (N111, N92, N5, N24, N72);
or OR4 (N112, N110, N46, N15, N3);
not NOT1 (N113, N111);
nand NAND2 (N114, N113, N1);
nor NOR3 (N115, N97, N62, N64);
nor NOR3 (N116, N115, N75, N49);
nor NOR2 (N117, N114, N61);
and AND4 (N118, N117, N109, N57, N48);
nor NOR3 (N119, N56, N4, N107);
or OR4 (N120, N42, N6, N71, N24);
and AND2 (N121, N120, N84);
and AND2 (N122, N106, N48);
or OR3 (N123, N119, N122, N112);
or OR3 (N124, N30, N120, N100);
or OR4 (N125, N2, N72, N61, N69);
not NOT1 (N126, N4);
xor XOR2 (N127, N123, N47);
xor XOR2 (N128, N124, N84);
buf BUF1 (N129, N127);
xor XOR2 (N130, N103, N124);
xor XOR2 (N131, N128, N90);
xor XOR2 (N132, N131, N43);
not NOT1 (N133, N121);
xor XOR2 (N134, N116, N60);
xor XOR2 (N135, N129, N20);
buf BUF1 (N136, N104);
or OR3 (N137, N118, N78, N42);
buf BUF1 (N138, N132);
and AND3 (N139, N133, N33, N118);
xor XOR2 (N140, N139, N113);
buf BUF1 (N141, N136);
buf BUF1 (N142, N134);
or OR3 (N143, N108, N8, N75);
nor NOR3 (N144, N140, N31, N8);
nor NOR2 (N145, N142, N122);
xor XOR2 (N146, N135, N18);
nand NAND3 (N147, N143, N72, N55);
nor NOR4 (N148, N146, N49, N91, N24);
not NOT1 (N149, N148);
nor NOR4 (N150, N125, N89, N38, N34);
and AND3 (N151, N145, N116, N38);
not NOT1 (N152, N147);
or OR2 (N153, N149, N70);
and AND2 (N154, N144, N4);
nor NOR4 (N155, N141, N124, N12, N100);
not NOT1 (N156, N126);
not NOT1 (N157, N138);
nor NOR3 (N158, N157, N139, N61);
not NOT1 (N159, N150);
xor XOR2 (N160, N151, N104);
or OR3 (N161, N137, N137, N35);
and AND3 (N162, N160, N94, N58);
and AND3 (N163, N159, N69, N10);
nor NOR3 (N164, N162, N129, N8);
not NOT1 (N165, N130);
nand NAND2 (N166, N165, N70);
and AND4 (N167, N152, N77, N77, N75);
nor NOR3 (N168, N167, N44, N155);
buf BUF1 (N169, N129);
nand NAND2 (N170, N164, N25);
not NOT1 (N171, N169);
or OR2 (N172, N171, N142);
or OR3 (N173, N156, N117, N36);
buf BUF1 (N174, N163);
nor NOR4 (N175, N153, N78, N49, N9);
nand NAND2 (N176, N172, N170);
buf BUF1 (N177, N172);
xor XOR2 (N178, N168, N10);
nor NOR2 (N179, N173, N32);
not NOT1 (N180, N176);
nand NAND2 (N181, N166, N99);
nand NAND3 (N182, N178, N78, N113);
not NOT1 (N183, N154);
or OR2 (N184, N183, N119);
and AND3 (N185, N177, N28, N19);
or OR2 (N186, N180, N106);
nor NOR2 (N187, N186, N11);
nor NOR2 (N188, N182, N16);
xor XOR2 (N189, N187, N117);
not NOT1 (N190, N184);
buf BUF1 (N191, N174);
and AND4 (N192, N190, N84, N117, N59);
nor NOR4 (N193, N192, N13, N159, N110);
buf BUF1 (N194, N181);
or OR2 (N195, N189, N101);
not NOT1 (N196, N158);
and AND3 (N197, N193, N57, N183);
and AND2 (N198, N195, N92);
and AND3 (N199, N194, N170, N174);
or OR2 (N200, N161, N104);
and AND2 (N201, N175, N165);
not NOT1 (N202, N198);
and AND3 (N203, N202, N18, N180);
not NOT1 (N204, N188);
and AND2 (N205, N200, N89);
or OR4 (N206, N205, N198, N19, N96);
xor XOR2 (N207, N185, N29);
or OR4 (N208, N197, N136, N190, N103);
xor XOR2 (N209, N199, N19);
and AND3 (N210, N206, N161, N84);
nand NAND3 (N211, N204, N126, N120);
and AND2 (N212, N203, N167);
or OR3 (N213, N179, N153, N66);
not NOT1 (N214, N213);
or OR3 (N215, N210, N29, N182);
or OR4 (N216, N196, N157, N130, N192);
nand NAND2 (N217, N216, N129);
buf BUF1 (N218, N191);
xor XOR2 (N219, N212, N113);
buf BUF1 (N220, N219);
xor XOR2 (N221, N209, N153);
not NOT1 (N222, N218);
nand NAND2 (N223, N220, N176);
nand NAND2 (N224, N223, N128);
buf BUF1 (N225, N214);
or OR3 (N226, N224, N154, N165);
not NOT1 (N227, N207);
xor XOR2 (N228, N208, N48);
not NOT1 (N229, N221);
and AND3 (N230, N227, N133, N21);
xor XOR2 (N231, N211, N208);
nor NOR2 (N232, N217, N1);
buf BUF1 (N233, N228);
nand NAND2 (N234, N230, N63);
nor NOR4 (N235, N225, N105, N81, N140);
not NOT1 (N236, N234);
nand NAND3 (N237, N201, N132, N51);
not NOT1 (N238, N231);
nand NAND3 (N239, N232, N230, N183);
not NOT1 (N240, N226);
xor XOR2 (N241, N215, N145);
buf BUF1 (N242, N235);
xor XOR2 (N243, N229, N62);
not NOT1 (N244, N233);
or OR4 (N245, N243, N93, N61, N126);
and AND2 (N246, N245, N60);
nand NAND3 (N247, N244, N206, N226);
xor XOR2 (N248, N247, N26);
xor XOR2 (N249, N241, N138);
or OR4 (N250, N246, N74, N246, N237);
buf BUF1 (N251, N2);
not NOT1 (N252, N240);
buf BUF1 (N253, N236);
nor NOR2 (N254, N253, N3);
buf BUF1 (N255, N251);
or OR4 (N256, N248, N51, N102, N62);
and AND4 (N257, N255, N132, N196, N168);
nor NOR2 (N258, N222, N117);
and AND2 (N259, N250, N54);
or OR4 (N260, N258, N136, N217, N179);
nor NOR3 (N261, N239, N42, N231);
nor NOR3 (N262, N261, N189, N13);
buf BUF1 (N263, N254);
or OR4 (N264, N249, N130, N256, N202);
or OR3 (N265, N80, N90, N121);
or OR2 (N266, N257, N184);
nor NOR2 (N267, N263, N203);
not NOT1 (N268, N242);
xor XOR2 (N269, N262, N200);
not NOT1 (N270, N238);
not NOT1 (N271, N259);
xor XOR2 (N272, N269, N253);
nand NAND3 (N273, N264, N179, N246);
or OR3 (N274, N273, N235, N261);
or OR2 (N275, N260, N94);
and AND2 (N276, N265, N251);
and AND4 (N277, N274, N116, N58, N169);
xor XOR2 (N278, N252, N75);
not NOT1 (N279, N271);
nand NAND3 (N280, N268, N191, N131);
xor XOR2 (N281, N278, N177);
buf BUF1 (N282, N270);
nor NOR4 (N283, N280, N160, N276, N204);
xor XOR2 (N284, N253, N77);
and AND2 (N285, N275, N250);
buf BUF1 (N286, N284);
and AND2 (N287, N266, N68);
nor NOR3 (N288, N267, N256, N235);
or OR2 (N289, N277, N146);
not NOT1 (N290, N288);
nand NAND4 (N291, N281, N96, N138, N276);
nand NAND3 (N292, N287, N279, N165);
xor XOR2 (N293, N283, N175);
xor XOR2 (N294, N159, N225);
buf BUF1 (N295, N292);
nand NAND2 (N296, N290, N214);
nor NOR4 (N297, N294, N171, N81, N118);
and AND3 (N298, N297, N195, N280);
buf BUF1 (N299, N296);
and AND3 (N300, N293, N100, N233);
not NOT1 (N301, N300);
and AND3 (N302, N282, N156, N196);
or OR3 (N303, N302, N287, N150);
buf BUF1 (N304, N291);
or OR4 (N305, N286, N169, N113, N100);
and AND2 (N306, N285, N233);
nand NAND3 (N307, N299, N24, N285);
not NOT1 (N308, N295);
nand NAND3 (N309, N289, N260, N65);
not NOT1 (N310, N301);
and AND3 (N311, N307, N196, N35);
or OR3 (N312, N310, N227, N84);
nor NOR4 (N313, N304, N310, N270, N311);
not NOT1 (N314, N88);
buf BUF1 (N315, N314);
xor XOR2 (N316, N306, N292);
buf BUF1 (N317, N309);
nand NAND4 (N318, N313, N17, N81, N296);
nand NAND3 (N319, N272, N38, N73);
and AND3 (N320, N312, N290, N222);
or OR2 (N321, N315, N276);
nor NOR2 (N322, N316, N231);
nor NOR3 (N323, N321, N78, N267);
buf BUF1 (N324, N303);
xor XOR2 (N325, N317, N140);
not NOT1 (N326, N322);
buf BUF1 (N327, N325);
nor NOR2 (N328, N305, N258);
and AND4 (N329, N327, N233, N102, N299);
or OR4 (N330, N320, N318, N211, N106);
or OR4 (N331, N220, N327, N315, N2);
and AND2 (N332, N308, N203);
nand NAND3 (N333, N328, N145, N187);
nand NAND3 (N334, N319, N171, N9);
nand NAND3 (N335, N331, N148, N72);
xor XOR2 (N336, N335, N95);
buf BUF1 (N337, N323);
not NOT1 (N338, N326);
not NOT1 (N339, N324);
nor NOR3 (N340, N337, N157, N137);
not NOT1 (N341, N334);
or OR4 (N342, N333, N184, N149, N174);
not NOT1 (N343, N340);
nand NAND4 (N344, N342, N107, N17, N301);
nand NAND2 (N345, N329, N187);
xor XOR2 (N346, N339, N253);
and AND3 (N347, N343, N60, N47);
not NOT1 (N348, N341);
buf BUF1 (N349, N347);
xor XOR2 (N350, N330, N201);
buf BUF1 (N351, N336);
buf BUF1 (N352, N351);
and AND2 (N353, N346, N37);
nand NAND4 (N354, N332, N291, N26, N139);
buf BUF1 (N355, N348);
xor XOR2 (N356, N298, N304);
nor NOR2 (N357, N355, N32);
xor XOR2 (N358, N349, N333);
and AND3 (N359, N353, N101, N197);
buf BUF1 (N360, N344);
nor NOR2 (N361, N360, N211);
and AND4 (N362, N352, N17, N97, N227);
or OR2 (N363, N362, N107);
nand NAND2 (N364, N363, N322);
not NOT1 (N365, N338);
nand NAND4 (N366, N357, N21, N140, N36);
and AND4 (N367, N361, N254, N200, N151);
nand NAND4 (N368, N356, N211, N53, N96);
buf BUF1 (N369, N365);
nand NAND2 (N370, N354, N224);
or OR3 (N371, N350, N249, N218);
and AND2 (N372, N371, N348);
and AND2 (N373, N358, N126);
nand NAND2 (N374, N368, N165);
nand NAND3 (N375, N359, N274, N374);
and AND4 (N376, N360, N77, N43, N316);
not NOT1 (N377, N376);
xor XOR2 (N378, N372, N167);
or OR3 (N379, N364, N373, N47);
or OR2 (N380, N239, N343);
not NOT1 (N381, N375);
and AND2 (N382, N379, N82);
nor NOR2 (N383, N366, N264);
or OR2 (N384, N383, N167);
or OR2 (N385, N378, N240);
not NOT1 (N386, N385);
nor NOR2 (N387, N367, N90);
and AND2 (N388, N386, N120);
nor NOR3 (N389, N380, N257, N226);
nand NAND3 (N390, N389, N197, N363);
xor XOR2 (N391, N382, N344);
not NOT1 (N392, N369);
nand NAND4 (N393, N377, N247, N333, N125);
buf BUF1 (N394, N391);
nand NAND4 (N395, N370, N20, N270, N113);
buf BUF1 (N396, N393);
nor NOR2 (N397, N384, N40);
nor NOR2 (N398, N396, N280);
nand NAND3 (N399, N397, N282, N290);
or OR2 (N400, N399, N131);
nor NOR4 (N401, N388, N13, N325, N226);
nor NOR2 (N402, N394, N318);
and AND3 (N403, N345, N303, N229);
xor XOR2 (N404, N390, N383);
buf BUF1 (N405, N404);
buf BUF1 (N406, N405);
not NOT1 (N407, N381);
nand NAND2 (N408, N401, N190);
not NOT1 (N409, N400);
nand NAND2 (N410, N398, N372);
and AND4 (N411, N403, N387, N345, N219);
or OR2 (N412, N161, N207);
not NOT1 (N413, N412);
xor XOR2 (N414, N408, N31);
xor XOR2 (N415, N413, N264);
nand NAND4 (N416, N409, N405, N191, N47);
or OR4 (N417, N411, N407, N343, N109);
nor NOR4 (N418, N279, N231, N31, N83);
or OR3 (N419, N414, N265, N131);
buf BUF1 (N420, N406);
buf BUF1 (N421, N410);
not NOT1 (N422, N420);
nor NOR3 (N423, N418, N222, N68);
buf BUF1 (N424, N423);
nand NAND4 (N425, N402, N255, N353, N226);
nor NOR2 (N426, N395, N114);
not NOT1 (N427, N426);
buf BUF1 (N428, N421);
buf BUF1 (N429, N424);
nor NOR4 (N430, N429, N291, N233, N145);
and AND3 (N431, N417, N21, N283);
xor XOR2 (N432, N428, N170);
not NOT1 (N433, N392);
and AND3 (N434, N430, N334, N120);
or OR4 (N435, N416, N18, N245, N208);
nand NAND2 (N436, N419, N249);
or OR4 (N437, N432, N185, N380, N290);
buf BUF1 (N438, N415);
not NOT1 (N439, N431);
xor XOR2 (N440, N437, N79);
xor XOR2 (N441, N439, N130);
nor NOR3 (N442, N422, N441, N375);
buf BUF1 (N443, N134);
not NOT1 (N444, N427);
nor NOR2 (N445, N435, N325);
or OR2 (N446, N443, N152);
or OR3 (N447, N433, N85, N407);
nor NOR3 (N448, N440, N170, N222);
and AND3 (N449, N442, N54, N177);
or OR3 (N450, N434, N305, N374);
or OR2 (N451, N436, N195);
and AND3 (N452, N445, N181, N150);
buf BUF1 (N453, N452);
not NOT1 (N454, N446);
xor XOR2 (N455, N450, N80);
and AND2 (N456, N451, N373);
nand NAND3 (N457, N454, N106, N27);
and AND4 (N458, N453, N420, N280, N51);
xor XOR2 (N459, N448, N219);
nor NOR2 (N460, N425, N69);
nor NOR2 (N461, N457, N341);
and AND2 (N462, N456, N271);
or OR4 (N463, N459, N249, N316, N2);
buf BUF1 (N464, N438);
buf BUF1 (N465, N458);
and AND3 (N466, N455, N129, N271);
not NOT1 (N467, N463);
not NOT1 (N468, N447);
or OR3 (N469, N461, N28, N12);
and AND3 (N470, N464, N181, N221);
nor NOR2 (N471, N444, N28);
nand NAND4 (N472, N449, N441, N183, N65);
nand NAND3 (N473, N469, N119, N60);
nand NAND4 (N474, N470, N378, N83, N340);
nand NAND3 (N475, N473, N83, N353);
not NOT1 (N476, N462);
not NOT1 (N477, N474);
xor XOR2 (N478, N466, N25);
nand NAND3 (N479, N467, N159, N53);
and AND4 (N480, N476, N103, N66, N76);
and AND2 (N481, N471, N74);
or OR3 (N482, N475, N411, N438);
xor XOR2 (N483, N460, N165);
xor XOR2 (N484, N465, N37);
xor XOR2 (N485, N484, N469);
nand NAND2 (N486, N485, N10);
and AND2 (N487, N468, N145);
nor NOR3 (N488, N472, N333, N16);
buf BUF1 (N489, N482);
nand NAND3 (N490, N487, N253, N330);
buf BUF1 (N491, N478);
or OR4 (N492, N480, N444, N87, N483);
not NOT1 (N493, N55);
and AND2 (N494, N490, N159);
nor NOR4 (N495, N491, N352, N448, N234);
buf BUF1 (N496, N481);
and AND4 (N497, N495, N355, N117, N317);
or OR2 (N498, N497, N70);
and AND2 (N499, N493, N222);
nand NAND4 (N500, N486, N8, N64, N42);
not NOT1 (N501, N477);
or OR2 (N502, N488, N39);
not NOT1 (N503, N494);
and AND4 (N504, N479, N1, N325, N294);
nand NAND4 (N505, N489, N160, N44, N484);
nor NOR3 (N506, N504, N93, N415);
xor XOR2 (N507, N506, N426);
or OR4 (N508, N500, N38, N474, N275);
nor NOR3 (N509, N492, N240, N195);
or OR2 (N510, N498, N387);
not NOT1 (N511, N505);
nor NOR3 (N512, N508, N408, N244);
or OR4 (N513, N511, N512, N80, N352);
not NOT1 (N514, N469);
and AND3 (N515, N496, N476, N168);
nor NOR2 (N516, N501, N252);
and AND2 (N517, N499, N489);
xor XOR2 (N518, N516, N102);
and AND4 (N519, N513, N17, N180, N341);
not NOT1 (N520, N514);
nand NAND2 (N521, N520, N423);
not NOT1 (N522, N517);
nand NAND2 (N523, N502, N219);
xor XOR2 (N524, N518, N401);
xor XOR2 (N525, N503, N212);
nor NOR2 (N526, N524, N356);
and AND4 (N527, N526, N482, N180, N43);
or OR3 (N528, N525, N449, N16);
not NOT1 (N529, N509);
or OR3 (N530, N521, N98, N21);
or OR4 (N531, N515, N190, N307, N156);
or OR2 (N532, N529, N352);
nand NAND3 (N533, N531, N222, N188);
nand NAND2 (N534, N507, N57);
not NOT1 (N535, N528);
nand NAND3 (N536, N519, N353, N346);
xor XOR2 (N537, N536, N26);
not NOT1 (N538, N535);
nand NAND2 (N539, N523, N208);
and AND4 (N540, N522, N65, N63, N448);
not NOT1 (N541, N510);
nor NOR4 (N542, N540, N346, N394, N396);
not NOT1 (N543, N542);
or OR2 (N544, N527, N99);
nand NAND3 (N545, N544, N110, N228);
xor XOR2 (N546, N530, N393);
nor NOR4 (N547, N534, N480, N464, N429);
or OR2 (N548, N543, N479);
nor NOR3 (N549, N548, N534, N212);
xor XOR2 (N550, N546, N528);
nand NAND2 (N551, N545, N427);
and AND3 (N552, N533, N157, N242);
not NOT1 (N553, N552);
and AND2 (N554, N537, N92);
nand NAND4 (N555, N550, N87, N256, N364);
not NOT1 (N556, N555);
nor NOR4 (N557, N549, N378, N251, N524);
or OR4 (N558, N538, N206, N438, N425);
not NOT1 (N559, N551);
or OR3 (N560, N556, N218, N97);
nor NOR4 (N561, N554, N60, N554, N79);
buf BUF1 (N562, N553);
buf BUF1 (N563, N561);
and AND3 (N564, N562, N385, N325);
nor NOR3 (N565, N559, N84, N192);
and AND4 (N566, N560, N481, N66, N292);
buf BUF1 (N567, N564);
xor XOR2 (N568, N532, N38);
nor NOR3 (N569, N563, N7, N290);
xor XOR2 (N570, N557, N9);
buf BUF1 (N571, N568);
nor NOR4 (N572, N571, N121, N429, N221);
nand NAND2 (N573, N572, N289);
and AND4 (N574, N565, N219, N482, N10);
xor XOR2 (N575, N574, N308);
nor NOR3 (N576, N566, N205, N304);
not NOT1 (N577, N570);
or OR4 (N578, N577, N347, N384, N118);
buf BUF1 (N579, N573);
buf BUF1 (N580, N539);
xor XOR2 (N581, N576, N345);
or OR3 (N582, N578, N52, N387);
buf BUF1 (N583, N547);
xor XOR2 (N584, N582, N496);
xor XOR2 (N585, N579, N485);
or OR2 (N586, N575, N230);
xor XOR2 (N587, N558, N562);
nor NOR3 (N588, N580, N37, N520);
buf BUF1 (N589, N584);
nand NAND3 (N590, N541, N395, N288);
or OR2 (N591, N586, N469);
nor NOR3 (N592, N569, N38, N252);
xor XOR2 (N593, N585, N98);
nor NOR4 (N594, N591, N206, N565, N462);
nor NOR3 (N595, N592, N471, N163);
xor XOR2 (N596, N590, N280);
and AND2 (N597, N567, N31);
and AND2 (N598, N595, N85);
not NOT1 (N599, N593);
and AND2 (N600, N587, N419);
and AND2 (N601, N594, N560);
or OR3 (N602, N589, N232, N485);
not NOT1 (N603, N602);
nand NAND2 (N604, N599, N50);
xor XOR2 (N605, N598, N198);
buf BUF1 (N606, N583);
buf BUF1 (N607, N588);
nand NAND2 (N608, N603, N339);
nor NOR3 (N609, N601, N294, N258);
nor NOR4 (N610, N606, N506, N110, N334);
not NOT1 (N611, N607);
nand NAND2 (N612, N597, N323);
or OR4 (N613, N600, N511, N228, N34);
not NOT1 (N614, N581);
or OR4 (N615, N613, N30, N411, N613);
nand NAND4 (N616, N611, N401, N22, N313);
xor XOR2 (N617, N614, N440);
or OR4 (N618, N604, N544, N40, N459);
nor NOR4 (N619, N612, N397, N552, N274);
or OR3 (N620, N615, N124, N288);
xor XOR2 (N621, N608, N164);
or OR3 (N622, N619, N414, N16);
nand NAND4 (N623, N609, N227, N385, N9);
nand NAND3 (N624, N618, N185, N500);
nor NOR2 (N625, N622, N191);
and AND4 (N626, N596, N445, N507, N199);
nor NOR2 (N627, N610, N239);
xor XOR2 (N628, N620, N543);
buf BUF1 (N629, N627);
not NOT1 (N630, N621);
buf BUF1 (N631, N628);
or OR4 (N632, N631, N531, N428, N287);
or OR3 (N633, N632, N623, N589);
not NOT1 (N634, N609);
buf BUF1 (N635, N629);
or OR2 (N636, N633, N233);
or OR4 (N637, N624, N145, N435, N265);
and AND3 (N638, N637, N636, N330);
or OR2 (N639, N529, N606);
nand NAND2 (N640, N634, N327);
xor XOR2 (N641, N616, N553);
nor NOR3 (N642, N630, N507, N444);
not NOT1 (N643, N639);
xor XOR2 (N644, N605, N69);
buf BUF1 (N645, N641);
nand NAND2 (N646, N644, N331);
or OR4 (N647, N626, N625, N512, N141);
nand NAND2 (N648, N561, N560);
or OR2 (N649, N617, N372);
not NOT1 (N650, N645);
and AND4 (N651, N650, N222, N12, N203);
nor NOR4 (N652, N651, N555, N70, N340);
nor NOR3 (N653, N635, N13, N219);
not NOT1 (N654, N648);
and AND3 (N655, N652, N278, N409);
nand NAND4 (N656, N642, N97, N498, N281);
and AND4 (N657, N647, N375, N181, N133);
and AND3 (N658, N638, N627, N568);
nor NOR2 (N659, N640, N499);
nor NOR3 (N660, N656, N132, N84);
or OR4 (N661, N643, N504, N424, N250);
or OR3 (N662, N661, N295, N308);
and AND3 (N663, N653, N134, N359);
nand NAND4 (N664, N655, N491, N302, N281);
or OR4 (N665, N658, N263, N100, N557);
and AND2 (N666, N649, N141);
or OR2 (N667, N662, N166);
or OR2 (N668, N660, N266);
or OR3 (N669, N657, N567, N589);
buf BUF1 (N670, N664);
or OR4 (N671, N646, N519, N402, N227);
xor XOR2 (N672, N666, N574);
not NOT1 (N673, N671);
not NOT1 (N674, N659);
or OR4 (N675, N669, N53, N165, N116);
nand NAND2 (N676, N667, N569);
buf BUF1 (N677, N663);
nor NOR3 (N678, N654, N384, N213);
buf BUF1 (N679, N668);
buf BUF1 (N680, N670);
xor XOR2 (N681, N665, N413);
and AND4 (N682, N675, N613, N648, N338);
nand NAND4 (N683, N681, N445, N199, N604);
or OR4 (N684, N679, N475, N683, N596);
xor XOR2 (N685, N271, N178);
xor XOR2 (N686, N676, N130);
or OR4 (N687, N674, N319, N110, N324);
buf BUF1 (N688, N682);
nor NOR4 (N689, N673, N673, N104, N561);
buf BUF1 (N690, N688);
buf BUF1 (N691, N687);
xor XOR2 (N692, N689, N560);
xor XOR2 (N693, N685, N173);
buf BUF1 (N694, N677);
buf BUF1 (N695, N694);
buf BUF1 (N696, N678);
nand NAND4 (N697, N686, N41, N558, N644);
buf BUF1 (N698, N695);
or OR2 (N699, N680, N574);
buf BUF1 (N700, N691);
buf BUF1 (N701, N698);
nand NAND4 (N702, N692, N45, N502, N218);
buf BUF1 (N703, N697);
buf BUF1 (N704, N684);
not NOT1 (N705, N703);
xor XOR2 (N706, N672, N641);
and AND2 (N707, N705, N380);
not NOT1 (N708, N701);
and AND3 (N709, N704, N37, N126);
not NOT1 (N710, N708);
or OR3 (N711, N709, N76, N73);
buf BUF1 (N712, N702);
nand NAND3 (N713, N690, N511, N534);
nor NOR3 (N714, N710, N204, N361);
nand NAND2 (N715, N696, N595);
nor NOR4 (N716, N700, N30, N493, N105);
nand NAND3 (N717, N706, N273, N60);
or OR4 (N718, N714, N443, N113, N312);
or OR3 (N719, N713, N662, N334);
and AND4 (N720, N717, N178, N658, N86);
not NOT1 (N721, N718);
buf BUF1 (N722, N711);
or OR3 (N723, N720, N586, N656);
xor XOR2 (N724, N716, N653);
buf BUF1 (N725, N699);
or OR2 (N726, N721, N72);
not NOT1 (N727, N693);
not NOT1 (N728, N715);
nand NAND2 (N729, N722, N494);
nand NAND4 (N730, N726, N53, N655, N212);
and AND4 (N731, N729, N311, N73, N369);
or OR2 (N732, N712, N713);
not NOT1 (N733, N723);
nand NAND4 (N734, N727, N630, N521, N304);
nor NOR2 (N735, N733, N687);
or OR3 (N736, N731, N141, N57);
and AND4 (N737, N719, N499, N146, N713);
and AND4 (N738, N732, N247, N447, N16);
and AND4 (N739, N707, N536, N161, N466);
nand NAND4 (N740, N734, N191, N106, N522);
or OR4 (N741, N737, N9, N498, N326);
buf BUF1 (N742, N738);
nand NAND4 (N743, N728, N657, N229, N404);
not NOT1 (N744, N725);
nand NAND2 (N745, N741, N230);
not NOT1 (N746, N740);
nor NOR2 (N747, N742, N690);
not NOT1 (N748, N744);
not NOT1 (N749, N746);
or OR3 (N750, N730, N401, N282);
nand NAND2 (N751, N747, N317);
nand NAND2 (N752, N748, N743);
nand NAND4 (N753, N580, N250, N185, N680);
xor XOR2 (N754, N749, N562);
and AND4 (N755, N736, N19, N663, N2);
not NOT1 (N756, N745);
and AND4 (N757, N751, N353, N243, N257);
buf BUF1 (N758, N754);
or OR3 (N759, N739, N27, N388);
or OR2 (N760, N755, N619);
xor XOR2 (N761, N759, N217);
and AND2 (N762, N752, N725);
not NOT1 (N763, N724);
and AND2 (N764, N735, N430);
and AND4 (N765, N753, N294, N273, N540);
buf BUF1 (N766, N764);
nor NOR2 (N767, N757, N178);
and AND2 (N768, N756, N157);
or OR4 (N769, N760, N126, N52, N660);
and AND4 (N770, N769, N675, N291, N442);
nor NOR3 (N771, N762, N217, N392);
nand NAND4 (N772, N771, N576, N29, N578);
not NOT1 (N773, N765);
xor XOR2 (N774, N768, N599);
nand NAND3 (N775, N770, N217, N275);
xor XOR2 (N776, N773, N752);
nor NOR2 (N777, N766, N90);
and AND4 (N778, N761, N524, N345, N585);
not NOT1 (N779, N763);
nor NOR4 (N780, N776, N741, N406, N415);
xor XOR2 (N781, N775, N136);
nand NAND4 (N782, N777, N489, N465, N182);
xor XOR2 (N783, N780, N11);
not NOT1 (N784, N779);
nor NOR4 (N785, N758, N649, N315, N404);
nand NAND4 (N786, N767, N386, N428, N484);
xor XOR2 (N787, N785, N237);
buf BUF1 (N788, N782);
buf BUF1 (N789, N786);
and AND2 (N790, N788, N770);
nor NOR3 (N791, N778, N488, N721);
and AND2 (N792, N750, N538);
nand NAND4 (N793, N783, N689, N278, N546);
not NOT1 (N794, N772);
xor XOR2 (N795, N784, N501);
xor XOR2 (N796, N795, N629);
nor NOR3 (N797, N790, N224, N361);
buf BUF1 (N798, N789);
buf BUF1 (N799, N791);
and AND4 (N800, N796, N345, N358, N440);
xor XOR2 (N801, N799, N599);
or OR4 (N802, N798, N33, N215, N466);
not NOT1 (N803, N793);
not NOT1 (N804, N787);
buf BUF1 (N805, N792);
or OR3 (N806, N803, N756, N75);
nand NAND3 (N807, N806, N171, N668);
nor NOR2 (N808, N797, N450);
xor XOR2 (N809, N781, N678);
xor XOR2 (N810, N800, N512);
xor XOR2 (N811, N809, N553);
not NOT1 (N812, N805);
nor NOR3 (N813, N811, N689, N251);
nand NAND2 (N814, N807, N580);
nand NAND3 (N815, N794, N790, N455);
nor NOR4 (N816, N814, N152, N644, N264);
xor XOR2 (N817, N804, N12);
and AND2 (N818, N801, N157);
nor NOR2 (N819, N818, N676);
or OR2 (N820, N815, N776);
nand NAND3 (N821, N808, N3, N39);
or OR2 (N822, N813, N113);
buf BUF1 (N823, N802);
not NOT1 (N824, N810);
and AND3 (N825, N817, N562, N568);
not NOT1 (N826, N820);
or OR2 (N827, N826, N294);
not NOT1 (N828, N821);
nor NOR2 (N829, N825, N471);
xor XOR2 (N830, N823, N178);
not NOT1 (N831, N830);
and AND4 (N832, N824, N260, N472, N235);
nor NOR2 (N833, N812, N625);
or OR4 (N834, N833, N98, N62, N318);
and AND2 (N835, N832, N357);
not NOT1 (N836, N834);
buf BUF1 (N837, N829);
buf BUF1 (N838, N828);
nor NOR4 (N839, N835, N251, N517, N217);
or OR3 (N840, N774, N29, N387);
or OR3 (N841, N838, N346, N609);
nand NAND2 (N842, N819, N538);
nand NAND3 (N843, N839, N778, N47);
not NOT1 (N844, N837);
not NOT1 (N845, N844);
xor XOR2 (N846, N843, N516);
or OR4 (N847, N841, N544, N147, N496);
and AND2 (N848, N847, N359);
buf BUF1 (N849, N845);
not NOT1 (N850, N842);
buf BUF1 (N851, N840);
not NOT1 (N852, N851);
buf BUF1 (N853, N836);
xor XOR2 (N854, N848, N330);
xor XOR2 (N855, N854, N499);
not NOT1 (N856, N852);
nand NAND2 (N857, N827, N773);
buf BUF1 (N858, N831);
not NOT1 (N859, N857);
buf BUF1 (N860, N856);
nor NOR4 (N861, N860, N826, N796, N739);
not NOT1 (N862, N858);
nor NOR2 (N863, N816, N11);
nor NOR4 (N864, N855, N516, N389, N475);
nor NOR4 (N865, N846, N35, N698, N333);
xor XOR2 (N866, N822, N827);
nor NOR4 (N867, N849, N710, N704, N452);
or OR4 (N868, N859, N579, N747, N787);
buf BUF1 (N869, N865);
nand NAND2 (N870, N868, N311);
not NOT1 (N871, N850);
or OR2 (N872, N871, N59);
not NOT1 (N873, N864);
nand NAND4 (N874, N869, N27, N485, N512);
nand NAND3 (N875, N862, N103, N264);
nand NAND4 (N876, N875, N402, N328, N831);
not NOT1 (N877, N870);
xor XOR2 (N878, N874, N105);
nand NAND3 (N879, N861, N470, N406);
nand NAND2 (N880, N866, N280);
or OR4 (N881, N872, N773, N854, N458);
not NOT1 (N882, N876);
xor XOR2 (N883, N878, N466);
and AND4 (N884, N867, N433, N95, N567);
buf BUF1 (N885, N880);
buf BUF1 (N886, N877);
xor XOR2 (N887, N884, N518);
nand NAND4 (N888, N882, N535, N549, N508);
and AND3 (N889, N885, N259, N553);
or OR2 (N890, N886, N427);
and AND4 (N891, N889, N98, N527, N537);
xor XOR2 (N892, N890, N74);
nor NOR2 (N893, N892, N389);
and AND3 (N894, N853, N459, N233);
buf BUF1 (N895, N863);
nor NOR4 (N896, N873, N254, N780, N854);
nor NOR3 (N897, N896, N259, N24);
or OR3 (N898, N891, N112, N374);
buf BUF1 (N899, N879);
and AND3 (N900, N893, N674, N430);
and AND3 (N901, N900, N858, N72);
xor XOR2 (N902, N895, N246);
nor NOR2 (N903, N883, N785);
not NOT1 (N904, N881);
nor NOR3 (N905, N888, N302, N220);
nand NAND4 (N906, N905, N235, N829, N854);
nor NOR3 (N907, N887, N491, N709);
buf BUF1 (N908, N898);
nand NAND4 (N909, N904, N798, N578, N806);
xor XOR2 (N910, N901, N489);
nor NOR2 (N911, N899, N459);
nor NOR2 (N912, N894, N623);
nand NAND3 (N913, N912, N537, N645);
nor NOR4 (N914, N910, N692, N276, N350);
nor NOR3 (N915, N913, N544, N210);
nand NAND2 (N916, N911, N314);
or OR3 (N917, N909, N393, N66);
buf BUF1 (N918, N906);
and AND2 (N919, N907, N232);
and AND3 (N920, N919, N224, N138);
buf BUF1 (N921, N897);
nor NOR4 (N922, N915, N637, N477, N437);
xor XOR2 (N923, N908, N234);
xor XOR2 (N924, N918, N298);
nor NOR4 (N925, N917, N845, N327, N733);
nor NOR3 (N926, N923, N490, N255);
buf BUF1 (N927, N902);
nand NAND2 (N928, N927, N236);
nor NOR3 (N929, N916, N789, N823);
nor NOR3 (N930, N914, N381, N768);
nand NAND3 (N931, N922, N749, N33);
buf BUF1 (N932, N926);
xor XOR2 (N933, N928, N454);
nand NAND2 (N934, N931, N566);
not NOT1 (N935, N933);
nor NOR3 (N936, N929, N138, N367);
or OR3 (N937, N935, N461, N126);
xor XOR2 (N938, N924, N472);
not NOT1 (N939, N930);
nor NOR4 (N940, N939, N311, N119, N493);
buf BUF1 (N941, N932);
or OR4 (N942, N941, N124, N861, N668);
xor XOR2 (N943, N940, N322);
and AND2 (N944, N920, N745);
nor NOR2 (N945, N921, N242);
nand NAND3 (N946, N925, N668, N884);
buf BUF1 (N947, N934);
and AND3 (N948, N937, N614, N170);
buf BUF1 (N949, N946);
buf BUF1 (N950, N948);
xor XOR2 (N951, N949, N313);
xor XOR2 (N952, N936, N742);
nand NAND3 (N953, N947, N289, N301);
or OR4 (N954, N953, N827, N822, N397);
nand NAND3 (N955, N938, N767, N449);
nand NAND2 (N956, N943, N877);
not NOT1 (N957, N954);
or OR4 (N958, N951, N755, N904, N306);
xor XOR2 (N959, N945, N850);
nor NOR2 (N960, N903, N88);
buf BUF1 (N961, N957);
buf BUF1 (N962, N944);
nand NAND2 (N963, N950, N675);
nor NOR3 (N964, N959, N657, N893);
buf BUF1 (N965, N955);
xor XOR2 (N966, N965, N257);
or OR4 (N967, N960, N36, N215, N71);
xor XOR2 (N968, N962, N411);
xor XOR2 (N969, N956, N337);
and AND3 (N970, N968, N158, N444);
buf BUF1 (N971, N964);
and AND2 (N972, N942, N43);
xor XOR2 (N973, N952, N298);
xor XOR2 (N974, N973, N108);
not NOT1 (N975, N970);
and AND4 (N976, N958, N347, N347, N800);
nand NAND2 (N977, N976, N905);
or OR3 (N978, N963, N681, N90);
or OR2 (N979, N971, N202);
and AND4 (N980, N961, N349, N336, N358);
xor XOR2 (N981, N972, N305);
xor XOR2 (N982, N974, N382);
buf BUF1 (N983, N981);
nor NOR2 (N984, N983, N554);
and AND4 (N985, N977, N552, N659, N422);
xor XOR2 (N986, N966, N379);
not NOT1 (N987, N978);
buf BUF1 (N988, N969);
nor NOR2 (N989, N967, N815);
nor NOR4 (N990, N975, N514, N859, N558);
nor NOR3 (N991, N982, N935, N762);
or OR2 (N992, N984, N489);
buf BUF1 (N993, N985);
nor NOR4 (N994, N979, N336, N464, N326);
nor NOR2 (N995, N986, N767);
xor XOR2 (N996, N980, N62);
nand NAND2 (N997, N994, N657);
xor XOR2 (N998, N990, N582);
nor NOR3 (N999, N997, N246, N294);
nor NOR2 (N1000, N992, N854);
or OR3 (N1001, N996, N602, N622);
or OR2 (N1002, N987, N775);
xor XOR2 (N1003, N998, N939);
buf BUF1 (N1004, N999);
xor XOR2 (N1005, N991, N425);
nor NOR4 (N1006, N1004, N137, N204, N812);
not NOT1 (N1007, N1005);
buf BUF1 (N1008, N1006);
not NOT1 (N1009, N1007);
or OR3 (N1010, N1009, N722, N941);
or OR2 (N1011, N1010, N333);
not NOT1 (N1012, N1011);
xor XOR2 (N1013, N1008, N207);
buf BUF1 (N1014, N988);
buf BUF1 (N1015, N1003);
and AND2 (N1016, N1002, N28);
nor NOR4 (N1017, N1015, N531, N21, N143);
nor NOR4 (N1018, N993, N496, N195, N37);
nand NAND2 (N1019, N1001, N562);
endmodule