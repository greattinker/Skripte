// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N1514,N1508,N1486,N1493,N1515,N1517,N1506,N1512,N1494,N1518;

or OR3 (N19, N8, N15, N13);
nand NAND3 (N20, N3, N5, N5);
not NOT1 (N21, N12);
buf BUF1 (N22, N14);
buf BUF1 (N23, N20);
not NOT1 (N24, N17);
nor NOR2 (N25, N9, N7);
nand NAND4 (N26, N14, N8, N11, N20);
buf BUF1 (N27, N7);
nor NOR3 (N28, N3, N3, N17);
xor XOR2 (N29, N27, N24);
or OR3 (N30, N29, N23, N24);
xor XOR2 (N31, N11, N2);
nand NAND2 (N32, N8, N30);
not NOT1 (N33, N31);
or OR3 (N34, N33, N22, N9);
or OR2 (N35, N8, N22);
xor XOR2 (N36, N10, N14);
not NOT1 (N37, N16);
nand NAND3 (N38, N37, N11, N5);
xor XOR2 (N39, N34, N4);
nor NOR4 (N40, N19, N33, N12, N22);
or OR3 (N41, N25, N19, N36);
and AND2 (N42, N28, N13);
not NOT1 (N43, N29);
and AND3 (N44, N35, N11, N39);
and AND4 (N45, N31, N41, N13, N31);
xor XOR2 (N46, N17, N18);
or OR2 (N47, N45, N37);
nand NAND3 (N48, N44, N39, N6);
and AND2 (N49, N43, N47);
nand NAND4 (N50, N23, N30, N2, N49);
and AND2 (N51, N26, N34);
not NOT1 (N52, N35);
xor XOR2 (N53, N46, N48);
not NOT1 (N54, N1);
and AND3 (N55, N38, N2, N15);
or OR3 (N56, N52, N43, N12);
and AND4 (N57, N53, N20, N48, N19);
buf BUF1 (N58, N32);
buf BUF1 (N59, N51);
or OR4 (N60, N58, N22, N54, N20);
and AND3 (N61, N40, N10, N17);
not NOT1 (N62, N48);
nor NOR2 (N63, N56, N21);
not NOT1 (N64, N1);
or OR2 (N65, N55, N2);
nor NOR4 (N66, N61, N64, N4, N30);
nand NAND2 (N67, N43, N55);
or OR2 (N68, N50, N21);
xor XOR2 (N69, N63, N2);
xor XOR2 (N70, N59, N29);
buf BUF1 (N71, N57);
buf BUF1 (N72, N70);
nand NAND3 (N73, N72, N53, N45);
buf BUF1 (N74, N60);
or OR3 (N75, N73, N55, N67);
buf BUF1 (N76, N51);
nor NOR4 (N77, N71, N43, N30, N1);
xor XOR2 (N78, N77, N29);
not NOT1 (N79, N78);
or OR4 (N80, N75, N47, N32, N30);
buf BUF1 (N81, N79);
buf BUF1 (N82, N80);
not NOT1 (N83, N69);
nand NAND3 (N84, N42, N65, N9);
and AND4 (N85, N49, N45, N51, N64);
or OR4 (N86, N74, N77, N15, N21);
nor NOR3 (N87, N83, N63, N41);
not NOT1 (N88, N81);
nor NOR4 (N89, N62, N12, N39, N32);
buf BUF1 (N90, N86);
nor NOR3 (N91, N66, N81, N74);
and AND2 (N92, N68, N70);
buf BUF1 (N93, N91);
nor NOR2 (N94, N76, N78);
nor NOR3 (N95, N84, N17, N25);
or OR4 (N96, N94, N5, N27, N75);
not NOT1 (N97, N88);
nor NOR4 (N98, N96, N20, N4, N74);
xor XOR2 (N99, N82, N31);
nand NAND3 (N100, N99, N61, N60);
nor NOR3 (N101, N95, N99, N11);
not NOT1 (N102, N85);
not NOT1 (N103, N92);
nand NAND3 (N104, N97, N95, N68);
not NOT1 (N105, N100);
or OR2 (N106, N98, N61);
not NOT1 (N107, N106);
not NOT1 (N108, N107);
or OR4 (N109, N103, N87, N42, N37);
buf BUF1 (N110, N24);
and AND2 (N111, N108, N55);
or OR3 (N112, N111, N18, N96);
not NOT1 (N113, N101);
nand NAND3 (N114, N104, N2, N54);
nor NOR2 (N115, N114, N21);
nand NAND3 (N116, N109, N55, N37);
and AND4 (N117, N89, N15, N43, N111);
nor NOR2 (N118, N105, N48);
nor NOR3 (N119, N117, N3, N9);
or OR4 (N120, N118, N61, N56, N59);
or OR4 (N121, N120, N50, N5, N91);
nor NOR2 (N122, N93, N74);
or OR3 (N123, N116, N29, N61);
buf BUF1 (N124, N110);
nand NAND4 (N125, N113, N80, N47, N13);
or OR4 (N126, N90, N90, N43, N51);
nand NAND4 (N127, N126, N93, N126, N37);
xor XOR2 (N128, N127, N72);
not NOT1 (N129, N121);
nand NAND3 (N130, N125, N28, N60);
nor NOR4 (N131, N119, N28, N75, N82);
buf BUF1 (N132, N124);
nor NOR3 (N133, N129, N13, N102);
buf BUF1 (N134, N92);
buf BUF1 (N135, N131);
buf BUF1 (N136, N123);
buf BUF1 (N137, N112);
nor NOR3 (N138, N115, N13, N129);
or OR3 (N139, N138, N73, N58);
or OR2 (N140, N136, N133);
nand NAND4 (N141, N93, N77, N82, N33);
or OR3 (N142, N130, N36, N108);
not NOT1 (N143, N139);
and AND4 (N144, N140, N82, N115, N122);
nor NOR2 (N145, N110, N104);
nor NOR4 (N146, N144, N37, N136, N103);
not NOT1 (N147, N141);
and AND2 (N148, N142, N85);
and AND2 (N149, N134, N64);
or OR3 (N150, N135, N10, N22);
and AND3 (N151, N145, N10, N41);
not NOT1 (N152, N150);
xor XOR2 (N153, N149, N84);
not NOT1 (N154, N151);
nand NAND3 (N155, N143, N38, N85);
xor XOR2 (N156, N155, N21);
buf BUF1 (N157, N132);
buf BUF1 (N158, N148);
not NOT1 (N159, N153);
buf BUF1 (N160, N158);
xor XOR2 (N161, N152, N53);
nand NAND3 (N162, N154, N129, N21);
nand NAND3 (N163, N147, N49, N2);
xor XOR2 (N164, N159, N70);
xor XOR2 (N165, N164, N153);
or OR2 (N166, N162, N79);
nand NAND3 (N167, N161, N26, N102);
nand NAND3 (N168, N157, N22, N57);
and AND2 (N169, N168, N21);
xor XOR2 (N170, N146, N165);
nand NAND2 (N171, N64, N68);
not NOT1 (N172, N156);
or OR3 (N173, N167, N63, N4);
nand NAND3 (N174, N171, N56, N26);
nor NOR3 (N175, N160, N10, N42);
xor XOR2 (N176, N169, N10);
buf BUF1 (N177, N128);
not NOT1 (N178, N173);
or OR2 (N179, N172, N70);
and AND4 (N180, N178, N53, N123, N25);
or OR4 (N181, N176, N99, N159, N1);
nor NOR3 (N182, N180, N181, N96);
not NOT1 (N183, N103);
buf BUF1 (N184, N177);
or OR2 (N185, N174, N180);
and AND4 (N186, N185, N181, N41, N2);
buf BUF1 (N187, N184);
nor NOR4 (N188, N186, N123, N42, N87);
nor NOR3 (N189, N183, N165, N112);
nor NOR2 (N190, N175, N182);
xor XOR2 (N191, N19, N94);
xor XOR2 (N192, N189, N106);
buf BUF1 (N193, N192);
xor XOR2 (N194, N193, N132);
buf BUF1 (N195, N170);
nor NOR3 (N196, N191, N162, N151);
buf BUF1 (N197, N166);
nand NAND2 (N198, N196, N51);
nand NAND4 (N199, N179, N193, N5, N109);
or OR2 (N200, N199, N100);
and AND4 (N201, N198, N33, N161, N16);
or OR2 (N202, N137, N127);
or OR4 (N203, N197, N26, N103, N109);
or OR2 (N204, N203, N123);
nor NOR3 (N205, N188, N80, N189);
nor NOR3 (N206, N195, N120, N100);
or OR3 (N207, N190, N56, N125);
nand NAND4 (N208, N205, N26, N147, N150);
and AND3 (N209, N207, N59, N186);
and AND4 (N210, N163, N72, N89, N3);
nand NAND3 (N211, N187, N42, N151);
buf BUF1 (N212, N201);
nor NOR3 (N213, N210, N174, N124);
and AND3 (N214, N204, N68, N93);
xor XOR2 (N215, N209, N87);
nor NOR2 (N216, N211, N127);
nor NOR2 (N217, N213, N140);
buf BUF1 (N218, N202);
nor NOR3 (N219, N215, N189, N215);
nand NAND4 (N220, N216, N183, N139, N42);
nand NAND2 (N221, N214, N190);
not NOT1 (N222, N194);
nand NAND3 (N223, N220, N95, N141);
or OR3 (N224, N223, N152, N20);
nor NOR2 (N225, N208, N25);
not NOT1 (N226, N218);
nand NAND4 (N227, N200, N194, N209, N220);
buf BUF1 (N228, N227);
xor XOR2 (N229, N219, N108);
nor NOR2 (N230, N226, N47);
and AND4 (N231, N228, N83, N100, N50);
not NOT1 (N232, N212);
not NOT1 (N233, N224);
or OR2 (N234, N231, N69);
or OR2 (N235, N232, N130);
nor NOR4 (N236, N234, N163, N70, N190);
nand NAND2 (N237, N217, N194);
buf BUF1 (N238, N206);
xor XOR2 (N239, N235, N29);
nor NOR4 (N240, N225, N191, N109, N70);
nand NAND3 (N241, N222, N39, N29);
xor XOR2 (N242, N240, N142);
buf BUF1 (N243, N229);
nor NOR3 (N244, N239, N123, N213);
xor XOR2 (N245, N230, N128);
and AND4 (N246, N241, N235, N232, N32);
not NOT1 (N247, N244);
nand NAND2 (N248, N237, N88);
and AND2 (N249, N247, N60);
nor NOR3 (N250, N248, N191, N63);
not NOT1 (N251, N242);
nor NOR3 (N252, N251, N2, N36);
xor XOR2 (N253, N238, N232);
and AND2 (N254, N250, N18);
and AND4 (N255, N252, N37, N150, N88);
buf BUF1 (N256, N253);
or OR4 (N257, N254, N120, N63, N95);
buf BUF1 (N258, N257);
and AND3 (N259, N258, N158, N228);
buf BUF1 (N260, N236);
not NOT1 (N261, N243);
xor XOR2 (N262, N245, N62);
or OR3 (N263, N262, N154, N123);
not NOT1 (N264, N256);
nand NAND3 (N265, N261, N45, N109);
or OR2 (N266, N221, N92);
xor XOR2 (N267, N264, N29);
and AND4 (N268, N267, N115, N114, N175);
and AND2 (N269, N263, N183);
nand NAND4 (N270, N260, N152, N233, N232);
or OR3 (N271, N192, N222, N26);
or OR3 (N272, N271, N237, N229);
not NOT1 (N273, N268);
xor XOR2 (N274, N265, N132);
nand NAND2 (N275, N272, N159);
nand NAND3 (N276, N266, N193, N29);
nand NAND2 (N277, N273, N92);
nor NOR3 (N278, N270, N263, N28);
not NOT1 (N279, N275);
not NOT1 (N280, N259);
and AND4 (N281, N274, N42, N126, N153);
and AND4 (N282, N279, N180, N236, N268);
or OR4 (N283, N280, N230, N166, N6);
nand NAND2 (N284, N278, N9);
xor XOR2 (N285, N246, N187);
or OR3 (N286, N269, N249, N105);
nor NOR4 (N287, N132, N21, N171, N84);
xor XOR2 (N288, N287, N237);
not NOT1 (N289, N284);
nand NAND4 (N290, N281, N78, N231, N238);
buf BUF1 (N291, N283);
not NOT1 (N292, N288);
and AND4 (N293, N291, N64, N169, N290);
nor NOR3 (N294, N189, N6, N9);
or OR4 (N295, N289, N2, N187, N110);
buf BUF1 (N296, N293);
or OR4 (N297, N286, N20, N98, N270);
or OR4 (N298, N276, N52, N264, N87);
or OR2 (N299, N277, N166);
nand NAND2 (N300, N285, N64);
and AND4 (N301, N299, N96, N228, N132);
or OR4 (N302, N297, N32, N272, N289);
nor NOR4 (N303, N298, N54, N262, N15);
and AND4 (N304, N302, N282, N201, N129);
nor NOR4 (N305, N41, N184, N186, N141);
buf BUF1 (N306, N296);
and AND4 (N307, N300, N244, N233, N210);
nand NAND3 (N308, N294, N182, N89);
or OR3 (N309, N255, N1, N66);
not NOT1 (N310, N305);
or OR2 (N311, N292, N26);
nor NOR3 (N312, N303, N228, N273);
buf BUF1 (N313, N310);
nand NAND2 (N314, N306, N4);
nor NOR3 (N315, N312, N314, N85);
not NOT1 (N316, N40);
nor NOR3 (N317, N304, N313, N289);
buf BUF1 (N318, N281);
not NOT1 (N319, N309);
or OR2 (N320, N307, N278);
not NOT1 (N321, N295);
xor XOR2 (N322, N316, N161);
nor NOR3 (N323, N318, N49, N160);
not NOT1 (N324, N321);
xor XOR2 (N325, N320, N91);
nor NOR3 (N326, N325, N273, N144);
nor NOR3 (N327, N319, N75, N231);
nor NOR3 (N328, N326, N89, N174);
xor XOR2 (N329, N315, N100);
and AND2 (N330, N322, N28);
buf BUF1 (N331, N317);
or OR3 (N332, N327, N212, N61);
not NOT1 (N333, N324);
xor XOR2 (N334, N333, N207);
nor NOR4 (N335, N330, N157, N177, N229);
or OR2 (N336, N332, N161);
nand NAND3 (N337, N336, N254, N179);
and AND3 (N338, N301, N8, N246);
nand NAND4 (N339, N311, N144, N299, N246);
or OR3 (N340, N328, N336, N196);
buf BUF1 (N341, N339);
not NOT1 (N342, N331);
buf BUF1 (N343, N342);
or OR3 (N344, N341, N89, N247);
buf BUF1 (N345, N334);
xor XOR2 (N346, N323, N123);
buf BUF1 (N347, N345);
nand NAND4 (N348, N335, N60, N90, N215);
nand NAND4 (N349, N337, N179, N301, N34);
or OR4 (N350, N346, N220, N37, N194);
buf BUF1 (N351, N350);
nor NOR4 (N352, N329, N193, N56, N100);
nand NAND3 (N353, N351, N213, N352);
or OR3 (N354, N296, N209, N70);
nor NOR4 (N355, N344, N99, N135, N145);
or OR2 (N356, N348, N54);
not NOT1 (N357, N338);
or OR4 (N358, N349, N133, N287, N110);
and AND4 (N359, N354, N47, N160, N16);
not NOT1 (N360, N355);
not NOT1 (N361, N343);
nand NAND4 (N362, N347, N17, N145, N252);
or OR3 (N363, N356, N361, N6);
and AND3 (N364, N186, N341, N47);
or OR3 (N365, N362, N181, N65);
and AND2 (N366, N357, N237);
and AND3 (N367, N308, N321, N320);
and AND2 (N368, N364, N335);
and AND4 (N369, N359, N227, N210, N97);
nor NOR2 (N370, N369, N357);
buf BUF1 (N371, N366);
or OR2 (N372, N363, N77);
buf BUF1 (N373, N371);
buf BUF1 (N374, N368);
and AND3 (N375, N340, N38, N195);
or OR4 (N376, N360, N190, N166, N129);
nor NOR3 (N377, N373, N232, N333);
or OR3 (N378, N367, N76, N190);
xor XOR2 (N379, N374, N127);
nand NAND2 (N380, N370, N260);
or OR2 (N381, N380, N146);
xor XOR2 (N382, N358, N324);
nor NOR2 (N383, N382, N268);
xor XOR2 (N384, N383, N154);
nand NAND3 (N385, N378, N306, N141);
not NOT1 (N386, N372);
nand NAND3 (N387, N385, N242, N370);
xor XOR2 (N388, N375, N314);
or OR4 (N389, N386, N299, N245, N147);
xor XOR2 (N390, N353, N126);
buf BUF1 (N391, N389);
nand NAND3 (N392, N379, N181, N182);
xor XOR2 (N393, N390, N45);
buf BUF1 (N394, N376);
or OR2 (N395, N387, N2);
nand NAND3 (N396, N394, N170, N191);
xor XOR2 (N397, N365, N326);
xor XOR2 (N398, N392, N148);
not NOT1 (N399, N393);
not NOT1 (N400, N391);
or OR3 (N401, N384, N356, N44);
nor NOR2 (N402, N388, N165);
nor NOR3 (N403, N381, N159, N188);
nor NOR4 (N404, N395, N323, N265, N283);
not NOT1 (N405, N400);
xor XOR2 (N406, N405, N351);
xor XOR2 (N407, N404, N21);
not NOT1 (N408, N398);
or OR2 (N409, N401, N151);
nand NAND3 (N410, N407, N136, N334);
and AND2 (N411, N399, N33);
not NOT1 (N412, N402);
xor XOR2 (N413, N410, N227);
buf BUF1 (N414, N408);
nor NOR3 (N415, N397, N315, N192);
nor NOR2 (N416, N414, N192);
nor NOR3 (N417, N412, N152, N332);
and AND3 (N418, N377, N305, N14);
or OR4 (N419, N416, N274, N33, N114);
not NOT1 (N420, N406);
buf BUF1 (N421, N418);
not NOT1 (N422, N421);
buf BUF1 (N423, N403);
nand NAND4 (N424, N411, N340, N383, N76);
nand NAND3 (N425, N396, N90, N118);
and AND3 (N426, N409, N92, N99);
not NOT1 (N427, N423);
or OR4 (N428, N413, N236, N34, N160);
nand NAND4 (N429, N422, N362, N302, N343);
nand NAND4 (N430, N429, N100, N393, N125);
or OR2 (N431, N419, N238);
and AND2 (N432, N417, N175);
nor NOR4 (N433, N415, N426, N92, N14);
xor XOR2 (N434, N284, N339);
not NOT1 (N435, N432);
buf BUF1 (N436, N425);
buf BUF1 (N437, N433);
or OR2 (N438, N435, N31);
or OR2 (N439, N430, N210);
nor NOR3 (N440, N438, N168, N122);
xor XOR2 (N441, N424, N71);
not NOT1 (N442, N434);
buf BUF1 (N443, N436);
or OR2 (N444, N439, N219);
or OR4 (N445, N442, N2, N432, N320);
not NOT1 (N446, N420);
and AND3 (N447, N443, N31, N60);
not NOT1 (N448, N428);
xor XOR2 (N449, N431, N215);
and AND3 (N450, N437, N134, N117);
and AND2 (N451, N449, N352);
nand NAND4 (N452, N451, N94, N233, N194);
buf BUF1 (N453, N445);
nor NOR2 (N454, N447, N424);
buf BUF1 (N455, N440);
or OR2 (N456, N450, N235);
and AND3 (N457, N454, N318, N353);
and AND4 (N458, N457, N350, N166, N429);
and AND4 (N459, N455, N368, N321, N204);
nand NAND4 (N460, N453, N72, N412, N52);
nor NOR3 (N461, N459, N240, N316);
buf BUF1 (N462, N456);
not NOT1 (N463, N448);
and AND4 (N464, N460, N288, N434, N117);
or OR2 (N465, N464, N326);
and AND3 (N466, N452, N287, N371);
nor NOR3 (N467, N446, N116, N198);
nand NAND4 (N468, N444, N100, N151, N294);
buf BUF1 (N469, N462);
or OR2 (N470, N466, N377);
xor XOR2 (N471, N468, N80);
nand NAND4 (N472, N427, N436, N378, N334);
not NOT1 (N473, N463);
or OR4 (N474, N458, N388, N425, N14);
nor NOR4 (N475, N474, N173, N283, N331);
not NOT1 (N476, N467);
and AND2 (N477, N465, N302);
or OR3 (N478, N477, N404, N224);
buf BUF1 (N479, N478);
xor XOR2 (N480, N470, N129);
nand NAND2 (N481, N479, N344);
not NOT1 (N482, N469);
nand NAND3 (N483, N461, N189, N439);
xor XOR2 (N484, N441, N332);
nand NAND3 (N485, N475, N281, N182);
nor NOR4 (N486, N473, N195, N428, N73);
nor NOR4 (N487, N481, N114, N430, N442);
or OR2 (N488, N482, N136);
nand NAND2 (N489, N488, N328);
and AND3 (N490, N486, N247, N319);
or OR4 (N491, N490, N372, N20, N193);
xor XOR2 (N492, N480, N144);
and AND2 (N493, N472, N26);
and AND4 (N494, N484, N433, N183, N310);
xor XOR2 (N495, N487, N444);
or OR2 (N496, N489, N440);
xor XOR2 (N497, N492, N69);
nand NAND4 (N498, N496, N256, N460, N90);
nor NOR3 (N499, N483, N69, N457);
buf BUF1 (N500, N476);
nor NOR4 (N501, N493, N20, N309, N87);
and AND2 (N502, N497, N113);
nor NOR3 (N503, N485, N328, N407);
not NOT1 (N504, N471);
not NOT1 (N505, N495);
xor XOR2 (N506, N499, N326);
xor XOR2 (N507, N494, N333);
nor NOR2 (N508, N500, N32);
not NOT1 (N509, N491);
xor XOR2 (N510, N498, N10);
and AND2 (N511, N503, N485);
nor NOR3 (N512, N501, N473, N123);
or OR4 (N513, N502, N362, N444, N109);
xor XOR2 (N514, N512, N142);
buf BUF1 (N515, N506);
nor NOR4 (N516, N505, N17, N324, N493);
nand NAND2 (N517, N515, N508);
or OR2 (N518, N244, N137);
xor XOR2 (N519, N514, N332);
nand NAND3 (N520, N513, N387, N219);
or OR4 (N521, N511, N152, N159, N79);
or OR3 (N522, N517, N94, N446);
not NOT1 (N523, N522);
buf BUF1 (N524, N510);
and AND3 (N525, N518, N233, N369);
not NOT1 (N526, N509);
or OR4 (N527, N516, N195, N33, N428);
or OR3 (N528, N525, N252, N217);
nand NAND2 (N529, N507, N80);
buf BUF1 (N530, N527);
not NOT1 (N531, N523);
xor XOR2 (N532, N531, N303);
or OR2 (N533, N532, N42);
buf BUF1 (N534, N504);
buf BUF1 (N535, N534);
and AND4 (N536, N520, N399, N477, N143);
not NOT1 (N537, N529);
xor XOR2 (N538, N528, N132);
not NOT1 (N539, N521);
not NOT1 (N540, N535);
xor XOR2 (N541, N533, N25);
nor NOR3 (N542, N539, N222, N212);
nor NOR3 (N543, N542, N130, N90);
nand NAND4 (N544, N519, N154, N174, N72);
nor NOR2 (N545, N544, N72);
nor NOR4 (N546, N541, N519, N249, N35);
xor XOR2 (N547, N537, N291);
not NOT1 (N548, N524);
and AND2 (N549, N545, N358);
buf BUF1 (N550, N547);
nand NAND3 (N551, N549, N263, N289);
not NOT1 (N552, N543);
and AND2 (N553, N536, N215);
nor NOR3 (N554, N550, N413, N452);
nor NOR2 (N555, N546, N218);
nor NOR3 (N556, N553, N138, N94);
or OR3 (N557, N552, N290, N527);
or OR2 (N558, N548, N184);
nor NOR4 (N559, N557, N348, N289, N105);
and AND4 (N560, N538, N194, N238, N433);
not NOT1 (N561, N559);
nor NOR2 (N562, N560, N148);
nor NOR3 (N563, N558, N331, N518);
or OR2 (N564, N551, N253);
nor NOR4 (N565, N561, N102, N290, N199);
nand NAND3 (N566, N563, N494, N296);
and AND3 (N567, N566, N62, N128);
not NOT1 (N568, N565);
not NOT1 (N569, N555);
nor NOR3 (N570, N569, N351, N37);
nand NAND3 (N571, N562, N136, N443);
nor NOR3 (N572, N564, N194, N210);
nand NAND3 (N573, N530, N518, N477);
not NOT1 (N574, N567);
nor NOR2 (N575, N573, N542);
nor NOR3 (N576, N574, N508, N141);
not NOT1 (N577, N540);
nor NOR3 (N578, N576, N474, N471);
xor XOR2 (N579, N578, N129);
not NOT1 (N580, N577);
or OR2 (N581, N579, N480);
not NOT1 (N582, N526);
nand NAND2 (N583, N581, N298);
not NOT1 (N584, N583);
nor NOR2 (N585, N572, N376);
or OR4 (N586, N571, N466, N178, N1);
nor NOR4 (N587, N580, N572, N219, N102);
and AND4 (N588, N568, N320, N235, N512);
and AND2 (N589, N586, N463);
or OR2 (N590, N588, N296);
nor NOR4 (N591, N584, N75, N392, N339);
nand NAND4 (N592, N585, N446, N555, N10);
xor XOR2 (N593, N582, N263);
nand NAND4 (N594, N593, N578, N572, N18);
buf BUF1 (N595, N591);
xor XOR2 (N596, N556, N276);
and AND2 (N597, N570, N235);
nor NOR2 (N598, N554, N147);
not NOT1 (N599, N595);
and AND4 (N600, N587, N186, N65, N53);
or OR3 (N601, N592, N388, N396);
xor XOR2 (N602, N601, N392);
xor XOR2 (N603, N590, N12);
not NOT1 (N604, N589);
nand NAND3 (N605, N597, N300, N199);
nand NAND3 (N606, N594, N519, N514);
nand NAND4 (N607, N600, N259, N520, N337);
nand NAND4 (N608, N575, N301, N321, N397);
and AND4 (N609, N598, N292, N578, N44);
nand NAND3 (N610, N606, N120, N137);
not NOT1 (N611, N604);
buf BUF1 (N612, N608);
nor NOR4 (N613, N603, N404, N451, N20);
xor XOR2 (N614, N610, N250);
or OR3 (N615, N612, N259, N68);
buf BUF1 (N616, N596);
nor NOR2 (N617, N607, N231);
or OR2 (N618, N602, N323);
xor XOR2 (N619, N618, N75);
xor XOR2 (N620, N615, N14);
and AND3 (N621, N619, N373, N308);
and AND2 (N622, N599, N538);
not NOT1 (N623, N614);
buf BUF1 (N624, N617);
or OR4 (N625, N613, N622, N398, N312);
nor NOR3 (N626, N169, N179, N227);
and AND2 (N627, N626, N512);
xor XOR2 (N628, N605, N20);
and AND2 (N629, N616, N266);
buf BUF1 (N630, N628);
buf BUF1 (N631, N621);
not NOT1 (N632, N627);
nor NOR2 (N633, N624, N362);
not NOT1 (N634, N620);
and AND4 (N635, N634, N181, N156, N81);
buf BUF1 (N636, N625);
buf BUF1 (N637, N609);
buf BUF1 (N638, N633);
xor XOR2 (N639, N638, N294);
xor XOR2 (N640, N632, N424);
buf BUF1 (N641, N630);
not NOT1 (N642, N636);
nand NAND4 (N643, N640, N472, N195, N48);
buf BUF1 (N644, N611);
buf BUF1 (N645, N641);
nand NAND2 (N646, N623, N32);
or OR3 (N647, N643, N357, N288);
nor NOR4 (N648, N629, N97, N351, N169);
nor NOR3 (N649, N631, N489, N59);
or OR3 (N650, N647, N40, N559);
nor NOR3 (N651, N642, N297, N373);
not NOT1 (N652, N637);
buf BUF1 (N653, N639);
nand NAND3 (N654, N649, N289, N70);
xor XOR2 (N655, N646, N32);
or OR4 (N656, N650, N477, N496, N304);
nand NAND4 (N657, N651, N14, N528, N270);
nor NOR4 (N658, N645, N30, N155, N454);
nand NAND2 (N659, N654, N167);
and AND3 (N660, N653, N437, N575);
xor XOR2 (N661, N656, N628);
nand NAND2 (N662, N658, N573);
not NOT1 (N663, N661);
nor NOR3 (N664, N648, N164, N498);
nor NOR2 (N665, N655, N481);
nand NAND3 (N666, N663, N435, N486);
or OR3 (N667, N657, N160, N639);
buf BUF1 (N668, N665);
and AND4 (N669, N666, N35, N408, N122);
xor XOR2 (N670, N635, N614);
or OR2 (N671, N664, N262);
buf BUF1 (N672, N670);
nand NAND2 (N673, N644, N331);
and AND4 (N674, N660, N575, N88, N105);
or OR3 (N675, N671, N477, N144);
and AND3 (N676, N668, N456, N616);
nor NOR3 (N677, N669, N121, N122);
or OR3 (N678, N675, N502, N339);
buf BUF1 (N679, N659);
not NOT1 (N680, N679);
xor XOR2 (N681, N662, N643);
not NOT1 (N682, N667);
and AND4 (N683, N652, N31, N84, N67);
or OR4 (N684, N680, N509, N261, N378);
and AND4 (N685, N672, N617, N263, N79);
and AND2 (N686, N677, N340);
not NOT1 (N687, N673);
nor NOR2 (N688, N674, N132);
nand NAND4 (N689, N682, N572, N327, N134);
nand NAND4 (N690, N685, N396, N497, N429);
and AND3 (N691, N689, N189, N16);
and AND4 (N692, N686, N149, N499, N573);
nor NOR4 (N693, N681, N329, N368, N204);
or OR4 (N694, N691, N448, N136, N636);
not NOT1 (N695, N688);
not NOT1 (N696, N676);
and AND2 (N697, N683, N159);
or OR4 (N698, N693, N476, N497, N604);
buf BUF1 (N699, N692);
or OR4 (N700, N678, N10, N532, N560);
xor XOR2 (N701, N698, N323);
and AND2 (N702, N687, N434);
not NOT1 (N703, N699);
and AND3 (N704, N684, N428, N202);
buf BUF1 (N705, N697);
buf BUF1 (N706, N694);
not NOT1 (N707, N690);
buf BUF1 (N708, N703);
nor NOR2 (N709, N707, N385);
nand NAND3 (N710, N696, N104, N203);
nor NOR4 (N711, N701, N261, N148, N231);
and AND3 (N712, N704, N288, N518);
or OR2 (N713, N705, N493);
buf BUF1 (N714, N712);
nand NAND3 (N715, N710, N686, N436);
or OR2 (N716, N714, N324);
or OR3 (N717, N708, N704, N119);
xor XOR2 (N718, N716, N674);
not NOT1 (N719, N718);
buf BUF1 (N720, N702);
nand NAND3 (N721, N711, N169, N85);
nor NOR2 (N722, N706, N182);
or OR2 (N723, N713, N427);
and AND2 (N724, N722, N360);
nand NAND4 (N725, N719, N563, N690, N679);
buf BUF1 (N726, N724);
and AND4 (N727, N723, N409, N374, N476);
buf BUF1 (N728, N720);
nand NAND4 (N729, N727, N207, N379, N273);
nor NOR4 (N730, N726, N221, N371, N452);
not NOT1 (N731, N728);
nor NOR4 (N732, N725, N201, N654, N565);
nand NAND4 (N733, N715, N284, N634, N12);
or OR3 (N734, N729, N74, N568);
nand NAND3 (N735, N700, N458, N637);
nor NOR3 (N736, N709, N584, N586);
buf BUF1 (N737, N735);
and AND2 (N738, N717, N5);
buf BUF1 (N739, N737);
buf BUF1 (N740, N730);
buf BUF1 (N741, N736);
or OR3 (N742, N741, N527, N260);
nand NAND2 (N743, N695, N294);
or OR2 (N744, N742, N636);
and AND3 (N745, N731, N376, N34);
buf BUF1 (N746, N743);
buf BUF1 (N747, N740);
and AND4 (N748, N747, N605, N217, N508);
xor XOR2 (N749, N734, N250);
nand NAND4 (N750, N733, N579, N452, N364);
nor NOR4 (N751, N750, N536, N209, N634);
nor NOR3 (N752, N721, N629, N517);
nor NOR3 (N753, N738, N175, N156);
and AND3 (N754, N751, N488, N101);
and AND3 (N755, N744, N719, N463);
buf BUF1 (N756, N754);
or OR2 (N757, N746, N404);
xor XOR2 (N758, N757, N150);
xor XOR2 (N759, N748, N478);
buf BUF1 (N760, N758);
and AND3 (N761, N749, N289, N90);
xor XOR2 (N762, N745, N591);
nor NOR2 (N763, N753, N612);
xor XOR2 (N764, N756, N503);
buf BUF1 (N765, N764);
or OR4 (N766, N765, N522, N46, N554);
or OR4 (N767, N762, N341, N299, N720);
and AND3 (N768, N752, N382, N135);
and AND2 (N769, N761, N326);
or OR2 (N770, N766, N109);
buf BUF1 (N771, N763);
xor XOR2 (N772, N732, N75);
xor XOR2 (N773, N760, N440);
and AND3 (N774, N759, N510, N426);
nand NAND3 (N775, N772, N635, N610);
not NOT1 (N776, N774);
and AND3 (N777, N755, N26, N421);
and AND3 (N778, N776, N381, N64);
xor XOR2 (N779, N777, N465);
and AND4 (N780, N768, N341, N674, N331);
not NOT1 (N781, N779);
xor XOR2 (N782, N773, N749);
and AND2 (N783, N778, N261);
not NOT1 (N784, N770);
nor NOR2 (N785, N767, N772);
nand NAND2 (N786, N784, N488);
not NOT1 (N787, N785);
xor XOR2 (N788, N786, N711);
xor XOR2 (N789, N782, N475);
and AND2 (N790, N775, N391);
not NOT1 (N791, N783);
not NOT1 (N792, N780);
not NOT1 (N793, N769);
and AND3 (N794, N739, N36, N786);
nand NAND4 (N795, N771, N15, N388, N370);
or OR3 (N796, N791, N45, N355);
xor XOR2 (N797, N796, N338);
or OR2 (N798, N787, N202);
or OR3 (N799, N781, N786, N586);
buf BUF1 (N800, N793);
and AND4 (N801, N799, N736, N495, N78);
not NOT1 (N802, N797);
nand NAND4 (N803, N790, N588, N265, N474);
nand NAND3 (N804, N798, N496, N49);
not NOT1 (N805, N792);
nor NOR4 (N806, N789, N586, N621, N598);
and AND2 (N807, N788, N697);
xor XOR2 (N808, N802, N162);
xor XOR2 (N809, N805, N445);
or OR2 (N810, N804, N636);
nand NAND3 (N811, N810, N720, N727);
and AND3 (N812, N794, N203, N766);
not NOT1 (N813, N808);
buf BUF1 (N814, N811);
nand NAND4 (N815, N801, N707, N27, N164);
or OR2 (N816, N806, N135);
buf BUF1 (N817, N809);
xor XOR2 (N818, N795, N50);
and AND4 (N819, N818, N466, N463, N479);
or OR3 (N820, N817, N757, N217);
nand NAND4 (N821, N814, N278, N506, N606);
not NOT1 (N822, N813);
not NOT1 (N823, N800);
and AND3 (N824, N819, N635, N635);
buf BUF1 (N825, N807);
and AND3 (N826, N820, N139, N793);
or OR3 (N827, N815, N399, N222);
nand NAND4 (N828, N826, N151, N139, N121);
nand NAND3 (N829, N825, N705, N364);
nor NOR2 (N830, N822, N534);
nand NAND4 (N831, N803, N246, N35, N110);
buf BUF1 (N832, N827);
xor XOR2 (N833, N812, N144);
not NOT1 (N834, N824);
and AND3 (N835, N828, N443, N168);
buf BUF1 (N836, N816);
and AND2 (N837, N832, N298);
nand NAND2 (N838, N831, N551);
or OR2 (N839, N834, N8);
not NOT1 (N840, N837);
or OR4 (N841, N838, N424, N806, N558);
buf BUF1 (N842, N821);
or OR2 (N843, N842, N220);
and AND2 (N844, N843, N566);
buf BUF1 (N845, N835);
nor NOR4 (N846, N840, N410, N316, N340);
xor XOR2 (N847, N841, N658);
buf BUF1 (N848, N845);
nor NOR3 (N849, N823, N589, N677);
xor XOR2 (N850, N848, N397);
nand NAND4 (N851, N850, N23, N14, N183);
nor NOR2 (N852, N851, N849);
or OR2 (N853, N367, N344);
and AND3 (N854, N833, N624, N397);
nand NAND2 (N855, N830, N293);
nand NAND2 (N856, N836, N782);
xor XOR2 (N857, N846, N90);
xor XOR2 (N858, N844, N231);
not NOT1 (N859, N847);
xor XOR2 (N860, N859, N782);
nor NOR3 (N861, N854, N735, N615);
nand NAND4 (N862, N853, N452, N488, N535);
nor NOR3 (N863, N829, N172, N104);
nor NOR2 (N864, N861, N273);
xor XOR2 (N865, N855, N259);
nor NOR4 (N866, N856, N499, N360, N185);
not NOT1 (N867, N862);
and AND4 (N868, N852, N235, N202, N338);
nor NOR2 (N869, N864, N531);
buf BUF1 (N870, N866);
buf BUF1 (N871, N858);
and AND4 (N872, N867, N801, N834, N212);
and AND2 (N873, N872, N529);
nor NOR2 (N874, N863, N171);
buf BUF1 (N875, N869);
not NOT1 (N876, N875);
nor NOR2 (N877, N868, N561);
not NOT1 (N878, N871);
buf BUF1 (N879, N839);
or OR3 (N880, N874, N646, N118);
xor XOR2 (N881, N865, N163);
buf BUF1 (N882, N857);
nand NAND2 (N883, N870, N430);
xor XOR2 (N884, N880, N795);
buf BUF1 (N885, N881);
not NOT1 (N886, N885);
nor NOR3 (N887, N882, N742, N264);
not NOT1 (N888, N878);
xor XOR2 (N889, N860, N493);
not NOT1 (N890, N889);
and AND2 (N891, N890, N653);
buf BUF1 (N892, N879);
not NOT1 (N893, N876);
nand NAND2 (N894, N886, N126);
nor NOR3 (N895, N887, N365, N774);
not NOT1 (N896, N893);
xor XOR2 (N897, N884, N510);
buf BUF1 (N898, N888);
and AND3 (N899, N894, N838, N117);
and AND3 (N900, N892, N254, N617);
or OR2 (N901, N891, N245);
or OR4 (N902, N897, N372, N154, N360);
and AND2 (N903, N899, N162);
or OR2 (N904, N901, N1);
nor NOR2 (N905, N902, N557);
xor XOR2 (N906, N905, N527);
xor XOR2 (N907, N896, N671);
not NOT1 (N908, N904);
nor NOR4 (N909, N883, N807, N903, N723);
not NOT1 (N910, N147);
nand NAND4 (N911, N895, N205, N106, N601);
xor XOR2 (N912, N908, N504);
and AND4 (N913, N910, N25, N309, N272);
or OR2 (N914, N877, N875);
nand NAND3 (N915, N900, N854, N386);
or OR2 (N916, N911, N403);
nor NOR4 (N917, N913, N706, N281, N540);
xor XOR2 (N918, N906, N713);
and AND3 (N919, N912, N524, N136);
nand NAND4 (N920, N915, N629, N661, N60);
and AND4 (N921, N907, N199, N569, N879);
and AND4 (N922, N898, N470, N364, N452);
buf BUF1 (N923, N922);
buf BUF1 (N924, N919);
buf BUF1 (N925, N909);
or OR2 (N926, N920, N869);
nand NAND2 (N927, N923, N881);
nand NAND4 (N928, N873, N408, N604, N412);
buf BUF1 (N929, N924);
or OR4 (N930, N916, N886, N332, N912);
nor NOR3 (N931, N929, N22, N733);
and AND2 (N932, N931, N639);
xor XOR2 (N933, N914, N638);
and AND2 (N934, N925, N244);
nor NOR3 (N935, N933, N71, N394);
nor NOR4 (N936, N918, N344, N155, N472);
not NOT1 (N937, N921);
and AND3 (N938, N917, N315, N329);
or OR3 (N939, N934, N305, N48);
xor XOR2 (N940, N926, N587);
or OR2 (N941, N939, N844);
not NOT1 (N942, N927);
and AND4 (N943, N932, N637, N426, N160);
not NOT1 (N944, N930);
or OR4 (N945, N943, N211, N203, N34);
and AND3 (N946, N941, N588, N939);
nand NAND3 (N947, N938, N280, N332);
and AND3 (N948, N940, N517, N476);
nand NAND3 (N949, N936, N635, N541);
not NOT1 (N950, N945);
nor NOR3 (N951, N937, N336, N523);
nand NAND3 (N952, N935, N245, N735);
buf BUF1 (N953, N950);
nor NOR3 (N954, N952, N852, N877);
or OR3 (N955, N949, N614, N839);
xor XOR2 (N956, N954, N11);
nand NAND4 (N957, N946, N571, N30, N58);
nor NOR2 (N958, N955, N645);
nand NAND3 (N959, N947, N920, N578);
xor XOR2 (N960, N928, N444);
buf BUF1 (N961, N944);
buf BUF1 (N962, N961);
or OR2 (N963, N962, N348);
nor NOR3 (N964, N957, N796, N919);
buf BUF1 (N965, N942);
not NOT1 (N966, N958);
nand NAND2 (N967, N965, N925);
nand NAND3 (N968, N951, N27, N554);
or OR4 (N969, N960, N869, N266, N355);
and AND4 (N970, N956, N943, N228, N95);
nor NOR4 (N971, N967, N62, N505, N93);
not NOT1 (N972, N969);
nand NAND2 (N973, N959, N670);
buf BUF1 (N974, N972);
or OR2 (N975, N948, N586);
nand NAND2 (N976, N963, N873);
nand NAND4 (N977, N966, N379, N52, N915);
xor XOR2 (N978, N974, N655);
nand NAND3 (N979, N973, N604, N444);
and AND4 (N980, N964, N551, N145, N948);
buf BUF1 (N981, N970);
or OR4 (N982, N976, N236, N727, N92);
not NOT1 (N983, N982);
or OR3 (N984, N980, N572, N600);
buf BUF1 (N985, N978);
not NOT1 (N986, N977);
or OR3 (N987, N984, N16, N280);
buf BUF1 (N988, N953);
and AND3 (N989, N985, N97, N174);
and AND3 (N990, N983, N478, N561);
nand NAND3 (N991, N979, N471, N283);
or OR3 (N992, N981, N211, N204);
buf BUF1 (N993, N991);
and AND4 (N994, N992, N942, N702, N379);
and AND3 (N995, N987, N297, N742);
nor NOR2 (N996, N988, N946);
not NOT1 (N997, N971);
not NOT1 (N998, N994);
buf BUF1 (N999, N998);
buf BUF1 (N1000, N995);
buf BUF1 (N1001, N999);
xor XOR2 (N1002, N986, N801);
and AND3 (N1003, N968, N897, N478);
buf BUF1 (N1004, N1000);
and AND4 (N1005, N1001, N274, N263, N690);
nor NOR4 (N1006, N1005, N461, N206, N317);
nor NOR2 (N1007, N975, N824);
and AND3 (N1008, N1007, N539, N128);
or OR3 (N1009, N1008, N757, N140);
not NOT1 (N1010, N997);
nor NOR4 (N1011, N1003, N591, N885, N107);
nor NOR2 (N1012, N996, N8);
nor NOR2 (N1013, N1006, N769);
not NOT1 (N1014, N1009);
xor XOR2 (N1015, N990, N984);
nand NAND4 (N1016, N1004, N757, N737, N133);
or OR3 (N1017, N1014, N5, N362);
not NOT1 (N1018, N1002);
not NOT1 (N1019, N1018);
buf BUF1 (N1020, N1010);
not NOT1 (N1021, N989);
or OR4 (N1022, N1011, N571, N60, N896);
or OR2 (N1023, N1020, N413);
buf BUF1 (N1024, N1012);
nand NAND4 (N1025, N993, N979, N73, N270);
or OR2 (N1026, N1022, N159);
xor XOR2 (N1027, N1016, N618);
buf BUF1 (N1028, N1013);
buf BUF1 (N1029, N1015);
and AND2 (N1030, N1024, N674);
not NOT1 (N1031, N1023);
buf BUF1 (N1032, N1021);
not NOT1 (N1033, N1029);
not NOT1 (N1034, N1019);
xor XOR2 (N1035, N1033, N985);
nor NOR2 (N1036, N1034, N47);
buf BUF1 (N1037, N1035);
buf BUF1 (N1038, N1031);
and AND3 (N1039, N1028, N258, N952);
xor XOR2 (N1040, N1037, N435);
not NOT1 (N1041, N1026);
buf BUF1 (N1042, N1038);
and AND4 (N1043, N1025, N678, N439, N391);
nor NOR3 (N1044, N1039, N932, N467);
nand NAND3 (N1045, N1040, N995, N29);
buf BUF1 (N1046, N1043);
or OR2 (N1047, N1042, N4);
and AND4 (N1048, N1030, N833, N984, N380);
buf BUF1 (N1049, N1032);
buf BUF1 (N1050, N1049);
buf BUF1 (N1051, N1048);
not NOT1 (N1052, N1017);
nor NOR3 (N1053, N1044, N814, N172);
xor XOR2 (N1054, N1046, N337);
buf BUF1 (N1055, N1041);
and AND3 (N1056, N1045, N54, N1001);
buf BUF1 (N1057, N1056);
nor NOR2 (N1058, N1054, N105);
xor XOR2 (N1059, N1058, N438);
and AND3 (N1060, N1050, N968, N683);
xor XOR2 (N1061, N1047, N396);
not NOT1 (N1062, N1052);
not NOT1 (N1063, N1057);
nor NOR3 (N1064, N1062, N748, N974);
xor XOR2 (N1065, N1051, N175);
nor NOR4 (N1066, N1059, N325, N735, N933);
or OR2 (N1067, N1053, N953);
xor XOR2 (N1068, N1067, N670);
and AND2 (N1069, N1055, N491);
nor NOR4 (N1070, N1060, N603, N888, N293);
xor XOR2 (N1071, N1065, N703);
not NOT1 (N1072, N1064);
buf BUF1 (N1073, N1027);
nand NAND4 (N1074, N1061, N446, N511, N502);
xor XOR2 (N1075, N1073, N121);
buf BUF1 (N1076, N1068);
xor XOR2 (N1077, N1066, N221);
not NOT1 (N1078, N1077);
buf BUF1 (N1079, N1063);
nor NOR4 (N1080, N1074, N160, N37, N736);
nor NOR2 (N1081, N1071, N521);
buf BUF1 (N1082, N1036);
nand NAND3 (N1083, N1082, N733, N523);
not NOT1 (N1084, N1076);
buf BUF1 (N1085, N1075);
or OR3 (N1086, N1080, N909, N616);
not NOT1 (N1087, N1084);
buf BUF1 (N1088, N1085);
xor XOR2 (N1089, N1079, N195);
buf BUF1 (N1090, N1088);
nand NAND3 (N1091, N1090, N287, N1074);
and AND2 (N1092, N1072, N171);
nand NAND4 (N1093, N1078, N930, N563, N468);
or OR2 (N1094, N1091, N241);
or OR3 (N1095, N1069, N736, N570);
nor NOR4 (N1096, N1081, N242, N770, N239);
not NOT1 (N1097, N1087);
and AND3 (N1098, N1092, N684, N621);
xor XOR2 (N1099, N1089, N361);
xor XOR2 (N1100, N1094, N713);
and AND3 (N1101, N1100, N908, N409);
or OR4 (N1102, N1086, N979, N431, N1027);
and AND3 (N1103, N1102, N862, N462);
nand NAND3 (N1104, N1070, N392, N204);
xor XOR2 (N1105, N1083, N556);
not NOT1 (N1106, N1104);
xor XOR2 (N1107, N1106, N632);
buf BUF1 (N1108, N1093);
xor XOR2 (N1109, N1097, N1080);
nand NAND4 (N1110, N1105, N407, N544, N100);
nand NAND3 (N1111, N1109, N465, N841);
buf BUF1 (N1112, N1108);
or OR4 (N1113, N1098, N744, N709, N1009);
buf BUF1 (N1114, N1111);
nor NOR3 (N1115, N1099, N611, N68);
not NOT1 (N1116, N1110);
not NOT1 (N1117, N1107);
not NOT1 (N1118, N1115);
nor NOR4 (N1119, N1113, N1004, N344, N289);
xor XOR2 (N1120, N1095, N1111);
or OR4 (N1121, N1112, N1068, N1013, N256);
and AND3 (N1122, N1116, N1115, N718);
and AND2 (N1123, N1121, N639);
buf BUF1 (N1124, N1122);
nand NAND4 (N1125, N1118, N66, N870, N824);
or OR2 (N1126, N1123, N742);
or OR3 (N1127, N1124, N463, N745);
buf BUF1 (N1128, N1119);
buf BUF1 (N1129, N1114);
not NOT1 (N1130, N1128);
or OR3 (N1131, N1096, N112, N647);
nand NAND2 (N1132, N1120, N745);
nand NAND4 (N1133, N1129, N705, N941, N323);
nand NAND3 (N1134, N1131, N335, N164);
or OR4 (N1135, N1132, N740, N279, N670);
xor XOR2 (N1136, N1127, N153);
buf BUF1 (N1137, N1103);
and AND3 (N1138, N1135, N803, N1128);
or OR3 (N1139, N1125, N373, N222);
xor XOR2 (N1140, N1134, N485);
and AND2 (N1141, N1137, N488);
not NOT1 (N1142, N1136);
not NOT1 (N1143, N1130);
xor XOR2 (N1144, N1133, N746);
and AND4 (N1145, N1101, N429, N188, N194);
or OR4 (N1146, N1126, N24, N983, N180);
nand NAND2 (N1147, N1140, N71);
not NOT1 (N1148, N1142);
nor NOR4 (N1149, N1143, N930, N333, N158);
or OR4 (N1150, N1138, N436, N760, N98);
xor XOR2 (N1151, N1149, N368);
xor XOR2 (N1152, N1141, N645);
nand NAND2 (N1153, N1150, N1092);
nor NOR3 (N1154, N1148, N1086, N982);
and AND4 (N1155, N1152, N1135, N1056, N864);
nor NOR3 (N1156, N1154, N269, N407);
not NOT1 (N1157, N1153);
nor NOR4 (N1158, N1145, N300, N481, N588);
nand NAND4 (N1159, N1155, N675, N854, N424);
xor XOR2 (N1160, N1158, N345);
nor NOR4 (N1161, N1157, N329, N958, N255);
or OR4 (N1162, N1139, N668, N927, N237);
xor XOR2 (N1163, N1151, N503);
nand NAND3 (N1164, N1146, N424, N678);
and AND2 (N1165, N1159, N770);
nand NAND2 (N1166, N1117, N454);
nor NOR3 (N1167, N1163, N930, N60);
not NOT1 (N1168, N1162);
and AND4 (N1169, N1147, N596, N352, N1024);
or OR2 (N1170, N1161, N969);
not NOT1 (N1171, N1168);
and AND3 (N1172, N1164, N888, N205);
nor NOR2 (N1173, N1169, N818);
buf BUF1 (N1174, N1156);
xor XOR2 (N1175, N1167, N698);
nand NAND4 (N1176, N1170, N614, N720, N647);
or OR3 (N1177, N1171, N799, N992);
and AND3 (N1178, N1172, N325, N188);
nor NOR2 (N1179, N1175, N357);
nor NOR3 (N1180, N1160, N915, N484);
and AND4 (N1181, N1144, N524, N823, N468);
nor NOR2 (N1182, N1181, N982);
not NOT1 (N1183, N1177);
xor XOR2 (N1184, N1182, N1181);
and AND2 (N1185, N1166, N423);
and AND4 (N1186, N1183, N172, N37, N137);
buf BUF1 (N1187, N1180);
or OR4 (N1188, N1178, N1041, N619, N1088);
and AND4 (N1189, N1187, N785, N777, N508);
and AND2 (N1190, N1184, N57);
nand NAND2 (N1191, N1165, N869);
or OR3 (N1192, N1186, N157, N488);
buf BUF1 (N1193, N1176);
not NOT1 (N1194, N1174);
nor NOR4 (N1195, N1192, N791, N484, N306);
not NOT1 (N1196, N1191);
and AND3 (N1197, N1194, N444, N513);
buf BUF1 (N1198, N1195);
xor XOR2 (N1199, N1197, N16);
nand NAND3 (N1200, N1185, N734, N508);
nand NAND3 (N1201, N1196, N48, N487);
or OR2 (N1202, N1200, N230);
and AND2 (N1203, N1189, N689);
not NOT1 (N1204, N1203);
and AND4 (N1205, N1199, N1121, N57, N344);
and AND2 (N1206, N1188, N815);
not NOT1 (N1207, N1193);
buf BUF1 (N1208, N1206);
not NOT1 (N1209, N1208);
buf BUF1 (N1210, N1205);
not NOT1 (N1211, N1210);
buf BUF1 (N1212, N1179);
nor NOR3 (N1213, N1202, N331, N1135);
and AND3 (N1214, N1207, N1167, N781);
not NOT1 (N1215, N1173);
not NOT1 (N1216, N1204);
buf BUF1 (N1217, N1216);
nor NOR3 (N1218, N1213, N9, N499);
xor XOR2 (N1219, N1217, N410);
not NOT1 (N1220, N1215);
buf BUF1 (N1221, N1201);
xor XOR2 (N1222, N1214, N1020);
nor NOR2 (N1223, N1222, N947);
nor NOR2 (N1224, N1190, N80);
or OR4 (N1225, N1224, N643, N461, N498);
nor NOR4 (N1226, N1198, N943, N1047, N214);
xor XOR2 (N1227, N1212, N680);
nor NOR2 (N1228, N1219, N872);
and AND2 (N1229, N1228, N846);
nor NOR3 (N1230, N1218, N657, N150);
buf BUF1 (N1231, N1221);
and AND4 (N1232, N1223, N1152, N88, N1024);
nand NAND2 (N1233, N1211, N154);
or OR4 (N1234, N1227, N332, N356, N837);
xor XOR2 (N1235, N1232, N479);
or OR2 (N1236, N1234, N379);
xor XOR2 (N1237, N1229, N323);
or OR4 (N1238, N1226, N588, N942, N967);
and AND3 (N1239, N1237, N206, N269);
nand NAND4 (N1240, N1220, N44, N1117, N886);
nand NAND3 (N1241, N1209, N653, N848);
xor XOR2 (N1242, N1238, N382);
xor XOR2 (N1243, N1233, N845);
or OR2 (N1244, N1242, N303);
buf BUF1 (N1245, N1240);
not NOT1 (N1246, N1235);
nand NAND3 (N1247, N1236, N187, N697);
nand NAND2 (N1248, N1247, N1209);
buf BUF1 (N1249, N1246);
buf BUF1 (N1250, N1248);
not NOT1 (N1251, N1239);
or OR3 (N1252, N1249, N418, N1207);
not NOT1 (N1253, N1231);
or OR2 (N1254, N1251, N99);
nand NAND3 (N1255, N1244, N53, N447);
not NOT1 (N1256, N1230);
xor XOR2 (N1257, N1255, N1251);
and AND2 (N1258, N1252, N282);
nand NAND3 (N1259, N1257, N91, N860);
and AND2 (N1260, N1250, N778);
nor NOR4 (N1261, N1253, N88, N989, N850);
or OR2 (N1262, N1259, N510);
buf BUF1 (N1263, N1260);
nand NAND3 (N1264, N1258, N899, N1241);
buf BUF1 (N1265, N152);
xor XOR2 (N1266, N1262, N1262);
nor NOR3 (N1267, N1261, N641, N557);
not NOT1 (N1268, N1245);
or OR3 (N1269, N1265, N257, N1048);
xor XOR2 (N1270, N1256, N883);
and AND4 (N1271, N1264, N856, N712, N810);
or OR4 (N1272, N1243, N591, N84, N851);
buf BUF1 (N1273, N1263);
xor XOR2 (N1274, N1266, N1225);
xor XOR2 (N1275, N1071, N229);
nand NAND2 (N1276, N1270, N170);
nand NAND3 (N1277, N1267, N758, N927);
nand NAND3 (N1278, N1269, N1136, N495);
buf BUF1 (N1279, N1276);
or OR3 (N1280, N1277, N608, N1212);
or OR3 (N1281, N1275, N950, N194);
not NOT1 (N1282, N1273);
xor XOR2 (N1283, N1278, N547);
not NOT1 (N1284, N1282);
nor NOR3 (N1285, N1280, N1226, N41);
not NOT1 (N1286, N1271);
or OR3 (N1287, N1286, N997, N211);
and AND3 (N1288, N1279, N658, N1188);
or OR3 (N1289, N1285, N23, N373);
or OR2 (N1290, N1287, N1192);
nand NAND3 (N1291, N1283, N1064, N1125);
xor XOR2 (N1292, N1290, N416);
xor XOR2 (N1293, N1274, N732);
nand NAND2 (N1294, N1272, N415);
xor XOR2 (N1295, N1254, N917);
not NOT1 (N1296, N1281);
xor XOR2 (N1297, N1293, N548);
nand NAND4 (N1298, N1294, N57, N970, N422);
and AND2 (N1299, N1288, N367);
xor XOR2 (N1300, N1299, N788);
buf BUF1 (N1301, N1284);
xor XOR2 (N1302, N1292, N19);
nand NAND4 (N1303, N1295, N669, N443, N1233);
not NOT1 (N1304, N1301);
and AND4 (N1305, N1304, N1185, N1097, N686);
nor NOR4 (N1306, N1302, N695, N698, N703);
not NOT1 (N1307, N1296);
xor XOR2 (N1308, N1305, N984);
nand NAND2 (N1309, N1291, N1007);
and AND4 (N1310, N1307, N645, N144, N28);
and AND3 (N1311, N1300, N1289, N340);
and AND4 (N1312, N524, N65, N1177, N1197);
buf BUF1 (N1313, N1310);
or OR2 (N1314, N1298, N347);
not NOT1 (N1315, N1268);
not NOT1 (N1316, N1314);
nor NOR2 (N1317, N1316, N1290);
not NOT1 (N1318, N1303);
nand NAND3 (N1319, N1315, N335, N1044);
xor XOR2 (N1320, N1317, N1297);
and AND3 (N1321, N947, N477, N1155);
nand NAND2 (N1322, N1318, N915);
and AND4 (N1323, N1320, N954, N139, N1093);
xor XOR2 (N1324, N1319, N627);
and AND3 (N1325, N1308, N796, N47);
nand NAND3 (N1326, N1312, N502, N312);
nor NOR2 (N1327, N1306, N527);
xor XOR2 (N1328, N1322, N143);
nand NAND2 (N1329, N1325, N220);
not NOT1 (N1330, N1321);
not NOT1 (N1331, N1313);
nor NOR2 (N1332, N1330, N749);
nand NAND3 (N1333, N1324, N1312, N125);
buf BUF1 (N1334, N1332);
nand NAND4 (N1335, N1323, N909, N1149, N767);
buf BUF1 (N1336, N1328);
nor NOR4 (N1337, N1335, N166, N87, N690);
buf BUF1 (N1338, N1309);
and AND4 (N1339, N1336, N1216, N938, N523);
nor NOR2 (N1340, N1326, N286);
nand NAND2 (N1341, N1333, N535);
not NOT1 (N1342, N1341);
and AND4 (N1343, N1334, N571, N11, N970);
and AND3 (N1344, N1338, N156, N223);
or OR2 (N1345, N1329, N46);
not NOT1 (N1346, N1337);
xor XOR2 (N1347, N1340, N216);
nand NAND3 (N1348, N1346, N1051, N437);
xor XOR2 (N1349, N1339, N107);
nor NOR2 (N1350, N1345, N18);
nor NOR4 (N1351, N1350, N236, N372, N844);
nor NOR3 (N1352, N1348, N700, N1104);
xor XOR2 (N1353, N1342, N1172);
and AND2 (N1354, N1343, N1176);
nand NAND4 (N1355, N1327, N964, N539, N85);
or OR2 (N1356, N1354, N597);
nor NOR2 (N1357, N1356, N1114);
not NOT1 (N1358, N1357);
and AND2 (N1359, N1349, N325);
and AND4 (N1360, N1352, N913, N1062, N1339);
not NOT1 (N1361, N1347);
nor NOR2 (N1362, N1331, N796);
nor NOR4 (N1363, N1351, N874, N298, N748);
or OR4 (N1364, N1362, N1091, N128, N493);
not NOT1 (N1365, N1364);
or OR4 (N1366, N1355, N578, N1200, N1301);
not NOT1 (N1367, N1311);
and AND3 (N1368, N1367, N179, N290);
buf BUF1 (N1369, N1366);
nor NOR2 (N1370, N1359, N321);
or OR2 (N1371, N1361, N915);
xor XOR2 (N1372, N1371, N1109);
not NOT1 (N1373, N1372);
xor XOR2 (N1374, N1370, N1190);
nand NAND4 (N1375, N1373, N1269, N1137, N1354);
buf BUF1 (N1376, N1374);
buf BUF1 (N1377, N1360);
nand NAND3 (N1378, N1363, N1203, N723);
buf BUF1 (N1379, N1353);
and AND2 (N1380, N1369, N375);
nor NOR4 (N1381, N1344, N339, N1001, N1039);
not NOT1 (N1382, N1377);
xor XOR2 (N1383, N1378, N992);
or OR2 (N1384, N1358, N163);
or OR2 (N1385, N1376, N1178);
nor NOR3 (N1386, N1382, N1014, N1025);
and AND2 (N1387, N1383, N189);
nand NAND4 (N1388, N1379, N401, N898, N355);
not NOT1 (N1389, N1387);
not NOT1 (N1390, N1380);
or OR4 (N1391, N1386, N885, N940, N156);
or OR3 (N1392, N1375, N172, N1358);
nand NAND2 (N1393, N1385, N797);
nand NAND3 (N1394, N1365, N9, N138);
not NOT1 (N1395, N1381);
nor NOR4 (N1396, N1384, N1081, N15, N425);
buf BUF1 (N1397, N1396);
buf BUF1 (N1398, N1390);
nand NAND4 (N1399, N1391, N1170, N1340, N1006);
xor XOR2 (N1400, N1398, N820);
or OR2 (N1401, N1389, N1229);
or OR2 (N1402, N1399, N635);
and AND2 (N1403, N1395, N324);
buf BUF1 (N1404, N1393);
nor NOR2 (N1405, N1400, N1199);
buf BUF1 (N1406, N1368);
or OR2 (N1407, N1405, N506);
nor NOR3 (N1408, N1397, N488, N934);
nor NOR3 (N1409, N1388, N381, N412);
xor XOR2 (N1410, N1408, N497);
nand NAND3 (N1411, N1410, N309, N803);
nand NAND2 (N1412, N1402, N1171);
xor XOR2 (N1413, N1403, N838);
nor NOR4 (N1414, N1406, N1122, N1030, N875);
and AND4 (N1415, N1412, N1119, N914, N627);
xor XOR2 (N1416, N1414, N357);
xor XOR2 (N1417, N1407, N912);
or OR4 (N1418, N1409, N739, N116, N1308);
or OR2 (N1419, N1394, N355);
or OR2 (N1420, N1413, N385);
or OR4 (N1421, N1401, N1261, N447, N798);
or OR2 (N1422, N1392, N153);
and AND3 (N1423, N1404, N299, N1409);
xor XOR2 (N1424, N1415, N175);
and AND3 (N1425, N1417, N556, N494);
nor NOR4 (N1426, N1419, N265, N1303, N1012);
or OR3 (N1427, N1411, N368, N1233);
nor NOR3 (N1428, N1418, N117, N1008);
nor NOR4 (N1429, N1428, N439, N654, N706);
nor NOR2 (N1430, N1424, N271);
nand NAND3 (N1431, N1422, N884, N1196);
xor XOR2 (N1432, N1429, N893);
and AND4 (N1433, N1430, N1400, N3, N361);
or OR3 (N1434, N1425, N257, N683);
or OR3 (N1435, N1433, N179, N1257);
nor NOR4 (N1436, N1416, N1019, N338, N949);
xor XOR2 (N1437, N1426, N32);
nand NAND3 (N1438, N1431, N364, N1054);
and AND3 (N1439, N1420, N31, N242);
nor NOR4 (N1440, N1439, N1217, N255, N1031);
buf BUF1 (N1441, N1427);
nor NOR4 (N1442, N1436, N70, N974, N1293);
nand NAND2 (N1443, N1437, N1243);
buf BUF1 (N1444, N1435);
not NOT1 (N1445, N1443);
or OR4 (N1446, N1441, N802, N1101, N903);
buf BUF1 (N1447, N1442);
not NOT1 (N1448, N1446);
nor NOR4 (N1449, N1432, N1129, N927, N197);
not NOT1 (N1450, N1449);
nor NOR4 (N1451, N1440, N937, N535, N632);
nor NOR2 (N1452, N1447, N176);
not NOT1 (N1453, N1450);
xor XOR2 (N1454, N1444, N207);
nand NAND3 (N1455, N1454, N538, N898);
buf BUF1 (N1456, N1423);
or OR2 (N1457, N1434, N224);
xor XOR2 (N1458, N1456, N1186);
nand NAND2 (N1459, N1421, N1128);
nor NOR2 (N1460, N1451, N1449);
xor XOR2 (N1461, N1448, N546);
nand NAND4 (N1462, N1445, N907, N34, N691);
xor XOR2 (N1463, N1438, N827);
or OR3 (N1464, N1458, N1301, N1097);
not NOT1 (N1465, N1452);
not NOT1 (N1466, N1462);
nor NOR3 (N1467, N1455, N647, N1377);
xor XOR2 (N1468, N1460, N603);
nand NAND4 (N1469, N1465, N1032, N1442, N700);
and AND2 (N1470, N1466, N764);
buf BUF1 (N1471, N1467);
xor XOR2 (N1472, N1457, N1239);
xor XOR2 (N1473, N1453, N1400);
xor XOR2 (N1474, N1459, N1316);
and AND3 (N1475, N1470, N862, N473);
or OR3 (N1476, N1464, N430, N951);
nand NAND3 (N1477, N1475, N62, N997);
or OR3 (N1478, N1463, N603, N762);
and AND2 (N1479, N1461, N1332);
nand NAND3 (N1480, N1474, N1367, N1078);
buf BUF1 (N1481, N1477);
nand NAND2 (N1482, N1473, N381);
nand NAND2 (N1483, N1478, N1461);
and AND2 (N1484, N1479, N58);
and AND4 (N1485, N1468, N368, N122, N1059);
not NOT1 (N1486, N1482);
or OR3 (N1487, N1472, N201, N40);
nand NAND2 (N1488, N1483, N160);
and AND2 (N1489, N1484, N165);
and AND3 (N1490, N1480, N1284, N923);
nand NAND2 (N1491, N1481, N125);
nand NAND3 (N1492, N1488, N213, N1348);
nor NOR4 (N1493, N1490, N644, N546, N146);
xor XOR2 (N1494, N1489, N664);
buf BUF1 (N1495, N1492);
and AND3 (N1496, N1476, N188, N2);
nand NAND4 (N1497, N1496, N440, N1298, N871);
buf BUF1 (N1498, N1491);
nor NOR4 (N1499, N1487, N1213, N934, N1205);
or OR3 (N1500, N1499, N1240, N441);
nand NAND2 (N1501, N1500, N611);
and AND4 (N1502, N1495, N1129, N691, N1249);
xor XOR2 (N1503, N1485, N500);
not NOT1 (N1504, N1497);
and AND4 (N1505, N1471, N443, N1475, N711);
buf BUF1 (N1506, N1503);
and AND4 (N1507, N1501, N836, N139, N466);
or OR2 (N1508, N1504, N71);
buf BUF1 (N1509, N1502);
not NOT1 (N1510, N1498);
nand NAND3 (N1511, N1469, N755, N1081);
or OR2 (N1512, N1509, N84);
and AND2 (N1513, N1510, N788);
not NOT1 (N1514, N1511);
buf BUF1 (N1515, N1507);
buf BUF1 (N1516, N1513);
nor NOR2 (N1517, N1505, N1081);
not NOT1 (N1518, N1516);
endmodule