// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N2017,N2020,N2021,N2015,N2007,N1997,N2002,N2018,N2008,N2022;

nor NOR3 (N23, N15, N9, N16);
and AND3 (N24, N12, N4, N5);
or OR4 (N25, N15, N20, N15, N5);
and AND3 (N26, N7, N15, N16);
not NOT1 (N27, N13);
or OR3 (N28, N24, N20, N19);
nor NOR2 (N29, N6, N18);
and AND4 (N30, N8, N18, N18, N12);
or OR3 (N31, N7, N11, N28);
xor XOR2 (N32, N20, N12);
buf BUF1 (N33, N13);
buf BUF1 (N34, N18);
or OR2 (N35, N32, N21);
nand NAND3 (N36, N27, N11, N30);
or OR2 (N37, N27, N36);
nand NAND4 (N38, N8, N8, N21, N18);
xor XOR2 (N39, N33, N24);
buf BUF1 (N40, N23);
nor NOR4 (N41, N35, N37, N8, N31);
or OR3 (N42, N41, N8, N37);
not NOT1 (N43, N25);
not NOT1 (N44, N15);
nand NAND3 (N45, N24, N20, N20);
nor NOR3 (N46, N45, N11, N38);
nand NAND3 (N47, N11, N32, N32);
or OR2 (N48, N44, N28);
and AND3 (N49, N43, N7, N45);
nor NOR2 (N50, N42, N16);
xor XOR2 (N51, N47, N32);
not NOT1 (N52, N39);
nor NOR3 (N53, N46, N37, N46);
nand NAND4 (N54, N48, N14, N46, N35);
nor NOR3 (N55, N52, N8, N20);
or OR3 (N56, N26, N17, N1);
or OR4 (N57, N56, N37, N37, N23);
buf BUF1 (N58, N57);
or OR3 (N59, N55, N10, N23);
nand NAND3 (N60, N54, N22, N2);
and AND4 (N61, N49, N56, N53, N2);
buf BUF1 (N62, N7);
buf BUF1 (N63, N50);
nand NAND2 (N64, N60, N35);
or OR2 (N65, N64, N13);
or OR2 (N66, N61, N65);
not NOT1 (N67, N66);
nand NAND3 (N68, N10, N27, N33);
xor XOR2 (N69, N34, N37);
buf BUF1 (N70, N58);
and AND4 (N71, N67, N49, N26, N27);
or OR2 (N72, N68, N23);
nand NAND3 (N73, N69, N52, N53);
nor NOR4 (N74, N51, N10, N13, N69);
and AND2 (N75, N70, N50);
not NOT1 (N76, N62);
not NOT1 (N77, N76);
xor XOR2 (N78, N75, N29);
nor NOR4 (N79, N43, N66, N52, N25);
and AND4 (N80, N40, N57, N20, N66);
buf BUF1 (N81, N80);
buf BUF1 (N82, N79);
or OR3 (N83, N81, N36, N73);
nor NOR4 (N84, N78, N20, N14, N11);
not NOT1 (N85, N79);
nand NAND2 (N86, N85, N50);
buf BUF1 (N87, N59);
nor NOR3 (N88, N74, N30, N52);
not NOT1 (N89, N84);
nand NAND2 (N90, N87, N72);
xor XOR2 (N91, N30, N14);
or OR3 (N92, N86, N66, N22);
xor XOR2 (N93, N77, N53);
nor NOR2 (N94, N82, N9);
xor XOR2 (N95, N90, N25);
buf BUF1 (N96, N88);
xor XOR2 (N97, N63, N61);
nand NAND3 (N98, N91, N61, N77);
and AND3 (N99, N94, N18, N29);
and AND2 (N100, N93, N67);
buf BUF1 (N101, N97);
and AND3 (N102, N71, N94, N38);
buf BUF1 (N103, N102);
nor NOR4 (N104, N103, N99, N26, N101);
xor XOR2 (N105, N12, N18);
nor NOR2 (N106, N21, N23);
or OR2 (N107, N96, N40);
buf BUF1 (N108, N105);
nor NOR2 (N109, N98, N72);
not NOT1 (N110, N83);
and AND3 (N111, N104, N44, N73);
nand NAND2 (N112, N106, N12);
buf BUF1 (N113, N100);
buf BUF1 (N114, N109);
or OR3 (N115, N108, N87, N10);
xor XOR2 (N116, N113, N113);
or OR4 (N117, N115, N19, N73, N40);
xor XOR2 (N118, N114, N95);
not NOT1 (N119, N118);
nand NAND3 (N120, N119, N117, N62);
and AND4 (N121, N10, N49, N94, N98);
buf BUF1 (N122, N22);
or OR4 (N123, N116, N39, N95, N15);
and AND2 (N124, N112, N33);
and AND2 (N125, N122, N10);
and AND3 (N126, N120, N37, N88);
or OR4 (N127, N126, N91, N101, N121);
and AND2 (N128, N74, N93);
or OR3 (N129, N107, N77, N126);
buf BUF1 (N130, N129);
not NOT1 (N131, N127);
nand NAND4 (N132, N124, N70, N45, N95);
not NOT1 (N133, N92);
or OR2 (N134, N125, N41);
buf BUF1 (N135, N123);
nand NAND4 (N136, N111, N133, N111, N113);
xor XOR2 (N137, N46, N68);
nor NOR2 (N138, N134, N121);
nor NOR2 (N139, N136, N94);
nor NOR2 (N140, N128, N5);
and AND2 (N141, N130, N106);
or OR2 (N142, N137, N19);
or OR3 (N143, N135, N130, N45);
nor NOR4 (N144, N142, N59, N100, N63);
nand NAND4 (N145, N131, N57, N40, N102);
and AND4 (N146, N144, N100, N57, N71);
or OR2 (N147, N132, N45);
xor XOR2 (N148, N140, N13);
nand NAND4 (N149, N147, N104, N97, N83);
nand NAND3 (N150, N143, N149, N18);
not NOT1 (N151, N145);
nor NOR2 (N152, N151, N13);
xor XOR2 (N153, N39, N69);
or OR2 (N154, N89, N30);
not NOT1 (N155, N150);
xor XOR2 (N156, N155, N3);
xor XOR2 (N157, N153, N59);
nand NAND3 (N158, N152, N86, N96);
buf BUF1 (N159, N157);
or OR3 (N160, N110, N86, N35);
nand NAND3 (N161, N139, N140, N112);
or OR4 (N162, N141, N17, N119, N37);
nand NAND4 (N163, N156, N70, N74, N144);
xor XOR2 (N164, N138, N131);
and AND2 (N165, N162, N66);
xor XOR2 (N166, N158, N23);
xor XOR2 (N167, N165, N92);
buf BUF1 (N168, N154);
not NOT1 (N169, N159);
or OR3 (N170, N148, N80, N154);
buf BUF1 (N171, N160);
nor NOR4 (N172, N171, N81, N77, N167);
and AND3 (N173, N168, N12, N100);
and AND4 (N174, N131, N171, N57, N31);
buf BUF1 (N175, N170);
nand NAND2 (N176, N175, N30);
or OR2 (N177, N163, N89);
buf BUF1 (N178, N169);
or OR3 (N179, N176, N59, N39);
nand NAND4 (N180, N172, N150, N95, N5);
buf BUF1 (N181, N180);
and AND3 (N182, N164, N156, N113);
and AND3 (N183, N181, N129, N22);
not NOT1 (N184, N161);
buf BUF1 (N185, N174);
and AND4 (N186, N182, N113, N50, N32);
xor XOR2 (N187, N146, N50);
buf BUF1 (N188, N179);
xor XOR2 (N189, N166, N172);
or OR2 (N190, N184, N114);
buf BUF1 (N191, N187);
nor NOR2 (N192, N183, N68);
nor NOR2 (N193, N189, N137);
buf BUF1 (N194, N173);
or OR3 (N195, N192, N123, N99);
or OR4 (N196, N177, N167, N104, N88);
buf BUF1 (N197, N195);
nand NAND2 (N198, N188, N126);
and AND2 (N199, N185, N3);
not NOT1 (N200, N186);
xor XOR2 (N201, N191, N3);
nor NOR4 (N202, N200, N75, N5, N142);
buf BUF1 (N203, N196);
and AND3 (N204, N202, N84, N178);
not NOT1 (N205, N137);
buf BUF1 (N206, N201);
xor XOR2 (N207, N197, N79);
not NOT1 (N208, N198);
not NOT1 (N209, N204);
or OR3 (N210, N203, N134, N44);
xor XOR2 (N211, N205, N16);
nor NOR3 (N212, N206, N129, N37);
or OR4 (N213, N208, N80, N129, N13);
buf BUF1 (N214, N190);
buf BUF1 (N215, N211);
nor NOR4 (N216, N193, N108, N191, N194);
nand NAND2 (N217, N59, N180);
not NOT1 (N218, N212);
nand NAND2 (N219, N213, N92);
or OR2 (N220, N214, N134);
and AND4 (N221, N218, N170, N182, N142);
nand NAND4 (N222, N199, N56, N201, N30);
or OR4 (N223, N217, N218, N90, N71);
nor NOR4 (N224, N216, N66, N145, N9);
nand NAND4 (N225, N221, N172, N68, N60);
not NOT1 (N226, N215);
nand NAND2 (N227, N220, N108);
and AND2 (N228, N224, N45);
nand NAND3 (N229, N210, N146, N24);
or OR2 (N230, N225, N192);
nand NAND2 (N231, N228, N28);
nand NAND4 (N232, N229, N32, N145, N226);
nor NOR3 (N233, N38, N169, N178);
and AND2 (N234, N209, N148);
nor NOR4 (N235, N227, N180, N85, N52);
nor NOR3 (N236, N223, N205, N64);
not NOT1 (N237, N207);
buf BUF1 (N238, N219);
buf BUF1 (N239, N234);
nor NOR3 (N240, N237, N132, N184);
buf BUF1 (N241, N238);
nand NAND4 (N242, N236, N189, N124, N22);
and AND2 (N243, N231, N27);
or OR2 (N244, N233, N194);
buf BUF1 (N245, N239);
and AND2 (N246, N230, N184);
xor XOR2 (N247, N235, N128);
xor XOR2 (N248, N246, N232);
and AND3 (N249, N178, N213, N115);
nand NAND2 (N250, N245, N2);
nor NOR4 (N251, N241, N144, N174, N125);
xor XOR2 (N252, N240, N136);
and AND3 (N253, N244, N206, N182);
and AND3 (N254, N248, N128, N215);
and AND3 (N255, N242, N183, N26);
nor NOR2 (N256, N253, N209);
or OR3 (N257, N249, N250, N220);
xor XOR2 (N258, N180, N28);
xor XOR2 (N259, N258, N141);
nand NAND4 (N260, N254, N118, N11, N129);
and AND3 (N261, N251, N257, N253);
buf BUF1 (N262, N28);
and AND2 (N263, N259, N257);
not NOT1 (N264, N260);
or OR2 (N265, N261, N129);
or OR4 (N266, N252, N155, N73, N219);
nand NAND3 (N267, N266, N11, N106);
nand NAND4 (N268, N243, N263, N1, N47);
not NOT1 (N269, N235);
nand NAND3 (N270, N222, N253, N249);
buf BUF1 (N271, N255);
or OR2 (N272, N247, N207);
nand NAND2 (N273, N265, N110);
not NOT1 (N274, N269);
xor XOR2 (N275, N256, N274);
and AND3 (N276, N192, N235, N231);
buf BUF1 (N277, N273);
not NOT1 (N278, N276);
buf BUF1 (N279, N267);
or OR3 (N280, N272, N107, N187);
and AND2 (N281, N275, N165);
and AND2 (N282, N279, N232);
buf BUF1 (N283, N268);
not NOT1 (N284, N262);
and AND2 (N285, N281, N85);
buf BUF1 (N286, N264);
xor XOR2 (N287, N286, N144);
xor XOR2 (N288, N284, N245);
not NOT1 (N289, N288);
not NOT1 (N290, N271);
buf BUF1 (N291, N280);
nand NAND2 (N292, N278, N118);
not NOT1 (N293, N290);
or OR4 (N294, N282, N68, N133, N79);
not NOT1 (N295, N292);
nor NOR3 (N296, N295, N190, N38);
buf BUF1 (N297, N294);
xor XOR2 (N298, N289, N36);
buf BUF1 (N299, N285);
nor NOR4 (N300, N297, N120, N175, N271);
not NOT1 (N301, N283);
nor NOR4 (N302, N298, N199, N149, N187);
nand NAND4 (N303, N293, N251, N42, N2);
not NOT1 (N304, N291);
nand NAND4 (N305, N304, N83, N214, N93);
xor XOR2 (N306, N300, N38);
nand NAND3 (N307, N299, N77, N70);
buf BUF1 (N308, N305);
buf BUF1 (N309, N306);
not NOT1 (N310, N301);
nor NOR4 (N311, N308, N162, N97, N55);
nor NOR2 (N312, N287, N44);
xor XOR2 (N313, N307, N299);
or OR4 (N314, N311, N160, N247, N162);
not NOT1 (N315, N309);
nor NOR4 (N316, N277, N277, N218, N125);
not NOT1 (N317, N296);
not NOT1 (N318, N317);
not NOT1 (N319, N314);
or OR3 (N320, N313, N108, N127);
not NOT1 (N321, N303);
xor XOR2 (N322, N320, N109);
xor XOR2 (N323, N310, N30);
or OR2 (N324, N321, N316);
buf BUF1 (N325, N175);
xor XOR2 (N326, N315, N67);
not NOT1 (N327, N325);
buf BUF1 (N328, N270);
nor NOR4 (N329, N324, N150, N167, N314);
not NOT1 (N330, N302);
nand NAND3 (N331, N322, N73, N191);
not NOT1 (N332, N318);
and AND2 (N333, N332, N39);
nor NOR3 (N334, N326, N122, N102);
nand NAND3 (N335, N330, N307, N102);
not NOT1 (N336, N334);
buf BUF1 (N337, N329);
and AND2 (N338, N331, N233);
or OR4 (N339, N338, N6, N338, N333);
not NOT1 (N340, N327);
xor XOR2 (N341, N281, N80);
nand NAND2 (N342, N337, N164);
and AND4 (N343, N336, N139, N153, N177);
nand NAND4 (N344, N312, N172, N103, N260);
not NOT1 (N345, N319);
and AND2 (N346, N340, N196);
nor NOR3 (N347, N346, N132, N299);
buf BUF1 (N348, N323);
buf BUF1 (N349, N344);
or OR3 (N350, N343, N218, N178);
nor NOR2 (N351, N347, N117);
or OR2 (N352, N342, N337);
nand NAND2 (N353, N350, N330);
nor NOR3 (N354, N335, N237, N238);
not NOT1 (N355, N349);
xor XOR2 (N356, N341, N284);
not NOT1 (N357, N339);
or OR3 (N358, N352, N351, N22);
xor XOR2 (N359, N277, N336);
buf BUF1 (N360, N358);
buf BUF1 (N361, N357);
nand NAND2 (N362, N354, N116);
nor NOR3 (N363, N359, N158, N315);
and AND4 (N364, N360, N244, N112, N55);
xor XOR2 (N365, N353, N70);
nand NAND2 (N366, N364, N147);
nor NOR2 (N367, N348, N229);
and AND4 (N368, N361, N362, N154, N296);
nor NOR3 (N369, N152, N263, N318);
and AND4 (N370, N363, N366, N229, N95);
not NOT1 (N371, N24);
not NOT1 (N372, N356);
xor XOR2 (N373, N370, N265);
buf BUF1 (N374, N371);
nand NAND2 (N375, N328, N326);
and AND3 (N376, N367, N60, N208);
or OR4 (N377, N373, N6, N62, N79);
buf BUF1 (N378, N345);
xor XOR2 (N379, N374, N376);
or OR4 (N380, N245, N318, N99, N172);
not NOT1 (N381, N375);
buf BUF1 (N382, N369);
buf BUF1 (N383, N372);
nand NAND4 (N384, N377, N46, N57, N125);
or OR4 (N385, N368, N224, N289, N317);
or OR2 (N386, N384, N227);
buf BUF1 (N387, N382);
nor NOR4 (N388, N383, N41, N214, N386);
xor XOR2 (N389, N333, N178);
xor XOR2 (N390, N355, N13);
xor XOR2 (N391, N385, N4);
nor NOR2 (N392, N365, N258);
and AND3 (N393, N379, N351, N136);
and AND3 (N394, N381, N344, N150);
nand NAND2 (N395, N378, N49);
xor XOR2 (N396, N392, N118);
xor XOR2 (N397, N387, N74);
not NOT1 (N398, N388);
or OR3 (N399, N391, N208, N235);
and AND3 (N400, N394, N190, N134);
and AND3 (N401, N389, N5, N217);
not NOT1 (N402, N400);
xor XOR2 (N403, N395, N386);
buf BUF1 (N404, N399);
or OR3 (N405, N380, N167, N258);
not NOT1 (N406, N398);
not NOT1 (N407, N397);
and AND4 (N408, N406, N236, N104, N148);
xor XOR2 (N409, N408, N172);
not NOT1 (N410, N393);
xor XOR2 (N411, N404, N320);
xor XOR2 (N412, N396, N372);
not NOT1 (N413, N412);
not NOT1 (N414, N402);
nand NAND4 (N415, N390, N357, N253, N41);
nand NAND3 (N416, N409, N378, N240);
or OR3 (N417, N415, N207, N404);
xor XOR2 (N418, N405, N71);
nand NAND4 (N419, N413, N170, N365, N277);
nor NOR4 (N420, N401, N103, N395, N104);
not NOT1 (N421, N419);
and AND3 (N422, N414, N179, N161);
nand NAND3 (N423, N407, N240, N327);
or OR3 (N424, N421, N300, N347);
not NOT1 (N425, N420);
nand NAND4 (N426, N418, N136, N116, N374);
and AND2 (N427, N426, N42);
nand NAND3 (N428, N424, N309, N316);
and AND2 (N429, N411, N309);
not NOT1 (N430, N416);
xor XOR2 (N431, N422, N4);
or OR3 (N432, N428, N399, N219);
nand NAND3 (N433, N425, N291, N360);
xor XOR2 (N434, N431, N197);
buf BUF1 (N435, N429);
not NOT1 (N436, N423);
xor XOR2 (N437, N436, N396);
nand NAND4 (N438, N433, N403, N137, N205);
or OR2 (N439, N61, N386);
or OR3 (N440, N438, N225, N225);
and AND3 (N441, N434, N133, N129);
not NOT1 (N442, N430);
buf BUF1 (N443, N410);
nor NOR4 (N444, N441, N251, N356, N32);
nand NAND3 (N445, N437, N234, N369);
nand NAND4 (N446, N444, N280, N222, N341);
xor XOR2 (N447, N442, N158);
buf BUF1 (N448, N443);
nand NAND3 (N449, N427, N136, N127);
or OR3 (N450, N447, N318, N383);
or OR4 (N451, N450, N44, N184, N233);
buf BUF1 (N452, N439);
not NOT1 (N453, N440);
nand NAND2 (N454, N451, N24);
nand NAND3 (N455, N446, N17, N73);
not NOT1 (N456, N432);
and AND4 (N457, N456, N266, N89, N389);
or OR3 (N458, N454, N164, N8);
and AND2 (N459, N449, N209);
not NOT1 (N460, N417);
nor NOR2 (N461, N459, N4);
and AND3 (N462, N455, N457, N53);
nor NOR2 (N463, N131, N48);
xor XOR2 (N464, N460, N95);
and AND4 (N465, N461, N304, N331, N153);
not NOT1 (N466, N463);
nor NOR3 (N467, N465, N185, N296);
nand NAND3 (N468, N453, N19, N297);
and AND2 (N469, N462, N213);
buf BUF1 (N470, N445);
not NOT1 (N471, N470);
not NOT1 (N472, N458);
nand NAND4 (N473, N448, N430, N347, N49);
nand NAND4 (N474, N471, N330, N454, N50);
buf BUF1 (N475, N435);
nand NAND4 (N476, N475, N304, N471, N144);
not NOT1 (N477, N474);
nor NOR2 (N478, N464, N45);
xor XOR2 (N479, N466, N217);
and AND3 (N480, N472, N18, N27);
xor XOR2 (N481, N473, N276);
nand NAND3 (N482, N480, N158, N455);
buf BUF1 (N483, N479);
and AND3 (N484, N478, N245, N293);
nor NOR2 (N485, N482, N354);
nand NAND3 (N486, N485, N451, N472);
buf BUF1 (N487, N481);
or OR3 (N488, N452, N431, N30);
not NOT1 (N489, N484);
nand NAND4 (N490, N468, N153, N163, N384);
nor NOR2 (N491, N469, N298);
or OR2 (N492, N489, N281);
nand NAND4 (N493, N490, N92, N127, N388);
nand NAND3 (N494, N486, N171, N123);
xor XOR2 (N495, N493, N43);
xor XOR2 (N496, N467, N451);
and AND2 (N497, N494, N6);
not NOT1 (N498, N476);
xor XOR2 (N499, N492, N245);
nand NAND3 (N500, N488, N175, N97);
or OR3 (N501, N496, N224, N396);
not NOT1 (N502, N498);
nor NOR3 (N503, N477, N238, N221);
buf BUF1 (N504, N501);
nor NOR2 (N505, N487, N429);
xor XOR2 (N506, N502, N404);
nand NAND2 (N507, N497, N250);
or OR4 (N508, N503, N196, N309, N359);
and AND4 (N509, N507, N133, N212, N18);
not NOT1 (N510, N495);
and AND4 (N511, N509, N500, N142, N506);
and AND2 (N512, N220, N446);
nand NAND2 (N513, N290, N432);
nor NOR4 (N514, N510, N105, N411, N442);
xor XOR2 (N515, N511, N258);
xor XOR2 (N516, N504, N209);
or OR3 (N517, N499, N455, N110);
or OR2 (N518, N513, N495);
or OR3 (N519, N514, N465, N163);
not NOT1 (N520, N483);
not NOT1 (N521, N491);
or OR2 (N522, N515, N67);
nand NAND2 (N523, N508, N467);
xor XOR2 (N524, N517, N389);
xor XOR2 (N525, N505, N295);
or OR3 (N526, N524, N101, N187);
or OR3 (N527, N525, N110, N470);
nand NAND2 (N528, N522, N146);
and AND2 (N529, N526, N115);
not NOT1 (N530, N520);
not NOT1 (N531, N527);
not NOT1 (N532, N531);
or OR4 (N533, N528, N401, N525, N219);
buf BUF1 (N534, N533);
xor XOR2 (N535, N532, N27);
and AND3 (N536, N518, N216, N160);
not NOT1 (N537, N530);
xor XOR2 (N538, N536, N331);
nand NAND4 (N539, N534, N345, N161, N261);
not NOT1 (N540, N538);
nor NOR2 (N541, N523, N391);
nor NOR2 (N542, N521, N532);
and AND4 (N543, N539, N22, N227, N23);
buf BUF1 (N544, N535);
nor NOR3 (N545, N529, N353, N24);
buf BUF1 (N546, N512);
not NOT1 (N547, N546);
xor XOR2 (N548, N544, N463);
not NOT1 (N549, N548);
xor XOR2 (N550, N547, N162);
or OR3 (N551, N516, N433, N323);
not NOT1 (N552, N540);
xor XOR2 (N553, N537, N498);
or OR2 (N554, N553, N438);
buf BUF1 (N555, N549);
xor XOR2 (N556, N545, N146);
buf BUF1 (N557, N551);
nor NOR3 (N558, N543, N129, N203);
xor XOR2 (N559, N542, N135);
buf BUF1 (N560, N555);
nor NOR2 (N561, N560, N419);
and AND3 (N562, N559, N166, N504);
nand NAND2 (N563, N554, N549);
nand NAND2 (N564, N558, N375);
xor XOR2 (N565, N561, N17);
nor NOR2 (N566, N563, N29);
buf BUF1 (N567, N565);
and AND3 (N568, N566, N240, N554);
nand NAND2 (N569, N556, N8);
buf BUF1 (N570, N562);
not NOT1 (N571, N564);
buf BUF1 (N572, N552);
nor NOR2 (N573, N571, N567);
not NOT1 (N574, N547);
or OR2 (N575, N557, N269);
or OR3 (N576, N519, N134, N82);
or OR3 (N577, N575, N476, N9);
not NOT1 (N578, N568);
or OR4 (N579, N572, N488, N135, N333);
and AND4 (N580, N577, N422, N22, N567);
nand NAND3 (N581, N574, N363, N505);
nand NAND2 (N582, N576, N240);
and AND3 (N583, N569, N504, N370);
nand NAND4 (N584, N583, N564, N577, N133);
xor XOR2 (N585, N584, N53);
xor XOR2 (N586, N580, N430);
or OR2 (N587, N579, N562);
nand NAND4 (N588, N550, N204, N192, N394);
nor NOR2 (N589, N581, N247);
buf BUF1 (N590, N570);
or OR2 (N591, N573, N486);
and AND4 (N592, N589, N4, N190, N301);
nand NAND3 (N593, N582, N569, N565);
nand NAND4 (N594, N593, N346, N463, N51);
buf BUF1 (N595, N592);
xor XOR2 (N596, N587, N355);
xor XOR2 (N597, N588, N49);
nor NOR4 (N598, N591, N480, N229, N374);
nor NOR2 (N599, N595, N110);
or OR2 (N600, N586, N329);
nor NOR2 (N601, N578, N492);
not NOT1 (N602, N598);
or OR4 (N603, N602, N15, N405, N116);
nor NOR2 (N604, N541, N424);
nand NAND4 (N605, N596, N56, N472, N307);
or OR3 (N606, N585, N292, N297);
buf BUF1 (N607, N600);
buf BUF1 (N608, N594);
and AND4 (N609, N601, N72, N390, N587);
buf BUF1 (N610, N608);
buf BUF1 (N611, N605);
not NOT1 (N612, N609);
buf BUF1 (N613, N610);
xor XOR2 (N614, N597, N394);
and AND2 (N615, N599, N518);
xor XOR2 (N616, N606, N74);
and AND4 (N617, N613, N287, N178, N553);
nand NAND3 (N618, N607, N346, N74);
not NOT1 (N619, N604);
xor XOR2 (N620, N614, N125);
not NOT1 (N621, N603);
nand NAND4 (N622, N619, N409, N340, N376);
buf BUF1 (N623, N615);
nand NAND3 (N624, N590, N489, N590);
nor NOR3 (N625, N621, N616, N309);
not NOT1 (N626, N558);
nor NOR3 (N627, N617, N577, N483);
xor XOR2 (N628, N620, N464);
or OR4 (N629, N623, N34, N58, N147);
and AND2 (N630, N625, N139);
nand NAND3 (N631, N612, N316, N330);
and AND3 (N632, N622, N390, N166);
xor XOR2 (N633, N631, N104);
nand NAND2 (N634, N611, N53);
xor XOR2 (N635, N633, N577);
and AND4 (N636, N632, N89, N96, N395);
buf BUF1 (N637, N618);
and AND3 (N638, N637, N247, N395);
and AND4 (N639, N627, N386, N542, N480);
and AND3 (N640, N624, N164, N596);
not NOT1 (N641, N634);
xor XOR2 (N642, N630, N619);
or OR3 (N643, N626, N268, N519);
buf BUF1 (N644, N635);
nor NOR4 (N645, N644, N532, N538, N496);
nand NAND4 (N646, N628, N352, N484, N579);
or OR4 (N647, N641, N475, N556, N338);
nand NAND4 (N648, N643, N582, N575, N360);
nand NAND3 (N649, N639, N199, N237);
nand NAND3 (N650, N645, N67, N418);
buf BUF1 (N651, N647);
and AND3 (N652, N646, N405, N457);
xor XOR2 (N653, N636, N10);
or OR2 (N654, N648, N155);
and AND4 (N655, N651, N494, N3, N151);
not NOT1 (N656, N654);
nor NOR2 (N657, N650, N264);
buf BUF1 (N658, N642);
buf BUF1 (N659, N629);
nor NOR3 (N660, N649, N496, N493);
nor NOR3 (N661, N652, N235, N459);
nand NAND4 (N662, N661, N651, N192, N139);
nor NOR2 (N663, N655, N441);
or OR4 (N664, N662, N249, N377, N182);
xor XOR2 (N665, N640, N466);
nand NAND3 (N666, N660, N360, N513);
xor XOR2 (N667, N666, N288);
buf BUF1 (N668, N664);
and AND2 (N669, N657, N634);
and AND3 (N670, N659, N624, N178);
xor XOR2 (N671, N653, N556);
xor XOR2 (N672, N663, N640);
or OR3 (N673, N656, N390, N262);
buf BUF1 (N674, N669);
nand NAND2 (N675, N672, N100);
nand NAND4 (N676, N670, N439, N248, N588);
not NOT1 (N677, N638);
not NOT1 (N678, N676);
and AND4 (N679, N674, N192, N383, N633);
not NOT1 (N680, N667);
not NOT1 (N681, N673);
nand NAND4 (N682, N668, N225, N619, N49);
nand NAND3 (N683, N680, N101, N113);
xor XOR2 (N684, N665, N240);
nor NOR4 (N685, N675, N457, N8, N499);
nand NAND2 (N686, N678, N182);
not NOT1 (N687, N658);
buf BUF1 (N688, N681);
buf BUF1 (N689, N679);
nand NAND2 (N690, N685, N286);
nand NAND4 (N691, N677, N133, N613, N175);
not NOT1 (N692, N684);
and AND3 (N693, N690, N60, N608);
nand NAND4 (N694, N683, N362, N15, N109);
nand NAND3 (N695, N687, N450, N411);
buf BUF1 (N696, N693);
xor XOR2 (N697, N682, N271);
not NOT1 (N698, N692);
not NOT1 (N699, N686);
buf BUF1 (N700, N691);
not NOT1 (N701, N700);
nand NAND2 (N702, N689, N58);
buf BUF1 (N703, N699);
or OR4 (N704, N694, N214, N692, N452);
and AND2 (N705, N702, N195);
xor XOR2 (N706, N705, N513);
buf BUF1 (N707, N695);
nor NOR4 (N708, N696, N209, N557, N332);
xor XOR2 (N709, N703, N548);
and AND2 (N710, N708, N106);
buf BUF1 (N711, N697);
nor NOR4 (N712, N688, N696, N566, N105);
not NOT1 (N713, N704);
and AND3 (N714, N706, N350, N283);
nand NAND4 (N715, N711, N422, N151, N506);
nor NOR2 (N716, N707, N8);
nor NOR4 (N717, N716, N181, N596, N633);
and AND4 (N718, N709, N624, N144, N138);
not NOT1 (N719, N713);
nor NOR2 (N720, N701, N305);
or OR4 (N721, N714, N636, N551, N704);
nand NAND3 (N722, N719, N526, N506);
xor XOR2 (N723, N712, N313);
nor NOR2 (N724, N671, N319);
or OR4 (N725, N720, N447, N705, N717);
and AND2 (N726, N119, N134);
xor XOR2 (N727, N718, N332);
nor NOR3 (N728, N724, N109, N437);
not NOT1 (N729, N721);
xor XOR2 (N730, N723, N323);
xor XOR2 (N731, N726, N464);
nand NAND2 (N732, N698, N603);
and AND4 (N733, N725, N411, N649, N648);
not NOT1 (N734, N727);
not NOT1 (N735, N734);
not NOT1 (N736, N735);
and AND2 (N737, N736, N118);
not NOT1 (N738, N730);
nand NAND2 (N739, N731, N677);
buf BUF1 (N740, N733);
buf BUF1 (N741, N728);
xor XOR2 (N742, N741, N419);
xor XOR2 (N743, N737, N472);
and AND2 (N744, N739, N215);
buf BUF1 (N745, N740);
not NOT1 (N746, N745);
and AND4 (N747, N742, N522, N526, N405);
nand NAND4 (N748, N729, N291, N87, N151);
and AND3 (N749, N748, N608, N4);
and AND3 (N750, N722, N60, N633);
not NOT1 (N751, N746);
not NOT1 (N752, N715);
not NOT1 (N753, N732);
nor NOR2 (N754, N743, N663);
and AND4 (N755, N747, N388, N656, N392);
nor NOR4 (N756, N751, N260, N679, N446);
or OR3 (N757, N749, N469, N509);
nand NAND2 (N758, N756, N636);
xor XOR2 (N759, N710, N255);
and AND2 (N760, N759, N296);
xor XOR2 (N761, N757, N655);
xor XOR2 (N762, N744, N632);
xor XOR2 (N763, N750, N609);
nand NAND2 (N764, N738, N137);
or OR3 (N765, N761, N51, N86);
not NOT1 (N766, N760);
or OR4 (N767, N766, N556, N231, N252);
and AND3 (N768, N764, N702, N328);
not NOT1 (N769, N767);
or OR3 (N770, N755, N350, N334);
buf BUF1 (N771, N758);
nand NAND2 (N772, N753, N440);
buf BUF1 (N773, N763);
not NOT1 (N774, N765);
xor XOR2 (N775, N771, N306);
buf BUF1 (N776, N754);
buf BUF1 (N777, N768);
xor XOR2 (N778, N770, N595);
or OR2 (N779, N775, N172);
and AND4 (N780, N776, N491, N390, N257);
nand NAND3 (N781, N780, N157, N55);
nor NOR3 (N782, N762, N699, N203);
nand NAND3 (N783, N782, N61, N756);
and AND4 (N784, N752, N268, N330, N583);
buf BUF1 (N785, N769);
or OR3 (N786, N781, N780, N236);
nand NAND2 (N787, N773, N637);
buf BUF1 (N788, N772);
not NOT1 (N789, N785);
buf BUF1 (N790, N784);
nand NAND3 (N791, N783, N31, N668);
buf BUF1 (N792, N779);
xor XOR2 (N793, N790, N74);
buf BUF1 (N794, N793);
buf BUF1 (N795, N792);
or OR4 (N796, N789, N528, N590, N648);
or OR4 (N797, N796, N136, N535, N400);
not NOT1 (N798, N791);
and AND2 (N799, N777, N684);
not NOT1 (N800, N794);
nor NOR4 (N801, N800, N48, N370, N327);
buf BUF1 (N802, N774);
xor XOR2 (N803, N801, N699);
buf BUF1 (N804, N786);
nor NOR4 (N805, N778, N601, N68, N244);
buf BUF1 (N806, N803);
buf BUF1 (N807, N799);
and AND3 (N808, N795, N773, N680);
nand NAND2 (N809, N798, N636);
xor XOR2 (N810, N802, N682);
buf BUF1 (N811, N808);
nand NAND3 (N812, N787, N141, N744);
nor NOR3 (N813, N810, N188, N27);
or OR3 (N814, N805, N774, N528);
nand NAND4 (N815, N812, N36, N630, N209);
or OR3 (N816, N815, N175, N352);
nand NAND2 (N817, N809, N163);
nand NAND4 (N818, N817, N511, N332, N45);
and AND3 (N819, N804, N437, N154);
nand NAND2 (N820, N806, N669);
and AND3 (N821, N797, N99, N262);
or OR3 (N822, N821, N378, N274);
and AND4 (N823, N816, N522, N340, N192);
not NOT1 (N824, N814);
xor XOR2 (N825, N819, N121);
or OR2 (N826, N813, N197);
or OR3 (N827, N788, N304, N11);
nor NOR2 (N828, N823, N219);
nor NOR3 (N829, N822, N458, N33);
xor XOR2 (N830, N811, N636);
nor NOR4 (N831, N829, N234, N266, N659);
and AND3 (N832, N828, N336, N684);
not NOT1 (N833, N826);
nor NOR4 (N834, N825, N97, N570, N283);
nand NAND3 (N835, N833, N237, N230);
xor XOR2 (N836, N807, N254);
nor NOR4 (N837, N830, N489, N299, N560);
or OR3 (N838, N832, N445, N281);
xor XOR2 (N839, N834, N266);
and AND4 (N840, N838, N534, N741, N717);
nor NOR2 (N841, N827, N595);
and AND4 (N842, N836, N540, N107, N123);
buf BUF1 (N843, N837);
nand NAND3 (N844, N835, N791, N481);
buf BUF1 (N845, N839);
xor XOR2 (N846, N840, N559);
xor XOR2 (N847, N846, N588);
and AND3 (N848, N818, N534, N94);
or OR4 (N849, N844, N806, N50, N698);
nand NAND4 (N850, N824, N173, N355, N359);
nor NOR4 (N851, N848, N517, N609, N379);
not NOT1 (N852, N820);
or OR4 (N853, N850, N364, N665, N839);
nand NAND4 (N854, N853, N818, N257, N831);
buf BUF1 (N855, N523);
nand NAND3 (N856, N843, N331, N815);
buf BUF1 (N857, N849);
or OR3 (N858, N841, N632, N677);
not NOT1 (N859, N845);
nor NOR3 (N860, N847, N677, N488);
not NOT1 (N861, N855);
xor XOR2 (N862, N858, N339);
nor NOR2 (N863, N857, N129);
or OR2 (N864, N863, N765);
and AND4 (N865, N864, N82, N851, N822);
not NOT1 (N866, N40);
or OR2 (N867, N852, N498);
nor NOR3 (N868, N866, N583, N854);
not NOT1 (N869, N309);
nor NOR3 (N870, N868, N87, N87);
and AND3 (N871, N860, N126, N464);
not NOT1 (N872, N871);
xor XOR2 (N873, N856, N241);
buf BUF1 (N874, N867);
nor NOR2 (N875, N872, N367);
xor XOR2 (N876, N875, N655);
not NOT1 (N877, N874);
not NOT1 (N878, N876);
xor XOR2 (N879, N873, N29);
nor NOR2 (N880, N861, N303);
nand NAND2 (N881, N869, N778);
or OR4 (N882, N862, N478, N309, N336);
nand NAND3 (N883, N842, N313, N90);
and AND2 (N884, N879, N262);
or OR3 (N885, N882, N705, N530);
or OR4 (N886, N859, N192, N782, N260);
xor XOR2 (N887, N870, N358);
buf BUF1 (N888, N877);
nor NOR4 (N889, N886, N311, N32, N540);
or OR4 (N890, N881, N452, N766, N102);
buf BUF1 (N891, N883);
xor XOR2 (N892, N885, N300);
nor NOR2 (N893, N865, N425);
not NOT1 (N894, N880);
nor NOR2 (N895, N884, N241);
not NOT1 (N896, N890);
nand NAND4 (N897, N893, N293, N584, N49);
nand NAND4 (N898, N888, N336, N802, N748);
xor XOR2 (N899, N895, N82);
xor XOR2 (N900, N896, N90);
xor XOR2 (N901, N900, N37);
not NOT1 (N902, N898);
xor XOR2 (N903, N902, N123);
xor XOR2 (N904, N889, N141);
and AND3 (N905, N904, N824, N512);
nand NAND4 (N906, N897, N524, N576, N380);
not NOT1 (N907, N891);
and AND3 (N908, N907, N624, N732);
or OR3 (N909, N905, N147, N20);
not NOT1 (N910, N909);
nand NAND4 (N911, N908, N407, N435, N144);
xor XOR2 (N912, N906, N155);
buf BUF1 (N913, N912);
or OR3 (N914, N911, N650, N881);
or OR2 (N915, N887, N890);
xor XOR2 (N916, N914, N334);
xor XOR2 (N917, N903, N224);
not NOT1 (N918, N878);
buf BUF1 (N919, N913);
and AND3 (N920, N901, N272, N323);
nand NAND4 (N921, N917, N449, N84, N753);
not NOT1 (N922, N915);
xor XOR2 (N923, N918, N24);
or OR2 (N924, N921, N716);
not NOT1 (N925, N923);
and AND3 (N926, N899, N621, N52);
and AND3 (N927, N926, N839, N473);
xor XOR2 (N928, N920, N717);
or OR3 (N929, N922, N757, N572);
and AND2 (N930, N924, N312);
not NOT1 (N931, N892);
nor NOR3 (N932, N929, N506, N715);
nand NAND3 (N933, N910, N879, N754);
buf BUF1 (N934, N894);
nor NOR4 (N935, N927, N759, N509, N933);
buf BUF1 (N936, N766);
and AND4 (N937, N934, N400, N657, N211);
xor XOR2 (N938, N931, N929);
not NOT1 (N939, N916);
and AND2 (N940, N935, N309);
and AND3 (N941, N939, N390, N445);
nand NAND3 (N942, N936, N921, N788);
and AND3 (N943, N942, N49, N70);
not NOT1 (N944, N925);
nor NOR3 (N945, N944, N215, N128);
xor XOR2 (N946, N943, N520);
not NOT1 (N947, N940);
or OR4 (N948, N932, N197, N834, N676);
xor XOR2 (N949, N919, N108);
or OR4 (N950, N946, N158, N216, N780);
buf BUF1 (N951, N945);
nand NAND3 (N952, N950, N606, N514);
xor XOR2 (N953, N948, N950);
buf BUF1 (N954, N949);
nand NAND4 (N955, N928, N183, N610, N732);
and AND2 (N956, N941, N35);
and AND4 (N957, N956, N90, N265, N406);
or OR2 (N958, N937, N523);
xor XOR2 (N959, N955, N777);
buf BUF1 (N960, N947);
not NOT1 (N961, N954);
or OR3 (N962, N957, N70, N468);
or OR2 (N963, N961, N78);
xor XOR2 (N964, N960, N217);
buf BUF1 (N965, N952);
or OR3 (N966, N965, N522, N563);
xor XOR2 (N967, N930, N812);
nand NAND4 (N968, N962, N276, N777, N851);
xor XOR2 (N969, N963, N127);
not NOT1 (N970, N958);
nor NOR2 (N971, N951, N47);
and AND3 (N972, N970, N679, N721);
nand NAND4 (N973, N968, N482, N430, N597);
not NOT1 (N974, N938);
xor XOR2 (N975, N967, N54);
and AND2 (N976, N966, N568);
and AND2 (N977, N973, N678);
nor NOR2 (N978, N976, N282);
nand NAND3 (N979, N978, N523, N331);
or OR4 (N980, N971, N928, N926, N890);
or OR4 (N981, N980, N541, N26, N59);
not NOT1 (N982, N969);
or OR4 (N983, N974, N463, N743, N125);
buf BUF1 (N984, N953);
not NOT1 (N985, N983);
xor XOR2 (N986, N964, N967);
nand NAND4 (N987, N972, N268, N485, N155);
xor XOR2 (N988, N986, N823);
or OR3 (N989, N985, N157, N589);
buf BUF1 (N990, N979);
nor NOR3 (N991, N990, N473, N714);
nand NAND2 (N992, N959, N305);
and AND3 (N993, N992, N161, N528);
nand NAND2 (N994, N993, N202);
buf BUF1 (N995, N984);
not NOT1 (N996, N975);
xor XOR2 (N997, N996, N232);
not NOT1 (N998, N988);
not NOT1 (N999, N995);
buf BUF1 (N1000, N991);
not NOT1 (N1001, N989);
buf BUF1 (N1002, N981);
and AND3 (N1003, N1001, N647, N669);
xor XOR2 (N1004, N998, N946);
nand NAND3 (N1005, N999, N784, N532);
nand NAND4 (N1006, N1005, N325, N545, N282);
nand NAND2 (N1007, N1000, N355);
nand NAND2 (N1008, N1004, N739);
not NOT1 (N1009, N1007);
nor NOR4 (N1010, N987, N178, N914, N56);
xor XOR2 (N1011, N1006, N597);
xor XOR2 (N1012, N1003, N10);
buf BUF1 (N1013, N1002);
buf BUF1 (N1014, N997);
xor XOR2 (N1015, N994, N674);
and AND2 (N1016, N977, N373);
buf BUF1 (N1017, N1014);
buf BUF1 (N1018, N1011);
nor NOR3 (N1019, N1009, N41, N176);
nor NOR3 (N1020, N1015, N294, N240);
or OR4 (N1021, N1017, N207, N95, N456);
not NOT1 (N1022, N1016);
nor NOR4 (N1023, N1019, N696, N78, N204);
buf BUF1 (N1024, N1012);
buf BUF1 (N1025, N1022);
and AND3 (N1026, N1010, N19, N964);
or OR4 (N1027, N1020, N152, N787, N712);
nor NOR2 (N1028, N1008, N505);
not NOT1 (N1029, N1021);
xor XOR2 (N1030, N1023, N771);
nand NAND3 (N1031, N1024, N393, N807);
xor XOR2 (N1032, N1030, N555);
or OR4 (N1033, N1025, N277, N311, N888);
nor NOR4 (N1034, N1029, N117, N878, N649);
nand NAND3 (N1035, N1013, N486, N242);
nand NAND2 (N1036, N1034, N748);
nand NAND4 (N1037, N1033, N312, N473, N57);
and AND2 (N1038, N1036, N605);
buf BUF1 (N1039, N1026);
buf BUF1 (N1040, N1018);
and AND4 (N1041, N1028, N16, N479, N488);
and AND2 (N1042, N1035, N936);
nand NAND3 (N1043, N1040, N67, N914);
nand NAND4 (N1044, N1038, N774, N303, N491);
and AND2 (N1045, N1042, N724);
or OR2 (N1046, N1031, N151);
nor NOR4 (N1047, N1037, N858, N688, N407);
xor XOR2 (N1048, N1041, N791);
nand NAND3 (N1049, N1046, N352, N906);
or OR2 (N1050, N1027, N6);
buf BUF1 (N1051, N1045);
buf BUF1 (N1052, N1051);
nand NAND3 (N1053, N1044, N31, N864);
or OR4 (N1054, N1052, N6, N749, N499);
nor NOR2 (N1055, N1039, N27);
nor NOR4 (N1056, N1047, N1017, N50, N364);
not NOT1 (N1057, N982);
nor NOR3 (N1058, N1043, N264, N483);
xor XOR2 (N1059, N1053, N740);
not NOT1 (N1060, N1055);
or OR2 (N1061, N1054, N371);
or OR3 (N1062, N1032, N64, N1048);
not NOT1 (N1063, N341);
xor XOR2 (N1064, N1057, N75);
nor NOR2 (N1065, N1061, N628);
not NOT1 (N1066, N1064);
not NOT1 (N1067, N1062);
nand NAND2 (N1068, N1059, N495);
not NOT1 (N1069, N1067);
nand NAND2 (N1070, N1056, N835);
and AND3 (N1071, N1060, N889, N557);
nand NAND3 (N1072, N1066, N210, N468);
not NOT1 (N1073, N1049);
and AND3 (N1074, N1071, N634, N866);
xor XOR2 (N1075, N1058, N226);
not NOT1 (N1076, N1074);
nand NAND2 (N1077, N1065, N955);
and AND4 (N1078, N1077, N501, N374, N678);
nand NAND4 (N1079, N1050, N105, N824, N390);
not NOT1 (N1080, N1076);
or OR4 (N1081, N1080, N403, N893, N241);
xor XOR2 (N1082, N1063, N1021);
not NOT1 (N1083, N1072);
or OR3 (N1084, N1075, N1020, N750);
not NOT1 (N1085, N1079);
nor NOR3 (N1086, N1068, N979, N729);
not NOT1 (N1087, N1081);
nand NAND3 (N1088, N1073, N979, N532);
not NOT1 (N1089, N1070);
buf BUF1 (N1090, N1088);
buf BUF1 (N1091, N1087);
xor XOR2 (N1092, N1091, N1020);
nor NOR2 (N1093, N1082, N904);
buf BUF1 (N1094, N1086);
nand NAND4 (N1095, N1090, N406, N546, N334);
nand NAND2 (N1096, N1089, N367);
xor XOR2 (N1097, N1085, N530);
nand NAND2 (N1098, N1092, N655);
buf BUF1 (N1099, N1069);
xor XOR2 (N1100, N1097, N341);
not NOT1 (N1101, N1094);
and AND3 (N1102, N1095, N172, N318);
not NOT1 (N1103, N1099);
xor XOR2 (N1104, N1096, N29);
buf BUF1 (N1105, N1093);
xor XOR2 (N1106, N1105, N408);
xor XOR2 (N1107, N1083, N168);
xor XOR2 (N1108, N1098, N1054);
xor XOR2 (N1109, N1101, N82);
nor NOR2 (N1110, N1108, N889);
nand NAND3 (N1111, N1109, N1034, N666);
buf BUF1 (N1112, N1078);
or OR2 (N1113, N1106, N46);
or OR3 (N1114, N1084, N785, N897);
nor NOR2 (N1115, N1114, N29);
nor NOR2 (N1116, N1100, N967);
not NOT1 (N1117, N1103);
nor NOR4 (N1118, N1111, N581, N543, N808);
xor XOR2 (N1119, N1102, N358);
or OR4 (N1120, N1115, N131, N861, N32);
buf BUF1 (N1121, N1116);
nor NOR4 (N1122, N1121, N650, N1038, N875);
xor XOR2 (N1123, N1119, N338);
or OR3 (N1124, N1112, N208, N568);
or OR3 (N1125, N1124, N989, N464);
nand NAND3 (N1126, N1122, N712, N454);
buf BUF1 (N1127, N1113);
buf BUF1 (N1128, N1123);
nand NAND3 (N1129, N1128, N762, N299);
xor XOR2 (N1130, N1120, N943);
nor NOR3 (N1131, N1125, N675, N737);
not NOT1 (N1132, N1129);
nand NAND3 (N1133, N1107, N662, N272);
or OR4 (N1134, N1127, N508, N351, N191);
buf BUF1 (N1135, N1130);
nor NOR3 (N1136, N1133, N22, N457);
buf BUF1 (N1137, N1118);
nand NAND2 (N1138, N1104, N34);
not NOT1 (N1139, N1134);
nand NAND2 (N1140, N1131, N310);
not NOT1 (N1141, N1136);
not NOT1 (N1142, N1110);
not NOT1 (N1143, N1141);
nor NOR2 (N1144, N1135, N800);
nor NOR3 (N1145, N1140, N684, N846);
not NOT1 (N1146, N1145);
nor NOR4 (N1147, N1139, N721, N115, N315);
nand NAND4 (N1148, N1137, N954, N387, N1104);
buf BUF1 (N1149, N1146);
and AND4 (N1150, N1138, N339, N588, N104);
xor XOR2 (N1151, N1132, N383);
xor XOR2 (N1152, N1150, N716);
buf BUF1 (N1153, N1142);
nand NAND3 (N1154, N1153, N463, N407);
nand NAND4 (N1155, N1151, N1114, N756, N962);
and AND2 (N1156, N1149, N857);
nand NAND2 (N1157, N1155, N379);
xor XOR2 (N1158, N1147, N641);
nor NOR3 (N1159, N1126, N663, N1080);
nor NOR3 (N1160, N1154, N639, N127);
nand NAND4 (N1161, N1152, N247, N1152, N640);
nand NAND3 (N1162, N1158, N231, N477);
nand NAND3 (N1163, N1156, N251, N641);
and AND2 (N1164, N1143, N736);
nand NAND3 (N1165, N1161, N613, N253);
buf BUF1 (N1166, N1148);
not NOT1 (N1167, N1163);
buf BUF1 (N1168, N1160);
or OR4 (N1169, N1162, N986, N748, N585);
not NOT1 (N1170, N1168);
nor NOR3 (N1171, N1165, N612, N1160);
nand NAND4 (N1172, N1171, N804, N622, N804);
nand NAND2 (N1173, N1117, N47);
nand NAND3 (N1174, N1172, N29, N192);
xor XOR2 (N1175, N1169, N172);
nand NAND3 (N1176, N1166, N212, N230);
not NOT1 (N1177, N1144);
not NOT1 (N1178, N1177);
or OR3 (N1179, N1175, N828, N324);
or OR2 (N1180, N1167, N526);
xor XOR2 (N1181, N1157, N1135);
not NOT1 (N1182, N1176);
xor XOR2 (N1183, N1178, N421);
not NOT1 (N1184, N1170);
not NOT1 (N1185, N1182);
nor NOR3 (N1186, N1174, N1004, N540);
or OR4 (N1187, N1180, N1091, N475, N374);
or OR2 (N1188, N1164, N984);
nor NOR3 (N1189, N1173, N527, N172);
nand NAND2 (N1190, N1186, N243);
not NOT1 (N1191, N1184);
xor XOR2 (N1192, N1185, N198);
or OR2 (N1193, N1192, N449);
nand NAND3 (N1194, N1191, N798, N121);
and AND4 (N1195, N1188, N8, N936, N581);
and AND2 (N1196, N1190, N582);
or OR2 (N1197, N1189, N188);
nand NAND3 (N1198, N1194, N1092, N447);
not NOT1 (N1199, N1179);
buf BUF1 (N1200, N1193);
nor NOR4 (N1201, N1196, N1078, N677, N409);
nor NOR2 (N1202, N1183, N837);
buf BUF1 (N1203, N1187);
and AND4 (N1204, N1200, N665, N302, N612);
or OR4 (N1205, N1204, N933, N129, N42);
buf BUF1 (N1206, N1159);
or OR4 (N1207, N1181, N807, N517, N842);
not NOT1 (N1208, N1195);
buf BUF1 (N1209, N1198);
nand NAND4 (N1210, N1203, N161, N93, N555);
nor NOR4 (N1211, N1206, N237, N395, N919);
nand NAND3 (N1212, N1199, N643, N648);
nand NAND3 (N1213, N1211, N1203, N843);
or OR2 (N1214, N1209, N1183);
or OR2 (N1215, N1214, N1147);
xor XOR2 (N1216, N1202, N256);
nand NAND2 (N1217, N1208, N90);
xor XOR2 (N1218, N1212, N1186);
not NOT1 (N1219, N1218);
and AND2 (N1220, N1219, N739);
nor NOR3 (N1221, N1213, N1080, N918);
not NOT1 (N1222, N1217);
or OR4 (N1223, N1210, N187, N461, N135);
not NOT1 (N1224, N1205);
and AND4 (N1225, N1215, N930, N1205, N686);
buf BUF1 (N1226, N1201);
buf BUF1 (N1227, N1224);
and AND3 (N1228, N1225, N1086, N610);
and AND3 (N1229, N1221, N861, N771);
nor NOR2 (N1230, N1227, N669);
buf BUF1 (N1231, N1226);
or OR2 (N1232, N1229, N728);
not NOT1 (N1233, N1207);
or OR2 (N1234, N1231, N1025);
xor XOR2 (N1235, N1234, N958);
nand NAND3 (N1236, N1233, N959, N1089);
and AND3 (N1237, N1220, N389, N347);
buf BUF1 (N1238, N1197);
nand NAND2 (N1239, N1228, N1018);
or OR3 (N1240, N1237, N588, N165);
or OR2 (N1241, N1240, N158);
buf BUF1 (N1242, N1223);
xor XOR2 (N1243, N1239, N1194);
nand NAND2 (N1244, N1243, N712);
xor XOR2 (N1245, N1242, N883);
nor NOR3 (N1246, N1235, N266, N14);
xor XOR2 (N1247, N1245, N312);
or OR3 (N1248, N1244, N167, N1095);
not NOT1 (N1249, N1241);
nor NOR4 (N1250, N1222, N308, N421, N1138);
and AND3 (N1251, N1232, N1156, N1137);
buf BUF1 (N1252, N1248);
nand NAND2 (N1253, N1249, N1224);
not NOT1 (N1254, N1238);
buf BUF1 (N1255, N1250);
not NOT1 (N1256, N1253);
or OR2 (N1257, N1252, N839);
not NOT1 (N1258, N1247);
nand NAND4 (N1259, N1256, N1195, N217, N374);
nor NOR2 (N1260, N1259, N113);
nand NAND4 (N1261, N1257, N877, N969, N232);
nand NAND2 (N1262, N1246, N102);
nand NAND4 (N1263, N1216, N356, N551, N829);
xor XOR2 (N1264, N1261, N428);
nor NOR4 (N1265, N1230, N155, N1190, N1141);
or OR3 (N1266, N1260, N641, N342);
or OR4 (N1267, N1251, N957, N206, N326);
or OR2 (N1268, N1266, N29);
not NOT1 (N1269, N1267);
xor XOR2 (N1270, N1236, N44);
and AND3 (N1271, N1262, N212, N28);
and AND4 (N1272, N1268, N382, N706, N1239);
or OR3 (N1273, N1272, N695, N137);
nor NOR3 (N1274, N1255, N762, N16);
and AND2 (N1275, N1274, N363);
or OR3 (N1276, N1273, N867, N532);
nand NAND2 (N1277, N1271, N728);
xor XOR2 (N1278, N1265, N1277);
or OR2 (N1279, N323, N790);
and AND2 (N1280, N1279, N1267);
buf BUF1 (N1281, N1276);
and AND3 (N1282, N1258, N1081, N829);
buf BUF1 (N1283, N1281);
nor NOR3 (N1284, N1275, N688, N1083);
nor NOR2 (N1285, N1283, N812);
nor NOR2 (N1286, N1282, N514);
buf BUF1 (N1287, N1280);
not NOT1 (N1288, N1254);
nand NAND4 (N1289, N1270, N1087, N1032, N112);
not NOT1 (N1290, N1287);
and AND4 (N1291, N1269, N567, N1064, N711);
buf BUF1 (N1292, N1278);
and AND3 (N1293, N1264, N792, N702);
nor NOR2 (N1294, N1263, N861);
xor XOR2 (N1295, N1291, N1263);
or OR2 (N1296, N1295, N825);
or OR3 (N1297, N1292, N238, N644);
not NOT1 (N1298, N1286);
buf BUF1 (N1299, N1284);
nor NOR2 (N1300, N1290, N372);
xor XOR2 (N1301, N1285, N453);
and AND3 (N1302, N1296, N310, N800);
or OR4 (N1303, N1298, N379, N39, N471);
nand NAND4 (N1304, N1303, N304, N1094, N467);
nand NAND2 (N1305, N1289, N438);
not NOT1 (N1306, N1300);
nand NAND4 (N1307, N1299, N139, N954, N1278);
nand NAND2 (N1308, N1288, N738);
nand NAND3 (N1309, N1307, N1276, N932);
buf BUF1 (N1310, N1304);
nand NAND2 (N1311, N1310, N949);
nand NAND4 (N1312, N1302, N418, N6, N467);
or OR2 (N1313, N1301, N471);
nor NOR2 (N1314, N1294, N2);
and AND2 (N1315, N1293, N838);
nand NAND2 (N1316, N1305, N644);
xor XOR2 (N1317, N1316, N326);
or OR4 (N1318, N1317, N1160, N85, N518);
nand NAND4 (N1319, N1315, N207, N1248, N54);
nor NOR3 (N1320, N1314, N724, N949);
buf BUF1 (N1321, N1319);
not NOT1 (N1322, N1297);
nor NOR2 (N1323, N1306, N335);
or OR3 (N1324, N1318, N808, N1115);
nand NAND4 (N1325, N1322, N770, N325, N1076);
nand NAND4 (N1326, N1311, N921, N933, N323);
buf BUF1 (N1327, N1313);
nor NOR4 (N1328, N1323, N128, N100, N516);
and AND4 (N1329, N1320, N1295, N339, N1081);
not NOT1 (N1330, N1321);
buf BUF1 (N1331, N1308);
or OR2 (N1332, N1328, N1255);
xor XOR2 (N1333, N1330, N220);
buf BUF1 (N1334, N1325);
nand NAND3 (N1335, N1332, N20, N549);
xor XOR2 (N1336, N1331, N691);
nand NAND4 (N1337, N1324, N431, N420, N4);
not NOT1 (N1338, N1337);
not NOT1 (N1339, N1326);
nand NAND3 (N1340, N1312, N1224, N1070);
nand NAND4 (N1341, N1335, N398, N723, N103);
buf BUF1 (N1342, N1334);
and AND4 (N1343, N1339, N737, N79, N379);
nand NAND4 (N1344, N1309, N991, N894, N774);
buf BUF1 (N1345, N1333);
and AND4 (N1346, N1327, N217, N882, N994);
nor NOR4 (N1347, N1340, N832, N828, N525);
or OR2 (N1348, N1344, N806);
or OR3 (N1349, N1347, N278, N622);
xor XOR2 (N1350, N1349, N1046);
buf BUF1 (N1351, N1343);
or OR3 (N1352, N1336, N130, N1069);
nand NAND2 (N1353, N1329, N21);
and AND3 (N1354, N1351, N433, N825);
or OR3 (N1355, N1342, N416, N368);
nand NAND4 (N1356, N1354, N1293, N776, N853);
not NOT1 (N1357, N1345);
buf BUF1 (N1358, N1338);
or OR3 (N1359, N1357, N68, N161);
or OR2 (N1360, N1350, N1076);
xor XOR2 (N1361, N1359, N1127);
nand NAND2 (N1362, N1346, N376);
xor XOR2 (N1363, N1355, N646);
or OR3 (N1364, N1353, N215, N946);
and AND3 (N1365, N1348, N94, N347);
nand NAND2 (N1366, N1352, N624);
nand NAND2 (N1367, N1365, N731);
buf BUF1 (N1368, N1363);
buf BUF1 (N1369, N1362);
xor XOR2 (N1370, N1356, N387);
buf BUF1 (N1371, N1368);
nor NOR3 (N1372, N1366, N687, N269);
buf BUF1 (N1373, N1370);
and AND2 (N1374, N1364, N111);
not NOT1 (N1375, N1358);
or OR4 (N1376, N1373, N196, N473, N362);
or OR2 (N1377, N1376, N367);
not NOT1 (N1378, N1371);
not NOT1 (N1379, N1361);
buf BUF1 (N1380, N1367);
or OR4 (N1381, N1372, N832, N104, N965);
or OR3 (N1382, N1360, N415, N1057);
nand NAND2 (N1383, N1379, N953);
not NOT1 (N1384, N1383);
not NOT1 (N1385, N1382);
not NOT1 (N1386, N1375);
or OR4 (N1387, N1381, N503, N654, N1129);
xor XOR2 (N1388, N1384, N193);
nor NOR3 (N1389, N1377, N159, N996);
not NOT1 (N1390, N1380);
buf BUF1 (N1391, N1390);
and AND3 (N1392, N1389, N1197, N947);
nor NOR4 (N1393, N1386, N541, N539, N1262);
and AND3 (N1394, N1385, N1216, N160);
and AND3 (N1395, N1393, N418, N731);
nand NAND2 (N1396, N1388, N1015);
and AND4 (N1397, N1396, N1312, N863, N543);
xor XOR2 (N1398, N1374, N780);
nor NOR3 (N1399, N1395, N1046, N1214);
nor NOR2 (N1400, N1397, N215);
not NOT1 (N1401, N1387);
xor XOR2 (N1402, N1378, N6);
buf BUF1 (N1403, N1401);
not NOT1 (N1404, N1399);
or OR4 (N1405, N1403, N1322, N1086, N1394);
and AND4 (N1406, N163, N1395, N504, N1143);
or OR2 (N1407, N1406, N248);
not NOT1 (N1408, N1398);
or OR3 (N1409, N1402, N375, N1265);
and AND2 (N1410, N1409, N521);
nand NAND4 (N1411, N1410, N1222, N1259, N1155);
not NOT1 (N1412, N1392);
buf BUF1 (N1413, N1412);
nand NAND3 (N1414, N1341, N1109, N1253);
buf BUF1 (N1415, N1413);
buf BUF1 (N1416, N1404);
not NOT1 (N1417, N1416);
xor XOR2 (N1418, N1414, N429);
nand NAND2 (N1419, N1408, N336);
or OR3 (N1420, N1405, N1352, N631);
nor NOR4 (N1421, N1411, N414, N491, N254);
xor XOR2 (N1422, N1407, N454);
buf BUF1 (N1423, N1418);
not NOT1 (N1424, N1400);
nor NOR2 (N1425, N1415, N895);
not NOT1 (N1426, N1425);
nor NOR2 (N1427, N1424, N924);
or OR2 (N1428, N1426, N472);
xor XOR2 (N1429, N1369, N61);
not NOT1 (N1430, N1427);
and AND4 (N1431, N1421, N953, N278, N169);
and AND2 (N1432, N1391, N276);
and AND3 (N1433, N1422, N267, N683);
and AND2 (N1434, N1430, N274);
or OR2 (N1435, N1420, N1196);
and AND4 (N1436, N1417, N684, N68, N164);
and AND3 (N1437, N1428, N1135, N375);
and AND3 (N1438, N1436, N674, N1216);
nand NAND3 (N1439, N1437, N156, N1155);
nor NOR3 (N1440, N1432, N1397, N1272);
nor NOR3 (N1441, N1435, N1095, N111);
buf BUF1 (N1442, N1423);
nand NAND3 (N1443, N1441, N888, N136);
and AND3 (N1444, N1439, N191, N532);
not NOT1 (N1445, N1429);
nand NAND3 (N1446, N1419, N415, N1248);
xor XOR2 (N1447, N1433, N390);
and AND4 (N1448, N1438, N134, N1172, N1380);
and AND3 (N1449, N1431, N510, N525);
nor NOR4 (N1450, N1446, N499, N885, N810);
and AND4 (N1451, N1443, N1228, N384, N1069);
and AND3 (N1452, N1442, N1159, N181);
or OR4 (N1453, N1444, N1287, N1331, N878);
or OR3 (N1454, N1448, N527, N965);
or OR4 (N1455, N1452, N9, N624, N602);
or OR3 (N1456, N1450, N21, N828);
and AND2 (N1457, N1445, N301);
xor XOR2 (N1458, N1447, N356);
xor XOR2 (N1459, N1451, N1434);
and AND4 (N1460, N629, N652, N1075, N849);
and AND2 (N1461, N1449, N409);
or OR2 (N1462, N1454, N1428);
not NOT1 (N1463, N1458);
and AND4 (N1464, N1453, N1422, N630, N892);
nor NOR2 (N1465, N1459, N769);
and AND2 (N1466, N1462, N837);
buf BUF1 (N1467, N1460);
xor XOR2 (N1468, N1464, N450);
nand NAND4 (N1469, N1457, N1387, N1303, N644);
or OR3 (N1470, N1463, N502, N538);
nor NOR4 (N1471, N1455, N1108, N661, N147);
nor NOR4 (N1472, N1465, N364, N100, N212);
nand NAND2 (N1473, N1466, N929);
and AND2 (N1474, N1472, N433);
xor XOR2 (N1475, N1469, N288);
nor NOR3 (N1476, N1467, N1040, N300);
not NOT1 (N1477, N1470);
not NOT1 (N1478, N1477);
nand NAND2 (N1479, N1475, N857);
and AND3 (N1480, N1440, N132, N293);
or OR3 (N1481, N1478, N482, N785);
buf BUF1 (N1482, N1481);
nor NOR3 (N1483, N1461, N1210, N1183);
nor NOR3 (N1484, N1480, N406, N409);
or OR3 (N1485, N1471, N738, N515);
or OR3 (N1486, N1456, N1138, N330);
and AND3 (N1487, N1474, N987, N587);
or OR4 (N1488, N1484, N974, N1352, N1361);
or OR3 (N1489, N1483, N358, N1065);
xor XOR2 (N1490, N1476, N1234);
or OR3 (N1491, N1490, N460, N145);
nor NOR3 (N1492, N1482, N877, N770);
xor XOR2 (N1493, N1491, N1434);
or OR3 (N1494, N1468, N1376, N784);
and AND4 (N1495, N1479, N1170, N985, N47);
and AND2 (N1496, N1487, N534);
not NOT1 (N1497, N1489);
or OR4 (N1498, N1494, N187, N601, N561);
and AND2 (N1499, N1495, N1247);
not NOT1 (N1500, N1493);
nand NAND4 (N1501, N1498, N870, N1073, N1063);
nor NOR4 (N1502, N1501, N1308, N1404, N755);
xor XOR2 (N1503, N1499, N610);
nand NAND4 (N1504, N1497, N1253, N1352, N558);
buf BUF1 (N1505, N1503);
xor XOR2 (N1506, N1492, N1433);
or OR2 (N1507, N1506, N1256);
and AND3 (N1508, N1486, N305, N1480);
buf BUF1 (N1509, N1505);
buf BUF1 (N1510, N1488);
nand NAND3 (N1511, N1500, N459, N370);
nor NOR2 (N1512, N1510, N938);
buf BUF1 (N1513, N1512);
or OR3 (N1514, N1485, N461, N212);
or OR4 (N1515, N1509, N1299, N787, N1117);
nand NAND3 (N1516, N1514, N904, N574);
xor XOR2 (N1517, N1496, N203);
or OR2 (N1518, N1515, N1001);
not NOT1 (N1519, N1513);
not NOT1 (N1520, N1473);
xor XOR2 (N1521, N1516, N87);
nand NAND2 (N1522, N1521, N1178);
nor NOR2 (N1523, N1518, N1277);
not NOT1 (N1524, N1507);
xor XOR2 (N1525, N1511, N827);
xor XOR2 (N1526, N1519, N398);
not NOT1 (N1527, N1522);
and AND2 (N1528, N1502, N799);
nand NAND4 (N1529, N1526, N1124, N1471, N639);
buf BUF1 (N1530, N1529);
not NOT1 (N1531, N1520);
not NOT1 (N1532, N1524);
xor XOR2 (N1533, N1531, N544);
and AND3 (N1534, N1533, N93, N1302);
or OR4 (N1535, N1523, N414, N1261, N835);
not NOT1 (N1536, N1508);
buf BUF1 (N1537, N1517);
and AND2 (N1538, N1530, N789);
xor XOR2 (N1539, N1535, N582);
not NOT1 (N1540, N1537);
buf BUF1 (N1541, N1532);
buf BUF1 (N1542, N1538);
not NOT1 (N1543, N1534);
nor NOR3 (N1544, N1525, N320, N768);
nor NOR2 (N1545, N1528, N883);
not NOT1 (N1546, N1542);
nor NOR2 (N1547, N1540, N198);
and AND3 (N1548, N1545, N84, N309);
or OR2 (N1549, N1543, N1491);
buf BUF1 (N1550, N1527);
nor NOR3 (N1551, N1547, N301, N60);
nand NAND2 (N1552, N1546, N534);
nand NAND2 (N1553, N1551, N292);
not NOT1 (N1554, N1550);
and AND2 (N1555, N1549, N221);
or OR4 (N1556, N1553, N994, N456, N918);
not NOT1 (N1557, N1539);
xor XOR2 (N1558, N1552, N1179);
nor NOR4 (N1559, N1555, N1286, N490, N517);
nand NAND4 (N1560, N1541, N489, N637, N419);
not NOT1 (N1561, N1559);
and AND3 (N1562, N1504, N890, N546);
or OR4 (N1563, N1558, N992, N920, N252);
or OR4 (N1564, N1544, N996, N552, N252);
nor NOR4 (N1565, N1548, N299, N491, N1116);
xor XOR2 (N1566, N1556, N1207);
not NOT1 (N1567, N1560);
nand NAND2 (N1568, N1564, N604);
or OR4 (N1569, N1557, N411, N640, N227);
buf BUF1 (N1570, N1563);
nand NAND3 (N1571, N1554, N223, N1271);
not NOT1 (N1572, N1561);
or OR2 (N1573, N1565, N133);
and AND3 (N1574, N1573, N895, N1206);
nor NOR3 (N1575, N1567, N703, N256);
not NOT1 (N1576, N1566);
xor XOR2 (N1577, N1562, N488);
nand NAND3 (N1578, N1569, N970, N1363);
and AND3 (N1579, N1571, N1334, N988);
xor XOR2 (N1580, N1578, N1144);
buf BUF1 (N1581, N1579);
xor XOR2 (N1582, N1570, N983);
nand NAND4 (N1583, N1582, N1259, N1283, N742);
and AND3 (N1584, N1583, N1443, N1195);
not NOT1 (N1585, N1584);
nor NOR3 (N1586, N1572, N155, N645);
buf BUF1 (N1587, N1577);
or OR3 (N1588, N1568, N203, N609);
buf BUF1 (N1589, N1581);
xor XOR2 (N1590, N1576, N1515);
or OR3 (N1591, N1580, N759, N478);
buf BUF1 (N1592, N1586);
or OR4 (N1593, N1575, N1469, N113, N1449);
xor XOR2 (N1594, N1574, N932);
not NOT1 (N1595, N1593);
buf BUF1 (N1596, N1595);
not NOT1 (N1597, N1588);
not NOT1 (N1598, N1591);
buf BUF1 (N1599, N1585);
xor XOR2 (N1600, N1594, N123);
and AND4 (N1601, N1592, N7, N1294, N704);
nand NAND4 (N1602, N1587, N192, N1052, N1489);
nand NAND4 (N1603, N1598, N329, N118, N200);
nand NAND2 (N1604, N1596, N1124);
nor NOR3 (N1605, N1601, N314, N975);
not NOT1 (N1606, N1603);
buf BUF1 (N1607, N1606);
and AND4 (N1608, N1604, N246, N1187, N1040);
not NOT1 (N1609, N1602);
not NOT1 (N1610, N1605);
xor XOR2 (N1611, N1610, N1083);
or OR4 (N1612, N1607, N1064, N823, N470);
buf BUF1 (N1613, N1608);
xor XOR2 (N1614, N1609, N1486);
buf BUF1 (N1615, N1600);
xor XOR2 (N1616, N1614, N1319);
not NOT1 (N1617, N1536);
and AND3 (N1618, N1616, N1031, N43);
and AND4 (N1619, N1617, N1174, N430, N952);
not NOT1 (N1620, N1611);
and AND2 (N1621, N1597, N580);
nor NOR3 (N1622, N1618, N1505, N935);
buf BUF1 (N1623, N1612);
nand NAND2 (N1624, N1619, N1104);
nor NOR4 (N1625, N1590, N1432, N728, N1397);
not NOT1 (N1626, N1589);
xor XOR2 (N1627, N1620, N1518);
nand NAND2 (N1628, N1626, N1505);
nand NAND4 (N1629, N1624, N863, N266, N1137);
or OR3 (N1630, N1622, N1043, N1214);
or OR3 (N1631, N1627, N1061, N971);
or OR3 (N1632, N1599, N83, N925);
nor NOR4 (N1633, N1632, N169, N1057, N617);
xor XOR2 (N1634, N1615, N1475);
nor NOR2 (N1635, N1628, N483);
xor XOR2 (N1636, N1629, N1326);
buf BUF1 (N1637, N1631);
not NOT1 (N1638, N1635);
xor XOR2 (N1639, N1630, N856);
and AND4 (N1640, N1625, N749, N1081, N718);
nand NAND4 (N1641, N1634, N1640, N1116, N76);
not NOT1 (N1642, N1481);
and AND3 (N1643, N1636, N106, N680);
not NOT1 (N1644, N1621);
not NOT1 (N1645, N1613);
buf BUF1 (N1646, N1643);
nand NAND3 (N1647, N1642, N1164, N128);
and AND2 (N1648, N1638, N1519);
not NOT1 (N1649, N1647);
xor XOR2 (N1650, N1623, N1631);
and AND2 (N1651, N1646, N874);
buf BUF1 (N1652, N1650);
or OR4 (N1653, N1645, N166, N1008, N1445);
xor XOR2 (N1654, N1641, N564);
buf BUF1 (N1655, N1651);
buf BUF1 (N1656, N1633);
nand NAND2 (N1657, N1648, N952);
not NOT1 (N1658, N1652);
nor NOR4 (N1659, N1657, N601, N1010, N541);
nand NAND2 (N1660, N1655, N792);
or OR3 (N1661, N1644, N45, N1288);
and AND4 (N1662, N1656, N1442, N1056, N1151);
nor NOR3 (N1663, N1653, N319, N1247);
buf BUF1 (N1664, N1637);
not NOT1 (N1665, N1663);
or OR2 (N1666, N1649, N1144);
xor XOR2 (N1667, N1660, N707);
nor NOR2 (N1668, N1666, N1562);
and AND4 (N1669, N1662, N805, N852, N695);
nor NOR3 (N1670, N1658, N1298, N1565);
xor XOR2 (N1671, N1661, N374);
buf BUF1 (N1672, N1664);
or OR4 (N1673, N1669, N1151, N803, N827);
xor XOR2 (N1674, N1673, N920);
and AND2 (N1675, N1672, N535);
nor NOR2 (N1676, N1674, N1069);
not NOT1 (N1677, N1654);
buf BUF1 (N1678, N1639);
not NOT1 (N1679, N1671);
or OR4 (N1680, N1667, N1611, N1401, N820);
and AND4 (N1681, N1670, N839, N985, N608);
buf BUF1 (N1682, N1680);
and AND4 (N1683, N1681, N1626, N1049, N1302);
xor XOR2 (N1684, N1668, N278);
or OR3 (N1685, N1683, N450, N846);
nand NAND4 (N1686, N1675, N761, N1089, N980);
nor NOR4 (N1687, N1682, N1583, N1527, N1518);
not NOT1 (N1688, N1687);
or OR4 (N1689, N1685, N545, N101, N1063);
or OR4 (N1690, N1688, N1231, N1113, N1010);
xor XOR2 (N1691, N1659, N1450);
buf BUF1 (N1692, N1678);
or OR4 (N1693, N1684, N274, N651, N500);
not NOT1 (N1694, N1691);
buf BUF1 (N1695, N1690);
nor NOR3 (N1696, N1686, N450, N293);
and AND3 (N1697, N1665, N1660, N1203);
xor XOR2 (N1698, N1694, N296);
and AND3 (N1699, N1677, N419, N467);
nor NOR2 (N1700, N1689, N201);
or OR3 (N1701, N1679, N108, N1381);
or OR4 (N1702, N1700, N842, N1496, N496);
nor NOR2 (N1703, N1698, N23);
not NOT1 (N1704, N1703);
nand NAND3 (N1705, N1695, N1617, N773);
not NOT1 (N1706, N1705);
nor NOR2 (N1707, N1701, N1172);
not NOT1 (N1708, N1676);
and AND4 (N1709, N1696, N481, N1225, N1473);
buf BUF1 (N1710, N1709);
and AND3 (N1711, N1710, N923, N364);
buf BUF1 (N1712, N1692);
not NOT1 (N1713, N1697);
nor NOR3 (N1714, N1706, N509, N1494);
xor XOR2 (N1715, N1714, N1097);
xor XOR2 (N1716, N1707, N493);
xor XOR2 (N1717, N1715, N75);
buf BUF1 (N1718, N1711);
and AND2 (N1719, N1699, N1130);
nand NAND4 (N1720, N1717, N1664, N1719, N526);
and AND4 (N1721, N957, N704, N1199, N643);
not NOT1 (N1722, N1702);
and AND3 (N1723, N1713, N225, N362);
or OR4 (N1724, N1716, N1318, N523, N309);
nand NAND3 (N1725, N1693, N338, N490);
nor NOR2 (N1726, N1722, N1017);
nand NAND2 (N1727, N1723, N560);
and AND2 (N1728, N1708, N665);
or OR2 (N1729, N1704, N15);
buf BUF1 (N1730, N1718);
or OR4 (N1731, N1730, N1479, N533, N1596);
and AND4 (N1732, N1725, N544, N259, N1192);
and AND3 (N1733, N1732, N223, N326);
nand NAND2 (N1734, N1721, N1491);
nand NAND3 (N1735, N1726, N661, N559);
buf BUF1 (N1736, N1728);
xor XOR2 (N1737, N1720, N1652);
xor XOR2 (N1738, N1712, N643);
or OR3 (N1739, N1724, N1442, N259);
xor XOR2 (N1740, N1736, N965);
or OR3 (N1741, N1737, N574, N1305);
buf BUF1 (N1742, N1731);
buf BUF1 (N1743, N1734);
or OR4 (N1744, N1742, N1248, N40, N104);
buf BUF1 (N1745, N1741);
not NOT1 (N1746, N1739);
nor NOR3 (N1747, N1733, N1625, N1031);
or OR2 (N1748, N1743, N56);
nand NAND2 (N1749, N1738, N1679);
or OR3 (N1750, N1749, N20, N158);
buf BUF1 (N1751, N1729);
nor NOR3 (N1752, N1747, N1501, N310);
nor NOR2 (N1753, N1746, N358);
nand NAND3 (N1754, N1740, N806, N1539);
xor XOR2 (N1755, N1735, N1052);
or OR3 (N1756, N1745, N1503, N1252);
or OR2 (N1757, N1751, N1699);
or OR4 (N1758, N1753, N968, N1634, N1636);
nand NAND4 (N1759, N1755, N1463, N202, N899);
not NOT1 (N1760, N1758);
nand NAND4 (N1761, N1754, N806, N1263, N1446);
and AND2 (N1762, N1752, N1515);
and AND2 (N1763, N1757, N925);
nand NAND2 (N1764, N1744, N1206);
nand NAND3 (N1765, N1727, N108, N979);
nand NAND2 (N1766, N1761, N1027);
or OR2 (N1767, N1756, N845);
buf BUF1 (N1768, N1750);
not NOT1 (N1769, N1759);
and AND3 (N1770, N1765, N1371, N1208);
xor XOR2 (N1771, N1770, N1243);
and AND4 (N1772, N1760, N757, N1183, N1728);
and AND4 (N1773, N1766, N640, N591, N987);
nand NAND4 (N1774, N1762, N199, N1748, N1307);
nand NAND3 (N1775, N1571, N243, N736);
and AND4 (N1776, N1775, N1699, N397, N425);
or OR2 (N1777, N1764, N1140);
or OR2 (N1778, N1774, N1223);
nand NAND2 (N1779, N1776, N152);
or OR3 (N1780, N1768, N630, N402);
nand NAND3 (N1781, N1779, N495, N386);
xor XOR2 (N1782, N1778, N665);
not NOT1 (N1783, N1782);
buf BUF1 (N1784, N1780);
and AND4 (N1785, N1784, N416, N1040, N734);
nand NAND4 (N1786, N1781, N836, N1358, N1588);
buf BUF1 (N1787, N1763);
nand NAND4 (N1788, N1783, N732, N1072, N721);
and AND4 (N1789, N1771, N133, N615, N687);
nand NAND3 (N1790, N1786, N1291, N860);
xor XOR2 (N1791, N1777, N261);
nand NAND4 (N1792, N1767, N267, N403, N990);
nand NAND3 (N1793, N1787, N1218, N1212);
or OR2 (N1794, N1773, N878);
or OR2 (N1795, N1772, N1414);
nor NOR2 (N1796, N1785, N448);
not NOT1 (N1797, N1792);
not NOT1 (N1798, N1788);
nand NAND3 (N1799, N1789, N1631, N639);
or OR3 (N1800, N1797, N163, N863);
nor NOR4 (N1801, N1798, N956, N28, N698);
xor XOR2 (N1802, N1799, N687);
buf BUF1 (N1803, N1796);
or OR2 (N1804, N1795, N1666);
nor NOR3 (N1805, N1793, N257, N1387);
xor XOR2 (N1806, N1804, N531);
xor XOR2 (N1807, N1802, N1582);
nand NAND4 (N1808, N1807, N1672, N1273, N1714);
and AND3 (N1809, N1806, N1490, N478);
or OR3 (N1810, N1809, N1789, N589);
not NOT1 (N1811, N1810);
not NOT1 (N1812, N1800);
not NOT1 (N1813, N1769);
or OR2 (N1814, N1812, N1797);
or OR2 (N1815, N1814, N879);
nand NAND4 (N1816, N1813, N506, N346, N700);
xor XOR2 (N1817, N1811, N206);
xor XOR2 (N1818, N1817, N1005);
nand NAND4 (N1819, N1803, N641, N129, N392);
buf BUF1 (N1820, N1801);
or OR4 (N1821, N1816, N816, N1168, N607);
nor NOR4 (N1822, N1808, N1539, N14, N1717);
xor XOR2 (N1823, N1805, N1031);
buf BUF1 (N1824, N1791);
or OR3 (N1825, N1819, N1333, N541);
xor XOR2 (N1826, N1818, N1359);
buf BUF1 (N1827, N1824);
and AND3 (N1828, N1821, N193, N1663);
nand NAND3 (N1829, N1815, N257, N1339);
and AND2 (N1830, N1827, N1369);
buf BUF1 (N1831, N1828);
xor XOR2 (N1832, N1830, N157);
xor XOR2 (N1833, N1829, N524);
nor NOR2 (N1834, N1833, N325);
or OR3 (N1835, N1820, N632, N1101);
nor NOR4 (N1836, N1825, N115, N938, N1063);
nor NOR3 (N1837, N1835, N241, N557);
nand NAND3 (N1838, N1826, N926, N207);
or OR3 (N1839, N1823, N903, N1191);
and AND4 (N1840, N1837, N1553, N736, N1759);
nand NAND3 (N1841, N1831, N18, N1249);
and AND4 (N1842, N1790, N34, N89, N955);
buf BUF1 (N1843, N1841);
nand NAND4 (N1844, N1834, N1231, N1162, N1224);
and AND2 (N1845, N1832, N1373);
and AND2 (N1846, N1839, N925);
xor XOR2 (N1847, N1840, N1347);
buf BUF1 (N1848, N1838);
buf BUF1 (N1849, N1847);
and AND4 (N1850, N1849, N804, N1258, N386);
nor NOR4 (N1851, N1842, N572, N1079, N1426);
and AND4 (N1852, N1846, N1033, N1667, N1353);
xor XOR2 (N1853, N1794, N770);
nand NAND3 (N1854, N1851, N183, N462);
or OR2 (N1855, N1836, N1723);
not NOT1 (N1856, N1848);
or OR3 (N1857, N1854, N404, N1028);
xor XOR2 (N1858, N1850, N1218);
or OR4 (N1859, N1858, N1810, N346, N777);
nand NAND2 (N1860, N1844, N1032);
buf BUF1 (N1861, N1845);
nor NOR4 (N1862, N1852, N1833, N769, N160);
or OR2 (N1863, N1856, N1639);
not NOT1 (N1864, N1855);
and AND4 (N1865, N1860, N1184, N595, N1044);
and AND4 (N1866, N1861, N608, N1840, N270);
buf BUF1 (N1867, N1862);
and AND2 (N1868, N1863, N633);
or OR3 (N1869, N1868, N156, N377);
buf BUF1 (N1870, N1853);
not NOT1 (N1871, N1857);
buf BUF1 (N1872, N1843);
xor XOR2 (N1873, N1872, N1371);
buf BUF1 (N1874, N1866);
nand NAND2 (N1875, N1822, N927);
xor XOR2 (N1876, N1859, N796);
not NOT1 (N1877, N1864);
nor NOR4 (N1878, N1874, N1104, N596, N1093);
xor XOR2 (N1879, N1875, N1620);
xor XOR2 (N1880, N1871, N1594);
not NOT1 (N1881, N1873);
nand NAND2 (N1882, N1878, N1659);
not NOT1 (N1883, N1869);
xor XOR2 (N1884, N1883, N13);
nand NAND2 (N1885, N1870, N1161);
nand NAND2 (N1886, N1884, N163);
nand NAND2 (N1887, N1877, N449);
not NOT1 (N1888, N1867);
xor XOR2 (N1889, N1886, N1847);
and AND2 (N1890, N1880, N599);
nor NOR3 (N1891, N1885, N989, N1136);
nand NAND4 (N1892, N1889, N170, N1507, N1086);
nand NAND4 (N1893, N1888, N1872, N1131, N791);
or OR2 (N1894, N1892, N123);
or OR4 (N1895, N1881, N925, N553, N816);
buf BUF1 (N1896, N1865);
and AND4 (N1897, N1896, N1403, N116, N1430);
nand NAND3 (N1898, N1895, N1883, N1092);
and AND4 (N1899, N1897, N1061, N1806, N1759);
xor XOR2 (N1900, N1893, N407);
and AND3 (N1901, N1890, N990, N1172);
or OR4 (N1902, N1876, N230, N1797, N949);
xor XOR2 (N1903, N1887, N33);
nor NOR2 (N1904, N1894, N1049);
nor NOR3 (N1905, N1882, N1690, N344);
not NOT1 (N1906, N1905);
or OR2 (N1907, N1901, N1131);
and AND2 (N1908, N1907, N287);
nand NAND2 (N1909, N1899, N1101);
or OR4 (N1910, N1908, N1820, N1386, N1669);
not NOT1 (N1911, N1906);
or OR4 (N1912, N1911, N1698, N438, N1734);
and AND4 (N1913, N1910, N506, N992, N1615);
or OR3 (N1914, N1902, N1039, N1775);
nor NOR3 (N1915, N1914, N1095, N1179);
and AND2 (N1916, N1903, N766);
or OR3 (N1917, N1900, N402, N88);
buf BUF1 (N1918, N1917);
nand NAND4 (N1919, N1879, N1309, N1853, N982);
not NOT1 (N1920, N1912);
nand NAND2 (N1921, N1918, N875);
nand NAND3 (N1922, N1904, N913, N1045);
nor NOR4 (N1923, N1891, N1405, N685, N568);
not NOT1 (N1924, N1898);
nor NOR4 (N1925, N1913, N799, N928, N1625);
or OR2 (N1926, N1921, N193);
and AND3 (N1927, N1926, N226, N875);
xor XOR2 (N1928, N1920, N1748);
xor XOR2 (N1929, N1925, N1248);
and AND3 (N1930, N1909, N104, N1331);
nand NAND3 (N1931, N1927, N1000, N1666);
and AND3 (N1932, N1919, N1209, N1068);
buf BUF1 (N1933, N1929);
and AND3 (N1934, N1924, N1228, N817);
nor NOR4 (N1935, N1923, N1553, N1400, N363);
not NOT1 (N1936, N1928);
nand NAND2 (N1937, N1931, N1823);
and AND4 (N1938, N1922, N467, N378, N256);
not NOT1 (N1939, N1916);
xor XOR2 (N1940, N1937, N1474);
not NOT1 (N1941, N1932);
not NOT1 (N1942, N1939);
or OR4 (N1943, N1940, N766, N823, N1209);
buf BUF1 (N1944, N1941);
nor NOR4 (N1945, N1934, N1493, N801, N766);
nor NOR2 (N1946, N1942, N614);
xor XOR2 (N1947, N1943, N1214);
and AND4 (N1948, N1946, N1238, N1394, N1829);
xor XOR2 (N1949, N1936, N1051);
not NOT1 (N1950, N1935);
xor XOR2 (N1951, N1933, N532);
and AND4 (N1952, N1951, N1205, N678, N1519);
buf BUF1 (N1953, N1945);
and AND4 (N1954, N1944, N1425, N1494, N1352);
or OR2 (N1955, N1947, N1230);
not NOT1 (N1956, N1954);
nor NOR3 (N1957, N1948, N545, N898);
or OR4 (N1958, N1957, N385, N1854, N381);
nand NAND2 (N1959, N1956, N752);
or OR2 (N1960, N1950, N1682);
xor XOR2 (N1961, N1952, N66);
nand NAND2 (N1962, N1949, N1533);
nand NAND3 (N1963, N1961, N1064, N1931);
buf BUF1 (N1964, N1958);
nand NAND2 (N1965, N1959, N1535);
nand NAND3 (N1966, N1915, N1357, N1826);
and AND2 (N1967, N1938, N249);
buf BUF1 (N1968, N1963);
nand NAND3 (N1969, N1965, N613, N217);
nand NAND4 (N1970, N1964, N1702, N46, N711);
or OR4 (N1971, N1968, N1417, N1355, N995);
buf BUF1 (N1972, N1971);
or OR4 (N1973, N1969, N998, N1496, N1429);
or OR4 (N1974, N1955, N791, N1803, N880);
or OR3 (N1975, N1960, N120, N534);
and AND2 (N1976, N1975, N9);
xor XOR2 (N1977, N1930, N220);
not NOT1 (N1978, N1977);
and AND2 (N1979, N1953, N1186);
xor XOR2 (N1980, N1966, N240);
xor XOR2 (N1981, N1979, N1933);
or OR3 (N1982, N1981, N1516, N28);
nor NOR4 (N1983, N1974, N536, N55, N284);
not NOT1 (N1984, N1978);
not NOT1 (N1985, N1976);
not NOT1 (N1986, N1980);
buf BUF1 (N1987, N1983);
buf BUF1 (N1988, N1984);
nand NAND3 (N1989, N1986, N920, N1652);
buf BUF1 (N1990, N1985);
xor XOR2 (N1991, N1973, N1094);
xor XOR2 (N1992, N1991, N874);
xor XOR2 (N1993, N1987, N589);
nand NAND3 (N1994, N1989, N1603, N54);
buf BUF1 (N1995, N1972);
xor XOR2 (N1996, N1993, N822);
not NOT1 (N1997, N1970);
nor NOR2 (N1998, N1988, N768);
buf BUF1 (N1999, N1996);
and AND4 (N2000, N1992, N535, N936, N779);
buf BUF1 (N2001, N1994);
xor XOR2 (N2002, N1995, N703);
not NOT1 (N2003, N1962);
nor NOR4 (N2004, N1998, N1263, N107, N1753);
or OR3 (N2005, N2001, N1518, N353);
nor NOR4 (N2006, N2000, N1321, N1811, N1999);
or OR2 (N2007, N1128, N131);
and AND4 (N2008, N2003, N241, N605, N1149);
nor NOR2 (N2009, N2004, N1269);
not NOT1 (N2010, N2005);
xor XOR2 (N2011, N2006, N1368);
nor NOR2 (N2012, N1990, N1999);
not NOT1 (N2013, N1982);
xor XOR2 (N2014, N2011, N1619);
nand NAND2 (N2015, N2009, N90);
nand NAND2 (N2016, N1967, N932);
not NOT1 (N2017, N2013);
and AND3 (N2018, N2016, N1089, N1594);
buf BUF1 (N2019, N2014);
nand NAND3 (N2020, N2010, N1229, N505);
nor NOR4 (N2021, N2012, N307, N480, N222);
nor NOR2 (N2022, N2019, N1642);
endmodule