// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N202,N208,N212,N169,N214,N198,N209,N201,N215,N216;

or OR3 (N17, N16, N15, N2);
or OR3 (N18, N14, N9, N8);
and AND2 (N19, N3, N13);
buf BUF1 (N20, N6);
buf BUF1 (N21, N18);
nand NAND4 (N22, N12, N14, N18, N3);
nor NOR2 (N23, N10, N11);
and AND3 (N24, N8, N11, N12);
xor XOR2 (N25, N15, N5);
nor NOR2 (N26, N24, N3);
and AND3 (N27, N2, N12, N1);
nand NAND4 (N28, N6, N25, N15, N2);
nor NOR4 (N29, N22, N19, N21, N6);
nand NAND3 (N30, N27, N20, N8);
buf BUF1 (N31, N13);
and AND4 (N32, N24, N8, N10, N20);
or OR4 (N33, N6, N12, N2, N26);
buf BUF1 (N34, N22);
or OR2 (N35, N3, N27);
buf BUF1 (N36, N29);
and AND2 (N37, N36, N6);
buf BUF1 (N38, N37);
nand NAND3 (N39, N30, N34, N38);
nand NAND4 (N40, N5, N12, N37, N25);
buf BUF1 (N41, N21);
nand NAND3 (N42, N23, N2, N15);
or OR4 (N43, N32, N19, N20, N3);
xor XOR2 (N44, N43, N18);
xor XOR2 (N45, N33, N27);
and AND2 (N46, N41, N38);
buf BUF1 (N47, N40);
not NOT1 (N48, N28);
not NOT1 (N49, N35);
not NOT1 (N50, N46);
nor NOR2 (N51, N45, N10);
nand NAND2 (N52, N39, N38);
buf BUF1 (N53, N47);
xor XOR2 (N54, N51, N37);
nor NOR3 (N55, N42, N28, N20);
xor XOR2 (N56, N55, N21);
nor NOR3 (N57, N49, N38, N45);
or OR3 (N58, N31, N53, N19);
and AND4 (N59, N9, N1, N22, N40);
nand NAND4 (N60, N44, N54, N36, N10);
buf BUF1 (N61, N22);
buf BUF1 (N62, N56);
nor NOR3 (N63, N59, N14, N37);
nor NOR3 (N64, N58, N32, N32);
and AND3 (N65, N62, N3, N8);
and AND4 (N66, N17, N35, N15, N45);
or OR3 (N67, N61, N55, N66);
nand NAND4 (N68, N63, N58, N51, N11);
buf BUF1 (N69, N68);
buf BUF1 (N70, N19);
not NOT1 (N71, N52);
xor XOR2 (N72, N50, N67);
not NOT1 (N73, N4);
not NOT1 (N74, N72);
or OR4 (N75, N64, N67, N5, N35);
or OR4 (N76, N57, N4, N1, N42);
xor XOR2 (N77, N65, N53);
nand NAND3 (N78, N69, N21, N33);
xor XOR2 (N79, N75, N23);
or OR4 (N80, N79, N65, N60, N4);
nor NOR4 (N81, N7, N33, N41, N23);
not NOT1 (N82, N76);
or OR4 (N83, N73, N57, N73, N79);
nand NAND3 (N84, N78, N72, N59);
nor NOR3 (N85, N82, N57, N13);
xor XOR2 (N86, N71, N47);
and AND4 (N87, N83, N1, N25, N55);
nand NAND4 (N88, N48, N69, N46, N34);
or OR2 (N89, N88, N30);
nand NAND2 (N90, N84, N59);
not NOT1 (N91, N90);
nand NAND3 (N92, N89, N22, N16);
and AND4 (N93, N86, N85, N50, N48);
not NOT1 (N94, N66);
nand NAND2 (N95, N92, N36);
not NOT1 (N96, N80);
or OR3 (N97, N95, N45, N30);
xor XOR2 (N98, N74, N13);
buf BUF1 (N99, N81);
xor XOR2 (N100, N97, N72);
nor NOR2 (N101, N100, N82);
or OR2 (N102, N70, N93);
nand NAND4 (N103, N49, N61, N78, N90);
nor NOR4 (N104, N102, N90, N28, N28);
buf BUF1 (N105, N104);
nand NAND4 (N106, N101, N1, N8, N53);
buf BUF1 (N107, N99);
buf BUF1 (N108, N107);
not NOT1 (N109, N98);
nand NAND4 (N110, N108, N18, N22, N89);
not NOT1 (N111, N106);
and AND2 (N112, N87, N11);
nor NOR2 (N113, N109, N38);
nor NOR4 (N114, N77, N21, N25, N70);
nor NOR2 (N115, N110, N107);
nand NAND2 (N116, N115, N41);
and AND4 (N117, N96, N82, N96, N104);
or OR3 (N118, N103, N55, N68);
xor XOR2 (N119, N116, N116);
xor XOR2 (N120, N112, N16);
buf BUF1 (N121, N111);
and AND3 (N122, N119, N17, N7);
buf BUF1 (N123, N113);
or OR3 (N124, N114, N122, N122);
xor XOR2 (N125, N83, N52);
nand NAND4 (N126, N94, N8, N12, N26);
and AND3 (N127, N91, N106, N89);
nor NOR3 (N128, N125, N20, N57);
nor NOR2 (N129, N118, N100);
nor NOR2 (N130, N123, N17);
nor NOR2 (N131, N126, N106);
not NOT1 (N132, N130);
not NOT1 (N133, N105);
and AND3 (N134, N120, N39, N123);
xor XOR2 (N135, N129, N117);
xor XOR2 (N136, N48, N109);
nand NAND4 (N137, N121, N97, N50, N100);
xor XOR2 (N138, N128, N43);
or OR3 (N139, N132, N2, N47);
and AND2 (N140, N131, N39);
or OR3 (N141, N140, N20, N5);
and AND3 (N142, N124, N116, N18);
not NOT1 (N143, N142);
nand NAND3 (N144, N133, N121, N84);
not NOT1 (N145, N137);
nand NAND2 (N146, N127, N67);
nand NAND2 (N147, N141, N113);
not NOT1 (N148, N146);
and AND3 (N149, N135, N76, N123);
nand NAND3 (N150, N139, N20, N113);
nor NOR2 (N151, N134, N82);
and AND4 (N152, N147, N28, N32, N136);
xor XOR2 (N153, N47, N9);
buf BUF1 (N154, N152);
xor XOR2 (N155, N149, N78);
not NOT1 (N156, N148);
buf BUF1 (N157, N138);
nand NAND3 (N158, N156, N42, N118);
and AND4 (N159, N153, N141, N142, N40);
xor XOR2 (N160, N143, N118);
buf BUF1 (N161, N158);
xor XOR2 (N162, N159, N44);
xor XOR2 (N163, N151, N50);
buf BUF1 (N164, N150);
and AND3 (N165, N160, N91, N23);
nand NAND3 (N166, N154, N140, N63);
not NOT1 (N167, N157);
nor NOR4 (N168, N165, N97, N132, N153);
xor XOR2 (N169, N168, N76);
nand NAND4 (N170, N162, N22, N123, N62);
nand NAND3 (N171, N155, N89, N72);
and AND2 (N172, N164, N17);
or OR4 (N173, N171, N149, N133, N94);
nand NAND3 (N174, N167, N11, N103);
or OR4 (N175, N144, N81, N141, N130);
not NOT1 (N176, N173);
xor XOR2 (N177, N174, N45);
nand NAND4 (N178, N176, N51, N68, N105);
not NOT1 (N179, N161);
nand NAND3 (N180, N178, N132, N173);
or OR4 (N181, N180, N82, N49, N161);
nor NOR4 (N182, N166, N27, N84, N102);
nand NAND4 (N183, N172, N5, N46, N117);
and AND4 (N184, N170, N111, N88, N131);
and AND3 (N185, N183, N135, N29);
and AND3 (N186, N184, N153, N178);
nand NAND4 (N187, N182, N133, N107, N69);
and AND2 (N188, N163, N150);
xor XOR2 (N189, N187, N159);
buf BUF1 (N190, N175);
nand NAND3 (N191, N185, N76, N162);
buf BUF1 (N192, N145);
not NOT1 (N193, N192);
xor XOR2 (N194, N179, N47);
buf BUF1 (N195, N186);
nor NOR2 (N196, N195, N92);
not NOT1 (N197, N189);
nand NAND3 (N198, N190, N79, N171);
buf BUF1 (N199, N197);
not NOT1 (N200, N177);
buf BUF1 (N201, N191);
buf BUF1 (N202, N181);
nor NOR4 (N203, N200, N188, N18, N107);
not NOT1 (N204, N143);
nor NOR3 (N205, N199, N28, N181);
buf BUF1 (N206, N205);
not NOT1 (N207, N194);
and AND4 (N208, N196, N58, N139, N37);
or OR3 (N209, N193, N125, N95);
buf BUF1 (N210, N203);
buf BUF1 (N211, N207);
xor XOR2 (N212, N204, N46);
or OR4 (N213, N206, N210, N149, N164);
and AND3 (N214, N131, N153, N138);
and AND3 (N215, N211, N113, N213);
not NOT1 (N216, N175);
endmodule