// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N1004,N1012,N1011,N983,N996,N1001,N1005,N1007,N1009,N1013;

not NOT1 (N14, N11);
not NOT1 (N15, N4);
nand NAND2 (N16, N10, N1);
or OR4 (N17, N10, N11, N10, N3);
and AND4 (N18, N4, N5, N16, N2);
or OR2 (N19, N7, N7);
and AND2 (N20, N5, N9);
nand NAND2 (N21, N16, N15);
not NOT1 (N22, N19);
buf BUF1 (N23, N12);
or OR3 (N24, N12, N9, N22);
nor NOR3 (N25, N4, N7, N18);
or OR4 (N26, N16, N7, N23, N6);
nor NOR3 (N27, N13, N8, N24);
nand NAND2 (N28, N7, N22);
buf BUF1 (N29, N18);
buf BUF1 (N30, N9);
xor XOR2 (N31, N25, N27);
and AND3 (N32, N16, N8, N25);
or OR2 (N33, N30, N30);
buf BUF1 (N34, N26);
and AND4 (N35, N17, N16, N16, N7);
buf BUF1 (N36, N21);
or OR2 (N37, N29, N13);
xor XOR2 (N38, N36, N10);
not NOT1 (N39, N37);
xor XOR2 (N40, N32, N28);
nand NAND2 (N41, N9, N28);
buf BUF1 (N42, N33);
nor NOR4 (N43, N42, N23, N12, N12);
not NOT1 (N44, N14);
buf BUF1 (N45, N39);
nor NOR3 (N46, N31, N16, N30);
buf BUF1 (N47, N40);
not NOT1 (N48, N20);
nor NOR2 (N49, N47, N7);
nand NAND4 (N50, N41, N31, N40, N19);
xor XOR2 (N51, N44, N19);
nand NAND2 (N52, N46, N5);
nor NOR4 (N53, N45, N6, N1, N14);
nand NAND3 (N54, N35, N23, N47);
xor XOR2 (N55, N52, N42);
or OR3 (N56, N38, N17, N7);
not NOT1 (N57, N54);
and AND3 (N58, N43, N50, N52);
xor XOR2 (N59, N3, N8);
not NOT1 (N60, N55);
and AND2 (N61, N34, N7);
buf BUF1 (N62, N53);
and AND2 (N63, N58, N58);
nand NAND4 (N64, N61, N41, N50, N56);
not NOT1 (N65, N20);
nand NAND3 (N66, N64, N12, N57);
and AND4 (N67, N49, N65, N49, N34);
not NOT1 (N68, N23);
not NOT1 (N69, N59);
or OR3 (N70, N21, N41, N65);
buf BUF1 (N71, N48);
xor XOR2 (N72, N69, N34);
and AND2 (N73, N63, N38);
nor NOR3 (N74, N66, N48, N37);
or OR4 (N75, N71, N60, N39, N8);
not NOT1 (N76, N20);
xor XOR2 (N77, N67, N73);
xor XOR2 (N78, N42, N57);
not NOT1 (N79, N74);
and AND3 (N80, N79, N67, N67);
or OR4 (N81, N70, N18, N67, N20);
or OR4 (N82, N78, N30, N71, N17);
or OR4 (N83, N80, N64, N64, N35);
nor NOR4 (N84, N76, N13, N11, N43);
not NOT1 (N85, N77);
nor NOR4 (N86, N75, N42, N67, N78);
and AND2 (N87, N85, N59);
xor XOR2 (N88, N83, N10);
not NOT1 (N89, N88);
nand NAND3 (N90, N82, N20, N59);
and AND3 (N91, N90, N82, N59);
not NOT1 (N92, N89);
and AND4 (N93, N68, N48, N83, N53);
and AND3 (N94, N91, N3, N13);
and AND4 (N95, N81, N24, N92, N68);
nor NOR3 (N96, N4, N48, N47);
xor XOR2 (N97, N84, N19);
nor NOR2 (N98, N51, N35);
or OR3 (N99, N72, N18, N69);
nor NOR4 (N100, N62, N75, N88, N33);
nor NOR4 (N101, N97, N31, N8, N95);
nor NOR3 (N102, N55, N94, N76);
not NOT1 (N103, N36);
or OR4 (N104, N103, N16, N89, N67);
buf BUF1 (N105, N98);
nand NAND4 (N106, N101, N7, N39, N60);
nand NAND4 (N107, N105, N40, N102, N87);
and AND4 (N108, N52, N43, N25, N16);
not NOT1 (N109, N95);
nand NAND3 (N110, N93, N59, N4);
buf BUF1 (N111, N99);
xor XOR2 (N112, N111, N99);
xor XOR2 (N113, N104, N74);
and AND2 (N114, N109, N108);
nand NAND4 (N115, N111, N22, N39, N98);
not NOT1 (N116, N86);
buf BUF1 (N117, N107);
nor NOR3 (N118, N114, N68, N47);
and AND4 (N119, N117, N96, N86, N61);
nor NOR3 (N120, N64, N94, N68);
and AND2 (N121, N112, N13);
or OR2 (N122, N100, N34);
nor NOR4 (N123, N116, N10, N82, N80);
and AND4 (N124, N123, N105, N112, N72);
not NOT1 (N125, N110);
buf BUF1 (N126, N115);
nand NAND2 (N127, N121, N68);
not NOT1 (N128, N127);
buf BUF1 (N129, N120);
buf BUF1 (N130, N113);
nand NAND2 (N131, N128, N17);
buf BUF1 (N132, N118);
nor NOR2 (N133, N131, N67);
and AND3 (N134, N125, N73, N122);
and AND4 (N135, N120, N41, N122, N8);
or OR4 (N136, N133, N54, N115, N105);
buf BUF1 (N137, N130);
not NOT1 (N138, N137);
or OR2 (N139, N126, N114);
nor NOR3 (N140, N139, N72, N83);
nand NAND3 (N141, N124, N54, N24);
or OR4 (N142, N135, N98, N67, N38);
or OR4 (N143, N134, N137, N70, N81);
nor NOR4 (N144, N106, N101, N116, N135);
buf BUF1 (N145, N140);
nand NAND3 (N146, N138, N58, N103);
not NOT1 (N147, N143);
and AND4 (N148, N147, N83, N74, N21);
nand NAND4 (N149, N132, N19, N48, N141);
and AND2 (N150, N132, N20);
buf BUF1 (N151, N148);
nand NAND2 (N152, N145, N57);
xor XOR2 (N153, N119, N55);
nand NAND3 (N154, N146, N94, N115);
xor XOR2 (N155, N151, N154);
not NOT1 (N156, N69);
or OR4 (N157, N142, N116, N132, N13);
buf BUF1 (N158, N153);
not NOT1 (N159, N156);
not NOT1 (N160, N157);
nor NOR3 (N161, N158, N33, N46);
nand NAND4 (N162, N160, N78, N105, N31);
nor NOR2 (N163, N152, N12);
and AND2 (N164, N161, N82);
and AND3 (N165, N162, N21, N57);
nor NOR3 (N166, N149, N112, N106);
not NOT1 (N167, N159);
xor XOR2 (N168, N136, N45);
nor NOR4 (N169, N167, N27, N6, N140);
or OR4 (N170, N169, N160, N85, N98);
nand NAND2 (N171, N168, N99);
or OR2 (N172, N163, N118);
nand NAND3 (N173, N172, N143, N165);
not NOT1 (N174, N101);
not NOT1 (N175, N164);
nand NAND4 (N176, N171, N155, N121, N90);
xor XOR2 (N177, N119, N172);
not NOT1 (N178, N175);
not NOT1 (N179, N170);
or OR3 (N180, N173, N162, N178);
or OR3 (N181, N12, N21, N152);
nand NAND2 (N182, N174, N29);
and AND4 (N183, N179, N178, N167, N27);
not NOT1 (N184, N150);
xor XOR2 (N185, N183, N141);
and AND4 (N186, N181, N81, N94, N133);
nand NAND2 (N187, N129, N84);
and AND4 (N188, N182, N69, N93, N27);
and AND2 (N189, N144, N45);
nand NAND3 (N190, N185, N58, N49);
and AND4 (N191, N188, N75, N74, N5);
nand NAND4 (N192, N189, N174, N140, N162);
not NOT1 (N193, N187);
nand NAND3 (N194, N186, N131, N138);
and AND4 (N195, N184, N106, N70, N114);
and AND4 (N196, N166, N111, N32, N182);
nor NOR3 (N197, N176, N77, N77);
and AND2 (N198, N197, N90);
not NOT1 (N199, N194);
and AND2 (N200, N196, N77);
nand NAND3 (N201, N195, N40, N108);
nor NOR2 (N202, N191, N47);
and AND4 (N203, N200, N173, N162, N151);
or OR4 (N204, N192, N103, N157, N102);
and AND2 (N205, N190, N175);
xor XOR2 (N206, N205, N109);
and AND2 (N207, N203, N52);
buf BUF1 (N208, N193);
nor NOR4 (N209, N202, N117, N79, N204);
nor NOR2 (N210, N152, N98);
not NOT1 (N211, N210);
nor NOR2 (N212, N211, N184);
nand NAND4 (N213, N201, N178, N167, N92);
buf BUF1 (N214, N180);
or OR2 (N215, N207, N42);
buf BUF1 (N216, N199);
xor XOR2 (N217, N215, N29);
nor NOR2 (N218, N198, N122);
or OR3 (N219, N177, N51, N150);
not NOT1 (N220, N209);
not NOT1 (N221, N206);
xor XOR2 (N222, N220, N217);
or OR2 (N223, N178, N152);
and AND4 (N224, N213, N180, N74, N106);
buf BUF1 (N225, N216);
nand NAND2 (N226, N222, N63);
nand NAND3 (N227, N208, N54, N204);
and AND4 (N228, N221, N35, N106, N145);
nor NOR4 (N229, N219, N103, N50, N165);
or OR3 (N230, N223, N129, N30);
nor NOR4 (N231, N228, N82, N130, N22);
or OR2 (N232, N225, N167);
nor NOR2 (N233, N227, N26);
not NOT1 (N234, N230);
nand NAND2 (N235, N218, N44);
not NOT1 (N236, N234);
nor NOR4 (N237, N235, N221, N116, N179);
nand NAND2 (N238, N237, N105);
or OR3 (N239, N232, N235, N234);
and AND4 (N240, N212, N190, N166, N97);
and AND2 (N241, N224, N129);
nor NOR3 (N242, N240, N112, N1);
not NOT1 (N243, N242);
not NOT1 (N244, N231);
nor NOR4 (N245, N214, N231, N70, N128);
buf BUF1 (N246, N244);
and AND2 (N247, N233, N159);
or OR4 (N248, N246, N121, N78, N9);
or OR4 (N249, N236, N58, N199, N87);
nor NOR3 (N250, N239, N35, N7);
xor XOR2 (N251, N245, N19);
and AND4 (N252, N238, N90, N246, N36);
buf BUF1 (N253, N241);
xor XOR2 (N254, N248, N101);
buf BUF1 (N255, N254);
buf BUF1 (N256, N251);
nor NOR4 (N257, N250, N134, N98, N66);
nor NOR2 (N258, N255, N60);
not NOT1 (N259, N229);
or OR4 (N260, N256, N57, N73, N80);
or OR4 (N261, N258, N74, N5, N58);
nor NOR3 (N262, N252, N35, N148);
xor XOR2 (N263, N261, N173);
and AND2 (N264, N247, N29);
nand NAND2 (N265, N257, N220);
and AND2 (N266, N263, N220);
nand NAND3 (N267, N266, N160, N194);
xor XOR2 (N268, N253, N65);
xor XOR2 (N269, N264, N36);
xor XOR2 (N270, N267, N99);
nor NOR2 (N271, N265, N151);
xor XOR2 (N272, N259, N174);
and AND4 (N273, N272, N171, N77, N75);
xor XOR2 (N274, N243, N222);
nand NAND4 (N275, N269, N108, N96, N60);
buf BUF1 (N276, N260);
nor NOR4 (N277, N274, N183, N7, N178);
nor NOR4 (N278, N262, N59, N157, N135);
nor NOR4 (N279, N249, N155, N222, N177);
and AND3 (N280, N268, N173, N54);
nand NAND3 (N281, N271, N164, N69);
or OR4 (N282, N277, N31, N84, N255);
or OR3 (N283, N270, N105, N133);
or OR2 (N284, N280, N172);
nand NAND4 (N285, N284, N201, N170, N193);
or OR2 (N286, N275, N44);
not NOT1 (N287, N273);
nor NOR3 (N288, N278, N25, N142);
nor NOR4 (N289, N276, N71, N232, N106);
xor XOR2 (N290, N287, N147);
buf BUF1 (N291, N281);
nor NOR2 (N292, N283, N197);
buf BUF1 (N293, N290);
nor NOR3 (N294, N285, N64, N15);
nor NOR3 (N295, N291, N76, N142);
buf BUF1 (N296, N293);
nor NOR2 (N297, N282, N108);
nor NOR2 (N298, N292, N217);
and AND2 (N299, N288, N41);
not NOT1 (N300, N296);
or OR4 (N301, N289, N193, N190, N122);
nand NAND3 (N302, N286, N59, N144);
or OR2 (N303, N301, N46);
xor XOR2 (N304, N303, N142);
nand NAND3 (N305, N298, N65, N199);
xor XOR2 (N306, N294, N290);
nand NAND2 (N307, N306, N239);
not NOT1 (N308, N302);
buf BUF1 (N309, N304);
nor NOR4 (N310, N308, N56, N176, N73);
and AND4 (N311, N297, N270, N254, N248);
or OR2 (N312, N310, N131);
nor NOR3 (N313, N279, N30, N218);
xor XOR2 (N314, N312, N132);
not NOT1 (N315, N295);
and AND2 (N316, N300, N59);
not NOT1 (N317, N305);
nor NOR3 (N318, N309, N34, N135);
xor XOR2 (N319, N313, N273);
not NOT1 (N320, N307);
nand NAND4 (N321, N318, N209, N202, N76);
xor XOR2 (N322, N319, N81);
or OR3 (N323, N322, N260, N67);
or OR2 (N324, N317, N182);
nand NAND2 (N325, N311, N96);
or OR2 (N326, N324, N146);
or OR3 (N327, N316, N51, N161);
buf BUF1 (N328, N326);
xor XOR2 (N329, N315, N280);
and AND3 (N330, N323, N221, N122);
xor XOR2 (N331, N321, N13);
not NOT1 (N332, N330);
not NOT1 (N333, N327);
xor XOR2 (N334, N329, N188);
xor XOR2 (N335, N325, N209);
buf BUF1 (N336, N299);
and AND3 (N337, N314, N93, N230);
not NOT1 (N338, N332);
and AND2 (N339, N337, N54);
xor XOR2 (N340, N328, N204);
or OR4 (N341, N338, N241, N25, N240);
nor NOR2 (N342, N320, N206);
nor NOR3 (N343, N333, N10, N177);
buf BUF1 (N344, N339);
or OR3 (N345, N336, N287, N90);
nor NOR3 (N346, N344, N99, N264);
not NOT1 (N347, N342);
xor XOR2 (N348, N340, N165);
and AND4 (N349, N346, N2, N307, N328);
nand NAND4 (N350, N349, N310, N34, N76);
nor NOR4 (N351, N341, N153, N101, N30);
or OR3 (N352, N334, N194, N65);
buf BUF1 (N353, N348);
nand NAND3 (N354, N226, N192, N83);
or OR4 (N355, N331, N255, N353, N327);
buf BUF1 (N356, N286);
not NOT1 (N357, N343);
not NOT1 (N358, N352);
and AND4 (N359, N351, N187, N306, N344);
or OR2 (N360, N359, N39);
buf BUF1 (N361, N357);
buf BUF1 (N362, N354);
buf BUF1 (N363, N335);
not NOT1 (N364, N350);
nand NAND2 (N365, N358, N345);
xor XOR2 (N366, N190, N241);
xor XOR2 (N367, N363, N267);
or OR3 (N368, N355, N328, N204);
not NOT1 (N369, N368);
nand NAND4 (N370, N364, N133, N304, N350);
and AND2 (N371, N365, N240);
nor NOR2 (N372, N361, N216);
not NOT1 (N373, N356);
and AND3 (N374, N367, N42, N122);
or OR4 (N375, N362, N215, N306, N89);
xor XOR2 (N376, N347, N359);
xor XOR2 (N377, N369, N360);
or OR2 (N378, N195, N359);
or OR2 (N379, N373, N248);
nand NAND3 (N380, N366, N131, N164);
and AND4 (N381, N377, N213, N159, N166);
nand NAND2 (N382, N374, N211);
xor XOR2 (N383, N380, N367);
buf BUF1 (N384, N370);
buf BUF1 (N385, N381);
not NOT1 (N386, N378);
not NOT1 (N387, N379);
xor XOR2 (N388, N375, N184);
xor XOR2 (N389, N371, N314);
xor XOR2 (N390, N372, N300);
buf BUF1 (N391, N389);
nand NAND3 (N392, N385, N103, N138);
buf BUF1 (N393, N391);
or OR2 (N394, N390, N392);
xor XOR2 (N395, N200, N120);
not NOT1 (N396, N394);
nor NOR3 (N397, N383, N38, N58);
or OR4 (N398, N376, N113, N36, N209);
and AND4 (N399, N397, N132, N108, N162);
or OR2 (N400, N399, N360);
nand NAND4 (N401, N396, N50, N58, N91);
nand NAND3 (N402, N386, N172, N104);
and AND3 (N403, N402, N38, N339);
not NOT1 (N404, N384);
xor XOR2 (N405, N401, N122);
nand NAND3 (N406, N388, N39, N101);
xor XOR2 (N407, N398, N289);
nor NOR4 (N408, N405, N67, N33, N83);
xor XOR2 (N409, N408, N163);
xor XOR2 (N410, N409, N283);
not NOT1 (N411, N382);
nand NAND4 (N412, N410, N104, N236, N237);
not NOT1 (N413, N395);
nand NAND2 (N414, N412, N51);
not NOT1 (N415, N403);
not NOT1 (N416, N411);
xor XOR2 (N417, N387, N51);
and AND3 (N418, N400, N253, N263);
xor XOR2 (N419, N415, N243);
not NOT1 (N420, N418);
nor NOR3 (N421, N414, N60, N81);
xor XOR2 (N422, N393, N118);
buf BUF1 (N423, N407);
nand NAND2 (N424, N404, N5);
xor XOR2 (N425, N422, N95);
nor NOR2 (N426, N413, N191);
not NOT1 (N427, N424);
xor XOR2 (N428, N426, N51);
buf BUF1 (N429, N417);
buf BUF1 (N430, N406);
xor XOR2 (N431, N425, N166);
buf BUF1 (N432, N428);
nor NOR3 (N433, N423, N285, N114);
buf BUF1 (N434, N430);
nand NAND2 (N435, N427, N174);
not NOT1 (N436, N435);
buf BUF1 (N437, N436);
nor NOR4 (N438, N419, N131, N220, N309);
or OR3 (N439, N431, N254, N369);
not NOT1 (N440, N434);
not NOT1 (N441, N432);
and AND4 (N442, N438, N138, N339, N231);
not NOT1 (N443, N433);
not NOT1 (N444, N421);
xor XOR2 (N445, N444, N420);
nand NAND3 (N446, N429, N371, N278);
xor XOR2 (N447, N160, N279);
xor XOR2 (N448, N437, N76);
buf BUF1 (N449, N443);
and AND3 (N450, N449, N419, N340);
nand NAND4 (N451, N446, N440, N194, N386);
buf BUF1 (N452, N64);
and AND2 (N453, N450, N222);
xor XOR2 (N454, N445, N379);
xor XOR2 (N455, N452, N113);
nor NOR3 (N456, N439, N349, N274);
not NOT1 (N457, N447);
buf BUF1 (N458, N453);
or OR3 (N459, N457, N31, N358);
nor NOR3 (N460, N454, N269, N76);
nand NAND2 (N461, N456, N57);
not NOT1 (N462, N448);
nand NAND4 (N463, N461, N124, N31, N270);
buf BUF1 (N464, N463);
and AND3 (N465, N455, N6, N209);
and AND3 (N466, N451, N253, N72);
xor XOR2 (N467, N441, N119);
and AND3 (N468, N458, N361, N195);
xor XOR2 (N469, N416, N450);
not NOT1 (N470, N468);
not NOT1 (N471, N462);
nor NOR3 (N472, N466, N202, N3);
or OR3 (N473, N470, N6, N418);
and AND2 (N474, N469, N378);
not NOT1 (N475, N464);
buf BUF1 (N476, N472);
or OR4 (N477, N473, N77, N312, N263);
not NOT1 (N478, N467);
nor NOR4 (N479, N465, N266, N167, N136);
nor NOR2 (N480, N460, N229);
and AND3 (N481, N474, N463, N410);
nor NOR2 (N482, N475, N38);
not NOT1 (N483, N479);
or OR2 (N484, N481, N465);
and AND2 (N485, N482, N58);
and AND4 (N486, N478, N276, N208, N13);
nor NOR4 (N487, N483, N48, N402, N453);
xor XOR2 (N488, N442, N486);
or OR2 (N489, N120, N244);
buf BUF1 (N490, N459);
and AND4 (N491, N488, N373, N488, N274);
buf BUF1 (N492, N471);
or OR3 (N493, N490, N64, N355);
nor NOR3 (N494, N492, N26, N314);
not NOT1 (N495, N493);
xor XOR2 (N496, N494, N201);
and AND2 (N497, N485, N445);
and AND4 (N498, N495, N11, N428, N292);
nand NAND3 (N499, N489, N436, N364);
buf BUF1 (N500, N499);
not NOT1 (N501, N498);
or OR4 (N502, N497, N438, N267, N8);
nand NAND4 (N503, N501, N143, N70, N68);
not NOT1 (N504, N487);
nand NAND4 (N505, N476, N333, N240, N5);
and AND3 (N506, N491, N378, N209);
xor XOR2 (N507, N477, N242);
nand NAND3 (N508, N496, N357, N315);
nor NOR4 (N509, N503, N287, N434, N92);
or OR4 (N510, N502, N475, N159, N76);
not NOT1 (N511, N505);
or OR3 (N512, N507, N401, N47);
nor NOR4 (N513, N506, N182, N218, N433);
nor NOR4 (N514, N512, N96, N489, N407);
not NOT1 (N515, N480);
nor NOR3 (N516, N511, N391, N299);
and AND2 (N517, N515, N318);
buf BUF1 (N518, N484);
buf BUF1 (N519, N509);
xor XOR2 (N520, N516, N362);
nor NOR4 (N521, N518, N101, N18, N481);
or OR2 (N522, N520, N374);
buf BUF1 (N523, N519);
not NOT1 (N524, N517);
or OR3 (N525, N513, N454, N130);
or OR2 (N526, N510, N206);
nand NAND3 (N527, N500, N216, N110);
nor NOR3 (N528, N523, N146, N19);
nor NOR4 (N529, N504, N326, N523, N57);
nand NAND4 (N530, N508, N214, N482, N347);
xor XOR2 (N531, N524, N107);
not NOT1 (N532, N531);
and AND4 (N533, N514, N127, N32, N168);
not NOT1 (N534, N529);
buf BUF1 (N535, N533);
and AND3 (N536, N522, N260, N401);
nor NOR3 (N537, N530, N251, N263);
buf BUF1 (N538, N534);
nor NOR3 (N539, N538, N49, N141);
nor NOR2 (N540, N525, N287);
nand NAND3 (N541, N539, N229, N361);
and AND3 (N542, N535, N527, N233);
nor NOR4 (N543, N16, N28, N136, N67);
not NOT1 (N544, N526);
or OR3 (N545, N537, N195, N23);
or OR3 (N546, N540, N432, N410);
not NOT1 (N547, N521);
nor NOR3 (N548, N546, N174, N270);
and AND3 (N549, N532, N7, N93);
nor NOR2 (N550, N548, N52);
nand NAND4 (N551, N536, N40, N226, N324);
buf BUF1 (N552, N551);
nor NOR4 (N553, N544, N491, N518, N472);
nor NOR2 (N554, N552, N186);
nand NAND3 (N555, N545, N528, N529);
nor NOR3 (N556, N555, N503, N490);
and AND2 (N557, N10, N501);
nor NOR4 (N558, N549, N426, N433, N458);
nor NOR3 (N559, N541, N521, N425);
and AND2 (N560, N543, N415);
xor XOR2 (N561, N556, N232);
and AND2 (N562, N560, N184);
nor NOR4 (N563, N547, N337, N13, N312);
buf BUF1 (N564, N554);
buf BUF1 (N565, N550);
and AND4 (N566, N557, N459, N327, N253);
or OR3 (N567, N566, N446, N438);
buf BUF1 (N568, N562);
nor NOR3 (N569, N542, N115, N525);
not NOT1 (N570, N558);
not NOT1 (N571, N565);
xor XOR2 (N572, N569, N311);
and AND3 (N573, N571, N183, N36);
nand NAND4 (N574, N573, N450, N350, N278);
and AND3 (N575, N568, N23, N440);
nor NOR4 (N576, N572, N148, N353, N239);
nor NOR2 (N577, N567, N397);
not NOT1 (N578, N577);
nor NOR2 (N579, N564, N91);
or OR3 (N580, N578, N486, N205);
not NOT1 (N581, N570);
nor NOR4 (N582, N580, N482, N376, N352);
buf BUF1 (N583, N579);
or OR2 (N584, N561, N415);
nor NOR2 (N585, N559, N198);
and AND3 (N586, N574, N168, N387);
nand NAND2 (N587, N586, N576);
or OR3 (N588, N342, N211, N159);
nor NOR2 (N589, N588, N311);
nand NAND2 (N590, N553, N59);
buf BUF1 (N591, N581);
or OR2 (N592, N563, N583);
or OR3 (N593, N246, N338, N115);
xor XOR2 (N594, N587, N185);
xor XOR2 (N595, N590, N381);
nand NAND3 (N596, N582, N73, N583);
xor XOR2 (N597, N595, N227);
not NOT1 (N598, N585);
and AND2 (N599, N597, N211);
nor NOR2 (N600, N584, N115);
and AND3 (N601, N589, N59, N476);
xor XOR2 (N602, N593, N274);
and AND2 (N603, N596, N52);
or OR2 (N604, N598, N511);
buf BUF1 (N605, N603);
buf BUF1 (N606, N575);
not NOT1 (N607, N601);
nor NOR4 (N608, N594, N147, N579, N415);
not NOT1 (N609, N605);
and AND4 (N610, N591, N332, N267, N337);
not NOT1 (N611, N609);
xor XOR2 (N612, N606, N449);
nor NOR4 (N613, N612, N179, N447, N593);
or OR3 (N614, N602, N311, N558);
buf BUF1 (N615, N614);
nand NAND2 (N616, N600, N240);
nand NAND3 (N617, N604, N33, N308);
and AND4 (N618, N615, N120, N570, N227);
xor XOR2 (N619, N616, N137);
nand NAND2 (N620, N611, N288);
and AND3 (N621, N610, N393, N295);
nand NAND3 (N622, N607, N352, N372);
or OR2 (N623, N618, N515);
and AND2 (N624, N608, N86);
xor XOR2 (N625, N617, N400);
xor XOR2 (N626, N624, N257);
not NOT1 (N627, N620);
and AND3 (N628, N625, N406, N76);
not NOT1 (N629, N622);
xor XOR2 (N630, N619, N524);
buf BUF1 (N631, N613);
and AND3 (N632, N599, N461, N518);
nand NAND2 (N633, N628, N235);
or OR3 (N634, N592, N276, N574);
buf BUF1 (N635, N630);
buf BUF1 (N636, N633);
buf BUF1 (N637, N632);
not NOT1 (N638, N627);
or OR4 (N639, N638, N98, N97, N117);
nand NAND2 (N640, N629, N265);
nand NAND3 (N641, N639, N532, N553);
not NOT1 (N642, N634);
and AND3 (N643, N631, N606, N521);
or OR3 (N644, N642, N360, N408);
xor XOR2 (N645, N641, N158);
xor XOR2 (N646, N635, N391);
nand NAND2 (N647, N645, N625);
nor NOR4 (N648, N621, N52, N608, N535);
nand NAND3 (N649, N646, N362, N399);
and AND3 (N650, N648, N261, N332);
nand NAND2 (N651, N647, N137);
not NOT1 (N652, N623);
not NOT1 (N653, N643);
nand NAND3 (N654, N626, N240, N266);
nor NOR2 (N655, N649, N113);
or OR3 (N656, N654, N593, N51);
or OR2 (N657, N640, N158);
and AND3 (N658, N637, N373, N34);
nand NAND3 (N659, N650, N576, N567);
nor NOR2 (N660, N655, N62);
nand NAND2 (N661, N656, N345);
or OR4 (N662, N636, N15, N58, N605);
buf BUF1 (N663, N653);
xor XOR2 (N664, N661, N260);
and AND3 (N665, N662, N253, N259);
nor NOR2 (N666, N660, N289);
or OR3 (N667, N666, N298, N657);
not NOT1 (N668, N67);
nand NAND3 (N669, N658, N37, N591);
buf BUF1 (N670, N664);
or OR3 (N671, N669, N546, N579);
buf BUF1 (N672, N665);
nor NOR2 (N673, N671, N122);
buf BUF1 (N674, N659);
and AND3 (N675, N644, N58, N95);
buf BUF1 (N676, N670);
xor XOR2 (N677, N663, N276);
nor NOR2 (N678, N672, N160);
nand NAND2 (N679, N677, N286);
nand NAND3 (N680, N674, N579, N371);
nor NOR2 (N681, N668, N583);
not NOT1 (N682, N652);
and AND4 (N683, N673, N556, N336, N664);
nand NAND4 (N684, N680, N160, N554, N212);
or OR2 (N685, N678, N306);
buf BUF1 (N686, N667);
not NOT1 (N687, N682);
or OR3 (N688, N683, N502, N94);
nor NOR2 (N689, N688, N362);
xor XOR2 (N690, N685, N75);
or OR2 (N691, N675, N482);
and AND3 (N692, N651, N518, N555);
not NOT1 (N693, N681);
or OR2 (N694, N690, N136);
nand NAND2 (N695, N684, N217);
buf BUF1 (N696, N691);
xor XOR2 (N697, N689, N504);
buf BUF1 (N698, N679);
xor XOR2 (N699, N693, N461);
xor XOR2 (N700, N699, N494);
xor XOR2 (N701, N695, N74);
or OR3 (N702, N698, N619, N478);
buf BUF1 (N703, N676);
or OR2 (N704, N701, N176);
nand NAND3 (N705, N694, N296, N57);
or OR2 (N706, N692, N149);
nand NAND4 (N707, N700, N518, N346, N117);
or OR4 (N708, N706, N499, N703, N598);
not NOT1 (N709, N399);
xor XOR2 (N710, N702, N90);
or OR2 (N711, N707, N550);
nand NAND4 (N712, N710, N518, N491, N276);
xor XOR2 (N713, N686, N514);
xor XOR2 (N714, N708, N544);
nor NOR3 (N715, N712, N463, N482);
buf BUF1 (N716, N714);
or OR2 (N717, N705, N503);
buf BUF1 (N718, N696);
or OR2 (N719, N687, N620);
nand NAND2 (N720, N697, N256);
buf BUF1 (N721, N720);
buf BUF1 (N722, N717);
nor NOR4 (N723, N709, N316, N127, N678);
or OR3 (N724, N711, N195, N489);
buf BUF1 (N725, N719);
and AND2 (N726, N722, N191);
or OR4 (N727, N704, N72, N649, N385);
not NOT1 (N728, N713);
not NOT1 (N729, N723);
nand NAND2 (N730, N724, N693);
xor XOR2 (N731, N727, N80);
or OR3 (N732, N718, N689, N708);
xor XOR2 (N733, N732, N422);
nand NAND3 (N734, N716, N316, N572);
buf BUF1 (N735, N733);
xor XOR2 (N736, N726, N466);
nand NAND4 (N737, N725, N412, N609, N181);
not NOT1 (N738, N737);
nor NOR2 (N739, N730, N131);
and AND4 (N740, N736, N697, N140, N534);
nor NOR3 (N741, N729, N43, N507);
buf BUF1 (N742, N741);
xor XOR2 (N743, N742, N401);
buf BUF1 (N744, N731);
and AND4 (N745, N744, N460, N513, N355);
nand NAND4 (N746, N740, N341, N326, N666);
nor NOR4 (N747, N721, N293, N559, N159);
nand NAND2 (N748, N745, N722);
and AND2 (N749, N735, N516);
xor XOR2 (N750, N739, N204);
or OR4 (N751, N728, N164, N525, N486);
xor XOR2 (N752, N747, N616);
nand NAND2 (N753, N746, N504);
buf BUF1 (N754, N750);
xor XOR2 (N755, N748, N414);
and AND2 (N756, N749, N666);
buf BUF1 (N757, N715);
or OR3 (N758, N757, N180, N555);
nand NAND4 (N759, N738, N167, N122, N511);
not NOT1 (N760, N759);
not NOT1 (N761, N753);
nor NOR4 (N762, N754, N411, N740, N419);
and AND2 (N763, N752, N433);
nand NAND2 (N764, N756, N151);
buf BUF1 (N765, N758);
and AND4 (N766, N734, N118, N28, N50);
xor XOR2 (N767, N751, N303);
not NOT1 (N768, N755);
nor NOR4 (N769, N766, N336, N286, N671);
xor XOR2 (N770, N761, N759);
buf BUF1 (N771, N743);
buf BUF1 (N772, N760);
and AND3 (N773, N768, N311, N614);
and AND4 (N774, N762, N673, N224, N319);
not NOT1 (N775, N765);
nor NOR4 (N776, N769, N533, N470, N709);
nor NOR3 (N777, N771, N465, N100);
or OR4 (N778, N774, N19, N326, N777);
xor XOR2 (N779, N175, N649);
nand NAND2 (N780, N778, N119);
not NOT1 (N781, N775);
or OR4 (N782, N779, N9, N276, N375);
nand NAND2 (N783, N780, N357);
not NOT1 (N784, N772);
nand NAND3 (N785, N763, N425, N779);
not NOT1 (N786, N764);
nand NAND4 (N787, N786, N665, N539, N588);
xor XOR2 (N788, N784, N471);
and AND2 (N789, N773, N775);
not NOT1 (N790, N782);
or OR3 (N791, N789, N408, N324);
buf BUF1 (N792, N788);
buf BUF1 (N793, N787);
nand NAND4 (N794, N781, N566, N146, N684);
xor XOR2 (N795, N770, N108);
and AND2 (N796, N795, N270);
nand NAND3 (N797, N767, N502, N779);
nand NAND3 (N798, N794, N540, N2);
nor NOR3 (N799, N798, N665, N7);
nand NAND4 (N800, N790, N791, N299, N465);
xor XOR2 (N801, N672, N75);
not NOT1 (N802, N796);
nand NAND3 (N803, N797, N123, N23);
not NOT1 (N804, N799);
buf BUF1 (N805, N776);
buf BUF1 (N806, N793);
or OR4 (N807, N800, N269, N166, N713);
nand NAND2 (N808, N804, N692);
or OR2 (N809, N808, N432);
and AND2 (N810, N792, N409);
buf BUF1 (N811, N805);
not NOT1 (N812, N807);
nand NAND3 (N813, N806, N84, N276);
nor NOR3 (N814, N801, N356, N720);
xor XOR2 (N815, N783, N50);
nor NOR3 (N816, N810, N271, N447);
xor XOR2 (N817, N813, N632);
not NOT1 (N818, N816);
or OR2 (N819, N815, N183);
nor NOR3 (N820, N809, N99, N591);
xor XOR2 (N821, N812, N777);
nor NOR4 (N822, N820, N318, N429, N117);
buf BUF1 (N823, N819);
not NOT1 (N824, N817);
xor XOR2 (N825, N803, N9);
buf BUF1 (N826, N818);
or OR3 (N827, N814, N327, N536);
not NOT1 (N828, N785);
not NOT1 (N829, N828);
nand NAND4 (N830, N811, N213, N682, N528);
and AND3 (N831, N826, N340, N99);
and AND3 (N832, N802, N589, N72);
buf BUF1 (N833, N824);
nand NAND4 (N834, N832, N407, N607, N176);
and AND3 (N835, N830, N35, N531);
xor XOR2 (N836, N821, N390);
not NOT1 (N837, N825);
nand NAND3 (N838, N834, N765, N163);
nor NOR3 (N839, N829, N423, N253);
nand NAND3 (N840, N835, N426, N538);
not NOT1 (N841, N836);
nand NAND4 (N842, N840, N705, N642, N547);
and AND3 (N843, N842, N142, N554);
not NOT1 (N844, N827);
nor NOR4 (N845, N843, N708, N562, N679);
not NOT1 (N846, N823);
nand NAND2 (N847, N845, N538);
nor NOR4 (N848, N837, N838, N544, N576);
buf BUF1 (N849, N235);
and AND3 (N850, N833, N315, N631);
nand NAND4 (N851, N849, N607, N665, N292);
not NOT1 (N852, N839);
or OR2 (N853, N850, N761);
nand NAND4 (N854, N841, N665, N397, N324);
xor XOR2 (N855, N854, N779);
buf BUF1 (N856, N848);
not NOT1 (N857, N856);
nor NOR3 (N858, N831, N747, N393);
buf BUF1 (N859, N851);
nor NOR4 (N860, N844, N680, N75, N281);
xor XOR2 (N861, N846, N256);
or OR2 (N862, N855, N4);
buf BUF1 (N863, N852);
not NOT1 (N864, N863);
not NOT1 (N865, N862);
nor NOR3 (N866, N865, N450, N697);
buf BUF1 (N867, N857);
or OR3 (N868, N864, N143, N2);
and AND2 (N869, N867, N84);
and AND3 (N870, N859, N97, N489);
and AND2 (N871, N847, N189);
buf BUF1 (N872, N822);
nor NOR4 (N873, N868, N381, N271, N846);
nand NAND2 (N874, N869, N159);
nand NAND3 (N875, N860, N99, N675);
nand NAND3 (N876, N872, N388, N656);
not NOT1 (N877, N873);
nand NAND3 (N878, N870, N176, N256);
buf BUF1 (N879, N876);
nor NOR3 (N880, N866, N598, N710);
not NOT1 (N881, N874);
nor NOR2 (N882, N881, N477);
xor XOR2 (N883, N880, N7);
nand NAND4 (N884, N853, N740, N431, N860);
not NOT1 (N885, N877);
and AND3 (N886, N882, N569, N449);
buf BUF1 (N887, N858);
or OR4 (N888, N875, N358, N334, N89);
and AND4 (N889, N886, N527, N635, N791);
buf BUF1 (N890, N885);
or OR2 (N891, N878, N439);
nand NAND2 (N892, N879, N756);
xor XOR2 (N893, N883, N555);
nor NOR4 (N894, N890, N104, N404, N809);
buf BUF1 (N895, N887);
xor XOR2 (N896, N888, N324);
and AND4 (N897, N891, N225, N384, N832);
xor XOR2 (N898, N895, N830);
xor XOR2 (N899, N894, N706);
not NOT1 (N900, N892);
nand NAND4 (N901, N900, N468, N801, N34);
xor XOR2 (N902, N889, N83);
and AND4 (N903, N901, N650, N275, N446);
xor XOR2 (N904, N897, N331);
and AND3 (N905, N884, N313, N122);
not NOT1 (N906, N904);
not NOT1 (N907, N902);
nor NOR3 (N908, N861, N828, N249);
and AND2 (N909, N907, N24);
nor NOR4 (N910, N899, N686, N824, N23);
nand NAND4 (N911, N906, N660, N42, N803);
nor NOR2 (N912, N911, N374);
xor XOR2 (N913, N903, N731);
xor XOR2 (N914, N913, N364);
nor NOR2 (N915, N908, N396);
not NOT1 (N916, N909);
nand NAND4 (N917, N915, N767, N453, N433);
or OR3 (N918, N914, N493, N691);
xor XOR2 (N919, N905, N190);
buf BUF1 (N920, N898);
nand NAND3 (N921, N896, N801, N167);
or OR3 (N922, N920, N432, N583);
nor NOR4 (N923, N893, N700, N691, N614);
buf BUF1 (N924, N917);
nor NOR4 (N925, N910, N794, N666, N639);
nand NAND4 (N926, N912, N155, N672, N168);
nor NOR3 (N927, N922, N490, N204);
and AND2 (N928, N916, N15);
buf BUF1 (N929, N925);
and AND4 (N930, N921, N854, N82, N387);
nand NAND4 (N931, N927, N120, N552, N440);
buf BUF1 (N932, N919);
xor XOR2 (N933, N928, N818);
and AND4 (N934, N932, N523, N367, N267);
or OR3 (N935, N929, N859, N199);
buf BUF1 (N936, N924);
xor XOR2 (N937, N936, N621);
nor NOR3 (N938, N926, N329, N816);
not NOT1 (N939, N934);
and AND3 (N940, N938, N56, N77);
and AND4 (N941, N933, N411, N821, N30);
buf BUF1 (N942, N937);
nand NAND3 (N943, N918, N235, N453);
buf BUF1 (N944, N943);
nand NAND3 (N945, N941, N940, N151);
not NOT1 (N946, N715);
and AND4 (N947, N931, N338, N744, N530);
nand NAND4 (N948, N946, N917, N579, N808);
and AND2 (N949, N939, N345);
nor NOR4 (N950, N947, N863, N267, N874);
and AND4 (N951, N930, N271, N407, N411);
or OR4 (N952, N871, N832, N878, N466);
buf BUF1 (N953, N945);
and AND4 (N954, N949, N568, N27, N434);
or OR2 (N955, N953, N512);
or OR3 (N956, N935, N509, N55);
xor XOR2 (N957, N950, N100);
nor NOR2 (N958, N952, N574);
or OR2 (N959, N955, N559);
xor XOR2 (N960, N954, N866);
not NOT1 (N961, N948);
nor NOR4 (N962, N942, N255, N487, N776);
xor XOR2 (N963, N923, N374);
and AND3 (N964, N956, N176, N350);
not NOT1 (N965, N964);
nand NAND4 (N966, N959, N88, N589, N861);
not NOT1 (N967, N961);
xor XOR2 (N968, N962, N211);
or OR4 (N969, N963, N642, N838, N362);
and AND3 (N970, N966, N385, N250);
or OR4 (N971, N969, N211, N221, N870);
and AND2 (N972, N967, N411);
and AND2 (N973, N965, N220);
not NOT1 (N974, N972);
and AND2 (N975, N944, N613);
buf BUF1 (N976, N960);
or OR4 (N977, N973, N514, N835, N171);
and AND2 (N978, N970, N287);
nor NOR2 (N979, N968, N293);
or OR4 (N980, N978, N301, N792, N502);
not NOT1 (N981, N980);
and AND2 (N982, N979, N363);
nor NOR4 (N983, N977, N229, N410, N123);
xor XOR2 (N984, N971, N800);
nor NOR2 (N985, N976, N527);
not NOT1 (N986, N975);
buf BUF1 (N987, N982);
and AND3 (N988, N985, N707, N374);
and AND4 (N989, N986, N120, N651, N79);
buf BUF1 (N990, N988);
not NOT1 (N991, N989);
nand NAND2 (N992, N987, N701);
xor XOR2 (N993, N992, N855);
nor NOR4 (N994, N990, N755, N100, N133);
nand NAND4 (N995, N958, N251, N169, N566);
xor XOR2 (N996, N995, N197);
not NOT1 (N997, N957);
nor NOR3 (N998, N997, N476, N616);
or OR4 (N999, N998, N393, N522, N699);
xor XOR2 (N1000, N991, N654);
nor NOR3 (N1001, N999, N666, N892);
nor NOR4 (N1002, N993, N807, N485, N998);
xor XOR2 (N1003, N1000, N836);
or OR4 (N1004, N981, N63, N37, N476);
buf BUF1 (N1005, N1003);
nand NAND2 (N1006, N974, N531);
and AND3 (N1007, N1002, N646, N598);
and AND2 (N1008, N994, N926);
not NOT1 (N1009, N951);
buf BUF1 (N1010, N984);
buf BUF1 (N1011, N1008);
nor NOR4 (N1012, N1010, N251, N184, N744);
or OR4 (N1013, N1006, N401, N85, N2);
endmodule