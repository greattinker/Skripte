// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N909,N888,N912,N894,N901,N911,N906,N903,N902,N913;

xor XOR2 (N14, N7, N8);
or OR2 (N15, N2, N11);
xor XOR2 (N16, N13, N15);
xor XOR2 (N17, N10, N5);
and AND3 (N18, N16, N15, N3);
nor NOR4 (N19, N14, N4, N8, N18);
and AND4 (N20, N16, N19, N12, N13);
and AND4 (N21, N3, N13, N14, N10);
or OR4 (N22, N21, N3, N13, N3);
not NOT1 (N23, N9);
nor NOR4 (N24, N2, N14, N1, N11);
buf BUF1 (N25, N5);
buf BUF1 (N26, N6);
or OR4 (N27, N1, N8, N14, N6);
nor NOR3 (N28, N17, N27, N18);
buf BUF1 (N29, N6);
xor XOR2 (N30, N15, N11);
xor XOR2 (N31, N7, N2);
not NOT1 (N32, N30);
xor XOR2 (N33, N29, N23);
or OR4 (N34, N22, N32, N17, N21);
xor XOR2 (N35, N26, N7);
buf BUF1 (N36, N22);
or OR3 (N37, N36, N2, N27);
or OR3 (N38, N15, N13, N10);
or OR2 (N39, N31, N19);
or OR4 (N40, N34, N31, N31, N19);
buf BUF1 (N41, N39);
nor NOR3 (N42, N41, N18, N10);
or OR2 (N43, N33, N41);
xor XOR2 (N44, N42, N41);
not NOT1 (N45, N35);
not NOT1 (N46, N45);
or OR2 (N47, N40, N4);
and AND2 (N48, N20, N15);
nor NOR3 (N49, N46, N47, N36);
nand NAND4 (N50, N27, N24, N29, N23);
nand NAND3 (N51, N45, N20, N46);
nand NAND2 (N52, N48, N24);
xor XOR2 (N53, N37, N52);
or OR4 (N54, N48, N47, N25, N33);
nor NOR2 (N55, N34, N5);
or OR2 (N56, N54, N48);
nand NAND3 (N57, N56, N55, N39);
or OR3 (N58, N36, N34, N18);
or OR3 (N59, N38, N22, N42);
nor NOR4 (N60, N57, N14, N7, N51);
and AND3 (N61, N59, N54, N30);
not NOT1 (N62, N5);
nand NAND2 (N63, N60, N16);
xor XOR2 (N64, N50, N50);
nand NAND3 (N65, N49, N35, N7);
and AND3 (N66, N28, N51, N21);
buf BUF1 (N67, N61);
buf BUF1 (N68, N67);
xor XOR2 (N69, N63, N32);
nor NOR3 (N70, N66, N31, N6);
or OR2 (N71, N53, N31);
and AND2 (N72, N68, N33);
xor XOR2 (N73, N62, N49);
xor XOR2 (N74, N69, N70);
or OR2 (N75, N66, N20);
or OR3 (N76, N72, N44, N61);
xor XOR2 (N77, N46, N33);
and AND2 (N78, N74, N74);
xor XOR2 (N79, N77, N39);
and AND2 (N80, N79, N51);
nand NAND2 (N81, N71, N46);
nand NAND4 (N82, N64, N2, N15, N45);
nand NAND3 (N83, N81, N11, N37);
buf BUF1 (N84, N58);
not NOT1 (N85, N82);
not NOT1 (N86, N84);
xor XOR2 (N87, N80, N52);
not NOT1 (N88, N85);
xor XOR2 (N89, N86, N4);
xor XOR2 (N90, N87, N19);
buf BUF1 (N91, N78);
or OR3 (N92, N73, N30, N6);
nor NOR4 (N93, N91, N23, N87, N6);
xor XOR2 (N94, N83, N85);
nor NOR4 (N95, N89, N5, N77, N91);
or OR3 (N96, N94, N71, N59);
nand NAND3 (N97, N92, N88, N43);
and AND3 (N98, N19, N69, N5);
or OR4 (N99, N67, N66, N47, N23);
xor XOR2 (N100, N96, N59);
nor NOR3 (N101, N98, N52, N52);
and AND2 (N102, N99, N8);
and AND4 (N103, N75, N7, N40, N14);
xor XOR2 (N104, N76, N75);
and AND2 (N105, N97, N83);
and AND2 (N106, N105, N89);
nand NAND2 (N107, N100, N58);
nor NOR3 (N108, N90, N59, N65);
nor NOR2 (N109, N72, N6);
and AND4 (N110, N95, N65, N85, N86);
nor NOR2 (N111, N104, N103);
xor XOR2 (N112, N48, N85);
and AND2 (N113, N106, N67);
not NOT1 (N114, N112);
nor NOR3 (N115, N110, N68, N91);
not NOT1 (N116, N114);
xor XOR2 (N117, N109, N51);
or OR2 (N118, N115, N34);
not NOT1 (N119, N93);
and AND3 (N120, N108, N114, N82);
not NOT1 (N121, N118);
nor NOR4 (N122, N121, N70, N121, N76);
not NOT1 (N123, N116);
not NOT1 (N124, N119);
nand NAND4 (N125, N113, N88, N63, N33);
nand NAND2 (N126, N117, N83);
buf BUF1 (N127, N122);
xor XOR2 (N128, N126, N9);
buf BUF1 (N129, N123);
nor NOR3 (N130, N125, N105, N101);
nor NOR3 (N131, N16, N68, N20);
buf BUF1 (N132, N130);
nand NAND4 (N133, N107, N65, N24, N5);
nand NAND4 (N134, N120, N34, N127, N69);
buf BUF1 (N135, N113);
nand NAND3 (N136, N102, N117, N87);
xor XOR2 (N137, N129, N67);
nand NAND3 (N138, N131, N102, N95);
nor NOR3 (N139, N134, N28, N122);
nand NAND4 (N140, N111, N31, N79, N55);
buf BUF1 (N141, N138);
nor NOR2 (N142, N132, N61);
nand NAND3 (N143, N141, N4, N110);
nor NOR2 (N144, N137, N83);
or OR4 (N145, N133, N55, N38, N134);
nor NOR4 (N146, N145, N4, N82, N12);
not NOT1 (N147, N128);
buf BUF1 (N148, N124);
or OR2 (N149, N143, N33);
or OR2 (N150, N149, N112);
or OR3 (N151, N135, N144, N149);
and AND3 (N152, N143, N34, N4);
or OR4 (N153, N139, N73, N72, N97);
nand NAND3 (N154, N146, N27, N135);
nand NAND3 (N155, N152, N48, N144);
not NOT1 (N156, N154);
and AND4 (N157, N147, N122, N130, N1);
buf BUF1 (N158, N136);
buf BUF1 (N159, N150);
nand NAND2 (N160, N155, N140);
nand NAND3 (N161, N22, N69, N42);
nor NOR4 (N162, N151, N52, N30, N95);
nor NOR3 (N163, N156, N33, N135);
xor XOR2 (N164, N159, N140);
not NOT1 (N165, N161);
or OR2 (N166, N148, N78);
not NOT1 (N167, N164);
buf BUF1 (N168, N158);
buf BUF1 (N169, N166);
buf BUF1 (N170, N142);
xor XOR2 (N171, N160, N35);
xor XOR2 (N172, N163, N119);
and AND2 (N173, N171, N22);
nand NAND3 (N174, N172, N5, N116);
and AND3 (N175, N173, N72, N8);
xor XOR2 (N176, N167, N39);
and AND4 (N177, N169, N149, N106, N141);
nand NAND3 (N178, N177, N61, N126);
not NOT1 (N179, N176);
nor NOR3 (N180, N162, N35, N48);
xor XOR2 (N181, N168, N80);
and AND2 (N182, N165, N113);
and AND4 (N183, N170, N60, N52, N48);
and AND2 (N184, N174, N152);
nor NOR3 (N185, N175, N57, N156);
or OR3 (N186, N182, N101, N91);
nand NAND2 (N187, N157, N53);
and AND3 (N188, N185, N76, N109);
not NOT1 (N189, N153);
or OR4 (N190, N188, N147, N27, N90);
nor NOR3 (N191, N181, N97, N64);
xor XOR2 (N192, N178, N117);
and AND2 (N193, N180, N107);
not NOT1 (N194, N190);
not NOT1 (N195, N189);
xor XOR2 (N196, N193, N105);
xor XOR2 (N197, N192, N176);
and AND2 (N198, N179, N191);
not NOT1 (N199, N112);
nor NOR2 (N200, N194, N50);
not NOT1 (N201, N197);
or OR2 (N202, N184, N121);
xor XOR2 (N203, N195, N106);
buf BUF1 (N204, N198);
and AND3 (N205, N187, N29, N78);
nand NAND4 (N206, N205, N181, N135, N153);
nand NAND4 (N207, N200, N89, N134, N5);
and AND3 (N208, N204, N104, N193);
buf BUF1 (N209, N202);
xor XOR2 (N210, N201, N137);
not NOT1 (N211, N196);
nand NAND4 (N212, N209, N205, N32, N46);
nand NAND3 (N213, N199, N87, N163);
buf BUF1 (N214, N213);
xor XOR2 (N215, N207, N108);
not NOT1 (N216, N214);
and AND3 (N217, N216, N77, N156);
or OR4 (N218, N203, N203, N167, N216);
nand NAND4 (N219, N210, N215, N92, N36);
nand NAND4 (N220, N212, N188, N80, N139);
and AND3 (N221, N214, N55, N30);
nor NOR3 (N222, N217, N105, N132);
or OR4 (N223, N222, N17, N210, N152);
and AND2 (N224, N220, N74);
xor XOR2 (N225, N186, N174);
buf BUF1 (N226, N219);
nor NOR2 (N227, N218, N32);
nand NAND2 (N228, N226, N40);
xor XOR2 (N229, N224, N56);
and AND2 (N230, N225, N138);
buf BUF1 (N231, N183);
and AND3 (N232, N206, N158, N211);
nor NOR2 (N233, N62, N56);
nor NOR4 (N234, N227, N41, N86, N95);
nand NAND2 (N235, N208, N202);
and AND3 (N236, N233, N60, N68);
and AND2 (N237, N235, N188);
or OR3 (N238, N232, N132, N85);
nor NOR3 (N239, N236, N29, N11);
buf BUF1 (N240, N239);
not NOT1 (N241, N240);
nand NAND3 (N242, N234, N34, N37);
not NOT1 (N243, N228);
nor NOR4 (N244, N231, N165, N228, N110);
or OR2 (N245, N241, N58);
not NOT1 (N246, N238);
nor NOR3 (N247, N245, N135, N42);
buf BUF1 (N248, N223);
and AND2 (N249, N242, N123);
buf BUF1 (N250, N248);
xor XOR2 (N251, N250, N88);
not NOT1 (N252, N247);
or OR4 (N253, N237, N92, N176, N81);
or OR4 (N254, N246, N139, N250, N253);
and AND4 (N255, N24, N166, N136, N90);
xor XOR2 (N256, N221, N228);
nor NOR4 (N257, N249, N66, N2, N239);
xor XOR2 (N258, N256, N230);
or OR4 (N259, N134, N121, N156, N123);
nor NOR2 (N260, N251, N214);
buf BUF1 (N261, N243);
nand NAND3 (N262, N260, N148, N250);
not NOT1 (N263, N229);
not NOT1 (N264, N257);
xor XOR2 (N265, N263, N163);
buf BUF1 (N266, N252);
nand NAND2 (N267, N255, N266);
not NOT1 (N268, N200);
buf BUF1 (N269, N267);
nand NAND2 (N270, N265, N94);
nand NAND2 (N271, N262, N249);
nor NOR2 (N272, N254, N71);
and AND2 (N273, N269, N118);
nor NOR3 (N274, N261, N77, N74);
not NOT1 (N275, N264);
not NOT1 (N276, N275);
not NOT1 (N277, N244);
not NOT1 (N278, N272);
nor NOR4 (N279, N276, N270, N110, N22);
nor NOR3 (N280, N213, N76, N254);
not NOT1 (N281, N274);
xor XOR2 (N282, N280, N75);
buf BUF1 (N283, N279);
or OR3 (N284, N268, N167, N73);
buf BUF1 (N285, N278);
nor NOR4 (N286, N281, N149, N96, N89);
and AND2 (N287, N283, N71);
nor NOR3 (N288, N284, N194, N78);
nand NAND2 (N289, N282, N225);
xor XOR2 (N290, N289, N180);
nor NOR3 (N291, N259, N234, N139);
xor XOR2 (N292, N271, N253);
nor NOR2 (N293, N292, N150);
not NOT1 (N294, N293);
and AND4 (N295, N273, N162, N61, N229);
nand NAND4 (N296, N277, N228, N169, N51);
or OR2 (N297, N290, N105);
or OR4 (N298, N285, N294, N89, N49);
nor NOR4 (N299, N76, N289, N11, N173);
xor XOR2 (N300, N297, N141);
and AND4 (N301, N286, N252, N34, N193);
xor XOR2 (N302, N300, N228);
not NOT1 (N303, N298);
xor XOR2 (N304, N303, N13);
and AND3 (N305, N258, N89, N189);
nand NAND4 (N306, N291, N161, N226, N239);
xor XOR2 (N307, N288, N11);
or OR3 (N308, N301, N5, N164);
nor NOR4 (N309, N304, N9, N269, N3);
nand NAND3 (N310, N299, N291, N29);
xor XOR2 (N311, N287, N143);
nor NOR3 (N312, N307, N42, N37);
nor NOR4 (N313, N311, N219, N125, N35);
not NOT1 (N314, N310);
buf BUF1 (N315, N308);
buf BUF1 (N316, N295);
nand NAND3 (N317, N312, N27, N187);
or OR2 (N318, N306, N143);
nand NAND2 (N319, N317, N11);
and AND2 (N320, N302, N271);
buf BUF1 (N321, N296);
or OR2 (N322, N305, N213);
not NOT1 (N323, N321);
not NOT1 (N324, N322);
and AND4 (N325, N323, N33, N311, N255);
and AND3 (N326, N316, N105, N116);
nor NOR2 (N327, N318, N267);
not NOT1 (N328, N320);
xor XOR2 (N329, N313, N48);
nand NAND3 (N330, N324, N232, N97);
or OR4 (N331, N329, N229, N218, N21);
and AND4 (N332, N314, N44, N167, N42);
not NOT1 (N333, N327);
buf BUF1 (N334, N315);
nor NOR3 (N335, N333, N163, N1);
nand NAND4 (N336, N309, N45, N296, N142);
nor NOR4 (N337, N331, N155, N95, N270);
xor XOR2 (N338, N337, N236);
and AND3 (N339, N335, N70, N293);
and AND4 (N340, N319, N285, N269, N205);
nand NAND2 (N341, N328, N294);
and AND2 (N342, N341, N108);
or OR2 (N343, N330, N280);
nand NAND3 (N344, N332, N196, N328);
xor XOR2 (N345, N339, N251);
or OR3 (N346, N336, N126, N242);
or OR2 (N347, N343, N214);
nand NAND3 (N348, N325, N344, N1);
xor XOR2 (N349, N42, N245);
not NOT1 (N350, N326);
nand NAND3 (N351, N350, N128, N126);
or OR4 (N352, N347, N31, N144, N16);
nand NAND4 (N353, N342, N27, N209, N155);
nand NAND3 (N354, N349, N257, N144);
nand NAND3 (N355, N348, N14, N22);
nor NOR3 (N356, N354, N305, N266);
xor XOR2 (N357, N338, N224);
not NOT1 (N358, N352);
or OR3 (N359, N353, N160, N307);
buf BUF1 (N360, N358);
nand NAND2 (N361, N360, N102);
buf BUF1 (N362, N359);
buf BUF1 (N363, N351);
not NOT1 (N364, N363);
buf BUF1 (N365, N340);
xor XOR2 (N366, N361, N243);
nand NAND2 (N367, N356, N261);
buf BUF1 (N368, N346);
and AND2 (N369, N357, N271);
nand NAND4 (N370, N366, N137, N202, N276);
xor XOR2 (N371, N362, N24);
buf BUF1 (N372, N355);
buf BUF1 (N373, N368);
and AND4 (N374, N365, N194, N208, N197);
nor NOR4 (N375, N345, N221, N176, N365);
nor NOR4 (N376, N375, N229, N232, N50);
nand NAND2 (N377, N373, N224);
xor XOR2 (N378, N364, N313);
nor NOR4 (N379, N377, N109, N301, N216);
buf BUF1 (N380, N370);
nor NOR4 (N381, N378, N70, N147, N296);
and AND2 (N382, N374, N250);
nand NAND4 (N383, N334, N218, N257, N281);
nor NOR2 (N384, N381, N157);
or OR2 (N385, N383, N59);
and AND3 (N386, N372, N165, N311);
and AND3 (N387, N380, N222, N158);
nor NOR2 (N388, N376, N7);
nand NAND2 (N389, N386, N365);
xor XOR2 (N390, N367, N367);
or OR2 (N391, N379, N338);
nor NOR4 (N392, N384, N376, N144, N52);
nor NOR3 (N393, N382, N290, N33);
nand NAND3 (N394, N388, N237, N67);
xor XOR2 (N395, N389, N95);
nor NOR2 (N396, N371, N53);
xor XOR2 (N397, N390, N186);
xor XOR2 (N398, N392, N28);
or OR4 (N399, N395, N225, N289, N127);
buf BUF1 (N400, N396);
and AND3 (N401, N387, N369, N297);
not NOT1 (N402, N230);
xor XOR2 (N403, N402, N178);
not NOT1 (N404, N403);
xor XOR2 (N405, N391, N361);
nand NAND4 (N406, N394, N316, N299, N29);
buf BUF1 (N407, N405);
nor NOR3 (N408, N407, N371, N143);
buf BUF1 (N409, N398);
not NOT1 (N410, N409);
and AND2 (N411, N406, N278);
nand NAND4 (N412, N401, N327, N373, N188);
nand NAND4 (N413, N410, N260, N219, N30);
not NOT1 (N414, N408);
nor NOR4 (N415, N414, N58, N83, N212);
or OR2 (N416, N404, N23);
nand NAND3 (N417, N397, N246, N101);
xor XOR2 (N418, N385, N415);
nor NOR4 (N419, N416, N274, N22, N65);
buf BUF1 (N420, N224);
xor XOR2 (N421, N411, N367);
or OR4 (N422, N400, N241, N223, N182);
and AND3 (N423, N399, N355, N415);
or OR3 (N424, N419, N157, N256);
nand NAND2 (N425, N420, N75);
xor XOR2 (N426, N418, N183);
and AND4 (N427, N421, N67, N125, N314);
and AND4 (N428, N426, N403, N80, N209);
and AND4 (N429, N417, N273, N409, N149);
buf BUF1 (N430, N425);
xor XOR2 (N431, N427, N359);
buf BUF1 (N432, N393);
not NOT1 (N433, N432);
and AND2 (N434, N433, N381);
and AND2 (N435, N428, N381);
not NOT1 (N436, N430);
xor XOR2 (N437, N436, N254);
buf BUF1 (N438, N437);
xor XOR2 (N439, N438, N95);
and AND2 (N440, N439, N428);
not NOT1 (N441, N412);
and AND2 (N442, N431, N122);
xor XOR2 (N443, N440, N46);
buf BUF1 (N444, N424);
and AND3 (N445, N443, N426, N416);
xor XOR2 (N446, N441, N103);
nor NOR4 (N447, N423, N342, N151, N231);
and AND3 (N448, N445, N288, N203);
not NOT1 (N449, N429);
xor XOR2 (N450, N434, N441);
or OR3 (N451, N447, N102, N170);
nor NOR4 (N452, N422, N438, N121, N281);
and AND2 (N453, N444, N224);
nor NOR4 (N454, N413, N194, N369, N412);
nor NOR4 (N455, N452, N183, N35, N388);
nor NOR2 (N456, N435, N293);
and AND3 (N457, N453, N331, N439);
nand NAND4 (N458, N448, N35, N152, N182);
and AND3 (N459, N446, N150, N206);
buf BUF1 (N460, N456);
and AND2 (N461, N442, N116);
and AND4 (N462, N461, N221, N277, N109);
or OR2 (N463, N462, N204);
buf BUF1 (N464, N458);
xor XOR2 (N465, N463, N307);
nor NOR3 (N466, N450, N411, N82);
nand NAND3 (N467, N460, N215, N69);
or OR4 (N468, N454, N341, N340, N14);
nand NAND4 (N469, N467, N331, N412, N371);
nand NAND4 (N470, N468, N97, N327, N129);
xor XOR2 (N471, N464, N179);
nor NOR3 (N472, N471, N327, N274);
or OR3 (N473, N457, N139, N212);
nand NAND2 (N474, N451, N448);
not NOT1 (N475, N472);
nor NOR2 (N476, N466, N137);
xor XOR2 (N477, N476, N333);
not NOT1 (N478, N470);
or OR4 (N479, N465, N42, N377, N307);
nand NAND2 (N480, N478, N222);
xor XOR2 (N481, N479, N136);
xor XOR2 (N482, N475, N129);
nand NAND2 (N483, N473, N417);
not NOT1 (N484, N480);
nor NOR4 (N485, N484, N177, N188, N156);
not NOT1 (N486, N449);
nand NAND2 (N487, N481, N18);
buf BUF1 (N488, N469);
nand NAND4 (N489, N455, N184, N404, N349);
nand NAND4 (N490, N486, N236, N488, N100);
and AND3 (N491, N389, N310, N202);
buf BUF1 (N492, N483);
nor NOR4 (N493, N459, N32, N137, N265);
nor NOR2 (N494, N487, N262);
nor NOR2 (N495, N489, N440);
xor XOR2 (N496, N494, N339);
buf BUF1 (N497, N482);
xor XOR2 (N498, N485, N375);
buf BUF1 (N499, N498);
or OR4 (N500, N491, N334, N462, N305);
nand NAND2 (N501, N477, N405);
buf BUF1 (N502, N492);
and AND2 (N503, N499, N208);
xor XOR2 (N504, N501, N59);
and AND3 (N505, N497, N469, N280);
not NOT1 (N506, N495);
or OR2 (N507, N504, N434);
and AND4 (N508, N507, N59, N262, N324);
xor XOR2 (N509, N500, N212);
xor XOR2 (N510, N503, N208);
and AND3 (N511, N505, N202, N98);
and AND4 (N512, N496, N432, N316, N471);
buf BUF1 (N513, N474);
or OR2 (N514, N490, N12);
buf BUF1 (N515, N493);
not NOT1 (N516, N511);
xor XOR2 (N517, N512, N374);
nor NOR3 (N518, N508, N354, N306);
buf BUF1 (N519, N502);
xor XOR2 (N520, N518, N440);
buf BUF1 (N521, N509);
nor NOR3 (N522, N515, N345, N365);
and AND4 (N523, N506, N97, N494, N82);
nand NAND3 (N524, N519, N202, N455);
nand NAND2 (N525, N517, N460);
and AND2 (N526, N525, N119);
xor XOR2 (N527, N510, N253);
or OR4 (N528, N513, N42, N161, N59);
buf BUF1 (N529, N514);
not NOT1 (N530, N524);
and AND3 (N531, N527, N12, N363);
not NOT1 (N532, N529);
nand NAND3 (N533, N528, N304, N140);
xor XOR2 (N534, N526, N529);
buf BUF1 (N535, N531);
and AND3 (N536, N520, N503, N72);
xor XOR2 (N537, N521, N67);
not NOT1 (N538, N533);
nor NOR4 (N539, N534, N363, N76, N108);
xor XOR2 (N540, N537, N39);
nand NAND4 (N541, N539, N10, N199, N33);
buf BUF1 (N542, N540);
buf BUF1 (N543, N538);
nand NAND3 (N544, N522, N280, N173);
nand NAND3 (N545, N523, N454, N409);
buf BUF1 (N546, N532);
nor NOR2 (N547, N543, N356);
nor NOR3 (N548, N535, N275, N303);
nor NOR4 (N549, N547, N499, N105, N175);
xor XOR2 (N550, N516, N294);
nand NAND3 (N551, N536, N349, N376);
and AND2 (N552, N548, N135);
nor NOR3 (N553, N541, N387, N101);
or OR2 (N554, N553, N275);
not NOT1 (N555, N552);
buf BUF1 (N556, N545);
not NOT1 (N557, N544);
nor NOR3 (N558, N550, N413, N159);
or OR4 (N559, N556, N295, N289, N220);
nor NOR3 (N560, N542, N447, N350);
buf BUF1 (N561, N530);
and AND2 (N562, N554, N316);
or OR3 (N563, N562, N64, N186);
buf BUF1 (N564, N555);
xor XOR2 (N565, N563, N74);
or OR2 (N566, N549, N406);
nand NAND2 (N567, N558, N383);
nand NAND2 (N568, N565, N562);
buf BUF1 (N569, N546);
nand NAND2 (N570, N564, N105);
and AND3 (N571, N566, N145, N346);
or OR4 (N572, N561, N505, N495, N531);
nor NOR3 (N573, N557, N205, N218);
nand NAND3 (N574, N567, N349, N176);
buf BUF1 (N575, N574);
nand NAND3 (N576, N560, N200, N75);
not NOT1 (N577, N569);
or OR4 (N578, N568, N68, N217, N256);
nor NOR4 (N579, N576, N68, N373, N569);
not NOT1 (N580, N571);
not NOT1 (N581, N579);
xor XOR2 (N582, N581, N426);
nand NAND2 (N583, N580, N325);
nor NOR2 (N584, N573, N360);
nand NAND4 (N585, N559, N52, N409, N494);
and AND4 (N586, N578, N439, N170, N171);
and AND4 (N587, N551, N28, N296, N245);
or OR4 (N588, N583, N384, N53, N378);
nor NOR2 (N589, N577, N125);
buf BUF1 (N590, N575);
and AND3 (N591, N572, N78, N195);
nand NAND4 (N592, N591, N187, N330, N113);
or OR3 (N593, N582, N327, N3);
not NOT1 (N594, N589);
and AND2 (N595, N586, N353);
nor NOR4 (N596, N593, N208, N271, N285);
nand NAND3 (N597, N595, N29, N429);
nand NAND4 (N598, N597, N595, N589, N125);
nand NAND4 (N599, N594, N318, N310, N491);
and AND3 (N600, N599, N247, N86);
xor XOR2 (N601, N584, N149);
xor XOR2 (N602, N590, N530);
nand NAND2 (N603, N602, N314);
buf BUF1 (N604, N600);
xor XOR2 (N605, N592, N540);
xor XOR2 (N606, N588, N167);
xor XOR2 (N607, N606, N59);
or OR2 (N608, N605, N581);
buf BUF1 (N609, N604);
nor NOR4 (N610, N585, N463, N59, N128);
buf BUF1 (N611, N603);
or OR2 (N612, N596, N421);
nand NAND3 (N613, N607, N35, N45);
not NOT1 (N614, N613);
not NOT1 (N615, N608);
buf BUF1 (N616, N611);
xor XOR2 (N617, N612, N493);
not NOT1 (N618, N598);
xor XOR2 (N619, N616, N151);
or OR4 (N620, N619, N102, N134, N272);
and AND2 (N621, N587, N614);
not NOT1 (N622, N165);
xor XOR2 (N623, N615, N147);
xor XOR2 (N624, N618, N158);
buf BUF1 (N625, N623);
not NOT1 (N626, N609);
and AND2 (N627, N625, N424);
or OR2 (N628, N601, N515);
xor XOR2 (N629, N624, N489);
buf BUF1 (N630, N629);
nand NAND3 (N631, N622, N342, N186);
nand NAND3 (N632, N630, N186, N436);
nand NAND4 (N633, N632, N507, N437, N175);
and AND2 (N634, N628, N98);
nand NAND2 (N635, N631, N103);
not NOT1 (N636, N627);
not NOT1 (N637, N633);
xor XOR2 (N638, N621, N209);
xor XOR2 (N639, N634, N352);
nand NAND3 (N640, N636, N18, N141);
or OR3 (N641, N637, N127, N240);
or OR3 (N642, N620, N496, N295);
or OR4 (N643, N639, N226, N509, N247);
not NOT1 (N644, N617);
nand NAND2 (N645, N570, N394);
xor XOR2 (N646, N644, N593);
and AND2 (N647, N635, N56);
buf BUF1 (N648, N646);
nand NAND3 (N649, N641, N99, N467);
or OR3 (N650, N610, N573, N342);
nand NAND3 (N651, N650, N194, N496);
or OR2 (N652, N626, N167);
xor XOR2 (N653, N647, N66);
xor XOR2 (N654, N643, N243);
xor XOR2 (N655, N654, N347);
xor XOR2 (N656, N645, N61);
nor NOR4 (N657, N656, N432, N63, N553);
not NOT1 (N658, N655);
nor NOR3 (N659, N638, N38, N405);
and AND3 (N660, N653, N282, N411);
xor XOR2 (N661, N648, N253);
nand NAND3 (N662, N657, N382, N411);
nand NAND4 (N663, N661, N197, N229, N501);
or OR2 (N664, N642, N372);
nand NAND4 (N665, N658, N393, N119, N346);
not NOT1 (N666, N652);
nand NAND4 (N667, N666, N125, N526, N277);
and AND3 (N668, N651, N68, N556);
not NOT1 (N669, N665);
nand NAND2 (N670, N640, N590);
and AND4 (N671, N668, N85, N498, N255);
not NOT1 (N672, N669);
xor XOR2 (N673, N663, N668);
and AND4 (N674, N659, N435, N8, N465);
or OR4 (N675, N664, N258, N564, N516);
nand NAND4 (N676, N675, N380, N324, N648);
and AND2 (N677, N673, N129);
and AND2 (N678, N676, N302);
xor XOR2 (N679, N671, N19);
nor NOR3 (N680, N672, N575, N484);
buf BUF1 (N681, N677);
nand NAND4 (N682, N679, N121, N255, N595);
not NOT1 (N683, N649);
xor XOR2 (N684, N660, N585);
or OR2 (N685, N681, N309);
and AND2 (N686, N685, N17);
and AND4 (N687, N674, N98, N295, N329);
not NOT1 (N688, N682);
xor XOR2 (N689, N680, N648);
nand NAND4 (N690, N684, N328, N25, N224);
or OR3 (N691, N686, N585, N200);
nand NAND2 (N692, N678, N315);
nor NOR4 (N693, N688, N342, N79, N125);
buf BUF1 (N694, N690);
nand NAND2 (N695, N691, N195);
not NOT1 (N696, N687);
nand NAND4 (N697, N683, N331, N34, N439);
buf BUF1 (N698, N693);
or OR2 (N699, N689, N586);
not NOT1 (N700, N696);
not NOT1 (N701, N667);
nor NOR3 (N702, N699, N406, N623);
xor XOR2 (N703, N694, N197);
nand NAND4 (N704, N700, N641, N2, N250);
nor NOR3 (N705, N662, N142, N195);
and AND2 (N706, N703, N284);
and AND3 (N707, N704, N9, N9);
and AND4 (N708, N695, N316, N106, N611);
and AND4 (N709, N697, N257, N247, N230);
and AND2 (N710, N702, N234);
nand NAND3 (N711, N706, N555, N185);
not NOT1 (N712, N705);
nor NOR4 (N713, N709, N659, N258, N708);
nand NAND4 (N714, N295, N662, N628, N218);
and AND2 (N715, N707, N373);
nand NAND4 (N716, N670, N25, N226, N242);
and AND2 (N717, N701, N167);
not NOT1 (N718, N712);
xor XOR2 (N719, N717, N420);
and AND3 (N720, N710, N33, N219);
and AND2 (N721, N716, N122);
nand NAND4 (N722, N719, N701, N238, N22);
xor XOR2 (N723, N698, N316);
nand NAND4 (N724, N711, N462, N20, N538);
not NOT1 (N725, N722);
xor XOR2 (N726, N713, N592);
nand NAND3 (N727, N692, N509, N547);
or OR2 (N728, N726, N311);
not NOT1 (N729, N718);
buf BUF1 (N730, N715);
and AND3 (N731, N729, N269, N611);
buf BUF1 (N732, N728);
not NOT1 (N733, N727);
not NOT1 (N734, N724);
not NOT1 (N735, N720);
xor XOR2 (N736, N714, N387);
not NOT1 (N737, N730);
and AND3 (N738, N734, N192, N245);
xor XOR2 (N739, N723, N534);
buf BUF1 (N740, N737);
nor NOR2 (N741, N732, N276);
nor NOR2 (N742, N721, N415);
nand NAND4 (N743, N741, N546, N51, N120);
not NOT1 (N744, N731);
xor XOR2 (N745, N740, N45);
or OR4 (N746, N744, N547, N360, N261);
xor XOR2 (N747, N733, N550);
nand NAND2 (N748, N742, N8);
nand NAND3 (N749, N725, N241, N457);
nand NAND2 (N750, N736, N533);
nand NAND2 (N751, N746, N444);
not NOT1 (N752, N738);
or OR3 (N753, N752, N241, N360);
or OR4 (N754, N748, N407, N706, N724);
not NOT1 (N755, N743);
nor NOR4 (N756, N755, N705, N441, N402);
buf BUF1 (N757, N747);
xor XOR2 (N758, N757, N308);
buf BUF1 (N759, N735);
nand NAND2 (N760, N749, N95);
buf BUF1 (N761, N753);
and AND3 (N762, N751, N295, N761);
or OR2 (N763, N446, N217);
not NOT1 (N764, N760);
buf BUF1 (N765, N759);
nand NAND2 (N766, N745, N487);
xor XOR2 (N767, N739, N95);
xor XOR2 (N768, N754, N329);
nor NOR3 (N769, N764, N4, N257);
and AND3 (N770, N767, N545, N378);
and AND4 (N771, N750, N269, N573, N129);
nand NAND4 (N772, N768, N137, N428, N651);
nor NOR4 (N773, N765, N179, N105, N485);
xor XOR2 (N774, N766, N312);
nand NAND3 (N775, N774, N347, N690);
nand NAND2 (N776, N756, N525);
or OR4 (N777, N772, N437, N249, N452);
not NOT1 (N778, N770);
nor NOR3 (N779, N776, N681, N557);
nor NOR2 (N780, N773, N24);
nand NAND2 (N781, N762, N340);
nand NAND2 (N782, N771, N258);
buf BUF1 (N783, N763);
buf BUF1 (N784, N781);
xor XOR2 (N785, N783, N153);
or OR2 (N786, N769, N681);
and AND3 (N787, N775, N212, N518);
xor XOR2 (N788, N784, N66);
xor XOR2 (N789, N785, N150);
buf BUF1 (N790, N789);
nor NOR3 (N791, N786, N719, N275);
nand NAND2 (N792, N780, N380);
or OR3 (N793, N758, N189, N11);
xor XOR2 (N794, N791, N635);
nor NOR3 (N795, N793, N429, N599);
not NOT1 (N796, N787);
nand NAND4 (N797, N795, N336, N676, N168);
or OR3 (N798, N777, N570, N578);
not NOT1 (N799, N792);
xor XOR2 (N800, N794, N316);
nor NOR4 (N801, N790, N90, N581, N667);
or OR2 (N802, N778, N798);
and AND3 (N803, N350, N204, N645);
buf BUF1 (N804, N799);
and AND2 (N805, N797, N37);
and AND2 (N806, N779, N697);
nand NAND3 (N807, N788, N686, N359);
and AND2 (N808, N800, N556);
not NOT1 (N809, N807);
or OR4 (N810, N803, N527, N745, N757);
buf BUF1 (N811, N809);
not NOT1 (N812, N808);
buf BUF1 (N813, N810);
nand NAND2 (N814, N802, N757);
xor XOR2 (N815, N806, N62);
or OR3 (N816, N805, N220, N750);
buf BUF1 (N817, N801);
and AND2 (N818, N804, N687);
xor XOR2 (N819, N813, N344);
nand NAND3 (N820, N811, N548, N442);
nand NAND2 (N821, N815, N443);
xor XOR2 (N822, N820, N806);
and AND2 (N823, N816, N76);
nor NOR2 (N824, N812, N88);
not NOT1 (N825, N817);
nor NOR3 (N826, N782, N490, N222);
not NOT1 (N827, N814);
nand NAND2 (N828, N825, N47);
xor XOR2 (N829, N827, N548);
nor NOR4 (N830, N829, N470, N538, N187);
or OR3 (N831, N796, N494, N494);
buf BUF1 (N832, N830);
not NOT1 (N833, N824);
xor XOR2 (N834, N821, N534);
xor XOR2 (N835, N833, N161);
or OR2 (N836, N819, N677);
and AND2 (N837, N822, N671);
buf BUF1 (N838, N835);
or OR3 (N839, N832, N310, N421);
and AND3 (N840, N826, N522, N499);
and AND4 (N841, N840, N188, N285, N41);
xor XOR2 (N842, N837, N694);
buf BUF1 (N843, N838);
or OR4 (N844, N842, N410, N121, N832);
xor XOR2 (N845, N818, N39);
buf BUF1 (N846, N845);
not NOT1 (N847, N843);
and AND3 (N848, N841, N526, N89);
and AND3 (N849, N846, N78, N296);
buf BUF1 (N850, N848);
and AND3 (N851, N847, N37, N619);
and AND2 (N852, N851, N106);
not NOT1 (N853, N849);
buf BUF1 (N854, N834);
buf BUF1 (N855, N831);
not NOT1 (N856, N836);
not NOT1 (N857, N850);
nor NOR2 (N858, N852, N506);
and AND4 (N859, N823, N257, N663, N590);
nand NAND2 (N860, N844, N214);
nor NOR4 (N861, N858, N85, N174, N367);
nand NAND2 (N862, N839, N35);
nor NOR4 (N863, N853, N134, N490, N10);
xor XOR2 (N864, N854, N58);
buf BUF1 (N865, N857);
nor NOR4 (N866, N865, N758, N74, N128);
xor XOR2 (N867, N859, N752);
or OR2 (N868, N855, N503);
or OR2 (N869, N861, N521);
nand NAND2 (N870, N860, N318);
buf BUF1 (N871, N828);
or OR4 (N872, N856, N747, N61, N661);
and AND4 (N873, N862, N445, N223, N869);
and AND4 (N874, N679, N73, N446, N729);
nand NAND4 (N875, N872, N760, N773, N46);
or OR2 (N876, N875, N578);
xor XOR2 (N877, N866, N518);
and AND4 (N878, N867, N650, N869, N132);
or OR4 (N879, N863, N582, N408, N810);
xor XOR2 (N880, N873, N553);
or OR2 (N881, N879, N307);
not NOT1 (N882, N878);
nand NAND4 (N883, N880, N606, N13, N745);
not NOT1 (N884, N874);
nand NAND4 (N885, N877, N187, N208, N401);
not NOT1 (N886, N884);
or OR4 (N887, N883, N375, N134, N533);
xor XOR2 (N888, N864, N519);
not NOT1 (N889, N887);
xor XOR2 (N890, N871, N653);
not NOT1 (N891, N868);
nor NOR2 (N892, N886, N779);
xor XOR2 (N893, N890, N457);
nand NAND3 (N894, N881, N789, N716);
not NOT1 (N895, N891);
not NOT1 (N896, N889);
buf BUF1 (N897, N870);
xor XOR2 (N898, N882, N495);
nor NOR3 (N899, N898, N841, N836);
xor XOR2 (N900, N893, N445);
not NOT1 (N901, N897);
xor XOR2 (N902, N896, N756);
xor XOR2 (N903, N876, N400);
nand NAND4 (N904, N900, N363, N713, N432);
xor XOR2 (N905, N899, N571);
or OR2 (N906, N904, N730);
and AND3 (N907, N892, N76, N231);
and AND4 (N908, N895, N891, N645, N75);
and AND4 (N909, N907, N486, N845, N224);
nor NOR3 (N910, N885, N489, N485);
and AND4 (N911, N905, N381, N276, N57);
or OR2 (N912, N910, N631);
and AND2 (N913, N908, N476);
endmodule