// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N597,N618,N613,N606,N612,N607,N617,N615,N619,N620;

buf BUF1 (N21, N18);
and AND2 (N22, N16, N12);
nand NAND4 (N23, N14, N6, N18, N1);
not NOT1 (N24, N8);
nor NOR3 (N25, N8, N24, N19);
not NOT1 (N26, N8);
or OR2 (N27, N16, N20);
nand NAND3 (N28, N18, N10, N2);
buf BUF1 (N29, N6);
xor XOR2 (N30, N28, N1);
or OR3 (N31, N18, N29, N11);
nand NAND4 (N32, N26, N1, N5, N20);
and AND2 (N33, N1, N10);
not NOT1 (N34, N18);
buf BUF1 (N35, N31);
not NOT1 (N36, N25);
xor XOR2 (N37, N21, N35);
buf BUF1 (N38, N20);
buf BUF1 (N39, N36);
or OR2 (N40, N39, N26);
and AND3 (N41, N38, N26, N39);
nand NAND4 (N42, N23, N10, N27, N29);
and AND2 (N43, N1, N38);
and AND2 (N44, N34, N32);
nand NAND2 (N45, N2, N29);
xor XOR2 (N46, N37, N29);
not NOT1 (N47, N30);
and AND2 (N48, N33, N8);
or OR2 (N49, N48, N15);
buf BUF1 (N50, N45);
nand NAND3 (N51, N43, N10, N40);
xor XOR2 (N52, N37, N49);
and AND3 (N53, N38, N7, N18);
xor XOR2 (N54, N44, N16);
or OR2 (N55, N50, N36);
buf BUF1 (N56, N41);
buf BUF1 (N57, N46);
nor NOR2 (N58, N56, N4);
nand NAND2 (N59, N42, N55);
xor XOR2 (N60, N46, N57);
xor XOR2 (N61, N35, N45);
buf BUF1 (N62, N61);
or OR4 (N63, N62, N27, N18, N38);
nand NAND3 (N64, N59, N38, N18);
not NOT1 (N65, N64);
and AND4 (N66, N47, N23, N43, N39);
nand NAND3 (N67, N58, N35, N31);
nor NOR3 (N68, N52, N38, N46);
nor NOR3 (N69, N65, N46, N54);
nor NOR3 (N70, N23, N11, N65);
nand NAND2 (N71, N22, N1);
or OR4 (N72, N63, N4, N43, N69);
xor XOR2 (N73, N20, N63);
and AND3 (N74, N51, N4, N25);
buf BUF1 (N75, N72);
or OR3 (N76, N53, N3, N51);
xor XOR2 (N77, N68, N65);
or OR4 (N78, N70, N31, N38, N21);
or OR2 (N79, N75, N71);
nand NAND2 (N80, N10, N30);
nor NOR3 (N81, N66, N24, N51);
not NOT1 (N82, N80);
nand NAND4 (N83, N76, N44, N16, N13);
not NOT1 (N84, N74);
xor XOR2 (N85, N77, N68);
nand NAND4 (N86, N83, N4, N66, N66);
and AND2 (N87, N78, N9);
buf BUF1 (N88, N85);
and AND4 (N89, N60, N18, N6, N10);
nor NOR4 (N90, N89, N51, N76, N80);
and AND3 (N91, N81, N37, N29);
not NOT1 (N92, N90);
buf BUF1 (N93, N88);
and AND2 (N94, N79, N2);
xor XOR2 (N95, N94, N39);
buf BUF1 (N96, N82);
buf BUF1 (N97, N92);
xor XOR2 (N98, N96, N73);
buf BUF1 (N99, N24);
nand NAND2 (N100, N93, N77);
buf BUF1 (N101, N98);
and AND2 (N102, N86, N1);
nand NAND2 (N103, N67, N29);
buf BUF1 (N104, N87);
not NOT1 (N105, N101);
nor NOR3 (N106, N100, N37, N41);
buf BUF1 (N107, N105);
xor XOR2 (N108, N99, N36);
and AND2 (N109, N103, N104);
buf BUF1 (N110, N35);
xor XOR2 (N111, N110, N9);
and AND2 (N112, N102, N29);
xor XOR2 (N113, N108, N16);
or OR2 (N114, N107, N23);
and AND2 (N115, N97, N99);
nor NOR2 (N116, N113, N39);
buf BUF1 (N117, N114);
xor XOR2 (N118, N112, N59);
buf BUF1 (N119, N106);
xor XOR2 (N120, N111, N42);
and AND3 (N121, N120, N120, N33);
buf BUF1 (N122, N116);
buf BUF1 (N123, N95);
nor NOR2 (N124, N115, N94);
buf BUF1 (N125, N84);
nor NOR3 (N126, N118, N13, N63);
nand NAND2 (N127, N117, N58);
nand NAND2 (N128, N126, N105);
xor XOR2 (N129, N122, N64);
and AND3 (N130, N91, N56, N94);
nor NOR3 (N131, N129, N108, N18);
and AND3 (N132, N119, N55, N107);
buf BUF1 (N133, N130);
not NOT1 (N134, N127);
xor XOR2 (N135, N121, N79);
or OR3 (N136, N132, N21, N118);
buf BUF1 (N137, N134);
nand NAND4 (N138, N135, N113, N109, N55);
not NOT1 (N139, N91);
nor NOR4 (N140, N128, N97, N101, N16);
xor XOR2 (N141, N133, N128);
nand NAND2 (N142, N136, N118);
or OR3 (N143, N138, N105, N63);
and AND4 (N144, N131, N16, N32, N24);
not NOT1 (N145, N137);
nand NAND2 (N146, N145, N123);
not NOT1 (N147, N132);
buf BUF1 (N148, N139);
not NOT1 (N149, N144);
nor NOR4 (N150, N140, N126, N48, N10);
buf BUF1 (N151, N124);
nor NOR2 (N152, N150, N38);
buf BUF1 (N153, N148);
and AND2 (N154, N147, N137);
or OR2 (N155, N143, N17);
nor NOR2 (N156, N142, N81);
not NOT1 (N157, N125);
buf BUF1 (N158, N152);
nor NOR2 (N159, N158, N51);
not NOT1 (N160, N157);
nand NAND2 (N161, N151, N103);
nand NAND4 (N162, N160, N110, N41, N113);
xor XOR2 (N163, N153, N84);
buf BUF1 (N164, N154);
not NOT1 (N165, N155);
not NOT1 (N166, N159);
nor NOR3 (N167, N162, N29, N133);
or OR2 (N168, N146, N164);
not NOT1 (N169, N81);
and AND3 (N170, N166, N55, N17);
or OR4 (N171, N161, N96, N146, N40);
buf BUF1 (N172, N167);
and AND4 (N173, N171, N122, N65, N127);
nand NAND2 (N174, N149, N65);
xor XOR2 (N175, N173, N46);
not NOT1 (N176, N170);
or OR2 (N177, N176, N44);
or OR2 (N178, N177, N111);
not NOT1 (N179, N178);
nor NOR2 (N180, N174, N36);
nor NOR3 (N181, N163, N133, N154);
not NOT1 (N182, N180);
xor XOR2 (N183, N179, N160);
buf BUF1 (N184, N183);
buf BUF1 (N185, N168);
nor NOR4 (N186, N141, N4, N171, N29);
nor NOR3 (N187, N185, N92, N168);
buf BUF1 (N188, N181);
not NOT1 (N189, N188);
nor NOR2 (N190, N184, N121);
not NOT1 (N191, N190);
not NOT1 (N192, N165);
or OR3 (N193, N172, N122, N84);
not NOT1 (N194, N193);
buf BUF1 (N195, N169);
buf BUF1 (N196, N192);
xor XOR2 (N197, N175, N113);
nand NAND4 (N198, N182, N85, N4, N139);
nand NAND4 (N199, N189, N105, N90, N65);
not NOT1 (N200, N156);
and AND3 (N201, N195, N129, N118);
xor XOR2 (N202, N199, N70);
not NOT1 (N203, N194);
or OR2 (N204, N203, N42);
and AND4 (N205, N200, N61, N36, N202);
or OR4 (N206, N28, N53, N179, N49);
not NOT1 (N207, N201);
nand NAND3 (N208, N191, N115, N45);
or OR3 (N209, N187, N49, N134);
and AND2 (N210, N197, N93);
nand NAND4 (N211, N186, N138, N34, N125);
nand NAND3 (N212, N198, N80, N57);
not NOT1 (N213, N207);
nor NOR4 (N214, N213, N47, N78, N9);
buf BUF1 (N215, N205);
and AND2 (N216, N204, N198);
and AND4 (N217, N208, N110, N177, N203);
buf BUF1 (N218, N196);
nor NOR4 (N219, N212, N70, N179, N207);
buf BUF1 (N220, N215);
not NOT1 (N221, N214);
nand NAND3 (N222, N220, N18, N14);
and AND3 (N223, N206, N37, N22);
not NOT1 (N224, N218);
xor XOR2 (N225, N211, N70);
nor NOR3 (N226, N222, N88, N122);
or OR3 (N227, N217, N90, N86);
nor NOR2 (N228, N223, N177);
nor NOR4 (N229, N210, N147, N156, N33);
nand NAND2 (N230, N209, N56);
nor NOR4 (N231, N230, N101, N69, N135);
buf BUF1 (N232, N227);
not NOT1 (N233, N224);
buf BUF1 (N234, N233);
nor NOR2 (N235, N229, N52);
nor NOR4 (N236, N231, N110, N53, N122);
and AND3 (N237, N225, N68, N170);
not NOT1 (N238, N237);
and AND2 (N239, N238, N153);
not NOT1 (N240, N219);
not NOT1 (N241, N226);
not NOT1 (N242, N236);
not NOT1 (N243, N240);
and AND2 (N244, N228, N113);
buf BUF1 (N245, N232);
and AND4 (N246, N241, N197, N182, N220);
or OR2 (N247, N242, N123);
nor NOR4 (N248, N235, N84, N114, N92);
nand NAND3 (N249, N221, N212, N231);
and AND3 (N250, N243, N47, N130);
nor NOR3 (N251, N246, N110, N191);
or OR4 (N252, N249, N85, N51, N169);
nand NAND2 (N253, N216, N67);
and AND2 (N254, N245, N94);
nor NOR2 (N255, N248, N102);
nand NAND2 (N256, N244, N21);
nor NOR2 (N257, N254, N5);
not NOT1 (N258, N251);
not NOT1 (N259, N253);
buf BUF1 (N260, N247);
nand NAND3 (N261, N255, N78, N5);
or OR2 (N262, N257, N72);
xor XOR2 (N263, N239, N231);
not NOT1 (N264, N258);
nand NAND4 (N265, N234, N6, N25, N84);
not NOT1 (N266, N259);
nand NAND4 (N267, N263, N162, N261, N237);
xor XOR2 (N268, N91, N155);
buf BUF1 (N269, N266);
or OR2 (N270, N264, N24);
nand NAND2 (N271, N252, N108);
not NOT1 (N272, N269);
or OR3 (N273, N268, N102, N10);
nor NOR4 (N274, N265, N102, N203, N263);
and AND3 (N275, N262, N100, N237);
or OR2 (N276, N271, N211);
not NOT1 (N277, N276);
nand NAND2 (N278, N250, N3);
buf BUF1 (N279, N272);
and AND3 (N280, N279, N103, N14);
and AND4 (N281, N256, N181, N188, N210);
or OR2 (N282, N260, N32);
not NOT1 (N283, N275);
nand NAND2 (N284, N277, N79);
xor XOR2 (N285, N274, N91);
or OR4 (N286, N282, N256, N15, N280);
and AND4 (N287, N74, N73, N44, N246);
nor NOR4 (N288, N283, N8, N92, N284);
buf BUF1 (N289, N253);
not NOT1 (N290, N285);
and AND2 (N291, N281, N181);
or OR2 (N292, N286, N84);
nor NOR4 (N293, N267, N238, N263, N265);
not NOT1 (N294, N292);
and AND4 (N295, N288, N192, N158, N162);
xor XOR2 (N296, N278, N229);
nand NAND4 (N297, N273, N194, N83, N29);
or OR3 (N298, N270, N72, N99);
and AND4 (N299, N289, N73, N98, N230);
xor XOR2 (N300, N299, N242);
buf BUF1 (N301, N287);
or OR4 (N302, N296, N265, N214, N223);
nand NAND2 (N303, N301, N172);
buf BUF1 (N304, N295);
buf BUF1 (N305, N303);
or OR2 (N306, N304, N81);
xor XOR2 (N307, N302, N71);
nor NOR3 (N308, N305, N299, N106);
buf BUF1 (N309, N293);
or OR3 (N310, N309, N54, N205);
nor NOR4 (N311, N300, N254, N19, N173);
not NOT1 (N312, N308);
and AND2 (N313, N310, N19);
nand NAND2 (N314, N311, N276);
or OR2 (N315, N294, N132);
nor NOR2 (N316, N290, N170);
or OR2 (N317, N316, N98);
or OR2 (N318, N313, N10);
and AND2 (N319, N297, N36);
nand NAND4 (N320, N315, N53, N181, N1);
nor NOR3 (N321, N291, N132, N305);
buf BUF1 (N322, N321);
not NOT1 (N323, N314);
not NOT1 (N324, N322);
nor NOR2 (N325, N307, N241);
not NOT1 (N326, N320);
nor NOR2 (N327, N318, N288);
nor NOR3 (N328, N319, N142, N112);
nand NAND3 (N329, N324, N190, N222);
buf BUF1 (N330, N328);
not NOT1 (N331, N323);
or OR3 (N332, N317, N241, N118);
nand NAND4 (N333, N327, N154, N44, N150);
nor NOR2 (N334, N298, N60);
and AND3 (N335, N330, N244, N247);
or OR4 (N336, N326, N115, N199, N61);
and AND4 (N337, N312, N330, N193, N224);
nor NOR4 (N338, N329, N155, N261, N186);
and AND3 (N339, N336, N276, N39);
not NOT1 (N340, N331);
and AND2 (N341, N333, N141);
xor XOR2 (N342, N339, N255);
nor NOR2 (N343, N337, N159);
nand NAND4 (N344, N340, N150, N26, N83);
not NOT1 (N345, N325);
or OR3 (N346, N341, N235, N217);
nor NOR2 (N347, N334, N50);
and AND2 (N348, N347, N60);
not NOT1 (N349, N348);
buf BUF1 (N350, N306);
nand NAND3 (N351, N335, N260, N31);
not NOT1 (N352, N342);
not NOT1 (N353, N349);
not NOT1 (N354, N338);
not NOT1 (N355, N345);
and AND4 (N356, N344, N220, N123, N186);
nand NAND2 (N357, N354, N201);
nand NAND2 (N358, N353, N74);
and AND3 (N359, N346, N180, N164);
and AND3 (N360, N357, N185, N218);
nand NAND2 (N361, N350, N56);
not NOT1 (N362, N352);
nand NAND2 (N363, N356, N291);
nor NOR2 (N364, N363, N43);
not NOT1 (N365, N359);
nor NOR3 (N366, N332, N103, N158);
and AND4 (N367, N343, N153, N101, N319);
nand NAND4 (N368, N366, N172, N187, N105);
xor XOR2 (N369, N361, N181);
nand NAND3 (N370, N362, N97, N215);
buf BUF1 (N371, N355);
nor NOR2 (N372, N365, N147);
not NOT1 (N373, N371);
nand NAND2 (N374, N364, N361);
nand NAND3 (N375, N370, N45, N303);
xor XOR2 (N376, N369, N228);
nor NOR2 (N377, N351, N234);
xor XOR2 (N378, N360, N323);
nand NAND3 (N379, N378, N342, N155);
or OR2 (N380, N379, N290);
xor XOR2 (N381, N376, N52);
nand NAND4 (N382, N368, N129, N376, N345);
nand NAND4 (N383, N375, N216, N378, N125);
and AND2 (N384, N381, N298);
not NOT1 (N385, N377);
and AND2 (N386, N385, N358);
nor NOR4 (N387, N113, N336, N361, N245);
nor NOR2 (N388, N373, N342);
or OR2 (N389, N380, N141);
not NOT1 (N390, N367);
or OR3 (N391, N383, N349, N154);
buf BUF1 (N392, N372);
and AND3 (N393, N389, N110, N374);
not NOT1 (N394, N100);
xor XOR2 (N395, N384, N95);
nand NAND2 (N396, N387, N112);
or OR3 (N397, N392, N286, N212);
and AND4 (N398, N395, N96, N145, N68);
nand NAND4 (N399, N386, N35, N332, N275);
xor XOR2 (N400, N398, N71);
or OR3 (N401, N396, N172, N307);
not NOT1 (N402, N388);
buf BUF1 (N403, N394);
buf BUF1 (N404, N400);
xor XOR2 (N405, N393, N129);
not NOT1 (N406, N382);
and AND3 (N407, N399, N40, N347);
not NOT1 (N408, N404);
nor NOR4 (N409, N403, N268, N279, N148);
or OR4 (N410, N390, N241, N123, N38);
xor XOR2 (N411, N402, N118);
nand NAND2 (N412, N409, N264);
not NOT1 (N413, N410);
not NOT1 (N414, N411);
xor XOR2 (N415, N405, N75);
xor XOR2 (N416, N397, N385);
and AND2 (N417, N413, N76);
nor NOR4 (N418, N412, N42, N74, N257);
not NOT1 (N419, N391);
xor XOR2 (N420, N401, N350);
not NOT1 (N421, N407);
and AND3 (N422, N417, N188, N168);
and AND4 (N423, N406, N3, N193, N19);
buf BUF1 (N424, N415);
nor NOR2 (N425, N408, N186);
not NOT1 (N426, N422);
xor XOR2 (N427, N420, N92);
or OR4 (N428, N423, N3, N317, N209);
nor NOR3 (N429, N418, N34, N57);
nand NAND4 (N430, N427, N45, N23, N84);
buf BUF1 (N431, N424);
not NOT1 (N432, N419);
or OR3 (N433, N429, N223, N199);
buf BUF1 (N434, N428);
not NOT1 (N435, N432);
nand NAND2 (N436, N414, N281);
xor XOR2 (N437, N434, N364);
and AND2 (N438, N433, N406);
nand NAND3 (N439, N416, N215, N117);
or OR2 (N440, N436, N192);
xor XOR2 (N441, N435, N177);
not NOT1 (N442, N421);
xor XOR2 (N443, N430, N291);
not NOT1 (N444, N439);
or OR3 (N445, N444, N310, N23);
buf BUF1 (N446, N425);
not NOT1 (N447, N437);
xor XOR2 (N448, N443, N247);
or OR4 (N449, N445, N66, N24, N370);
nand NAND4 (N450, N440, N238, N359, N83);
and AND4 (N451, N442, N20, N247, N322);
not NOT1 (N452, N448);
and AND2 (N453, N451, N237);
nand NAND2 (N454, N446, N400);
xor XOR2 (N455, N452, N136);
and AND2 (N456, N453, N220);
not NOT1 (N457, N450);
nor NOR4 (N458, N431, N87, N311, N289);
nand NAND4 (N459, N457, N346, N128, N45);
nor NOR4 (N460, N447, N215, N29, N191);
and AND3 (N461, N441, N425, N396);
not NOT1 (N462, N461);
not NOT1 (N463, N459);
buf BUF1 (N464, N462);
nand NAND3 (N465, N458, N198, N75);
nor NOR3 (N466, N449, N170, N141);
buf BUF1 (N467, N455);
or OR4 (N468, N456, N260, N107, N81);
or OR3 (N469, N460, N13, N123);
or OR4 (N470, N469, N423, N24, N177);
or OR3 (N471, N468, N373, N90);
nand NAND3 (N472, N470, N111, N203);
xor XOR2 (N473, N465, N151);
xor XOR2 (N474, N464, N129);
xor XOR2 (N475, N474, N153);
not NOT1 (N476, N473);
nor NOR3 (N477, N454, N305, N92);
not NOT1 (N478, N475);
or OR4 (N479, N478, N188, N424, N388);
nor NOR4 (N480, N476, N217, N37, N309);
not NOT1 (N481, N463);
nor NOR4 (N482, N426, N466, N360, N297);
and AND2 (N483, N336, N389);
and AND3 (N484, N471, N188, N254);
nor NOR3 (N485, N479, N274, N251);
not NOT1 (N486, N477);
nand NAND3 (N487, N482, N170, N341);
nor NOR4 (N488, N484, N248, N265, N204);
xor XOR2 (N489, N487, N154);
xor XOR2 (N490, N467, N95);
or OR4 (N491, N480, N382, N35, N318);
buf BUF1 (N492, N485);
buf BUF1 (N493, N490);
and AND4 (N494, N491, N310, N412, N239);
not NOT1 (N495, N488);
nand NAND2 (N496, N486, N297);
nor NOR2 (N497, N492, N473);
not NOT1 (N498, N481);
xor XOR2 (N499, N497, N491);
buf BUF1 (N500, N483);
xor XOR2 (N501, N472, N344);
not NOT1 (N502, N500);
and AND4 (N503, N489, N382, N355, N320);
nand NAND3 (N504, N438, N308, N204);
nand NAND4 (N505, N493, N185, N491, N48);
nor NOR4 (N506, N504, N426, N301, N213);
buf BUF1 (N507, N494);
nor NOR2 (N508, N502, N251);
xor XOR2 (N509, N507, N292);
buf BUF1 (N510, N498);
nor NOR3 (N511, N503, N441, N57);
nand NAND2 (N512, N499, N269);
nand NAND4 (N513, N511, N163, N266, N95);
not NOT1 (N514, N508);
nor NOR4 (N515, N495, N48, N478, N341);
buf BUF1 (N516, N505);
nor NOR2 (N517, N515, N398);
not NOT1 (N518, N496);
nor NOR4 (N519, N512, N57, N441, N463);
nor NOR4 (N520, N517, N397, N318, N327);
or OR3 (N521, N501, N508, N50);
or OR2 (N522, N520, N379);
nand NAND2 (N523, N519, N272);
xor XOR2 (N524, N522, N75);
and AND2 (N525, N523, N102);
nand NAND4 (N526, N518, N17, N251, N193);
buf BUF1 (N527, N516);
and AND3 (N528, N526, N442, N378);
or OR4 (N529, N527, N378, N526, N309);
xor XOR2 (N530, N510, N235);
xor XOR2 (N531, N513, N313);
or OR4 (N532, N530, N374, N145, N59);
nor NOR4 (N533, N506, N270, N284, N509);
nor NOR2 (N534, N482, N147);
buf BUF1 (N535, N528);
or OR2 (N536, N524, N34);
and AND2 (N537, N514, N487);
not NOT1 (N538, N531);
not NOT1 (N539, N525);
nand NAND2 (N540, N521, N417);
nand NAND3 (N541, N540, N225, N119);
xor XOR2 (N542, N538, N31);
and AND2 (N543, N536, N236);
or OR4 (N544, N529, N396, N271, N406);
and AND3 (N545, N535, N235, N469);
or OR2 (N546, N542, N175);
nor NOR3 (N547, N543, N307, N282);
buf BUF1 (N548, N532);
or OR2 (N549, N541, N261);
nand NAND2 (N550, N544, N440);
not NOT1 (N551, N545);
nor NOR4 (N552, N537, N382, N111, N226);
or OR4 (N553, N552, N37, N194, N227);
or OR3 (N554, N534, N351, N333);
buf BUF1 (N555, N539);
nand NAND2 (N556, N554, N544);
or OR4 (N557, N551, N439, N108, N215);
buf BUF1 (N558, N553);
and AND4 (N559, N548, N46, N424, N157);
nand NAND4 (N560, N549, N185, N101, N373);
or OR3 (N561, N555, N105, N226);
buf BUF1 (N562, N558);
xor XOR2 (N563, N562, N68);
xor XOR2 (N564, N563, N89);
nor NOR2 (N565, N560, N218);
xor XOR2 (N566, N559, N301);
not NOT1 (N567, N566);
or OR3 (N568, N546, N280, N110);
nor NOR2 (N569, N557, N508);
nand NAND2 (N570, N564, N186);
nor NOR4 (N571, N567, N340, N80, N535);
nand NAND4 (N572, N565, N174, N239, N78);
nor NOR4 (N573, N533, N192, N346, N127);
buf BUF1 (N574, N561);
and AND4 (N575, N556, N44, N469, N131);
not NOT1 (N576, N573);
or OR2 (N577, N570, N523);
nand NAND2 (N578, N547, N20);
buf BUF1 (N579, N550);
or OR3 (N580, N572, N259, N489);
buf BUF1 (N581, N576);
buf BUF1 (N582, N571);
buf BUF1 (N583, N581);
nand NAND3 (N584, N580, N540, N440);
or OR3 (N585, N575, N427, N324);
and AND2 (N586, N577, N462);
nand NAND2 (N587, N578, N137);
nand NAND4 (N588, N586, N417, N401, N108);
not NOT1 (N589, N569);
xor XOR2 (N590, N589, N478);
xor XOR2 (N591, N587, N284);
not NOT1 (N592, N574);
or OR3 (N593, N583, N282, N117);
buf BUF1 (N594, N585);
not NOT1 (N595, N590);
nand NAND4 (N596, N594, N386, N333, N5);
and AND4 (N597, N596, N207, N527, N261);
or OR2 (N598, N592, N528);
nand NAND4 (N599, N579, N586, N519, N253);
not NOT1 (N600, N591);
not NOT1 (N601, N598);
and AND4 (N602, N601, N566, N398, N5);
or OR3 (N603, N599, N209, N580);
xor XOR2 (N604, N568, N11);
nand NAND3 (N605, N582, N91, N421);
not NOT1 (N606, N600);
nand NAND3 (N607, N588, N283, N443);
buf BUF1 (N608, N584);
and AND3 (N609, N604, N89, N456);
nor NOR3 (N610, N608, N90, N238);
xor XOR2 (N611, N602, N121);
not NOT1 (N612, N593);
not NOT1 (N613, N609);
or OR4 (N614, N595, N47, N510, N314);
nor NOR2 (N615, N611, N548);
and AND3 (N616, N614, N421, N240);
nor NOR2 (N617, N616, N177);
buf BUF1 (N618, N610);
or OR3 (N619, N603, N142, N151);
buf BUF1 (N620, N605);
endmodule