// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N1510,N1514,N1516,N1512,N1508,N1509,N1501,N1503,N1506,N1517;

not NOT1 (N18, N4);
and AND4 (N19, N16, N18, N3, N2);
and AND2 (N20, N16, N14);
nor NOR4 (N21, N11, N19, N12, N15);
and AND2 (N22, N11, N13);
not NOT1 (N23, N21);
or OR4 (N24, N23, N17, N7, N21);
nand NAND3 (N25, N7, N6, N9);
and AND2 (N26, N3, N25);
not NOT1 (N27, N23);
or OR3 (N28, N20, N14, N14);
not NOT1 (N29, N25);
not NOT1 (N30, N28);
xor XOR2 (N31, N5, N21);
xor XOR2 (N32, N23, N1);
and AND2 (N33, N14, N2);
or OR3 (N34, N9, N18, N6);
and AND4 (N35, N33, N21, N10, N13);
nand NAND4 (N36, N22, N32, N24, N11);
xor XOR2 (N37, N1, N32);
xor XOR2 (N38, N18, N12);
nand NAND3 (N39, N38, N13, N38);
xor XOR2 (N40, N26, N29);
nand NAND3 (N41, N34, N16, N1);
nand NAND2 (N42, N22, N41);
nor NOR3 (N43, N40, N25, N1);
nand NAND2 (N44, N26, N16);
or OR2 (N45, N35, N20);
nor NOR4 (N46, N44, N4, N22, N40);
not NOT1 (N47, N45);
or OR2 (N48, N43, N13);
not NOT1 (N49, N37);
nand NAND3 (N50, N48, N24, N41);
nand NAND4 (N51, N39, N17, N2, N42);
nor NOR4 (N52, N7, N47, N46, N11);
buf BUF1 (N53, N44);
nor NOR2 (N54, N18, N48);
buf BUF1 (N55, N51);
nor NOR2 (N56, N31, N35);
not NOT1 (N57, N53);
xor XOR2 (N58, N36, N21);
not NOT1 (N59, N30);
nand NAND4 (N60, N58, N12, N4, N56);
not NOT1 (N61, N15);
buf BUF1 (N62, N61);
nand NAND2 (N63, N54, N6);
nor NOR3 (N64, N27, N8, N12);
or OR2 (N65, N64, N41);
or OR3 (N66, N60, N34, N62);
xor XOR2 (N67, N40, N33);
xor XOR2 (N68, N49, N42);
nor NOR2 (N69, N59, N51);
xor XOR2 (N70, N65, N28);
nor NOR2 (N71, N68, N8);
nand NAND4 (N72, N71, N45, N69, N9);
nor NOR2 (N73, N33, N72);
or OR3 (N74, N47, N55, N63);
and AND2 (N75, N18, N47);
or OR4 (N76, N74, N19, N57, N47);
buf BUF1 (N77, N10);
nor NOR4 (N78, N11, N1, N58, N6);
or OR2 (N79, N52, N26);
buf BUF1 (N80, N67);
and AND2 (N81, N77, N53);
nand NAND4 (N82, N70, N45, N66, N28);
or OR2 (N83, N1, N5);
nand NAND3 (N84, N80, N51, N12);
buf BUF1 (N85, N76);
and AND4 (N86, N85, N58, N48, N34);
nor NOR4 (N87, N84, N67, N65, N63);
buf BUF1 (N88, N86);
or OR2 (N89, N87, N13);
or OR2 (N90, N50, N21);
nor NOR3 (N91, N89, N20, N72);
and AND2 (N92, N78, N52);
nor NOR3 (N93, N88, N76, N64);
xor XOR2 (N94, N92, N11);
not NOT1 (N95, N83);
nand NAND4 (N96, N93, N5, N35, N52);
not NOT1 (N97, N82);
nand NAND4 (N98, N90, N43, N36, N71);
nand NAND3 (N99, N91, N95, N22);
buf BUF1 (N100, N96);
or OR2 (N101, N68, N68);
or OR3 (N102, N98, N90, N65);
nor NOR2 (N103, N79, N36);
buf BUF1 (N104, N99);
and AND2 (N105, N81, N103);
nor NOR2 (N106, N70, N41);
and AND4 (N107, N105, N32, N35, N67);
xor XOR2 (N108, N94, N96);
xor XOR2 (N109, N101, N82);
or OR4 (N110, N73, N87, N31, N15);
nand NAND3 (N111, N107, N29, N8);
nand NAND2 (N112, N109, N83);
not NOT1 (N113, N100);
and AND2 (N114, N106, N98);
buf BUF1 (N115, N110);
not NOT1 (N116, N104);
not NOT1 (N117, N102);
xor XOR2 (N118, N113, N75);
or OR4 (N119, N87, N72, N21, N88);
nor NOR3 (N120, N112, N65, N69);
not NOT1 (N121, N97);
xor XOR2 (N122, N119, N18);
buf BUF1 (N123, N118);
xor XOR2 (N124, N122, N73);
nor NOR2 (N125, N111, N119);
nand NAND3 (N126, N120, N71, N63);
not NOT1 (N127, N117);
nor NOR2 (N128, N125, N58);
nor NOR2 (N129, N127, N66);
xor XOR2 (N130, N116, N101);
xor XOR2 (N131, N123, N39);
xor XOR2 (N132, N126, N83);
not NOT1 (N133, N124);
buf BUF1 (N134, N133);
nor NOR4 (N135, N130, N120, N11, N18);
or OR4 (N136, N129, N69, N46, N132);
buf BUF1 (N137, N67);
or OR3 (N138, N114, N115, N130);
and AND2 (N139, N55, N29);
buf BUF1 (N140, N139);
xor XOR2 (N141, N121, N94);
or OR2 (N142, N128, N58);
or OR4 (N143, N138, N71, N44, N14);
not NOT1 (N144, N140);
and AND3 (N145, N135, N63, N88);
and AND2 (N146, N141, N60);
xor XOR2 (N147, N134, N88);
not NOT1 (N148, N108);
buf BUF1 (N149, N145);
and AND4 (N150, N149, N94, N76, N9);
nor NOR2 (N151, N136, N18);
and AND3 (N152, N144, N63, N115);
or OR2 (N153, N146, N136);
nand NAND3 (N154, N131, N54, N150);
not NOT1 (N155, N106);
and AND4 (N156, N148, N107, N26, N82);
nor NOR3 (N157, N152, N31, N20);
and AND2 (N158, N157, N136);
nand NAND2 (N159, N137, N96);
and AND4 (N160, N147, N97, N125, N123);
buf BUF1 (N161, N159);
not NOT1 (N162, N158);
nand NAND3 (N163, N153, N98, N94);
or OR4 (N164, N156, N20, N154, N117);
nor NOR4 (N165, N67, N155, N116, N85);
xor XOR2 (N166, N102, N115);
not NOT1 (N167, N163);
not NOT1 (N168, N161);
or OR2 (N169, N168, N44);
and AND3 (N170, N169, N125, N35);
buf BUF1 (N171, N151);
and AND2 (N172, N171, N57);
not NOT1 (N173, N160);
and AND3 (N174, N173, N128, N86);
nand NAND2 (N175, N164, N70);
buf BUF1 (N176, N175);
nand NAND4 (N177, N165, N99, N77, N64);
buf BUF1 (N178, N166);
nor NOR4 (N179, N177, N177, N70, N89);
xor XOR2 (N180, N162, N111);
nor NOR3 (N181, N180, N2, N34);
or OR3 (N182, N167, N23, N101);
xor XOR2 (N183, N143, N64);
nor NOR2 (N184, N172, N33);
xor XOR2 (N185, N184, N112);
and AND4 (N186, N182, N159, N39, N59);
and AND4 (N187, N181, N186, N12, N12);
nand NAND4 (N188, N34, N60, N170, N91);
not NOT1 (N189, N45);
not NOT1 (N190, N179);
nand NAND4 (N191, N188, N107, N120, N97);
and AND2 (N192, N183, N13);
or OR3 (N193, N192, N82, N61);
and AND4 (N194, N176, N69, N190, N137);
buf BUF1 (N195, N53);
not NOT1 (N196, N193);
xor XOR2 (N197, N178, N83);
xor XOR2 (N198, N174, N13);
not NOT1 (N199, N195);
nor NOR2 (N200, N142, N94);
and AND3 (N201, N185, N83, N109);
or OR2 (N202, N201, N92);
buf BUF1 (N203, N191);
not NOT1 (N204, N200);
buf BUF1 (N205, N202);
xor XOR2 (N206, N204, N172);
not NOT1 (N207, N206);
or OR4 (N208, N198, N7, N180, N79);
nor NOR2 (N209, N187, N26);
nor NOR2 (N210, N205, N27);
or OR2 (N211, N208, N101);
xor XOR2 (N212, N210, N147);
nand NAND2 (N213, N212, N112);
and AND4 (N214, N189, N139, N189, N28);
nor NOR4 (N215, N214, N126, N194, N132);
nor NOR4 (N216, N160, N56, N8, N52);
nand NAND4 (N217, N216, N185, N102, N58);
not NOT1 (N218, N199);
nand NAND2 (N219, N218, N101);
nand NAND3 (N220, N207, N56, N122);
nor NOR3 (N221, N196, N112, N45);
and AND3 (N222, N217, N52, N89);
nor NOR2 (N223, N215, N206);
nand NAND4 (N224, N209, N54, N17, N215);
or OR2 (N225, N222, N26);
nor NOR2 (N226, N224, N166);
buf BUF1 (N227, N220);
xor XOR2 (N228, N197, N163);
not NOT1 (N229, N225);
not NOT1 (N230, N203);
buf BUF1 (N231, N227);
nor NOR4 (N232, N223, N204, N153, N115);
not NOT1 (N233, N221);
buf BUF1 (N234, N226);
nand NAND3 (N235, N228, N185, N205);
not NOT1 (N236, N234);
not NOT1 (N237, N219);
not NOT1 (N238, N230);
nand NAND3 (N239, N235, N178, N187);
xor XOR2 (N240, N232, N100);
xor XOR2 (N241, N239, N196);
not NOT1 (N242, N240);
buf BUF1 (N243, N241);
and AND4 (N244, N242, N99, N53, N172);
xor XOR2 (N245, N213, N42);
and AND4 (N246, N229, N19, N171, N43);
buf BUF1 (N247, N244);
nor NOR2 (N248, N247, N43);
and AND4 (N249, N248, N99, N159, N142);
or OR4 (N250, N231, N63, N175, N168);
nor NOR3 (N251, N236, N135, N14);
xor XOR2 (N252, N243, N228);
nand NAND4 (N253, N252, N64, N179, N16);
xor XOR2 (N254, N238, N40);
nand NAND2 (N255, N233, N148);
xor XOR2 (N256, N254, N177);
nor NOR4 (N257, N250, N146, N17, N102);
and AND3 (N258, N237, N32, N208);
not NOT1 (N259, N253);
and AND4 (N260, N249, N15, N82, N11);
nand NAND4 (N261, N211, N130, N109, N5);
nand NAND2 (N262, N255, N199);
not NOT1 (N263, N246);
buf BUF1 (N264, N262);
or OR3 (N265, N258, N243, N71);
not NOT1 (N266, N256);
buf BUF1 (N267, N245);
nand NAND4 (N268, N265, N1, N209, N213);
and AND2 (N269, N267, N222);
not NOT1 (N270, N269);
and AND4 (N271, N270, N136, N15, N208);
nor NOR2 (N272, N264, N48);
nor NOR4 (N273, N271, N116, N147, N96);
nand NAND2 (N274, N268, N215);
nor NOR2 (N275, N260, N9);
nor NOR4 (N276, N251, N111, N82, N247);
xor XOR2 (N277, N261, N225);
or OR4 (N278, N266, N198, N205, N159);
nand NAND4 (N279, N272, N77, N101, N109);
or OR4 (N280, N274, N16, N133, N138);
or OR2 (N281, N276, N134);
and AND4 (N282, N281, N189, N56, N90);
buf BUF1 (N283, N279);
nand NAND2 (N284, N280, N115);
and AND2 (N285, N284, N105);
buf BUF1 (N286, N277);
nand NAND4 (N287, N282, N218, N202, N230);
not NOT1 (N288, N257);
buf BUF1 (N289, N286);
nand NAND3 (N290, N289, N45, N22);
nor NOR4 (N291, N263, N207, N62, N274);
nand NAND4 (N292, N291, N80, N12, N245);
or OR3 (N293, N290, N228, N56);
xor XOR2 (N294, N275, N57);
xor XOR2 (N295, N285, N153);
nand NAND2 (N296, N294, N244);
nor NOR2 (N297, N296, N197);
not NOT1 (N298, N293);
and AND4 (N299, N287, N220, N126, N19);
nand NAND2 (N300, N273, N207);
nor NOR4 (N301, N295, N30, N60, N24);
xor XOR2 (N302, N259, N206);
nor NOR2 (N303, N288, N34);
nor NOR2 (N304, N303, N81);
buf BUF1 (N305, N299);
xor XOR2 (N306, N305, N157);
not NOT1 (N307, N306);
and AND3 (N308, N301, N198, N136);
nand NAND4 (N309, N298, N242, N179, N20);
buf BUF1 (N310, N302);
buf BUF1 (N311, N304);
nand NAND4 (N312, N300, N256, N265, N8);
or OR3 (N313, N308, N285, N282);
xor XOR2 (N314, N283, N166);
buf BUF1 (N315, N292);
buf BUF1 (N316, N278);
xor XOR2 (N317, N312, N111);
nand NAND3 (N318, N314, N291, N162);
xor XOR2 (N319, N318, N148);
buf BUF1 (N320, N297);
nor NOR3 (N321, N307, N310, N175);
buf BUF1 (N322, N216);
nand NAND3 (N323, N319, N178, N163);
nor NOR2 (N324, N323, N54);
and AND3 (N325, N322, N269, N190);
buf BUF1 (N326, N309);
or OR4 (N327, N320, N286, N129, N33);
xor XOR2 (N328, N327, N307);
buf BUF1 (N329, N315);
buf BUF1 (N330, N313);
nor NOR4 (N331, N317, N122, N241, N303);
or OR4 (N332, N311, N134, N290, N11);
nand NAND2 (N333, N325, N166);
nor NOR4 (N334, N324, N215, N140, N309);
nor NOR3 (N335, N321, N51, N38);
nor NOR4 (N336, N331, N149, N18, N206);
and AND3 (N337, N333, N320, N5);
xor XOR2 (N338, N329, N257);
and AND3 (N339, N332, N133, N210);
nand NAND3 (N340, N334, N44, N226);
nor NOR3 (N341, N340, N111, N123);
and AND4 (N342, N336, N147, N139, N157);
and AND4 (N343, N342, N28, N132, N154);
nand NAND4 (N344, N337, N237, N298, N19);
nand NAND4 (N345, N343, N41, N220, N165);
not NOT1 (N346, N341);
nand NAND2 (N347, N346, N110);
and AND3 (N348, N338, N326, N54);
and AND2 (N349, N290, N45);
buf BUF1 (N350, N335);
buf BUF1 (N351, N345);
buf BUF1 (N352, N330);
xor XOR2 (N353, N352, N347);
buf BUF1 (N354, N188);
nand NAND2 (N355, N344, N341);
not NOT1 (N356, N328);
not NOT1 (N357, N350);
and AND4 (N358, N356, N51, N56, N63);
and AND4 (N359, N351, N217, N75, N158);
nor NOR4 (N360, N353, N303, N249, N303);
or OR4 (N361, N359, N86, N22, N83);
buf BUF1 (N362, N358);
not NOT1 (N363, N357);
buf BUF1 (N364, N349);
xor XOR2 (N365, N348, N79);
nor NOR4 (N366, N362, N34, N130, N149);
nor NOR2 (N367, N365, N308);
xor XOR2 (N368, N361, N345);
not NOT1 (N369, N354);
nand NAND3 (N370, N363, N19, N271);
and AND3 (N371, N339, N340, N210);
not NOT1 (N372, N368);
nor NOR4 (N373, N360, N169, N192, N194);
not NOT1 (N374, N355);
or OR2 (N375, N374, N200);
nor NOR3 (N376, N364, N313, N210);
not NOT1 (N377, N366);
nor NOR3 (N378, N373, N14, N205);
nand NAND2 (N379, N372, N214);
and AND3 (N380, N375, N185, N290);
not NOT1 (N381, N378);
buf BUF1 (N382, N316);
xor XOR2 (N383, N369, N183);
and AND2 (N384, N367, N269);
not NOT1 (N385, N383);
and AND3 (N386, N385, N368, N271);
nor NOR4 (N387, N382, N78, N67, N44);
and AND3 (N388, N380, N317, N164);
nor NOR2 (N389, N387, N356);
buf BUF1 (N390, N381);
buf BUF1 (N391, N371);
buf BUF1 (N392, N388);
nor NOR4 (N393, N386, N119, N326, N166);
and AND3 (N394, N377, N343, N121);
or OR2 (N395, N370, N19);
or OR2 (N396, N394, N265);
nand NAND4 (N397, N390, N267, N244, N41);
or OR4 (N398, N395, N393, N61, N291);
not NOT1 (N399, N71);
nor NOR2 (N400, N392, N64);
and AND4 (N401, N397, N109, N126, N196);
not NOT1 (N402, N400);
and AND4 (N403, N376, N150, N361, N3);
nor NOR2 (N404, N379, N384);
and AND4 (N405, N90, N360, N89, N343);
nor NOR3 (N406, N391, N398, N144);
buf BUF1 (N407, N37);
buf BUF1 (N408, N396);
xor XOR2 (N409, N402, N176);
or OR2 (N410, N403, N319);
buf BUF1 (N411, N406);
nand NAND2 (N412, N389, N407);
nor NOR3 (N413, N114, N179, N408);
xor XOR2 (N414, N384, N51);
and AND2 (N415, N412, N185);
buf BUF1 (N416, N401);
and AND3 (N417, N405, N178, N340);
nand NAND4 (N418, N416, N276, N252, N241);
or OR3 (N419, N399, N188, N401);
not NOT1 (N420, N404);
or OR3 (N421, N417, N409, N146);
nand NAND2 (N422, N101, N178);
or OR2 (N423, N421, N212);
or OR3 (N424, N420, N289, N349);
or OR3 (N425, N413, N111, N376);
not NOT1 (N426, N410);
nor NOR4 (N427, N414, N60, N258, N337);
nor NOR3 (N428, N418, N362, N224);
xor XOR2 (N429, N415, N295);
not NOT1 (N430, N424);
xor XOR2 (N431, N422, N387);
buf BUF1 (N432, N411);
nor NOR3 (N433, N419, N42, N29);
buf BUF1 (N434, N431);
not NOT1 (N435, N432);
xor XOR2 (N436, N433, N410);
nor NOR4 (N437, N426, N410, N145, N256);
or OR2 (N438, N425, N308);
buf BUF1 (N439, N436);
and AND4 (N440, N430, N296, N92, N6);
not NOT1 (N441, N428);
not NOT1 (N442, N441);
or OR2 (N443, N429, N73);
xor XOR2 (N444, N442, N372);
or OR4 (N445, N437, N334, N311, N140);
nor NOR4 (N446, N445, N374, N24, N429);
buf BUF1 (N447, N434);
not NOT1 (N448, N440);
xor XOR2 (N449, N444, N69);
not NOT1 (N450, N427);
not NOT1 (N451, N446);
buf BUF1 (N452, N443);
buf BUF1 (N453, N448);
not NOT1 (N454, N439);
and AND2 (N455, N452, N410);
nor NOR3 (N456, N447, N389, N132);
xor XOR2 (N457, N449, N329);
or OR4 (N458, N450, N305, N40, N50);
xor XOR2 (N459, N454, N151);
and AND3 (N460, N423, N314, N406);
and AND3 (N461, N459, N134, N206);
or OR2 (N462, N438, N440);
buf BUF1 (N463, N462);
xor XOR2 (N464, N453, N135);
xor XOR2 (N465, N460, N263);
nand NAND4 (N466, N451, N143, N430, N264);
not NOT1 (N467, N435);
and AND4 (N468, N455, N229, N233, N387);
or OR4 (N469, N463, N439, N356, N184);
nor NOR3 (N470, N468, N196, N361);
buf BUF1 (N471, N469);
buf BUF1 (N472, N464);
and AND4 (N473, N456, N248, N62, N415);
buf BUF1 (N474, N465);
nor NOR4 (N475, N474, N330, N395, N95);
nand NAND3 (N476, N473, N24, N455);
or OR2 (N477, N475, N418);
and AND4 (N478, N457, N255, N206, N282);
xor XOR2 (N479, N470, N374);
or OR4 (N480, N467, N229, N98, N104);
nand NAND2 (N481, N479, N364);
not NOT1 (N482, N471);
buf BUF1 (N483, N461);
nand NAND3 (N484, N478, N303, N128);
and AND2 (N485, N476, N235);
xor XOR2 (N486, N458, N130);
nand NAND4 (N487, N480, N401, N249, N269);
and AND4 (N488, N466, N416, N94, N91);
nor NOR4 (N489, N487, N281, N101, N425);
buf BUF1 (N490, N485);
and AND3 (N491, N484, N223, N104);
nand NAND3 (N492, N482, N177, N14);
or OR2 (N493, N481, N272);
not NOT1 (N494, N483);
and AND2 (N495, N493, N18);
nand NAND4 (N496, N491, N164, N407, N245);
buf BUF1 (N497, N495);
nor NOR4 (N498, N477, N483, N283, N440);
nand NAND3 (N499, N489, N394, N223);
and AND2 (N500, N486, N452);
or OR2 (N501, N498, N271);
or OR3 (N502, N500, N157, N234);
buf BUF1 (N503, N499);
nor NOR3 (N504, N494, N80, N344);
nor NOR4 (N505, N488, N348, N229, N332);
nand NAND4 (N506, N472, N205, N12, N485);
buf BUF1 (N507, N505);
or OR2 (N508, N497, N503);
or OR2 (N509, N374, N458);
not NOT1 (N510, N492);
buf BUF1 (N511, N501);
and AND3 (N512, N504, N225, N55);
nor NOR3 (N513, N507, N214, N502);
buf BUF1 (N514, N45);
or OR2 (N515, N509, N238);
not NOT1 (N516, N496);
nand NAND4 (N517, N514, N26, N308, N117);
xor XOR2 (N518, N511, N436);
nand NAND2 (N519, N490, N86);
buf BUF1 (N520, N513);
nand NAND4 (N521, N515, N402, N63, N359);
or OR4 (N522, N520, N449, N511, N301);
and AND4 (N523, N518, N196, N4, N76);
xor XOR2 (N524, N506, N419);
or OR4 (N525, N516, N216, N190, N444);
nor NOR2 (N526, N510, N212);
xor XOR2 (N527, N521, N135);
and AND4 (N528, N525, N145, N449, N261);
xor XOR2 (N529, N522, N274);
not NOT1 (N530, N528);
not NOT1 (N531, N530);
buf BUF1 (N532, N512);
nand NAND2 (N533, N531, N137);
and AND3 (N534, N523, N21, N42);
nor NOR3 (N535, N534, N401, N197);
xor XOR2 (N536, N533, N334);
nand NAND4 (N537, N536, N529, N495, N444);
buf BUF1 (N538, N110);
or OR2 (N539, N537, N194);
nor NOR2 (N540, N519, N472);
xor XOR2 (N541, N532, N285);
buf BUF1 (N542, N526);
nand NAND3 (N543, N541, N67, N69);
and AND3 (N544, N538, N94, N123);
and AND2 (N545, N535, N516);
nand NAND2 (N546, N524, N278);
nor NOR4 (N547, N544, N365, N241, N17);
not NOT1 (N548, N546);
nor NOR3 (N549, N545, N502, N357);
or OR4 (N550, N517, N443, N103, N368);
xor XOR2 (N551, N548, N5);
not NOT1 (N552, N543);
or OR3 (N553, N552, N541, N28);
or OR3 (N554, N540, N290, N20);
not NOT1 (N555, N550);
or OR4 (N556, N542, N62, N440, N104);
nor NOR2 (N557, N554, N40);
and AND3 (N558, N553, N474, N179);
buf BUF1 (N559, N551);
xor XOR2 (N560, N555, N79);
or OR3 (N561, N558, N264, N416);
not NOT1 (N562, N559);
nor NOR2 (N563, N508, N259);
nand NAND3 (N564, N549, N195, N334);
xor XOR2 (N565, N557, N168);
xor XOR2 (N566, N565, N88);
buf BUF1 (N567, N562);
buf BUF1 (N568, N566);
and AND2 (N569, N560, N31);
not NOT1 (N570, N556);
or OR4 (N571, N539, N99, N231, N102);
not NOT1 (N572, N547);
buf BUF1 (N573, N567);
or OR3 (N574, N569, N171, N103);
and AND2 (N575, N571, N85);
or OR3 (N576, N573, N24, N538);
or OR2 (N577, N568, N439);
or OR3 (N578, N561, N271, N275);
and AND2 (N579, N564, N160);
buf BUF1 (N580, N574);
nand NAND3 (N581, N578, N416, N246);
not NOT1 (N582, N527);
not NOT1 (N583, N580);
or OR3 (N584, N572, N368, N207);
and AND2 (N585, N582, N443);
not NOT1 (N586, N584);
buf BUF1 (N587, N570);
and AND4 (N588, N585, N206, N261, N309);
nand NAND4 (N589, N583, N567, N19, N121);
buf BUF1 (N590, N588);
xor XOR2 (N591, N579, N503);
nand NAND2 (N592, N577, N543);
not NOT1 (N593, N586);
buf BUF1 (N594, N590);
nand NAND2 (N595, N592, N38);
xor XOR2 (N596, N587, N33);
buf BUF1 (N597, N575);
buf BUF1 (N598, N596);
nand NAND4 (N599, N594, N112, N181, N190);
or OR4 (N600, N576, N378, N469, N126);
nand NAND2 (N601, N597, N317);
xor XOR2 (N602, N595, N272);
not NOT1 (N603, N593);
not NOT1 (N604, N600);
nand NAND4 (N605, N603, N594, N379, N173);
and AND3 (N606, N599, N265, N25);
nand NAND3 (N607, N591, N223, N530);
nor NOR3 (N608, N601, N15, N473);
not NOT1 (N609, N581);
and AND3 (N610, N598, N533, N402);
xor XOR2 (N611, N605, N483);
nand NAND2 (N612, N611, N302);
nand NAND2 (N613, N602, N60);
nor NOR4 (N614, N606, N351, N426, N266);
not NOT1 (N615, N612);
xor XOR2 (N616, N607, N291);
xor XOR2 (N617, N563, N143);
nor NOR3 (N618, N614, N8, N602);
nor NOR3 (N619, N618, N600, N371);
nor NOR3 (N620, N589, N129, N204);
nand NAND3 (N621, N613, N104, N505);
nand NAND3 (N622, N615, N612, N233);
and AND4 (N623, N621, N534, N369, N112);
buf BUF1 (N624, N622);
buf BUF1 (N625, N623);
or OR3 (N626, N619, N240, N470);
nand NAND4 (N627, N616, N351, N493, N228);
buf BUF1 (N628, N625);
and AND3 (N629, N610, N145, N276);
nor NOR4 (N630, N626, N448, N1, N381);
nand NAND4 (N631, N630, N450, N24, N501);
nor NOR2 (N632, N628, N518);
xor XOR2 (N633, N632, N8);
xor XOR2 (N634, N627, N238);
not NOT1 (N635, N624);
and AND3 (N636, N635, N212, N230);
xor XOR2 (N637, N609, N633);
xor XOR2 (N638, N62, N200);
and AND3 (N639, N634, N66, N147);
not NOT1 (N640, N620);
or OR4 (N641, N639, N527, N350, N370);
not NOT1 (N642, N640);
xor XOR2 (N643, N631, N496);
and AND3 (N644, N608, N311, N159);
not NOT1 (N645, N617);
xor XOR2 (N646, N643, N357);
or OR3 (N647, N646, N84, N211);
and AND4 (N648, N604, N125, N266, N306);
and AND4 (N649, N637, N184, N545, N126);
not NOT1 (N650, N645);
or OR2 (N651, N644, N103);
and AND3 (N652, N629, N577, N495);
nand NAND2 (N653, N649, N414);
and AND2 (N654, N652, N17);
or OR3 (N655, N638, N172, N317);
not NOT1 (N656, N641);
and AND3 (N657, N636, N429, N478);
nand NAND2 (N658, N642, N35);
nand NAND3 (N659, N654, N209, N480);
or OR3 (N660, N650, N498, N30);
xor XOR2 (N661, N660, N170);
nand NAND4 (N662, N655, N494, N353, N268);
nand NAND4 (N663, N647, N383, N335, N193);
buf BUF1 (N664, N663);
and AND3 (N665, N658, N107, N251);
buf BUF1 (N666, N662);
nor NOR3 (N667, N661, N592, N560);
and AND2 (N668, N651, N309);
not NOT1 (N669, N667);
not NOT1 (N670, N668);
not NOT1 (N671, N664);
nor NOR3 (N672, N656, N601, N386);
nand NAND4 (N673, N657, N401, N39, N80);
and AND3 (N674, N672, N415, N56);
nand NAND3 (N675, N670, N248, N148);
nor NOR2 (N676, N673, N403);
nand NAND4 (N677, N648, N443, N132, N489);
nor NOR4 (N678, N676, N241, N478, N434);
xor XOR2 (N679, N674, N247);
or OR2 (N680, N675, N321);
xor XOR2 (N681, N669, N493);
not NOT1 (N682, N671);
nand NAND4 (N683, N682, N35, N610, N360);
xor XOR2 (N684, N678, N483);
buf BUF1 (N685, N666);
and AND3 (N686, N677, N404, N643);
nand NAND2 (N687, N659, N176);
nand NAND4 (N688, N684, N553, N226, N545);
and AND4 (N689, N683, N618, N503, N233);
buf BUF1 (N690, N688);
not NOT1 (N691, N653);
nand NAND3 (N692, N665, N174, N471);
nor NOR2 (N693, N685, N578);
and AND3 (N694, N691, N114, N620);
and AND4 (N695, N687, N640, N150, N251);
not NOT1 (N696, N693);
buf BUF1 (N697, N695);
and AND4 (N698, N689, N106, N71, N141);
or OR3 (N699, N679, N322, N471);
nand NAND2 (N700, N681, N292);
xor XOR2 (N701, N690, N381);
or OR2 (N702, N697, N478);
buf BUF1 (N703, N700);
nor NOR3 (N704, N692, N309, N314);
or OR3 (N705, N694, N254, N523);
not NOT1 (N706, N703);
nor NOR2 (N707, N696, N559);
not NOT1 (N708, N707);
nor NOR3 (N709, N698, N440, N192);
nand NAND3 (N710, N706, N332, N457);
buf BUF1 (N711, N705);
not NOT1 (N712, N709);
nand NAND2 (N713, N699, N424);
nand NAND4 (N714, N704, N58, N442, N34);
nor NOR2 (N715, N701, N458);
nand NAND3 (N716, N710, N523, N153);
not NOT1 (N717, N714);
xor XOR2 (N718, N702, N258);
or OR4 (N719, N686, N454, N372, N574);
xor XOR2 (N720, N711, N118);
or OR2 (N721, N708, N503);
nor NOR3 (N722, N721, N573, N498);
and AND4 (N723, N722, N514, N195, N558);
nor NOR4 (N724, N680, N195, N391, N598);
nand NAND3 (N725, N723, N675, N194);
and AND3 (N726, N715, N582, N186);
and AND3 (N727, N719, N470, N567);
xor XOR2 (N728, N718, N265);
or OR3 (N729, N727, N328, N447);
nand NAND2 (N730, N729, N77);
xor XOR2 (N731, N725, N507);
xor XOR2 (N732, N724, N249);
or OR4 (N733, N728, N46, N596, N663);
nand NAND2 (N734, N712, N545);
buf BUF1 (N735, N726);
xor XOR2 (N736, N732, N382);
or OR3 (N737, N731, N601, N321);
and AND3 (N738, N716, N540, N421);
or OR3 (N739, N737, N139, N119);
buf BUF1 (N740, N713);
and AND4 (N741, N730, N331, N605, N258);
and AND2 (N742, N733, N214);
xor XOR2 (N743, N739, N267);
buf BUF1 (N744, N717);
or OR3 (N745, N736, N650, N652);
buf BUF1 (N746, N734);
or OR3 (N747, N720, N505, N158);
or OR3 (N748, N746, N4, N577);
nor NOR3 (N749, N741, N433, N300);
buf BUF1 (N750, N747);
not NOT1 (N751, N740);
nand NAND2 (N752, N750, N118);
and AND2 (N753, N738, N605);
and AND3 (N754, N743, N543, N110);
nor NOR2 (N755, N752, N687);
xor XOR2 (N756, N749, N344);
not NOT1 (N757, N748);
and AND3 (N758, N735, N585, N346);
or OR3 (N759, N756, N332, N288);
nand NAND3 (N760, N744, N670, N267);
and AND4 (N761, N751, N336, N318, N279);
or OR3 (N762, N745, N199, N401);
nand NAND2 (N763, N742, N173);
or OR3 (N764, N763, N316, N258);
or OR3 (N765, N760, N438, N148);
xor XOR2 (N766, N762, N130);
xor XOR2 (N767, N759, N579);
nor NOR4 (N768, N764, N142, N325, N147);
and AND4 (N769, N755, N270, N344, N367);
xor XOR2 (N770, N765, N749);
nand NAND3 (N771, N754, N237, N355);
xor XOR2 (N772, N770, N169);
or OR3 (N773, N761, N727, N54);
xor XOR2 (N774, N753, N255);
buf BUF1 (N775, N773);
buf BUF1 (N776, N772);
xor XOR2 (N777, N768, N385);
nor NOR4 (N778, N776, N299, N359, N89);
buf BUF1 (N779, N775);
buf BUF1 (N780, N766);
or OR2 (N781, N769, N523);
nand NAND4 (N782, N771, N754, N591, N34);
nand NAND3 (N783, N780, N658, N414);
not NOT1 (N784, N778);
or OR4 (N785, N757, N633, N324, N272);
and AND3 (N786, N777, N485, N742);
or OR4 (N787, N779, N748, N600, N362);
nor NOR4 (N788, N785, N66, N724, N540);
or OR4 (N789, N787, N60, N327, N181);
nor NOR4 (N790, N786, N778, N706, N266);
or OR3 (N791, N784, N434, N540);
xor XOR2 (N792, N781, N439);
or OR2 (N793, N767, N263);
and AND2 (N794, N792, N410);
not NOT1 (N795, N794);
not NOT1 (N796, N791);
or OR2 (N797, N788, N520);
and AND4 (N798, N774, N405, N81, N2);
buf BUF1 (N799, N789);
nand NAND2 (N800, N799, N477);
and AND4 (N801, N797, N779, N54, N115);
or OR2 (N802, N795, N390);
xor XOR2 (N803, N801, N208);
xor XOR2 (N804, N803, N272);
xor XOR2 (N805, N804, N533);
nor NOR3 (N806, N805, N91, N710);
or OR2 (N807, N793, N628);
not NOT1 (N808, N807);
nor NOR2 (N809, N790, N288);
buf BUF1 (N810, N758);
xor XOR2 (N811, N802, N538);
not NOT1 (N812, N800);
or OR3 (N813, N810, N228, N242);
buf BUF1 (N814, N809);
or OR2 (N815, N814, N42);
nand NAND2 (N816, N782, N560);
nor NOR2 (N817, N808, N374);
nor NOR4 (N818, N806, N181, N752, N708);
xor XOR2 (N819, N798, N333);
not NOT1 (N820, N796);
xor XOR2 (N821, N819, N216);
nand NAND2 (N822, N821, N508);
not NOT1 (N823, N783);
and AND4 (N824, N820, N301, N211, N123);
nand NAND4 (N825, N823, N168, N234, N682);
or OR3 (N826, N824, N396, N455);
not NOT1 (N827, N817);
and AND2 (N828, N811, N653);
xor XOR2 (N829, N822, N346);
or OR4 (N830, N818, N501, N553, N479);
nor NOR3 (N831, N826, N704, N762);
nand NAND2 (N832, N812, N761);
and AND3 (N833, N825, N492, N239);
nand NAND4 (N834, N829, N353, N3, N200);
not NOT1 (N835, N815);
buf BUF1 (N836, N833);
nor NOR2 (N837, N830, N625);
nor NOR2 (N838, N835, N243);
nand NAND3 (N839, N831, N92, N657);
and AND2 (N840, N838, N806);
or OR2 (N841, N827, N80);
or OR2 (N842, N841, N380);
nor NOR3 (N843, N836, N585, N72);
or OR4 (N844, N834, N585, N500, N826);
not NOT1 (N845, N843);
nand NAND3 (N846, N839, N789, N656);
and AND2 (N847, N842, N275);
not NOT1 (N848, N845);
xor XOR2 (N849, N828, N91);
and AND2 (N850, N813, N176);
or OR4 (N851, N840, N788, N310, N354);
and AND2 (N852, N832, N553);
or OR4 (N853, N837, N787, N526, N687);
nor NOR4 (N854, N849, N552, N298, N664);
xor XOR2 (N855, N847, N548);
nand NAND2 (N856, N852, N678);
nand NAND3 (N857, N816, N182, N269);
not NOT1 (N858, N857);
xor XOR2 (N859, N854, N584);
and AND2 (N860, N844, N285);
buf BUF1 (N861, N853);
not NOT1 (N862, N848);
not NOT1 (N863, N860);
xor XOR2 (N864, N862, N246);
or OR4 (N865, N850, N490, N735, N684);
nor NOR2 (N866, N851, N315);
not NOT1 (N867, N855);
and AND3 (N868, N863, N401, N200);
buf BUF1 (N869, N846);
and AND2 (N870, N861, N448);
or OR4 (N871, N864, N718, N180, N801);
nand NAND3 (N872, N871, N625, N620);
and AND2 (N873, N866, N119);
or OR4 (N874, N856, N159, N254, N422);
xor XOR2 (N875, N867, N516);
buf BUF1 (N876, N858);
nor NOR3 (N877, N859, N270, N205);
nand NAND4 (N878, N875, N216, N201, N695);
xor XOR2 (N879, N870, N503);
xor XOR2 (N880, N868, N121);
buf BUF1 (N881, N880);
xor XOR2 (N882, N876, N855);
and AND4 (N883, N879, N863, N768, N739);
and AND3 (N884, N881, N748, N2);
xor XOR2 (N885, N882, N192);
nand NAND4 (N886, N884, N411, N860, N175);
nor NOR2 (N887, N872, N885);
nand NAND2 (N888, N856, N17);
nor NOR4 (N889, N877, N550, N870, N424);
xor XOR2 (N890, N865, N722);
nor NOR2 (N891, N874, N159);
or OR2 (N892, N889, N82);
nand NAND2 (N893, N873, N174);
not NOT1 (N894, N890);
nand NAND2 (N895, N888, N665);
buf BUF1 (N896, N883);
nor NOR4 (N897, N894, N655, N543, N242);
not NOT1 (N898, N895);
not NOT1 (N899, N886);
not NOT1 (N900, N887);
nand NAND3 (N901, N896, N20, N516);
and AND4 (N902, N893, N284, N32, N771);
nor NOR3 (N903, N901, N381, N119);
buf BUF1 (N904, N869);
not NOT1 (N905, N891);
xor XOR2 (N906, N878, N178);
and AND2 (N907, N906, N726);
nand NAND4 (N908, N897, N100, N512, N814);
xor XOR2 (N909, N892, N747);
xor XOR2 (N910, N898, N644);
xor XOR2 (N911, N902, N344);
buf BUF1 (N912, N907);
not NOT1 (N913, N912);
buf BUF1 (N914, N913);
nand NAND4 (N915, N914, N622, N240, N467);
xor XOR2 (N916, N908, N364);
nand NAND3 (N917, N903, N734, N375);
not NOT1 (N918, N915);
buf BUF1 (N919, N904);
buf BUF1 (N920, N919);
nand NAND4 (N921, N905, N327, N764, N678);
or OR2 (N922, N916, N100);
buf BUF1 (N923, N921);
nand NAND4 (N924, N917, N916, N440, N89);
nor NOR3 (N925, N923, N534, N133);
nand NAND4 (N926, N925, N751, N205, N364);
not NOT1 (N927, N899);
nand NAND4 (N928, N918, N194, N526, N299);
buf BUF1 (N929, N926);
nand NAND3 (N930, N911, N449, N653);
and AND3 (N931, N920, N389, N216);
or OR3 (N932, N927, N742, N10);
and AND3 (N933, N928, N547, N541);
and AND4 (N934, N910, N886, N526, N836);
nand NAND3 (N935, N929, N154, N409);
not NOT1 (N936, N900);
nand NAND2 (N937, N936, N776);
buf BUF1 (N938, N909);
and AND2 (N939, N924, N843);
not NOT1 (N940, N939);
and AND4 (N941, N933, N772, N539, N342);
and AND2 (N942, N937, N430);
not NOT1 (N943, N931);
xor XOR2 (N944, N943, N317);
not NOT1 (N945, N935);
and AND4 (N946, N940, N867, N555, N234);
buf BUF1 (N947, N932);
nor NOR4 (N948, N938, N307, N328, N703);
nor NOR3 (N949, N934, N561, N891);
buf BUF1 (N950, N922);
not NOT1 (N951, N947);
or OR3 (N952, N951, N51, N298);
not NOT1 (N953, N941);
not NOT1 (N954, N944);
or OR3 (N955, N954, N186, N467);
buf BUF1 (N956, N950);
nor NOR3 (N957, N945, N212, N313);
xor XOR2 (N958, N957, N328);
not NOT1 (N959, N942);
not NOT1 (N960, N946);
nor NOR3 (N961, N958, N500, N546);
nand NAND3 (N962, N948, N151, N399);
not NOT1 (N963, N961);
or OR4 (N964, N956, N806, N81, N703);
not NOT1 (N965, N952);
and AND3 (N966, N962, N531, N360);
nor NOR4 (N967, N960, N637, N509, N381);
and AND4 (N968, N967, N778, N116, N675);
nor NOR4 (N969, N966, N214, N898, N780);
not NOT1 (N970, N953);
and AND2 (N971, N969, N489);
buf BUF1 (N972, N968);
and AND3 (N973, N949, N249, N330);
xor XOR2 (N974, N964, N121);
nor NOR2 (N975, N973, N337);
and AND4 (N976, N974, N721, N344, N960);
xor XOR2 (N977, N976, N79);
nand NAND2 (N978, N965, N229);
not NOT1 (N979, N955);
not NOT1 (N980, N970);
and AND3 (N981, N971, N20, N29);
nor NOR2 (N982, N972, N311);
nor NOR3 (N983, N982, N668, N233);
xor XOR2 (N984, N983, N870);
xor XOR2 (N985, N979, N558);
not NOT1 (N986, N930);
xor XOR2 (N987, N959, N162);
or OR2 (N988, N987, N495);
and AND3 (N989, N988, N723, N709);
not NOT1 (N990, N985);
xor XOR2 (N991, N975, N304);
nor NOR4 (N992, N990, N116, N891, N771);
xor XOR2 (N993, N992, N822);
buf BUF1 (N994, N989);
xor XOR2 (N995, N993, N312);
and AND4 (N996, N995, N502, N584, N658);
and AND2 (N997, N986, N858);
nand NAND2 (N998, N963, N972);
xor XOR2 (N999, N997, N349);
xor XOR2 (N1000, N991, N642);
not NOT1 (N1001, N980);
nor NOR4 (N1002, N981, N609, N139, N446);
or OR4 (N1003, N1001, N303, N167, N678);
and AND4 (N1004, N984, N770, N575, N207);
and AND3 (N1005, N998, N323, N1001);
not NOT1 (N1006, N996);
nand NAND2 (N1007, N1004, N110);
and AND4 (N1008, N1005, N594, N656, N869);
or OR3 (N1009, N994, N776, N751);
xor XOR2 (N1010, N1006, N672);
and AND3 (N1011, N1009, N248, N819);
nor NOR4 (N1012, N1011, N17, N837, N642);
xor XOR2 (N1013, N1002, N105);
nor NOR4 (N1014, N1010, N456, N919, N88);
xor XOR2 (N1015, N1014, N862);
buf BUF1 (N1016, N978);
or OR2 (N1017, N1013, N619);
nand NAND3 (N1018, N1007, N781, N79);
not NOT1 (N1019, N1015);
nand NAND3 (N1020, N999, N7, N969);
buf BUF1 (N1021, N1016);
or OR4 (N1022, N1021, N588, N430, N794);
buf BUF1 (N1023, N1017);
buf BUF1 (N1024, N1023);
or OR2 (N1025, N1003, N550);
buf BUF1 (N1026, N1022);
buf BUF1 (N1027, N1000);
or OR2 (N1028, N1018, N372);
and AND3 (N1029, N1028, N585, N254);
and AND3 (N1030, N1025, N952, N308);
and AND3 (N1031, N1027, N917, N239);
xor XOR2 (N1032, N1024, N449);
nor NOR3 (N1033, N1012, N800, N965);
buf BUF1 (N1034, N1019);
buf BUF1 (N1035, N1026);
xor XOR2 (N1036, N1030, N950);
buf BUF1 (N1037, N1032);
nand NAND2 (N1038, N1031, N639);
xor XOR2 (N1039, N1033, N228);
nand NAND3 (N1040, N1038, N643, N341);
nor NOR2 (N1041, N977, N354);
and AND2 (N1042, N1029, N80);
or OR2 (N1043, N1020, N333);
or OR4 (N1044, N1036, N122, N852, N35);
not NOT1 (N1045, N1043);
or OR2 (N1046, N1008, N757);
and AND4 (N1047, N1039, N679, N391, N828);
not NOT1 (N1048, N1037);
xor XOR2 (N1049, N1034, N847);
not NOT1 (N1050, N1049);
and AND4 (N1051, N1050, N733, N409, N786);
buf BUF1 (N1052, N1040);
or OR3 (N1053, N1045, N196, N108);
nor NOR3 (N1054, N1046, N749, N684);
nand NAND3 (N1055, N1044, N885, N334);
not NOT1 (N1056, N1052);
nand NAND4 (N1057, N1042, N239, N17, N967);
xor XOR2 (N1058, N1053, N816);
or OR2 (N1059, N1057, N703);
or OR3 (N1060, N1041, N303, N907);
nor NOR4 (N1061, N1051, N433, N953, N1038);
nand NAND3 (N1062, N1048, N184, N20);
buf BUF1 (N1063, N1054);
buf BUF1 (N1064, N1047);
nor NOR2 (N1065, N1063, N866);
and AND3 (N1066, N1064, N312, N542);
buf BUF1 (N1067, N1056);
not NOT1 (N1068, N1066);
nand NAND3 (N1069, N1055, N107, N458);
not NOT1 (N1070, N1058);
not NOT1 (N1071, N1069);
not NOT1 (N1072, N1068);
or OR3 (N1073, N1061, N696, N807);
or OR4 (N1074, N1060, N347, N1043, N257);
or OR3 (N1075, N1035, N1064, N235);
not NOT1 (N1076, N1072);
buf BUF1 (N1077, N1067);
xor XOR2 (N1078, N1073, N440);
not NOT1 (N1079, N1071);
or OR3 (N1080, N1078, N209, N779);
nor NOR2 (N1081, N1062, N840);
buf BUF1 (N1082, N1077);
nor NOR2 (N1083, N1076, N342);
and AND3 (N1084, N1083, N407, N206);
nand NAND3 (N1085, N1059, N342, N760);
buf BUF1 (N1086, N1080);
or OR4 (N1087, N1075, N171, N267, N421);
nand NAND4 (N1088, N1081, N385, N693, N328);
and AND4 (N1089, N1082, N127, N382, N549);
not NOT1 (N1090, N1085);
xor XOR2 (N1091, N1065, N438);
and AND2 (N1092, N1074, N41);
not NOT1 (N1093, N1088);
nand NAND2 (N1094, N1093, N880);
or OR4 (N1095, N1092, N847, N611, N387);
buf BUF1 (N1096, N1089);
not NOT1 (N1097, N1096);
buf BUF1 (N1098, N1084);
nand NAND4 (N1099, N1098, N560, N403, N102);
or OR2 (N1100, N1086, N1059);
xor XOR2 (N1101, N1090, N900);
or OR4 (N1102, N1097, N50, N596, N562);
nor NOR4 (N1103, N1100, N570, N734, N263);
not NOT1 (N1104, N1095);
xor XOR2 (N1105, N1079, N359);
or OR4 (N1106, N1102, N527, N511, N865);
nand NAND4 (N1107, N1099, N439, N681, N29);
and AND3 (N1108, N1105, N906, N850);
not NOT1 (N1109, N1094);
nor NOR2 (N1110, N1109, N1013);
or OR4 (N1111, N1070, N940, N218, N609);
not NOT1 (N1112, N1104);
not NOT1 (N1113, N1112);
nand NAND4 (N1114, N1107, N1012, N467, N1083);
and AND3 (N1115, N1106, N999, N42);
xor XOR2 (N1116, N1110, N1098);
buf BUF1 (N1117, N1115);
or OR3 (N1118, N1103, N466, N420);
nor NOR2 (N1119, N1101, N999);
xor XOR2 (N1120, N1108, N20);
buf BUF1 (N1121, N1118);
not NOT1 (N1122, N1114);
nor NOR2 (N1123, N1111, N1107);
or OR2 (N1124, N1122, N893);
xor XOR2 (N1125, N1116, N246);
nand NAND4 (N1126, N1123, N902, N265, N1003);
buf BUF1 (N1127, N1091);
nor NOR4 (N1128, N1126, N1, N796, N975);
or OR4 (N1129, N1125, N534, N561, N728);
or OR4 (N1130, N1087, N1026, N264, N422);
buf BUF1 (N1131, N1129);
nand NAND4 (N1132, N1121, N375, N628, N157);
nand NAND3 (N1133, N1119, N122, N1054);
or OR4 (N1134, N1130, N341, N1109, N243);
and AND3 (N1135, N1120, N1085, N1022);
and AND3 (N1136, N1132, N64, N913);
buf BUF1 (N1137, N1135);
nor NOR2 (N1138, N1131, N417);
or OR4 (N1139, N1113, N183, N523, N79);
nand NAND3 (N1140, N1127, N122, N961);
or OR4 (N1141, N1138, N571, N625, N158);
not NOT1 (N1142, N1128);
nand NAND3 (N1143, N1136, N480, N866);
and AND4 (N1144, N1133, N348, N571, N281);
xor XOR2 (N1145, N1134, N72);
buf BUF1 (N1146, N1143);
and AND2 (N1147, N1137, N417);
buf BUF1 (N1148, N1140);
buf BUF1 (N1149, N1139);
not NOT1 (N1150, N1147);
xor XOR2 (N1151, N1142, N1011);
not NOT1 (N1152, N1117);
and AND2 (N1153, N1148, N935);
and AND4 (N1154, N1124, N97, N461, N622);
nand NAND3 (N1155, N1150, N1080, N4);
nor NOR2 (N1156, N1155, N697);
not NOT1 (N1157, N1145);
xor XOR2 (N1158, N1156, N465);
nand NAND4 (N1159, N1152, N755, N248, N98);
nor NOR2 (N1160, N1149, N433);
and AND3 (N1161, N1158, N73, N990);
and AND4 (N1162, N1161, N156, N100, N505);
xor XOR2 (N1163, N1159, N544);
buf BUF1 (N1164, N1153);
nor NOR4 (N1165, N1154, N61, N506, N703);
not NOT1 (N1166, N1141);
or OR3 (N1167, N1157, N268, N412);
and AND2 (N1168, N1160, N119);
nor NOR3 (N1169, N1166, N524, N1160);
nor NOR3 (N1170, N1162, N470, N554);
nand NAND4 (N1171, N1169, N596, N1046, N906);
nand NAND4 (N1172, N1164, N636, N178, N117);
not NOT1 (N1173, N1168);
buf BUF1 (N1174, N1173);
buf BUF1 (N1175, N1151);
not NOT1 (N1176, N1171);
nor NOR4 (N1177, N1167, N177, N1093, N927);
nand NAND2 (N1178, N1170, N179);
nor NOR3 (N1179, N1178, N427, N1135);
buf BUF1 (N1180, N1146);
xor XOR2 (N1181, N1179, N1148);
and AND2 (N1182, N1172, N982);
nor NOR3 (N1183, N1144, N322, N659);
nand NAND4 (N1184, N1176, N980, N350, N522);
xor XOR2 (N1185, N1174, N682);
not NOT1 (N1186, N1183);
not NOT1 (N1187, N1180);
not NOT1 (N1188, N1186);
xor XOR2 (N1189, N1187, N367);
not NOT1 (N1190, N1181);
nand NAND3 (N1191, N1189, N676, N83);
and AND3 (N1192, N1184, N1180, N67);
buf BUF1 (N1193, N1185);
nor NOR3 (N1194, N1192, N785, N1076);
or OR2 (N1195, N1188, N459);
nor NOR3 (N1196, N1182, N868, N776);
not NOT1 (N1197, N1191);
nor NOR4 (N1198, N1163, N429, N299, N50);
xor XOR2 (N1199, N1190, N805);
buf BUF1 (N1200, N1196);
xor XOR2 (N1201, N1198, N237);
and AND2 (N1202, N1175, N1046);
buf BUF1 (N1203, N1194);
or OR3 (N1204, N1193, N266, N772);
and AND2 (N1205, N1177, N400);
buf BUF1 (N1206, N1205);
or OR4 (N1207, N1204, N861, N705, N484);
and AND2 (N1208, N1207, N372);
nand NAND4 (N1209, N1195, N927, N312, N586);
and AND4 (N1210, N1206, N743, N546, N383);
buf BUF1 (N1211, N1165);
not NOT1 (N1212, N1211);
buf BUF1 (N1213, N1201);
not NOT1 (N1214, N1200);
xor XOR2 (N1215, N1202, N31);
xor XOR2 (N1216, N1215, N390);
not NOT1 (N1217, N1203);
xor XOR2 (N1218, N1197, N1079);
buf BUF1 (N1219, N1212);
nor NOR4 (N1220, N1199, N1152, N594, N315);
buf BUF1 (N1221, N1213);
not NOT1 (N1222, N1217);
and AND4 (N1223, N1218, N681, N1200, N506);
not NOT1 (N1224, N1216);
buf BUF1 (N1225, N1223);
and AND3 (N1226, N1222, N1109, N798);
nor NOR3 (N1227, N1208, N31, N288);
nand NAND3 (N1228, N1224, N691, N215);
nand NAND3 (N1229, N1214, N778, N289);
xor XOR2 (N1230, N1219, N625);
buf BUF1 (N1231, N1221);
not NOT1 (N1232, N1220);
or OR3 (N1233, N1229, N795, N1035);
nor NOR3 (N1234, N1231, N305, N233);
xor XOR2 (N1235, N1234, N321);
buf BUF1 (N1236, N1232);
or OR2 (N1237, N1209, N1009);
buf BUF1 (N1238, N1210);
or OR3 (N1239, N1235, N1009, N1061);
nor NOR3 (N1240, N1230, N636, N1101);
nor NOR3 (N1241, N1227, N361, N622);
and AND4 (N1242, N1238, N61, N693, N152);
nand NAND3 (N1243, N1226, N820, N438);
not NOT1 (N1244, N1228);
and AND3 (N1245, N1241, N1109, N135);
not NOT1 (N1246, N1243);
and AND2 (N1247, N1244, N820);
not NOT1 (N1248, N1246);
nor NOR4 (N1249, N1239, N1119, N888, N108);
nor NOR4 (N1250, N1233, N1064, N912, N132);
nor NOR4 (N1251, N1245, N462, N345, N1144);
xor XOR2 (N1252, N1248, N543);
not NOT1 (N1253, N1240);
nand NAND2 (N1254, N1247, N937);
nand NAND3 (N1255, N1236, N352, N1232);
or OR2 (N1256, N1225, N1033);
and AND3 (N1257, N1251, N1120, N59);
nand NAND3 (N1258, N1257, N306, N422);
or OR3 (N1259, N1242, N835, N268);
not NOT1 (N1260, N1249);
or OR2 (N1261, N1253, N1189);
and AND2 (N1262, N1252, N966);
or OR4 (N1263, N1258, N1140, N893, N331);
buf BUF1 (N1264, N1259);
buf BUF1 (N1265, N1237);
and AND3 (N1266, N1255, N219, N1231);
buf BUF1 (N1267, N1262);
buf BUF1 (N1268, N1261);
nor NOR2 (N1269, N1265, N227);
nor NOR4 (N1270, N1263, N1124, N431, N567);
nor NOR4 (N1271, N1256, N601, N759, N358);
nand NAND4 (N1272, N1264, N10, N26, N1246);
not NOT1 (N1273, N1266);
not NOT1 (N1274, N1254);
xor XOR2 (N1275, N1273, N408);
nand NAND2 (N1276, N1270, N1248);
xor XOR2 (N1277, N1260, N362);
not NOT1 (N1278, N1250);
xor XOR2 (N1279, N1275, N616);
not NOT1 (N1280, N1269);
and AND2 (N1281, N1279, N1089);
nand NAND4 (N1282, N1278, N627, N1244, N216);
buf BUF1 (N1283, N1268);
not NOT1 (N1284, N1280);
nor NOR3 (N1285, N1277, N343, N230);
buf BUF1 (N1286, N1267);
nand NAND2 (N1287, N1285, N571);
nor NOR4 (N1288, N1281, N787, N159, N1105);
buf BUF1 (N1289, N1287);
and AND4 (N1290, N1272, N403, N474, N806);
xor XOR2 (N1291, N1289, N309);
buf BUF1 (N1292, N1284);
nor NOR4 (N1293, N1288, N1048, N1264, N144);
nor NOR2 (N1294, N1274, N782);
not NOT1 (N1295, N1293);
not NOT1 (N1296, N1282);
and AND3 (N1297, N1291, N310, N1098);
nor NOR2 (N1298, N1283, N829);
buf BUF1 (N1299, N1295);
not NOT1 (N1300, N1271);
xor XOR2 (N1301, N1276, N665);
and AND4 (N1302, N1296, N1022, N227, N508);
not NOT1 (N1303, N1294);
nand NAND2 (N1304, N1301, N793);
xor XOR2 (N1305, N1302, N758);
nor NOR3 (N1306, N1299, N1149, N498);
not NOT1 (N1307, N1297);
or OR2 (N1308, N1305, N861);
not NOT1 (N1309, N1307);
nand NAND4 (N1310, N1286, N676, N1219, N221);
xor XOR2 (N1311, N1292, N511);
xor XOR2 (N1312, N1303, N204);
buf BUF1 (N1313, N1308);
not NOT1 (N1314, N1310);
and AND3 (N1315, N1304, N644, N487);
or OR3 (N1316, N1300, N689, N1278);
and AND4 (N1317, N1313, N163, N268, N834);
or OR4 (N1318, N1298, N67, N1004, N568);
nand NAND2 (N1319, N1309, N812);
buf BUF1 (N1320, N1306);
nor NOR4 (N1321, N1320, N1218, N808, N985);
nand NAND3 (N1322, N1316, N369, N11);
or OR3 (N1323, N1318, N988, N349);
nand NAND3 (N1324, N1322, N660, N1092);
xor XOR2 (N1325, N1321, N1256);
or OR4 (N1326, N1323, N579, N934, N914);
nor NOR2 (N1327, N1319, N1239);
or OR4 (N1328, N1312, N45, N702, N1231);
and AND3 (N1329, N1326, N837, N501);
or OR4 (N1330, N1315, N1247, N441, N738);
and AND2 (N1331, N1330, N1257);
nand NAND4 (N1332, N1331, N395, N31, N138);
buf BUF1 (N1333, N1317);
buf BUF1 (N1334, N1325);
and AND4 (N1335, N1311, N1333, N1182, N1258);
not NOT1 (N1336, N16);
not NOT1 (N1337, N1327);
and AND3 (N1338, N1336, N163, N1188);
and AND3 (N1339, N1332, N904, N744);
buf BUF1 (N1340, N1290);
not NOT1 (N1341, N1329);
and AND3 (N1342, N1337, N1233, N456);
buf BUF1 (N1343, N1338);
not NOT1 (N1344, N1343);
nor NOR4 (N1345, N1324, N431, N1288, N31);
xor XOR2 (N1346, N1314, N1260);
buf BUF1 (N1347, N1346);
xor XOR2 (N1348, N1335, N488);
xor XOR2 (N1349, N1341, N470);
not NOT1 (N1350, N1328);
not NOT1 (N1351, N1344);
not NOT1 (N1352, N1347);
or OR4 (N1353, N1352, N496, N392, N659);
not NOT1 (N1354, N1334);
nand NAND4 (N1355, N1345, N1094, N1069, N445);
xor XOR2 (N1356, N1355, N116);
and AND2 (N1357, N1356, N1316);
buf BUF1 (N1358, N1348);
nor NOR3 (N1359, N1354, N206, N46);
xor XOR2 (N1360, N1342, N894);
nand NAND3 (N1361, N1350, N684, N711);
and AND2 (N1362, N1353, N421);
buf BUF1 (N1363, N1357);
and AND3 (N1364, N1358, N722, N941);
nor NOR2 (N1365, N1349, N1074);
not NOT1 (N1366, N1363);
or OR3 (N1367, N1340, N1338, N587);
nand NAND3 (N1368, N1339, N745, N978);
xor XOR2 (N1369, N1367, N111);
or OR2 (N1370, N1351, N784);
nor NOR2 (N1371, N1361, N658);
nor NOR2 (N1372, N1370, N262);
xor XOR2 (N1373, N1360, N396);
or OR2 (N1374, N1366, N956);
or OR2 (N1375, N1368, N1003);
nand NAND4 (N1376, N1365, N928, N546, N488);
nand NAND4 (N1377, N1371, N1144, N486, N710);
buf BUF1 (N1378, N1373);
nand NAND2 (N1379, N1362, N827);
nand NAND3 (N1380, N1375, N694, N271);
buf BUF1 (N1381, N1369);
xor XOR2 (N1382, N1372, N398);
or OR4 (N1383, N1364, N279, N418, N10);
nor NOR4 (N1384, N1359, N292, N1304, N431);
nand NAND3 (N1385, N1376, N928, N1342);
and AND4 (N1386, N1381, N1205, N1231, N836);
or OR4 (N1387, N1384, N1033, N308, N1028);
or OR2 (N1388, N1385, N1092);
not NOT1 (N1389, N1383);
nor NOR2 (N1390, N1380, N493);
nor NOR4 (N1391, N1378, N732, N69, N264);
nor NOR3 (N1392, N1389, N902, N691);
xor XOR2 (N1393, N1387, N1149);
and AND2 (N1394, N1374, N264);
or OR4 (N1395, N1390, N668, N847, N1005);
or OR4 (N1396, N1386, N1247, N330, N426);
nand NAND2 (N1397, N1377, N1349);
or OR4 (N1398, N1393, N803, N645, N839);
or OR2 (N1399, N1397, N664);
nor NOR4 (N1400, N1379, N1229, N163, N104);
not NOT1 (N1401, N1395);
buf BUF1 (N1402, N1396);
or OR4 (N1403, N1394, N614, N1079, N683);
and AND3 (N1404, N1388, N928, N497);
xor XOR2 (N1405, N1402, N53);
or OR2 (N1406, N1404, N139);
and AND4 (N1407, N1399, N580, N339, N1142);
and AND2 (N1408, N1382, N621);
and AND4 (N1409, N1407, N1309, N609, N936);
nor NOR3 (N1410, N1400, N869, N219);
not NOT1 (N1411, N1401);
not NOT1 (N1412, N1405);
buf BUF1 (N1413, N1391);
nand NAND4 (N1414, N1410, N86, N808, N1251);
and AND2 (N1415, N1409, N137);
nor NOR3 (N1416, N1412, N317, N1046);
not NOT1 (N1417, N1416);
buf BUF1 (N1418, N1413);
nor NOR4 (N1419, N1417, N253, N74, N261);
nand NAND3 (N1420, N1411, N1043, N144);
nor NOR2 (N1421, N1403, N1148);
xor XOR2 (N1422, N1419, N762);
nand NAND4 (N1423, N1414, N584, N1056, N786);
buf BUF1 (N1424, N1418);
xor XOR2 (N1425, N1415, N1408);
buf BUF1 (N1426, N142);
nor NOR4 (N1427, N1426, N724, N746, N466);
not NOT1 (N1428, N1427);
nor NOR4 (N1429, N1392, N108, N146, N15);
nand NAND4 (N1430, N1406, N1357, N1401, N373);
nand NAND2 (N1431, N1422, N574);
and AND2 (N1432, N1423, N652);
not NOT1 (N1433, N1420);
buf BUF1 (N1434, N1429);
and AND2 (N1435, N1398, N750);
xor XOR2 (N1436, N1431, N304);
not NOT1 (N1437, N1421);
nor NOR3 (N1438, N1432, N982, N1353);
nor NOR2 (N1439, N1428, N11);
nand NAND2 (N1440, N1430, N590);
or OR2 (N1441, N1435, N895);
nand NAND4 (N1442, N1438, N1078, N388, N44);
nor NOR2 (N1443, N1442, N384);
or OR3 (N1444, N1436, N291, N1205);
nor NOR3 (N1445, N1433, N1396, N1157);
buf BUF1 (N1446, N1437);
nor NOR4 (N1447, N1445, N805, N813, N1172);
nand NAND4 (N1448, N1424, N151, N1325, N892);
buf BUF1 (N1449, N1434);
xor XOR2 (N1450, N1440, N834);
nand NAND4 (N1451, N1441, N1008, N1161, N952);
not NOT1 (N1452, N1451);
buf BUF1 (N1453, N1439);
buf BUF1 (N1454, N1425);
buf BUF1 (N1455, N1444);
or OR3 (N1456, N1446, N723, N1263);
xor XOR2 (N1457, N1456, N1394);
nor NOR3 (N1458, N1453, N1336, N849);
xor XOR2 (N1459, N1454, N1045);
and AND2 (N1460, N1447, N572);
not NOT1 (N1461, N1457);
or OR3 (N1462, N1455, N1088, N1166);
nor NOR2 (N1463, N1459, N772);
nand NAND2 (N1464, N1458, N497);
nand NAND2 (N1465, N1448, N426);
or OR2 (N1466, N1450, N85);
or OR4 (N1467, N1465, N786, N221, N1002);
xor XOR2 (N1468, N1443, N483);
nand NAND4 (N1469, N1462, N564, N1378, N1125);
and AND4 (N1470, N1463, N1438, N925, N394);
not NOT1 (N1471, N1460);
nor NOR4 (N1472, N1452, N1006, N816, N1434);
buf BUF1 (N1473, N1471);
xor XOR2 (N1474, N1466, N793);
nor NOR3 (N1475, N1470, N1096, N747);
nor NOR2 (N1476, N1461, N945);
nor NOR4 (N1477, N1475, N1455, N39, N749);
nand NAND2 (N1478, N1477, N440);
not NOT1 (N1479, N1478);
or OR3 (N1480, N1468, N225, N45);
not NOT1 (N1481, N1479);
nor NOR2 (N1482, N1480, N1455);
nor NOR3 (N1483, N1481, N212, N249);
nor NOR2 (N1484, N1482, N108);
or OR4 (N1485, N1467, N323, N431, N689);
xor XOR2 (N1486, N1483, N1457);
not NOT1 (N1487, N1486);
not NOT1 (N1488, N1474);
buf BUF1 (N1489, N1473);
buf BUF1 (N1490, N1449);
nor NOR2 (N1491, N1490, N117);
and AND3 (N1492, N1487, N310, N1466);
nand NAND2 (N1493, N1472, N734);
and AND2 (N1494, N1493, N146);
and AND4 (N1495, N1469, N352, N123, N1223);
buf BUF1 (N1496, N1488);
not NOT1 (N1497, N1491);
nor NOR3 (N1498, N1464, N816, N130);
nor NOR2 (N1499, N1485, N631);
or OR4 (N1500, N1494, N1181, N1275, N1434);
or OR3 (N1501, N1498, N20, N876);
and AND3 (N1502, N1492, N1386, N1094);
nor NOR4 (N1503, N1484, N411, N1375, N33);
buf BUF1 (N1504, N1496);
buf BUF1 (N1505, N1476);
xor XOR2 (N1506, N1505, N747);
and AND2 (N1507, N1504, N1316);
nand NAND2 (N1508, N1499, N832);
and AND2 (N1509, N1497, N810);
nand NAND4 (N1510, N1489, N280, N1176, N1413);
and AND3 (N1511, N1495, N853, N1438);
buf BUF1 (N1512, N1511);
buf BUF1 (N1513, N1507);
and AND3 (N1514, N1500, N68, N349);
nor NOR3 (N1515, N1513, N811, N528);
not NOT1 (N1516, N1502);
or OR3 (N1517, N1515, N787, N580);
endmodule