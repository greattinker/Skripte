// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N890,N910,N906,N918,N915,N919,N917,N913,N916,N920;

nand NAND3 (N21, N12, N4, N18);
not NOT1 (N22, N13);
xor XOR2 (N23, N17, N8);
and AND4 (N24, N1, N12, N23, N8);
nand NAND3 (N25, N22, N24, N1);
and AND3 (N26, N12, N20, N3);
and AND4 (N27, N7, N21, N24, N6);
buf BUF1 (N28, N9);
nor NOR3 (N29, N6, N9, N15);
nand NAND3 (N30, N18, N28, N16);
buf BUF1 (N31, N9);
not NOT1 (N32, N3);
buf BUF1 (N33, N22);
or OR3 (N34, N13, N17, N17);
or OR2 (N35, N33, N10);
not NOT1 (N36, N16);
xor XOR2 (N37, N30, N20);
not NOT1 (N38, N35);
not NOT1 (N39, N29);
xor XOR2 (N40, N39, N24);
xor XOR2 (N41, N25, N6);
xor XOR2 (N42, N26, N38);
xor XOR2 (N43, N37, N30);
and AND2 (N44, N2, N27);
buf BUF1 (N45, N21);
and AND2 (N46, N40, N3);
nor NOR2 (N47, N32, N39);
nor NOR2 (N48, N45, N30);
nand NAND4 (N49, N42, N42, N8, N35);
not NOT1 (N50, N46);
or OR3 (N51, N44, N4, N18);
and AND2 (N52, N51, N23);
buf BUF1 (N53, N47);
not NOT1 (N54, N49);
not NOT1 (N55, N43);
nand NAND4 (N56, N48, N44, N41, N42);
not NOT1 (N57, N34);
not NOT1 (N58, N46);
nor NOR2 (N59, N57, N36);
xor XOR2 (N60, N21, N36);
not NOT1 (N61, N52);
and AND4 (N62, N54, N12, N39, N1);
nor NOR4 (N63, N61, N14, N16, N44);
not NOT1 (N64, N63);
not NOT1 (N65, N60);
not NOT1 (N66, N56);
xor XOR2 (N67, N50, N7);
xor XOR2 (N68, N55, N31);
not NOT1 (N69, N14);
nand NAND2 (N70, N65, N52);
not NOT1 (N71, N59);
nand NAND4 (N72, N64, N33, N69, N34);
xor XOR2 (N73, N67, N36);
and AND4 (N74, N31, N71, N59, N72);
xor XOR2 (N75, N52, N39);
nor NOR2 (N76, N11, N42);
and AND2 (N77, N76, N2);
xor XOR2 (N78, N77, N76);
or OR3 (N79, N73, N34, N44);
or OR2 (N80, N70, N36);
buf BUF1 (N81, N80);
xor XOR2 (N82, N53, N60);
or OR4 (N83, N79, N67, N73, N37);
xor XOR2 (N84, N75, N72);
nor NOR2 (N85, N84, N64);
or OR3 (N86, N66, N70, N52);
xor XOR2 (N87, N85, N18);
and AND2 (N88, N83, N41);
xor XOR2 (N89, N81, N36);
nand NAND4 (N90, N89, N83, N49, N84);
buf BUF1 (N91, N88);
not NOT1 (N92, N86);
not NOT1 (N93, N92);
nand NAND2 (N94, N87, N81);
or OR2 (N95, N62, N5);
xor XOR2 (N96, N95, N38);
not NOT1 (N97, N96);
xor XOR2 (N98, N82, N20);
not NOT1 (N99, N94);
xor XOR2 (N100, N91, N38);
and AND4 (N101, N78, N18, N6, N61);
not NOT1 (N102, N101);
buf BUF1 (N103, N93);
or OR4 (N104, N90, N13, N99, N54);
not NOT1 (N105, N80);
and AND3 (N106, N100, N46, N43);
nand NAND3 (N107, N68, N57, N51);
and AND4 (N108, N98, N33, N33, N102);
not NOT1 (N109, N6);
xor XOR2 (N110, N58, N11);
xor XOR2 (N111, N105, N110);
nor NOR3 (N112, N110, N44, N55);
nor NOR4 (N113, N112, N71, N25, N54);
xor XOR2 (N114, N111, N82);
nand NAND3 (N115, N109, N20, N41);
nor NOR3 (N116, N108, N5, N113);
nand NAND3 (N117, N48, N24, N27);
and AND2 (N118, N115, N103);
nor NOR3 (N119, N74, N70, N56);
and AND4 (N120, N91, N40, N92, N104);
or OR3 (N121, N90, N71, N75);
nor NOR4 (N122, N116, N106, N1, N50);
xor XOR2 (N123, N39, N80);
buf BUF1 (N124, N117);
xor XOR2 (N125, N107, N87);
nor NOR4 (N126, N119, N73, N33, N116);
nor NOR3 (N127, N118, N111, N48);
xor XOR2 (N128, N97, N72);
and AND4 (N129, N126, N16, N11, N105);
not NOT1 (N130, N121);
nor NOR4 (N131, N122, N69, N100, N19);
nand NAND3 (N132, N125, N111, N65);
and AND2 (N133, N127, N49);
or OR3 (N134, N129, N25, N81);
nand NAND3 (N135, N128, N126, N34);
nor NOR2 (N136, N132, N66);
buf BUF1 (N137, N130);
not NOT1 (N138, N124);
not NOT1 (N139, N136);
nand NAND2 (N140, N123, N24);
or OR2 (N141, N134, N108);
not NOT1 (N142, N131);
xor XOR2 (N143, N140, N126);
nor NOR2 (N144, N142, N4);
nand NAND3 (N145, N137, N70, N101);
or OR3 (N146, N120, N101, N114);
nand NAND3 (N147, N1, N136, N137);
not NOT1 (N148, N147);
or OR4 (N149, N138, N137, N121, N59);
nand NAND4 (N150, N135, N135, N77, N135);
nor NOR3 (N151, N143, N9, N116);
or OR2 (N152, N148, N147);
xor XOR2 (N153, N146, N117);
and AND4 (N154, N145, N119, N56, N40);
or OR4 (N155, N152, N39, N26, N147);
nand NAND2 (N156, N153, N138);
and AND2 (N157, N156, N22);
buf BUF1 (N158, N151);
nand NAND4 (N159, N139, N9, N76, N5);
nor NOR3 (N160, N149, N56, N69);
xor XOR2 (N161, N157, N29);
or OR3 (N162, N150, N2, N81);
or OR4 (N163, N158, N111, N26, N112);
or OR2 (N164, N159, N155);
not NOT1 (N165, N159);
nor NOR4 (N166, N160, N59, N152, N150);
xor XOR2 (N167, N165, N84);
or OR3 (N168, N164, N27, N77);
nand NAND2 (N169, N166, N3);
and AND2 (N170, N167, N147);
nor NOR3 (N171, N163, N57, N128);
or OR3 (N172, N133, N71, N128);
not NOT1 (N173, N169);
nor NOR4 (N174, N154, N63, N86, N130);
or OR2 (N175, N171, N165);
or OR4 (N176, N174, N34, N7, N170);
and AND4 (N177, N129, N175, N153, N169);
nand NAND4 (N178, N102, N112, N122, N47);
xor XOR2 (N179, N141, N119);
or OR4 (N180, N173, N73, N154, N74);
nor NOR4 (N181, N168, N106, N53, N127);
or OR2 (N182, N176, N133);
xor XOR2 (N183, N178, N1);
and AND2 (N184, N162, N1);
nor NOR3 (N185, N184, N6, N58);
or OR3 (N186, N179, N145, N77);
xor XOR2 (N187, N185, N74);
not NOT1 (N188, N177);
nor NOR3 (N189, N144, N1, N142);
or OR2 (N190, N187, N152);
not NOT1 (N191, N181);
or OR2 (N192, N180, N151);
xor XOR2 (N193, N172, N162);
not NOT1 (N194, N182);
nor NOR4 (N195, N194, N97, N3, N127);
or OR2 (N196, N192, N129);
nand NAND3 (N197, N186, N20, N57);
and AND3 (N198, N161, N28, N56);
nor NOR2 (N199, N195, N167);
or OR4 (N200, N199, N41, N137, N60);
not NOT1 (N201, N196);
nor NOR2 (N202, N198, N52);
and AND3 (N203, N202, N193, N3);
not NOT1 (N204, N153);
nor NOR3 (N205, N203, N101, N51);
or OR4 (N206, N191, N54, N15, N132);
or OR2 (N207, N188, N174);
and AND2 (N208, N183, N36);
nand NAND4 (N209, N197, N19, N194, N123);
xor XOR2 (N210, N207, N5);
nand NAND4 (N211, N189, N103, N173, N136);
buf BUF1 (N212, N201);
buf BUF1 (N213, N211);
buf BUF1 (N214, N209);
xor XOR2 (N215, N204, N190);
buf BUF1 (N216, N155);
nand NAND4 (N217, N208, N148, N58, N49);
xor XOR2 (N218, N216, N185);
xor XOR2 (N219, N210, N96);
or OR3 (N220, N217, N8, N38);
not NOT1 (N221, N206);
nor NOR2 (N222, N200, N71);
nand NAND3 (N223, N214, N149, N72);
or OR4 (N224, N205, N157, N11, N216);
buf BUF1 (N225, N220);
xor XOR2 (N226, N224, N90);
buf BUF1 (N227, N218);
nor NOR3 (N228, N223, N96, N117);
nand NAND4 (N229, N215, N64, N16, N211);
xor XOR2 (N230, N225, N45);
nand NAND4 (N231, N228, N205, N135, N22);
and AND3 (N232, N213, N123, N18);
or OR4 (N233, N221, N214, N27, N86);
nand NAND2 (N234, N231, N167);
not NOT1 (N235, N234);
xor XOR2 (N236, N235, N196);
not NOT1 (N237, N219);
not NOT1 (N238, N237);
not NOT1 (N239, N236);
buf BUF1 (N240, N227);
nor NOR2 (N241, N229, N116);
xor XOR2 (N242, N222, N108);
buf BUF1 (N243, N238);
not NOT1 (N244, N212);
not NOT1 (N245, N241);
not NOT1 (N246, N240);
buf BUF1 (N247, N233);
not NOT1 (N248, N239);
xor XOR2 (N249, N245, N225);
or OR2 (N250, N232, N197);
buf BUF1 (N251, N244);
or OR3 (N252, N243, N144, N22);
nor NOR4 (N253, N248, N92, N93, N175);
nor NOR4 (N254, N246, N211, N55, N99);
xor XOR2 (N255, N230, N245);
nand NAND3 (N256, N226, N194, N179);
xor XOR2 (N257, N250, N81);
nor NOR4 (N258, N255, N115, N179, N233);
buf BUF1 (N259, N251);
not NOT1 (N260, N253);
buf BUF1 (N261, N259);
nand NAND2 (N262, N252, N2);
or OR4 (N263, N258, N242, N101, N32);
and AND4 (N264, N137, N152, N71, N241);
nand NAND3 (N265, N257, N122, N239);
not NOT1 (N266, N263);
nand NAND3 (N267, N249, N166, N142);
nand NAND4 (N268, N254, N127, N18, N250);
buf BUF1 (N269, N260);
nand NAND4 (N270, N268, N99, N124, N197);
and AND4 (N271, N269, N210, N218, N12);
nor NOR3 (N272, N266, N271, N22);
not NOT1 (N273, N225);
buf BUF1 (N274, N256);
buf BUF1 (N275, N272);
xor XOR2 (N276, N261, N272);
nand NAND3 (N277, N267, N127, N267);
or OR2 (N278, N270, N153);
and AND4 (N279, N274, N25, N250, N218);
nor NOR4 (N280, N276, N14, N203, N88);
nor NOR3 (N281, N273, N218, N65);
xor XOR2 (N282, N275, N138);
not NOT1 (N283, N262);
buf BUF1 (N284, N279);
xor XOR2 (N285, N282, N139);
nor NOR3 (N286, N278, N37, N133);
or OR4 (N287, N277, N2, N13, N76);
not NOT1 (N288, N281);
nand NAND4 (N289, N264, N186, N112, N157);
or OR3 (N290, N284, N22, N247);
buf BUF1 (N291, N288);
not NOT1 (N292, N157);
buf BUF1 (N293, N286);
buf BUF1 (N294, N280);
xor XOR2 (N295, N285, N159);
nand NAND4 (N296, N290, N11, N146, N286);
nand NAND3 (N297, N289, N239, N10);
xor XOR2 (N298, N294, N280);
nand NAND2 (N299, N297, N34);
or OR4 (N300, N299, N24, N299, N112);
not NOT1 (N301, N296);
xor XOR2 (N302, N300, N125);
or OR3 (N303, N287, N61, N238);
xor XOR2 (N304, N293, N190);
nand NAND2 (N305, N298, N267);
not NOT1 (N306, N292);
xor XOR2 (N307, N302, N159);
not NOT1 (N308, N305);
or OR2 (N309, N303, N171);
nor NOR4 (N310, N295, N159, N138, N24);
nor NOR2 (N311, N265, N93);
or OR3 (N312, N310, N96, N15);
and AND2 (N313, N304, N242);
nor NOR3 (N314, N312, N92, N62);
or OR2 (N315, N314, N288);
nand NAND3 (N316, N301, N260, N193);
nor NOR2 (N317, N315, N71);
xor XOR2 (N318, N283, N130);
nand NAND3 (N319, N316, N197, N16);
nor NOR2 (N320, N306, N258);
nor NOR3 (N321, N320, N220, N266);
xor XOR2 (N322, N307, N201);
xor XOR2 (N323, N318, N246);
nor NOR4 (N324, N323, N117, N74, N18);
not NOT1 (N325, N319);
nand NAND4 (N326, N325, N276, N184, N72);
buf BUF1 (N327, N291);
nor NOR2 (N328, N308, N40);
nor NOR3 (N329, N322, N86, N85);
buf BUF1 (N330, N326);
or OR2 (N331, N328, N150);
nand NAND4 (N332, N329, N259, N39, N160);
nand NAND2 (N333, N327, N160);
xor XOR2 (N334, N324, N31);
nor NOR2 (N335, N331, N76);
nand NAND3 (N336, N333, N162, N190);
buf BUF1 (N337, N313);
buf BUF1 (N338, N332);
nand NAND2 (N339, N330, N114);
and AND2 (N340, N311, N200);
nor NOR4 (N341, N334, N160, N175, N48);
and AND3 (N342, N336, N260, N313);
nand NAND4 (N343, N338, N62, N103, N206);
nor NOR4 (N344, N341, N46, N204, N279);
or OR4 (N345, N342, N253, N92, N248);
nand NAND4 (N346, N344, N74, N199, N139);
nand NAND4 (N347, N337, N271, N138, N58);
not NOT1 (N348, N339);
not NOT1 (N349, N321);
not NOT1 (N350, N346);
or OR4 (N351, N345, N339, N129, N226);
buf BUF1 (N352, N351);
buf BUF1 (N353, N350);
nor NOR4 (N354, N309, N106, N46, N242);
nand NAND2 (N355, N348, N221);
buf BUF1 (N356, N354);
and AND2 (N357, N356, N119);
or OR4 (N358, N317, N262, N350, N216);
nor NOR2 (N359, N357, N157);
not NOT1 (N360, N335);
and AND4 (N361, N343, N177, N240, N69);
xor XOR2 (N362, N349, N286);
and AND3 (N363, N361, N182, N40);
xor XOR2 (N364, N355, N287);
or OR3 (N365, N358, N274, N90);
and AND4 (N366, N340, N64, N320, N99);
xor XOR2 (N367, N347, N251);
and AND4 (N368, N353, N293, N164, N276);
xor XOR2 (N369, N366, N64);
xor XOR2 (N370, N362, N295);
or OR4 (N371, N360, N294, N146, N289);
xor XOR2 (N372, N368, N262);
nor NOR4 (N373, N365, N304, N254, N360);
nand NAND4 (N374, N372, N152, N160, N230);
nand NAND2 (N375, N374, N66);
xor XOR2 (N376, N375, N234);
or OR4 (N377, N369, N330, N89, N296);
nand NAND4 (N378, N371, N206, N98, N20);
xor XOR2 (N379, N377, N212);
not NOT1 (N380, N363);
and AND3 (N381, N370, N239, N209);
and AND3 (N382, N373, N150, N114);
not NOT1 (N383, N376);
nor NOR2 (N384, N380, N376);
not NOT1 (N385, N384);
not NOT1 (N386, N364);
xor XOR2 (N387, N383, N278);
not NOT1 (N388, N359);
xor XOR2 (N389, N388, N301);
buf BUF1 (N390, N389);
or OR4 (N391, N367, N287, N344, N64);
nor NOR2 (N392, N379, N10);
or OR2 (N393, N378, N318);
nand NAND4 (N394, N387, N27, N7, N340);
and AND2 (N395, N385, N71);
not NOT1 (N396, N393);
nand NAND3 (N397, N392, N212, N308);
xor XOR2 (N398, N382, N145);
nor NOR4 (N399, N396, N226, N332, N310);
nand NAND2 (N400, N394, N231);
nor NOR4 (N401, N386, N38, N334, N92);
not NOT1 (N402, N401);
or OR3 (N403, N381, N25, N61);
buf BUF1 (N404, N352);
or OR4 (N405, N404, N307, N68, N274);
nor NOR3 (N406, N390, N359, N384);
nand NAND4 (N407, N405, N157, N149, N387);
nor NOR2 (N408, N395, N197);
nand NAND4 (N409, N402, N325, N203, N239);
or OR3 (N410, N408, N36, N299);
xor XOR2 (N411, N406, N98);
not NOT1 (N412, N400);
not NOT1 (N413, N403);
xor XOR2 (N414, N413, N104);
or OR3 (N415, N407, N120, N172);
and AND2 (N416, N412, N89);
nand NAND4 (N417, N397, N371, N327, N239);
or OR3 (N418, N399, N414, N213);
not NOT1 (N419, N403);
nand NAND4 (N420, N411, N270, N74, N162);
or OR4 (N421, N415, N222, N377, N199);
nand NAND2 (N422, N421, N173);
nand NAND4 (N423, N418, N296, N271, N66);
xor XOR2 (N424, N422, N81);
or OR3 (N425, N398, N32, N83);
nor NOR2 (N426, N425, N249);
or OR3 (N427, N424, N128, N236);
xor XOR2 (N428, N409, N330);
buf BUF1 (N429, N426);
not NOT1 (N430, N423);
or OR3 (N431, N428, N94, N112);
xor XOR2 (N432, N417, N166);
xor XOR2 (N433, N420, N58);
buf BUF1 (N434, N433);
buf BUF1 (N435, N416);
buf BUF1 (N436, N432);
and AND2 (N437, N436, N231);
nor NOR4 (N438, N410, N107, N81, N233);
xor XOR2 (N439, N438, N385);
nor NOR3 (N440, N427, N428, N354);
not NOT1 (N441, N391);
or OR4 (N442, N437, N348, N24, N104);
and AND2 (N443, N419, N237);
xor XOR2 (N444, N434, N432);
xor XOR2 (N445, N431, N16);
nand NAND2 (N446, N444, N40);
buf BUF1 (N447, N441);
xor XOR2 (N448, N445, N441);
buf BUF1 (N449, N439);
nand NAND4 (N450, N440, N292, N359, N312);
or OR4 (N451, N429, N370, N189, N1);
xor XOR2 (N452, N435, N151);
xor XOR2 (N453, N451, N372);
or OR4 (N454, N452, N372, N280, N380);
nand NAND4 (N455, N443, N221, N55, N329);
nand NAND3 (N456, N442, N217, N241);
xor XOR2 (N457, N456, N188);
and AND4 (N458, N449, N207, N228, N45);
buf BUF1 (N459, N455);
xor XOR2 (N460, N430, N259);
and AND2 (N461, N448, N149);
nor NOR4 (N462, N459, N21, N454, N316);
or OR3 (N463, N363, N132, N152);
nand NAND4 (N464, N460, N319, N138, N255);
xor XOR2 (N465, N453, N431);
nand NAND4 (N466, N461, N20, N8, N169);
or OR2 (N467, N458, N411);
nand NAND3 (N468, N446, N209, N417);
nor NOR4 (N469, N463, N137, N3, N273);
or OR2 (N470, N457, N361);
buf BUF1 (N471, N462);
or OR2 (N472, N447, N191);
nor NOR3 (N473, N472, N72, N267);
or OR3 (N474, N471, N30, N126);
or OR2 (N475, N474, N190);
buf BUF1 (N476, N466);
or OR4 (N477, N465, N417, N260, N273);
and AND3 (N478, N473, N391, N384);
and AND2 (N479, N469, N252);
buf BUF1 (N480, N478);
and AND3 (N481, N470, N411, N194);
not NOT1 (N482, N468);
nand NAND3 (N483, N475, N146, N42);
and AND2 (N484, N450, N111);
and AND2 (N485, N484, N476);
not NOT1 (N486, N481);
nand NAND2 (N487, N320, N261);
nand NAND3 (N488, N479, N102, N436);
buf BUF1 (N489, N483);
and AND3 (N490, N485, N152, N433);
not NOT1 (N491, N467);
buf BUF1 (N492, N482);
not NOT1 (N493, N464);
buf BUF1 (N494, N487);
and AND3 (N495, N488, N383, N73);
buf BUF1 (N496, N489);
or OR4 (N497, N480, N473, N159, N9);
xor XOR2 (N498, N477, N216);
or OR3 (N499, N493, N367, N179);
xor XOR2 (N500, N499, N193);
buf BUF1 (N501, N500);
xor XOR2 (N502, N495, N349);
xor XOR2 (N503, N490, N260);
nor NOR3 (N504, N501, N324, N400);
xor XOR2 (N505, N502, N467);
xor XOR2 (N506, N494, N290);
nor NOR2 (N507, N506, N425);
not NOT1 (N508, N505);
and AND2 (N509, N504, N293);
and AND4 (N510, N492, N483, N306, N160);
buf BUF1 (N511, N508);
and AND4 (N512, N496, N174, N502, N374);
or OR4 (N513, N511, N225, N223, N280);
buf BUF1 (N514, N503);
or OR2 (N515, N514, N410);
nand NAND3 (N516, N513, N428, N109);
xor XOR2 (N517, N498, N347);
xor XOR2 (N518, N515, N35);
buf BUF1 (N519, N509);
and AND4 (N520, N519, N56, N265, N243);
xor XOR2 (N521, N486, N256);
nand NAND4 (N522, N507, N63, N153, N249);
xor XOR2 (N523, N520, N441);
nor NOR4 (N524, N522, N327, N463, N518);
buf BUF1 (N525, N320);
nor NOR3 (N526, N525, N15, N401);
and AND3 (N527, N512, N212, N182);
nor NOR4 (N528, N524, N290, N24, N397);
nand NAND4 (N529, N510, N450, N98, N314);
and AND2 (N530, N497, N1);
nor NOR2 (N531, N521, N255);
or OR3 (N532, N523, N5, N485);
or OR2 (N533, N526, N111);
nor NOR2 (N534, N533, N531);
or OR4 (N535, N144, N342, N44, N107);
buf BUF1 (N536, N534);
buf BUF1 (N537, N532);
nor NOR3 (N538, N517, N332, N439);
or OR4 (N539, N530, N265, N302, N494);
xor XOR2 (N540, N536, N106);
buf BUF1 (N541, N539);
or OR4 (N542, N540, N458, N493, N131);
xor XOR2 (N543, N537, N97);
buf BUF1 (N544, N527);
nor NOR2 (N545, N544, N13);
or OR2 (N546, N543, N388);
not NOT1 (N547, N546);
nand NAND3 (N548, N545, N238, N5);
or OR2 (N549, N541, N252);
nand NAND2 (N550, N516, N8);
and AND3 (N551, N547, N93, N252);
xor XOR2 (N552, N529, N18);
and AND2 (N553, N535, N292);
or OR3 (N554, N549, N62, N203);
nand NAND4 (N555, N551, N535, N157, N547);
xor XOR2 (N556, N548, N498);
or OR3 (N557, N550, N57, N166);
or OR4 (N558, N528, N511, N267, N348);
or OR4 (N559, N557, N416, N88, N60);
buf BUF1 (N560, N542);
or OR3 (N561, N553, N153, N184);
nand NAND3 (N562, N559, N236, N37);
and AND4 (N563, N558, N302, N455, N34);
and AND4 (N564, N561, N124, N526, N136);
xor XOR2 (N565, N564, N20);
and AND3 (N566, N562, N159, N289);
nor NOR4 (N567, N555, N340, N359, N535);
nor NOR2 (N568, N491, N560);
not NOT1 (N569, N314);
or OR4 (N570, N567, N498, N491, N560);
nor NOR3 (N571, N569, N555, N235);
buf BUF1 (N572, N568);
nor NOR4 (N573, N554, N12, N33, N128);
buf BUF1 (N574, N565);
not NOT1 (N575, N574);
nor NOR3 (N576, N563, N200, N415);
nor NOR2 (N577, N575, N151);
not NOT1 (N578, N577);
nor NOR3 (N579, N572, N348, N291);
and AND2 (N580, N566, N459);
and AND4 (N581, N578, N160, N201, N312);
buf BUF1 (N582, N580);
or OR4 (N583, N538, N99, N207, N377);
buf BUF1 (N584, N571);
nor NOR4 (N585, N570, N89, N350, N133);
xor XOR2 (N586, N579, N414);
nand NAND4 (N587, N573, N221, N183, N308);
or OR4 (N588, N556, N78, N96, N252);
buf BUF1 (N589, N584);
not NOT1 (N590, N552);
buf BUF1 (N591, N590);
not NOT1 (N592, N585);
buf BUF1 (N593, N586);
xor XOR2 (N594, N588, N315);
not NOT1 (N595, N591);
not NOT1 (N596, N595);
buf BUF1 (N597, N589);
and AND4 (N598, N576, N72, N98, N67);
and AND3 (N599, N594, N82, N143);
buf BUF1 (N600, N581);
not NOT1 (N601, N593);
nand NAND2 (N602, N599, N585);
and AND2 (N603, N601, N455);
nand NAND4 (N604, N583, N578, N374, N32);
xor XOR2 (N605, N592, N260);
nand NAND4 (N606, N605, N53, N463, N56);
buf BUF1 (N607, N598);
nor NOR4 (N608, N607, N342, N601, N551);
buf BUF1 (N609, N597);
xor XOR2 (N610, N603, N180);
xor XOR2 (N611, N582, N475);
nor NOR3 (N612, N587, N220, N274);
not NOT1 (N613, N602);
not NOT1 (N614, N604);
not NOT1 (N615, N612);
nor NOR4 (N616, N609, N290, N46, N25);
xor XOR2 (N617, N613, N207);
and AND3 (N618, N610, N41, N200);
buf BUF1 (N619, N615);
or OR4 (N620, N611, N514, N358, N533);
nor NOR4 (N621, N616, N489, N557, N439);
nand NAND2 (N622, N618, N502);
or OR3 (N623, N614, N445, N406);
nand NAND4 (N624, N623, N140, N289, N237);
and AND3 (N625, N608, N363, N241);
buf BUF1 (N626, N617);
xor XOR2 (N627, N619, N599);
xor XOR2 (N628, N622, N173);
and AND3 (N629, N621, N22, N604);
xor XOR2 (N630, N606, N336);
xor XOR2 (N631, N596, N569);
buf BUF1 (N632, N627);
nand NAND2 (N633, N624, N345);
nor NOR4 (N634, N630, N539, N285, N490);
nand NAND2 (N635, N632, N525);
and AND2 (N636, N600, N468);
nand NAND3 (N637, N625, N435, N31);
buf BUF1 (N638, N626);
or OR4 (N639, N631, N77, N365, N397);
nand NAND3 (N640, N638, N355, N283);
buf BUF1 (N641, N620);
nand NAND2 (N642, N635, N125);
not NOT1 (N643, N637);
not NOT1 (N644, N633);
not NOT1 (N645, N628);
nand NAND3 (N646, N640, N69, N454);
nor NOR3 (N647, N634, N32, N371);
and AND4 (N648, N646, N257, N629, N124);
xor XOR2 (N649, N156, N288);
not NOT1 (N650, N644);
or OR4 (N651, N641, N46, N304, N482);
nand NAND2 (N652, N649, N615);
buf BUF1 (N653, N650);
nand NAND4 (N654, N642, N266, N585, N607);
buf BUF1 (N655, N648);
nor NOR4 (N656, N639, N350, N495, N588);
nor NOR4 (N657, N653, N656, N568, N411);
nand NAND4 (N658, N83, N295, N387, N128);
buf BUF1 (N659, N657);
or OR4 (N660, N645, N534, N157, N366);
buf BUF1 (N661, N636);
or OR2 (N662, N643, N338);
nor NOR3 (N663, N655, N219, N481);
and AND4 (N664, N661, N232, N375, N178);
nor NOR4 (N665, N663, N482, N146, N360);
not NOT1 (N666, N658);
and AND2 (N667, N652, N25);
buf BUF1 (N668, N665);
or OR4 (N669, N651, N198, N258, N33);
xor XOR2 (N670, N667, N101);
not NOT1 (N671, N647);
and AND3 (N672, N668, N475, N410);
and AND2 (N673, N664, N304);
nor NOR4 (N674, N654, N621, N30, N255);
nand NAND4 (N675, N666, N669, N620, N247);
not NOT1 (N676, N230);
or OR3 (N677, N676, N563, N501);
xor XOR2 (N678, N671, N504);
not NOT1 (N679, N660);
or OR3 (N680, N679, N350, N596);
nor NOR3 (N681, N680, N361, N663);
and AND2 (N682, N677, N96);
nand NAND2 (N683, N670, N608);
nand NAND2 (N684, N662, N607);
xor XOR2 (N685, N672, N668);
and AND2 (N686, N674, N82);
buf BUF1 (N687, N681);
buf BUF1 (N688, N684);
xor XOR2 (N689, N678, N347);
buf BUF1 (N690, N673);
buf BUF1 (N691, N659);
nor NOR4 (N692, N687, N283, N600, N97);
nand NAND4 (N693, N691, N380, N38, N277);
buf BUF1 (N694, N686);
buf BUF1 (N695, N675);
not NOT1 (N696, N694);
or OR3 (N697, N690, N33, N679);
or OR4 (N698, N693, N281, N606, N12);
buf BUF1 (N699, N695);
not NOT1 (N700, N689);
not NOT1 (N701, N699);
not NOT1 (N702, N701);
nor NOR3 (N703, N685, N254, N699);
buf BUF1 (N704, N682);
or OR4 (N705, N698, N317, N438, N396);
and AND2 (N706, N702, N624);
or OR2 (N707, N703, N550);
nand NAND2 (N708, N707, N246);
buf BUF1 (N709, N700);
and AND3 (N710, N708, N162, N291);
and AND4 (N711, N705, N214, N512, N211);
xor XOR2 (N712, N696, N27);
nor NOR2 (N713, N711, N621);
nor NOR3 (N714, N704, N304, N669);
or OR2 (N715, N714, N298);
and AND3 (N716, N692, N301, N611);
xor XOR2 (N717, N706, N706);
or OR2 (N718, N713, N665);
nand NAND4 (N719, N717, N180, N207, N700);
and AND3 (N720, N710, N401, N69);
not NOT1 (N721, N688);
nor NOR4 (N722, N720, N581, N29, N32);
and AND4 (N723, N715, N444, N504, N697);
and AND3 (N724, N634, N40, N66);
and AND2 (N725, N683, N338);
and AND3 (N726, N723, N710, N500);
nand NAND2 (N727, N721, N184);
and AND4 (N728, N725, N243, N645, N543);
and AND3 (N729, N728, N43, N476);
nor NOR2 (N730, N719, N663);
buf BUF1 (N731, N727);
not NOT1 (N732, N729);
and AND4 (N733, N724, N338, N269, N633);
xor XOR2 (N734, N726, N199);
nand NAND4 (N735, N732, N676, N44, N710);
nand NAND3 (N736, N730, N517, N442);
xor XOR2 (N737, N718, N633);
not NOT1 (N738, N722);
and AND2 (N739, N737, N227);
not NOT1 (N740, N733);
buf BUF1 (N741, N716);
not NOT1 (N742, N735);
not NOT1 (N743, N738);
and AND2 (N744, N712, N202);
and AND3 (N745, N709, N334, N483);
buf BUF1 (N746, N734);
nor NOR2 (N747, N739, N230);
and AND4 (N748, N731, N220, N366, N331);
not NOT1 (N749, N746);
or OR2 (N750, N749, N249);
buf BUF1 (N751, N741);
or OR4 (N752, N742, N523, N645, N611);
nand NAND2 (N753, N751, N152);
nand NAND2 (N754, N750, N722);
nor NOR2 (N755, N747, N94);
nor NOR3 (N756, N754, N365, N560);
not NOT1 (N757, N756);
and AND3 (N758, N757, N651, N475);
nand NAND3 (N759, N744, N621, N472);
not NOT1 (N760, N743);
or OR3 (N761, N755, N505, N707);
xor XOR2 (N762, N759, N460);
buf BUF1 (N763, N761);
buf BUF1 (N764, N753);
nor NOR2 (N765, N740, N117);
or OR3 (N766, N752, N467, N587);
or OR3 (N767, N763, N534, N317);
buf BUF1 (N768, N762);
and AND3 (N769, N745, N537, N617);
not NOT1 (N770, N748);
nand NAND2 (N771, N758, N23);
xor XOR2 (N772, N768, N198);
xor XOR2 (N773, N760, N432);
nand NAND3 (N774, N773, N492, N88);
xor XOR2 (N775, N770, N476);
and AND2 (N776, N774, N83);
xor XOR2 (N777, N766, N730);
xor XOR2 (N778, N777, N295);
nor NOR2 (N779, N775, N604);
and AND2 (N780, N764, N611);
buf BUF1 (N781, N776);
nand NAND3 (N782, N780, N545, N439);
or OR3 (N783, N782, N103, N533);
xor XOR2 (N784, N769, N557);
or OR3 (N785, N736, N375, N574);
and AND3 (N786, N784, N773, N385);
buf BUF1 (N787, N785);
xor XOR2 (N788, N787, N753);
xor XOR2 (N789, N771, N269);
or OR4 (N790, N788, N367, N23, N266);
buf BUF1 (N791, N789);
nand NAND3 (N792, N786, N158, N484);
nor NOR4 (N793, N791, N658, N443, N460);
nand NAND4 (N794, N767, N462, N189, N250);
buf BUF1 (N795, N790);
or OR2 (N796, N778, N5);
nand NAND3 (N797, N792, N177, N660);
nor NOR2 (N798, N781, N575);
and AND4 (N799, N797, N128, N164, N484);
and AND4 (N800, N779, N590, N626, N498);
not NOT1 (N801, N795);
and AND3 (N802, N783, N77, N139);
and AND2 (N803, N772, N482);
nor NOR3 (N804, N803, N263, N188);
not NOT1 (N805, N793);
and AND2 (N806, N794, N280);
or OR4 (N807, N801, N221, N366, N331);
xor XOR2 (N808, N802, N525);
nor NOR3 (N809, N765, N427, N629);
buf BUF1 (N810, N809);
nand NAND2 (N811, N810, N383);
buf BUF1 (N812, N808);
buf BUF1 (N813, N811);
xor XOR2 (N814, N807, N199);
or OR3 (N815, N798, N704, N526);
nand NAND3 (N816, N800, N415, N42);
and AND2 (N817, N813, N325);
nor NOR3 (N818, N817, N390, N496);
buf BUF1 (N819, N818);
nand NAND3 (N820, N819, N594, N489);
nand NAND3 (N821, N799, N322, N810);
buf BUF1 (N822, N815);
not NOT1 (N823, N805);
nand NAND4 (N824, N796, N387, N634, N439);
and AND2 (N825, N814, N813);
or OR2 (N826, N816, N282);
nor NOR3 (N827, N812, N495, N49);
nand NAND4 (N828, N822, N641, N816, N593);
and AND4 (N829, N824, N370, N797, N628);
nand NAND4 (N830, N828, N112, N497, N399);
buf BUF1 (N831, N830);
not NOT1 (N832, N821);
buf BUF1 (N833, N804);
nand NAND4 (N834, N823, N49, N378, N233);
not NOT1 (N835, N826);
nand NAND4 (N836, N833, N370, N201, N578);
or OR3 (N837, N829, N479, N407);
nor NOR4 (N838, N834, N216, N524, N809);
nor NOR4 (N839, N837, N219, N212, N274);
nor NOR2 (N840, N839, N360);
nor NOR4 (N841, N840, N325, N372, N636);
nor NOR2 (N842, N825, N720);
nor NOR4 (N843, N836, N322, N50, N4);
and AND3 (N844, N841, N251, N626);
and AND4 (N845, N835, N788, N635, N150);
nand NAND4 (N846, N832, N425, N591, N341);
and AND4 (N847, N843, N65, N313, N518);
not NOT1 (N848, N842);
not NOT1 (N849, N838);
and AND2 (N850, N806, N752);
and AND4 (N851, N847, N5, N210, N171);
xor XOR2 (N852, N846, N160);
and AND4 (N853, N845, N65, N43, N228);
nand NAND2 (N854, N850, N730);
or OR3 (N855, N852, N141, N105);
nand NAND2 (N856, N851, N704);
or OR3 (N857, N855, N756, N716);
and AND2 (N858, N854, N327);
or OR2 (N859, N856, N794);
not NOT1 (N860, N853);
or OR4 (N861, N848, N426, N46, N122);
buf BUF1 (N862, N859);
nand NAND4 (N863, N858, N57, N475, N615);
or OR4 (N864, N831, N337, N524, N354);
nor NOR2 (N865, N864, N841);
buf BUF1 (N866, N849);
not NOT1 (N867, N863);
and AND3 (N868, N844, N599, N845);
xor XOR2 (N869, N867, N680);
and AND3 (N870, N865, N201, N319);
buf BUF1 (N871, N866);
or OR3 (N872, N857, N693, N59);
or OR4 (N873, N872, N441, N554, N732);
nor NOR2 (N874, N820, N794);
and AND4 (N875, N868, N706, N69, N845);
not NOT1 (N876, N827);
nand NAND3 (N877, N876, N431, N291);
buf BUF1 (N878, N862);
nor NOR3 (N879, N869, N420, N863);
and AND2 (N880, N879, N1);
not NOT1 (N881, N878);
and AND3 (N882, N871, N97, N768);
buf BUF1 (N883, N877);
and AND4 (N884, N873, N162, N18, N713);
xor XOR2 (N885, N860, N576);
buf BUF1 (N886, N883);
or OR4 (N887, N886, N201, N442, N270);
xor XOR2 (N888, N874, N169);
xor XOR2 (N889, N885, N587);
buf BUF1 (N890, N880);
nand NAND4 (N891, N888, N10, N105, N385);
xor XOR2 (N892, N881, N639);
nand NAND2 (N893, N887, N447);
or OR3 (N894, N882, N612, N543);
not NOT1 (N895, N875);
buf BUF1 (N896, N870);
not NOT1 (N897, N889);
xor XOR2 (N898, N892, N533);
not NOT1 (N899, N898);
and AND3 (N900, N884, N350, N70);
or OR4 (N901, N900, N661, N584, N625);
nand NAND4 (N902, N895, N368, N202, N657);
or OR2 (N903, N899, N511);
nand NAND4 (N904, N903, N585, N16, N308);
nor NOR2 (N905, N896, N802);
not NOT1 (N906, N891);
nand NAND3 (N907, N894, N435, N712);
nand NAND2 (N908, N904, N124);
not NOT1 (N909, N907);
or OR4 (N910, N861, N647, N511, N400);
nor NOR3 (N911, N908, N216, N245);
nor NOR2 (N912, N901, N681);
not NOT1 (N913, N905);
buf BUF1 (N914, N911);
nor NOR4 (N915, N909, N203, N554, N787);
nand NAND2 (N916, N897, N351);
and AND3 (N917, N893, N674, N181);
and AND2 (N918, N902, N895);
not NOT1 (N919, N914);
and AND3 (N920, N912, N451, N541);
endmodule