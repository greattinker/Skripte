// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N819,N814,N820,N803,N810,N786,N821,N812,N815,N822;

and AND2 (N23, N3, N18);
and AND3 (N24, N16, N11, N22);
nor NOR2 (N25, N18, N14);
and AND4 (N26, N18, N3, N22, N16);
or OR3 (N27, N5, N10, N3);
xor XOR2 (N28, N11, N7);
and AND2 (N29, N12, N10);
buf BUF1 (N30, N15);
not NOT1 (N31, N4);
or OR4 (N32, N4, N9, N28, N27);
and AND3 (N33, N7, N12, N14);
nor NOR3 (N34, N30, N28, N10);
buf BUF1 (N35, N4);
nor NOR2 (N36, N23, N7);
nor NOR2 (N37, N25, N26);
or OR3 (N38, N24, N4, N33);
nand NAND4 (N39, N2, N16, N17, N28);
nor NOR4 (N40, N17, N38, N29, N13);
or OR3 (N41, N17, N5, N25);
and AND2 (N42, N29, N6);
and AND2 (N43, N31, N12);
nand NAND4 (N44, N39, N3, N17, N12);
or OR2 (N45, N42, N35);
nand NAND2 (N46, N26, N31);
nor NOR3 (N47, N36, N31, N39);
or OR3 (N48, N40, N15, N31);
not NOT1 (N49, N41);
xor XOR2 (N50, N37, N37);
or OR2 (N51, N46, N16);
or OR3 (N52, N50, N34, N17);
not NOT1 (N53, N13);
not NOT1 (N54, N47);
xor XOR2 (N55, N44, N49);
buf BUF1 (N56, N35);
nor NOR3 (N57, N48, N44, N15);
or OR3 (N58, N56, N49, N32);
xor XOR2 (N59, N49, N50);
or OR3 (N60, N58, N54, N23);
nor NOR2 (N61, N8, N20);
xor XOR2 (N62, N51, N22);
buf BUF1 (N63, N57);
not NOT1 (N64, N60);
or OR4 (N65, N53, N18, N8, N9);
and AND3 (N66, N55, N29, N25);
buf BUF1 (N67, N65);
nand NAND2 (N68, N61, N3);
nor NOR4 (N69, N59, N16, N43, N45);
nand NAND3 (N70, N16, N12, N14);
xor XOR2 (N71, N14, N3);
xor XOR2 (N72, N62, N50);
nand NAND3 (N73, N63, N3, N21);
not NOT1 (N74, N71);
buf BUF1 (N75, N67);
and AND3 (N76, N52, N53, N61);
nand NAND2 (N77, N70, N18);
or OR2 (N78, N64, N14);
nand NAND4 (N79, N76, N46, N7, N44);
not NOT1 (N80, N78);
not NOT1 (N81, N79);
nor NOR2 (N82, N75, N14);
not NOT1 (N83, N81);
buf BUF1 (N84, N73);
nand NAND4 (N85, N72, N10, N36, N15);
or OR3 (N86, N83, N46, N33);
nor NOR3 (N87, N74, N7, N44);
buf BUF1 (N88, N69);
xor XOR2 (N89, N85, N38);
or OR4 (N90, N68, N12, N61, N12);
xor XOR2 (N91, N89, N73);
xor XOR2 (N92, N88, N73);
nand NAND4 (N93, N86, N37, N90, N24);
buf BUF1 (N94, N57);
buf BUF1 (N95, N77);
nor NOR4 (N96, N66, N27, N28, N62);
or OR3 (N97, N91, N32, N91);
not NOT1 (N98, N94);
buf BUF1 (N99, N95);
buf BUF1 (N100, N92);
nor NOR2 (N101, N98, N1);
and AND3 (N102, N82, N54, N100);
buf BUF1 (N103, N14);
and AND3 (N104, N101, N12, N28);
and AND2 (N105, N84, N77);
xor XOR2 (N106, N99, N76);
and AND3 (N107, N103, N44, N50);
or OR3 (N108, N105, N51, N57);
buf BUF1 (N109, N102);
nor NOR2 (N110, N93, N62);
nand NAND4 (N111, N96, N109, N58, N41);
xor XOR2 (N112, N89, N60);
nor NOR3 (N113, N108, N81, N51);
and AND2 (N114, N104, N85);
xor XOR2 (N115, N111, N59);
nand NAND3 (N116, N114, N114, N97);
or OR4 (N117, N80, N48, N61, N34);
nand NAND4 (N118, N34, N81, N50, N98);
xor XOR2 (N119, N118, N77);
buf BUF1 (N120, N113);
buf BUF1 (N121, N116);
not NOT1 (N122, N121);
nor NOR2 (N123, N120, N27);
nor NOR4 (N124, N117, N53, N85, N76);
xor XOR2 (N125, N124, N54);
or OR4 (N126, N87, N32, N45, N55);
nor NOR3 (N127, N122, N124, N56);
nor NOR3 (N128, N127, N47, N122);
buf BUF1 (N129, N128);
or OR3 (N130, N129, N17, N99);
nand NAND3 (N131, N130, N83, N68);
nor NOR2 (N132, N131, N50);
nor NOR2 (N133, N107, N48);
and AND2 (N134, N112, N124);
buf BUF1 (N135, N106);
or OR2 (N136, N125, N29);
not NOT1 (N137, N136);
xor XOR2 (N138, N134, N72);
nor NOR3 (N139, N138, N55, N1);
or OR2 (N140, N119, N10);
xor XOR2 (N141, N126, N46);
buf BUF1 (N142, N140);
nand NAND3 (N143, N137, N95, N34);
or OR3 (N144, N139, N8, N143);
buf BUF1 (N145, N74);
and AND3 (N146, N141, N138, N86);
or OR2 (N147, N110, N123);
not NOT1 (N148, N47);
nand NAND4 (N149, N142, N132, N88, N114);
buf BUF1 (N150, N140);
or OR2 (N151, N115, N100);
nand NAND2 (N152, N149, N140);
nor NOR3 (N153, N145, N131, N14);
and AND2 (N154, N152, N89);
nor NOR4 (N155, N148, N53, N110, N141);
or OR2 (N156, N153, N64);
not NOT1 (N157, N150);
not NOT1 (N158, N154);
nand NAND4 (N159, N135, N62, N68, N84);
not NOT1 (N160, N155);
or OR2 (N161, N144, N8);
or OR3 (N162, N156, N97, N92);
buf BUF1 (N163, N147);
and AND4 (N164, N158, N121, N68, N140);
nand NAND2 (N165, N163, N144);
not NOT1 (N166, N162);
and AND3 (N167, N165, N108, N2);
buf BUF1 (N168, N146);
and AND4 (N169, N161, N110, N66, N155);
and AND4 (N170, N160, N44, N113, N95);
or OR2 (N171, N169, N151);
nor NOR4 (N172, N125, N42, N65, N49);
nor NOR4 (N173, N171, N10, N168, N144);
or OR2 (N174, N54, N87);
not NOT1 (N175, N157);
nor NOR4 (N176, N170, N33, N83, N160);
nand NAND4 (N177, N175, N136, N13, N98);
buf BUF1 (N178, N167);
buf BUF1 (N179, N166);
xor XOR2 (N180, N177, N52);
xor XOR2 (N181, N164, N96);
nand NAND3 (N182, N176, N171, N123);
not NOT1 (N183, N133);
nand NAND2 (N184, N172, N170);
or OR4 (N185, N159, N104, N18, N81);
buf BUF1 (N186, N179);
xor XOR2 (N187, N184, N105);
and AND4 (N188, N183, N128, N15, N2);
buf BUF1 (N189, N178);
and AND2 (N190, N189, N74);
nor NOR2 (N191, N181, N185);
nor NOR4 (N192, N47, N162, N117, N111);
buf BUF1 (N193, N180);
or OR3 (N194, N192, N126, N70);
or OR4 (N195, N182, N140, N143, N185);
nor NOR4 (N196, N194, N169, N161, N160);
not NOT1 (N197, N187);
nand NAND4 (N198, N197, N178, N22, N108);
nor NOR3 (N199, N198, N158, N76);
nand NAND3 (N200, N186, N50, N199);
nor NOR3 (N201, N107, N124, N193);
xor XOR2 (N202, N120, N23);
not NOT1 (N203, N196);
buf BUF1 (N204, N203);
buf BUF1 (N205, N200);
and AND4 (N206, N201, N91, N143, N128);
nor NOR2 (N207, N174, N103);
buf BUF1 (N208, N205);
and AND4 (N209, N206, N157, N14, N66);
xor XOR2 (N210, N208, N16);
nor NOR2 (N211, N191, N194);
nand NAND4 (N212, N202, N194, N117, N88);
nor NOR4 (N213, N190, N1, N195, N163);
or OR2 (N214, N148, N51);
and AND4 (N215, N214, N28, N40, N129);
nor NOR4 (N216, N207, N37, N42, N103);
nor NOR4 (N217, N173, N82, N45, N1);
and AND3 (N218, N217, N2, N29);
xor XOR2 (N219, N215, N127);
buf BUF1 (N220, N212);
and AND3 (N221, N188, N203, N149);
nand NAND4 (N222, N210, N4, N213, N27);
nor NOR2 (N223, N60, N163);
or OR4 (N224, N218, N40, N93, N44);
nand NAND4 (N225, N220, N162, N18, N129);
nand NAND2 (N226, N219, N21);
not NOT1 (N227, N223);
buf BUF1 (N228, N225);
xor XOR2 (N229, N221, N219);
nor NOR4 (N230, N229, N191, N68, N103);
not NOT1 (N231, N226);
and AND4 (N232, N211, N144, N140, N103);
not NOT1 (N233, N231);
or OR2 (N234, N224, N151);
xor XOR2 (N235, N204, N173);
nand NAND4 (N236, N222, N189, N89, N200);
or OR2 (N237, N234, N79);
nand NAND4 (N238, N235, N41, N177, N129);
buf BUF1 (N239, N227);
nand NAND2 (N240, N239, N226);
xor XOR2 (N241, N236, N34);
and AND2 (N242, N228, N183);
and AND4 (N243, N238, N68, N157, N17);
not NOT1 (N244, N209);
nand NAND4 (N245, N230, N189, N192, N141);
or OR4 (N246, N232, N39, N217, N216);
xor XOR2 (N247, N172, N176);
nor NOR4 (N248, N240, N195, N143, N219);
buf BUF1 (N249, N246);
xor XOR2 (N250, N243, N6);
buf BUF1 (N251, N245);
nor NOR3 (N252, N233, N172, N53);
xor XOR2 (N253, N242, N20);
not NOT1 (N254, N250);
and AND4 (N255, N247, N27, N239, N47);
xor XOR2 (N256, N244, N91);
or OR4 (N257, N252, N97, N197, N212);
and AND3 (N258, N256, N84, N104);
xor XOR2 (N259, N258, N85);
or OR3 (N260, N241, N110, N3);
not NOT1 (N261, N257);
nand NAND3 (N262, N259, N237, N76);
nand NAND3 (N263, N177, N106, N238);
nand NAND4 (N264, N248, N33, N136, N224);
nor NOR2 (N265, N255, N34);
and AND3 (N266, N251, N150, N193);
nor NOR3 (N267, N266, N258, N96);
buf BUF1 (N268, N263);
xor XOR2 (N269, N253, N248);
nor NOR3 (N270, N267, N193, N95);
buf BUF1 (N271, N264);
xor XOR2 (N272, N268, N153);
buf BUF1 (N273, N249);
not NOT1 (N274, N265);
not NOT1 (N275, N262);
buf BUF1 (N276, N270);
nand NAND2 (N277, N260, N184);
nand NAND2 (N278, N269, N23);
nand NAND2 (N279, N272, N185);
nand NAND3 (N280, N279, N150, N273);
buf BUF1 (N281, N124);
nor NOR2 (N282, N271, N249);
nor NOR3 (N283, N278, N275, N144);
not NOT1 (N284, N110);
and AND3 (N285, N254, N156, N271);
xor XOR2 (N286, N282, N257);
nand NAND2 (N287, N281, N188);
not NOT1 (N288, N285);
nor NOR3 (N289, N286, N78, N278);
nand NAND4 (N290, N288, N177, N26, N278);
and AND4 (N291, N284, N239, N178, N1);
or OR3 (N292, N283, N196, N98);
and AND3 (N293, N280, N283, N2);
or OR4 (N294, N276, N263, N282, N84);
or OR2 (N295, N292, N285);
buf BUF1 (N296, N287);
xor XOR2 (N297, N293, N79);
and AND3 (N298, N291, N227, N173);
nand NAND3 (N299, N277, N175, N142);
buf BUF1 (N300, N289);
nand NAND2 (N301, N294, N107);
or OR2 (N302, N290, N301);
buf BUF1 (N303, N144);
buf BUF1 (N304, N298);
buf BUF1 (N305, N297);
not NOT1 (N306, N302);
buf BUF1 (N307, N299);
nand NAND3 (N308, N305, N32, N169);
xor XOR2 (N309, N295, N287);
or OR4 (N310, N303, N128, N72, N165);
buf BUF1 (N311, N309);
nand NAND3 (N312, N300, N187, N172);
not NOT1 (N313, N310);
or OR2 (N314, N311, N7);
nor NOR3 (N315, N313, N100, N28);
and AND2 (N316, N274, N196);
or OR3 (N317, N315, N312, N192);
buf BUF1 (N318, N28);
xor XOR2 (N319, N304, N160);
or OR2 (N320, N314, N219);
nor NOR3 (N321, N319, N87, N252);
and AND2 (N322, N320, N132);
nor NOR4 (N323, N296, N60, N68, N131);
xor XOR2 (N324, N323, N83);
or OR3 (N325, N308, N282, N86);
nor NOR4 (N326, N306, N289, N197, N319);
not NOT1 (N327, N326);
nor NOR3 (N328, N317, N311, N152);
and AND2 (N329, N322, N68);
xor XOR2 (N330, N307, N319);
xor XOR2 (N331, N330, N132);
nor NOR2 (N332, N325, N296);
not NOT1 (N333, N332);
and AND2 (N334, N261, N287);
xor XOR2 (N335, N333, N198);
buf BUF1 (N336, N334);
not NOT1 (N337, N335);
nor NOR2 (N338, N321, N143);
nor NOR4 (N339, N328, N193, N218, N233);
nand NAND2 (N340, N339, N213);
or OR2 (N341, N340, N330);
buf BUF1 (N342, N331);
and AND3 (N343, N336, N87, N318);
nor NOR4 (N344, N118, N109, N166, N258);
or OR4 (N345, N341, N52, N334, N322);
buf BUF1 (N346, N329);
buf BUF1 (N347, N343);
nand NAND4 (N348, N327, N287, N319, N279);
buf BUF1 (N349, N337);
buf BUF1 (N350, N316);
not NOT1 (N351, N349);
and AND4 (N352, N348, N210, N270, N158);
and AND4 (N353, N338, N205, N52, N257);
not NOT1 (N354, N345);
not NOT1 (N355, N342);
xor XOR2 (N356, N351, N322);
nand NAND2 (N357, N352, N195);
not NOT1 (N358, N354);
not NOT1 (N359, N347);
or OR4 (N360, N350, N110, N230, N112);
nand NAND4 (N361, N356, N282, N75, N302);
not NOT1 (N362, N324);
not NOT1 (N363, N360);
or OR3 (N364, N362, N52, N335);
or OR3 (N365, N363, N55, N121);
nand NAND2 (N366, N359, N288);
and AND3 (N367, N346, N289, N111);
not NOT1 (N368, N364);
nor NOR2 (N369, N357, N149);
xor XOR2 (N370, N365, N15);
xor XOR2 (N371, N370, N81);
not NOT1 (N372, N366);
not NOT1 (N373, N367);
xor XOR2 (N374, N344, N30);
not NOT1 (N375, N358);
or OR4 (N376, N368, N292, N101, N269);
xor XOR2 (N377, N361, N270);
xor XOR2 (N378, N374, N173);
buf BUF1 (N379, N375);
buf BUF1 (N380, N373);
not NOT1 (N381, N377);
and AND2 (N382, N381, N150);
xor XOR2 (N383, N371, N234);
and AND3 (N384, N376, N132, N197);
nand NAND3 (N385, N369, N382, N67);
nand NAND2 (N386, N123, N61);
buf BUF1 (N387, N355);
nor NOR3 (N388, N372, N201, N323);
and AND4 (N389, N384, N386, N11, N189);
nand NAND2 (N390, N43, N97);
and AND2 (N391, N378, N299);
nand NAND4 (N392, N390, N375, N64, N299);
not NOT1 (N393, N392);
not NOT1 (N394, N388);
xor XOR2 (N395, N385, N326);
xor XOR2 (N396, N389, N34);
xor XOR2 (N397, N383, N180);
not NOT1 (N398, N397);
nor NOR4 (N399, N396, N192, N313, N100);
xor XOR2 (N400, N398, N200);
or OR3 (N401, N399, N309, N355);
and AND2 (N402, N380, N49);
nor NOR3 (N403, N400, N104, N47);
nor NOR2 (N404, N353, N276);
nor NOR3 (N405, N393, N373, N87);
nand NAND3 (N406, N395, N164, N107);
or OR3 (N407, N404, N63, N52);
xor XOR2 (N408, N379, N205);
nand NAND4 (N409, N408, N325, N52, N90);
not NOT1 (N410, N402);
and AND3 (N411, N394, N66, N357);
buf BUF1 (N412, N401);
xor XOR2 (N413, N391, N164);
xor XOR2 (N414, N413, N119);
xor XOR2 (N415, N414, N363);
and AND3 (N416, N387, N166, N286);
or OR3 (N417, N410, N296, N20);
and AND3 (N418, N411, N104, N56);
nand NAND2 (N419, N416, N374);
not NOT1 (N420, N405);
nor NOR3 (N421, N418, N407, N363);
not NOT1 (N422, N179);
or OR2 (N423, N421, N24);
not NOT1 (N424, N409);
nand NAND2 (N425, N422, N387);
nor NOR2 (N426, N424, N289);
and AND2 (N427, N415, N133);
or OR3 (N428, N406, N310, N234);
or OR2 (N429, N420, N65);
not NOT1 (N430, N427);
nand NAND3 (N431, N429, N236, N387);
not NOT1 (N432, N417);
or OR4 (N433, N426, N277, N161, N101);
nand NAND4 (N434, N425, N294, N276, N89);
not NOT1 (N435, N431);
xor XOR2 (N436, N423, N387);
or OR4 (N437, N432, N43, N141, N170);
nor NOR3 (N438, N403, N85, N67);
and AND2 (N439, N437, N18);
not NOT1 (N440, N439);
xor XOR2 (N441, N436, N24);
or OR2 (N442, N441, N82);
and AND4 (N443, N442, N147, N376, N267);
not NOT1 (N444, N430);
not NOT1 (N445, N443);
not NOT1 (N446, N435);
and AND3 (N447, N428, N43, N351);
and AND3 (N448, N444, N242, N106);
or OR4 (N449, N434, N270, N105, N145);
not NOT1 (N450, N433);
not NOT1 (N451, N419);
nand NAND2 (N452, N449, N451);
nand NAND2 (N453, N216, N308);
nor NOR3 (N454, N452, N289, N304);
buf BUF1 (N455, N450);
nor NOR4 (N456, N445, N65, N154, N133);
nand NAND2 (N457, N453, N228);
buf BUF1 (N458, N446);
nand NAND3 (N459, N412, N181, N207);
or OR3 (N460, N448, N328, N285);
nand NAND3 (N461, N460, N39, N144);
xor XOR2 (N462, N458, N345);
xor XOR2 (N463, N455, N183);
not NOT1 (N464, N456);
buf BUF1 (N465, N463);
nand NAND2 (N466, N459, N139);
not NOT1 (N467, N461);
or OR3 (N468, N457, N416, N9);
or OR4 (N469, N464, N264, N131, N327);
nand NAND3 (N470, N438, N257, N456);
or OR4 (N471, N447, N185, N319, N217);
nand NAND4 (N472, N462, N357, N245, N85);
xor XOR2 (N473, N466, N44);
or OR4 (N474, N465, N352, N116, N146);
or OR4 (N475, N471, N71, N172, N351);
nand NAND4 (N476, N474, N387, N237, N255);
and AND3 (N477, N472, N343, N137);
not NOT1 (N478, N477);
xor XOR2 (N479, N467, N310);
buf BUF1 (N480, N479);
and AND3 (N481, N478, N139, N323);
buf BUF1 (N482, N480);
nor NOR2 (N483, N454, N191);
not NOT1 (N484, N476);
and AND2 (N485, N481, N241);
not NOT1 (N486, N469);
and AND2 (N487, N484, N212);
buf BUF1 (N488, N486);
nor NOR4 (N489, N468, N176, N318, N93);
not NOT1 (N490, N440);
or OR4 (N491, N475, N227, N354, N69);
nor NOR4 (N492, N489, N124, N414, N273);
buf BUF1 (N493, N470);
buf BUF1 (N494, N473);
nand NAND2 (N495, N492, N221);
and AND2 (N496, N482, N175);
and AND3 (N497, N494, N114, N169);
or OR3 (N498, N488, N95, N262);
nand NAND3 (N499, N497, N179, N171);
not NOT1 (N500, N487);
xor XOR2 (N501, N495, N494);
xor XOR2 (N502, N493, N81);
nand NAND3 (N503, N496, N215, N101);
not NOT1 (N504, N490);
nand NAND4 (N505, N500, N376, N246, N326);
xor XOR2 (N506, N503, N95);
and AND4 (N507, N506, N443, N317, N153);
buf BUF1 (N508, N501);
or OR2 (N509, N508, N505);
nand NAND2 (N510, N136, N401);
buf BUF1 (N511, N483);
nand NAND2 (N512, N504, N189);
and AND3 (N513, N510, N127, N266);
not NOT1 (N514, N507);
and AND4 (N515, N498, N312, N396, N467);
buf BUF1 (N516, N515);
and AND4 (N517, N502, N350, N51, N477);
nor NOR3 (N518, N512, N424, N338);
buf BUF1 (N519, N516);
or OR2 (N520, N491, N398);
buf BUF1 (N521, N509);
xor XOR2 (N522, N514, N16);
or OR3 (N523, N521, N193, N45);
nor NOR3 (N524, N511, N65, N55);
nand NAND3 (N525, N513, N296, N516);
not NOT1 (N526, N499);
not NOT1 (N527, N522);
or OR3 (N528, N527, N194, N1);
xor XOR2 (N529, N520, N145);
xor XOR2 (N530, N526, N340);
xor XOR2 (N531, N529, N44);
or OR4 (N532, N530, N351, N132, N111);
nand NAND3 (N533, N525, N142, N379);
nor NOR3 (N534, N485, N35, N396);
buf BUF1 (N535, N517);
or OR4 (N536, N524, N171, N202, N522);
nand NAND3 (N537, N531, N131, N399);
buf BUF1 (N538, N518);
not NOT1 (N539, N535);
or OR4 (N540, N538, N405, N164, N240);
nand NAND4 (N541, N536, N405, N352, N484);
nand NAND3 (N542, N532, N501, N369);
nand NAND4 (N543, N542, N169, N85, N159);
xor XOR2 (N544, N519, N306);
buf BUF1 (N545, N543);
or OR4 (N546, N534, N476, N537, N209);
xor XOR2 (N547, N509, N74);
nand NAND3 (N548, N539, N285, N281);
nor NOR4 (N549, N545, N219, N508, N4);
not NOT1 (N550, N546);
buf BUF1 (N551, N541);
not NOT1 (N552, N549);
and AND2 (N553, N551, N34);
xor XOR2 (N554, N550, N344);
nor NOR2 (N555, N548, N107);
nand NAND2 (N556, N552, N419);
or OR2 (N557, N533, N378);
not NOT1 (N558, N555);
nand NAND4 (N559, N557, N221, N55, N373);
nand NAND2 (N560, N540, N249);
not NOT1 (N561, N554);
not NOT1 (N562, N553);
xor XOR2 (N563, N562, N519);
xor XOR2 (N564, N561, N450);
and AND4 (N565, N564, N11, N125, N146);
nand NAND2 (N566, N544, N441);
and AND4 (N567, N547, N222, N549, N479);
nand NAND3 (N568, N523, N266, N434);
nand NAND3 (N569, N560, N241, N67);
buf BUF1 (N570, N565);
nand NAND4 (N571, N559, N440, N502, N255);
nand NAND3 (N572, N570, N1, N430);
buf BUF1 (N573, N568);
xor XOR2 (N574, N556, N126);
not NOT1 (N575, N573);
and AND3 (N576, N574, N558, N345);
and AND2 (N577, N559, N261);
and AND4 (N578, N566, N29, N110, N310);
or OR3 (N579, N577, N359, N465);
xor XOR2 (N580, N576, N149);
nand NAND3 (N581, N528, N367, N112);
or OR4 (N582, N581, N9, N162, N541);
or OR4 (N583, N580, N329, N250, N450);
or OR3 (N584, N571, N73, N457);
not NOT1 (N585, N567);
xor XOR2 (N586, N578, N203);
buf BUF1 (N587, N582);
not NOT1 (N588, N586);
nor NOR3 (N589, N563, N428, N46);
xor XOR2 (N590, N579, N353);
buf BUF1 (N591, N572);
nor NOR4 (N592, N583, N261, N81, N302);
xor XOR2 (N593, N585, N426);
buf BUF1 (N594, N569);
buf BUF1 (N595, N592);
nor NOR4 (N596, N588, N370, N494, N111);
buf BUF1 (N597, N591);
and AND4 (N598, N595, N46, N53, N278);
and AND3 (N599, N594, N442, N32);
buf BUF1 (N600, N593);
not NOT1 (N601, N589);
or OR3 (N602, N587, N466, N221);
not NOT1 (N603, N596);
not NOT1 (N604, N600);
buf BUF1 (N605, N602);
not NOT1 (N606, N584);
or OR3 (N607, N603, N568, N187);
or OR4 (N608, N590, N228, N8, N588);
nand NAND3 (N609, N575, N102, N340);
not NOT1 (N610, N598);
nor NOR3 (N611, N605, N150, N132);
nand NAND4 (N612, N611, N99, N321, N127);
or OR3 (N613, N610, N37, N383);
or OR3 (N614, N607, N297, N540);
nor NOR3 (N615, N601, N12, N306);
not NOT1 (N616, N604);
nand NAND4 (N617, N616, N54, N606, N287);
not NOT1 (N618, N482);
xor XOR2 (N619, N614, N287);
buf BUF1 (N620, N618);
xor XOR2 (N621, N599, N264);
or OR4 (N622, N612, N333, N575, N309);
nand NAND2 (N623, N597, N185);
xor XOR2 (N624, N622, N107);
nor NOR3 (N625, N619, N356, N193);
or OR4 (N626, N615, N195, N345, N599);
or OR2 (N627, N623, N282);
not NOT1 (N628, N621);
nor NOR3 (N629, N620, N590, N512);
or OR2 (N630, N627, N111);
nand NAND4 (N631, N624, N109, N356, N275);
nand NAND4 (N632, N631, N215, N378, N367);
not NOT1 (N633, N630);
buf BUF1 (N634, N632);
and AND2 (N635, N617, N42);
nand NAND4 (N636, N613, N486, N297, N541);
not NOT1 (N637, N608);
and AND2 (N638, N625, N494);
or OR3 (N639, N626, N536, N317);
not NOT1 (N640, N637);
xor XOR2 (N641, N609, N116);
and AND2 (N642, N636, N582);
xor XOR2 (N643, N639, N348);
not NOT1 (N644, N640);
nand NAND3 (N645, N643, N32, N531);
buf BUF1 (N646, N635);
nand NAND3 (N647, N641, N94, N44);
and AND4 (N648, N633, N51, N285, N400);
nor NOR4 (N649, N628, N132, N12, N182);
and AND4 (N650, N638, N628, N393, N636);
nand NAND3 (N651, N647, N234, N574);
buf BUF1 (N652, N644);
nor NOR3 (N653, N629, N230, N110);
nor NOR2 (N654, N653, N541);
xor XOR2 (N655, N634, N483);
nor NOR3 (N656, N645, N229, N43);
or OR4 (N657, N652, N590, N452, N230);
or OR4 (N658, N646, N448, N291, N420);
nand NAND2 (N659, N655, N596);
nor NOR4 (N660, N651, N393, N559, N494);
and AND2 (N661, N656, N603);
not NOT1 (N662, N658);
and AND4 (N663, N661, N123, N23, N93);
not NOT1 (N664, N657);
xor XOR2 (N665, N660, N411);
and AND2 (N666, N664, N27);
buf BUF1 (N667, N662);
and AND3 (N668, N659, N102, N118);
buf BUF1 (N669, N667);
xor XOR2 (N670, N665, N466);
xor XOR2 (N671, N669, N603);
xor XOR2 (N672, N666, N12);
or OR3 (N673, N670, N418, N274);
nand NAND2 (N674, N668, N143);
nand NAND3 (N675, N672, N5, N120);
xor XOR2 (N676, N654, N53);
xor XOR2 (N677, N648, N632);
and AND3 (N678, N650, N373, N523);
or OR3 (N679, N678, N655, N293);
xor XOR2 (N680, N677, N573);
not NOT1 (N681, N663);
not NOT1 (N682, N642);
or OR4 (N683, N673, N174, N338, N536);
and AND4 (N684, N676, N446, N373, N221);
buf BUF1 (N685, N680);
or OR2 (N686, N674, N494);
not NOT1 (N687, N675);
nand NAND3 (N688, N671, N177, N300);
nor NOR4 (N689, N688, N611, N635, N362);
buf BUF1 (N690, N685);
not NOT1 (N691, N686);
not NOT1 (N692, N684);
nor NOR3 (N693, N689, N62, N361);
xor XOR2 (N694, N679, N3);
not NOT1 (N695, N694);
or OR4 (N696, N649, N482, N407, N601);
nand NAND3 (N697, N692, N307, N431);
and AND3 (N698, N695, N248, N637);
not NOT1 (N699, N687);
and AND3 (N700, N682, N123, N94);
not NOT1 (N701, N690);
buf BUF1 (N702, N698);
and AND3 (N703, N699, N49, N352);
buf BUF1 (N704, N693);
nor NOR4 (N705, N696, N684, N289, N679);
nor NOR3 (N706, N704, N135, N401);
buf BUF1 (N707, N691);
nor NOR4 (N708, N683, N252, N82, N239);
buf BUF1 (N709, N707);
buf BUF1 (N710, N705);
nand NAND2 (N711, N697, N187);
not NOT1 (N712, N710);
xor XOR2 (N713, N708, N218);
nor NOR3 (N714, N703, N377, N583);
nand NAND3 (N715, N701, N705, N340);
not NOT1 (N716, N715);
not NOT1 (N717, N714);
xor XOR2 (N718, N681, N365);
nand NAND2 (N719, N718, N299);
xor XOR2 (N720, N719, N540);
buf BUF1 (N721, N720);
or OR4 (N722, N711, N676, N424, N515);
not NOT1 (N723, N721);
or OR4 (N724, N723, N630, N421, N679);
and AND3 (N725, N709, N239, N696);
nand NAND3 (N726, N700, N464, N340);
and AND4 (N727, N713, N189, N466, N467);
nor NOR3 (N728, N726, N586, N144);
and AND2 (N729, N702, N345);
or OR2 (N730, N724, N217);
and AND2 (N731, N706, N301);
or OR2 (N732, N727, N341);
not NOT1 (N733, N725);
and AND3 (N734, N712, N561, N169);
nor NOR3 (N735, N716, N725, N3);
buf BUF1 (N736, N730);
nand NAND3 (N737, N722, N173, N637);
or OR2 (N738, N735, N310);
nor NOR2 (N739, N729, N422);
or OR4 (N740, N734, N553, N271, N637);
not NOT1 (N741, N739);
buf BUF1 (N742, N740);
xor XOR2 (N743, N742, N184);
buf BUF1 (N744, N728);
nor NOR2 (N745, N732, N539);
nand NAND4 (N746, N736, N483, N630, N86);
and AND2 (N747, N733, N9);
xor XOR2 (N748, N744, N540);
or OR3 (N749, N746, N313, N368);
buf BUF1 (N750, N749);
buf BUF1 (N751, N717);
not NOT1 (N752, N751);
buf BUF1 (N753, N737);
or OR3 (N754, N741, N144, N693);
and AND4 (N755, N738, N113, N618, N537);
nor NOR2 (N756, N750, N96);
buf BUF1 (N757, N756);
nor NOR2 (N758, N753, N194);
not NOT1 (N759, N752);
nor NOR3 (N760, N757, N700, N385);
buf BUF1 (N761, N754);
nand NAND4 (N762, N743, N752, N388, N720);
nand NAND2 (N763, N758, N526);
not NOT1 (N764, N755);
buf BUF1 (N765, N762);
nand NAND2 (N766, N745, N196);
nor NOR3 (N767, N747, N434, N360);
nor NOR4 (N768, N731, N309, N252, N592);
buf BUF1 (N769, N768);
buf BUF1 (N770, N767);
buf BUF1 (N771, N770);
and AND2 (N772, N771, N204);
nor NOR2 (N773, N759, N27);
buf BUF1 (N774, N773);
nor NOR2 (N775, N764, N101);
xor XOR2 (N776, N766, N611);
nand NAND4 (N777, N776, N572, N455, N270);
and AND2 (N778, N775, N714);
nand NAND2 (N779, N778, N373);
nor NOR2 (N780, N779, N706);
nor NOR3 (N781, N763, N188, N707);
nor NOR3 (N782, N777, N696, N200);
nand NAND3 (N783, N780, N376, N252);
xor XOR2 (N784, N748, N239);
xor XOR2 (N785, N765, N394);
nand NAND3 (N786, N760, N162, N56);
or OR4 (N787, N782, N375, N100, N627);
buf BUF1 (N788, N769);
buf BUF1 (N789, N787);
not NOT1 (N790, N785);
nand NAND2 (N791, N790, N134);
not NOT1 (N792, N781);
not NOT1 (N793, N791);
xor XOR2 (N794, N792, N669);
nand NAND3 (N795, N789, N45, N726);
xor XOR2 (N796, N788, N626);
nor NOR2 (N797, N783, N791);
xor XOR2 (N798, N793, N788);
and AND3 (N799, N797, N340, N57);
nand NAND4 (N800, N761, N344, N206, N733);
nor NOR2 (N801, N772, N797);
buf BUF1 (N802, N794);
not NOT1 (N803, N784);
xor XOR2 (N804, N798, N336);
xor XOR2 (N805, N804, N335);
not NOT1 (N806, N805);
nand NAND3 (N807, N802, N97, N132);
buf BUF1 (N808, N799);
xor XOR2 (N809, N807, N796);
nor NOR3 (N810, N545, N236, N571);
xor XOR2 (N811, N774, N673);
not NOT1 (N812, N811);
or OR4 (N813, N795, N713, N214, N626);
buf BUF1 (N814, N800);
buf BUF1 (N815, N809);
nand NAND4 (N816, N813, N10, N794, N595);
nand NAND3 (N817, N806, N40, N55);
or OR4 (N818, N816, N402, N69, N785);
and AND4 (N819, N817, N343, N641, N55);
xor XOR2 (N820, N801, N129);
nand NAND2 (N821, N808, N186);
nor NOR2 (N822, N818, N757);
endmodule