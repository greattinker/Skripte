// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N399,N393,N403,N407,N411,N413,N405,N409,N410,N414;

not NOT1 (N15, N12);
nand NAND4 (N16, N3, N10, N4, N14);
buf BUF1 (N17, N11);
or OR2 (N18, N17, N3);
nand NAND2 (N19, N17, N4);
buf BUF1 (N20, N8);
and AND4 (N21, N7, N6, N11, N2);
xor XOR2 (N22, N19, N11);
nor NOR4 (N23, N7, N6, N1, N22);
nand NAND4 (N24, N18, N2, N1, N18);
buf BUF1 (N25, N20);
nor NOR2 (N26, N18, N21);
and AND4 (N27, N21, N15, N25, N26);
buf BUF1 (N28, N15);
xor XOR2 (N29, N28, N23);
or OR3 (N30, N29, N13, N9);
nand NAND4 (N31, N8, N12, N14, N23);
and AND2 (N32, N2, N31);
or OR2 (N33, N23, N29);
xor XOR2 (N34, N32, N14);
or OR4 (N35, N11, N20, N29, N19);
and AND4 (N36, N30, N35, N9, N1);
xor XOR2 (N37, N27, N14);
nor NOR4 (N38, N23, N9, N4, N5);
and AND3 (N39, N37, N22, N4);
xor XOR2 (N40, N32, N28);
not NOT1 (N41, N4);
nor NOR3 (N42, N8, N22, N16);
nor NOR4 (N43, N30, N30, N34, N1);
xor XOR2 (N44, N11, N6);
xor XOR2 (N45, N41, N15);
nor NOR4 (N46, N24, N13, N6, N41);
and AND3 (N47, N36, N6, N46);
nor NOR4 (N48, N7, N2, N21, N8);
xor XOR2 (N49, N33, N16);
not NOT1 (N50, N42);
nor NOR4 (N51, N43, N11, N19, N13);
nand NAND3 (N52, N39, N2, N23);
xor XOR2 (N53, N49, N34);
xor XOR2 (N54, N51, N43);
nand NAND3 (N55, N44, N43, N34);
or OR3 (N56, N48, N54, N28);
nor NOR2 (N57, N33, N56);
xor XOR2 (N58, N55, N44);
buf BUF1 (N59, N57);
not NOT1 (N60, N58);
nand NAND4 (N61, N24, N48, N35, N12);
xor XOR2 (N62, N60, N19);
nor NOR2 (N63, N53, N47);
xor XOR2 (N64, N58, N44);
xor XOR2 (N65, N62, N21);
buf BUF1 (N66, N52);
nand NAND4 (N67, N40, N1, N22, N54);
nand NAND4 (N68, N38, N8, N22, N12);
nand NAND2 (N69, N59, N33);
nor NOR3 (N70, N50, N65, N45);
nand NAND3 (N71, N13, N63, N56);
or OR2 (N72, N45, N25);
buf BUF1 (N73, N45);
or OR4 (N74, N67, N5, N70, N7);
not NOT1 (N75, N29);
or OR2 (N76, N68, N19);
nor NOR2 (N77, N73, N7);
nor NOR4 (N78, N75, N34, N52, N57);
nor NOR3 (N79, N64, N49, N10);
or OR2 (N80, N79, N15);
xor XOR2 (N81, N80, N8);
not NOT1 (N82, N78);
and AND4 (N83, N72, N69, N76, N75);
or OR2 (N84, N73, N13);
nand NAND4 (N85, N2, N14, N24, N65);
buf BUF1 (N86, N71);
nor NOR3 (N87, N83, N38, N36);
buf BUF1 (N88, N66);
and AND4 (N89, N86, N29, N15, N80);
nor NOR3 (N90, N77, N12, N41);
nand NAND4 (N91, N74, N12, N22, N66);
nor NOR4 (N92, N90, N80, N79, N27);
not NOT1 (N93, N81);
xor XOR2 (N94, N92, N63);
nor NOR3 (N95, N61, N93, N82);
nand NAND2 (N96, N57, N2);
nand NAND3 (N97, N17, N75, N16);
or OR2 (N98, N97, N64);
not NOT1 (N99, N89);
xor XOR2 (N100, N99, N65);
and AND4 (N101, N96, N82, N49, N7);
nand NAND2 (N102, N100, N60);
or OR3 (N103, N94, N22, N98);
not NOT1 (N104, N25);
or OR2 (N105, N103, N35);
and AND4 (N106, N101, N46, N57, N26);
nor NOR2 (N107, N88, N5);
or OR4 (N108, N95, N3, N24, N105);
not NOT1 (N109, N79);
or OR4 (N110, N84, N77, N32, N106);
nor NOR2 (N111, N82, N44);
and AND2 (N112, N111, N72);
xor XOR2 (N113, N109, N32);
not NOT1 (N114, N113);
buf BUF1 (N115, N85);
and AND3 (N116, N91, N105, N68);
and AND4 (N117, N114, N38, N63, N33);
nand NAND2 (N118, N117, N4);
xor XOR2 (N119, N87, N108);
not NOT1 (N120, N96);
buf BUF1 (N121, N120);
and AND3 (N122, N102, N35, N75);
and AND2 (N123, N107, N103);
buf BUF1 (N124, N119);
nor NOR2 (N125, N118, N118);
xor XOR2 (N126, N115, N101);
nand NAND2 (N127, N125, N48);
or OR4 (N128, N124, N36, N56, N127);
not NOT1 (N129, N67);
xor XOR2 (N130, N112, N3);
and AND2 (N131, N126, N70);
not NOT1 (N132, N110);
xor XOR2 (N133, N104, N58);
nand NAND4 (N134, N133, N33, N10, N14);
nor NOR3 (N135, N123, N80, N113);
not NOT1 (N136, N134);
not NOT1 (N137, N131);
buf BUF1 (N138, N137);
or OR2 (N139, N128, N39);
not NOT1 (N140, N139);
or OR4 (N141, N130, N116, N125, N85);
buf BUF1 (N142, N56);
nand NAND4 (N143, N132, N115, N64, N91);
nor NOR4 (N144, N141, N18, N42, N5);
and AND3 (N145, N140, N18, N143);
and AND2 (N146, N117, N138);
buf BUF1 (N147, N3);
not NOT1 (N148, N135);
xor XOR2 (N149, N147, N108);
not NOT1 (N150, N146);
or OR3 (N151, N144, N89, N92);
nand NAND2 (N152, N142, N29);
or OR4 (N153, N145, N140, N19, N55);
nand NAND2 (N154, N150, N79);
nand NAND2 (N155, N148, N41);
not NOT1 (N156, N121);
xor XOR2 (N157, N155, N138);
buf BUF1 (N158, N129);
xor XOR2 (N159, N122, N68);
nor NOR4 (N160, N136, N121, N23, N42);
nor NOR4 (N161, N160, N132, N88, N130);
buf BUF1 (N162, N151);
buf BUF1 (N163, N158);
not NOT1 (N164, N162);
not NOT1 (N165, N164);
nor NOR4 (N166, N165, N38, N2, N74);
xor XOR2 (N167, N163, N81);
xor XOR2 (N168, N157, N78);
or OR4 (N169, N152, N84, N48, N81);
or OR3 (N170, N149, N42, N21);
xor XOR2 (N171, N170, N117);
buf BUF1 (N172, N166);
nor NOR2 (N173, N169, N14);
nor NOR4 (N174, N156, N159, N26, N15);
nor NOR2 (N175, N19, N84);
nand NAND3 (N176, N175, N37, N141);
not NOT1 (N177, N171);
buf BUF1 (N178, N168);
nand NAND2 (N179, N174, N58);
nor NOR3 (N180, N176, N153, N99);
nor NOR2 (N181, N142, N106);
and AND2 (N182, N178, N100);
buf BUF1 (N183, N173);
nand NAND3 (N184, N181, N7, N56);
buf BUF1 (N185, N180);
or OR4 (N186, N184, N136, N115, N100);
buf BUF1 (N187, N154);
xor XOR2 (N188, N185, N85);
not NOT1 (N189, N167);
xor XOR2 (N190, N172, N44);
buf BUF1 (N191, N186);
nand NAND4 (N192, N183, N136, N110, N82);
or OR4 (N193, N182, N69, N38, N144);
or OR4 (N194, N187, N140, N4, N26);
not NOT1 (N195, N179);
not NOT1 (N196, N161);
nand NAND2 (N197, N193, N186);
not NOT1 (N198, N189);
nor NOR4 (N199, N198, N190, N171, N101);
not NOT1 (N200, N172);
not NOT1 (N201, N196);
and AND2 (N202, N199, N100);
nor NOR3 (N203, N201, N25, N89);
not NOT1 (N204, N200);
not NOT1 (N205, N202);
or OR4 (N206, N205, N120, N139, N144);
or OR3 (N207, N197, N186, N127);
not NOT1 (N208, N188);
nor NOR3 (N209, N194, N162, N204);
xor XOR2 (N210, N65, N104);
nor NOR3 (N211, N206, N195, N64);
buf BUF1 (N212, N40);
and AND2 (N213, N211, N85);
buf BUF1 (N214, N203);
or OR2 (N215, N213, N168);
not NOT1 (N216, N210);
nor NOR3 (N217, N208, N151, N69);
nand NAND4 (N218, N216, N146, N67, N194);
and AND2 (N219, N218, N178);
or OR2 (N220, N177, N149);
or OR2 (N221, N215, N156);
or OR2 (N222, N217, N185);
nand NAND3 (N223, N212, N88, N164);
and AND3 (N224, N219, N153, N65);
buf BUF1 (N225, N224);
nand NAND2 (N226, N221, N186);
not NOT1 (N227, N220);
nand NAND4 (N228, N209, N92, N121, N111);
and AND4 (N229, N214, N129, N167, N35);
xor XOR2 (N230, N226, N183);
buf BUF1 (N231, N225);
or OR3 (N232, N227, N104, N187);
nand NAND4 (N233, N229, N100, N42, N150);
not NOT1 (N234, N223);
or OR2 (N235, N222, N85);
buf BUF1 (N236, N207);
not NOT1 (N237, N231);
buf BUF1 (N238, N233);
and AND3 (N239, N232, N96, N2);
and AND3 (N240, N228, N206, N174);
nor NOR4 (N241, N191, N133, N239, N159);
and AND4 (N242, N28, N121, N99, N128);
not NOT1 (N243, N237);
and AND2 (N244, N240, N128);
or OR3 (N245, N230, N116, N54);
and AND4 (N246, N243, N115, N234, N184);
xor XOR2 (N247, N168, N101);
xor XOR2 (N248, N246, N114);
nand NAND2 (N249, N248, N194);
and AND3 (N250, N242, N107, N66);
or OR2 (N251, N192, N186);
nand NAND2 (N252, N250, N204);
or OR4 (N253, N247, N39, N95, N64);
not NOT1 (N254, N245);
xor XOR2 (N255, N252, N170);
nor NOR3 (N256, N253, N144, N208);
nand NAND3 (N257, N241, N180, N162);
xor XOR2 (N258, N257, N94);
not NOT1 (N259, N255);
nor NOR2 (N260, N254, N66);
or OR4 (N261, N259, N18, N122, N196);
buf BUF1 (N262, N238);
nand NAND4 (N263, N256, N26, N47, N258);
and AND3 (N264, N34, N132, N211);
nor NOR3 (N265, N261, N168, N11);
not NOT1 (N266, N236);
nand NAND3 (N267, N251, N168, N78);
not NOT1 (N268, N266);
or OR4 (N269, N267, N88, N226, N88);
not NOT1 (N270, N269);
nand NAND2 (N271, N244, N57);
xor XOR2 (N272, N235, N66);
not NOT1 (N273, N270);
not NOT1 (N274, N260);
buf BUF1 (N275, N262);
and AND3 (N276, N265, N148, N10);
buf BUF1 (N277, N249);
and AND3 (N278, N271, N48, N125);
xor XOR2 (N279, N264, N272);
and AND4 (N280, N242, N86, N240, N12);
xor XOR2 (N281, N279, N178);
nand NAND4 (N282, N277, N134, N62, N86);
not NOT1 (N283, N268);
nand NAND3 (N284, N282, N275, N121);
or OR4 (N285, N47, N79, N3, N135);
nand NAND4 (N286, N263, N5, N211, N166);
xor XOR2 (N287, N283, N18);
xor XOR2 (N288, N287, N93);
xor XOR2 (N289, N278, N236);
buf BUF1 (N290, N281);
nor NOR3 (N291, N280, N249, N174);
not NOT1 (N292, N286);
buf BUF1 (N293, N285);
and AND3 (N294, N288, N153, N63);
and AND4 (N295, N294, N128, N238, N191);
nor NOR3 (N296, N284, N247, N213);
xor XOR2 (N297, N293, N240);
and AND4 (N298, N292, N125, N12, N281);
not NOT1 (N299, N290);
and AND3 (N300, N299, N250, N152);
and AND4 (N301, N289, N266, N263, N103);
not NOT1 (N302, N300);
nor NOR4 (N303, N273, N134, N243, N139);
or OR2 (N304, N274, N205);
nand NAND2 (N305, N295, N293);
nor NOR2 (N306, N304, N3);
nor NOR3 (N307, N305, N188, N220);
and AND2 (N308, N306, N107);
and AND2 (N309, N298, N183);
nand NAND2 (N310, N303, N200);
xor XOR2 (N311, N310, N148);
buf BUF1 (N312, N297);
or OR4 (N313, N312, N157, N163, N104);
nor NOR4 (N314, N309, N12, N145, N208);
nor NOR2 (N315, N291, N171);
nand NAND4 (N316, N301, N223, N181, N177);
or OR3 (N317, N311, N17, N256);
xor XOR2 (N318, N313, N173);
nor NOR3 (N319, N308, N260, N212);
buf BUF1 (N320, N296);
nand NAND2 (N321, N315, N295);
nor NOR4 (N322, N321, N107, N248, N312);
nor NOR3 (N323, N318, N88, N153);
xor XOR2 (N324, N314, N16);
buf BUF1 (N325, N276);
xor XOR2 (N326, N320, N146);
buf BUF1 (N327, N324);
nand NAND4 (N328, N327, N218, N216, N216);
not NOT1 (N329, N326);
buf BUF1 (N330, N329);
nand NAND3 (N331, N302, N272, N93);
xor XOR2 (N332, N307, N132);
or OR2 (N333, N330, N85);
not NOT1 (N334, N331);
nor NOR4 (N335, N323, N169, N118, N318);
xor XOR2 (N336, N322, N297);
and AND4 (N337, N325, N40, N266, N150);
xor XOR2 (N338, N335, N217);
nand NAND4 (N339, N336, N280, N114, N123);
or OR2 (N340, N328, N173);
nand NAND2 (N341, N340, N135);
not NOT1 (N342, N332);
not NOT1 (N343, N319);
nand NAND3 (N344, N337, N301, N253);
or OR2 (N345, N339, N74);
buf BUF1 (N346, N334);
and AND4 (N347, N344, N329, N323, N189);
nand NAND2 (N348, N342, N210);
or OR2 (N349, N347, N31);
not NOT1 (N350, N316);
xor XOR2 (N351, N317, N328);
buf BUF1 (N352, N351);
nand NAND3 (N353, N341, N137, N108);
and AND3 (N354, N348, N200, N197);
and AND2 (N355, N350, N310);
nor NOR2 (N356, N349, N40);
nor NOR4 (N357, N352, N112, N9, N136);
not NOT1 (N358, N346);
nand NAND4 (N359, N343, N356, N69, N57);
not NOT1 (N360, N213);
not NOT1 (N361, N358);
nor NOR2 (N362, N360, N235);
buf BUF1 (N363, N359);
nor NOR4 (N364, N353, N200, N183, N180);
nor NOR4 (N365, N364, N287, N241, N170);
or OR2 (N366, N365, N200);
or OR4 (N367, N366, N361, N136, N95);
and AND2 (N368, N257, N245);
or OR2 (N369, N333, N283);
nor NOR3 (N370, N363, N207, N54);
not NOT1 (N371, N355);
or OR2 (N372, N338, N110);
buf BUF1 (N373, N345);
xor XOR2 (N374, N371, N273);
not NOT1 (N375, N373);
or OR3 (N376, N374, N300, N312);
buf BUF1 (N377, N367);
not NOT1 (N378, N354);
nor NOR3 (N379, N378, N283, N160);
xor XOR2 (N380, N376, N67);
nand NAND2 (N381, N372, N226);
and AND2 (N382, N377, N286);
buf BUF1 (N383, N362);
not NOT1 (N384, N383);
not NOT1 (N385, N381);
xor XOR2 (N386, N380, N61);
nand NAND2 (N387, N386, N249);
not NOT1 (N388, N384);
buf BUF1 (N389, N387);
or OR4 (N390, N369, N190, N110, N214);
and AND3 (N391, N370, N382, N306);
nand NAND4 (N392, N311, N204, N370, N208);
not NOT1 (N393, N392);
buf BUF1 (N394, N375);
not NOT1 (N395, N357);
not NOT1 (N396, N368);
buf BUF1 (N397, N390);
xor XOR2 (N398, N389, N283);
buf BUF1 (N399, N398);
not NOT1 (N400, N394);
xor XOR2 (N401, N395, N281);
nand NAND4 (N402, N397, N305, N326, N110);
not NOT1 (N403, N401);
xor XOR2 (N404, N402, N301);
or OR2 (N405, N388, N315);
nor NOR4 (N406, N391, N292, N291, N265);
not NOT1 (N407, N404);
nand NAND2 (N408, N379, N91);
buf BUF1 (N409, N396);
xor XOR2 (N410, N385, N175);
and AND2 (N411, N406, N63);
nor NOR2 (N412, N400, N254);
or OR2 (N413, N408, N178);
nand NAND2 (N414, N412, N38);
endmodule