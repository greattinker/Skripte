// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N1511,N1518,N1522,N1499,N1519,N1507,N1504,N1520,N1516,N1523;

nand NAND4 (N24, N11, N13, N22, N16);
and AND2 (N25, N15, N1);
xor XOR2 (N26, N20, N11);
and AND2 (N27, N12, N10);
nand NAND4 (N28, N15, N15, N5, N21);
or OR2 (N29, N19, N26);
and AND2 (N30, N8, N12);
nand NAND4 (N31, N25, N21, N7, N3);
not NOT1 (N32, N20);
nor NOR3 (N33, N30, N21, N32);
nor NOR4 (N34, N12, N27, N22, N22);
not NOT1 (N35, N6);
nand NAND3 (N36, N32, N27, N15);
and AND3 (N37, N26, N28, N28);
and AND4 (N38, N30, N33, N26, N28);
or OR4 (N39, N12, N23, N35, N18);
not NOT1 (N40, N2);
or OR4 (N41, N20, N5, N16, N27);
or OR2 (N42, N24, N16);
nand NAND4 (N43, N41, N34, N31, N15);
not NOT1 (N44, N31);
not NOT1 (N45, N1);
and AND3 (N46, N43, N36, N33);
and AND3 (N47, N36, N39, N17);
xor XOR2 (N48, N10, N28);
nand NAND2 (N49, N48, N48);
or OR4 (N50, N42, N18, N15, N18);
and AND4 (N51, N38, N7, N31, N23);
nor NOR3 (N52, N50, N39, N24);
or OR3 (N53, N51, N37, N51);
or OR4 (N54, N27, N3, N52, N14);
and AND4 (N55, N3, N25, N9, N14);
xor XOR2 (N56, N29, N16);
or OR4 (N57, N47, N53, N3, N36);
xor XOR2 (N58, N15, N28);
and AND3 (N59, N56, N34, N57);
xor XOR2 (N60, N48, N59);
not NOT1 (N61, N54);
nand NAND4 (N62, N40, N61, N49, N2);
nor NOR4 (N63, N46, N27, N29, N45);
buf BUF1 (N64, N22);
xor XOR2 (N65, N8, N53);
nand NAND4 (N66, N63, N18, N55, N11);
nand NAND2 (N67, N53, N24);
not NOT1 (N68, N66);
buf BUF1 (N69, N11);
xor XOR2 (N70, N11, N20);
buf BUF1 (N71, N64);
or OR4 (N72, N68, N20, N17, N10);
not NOT1 (N73, N44);
buf BUF1 (N74, N62);
and AND2 (N75, N71, N54);
and AND3 (N76, N67, N74, N10);
xor XOR2 (N77, N36, N55);
nor NOR4 (N78, N70, N37, N62, N21);
nand NAND4 (N79, N77, N24, N69, N11);
not NOT1 (N80, N49);
not NOT1 (N81, N73);
nand NAND3 (N82, N65, N52, N8);
nor NOR2 (N83, N78, N5);
xor XOR2 (N84, N79, N51);
nor NOR4 (N85, N72, N1, N26, N51);
buf BUF1 (N86, N83);
or OR2 (N87, N86, N14);
and AND4 (N88, N60, N40, N23, N53);
or OR2 (N89, N82, N9);
buf BUF1 (N90, N80);
xor XOR2 (N91, N88, N76);
buf BUF1 (N92, N91);
or OR2 (N93, N79, N6);
nand NAND2 (N94, N93, N83);
nor NOR2 (N95, N58, N40);
xor XOR2 (N96, N87, N53);
or OR2 (N97, N84, N69);
and AND2 (N98, N90, N79);
nand NAND4 (N99, N98, N14, N18, N85);
nand NAND4 (N100, N10, N2, N84, N55);
xor XOR2 (N101, N99, N79);
nand NAND3 (N102, N89, N65, N19);
xor XOR2 (N103, N75, N88);
or OR3 (N104, N103, N79, N93);
nor NOR2 (N105, N81, N60);
xor XOR2 (N106, N105, N25);
not NOT1 (N107, N95);
buf BUF1 (N108, N102);
nand NAND2 (N109, N92, N67);
and AND4 (N110, N94, N41, N24, N31);
nor NOR3 (N111, N96, N96, N89);
nor NOR2 (N112, N111, N56);
buf BUF1 (N113, N97);
buf BUF1 (N114, N110);
nand NAND2 (N115, N100, N80);
xor XOR2 (N116, N109, N43);
nand NAND4 (N117, N113, N41, N13, N22);
xor XOR2 (N118, N112, N78);
nor NOR3 (N119, N116, N97, N36);
buf BUF1 (N120, N101);
nor NOR4 (N121, N119, N103, N79, N14);
buf BUF1 (N122, N107);
nand NAND2 (N123, N118, N111);
buf BUF1 (N124, N104);
buf BUF1 (N125, N106);
xor XOR2 (N126, N121, N44);
xor XOR2 (N127, N108, N106);
nand NAND4 (N128, N124, N19, N2, N36);
or OR3 (N129, N122, N23, N60);
not NOT1 (N130, N129);
buf BUF1 (N131, N120);
buf BUF1 (N132, N128);
nor NOR3 (N133, N115, N62, N44);
xor XOR2 (N134, N127, N14);
nand NAND2 (N135, N114, N85);
nand NAND2 (N136, N125, N30);
nand NAND2 (N137, N132, N86);
buf BUF1 (N138, N126);
and AND4 (N139, N138, N18, N59, N64);
and AND2 (N140, N135, N139);
and AND2 (N141, N131, N110);
xor XOR2 (N142, N89, N58);
or OR4 (N143, N142, N100, N61, N4);
xor XOR2 (N144, N141, N21);
and AND4 (N145, N117, N7, N31, N110);
nor NOR2 (N146, N130, N103);
nand NAND2 (N147, N136, N141);
or OR3 (N148, N133, N29, N99);
and AND4 (N149, N143, N18, N90, N105);
nor NOR2 (N150, N145, N75);
and AND4 (N151, N150, N129, N130, N11);
nor NOR3 (N152, N147, N40, N36);
buf BUF1 (N153, N148);
and AND2 (N154, N153, N83);
not NOT1 (N155, N149);
xor XOR2 (N156, N146, N38);
not NOT1 (N157, N140);
nor NOR4 (N158, N156, N7, N77, N54);
and AND3 (N159, N155, N100, N88);
xor XOR2 (N160, N159, N41);
or OR2 (N161, N157, N16);
buf BUF1 (N162, N158);
or OR2 (N163, N161, N133);
buf BUF1 (N164, N123);
or OR3 (N165, N151, N144, N10);
xor XOR2 (N166, N20, N154);
or OR4 (N167, N18, N99, N92, N37);
nand NAND4 (N168, N166, N113, N103, N22);
xor XOR2 (N169, N152, N131);
nand NAND4 (N170, N163, N87, N22, N73);
or OR2 (N171, N169, N24);
not NOT1 (N172, N137);
and AND3 (N173, N165, N120, N80);
nand NAND4 (N174, N173, N120, N100, N108);
or OR4 (N175, N162, N129, N131, N156);
nor NOR3 (N176, N171, N96, N164);
nor NOR3 (N177, N131, N130, N104);
not NOT1 (N178, N174);
xor XOR2 (N179, N178, N52);
and AND2 (N180, N167, N70);
and AND2 (N181, N172, N20);
and AND2 (N182, N181, N58);
nor NOR4 (N183, N134, N33, N127, N179);
buf BUF1 (N184, N20);
nand NAND3 (N185, N184, N156, N51);
buf BUF1 (N186, N177);
and AND3 (N187, N176, N86, N2);
xor XOR2 (N188, N183, N105);
xor XOR2 (N189, N175, N54);
not NOT1 (N190, N160);
nor NOR2 (N191, N187, N117);
xor XOR2 (N192, N190, N171);
or OR4 (N193, N191, N20, N37, N178);
nor NOR3 (N194, N188, N57, N190);
not NOT1 (N195, N180);
buf BUF1 (N196, N189);
nor NOR2 (N197, N193, N15);
nand NAND3 (N198, N197, N132, N102);
buf BUF1 (N199, N196);
nor NOR2 (N200, N198, N191);
or OR4 (N201, N185, N43, N151, N75);
not NOT1 (N202, N186);
nor NOR2 (N203, N202, N108);
not NOT1 (N204, N199);
not NOT1 (N205, N182);
nand NAND2 (N206, N194, N165);
and AND3 (N207, N203, N20, N196);
or OR4 (N208, N206, N154, N141, N164);
not NOT1 (N209, N204);
and AND2 (N210, N201, N198);
xor XOR2 (N211, N170, N33);
not NOT1 (N212, N205);
or OR4 (N213, N210, N4, N75, N197);
or OR2 (N214, N195, N13);
nor NOR4 (N215, N214, N170, N156, N4);
nor NOR2 (N216, N213, N131);
or OR4 (N217, N212, N86, N93, N126);
not NOT1 (N218, N200);
xor XOR2 (N219, N211, N101);
xor XOR2 (N220, N219, N190);
or OR4 (N221, N220, N175, N143, N126);
nor NOR3 (N222, N208, N193, N22);
xor XOR2 (N223, N222, N95);
and AND2 (N224, N207, N209);
not NOT1 (N225, N206);
nor NOR3 (N226, N192, N199, N137);
or OR4 (N227, N168, N173, N55, N90);
buf BUF1 (N228, N223);
not NOT1 (N229, N221);
nor NOR2 (N230, N226, N148);
buf BUF1 (N231, N228);
nand NAND2 (N232, N217, N127);
buf BUF1 (N233, N218);
and AND4 (N234, N231, N97, N163, N58);
xor XOR2 (N235, N225, N76);
not NOT1 (N236, N216);
not NOT1 (N237, N234);
nor NOR4 (N238, N230, N156, N136, N185);
nand NAND4 (N239, N236, N2, N134, N166);
and AND3 (N240, N237, N172, N25);
buf BUF1 (N241, N238);
buf BUF1 (N242, N227);
nor NOR2 (N243, N229, N204);
xor XOR2 (N244, N232, N100);
not NOT1 (N245, N240);
or OR3 (N246, N241, N197, N50);
nand NAND4 (N247, N244, N84, N33, N233);
nor NOR4 (N248, N90, N29, N34, N157);
or OR4 (N249, N245, N141, N162, N153);
nand NAND3 (N250, N247, N218, N42);
or OR2 (N251, N246, N145);
and AND3 (N252, N251, N175, N139);
and AND3 (N253, N252, N146, N89);
or OR2 (N254, N215, N250);
not NOT1 (N255, N166);
nor NOR2 (N256, N243, N1);
buf BUF1 (N257, N248);
not NOT1 (N258, N255);
xor XOR2 (N259, N242, N165);
or OR4 (N260, N224, N101, N203, N52);
not NOT1 (N261, N258);
nand NAND4 (N262, N253, N8, N154, N141);
nand NAND4 (N263, N260, N124, N253, N78);
and AND2 (N264, N261, N70);
nor NOR4 (N265, N259, N201, N163, N125);
and AND2 (N266, N257, N203);
nand NAND3 (N267, N254, N175, N229);
nand NAND3 (N268, N256, N166, N38);
not NOT1 (N269, N262);
and AND2 (N270, N268, N127);
buf BUF1 (N271, N263);
buf BUF1 (N272, N270);
or OR3 (N273, N264, N231, N26);
or OR3 (N274, N273, N173, N11);
or OR4 (N275, N266, N212, N274, N230);
or OR3 (N276, N195, N73, N12);
nor NOR3 (N277, N235, N176, N64);
nor NOR3 (N278, N271, N129, N80);
not NOT1 (N279, N275);
and AND3 (N280, N267, N22, N25);
or OR4 (N281, N265, N190, N264, N220);
buf BUF1 (N282, N269);
not NOT1 (N283, N278);
and AND4 (N284, N272, N53, N139, N71);
xor XOR2 (N285, N279, N195);
or OR2 (N286, N283, N255);
nand NAND2 (N287, N249, N81);
and AND3 (N288, N239, N55, N153);
or OR3 (N289, N281, N216, N167);
xor XOR2 (N290, N277, N95);
nor NOR3 (N291, N282, N15, N124);
not NOT1 (N292, N287);
not NOT1 (N293, N284);
or OR3 (N294, N276, N152, N150);
and AND4 (N295, N294, N31, N207, N127);
nor NOR4 (N296, N285, N178, N235, N52);
nand NAND4 (N297, N292, N59, N33, N133);
nand NAND2 (N298, N291, N257);
buf BUF1 (N299, N289);
buf BUF1 (N300, N286);
not NOT1 (N301, N299);
or OR2 (N302, N288, N260);
xor XOR2 (N303, N300, N262);
xor XOR2 (N304, N290, N197);
not NOT1 (N305, N296);
and AND3 (N306, N295, N245, N80);
and AND2 (N307, N302, N68);
nor NOR3 (N308, N298, N185, N125);
xor XOR2 (N309, N280, N60);
xor XOR2 (N310, N303, N143);
or OR2 (N311, N307, N114);
nor NOR3 (N312, N301, N151, N146);
and AND3 (N313, N297, N119, N42);
or OR2 (N314, N312, N262);
or OR3 (N315, N311, N150, N208);
not NOT1 (N316, N308);
nor NOR2 (N317, N304, N104);
xor XOR2 (N318, N310, N212);
nand NAND3 (N319, N318, N316, N256);
or OR4 (N320, N65, N316, N296, N205);
or OR4 (N321, N313, N147, N30, N38);
nor NOR3 (N322, N309, N120, N186);
not NOT1 (N323, N293);
xor XOR2 (N324, N321, N68);
not NOT1 (N325, N315);
xor XOR2 (N326, N314, N298);
nand NAND2 (N327, N322, N51);
or OR4 (N328, N317, N50, N291, N54);
or OR4 (N329, N306, N165, N159, N5);
buf BUF1 (N330, N325);
or OR2 (N331, N327, N130);
xor XOR2 (N332, N305, N308);
buf BUF1 (N333, N323);
not NOT1 (N334, N328);
buf BUF1 (N335, N320);
and AND2 (N336, N334, N227);
nor NOR2 (N337, N336, N84);
buf BUF1 (N338, N333);
buf BUF1 (N339, N335);
buf BUF1 (N340, N337);
nor NOR2 (N341, N338, N128);
nand NAND2 (N342, N339, N24);
buf BUF1 (N343, N326);
and AND4 (N344, N319, N314, N71, N146);
nand NAND2 (N345, N330, N341);
not NOT1 (N346, N224);
and AND4 (N347, N324, N191, N257, N102);
buf BUF1 (N348, N342);
xor XOR2 (N349, N345, N219);
buf BUF1 (N350, N332);
nor NOR2 (N351, N350, N269);
nor NOR3 (N352, N329, N208, N298);
or OR2 (N353, N340, N29);
or OR2 (N354, N347, N307);
and AND4 (N355, N331, N178, N203, N336);
xor XOR2 (N356, N351, N216);
nand NAND2 (N357, N354, N320);
xor XOR2 (N358, N343, N240);
not NOT1 (N359, N344);
xor XOR2 (N360, N349, N20);
not NOT1 (N361, N355);
or OR3 (N362, N359, N16, N152);
and AND4 (N363, N361, N147, N71, N20);
buf BUF1 (N364, N356);
nand NAND4 (N365, N360, N254, N362, N152);
nand NAND2 (N366, N148, N127);
or OR2 (N367, N346, N125);
and AND4 (N368, N352, N298, N196, N31);
nor NOR3 (N369, N365, N275, N195);
nor NOR4 (N370, N357, N228, N320, N214);
and AND4 (N371, N370, N254, N305, N187);
and AND2 (N372, N358, N264);
not NOT1 (N373, N353);
nand NAND2 (N374, N368, N282);
xor XOR2 (N375, N364, N350);
or OR2 (N376, N372, N351);
not NOT1 (N377, N374);
and AND4 (N378, N371, N249, N16, N125);
not NOT1 (N379, N366);
xor XOR2 (N380, N375, N241);
buf BUF1 (N381, N376);
buf BUF1 (N382, N381);
nand NAND2 (N383, N378, N59);
not NOT1 (N384, N383);
and AND2 (N385, N369, N52);
or OR4 (N386, N380, N75, N380, N173);
not NOT1 (N387, N348);
not NOT1 (N388, N373);
not NOT1 (N389, N385);
or OR4 (N390, N386, N356, N23, N310);
buf BUF1 (N391, N367);
nand NAND3 (N392, N379, N390, N23);
not NOT1 (N393, N299);
and AND3 (N394, N391, N219, N51);
or OR2 (N395, N389, N5);
buf BUF1 (N396, N387);
or OR4 (N397, N395, N300, N304, N208);
nand NAND4 (N398, N384, N24, N198, N392);
nand NAND2 (N399, N216, N105);
nor NOR2 (N400, N388, N55);
not NOT1 (N401, N393);
nand NAND2 (N402, N396, N293);
not NOT1 (N403, N401);
nand NAND3 (N404, N363, N134, N237);
buf BUF1 (N405, N382);
nor NOR2 (N406, N398, N385);
nand NAND4 (N407, N377, N338, N32, N383);
or OR4 (N408, N402, N96, N22, N128);
and AND3 (N409, N404, N365, N292);
nor NOR4 (N410, N409, N113, N353, N153);
xor XOR2 (N411, N410, N58);
or OR3 (N412, N394, N406, N357);
nor NOR2 (N413, N136, N390);
buf BUF1 (N414, N400);
and AND4 (N415, N397, N67, N254, N396);
and AND3 (N416, N399, N385, N288);
nor NOR2 (N417, N415, N330);
not NOT1 (N418, N403);
buf BUF1 (N419, N414);
xor XOR2 (N420, N413, N27);
buf BUF1 (N421, N416);
not NOT1 (N422, N417);
buf BUF1 (N423, N408);
not NOT1 (N424, N411);
nand NAND3 (N425, N422, N112, N388);
and AND3 (N426, N425, N45, N222);
xor XOR2 (N427, N421, N423);
nand NAND3 (N428, N298, N324, N9);
and AND2 (N429, N419, N238);
nand NAND3 (N430, N428, N415, N8);
buf BUF1 (N431, N430);
not NOT1 (N432, N429);
xor XOR2 (N433, N412, N237);
nand NAND2 (N434, N424, N261);
xor XOR2 (N435, N426, N185);
not NOT1 (N436, N427);
and AND3 (N437, N405, N33, N349);
and AND2 (N438, N433, N58);
nor NOR2 (N439, N435, N278);
xor XOR2 (N440, N436, N169);
nor NOR3 (N441, N432, N146, N406);
not NOT1 (N442, N407);
not NOT1 (N443, N439);
nand NAND3 (N444, N440, N425, N40);
and AND3 (N445, N441, N425, N38);
xor XOR2 (N446, N434, N417);
or OR4 (N447, N445, N44, N109, N265);
not NOT1 (N448, N437);
xor XOR2 (N449, N448, N288);
or OR3 (N450, N443, N104, N69);
buf BUF1 (N451, N447);
and AND2 (N452, N451, N382);
buf BUF1 (N453, N450);
nor NOR2 (N454, N438, N205);
buf BUF1 (N455, N420);
buf BUF1 (N456, N453);
buf BUF1 (N457, N418);
nor NOR2 (N458, N457, N289);
nor NOR3 (N459, N444, N424, N212);
buf BUF1 (N460, N446);
xor XOR2 (N461, N459, N295);
or OR2 (N462, N442, N7);
and AND2 (N463, N431, N352);
nor NOR4 (N464, N452, N226, N205, N110);
or OR3 (N465, N458, N387, N224);
or OR3 (N466, N461, N297, N290);
or OR2 (N467, N465, N146);
xor XOR2 (N468, N456, N243);
and AND3 (N469, N464, N274, N102);
or OR3 (N470, N449, N17, N346);
nand NAND4 (N471, N462, N147, N220, N387);
buf BUF1 (N472, N468);
nand NAND4 (N473, N467, N193, N62, N394);
buf BUF1 (N474, N466);
nand NAND4 (N475, N455, N132, N32, N374);
and AND3 (N476, N460, N136, N292);
nor NOR4 (N477, N472, N419, N310, N27);
buf BUF1 (N478, N476);
and AND4 (N479, N477, N452, N466, N184);
nor NOR3 (N480, N478, N321, N442);
not NOT1 (N481, N454);
not NOT1 (N482, N469);
nand NAND3 (N483, N481, N86, N43);
nor NOR2 (N484, N470, N263);
or OR4 (N485, N474, N308, N356, N78);
not NOT1 (N486, N485);
nand NAND3 (N487, N484, N417, N147);
buf BUF1 (N488, N482);
or OR4 (N489, N483, N246, N233, N57);
nand NAND4 (N490, N489, N43, N143, N471);
buf BUF1 (N491, N338);
xor XOR2 (N492, N463, N444);
buf BUF1 (N493, N490);
nor NOR3 (N494, N473, N153, N342);
nor NOR2 (N495, N487, N469);
and AND2 (N496, N486, N478);
nand NAND2 (N497, N480, N70);
nor NOR2 (N498, N491, N310);
and AND4 (N499, N488, N454, N281, N297);
and AND4 (N500, N479, N377, N285, N229);
nor NOR3 (N501, N497, N453, N432);
xor XOR2 (N502, N494, N163);
or OR3 (N503, N492, N207, N273);
and AND2 (N504, N502, N424);
nand NAND3 (N505, N500, N440, N455);
buf BUF1 (N506, N499);
nand NAND2 (N507, N493, N245);
xor XOR2 (N508, N501, N181);
not NOT1 (N509, N503);
nor NOR3 (N510, N498, N291, N27);
nand NAND4 (N511, N507, N506, N484, N318);
buf BUF1 (N512, N37);
xor XOR2 (N513, N495, N162);
nand NAND3 (N514, N496, N69, N333);
not NOT1 (N515, N514);
and AND2 (N516, N511, N174);
nand NAND2 (N517, N508, N158);
buf BUF1 (N518, N512);
nand NAND3 (N519, N515, N476, N471);
or OR2 (N520, N517, N56);
buf BUF1 (N521, N475);
or OR4 (N522, N518, N339, N509, N113);
and AND4 (N523, N315, N300, N169, N250);
nor NOR4 (N524, N519, N329, N448, N355);
buf BUF1 (N525, N523);
xor XOR2 (N526, N505, N262);
buf BUF1 (N527, N510);
nand NAND3 (N528, N504, N35, N304);
or OR3 (N529, N528, N230, N73);
and AND2 (N530, N525, N325);
xor XOR2 (N531, N524, N318);
or OR2 (N532, N530, N482);
not NOT1 (N533, N529);
and AND4 (N534, N513, N8, N495, N278);
buf BUF1 (N535, N526);
not NOT1 (N536, N522);
nand NAND4 (N537, N520, N404, N255, N286);
not NOT1 (N538, N531);
not NOT1 (N539, N521);
nor NOR2 (N540, N539, N426);
buf BUF1 (N541, N535);
nand NAND4 (N542, N538, N7, N428, N62);
xor XOR2 (N543, N537, N205);
and AND4 (N544, N542, N448, N393, N81);
buf BUF1 (N545, N536);
nand NAND4 (N546, N533, N351, N141, N389);
nand NAND2 (N547, N532, N274);
nand NAND2 (N548, N527, N179);
and AND3 (N549, N544, N234, N252);
buf BUF1 (N550, N540);
nor NOR3 (N551, N549, N409, N452);
not NOT1 (N552, N534);
and AND4 (N553, N548, N129, N314, N514);
xor XOR2 (N554, N545, N155);
nor NOR3 (N555, N543, N369, N90);
or OR4 (N556, N554, N30, N207, N254);
and AND2 (N557, N555, N281);
xor XOR2 (N558, N547, N238);
not NOT1 (N559, N557);
and AND4 (N560, N516, N274, N265, N539);
or OR2 (N561, N541, N452);
nand NAND3 (N562, N553, N137, N356);
nand NAND3 (N563, N561, N279, N486);
not NOT1 (N564, N550);
not NOT1 (N565, N562);
nand NAND3 (N566, N559, N285, N183);
not NOT1 (N567, N546);
or OR4 (N568, N556, N339, N172, N449);
buf BUF1 (N569, N568);
buf BUF1 (N570, N566);
nand NAND2 (N571, N564, N56);
not NOT1 (N572, N570);
or OR3 (N573, N571, N226, N26);
nor NOR3 (N574, N573, N415, N384);
or OR4 (N575, N552, N330, N271, N348);
nor NOR4 (N576, N567, N273, N501, N434);
nor NOR2 (N577, N563, N411);
xor XOR2 (N578, N551, N575);
nand NAND2 (N579, N381, N298);
not NOT1 (N580, N574);
and AND3 (N581, N572, N169, N376);
xor XOR2 (N582, N581, N116);
and AND2 (N583, N579, N73);
and AND4 (N584, N560, N220, N8, N228);
nor NOR3 (N585, N583, N381, N242);
nand NAND2 (N586, N577, N503);
and AND4 (N587, N580, N167, N87, N519);
or OR4 (N588, N582, N119, N362, N241);
nand NAND4 (N589, N588, N76, N203, N558);
and AND3 (N590, N525, N410, N200);
and AND4 (N591, N576, N393, N12, N1);
nand NAND3 (N592, N584, N94, N450);
not NOT1 (N593, N578);
xor XOR2 (N594, N586, N223);
not NOT1 (N595, N589);
or OR4 (N596, N594, N306, N79, N374);
not NOT1 (N597, N587);
xor XOR2 (N598, N597, N127);
or OR4 (N599, N598, N156, N246, N355);
or OR3 (N600, N569, N107, N462);
buf BUF1 (N601, N585);
not NOT1 (N602, N596);
not NOT1 (N603, N600);
and AND3 (N604, N591, N558, N48);
or OR3 (N605, N593, N362, N124);
and AND2 (N606, N599, N82);
or OR3 (N607, N606, N379, N556);
not NOT1 (N608, N601);
not NOT1 (N609, N565);
xor XOR2 (N610, N605, N177);
or OR4 (N611, N609, N196, N430, N607);
nor NOR4 (N612, N301, N420, N68, N336);
and AND4 (N613, N608, N170, N612, N190);
or OR2 (N614, N151, N238);
not NOT1 (N615, N613);
not NOT1 (N616, N604);
not NOT1 (N617, N602);
nand NAND2 (N618, N611, N585);
not NOT1 (N619, N592);
buf BUF1 (N620, N595);
nand NAND3 (N621, N619, N152, N620);
nor NOR3 (N622, N114, N508, N32);
xor XOR2 (N623, N590, N497);
nor NOR3 (N624, N614, N144, N22);
xor XOR2 (N625, N623, N550);
nor NOR2 (N626, N624, N378);
and AND2 (N627, N626, N598);
not NOT1 (N628, N617);
and AND4 (N629, N610, N506, N559, N184);
nand NAND2 (N630, N618, N489);
nand NAND2 (N631, N621, N61);
buf BUF1 (N632, N603);
or OR3 (N633, N630, N630, N575);
xor XOR2 (N634, N631, N287);
xor XOR2 (N635, N633, N508);
nor NOR3 (N636, N628, N558, N83);
or OR2 (N637, N636, N628);
and AND2 (N638, N622, N419);
or OR4 (N639, N637, N285, N309, N313);
or OR4 (N640, N629, N601, N416, N606);
nand NAND4 (N641, N639, N636, N285, N564);
or OR3 (N642, N634, N598, N317);
or OR3 (N643, N627, N619, N261);
or OR3 (N644, N640, N612, N435);
nand NAND3 (N645, N642, N252, N473);
not NOT1 (N646, N632);
xor XOR2 (N647, N625, N625);
nand NAND3 (N648, N643, N136, N489);
not NOT1 (N649, N641);
not NOT1 (N650, N647);
buf BUF1 (N651, N648);
and AND2 (N652, N651, N101);
xor XOR2 (N653, N644, N372);
buf BUF1 (N654, N635);
buf BUF1 (N655, N638);
nor NOR2 (N656, N652, N139);
and AND2 (N657, N615, N314);
buf BUF1 (N658, N650);
xor XOR2 (N659, N646, N72);
or OR3 (N660, N656, N580, N633);
or OR4 (N661, N657, N181, N660, N564);
nand NAND3 (N662, N186, N481, N108);
not NOT1 (N663, N645);
nor NOR4 (N664, N616, N589, N594, N603);
and AND2 (N665, N653, N124);
nand NAND3 (N666, N655, N374, N77);
xor XOR2 (N667, N659, N298);
nand NAND4 (N668, N667, N620, N337, N448);
xor XOR2 (N669, N664, N178);
buf BUF1 (N670, N668);
nor NOR4 (N671, N669, N576, N656, N670);
nor NOR2 (N672, N219, N483);
nand NAND4 (N673, N654, N324, N490, N274);
xor XOR2 (N674, N666, N28);
buf BUF1 (N675, N671);
and AND3 (N676, N675, N164, N206);
nand NAND2 (N677, N658, N613);
and AND4 (N678, N673, N473, N509, N110);
buf BUF1 (N679, N661);
buf BUF1 (N680, N665);
xor XOR2 (N681, N676, N199);
nor NOR4 (N682, N674, N341, N320, N124);
nor NOR4 (N683, N649, N230, N358, N269);
nor NOR4 (N684, N683, N493, N412, N527);
xor XOR2 (N685, N663, N129);
not NOT1 (N686, N678);
nand NAND2 (N687, N682, N327);
and AND3 (N688, N681, N475, N586);
xor XOR2 (N689, N672, N88);
nor NOR2 (N690, N685, N225);
not NOT1 (N691, N662);
xor XOR2 (N692, N687, N488);
xor XOR2 (N693, N692, N585);
not NOT1 (N694, N679);
xor XOR2 (N695, N690, N182);
and AND3 (N696, N691, N374, N616);
xor XOR2 (N697, N686, N72);
buf BUF1 (N698, N688);
buf BUF1 (N699, N698);
nor NOR3 (N700, N684, N517, N367);
nand NAND2 (N701, N689, N332);
nor NOR3 (N702, N695, N471, N257);
xor XOR2 (N703, N677, N589);
nor NOR2 (N704, N697, N421);
xor XOR2 (N705, N696, N302);
and AND3 (N706, N694, N637, N132);
not NOT1 (N707, N705);
buf BUF1 (N708, N701);
and AND4 (N709, N700, N383, N88, N6);
buf BUF1 (N710, N702);
and AND3 (N711, N704, N377, N244);
buf BUF1 (N712, N706);
nor NOR2 (N713, N707, N161);
nor NOR3 (N714, N699, N242, N713);
nand NAND2 (N715, N151, N536);
xor XOR2 (N716, N711, N248);
xor XOR2 (N717, N693, N277);
nand NAND4 (N718, N712, N379, N201, N209);
xor XOR2 (N719, N716, N704);
nand NAND3 (N720, N714, N30, N468);
xor XOR2 (N721, N719, N104);
xor XOR2 (N722, N715, N560);
nor NOR3 (N723, N710, N419, N274);
nand NAND3 (N724, N703, N651, N454);
buf BUF1 (N725, N718);
nor NOR2 (N726, N723, N568);
not NOT1 (N727, N722);
xor XOR2 (N728, N680, N240);
or OR2 (N729, N726, N706);
nand NAND4 (N730, N720, N487, N530, N236);
nor NOR3 (N731, N724, N222, N168);
nor NOR4 (N732, N731, N58, N215, N168);
and AND3 (N733, N728, N395, N671);
xor XOR2 (N734, N727, N201);
xor XOR2 (N735, N721, N636);
nor NOR2 (N736, N733, N197);
or OR2 (N737, N708, N310);
not NOT1 (N738, N730);
and AND3 (N739, N717, N529, N149);
and AND4 (N740, N738, N82, N705, N248);
xor XOR2 (N741, N709, N11);
and AND3 (N742, N734, N603, N538);
not NOT1 (N743, N742);
xor XOR2 (N744, N729, N595);
or OR3 (N745, N744, N646, N723);
not NOT1 (N746, N743);
and AND3 (N747, N732, N363, N730);
nand NAND3 (N748, N746, N479, N151);
buf BUF1 (N749, N740);
or OR2 (N750, N739, N7);
buf BUF1 (N751, N736);
buf BUF1 (N752, N725);
not NOT1 (N753, N737);
nand NAND4 (N754, N735, N69, N687, N407);
xor XOR2 (N755, N741, N388);
nand NAND4 (N756, N750, N24, N64, N210);
buf BUF1 (N757, N747);
and AND4 (N758, N753, N195, N126, N137);
and AND4 (N759, N751, N82, N534, N338);
xor XOR2 (N760, N758, N241);
not NOT1 (N761, N748);
or OR4 (N762, N760, N589, N438, N594);
nor NOR3 (N763, N757, N260, N596);
and AND3 (N764, N756, N206, N385);
not NOT1 (N765, N759);
or OR4 (N766, N749, N469, N438, N300);
or OR3 (N767, N755, N654, N443);
nor NOR2 (N768, N763, N668);
not NOT1 (N769, N762);
not NOT1 (N770, N768);
nor NOR4 (N771, N770, N338, N525, N193);
not NOT1 (N772, N766);
xor XOR2 (N773, N771, N61);
buf BUF1 (N774, N767);
buf BUF1 (N775, N769);
buf BUF1 (N776, N774);
not NOT1 (N777, N773);
not NOT1 (N778, N777);
nand NAND3 (N779, N761, N8, N92);
buf BUF1 (N780, N776);
xor XOR2 (N781, N764, N112);
nand NAND4 (N782, N775, N351, N496, N154);
or OR2 (N783, N745, N584);
xor XOR2 (N784, N779, N196);
or OR3 (N785, N765, N199, N696);
xor XOR2 (N786, N784, N273);
xor XOR2 (N787, N782, N504);
not NOT1 (N788, N787);
or OR2 (N789, N780, N772);
nor NOR3 (N790, N433, N114, N299);
nor NOR3 (N791, N786, N71, N503);
or OR4 (N792, N783, N210, N769, N240);
nand NAND2 (N793, N788, N28);
buf BUF1 (N794, N793);
xor XOR2 (N795, N794, N454);
not NOT1 (N796, N792);
not NOT1 (N797, N791);
or OR3 (N798, N790, N329, N201);
and AND4 (N799, N781, N200, N126, N37);
nor NOR2 (N800, N797, N149);
nor NOR3 (N801, N789, N770, N76);
xor XOR2 (N802, N796, N199);
nor NOR3 (N803, N754, N62, N63);
or OR3 (N804, N798, N426, N275);
xor XOR2 (N805, N752, N783);
xor XOR2 (N806, N801, N648);
or OR4 (N807, N805, N199, N552, N751);
not NOT1 (N808, N804);
or OR4 (N809, N806, N433, N646, N609);
xor XOR2 (N810, N778, N748);
or OR4 (N811, N799, N625, N347, N785);
buf BUF1 (N812, N353);
xor XOR2 (N813, N803, N380);
buf BUF1 (N814, N812);
or OR3 (N815, N814, N89, N18);
or OR3 (N816, N800, N461, N145);
or OR2 (N817, N815, N294);
not NOT1 (N818, N795);
xor XOR2 (N819, N817, N205);
buf BUF1 (N820, N816);
xor XOR2 (N821, N818, N549);
not NOT1 (N822, N821);
xor XOR2 (N823, N807, N553);
xor XOR2 (N824, N823, N529);
nand NAND3 (N825, N808, N725, N196);
xor XOR2 (N826, N820, N261);
not NOT1 (N827, N810);
not NOT1 (N828, N827);
and AND3 (N829, N822, N405, N186);
not NOT1 (N830, N802);
or OR3 (N831, N830, N317, N339);
not NOT1 (N832, N811);
nor NOR4 (N833, N831, N181, N75, N393);
buf BUF1 (N834, N825);
or OR3 (N835, N819, N550, N346);
and AND3 (N836, N835, N123, N134);
xor XOR2 (N837, N813, N418);
nand NAND2 (N838, N834, N80);
and AND3 (N839, N833, N482, N436);
or OR4 (N840, N838, N264, N73, N489);
and AND3 (N841, N832, N268, N64);
nor NOR2 (N842, N829, N745);
nand NAND2 (N843, N824, N162);
not NOT1 (N844, N840);
and AND2 (N845, N844, N233);
nor NOR2 (N846, N841, N254);
xor XOR2 (N847, N809, N515);
not NOT1 (N848, N828);
not NOT1 (N849, N842);
or OR2 (N850, N848, N844);
buf BUF1 (N851, N837);
and AND4 (N852, N846, N558, N577, N745);
nor NOR3 (N853, N849, N494, N43);
and AND2 (N854, N826, N141);
xor XOR2 (N855, N847, N333);
buf BUF1 (N856, N850);
or OR2 (N857, N855, N138);
and AND2 (N858, N839, N385);
nor NOR4 (N859, N858, N537, N466, N610);
buf BUF1 (N860, N845);
xor XOR2 (N861, N857, N105);
xor XOR2 (N862, N851, N636);
not NOT1 (N863, N861);
nand NAND2 (N864, N852, N76);
not NOT1 (N865, N863);
or OR3 (N866, N859, N767, N179);
buf BUF1 (N867, N856);
and AND4 (N868, N862, N361, N715, N243);
not NOT1 (N869, N864);
buf BUF1 (N870, N865);
nand NAND2 (N871, N869, N691);
nor NOR3 (N872, N836, N384, N458);
nand NAND3 (N873, N867, N846, N802);
not NOT1 (N874, N873);
xor XOR2 (N875, N866, N721);
not NOT1 (N876, N874);
and AND2 (N877, N871, N563);
or OR2 (N878, N875, N143);
nand NAND2 (N879, N843, N735);
and AND3 (N880, N879, N3, N267);
and AND4 (N881, N878, N233, N591, N17);
xor XOR2 (N882, N853, N860);
xor XOR2 (N883, N454, N726);
buf BUF1 (N884, N883);
buf BUF1 (N885, N881);
buf BUF1 (N886, N877);
xor XOR2 (N887, N886, N501);
not NOT1 (N888, N872);
not NOT1 (N889, N854);
xor XOR2 (N890, N876, N156);
xor XOR2 (N891, N885, N477);
nor NOR4 (N892, N870, N12, N85, N368);
not NOT1 (N893, N888);
buf BUF1 (N894, N882);
nor NOR2 (N895, N892, N267);
not NOT1 (N896, N887);
or OR3 (N897, N890, N811, N281);
nor NOR4 (N898, N895, N511, N536, N296);
buf BUF1 (N899, N891);
buf BUF1 (N900, N893);
nand NAND4 (N901, N884, N718, N191, N531);
and AND2 (N902, N894, N182);
not NOT1 (N903, N899);
xor XOR2 (N904, N897, N141);
xor XOR2 (N905, N896, N659);
buf BUF1 (N906, N904);
xor XOR2 (N907, N903, N650);
nand NAND2 (N908, N880, N710);
xor XOR2 (N909, N908, N815);
and AND4 (N910, N898, N671, N381, N499);
buf BUF1 (N911, N868);
nor NOR2 (N912, N902, N711);
and AND2 (N913, N907, N179);
or OR2 (N914, N910, N228);
nand NAND3 (N915, N914, N847, N194);
or OR2 (N916, N905, N337);
not NOT1 (N917, N915);
or OR3 (N918, N909, N195, N362);
or OR4 (N919, N911, N682, N547, N599);
xor XOR2 (N920, N916, N185);
or OR2 (N921, N917, N449);
xor XOR2 (N922, N921, N556);
nor NOR3 (N923, N913, N902, N663);
or OR2 (N924, N889, N57);
buf BUF1 (N925, N901);
nand NAND4 (N926, N906, N124, N641, N55);
not NOT1 (N927, N918);
or OR3 (N928, N912, N915, N486);
nor NOR2 (N929, N919, N573);
nand NAND2 (N930, N928, N296);
and AND2 (N931, N926, N257);
not NOT1 (N932, N924);
nand NAND3 (N933, N922, N355, N139);
xor XOR2 (N934, N930, N484);
and AND3 (N935, N900, N832, N830);
nand NAND3 (N936, N920, N517, N219);
xor XOR2 (N937, N923, N557);
and AND3 (N938, N937, N792, N71);
xor XOR2 (N939, N934, N196);
xor XOR2 (N940, N933, N295);
not NOT1 (N941, N929);
or OR2 (N942, N940, N378);
buf BUF1 (N943, N925);
nand NAND2 (N944, N943, N43);
not NOT1 (N945, N938);
nor NOR4 (N946, N941, N360, N469, N877);
or OR2 (N947, N931, N559);
nor NOR4 (N948, N947, N757, N107, N896);
buf BUF1 (N949, N927);
nand NAND3 (N950, N948, N664, N758);
or OR2 (N951, N946, N861);
nor NOR2 (N952, N939, N71);
nor NOR2 (N953, N951, N819);
buf BUF1 (N954, N936);
nand NAND4 (N955, N954, N653, N601, N95);
nand NAND2 (N956, N949, N786);
not NOT1 (N957, N952);
nand NAND4 (N958, N942, N269, N857, N37);
xor XOR2 (N959, N950, N820);
or OR4 (N960, N957, N273, N717, N866);
nand NAND4 (N961, N959, N513, N572, N386);
or OR3 (N962, N961, N166, N237);
nand NAND4 (N963, N955, N656, N180, N20);
and AND3 (N964, N932, N505, N271);
xor XOR2 (N965, N945, N618);
nor NOR2 (N966, N960, N492);
nor NOR3 (N967, N964, N767, N746);
nor NOR4 (N968, N967, N270, N666, N962);
nand NAND4 (N969, N528, N718, N19, N872);
and AND2 (N970, N944, N253);
not NOT1 (N971, N969);
nand NAND2 (N972, N970, N160);
not NOT1 (N973, N966);
or OR4 (N974, N965, N109, N505, N380);
or OR4 (N975, N956, N544, N184, N39);
and AND3 (N976, N971, N234, N637);
nor NOR3 (N977, N968, N530, N275);
and AND3 (N978, N976, N163, N613);
xor XOR2 (N979, N963, N650);
xor XOR2 (N980, N958, N618);
buf BUF1 (N981, N978);
or OR4 (N982, N973, N9, N628, N713);
xor XOR2 (N983, N979, N191);
buf BUF1 (N984, N974);
xor XOR2 (N985, N984, N645);
or OR2 (N986, N977, N108);
xor XOR2 (N987, N980, N46);
xor XOR2 (N988, N953, N150);
buf BUF1 (N989, N972);
xor XOR2 (N990, N975, N743);
or OR4 (N991, N982, N85, N327, N150);
xor XOR2 (N992, N983, N891);
nand NAND4 (N993, N986, N83, N934, N96);
buf BUF1 (N994, N990);
buf BUF1 (N995, N991);
nor NOR4 (N996, N989, N794, N31, N27);
xor XOR2 (N997, N993, N125);
nand NAND2 (N998, N985, N912);
nand NAND4 (N999, N998, N597, N596, N324);
and AND4 (N1000, N994, N741, N288, N310);
nor NOR3 (N1001, N935, N971, N953);
not NOT1 (N1002, N995);
not NOT1 (N1003, N988);
or OR4 (N1004, N987, N43, N69, N320);
not NOT1 (N1005, N992);
xor XOR2 (N1006, N1002, N277);
buf BUF1 (N1007, N1001);
buf BUF1 (N1008, N997);
or OR3 (N1009, N981, N388, N399);
nand NAND3 (N1010, N1007, N951, N601);
nand NAND4 (N1011, N1006, N738, N76, N882);
or OR4 (N1012, N999, N835, N950, N867);
or OR4 (N1013, N1012, N262, N153, N107);
nor NOR3 (N1014, N1008, N696, N213);
not NOT1 (N1015, N1014);
or OR3 (N1016, N1013, N604, N124);
nor NOR2 (N1017, N1004, N301);
and AND4 (N1018, N1000, N537, N378, N440);
or OR4 (N1019, N1018, N127, N763, N639);
xor XOR2 (N1020, N1015, N413);
and AND4 (N1021, N1019, N820, N28, N86);
xor XOR2 (N1022, N1021, N865);
buf BUF1 (N1023, N1003);
or OR4 (N1024, N1005, N678, N274, N6);
nor NOR3 (N1025, N1010, N663, N280);
nor NOR2 (N1026, N1016, N977);
buf BUF1 (N1027, N1020);
xor XOR2 (N1028, N1025, N784);
and AND2 (N1029, N1011, N942);
nand NAND3 (N1030, N1028, N470, N566);
nand NAND2 (N1031, N1024, N852);
xor XOR2 (N1032, N1009, N246);
nand NAND2 (N1033, N1022, N853);
buf BUF1 (N1034, N1023);
and AND4 (N1035, N1029, N630, N952, N913);
or OR2 (N1036, N1034, N113);
buf BUF1 (N1037, N1027);
buf BUF1 (N1038, N1030);
nand NAND2 (N1039, N1035, N493);
not NOT1 (N1040, N1038);
and AND3 (N1041, N1017, N204, N886);
nand NAND2 (N1042, N996, N936);
or OR4 (N1043, N1041, N65, N789, N945);
not NOT1 (N1044, N1032);
nor NOR2 (N1045, N1031, N463);
and AND2 (N1046, N1039, N619);
buf BUF1 (N1047, N1042);
xor XOR2 (N1048, N1045, N673);
and AND2 (N1049, N1040, N359);
buf BUF1 (N1050, N1049);
buf BUF1 (N1051, N1044);
xor XOR2 (N1052, N1037, N334);
xor XOR2 (N1053, N1043, N699);
and AND4 (N1054, N1033, N546, N1036, N641);
buf BUF1 (N1055, N275);
xor XOR2 (N1056, N1047, N965);
not NOT1 (N1057, N1056);
xor XOR2 (N1058, N1052, N697);
and AND2 (N1059, N1050, N474);
and AND4 (N1060, N1046, N830, N682, N39);
xor XOR2 (N1061, N1059, N1025);
not NOT1 (N1062, N1053);
nor NOR3 (N1063, N1061, N632, N960);
and AND2 (N1064, N1062, N1037);
nor NOR4 (N1065, N1054, N777, N601, N416);
xor XOR2 (N1066, N1051, N848);
and AND3 (N1067, N1055, N613, N35);
xor XOR2 (N1068, N1066, N314);
not NOT1 (N1069, N1068);
not NOT1 (N1070, N1057);
buf BUF1 (N1071, N1048);
not NOT1 (N1072, N1071);
or OR2 (N1073, N1072, N971);
and AND4 (N1074, N1073, N1019, N512, N647);
nand NAND3 (N1075, N1067, N597, N327);
or OR4 (N1076, N1026, N271, N862, N812);
nand NAND3 (N1077, N1069, N81, N625);
not NOT1 (N1078, N1075);
not NOT1 (N1079, N1070);
nand NAND3 (N1080, N1063, N1041, N551);
nand NAND4 (N1081, N1077, N275, N994, N212);
buf BUF1 (N1082, N1065);
buf BUF1 (N1083, N1058);
or OR2 (N1084, N1076, N1046);
or OR2 (N1085, N1080, N963);
not NOT1 (N1086, N1060);
nand NAND2 (N1087, N1084, N497);
not NOT1 (N1088, N1083);
nand NAND2 (N1089, N1081, N488);
or OR4 (N1090, N1085, N1073, N359, N829);
or OR2 (N1091, N1089, N746);
nand NAND4 (N1092, N1064, N43, N355, N623);
and AND2 (N1093, N1090, N569);
xor XOR2 (N1094, N1092, N74);
nor NOR4 (N1095, N1078, N506, N298, N1093);
and AND2 (N1096, N817, N1077);
and AND3 (N1097, N1094, N875, N240);
xor XOR2 (N1098, N1096, N699);
xor XOR2 (N1099, N1091, N462);
or OR3 (N1100, N1079, N1028, N742);
nor NOR4 (N1101, N1099, N622, N597, N892);
buf BUF1 (N1102, N1100);
buf BUF1 (N1103, N1087);
or OR2 (N1104, N1086, N855);
and AND3 (N1105, N1102, N813, N885);
and AND4 (N1106, N1074, N861, N11, N296);
or OR2 (N1107, N1104, N410);
and AND3 (N1108, N1095, N642, N610);
nand NAND2 (N1109, N1105, N782);
or OR3 (N1110, N1108, N330, N540);
or OR4 (N1111, N1109, N820, N981, N854);
xor XOR2 (N1112, N1082, N33);
nand NAND2 (N1113, N1097, N412);
and AND2 (N1114, N1101, N365);
nor NOR3 (N1115, N1114, N442, N244);
xor XOR2 (N1116, N1103, N263);
or OR4 (N1117, N1115, N947, N854, N143);
or OR2 (N1118, N1113, N125);
not NOT1 (N1119, N1118);
nand NAND2 (N1120, N1088, N1103);
and AND2 (N1121, N1120, N1053);
nand NAND3 (N1122, N1121, N93, N439);
and AND4 (N1123, N1122, N583, N584, N471);
and AND2 (N1124, N1112, N736);
xor XOR2 (N1125, N1106, N949);
nor NOR3 (N1126, N1098, N656, N705);
xor XOR2 (N1127, N1126, N257);
nor NOR4 (N1128, N1125, N921, N476, N806);
or OR2 (N1129, N1111, N508);
buf BUF1 (N1130, N1107);
nor NOR4 (N1131, N1127, N665, N916, N275);
xor XOR2 (N1132, N1119, N784);
buf BUF1 (N1133, N1123);
not NOT1 (N1134, N1133);
buf BUF1 (N1135, N1132);
and AND3 (N1136, N1129, N186, N1114);
and AND4 (N1137, N1135, N373, N769, N569);
and AND3 (N1138, N1134, N29, N178);
and AND4 (N1139, N1131, N877, N43, N554);
buf BUF1 (N1140, N1136);
not NOT1 (N1141, N1116);
not NOT1 (N1142, N1141);
nor NOR3 (N1143, N1139, N322, N864);
and AND4 (N1144, N1138, N1070, N337, N740);
not NOT1 (N1145, N1142);
and AND2 (N1146, N1143, N169);
buf BUF1 (N1147, N1117);
nor NOR3 (N1148, N1128, N1010, N688);
or OR2 (N1149, N1148, N34);
and AND2 (N1150, N1124, N814);
xor XOR2 (N1151, N1137, N180);
or OR3 (N1152, N1110, N337, N412);
not NOT1 (N1153, N1151);
or OR4 (N1154, N1150, N370, N1070, N1021);
nor NOR3 (N1155, N1152, N207, N803);
nor NOR3 (N1156, N1146, N682, N997);
and AND4 (N1157, N1140, N248, N909, N208);
nor NOR4 (N1158, N1130, N790, N813, N549);
nand NAND3 (N1159, N1157, N112, N287);
nor NOR4 (N1160, N1159, N736, N444, N45);
nand NAND2 (N1161, N1145, N773);
or OR3 (N1162, N1149, N1135, N492);
buf BUF1 (N1163, N1160);
buf BUF1 (N1164, N1154);
xor XOR2 (N1165, N1155, N207);
nand NAND2 (N1166, N1156, N685);
xor XOR2 (N1167, N1144, N540);
not NOT1 (N1168, N1162);
not NOT1 (N1169, N1164);
nand NAND4 (N1170, N1161, N292, N85, N551);
nand NAND2 (N1171, N1167, N931);
xor XOR2 (N1172, N1147, N150);
nor NOR4 (N1173, N1171, N580, N933, N826);
nor NOR4 (N1174, N1170, N371, N68, N357);
buf BUF1 (N1175, N1168);
xor XOR2 (N1176, N1174, N496);
nand NAND4 (N1177, N1158, N266, N422, N968);
nand NAND3 (N1178, N1166, N519, N289);
buf BUF1 (N1179, N1169);
not NOT1 (N1180, N1176);
or OR3 (N1181, N1153, N558, N255);
or OR4 (N1182, N1178, N404, N37, N726);
xor XOR2 (N1183, N1165, N140);
buf BUF1 (N1184, N1180);
and AND2 (N1185, N1179, N988);
xor XOR2 (N1186, N1173, N355);
nand NAND3 (N1187, N1175, N988, N421);
and AND3 (N1188, N1185, N60, N677);
and AND2 (N1189, N1182, N237);
or OR2 (N1190, N1172, N1058);
and AND2 (N1191, N1189, N393);
and AND2 (N1192, N1163, N1063);
buf BUF1 (N1193, N1190);
xor XOR2 (N1194, N1191, N526);
xor XOR2 (N1195, N1194, N58);
nor NOR2 (N1196, N1181, N41);
nor NOR4 (N1197, N1196, N1062, N348, N711);
and AND2 (N1198, N1192, N544);
and AND4 (N1199, N1188, N895, N433, N665);
nor NOR3 (N1200, N1193, N288, N745);
not NOT1 (N1201, N1199);
and AND4 (N1202, N1187, N483, N1134, N1039);
or OR4 (N1203, N1177, N983, N1079, N540);
xor XOR2 (N1204, N1197, N840);
nor NOR4 (N1205, N1195, N131, N1079, N378);
nand NAND2 (N1206, N1184, N814);
not NOT1 (N1207, N1186);
nor NOR2 (N1208, N1201, N534);
nor NOR4 (N1209, N1203, N6, N547, N1105);
and AND2 (N1210, N1202, N737);
xor XOR2 (N1211, N1208, N527);
xor XOR2 (N1212, N1205, N1184);
xor XOR2 (N1213, N1204, N659);
nand NAND3 (N1214, N1206, N1188, N592);
nand NAND3 (N1215, N1207, N1051, N735);
nor NOR2 (N1216, N1213, N395);
and AND3 (N1217, N1209, N955, N73);
and AND4 (N1218, N1198, N1147, N644, N568);
buf BUF1 (N1219, N1216);
nor NOR4 (N1220, N1214, N875, N344, N98);
or OR3 (N1221, N1211, N1067, N776);
or OR2 (N1222, N1219, N115);
buf BUF1 (N1223, N1200);
xor XOR2 (N1224, N1222, N846);
xor XOR2 (N1225, N1224, N13);
nor NOR4 (N1226, N1225, N293, N505, N928);
and AND2 (N1227, N1218, N644);
nand NAND3 (N1228, N1212, N631, N1116);
nor NOR4 (N1229, N1220, N1196, N615, N358);
nand NAND2 (N1230, N1228, N550);
nand NAND4 (N1231, N1229, N172, N1188, N347);
and AND2 (N1232, N1183, N1207);
not NOT1 (N1233, N1210);
and AND3 (N1234, N1215, N844, N750);
nor NOR2 (N1235, N1227, N673);
buf BUF1 (N1236, N1230);
xor XOR2 (N1237, N1223, N208);
buf BUF1 (N1238, N1237);
or OR4 (N1239, N1231, N158, N913, N472);
not NOT1 (N1240, N1233);
nand NAND2 (N1241, N1226, N317);
buf BUF1 (N1242, N1235);
and AND3 (N1243, N1241, N987, N1241);
and AND3 (N1244, N1217, N1056, N379);
nand NAND2 (N1245, N1234, N611);
nor NOR2 (N1246, N1244, N702);
xor XOR2 (N1247, N1245, N1067);
buf BUF1 (N1248, N1239);
or OR2 (N1249, N1247, N328);
xor XOR2 (N1250, N1243, N1116);
and AND3 (N1251, N1232, N1086, N703);
buf BUF1 (N1252, N1236);
buf BUF1 (N1253, N1250);
or OR2 (N1254, N1248, N115);
xor XOR2 (N1255, N1251, N1199);
buf BUF1 (N1256, N1254);
not NOT1 (N1257, N1249);
nand NAND2 (N1258, N1240, N1165);
and AND4 (N1259, N1258, N645, N968, N446);
nor NOR4 (N1260, N1255, N809, N474, N464);
nor NOR4 (N1261, N1221, N374, N1248, N426);
nor NOR3 (N1262, N1252, N1084, N229);
nor NOR3 (N1263, N1246, N211, N327);
not NOT1 (N1264, N1262);
nor NOR4 (N1265, N1242, N839, N965, N1114);
xor XOR2 (N1266, N1238, N113);
or OR4 (N1267, N1253, N896, N441, N949);
nand NAND3 (N1268, N1263, N86, N459);
nand NAND3 (N1269, N1259, N154, N436);
and AND3 (N1270, N1265, N867, N896);
nor NOR2 (N1271, N1269, N1026);
or OR3 (N1272, N1266, N1176, N971);
not NOT1 (N1273, N1261);
not NOT1 (N1274, N1272);
not NOT1 (N1275, N1267);
nor NOR2 (N1276, N1257, N137);
not NOT1 (N1277, N1274);
buf BUF1 (N1278, N1277);
buf BUF1 (N1279, N1268);
and AND2 (N1280, N1271, N435);
not NOT1 (N1281, N1256);
buf BUF1 (N1282, N1275);
buf BUF1 (N1283, N1278);
xor XOR2 (N1284, N1264, N1194);
or OR2 (N1285, N1270, N972);
and AND4 (N1286, N1285, N1078, N6, N486);
not NOT1 (N1287, N1284);
nand NAND3 (N1288, N1281, N385, N1207);
or OR2 (N1289, N1288, N361);
xor XOR2 (N1290, N1273, N762);
nand NAND2 (N1291, N1289, N639);
or OR2 (N1292, N1279, N953);
nor NOR3 (N1293, N1292, N166, N1110);
xor XOR2 (N1294, N1293, N472);
nand NAND3 (N1295, N1283, N247, N261);
not NOT1 (N1296, N1287);
or OR4 (N1297, N1291, N919, N1261, N764);
not NOT1 (N1298, N1296);
nor NOR4 (N1299, N1280, N925, N780, N464);
or OR3 (N1300, N1299, N963, N403);
xor XOR2 (N1301, N1286, N975);
xor XOR2 (N1302, N1297, N923);
or OR3 (N1303, N1282, N1195, N739);
and AND2 (N1304, N1276, N438);
or OR4 (N1305, N1304, N154, N657, N287);
buf BUF1 (N1306, N1290);
nand NAND2 (N1307, N1301, N862);
nor NOR4 (N1308, N1260, N659, N125, N1033);
nor NOR2 (N1309, N1305, N234);
or OR2 (N1310, N1307, N1263);
not NOT1 (N1311, N1308);
not NOT1 (N1312, N1295);
buf BUF1 (N1313, N1306);
not NOT1 (N1314, N1309);
not NOT1 (N1315, N1314);
not NOT1 (N1316, N1303);
buf BUF1 (N1317, N1316);
not NOT1 (N1318, N1313);
not NOT1 (N1319, N1302);
xor XOR2 (N1320, N1317, N295);
nand NAND2 (N1321, N1298, N5);
and AND4 (N1322, N1294, N348, N265, N385);
buf BUF1 (N1323, N1322);
xor XOR2 (N1324, N1321, N216);
nand NAND4 (N1325, N1312, N1008, N1197, N1025);
and AND3 (N1326, N1323, N219, N33);
nand NAND4 (N1327, N1300, N64, N1302, N815);
or OR4 (N1328, N1318, N1178, N1120, N396);
buf BUF1 (N1329, N1310);
xor XOR2 (N1330, N1315, N633);
or OR2 (N1331, N1311, N966);
not NOT1 (N1332, N1319);
xor XOR2 (N1333, N1325, N58);
nand NAND3 (N1334, N1324, N1094, N1104);
nor NOR2 (N1335, N1326, N603);
and AND2 (N1336, N1327, N1198);
nor NOR2 (N1337, N1332, N806);
or OR4 (N1338, N1337, N406, N159, N569);
nand NAND2 (N1339, N1333, N403);
nand NAND4 (N1340, N1338, N1012, N521, N1142);
xor XOR2 (N1341, N1330, N418);
and AND3 (N1342, N1336, N104, N1154);
nand NAND4 (N1343, N1340, N1305, N381, N1314);
xor XOR2 (N1344, N1329, N465);
or OR3 (N1345, N1344, N344, N783);
not NOT1 (N1346, N1343);
or OR3 (N1347, N1341, N801, N1229);
and AND2 (N1348, N1334, N455);
nor NOR4 (N1349, N1345, N661, N1153, N515);
nor NOR2 (N1350, N1348, N402);
xor XOR2 (N1351, N1335, N362);
and AND3 (N1352, N1328, N177, N544);
nand NAND3 (N1353, N1350, N382, N1129);
xor XOR2 (N1354, N1346, N238);
nor NOR2 (N1355, N1339, N963);
xor XOR2 (N1356, N1320, N1305);
nor NOR2 (N1357, N1351, N71);
nor NOR4 (N1358, N1357, N1088, N309, N842);
nor NOR2 (N1359, N1342, N514);
or OR3 (N1360, N1352, N783, N738);
nand NAND3 (N1361, N1354, N981, N1241);
nor NOR3 (N1362, N1349, N218, N748);
xor XOR2 (N1363, N1360, N300);
nor NOR3 (N1364, N1363, N413, N137);
buf BUF1 (N1365, N1331);
or OR2 (N1366, N1359, N1310);
nand NAND4 (N1367, N1353, N1090, N1124, N1187);
xor XOR2 (N1368, N1367, N601);
nor NOR4 (N1369, N1361, N74, N1265, N164);
and AND4 (N1370, N1364, N814, N1134, N275);
not NOT1 (N1371, N1369);
xor XOR2 (N1372, N1358, N713);
nor NOR3 (N1373, N1355, N37, N607);
nand NAND3 (N1374, N1371, N985, N83);
and AND2 (N1375, N1370, N289);
and AND3 (N1376, N1372, N1147, N1165);
nor NOR4 (N1377, N1362, N1297, N698, N159);
or OR4 (N1378, N1374, N393, N141, N115);
or OR4 (N1379, N1377, N188, N850, N854);
nand NAND3 (N1380, N1365, N299, N598);
and AND4 (N1381, N1378, N835, N603, N69);
or OR2 (N1382, N1373, N129);
nor NOR3 (N1383, N1375, N1341, N1002);
or OR3 (N1384, N1376, N199, N983);
and AND2 (N1385, N1356, N138);
buf BUF1 (N1386, N1385);
and AND4 (N1387, N1347, N1031, N28, N49);
xor XOR2 (N1388, N1386, N914);
nand NAND3 (N1389, N1387, N531, N1245);
nor NOR2 (N1390, N1368, N727);
and AND2 (N1391, N1379, N1031);
xor XOR2 (N1392, N1381, N1186);
xor XOR2 (N1393, N1392, N42);
nand NAND4 (N1394, N1389, N79, N1189, N401);
not NOT1 (N1395, N1388);
nand NAND4 (N1396, N1390, N942, N541, N500);
not NOT1 (N1397, N1382);
nor NOR2 (N1398, N1391, N949);
nor NOR3 (N1399, N1393, N865, N478);
not NOT1 (N1400, N1380);
buf BUF1 (N1401, N1398);
nor NOR2 (N1402, N1401, N913);
not NOT1 (N1403, N1402);
nor NOR3 (N1404, N1395, N1108, N1059);
nand NAND2 (N1405, N1366, N989);
nand NAND2 (N1406, N1403, N86);
not NOT1 (N1407, N1404);
nor NOR2 (N1408, N1397, N1321);
nor NOR3 (N1409, N1408, N1058, N182);
nand NAND2 (N1410, N1383, N1364);
buf BUF1 (N1411, N1400);
or OR3 (N1412, N1394, N300, N133);
or OR4 (N1413, N1405, N602, N1412, N1201);
buf BUF1 (N1414, N726);
buf BUF1 (N1415, N1384);
not NOT1 (N1416, N1411);
not NOT1 (N1417, N1407);
or OR2 (N1418, N1417, N1374);
or OR4 (N1419, N1413, N870, N170, N467);
and AND3 (N1420, N1419, N1328, N253);
xor XOR2 (N1421, N1416, N1338);
and AND3 (N1422, N1420, N985, N570);
nand NAND3 (N1423, N1418, N444, N254);
nand NAND2 (N1424, N1396, N550);
and AND2 (N1425, N1423, N374);
buf BUF1 (N1426, N1414);
not NOT1 (N1427, N1399);
xor XOR2 (N1428, N1410, N480);
not NOT1 (N1429, N1426);
and AND4 (N1430, N1406, N430, N11, N386);
or OR3 (N1431, N1424, N21, N1174);
and AND3 (N1432, N1415, N554, N689);
not NOT1 (N1433, N1431);
and AND4 (N1434, N1429, N944, N656, N718);
and AND2 (N1435, N1428, N1357);
and AND2 (N1436, N1409, N622);
xor XOR2 (N1437, N1427, N361);
or OR4 (N1438, N1436, N1276, N216, N1406);
buf BUF1 (N1439, N1433);
nor NOR2 (N1440, N1421, N1283);
or OR2 (N1441, N1434, N318);
xor XOR2 (N1442, N1430, N423);
nor NOR4 (N1443, N1435, N1352, N561, N981);
nor NOR3 (N1444, N1442, N181, N1245);
nand NAND4 (N1445, N1437, N1109, N483, N1367);
nor NOR4 (N1446, N1440, N885, N1004, N803);
or OR3 (N1447, N1439, N921, N1021);
and AND3 (N1448, N1443, N551, N4);
nor NOR3 (N1449, N1445, N648, N1244);
and AND3 (N1450, N1438, N429, N960);
not NOT1 (N1451, N1446);
not NOT1 (N1452, N1448);
and AND2 (N1453, N1450, N1238);
and AND4 (N1454, N1452, N111, N128, N223);
nand NAND2 (N1455, N1454, N209);
and AND3 (N1456, N1425, N349, N678);
and AND4 (N1457, N1444, N725, N595, N1041);
not NOT1 (N1458, N1422);
buf BUF1 (N1459, N1458);
nor NOR3 (N1460, N1457, N1387, N1055);
nand NAND3 (N1461, N1449, N423, N886);
or OR3 (N1462, N1441, N533, N230);
nand NAND2 (N1463, N1456, N1436);
nor NOR3 (N1464, N1455, N696, N1373);
nand NAND2 (N1465, N1459, N906);
xor XOR2 (N1466, N1461, N1074);
nor NOR4 (N1467, N1465, N162, N55, N1397);
and AND3 (N1468, N1467, N1466, N1193);
xor XOR2 (N1469, N1291, N923);
not NOT1 (N1470, N1469);
and AND4 (N1471, N1447, N1004, N126, N181);
and AND3 (N1472, N1471, N574, N864);
or OR4 (N1473, N1451, N135, N1144, N1283);
and AND2 (N1474, N1473, N698);
not NOT1 (N1475, N1463);
or OR3 (N1476, N1432, N92, N1193);
and AND3 (N1477, N1468, N522, N1264);
not NOT1 (N1478, N1472);
buf BUF1 (N1479, N1464);
nand NAND2 (N1480, N1453, N1133);
or OR2 (N1481, N1460, N1023);
or OR3 (N1482, N1462, N1165, N474);
and AND3 (N1483, N1474, N1057, N910);
or OR3 (N1484, N1475, N1103, N204);
xor XOR2 (N1485, N1470, N237);
xor XOR2 (N1486, N1482, N651);
nor NOR2 (N1487, N1477, N893);
or OR2 (N1488, N1484, N875);
buf BUF1 (N1489, N1485);
nor NOR2 (N1490, N1486, N1389);
buf BUF1 (N1491, N1490);
xor XOR2 (N1492, N1478, N630);
xor XOR2 (N1493, N1487, N653);
not NOT1 (N1494, N1481);
or OR4 (N1495, N1488, N1155, N427, N1052);
not NOT1 (N1496, N1489);
nand NAND3 (N1497, N1476, N1178, N997);
xor XOR2 (N1498, N1493, N1257);
not NOT1 (N1499, N1498);
not NOT1 (N1500, N1491);
xor XOR2 (N1501, N1480, N1441);
xor XOR2 (N1502, N1496, N1336);
or OR4 (N1503, N1500, N805, N644, N950);
not NOT1 (N1504, N1503);
nand NAND4 (N1505, N1483, N211, N217, N1305);
nor NOR4 (N1506, N1505, N1317, N126, N880);
or OR2 (N1507, N1492, N1289);
nor NOR2 (N1508, N1497, N278);
or OR4 (N1509, N1508, N445, N1084, N1036);
not NOT1 (N1510, N1502);
buf BUF1 (N1511, N1510);
nor NOR3 (N1512, N1494, N224, N199);
and AND3 (N1513, N1512, N770, N1098);
nand NAND3 (N1514, N1506, N1356, N1142);
xor XOR2 (N1515, N1501, N380);
buf BUF1 (N1516, N1479);
and AND4 (N1517, N1514, N1394, N282, N1273);
nand NAND3 (N1518, N1515, N48, N763);
or OR2 (N1519, N1495, N257);
and AND4 (N1520, N1517, N1127, N74, N1035);
nand NAND4 (N1521, N1513, N336, N713, N75);
buf BUF1 (N1522, N1521);
nor NOR4 (N1523, N1509, N113, N10, N748);
endmodule