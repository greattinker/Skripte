// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N511,N514,N512,N513,N495,N508,N515,N503,N506,N516;

and AND4 (N17, N6, N9, N14, N3);
nor NOR3 (N18, N4, N8, N9);
nor NOR4 (N19, N15, N7, N18, N1);
nor NOR4 (N20, N12, N9, N19, N2);
xor XOR2 (N21, N9, N14);
not NOT1 (N22, N12);
xor XOR2 (N23, N15, N1);
and AND4 (N24, N11, N17, N9, N11);
or OR2 (N25, N8, N19);
and AND3 (N26, N12, N4, N24);
nand NAND2 (N27, N6, N13);
not NOT1 (N28, N24);
not NOT1 (N29, N5);
or OR4 (N30, N26, N24, N19, N3);
not NOT1 (N31, N3);
buf BUF1 (N32, N21);
or OR3 (N33, N29, N16, N21);
nor NOR2 (N34, N31, N27);
nor NOR2 (N35, N11, N8);
nor NOR4 (N36, N30, N35, N5, N19);
and AND2 (N37, N32, N17);
xor XOR2 (N38, N13, N12);
nor NOR2 (N39, N22, N24);
nor NOR3 (N40, N38, N12, N24);
and AND3 (N41, N34, N34, N30);
nand NAND3 (N42, N20, N15, N7);
and AND3 (N43, N37, N33, N16);
nand NAND3 (N44, N27, N5, N5);
buf BUF1 (N45, N28);
xor XOR2 (N46, N40, N8);
not NOT1 (N47, N36);
or OR4 (N48, N47, N38, N31, N20);
nand NAND3 (N49, N44, N44, N15);
nand NAND2 (N50, N41, N8);
xor XOR2 (N51, N42, N26);
buf BUF1 (N52, N48);
not NOT1 (N53, N25);
nand NAND2 (N54, N53, N3);
buf BUF1 (N55, N52);
nor NOR3 (N56, N39, N28, N53);
xor XOR2 (N57, N51, N3);
or OR4 (N58, N54, N33, N38, N8);
or OR2 (N59, N46, N35);
nor NOR4 (N60, N59, N21, N6, N17);
and AND3 (N61, N49, N6, N41);
and AND3 (N62, N50, N34, N21);
not NOT1 (N63, N45);
nor NOR3 (N64, N23, N8, N51);
nand NAND4 (N65, N61, N50, N59, N9);
nor NOR3 (N66, N65, N64, N4);
and AND3 (N67, N22, N54, N10);
nor NOR3 (N68, N62, N67, N60);
nor NOR3 (N69, N48, N57, N7);
not NOT1 (N70, N51);
nand NAND4 (N71, N20, N28, N36, N27);
nand NAND2 (N72, N66, N18);
and AND3 (N73, N71, N58, N36);
not NOT1 (N74, N6);
xor XOR2 (N75, N68, N40);
or OR2 (N76, N63, N37);
or OR2 (N77, N75, N66);
buf BUF1 (N78, N74);
nor NOR2 (N79, N70, N18);
buf BUF1 (N80, N55);
nand NAND3 (N81, N69, N43, N22);
xor XOR2 (N82, N23, N32);
not NOT1 (N83, N79);
buf BUF1 (N84, N72);
not NOT1 (N85, N76);
or OR3 (N86, N81, N13, N72);
or OR4 (N87, N80, N11, N30, N77);
buf BUF1 (N88, N30);
buf BUF1 (N89, N86);
not NOT1 (N90, N82);
or OR2 (N91, N89, N80);
xor XOR2 (N92, N85, N49);
xor XOR2 (N93, N87, N80);
buf BUF1 (N94, N73);
and AND2 (N95, N91, N63);
or OR3 (N96, N83, N16, N52);
nor NOR3 (N97, N90, N83, N25);
buf BUF1 (N98, N93);
buf BUF1 (N99, N97);
xor XOR2 (N100, N56, N70);
buf BUF1 (N101, N95);
nand NAND2 (N102, N88, N70);
xor XOR2 (N103, N78, N58);
and AND3 (N104, N101, N96, N103);
buf BUF1 (N105, N95);
not NOT1 (N106, N64);
buf BUF1 (N107, N105);
buf BUF1 (N108, N98);
nor NOR4 (N109, N100, N46, N48, N76);
not NOT1 (N110, N92);
buf BUF1 (N111, N108);
or OR4 (N112, N110, N35, N7, N2);
and AND4 (N113, N112, N92, N58, N85);
or OR2 (N114, N84, N55);
nand NAND2 (N115, N99, N41);
xor XOR2 (N116, N107, N32);
buf BUF1 (N117, N106);
and AND3 (N118, N102, N105, N84);
and AND2 (N119, N117, N35);
and AND2 (N120, N113, N93);
and AND4 (N121, N111, N48, N20, N85);
buf BUF1 (N122, N109);
and AND2 (N123, N116, N29);
nor NOR4 (N124, N114, N76, N88, N89);
and AND2 (N125, N119, N59);
buf BUF1 (N126, N124);
not NOT1 (N127, N122);
xor XOR2 (N128, N126, N84);
xor XOR2 (N129, N121, N18);
or OR3 (N130, N104, N59, N78);
nand NAND4 (N131, N118, N27, N5, N55);
nand NAND3 (N132, N130, N16, N50);
xor XOR2 (N133, N128, N74);
not NOT1 (N134, N133);
xor XOR2 (N135, N115, N68);
and AND3 (N136, N125, N63, N21);
nor NOR3 (N137, N120, N104, N90);
nor NOR4 (N138, N131, N117, N127, N123);
nor NOR4 (N139, N38, N42, N30, N73);
buf BUF1 (N140, N68);
or OR2 (N141, N134, N128);
xor XOR2 (N142, N135, N26);
or OR3 (N143, N129, N57, N48);
and AND2 (N144, N143, N70);
nor NOR4 (N145, N138, N54, N24, N134);
and AND3 (N146, N140, N67, N121);
not NOT1 (N147, N144);
xor XOR2 (N148, N142, N135);
nor NOR3 (N149, N137, N119, N69);
and AND3 (N150, N147, N41, N102);
or OR3 (N151, N94, N89, N149);
nand NAND4 (N152, N126, N64, N105, N146);
nor NOR3 (N153, N104, N98, N66);
or OR2 (N154, N153, N139);
xor XOR2 (N155, N81, N45);
xor XOR2 (N156, N155, N85);
or OR2 (N157, N132, N38);
buf BUF1 (N158, N151);
or OR4 (N159, N152, N107, N93, N81);
or OR2 (N160, N154, N86);
or OR4 (N161, N148, N69, N1, N138);
xor XOR2 (N162, N157, N124);
buf BUF1 (N163, N161);
nor NOR2 (N164, N141, N18);
and AND2 (N165, N150, N150);
xor XOR2 (N166, N156, N53);
buf BUF1 (N167, N165);
buf BUF1 (N168, N163);
nor NOR4 (N169, N136, N114, N50, N62);
xor XOR2 (N170, N169, N31);
buf BUF1 (N171, N166);
buf BUF1 (N172, N168);
buf BUF1 (N173, N170);
nor NOR4 (N174, N173, N44, N143, N122);
xor XOR2 (N175, N162, N65);
or OR3 (N176, N174, N33, N110);
not NOT1 (N177, N145);
not NOT1 (N178, N158);
nand NAND2 (N179, N171, N43);
xor XOR2 (N180, N177, N76);
and AND3 (N181, N175, N171, N160);
not NOT1 (N182, N177);
nand NAND2 (N183, N167, N27);
buf BUF1 (N184, N181);
or OR3 (N185, N184, N57, N78);
or OR3 (N186, N176, N88, N150);
nand NAND2 (N187, N179, N89);
not NOT1 (N188, N186);
and AND4 (N189, N183, N21, N180, N126);
xor XOR2 (N190, N186, N21);
and AND3 (N191, N159, N116, N118);
or OR3 (N192, N172, N63, N151);
and AND3 (N193, N178, N120, N118);
not NOT1 (N194, N191);
not NOT1 (N195, N190);
or OR3 (N196, N193, N47, N44);
buf BUF1 (N197, N182);
xor XOR2 (N198, N195, N42);
and AND3 (N199, N196, N169, N179);
or OR4 (N200, N198, N74, N166, N103);
or OR2 (N201, N199, N54);
xor XOR2 (N202, N164, N124);
or OR4 (N203, N189, N144, N201, N93);
xor XOR2 (N204, N69, N145);
buf BUF1 (N205, N204);
buf BUF1 (N206, N185);
buf BUF1 (N207, N200);
xor XOR2 (N208, N187, N10);
buf BUF1 (N209, N202);
buf BUF1 (N210, N207);
or OR4 (N211, N203, N199, N172, N55);
not NOT1 (N212, N188);
nand NAND2 (N213, N212, N140);
nor NOR4 (N214, N206, N127, N104, N179);
and AND4 (N215, N197, N37, N26, N25);
not NOT1 (N216, N194);
buf BUF1 (N217, N208);
or OR2 (N218, N215, N42);
buf BUF1 (N219, N218);
xor XOR2 (N220, N192, N65);
buf BUF1 (N221, N217);
buf BUF1 (N222, N220);
buf BUF1 (N223, N210);
nand NAND3 (N224, N205, N62, N158);
nor NOR4 (N225, N216, N214, N93, N96);
nand NAND3 (N226, N77, N12, N82);
xor XOR2 (N227, N226, N165);
buf BUF1 (N228, N227);
nor NOR4 (N229, N224, N73, N129, N221);
nor NOR4 (N230, N184, N145, N21, N134);
and AND3 (N231, N225, N1, N26);
buf BUF1 (N232, N211);
buf BUF1 (N233, N230);
xor XOR2 (N234, N209, N130);
xor XOR2 (N235, N234, N116);
nor NOR2 (N236, N229, N158);
nor NOR2 (N237, N213, N176);
not NOT1 (N238, N228);
nor NOR3 (N239, N237, N142, N220);
nand NAND2 (N240, N236, N125);
buf BUF1 (N241, N222);
or OR2 (N242, N233, N200);
nor NOR4 (N243, N242, N135, N95, N233);
and AND4 (N244, N243, N243, N221, N188);
nor NOR4 (N245, N238, N176, N202, N20);
not NOT1 (N246, N223);
or OR2 (N247, N241, N209);
xor XOR2 (N248, N247, N123);
nor NOR3 (N249, N219, N22, N6);
nor NOR4 (N250, N231, N28, N178, N158);
and AND3 (N251, N239, N102, N154);
xor XOR2 (N252, N244, N176);
not NOT1 (N253, N246);
buf BUF1 (N254, N252);
and AND4 (N255, N248, N242, N15, N97);
not NOT1 (N256, N253);
buf BUF1 (N257, N250);
buf BUF1 (N258, N235);
not NOT1 (N259, N254);
buf BUF1 (N260, N259);
not NOT1 (N261, N256);
nor NOR3 (N262, N251, N121, N44);
buf BUF1 (N263, N261);
or OR4 (N264, N263, N53, N168, N142);
not NOT1 (N265, N245);
xor XOR2 (N266, N232, N100);
nand NAND2 (N267, N255, N262);
nand NAND2 (N268, N119, N227);
or OR4 (N269, N260, N87, N240, N140);
or OR4 (N270, N9, N256, N74, N126);
buf BUF1 (N271, N267);
buf BUF1 (N272, N264);
nor NOR4 (N273, N257, N64, N183, N193);
or OR3 (N274, N273, N186, N217);
buf BUF1 (N275, N265);
xor XOR2 (N276, N272, N215);
nor NOR4 (N277, N270, N119, N127, N37);
and AND3 (N278, N276, N34, N137);
not NOT1 (N279, N269);
nand NAND3 (N280, N268, N177, N246);
xor XOR2 (N281, N280, N64);
nand NAND4 (N282, N278, N248, N71, N55);
xor XOR2 (N283, N281, N5);
nand NAND3 (N284, N277, N261, N44);
xor XOR2 (N285, N284, N8);
buf BUF1 (N286, N258);
and AND4 (N287, N274, N57, N225, N215);
xor XOR2 (N288, N249, N102);
nor NOR4 (N289, N275, N107, N43, N79);
or OR3 (N290, N287, N69, N45);
xor XOR2 (N291, N266, N216);
nor NOR2 (N292, N286, N274);
not NOT1 (N293, N279);
xor XOR2 (N294, N285, N181);
not NOT1 (N295, N292);
nor NOR3 (N296, N290, N64, N212);
nor NOR3 (N297, N271, N244, N237);
and AND3 (N298, N291, N108, N105);
or OR2 (N299, N297, N171);
and AND4 (N300, N299, N284, N25, N191);
not NOT1 (N301, N289);
or OR4 (N302, N295, N299, N152, N301);
or OR2 (N303, N107, N160);
not NOT1 (N304, N298);
or OR3 (N305, N293, N10, N29);
or OR3 (N306, N305, N139, N170);
nand NAND2 (N307, N283, N285);
buf BUF1 (N308, N304);
xor XOR2 (N309, N307, N202);
buf BUF1 (N310, N300);
not NOT1 (N311, N282);
not NOT1 (N312, N294);
and AND2 (N313, N302, N17);
xor XOR2 (N314, N303, N83);
not NOT1 (N315, N296);
buf BUF1 (N316, N288);
and AND4 (N317, N312, N187, N210, N215);
not NOT1 (N318, N315);
xor XOR2 (N319, N308, N50);
or OR4 (N320, N310, N63, N236, N309);
nor NOR3 (N321, N194, N133, N79);
nor NOR3 (N322, N321, N267, N108);
nor NOR2 (N323, N306, N132);
xor XOR2 (N324, N318, N252);
or OR4 (N325, N316, N77, N223, N48);
not NOT1 (N326, N322);
buf BUF1 (N327, N325);
or OR2 (N328, N327, N198);
not NOT1 (N329, N326);
not NOT1 (N330, N329);
and AND3 (N331, N314, N167, N275);
nand NAND4 (N332, N320, N306, N155, N24);
not NOT1 (N333, N317);
xor XOR2 (N334, N330, N260);
nand NAND3 (N335, N323, N12, N165);
or OR2 (N336, N328, N222);
not NOT1 (N337, N336);
or OR4 (N338, N333, N57, N110, N145);
nor NOR3 (N339, N332, N6, N18);
and AND4 (N340, N334, N230, N14, N65);
and AND3 (N341, N331, N18, N56);
nor NOR2 (N342, N313, N55);
buf BUF1 (N343, N342);
or OR3 (N344, N340, N157, N195);
xor XOR2 (N345, N311, N240);
xor XOR2 (N346, N337, N270);
or OR3 (N347, N324, N196, N271);
xor XOR2 (N348, N338, N57);
nand NAND3 (N349, N348, N34, N58);
nor NOR3 (N350, N335, N193, N178);
xor XOR2 (N351, N343, N271);
buf BUF1 (N352, N349);
nor NOR3 (N353, N344, N77, N223);
or OR3 (N354, N350, N171, N346);
xor XOR2 (N355, N131, N61);
and AND3 (N356, N345, N216, N228);
xor XOR2 (N357, N351, N184);
nand NAND4 (N358, N356, N72, N170, N201);
and AND3 (N359, N341, N245, N210);
and AND3 (N360, N354, N249, N353);
nand NAND4 (N361, N354, N195, N140, N216);
xor XOR2 (N362, N319, N274);
or OR4 (N363, N347, N163, N13, N277);
or OR4 (N364, N360, N173, N124, N225);
buf BUF1 (N365, N358);
not NOT1 (N366, N361);
nand NAND2 (N367, N363, N238);
nor NOR2 (N368, N367, N218);
xor XOR2 (N369, N352, N217);
or OR3 (N370, N369, N80, N92);
nand NAND4 (N371, N339, N123, N11, N142);
or OR4 (N372, N355, N281, N365, N32);
buf BUF1 (N373, N333);
xor XOR2 (N374, N370, N21);
and AND2 (N375, N362, N75);
nand NAND4 (N376, N368, N255, N216, N267);
not NOT1 (N377, N366);
xor XOR2 (N378, N364, N306);
nand NAND4 (N379, N377, N105, N9, N266);
or OR2 (N380, N374, N226);
or OR3 (N381, N371, N272, N4);
nor NOR2 (N382, N373, N314);
xor XOR2 (N383, N372, N278);
or OR3 (N384, N379, N61, N209);
xor XOR2 (N385, N375, N233);
buf BUF1 (N386, N384);
nor NOR3 (N387, N383, N56, N106);
and AND2 (N388, N381, N300);
or OR2 (N389, N380, N115);
nor NOR3 (N390, N389, N166, N177);
and AND2 (N391, N378, N197);
buf BUF1 (N392, N390);
nand NAND3 (N393, N388, N328, N148);
and AND4 (N394, N359, N210, N363, N91);
buf BUF1 (N395, N393);
nor NOR3 (N396, N392, N94, N193);
and AND3 (N397, N357, N45, N204);
nor NOR2 (N398, N391, N198);
buf BUF1 (N399, N394);
and AND3 (N400, N397, N180, N349);
not NOT1 (N401, N398);
or OR3 (N402, N382, N376, N117);
buf BUF1 (N403, N174);
nor NOR3 (N404, N400, N229, N335);
buf BUF1 (N405, N399);
or OR4 (N406, N404, N368, N147, N45);
nand NAND4 (N407, N405, N61, N319, N137);
nor NOR2 (N408, N387, N239);
buf BUF1 (N409, N402);
xor XOR2 (N410, N406, N51);
not NOT1 (N411, N403);
xor XOR2 (N412, N401, N133);
buf BUF1 (N413, N411);
xor XOR2 (N414, N395, N34);
xor XOR2 (N415, N409, N180);
nand NAND2 (N416, N386, N85);
xor XOR2 (N417, N396, N1);
nand NAND3 (N418, N385, N290, N234);
nor NOR4 (N419, N418, N65, N33, N196);
nand NAND2 (N420, N413, N194);
nand NAND4 (N421, N408, N56, N3, N246);
not NOT1 (N422, N412);
and AND4 (N423, N414, N62, N359, N197);
nand NAND2 (N424, N423, N80);
and AND2 (N425, N419, N190);
buf BUF1 (N426, N410);
nand NAND3 (N427, N421, N299, N345);
nor NOR3 (N428, N416, N235, N47);
buf BUF1 (N429, N424);
nand NAND2 (N430, N420, N199);
not NOT1 (N431, N415);
and AND3 (N432, N427, N237, N81);
nand NAND4 (N433, N429, N339, N140, N121);
or OR2 (N434, N433, N358);
or OR4 (N435, N426, N274, N100, N211);
or OR3 (N436, N434, N181, N207);
or OR2 (N437, N425, N192);
not NOT1 (N438, N437);
and AND2 (N439, N431, N176);
xor XOR2 (N440, N428, N258);
not NOT1 (N441, N440);
nor NOR2 (N442, N439, N19);
xor XOR2 (N443, N407, N47);
not NOT1 (N444, N430);
buf BUF1 (N445, N442);
xor XOR2 (N446, N445, N32);
nor NOR2 (N447, N432, N62);
xor XOR2 (N448, N447, N371);
and AND2 (N449, N438, N123);
xor XOR2 (N450, N448, N4);
and AND4 (N451, N450, N213, N18, N170);
buf BUF1 (N452, N451);
xor XOR2 (N453, N441, N141);
xor XOR2 (N454, N449, N354);
and AND3 (N455, N443, N358, N74);
and AND2 (N456, N446, N277);
buf BUF1 (N457, N444);
not NOT1 (N458, N452);
xor XOR2 (N459, N417, N295);
or OR2 (N460, N457, N248);
nor NOR3 (N461, N454, N22, N203);
not NOT1 (N462, N459);
nand NAND2 (N463, N455, N46);
xor XOR2 (N464, N456, N181);
buf BUF1 (N465, N461);
and AND3 (N466, N460, N59, N255);
xor XOR2 (N467, N466, N365);
and AND2 (N468, N453, N424);
nand NAND2 (N469, N463, N462);
and AND2 (N470, N357, N16);
nand NAND2 (N471, N469, N40);
nor NOR2 (N472, N471, N127);
xor XOR2 (N473, N464, N87);
nor NOR2 (N474, N435, N32);
and AND2 (N475, N473, N374);
or OR4 (N476, N475, N63, N369, N469);
or OR3 (N477, N422, N218, N421);
xor XOR2 (N478, N470, N474);
not NOT1 (N479, N262);
and AND2 (N480, N479, N90);
or OR3 (N481, N477, N5, N180);
and AND2 (N482, N472, N282);
or OR4 (N483, N467, N277, N193, N219);
nor NOR4 (N484, N468, N449, N140, N407);
not NOT1 (N485, N482);
nand NAND3 (N486, N478, N456, N469);
xor XOR2 (N487, N486, N194);
buf BUF1 (N488, N487);
xor XOR2 (N489, N480, N389);
nand NAND3 (N490, N484, N18, N106);
nor NOR2 (N491, N465, N373);
not NOT1 (N492, N483);
nor NOR2 (N493, N485, N309);
or OR2 (N494, N489, N121);
buf BUF1 (N495, N492);
buf BUF1 (N496, N491);
not NOT1 (N497, N488);
not NOT1 (N498, N497);
or OR2 (N499, N476, N474);
not NOT1 (N500, N499);
or OR4 (N501, N458, N72, N156, N295);
and AND3 (N502, N500, N479, N38);
nand NAND3 (N503, N498, N391, N216);
or OR4 (N504, N436, N349, N496, N352);
not NOT1 (N505, N2);
xor XOR2 (N506, N501, N465);
xor XOR2 (N507, N502, N336);
nand NAND3 (N508, N481, N121, N339);
nand NAND2 (N509, N493, N390);
or OR3 (N510, N504, N163, N439);
nor NOR2 (N511, N509, N118);
and AND3 (N512, N490, N492, N312);
or OR4 (N513, N494, N318, N510, N180);
nor NOR2 (N514, N163, N428);
nand NAND3 (N515, N505, N119, N43);
or OR3 (N516, N507, N231, N421);
endmodule