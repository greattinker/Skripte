// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N118,N113,N98,N122,N111,N117,N120,N115,N114,N123;

nand NAND4 (N24, N6, N3, N1, N16);
nor NOR3 (N25, N14, N20, N1);
or OR2 (N26, N18, N25);
xor XOR2 (N27, N8, N23);
not NOT1 (N28, N22);
not NOT1 (N29, N26);
not NOT1 (N30, N19);
not NOT1 (N31, N29);
and AND2 (N32, N30, N13);
nor NOR3 (N33, N24, N20, N22);
nand NAND2 (N34, N17, N16);
buf BUF1 (N35, N34);
or OR4 (N36, N34, N25, N27, N14);
not NOT1 (N37, N8);
nor NOR4 (N38, N11, N33, N22, N15);
nand NAND3 (N39, N28, N25, N21);
or OR4 (N40, N6, N15, N17, N5);
nand NAND3 (N41, N38, N40, N35);
not NOT1 (N42, N12);
nand NAND4 (N43, N26, N22, N24, N41);
buf BUF1 (N44, N32);
and AND3 (N45, N4, N21, N8);
or OR4 (N46, N3, N17, N9, N40);
and AND2 (N47, N37, N7);
xor XOR2 (N48, N14, N34);
buf BUF1 (N49, N47);
buf BUF1 (N50, N36);
nor NOR2 (N51, N49, N47);
and AND3 (N52, N46, N33, N31);
xor XOR2 (N53, N16, N20);
nand NAND4 (N54, N53, N5, N19, N53);
buf BUF1 (N55, N50);
buf BUF1 (N56, N44);
and AND2 (N57, N45, N37);
not NOT1 (N58, N48);
not NOT1 (N59, N51);
not NOT1 (N60, N39);
xor XOR2 (N61, N57, N48);
nand NAND4 (N62, N61, N21, N28, N26);
and AND4 (N63, N43, N57, N53, N13);
or OR2 (N64, N55, N62);
buf BUF1 (N65, N26);
and AND4 (N66, N54, N58, N13, N29);
not NOT1 (N67, N13);
nand NAND3 (N68, N64, N60, N61);
not NOT1 (N69, N52);
and AND4 (N70, N36, N39, N10, N10);
or OR4 (N71, N42, N11, N28, N37);
buf BUF1 (N72, N69);
and AND3 (N73, N70, N13, N68);
and AND2 (N74, N35, N52);
nand NAND2 (N75, N66, N38);
nor NOR3 (N76, N63, N25, N12);
not NOT1 (N77, N75);
nor NOR2 (N78, N72, N19);
nor NOR4 (N79, N56, N43, N15, N14);
or OR2 (N80, N67, N33);
xor XOR2 (N81, N71, N3);
not NOT1 (N82, N80);
not NOT1 (N83, N79);
and AND3 (N84, N81, N46, N37);
buf BUF1 (N85, N73);
buf BUF1 (N86, N59);
or OR3 (N87, N84, N57, N86);
nor NOR2 (N88, N45, N11);
not NOT1 (N89, N85);
or OR4 (N90, N77, N31, N78, N80);
buf BUF1 (N91, N37);
and AND2 (N92, N89, N52);
buf BUF1 (N93, N91);
nor NOR3 (N94, N88, N53, N35);
buf BUF1 (N95, N93);
xor XOR2 (N96, N95, N85);
nand NAND2 (N97, N74, N6);
not NOT1 (N98, N83);
xor XOR2 (N99, N82, N64);
xor XOR2 (N100, N94, N1);
and AND3 (N101, N97, N68, N26);
xor XOR2 (N102, N76, N88);
nor NOR3 (N103, N101, N30, N9);
buf BUF1 (N104, N65);
not NOT1 (N105, N87);
or OR4 (N106, N90, N61, N81, N21);
and AND2 (N107, N105, N94);
and AND2 (N108, N106, N56);
buf BUF1 (N109, N103);
or OR2 (N110, N102, N69);
xor XOR2 (N111, N96, N10);
nor NOR3 (N112, N92, N58, N105);
nand NAND3 (N113, N104, N89, N112);
nor NOR2 (N114, N65, N100);
and AND2 (N115, N79, N57);
not NOT1 (N116, N109);
xor XOR2 (N117, N107, N30);
nor NOR4 (N118, N99, N29, N99, N94);
not NOT1 (N119, N110);
and AND2 (N120, N119, N54);
nor NOR3 (N121, N108, N96, N103);
xor XOR2 (N122, N116, N96);
nor NOR4 (N123, N121, N46, N59, N13);
endmodule