// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N805,N815,N811,N797,N820,N801,N817,N814,N816,N821;

or OR3 (N22, N9, N9, N17);
not NOT1 (N23, N7);
and AND3 (N24, N22, N8, N23);
buf BUF1 (N25, N21);
xor XOR2 (N26, N18, N1);
or OR2 (N27, N20, N19);
nand NAND2 (N28, N16, N4);
or OR3 (N29, N7, N9, N13);
xor XOR2 (N30, N29, N10);
not NOT1 (N31, N11);
and AND4 (N32, N23, N18, N24, N29);
and AND3 (N33, N28, N14, N1);
xor XOR2 (N34, N15, N27);
not NOT1 (N35, N20);
xor XOR2 (N36, N30, N15);
nand NAND4 (N37, N6, N31, N33, N32);
buf BUF1 (N38, N27);
nand NAND2 (N39, N35, N20);
or OR2 (N40, N36, N21);
not NOT1 (N41, N16);
and AND3 (N42, N33, N41, N24);
or OR3 (N43, N25, N11, N35);
xor XOR2 (N44, N30, N38);
nor NOR4 (N45, N19, N29, N5, N43);
nand NAND3 (N46, N14, N25, N29);
nor NOR3 (N47, N1, N26, N40);
nand NAND2 (N48, N15, N39);
not NOT1 (N49, N27);
and AND4 (N50, N20, N47, N6, N16);
not NOT1 (N51, N33);
not NOT1 (N52, N45);
nand NAND4 (N53, N37, N41, N39, N31);
xor XOR2 (N54, N51, N49);
not NOT1 (N55, N11);
buf BUF1 (N56, N42);
xor XOR2 (N57, N48, N44);
and AND2 (N58, N20, N11);
and AND2 (N59, N50, N11);
not NOT1 (N60, N52);
nand NAND4 (N61, N60, N25, N6, N20);
nor NOR2 (N62, N46, N38);
or OR4 (N63, N56, N43, N21, N7);
and AND3 (N64, N61, N31, N41);
buf BUF1 (N65, N62);
not NOT1 (N66, N54);
buf BUF1 (N67, N55);
xor XOR2 (N68, N34, N38);
or OR3 (N69, N65, N8, N8);
and AND4 (N70, N57, N36, N16, N69);
nand NAND3 (N71, N48, N67, N2);
nand NAND4 (N72, N37, N45, N60, N64);
buf BUF1 (N73, N27);
buf BUF1 (N74, N58);
nand NAND2 (N75, N74, N54);
and AND3 (N76, N53, N39, N54);
buf BUF1 (N77, N72);
buf BUF1 (N78, N66);
or OR4 (N79, N77, N77, N21, N77);
xor XOR2 (N80, N59, N24);
nor NOR2 (N81, N79, N58);
not NOT1 (N82, N78);
not NOT1 (N83, N70);
buf BUF1 (N84, N71);
not NOT1 (N85, N82);
and AND3 (N86, N81, N82, N84);
not NOT1 (N87, N36);
nor NOR2 (N88, N75, N22);
xor XOR2 (N89, N76, N30);
nor NOR2 (N90, N87, N34);
or OR3 (N91, N86, N13, N41);
and AND3 (N92, N89, N51, N54);
buf BUF1 (N93, N85);
buf BUF1 (N94, N73);
not NOT1 (N95, N92);
nand NAND3 (N96, N63, N43, N74);
and AND4 (N97, N95, N50, N58, N19);
nand NAND2 (N98, N91, N32);
buf BUF1 (N99, N68);
and AND4 (N100, N90, N67, N34, N12);
not NOT1 (N101, N93);
or OR2 (N102, N96, N18);
nor NOR2 (N103, N88, N62);
nand NAND3 (N104, N98, N75, N2);
nand NAND2 (N105, N94, N21);
or OR3 (N106, N83, N49, N59);
or OR2 (N107, N106, N98);
nand NAND3 (N108, N101, N6, N59);
buf BUF1 (N109, N80);
nand NAND4 (N110, N100, N24, N97, N73);
xor XOR2 (N111, N68, N64);
buf BUF1 (N112, N108);
nor NOR3 (N113, N107, N107, N62);
nor NOR3 (N114, N102, N22, N49);
not NOT1 (N115, N114);
nand NAND2 (N116, N99, N49);
buf BUF1 (N117, N110);
not NOT1 (N118, N103);
nand NAND3 (N119, N118, N100, N83);
not NOT1 (N120, N113);
or OR2 (N121, N119, N80);
nand NAND2 (N122, N109, N74);
nor NOR3 (N123, N117, N26, N38);
nand NAND3 (N124, N122, N61, N108);
nor NOR4 (N125, N104, N100, N6, N109);
buf BUF1 (N126, N121);
and AND4 (N127, N111, N118, N76, N125);
nand NAND3 (N128, N51, N37, N49);
or OR4 (N129, N123, N92, N9, N126);
buf BUF1 (N130, N24);
not NOT1 (N131, N116);
nand NAND3 (N132, N128, N67, N93);
nand NAND3 (N133, N129, N52, N70);
and AND2 (N134, N127, N23);
not NOT1 (N135, N132);
or OR3 (N136, N131, N68, N126);
xor XOR2 (N137, N112, N57);
not NOT1 (N138, N124);
and AND4 (N139, N134, N14, N83, N10);
nand NAND2 (N140, N130, N97);
buf BUF1 (N141, N133);
and AND2 (N142, N140, N34);
or OR2 (N143, N136, N100);
xor XOR2 (N144, N142, N34);
nand NAND3 (N145, N138, N57, N120);
xor XOR2 (N146, N73, N58);
nand NAND2 (N147, N145, N9);
and AND3 (N148, N137, N125, N43);
not NOT1 (N149, N141);
nand NAND2 (N150, N146, N149);
xor XOR2 (N151, N115, N60);
or OR2 (N152, N40, N62);
or OR3 (N153, N135, N113, N2);
nand NAND2 (N154, N144, N150);
nor NOR2 (N155, N36, N9);
nand NAND2 (N156, N153, N105);
nor NOR2 (N157, N109, N17);
xor XOR2 (N158, N157, N21);
nand NAND4 (N159, N155, N56, N45, N139);
or OR2 (N160, N147, N97);
not NOT1 (N161, N20);
xor XOR2 (N162, N160, N112);
nor NOR4 (N163, N161, N86, N116, N1);
not NOT1 (N164, N151);
and AND4 (N165, N159, N148, N117, N110);
not NOT1 (N166, N39);
buf BUF1 (N167, N154);
or OR4 (N168, N162, N160, N126, N4);
and AND3 (N169, N163, N75, N2);
xor XOR2 (N170, N167, N18);
nand NAND2 (N171, N164, N25);
nor NOR3 (N172, N168, N136, N159);
nor NOR2 (N173, N165, N168);
and AND4 (N174, N158, N166, N134, N49);
or OR4 (N175, N57, N44, N49, N157);
and AND3 (N176, N170, N150, N5);
buf BUF1 (N177, N152);
nor NOR4 (N178, N174, N5, N163, N85);
not NOT1 (N179, N171);
nor NOR2 (N180, N169, N146);
buf BUF1 (N181, N156);
nand NAND2 (N182, N176, N35);
nor NOR4 (N183, N173, N32, N109, N35);
and AND3 (N184, N179, N16, N45);
xor XOR2 (N185, N177, N146);
nor NOR3 (N186, N185, N185, N19);
or OR4 (N187, N181, N34, N50, N58);
and AND2 (N188, N187, N96);
nor NOR4 (N189, N178, N65, N182, N20);
and AND2 (N190, N115, N80);
or OR3 (N191, N175, N89, N126);
nor NOR3 (N192, N183, N40, N107);
or OR4 (N193, N190, N105, N130, N124);
nand NAND3 (N194, N192, N69, N112);
xor XOR2 (N195, N191, N159);
not NOT1 (N196, N172);
nand NAND3 (N197, N184, N12, N138);
not NOT1 (N198, N194);
nor NOR4 (N199, N180, N106, N64, N139);
and AND3 (N200, N189, N19, N76);
nor NOR3 (N201, N199, N140, N155);
or OR3 (N202, N197, N53, N42);
or OR3 (N203, N143, N53, N84);
nor NOR4 (N204, N196, N39, N49, N29);
buf BUF1 (N205, N188);
not NOT1 (N206, N205);
not NOT1 (N207, N186);
and AND4 (N208, N202, N69, N149, N56);
and AND2 (N209, N201, N202);
not NOT1 (N210, N206);
not NOT1 (N211, N200);
nand NAND4 (N212, N198, N192, N89, N72);
xor XOR2 (N213, N208, N76);
buf BUF1 (N214, N209);
buf BUF1 (N215, N212);
buf BUF1 (N216, N207);
nor NOR2 (N217, N213, N153);
nand NAND2 (N218, N214, N177);
nand NAND4 (N219, N216, N180, N7, N77);
nand NAND4 (N220, N219, N90, N59, N211);
nor NOR2 (N221, N21, N186);
not NOT1 (N222, N217);
xor XOR2 (N223, N193, N155);
buf BUF1 (N224, N203);
and AND4 (N225, N195, N115, N172, N113);
not NOT1 (N226, N220);
nand NAND2 (N227, N223, N10);
or OR2 (N228, N210, N198);
not NOT1 (N229, N224);
and AND2 (N230, N225, N122);
and AND2 (N231, N229, N125);
and AND2 (N232, N228, N7);
xor XOR2 (N233, N232, N76);
buf BUF1 (N234, N215);
nand NAND4 (N235, N226, N99, N178, N221);
buf BUF1 (N236, N173);
buf BUF1 (N237, N234);
nand NAND3 (N238, N222, N19, N126);
nor NOR3 (N239, N227, N130, N29);
not NOT1 (N240, N233);
nor NOR2 (N241, N239, N136);
not NOT1 (N242, N240);
and AND3 (N243, N236, N99, N128);
not NOT1 (N244, N230);
not NOT1 (N245, N218);
and AND4 (N246, N204, N3, N206, N152);
and AND2 (N247, N237, N77);
not NOT1 (N248, N247);
buf BUF1 (N249, N244);
buf BUF1 (N250, N249);
xor XOR2 (N251, N238, N238);
not NOT1 (N252, N251);
or OR2 (N253, N252, N156);
or OR3 (N254, N253, N188, N88);
or OR3 (N255, N231, N111, N99);
not NOT1 (N256, N243);
not NOT1 (N257, N242);
nand NAND2 (N258, N246, N80);
not NOT1 (N259, N250);
nor NOR3 (N260, N235, N86, N79);
xor XOR2 (N261, N258, N44);
and AND3 (N262, N248, N17, N48);
or OR3 (N263, N259, N90, N177);
xor XOR2 (N264, N263, N31);
and AND2 (N265, N256, N209);
nand NAND2 (N266, N262, N124);
nand NAND2 (N267, N261, N231);
nor NOR3 (N268, N241, N212, N142);
buf BUF1 (N269, N257);
or OR3 (N270, N268, N53, N182);
and AND4 (N271, N264, N18, N216, N58);
buf BUF1 (N272, N254);
buf BUF1 (N273, N260);
nand NAND2 (N274, N270, N52);
not NOT1 (N275, N265);
buf BUF1 (N276, N272);
nor NOR4 (N277, N276, N233, N208, N102);
xor XOR2 (N278, N269, N15);
xor XOR2 (N279, N277, N46);
or OR4 (N280, N266, N110, N211, N246);
nand NAND3 (N281, N280, N20, N75);
and AND4 (N282, N273, N215, N97, N222);
xor XOR2 (N283, N255, N270);
nor NOR2 (N284, N245, N224);
nor NOR4 (N285, N278, N257, N167, N55);
and AND2 (N286, N275, N23);
or OR3 (N287, N279, N281, N87);
nand NAND4 (N288, N175, N92, N85, N44);
xor XOR2 (N289, N286, N89);
and AND3 (N290, N285, N114, N97);
or OR4 (N291, N274, N46, N200, N275);
not NOT1 (N292, N289);
xor XOR2 (N293, N287, N114);
xor XOR2 (N294, N292, N225);
nand NAND4 (N295, N283, N289, N123, N248);
xor XOR2 (N296, N294, N49);
and AND4 (N297, N296, N233, N18, N269);
nand NAND4 (N298, N284, N262, N198, N181);
nor NOR2 (N299, N267, N133);
buf BUF1 (N300, N297);
nor NOR4 (N301, N288, N58, N80, N257);
xor XOR2 (N302, N301, N182);
not NOT1 (N303, N291);
and AND2 (N304, N282, N63);
nand NAND4 (N305, N298, N191, N245, N247);
buf BUF1 (N306, N271);
xor XOR2 (N307, N293, N284);
and AND2 (N308, N303, N123);
nand NAND4 (N309, N295, N32, N34, N196);
not NOT1 (N310, N302);
xor XOR2 (N311, N300, N48);
nor NOR3 (N312, N290, N131, N133);
or OR3 (N313, N310, N116, N286);
buf BUF1 (N314, N312);
not NOT1 (N315, N304);
nor NOR4 (N316, N308, N22, N40, N124);
buf BUF1 (N317, N299);
or OR4 (N318, N315, N180, N316, N219);
buf BUF1 (N319, N263);
buf BUF1 (N320, N309);
and AND2 (N321, N305, N172);
or OR2 (N322, N320, N115);
nand NAND3 (N323, N317, N203, N124);
and AND3 (N324, N323, N270, N136);
not NOT1 (N325, N321);
nor NOR4 (N326, N319, N293, N325, N49);
xor XOR2 (N327, N49, N20);
nor NOR3 (N328, N311, N199, N116);
or OR4 (N329, N313, N1, N327, N134);
nor NOR3 (N330, N260, N297, N134);
and AND2 (N331, N328, N279);
nand NAND4 (N332, N322, N303, N225, N45);
and AND4 (N333, N332, N94, N204, N257);
buf BUF1 (N334, N331);
nor NOR3 (N335, N314, N163, N31);
nor NOR2 (N336, N334, N22);
and AND3 (N337, N329, N199, N298);
nor NOR3 (N338, N330, N162, N120);
nand NAND3 (N339, N324, N99, N227);
xor XOR2 (N340, N333, N118);
nand NAND3 (N341, N340, N239, N69);
nand NAND3 (N342, N306, N139, N16);
and AND2 (N343, N318, N282);
or OR2 (N344, N307, N113);
nor NOR3 (N345, N337, N310, N327);
nand NAND3 (N346, N344, N50, N330);
xor XOR2 (N347, N339, N262);
not NOT1 (N348, N347);
and AND3 (N349, N338, N219, N243);
xor XOR2 (N350, N341, N127);
nand NAND4 (N351, N342, N67, N219, N150);
or OR4 (N352, N335, N58, N21, N178);
nand NAND4 (N353, N351, N130, N258, N42);
not NOT1 (N354, N343);
not NOT1 (N355, N353);
nand NAND3 (N356, N345, N269, N293);
or OR4 (N357, N355, N207, N179, N102);
not NOT1 (N358, N352);
nand NAND4 (N359, N354, N163, N315, N210);
buf BUF1 (N360, N349);
nor NOR2 (N361, N360, N234);
or OR4 (N362, N361, N292, N129, N343);
xor XOR2 (N363, N346, N324);
and AND3 (N364, N357, N281, N47);
nor NOR3 (N365, N359, N286, N108);
not NOT1 (N366, N326);
nand NAND2 (N367, N365, N301);
not NOT1 (N368, N336);
buf BUF1 (N369, N367);
and AND4 (N370, N366, N163, N106, N159);
or OR4 (N371, N350, N325, N169, N48);
or OR2 (N372, N348, N255);
nand NAND4 (N373, N364, N367, N23, N182);
nor NOR4 (N374, N370, N10, N327, N332);
or OR3 (N375, N374, N53, N212);
xor XOR2 (N376, N375, N20);
and AND4 (N377, N369, N80, N249, N229);
and AND2 (N378, N372, N168);
buf BUF1 (N379, N356);
or OR4 (N380, N373, N164, N74, N268);
or OR2 (N381, N358, N278);
nand NAND4 (N382, N381, N228, N13, N60);
or OR3 (N383, N379, N231, N296);
nand NAND2 (N384, N362, N99);
not NOT1 (N385, N378);
or OR3 (N386, N383, N303, N18);
not NOT1 (N387, N371);
nor NOR2 (N388, N376, N327);
buf BUF1 (N389, N382);
nand NAND2 (N390, N363, N363);
buf BUF1 (N391, N389);
xor XOR2 (N392, N385, N381);
buf BUF1 (N393, N380);
and AND3 (N394, N391, N142, N71);
buf BUF1 (N395, N386);
buf BUF1 (N396, N394);
buf BUF1 (N397, N368);
nand NAND4 (N398, N390, N327, N341, N385);
or OR2 (N399, N397, N110);
and AND3 (N400, N395, N289, N356);
xor XOR2 (N401, N392, N43);
buf BUF1 (N402, N384);
nand NAND2 (N403, N398, N355);
buf BUF1 (N404, N401);
xor XOR2 (N405, N400, N24);
nand NAND2 (N406, N387, N249);
nor NOR3 (N407, N406, N328, N270);
buf BUF1 (N408, N403);
nor NOR2 (N409, N393, N20);
not NOT1 (N410, N377);
nor NOR4 (N411, N399, N397, N192, N90);
buf BUF1 (N412, N404);
nand NAND3 (N413, N388, N92, N308);
not NOT1 (N414, N412);
not NOT1 (N415, N409);
nand NAND4 (N416, N402, N399, N107, N208);
nor NOR2 (N417, N408, N9);
buf BUF1 (N418, N416);
buf BUF1 (N419, N411);
nor NOR3 (N420, N410, N330, N352);
not NOT1 (N421, N414);
buf BUF1 (N422, N415);
nand NAND3 (N423, N420, N79, N60);
nand NAND4 (N424, N421, N274, N43, N293);
nand NAND2 (N425, N405, N149);
or OR2 (N426, N407, N345);
or OR3 (N427, N424, N287, N392);
xor XOR2 (N428, N423, N61);
not NOT1 (N429, N413);
and AND4 (N430, N419, N290, N18, N308);
not NOT1 (N431, N425);
buf BUF1 (N432, N426);
and AND4 (N433, N418, N234, N285, N362);
buf BUF1 (N434, N417);
buf BUF1 (N435, N434);
and AND2 (N436, N422, N169);
nand NAND2 (N437, N429, N393);
nand NAND4 (N438, N427, N53, N203, N248);
nor NOR4 (N439, N437, N171, N47, N356);
not NOT1 (N440, N431);
buf BUF1 (N441, N433);
buf BUF1 (N442, N439);
nor NOR4 (N443, N432, N416, N379, N164);
buf BUF1 (N444, N443);
xor XOR2 (N445, N396, N186);
or OR2 (N446, N438, N365);
and AND4 (N447, N435, N66, N122, N307);
xor XOR2 (N448, N445, N248);
buf BUF1 (N449, N428);
xor XOR2 (N450, N449, N116);
nand NAND3 (N451, N436, N38, N131);
xor XOR2 (N452, N451, N156);
and AND2 (N453, N440, N77);
and AND4 (N454, N450, N18, N374, N313);
nor NOR2 (N455, N453, N2);
xor XOR2 (N456, N430, N353);
nor NOR3 (N457, N444, N244, N88);
xor XOR2 (N458, N442, N446);
buf BUF1 (N459, N438);
nand NAND4 (N460, N458, N185, N434, N133);
nor NOR4 (N461, N454, N163, N255, N175);
and AND4 (N462, N441, N397, N446, N368);
and AND4 (N463, N459, N364, N456, N163);
and AND4 (N464, N347, N292, N124, N29);
and AND4 (N465, N461, N233, N161, N110);
xor XOR2 (N466, N465, N407);
buf BUF1 (N467, N460);
buf BUF1 (N468, N462);
buf BUF1 (N469, N466);
and AND2 (N470, N452, N7);
or OR2 (N471, N463, N403);
nand NAND3 (N472, N457, N454, N140);
nand NAND4 (N473, N469, N62, N308, N264);
not NOT1 (N474, N464);
not NOT1 (N475, N448);
or OR3 (N476, N471, N42, N124);
nor NOR4 (N477, N470, N362, N264, N19);
and AND3 (N478, N455, N321, N391);
or OR4 (N479, N474, N281, N128, N8);
or OR4 (N480, N447, N248, N255, N356);
not NOT1 (N481, N476);
or OR2 (N482, N480, N404);
xor XOR2 (N483, N479, N35);
xor XOR2 (N484, N472, N161);
and AND2 (N485, N475, N160);
nand NAND2 (N486, N481, N347);
buf BUF1 (N487, N485);
not NOT1 (N488, N467);
xor XOR2 (N489, N477, N149);
nand NAND4 (N490, N482, N414, N296, N200);
nor NOR4 (N491, N483, N384, N295, N395);
nor NOR3 (N492, N488, N255, N397);
buf BUF1 (N493, N478);
not NOT1 (N494, N489);
not NOT1 (N495, N486);
and AND3 (N496, N492, N45, N479);
buf BUF1 (N497, N484);
xor XOR2 (N498, N487, N275);
nor NOR2 (N499, N498, N223);
or OR2 (N500, N497, N249);
or OR2 (N501, N499, N105);
xor XOR2 (N502, N490, N192);
not NOT1 (N503, N502);
and AND3 (N504, N501, N439, N42);
or OR4 (N505, N468, N436, N469, N88);
xor XOR2 (N506, N495, N181);
nor NOR3 (N507, N494, N202, N227);
xor XOR2 (N508, N491, N188);
buf BUF1 (N509, N507);
not NOT1 (N510, N500);
nor NOR2 (N511, N504, N463);
xor XOR2 (N512, N473, N277);
and AND3 (N513, N510, N372, N439);
or OR2 (N514, N506, N4);
buf BUF1 (N515, N493);
or OR3 (N516, N503, N461, N135);
xor XOR2 (N517, N505, N44);
nand NAND2 (N518, N517, N370);
not NOT1 (N519, N514);
nand NAND4 (N520, N496, N502, N154, N324);
not NOT1 (N521, N508);
xor XOR2 (N522, N509, N292);
or OR4 (N523, N516, N59, N348, N383);
not NOT1 (N524, N515);
nor NOR4 (N525, N521, N481, N337, N262);
buf BUF1 (N526, N523);
not NOT1 (N527, N513);
not NOT1 (N528, N520);
nor NOR2 (N529, N526, N235);
xor XOR2 (N530, N511, N426);
nor NOR2 (N531, N530, N301);
and AND4 (N532, N527, N407, N215, N48);
nor NOR2 (N533, N532, N504);
nand NAND2 (N534, N531, N251);
not NOT1 (N535, N524);
nand NAND2 (N536, N522, N360);
buf BUF1 (N537, N518);
buf BUF1 (N538, N528);
and AND4 (N539, N536, N37, N92, N126);
or OR4 (N540, N519, N62, N260, N442);
buf BUF1 (N541, N534);
nor NOR2 (N542, N533, N254);
xor XOR2 (N543, N525, N128);
or OR2 (N544, N535, N510);
not NOT1 (N545, N512);
nand NAND2 (N546, N539, N345);
or OR4 (N547, N529, N425, N263, N194);
xor XOR2 (N548, N543, N125);
and AND2 (N549, N544, N64);
not NOT1 (N550, N545);
buf BUF1 (N551, N548);
nand NAND4 (N552, N537, N21, N35, N526);
and AND4 (N553, N552, N157, N116, N304);
or OR4 (N554, N546, N207, N337, N253);
xor XOR2 (N555, N538, N97);
and AND2 (N556, N549, N35);
or OR3 (N557, N555, N334, N102);
or OR2 (N558, N540, N428);
or OR2 (N559, N557, N145);
or OR3 (N560, N547, N543, N109);
nand NAND3 (N561, N550, N315, N151);
nor NOR2 (N562, N542, N449);
or OR2 (N563, N560, N546);
buf BUF1 (N564, N562);
and AND3 (N565, N553, N471, N547);
xor XOR2 (N566, N565, N528);
not NOT1 (N567, N541);
not NOT1 (N568, N551);
not NOT1 (N569, N564);
nand NAND4 (N570, N554, N155, N43, N84);
buf BUF1 (N571, N561);
not NOT1 (N572, N558);
nor NOR4 (N573, N571, N171, N327, N109);
not NOT1 (N574, N566);
nand NAND3 (N575, N574, N305, N283);
xor XOR2 (N576, N568, N360);
nor NOR3 (N577, N575, N92, N47);
and AND4 (N578, N577, N414, N215, N120);
and AND3 (N579, N572, N34, N182);
not NOT1 (N580, N579);
xor XOR2 (N581, N559, N70);
nor NOR3 (N582, N576, N456, N122);
or OR4 (N583, N581, N71, N416, N167);
xor XOR2 (N584, N569, N468);
buf BUF1 (N585, N580);
and AND2 (N586, N556, N119);
nand NAND2 (N587, N567, N436);
or OR4 (N588, N570, N552, N306, N509);
or OR4 (N589, N578, N374, N100, N361);
nor NOR4 (N590, N586, N63, N436, N35);
not NOT1 (N591, N582);
and AND4 (N592, N563, N359, N454, N552);
and AND3 (N593, N584, N103, N303);
and AND4 (N594, N591, N477, N405, N572);
and AND3 (N595, N590, N33, N101);
and AND2 (N596, N585, N85);
or OR2 (N597, N594, N563);
and AND4 (N598, N595, N80, N409, N234);
or OR3 (N599, N588, N416, N373);
nand NAND4 (N600, N573, N56, N288, N247);
not NOT1 (N601, N593);
buf BUF1 (N602, N598);
not NOT1 (N603, N602);
nor NOR2 (N604, N583, N285);
and AND2 (N605, N599, N53);
buf BUF1 (N606, N596);
nand NAND4 (N607, N606, N5, N190, N355);
xor XOR2 (N608, N592, N245);
xor XOR2 (N609, N601, N466);
and AND2 (N610, N605, N155);
nand NAND4 (N611, N589, N320, N316, N100);
or OR2 (N612, N604, N465);
xor XOR2 (N613, N611, N556);
and AND2 (N614, N587, N251);
and AND3 (N615, N610, N116, N159);
nand NAND4 (N616, N614, N11, N577, N288);
nor NOR3 (N617, N612, N506, N246);
xor XOR2 (N618, N608, N433);
or OR2 (N619, N600, N569);
nand NAND4 (N620, N615, N357, N444, N3);
not NOT1 (N621, N617);
or OR4 (N622, N613, N346, N520, N158);
buf BUF1 (N623, N618);
and AND2 (N624, N597, N447);
nor NOR2 (N625, N622, N526);
nand NAND3 (N626, N616, N439, N68);
nor NOR3 (N627, N625, N57, N282);
and AND2 (N628, N607, N270);
buf BUF1 (N629, N624);
or OR3 (N630, N620, N293, N171);
or OR2 (N631, N619, N238);
nand NAND3 (N632, N631, N507, N575);
and AND3 (N633, N623, N505, N392);
nand NAND2 (N634, N630, N435);
xor XOR2 (N635, N626, N417);
xor XOR2 (N636, N632, N34);
nand NAND2 (N637, N609, N221);
or OR4 (N638, N629, N216, N249, N477);
nor NOR3 (N639, N634, N422, N385);
and AND3 (N640, N636, N217, N538);
and AND2 (N641, N628, N162);
nand NAND2 (N642, N621, N308);
not NOT1 (N643, N627);
and AND4 (N644, N642, N384, N224, N560);
nand NAND3 (N645, N638, N472, N593);
not NOT1 (N646, N641);
buf BUF1 (N647, N633);
not NOT1 (N648, N635);
nand NAND3 (N649, N644, N31, N580);
or OR3 (N650, N647, N160, N343);
nor NOR3 (N651, N649, N97, N342);
buf BUF1 (N652, N643);
nand NAND2 (N653, N603, N94);
or OR3 (N654, N646, N17, N252);
nand NAND4 (N655, N651, N162, N32, N428);
not NOT1 (N656, N637);
nand NAND3 (N657, N640, N439, N242);
nand NAND4 (N658, N657, N28, N288, N105);
nor NOR4 (N659, N654, N134, N396, N325);
nor NOR2 (N660, N655, N659);
nor NOR2 (N661, N162, N441);
or OR4 (N662, N656, N365, N217, N87);
nand NAND3 (N663, N648, N249, N568);
nor NOR2 (N664, N663, N332);
not NOT1 (N665, N661);
or OR4 (N666, N652, N650, N52, N528);
buf BUF1 (N667, N354);
nor NOR3 (N668, N653, N406, N205);
nor NOR4 (N669, N662, N112, N181, N381);
xor XOR2 (N670, N639, N187);
xor XOR2 (N671, N667, N90);
nor NOR2 (N672, N666, N338);
buf BUF1 (N673, N664);
and AND3 (N674, N658, N532, N44);
xor XOR2 (N675, N645, N403);
nand NAND2 (N676, N669, N367);
nand NAND2 (N677, N668, N554);
nand NAND2 (N678, N675, N172);
or OR3 (N679, N676, N147, N105);
and AND3 (N680, N673, N280, N597);
nand NAND3 (N681, N679, N430, N344);
nor NOR4 (N682, N671, N426, N124, N507);
not NOT1 (N683, N680);
buf BUF1 (N684, N672);
xor XOR2 (N685, N677, N445);
and AND2 (N686, N670, N191);
nor NOR2 (N687, N678, N462);
nor NOR3 (N688, N674, N110, N652);
not NOT1 (N689, N665);
and AND3 (N690, N683, N140, N149);
nand NAND3 (N691, N687, N186, N1);
nand NAND4 (N692, N685, N158, N445, N147);
nand NAND4 (N693, N688, N298, N349, N411);
or OR4 (N694, N692, N202, N11, N23);
and AND2 (N695, N694, N397);
nand NAND3 (N696, N684, N173, N299);
xor XOR2 (N697, N691, N459);
buf BUF1 (N698, N682);
not NOT1 (N699, N695);
not NOT1 (N700, N693);
nand NAND2 (N701, N697, N451);
xor XOR2 (N702, N700, N40);
nor NOR2 (N703, N699, N671);
not NOT1 (N704, N703);
xor XOR2 (N705, N701, N160);
or OR4 (N706, N704, N144, N637, N232);
or OR3 (N707, N686, N368, N327);
buf BUF1 (N708, N698);
nor NOR2 (N709, N690, N703);
xor XOR2 (N710, N696, N43);
nand NAND3 (N711, N710, N601, N611);
or OR4 (N712, N681, N355, N384, N275);
buf BUF1 (N713, N709);
nand NAND3 (N714, N712, N493, N321);
nand NAND3 (N715, N707, N68, N392);
not NOT1 (N716, N708);
or OR3 (N717, N713, N465, N147);
buf BUF1 (N718, N705);
nor NOR3 (N719, N689, N345, N442);
xor XOR2 (N720, N660, N631);
nand NAND3 (N721, N714, N527, N608);
buf BUF1 (N722, N720);
and AND3 (N723, N721, N482, N434);
nand NAND4 (N724, N711, N414, N412, N354);
not NOT1 (N725, N717);
nand NAND2 (N726, N722, N150);
not NOT1 (N727, N723);
not NOT1 (N728, N727);
nand NAND3 (N729, N715, N389, N700);
buf BUF1 (N730, N718);
and AND3 (N731, N728, N126, N372);
and AND4 (N732, N731, N59, N305, N330);
xor XOR2 (N733, N725, N412);
nor NOR2 (N734, N706, N654);
nand NAND4 (N735, N716, N177, N488, N91);
buf BUF1 (N736, N730);
nor NOR4 (N737, N724, N194, N67, N439);
xor XOR2 (N738, N732, N85);
xor XOR2 (N739, N738, N303);
xor XOR2 (N740, N729, N139);
xor XOR2 (N741, N719, N251);
or OR3 (N742, N735, N255, N714);
xor XOR2 (N743, N740, N620);
xor XOR2 (N744, N737, N592);
xor XOR2 (N745, N726, N437);
buf BUF1 (N746, N702);
buf BUF1 (N747, N741);
buf BUF1 (N748, N746);
or OR4 (N749, N748, N329, N552, N319);
nand NAND2 (N750, N733, N337);
not NOT1 (N751, N747);
or OR3 (N752, N745, N682, N40);
nand NAND3 (N753, N744, N589, N449);
nor NOR4 (N754, N742, N13, N41, N146);
or OR3 (N755, N734, N213, N599);
or OR3 (N756, N752, N323, N474);
nand NAND4 (N757, N750, N379, N208, N314);
nor NOR3 (N758, N751, N134, N617);
nor NOR2 (N759, N755, N2);
buf BUF1 (N760, N759);
not NOT1 (N761, N753);
nand NAND2 (N762, N739, N397);
and AND3 (N763, N743, N415, N565);
or OR2 (N764, N763, N569);
or OR2 (N765, N736, N341);
not NOT1 (N766, N762);
and AND3 (N767, N761, N79, N588);
nor NOR4 (N768, N756, N71, N162, N757);
xor XOR2 (N769, N227, N626);
buf BUF1 (N770, N765);
nand NAND3 (N771, N749, N626, N9);
and AND2 (N772, N769, N385);
and AND4 (N773, N770, N431, N59, N334);
and AND2 (N774, N772, N23);
or OR2 (N775, N768, N586);
not NOT1 (N776, N767);
not NOT1 (N777, N773);
xor XOR2 (N778, N758, N435);
xor XOR2 (N779, N778, N354);
and AND4 (N780, N776, N762, N770, N452);
not NOT1 (N781, N754);
xor XOR2 (N782, N777, N413);
xor XOR2 (N783, N782, N499);
not NOT1 (N784, N771);
or OR3 (N785, N764, N770, N487);
nor NOR2 (N786, N766, N394);
nor NOR2 (N787, N783, N381);
nand NAND3 (N788, N781, N531, N131);
xor XOR2 (N789, N785, N244);
buf BUF1 (N790, N774);
nor NOR3 (N791, N786, N33, N149);
not NOT1 (N792, N775);
buf BUF1 (N793, N788);
xor XOR2 (N794, N784, N487);
nand NAND3 (N795, N791, N230, N500);
xor XOR2 (N796, N760, N370);
nand NAND4 (N797, N787, N285, N213, N157);
xor XOR2 (N798, N794, N793);
not NOT1 (N799, N180);
or OR3 (N800, N799, N674, N267);
nand NAND4 (N801, N795, N130, N98, N421);
not NOT1 (N802, N798);
xor XOR2 (N803, N789, N50);
not NOT1 (N804, N800);
or OR3 (N805, N779, N566, N160);
or OR3 (N806, N792, N716, N784);
xor XOR2 (N807, N806, N435);
and AND3 (N808, N807, N779, N192);
and AND4 (N809, N802, N714, N670, N660);
nand NAND3 (N810, N780, N790, N352);
not NOT1 (N811, N387);
xor XOR2 (N812, N796, N300);
and AND4 (N813, N808, N113, N482, N441);
or OR2 (N814, N809, N170);
not NOT1 (N815, N803);
xor XOR2 (N816, N804, N813);
or OR3 (N817, N4, N712, N433);
nor NOR4 (N818, N812, N246, N1, N238);
not NOT1 (N819, N818);
nor NOR3 (N820, N810, N94, N46);
xor XOR2 (N821, N819, N622);
endmodule