// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N915,N908,N913,N921,N916,N919,N911,N920,N917,N922;

nor NOR4 (N23, N13, N5, N12, N21);
or OR2 (N24, N6, N3);
and AND2 (N25, N8, N20);
or OR4 (N26, N16, N24, N15, N15);
nor NOR2 (N27, N11, N13);
and AND4 (N28, N14, N8, N2, N7);
and AND4 (N29, N24, N4, N13, N28);
nor NOR4 (N30, N5, N7, N29, N2);
nor NOR4 (N31, N9, N14, N23, N16);
buf BUF1 (N32, N22);
not NOT1 (N33, N20);
buf BUF1 (N34, N32);
nand NAND4 (N35, N19, N20, N28, N28);
xor XOR2 (N36, N31, N20);
xor XOR2 (N37, N19, N24);
or OR2 (N38, N35, N16);
nand NAND4 (N39, N25, N21, N1, N38);
not NOT1 (N40, N6);
buf BUF1 (N41, N35);
buf BUF1 (N42, N36);
and AND2 (N43, N27, N33);
or OR4 (N44, N7, N1, N11, N5);
nand NAND3 (N45, N39, N17, N10);
not NOT1 (N46, N41);
buf BUF1 (N47, N30);
buf BUF1 (N48, N40);
and AND3 (N49, N45, N31, N47);
nand NAND2 (N50, N2, N2);
and AND2 (N51, N49, N37);
not NOT1 (N52, N45);
or OR4 (N53, N51, N18, N51, N2);
nor NOR4 (N54, N42, N15, N49, N45);
nor NOR2 (N55, N26, N35);
xor XOR2 (N56, N55, N34);
not NOT1 (N57, N35);
not NOT1 (N58, N54);
nand NAND3 (N59, N56, N16, N18);
not NOT1 (N60, N43);
xor XOR2 (N61, N50, N16);
not NOT1 (N62, N52);
nand NAND3 (N63, N59, N60, N18);
not NOT1 (N64, N38);
or OR4 (N65, N63, N59, N50, N28);
or OR2 (N66, N57, N63);
nand NAND4 (N67, N65, N46, N26, N20);
nand NAND3 (N68, N38, N54, N17);
buf BUF1 (N69, N61);
and AND2 (N70, N53, N57);
buf BUF1 (N71, N67);
and AND4 (N72, N69, N10, N1, N3);
buf BUF1 (N73, N71);
buf BUF1 (N74, N48);
nor NOR4 (N75, N44, N37, N10, N17);
buf BUF1 (N76, N75);
xor XOR2 (N77, N74, N71);
not NOT1 (N78, N72);
nand NAND2 (N79, N58, N76);
buf BUF1 (N80, N53);
xor XOR2 (N81, N79, N46);
buf BUF1 (N82, N78);
or OR4 (N83, N81, N79, N16, N76);
nand NAND4 (N84, N82, N17, N45, N32);
nor NOR2 (N85, N68, N22);
not NOT1 (N86, N80);
buf BUF1 (N87, N83);
buf BUF1 (N88, N66);
buf BUF1 (N89, N64);
nor NOR2 (N90, N88, N86);
or OR4 (N91, N42, N30, N89, N10);
nor NOR2 (N92, N35, N60);
and AND4 (N93, N90, N21, N67, N84);
or OR4 (N94, N17, N14, N10, N55);
nor NOR4 (N95, N62, N90, N68, N38);
nand NAND4 (N96, N73, N64, N47, N10);
or OR4 (N97, N87, N80, N51, N73);
not NOT1 (N98, N85);
and AND3 (N99, N92, N77, N40);
and AND2 (N100, N41, N80);
buf BUF1 (N101, N93);
xor XOR2 (N102, N70, N52);
xor XOR2 (N103, N95, N19);
buf BUF1 (N104, N103);
buf BUF1 (N105, N91);
nor NOR2 (N106, N96, N50);
buf BUF1 (N107, N99);
and AND2 (N108, N100, N86);
and AND3 (N109, N107, N30, N16);
nor NOR3 (N110, N97, N68, N3);
and AND4 (N111, N102, N39, N56, N14);
xor XOR2 (N112, N111, N82);
not NOT1 (N113, N94);
and AND3 (N114, N113, N66, N19);
buf BUF1 (N115, N112);
xor XOR2 (N116, N105, N73);
not NOT1 (N117, N98);
and AND3 (N118, N117, N44, N53);
xor XOR2 (N119, N114, N32);
not NOT1 (N120, N119);
buf BUF1 (N121, N116);
xor XOR2 (N122, N118, N10);
xor XOR2 (N123, N110, N49);
nor NOR4 (N124, N109, N12, N22, N37);
nor NOR4 (N125, N122, N102, N59, N21);
xor XOR2 (N126, N106, N105);
xor XOR2 (N127, N124, N32);
nand NAND3 (N128, N123, N107, N68);
buf BUF1 (N129, N128);
nor NOR3 (N130, N129, N53, N80);
or OR2 (N131, N121, N79);
nor NOR3 (N132, N104, N112, N24);
buf BUF1 (N133, N120);
nand NAND3 (N134, N115, N16, N3);
xor XOR2 (N135, N101, N56);
nor NOR2 (N136, N134, N40);
buf BUF1 (N137, N133);
buf BUF1 (N138, N132);
or OR4 (N139, N137, N84, N128, N63);
xor XOR2 (N140, N139, N134);
buf BUF1 (N141, N138);
and AND4 (N142, N126, N47, N85, N132);
buf BUF1 (N143, N108);
xor XOR2 (N144, N141, N55);
nand NAND3 (N145, N136, N4, N118);
not NOT1 (N146, N140);
buf BUF1 (N147, N125);
buf BUF1 (N148, N135);
not NOT1 (N149, N131);
buf BUF1 (N150, N147);
or OR4 (N151, N145, N64, N5, N134);
not NOT1 (N152, N149);
or OR2 (N153, N130, N20);
nor NOR3 (N154, N148, N116, N95);
or OR3 (N155, N152, N149, N46);
buf BUF1 (N156, N155);
buf BUF1 (N157, N154);
not NOT1 (N158, N143);
nor NOR3 (N159, N150, N115, N95);
or OR4 (N160, N153, N158, N18, N9);
nand NAND2 (N161, N9, N71);
and AND4 (N162, N127, N29, N105, N148);
nand NAND2 (N163, N159, N125);
nand NAND3 (N164, N146, N48, N89);
or OR3 (N165, N151, N105, N35);
nand NAND2 (N166, N160, N155);
not NOT1 (N167, N162);
not NOT1 (N168, N157);
nor NOR4 (N169, N163, N16, N52, N87);
and AND3 (N170, N164, N158, N97);
nand NAND3 (N171, N169, N164, N81);
or OR3 (N172, N161, N152, N99);
or OR4 (N173, N167, N120, N40, N122);
nor NOR2 (N174, N173, N1);
nor NOR2 (N175, N156, N8);
and AND4 (N176, N172, N101, N167, N83);
not NOT1 (N177, N142);
nor NOR4 (N178, N168, N120, N50, N39);
buf BUF1 (N179, N176);
nor NOR3 (N180, N165, N25, N116);
or OR2 (N181, N180, N168);
not NOT1 (N182, N178);
nand NAND2 (N183, N179, N28);
or OR4 (N184, N174, N76, N106, N70);
not NOT1 (N185, N144);
and AND3 (N186, N184, N21, N88);
not NOT1 (N187, N185);
not NOT1 (N188, N183);
not NOT1 (N189, N187);
nor NOR4 (N190, N175, N189, N89, N114);
nor NOR3 (N191, N128, N141, N179);
or OR4 (N192, N186, N29, N54, N175);
not NOT1 (N193, N177);
or OR4 (N194, N193, N21, N38, N90);
or OR2 (N195, N191, N131);
xor XOR2 (N196, N194, N189);
xor XOR2 (N197, N166, N195);
not NOT1 (N198, N90);
not NOT1 (N199, N171);
nor NOR2 (N200, N170, N151);
xor XOR2 (N201, N192, N23);
xor XOR2 (N202, N199, N37);
or OR3 (N203, N198, N45, N65);
nand NAND2 (N204, N182, N4);
or OR3 (N205, N188, N58, N120);
buf BUF1 (N206, N205);
buf BUF1 (N207, N206);
not NOT1 (N208, N200);
nand NAND3 (N209, N207, N12, N46);
buf BUF1 (N210, N204);
or OR3 (N211, N196, N110, N158);
buf BUF1 (N212, N202);
or OR3 (N213, N209, N44, N51);
not NOT1 (N214, N213);
and AND3 (N215, N181, N67, N48);
or OR2 (N216, N210, N70);
buf BUF1 (N217, N197);
buf BUF1 (N218, N201);
xor XOR2 (N219, N215, N66);
nor NOR3 (N220, N208, N139, N170);
xor XOR2 (N221, N216, N134);
buf BUF1 (N222, N219);
not NOT1 (N223, N214);
xor XOR2 (N224, N220, N5);
not NOT1 (N225, N222);
buf BUF1 (N226, N221);
or OR4 (N227, N203, N222, N8, N188);
nand NAND2 (N228, N226, N10);
xor XOR2 (N229, N227, N63);
not NOT1 (N230, N217);
or OR3 (N231, N223, N39, N163);
and AND3 (N232, N224, N186, N79);
nand NAND4 (N233, N232, N21, N60, N97);
nand NAND4 (N234, N233, N20, N223, N141);
buf BUF1 (N235, N218);
nand NAND4 (N236, N190, N150, N170, N9);
nand NAND4 (N237, N230, N187, N115, N46);
buf BUF1 (N238, N211);
buf BUF1 (N239, N234);
nor NOR2 (N240, N229, N57);
or OR2 (N241, N236, N111);
or OR4 (N242, N240, N234, N190, N25);
nor NOR3 (N243, N241, N205, N192);
and AND2 (N244, N231, N235);
buf BUF1 (N245, N40);
and AND2 (N246, N244, N160);
not NOT1 (N247, N237);
not NOT1 (N248, N239);
and AND2 (N249, N248, N51);
buf BUF1 (N250, N246);
nand NAND2 (N251, N228, N210);
xor XOR2 (N252, N242, N44);
xor XOR2 (N253, N245, N36);
and AND3 (N254, N251, N250, N203);
xor XOR2 (N255, N117, N200);
not NOT1 (N256, N243);
nor NOR4 (N257, N254, N247, N97, N77);
and AND3 (N258, N92, N1, N245);
buf BUF1 (N259, N253);
and AND3 (N260, N258, N83, N231);
or OR3 (N261, N255, N153, N65);
nand NAND3 (N262, N212, N152, N36);
or OR3 (N263, N257, N14, N249);
xor XOR2 (N264, N174, N115);
nand NAND3 (N265, N256, N227, N189);
buf BUF1 (N266, N263);
nor NOR3 (N267, N266, N252, N143);
xor XOR2 (N268, N116, N256);
and AND2 (N269, N238, N161);
buf BUF1 (N270, N261);
nor NOR2 (N271, N262, N94);
not NOT1 (N272, N265);
and AND2 (N273, N259, N164);
not NOT1 (N274, N273);
buf BUF1 (N275, N260);
xor XOR2 (N276, N268, N13);
nor NOR2 (N277, N272, N227);
not NOT1 (N278, N269);
nand NAND2 (N279, N276, N85);
nand NAND3 (N280, N279, N99, N126);
nand NAND4 (N281, N275, N82, N57, N93);
buf BUF1 (N282, N271);
nor NOR3 (N283, N281, N107, N43);
or OR2 (N284, N283, N211);
not NOT1 (N285, N278);
nand NAND4 (N286, N284, N46, N204, N258);
and AND4 (N287, N280, N86, N16, N218);
buf BUF1 (N288, N225);
nor NOR2 (N289, N286, N276);
or OR2 (N290, N274, N204);
buf BUF1 (N291, N277);
or OR2 (N292, N287, N44);
xor XOR2 (N293, N289, N112);
nor NOR3 (N294, N267, N116, N141);
or OR3 (N295, N288, N231, N200);
and AND2 (N296, N293, N19);
not NOT1 (N297, N270);
nand NAND4 (N298, N264, N66, N134, N182);
or OR2 (N299, N285, N246);
not NOT1 (N300, N297);
or OR3 (N301, N298, N94, N35);
and AND2 (N302, N295, N265);
nor NOR3 (N303, N291, N83, N13);
nand NAND4 (N304, N296, N162, N40, N13);
nor NOR3 (N305, N303, N270, N152);
nand NAND3 (N306, N300, N114, N153);
nor NOR2 (N307, N305, N49);
and AND2 (N308, N302, N279);
nor NOR4 (N309, N294, N225, N209, N9);
and AND2 (N310, N301, N91);
nor NOR3 (N311, N290, N241, N10);
or OR2 (N312, N282, N23);
buf BUF1 (N313, N307);
and AND2 (N314, N310, N122);
buf BUF1 (N315, N314);
nor NOR3 (N316, N306, N264, N264);
and AND2 (N317, N311, N32);
or OR3 (N318, N316, N203, N48);
xor XOR2 (N319, N313, N1);
xor XOR2 (N320, N309, N243);
xor XOR2 (N321, N318, N75);
xor XOR2 (N322, N315, N200);
nand NAND3 (N323, N312, N207, N251);
and AND3 (N324, N322, N287, N52);
and AND3 (N325, N323, N193, N236);
nand NAND4 (N326, N324, N31, N226, N236);
buf BUF1 (N327, N292);
buf BUF1 (N328, N325);
buf BUF1 (N329, N319);
not NOT1 (N330, N317);
xor XOR2 (N331, N330, N297);
nor NOR3 (N332, N308, N97, N276);
nor NOR3 (N333, N329, N207, N302);
and AND3 (N334, N328, N22, N152);
and AND3 (N335, N299, N154, N250);
not NOT1 (N336, N321);
and AND3 (N337, N336, N206, N35);
nor NOR2 (N338, N333, N79);
and AND4 (N339, N335, N37, N225, N171);
or OR4 (N340, N304, N314, N157, N176);
xor XOR2 (N341, N337, N112);
nor NOR2 (N342, N334, N94);
not NOT1 (N343, N327);
not NOT1 (N344, N342);
nand NAND4 (N345, N344, N162, N23, N53);
nor NOR2 (N346, N341, N326);
and AND3 (N347, N208, N279, N139);
and AND2 (N348, N339, N85);
nand NAND4 (N349, N332, N297, N305, N215);
or OR3 (N350, N348, N349, N341);
not NOT1 (N351, N99);
buf BUF1 (N352, N340);
and AND2 (N353, N346, N158);
or OR4 (N354, N320, N226, N142, N29);
or OR2 (N355, N338, N93);
and AND4 (N356, N355, N306, N277, N275);
xor XOR2 (N357, N352, N243);
nand NAND4 (N358, N356, N1, N137, N336);
and AND4 (N359, N354, N99, N212, N177);
nand NAND2 (N360, N345, N134);
or OR4 (N361, N347, N33, N31, N289);
and AND3 (N362, N343, N263, N319);
nand NAND2 (N363, N359, N5);
buf BUF1 (N364, N358);
and AND2 (N365, N353, N238);
and AND3 (N366, N351, N248, N301);
not NOT1 (N367, N357);
buf BUF1 (N368, N366);
and AND3 (N369, N365, N42, N94);
nor NOR2 (N370, N331, N204);
buf BUF1 (N371, N363);
nor NOR4 (N372, N364, N189, N62, N328);
nand NAND2 (N373, N367, N293);
or OR3 (N374, N361, N55, N32);
and AND3 (N375, N370, N304, N3);
and AND4 (N376, N350, N276, N126, N97);
nor NOR4 (N377, N368, N288, N291, N228);
nand NAND4 (N378, N376, N342, N113, N135);
not NOT1 (N379, N369);
not NOT1 (N380, N375);
xor XOR2 (N381, N362, N378);
xor XOR2 (N382, N80, N304);
or OR2 (N383, N380, N224);
buf BUF1 (N384, N383);
buf BUF1 (N385, N373);
nand NAND2 (N386, N374, N73);
and AND3 (N387, N386, N297, N109);
or OR2 (N388, N381, N97);
nor NOR4 (N389, N379, N278, N165, N105);
and AND2 (N390, N387, N92);
nand NAND3 (N391, N385, N390, N380);
buf BUF1 (N392, N231);
nand NAND2 (N393, N371, N347);
and AND3 (N394, N384, N72, N12);
not NOT1 (N395, N393);
or OR2 (N396, N395, N6);
not NOT1 (N397, N391);
buf BUF1 (N398, N396);
not NOT1 (N399, N398);
nor NOR3 (N400, N389, N330, N86);
not NOT1 (N401, N388);
buf BUF1 (N402, N400);
not NOT1 (N403, N382);
buf BUF1 (N404, N360);
buf BUF1 (N405, N402);
xor XOR2 (N406, N372, N291);
and AND4 (N407, N404, N118, N181, N222);
nand NAND2 (N408, N403, N204);
and AND3 (N409, N399, N358, N375);
nand NAND3 (N410, N409, N41, N107);
xor XOR2 (N411, N405, N118);
buf BUF1 (N412, N406);
not NOT1 (N413, N377);
not NOT1 (N414, N408);
not NOT1 (N415, N401);
or OR4 (N416, N407, N375, N248, N320);
and AND2 (N417, N411, N11);
not NOT1 (N418, N416);
buf BUF1 (N419, N414);
not NOT1 (N420, N413);
and AND2 (N421, N415, N134);
or OR3 (N422, N410, N40, N242);
buf BUF1 (N423, N420);
or OR4 (N424, N392, N306, N23, N148);
xor XOR2 (N425, N394, N126);
xor XOR2 (N426, N418, N148);
and AND2 (N427, N421, N118);
xor XOR2 (N428, N425, N375);
nor NOR4 (N429, N423, N73, N422, N113);
nor NOR4 (N430, N286, N188, N31, N360);
nand NAND3 (N431, N397, N258, N287);
nor NOR2 (N432, N430, N22);
nand NAND2 (N433, N417, N233);
not NOT1 (N434, N433);
buf BUF1 (N435, N427);
not NOT1 (N436, N429);
not NOT1 (N437, N432);
and AND4 (N438, N412, N250, N353, N127);
nor NOR4 (N439, N431, N63, N139, N277);
xor XOR2 (N440, N434, N404);
nor NOR3 (N441, N438, N191, N40);
nor NOR4 (N442, N419, N99, N409, N111);
and AND4 (N443, N436, N375, N390, N72);
not NOT1 (N444, N435);
xor XOR2 (N445, N428, N167);
buf BUF1 (N446, N426);
nand NAND3 (N447, N442, N21, N312);
buf BUF1 (N448, N446);
not NOT1 (N449, N444);
not NOT1 (N450, N448);
or OR4 (N451, N445, N429, N407, N24);
nand NAND2 (N452, N451, N49);
or OR3 (N453, N452, N130, N417);
nor NOR3 (N454, N443, N201, N352);
xor XOR2 (N455, N454, N446);
and AND3 (N456, N453, N453, N149);
not NOT1 (N457, N447);
nand NAND3 (N458, N424, N113, N395);
buf BUF1 (N459, N437);
and AND2 (N460, N441, N250);
buf BUF1 (N461, N440);
or OR3 (N462, N460, N206, N111);
xor XOR2 (N463, N459, N393);
xor XOR2 (N464, N449, N59);
and AND4 (N465, N463, N399, N39, N356);
nor NOR2 (N466, N458, N146);
xor XOR2 (N467, N462, N353);
nor NOR4 (N468, N467, N322, N14, N315);
not NOT1 (N469, N455);
nor NOR2 (N470, N468, N121);
or OR3 (N471, N450, N207, N329);
nand NAND3 (N472, N465, N446, N409);
and AND4 (N473, N439, N241, N116, N262);
or OR3 (N474, N461, N279, N1);
xor XOR2 (N475, N466, N146);
not NOT1 (N476, N457);
nor NOR3 (N477, N472, N158, N438);
xor XOR2 (N478, N477, N236);
not NOT1 (N479, N456);
buf BUF1 (N480, N478);
nand NAND3 (N481, N475, N242, N284);
buf BUF1 (N482, N474);
buf BUF1 (N483, N476);
not NOT1 (N484, N473);
and AND2 (N485, N480, N146);
buf BUF1 (N486, N483);
nand NAND3 (N487, N482, N56, N41);
buf BUF1 (N488, N479);
and AND3 (N489, N484, N198, N6);
nor NOR4 (N490, N488, N13, N436, N150);
nand NAND3 (N491, N469, N338, N131);
nand NAND3 (N492, N464, N273, N468);
buf BUF1 (N493, N470);
xor XOR2 (N494, N471, N12);
nor NOR3 (N495, N491, N412, N216);
nor NOR4 (N496, N493, N364, N292, N145);
buf BUF1 (N497, N496);
buf BUF1 (N498, N492);
nand NAND2 (N499, N485, N77);
nand NAND3 (N500, N490, N210, N159);
buf BUF1 (N501, N495);
nand NAND2 (N502, N498, N80);
nor NOR3 (N503, N489, N327, N208);
not NOT1 (N504, N503);
or OR3 (N505, N494, N469, N501);
not NOT1 (N506, N242);
nor NOR2 (N507, N497, N418);
buf BUF1 (N508, N481);
nor NOR3 (N509, N499, N507, N18);
nor NOR3 (N510, N59, N175, N15);
or OR2 (N511, N508, N439);
buf BUF1 (N512, N502);
nor NOR4 (N513, N512, N100, N104, N500);
not NOT1 (N514, N335);
or OR4 (N515, N506, N11, N3, N414);
nor NOR4 (N516, N504, N22, N41, N355);
nand NAND2 (N517, N516, N157);
and AND4 (N518, N510, N517, N451, N263);
nand NAND2 (N519, N68, N186);
nor NOR4 (N520, N505, N222, N192, N270);
not NOT1 (N521, N487);
nor NOR2 (N522, N513, N505);
nor NOR4 (N523, N519, N256, N475, N259);
buf BUF1 (N524, N509);
not NOT1 (N525, N522);
xor XOR2 (N526, N518, N335);
and AND2 (N527, N520, N488);
nor NOR4 (N528, N514, N368, N180, N125);
buf BUF1 (N529, N511);
buf BUF1 (N530, N528);
and AND2 (N531, N524, N147);
or OR3 (N532, N523, N93, N305);
xor XOR2 (N533, N526, N262);
buf BUF1 (N534, N521);
xor XOR2 (N535, N529, N461);
nor NOR3 (N536, N531, N38, N465);
and AND4 (N537, N486, N423, N230, N275);
xor XOR2 (N538, N515, N190);
nand NAND2 (N539, N530, N447);
or OR2 (N540, N533, N408);
nor NOR4 (N541, N532, N455, N81, N252);
and AND3 (N542, N525, N314, N282);
nand NAND4 (N543, N541, N368, N293, N417);
not NOT1 (N544, N534);
or OR4 (N545, N544, N281, N86, N20);
or OR2 (N546, N539, N380);
and AND2 (N547, N545, N126);
or OR4 (N548, N535, N220, N510, N166);
nand NAND3 (N549, N542, N455, N277);
not NOT1 (N550, N536);
nor NOR3 (N551, N543, N499, N369);
buf BUF1 (N552, N551);
not NOT1 (N553, N552);
or OR4 (N554, N538, N110, N464, N98);
or OR3 (N555, N546, N138, N409);
and AND2 (N556, N540, N496);
xor XOR2 (N557, N547, N60);
not NOT1 (N558, N549);
nor NOR4 (N559, N555, N315, N78, N543);
buf BUF1 (N560, N557);
xor XOR2 (N561, N527, N408);
nand NAND2 (N562, N559, N67);
xor XOR2 (N563, N562, N528);
and AND4 (N564, N553, N134, N167, N34);
buf BUF1 (N565, N548);
xor XOR2 (N566, N537, N456);
and AND3 (N567, N558, N503, N392);
nand NAND3 (N568, N554, N69, N331);
nor NOR2 (N569, N556, N81);
nor NOR3 (N570, N565, N151, N207);
not NOT1 (N571, N569);
nand NAND3 (N572, N560, N470, N437);
or OR4 (N573, N564, N327, N512, N332);
nor NOR3 (N574, N563, N539, N194);
and AND2 (N575, N568, N312);
or OR3 (N576, N561, N559, N45);
xor XOR2 (N577, N572, N116);
nor NOR2 (N578, N567, N524);
and AND4 (N579, N550, N101, N329, N256);
and AND3 (N580, N575, N97, N65);
not NOT1 (N581, N578);
xor XOR2 (N582, N566, N280);
buf BUF1 (N583, N570);
xor XOR2 (N584, N582, N540);
not NOT1 (N585, N580);
or OR2 (N586, N573, N492);
and AND2 (N587, N581, N203);
buf BUF1 (N588, N574);
nand NAND2 (N589, N576, N142);
buf BUF1 (N590, N588);
and AND4 (N591, N590, N403, N411, N478);
and AND3 (N592, N591, N232, N242);
nor NOR4 (N593, N577, N529, N253, N331);
or OR4 (N594, N585, N362, N106, N449);
nor NOR2 (N595, N571, N536);
nand NAND3 (N596, N579, N202, N169);
nand NAND2 (N597, N594, N72);
buf BUF1 (N598, N595);
and AND4 (N599, N593, N73, N572, N70);
and AND4 (N600, N598, N324, N480, N478);
not NOT1 (N601, N584);
or OR4 (N602, N596, N133, N75, N450);
buf BUF1 (N603, N597);
and AND2 (N604, N592, N360);
or OR4 (N605, N601, N195, N532, N114);
xor XOR2 (N606, N589, N245);
not NOT1 (N607, N604);
not NOT1 (N608, N599);
nand NAND3 (N609, N602, N271, N411);
nand NAND2 (N610, N607, N9);
xor XOR2 (N611, N600, N196);
xor XOR2 (N612, N603, N399);
or OR4 (N613, N606, N117, N368, N171);
not NOT1 (N614, N605);
buf BUF1 (N615, N613);
xor XOR2 (N616, N614, N66);
not NOT1 (N617, N587);
nand NAND2 (N618, N609, N523);
or OR2 (N619, N610, N203);
nand NAND4 (N620, N608, N325, N28, N375);
buf BUF1 (N621, N586);
not NOT1 (N622, N618);
not NOT1 (N623, N611);
not NOT1 (N624, N622);
not NOT1 (N625, N624);
xor XOR2 (N626, N620, N40);
nand NAND2 (N627, N626, N228);
xor XOR2 (N628, N617, N5);
or OR4 (N629, N628, N467, N400, N369);
buf BUF1 (N630, N621);
not NOT1 (N631, N616);
buf BUF1 (N632, N615);
xor XOR2 (N633, N619, N178);
buf BUF1 (N634, N625);
and AND3 (N635, N612, N128, N348);
buf BUF1 (N636, N631);
buf BUF1 (N637, N635);
not NOT1 (N638, N630);
xor XOR2 (N639, N634, N268);
and AND2 (N640, N623, N495);
nand NAND3 (N641, N636, N398, N35);
or OR2 (N642, N637, N418);
and AND3 (N643, N632, N199, N78);
or OR3 (N644, N642, N66, N156);
nor NOR3 (N645, N633, N608, N394);
nor NOR4 (N646, N629, N276, N75, N3);
and AND3 (N647, N641, N462, N396);
nand NAND4 (N648, N638, N100, N270, N281);
and AND3 (N649, N643, N96, N184);
or OR3 (N650, N648, N532, N363);
xor XOR2 (N651, N645, N285);
or OR2 (N652, N640, N303);
nand NAND3 (N653, N583, N1, N451);
buf BUF1 (N654, N639);
or OR2 (N655, N651, N305);
nor NOR4 (N656, N646, N364, N56, N38);
and AND2 (N657, N649, N377);
xor XOR2 (N658, N657, N407);
or OR2 (N659, N650, N414);
buf BUF1 (N660, N647);
nand NAND2 (N661, N627, N315);
not NOT1 (N662, N655);
buf BUF1 (N663, N659);
or OR4 (N664, N644, N289, N24, N319);
not NOT1 (N665, N656);
not NOT1 (N666, N658);
and AND3 (N667, N652, N440, N41);
xor XOR2 (N668, N666, N602);
not NOT1 (N669, N653);
and AND3 (N670, N669, N616, N389);
and AND2 (N671, N668, N569);
not NOT1 (N672, N663);
not NOT1 (N673, N660);
not NOT1 (N674, N672);
buf BUF1 (N675, N654);
not NOT1 (N676, N661);
or OR4 (N677, N676, N302, N354, N179);
not NOT1 (N678, N667);
not NOT1 (N679, N670);
nand NAND2 (N680, N679, N558);
nand NAND2 (N681, N678, N358);
and AND2 (N682, N671, N183);
nand NAND2 (N683, N680, N661);
nor NOR3 (N684, N665, N426, N294);
xor XOR2 (N685, N673, N566);
not NOT1 (N686, N682);
nor NOR2 (N687, N684, N398);
xor XOR2 (N688, N677, N129);
xor XOR2 (N689, N688, N360);
or OR4 (N690, N687, N88, N448, N197);
and AND2 (N691, N675, N3);
and AND4 (N692, N683, N34, N626, N487);
or OR3 (N693, N681, N404, N8);
buf BUF1 (N694, N689);
nand NAND2 (N695, N674, N67);
xor XOR2 (N696, N685, N573);
nand NAND2 (N697, N690, N643);
not NOT1 (N698, N691);
not NOT1 (N699, N664);
and AND3 (N700, N699, N633, N215);
xor XOR2 (N701, N696, N612);
buf BUF1 (N702, N695);
not NOT1 (N703, N702);
not NOT1 (N704, N701);
or OR3 (N705, N694, N140, N288);
or OR2 (N706, N662, N392);
and AND2 (N707, N693, N295);
or OR4 (N708, N706, N307, N296, N36);
nand NAND2 (N709, N705, N279);
nand NAND2 (N710, N704, N673);
nand NAND3 (N711, N709, N617, N434);
xor XOR2 (N712, N710, N199);
nand NAND2 (N713, N700, N706);
nand NAND4 (N714, N713, N182, N42, N533);
nor NOR2 (N715, N686, N530);
and AND3 (N716, N711, N37, N596);
xor XOR2 (N717, N714, N198);
nand NAND4 (N718, N707, N82, N499, N643);
or OR3 (N719, N716, N308, N291);
not NOT1 (N720, N719);
and AND2 (N721, N717, N325);
buf BUF1 (N722, N715);
and AND2 (N723, N712, N454);
or OR2 (N724, N718, N25);
xor XOR2 (N725, N724, N679);
xor XOR2 (N726, N708, N160);
xor XOR2 (N727, N697, N131);
nor NOR4 (N728, N726, N626, N106, N505);
nand NAND4 (N729, N703, N506, N505, N295);
not NOT1 (N730, N729);
or OR4 (N731, N727, N580, N60, N421);
nor NOR3 (N732, N728, N95, N148);
xor XOR2 (N733, N732, N482);
nand NAND3 (N734, N722, N319, N364);
xor XOR2 (N735, N698, N281);
or OR2 (N736, N692, N581);
or OR2 (N737, N720, N703);
buf BUF1 (N738, N723);
nand NAND2 (N739, N738, N5);
and AND2 (N740, N721, N119);
xor XOR2 (N741, N725, N663);
buf BUF1 (N742, N740);
not NOT1 (N743, N737);
xor XOR2 (N744, N730, N598);
nand NAND4 (N745, N731, N136, N256, N144);
not NOT1 (N746, N742);
or OR3 (N747, N733, N42, N470);
or OR4 (N748, N745, N642, N642, N612);
xor XOR2 (N749, N736, N153);
buf BUF1 (N750, N744);
nand NAND4 (N751, N735, N470, N225, N117);
buf BUF1 (N752, N743);
xor XOR2 (N753, N739, N504);
or OR2 (N754, N752, N304);
xor XOR2 (N755, N748, N590);
nand NAND4 (N756, N746, N240, N727, N220);
nand NAND3 (N757, N755, N632, N387);
nand NAND3 (N758, N754, N103, N229);
nor NOR3 (N759, N741, N141, N241);
and AND4 (N760, N747, N671, N602, N431);
not NOT1 (N761, N758);
xor XOR2 (N762, N734, N408);
nor NOR3 (N763, N759, N699, N695);
or OR2 (N764, N761, N2);
not NOT1 (N765, N749);
xor XOR2 (N766, N753, N122);
or OR2 (N767, N766, N696);
and AND3 (N768, N751, N503, N162);
or OR2 (N769, N767, N439);
nor NOR2 (N770, N769, N198);
or OR4 (N771, N762, N724, N33, N376);
nor NOR4 (N772, N750, N39, N561, N572);
or OR4 (N773, N771, N214, N224, N324);
buf BUF1 (N774, N757);
or OR2 (N775, N773, N29);
not NOT1 (N776, N774);
buf BUF1 (N777, N770);
xor XOR2 (N778, N760, N540);
or OR3 (N779, N763, N16, N258);
xor XOR2 (N780, N764, N96);
xor XOR2 (N781, N779, N564);
xor XOR2 (N782, N781, N309);
and AND2 (N783, N772, N486);
and AND3 (N784, N775, N481, N297);
not NOT1 (N785, N782);
nand NAND3 (N786, N756, N312, N427);
nor NOR3 (N787, N777, N88, N180);
not NOT1 (N788, N778);
nand NAND4 (N789, N788, N557, N659, N276);
nand NAND3 (N790, N784, N718, N298);
buf BUF1 (N791, N776);
or OR3 (N792, N785, N548, N778);
buf BUF1 (N793, N780);
or OR3 (N794, N791, N585, N463);
xor XOR2 (N795, N787, N719);
and AND2 (N796, N765, N251);
nor NOR2 (N797, N796, N757);
or OR4 (N798, N789, N585, N524, N258);
not NOT1 (N799, N768);
xor XOR2 (N800, N797, N350);
nor NOR2 (N801, N800, N483);
xor XOR2 (N802, N795, N113);
xor XOR2 (N803, N802, N13);
or OR4 (N804, N798, N661, N102, N81);
not NOT1 (N805, N804);
or OR4 (N806, N799, N479, N707, N804);
nand NAND4 (N807, N792, N627, N491, N684);
and AND3 (N808, N783, N152, N281);
and AND4 (N809, N790, N206, N762, N194);
nand NAND4 (N810, N794, N642, N160, N24);
buf BUF1 (N811, N807);
xor XOR2 (N812, N809, N318);
nor NOR4 (N813, N786, N362, N217, N235);
xor XOR2 (N814, N793, N133);
buf BUF1 (N815, N814);
or OR2 (N816, N808, N697);
xor XOR2 (N817, N816, N468);
not NOT1 (N818, N803);
not NOT1 (N819, N811);
not NOT1 (N820, N818);
not NOT1 (N821, N812);
nand NAND3 (N822, N819, N750, N779);
nand NAND3 (N823, N805, N370, N744);
buf BUF1 (N824, N813);
and AND3 (N825, N820, N484, N648);
nor NOR3 (N826, N810, N105, N2);
nor NOR4 (N827, N815, N732, N232, N820);
xor XOR2 (N828, N824, N630);
buf BUF1 (N829, N822);
xor XOR2 (N830, N828, N291);
nand NAND4 (N831, N829, N683, N813, N640);
xor XOR2 (N832, N801, N514);
buf BUF1 (N833, N825);
buf BUF1 (N834, N826);
buf BUF1 (N835, N821);
and AND3 (N836, N835, N632, N341);
nor NOR3 (N837, N823, N430, N133);
and AND2 (N838, N830, N312);
buf BUF1 (N839, N806);
nand NAND3 (N840, N839, N397, N550);
not NOT1 (N841, N834);
nand NAND2 (N842, N836, N168);
not NOT1 (N843, N837);
nor NOR4 (N844, N843, N406, N496, N672);
xor XOR2 (N845, N817, N799);
and AND2 (N846, N840, N91);
or OR3 (N847, N832, N806, N135);
and AND4 (N848, N846, N273, N679, N211);
nand NAND3 (N849, N844, N487, N104);
xor XOR2 (N850, N833, N13);
nor NOR3 (N851, N847, N569, N806);
nor NOR2 (N852, N851, N296);
xor XOR2 (N853, N845, N320);
and AND4 (N854, N853, N326, N142, N605);
xor XOR2 (N855, N841, N634);
xor XOR2 (N856, N827, N432);
and AND3 (N857, N849, N576, N590);
nor NOR3 (N858, N838, N583, N117);
not NOT1 (N859, N858);
nor NOR3 (N860, N842, N667, N243);
not NOT1 (N861, N848);
or OR2 (N862, N831, N607);
buf BUF1 (N863, N854);
or OR3 (N864, N852, N623, N562);
not NOT1 (N865, N856);
buf BUF1 (N866, N850);
or OR2 (N867, N860, N236);
nand NAND4 (N868, N865, N594, N613, N404);
and AND3 (N869, N862, N750, N858);
not NOT1 (N870, N864);
or OR2 (N871, N855, N483);
xor XOR2 (N872, N869, N251);
or OR2 (N873, N866, N131);
and AND4 (N874, N871, N180, N853, N687);
buf BUF1 (N875, N861);
xor XOR2 (N876, N863, N32);
nor NOR3 (N877, N876, N79, N76);
and AND4 (N878, N868, N406, N424, N578);
and AND2 (N879, N872, N80);
xor XOR2 (N880, N873, N578);
not NOT1 (N881, N867);
nor NOR3 (N882, N870, N690, N616);
buf BUF1 (N883, N879);
nor NOR4 (N884, N877, N276, N396, N729);
nand NAND2 (N885, N875, N855);
nand NAND4 (N886, N885, N385, N876, N73);
buf BUF1 (N887, N881);
or OR2 (N888, N857, N862);
nor NOR4 (N889, N878, N374, N529, N656);
xor XOR2 (N890, N887, N661);
buf BUF1 (N891, N888);
or OR4 (N892, N891, N823, N60, N63);
nand NAND2 (N893, N880, N142);
buf BUF1 (N894, N893);
nand NAND3 (N895, N883, N520, N316);
nand NAND3 (N896, N892, N742, N444);
nor NOR4 (N897, N894, N149, N666, N705);
nor NOR2 (N898, N886, N817);
or OR2 (N899, N859, N793);
nand NAND4 (N900, N899, N296, N354, N391);
nor NOR2 (N901, N898, N755);
and AND2 (N902, N890, N438);
and AND3 (N903, N901, N396, N674);
xor XOR2 (N904, N897, N553);
not NOT1 (N905, N884);
buf BUF1 (N906, N903);
xor XOR2 (N907, N882, N380);
nor NOR3 (N908, N896, N906, N628);
nand NAND2 (N909, N510, N679);
buf BUF1 (N910, N905);
not NOT1 (N911, N902);
nor NOR2 (N912, N889, N614);
nand NAND2 (N913, N907, N539);
or OR2 (N914, N909, N583);
or OR2 (N915, N900, N570);
nor NOR2 (N916, N904, N212);
nor NOR2 (N917, N914, N771);
not NOT1 (N918, N910);
and AND4 (N919, N918, N160, N247, N613);
xor XOR2 (N920, N895, N906);
nand NAND3 (N921, N874, N562, N185);
and AND3 (N922, N912, N302, N708);
endmodule