// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N2510,N2497,N2504,N2517,N2515,N2512,N2513,N2503,N2516,N2518;

nand NAND4 (N19, N9, N9, N5, N11);
buf BUF1 (N20, N9);
not NOT1 (N21, N15);
buf BUF1 (N22, N10);
nor NOR2 (N23, N13, N6);
nand NAND4 (N24, N2, N10, N12, N6);
buf BUF1 (N25, N14);
and AND2 (N26, N16, N12);
and AND3 (N27, N25, N21, N22);
not NOT1 (N28, N16);
not NOT1 (N29, N13);
not NOT1 (N30, N23);
nor NOR4 (N31, N15, N13, N27, N18);
not NOT1 (N32, N8);
and AND3 (N33, N29, N2, N4);
buf BUF1 (N34, N31);
xor XOR2 (N35, N25, N23);
nor NOR4 (N36, N33, N34, N9, N34);
buf BUF1 (N37, N21);
and AND2 (N38, N26, N37);
nand NAND2 (N39, N35, N6);
nor NOR4 (N40, N34, N26, N22, N16);
xor XOR2 (N41, N40, N1);
nor NOR3 (N42, N19, N29, N4);
and AND4 (N43, N42, N3, N24, N32);
xor XOR2 (N44, N6, N4);
nand NAND2 (N45, N9, N32);
and AND2 (N46, N38, N6);
nor NOR4 (N47, N36, N21, N3, N34);
or OR4 (N48, N47, N25, N28, N14);
xor XOR2 (N49, N12, N34);
nor NOR2 (N50, N45, N44);
and AND4 (N51, N49, N15, N50, N3);
or OR2 (N52, N17, N36);
and AND3 (N53, N15, N31, N39);
buf BUF1 (N54, N29);
nor NOR4 (N55, N54, N17, N10, N4);
xor XOR2 (N56, N46, N30);
nand NAND4 (N57, N39, N33, N48, N21);
not NOT1 (N58, N36);
buf BUF1 (N59, N41);
and AND3 (N60, N55, N44, N41);
xor XOR2 (N61, N60, N10);
nand NAND2 (N62, N61, N35);
nor NOR3 (N63, N59, N15, N23);
buf BUF1 (N64, N20);
or OR2 (N65, N57, N52);
not NOT1 (N66, N64);
nand NAND2 (N67, N41, N33);
nand NAND3 (N68, N51, N67, N6);
not NOT1 (N69, N12);
and AND3 (N70, N63, N65, N34);
buf BUF1 (N71, N10);
xor XOR2 (N72, N71, N2);
nand NAND3 (N73, N72, N19, N57);
xor XOR2 (N74, N43, N14);
and AND3 (N75, N68, N21, N44);
buf BUF1 (N76, N70);
and AND3 (N77, N62, N9, N71);
xor XOR2 (N78, N74, N14);
buf BUF1 (N79, N53);
buf BUF1 (N80, N77);
or OR4 (N81, N80, N59, N73, N35);
and AND4 (N82, N28, N21, N45, N14);
buf BUF1 (N83, N66);
nor NOR4 (N84, N56, N64, N26, N66);
nand NAND3 (N85, N69, N59, N77);
and AND3 (N86, N78, N43, N23);
nand NAND2 (N87, N84, N30);
xor XOR2 (N88, N82, N31);
xor XOR2 (N89, N76, N50);
not NOT1 (N90, N88);
nor NOR2 (N91, N90, N90);
buf BUF1 (N92, N85);
buf BUF1 (N93, N89);
not NOT1 (N94, N83);
and AND2 (N95, N92, N32);
not NOT1 (N96, N81);
buf BUF1 (N97, N79);
nor NOR2 (N98, N94, N39);
buf BUF1 (N99, N75);
or OR2 (N100, N93, N12);
or OR4 (N101, N91, N48, N75, N26);
or OR4 (N102, N95, N89, N73, N8);
nor NOR2 (N103, N58, N31);
or OR3 (N104, N102, N75, N49);
buf BUF1 (N105, N104);
nor NOR4 (N106, N103, N14, N15, N86);
xor XOR2 (N107, N79, N68);
buf BUF1 (N108, N97);
buf BUF1 (N109, N108);
buf BUF1 (N110, N98);
and AND3 (N111, N110, N105, N60);
nand NAND3 (N112, N3, N72, N98);
or OR4 (N113, N111, N65, N11, N96);
or OR4 (N114, N71, N110, N66, N42);
xor XOR2 (N115, N107, N72);
buf BUF1 (N116, N109);
xor XOR2 (N117, N114, N22);
xor XOR2 (N118, N112, N53);
and AND4 (N119, N113, N62, N35, N99);
buf BUF1 (N120, N57);
and AND3 (N121, N116, N7, N99);
nor NOR3 (N122, N118, N89, N18);
not NOT1 (N123, N100);
not NOT1 (N124, N122);
xor XOR2 (N125, N87, N32);
and AND3 (N126, N123, N111, N106);
not NOT1 (N127, N118);
nand NAND2 (N128, N127, N84);
or OR4 (N129, N115, N22, N47, N83);
buf BUF1 (N130, N119);
nor NOR2 (N131, N129, N81);
buf BUF1 (N132, N117);
nor NOR2 (N133, N121, N50);
and AND4 (N134, N133, N55, N10, N20);
not NOT1 (N135, N130);
nor NOR4 (N136, N101, N61, N61, N52);
and AND4 (N137, N134, N80, N94, N93);
not NOT1 (N138, N131);
and AND3 (N139, N138, N29, N68);
or OR3 (N140, N135, N105, N135);
nor NOR4 (N141, N124, N39, N91, N107);
and AND3 (N142, N137, N17, N120);
or OR3 (N143, N55, N3, N48);
xor XOR2 (N144, N132, N28);
and AND3 (N145, N141, N126, N62);
or OR3 (N146, N50, N111, N61);
not NOT1 (N147, N136);
nand NAND2 (N148, N145, N96);
nand NAND4 (N149, N125, N140, N19, N86);
buf BUF1 (N150, N145);
xor XOR2 (N151, N143, N150);
buf BUF1 (N152, N13);
buf BUF1 (N153, N142);
not NOT1 (N154, N128);
xor XOR2 (N155, N147, N153);
nand NAND4 (N156, N65, N139, N7, N125);
xor XOR2 (N157, N145, N150);
nor NOR3 (N158, N144, N140, N9);
xor XOR2 (N159, N154, N90);
nor NOR3 (N160, N151, N56, N112);
nand NAND3 (N161, N159, N146, N66);
and AND2 (N162, N103, N150);
or OR4 (N163, N155, N72, N38, N28);
xor XOR2 (N164, N157, N104);
nand NAND2 (N165, N164, N81);
nand NAND4 (N166, N156, N140, N44, N9);
not NOT1 (N167, N163);
buf BUF1 (N168, N149);
and AND3 (N169, N152, N47, N59);
xor XOR2 (N170, N169, N54);
xor XOR2 (N171, N165, N12);
xor XOR2 (N172, N168, N60);
buf BUF1 (N173, N170);
not NOT1 (N174, N173);
or OR3 (N175, N171, N82, N98);
nor NOR2 (N176, N166, N72);
buf BUF1 (N177, N175);
buf BUF1 (N178, N148);
and AND3 (N179, N160, N135, N90);
or OR4 (N180, N158, N103, N128, N22);
not NOT1 (N181, N180);
xor XOR2 (N182, N162, N107);
nand NAND2 (N183, N172, N114);
xor XOR2 (N184, N174, N111);
or OR4 (N185, N184, N55, N37, N167);
nor NOR2 (N186, N71, N66);
buf BUF1 (N187, N176);
or OR3 (N188, N177, N121, N151);
buf BUF1 (N189, N187);
nand NAND4 (N190, N178, N36, N148, N163);
nor NOR4 (N191, N179, N118, N60, N23);
not NOT1 (N192, N185);
or OR3 (N193, N192, N174, N1);
nor NOR3 (N194, N193, N91, N124);
and AND3 (N195, N189, N161, N165);
nor NOR3 (N196, N28, N31, N74);
not NOT1 (N197, N188);
nor NOR2 (N198, N196, N83);
and AND4 (N199, N183, N32, N168, N54);
xor XOR2 (N200, N195, N37);
buf BUF1 (N201, N200);
and AND2 (N202, N199, N13);
or OR3 (N203, N198, N54, N53);
buf BUF1 (N204, N203);
or OR3 (N205, N190, N202, N83);
xor XOR2 (N206, N67, N51);
and AND3 (N207, N194, N167, N5);
nor NOR4 (N208, N207, N52, N27, N112);
xor XOR2 (N209, N204, N126);
nand NAND4 (N210, N201, N91, N120, N16);
xor XOR2 (N211, N186, N158);
or OR3 (N212, N209, N205, N167);
not NOT1 (N213, N144);
and AND3 (N214, N182, N45, N55);
and AND2 (N215, N208, N200);
nand NAND3 (N216, N211, N175, N59);
nand NAND2 (N217, N212, N136);
not NOT1 (N218, N217);
nor NOR2 (N219, N181, N18);
and AND4 (N220, N210, N207, N135, N74);
and AND2 (N221, N214, N76);
not NOT1 (N222, N221);
and AND2 (N223, N218, N153);
nand NAND3 (N224, N197, N105, N110);
nand NAND2 (N225, N223, N2);
or OR4 (N226, N224, N31, N219, N163);
buf BUF1 (N227, N34);
buf BUF1 (N228, N220);
and AND2 (N229, N215, N58);
buf BUF1 (N230, N213);
buf BUF1 (N231, N226);
xor XOR2 (N232, N230, N9);
xor XOR2 (N233, N232, N153);
not NOT1 (N234, N227);
nor NOR2 (N235, N229, N11);
buf BUF1 (N236, N228);
and AND2 (N237, N191, N99);
not NOT1 (N238, N206);
buf BUF1 (N239, N237);
xor XOR2 (N240, N235, N34);
xor XOR2 (N241, N234, N6);
buf BUF1 (N242, N239);
xor XOR2 (N243, N222, N226);
not NOT1 (N244, N236);
and AND2 (N245, N241, N123);
and AND2 (N246, N240, N39);
xor XOR2 (N247, N245, N12);
buf BUF1 (N248, N238);
xor XOR2 (N249, N246, N100);
or OR3 (N250, N243, N196, N203);
not NOT1 (N251, N242);
or OR2 (N252, N247, N119);
nor NOR4 (N253, N216, N37, N198, N82);
or OR3 (N254, N231, N23, N174);
not NOT1 (N255, N225);
buf BUF1 (N256, N254);
nand NAND4 (N257, N252, N78, N247, N44);
nor NOR4 (N258, N251, N50, N65, N143);
not NOT1 (N259, N256);
not NOT1 (N260, N233);
or OR2 (N261, N249, N59);
nand NAND3 (N262, N261, N133, N138);
or OR4 (N263, N258, N233, N170, N48);
nand NAND3 (N264, N248, N188, N27);
buf BUF1 (N265, N255);
nor NOR4 (N266, N244, N203, N164, N236);
not NOT1 (N267, N257);
xor XOR2 (N268, N264, N265);
xor XOR2 (N269, N65, N181);
buf BUF1 (N270, N268);
not NOT1 (N271, N269);
and AND3 (N272, N259, N125, N39);
buf BUF1 (N273, N267);
not NOT1 (N274, N263);
and AND4 (N275, N272, N87, N189, N228);
and AND4 (N276, N266, N222, N109, N245);
or OR3 (N277, N250, N45, N129);
or OR2 (N278, N260, N35);
not NOT1 (N279, N273);
not NOT1 (N280, N279);
buf BUF1 (N281, N280);
buf BUF1 (N282, N275);
or OR3 (N283, N253, N262, N86);
xor XOR2 (N284, N196, N92);
buf BUF1 (N285, N270);
not NOT1 (N286, N281);
not NOT1 (N287, N271);
and AND3 (N288, N282, N149, N13);
and AND4 (N289, N277, N103, N266, N87);
buf BUF1 (N290, N276);
or OR4 (N291, N287, N215, N254, N228);
xor XOR2 (N292, N289, N37);
or OR4 (N293, N285, N147, N239, N210);
and AND3 (N294, N284, N287, N146);
nor NOR4 (N295, N286, N91, N185, N99);
nand NAND4 (N296, N295, N36, N71, N204);
nand NAND3 (N297, N283, N280, N236);
buf BUF1 (N298, N278);
and AND2 (N299, N294, N134);
buf BUF1 (N300, N298);
and AND2 (N301, N300, N264);
or OR4 (N302, N297, N220, N273, N175);
nand NAND3 (N303, N293, N268, N47);
buf BUF1 (N304, N274);
buf BUF1 (N305, N292);
and AND4 (N306, N288, N148, N74, N304);
nand NAND4 (N307, N40, N279, N293, N50);
xor XOR2 (N308, N296, N19);
or OR4 (N309, N302, N68, N140, N297);
or OR4 (N310, N308, N217, N148, N196);
nand NAND3 (N311, N306, N31, N224);
nor NOR4 (N312, N309, N208, N64, N232);
not NOT1 (N313, N301);
and AND4 (N314, N313, N156, N93, N169);
buf BUF1 (N315, N290);
nand NAND2 (N316, N305, N51);
xor XOR2 (N317, N316, N316);
nand NAND3 (N318, N303, N254, N257);
and AND4 (N319, N307, N13, N299, N22);
xor XOR2 (N320, N237, N68);
xor XOR2 (N321, N291, N280);
and AND4 (N322, N312, N172, N9, N92);
xor XOR2 (N323, N310, N214);
xor XOR2 (N324, N315, N314);
or OR4 (N325, N106, N59, N318, N144);
nand NAND3 (N326, N238, N308, N131);
and AND4 (N327, N326, N13, N16, N107);
not NOT1 (N328, N319);
not NOT1 (N329, N322);
xor XOR2 (N330, N324, N160);
nor NOR3 (N331, N328, N274, N189);
buf BUF1 (N332, N311);
not NOT1 (N333, N330);
buf BUF1 (N334, N327);
and AND4 (N335, N329, N280, N95, N271);
buf BUF1 (N336, N335);
and AND3 (N337, N317, N159, N142);
buf BUF1 (N338, N332);
not NOT1 (N339, N331);
or OR2 (N340, N323, N244);
not NOT1 (N341, N334);
buf BUF1 (N342, N336);
nor NOR2 (N343, N341, N85);
and AND4 (N344, N343, N15, N278, N341);
and AND4 (N345, N340, N275, N164, N113);
nand NAND2 (N346, N338, N213);
and AND2 (N347, N344, N343);
and AND2 (N348, N337, N265);
and AND3 (N349, N347, N124, N181);
buf BUF1 (N350, N349);
nor NOR4 (N351, N339, N222, N191, N74);
not NOT1 (N352, N325);
nor NOR3 (N353, N352, N235, N259);
or OR2 (N354, N353, N126);
not NOT1 (N355, N333);
nand NAND2 (N356, N351, N134);
nand NAND2 (N357, N348, N319);
nand NAND3 (N358, N345, N161, N264);
nor NOR4 (N359, N342, N180, N317, N30);
xor XOR2 (N360, N320, N89);
buf BUF1 (N361, N358);
nand NAND2 (N362, N359, N186);
and AND3 (N363, N354, N243, N239);
not NOT1 (N364, N356);
not NOT1 (N365, N321);
and AND4 (N366, N361, N157, N89, N347);
or OR4 (N367, N355, N293, N21, N300);
nand NAND2 (N368, N350, N227);
not NOT1 (N369, N364);
xor XOR2 (N370, N365, N148);
not NOT1 (N371, N357);
nand NAND2 (N372, N367, N63);
xor XOR2 (N373, N369, N76);
nand NAND2 (N374, N368, N9);
or OR4 (N375, N360, N125, N99, N195);
nor NOR2 (N376, N374, N221);
xor XOR2 (N377, N373, N354);
buf BUF1 (N378, N371);
xor XOR2 (N379, N362, N80);
or OR3 (N380, N370, N302, N333);
nand NAND4 (N381, N376, N142, N3, N168);
xor XOR2 (N382, N379, N160);
nor NOR3 (N383, N381, N281, N312);
and AND3 (N384, N383, N267, N97);
not NOT1 (N385, N380);
nor NOR2 (N386, N382, N356);
not NOT1 (N387, N366);
or OR4 (N388, N375, N379, N123, N322);
nor NOR4 (N389, N346, N55, N235, N70);
not NOT1 (N390, N385);
nor NOR4 (N391, N384, N119, N340, N269);
not NOT1 (N392, N390);
or OR2 (N393, N386, N226);
not NOT1 (N394, N391);
buf BUF1 (N395, N392);
xor XOR2 (N396, N387, N228);
buf BUF1 (N397, N393);
buf BUF1 (N398, N397);
xor XOR2 (N399, N372, N184);
not NOT1 (N400, N398);
not NOT1 (N401, N377);
nand NAND4 (N402, N400, N311, N115, N364);
and AND3 (N403, N395, N365, N77);
or OR2 (N404, N363, N147);
xor XOR2 (N405, N388, N2);
buf BUF1 (N406, N404);
nor NOR4 (N407, N406, N95, N80, N6);
nor NOR3 (N408, N402, N365, N131);
or OR4 (N409, N399, N127, N231, N25);
xor XOR2 (N410, N394, N269);
xor XOR2 (N411, N407, N282);
not NOT1 (N412, N410);
nand NAND2 (N413, N412, N316);
xor XOR2 (N414, N389, N387);
and AND3 (N415, N413, N176, N13);
nor NOR2 (N416, N396, N125);
nand NAND4 (N417, N403, N384, N95, N309);
xor XOR2 (N418, N415, N143);
not NOT1 (N419, N401);
or OR2 (N420, N405, N137);
and AND2 (N421, N419, N34);
or OR3 (N422, N409, N371, N358);
nand NAND3 (N423, N417, N110, N60);
buf BUF1 (N424, N420);
and AND3 (N425, N418, N328, N401);
or OR4 (N426, N423, N216, N315, N59);
nand NAND2 (N427, N408, N426);
xor XOR2 (N428, N266, N186);
buf BUF1 (N429, N427);
and AND4 (N430, N414, N10, N177, N122);
nor NOR3 (N431, N425, N285, N163);
buf BUF1 (N432, N422);
or OR3 (N433, N411, N369, N304);
xor XOR2 (N434, N429, N253);
buf BUF1 (N435, N378);
nand NAND2 (N436, N430, N270);
not NOT1 (N437, N435);
xor XOR2 (N438, N421, N298);
xor XOR2 (N439, N431, N25);
and AND3 (N440, N437, N147, N161);
and AND4 (N441, N428, N435, N390, N432);
xor XOR2 (N442, N22, N132);
nand NAND2 (N443, N441, N76);
and AND3 (N444, N442, N434, N281);
nor NOR3 (N445, N346, N398, N288);
nand NAND4 (N446, N440, N429, N167, N36);
buf BUF1 (N447, N416);
not NOT1 (N448, N438);
and AND3 (N449, N439, N209, N309);
or OR2 (N450, N443, N204);
nand NAND3 (N451, N449, N373, N375);
nor NOR3 (N452, N444, N294, N256);
xor XOR2 (N453, N436, N73);
and AND3 (N454, N446, N11, N422);
buf BUF1 (N455, N452);
not NOT1 (N456, N447);
nor NOR2 (N457, N450, N92);
nand NAND4 (N458, N454, N279, N341, N413);
and AND3 (N459, N433, N420, N121);
or OR3 (N460, N458, N175, N443);
xor XOR2 (N461, N457, N393);
xor XOR2 (N462, N461, N234);
nand NAND3 (N463, N455, N418, N76);
nor NOR4 (N464, N456, N376, N393, N272);
not NOT1 (N465, N460);
not NOT1 (N466, N465);
xor XOR2 (N467, N463, N22);
nor NOR2 (N468, N467, N213);
nand NAND3 (N469, N424, N141, N374);
nand NAND2 (N470, N451, N277);
or OR2 (N471, N469, N43);
buf BUF1 (N472, N448);
nor NOR2 (N473, N468, N449);
and AND3 (N474, N466, N166, N456);
and AND3 (N475, N473, N318, N20);
xor XOR2 (N476, N470, N395);
nor NOR3 (N477, N475, N375, N288);
buf BUF1 (N478, N453);
or OR3 (N479, N464, N163, N392);
nor NOR3 (N480, N462, N300, N348);
nand NAND3 (N481, N477, N44, N420);
nor NOR4 (N482, N481, N395, N367, N458);
xor XOR2 (N483, N474, N196);
buf BUF1 (N484, N479);
nand NAND4 (N485, N483, N244, N380, N316);
not NOT1 (N486, N445);
or OR3 (N487, N486, N213, N250);
nor NOR4 (N488, N480, N323, N43, N282);
xor XOR2 (N489, N472, N136);
xor XOR2 (N490, N471, N400);
nor NOR3 (N491, N485, N361, N265);
xor XOR2 (N492, N482, N25);
nor NOR4 (N493, N487, N353, N313, N73);
or OR2 (N494, N476, N135);
not NOT1 (N495, N484);
nand NAND2 (N496, N491, N50);
buf BUF1 (N497, N494);
buf BUF1 (N498, N496);
or OR3 (N499, N492, N126, N62);
xor XOR2 (N500, N499, N397);
xor XOR2 (N501, N493, N308);
buf BUF1 (N502, N500);
or OR4 (N503, N501, N483, N408, N337);
buf BUF1 (N504, N488);
buf BUF1 (N505, N504);
and AND3 (N506, N478, N320, N107);
not NOT1 (N507, N495);
buf BUF1 (N508, N498);
nand NAND4 (N509, N497, N312, N403, N8);
not NOT1 (N510, N502);
or OR4 (N511, N510, N438, N292, N48);
nand NAND2 (N512, N511, N148);
buf BUF1 (N513, N489);
and AND4 (N514, N506, N78, N100, N26);
and AND4 (N515, N508, N133, N245, N152);
nor NOR2 (N516, N503, N186);
nand NAND4 (N517, N507, N51, N368, N508);
nand NAND3 (N518, N490, N301, N486);
and AND4 (N519, N514, N155, N142, N402);
or OR4 (N520, N519, N221, N242, N12);
not NOT1 (N521, N520);
nand NAND2 (N522, N516, N250);
not NOT1 (N523, N459);
buf BUF1 (N524, N521);
nor NOR4 (N525, N517, N426, N443, N414);
or OR2 (N526, N513, N71);
and AND3 (N527, N525, N101, N327);
or OR2 (N528, N509, N40);
buf BUF1 (N529, N528);
and AND3 (N530, N529, N218, N91);
nand NAND3 (N531, N526, N488, N261);
nor NOR2 (N532, N518, N526);
buf BUF1 (N533, N523);
or OR2 (N534, N533, N5);
not NOT1 (N535, N530);
xor XOR2 (N536, N535, N90);
buf BUF1 (N537, N515);
and AND3 (N538, N536, N230, N38);
and AND4 (N539, N537, N263, N16, N8);
or OR4 (N540, N522, N194, N187, N220);
buf BUF1 (N541, N531);
buf BUF1 (N542, N538);
not NOT1 (N543, N505);
nand NAND2 (N544, N532, N492);
buf BUF1 (N545, N534);
buf BUF1 (N546, N527);
nor NOR3 (N547, N539, N378, N448);
xor XOR2 (N548, N545, N130);
or OR3 (N549, N544, N512, N123);
and AND4 (N550, N329, N143, N433, N69);
and AND3 (N551, N550, N403, N192);
xor XOR2 (N552, N546, N306);
xor XOR2 (N553, N541, N238);
not NOT1 (N554, N549);
buf BUF1 (N555, N543);
xor XOR2 (N556, N542, N502);
nor NOR3 (N557, N551, N305, N241);
buf BUF1 (N558, N547);
nand NAND2 (N559, N540, N90);
nor NOR2 (N560, N559, N109);
or OR4 (N561, N553, N508, N104, N181);
not NOT1 (N562, N524);
and AND2 (N563, N556, N60);
and AND2 (N564, N555, N421);
not NOT1 (N565, N548);
nor NOR3 (N566, N564, N539, N481);
not NOT1 (N567, N558);
and AND3 (N568, N566, N34, N214);
not NOT1 (N569, N568);
nor NOR4 (N570, N552, N313, N171, N541);
and AND2 (N571, N557, N432);
buf BUF1 (N572, N569);
nand NAND3 (N573, N554, N112, N244);
or OR2 (N574, N571, N197);
buf BUF1 (N575, N572);
nand NAND3 (N576, N561, N179, N554);
xor XOR2 (N577, N573, N541);
nor NOR4 (N578, N574, N426, N55, N571);
xor XOR2 (N579, N576, N567);
buf BUF1 (N580, N126);
and AND4 (N581, N570, N187, N226, N59);
and AND3 (N582, N580, N54, N2);
or OR2 (N583, N581, N154);
buf BUF1 (N584, N578);
nor NOR2 (N585, N577, N81);
buf BUF1 (N586, N565);
nor NOR4 (N587, N584, N521, N185, N134);
buf BUF1 (N588, N563);
and AND4 (N589, N560, N113, N260, N223);
xor XOR2 (N590, N582, N180);
nor NOR2 (N591, N579, N203);
nand NAND3 (N592, N588, N545, N85);
not NOT1 (N593, N562);
or OR3 (N594, N591, N221, N303);
buf BUF1 (N595, N586);
or OR3 (N596, N589, N457, N504);
xor XOR2 (N597, N575, N236);
buf BUF1 (N598, N596);
nand NAND3 (N599, N585, N252, N203);
not NOT1 (N600, N593);
nand NAND4 (N601, N600, N472, N233, N195);
not NOT1 (N602, N595);
or OR2 (N603, N590, N516);
or OR4 (N604, N597, N139, N268, N111);
and AND2 (N605, N604, N316);
not NOT1 (N606, N583);
or OR3 (N607, N601, N297, N474);
nor NOR2 (N608, N594, N343);
or OR2 (N609, N599, N557);
or OR2 (N610, N603, N257);
nand NAND3 (N611, N587, N582, N128);
xor XOR2 (N612, N605, N297);
or OR4 (N613, N608, N557, N379, N605);
nor NOR3 (N614, N592, N326, N49);
nor NOR4 (N615, N609, N18, N59, N370);
nand NAND2 (N616, N612, N173);
or OR4 (N617, N610, N236, N570, N313);
nand NAND2 (N618, N602, N131);
not NOT1 (N619, N615);
not NOT1 (N620, N614);
xor XOR2 (N621, N617, N290);
and AND4 (N622, N616, N463, N611, N527);
nand NAND2 (N623, N222, N171);
or OR2 (N624, N620, N471);
and AND3 (N625, N606, N102, N106);
nor NOR4 (N626, N607, N609, N389, N7);
nor NOR3 (N627, N624, N204, N94);
not NOT1 (N628, N622);
and AND4 (N629, N598, N376, N573, N123);
buf BUF1 (N630, N619);
and AND4 (N631, N626, N504, N462, N454);
or OR2 (N632, N628, N601);
xor XOR2 (N633, N632, N116);
xor XOR2 (N634, N623, N6);
and AND4 (N635, N621, N254, N429, N271);
nor NOR2 (N636, N630, N489);
buf BUF1 (N637, N634);
not NOT1 (N638, N613);
nor NOR3 (N639, N631, N119, N441);
and AND2 (N640, N633, N319);
xor XOR2 (N641, N625, N617);
buf BUF1 (N642, N640);
nand NAND4 (N643, N641, N296, N376, N298);
xor XOR2 (N644, N642, N132);
buf BUF1 (N645, N627);
buf BUF1 (N646, N638);
not NOT1 (N647, N645);
or OR4 (N648, N618, N430, N103, N539);
or OR3 (N649, N643, N473, N89);
not NOT1 (N650, N637);
xor XOR2 (N651, N650, N315);
buf BUF1 (N652, N636);
xor XOR2 (N653, N646, N22);
not NOT1 (N654, N635);
nand NAND4 (N655, N651, N578, N652, N197);
buf BUF1 (N656, N577);
and AND3 (N657, N644, N283, N281);
xor XOR2 (N658, N629, N421);
nand NAND4 (N659, N647, N539, N354, N254);
and AND4 (N660, N658, N248, N591, N240);
buf BUF1 (N661, N648);
not NOT1 (N662, N649);
not NOT1 (N663, N661);
or OR3 (N664, N659, N393, N129);
xor XOR2 (N665, N656, N620);
buf BUF1 (N666, N660);
buf BUF1 (N667, N654);
and AND4 (N668, N665, N17, N293, N330);
nand NAND2 (N669, N657, N263);
buf BUF1 (N670, N662);
not NOT1 (N671, N670);
buf BUF1 (N672, N666);
and AND2 (N673, N653, N461);
buf BUF1 (N674, N639);
xor XOR2 (N675, N672, N241);
nand NAND2 (N676, N663, N42);
nor NOR2 (N677, N667, N336);
nor NOR2 (N678, N671, N188);
not NOT1 (N679, N674);
and AND4 (N680, N675, N663, N415, N182);
or OR2 (N681, N677, N97);
nand NAND4 (N682, N668, N96, N274, N146);
xor XOR2 (N683, N669, N120);
not NOT1 (N684, N678);
and AND3 (N685, N681, N375, N432);
xor XOR2 (N686, N676, N309);
and AND4 (N687, N684, N102, N538, N375);
and AND4 (N688, N685, N73, N59, N235);
or OR2 (N689, N686, N602);
and AND2 (N690, N689, N178);
buf BUF1 (N691, N673);
nand NAND3 (N692, N683, N99, N193);
nor NOR4 (N693, N680, N388, N688, N456);
not NOT1 (N694, N249);
xor XOR2 (N695, N692, N225);
and AND4 (N696, N687, N593, N523, N301);
or OR3 (N697, N682, N97, N527);
and AND4 (N698, N691, N16, N34, N656);
and AND3 (N699, N690, N226, N644);
xor XOR2 (N700, N664, N537);
nor NOR2 (N701, N700, N686);
buf BUF1 (N702, N695);
nor NOR2 (N703, N655, N404);
nor NOR3 (N704, N694, N211, N280);
nor NOR3 (N705, N703, N26, N603);
xor XOR2 (N706, N696, N464);
buf BUF1 (N707, N705);
nand NAND3 (N708, N704, N46, N175);
buf BUF1 (N709, N708);
nor NOR2 (N710, N698, N388);
and AND2 (N711, N679, N596);
not NOT1 (N712, N693);
or OR2 (N713, N706, N289);
nor NOR2 (N714, N701, N456);
nand NAND3 (N715, N711, N122, N37);
and AND4 (N716, N707, N359, N558, N307);
nor NOR4 (N717, N715, N579, N568, N171);
or OR3 (N718, N713, N161, N43);
and AND4 (N719, N717, N580, N13, N677);
nand NAND2 (N720, N718, N499);
nand NAND3 (N721, N714, N677, N71);
nand NAND3 (N722, N716, N24, N188);
not NOT1 (N723, N702);
not NOT1 (N724, N723);
nand NAND4 (N725, N722, N521, N289, N79);
nor NOR4 (N726, N710, N123, N407, N58);
xor XOR2 (N727, N697, N460);
nand NAND4 (N728, N724, N396, N114, N268);
not NOT1 (N729, N728);
xor XOR2 (N730, N712, N340);
nor NOR3 (N731, N720, N523, N439);
or OR3 (N732, N726, N711, N153);
xor XOR2 (N733, N709, N188);
nor NOR3 (N734, N725, N732, N65);
and AND2 (N735, N14, N711);
not NOT1 (N736, N733);
xor XOR2 (N737, N727, N386);
buf BUF1 (N738, N731);
and AND3 (N739, N721, N378, N78);
nand NAND4 (N740, N739, N176, N617, N539);
and AND3 (N741, N734, N537, N627);
or OR3 (N742, N729, N534, N643);
xor XOR2 (N743, N742, N653);
or OR3 (N744, N737, N543, N120);
buf BUF1 (N745, N736);
or OR4 (N746, N735, N290, N694, N17);
not NOT1 (N747, N740);
nor NOR2 (N748, N745, N191);
xor XOR2 (N749, N699, N439);
or OR3 (N750, N730, N744, N364);
and AND2 (N751, N5, N248);
not NOT1 (N752, N747);
nand NAND4 (N753, N750, N691, N247, N690);
xor XOR2 (N754, N719, N255);
not NOT1 (N755, N752);
nand NAND3 (N756, N754, N527, N129);
and AND2 (N757, N756, N756);
and AND4 (N758, N753, N616, N344, N577);
not NOT1 (N759, N755);
buf BUF1 (N760, N746);
not NOT1 (N761, N738);
buf BUF1 (N762, N749);
buf BUF1 (N763, N741);
nand NAND4 (N764, N760, N673, N654, N414);
and AND4 (N765, N761, N651, N376, N668);
and AND3 (N766, N762, N337, N724);
nand NAND2 (N767, N748, N130);
nand NAND3 (N768, N743, N198, N363);
xor XOR2 (N769, N766, N267);
not NOT1 (N770, N763);
and AND3 (N771, N765, N88, N151);
buf BUF1 (N772, N770);
not NOT1 (N773, N764);
and AND3 (N774, N768, N668, N369);
not NOT1 (N775, N772);
nand NAND2 (N776, N758, N382);
xor XOR2 (N777, N773, N531);
nand NAND4 (N778, N774, N771, N131, N130);
buf BUF1 (N779, N164);
or OR3 (N780, N776, N346, N413);
nor NOR3 (N781, N780, N690, N419);
buf BUF1 (N782, N767);
or OR3 (N783, N779, N209, N581);
xor XOR2 (N784, N782, N186);
buf BUF1 (N785, N783);
and AND3 (N786, N778, N611, N695);
nor NOR3 (N787, N785, N90, N359);
or OR3 (N788, N777, N541, N55);
not NOT1 (N789, N751);
or OR2 (N790, N784, N347);
not NOT1 (N791, N789);
nor NOR3 (N792, N759, N399, N736);
and AND4 (N793, N757, N174, N110, N65);
and AND2 (N794, N769, N296);
xor XOR2 (N795, N791, N444);
nor NOR4 (N796, N786, N373, N430, N459);
xor XOR2 (N797, N775, N199);
nand NAND3 (N798, N788, N326, N254);
buf BUF1 (N799, N795);
buf BUF1 (N800, N793);
or OR4 (N801, N792, N591, N257, N3);
and AND4 (N802, N781, N330, N171, N725);
buf BUF1 (N803, N790);
nand NAND2 (N804, N787, N206);
xor XOR2 (N805, N803, N462);
nor NOR3 (N806, N801, N469, N490);
not NOT1 (N807, N796);
xor XOR2 (N808, N805, N465);
xor XOR2 (N809, N799, N56);
nor NOR4 (N810, N806, N634, N715, N149);
and AND3 (N811, N809, N702, N187);
nand NAND4 (N812, N808, N706, N574, N216);
nor NOR4 (N813, N811, N747, N314, N548);
not NOT1 (N814, N812);
not NOT1 (N815, N804);
xor XOR2 (N816, N807, N707);
not NOT1 (N817, N810);
not NOT1 (N818, N797);
nand NAND2 (N819, N802, N407);
nand NAND3 (N820, N818, N138, N677);
nand NAND2 (N821, N816, N324);
and AND3 (N822, N813, N389, N58);
or OR4 (N823, N798, N166, N790, N90);
or OR3 (N824, N819, N710, N789);
nor NOR2 (N825, N822, N583);
and AND4 (N826, N815, N323, N202, N550);
nor NOR4 (N827, N800, N437, N774, N583);
xor XOR2 (N828, N794, N252);
xor XOR2 (N829, N825, N340);
nor NOR2 (N830, N817, N362);
not NOT1 (N831, N829);
not NOT1 (N832, N827);
nand NAND4 (N833, N828, N477, N191, N107);
xor XOR2 (N834, N832, N182);
or OR3 (N835, N830, N693, N604);
nand NAND4 (N836, N820, N437, N715, N798);
nor NOR2 (N837, N835, N64);
buf BUF1 (N838, N831);
nand NAND3 (N839, N834, N276, N335);
nor NOR2 (N840, N839, N5);
xor XOR2 (N841, N840, N249);
xor XOR2 (N842, N838, N663);
nand NAND3 (N843, N826, N477, N65);
nand NAND2 (N844, N824, N350);
nand NAND4 (N845, N842, N621, N358, N774);
or OR4 (N846, N823, N662, N477, N570);
nand NAND2 (N847, N845, N519);
xor XOR2 (N848, N846, N548);
nor NOR4 (N849, N843, N808, N434, N475);
and AND2 (N850, N836, N64);
buf BUF1 (N851, N850);
xor XOR2 (N852, N821, N268);
or OR4 (N853, N814, N833, N760, N401);
buf BUF1 (N854, N300);
nor NOR4 (N855, N854, N289, N215, N105);
nand NAND3 (N856, N848, N793, N293);
nor NOR4 (N857, N852, N201, N98, N536);
nor NOR3 (N858, N844, N465, N839);
not NOT1 (N859, N841);
not NOT1 (N860, N857);
and AND4 (N861, N853, N574, N624, N693);
and AND4 (N862, N851, N533, N69, N813);
not NOT1 (N863, N858);
not NOT1 (N864, N849);
nor NOR2 (N865, N856, N210);
nand NAND4 (N866, N847, N700, N82, N554);
or OR4 (N867, N866, N493, N725, N440);
xor XOR2 (N868, N867, N790);
or OR4 (N869, N861, N602, N601, N549);
buf BUF1 (N870, N869);
nand NAND2 (N871, N865, N454);
or OR4 (N872, N859, N268, N311, N548);
nand NAND3 (N873, N837, N14, N602);
nor NOR4 (N874, N871, N153, N351, N174);
and AND2 (N875, N870, N334);
not NOT1 (N876, N855);
not NOT1 (N877, N864);
buf BUF1 (N878, N875);
xor XOR2 (N879, N874, N625);
not NOT1 (N880, N860);
nor NOR4 (N881, N878, N50, N822, N650);
buf BUF1 (N882, N862);
not NOT1 (N883, N879);
xor XOR2 (N884, N881, N252);
nor NOR3 (N885, N868, N555, N44);
nand NAND4 (N886, N883, N417, N823, N450);
xor XOR2 (N887, N882, N105);
nor NOR4 (N888, N876, N770, N359, N724);
xor XOR2 (N889, N863, N349);
buf BUF1 (N890, N880);
and AND2 (N891, N877, N534);
buf BUF1 (N892, N873);
nor NOR3 (N893, N872, N502, N596);
not NOT1 (N894, N888);
or OR4 (N895, N889, N584, N801, N494);
buf BUF1 (N896, N887);
not NOT1 (N897, N891);
nand NAND3 (N898, N897, N680, N37);
nand NAND2 (N899, N895, N71);
and AND4 (N900, N892, N155, N126, N82);
and AND3 (N901, N884, N727, N694);
not NOT1 (N902, N894);
xor XOR2 (N903, N896, N322);
nand NAND2 (N904, N890, N320);
nor NOR4 (N905, N886, N133, N555, N144);
nor NOR2 (N906, N885, N502);
not NOT1 (N907, N893);
or OR4 (N908, N906, N561, N829, N246);
or OR4 (N909, N907, N447, N905, N373);
xor XOR2 (N910, N415, N126);
buf BUF1 (N911, N910);
and AND3 (N912, N901, N15, N16);
buf BUF1 (N913, N912);
or OR3 (N914, N904, N44, N803);
nor NOR3 (N915, N902, N600, N227);
or OR3 (N916, N899, N550, N309);
xor XOR2 (N917, N898, N677);
or OR4 (N918, N915, N118, N550, N40);
xor XOR2 (N919, N918, N662);
xor XOR2 (N920, N913, N684);
and AND4 (N921, N920, N267, N38, N307);
or OR4 (N922, N908, N142, N427, N75);
and AND3 (N923, N909, N578, N5);
and AND3 (N924, N916, N624, N520);
or OR2 (N925, N923, N247);
not NOT1 (N926, N911);
or OR2 (N927, N900, N386);
or OR2 (N928, N917, N240);
nor NOR3 (N929, N922, N476, N16);
buf BUF1 (N930, N921);
or OR2 (N931, N930, N570);
or OR4 (N932, N926, N609, N231, N727);
xor XOR2 (N933, N903, N463);
buf BUF1 (N934, N919);
buf BUF1 (N935, N933);
not NOT1 (N936, N931);
nor NOR2 (N937, N925, N111);
xor XOR2 (N938, N937, N136);
or OR3 (N939, N936, N675, N909);
nor NOR3 (N940, N932, N458, N504);
nor NOR2 (N941, N928, N760);
not NOT1 (N942, N940);
xor XOR2 (N943, N927, N411);
nand NAND2 (N944, N934, N547);
nand NAND3 (N945, N943, N825, N544);
not NOT1 (N946, N944);
nor NOR2 (N947, N914, N102);
and AND3 (N948, N942, N585, N531);
xor XOR2 (N949, N947, N593);
not NOT1 (N950, N939);
and AND3 (N951, N935, N313, N865);
nand NAND3 (N952, N938, N662, N77);
nor NOR3 (N953, N950, N542, N807);
buf BUF1 (N954, N952);
or OR2 (N955, N954, N316);
and AND3 (N956, N948, N353, N610);
not NOT1 (N957, N953);
buf BUF1 (N958, N956);
buf BUF1 (N959, N929);
buf BUF1 (N960, N958);
and AND2 (N961, N949, N672);
or OR3 (N962, N941, N600, N493);
not NOT1 (N963, N924);
buf BUF1 (N964, N963);
buf BUF1 (N965, N951);
nand NAND3 (N966, N945, N755, N108);
nor NOR2 (N967, N955, N912);
or OR4 (N968, N965, N630, N849, N817);
nand NAND3 (N969, N946, N763, N326);
nand NAND3 (N970, N962, N458, N589);
and AND3 (N971, N968, N522, N324);
not NOT1 (N972, N970);
not NOT1 (N973, N972);
not NOT1 (N974, N957);
nand NAND2 (N975, N961, N972);
nor NOR4 (N976, N966, N730, N586, N304);
nand NAND3 (N977, N974, N526, N288);
nor NOR2 (N978, N971, N209);
not NOT1 (N979, N975);
or OR2 (N980, N964, N292);
not NOT1 (N981, N959);
and AND3 (N982, N976, N214, N909);
nor NOR2 (N983, N973, N980);
xor XOR2 (N984, N227, N221);
buf BUF1 (N985, N982);
or OR4 (N986, N977, N791, N222, N144);
and AND3 (N987, N967, N722, N254);
or OR3 (N988, N983, N475, N711);
or OR2 (N989, N985, N898);
nand NAND3 (N990, N984, N260, N278);
or OR2 (N991, N987, N979);
and AND4 (N992, N550, N772, N984, N331);
buf BUF1 (N993, N981);
not NOT1 (N994, N991);
and AND3 (N995, N990, N46, N878);
and AND4 (N996, N969, N152, N193, N478);
and AND2 (N997, N989, N56);
or OR2 (N998, N988, N324);
or OR4 (N999, N992, N574, N41, N893);
xor XOR2 (N1000, N960, N617);
not NOT1 (N1001, N1000);
nand NAND4 (N1002, N998, N778, N383, N839);
and AND3 (N1003, N978, N121, N78);
xor XOR2 (N1004, N1002, N47);
buf BUF1 (N1005, N1004);
not NOT1 (N1006, N999);
nand NAND3 (N1007, N986, N776, N259);
or OR2 (N1008, N996, N819);
buf BUF1 (N1009, N993);
not NOT1 (N1010, N1008);
nand NAND3 (N1011, N997, N252, N790);
not NOT1 (N1012, N1007);
buf BUF1 (N1013, N1012);
nor NOR4 (N1014, N1005, N610, N703, N819);
and AND2 (N1015, N1013, N276);
and AND3 (N1016, N1010, N745, N226);
or OR2 (N1017, N1003, N612);
not NOT1 (N1018, N1016);
nand NAND3 (N1019, N995, N498, N944);
nor NOR2 (N1020, N1018, N502);
and AND2 (N1021, N994, N977);
xor XOR2 (N1022, N1020, N158);
nand NAND3 (N1023, N1009, N353, N241);
nand NAND2 (N1024, N1022, N66);
buf BUF1 (N1025, N1021);
and AND3 (N1026, N1025, N940, N906);
not NOT1 (N1027, N1014);
not NOT1 (N1028, N1011);
or OR2 (N1029, N1017, N668);
nor NOR4 (N1030, N1028, N97, N67, N669);
or OR4 (N1031, N1006, N36, N433, N372);
buf BUF1 (N1032, N1030);
not NOT1 (N1033, N1029);
nor NOR4 (N1034, N1024, N1019, N603, N388);
buf BUF1 (N1035, N554);
xor XOR2 (N1036, N1033, N632);
nor NOR2 (N1037, N1026, N138);
nand NAND2 (N1038, N1037, N167);
nand NAND4 (N1039, N1031, N339, N107, N856);
xor XOR2 (N1040, N1038, N706);
or OR2 (N1041, N1032, N955);
nor NOR2 (N1042, N1023, N621);
and AND3 (N1043, N1036, N390, N976);
and AND4 (N1044, N1015, N671, N780, N527);
nand NAND3 (N1045, N1044, N788, N1040);
and AND2 (N1046, N589, N820);
nor NOR4 (N1047, N1042, N479, N298, N845);
nand NAND3 (N1048, N1039, N1036, N335);
nand NAND4 (N1049, N1001, N568, N36, N990);
nand NAND2 (N1050, N1049, N726);
xor XOR2 (N1051, N1043, N687);
not NOT1 (N1052, N1034);
not NOT1 (N1053, N1041);
buf BUF1 (N1054, N1053);
and AND2 (N1055, N1047, N1005);
not NOT1 (N1056, N1052);
buf BUF1 (N1057, N1055);
not NOT1 (N1058, N1057);
nand NAND3 (N1059, N1056, N328, N667);
buf BUF1 (N1060, N1059);
xor XOR2 (N1061, N1058, N291);
xor XOR2 (N1062, N1050, N1057);
nand NAND2 (N1063, N1061, N381);
nor NOR2 (N1064, N1062, N899);
nand NAND2 (N1065, N1060, N887);
nand NAND3 (N1066, N1063, N621, N964);
buf BUF1 (N1067, N1046);
nand NAND3 (N1068, N1054, N500, N868);
buf BUF1 (N1069, N1035);
nor NOR3 (N1070, N1064, N682, N114);
and AND4 (N1071, N1070, N499, N265, N272);
xor XOR2 (N1072, N1048, N261);
xor XOR2 (N1073, N1066, N671);
buf BUF1 (N1074, N1067);
or OR4 (N1075, N1068, N1024, N899, N699);
buf BUF1 (N1076, N1069);
buf BUF1 (N1077, N1072);
xor XOR2 (N1078, N1074, N497);
nor NOR2 (N1079, N1051, N1);
nor NOR2 (N1080, N1027, N337);
xor XOR2 (N1081, N1076, N943);
and AND2 (N1082, N1081, N263);
buf BUF1 (N1083, N1071);
buf BUF1 (N1084, N1045);
buf BUF1 (N1085, N1082);
buf BUF1 (N1086, N1080);
xor XOR2 (N1087, N1078, N1034);
or OR3 (N1088, N1075, N331, N366);
or OR4 (N1089, N1065, N486, N924, N358);
nor NOR2 (N1090, N1084, N959);
buf BUF1 (N1091, N1090);
buf BUF1 (N1092, N1073);
not NOT1 (N1093, N1089);
or OR2 (N1094, N1086, N650);
nor NOR3 (N1095, N1088, N652, N1052);
xor XOR2 (N1096, N1095, N783);
nor NOR2 (N1097, N1094, N207);
buf BUF1 (N1098, N1097);
buf BUF1 (N1099, N1077);
buf BUF1 (N1100, N1092);
not NOT1 (N1101, N1085);
or OR2 (N1102, N1079, N457);
not NOT1 (N1103, N1099);
nand NAND3 (N1104, N1100, N317, N771);
xor XOR2 (N1105, N1101, N493);
nand NAND2 (N1106, N1104, N50);
xor XOR2 (N1107, N1093, N197);
buf BUF1 (N1108, N1098);
not NOT1 (N1109, N1096);
and AND3 (N1110, N1091, N997, N650);
nand NAND4 (N1111, N1105, N986, N1044, N1064);
not NOT1 (N1112, N1102);
and AND4 (N1113, N1083, N748, N1002, N882);
or OR4 (N1114, N1110, N733, N298, N782);
or OR4 (N1115, N1113, N625, N578, N325);
or OR4 (N1116, N1109, N621, N357, N537);
nand NAND3 (N1117, N1106, N317, N908);
or OR2 (N1118, N1114, N699);
xor XOR2 (N1119, N1115, N210);
not NOT1 (N1120, N1119);
buf BUF1 (N1121, N1108);
and AND3 (N1122, N1116, N478, N66);
nor NOR2 (N1123, N1121, N987);
buf BUF1 (N1124, N1107);
and AND3 (N1125, N1123, N1053, N354);
nand NAND2 (N1126, N1124, N84);
not NOT1 (N1127, N1125);
xor XOR2 (N1128, N1087, N239);
and AND3 (N1129, N1112, N902, N984);
nand NAND2 (N1130, N1122, N747);
nor NOR3 (N1131, N1120, N764, N456);
nor NOR4 (N1132, N1118, N528, N50, N452);
or OR3 (N1133, N1129, N164, N324);
nor NOR2 (N1134, N1132, N973);
buf BUF1 (N1135, N1111);
buf BUF1 (N1136, N1117);
xor XOR2 (N1137, N1127, N755);
and AND2 (N1138, N1128, N787);
not NOT1 (N1139, N1103);
and AND2 (N1140, N1130, N452);
or OR3 (N1141, N1137, N481, N398);
nor NOR2 (N1142, N1131, N660);
nor NOR2 (N1143, N1136, N1003);
or OR2 (N1144, N1133, N712);
and AND2 (N1145, N1140, N61);
or OR3 (N1146, N1145, N974, N65);
and AND2 (N1147, N1139, N192);
nand NAND2 (N1148, N1141, N166);
xor XOR2 (N1149, N1134, N292);
nor NOR4 (N1150, N1149, N867, N973, N509);
nand NAND3 (N1151, N1148, N597, N90);
buf BUF1 (N1152, N1126);
and AND4 (N1153, N1150, N420, N1022, N853);
nor NOR2 (N1154, N1146, N477);
nor NOR2 (N1155, N1135, N358);
or OR2 (N1156, N1143, N495);
not NOT1 (N1157, N1152);
buf BUF1 (N1158, N1144);
not NOT1 (N1159, N1142);
nand NAND2 (N1160, N1158, N216);
and AND3 (N1161, N1160, N154, N515);
or OR2 (N1162, N1153, N1148);
buf BUF1 (N1163, N1156);
and AND3 (N1164, N1151, N144, N80);
not NOT1 (N1165, N1162);
buf BUF1 (N1166, N1138);
not NOT1 (N1167, N1165);
nor NOR3 (N1168, N1161, N410, N300);
buf BUF1 (N1169, N1157);
nand NAND2 (N1170, N1164, N986);
buf BUF1 (N1171, N1166);
and AND2 (N1172, N1171, N98);
buf BUF1 (N1173, N1167);
not NOT1 (N1174, N1163);
nor NOR2 (N1175, N1170, N513);
nor NOR3 (N1176, N1173, N342, N672);
nor NOR3 (N1177, N1168, N777, N141);
xor XOR2 (N1178, N1172, N418);
nor NOR3 (N1179, N1154, N4, N1031);
xor XOR2 (N1180, N1178, N55);
nor NOR2 (N1181, N1147, N91);
xor XOR2 (N1182, N1180, N651);
nor NOR4 (N1183, N1179, N423, N1123, N306);
nand NAND4 (N1184, N1183, N1090, N703, N231);
and AND2 (N1185, N1176, N608);
buf BUF1 (N1186, N1155);
buf BUF1 (N1187, N1169);
nand NAND4 (N1188, N1181, N431, N1121, N739);
xor XOR2 (N1189, N1175, N961);
and AND2 (N1190, N1177, N490);
or OR4 (N1191, N1186, N686, N951, N118);
not NOT1 (N1192, N1187);
not NOT1 (N1193, N1190);
and AND2 (N1194, N1188, N1095);
not NOT1 (N1195, N1184);
and AND4 (N1196, N1192, N468, N47, N213);
buf BUF1 (N1197, N1189);
not NOT1 (N1198, N1196);
or OR2 (N1199, N1191, N30);
buf BUF1 (N1200, N1159);
xor XOR2 (N1201, N1199, N1064);
buf BUF1 (N1202, N1195);
nand NAND2 (N1203, N1182, N436);
not NOT1 (N1204, N1185);
nor NOR3 (N1205, N1203, N1054, N1193);
xor XOR2 (N1206, N946, N1088);
and AND2 (N1207, N1204, N889);
or OR2 (N1208, N1197, N476);
buf BUF1 (N1209, N1198);
not NOT1 (N1210, N1201);
not NOT1 (N1211, N1210);
and AND4 (N1212, N1174, N1092, N312, N386);
not NOT1 (N1213, N1205);
nand NAND3 (N1214, N1208, N932, N639);
buf BUF1 (N1215, N1202);
or OR2 (N1216, N1214, N480);
xor XOR2 (N1217, N1215, N682);
or OR3 (N1218, N1217, N1042, N310);
and AND2 (N1219, N1213, N904);
buf BUF1 (N1220, N1207);
nor NOR3 (N1221, N1194, N530, N671);
or OR2 (N1222, N1216, N1060);
nor NOR4 (N1223, N1222, N430, N222, N529);
xor XOR2 (N1224, N1209, N859);
not NOT1 (N1225, N1223);
and AND2 (N1226, N1220, N1187);
or OR2 (N1227, N1211, N365);
or OR3 (N1228, N1224, N6, N824);
xor XOR2 (N1229, N1227, N511);
or OR2 (N1230, N1226, N1005);
nor NOR4 (N1231, N1219, N665, N1039, N531);
not NOT1 (N1232, N1229);
or OR4 (N1233, N1206, N74, N1177, N497);
nor NOR3 (N1234, N1218, N217, N891);
nand NAND4 (N1235, N1221, N930, N1123, N390);
xor XOR2 (N1236, N1212, N73);
nand NAND2 (N1237, N1235, N368);
nand NAND3 (N1238, N1225, N1156, N1153);
nor NOR4 (N1239, N1233, N865, N701, N41);
not NOT1 (N1240, N1232);
xor XOR2 (N1241, N1236, N99);
xor XOR2 (N1242, N1228, N1035);
or OR2 (N1243, N1242, N1051);
xor XOR2 (N1244, N1240, N153);
nor NOR4 (N1245, N1243, N552, N86, N833);
nor NOR2 (N1246, N1244, N744);
nand NAND4 (N1247, N1237, N186, N474, N306);
not NOT1 (N1248, N1241);
nor NOR3 (N1249, N1247, N202, N453);
and AND4 (N1250, N1239, N1000, N887, N591);
buf BUF1 (N1251, N1245);
not NOT1 (N1252, N1200);
xor XOR2 (N1253, N1234, N603);
and AND3 (N1254, N1250, N215, N469);
nand NAND2 (N1255, N1254, N636);
buf BUF1 (N1256, N1246);
and AND4 (N1257, N1230, N914, N1090, N827);
not NOT1 (N1258, N1248);
and AND2 (N1259, N1255, N1);
buf BUF1 (N1260, N1253);
nand NAND3 (N1261, N1249, N809, N499);
not NOT1 (N1262, N1257);
buf BUF1 (N1263, N1259);
buf BUF1 (N1264, N1231);
nor NOR2 (N1265, N1238, N639);
or OR4 (N1266, N1262, N1100, N538, N54);
buf BUF1 (N1267, N1256);
nor NOR2 (N1268, N1267, N624);
or OR4 (N1269, N1252, N684, N403, N854);
not NOT1 (N1270, N1258);
nor NOR4 (N1271, N1265, N51, N891, N15);
or OR2 (N1272, N1268, N790);
nor NOR2 (N1273, N1271, N244);
buf BUF1 (N1274, N1269);
or OR4 (N1275, N1272, N496, N637, N119);
nor NOR3 (N1276, N1273, N604, N178);
not NOT1 (N1277, N1276);
not NOT1 (N1278, N1264);
nand NAND3 (N1279, N1251, N352, N268);
and AND2 (N1280, N1263, N573);
not NOT1 (N1281, N1260);
xor XOR2 (N1282, N1275, N684);
xor XOR2 (N1283, N1282, N173);
or OR4 (N1284, N1266, N117, N177, N994);
or OR3 (N1285, N1281, N984, N927);
nand NAND3 (N1286, N1274, N481, N665);
not NOT1 (N1287, N1270);
not NOT1 (N1288, N1286);
xor XOR2 (N1289, N1283, N432);
xor XOR2 (N1290, N1287, N14);
and AND4 (N1291, N1278, N1148, N305, N1283);
not NOT1 (N1292, N1285);
buf BUF1 (N1293, N1277);
nor NOR3 (N1294, N1290, N866, N255);
buf BUF1 (N1295, N1291);
or OR2 (N1296, N1289, N1136);
or OR4 (N1297, N1296, N469, N1146, N962);
buf BUF1 (N1298, N1284);
nor NOR4 (N1299, N1295, N396, N1105, N1114);
nor NOR4 (N1300, N1297, N889, N1247, N470);
not NOT1 (N1301, N1298);
not NOT1 (N1302, N1301);
not NOT1 (N1303, N1261);
or OR2 (N1304, N1288, N246);
nand NAND3 (N1305, N1280, N80, N328);
xor XOR2 (N1306, N1292, N996);
buf BUF1 (N1307, N1299);
not NOT1 (N1308, N1293);
xor XOR2 (N1309, N1294, N529);
nand NAND4 (N1310, N1304, N1228, N7, N240);
xor XOR2 (N1311, N1300, N124);
and AND4 (N1312, N1307, N847, N1309, N313);
nor NOR4 (N1313, N387, N248, N953, N229);
not NOT1 (N1314, N1312);
xor XOR2 (N1315, N1302, N510);
nor NOR2 (N1316, N1306, N1230);
nand NAND4 (N1317, N1308, N191, N351, N1272);
buf BUF1 (N1318, N1303);
not NOT1 (N1319, N1313);
nand NAND2 (N1320, N1314, N90);
or OR3 (N1321, N1279, N1291, N59);
or OR4 (N1322, N1319, N320, N829, N163);
not NOT1 (N1323, N1310);
nor NOR2 (N1324, N1320, N407);
not NOT1 (N1325, N1324);
xor XOR2 (N1326, N1322, N1316);
not NOT1 (N1327, N728);
nand NAND4 (N1328, N1321, N77, N185, N495);
or OR4 (N1329, N1326, N1195, N912, N1209);
not NOT1 (N1330, N1315);
not NOT1 (N1331, N1305);
or OR2 (N1332, N1323, N283);
nor NOR4 (N1333, N1329, N891, N739, N1000);
xor XOR2 (N1334, N1330, N863);
xor XOR2 (N1335, N1334, N1133);
buf BUF1 (N1336, N1332);
or OR2 (N1337, N1325, N472);
not NOT1 (N1338, N1317);
or OR2 (N1339, N1337, N800);
xor XOR2 (N1340, N1311, N1203);
buf BUF1 (N1341, N1338);
xor XOR2 (N1342, N1335, N805);
xor XOR2 (N1343, N1339, N475);
nor NOR4 (N1344, N1340, N214, N1159, N432);
or OR2 (N1345, N1327, N239);
buf BUF1 (N1346, N1328);
and AND4 (N1347, N1344, N628, N210, N173);
xor XOR2 (N1348, N1341, N268);
or OR4 (N1349, N1331, N1193, N704, N643);
buf BUF1 (N1350, N1346);
nor NOR3 (N1351, N1347, N385, N714);
nand NAND4 (N1352, N1342, N285, N803, N390);
not NOT1 (N1353, N1333);
xor XOR2 (N1354, N1343, N1);
nor NOR4 (N1355, N1351, N756, N390, N1303);
not NOT1 (N1356, N1352);
xor XOR2 (N1357, N1356, N721);
nor NOR2 (N1358, N1357, N649);
nor NOR2 (N1359, N1354, N1094);
not NOT1 (N1360, N1349);
buf BUF1 (N1361, N1345);
or OR2 (N1362, N1353, N457);
or OR4 (N1363, N1336, N989, N1260, N836);
and AND3 (N1364, N1358, N324, N1026);
or OR3 (N1365, N1362, N1330, N819);
xor XOR2 (N1366, N1360, N146);
nor NOR2 (N1367, N1364, N123);
not NOT1 (N1368, N1361);
nor NOR2 (N1369, N1367, N888);
nor NOR2 (N1370, N1348, N233);
nand NAND2 (N1371, N1366, N132);
not NOT1 (N1372, N1359);
or OR2 (N1373, N1370, N1352);
nand NAND3 (N1374, N1363, N1250, N349);
buf BUF1 (N1375, N1374);
not NOT1 (N1376, N1350);
and AND3 (N1377, N1368, N278, N878);
nor NOR4 (N1378, N1371, N1049, N440, N928);
or OR2 (N1379, N1372, N429);
xor XOR2 (N1380, N1377, N131);
buf BUF1 (N1381, N1375);
not NOT1 (N1382, N1381);
xor XOR2 (N1383, N1369, N915);
buf BUF1 (N1384, N1378);
not NOT1 (N1385, N1379);
nand NAND4 (N1386, N1355, N205, N844, N388);
and AND2 (N1387, N1376, N933);
nor NOR2 (N1388, N1387, N744);
or OR2 (N1389, N1384, N1130);
nand NAND4 (N1390, N1373, N48, N717, N113);
and AND4 (N1391, N1365, N1243, N212, N813);
and AND3 (N1392, N1318, N438, N1374);
buf BUF1 (N1393, N1383);
and AND2 (N1394, N1393, N1140);
not NOT1 (N1395, N1386);
nand NAND2 (N1396, N1391, N908);
xor XOR2 (N1397, N1389, N307);
and AND4 (N1398, N1382, N999, N1181, N822);
or OR4 (N1399, N1397, N1007, N305, N616);
nor NOR2 (N1400, N1380, N336);
or OR3 (N1401, N1388, N1390, N484);
or OR4 (N1402, N614, N1120, N428, N1394);
xor XOR2 (N1403, N726, N303);
not NOT1 (N1404, N1392);
and AND3 (N1405, N1401, N1147, N413);
or OR3 (N1406, N1398, N616, N202);
not NOT1 (N1407, N1396);
not NOT1 (N1408, N1406);
and AND2 (N1409, N1407, N1303);
buf BUF1 (N1410, N1395);
buf BUF1 (N1411, N1409);
buf BUF1 (N1412, N1405);
or OR3 (N1413, N1403, N79, N759);
buf BUF1 (N1414, N1412);
buf BUF1 (N1415, N1414);
not NOT1 (N1416, N1400);
buf BUF1 (N1417, N1399);
xor XOR2 (N1418, N1416, N959);
and AND3 (N1419, N1418, N624, N60);
nand NAND2 (N1420, N1413, N935);
nor NOR3 (N1421, N1417, N118, N1188);
nand NAND3 (N1422, N1420, N415, N895);
and AND4 (N1423, N1408, N143, N5, N1172);
nand NAND2 (N1424, N1423, N135);
or OR4 (N1425, N1424, N942, N445, N1264);
nor NOR3 (N1426, N1385, N147, N1103);
not NOT1 (N1427, N1415);
not NOT1 (N1428, N1422);
not NOT1 (N1429, N1428);
not NOT1 (N1430, N1427);
buf BUF1 (N1431, N1404);
nor NOR4 (N1432, N1430, N551, N1252, N1424);
and AND2 (N1433, N1426, N1156);
xor XOR2 (N1434, N1419, N977);
or OR4 (N1435, N1410, N636, N260, N984);
nand NAND2 (N1436, N1435, N1256);
buf BUF1 (N1437, N1433);
and AND4 (N1438, N1437, N1004, N1433, N1058);
buf BUF1 (N1439, N1431);
buf BUF1 (N1440, N1425);
buf BUF1 (N1441, N1438);
not NOT1 (N1442, N1441);
xor XOR2 (N1443, N1402, N191);
xor XOR2 (N1444, N1421, N69);
not NOT1 (N1445, N1440);
nor NOR2 (N1446, N1439, N1235);
xor XOR2 (N1447, N1434, N118);
nor NOR4 (N1448, N1411, N1143, N757, N619);
buf BUF1 (N1449, N1436);
or OR4 (N1450, N1448, N312, N778, N138);
nor NOR2 (N1451, N1432, N204);
not NOT1 (N1452, N1429);
or OR3 (N1453, N1452, N239, N432);
not NOT1 (N1454, N1449);
nor NOR3 (N1455, N1451, N1000, N1379);
not NOT1 (N1456, N1442);
and AND3 (N1457, N1456, N941, N580);
or OR3 (N1458, N1447, N97, N1333);
nand NAND2 (N1459, N1446, N821);
buf BUF1 (N1460, N1450);
nand NAND4 (N1461, N1454, N1355, N315, N1019);
or OR3 (N1462, N1453, N337, N672);
buf BUF1 (N1463, N1443);
nand NAND3 (N1464, N1460, N464, N848);
nand NAND2 (N1465, N1457, N813);
buf BUF1 (N1466, N1455);
xor XOR2 (N1467, N1466, N533);
nor NOR2 (N1468, N1462, N958);
buf BUF1 (N1469, N1463);
nand NAND4 (N1470, N1445, N587, N431, N992);
or OR2 (N1471, N1461, N1149);
buf BUF1 (N1472, N1459);
nand NAND2 (N1473, N1444, N1322);
or OR3 (N1474, N1470, N623, N604);
not NOT1 (N1475, N1473);
nor NOR3 (N1476, N1475, N1088, N1091);
buf BUF1 (N1477, N1458);
or OR4 (N1478, N1465, N1160, N799, N369);
or OR4 (N1479, N1476, N1067, N461, N1443);
or OR4 (N1480, N1471, N558, N507, N809);
or OR3 (N1481, N1478, N464, N1419);
not NOT1 (N1482, N1472);
nand NAND3 (N1483, N1482, N120, N967);
not NOT1 (N1484, N1480);
not NOT1 (N1485, N1481);
nand NAND3 (N1486, N1484, N748, N1339);
buf BUF1 (N1487, N1467);
buf BUF1 (N1488, N1468);
xor XOR2 (N1489, N1488, N404);
or OR4 (N1490, N1477, N230, N1168, N420);
not NOT1 (N1491, N1489);
buf BUF1 (N1492, N1487);
xor XOR2 (N1493, N1492, N515);
or OR4 (N1494, N1464, N1169, N721, N927);
or OR3 (N1495, N1479, N304, N1492);
and AND2 (N1496, N1469, N1000);
not NOT1 (N1497, N1493);
not NOT1 (N1498, N1474);
or OR2 (N1499, N1486, N232);
not NOT1 (N1500, N1495);
xor XOR2 (N1501, N1494, N1195);
not NOT1 (N1502, N1500);
and AND3 (N1503, N1501, N89, N988);
buf BUF1 (N1504, N1503);
or OR3 (N1505, N1490, N894, N100);
not NOT1 (N1506, N1497);
nor NOR3 (N1507, N1496, N398, N624);
buf BUF1 (N1508, N1506);
xor XOR2 (N1509, N1508, N946);
and AND3 (N1510, N1504, N488, N427);
and AND3 (N1511, N1499, N776, N1441);
nor NOR3 (N1512, N1491, N1325, N706);
and AND3 (N1513, N1510, N645, N143);
nand NAND3 (N1514, N1511, N1101, N676);
not NOT1 (N1515, N1505);
or OR3 (N1516, N1512, N617, N735);
not NOT1 (N1517, N1513);
not NOT1 (N1518, N1514);
buf BUF1 (N1519, N1515);
or OR4 (N1520, N1498, N511, N1065, N1493);
nor NOR3 (N1521, N1507, N1048, N1378);
or OR2 (N1522, N1485, N89);
or OR4 (N1523, N1522, N285, N912, N1040);
xor XOR2 (N1524, N1521, N1389);
nand NAND2 (N1525, N1502, N399);
nor NOR4 (N1526, N1524, N255, N491, N536);
and AND3 (N1527, N1483, N1221, N470);
not NOT1 (N1528, N1520);
nor NOR3 (N1529, N1528, N444, N10);
nor NOR2 (N1530, N1527, N488);
buf BUF1 (N1531, N1518);
not NOT1 (N1532, N1526);
nor NOR2 (N1533, N1532, N1378);
nor NOR3 (N1534, N1529, N321, N1328);
xor XOR2 (N1535, N1533, N247);
nand NAND4 (N1536, N1534, N269, N95, N577);
nand NAND2 (N1537, N1536, N630);
xor XOR2 (N1538, N1523, N1248);
not NOT1 (N1539, N1517);
xor XOR2 (N1540, N1535, N207);
or OR3 (N1541, N1530, N357, N26);
xor XOR2 (N1542, N1541, N1478);
not NOT1 (N1543, N1525);
and AND4 (N1544, N1539, N943, N785, N1483);
xor XOR2 (N1545, N1531, N98);
buf BUF1 (N1546, N1543);
xor XOR2 (N1547, N1537, N1259);
and AND4 (N1548, N1519, N190, N337, N962);
xor XOR2 (N1549, N1548, N1428);
nand NAND3 (N1550, N1509, N436, N1000);
nand NAND4 (N1551, N1516, N1060, N419, N1204);
buf BUF1 (N1552, N1546);
nand NAND4 (N1553, N1545, N1226, N792, N1000);
and AND3 (N1554, N1552, N219, N412);
nor NOR2 (N1555, N1544, N819);
xor XOR2 (N1556, N1550, N1340);
nor NOR3 (N1557, N1554, N995, N613);
nor NOR3 (N1558, N1540, N1024, N39);
xor XOR2 (N1559, N1558, N1186);
nor NOR3 (N1560, N1555, N1534, N594);
nand NAND4 (N1561, N1551, N1018, N753, N611);
nor NOR3 (N1562, N1553, N1182, N873);
xor XOR2 (N1563, N1538, N226);
nand NAND2 (N1564, N1547, N143);
and AND4 (N1565, N1557, N365, N1392, N1151);
and AND4 (N1566, N1559, N1214, N1327, N488);
nor NOR4 (N1567, N1565, N165, N456, N568);
or OR3 (N1568, N1566, N1324, N655);
nor NOR3 (N1569, N1560, N650, N780);
not NOT1 (N1570, N1562);
nand NAND2 (N1571, N1561, N631);
or OR3 (N1572, N1569, N1197, N1165);
not NOT1 (N1573, N1567);
or OR2 (N1574, N1570, N26);
or OR3 (N1575, N1573, N835, N1540);
and AND4 (N1576, N1568, N539, N1419, N1119);
and AND3 (N1577, N1542, N749, N1268);
not NOT1 (N1578, N1564);
nor NOR4 (N1579, N1576, N1450, N351, N154);
buf BUF1 (N1580, N1549);
and AND3 (N1581, N1580, N902, N1540);
buf BUF1 (N1582, N1571);
or OR3 (N1583, N1577, N343, N218);
buf BUF1 (N1584, N1556);
nand NAND4 (N1585, N1582, N1240, N931, N881);
buf BUF1 (N1586, N1572);
not NOT1 (N1587, N1586);
nor NOR4 (N1588, N1587, N452, N575, N506);
buf BUF1 (N1589, N1575);
nand NAND3 (N1590, N1585, N1374, N861);
nand NAND2 (N1591, N1584, N1195);
or OR4 (N1592, N1583, N721, N297, N1451);
and AND4 (N1593, N1563, N1071, N259, N729);
not NOT1 (N1594, N1579);
xor XOR2 (N1595, N1588, N388);
buf BUF1 (N1596, N1594);
not NOT1 (N1597, N1591);
and AND4 (N1598, N1574, N411, N1236, N258);
nor NOR4 (N1599, N1589, N758, N1174, N1255);
or OR4 (N1600, N1590, N1570, N104, N348);
nor NOR3 (N1601, N1593, N740, N124);
or OR3 (N1602, N1597, N78, N742);
buf BUF1 (N1603, N1578);
and AND3 (N1604, N1600, N97, N205);
and AND2 (N1605, N1602, N1108);
nand NAND4 (N1606, N1604, N152, N1290, N118);
buf BUF1 (N1607, N1595);
nand NAND4 (N1608, N1601, N1092, N1361, N1067);
xor XOR2 (N1609, N1607, N1467);
nor NOR2 (N1610, N1608, N102);
buf BUF1 (N1611, N1605);
buf BUF1 (N1612, N1609);
and AND4 (N1613, N1592, N939, N73, N1004);
nand NAND3 (N1614, N1611, N412, N228);
not NOT1 (N1615, N1613);
not NOT1 (N1616, N1612);
xor XOR2 (N1617, N1596, N961);
nor NOR3 (N1618, N1615, N1173, N610);
xor XOR2 (N1619, N1581, N184);
nor NOR3 (N1620, N1614, N704, N835);
and AND4 (N1621, N1617, N775, N611, N652);
or OR3 (N1622, N1610, N1074, N1419);
and AND3 (N1623, N1619, N175, N1079);
xor XOR2 (N1624, N1603, N710);
xor XOR2 (N1625, N1618, N1348);
or OR4 (N1626, N1621, N688, N1445, N456);
and AND3 (N1627, N1598, N760, N843);
or OR3 (N1628, N1626, N287, N636);
and AND4 (N1629, N1623, N565, N1042, N696);
buf BUF1 (N1630, N1629);
nor NOR2 (N1631, N1599, N1607);
xor XOR2 (N1632, N1622, N120);
nor NOR3 (N1633, N1616, N698, N1103);
nand NAND2 (N1634, N1628, N108);
or OR4 (N1635, N1606, N1600, N1504, N320);
and AND2 (N1636, N1620, N1104);
and AND2 (N1637, N1627, N565);
and AND2 (N1638, N1635, N1503);
not NOT1 (N1639, N1624);
and AND2 (N1640, N1636, N1137);
buf BUF1 (N1641, N1633);
nor NOR2 (N1642, N1637, N76);
nor NOR3 (N1643, N1642, N774, N277);
nor NOR2 (N1644, N1640, N561);
xor XOR2 (N1645, N1644, N845);
not NOT1 (N1646, N1641);
not NOT1 (N1647, N1625);
buf BUF1 (N1648, N1631);
xor XOR2 (N1649, N1643, N828);
not NOT1 (N1650, N1634);
or OR4 (N1651, N1639, N401, N1566, N164);
xor XOR2 (N1652, N1632, N1416);
not NOT1 (N1653, N1648);
and AND4 (N1654, N1630, N1394, N451, N360);
nor NOR4 (N1655, N1653, N1180, N616, N490);
buf BUF1 (N1656, N1638);
buf BUF1 (N1657, N1656);
buf BUF1 (N1658, N1650);
xor XOR2 (N1659, N1651, N1607);
or OR3 (N1660, N1657, N641, N1636);
and AND2 (N1661, N1655, N1248);
and AND3 (N1662, N1660, N1025, N1219);
nand NAND2 (N1663, N1654, N738);
nand NAND4 (N1664, N1646, N84, N440, N24);
buf BUF1 (N1665, N1659);
nand NAND4 (N1666, N1649, N934, N654, N998);
buf BUF1 (N1667, N1647);
and AND2 (N1668, N1658, N1549);
nor NOR2 (N1669, N1665, N89);
buf BUF1 (N1670, N1669);
and AND2 (N1671, N1668, N769);
and AND4 (N1672, N1645, N271, N1241, N86);
nand NAND3 (N1673, N1671, N456, N1514);
nand NAND4 (N1674, N1673, N898, N336, N1091);
nor NOR4 (N1675, N1667, N935, N1131, N397);
and AND4 (N1676, N1666, N878, N1342, N352);
not NOT1 (N1677, N1661);
nor NOR3 (N1678, N1662, N1274, N797);
buf BUF1 (N1679, N1676);
nor NOR4 (N1680, N1674, N304, N922, N1012);
nand NAND2 (N1681, N1677, N488);
or OR4 (N1682, N1670, N560, N738, N730);
or OR4 (N1683, N1679, N309, N313, N1051);
not NOT1 (N1684, N1683);
nand NAND3 (N1685, N1678, N1510, N533);
nand NAND2 (N1686, N1672, N819);
xor XOR2 (N1687, N1685, N923);
nand NAND4 (N1688, N1675, N875, N1110, N1075);
nand NAND3 (N1689, N1681, N1679, N370);
or OR4 (N1690, N1689, N652, N451, N1307);
not NOT1 (N1691, N1652);
buf BUF1 (N1692, N1691);
nand NAND3 (N1693, N1690, N7, N577);
nor NOR4 (N1694, N1687, N577, N854, N452);
buf BUF1 (N1695, N1682);
or OR4 (N1696, N1686, N202, N259, N463);
xor XOR2 (N1697, N1694, N934);
not NOT1 (N1698, N1693);
nor NOR3 (N1699, N1692, N129, N815);
buf BUF1 (N1700, N1695);
not NOT1 (N1701, N1696);
not NOT1 (N1702, N1700);
xor XOR2 (N1703, N1684, N913);
xor XOR2 (N1704, N1680, N184);
and AND4 (N1705, N1704, N1415, N1511, N572);
xor XOR2 (N1706, N1698, N714);
nor NOR2 (N1707, N1701, N153);
nand NAND3 (N1708, N1697, N1330, N1704);
or OR4 (N1709, N1688, N739, N1229, N1180);
not NOT1 (N1710, N1709);
buf BUF1 (N1711, N1699);
or OR3 (N1712, N1664, N192, N1503);
nand NAND2 (N1713, N1706, N208);
and AND4 (N1714, N1712, N1302, N1479, N1624);
and AND2 (N1715, N1710, N1043);
buf BUF1 (N1716, N1713);
not NOT1 (N1717, N1708);
and AND3 (N1718, N1711, N140, N1625);
or OR2 (N1719, N1663, N1502);
and AND2 (N1720, N1703, N54);
buf BUF1 (N1721, N1705);
xor XOR2 (N1722, N1715, N1518);
or OR4 (N1723, N1716, N1430, N1344, N1229);
or OR2 (N1724, N1720, N259);
not NOT1 (N1725, N1702);
not NOT1 (N1726, N1714);
buf BUF1 (N1727, N1724);
buf BUF1 (N1728, N1707);
and AND4 (N1729, N1725, N1162, N1020, N187);
buf BUF1 (N1730, N1719);
not NOT1 (N1731, N1726);
or OR3 (N1732, N1729, N1107, N589);
nand NAND3 (N1733, N1728, N350, N1600);
nand NAND3 (N1734, N1722, N303, N1336);
xor XOR2 (N1735, N1732, N951);
or OR2 (N1736, N1723, N1075);
not NOT1 (N1737, N1718);
and AND2 (N1738, N1727, N1354);
nor NOR4 (N1739, N1730, N1698, N694, N956);
xor XOR2 (N1740, N1717, N1728);
nand NAND4 (N1741, N1735, N1694, N842, N846);
not NOT1 (N1742, N1737);
and AND4 (N1743, N1741, N1549, N362, N130);
xor XOR2 (N1744, N1721, N729);
nor NOR3 (N1745, N1731, N1218, N1609);
or OR2 (N1746, N1738, N1273);
and AND4 (N1747, N1733, N1647, N1517, N837);
or OR2 (N1748, N1745, N510);
buf BUF1 (N1749, N1743);
nand NAND3 (N1750, N1744, N358, N1611);
nand NAND2 (N1751, N1749, N377);
buf BUF1 (N1752, N1740);
or OR2 (N1753, N1746, N53);
xor XOR2 (N1754, N1736, N1308);
or OR2 (N1755, N1734, N1099);
xor XOR2 (N1756, N1751, N121);
nor NOR2 (N1757, N1739, N1608);
nand NAND4 (N1758, N1757, N1464, N1672, N1707);
not NOT1 (N1759, N1753);
xor XOR2 (N1760, N1748, N1728);
and AND3 (N1761, N1752, N380, N1319);
nor NOR2 (N1762, N1760, N1162);
not NOT1 (N1763, N1762);
not NOT1 (N1764, N1758);
buf BUF1 (N1765, N1756);
not NOT1 (N1766, N1764);
or OR4 (N1767, N1765, N475, N1736, N185);
nand NAND4 (N1768, N1766, N1686, N1707, N531);
buf BUF1 (N1769, N1747);
and AND2 (N1770, N1763, N1750);
xor XOR2 (N1771, N1030, N1380);
nor NOR2 (N1772, N1742, N1613);
nor NOR2 (N1773, N1768, N288);
buf BUF1 (N1774, N1754);
xor XOR2 (N1775, N1774, N1282);
not NOT1 (N1776, N1767);
buf BUF1 (N1777, N1755);
and AND2 (N1778, N1777, N322);
or OR3 (N1779, N1775, N1277, N1699);
xor XOR2 (N1780, N1772, N958);
or OR3 (N1781, N1780, N430, N891);
and AND3 (N1782, N1769, N208, N745);
buf BUF1 (N1783, N1781);
buf BUF1 (N1784, N1776);
or OR2 (N1785, N1778, N987);
buf BUF1 (N1786, N1771);
nor NOR3 (N1787, N1786, N1101, N1117);
nand NAND2 (N1788, N1770, N431);
not NOT1 (N1789, N1788);
xor XOR2 (N1790, N1782, N1756);
not NOT1 (N1791, N1785);
and AND4 (N1792, N1773, N1250, N876, N878);
nand NAND3 (N1793, N1761, N946, N1761);
nor NOR3 (N1794, N1793, N1359, N790);
buf BUF1 (N1795, N1794);
and AND4 (N1796, N1784, N1305, N1044, N292);
or OR4 (N1797, N1783, N841, N1238, N1549);
and AND4 (N1798, N1787, N753, N1522, N607);
buf BUF1 (N1799, N1779);
xor XOR2 (N1800, N1792, N678);
nand NAND2 (N1801, N1759, N973);
nor NOR2 (N1802, N1790, N155);
not NOT1 (N1803, N1801);
buf BUF1 (N1804, N1796);
and AND4 (N1805, N1795, N706, N1713, N1787);
buf BUF1 (N1806, N1797);
buf BUF1 (N1807, N1799);
not NOT1 (N1808, N1804);
not NOT1 (N1809, N1803);
nor NOR2 (N1810, N1789, N381);
nor NOR4 (N1811, N1808, N599, N1049, N1331);
xor XOR2 (N1812, N1802, N14);
buf BUF1 (N1813, N1805);
or OR4 (N1814, N1811, N368, N1763, N1442);
xor XOR2 (N1815, N1806, N1173);
and AND4 (N1816, N1815, N880, N1179, N644);
or OR4 (N1817, N1809, N1076, N1191, N1455);
or OR3 (N1818, N1791, N1653, N368);
not NOT1 (N1819, N1800);
not NOT1 (N1820, N1807);
xor XOR2 (N1821, N1813, N849);
xor XOR2 (N1822, N1821, N1519);
xor XOR2 (N1823, N1816, N1495);
nand NAND4 (N1824, N1822, N333, N1327, N479);
and AND4 (N1825, N1810, N1360, N359, N287);
or OR4 (N1826, N1825, N1218, N431, N1220);
and AND4 (N1827, N1820, N1001, N1289, N712);
and AND2 (N1828, N1826, N715);
nor NOR3 (N1829, N1824, N1234, N487);
buf BUF1 (N1830, N1828);
buf BUF1 (N1831, N1827);
or OR4 (N1832, N1812, N944, N617, N1769);
nor NOR2 (N1833, N1818, N1137);
buf BUF1 (N1834, N1823);
or OR2 (N1835, N1819, N1283);
nand NAND3 (N1836, N1834, N16, N1045);
or OR2 (N1837, N1829, N658);
nand NAND4 (N1838, N1817, N356, N1370, N201);
not NOT1 (N1839, N1833);
nor NOR4 (N1840, N1814, N1816, N193, N1134);
and AND4 (N1841, N1835, N1464, N1545, N178);
buf BUF1 (N1842, N1832);
buf BUF1 (N1843, N1830);
and AND4 (N1844, N1840, N1019, N685, N276);
nor NOR2 (N1845, N1838, N204);
and AND4 (N1846, N1845, N199, N1672, N1759);
nor NOR2 (N1847, N1837, N452);
nor NOR3 (N1848, N1847, N2, N1788);
xor XOR2 (N1849, N1843, N492);
not NOT1 (N1850, N1798);
buf BUF1 (N1851, N1836);
nor NOR3 (N1852, N1841, N267, N31);
buf BUF1 (N1853, N1850);
nand NAND2 (N1854, N1851, N407);
xor XOR2 (N1855, N1839, N201);
nor NOR4 (N1856, N1852, N577, N526, N1080);
xor XOR2 (N1857, N1831, N356);
xor XOR2 (N1858, N1844, N1141);
buf BUF1 (N1859, N1846);
nand NAND2 (N1860, N1859, N482);
buf BUF1 (N1861, N1856);
not NOT1 (N1862, N1860);
xor XOR2 (N1863, N1857, N1367);
xor XOR2 (N1864, N1842, N1027);
nand NAND3 (N1865, N1849, N200, N83);
nor NOR2 (N1866, N1863, N1091);
or OR2 (N1867, N1862, N782);
not NOT1 (N1868, N1867);
or OR3 (N1869, N1858, N33, N583);
or OR2 (N1870, N1848, N1011);
nand NAND4 (N1871, N1869, N901, N21, N241);
or OR4 (N1872, N1870, N331, N1022, N1090);
not NOT1 (N1873, N1872);
nor NOR3 (N1874, N1873, N1338, N1043);
xor XOR2 (N1875, N1871, N1798);
buf BUF1 (N1876, N1853);
or OR3 (N1877, N1854, N1532, N1761);
nand NAND2 (N1878, N1875, N610);
nand NAND2 (N1879, N1855, N274);
or OR2 (N1880, N1876, N1160);
xor XOR2 (N1881, N1864, N1345);
and AND2 (N1882, N1866, N16);
nor NOR4 (N1883, N1882, N1473, N1628, N1750);
and AND3 (N1884, N1883, N1565, N1135);
nor NOR3 (N1885, N1880, N1460, N1733);
or OR2 (N1886, N1868, N1186);
xor XOR2 (N1887, N1865, N896);
and AND4 (N1888, N1885, N999, N1188, N125);
buf BUF1 (N1889, N1878);
not NOT1 (N1890, N1877);
nor NOR4 (N1891, N1887, N815, N444, N951);
nor NOR4 (N1892, N1879, N214, N262, N818);
not NOT1 (N1893, N1884);
or OR3 (N1894, N1892, N1314, N1797);
buf BUF1 (N1895, N1881);
nor NOR3 (N1896, N1894, N388, N1099);
buf BUF1 (N1897, N1889);
and AND2 (N1898, N1897, N593);
and AND3 (N1899, N1896, N1304, N954);
buf BUF1 (N1900, N1874);
nand NAND4 (N1901, N1900, N847, N1790, N379);
nand NAND4 (N1902, N1901, N1037, N1829, N1768);
or OR3 (N1903, N1893, N1703, N1217);
or OR2 (N1904, N1886, N294);
xor XOR2 (N1905, N1903, N1300);
buf BUF1 (N1906, N1898);
nand NAND4 (N1907, N1890, N807, N635, N1295);
not NOT1 (N1908, N1902);
not NOT1 (N1909, N1891);
and AND4 (N1910, N1907, N887, N1280, N355);
or OR3 (N1911, N1906, N635, N1712);
nor NOR4 (N1912, N1904, N1482, N579, N1563);
not NOT1 (N1913, N1912);
or OR4 (N1914, N1910, N1807, N763, N431);
and AND3 (N1915, N1895, N1480, N93);
nand NAND3 (N1916, N1915, N953, N915);
and AND3 (N1917, N1916, N1658, N1063);
buf BUF1 (N1918, N1917);
and AND3 (N1919, N1905, N541, N916);
xor XOR2 (N1920, N1918, N1711);
buf BUF1 (N1921, N1919);
nand NAND4 (N1922, N1908, N241, N1812, N103);
xor XOR2 (N1923, N1899, N1279);
nand NAND3 (N1924, N1909, N478, N1873);
not NOT1 (N1925, N1911);
and AND3 (N1926, N1920, N823, N1041);
xor XOR2 (N1927, N1888, N4);
and AND2 (N1928, N1913, N1431);
buf BUF1 (N1929, N1928);
nor NOR2 (N1930, N1925, N1763);
not NOT1 (N1931, N1923);
or OR4 (N1932, N1929, N21, N863, N90);
nor NOR4 (N1933, N1921, N975, N1415, N1752);
nand NAND4 (N1934, N1930, N1226, N1779, N103);
xor XOR2 (N1935, N1914, N680);
nor NOR2 (N1936, N1932, N813);
and AND2 (N1937, N1936, N251);
xor XOR2 (N1938, N1926, N1730);
nor NOR2 (N1939, N1931, N455);
xor XOR2 (N1940, N1922, N1456);
not NOT1 (N1941, N1933);
and AND4 (N1942, N1939, N1828, N1860, N943);
and AND4 (N1943, N1940, N1719, N1766, N301);
not NOT1 (N1944, N1938);
buf BUF1 (N1945, N1937);
or OR3 (N1946, N1944, N1503, N761);
nand NAND2 (N1947, N1941, N210);
nand NAND3 (N1948, N1861, N1703, N1165);
nor NOR2 (N1949, N1946, N1424);
and AND3 (N1950, N1948, N1597, N120);
and AND4 (N1951, N1947, N1298, N1195, N1813);
nor NOR2 (N1952, N1943, N1511);
and AND2 (N1953, N1927, N1366);
xor XOR2 (N1954, N1934, N1151);
xor XOR2 (N1955, N1945, N669);
buf BUF1 (N1956, N1935);
not NOT1 (N1957, N1955);
nor NOR2 (N1958, N1949, N77);
not NOT1 (N1959, N1942);
and AND4 (N1960, N1950, N190, N166, N1939);
nor NOR2 (N1961, N1951, N1047);
buf BUF1 (N1962, N1952);
or OR2 (N1963, N1953, N1684);
and AND2 (N1964, N1961, N604);
and AND4 (N1965, N1964, N1529, N225, N1335);
buf BUF1 (N1966, N1959);
or OR2 (N1967, N1924, N469);
nand NAND3 (N1968, N1962, N1622, N981);
nor NOR2 (N1969, N1963, N664);
and AND2 (N1970, N1967, N1006);
and AND2 (N1971, N1966, N644);
nand NAND4 (N1972, N1954, N92, N1133, N1367);
and AND4 (N1973, N1970, N891, N179, N1889);
not NOT1 (N1974, N1960);
nand NAND2 (N1975, N1974, N166);
not NOT1 (N1976, N1968);
nor NOR2 (N1977, N1971, N271);
and AND3 (N1978, N1957, N319, N1471);
not NOT1 (N1979, N1973);
and AND3 (N1980, N1978, N1260, N978);
xor XOR2 (N1981, N1975, N230);
xor XOR2 (N1982, N1969, N1955);
or OR2 (N1983, N1977, N599);
buf BUF1 (N1984, N1980);
xor XOR2 (N1985, N1956, N408);
and AND2 (N1986, N1985, N871);
xor XOR2 (N1987, N1972, N1005);
nor NOR3 (N1988, N1965, N1238, N1290);
not NOT1 (N1989, N1976);
nor NOR2 (N1990, N1989, N1832);
buf BUF1 (N1991, N1983);
buf BUF1 (N1992, N1986);
not NOT1 (N1993, N1992);
xor XOR2 (N1994, N1993, N1316);
nand NAND2 (N1995, N1982, N803);
xor XOR2 (N1996, N1988, N1607);
nand NAND4 (N1997, N1996, N274, N268, N92);
nand NAND2 (N1998, N1987, N1974);
not NOT1 (N1999, N1990);
or OR2 (N2000, N1994, N1226);
not NOT1 (N2001, N1991);
nor NOR3 (N2002, N1997, N272, N1386);
not NOT1 (N2003, N1995);
and AND4 (N2004, N2002, N222, N1019, N43);
nand NAND2 (N2005, N1984, N100);
or OR2 (N2006, N2003, N510);
or OR2 (N2007, N2004, N1269);
buf BUF1 (N2008, N1999);
nand NAND2 (N2009, N2008, N1504);
nand NAND2 (N2010, N2009, N1629);
nand NAND4 (N2011, N2007, N603, N431, N419);
nand NAND2 (N2012, N2006, N360);
not NOT1 (N2013, N2011);
or OR4 (N2014, N1998, N1152, N675, N1411);
not NOT1 (N2015, N1979);
buf BUF1 (N2016, N2015);
not NOT1 (N2017, N2012);
nand NAND2 (N2018, N2016, N1531);
nor NOR3 (N2019, N2005, N1881, N1696);
nor NOR3 (N2020, N2019, N1299, N844);
and AND4 (N2021, N2010, N1108, N45, N1618);
xor XOR2 (N2022, N1981, N1504);
buf BUF1 (N2023, N2021);
buf BUF1 (N2024, N2023);
or OR2 (N2025, N2018, N1034);
or OR2 (N2026, N2013, N1013);
and AND3 (N2027, N2014, N698, N30);
buf BUF1 (N2028, N2027);
or OR4 (N2029, N1958, N547, N1034, N614);
nand NAND4 (N2030, N2000, N491, N1530, N1092);
or OR4 (N2031, N2030, N1140, N1166, N888);
or OR2 (N2032, N2024, N818);
nor NOR3 (N2033, N2031, N1208, N913);
nand NAND2 (N2034, N2028, N1098);
nor NOR4 (N2035, N2001, N1903, N1188, N1995);
not NOT1 (N2036, N2029);
nor NOR4 (N2037, N2020, N84, N1583, N56);
or OR3 (N2038, N2026, N395, N1572);
nand NAND3 (N2039, N2033, N239, N1455);
not NOT1 (N2040, N2036);
not NOT1 (N2041, N2037);
and AND2 (N2042, N2017, N1841);
not NOT1 (N2043, N2025);
buf BUF1 (N2044, N2022);
nor NOR4 (N2045, N2039, N798, N1404, N1974);
nor NOR3 (N2046, N2038, N1095, N1159);
xor XOR2 (N2047, N2041, N1640);
not NOT1 (N2048, N2047);
xor XOR2 (N2049, N2042, N1724);
buf BUF1 (N2050, N2048);
or OR2 (N2051, N2032, N1511);
nor NOR2 (N2052, N2050, N1890);
not NOT1 (N2053, N2044);
buf BUF1 (N2054, N2052);
and AND2 (N2055, N2043, N841);
nor NOR4 (N2056, N2040, N1210, N1425, N1684);
nor NOR3 (N2057, N2056, N469, N635);
nor NOR4 (N2058, N2049, N1975, N44, N490);
buf BUF1 (N2059, N2054);
nand NAND2 (N2060, N2057, N731);
and AND2 (N2061, N2060, N1677);
nor NOR2 (N2062, N2053, N1117);
nor NOR4 (N2063, N2061, N57, N456, N106);
nor NOR3 (N2064, N2045, N2052, N425);
xor XOR2 (N2065, N2059, N1002);
xor XOR2 (N2066, N2065, N597);
and AND3 (N2067, N2058, N1550, N803);
and AND2 (N2068, N2051, N1079);
not NOT1 (N2069, N2034);
or OR2 (N2070, N2068, N901);
xor XOR2 (N2071, N2066, N1031);
buf BUF1 (N2072, N2064);
xor XOR2 (N2073, N2062, N1820);
buf BUF1 (N2074, N2072);
or OR3 (N2075, N2073, N1872, N1940);
nand NAND3 (N2076, N2035, N150, N1002);
nor NOR4 (N2077, N2069, N1882, N1100, N1681);
buf BUF1 (N2078, N2070);
buf BUF1 (N2079, N2077);
or OR3 (N2080, N2074, N1240, N79);
xor XOR2 (N2081, N2075, N1515);
and AND2 (N2082, N2080, N960);
or OR4 (N2083, N2055, N1871, N964, N14);
not NOT1 (N2084, N2078);
buf BUF1 (N2085, N2083);
nor NOR3 (N2086, N2046, N1514, N1473);
nor NOR4 (N2087, N2081, N1021, N1936, N1225);
nand NAND2 (N2088, N2071, N2067);
xor XOR2 (N2089, N1664, N518);
and AND3 (N2090, N2082, N258, N1217);
and AND3 (N2091, N2090, N950, N1460);
buf BUF1 (N2092, N2086);
or OR2 (N2093, N2088, N1639);
buf BUF1 (N2094, N2079);
nor NOR3 (N2095, N2089, N823, N2047);
not NOT1 (N2096, N2091);
nor NOR2 (N2097, N2063, N827);
nor NOR4 (N2098, N2085, N1430, N1902, N2066);
nor NOR3 (N2099, N2087, N1934, N1806);
and AND3 (N2100, N2084, N731, N1951);
nand NAND3 (N2101, N2094, N1907, N2058);
buf BUF1 (N2102, N2096);
nor NOR3 (N2103, N2102, N587, N1296);
buf BUF1 (N2104, N2095);
nor NOR4 (N2105, N2104, N1181, N1171, N874);
buf BUF1 (N2106, N2093);
nor NOR4 (N2107, N2103, N1148, N1450, N1905);
nor NOR2 (N2108, N2098, N248);
or OR2 (N2109, N2076, N1095);
xor XOR2 (N2110, N2109, N1129);
nor NOR3 (N2111, N2107, N360, N222);
not NOT1 (N2112, N2092);
and AND2 (N2113, N2110, N1863);
buf BUF1 (N2114, N2100);
xor XOR2 (N2115, N2108, N91);
buf BUF1 (N2116, N2114);
buf BUF1 (N2117, N2105);
buf BUF1 (N2118, N2101);
xor XOR2 (N2119, N2117, N487);
nand NAND3 (N2120, N2099, N2014, N147);
buf BUF1 (N2121, N2111);
nor NOR4 (N2122, N2112, N933, N891, N1374);
nor NOR2 (N2123, N2115, N899);
or OR4 (N2124, N2120, N1356, N676, N1315);
xor XOR2 (N2125, N2116, N1078);
not NOT1 (N2126, N2106);
buf BUF1 (N2127, N2125);
nor NOR2 (N2128, N2122, N444);
and AND3 (N2129, N2119, N2026, N46);
not NOT1 (N2130, N2123);
nor NOR3 (N2131, N2121, N965, N791);
or OR4 (N2132, N2097, N771, N246, N104);
or OR2 (N2133, N2124, N1613);
nand NAND3 (N2134, N2126, N82, N1930);
or OR3 (N2135, N2113, N546, N1811);
not NOT1 (N2136, N2132);
or OR4 (N2137, N2127, N1218, N350, N2083);
buf BUF1 (N2138, N2130);
buf BUF1 (N2139, N2136);
nand NAND2 (N2140, N2128, N1308);
nor NOR3 (N2141, N2134, N494, N123);
not NOT1 (N2142, N2138);
not NOT1 (N2143, N2129);
and AND4 (N2144, N2133, N1107, N862, N1660);
and AND3 (N2145, N2141, N330, N1014);
nor NOR2 (N2146, N2142, N1137);
or OR4 (N2147, N2146, N454, N1860, N338);
nor NOR2 (N2148, N2145, N597);
buf BUF1 (N2149, N2131);
buf BUF1 (N2150, N2149);
or OR4 (N2151, N2139, N1325, N1113, N934);
buf BUF1 (N2152, N2151);
or OR3 (N2153, N2143, N1872, N149);
nor NOR3 (N2154, N2147, N1516, N88);
xor XOR2 (N2155, N2135, N1589);
buf BUF1 (N2156, N2144);
xor XOR2 (N2157, N2152, N2091);
or OR2 (N2158, N2157, N1783);
nand NAND3 (N2159, N2137, N1969, N87);
nand NAND2 (N2160, N2159, N862);
nor NOR4 (N2161, N2158, N1994, N2083, N1490);
buf BUF1 (N2162, N2140);
not NOT1 (N2163, N2156);
not NOT1 (N2164, N2150);
xor XOR2 (N2165, N2118, N747);
and AND4 (N2166, N2153, N743, N784, N1744);
buf BUF1 (N2167, N2160);
nand NAND3 (N2168, N2161, N696, N15);
xor XOR2 (N2169, N2163, N1796);
nor NOR3 (N2170, N2154, N642, N181);
not NOT1 (N2171, N2167);
nand NAND3 (N2172, N2155, N1592, N900);
and AND2 (N2173, N2172, N916);
and AND2 (N2174, N2170, N454);
or OR4 (N2175, N2169, N562, N2025, N757);
or OR4 (N2176, N2173, N1210, N513, N981);
not NOT1 (N2177, N2165);
buf BUF1 (N2178, N2174);
not NOT1 (N2179, N2164);
or OR4 (N2180, N2175, N2146, N1253, N1993);
not NOT1 (N2181, N2148);
nand NAND4 (N2182, N2179, N111, N391, N1620);
or OR4 (N2183, N2181, N127, N851, N102);
xor XOR2 (N2184, N2180, N2005);
xor XOR2 (N2185, N2166, N642);
or OR4 (N2186, N2162, N1052, N2067, N1592);
and AND3 (N2187, N2183, N1231, N1808);
nor NOR3 (N2188, N2178, N1711, N2144);
xor XOR2 (N2189, N2176, N2085);
xor XOR2 (N2190, N2184, N1328);
nand NAND4 (N2191, N2189, N1948, N1646, N258);
or OR2 (N2192, N2190, N1028);
nor NOR3 (N2193, N2186, N1086, N674);
xor XOR2 (N2194, N2191, N158);
xor XOR2 (N2195, N2168, N1243);
not NOT1 (N2196, N2185);
not NOT1 (N2197, N2193);
buf BUF1 (N2198, N2197);
not NOT1 (N2199, N2187);
not NOT1 (N2200, N2194);
not NOT1 (N2201, N2199);
xor XOR2 (N2202, N2196, N65);
nor NOR3 (N2203, N2200, N408, N785);
nand NAND3 (N2204, N2188, N253, N659);
nor NOR4 (N2205, N2192, N327, N503, N578);
nand NAND4 (N2206, N2182, N1257, N1763, N627);
nand NAND3 (N2207, N2177, N1865, N1944);
not NOT1 (N2208, N2205);
xor XOR2 (N2209, N2202, N710);
or OR3 (N2210, N2201, N507, N1303);
not NOT1 (N2211, N2204);
not NOT1 (N2212, N2198);
and AND3 (N2213, N2209, N62, N208);
not NOT1 (N2214, N2203);
nor NOR4 (N2215, N2208, N20, N1256, N1015);
nor NOR2 (N2216, N2206, N1797);
xor XOR2 (N2217, N2195, N1106);
xor XOR2 (N2218, N2213, N1066);
nand NAND3 (N2219, N2212, N665, N1234);
or OR4 (N2220, N2214, N1159, N1918, N169);
nor NOR2 (N2221, N2207, N1011);
not NOT1 (N2222, N2210);
not NOT1 (N2223, N2215);
nand NAND3 (N2224, N2219, N1874, N245);
nor NOR2 (N2225, N2211, N1339);
nor NOR4 (N2226, N2220, N2209, N875, N1907);
and AND4 (N2227, N2217, N2128, N700, N848);
or OR2 (N2228, N2218, N1909);
buf BUF1 (N2229, N2222);
nor NOR4 (N2230, N2223, N1094, N959, N1263);
and AND4 (N2231, N2171, N1861, N1803, N151);
or OR3 (N2232, N2221, N953, N970);
xor XOR2 (N2233, N2229, N1592);
nand NAND3 (N2234, N2216, N1575, N2147);
buf BUF1 (N2235, N2225);
or OR2 (N2236, N2233, N2015);
not NOT1 (N2237, N2231);
and AND2 (N2238, N2235, N1951);
xor XOR2 (N2239, N2234, N1154);
not NOT1 (N2240, N2228);
not NOT1 (N2241, N2224);
or OR3 (N2242, N2230, N1769, N1957);
or OR2 (N2243, N2239, N2081);
not NOT1 (N2244, N2232);
or OR3 (N2245, N2227, N1855, N1059);
xor XOR2 (N2246, N2238, N167);
nor NOR2 (N2247, N2244, N1994);
not NOT1 (N2248, N2245);
xor XOR2 (N2249, N2226, N418);
not NOT1 (N2250, N2246);
not NOT1 (N2251, N2241);
nand NAND4 (N2252, N2250, N1408, N2212, N1054);
xor XOR2 (N2253, N2243, N1693);
nand NAND2 (N2254, N2253, N1808);
not NOT1 (N2255, N2254);
nor NOR3 (N2256, N2255, N584, N243);
xor XOR2 (N2257, N2240, N867);
or OR4 (N2258, N2249, N1894, N974, N175);
nor NOR2 (N2259, N2256, N1907);
buf BUF1 (N2260, N2237);
nand NAND4 (N2261, N2236, N2220, N1978, N1415);
buf BUF1 (N2262, N2242);
not NOT1 (N2263, N2262);
or OR4 (N2264, N2260, N1491, N223, N1407);
nand NAND2 (N2265, N2259, N860);
xor XOR2 (N2266, N2263, N283);
and AND3 (N2267, N2247, N2156, N492);
nor NOR3 (N2268, N2252, N30, N659);
xor XOR2 (N2269, N2261, N1002);
or OR3 (N2270, N2264, N660, N2224);
or OR4 (N2271, N2268, N1258, N2212, N1844);
or OR4 (N2272, N2258, N2174, N1319, N2024);
buf BUF1 (N2273, N2267);
and AND4 (N2274, N2266, N1880, N502, N2247);
buf BUF1 (N2275, N2257);
nor NOR3 (N2276, N2271, N822, N322);
nor NOR4 (N2277, N2274, N1770, N777, N1160);
not NOT1 (N2278, N2270);
nor NOR3 (N2279, N2251, N1097, N10);
not NOT1 (N2280, N2265);
nand NAND3 (N2281, N2280, N1045, N504);
or OR2 (N2282, N2279, N1725);
buf BUF1 (N2283, N2276);
or OR3 (N2284, N2281, N1662, N1150);
buf BUF1 (N2285, N2248);
and AND4 (N2286, N2285, N476, N1737, N1591);
nand NAND3 (N2287, N2286, N767, N304);
or OR3 (N2288, N2273, N590, N1844);
buf BUF1 (N2289, N2269);
nor NOR3 (N2290, N2287, N187, N276);
xor XOR2 (N2291, N2289, N1041);
xor XOR2 (N2292, N2288, N1473);
xor XOR2 (N2293, N2277, N965);
xor XOR2 (N2294, N2272, N922);
buf BUF1 (N2295, N2291);
nand NAND4 (N2296, N2292, N2046, N941, N1846);
xor XOR2 (N2297, N2275, N1100);
and AND4 (N2298, N2278, N2236, N1100, N716);
not NOT1 (N2299, N2298);
not NOT1 (N2300, N2283);
xor XOR2 (N2301, N2282, N1513);
buf BUF1 (N2302, N2295);
or OR4 (N2303, N2301, N734, N1600, N2271);
xor XOR2 (N2304, N2299, N417);
xor XOR2 (N2305, N2293, N337);
and AND2 (N2306, N2304, N1842);
nand NAND4 (N2307, N2305, N1487, N2084, N1668);
buf BUF1 (N2308, N2302);
nand NAND3 (N2309, N2303, N1767, N1333);
not NOT1 (N2310, N2297);
and AND3 (N2311, N2284, N1958, N2279);
xor XOR2 (N2312, N2294, N1115);
not NOT1 (N2313, N2312);
or OR2 (N2314, N2310, N1926);
nand NAND3 (N2315, N2307, N1145, N468);
nor NOR2 (N2316, N2315, N702);
xor XOR2 (N2317, N2308, N2135);
nand NAND4 (N2318, N2313, N1498, N783, N289);
or OR4 (N2319, N2290, N40, N1875, N1909);
or OR4 (N2320, N2306, N194, N625, N206);
or OR3 (N2321, N2320, N1953, N634);
nand NAND4 (N2322, N2296, N835, N1661, N1740);
nand NAND2 (N2323, N2314, N515);
nor NOR3 (N2324, N2309, N491, N2172);
not NOT1 (N2325, N2323);
nand NAND4 (N2326, N2324, N160, N1081, N1605);
or OR3 (N2327, N2318, N1227, N1732);
nand NAND4 (N2328, N2326, N398, N1261, N549);
or OR4 (N2329, N2327, N2284, N400, N491);
buf BUF1 (N2330, N2328);
buf BUF1 (N2331, N2322);
nor NOR4 (N2332, N2316, N1218, N1882, N2009);
buf BUF1 (N2333, N2325);
or OR4 (N2334, N2332, N112, N1772, N63);
nand NAND3 (N2335, N2334, N1345, N2229);
nor NOR2 (N2336, N2319, N1929);
xor XOR2 (N2337, N2311, N545);
nand NAND3 (N2338, N2337, N1345, N1755);
buf BUF1 (N2339, N2333);
or OR4 (N2340, N2300, N196, N1124, N282);
or OR2 (N2341, N2338, N1645);
or OR2 (N2342, N2321, N262);
or OR3 (N2343, N2317, N279, N1586);
buf BUF1 (N2344, N2335);
xor XOR2 (N2345, N2329, N1105);
or OR2 (N2346, N2345, N284);
buf BUF1 (N2347, N2330);
nor NOR4 (N2348, N2346, N125, N131, N924);
not NOT1 (N2349, N2343);
nand NAND3 (N2350, N2349, N1246, N2091);
and AND2 (N2351, N2341, N1160);
buf BUF1 (N2352, N2339);
nor NOR3 (N2353, N2336, N12, N2189);
nor NOR2 (N2354, N2353, N1736);
xor XOR2 (N2355, N2347, N752);
nor NOR4 (N2356, N2342, N2149, N1566, N1146);
nor NOR3 (N2357, N2348, N619, N320);
nand NAND4 (N2358, N2340, N1961, N1691, N90);
buf BUF1 (N2359, N2344);
and AND3 (N2360, N2356, N1433, N1281);
xor XOR2 (N2361, N2351, N306);
xor XOR2 (N2362, N2357, N349);
and AND3 (N2363, N2359, N316, N1639);
xor XOR2 (N2364, N2362, N709);
or OR2 (N2365, N2331, N1801);
or OR2 (N2366, N2358, N1203);
or OR4 (N2367, N2352, N2003, N2335, N558);
or OR2 (N2368, N2366, N583);
buf BUF1 (N2369, N2367);
or OR2 (N2370, N2369, N1446);
xor XOR2 (N2371, N2360, N2213);
and AND2 (N2372, N2365, N2353);
not NOT1 (N2373, N2368);
not NOT1 (N2374, N2355);
nor NOR2 (N2375, N2350, N365);
xor XOR2 (N2376, N2363, N677);
not NOT1 (N2377, N2354);
not NOT1 (N2378, N2377);
nor NOR2 (N2379, N2375, N251);
buf BUF1 (N2380, N2371);
xor XOR2 (N2381, N2378, N23);
buf BUF1 (N2382, N2374);
and AND3 (N2383, N2364, N448, N363);
nand NAND4 (N2384, N2379, N1288, N2350, N454);
xor XOR2 (N2385, N2384, N296);
or OR2 (N2386, N2382, N1912);
nand NAND4 (N2387, N2386, N432, N180, N679);
not NOT1 (N2388, N2376);
or OR2 (N2389, N2373, N2346);
and AND4 (N2390, N2385, N948, N204, N1836);
or OR2 (N2391, N2390, N2315);
xor XOR2 (N2392, N2389, N1490);
nand NAND3 (N2393, N2361, N1931, N838);
not NOT1 (N2394, N2387);
xor XOR2 (N2395, N2370, N1770);
xor XOR2 (N2396, N2395, N1366);
nor NOR3 (N2397, N2392, N1609, N1577);
not NOT1 (N2398, N2372);
or OR3 (N2399, N2380, N899, N1677);
xor XOR2 (N2400, N2396, N1230);
nor NOR3 (N2401, N2399, N122, N1213);
or OR3 (N2402, N2398, N802, N2095);
xor XOR2 (N2403, N2391, N1097);
nor NOR4 (N2404, N2397, N1761, N1251, N2289);
xor XOR2 (N2405, N2394, N1464);
xor XOR2 (N2406, N2405, N91);
nand NAND4 (N2407, N2400, N312, N304, N1231);
or OR2 (N2408, N2388, N933);
nand NAND4 (N2409, N2393, N1685, N2307, N267);
and AND2 (N2410, N2406, N2023);
xor XOR2 (N2411, N2409, N1146);
xor XOR2 (N2412, N2403, N463);
xor XOR2 (N2413, N2412, N739);
not NOT1 (N2414, N2413);
xor XOR2 (N2415, N2407, N1162);
not NOT1 (N2416, N2383);
xor XOR2 (N2417, N2414, N2092);
nor NOR2 (N2418, N2408, N1866);
nand NAND4 (N2419, N2381, N2097, N1593, N2276);
or OR2 (N2420, N2411, N1984);
xor XOR2 (N2421, N2415, N1082);
xor XOR2 (N2422, N2418, N2324);
or OR4 (N2423, N2417, N431, N1516, N1077);
and AND4 (N2424, N2410, N1097, N633, N1546);
or OR2 (N2425, N2421, N571);
not NOT1 (N2426, N2416);
nor NOR2 (N2427, N2422, N1250);
or OR3 (N2428, N2423, N171, N82);
and AND2 (N2429, N2402, N1923);
not NOT1 (N2430, N2401);
xor XOR2 (N2431, N2420, N900);
buf BUF1 (N2432, N2425);
xor XOR2 (N2433, N2404, N1524);
xor XOR2 (N2434, N2424, N2007);
buf BUF1 (N2435, N2426);
nand NAND4 (N2436, N2427, N323, N21, N934);
not NOT1 (N2437, N2428);
xor XOR2 (N2438, N2435, N1651);
and AND4 (N2439, N2432, N281, N1841, N1585);
nor NOR2 (N2440, N2439, N736);
nand NAND4 (N2441, N2440, N2227, N2295, N685);
nor NOR2 (N2442, N2429, N1676);
not NOT1 (N2443, N2431);
xor XOR2 (N2444, N2436, N1350);
or OR2 (N2445, N2430, N1828);
or OR3 (N2446, N2443, N1146, N605);
or OR2 (N2447, N2446, N2122);
nand NAND4 (N2448, N2444, N951, N56, N432);
and AND4 (N2449, N2433, N31, N186, N619);
and AND3 (N2450, N2434, N2070, N2018);
nor NOR4 (N2451, N2441, N1574, N1424, N1055);
or OR3 (N2452, N2442, N1356, N16);
nand NAND4 (N2453, N2450, N1369, N347, N132);
xor XOR2 (N2454, N2453, N1403);
nor NOR4 (N2455, N2449, N1869, N365, N248);
xor XOR2 (N2456, N2419, N705);
or OR2 (N2457, N2448, N842);
buf BUF1 (N2458, N2451);
nand NAND3 (N2459, N2457, N1058, N2405);
nand NAND4 (N2460, N2445, N1738, N2397, N835);
buf BUF1 (N2461, N2460);
not NOT1 (N2462, N2459);
nor NOR3 (N2463, N2455, N755, N249);
nor NOR4 (N2464, N2462, N1884, N341, N1458);
or OR4 (N2465, N2463, N2306, N1795, N2391);
nand NAND4 (N2466, N2461, N2260, N945, N2);
nor NOR3 (N2467, N2466, N126, N2368);
and AND3 (N2468, N2438, N1330, N95);
nor NOR3 (N2469, N2468, N2231, N1579);
and AND4 (N2470, N2458, N1653, N709, N990);
nor NOR2 (N2471, N2447, N1098);
xor XOR2 (N2472, N2456, N2025);
nor NOR3 (N2473, N2454, N1327, N1089);
buf BUF1 (N2474, N2452);
nor NOR4 (N2475, N2474, N1213, N1071, N2108);
and AND4 (N2476, N2437, N1603, N1135, N1913);
not NOT1 (N2477, N2464);
xor XOR2 (N2478, N2470, N1964);
xor XOR2 (N2479, N2473, N2345);
and AND4 (N2480, N2467, N563, N731, N2062);
xor XOR2 (N2481, N2480, N1292);
or OR2 (N2482, N2479, N2329);
nand NAND2 (N2483, N2471, N228);
nor NOR3 (N2484, N2469, N369, N1271);
or OR4 (N2485, N2482, N60, N685, N2128);
not NOT1 (N2486, N2484);
nand NAND2 (N2487, N2485, N493);
xor XOR2 (N2488, N2475, N643);
or OR2 (N2489, N2476, N957);
nor NOR3 (N2490, N2481, N1484, N1756);
xor XOR2 (N2491, N2465, N70);
not NOT1 (N2492, N2489);
nor NOR4 (N2493, N2477, N857, N691, N570);
xor XOR2 (N2494, N2490, N2169);
xor XOR2 (N2495, N2494, N32);
not NOT1 (N2496, N2488);
buf BUF1 (N2497, N2483);
buf BUF1 (N2498, N2486);
or OR3 (N2499, N2478, N2369, N1856);
xor XOR2 (N2500, N2499, N1767);
and AND2 (N2501, N2487, N366);
and AND3 (N2502, N2498, N1952, N1875);
nand NAND3 (N2503, N2492, N2117, N1799);
or OR3 (N2504, N2491, N1579, N1797);
nor NOR3 (N2505, N2495, N1810, N1616);
not NOT1 (N2506, N2472);
not NOT1 (N2507, N2493);
or OR4 (N2508, N2502, N2268, N1204, N928);
xor XOR2 (N2509, N2508, N1535);
nor NOR2 (N2510, N2507, N246);
and AND2 (N2511, N2506, N1287);
nand NAND2 (N2512, N2500, N28);
buf BUF1 (N2513, N2496);
and AND3 (N2514, N2501, N2412, N1189);
nand NAND3 (N2515, N2505, N162, N91);
or OR2 (N2516, N2514, N857);
xor XOR2 (N2517, N2509, N2040);
buf BUF1 (N2518, N2511);
endmodule