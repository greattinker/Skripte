// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N809,N819,N817,N812,N816,N801,N818,N807,N791,N820;

buf BUF1 (N21, N16);
or OR2 (N22, N5, N20);
not NOT1 (N23, N13);
nor NOR2 (N24, N4, N13);
xor XOR2 (N25, N10, N19);
buf BUF1 (N26, N20);
or OR4 (N27, N10, N6, N23, N12);
buf BUF1 (N28, N1);
not NOT1 (N29, N19);
not NOT1 (N30, N25);
or OR4 (N31, N24, N9, N24, N28);
xor XOR2 (N32, N12, N9);
xor XOR2 (N33, N26, N6);
xor XOR2 (N34, N2, N16);
buf BUF1 (N35, N17);
and AND4 (N36, N27, N13, N34, N15);
and AND2 (N37, N5, N32);
and AND3 (N38, N6, N10, N24);
nor NOR2 (N39, N33, N30);
or OR3 (N40, N26, N19, N1);
or OR3 (N41, N39, N20, N28);
xor XOR2 (N42, N36, N23);
and AND3 (N43, N21, N16, N18);
buf BUF1 (N44, N40);
nand NAND2 (N45, N22, N25);
buf BUF1 (N46, N31);
nor NOR2 (N47, N41, N35);
and AND4 (N48, N18, N1, N12, N9);
not NOT1 (N49, N37);
and AND4 (N50, N48, N35, N4, N6);
or OR2 (N51, N42, N6);
buf BUF1 (N52, N51);
not NOT1 (N53, N29);
nand NAND3 (N54, N38, N23, N1);
xor XOR2 (N55, N52, N4);
xor XOR2 (N56, N55, N44);
and AND3 (N57, N51, N9, N34);
xor XOR2 (N58, N46, N22);
or OR2 (N59, N45, N32);
and AND4 (N60, N54, N59, N54, N23);
or OR2 (N61, N45, N5);
nand NAND4 (N62, N60, N6, N21, N34);
nor NOR2 (N63, N49, N46);
not NOT1 (N64, N56);
or OR3 (N65, N53, N7, N60);
nor NOR3 (N66, N65, N10, N33);
or OR2 (N67, N63, N28);
not NOT1 (N68, N43);
nor NOR4 (N69, N68, N36, N42, N21);
and AND2 (N70, N64, N26);
nor NOR4 (N71, N70, N35, N36, N44);
and AND4 (N72, N57, N56, N18, N11);
or OR2 (N73, N50, N43);
nor NOR2 (N74, N58, N19);
or OR2 (N75, N74, N69);
nand NAND3 (N76, N7, N49, N64);
xor XOR2 (N77, N71, N18);
not NOT1 (N78, N77);
nor NOR2 (N79, N61, N63);
and AND4 (N80, N78, N26, N3, N70);
buf BUF1 (N81, N72);
nor NOR2 (N82, N47, N5);
buf BUF1 (N83, N73);
and AND4 (N84, N81, N51, N19, N43);
nor NOR4 (N85, N66, N51, N74, N48);
nor NOR4 (N86, N76, N59, N11, N14);
xor XOR2 (N87, N80, N50);
or OR2 (N88, N62, N44);
and AND3 (N89, N84, N35, N75);
or OR4 (N90, N59, N12, N61, N10);
not NOT1 (N91, N79);
or OR4 (N92, N90, N64, N46, N88);
buf BUF1 (N93, N4);
nand NAND2 (N94, N83, N7);
nor NOR2 (N95, N93, N81);
not NOT1 (N96, N94);
not NOT1 (N97, N82);
xor XOR2 (N98, N95, N85);
not NOT1 (N99, N58);
buf BUF1 (N100, N86);
not NOT1 (N101, N87);
and AND3 (N102, N98, N99, N83);
xor XOR2 (N103, N43, N69);
nand NAND2 (N104, N101, N20);
not NOT1 (N105, N104);
not NOT1 (N106, N89);
nand NAND3 (N107, N97, N52, N14);
buf BUF1 (N108, N91);
xor XOR2 (N109, N108, N30);
nor NOR3 (N110, N96, N63, N97);
buf BUF1 (N111, N107);
or OR2 (N112, N102, N52);
not NOT1 (N113, N109);
buf BUF1 (N114, N110);
or OR4 (N115, N92, N87, N31, N69);
not NOT1 (N116, N112);
xor XOR2 (N117, N67, N25);
xor XOR2 (N118, N106, N104);
nor NOR2 (N119, N100, N98);
buf BUF1 (N120, N103);
not NOT1 (N121, N111);
xor XOR2 (N122, N119, N2);
nand NAND4 (N123, N121, N114, N72, N75);
xor XOR2 (N124, N95, N61);
buf BUF1 (N125, N113);
and AND2 (N126, N122, N12);
nand NAND4 (N127, N115, N105, N108, N19);
buf BUF1 (N128, N42);
xor XOR2 (N129, N118, N65);
or OR3 (N130, N127, N82, N2);
nor NOR4 (N131, N128, N99, N60, N104);
or OR2 (N132, N124, N113);
or OR4 (N133, N130, N74, N71, N68);
or OR4 (N134, N131, N88, N61, N66);
and AND2 (N135, N116, N115);
not NOT1 (N136, N133);
and AND4 (N137, N126, N71, N21, N124);
not NOT1 (N138, N123);
buf BUF1 (N139, N129);
nand NAND2 (N140, N135, N109);
and AND3 (N141, N125, N122, N20);
nor NOR2 (N142, N134, N88);
and AND4 (N143, N136, N55, N91, N103);
nand NAND3 (N144, N120, N128, N105);
not NOT1 (N145, N140);
buf BUF1 (N146, N138);
buf BUF1 (N147, N146);
buf BUF1 (N148, N132);
or OR4 (N149, N143, N74, N76, N118);
xor XOR2 (N150, N137, N14);
not NOT1 (N151, N149);
buf BUF1 (N152, N141);
xor XOR2 (N153, N152, N124);
and AND3 (N154, N144, N80, N61);
nand NAND4 (N155, N153, N111, N139, N34);
nand NAND2 (N156, N133, N63);
or OR3 (N157, N147, N32, N1);
not NOT1 (N158, N117);
nand NAND3 (N159, N150, N64, N108);
or OR2 (N160, N151, N109);
nand NAND4 (N161, N154, N112, N24, N17);
nor NOR3 (N162, N157, N27, N142);
nand NAND3 (N163, N143, N10, N155);
xor XOR2 (N164, N117, N110);
nor NOR4 (N165, N145, N138, N75, N44);
nor NOR3 (N166, N158, N63, N152);
nor NOR3 (N167, N162, N64, N119);
and AND2 (N168, N167, N42);
not NOT1 (N169, N165);
and AND3 (N170, N168, N140, N48);
and AND3 (N171, N148, N122, N7);
nor NOR4 (N172, N166, N103, N72, N53);
or OR3 (N173, N161, N152, N125);
or OR2 (N174, N170, N22);
xor XOR2 (N175, N156, N121);
nor NOR2 (N176, N172, N160);
nand NAND4 (N177, N113, N90, N32, N62);
buf BUF1 (N178, N164);
nand NAND2 (N179, N176, N170);
and AND3 (N180, N177, N124, N157);
or OR4 (N181, N163, N162, N143, N22);
buf BUF1 (N182, N181);
buf BUF1 (N183, N178);
not NOT1 (N184, N159);
and AND3 (N185, N180, N133, N78);
nand NAND4 (N186, N174, N58, N78, N28);
or OR2 (N187, N185, N162);
buf BUF1 (N188, N182);
or OR4 (N189, N188, N110, N72, N111);
not NOT1 (N190, N169);
nand NAND3 (N191, N171, N59, N103);
xor XOR2 (N192, N190, N15);
xor XOR2 (N193, N192, N90);
xor XOR2 (N194, N183, N122);
or OR2 (N195, N175, N191);
nor NOR2 (N196, N70, N117);
not NOT1 (N197, N184);
or OR4 (N198, N197, N70, N23, N28);
and AND2 (N199, N173, N93);
nand NAND4 (N200, N187, N69, N70, N5);
buf BUF1 (N201, N200);
not NOT1 (N202, N179);
nand NAND4 (N203, N198, N63, N95, N128);
or OR3 (N204, N202, N185, N130);
or OR2 (N205, N199, N34);
nor NOR2 (N206, N189, N11);
nand NAND2 (N207, N204, N160);
nand NAND2 (N208, N205, N152);
nand NAND4 (N209, N207, N100, N91, N193);
nor NOR4 (N210, N147, N77, N12, N82);
nor NOR2 (N211, N195, N78);
and AND4 (N212, N196, N7, N61, N27);
nor NOR2 (N213, N208, N185);
xor XOR2 (N214, N213, N50);
nand NAND4 (N215, N206, N104, N84, N155);
xor XOR2 (N216, N211, N203);
xor XOR2 (N217, N121, N207);
xor XOR2 (N218, N216, N49);
not NOT1 (N219, N201);
or OR2 (N220, N217, N138);
and AND3 (N221, N186, N20, N165);
or OR3 (N222, N194, N155, N210);
and AND4 (N223, N10, N114, N102, N66);
buf BUF1 (N224, N219);
or OR4 (N225, N214, N114, N38, N194);
xor XOR2 (N226, N209, N85);
not NOT1 (N227, N223);
nand NAND2 (N228, N227, N56);
not NOT1 (N229, N221);
xor XOR2 (N230, N215, N70);
and AND4 (N231, N220, N188, N183, N100);
or OR3 (N232, N222, N10, N192);
buf BUF1 (N233, N225);
nor NOR4 (N234, N230, N215, N124, N213);
buf BUF1 (N235, N218);
or OR2 (N236, N229, N11);
or OR4 (N237, N226, N8, N17, N189);
buf BUF1 (N238, N236);
nand NAND4 (N239, N235, N18, N79, N200);
and AND3 (N240, N237, N139, N128);
nor NOR2 (N241, N234, N161);
nor NOR3 (N242, N238, N123, N213);
not NOT1 (N243, N231);
nand NAND2 (N244, N232, N80);
nor NOR4 (N245, N242, N81, N230, N244);
not NOT1 (N246, N108);
nand NAND4 (N247, N228, N33, N177, N165);
not NOT1 (N248, N212);
nor NOR3 (N249, N241, N190, N186);
xor XOR2 (N250, N249, N244);
not NOT1 (N251, N248);
xor XOR2 (N252, N251, N79);
xor XOR2 (N253, N224, N33);
xor XOR2 (N254, N240, N145);
not NOT1 (N255, N233);
not NOT1 (N256, N250);
and AND2 (N257, N245, N168);
nor NOR3 (N258, N239, N80, N146);
and AND4 (N259, N255, N164, N257, N20);
nor NOR2 (N260, N233, N94);
nand NAND4 (N261, N254, N137, N240, N230);
buf BUF1 (N262, N252);
nor NOR3 (N263, N260, N12, N210);
buf BUF1 (N264, N243);
and AND3 (N265, N261, N111, N127);
or OR3 (N266, N253, N202, N227);
nor NOR2 (N267, N263, N46);
nor NOR3 (N268, N246, N80, N246);
nand NAND2 (N269, N262, N52);
buf BUF1 (N270, N256);
xor XOR2 (N271, N265, N254);
and AND4 (N272, N271, N240, N166, N233);
nor NOR2 (N273, N272, N173);
nor NOR2 (N274, N259, N122);
and AND2 (N275, N274, N226);
not NOT1 (N276, N273);
not NOT1 (N277, N267);
not NOT1 (N278, N266);
nand NAND4 (N279, N276, N64, N43, N47);
nor NOR2 (N280, N269, N68);
nand NAND3 (N281, N277, N109, N245);
buf BUF1 (N282, N281);
nor NOR2 (N283, N270, N70);
and AND4 (N284, N280, N276, N102, N268);
nor NOR2 (N285, N112, N49);
nand NAND3 (N286, N283, N222, N116);
xor XOR2 (N287, N278, N1);
not NOT1 (N288, N264);
buf BUF1 (N289, N258);
or OR4 (N290, N285, N279, N278, N104);
or OR3 (N291, N283, N186, N44);
nand NAND3 (N292, N287, N41, N130);
nand NAND2 (N293, N290, N59);
xor XOR2 (N294, N292, N182);
not NOT1 (N295, N247);
nand NAND2 (N296, N293, N85);
nor NOR3 (N297, N284, N19, N15);
not NOT1 (N298, N288);
buf BUF1 (N299, N297);
not NOT1 (N300, N294);
buf BUF1 (N301, N289);
xor XOR2 (N302, N295, N255);
nand NAND2 (N303, N301, N204);
nand NAND3 (N304, N296, N129, N227);
buf BUF1 (N305, N298);
buf BUF1 (N306, N299);
buf BUF1 (N307, N275);
xor XOR2 (N308, N282, N217);
buf BUF1 (N309, N291);
buf BUF1 (N310, N304);
and AND3 (N311, N307, N85, N11);
nor NOR2 (N312, N310, N226);
xor XOR2 (N313, N312, N108);
buf BUF1 (N314, N313);
buf BUF1 (N315, N314);
or OR2 (N316, N302, N187);
not NOT1 (N317, N309);
and AND4 (N318, N300, N173, N64, N305);
nor NOR3 (N319, N7, N173, N148);
or OR4 (N320, N286, N307, N47, N272);
or OR2 (N321, N311, N134);
or OR3 (N322, N319, N220, N236);
buf BUF1 (N323, N303);
not NOT1 (N324, N308);
not NOT1 (N325, N317);
nand NAND2 (N326, N316, N127);
nand NAND2 (N327, N324, N98);
not NOT1 (N328, N320);
xor XOR2 (N329, N327, N266);
not NOT1 (N330, N328);
xor XOR2 (N331, N323, N138);
nor NOR2 (N332, N315, N130);
not NOT1 (N333, N330);
xor XOR2 (N334, N331, N25);
and AND2 (N335, N333, N183);
not NOT1 (N336, N332);
or OR4 (N337, N326, N246, N321, N48);
nor NOR2 (N338, N21, N164);
nand NAND4 (N339, N329, N136, N338, N313);
not NOT1 (N340, N70);
and AND3 (N341, N334, N210, N20);
buf BUF1 (N342, N337);
not NOT1 (N343, N341);
and AND3 (N344, N318, N137, N108);
buf BUF1 (N345, N344);
not NOT1 (N346, N345);
nand NAND4 (N347, N340, N226, N314, N331);
nor NOR4 (N348, N325, N315, N325, N214);
or OR3 (N349, N322, N322, N283);
xor XOR2 (N350, N342, N12);
nand NAND3 (N351, N349, N151, N258);
nor NOR3 (N352, N306, N263, N238);
and AND2 (N353, N352, N78);
nand NAND4 (N354, N339, N62, N174, N15);
or OR3 (N355, N350, N279, N326);
nand NAND2 (N356, N335, N127);
nand NAND3 (N357, N356, N321, N220);
nand NAND2 (N358, N357, N209);
nor NOR3 (N359, N351, N152, N78);
nand NAND4 (N360, N347, N251, N185, N100);
nor NOR2 (N361, N348, N11);
or OR3 (N362, N353, N282, N151);
and AND3 (N363, N336, N38, N157);
or OR3 (N364, N358, N249, N207);
buf BUF1 (N365, N362);
nor NOR2 (N366, N363, N24);
or OR4 (N367, N346, N229, N115, N290);
xor XOR2 (N368, N343, N100);
buf BUF1 (N369, N361);
or OR4 (N370, N359, N350, N294, N184);
buf BUF1 (N371, N367);
nor NOR3 (N372, N355, N92, N277);
not NOT1 (N373, N354);
not NOT1 (N374, N369);
or OR2 (N375, N370, N57);
nand NAND2 (N376, N372, N367);
nand NAND4 (N377, N364, N323, N121, N231);
and AND2 (N378, N360, N281);
not NOT1 (N379, N378);
and AND2 (N380, N377, N185);
nor NOR4 (N381, N376, N312, N350, N96);
xor XOR2 (N382, N366, N6);
buf BUF1 (N383, N381);
xor XOR2 (N384, N368, N47);
or OR4 (N385, N375, N47, N208, N340);
xor XOR2 (N386, N380, N14);
not NOT1 (N387, N371);
nand NAND4 (N388, N374, N290, N205, N199);
nor NOR2 (N389, N383, N210);
buf BUF1 (N390, N388);
or OR2 (N391, N389, N179);
and AND4 (N392, N373, N387, N169, N113);
and AND2 (N393, N324, N350);
or OR3 (N394, N382, N241, N202);
xor XOR2 (N395, N391, N113);
buf BUF1 (N396, N393);
nor NOR4 (N397, N396, N205, N239, N134);
nor NOR4 (N398, N365, N273, N205, N53);
and AND4 (N399, N392, N321, N191, N111);
nor NOR2 (N400, N386, N33);
not NOT1 (N401, N394);
nand NAND4 (N402, N384, N27, N309, N156);
nand NAND2 (N403, N402, N43);
or OR4 (N404, N403, N109, N174, N124);
and AND4 (N405, N398, N15, N199, N260);
or OR2 (N406, N404, N294);
nor NOR2 (N407, N401, N373);
or OR4 (N408, N405, N180, N230, N34);
buf BUF1 (N409, N385);
or OR4 (N410, N397, N350, N180, N191);
and AND2 (N411, N406, N27);
nor NOR4 (N412, N410, N97, N228, N315);
nand NAND3 (N413, N409, N362, N65);
buf BUF1 (N414, N395);
nor NOR4 (N415, N407, N50, N121, N26);
or OR4 (N416, N412, N33, N122, N201);
not NOT1 (N417, N416);
not NOT1 (N418, N399);
or OR3 (N419, N414, N264, N64);
buf BUF1 (N420, N400);
nor NOR2 (N421, N413, N151);
or OR4 (N422, N420, N257, N393, N91);
not NOT1 (N423, N422);
and AND3 (N424, N390, N165, N122);
buf BUF1 (N425, N415);
buf BUF1 (N426, N418);
xor XOR2 (N427, N408, N169);
and AND4 (N428, N411, N74, N216, N106);
buf BUF1 (N429, N417);
buf BUF1 (N430, N423);
xor XOR2 (N431, N424, N163);
nor NOR4 (N432, N425, N409, N31, N153);
and AND2 (N433, N430, N294);
xor XOR2 (N434, N432, N330);
or OR2 (N435, N379, N367);
buf BUF1 (N436, N429);
not NOT1 (N437, N431);
not NOT1 (N438, N435);
buf BUF1 (N439, N434);
and AND3 (N440, N433, N142, N46);
and AND4 (N441, N426, N50, N176, N378);
or OR3 (N442, N436, N303, N316);
or OR4 (N443, N442, N354, N405, N132);
nor NOR2 (N444, N437, N200);
and AND2 (N445, N428, N389);
and AND4 (N446, N419, N27, N393, N267);
xor XOR2 (N447, N445, N67);
xor XOR2 (N448, N421, N258);
xor XOR2 (N449, N441, N339);
xor XOR2 (N450, N444, N115);
or OR2 (N451, N448, N219);
not NOT1 (N452, N440);
nor NOR3 (N453, N449, N87, N327);
nand NAND4 (N454, N451, N447, N231, N377);
xor XOR2 (N455, N165, N247);
xor XOR2 (N456, N443, N101);
not NOT1 (N457, N450);
not NOT1 (N458, N455);
not NOT1 (N459, N453);
and AND4 (N460, N457, N92, N78, N74);
buf BUF1 (N461, N446);
and AND4 (N462, N454, N361, N227, N339);
not NOT1 (N463, N458);
nor NOR4 (N464, N438, N346, N443, N402);
buf BUF1 (N465, N460);
nand NAND2 (N466, N459, N80);
and AND2 (N467, N427, N428);
or OR2 (N468, N467, N337);
xor XOR2 (N469, N465, N347);
nor NOR2 (N470, N468, N252);
not NOT1 (N471, N464);
and AND4 (N472, N439, N333, N50, N386);
xor XOR2 (N473, N470, N332);
or OR4 (N474, N466, N453, N311, N310);
not NOT1 (N475, N473);
or OR3 (N476, N472, N421, N131);
not NOT1 (N477, N462);
nand NAND4 (N478, N452, N220, N448, N415);
or OR3 (N479, N477, N217, N163);
and AND4 (N480, N463, N290, N264, N248);
nand NAND3 (N481, N456, N42, N439);
nor NOR4 (N482, N471, N232, N441, N297);
nor NOR4 (N483, N461, N283, N241, N393);
nand NAND2 (N484, N479, N103);
not NOT1 (N485, N478);
not NOT1 (N486, N482);
nor NOR2 (N487, N469, N450);
xor XOR2 (N488, N486, N468);
nor NOR3 (N489, N474, N259, N262);
nand NAND2 (N490, N475, N51);
xor XOR2 (N491, N481, N350);
not NOT1 (N492, N489);
or OR2 (N493, N492, N104);
buf BUF1 (N494, N487);
or OR2 (N495, N494, N332);
xor XOR2 (N496, N488, N416);
xor XOR2 (N497, N476, N111);
nor NOR3 (N498, N493, N260, N12);
nand NAND2 (N499, N480, N457);
nand NAND4 (N500, N490, N421, N421, N36);
not NOT1 (N501, N484);
nand NAND4 (N502, N498, N68, N136, N33);
buf BUF1 (N503, N500);
buf BUF1 (N504, N499);
not NOT1 (N505, N497);
nor NOR4 (N506, N483, N71, N267, N143);
nand NAND3 (N507, N506, N425, N287);
and AND4 (N508, N495, N117, N166, N468);
or OR2 (N509, N502, N469);
and AND3 (N510, N503, N319, N478);
not NOT1 (N511, N504);
xor XOR2 (N512, N510, N486);
or OR2 (N513, N508, N20);
nor NOR3 (N514, N513, N422, N490);
nor NOR2 (N515, N514, N362);
or OR3 (N516, N501, N26, N73);
not NOT1 (N517, N505);
buf BUF1 (N518, N515);
buf BUF1 (N519, N517);
not NOT1 (N520, N518);
buf BUF1 (N521, N512);
or OR2 (N522, N496, N285);
xor XOR2 (N523, N491, N260);
and AND2 (N524, N485, N26);
buf BUF1 (N525, N523);
buf BUF1 (N526, N522);
xor XOR2 (N527, N526, N329);
xor XOR2 (N528, N521, N519);
buf BUF1 (N529, N161);
buf BUF1 (N530, N529);
xor XOR2 (N531, N530, N338);
buf BUF1 (N532, N525);
or OR3 (N533, N509, N520, N356);
xor XOR2 (N534, N53, N132);
nand NAND3 (N535, N531, N276, N378);
and AND3 (N536, N535, N332, N119);
xor XOR2 (N537, N533, N364);
and AND3 (N538, N536, N261, N370);
xor XOR2 (N539, N538, N330);
nand NAND2 (N540, N537, N345);
not NOT1 (N541, N507);
not NOT1 (N542, N516);
and AND2 (N543, N532, N309);
xor XOR2 (N544, N511, N425);
xor XOR2 (N545, N527, N417);
and AND4 (N546, N539, N233, N266, N307);
not NOT1 (N547, N545);
and AND3 (N548, N534, N132, N531);
and AND2 (N549, N543, N497);
and AND2 (N550, N547, N174);
nand NAND2 (N551, N541, N72);
not NOT1 (N552, N524);
nor NOR2 (N553, N551, N31);
nor NOR4 (N554, N542, N87, N327, N545);
xor XOR2 (N555, N528, N472);
or OR2 (N556, N548, N136);
and AND4 (N557, N553, N514, N373, N324);
nor NOR3 (N558, N556, N545, N381);
xor XOR2 (N559, N549, N266);
and AND2 (N560, N555, N92);
buf BUF1 (N561, N560);
nand NAND4 (N562, N559, N316, N125, N205);
nand NAND4 (N563, N561, N99, N431, N527);
or OR3 (N564, N552, N267, N407);
nand NAND4 (N565, N562, N562, N55, N261);
and AND3 (N566, N544, N394, N533);
nor NOR4 (N567, N563, N141, N386, N100);
nor NOR3 (N568, N567, N426, N385);
or OR2 (N569, N564, N482);
not NOT1 (N570, N569);
nor NOR3 (N571, N566, N412, N408);
and AND4 (N572, N571, N566, N12, N300);
nor NOR4 (N573, N550, N314, N475, N566);
xor XOR2 (N574, N565, N264);
not NOT1 (N575, N574);
buf BUF1 (N576, N557);
not NOT1 (N577, N568);
or OR2 (N578, N540, N538);
nor NOR4 (N579, N558, N496, N564, N142);
and AND4 (N580, N578, N233, N545, N455);
nor NOR3 (N581, N546, N270, N435);
and AND4 (N582, N573, N407, N2, N491);
not NOT1 (N583, N575);
or OR4 (N584, N577, N207, N274, N561);
and AND4 (N585, N554, N61, N29, N20);
nor NOR2 (N586, N584, N175);
nand NAND2 (N587, N581, N438);
buf BUF1 (N588, N586);
nand NAND2 (N589, N572, N243);
xor XOR2 (N590, N582, N58);
and AND4 (N591, N588, N236, N181, N365);
xor XOR2 (N592, N570, N370);
or OR2 (N593, N576, N503);
not NOT1 (N594, N585);
nand NAND4 (N595, N591, N322, N355, N256);
and AND4 (N596, N594, N551, N157, N359);
nor NOR4 (N597, N596, N468, N435, N112);
nand NAND2 (N598, N587, N460);
not NOT1 (N599, N590);
nand NAND4 (N600, N583, N10, N581, N476);
not NOT1 (N601, N592);
nand NAND4 (N602, N601, N537, N291, N25);
buf BUF1 (N603, N600);
or OR4 (N604, N599, N555, N204, N530);
xor XOR2 (N605, N597, N201);
or OR2 (N606, N589, N143);
and AND2 (N607, N606, N80);
xor XOR2 (N608, N605, N298);
buf BUF1 (N609, N607);
nor NOR4 (N610, N593, N584, N67, N323);
nor NOR2 (N611, N595, N195);
and AND2 (N612, N604, N201);
nand NAND4 (N613, N612, N428, N31, N60);
buf BUF1 (N614, N611);
nor NOR4 (N615, N613, N599, N518, N430);
or OR4 (N616, N603, N234, N244, N343);
not NOT1 (N617, N609);
nand NAND2 (N618, N614, N435);
not NOT1 (N619, N598);
nor NOR4 (N620, N608, N425, N447, N481);
and AND4 (N621, N617, N402, N151, N100);
nand NAND2 (N622, N602, N293);
nand NAND4 (N623, N616, N577, N297, N184);
nor NOR3 (N624, N580, N342, N139);
nand NAND3 (N625, N579, N124, N582);
nand NAND4 (N626, N619, N339, N231, N58);
nor NOR3 (N627, N622, N156, N10);
xor XOR2 (N628, N627, N435);
or OR4 (N629, N615, N327, N397, N55);
or OR2 (N630, N626, N355);
and AND4 (N631, N618, N341, N352, N340);
nor NOR3 (N632, N624, N520, N562);
and AND4 (N633, N628, N280, N1, N474);
xor XOR2 (N634, N610, N35);
or OR3 (N635, N620, N314, N493);
xor XOR2 (N636, N633, N487);
nor NOR3 (N637, N632, N351, N314);
and AND4 (N638, N636, N544, N458, N94);
nor NOR3 (N639, N634, N23, N546);
nor NOR2 (N640, N625, N426);
xor XOR2 (N641, N635, N548);
xor XOR2 (N642, N623, N379);
nand NAND4 (N643, N629, N474, N564, N579);
or OR3 (N644, N630, N62, N237);
and AND2 (N645, N644, N75);
nor NOR4 (N646, N639, N75, N196, N431);
buf BUF1 (N647, N646);
nand NAND4 (N648, N638, N79, N236, N275);
and AND3 (N649, N631, N461, N636);
not NOT1 (N650, N645);
and AND4 (N651, N621, N595, N185, N287);
not NOT1 (N652, N649);
nand NAND4 (N653, N637, N461, N382, N239);
or OR2 (N654, N643, N278);
nor NOR4 (N655, N654, N152, N397, N468);
buf BUF1 (N656, N652);
buf BUF1 (N657, N655);
buf BUF1 (N658, N656);
or OR2 (N659, N642, N552);
xor XOR2 (N660, N658, N373);
or OR4 (N661, N653, N61, N64, N551);
nand NAND4 (N662, N660, N287, N223, N455);
not NOT1 (N663, N651);
and AND2 (N664, N648, N112);
buf BUF1 (N665, N650);
or OR3 (N666, N641, N521, N317);
not NOT1 (N667, N665);
or OR3 (N668, N657, N57, N417);
and AND2 (N669, N659, N131);
buf BUF1 (N670, N647);
and AND4 (N671, N667, N232, N646, N212);
xor XOR2 (N672, N661, N288);
and AND4 (N673, N664, N129, N141, N121);
buf BUF1 (N674, N670);
xor XOR2 (N675, N671, N249);
xor XOR2 (N676, N669, N75);
nor NOR3 (N677, N674, N573, N420);
xor XOR2 (N678, N666, N632);
nor NOR3 (N679, N677, N678, N317);
buf BUF1 (N680, N202);
buf BUF1 (N681, N679);
and AND3 (N682, N673, N440, N30);
and AND3 (N683, N681, N678, N534);
buf BUF1 (N684, N640);
nand NAND4 (N685, N668, N669, N665, N392);
buf BUF1 (N686, N672);
buf BUF1 (N687, N680);
buf BUF1 (N688, N663);
buf BUF1 (N689, N684);
xor XOR2 (N690, N686, N401);
nand NAND3 (N691, N683, N626, N181);
xor XOR2 (N692, N675, N285);
buf BUF1 (N693, N690);
nor NOR3 (N694, N662, N317, N365);
buf BUF1 (N695, N682);
and AND2 (N696, N691, N163);
nor NOR3 (N697, N688, N22, N371);
nand NAND4 (N698, N693, N653, N334, N579);
nand NAND3 (N699, N698, N566, N274);
and AND4 (N700, N692, N97, N204, N336);
not NOT1 (N701, N689);
nor NOR2 (N702, N696, N187);
nor NOR2 (N703, N697, N79);
nor NOR4 (N704, N687, N166, N92, N438);
not NOT1 (N705, N702);
nor NOR4 (N706, N685, N45, N648, N544);
and AND3 (N707, N700, N30, N216);
buf BUF1 (N708, N703);
nand NAND4 (N709, N676, N619, N494, N364);
nor NOR4 (N710, N694, N175, N282, N530);
not NOT1 (N711, N704);
nor NOR3 (N712, N695, N360, N493);
nand NAND4 (N713, N699, N108, N290, N125);
nand NAND4 (N714, N711, N202, N273, N355);
or OR2 (N715, N714, N486);
buf BUF1 (N716, N705);
not NOT1 (N717, N716);
not NOT1 (N718, N717);
xor XOR2 (N719, N708, N535);
xor XOR2 (N720, N706, N291);
and AND4 (N721, N718, N68, N139, N190);
buf BUF1 (N722, N721);
or OR2 (N723, N707, N214);
xor XOR2 (N724, N719, N685);
not NOT1 (N725, N709);
or OR3 (N726, N722, N209, N118);
or OR2 (N727, N710, N697);
nor NOR3 (N728, N715, N491, N324);
or OR3 (N729, N701, N410, N607);
not NOT1 (N730, N720);
or OR4 (N731, N723, N613, N706, N23);
nand NAND3 (N732, N725, N335, N163);
nand NAND4 (N733, N732, N146, N441, N230);
and AND2 (N734, N712, N141);
and AND2 (N735, N727, N202);
nor NOR2 (N736, N713, N379);
or OR3 (N737, N734, N151, N2);
nand NAND3 (N738, N726, N581, N220);
xor XOR2 (N739, N724, N334);
or OR4 (N740, N728, N238, N313, N5);
nor NOR4 (N741, N740, N492, N507, N720);
nor NOR3 (N742, N739, N711, N71);
and AND4 (N743, N741, N629, N193, N645);
nor NOR3 (N744, N743, N152, N609);
nor NOR4 (N745, N742, N304, N300, N401);
nand NAND4 (N746, N735, N660, N434, N221);
not NOT1 (N747, N744);
nand NAND2 (N748, N736, N294);
nand NAND2 (N749, N738, N345);
not NOT1 (N750, N737);
nand NAND3 (N751, N733, N95, N102);
nand NAND4 (N752, N751, N2, N485, N534);
nand NAND3 (N753, N748, N255, N449);
or OR3 (N754, N749, N177, N333);
and AND3 (N755, N750, N637, N94);
and AND3 (N756, N752, N139, N23);
or OR4 (N757, N730, N210, N136, N558);
nand NAND2 (N758, N756, N275);
and AND3 (N759, N747, N679, N624);
nand NAND4 (N760, N757, N534, N532, N718);
nor NOR2 (N761, N746, N36);
nand NAND2 (N762, N745, N117);
nand NAND3 (N763, N762, N417, N337);
or OR3 (N764, N763, N151, N761);
and AND4 (N765, N438, N63, N286, N273);
nor NOR3 (N766, N731, N624, N175);
and AND4 (N767, N729, N485, N356, N422);
xor XOR2 (N768, N758, N557);
nand NAND3 (N769, N768, N266, N623);
not NOT1 (N770, N764);
nand NAND3 (N771, N754, N222, N394);
xor XOR2 (N772, N759, N507);
buf BUF1 (N773, N767);
xor XOR2 (N774, N765, N213);
or OR2 (N775, N770, N688);
or OR3 (N776, N766, N239, N565);
nand NAND3 (N777, N774, N592, N212);
nand NAND4 (N778, N772, N58, N700, N667);
xor XOR2 (N779, N776, N169);
not NOT1 (N780, N755);
and AND2 (N781, N780, N41);
not NOT1 (N782, N777);
not NOT1 (N783, N771);
buf BUF1 (N784, N778);
buf BUF1 (N785, N775);
and AND4 (N786, N779, N590, N330, N576);
and AND2 (N787, N785, N564);
nand NAND4 (N788, N773, N417, N748, N651);
not NOT1 (N789, N788);
nor NOR2 (N790, N781, N691);
or OR3 (N791, N787, N360, N340);
xor XOR2 (N792, N753, N601);
xor XOR2 (N793, N783, N300);
or OR3 (N794, N782, N690, N170);
or OR3 (N795, N792, N434, N19);
buf BUF1 (N796, N793);
not NOT1 (N797, N760);
xor XOR2 (N798, N796, N693);
nand NAND3 (N799, N794, N426, N670);
or OR3 (N800, N798, N386, N790);
and AND3 (N801, N525, N750, N556);
nand NAND3 (N802, N799, N11, N302);
or OR3 (N803, N795, N454, N514);
and AND3 (N804, N800, N484, N110);
buf BUF1 (N805, N769);
and AND4 (N806, N786, N64, N572, N743);
nor NOR3 (N807, N789, N724, N712);
and AND2 (N808, N784, N794);
xor XOR2 (N809, N797, N559);
and AND4 (N810, N802, N609, N565, N450);
not NOT1 (N811, N804);
nor NOR2 (N812, N808, N578);
nand NAND4 (N813, N806, N496, N388, N428);
nor NOR3 (N814, N810, N334, N512);
or OR2 (N815, N814, N155);
xor XOR2 (N816, N803, N665);
or OR3 (N817, N811, N532, N14);
not NOT1 (N818, N813);
or OR3 (N819, N805, N114, N204);
not NOT1 (N820, N815);
endmodule