// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N1600,N1613,N1618,N1617,N1610,N1585,N1616,N1596,N1619,N1620;

buf BUF1 (N21, N20);
not NOT1 (N22, N2);
nor NOR2 (N23, N2, N15);
nand NAND3 (N24, N22, N12, N9);
nor NOR4 (N25, N11, N6, N1, N16);
not NOT1 (N26, N8);
buf BUF1 (N27, N17);
not NOT1 (N28, N26);
nor NOR3 (N29, N3, N1, N16);
nand NAND2 (N30, N21, N23);
xor XOR2 (N31, N21, N16);
xor XOR2 (N32, N17, N5);
not NOT1 (N33, N27);
not NOT1 (N34, N32);
not NOT1 (N35, N2);
not NOT1 (N36, N32);
and AND3 (N37, N30, N5, N36);
xor XOR2 (N38, N6, N36);
not NOT1 (N39, N33);
xor XOR2 (N40, N31, N24);
nor NOR3 (N41, N34, N4, N18);
nor NOR4 (N42, N30, N11, N4, N6);
and AND2 (N43, N29, N19);
not NOT1 (N44, N38);
xor XOR2 (N45, N41, N9);
nor NOR2 (N46, N37, N1);
and AND4 (N47, N44, N37, N37, N3);
xor XOR2 (N48, N40, N18);
buf BUF1 (N49, N39);
nand NAND2 (N50, N42, N26);
not NOT1 (N51, N50);
nand NAND2 (N52, N48, N6);
nand NAND4 (N53, N45, N16, N34, N3);
buf BUF1 (N54, N35);
nand NAND2 (N55, N46, N51);
nand NAND2 (N56, N40, N9);
xor XOR2 (N57, N49, N48);
buf BUF1 (N58, N53);
and AND3 (N59, N57, N12, N6);
nor NOR4 (N60, N58, N23, N11, N9);
nor NOR3 (N61, N52, N15, N22);
buf BUF1 (N62, N60);
not NOT1 (N63, N47);
xor XOR2 (N64, N54, N37);
buf BUF1 (N65, N43);
or OR4 (N66, N65, N52, N41, N27);
nand NAND4 (N67, N56, N21, N5, N29);
and AND3 (N68, N28, N10, N38);
and AND2 (N69, N63, N3);
and AND4 (N70, N62, N9, N23, N11);
not NOT1 (N71, N69);
not NOT1 (N72, N64);
or OR4 (N73, N70, N70, N44, N18);
buf BUF1 (N74, N66);
not NOT1 (N75, N73);
xor XOR2 (N76, N67, N58);
nand NAND2 (N77, N25, N48);
and AND3 (N78, N61, N44, N54);
buf BUF1 (N79, N72);
nor NOR2 (N80, N76, N23);
nand NAND3 (N81, N59, N9, N6);
xor XOR2 (N82, N80, N16);
xor XOR2 (N83, N79, N65);
or OR4 (N84, N82, N31, N83, N47);
buf BUF1 (N85, N55);
not NOT1 (N86, N21);
and AND3 (N87, N85, N78, N51);
nor NOR3 (N88, N76, N66, N47);
or OR3 (N89, N81, N48, N49);
not NOT1 (N90, N86);
nor NOR4 (N91, N87, N18, N59, N67);
not NOT1 (N92, N68);
and AND2 (N93, N77, N51);
and AND2 (N94, N91, N24);
not NOT1 (N95, N71);
buf BUF1 (N96, N74);
or OR2 (N97, N96, N49);
xor XOR2 (N98, N92, N82);
nor NOR4 (N99, N84, N80, N4, N23);
or OR4 (N100, N75, N53, N17, N62);
nand NAND2 (N101, N98, N58);
nor NOR4 (N102, N89, N79, N15, N12);
buf BUF1 (N103, N100);
buf BUF1 (N104, N90);
buf BUF1 (N105, N99);
not NOT1 (N106, N94);
or OR4 (N107, N95, N84, N16, N41);
buf BUF1 (N108, N93);
nand NAND2 (N109, N107, N93);
buf BUF1 (N110, N103);
not NOT1 (N111, N88);
nor NOR4 (N112, N102, N29, N57, N3);
buf BUF1 (N113, N111);
xor XOR2 (N114, N104, N73);
nand NAND4 (N115, N109, N82, N41, N39);
nand NAND4 (N116, N108, N91, N5, N64);
nand NAND4 (N117, N106, N7, N29, N19);
and AND3 (N118, N101, N68, N116);
buf BUF1 (N119, N38);
and AND4 (N120, N97, N31, N45, N22);
or OR2 (N121, N112, N44);
xor XOR2 (N122, N117, N75);
and AND3 (N123, N121, N11, N120);
buf BUF1 (N124, N14);
buf BUF1 (N125, N124);
or OR4 (N126, N113, N18, N107, N2);
or OR2 (N127, N115, N45);
buf BUF1 (N128, N126);
xor XOR2 (N129, N127, N91);
or OR4 (N130, N119, N14, N26, N127);
xor XOR2 (N131, N122, N8);
buf BUF1 (N132, N128);
xor XOR2 (N133, N123, N69);
xor XOR2 (N134, N131, N94);
xor XOR2 (N135, N129, N85);
xor XOR2 (N136, N118, N75);
nand NAND4 (N137, N132, N80, N134, N92);
not NOT1 (N138, N111);
not NOT1 (N139, N105);
and AND2 (N140, N125, N35);
buf BUF1 (N141, N135);
and AND2 (N142, N137, N117);
and AND4 (N143, N110, N138, N15, N103);
xor XOR2 (N144, N120, N91);
nand NAND3 (N145, N142, N142, N1);
nand NAND2 (N146, N136, N128);
not NOT1 (N147, N139);
xor XOR2 (N148, N141, N8);
buf BUF1 (N149, N140);
nand NAND3 (N150, N147, N114, N116);
and AND3 (N151, N41, N110, N71);
xor XOR2 (N152, N133, N127);
and AND2 (N153, N152, N87);
nand NAND2 (N154, N144, N115);
nand NAND2 (N155, N146, N63);
xor XOR2 (N156, N150, N69);
nand NAND4 (N157, N155, N151, N87, N75);
nor NOR3 (N158, N150, N69, N140);
and AND2 (N159, N157, N3);
nor NOR2 (N160, N149, N80);
nand NAND2 (N161, N158, N155);
and AND4 (N162, N148, N59, N20, N126);
buf BUF1 (N163, N161);
and AND3 (N164, N159, N74, N13);
xor XOR2 (N165, N160, N154);
nand NAND2 (N166, N32, N52);
and AND3 (N167, N156, N59, N44);
nor NOR4 (N168, N164, N140, N13, N61);
nand NAND2 (N169, N166, N50);
and AND4 (N170, N163, N119, N86, N83);
or OR3 (N171, N153, N116, N165);
buf BUF1 (N172, N56);
and AND3 (N173, N167, N54, N32);
buf BUF1 (N174, N168);
xor XOR2 (N175, N169, N67);
or OR2 (N176, N171, N86);
nor NOR2 (N177, N173, N163);
or OR4 (N178, N176, N177, N15, N126);
nor NOR3 (N179, N137, N105, N119);
and AND2 (N180, N130, N154);
xor XOR2 (N181, N174, N110);
xor XOR2 (N182, N145, N139);
or OR2 (N183, N172, N114);
and AND4 (N184, N162, N149, N182, N158);
xor XOR2 (N185, N33, N131);
or OR2 (N186, N184, N90);
nor NOR4 (N187, N181, N71, N60, N138);
buf BUF1 (N188, N179);
buf BUF1 (N189, N170);
nor NOR2 (N190, N185, N87);
and AND4 (N191, N187, N8, N46, N30);
or OR3 (N192, N183, N74, N110);
or OR3 (N193, N188, N145, N45);
nor NOR3 (N194, N175, N89, N15);
buf BUF1 (N195, N193);
buf BUF1 (N196, N186);
nand NAND4 (N197, N190, N29, N78, N91);
and AND2 (N198, N143, N147);
nand NAND4 (N199, N197, N9, N130, N132);
not NOT1 (N200, N194);
or OR4 (N201, N192, N92, N22, N31);
not NOT1 (N202, N201);
buf BUF1 (N203, N202);
nor NOR3 (N204, N199, N169, N91);
or OR3 (N205, N180, N7, N21);
and AND2 (N206, N191, N109);
and AND4 (N207, N200, N184, N154, N121);
buf BUF1 (N208, N207);
nand NAND3 (N209, N208, N65, N102);
nor NOR4 (N210, N195, N71, N76, N198);
or OR2 (N211, N87, N33);
xor XOR2 (N212, N210, N81);
buf BUF1 (N213, N206);
and AND4 (N214, N189, N6, N97, N92);
or OR4 (N215, N205, N3, N19, N30);
not NOT1 (N216, N212);
or OR2 (N217, N214, N8);
nand NAND4 (N218, N216, N64, N58, N113);
nor NOR3 (N219, N178, N215, N6);
or OR3 (N220, N199, N71, N174);
nor NOR3 (N221, N213, N188, N181);
and AND3 (N222, N221, N88, N199);
xor XOR2 (N223, N196, N104);
nor NOR3 (N224, N204, N16, N174);
or OR4 (N225, N223, N207, N83, N69);
xor XOR2 (N226, N218, N3);
buf BUF1 (N227, N211);
buf BUF1 (N228, N227);
and AND2 (N229, N219, N87);
buf BUF1 (N230, N220);
buf BUF1 (N231, N224);
buf BUF1 (N232, N203);
xor XOR2 (N233, N222, N200);
not NOT1 (N234, N228);
or OR2 (N235, N230, N212);
xor XOR2 (N236, N231, N102);
buf BUF1 (N237, N232);
nor NOR2 (N238, N225, N120);
nand NAND2 (N239, N233, N128);
nand NAND4 (N240, N234, N2, N233, N86);
xor XOR2 (N241, N239, N89);
nand NAND2 (N242, N238, N119);
buf BUF1 (N243, N229);
or OR2 (N244, N236, N212);
not NOT1 (N245, N243);
buf BUF1 (N246, N217);
nand NAND4 (N247, N246, N114, N149, N166);
xor XOR2 (N248, N247, N48);
buf BUF1 (N249, N209);
or OR4 (N250, N237, N108, N122, N160);
nand NAND4 (N251, N226, N235, N36, N218);
and AND2 (N252, N236, N165);
xor XOR2 (N253, N252, N178);
xor XOR2 (N254, N240, N54);
not NOT1 (N255, N241);
and AND2 (N256, N253, N50);
xor XOR2 (N257, N250, N98);
nor NOR3 (N258, N245, N122, N109);
not NOT1 (N259, N255);
nor NOR2 (N260, N256, N117);
nor NOR4 (N261, N251, N258, N243, N105);
xor XOR2 (N262, N125, N154);
or OR2 (N263, N259, N135);
and AND3 (N264, N262, N194, N146);
or OR2 (N265, N260, N103);
nand NAND4 (N266, N244, N71, N76, N227);
nand NAND2 (N267, N249, N57);
xor XOR2 (N268, N266, N152);
xor XOR2 (N269, N268, N257);
xor XOR2 (N270, N192, N159);
xor XOR2 (N271, N269, N132);
buf BUF1 (N272, N261);
not NOT1 (N273, N263);
not NOT1 (N274, N265);
not NOT1 (N275, N272);
buf BUF1 (N276, N254);
xor XOR2 (N277, N248, N91);
or OR4 (N278, N264, N18, N93, N227);
buf BUF1 (N279, N273);
not NOT1 (N280, N267);
nand NAND4 (N281, N279, N80, N151, N125);
or OR4 (N282, N277, N270, N226, N185);
or OR2 (N283, N230, N155);
xor XOR2 (N284, N275, N68);
or OR3 (N285, N278, N240, N108);
or OR2 (N286, N281, N140);
nor NOR4 (N287, N284, N270, N166, N106);
and AND4 (N288, N274, N67, N72, N247);
or OR2 (N289, N271, N17);
nor NOR2 (N290, N289, N48);
not NOT1 (N291, N282);
not NOT1 (N292, N288);
or OR4 (N293, N292, N19, N178, N192);
nand NAND3 (N294, N283, N33, N283);
not NOT1 (N295, N294);
nor NOR4 (N296, N295, N46, N158, N74);
nor NOR2 (N297, N290, N138);
buf BUF1 (N298, N287);
not NOT1 (N299, N276);
and AND4 (N300, N293, N221, N98, N236);
and AND3 (N301, N286, N178, N79);
not NOT1 (N302, N301);
nor NOR3 (N303, N242, N249, N285);
or OR2 (N304, N124, N297);
xor XOR2 (N305, N209, N171);
and AND2 (N306, N296, N305);
xor XOR2 (N307, N104, N214);
or OR3 (N308, N300, N1, N245);
not NOT1 (N309, N308);
nand NAND4 (N310, N306, N251, N207, N157);
not NOT1 (N311, N298);
nor NOR3 (N312, N299, N107, N257);
nor NOR2 (N313, N309, N259);
xor XOR2 (N314, N302, N218);
buf BUF1 (N315, N312);
xor XOR2 (N316, N310, N9);
xor XOR2 (N317, N291, N8);
xor XOR2 (N318, N316, N155);
and AND3 (N319, N313, N196, N187);
or OR3 (N320, N317, N245, N128);
xor XOR2 (N321, N307, N84);
nor NOR3 (N322, N319, N174, N65);
nor NOR4 (N323, N311, N176, N9, N175);
and AND4 (N324, N314, N1, N146, N188);
not NOT1 (N325, N324);
buf BUF1 (N326, N303);
and AND4 (N327, N315, N166, N235, N245);
xor XOR2 (N328, N326, N293);
and AND3 (N329, N322, N87, N129);
nand NAND2 (N330, N329, N191);
and AND3 (N331, N325, N184, N290);
xor XOR2 (N332, N321, N128);
nor NOR4 (N333, N320, N214, N114, N277);
nand NAND3 (N334, N323, N269, N187);
xor XOR2 (N335, N318, N131);
nor NOR4 (N336, N304, N166, N266, N165);
nand NAND3 (N337, N335, N160, N71);
buf BUF1 (N338, N331);
nor NOR2 (N339, N337, N158);
nand NAND2 (N340, N328, N31);
nand NAND2 (N341, N333, N76);
not NOT1 (N342, N330);
or OR3 (N343, N334, N218, N321);
nand NAND3 (N344, N332, N131, N331);
not NOT1 (N345, N336);
or OR4 (N346, N342, N235, N228, N89);
not NOT1 (N347, N339);
nor NOR4 (N348, N280, N322, N318, N21);
and AND3 (N349, N340, N66, N320);
buf BUF1 (N350, N344);
nor NOR2 (N351, N341, N175);
nand NAND3 (N352, N348, N287, N261);
xor XOR2 (N353, N346, N75);
buf BUF1 (N354, N352);
nor NOR3 (N355, N351, N69, N204);
or OR3 (N356, N347, N335, N91);
xor XOR2 (N357, N338, N343);
or OR3 (N358, N37, N328, N126);
xor XOR2 (N359, N350, N222);
xor XOR2 (N360, N354, N256);
nor NOR4 (N361, N358, N178, N149, N43);
nor NOR4 (N362, N356, N32, N290, N110);
buf BUF1 (N363, N355);
and AND2 (N364, N357, N280);
xor XOR2 (N365, N359, N7);
nor NOR3 (N366, N349, N189, N353);
and AND2 (N367, N39, N224);
nand NAND4 (N368, N363, N168, N232, N270);
and AND2 (N369, N366, N148);
nand NAND3 (N370, N365, N161, N134);
xor XOR2 (N371, N370, N87);
nand NAND2 (N372, N371, N131);
and AND2 (N373, N364, N303);
nor NOR3 (N374, N361, N138, N338);
and AND3 (N375, N360, N315, N278);
xor XOR2 (N376, N375, N196);
and AND3 (N377, N327, N274, N77);
and AND3 (N378, N373, N114, N321);
and AND2 (N379, N377, N192);
buf BUF1 (N380, N379);
or OR4 (N381, N345, N64, N362, N70);
not NOT1 (N382, N325);
or OR2 (N383, N372, N147);
buf BUF1 (N384, N367);
nand NAND4 (N385, N380, N294, N2, N82);
and AND2 (N386, N376, N10);
not NOT1 (N387, N384);
not NOT1 (N388, N385);
or OR2 (N389, N369, N148);
not NOT1 (N390, N383);
nand NAND3 (N391, N390, N319, N124);
xor XOR2 (N392, N387, N220);
and AND2 (N393, N368, N243);
nor NOR4 (N394, N386, N30, N374, N205);
not NOT1 (N395, N304);
nor NOR4 (N396, N391, N79, N53, N113);
buf BUF1 (N397, N389);
buf BUF1 (N398, N394);
or OR3 (N399, N393, N322, N26);
and AND4 (N400, N395, N212, N117, N38);
not NOT1 (N401, N382);
nor NOR3 (N402, N378, N47, N146);
buf BUF1 (N403, N398);
or OR3 (N404, N381, N38, N355);
not NOT1 (N405, N401);
nor NOR2 (N406, N403, N181);
xor XOR2 (N407, N396, N312);
not NOT1 (N408, N392);
buf BUF1 (N409, N400);
nor NOR4 (N410, N406, N147, N142, N174);
or OR3 (N411, N397, N183, N156);
nor NOR2 (N412, N410, N60);
not NOT1 (N413, N412);
and AND2 (N414, N409, N360);
xor XOR2 (N415, N413, N174);
nor NOR2 (N416, N402, N244);
or OR3 (N417, N408, N390, N310);
buf BUF1 (N418, N388);
not NOT1 (N419, N399);
and AND2 (N420, N415, N211);
xor XOR2 (N421, N418, N225);
and AND4 (N422, N404, N23, N123, N167);
nor NOR4 (N423, N414, N157, N285, N324);
and AND3 (N424, N405, N229, N265);
not NOT1 (N425, N416);
buf BUF1 (N426, N424);
xor XOR2 (N427, N419, N183);
or OR4 (N428, N426, N40, N5, N5);
not NOT1 (N429, N411);
and AND4 (N430, N422, N145, N147, N118);
and AND4 (N431, N407, N48, N278, N4);
and AND2 (N432, N420, N302);
not NOT1 (N433, N425);
nor NOR2 (N434, N429, N372);
and AND2 (N435, N430, N146);
xor XOR2 (N436, N434, N399);
buf BUF1 (N437, N427);
xor XOR2 (N438, N432, N30);
or OR3 (N439, N428, N24, N36);
nand NAND3 (N440, N435, N179, N343);
nand NAND4 (N441, N436, N132, N41, N284);
nand NAND4 (N442, N417, N120, N305, N153);
or OR2 (N443, N442, N14);
or OR2 (N444, N437, N170);
buf BUF1 (N445, N433);
nand NAND2 (N446, N445, N206);
nor NOR2 (N447, N421, N36);
and AND2 (N448, N444, N162);
buf BUF1 (N449, N438);
nand NAND2 (N450, N431, N126);
and AND4 (N451, N447, N313, N86, N3);
not NOT1 (N452, N450);
buf BUF1 (N453, N446);
and AND4 (N454, N451, N269, N147, N176);
xor XOR2 (N455, N449, N363);
or OR3 (N456, N440, N255, N391);
nand NAND2 (N457, N454, N354);
or OR2 (N458, N452, N220);
and AND4 (N459, N423, N434, N209, N399);
buf BUF1 (N460, N443);
nor NOR2 (N461, N439, N369);
and AND3 (N462, N456, N53, N205);
nand NAND2 (N463, N458, N272);
xor XOR2 (N464, N455, N168);
xor XOR2 (N465, N460, N381);
nor NOR4 (N466, N448, N228, N334, N83);
xor XOR2 (N467, N461, N89);
nand NAND4 (N468, N463, N315, N4, N55);
and AND2 (N469, N466, N26);
xor XOR2 (N470, N441, N7);
and AND4 (N471, N462, N434, N8, N206);
not NOT1 (N472, N464);
buf BUF1 (N473, N470);
nor NOR2 (N474, N469, N404);
xor XOR2 (N475, N467, N72);
nand NAND2 (N476, N473, N445);
xor XOR2 (N477, N476, N416);
nand NAND3 (N478, N472, N231, N211);
buf BUF1 (N479, N471);
nand NAND2 (N480, N475, N254);
buf BUF1 (N481, N453);
xor XOR2 (N482, N457, N263);
nand NAND2 (N483, N482, N57);
nand NAND3 (N484, N481, N137, N197);
xor XOR2 (N485, N480, N241);
nand NAND3 (N486, N474, N478, N243);
or OR4 (N487, N396, N265, N144, N406);
or OR3 (N488, N483, N452, N264);
xor XOR2 (N489, N465, N433);
nand NAND3 (N490, N488, N261, N194);
not NOT1 (N491, N485);
and AND2 (N492, N479, N453);
or OR4 (N493, N489, N120, N172, N70);
xor XOR2 (N494, N492, N451);
buf BUF1 (N495, N459);
buf BUF1 (N496, N477);
not NOT1 (N497, N494);
buf BUF1 (N498, N486);
nand NAND2 (N499, N468, N458);
buf BUF1 (N500, N491);
and AND3 (N501, N490, N33, N81);
and AND4 (N502, N487, N460, N191, N441);
and AND2 (N503, N497, N353);
nor NOR2 (N504, N501, N488);
buf BUF1 (N505, N500);
nand NAND3 (N506, N495, N292, N44);
or OR3 (N507, N505, N261, N474);
xor XOR2 (N508, N493, N477);
nor NOR3 (N509, N507, N243, N188);
xor XOR2 (N510, N504, N253);
and AND2 (N511, N503, N263);
not NOT1 (N512, N510);
nand NAND4 (N513, N509, N103, N316, N76);
xor XOR2 (N514, N498, N122);
xor XOR2 (N515, N496, N325);
buf BUF1 (N516, N499);
or OR2 (N517, N511, N2);
nand NAND4 (N518, N516, N477, N57, N147);
nand NAND4 (N519, N502, N248, N460, N504);
nand NAND3 (N520, N518, N166, N114);
xor XOR2 (N521, N513, N114);
nor NOR3 (N522, N521, N228, N441);
and AND3 (N523, N520, N146, N179);
nand NAND3 (N524, N515, N522, N328);
xor XOR2 (N525, N140, N72);
buf BUF1 (N526, N506);
nor NOR2 (N527, N525, N204);
not NOT1 (N528, N512);
buf BUF1 (N529, N527);
buf BUF1 (N530, N519);
xor XOR2 (N531, N517, N430);
not NOT1 (N532, N523);
nor NOR2 (N533, N526, N442);
nor NOR4 (N534, N531, N77, N495, N378);
or OR3 (N535, N524, N394, N239);
nand NAND2 (N536, N533, N440);
nand NAND4 (N537, N484, N106, N30, N389);
buf BUF1 (N538, N529);
and AND2 (N539, N535, N341);
xor XOR2 (N540, N538, N160);
or OR3 (N541, N532, N241, N268);
or OR4 (N542, N534, N513, N72, N250);
nand NAND2 (N543, N540, N130);
nor NOR3 (N544, N528, N357, N112);
nor NOR3 (N545, N544, N56, N300);
xor XOR2 (N546, N543, N175);
buf BUF1 (N547, N545);
nor NOR2 (N548, N546, N100);
nand NAND4 (N549, N548, N61, N394, N447);
or OR4 (N550, N539, N220, N366, N437);
xor XOR2 (N551, N536, N409);
buf BUF1 (N552, N514);
nand NAND2 (N553, N547, N12);
or OR3 (N554, N553, N265, N389);
or OR4 (N555, N549, N127, N237, N70);
buf BUF1 (N556, N530);
nor NOR4 (N557, N542, N217, N316, N83);
not NOT1 (N558, N556);
or OR2 (N559, N555, N97);
buf BUF1 (N560, N558);
and AND2 (N561, N552, N153);
buf BUF1 (N562, N554);
or OR3 (N563, N561, N307, N237);
buf BUF1 (N564, N551);
buf BUF1 (N565, N541);
xor XOR2 (N566, N559, N57);
not NOT1 (N567, N566);
or OR4 (N568, N562, N33, N37, N98);
not NOT1 (N569, N557);
not NOT1 (N570, N564);
nor NOR3 (N571, N569, N373, N312);
buf BUF1 (N572, N563);
and AND3 (N573, N567, N531, N301);
nand NAND2 (N574, N508, N222);
buf BUF1 (N575, N572);
and AND2 (N576, N560, N354);
not NOT1 (N577, N550);
xor XOR2 (N578, N574, N208);
not NOT1 (N579, N577);
nand NAND3 (N580, N568, N562, N97);
and AND4 (N581, N571, N479, N56, N145);
or OR3 (N582, N575, N294, N371);
and AND3 (N583, N576, N95, N495);
xor XOR2 (N584, N582, N63);
xor XOR2 (N585, N583, N408);
buf BUF1 (N586, N584);
nor NOR2 (N587, N585, N415);
nor NOR3 (N588, N570, N87, N358);
and AND2 (N589, N579, N199);
xor XOR2 (N590, N589, N139);
nand NAND3 (N591, N565, N547, N448);
and AND4 (N592, N590, N121, N169, N509);
buf BUF1 (N593, N587);
nand NAND4 (N594, N588, N239, N555, N476);
nand NAND3 (N595, N580, N554, N310);
not NOT1 (N596, N591);
nor NOR3 (N597, N593, N158, N137);
nand NAND3 (N598, N573, N98, N320);
nand NAND3 (N599, N595, N172, N121);
xor XOR2 (N600, N599, N335);
buf BUF1 (N601, N596);
or OR3 (N602, N594, N203, N267);
not NOT1 (N603, N586);
nand NAND2 (N604, N597, N241);
nand NAND3 (N605, N600, N63, N23);
nor NOR3 (N606, N604, N60, N79);
nand NAND3 (N607, N581, N450, N446);
xor XOR2 (N608, N578, N137);
not NOT1 (N609, N606);
and AND2 (N610, N609, N300);
nor NOR4 (N611, N598, N108, N357, N320);
nand NAND2 (N612, N607, N136);
and AND3 (N613, N612, N593, N21);
xor XOR2 (N614, N537, N368);
nor NOR3 (N615, N614, N40, N220);
not NOT1 (N616, N608);
nor NOR3 (N617, N615, N82, N260);
xor XOR2 (N618, N613, N75);
nand NAND2 (N619, N602, N422);
or OR2 (N620, N616, N379);
and AND4 (N621, N617, N401, N523, N43);
or OR2 (N622, N621, N489);
nand NAND4 (N623, N605, N276, N444, N496);
nor NOR4 (N624, N622, N154, N561, N132);
nor NOR4 (N625, N618, N454, N321, N374);
not NOT1 (N626, N623);
buf BUF1 (N627, N619);
not NOT1 (N628, N627);
xor XOR2 (N629, N610, N570);
nor NOR2 (N630, N629, N104);
nand NAND4 (N631, N601, N67, N79, N62);
or OR3 (N632, N592, N187, N397);
buf BUF1 (N633, N628);
not NOT1 (N634, N630);
not NOT1 (N635, N620);
buf BUF1 (N636, N633);
not NOT1 (N637, N634);
and AND2 (N638, N632, N569);
nand NAND2 (N639, N625, N268);
and AND3 (N640, N631, N555, N380);
or OR2 (N641, N639, N282);
nand NAND2 (N642, N636, N68);
not NOT1 (N643, N637);
xor XOR2 (N644, N603, N175);
nand NAND3 (N645, N644, N127, N12);
xor XOR2 (N646, N642, N206);
xor XOR2 (N647, N641, N454);
buf BUF1 (N648, N640);
nor NOR2 (N649, N643, N215);
not NOT1 (N650, N626);
and AND2 (N651, N647, N555);
not NOT1 (N652, N611);
nor NOR4 (N653, N652, N625, N500, N205);
nor NOR4 (N654, N645, N614, N324, N289);
not NOT1 (N655, N635);
and AND4 (N656, N624, N7, N113, N425);
xor XOR2 (N657, N653, N452);
xor XOR2 (N658, N654, N420);
or OR3 (N659, N650, N654, N645);
and AND2 (N660, N655, N267);
nor NOR3 (N661, N657, N476, N569);
xor XOR2 (N662, N646, N409);
nor NOR2 (N663, N660, N478);
not NOT1 (N664, N658);
xor XOR2 (N665, N661, N539);
nand NAND4 (N666, N649, N589, N28, N437);
buf BUF1 (N667, N664);
xor XOR2 (N668, N651, N379);
and AND3 (N669, N668, N589, N441);
or OR2 (N670, N656, N238);
xor XOR2 (N671, N670, N595);
nand NAND2 (N672, N665, N666);
nor NOR3 (N673, N531, N308, N6);
buf BUF1 (N674, N667);
nand NAND4 (N675, N674, N459, N460, N214);
buf BUF1 (N676, N671);
nand NAND4 (N677, N675, N77, N635, N129);
or OR2 (N678, N672, N153);
nand NAND4 (N679, N663, N594, N58, N505);
and AND4 (N680, N673, N274, N81, N337);
nor NOR3 (N681, N680, N391, N574);
nand NAND3 (N682, N679, N61, N60);
buf BUF1 (N683, N638);
buf BUF1 (N684, N677);
nor NOR4 (N685, N648, N77, N13, N27);
and AND2 (N686, N681, N181);
nand NAND4 (N687, N682, N461, N75, N342);
not NOT1 (N688, N683);
xor XOR2 (N689, N669, N466);
buf BUF1 (N690, N689);
and AND3 (N691, N687, N649, N203);
and AND4 (N692, N690, N190, N299, N99);
not NOT1 (N693, N676);
xor XOR2 (N694, N688, N574);
not NOT1 (N695, N662);
buf BUF1 (N696, N678);
buf BUF1 (N697, N685);
xor XOR2 (N698, N686, N482);
xor XOR2 (N699, N691, N130);
nand NAND2 (N700, N684, N40);
nor NOR2 (N701, N692, N119);
buf BUF1 (N702, N696);
or OR2 (N703, N702, N354);
not NOT1 (N704, N695);
xor XOR2 (N705, N699, N95);
xor XOR2 (N706, N694, N132);
xor XOR2 (N707, N700, N171);
or OR4 (N708, N707, N687, N669, N322);
xor XOR2 (N709, N659, N222);
nor NOR3 (N710, N704, N624, N484);
nand NAND4 (N711, N706, N629, N705, N362);
not NOT1 (N712, N364);
nand NAND2 (N713, N697, N372);
and AND3 (N714, N708, N146, N261);
buf BUF1 (N715, N713);
nor NOR3 (N716, N698, N3, N143);
xor XOR2 (N717, N710, N289);
xor XOR2 (N718, N715, N183);
xor XOR2 (N719, N717, N654);
xor XOR2 (N720, N693, N103);
xor XOR2 (N721, N701, N417);
nand NAND3 (N722, N718, N718, N123);
buf BUF1 (N723, N719);
and AND3 (N724, N712, N295, N687);
and AND4 (N725, N709, N92, N158, N165);
xor XOR2 (N726, N711, N478);
or OR4 (N727, N725, N94, N519, N102);
nor NOR2 (N728, N720, N721);
nor NOR3 (N729, N89, N441, N456);
not NOT1 (N730, N729);
not NOT1 (N731, N726);
buf BUF1 (N732, N722);
not NOT1 (N733, N731);
nor NOR3 (N734, N716, N618, N428);
xor XOR2 (N735, N730, N476);
nor NOR3 (N736, N714, N25, N512);
nor NOR2 (N737, N733, N266);
not NOT1 (N738, N736);
or OR4 (N739, N728, N394, N270, N62);
xor XOR2 (N740, N723, N660);
and AND4 (N741, N732, N359, N423, N299);
or OR2 (N742, N727, N140);
or OR4 (N743, N740, N177, N582, N607);
xor XOR2 (N744, N724, N308);
and AND4 (N745, N703, N712, N349, N69);
not NOT1 (N746, N744);
or OR2 (N747, N741, N46);
nor NOR4 (N748, N739, N499, N400, N554);
xor XOR2 (N749, N737, N615);
not NOT1 (N750, N748);
or OR2 (N751, N746, N711);
buf BUF1 (N752, N738);
nand NAND3 (N753, N747, N69, N116);
nor NOR2 (N754, N742, N462);
not NOT1 (N755, N745);
buf BUF1 (N756, N735);
not NOT1 (N757, N756);
or OR4 (N758, N751, N190, N581, N235);
buf BUF1 (N759, N750);
nand NAND2 (N760, N755, N101);
buf BUF1 (N761, N760);
or OR3 (N762, N754, N31, N423);
not NOT1 (N763, N749);
or OR3 (N764, N752, N445, N72);
and AND2 (N765, N743, N238);
nand NAND3 (N766, N759, N133, N394);
or OR2 (N767, N762, N97);
or OR2 (N768, N766, N506);
buf BUF1 (N769, N753);
nand NAND2 (N770, N765, N134);
or OR3 (N771, N768, N265, N239);
nor NOR3 (N772, N769, N696, N485);
or OR4 (N773, N767, N230, N377, N743);
and AND3 (N774, N763, N340, N30);
or OR2 (N775, N734, N23);
or OR2 (N776, N773, N753);
not NOT1 (N777, N758);
not NOT1 (N778, N764);
not NOT1 (N779, N772);
not NOT1 (N780, N757);
nand NAND4 (N781, N770, N190, N211, N373);
and AND2 (N782, N776, N477);
xor XOR2 (N783, N779, N297);
nor NOR2 (N784, N771, N768);
or OR4 (N785, N778, N90, N205, N752);
buf BUF1 (N786, N785);
xor XOR2 (N787, N761, N333);
not NOT1 (N788, N787);
or OR3 (N789, N784, N772, N599);
buf BUF1 (N790, N774);
xor XOR2 (N791, N781, N615);
or OR2 (N792, N777, N444);
nor NOR2 (N793, N780, N474);
xor XOR2 (N794, N790, N511);
buf BUF1 (N795, N782);
or OR3 (N796, N789, N421, N69);
not NOT1 (N797, N786);
or OR3 (N798, N797, N778, N25);
or OR3 (N799, N791, N122, N363);
nand NAND2 (N800, N799, N592);
or OR3 (N801, N798, N735, N583);
buf BUF1 (N802, N794);
not NOT1 (N803, N792);
nor NOR2 (N804, N793, N115);
or OR3 (N805, N796, N315, N27);
buf BUF1 (N806, N801);
or OR3 (N807, N795, N471, N791);
xor XOR2 (N808, N788, N132);
not NOT1 (N809, N804);
xor XOR2 (N810, N802, N624);
not NOT1 (N811, N775);
or OR4 (N812, N810, N16, N185, N568);
or OR2 (N813, N805, N767);
or OR4 (N814, N800, N4, N715, N324);
nand NAND2 (N815, N809, N410);
xor XOR2 (N816, N807, N30);
not NOT1 (N817, N806);
not NOT1 (N818, N814);
nor NOR2 (N819, N816, N729);
not NOT1 (N820, N811);
xor XOR2 (N821, N820, N403);
nand NAND3 (N822, N783, N297, N700);
and AND3 (N823, N818, N395, N816);
nand NAND2 (N824, N813, N664);
xor XOR2 (N825, N821, N398);
xor XOR2 (N826, N825, N699);
nor NOR3 (N827, N803, N498, N369);
and AND4 (N828, N827, N358, N777, N673);
nor NOR3 (N829, N822, N668, N177);
nand NAND4 (N830, N828, N314, N669, N758);
buf BUF1 (N831, N808);
nand NAND4 (N832, N830, N167, N532, N742);
or OR4 (N833, N832, N809, N204, N5);
or OR2 (N834, N833, N137);
xor XOR2 (N835, N819, N29);
nand NAND2 (N836, N824, N243);
xor XOR2 (N837, N817, N374);
buf BUF1 (N838, N826);
xor XOR2 (N839, N834, N683);
buf BUF1 (N840, N812);
not NOT1 (N841, N839);
nor NOR2 (N842, N840, N704);
and AND4 (N843, N831, N730, N358, N221);
nor NOR3 (N844, N838, N95, N535);
xor XOR2 (N845, N823, N523);
nor NOR2 (N846, N844, N513);
xor XOR2 (N847, N841, N133);
buf BUF1 (N848, N836);
xor XOR2 (N849, N842, N635);
not NOT1 (N850, N815);
nand NAND3 (N851, N845, N106, N284);
xor XOR2 (N852, N850, N847);
and AND2 (N853, N296, N830);
or OR3 (N854, N843, N611, N290);
xor XOR2 (N855, N837, N749);
nor NOR2 (N856, N853, N662);
xor XOR2 (N857, N849, N223);
buf BUF1 (N858, N829);
xor XOR2 (N859, N857, N320);
xor XOR2 (N860, N856, N801);
or OR4 (N861, N848, N215, N364, N97);
nor NOR2 (N862, N860, N622);
not NOT1 (N863, N846);
not NOT1 (N864, N861);
nand NAND3 (N865, N858, N672, N640);
xor XOR2 (N866, N851, N601);
nor NOR4 (N867, N864, N843, N564, N808);
xor XOR2 (N868, N866, N715);
not NOT1 (N869, N862);
and AND2 (N870, N852, N795);
buf BUF1 (N871, N869);
buf BUF1 (N872, N867);
xor XOR2 (N873, N872, N769);
nor NOR4 (N874, N863, N348, N357, N527);
nand NAND3 (N875, N871, N430, N777);
buf BUF1 (N876, N868);
nand NAND4 (N877, N875, N357, N209, N562);
and AND3 (N878, N870, N209, N494);
nor NOR2 (N879, N877, N621);
buf BUF1 (N880, N835);
and AND3 (N881, N859, N423, N777);
nand NAND4 (N882, N879, N474, N608, N438);
or OR3 (N883, N874, N789, N112);
or OR2 (N884, N873, N565);
or OR3 (N885, N878, N857, N538);
nand NAND3 (N886, N882, N684, N607);
buf BUF1 (N887, N881);
or OR3 (N888, N876, N557, N58);
not NOT1 (N889, N865);
nand NAND4 (N890, N880, N395, N205, N672);
not NOT1 (N891, N885);
not NOT1 (N892, N883);
or OR2 (N893, N888, N243);
and AND2 (N894, N893, N550);
not NOT1 (N895, N894);
buf BUF1 (N896, N854);
xor XOR2 (N897, N884, N115);
buf BUF1 (N898, N889);
not NOT1 (N899, N887);
nor NOR2 (N900, N891, N264);
nor NOR4 (N901, N898, N144, N564, N667);
nor NOR4 (N902, N896, N181, N748, N615);
or OR2 (N903, N900, N495);
buf BUF1 (N904, N902);
buf BUF1 (N905, N855);
not NOT1 (N906, N890);
or OR3 (N907, N897, N54, N749);
xor XOR2 (N908, N907, N22);
and AND2 (N909, N892, N393);
or OR2 (N910, N906, N890);
nand NAND4 (N911, N910, N488, N871, N226);
not NOT1 (N912, N908);
buf BUF1 (N913, N911);
nor NOR4 (N914, N905, N213, N718, N617);
xor XOR2 (N915, N903, N534);
nand NAND3 (N916, N886, N416, N635);
or OR2 (N917, N901, N743);
nand NAND3 (N918, N914, N818, N508);
buf BUF1 (N919, N912);
buf BUF1 (N920, N895);
nor NOR3 (N921, N919, N524, N586);
xor XOR2 (N922, N899, N185);
not NOT1 (N923, N904);
not NOT1 (N924, N922);
and AND2 (N925, N915, N608);
nor NOR3 (N926, N917, N185, N324);
and AND2 (N927, N926, N888);
not NOT1 (N928, N924);
nand NAND4 (N929, N927, N173, N505, N78);
not NOT1 (N930, N918);
and AND2 (N931, N913, N345);
not NOT1 (N932, N931);
nor NOR3 (N933, N929, N547, N450);
xor XOR2 (N934, N920, N728);
nand NAND3 (N935, N933, N886, N555);
not NOT1 (N936, N932);
and AND2 (N937, N925, N50);
nor NOR4 (N938, N934, N852, N767, N684);
buf BUF1 (N939, N909);
or OR2 (N940, N930, N726);
nor NOR2 (N941, N940, N835);
nand NAND2 (N942, N921, N128);
or OR4 (N943, N939, N443, N371, N583);
buf BUF1 (N944, N923);
nand NAND4 (N945, N935, N933, N180, N259);
xor XOR2 (N946, N928, N943);
nand NAND2 (N947, N63, N311);
xor XOR2 (N948, N947, N49);
or OR4 (N949, N944, N851, N901, N424);
buf BUF1 (N950, N942);
xor XOR2 (N951, N916, N62);
not NOT1 (N952, N936);
or OR3 (N953, N952, N906, N128);
nand NAND4 (N954, N946, N948, N597, N364);
nor NOR2 (N955, N812, N476);
not NOT1 (N956, N950);
xor XOR2 (N957, N945, N356);
nor NOR4 (N958, N957, N900, N565, N625);
xor XOR2 (N959, N949, N927);
or OR3 (N960, N951, N590, N395);
xor XOR2 (N961, N960, N519);
nand NAND3 (N962, N937, N690, N906);
xor XOR2 (N963, N955, N37);
nand NAND4 (N964, N953, N907, N669, N762);
and AND3 (N965, N962, N471, N745);
xor XOR2 (N966, N938, N960);
xor XOR2 (N967, N941, N229);
xor XOR2 (N968, N963, N49);
not NOT1 (N969, N968);
nand NAND3 (N970, N958, N325, N526);
nand NAND4 (N971, N964, N796, N360, N292);
xor XOR2 (N972, N965, N260);
nor NOR2 (N973, N956, N933);
nor NOR3 (N974, N966, N67, N229);
not NOT1 (N975, N974);
and AND3 (N976, N973, N718, N913);
not NOT1 (N977, N967);
nand NAND3 (N978, N954, N727, N594);
xor XOR2 (N979, N977, N892);
not NOT1 (N980, N979);
buf BUF1 (N981, N980);
or OR2 (N982, N959, N470);
and AND3 (N983, N961, N175, N446);
nand NAND2 (N984, N969, N979);
xor XOR2 (N985, N981, N480);
buf BUF1 (N986, N984);
xor XOR2 (N987, N975, N700);
not NOT1 (N988, N983);
and AND2 (N989, N970, N737);
nand NAND3 (N990, N976, N212, N920);
or OR2 (N991, N971, N197);
not NOT1 (N992, N987);
nand NAND2 (N993, N982, N695);
and AND4 (N994, N989, N585, N286, N358);
nor NOR4 (N995, N988, N334, N471, N550);
not NOT1 (N996, N995);
and AND3 (N997, N992, N401, N121);
buf BUF1 (N998, N986);
not NOT1 (N999, N978);
buf BUF1 (N1000, N990);
and AND3 (N1001, N985, N747, N39);
buf BUF1 (N1002, N1001);
nor NOR2 (N1003, N1002, N977);
buf BUF1 (N1004, N997);
buf BUF1 (N1005, N972);
nand NAND2 (N1006, N996, N132);
buf BUF1 (N1007, N1003);
nand NAND3 (N1008, N1006, N1002, N237);
nor NOR4 (N1009, N998, N332, N17, N859);
xor XOR2 (N1010, N1007, N504);
nor NOR2 (N1011, N994, N960);
and AND4 (N1012, N991, N964, N733, N235);
and AND2 (N1013, N1000, N903);
not NOT1 (N1014, N1004);
buf BUF1 (N1015, N1011);
and AND2 (N1016, N1015, N390);
nand NAND2 (N1017, N1005, N1015);
and AND3 (N1018, N1014, N354, N880);
nand NAND2 (N1019, N1018, N108);
buf BUF1 (N1020, N999);
nor NOR2 (N1021, N1010, N1006);
or OR3 (N1022, N1020, N225, N88);
nand NAND2 (N1023, N993, N149);
and AND2 (N1024, N1019, N592);
nand NAND2 (N1025, N1012, N215);
xor XOR2 (N1026, N1008, N928);
xor XOR2 (N1027, N1022, N81);
xor XOR2 (N1028, N1026, N532);
nand NAND2 (N1029, N1028, N59);
xor XOR2 (N1030, N1027, N503);
or OR3 (N1031, N1013, N367, N342);
and AND2 (N1032, N1030, N296);
buf BUF1 (N1033, N1023);
not NOT1 (N1034, N1024);
nand NAND4 (N1035, N1009, N94, N740, N1);
and AND2 (N1036, N1034, N957);
xor XOR2 (N1037, N1017, N260);
nand NAND3 (N1038, N1035, N348, N158);
not NOT1 (N1039, N1021);
not NOT1 (N1040, N1032);
and AND3 (N1041, N1036, N704, N953);
nor NOR2 (N1042, N1033, N337);
or OR4 (N1043, N1042, N609, N936, N61);
nand NAND4 (N1044, N1039, N355, N77, N858);
buf BUF1 (N1045, N1025);
nand NAND4 (N1046, N1037, N796, N485, N489);
or OR2 (N1047, N1029, N756);
not NOT1 (N1048, N1046);
xor XOR2 (N1049, N1016, N122);
not NOT1 (N1050, N1049);
or OR3 (N1051, N1038, N16, N634);
nand NAND3 (N1052, N1047, N374, N659);
and AND2 (N1053, N1044, N307);
xor XOR2 (N1054, N1043, N256);
nand NAND2 (N1055, N1051, N130);
nor NOR3 (N1056, N1055, N986, N870);
xor XOR2 (N1057, N1040, N1048);
buf BUF1 (N1058, N531);
xor XOR2 (N1059, N1052, N604);
xor XOR2 (N1060, N1050, N642);
xor XOR2 (N1061, N1045, N1005);
or OR3 (N1062, N1041, N855, N563);
buf BUF1 (N1063, N1056);
not NOT1 (N1064, N1031);
nor NOR4 (N1065, N1057, N1009, N594, N340);
and AND3 (N1066, N1060, N1009, N947);
and AND4 (N1067, N1063, N963, N148, N655);
xor XOR2 (N1068, N1067, N119);
xor XOR2 (N1069, N1062, N921);
and AND4 (N1070, N1068, N899, N1046, N338);
buf BUF1 (N1071, N1061);
nor NOR2 (N1072, N1071, N574);
or OR3 (N1073, N1066, N324, N195);
xor XOR2 (N1074, N1072, N17);
and AND2 (N1075, N1064, N672);
buf BUF1 (N1076, N1053);
and AND3 (N1077, N1074, N534, N591);
nor NOR4 (N1078, N1058, N763, N783, N41);
or OR2 (N1079, N1075, N394);
xor XOR2 (N1080, N1078, N150);
not NOT1 (N1081, N1077);
xor XOR2 (N1082, N1070, N289);
nand NAND2 (N1083, N1082, N410);
nand NAND3 (N1084, N1080, N811, N680);
nor NOR2 (N1085, N1079, N312);
or OR3 (N1086, N1065, N434, N575);
xor XOR2 (N1087, N1069, N159);
nand NAND2 (N1088, N1054, N709);
xor XOR2 (N1089, N1076, N675);
buf BUF1 (N1090, N1083);
or OR4 (N1091, N1087, N526, N278, N114);
xor XOR2 (N1092, N1081, N380);
buf BUF1 (N1093, N1089);
nor NOR2 (N1094, N1084, N563);
nor NOR4 (N1095, N1091, N352, N280, N107);
or OR3 (N1096, N1059, N972, N502);
or OR2 (N1097, N1092, N194);
or OR3 (N1098, N1088, N545, N1082);
not NOT1 (N1099, N1086);
and AND4 (N1100, N1097, N717, N446, N1061);
or OR2 (N1101, N1099, N713);
buf BUF1 (N1102, N1096);
nand NAND3 (N1103, N1094, N132, N459);
xor XOR2 (N1104, N1098, N344);
nand NAND3 (N1105, N1101, N359, N244);
not NOT1 (N1106, N1090);
not NOT1 (N1107, N1100);
nand NAND2 (N1108, N1085, N390);
nand NAND4 (N1109, N1103, N447, N348, N1017);
buf BUF1 (N1110, N1108);
not NOT1 (N1111, N1073);
not NOT1 (N1112, N1102);
not NOT1 (N1113, N1106);
nor NOR2 (N1114, N1112, N136);
xor XOR2 (N1115, N1109, N658);
not NOT1 (N1116, N1114);
or OR4 (N1117, N1093, N612, N1072, N423);
buf BUF1 (N1118, N1110);
nand NAND3 (N1119, N1113, N58, N1018);
buf BUF1 (N1120, N1118);
nor NOR4 (N1121, N1095, N827, N980, N167);
or OR4 (N1122, N1115, N1029, N497, N922);
or OR4 (N1123, N1121, N1020, N391, N749);
and AND4 (N1124, N1123, N253, N309, N335);
or OR4 (N1125, N1122, N1043, N678, N350);
nand NAND4 (N1126, N1124, N1026, N856, N298);
xor XOR2 (N1127, N1111, N924);
and AND3 (N1128, N1116, N76, N313);
nand NAND2 (N1129, N1125, N193);
nor NOR3 (N1130, N1126, N328, N718);
buf BUF1 (N1131, N1129);
nand NAND4 (N1132, N1104, N960, N166, N1013);
xor XOR2 (N1133, N1132, N436);
or OR4 (N1134, N1130, N347, N279, N653);
nor NOR2 (N1135, N1133, N655);
nand NAND2 (N1136, N1105, N860);
not NOT1 (N1137, N1128);
xor XOR2 (N1138, N1120, N865);
xor XOR2 (N1139, N1134, N1102);
and AND2 (N1140, N1117, N366);
buf BUF1 (N1141, N1136);
and AND2 (N1142, N1141, N530);
nor NOR2 (N1143, N1140, N313);
nor NOR2 (N1144, N1137, N924);
or OR3 (N1145, N1131, N786, N262);
nand NAND2 (N1146, N1143, N74);
or OR2 (N1147, N1139, N28);
buf BUF1 (N1148, N1144);
nor NOR2 (N1149, N1135, N455);
nor NOR2 (N1150, N1147, N640);
and AND3 (N1151, N1146, N765, N352);
nand NAND4 (N1152, N1151, N881, N823, N483);
nand NAND4 (N1153, N1152, N1084, N181, N1050);
or OR3 (N1154, N1145, N642, N601);
buf BUF1 (N1155, N1107);
nand NAND4 (N1156, N1155, N866, N86, N12);
and AND2 (N1157, N1150, N558);
not NOT1 (N1158, N1154);
nor NOR2 (N1159, N1119, N835);
and AND4 (N1160, N1148, N995, N977, N285);
not NOT1 (N1161, N1153);
not NOT1 (N1162, N1138);
nor NOR3 (N1163, N1149, N216, N1051);
buf BUF1 (N1164, N1163);
not NOT1 (N1165, N1164);
nand NAND2 (N1166, N1161, N26);
buf BUF1 (N1167, N1158);
nand NAND2 (N1168, N1127, N657);
and AND2 (N1169, N1166, N240);
nand NAND2 (N1170, N1142, N718);
not NOT1 (N1171, N1167);
nand NAND3 (N1172, N1170, N865, N324);
nor NOR2 (N1173, N1169, N1096);
nand NAND2 (N1174, N1165, N62);
or OR3 (N1175, N1156, N951, N993);
buf BUF1 (N1176, N1162);
or OR4 (N1177, N1171, N621, N376, N852);
buf BUF1 (N1178, N1173);
buf BUF1 (N1179, N1177);
buf BUF1 (N1180, N1175);
nand NAND2 (N1181, N1179, N155);
nand NAND4 (N1182, N1168, N57, N137, N912);
buf BUF1 (N1183, N1180);
nand NAND3 (N1184, N1183, N717, N1148);
and AND2 (N1185, N1176, N243);
nand NAND3 (N1186, N1159, N747, N377);
xor XOR2 (N1187, N1172, N658);
nor NOR3 (N1188, N1186, N140, N794);
nor NOR3 (N1189, N1188, N1107, N657);
nor NOR3 (N1190, N1181, N337, N1013);
buf BUF1 (N1191, N1160);
xor XOR2 (N1192, N1157, N384);
buf BUF1 (N1193, N1178);
nor NOR3 (N1194, N1184, N717, N960);
nand NAND3 (N1195, N1185, N444, N1131);
nand NAND2 (N1196, N1193, N279);
or OR3 (N1197, N1195, N1083, N309);
nand NAND3 (N1198, N1191, N50, N801);
nor NOR4 (N1199, N1194, N326, N25, N1139);
buf BUF1 (N1200, N1187);
not NOT1 (N1201, N1190);
and AND2 (N1202, N1196, N303);
nand NAND2 (N1203, N1189, N513);
buf BUF1 (N1204, N1197);
xor XOR2 (N1205, N1182, N373);
nor NOR2 (N1206, N1203, N116);
or OR4 (N1207, N1200, N88, N1093, N737);
buf BUF1 (N1208, N1205);
or OR3 (N1209, N1208, N757, N666);
and AND2 (N1210, N1201, N814);
xor XOR2 (N1211, N1207, N1033);
buf BUF1 (N1212, N1204);
not NOT1 (N1213, N1192);
and AND3 (N1214, N1210, N1095, N614);
and AND3 (N1215, N1209, N1153, N17);
not NOT1 (N1216, N1202);
xor XOR2 (N1217, N1211, N742);
nor NOR3 (N1218, N1174, N816, N496);
xor XOR2 (N1219, N1213, N1055);
buf BUF1 (N1220, N1215);
not NOT1 (N1221, N1217);
nor NOR4 (N1222, N1220, N1146, N976, N1062);
and AND4 (N1223, N1212, N353, N68, N984);
buf BUF1 (N1224, N1221);
buf BUF1 (N1225, N1222);
xor XOR2 (N1226, N1224, N948);
buf BUF1 (N1227, N1223);
buf BUF1 (N1228, N1227);
nor NOR3 (N1229, N1228, N1208, N209);
buf BUF1 (N1230, N1225);
or OR2 (N1231, N1219, N470);
not NOT1 (N1232, N1216);
not NOT1 (N1233, N1199);
buf BUF1 (N1234, N1232);
and AND2 (N1235, N1218, N165);
buf BUF1 (N1236, N1206);
buf BUF1 (N1237, N1229);
or OR3 (N1238, N1230, N182, N251);
and AND3 (N1239, N1233, N1178, N163);
nor NOR4 (N1240, N1226, N180, N1189, N219);
buf BUF1 (N1241, N1240);
not NOT1 (N1242, N1239);
xor XOR2 (N1243, N1234, N978);
nor NOR4 (N1244, N1238, N342, N323, N337);
nor NOR3 (N1245, N1235, N785, N988);
nand NAND2 (N1246, N1214, N459);
not NOT1 (N1247, N1241);
and AND2 (N1248, N1237, N264);
nand NAND2 (N1249, N1244, N339);
xor XOR2 (N1250, N1231, N355);
or OR4 (N1251, N1249, N423, N280, N652);
xor XOR2 (N1252, N1246, N161);
or OR3 (N1253, N1245, N1238, N453);
and AND2 (N1254, N1242, N508);
not NOT1 (N1255, N1252);
not NOT1 (N1256, N1198);
nand NAND3 (N1257, N1243, N985, N876);
not NOT1 (N1258, N1247);
not NOT1 (N1259, N1236);
not NOT1 (N1260, N1255);
or OR2 (N1261, N1258, N618);
xor XOR2 (N1262, N1257, N1155);
or OR4 (N1263, N1253, N1032, N868, N428);
or OR4 (N1264, N1259, N29, N208, N486);
and AND4 (N1265, N1250, N1170, N718, N1057);
nor NOR2 (N1266, N1248, N545);
or OR2 (N1267, N1254, N520);
and AND2 (N1268, N1265, N137);
and AND3 (N1269, N1261, N402, N357);
or OR3 (N1270, N1264, N334, N70);
nand NAND2 (N1271, N1263, N310);
xor XOR2 (N1272, N1271, N360);
nor NOR2 (N1273, N1251, N358);
xor XOR2 (N1274, N1268, N908);
nand NAND3 (N1275, N1260, N1220, N448);
nand NAND3 (N1276, N1275, N1064, N1071);
buf BUF1 (N1277, N1267);
not NOT1 (N1278, N1274);
or OR2 (N1279, N1272, N1172);
and AND2 (N1280, N1278, N168);
nand NAND2 (N1281, N1276, N11);
xor XOR2 (N1282, N1273, N184);
nor NOR3 (N1283, N1282, N1123, N992);
nor NOR4 (N1284, N1266, N626, N1095, N1267);
xor XOR2 (N1285, N1270, N279);
not NOT1 (N1286, N1281);
or OR2 (N1287, N1284, N479);
nor NOR2 (N1288, N1283, N722);
or OR4 (N1289, N1256, N551, N134, N143);
or OR2 (N1290, N1285, N797);
or OR2 (N1291, N1287, N1088);
buf BUF1 (N1292, N1289);
not NOT1 (N1293, N1291);
and AND3 (N1294, N1292, N447, N798);
nand NAND4 (N1295, N1286, N270, N597, N69);
not NOT1 (N1296, N1290);
or OR2 (N1297, N1269, N972);
or OR3 (N1298, N1280, N241, N829);
nor NOR2 (N1299, N1293, N927);
not NOT1 (N1300, N1298);
nor NOR3 (N1301, N1297, N834, N136);
xor XOR2 (N1302, N1300, N123);
buf BUF1 (N1303, N1295);
nand NAND3 (N1304, N1296, N707, N216);
not NOT1 (N1305, N1299);
or OR4 (N1306, N1304, N767, N725, N253);
or OR3 (N1307, N1279, N627, N271);
not NOT1 (N1308, N1307);
or OR2 (N1309, N1306, N847);
nand NAND3 (N1310, N1301, N680, N76);
and AND3 (N1311, N1277, N841, N209);
nand NAND4 (N1312, N1303, N1094, N957, N1185);
nor NOR3 (N1313, N1310, N532, N670);
xor XOR2 (N1314, N1308, N1308);
or OR4 (N1315, N1309, N1272, N517, N1134);
and AND3 (N1316, N1314, N1130, N738);
and AND4 (N1317, N1288, N1272, N653, N804);
nor NOR2 (N1318, N1316, N659);
or OR2 (N1319, N1318, N475);
xor XOR2 (N1320, N1302, N864);
nand NAND2 (N1321, N1315, N57);
or OR3 (N1322, N1317, N549, N1025);
not NOT1 (N1323, N1313);
not NOT1 (N1324, N1294);
buf BUF1 (N1325, N1323);
and AND2 (N1326, N1319, N373);
buf BUF1 (N1327, N1320);
nand NAND3 (N1328, N1305, N159, N686);
xor XOR2 (N1329, N1311, N216);
xor XOR2 (N1330, N1321, N130);
buf BUF1 (N1331, N1325);
nor NOR4 (N1332, N1262, N1, N1037, N1323);
xor XOR2 (N1333, N1328, N906);
xor XOR2 (N1334, N1322, N827);
and AND4 (N1335, N1333, N724, N1055, N795);
and AND3 (N1336, N1334, N634, N1233);
buf BUF1 (N1337, N1329);
not NOT1 (N1338, N1332);
nand NAND4 (N1339, N1326, N1182, N392, N61);
or OR2 (N1340, N1312, N465);
nor NOR2 (N1341, N1338, N433);
xor XOR2 (N1342, N1327, N697);
nor NOR3 (N1343, N1336, N1313, N324);
and AND3 (N1344, N1337, N947, N1191);
or OR3 (N1345, N1341, N792, N92);
nor NOR3 (N1346, N1342, N618, N689);
and AND2 (N1347, N1331, N796);
nand NAND4 (N1348, N1344, N1223, N1334, N1017);
nor NOR2 (N1349, N1345, N738);
or OR2 (N1350, N1339, N961);
nand NAND2 (N1351, N1346, N1317);
or OR2 (N1352, N1340, N326);
buf BUF1 (N1353, N1335);
or OR2 (N1354, N1348, N764);
nand NAND2 (N1355, N1347, N265);
or OR4 (N1356, N1343, N840, N1055, N56);
or OR4 (N1357, N1352, N1198, N601, N24);
and AND3 (N1358, N1351, N182, N616);
nor NOR2 (N1359, N1356, N356);
and AND4 (N1360, N1350, N1292, N992, N390);
xor XOR2 (N1361, N1353, N102);
xor XOR2 (N1362, N1330, N614);
or OR3 (N1363, N1357, N1151, N856);
not NOT1 (N1364, N1354);
xor XOR2 (N1365, N1361, N44);
nor NOR2 (N1366, N1358, N976);
buf BUF1 (N1367, N1349);
xor XOR2 (N1368, N1359, N1006);
xor XOR2 (N1369, N1363, N1300);
nor NOR3 (N1370, N1365, N1097, N834);
or OR2 (N1371, N1360, N8);
or OR2 (N1372, N1366, N437);
buf BUF1 (N1373, N1324);
nor NOR3 (N1374, N1369, N113, N492);
not NOT1 (N1375, N1368);
nand NAND4 (N1376, N1371, N907, N797, N427);
and AND4 (N1377, N1367, N48, N612, N496);
nand NAND2 (N1378, N1364, N402);
not NOT1 (N1379, N1355);
buf BUF1 (N1380, N1374);
nor NOR3 (N1381, N1376, N1161, N284);
or OR4 (N1382, N1380, N1076, N141, N15);
buf BUF1 (N1383, N1378);
nand NAND2 (N1384, N1375, N139);
buf BUF1 (N1385, N1362);
not NOT1 (N1386, N1377);
buf BUF1 (N1387, N1384);
nand NAND2 (N1388, N1382, N155);
buf BUF1 (N1389, N1383);
xor XOR2 (N1390, N1385, N649);
and AND4 (N1391, N1379, N1341, N1203, N36);
and AND3 (N1392, N1386, N1107, N542);
buf BUF1 (N1393, N1381);
buf BUF1 (N1394, N1389);
buf BUF1 (N1395, N1391);
nand NAND3 (N1396, N1388, N350, N759);
not NOT1 (N1397, N1390);
and AND2 (N1398, N1372, N435);
not NOT1 (N1399, N1397);
or OR3 (N1400, N1393, N171, N372);
or OR4 (N1401, N1392, N471, N432, N1204);
nor NOR4 (N1402, N1395, N1228, N199, N1368);
not NOT1 (N1403, N1394);
nor NOR2 (N1404, N1402, N1216);
not NOT1 (N1405, N1400);
or OR3 (N1406, N1398, N684, N654);
not NOT1 (N1407, N1370);
nand NAND2 (N1408, N1403, N241);
and AND2 (N1409, N1404, N163);
and AND2 (N1410, N1407, N282);
nand NAND2 (N1411, N1396, N908);
nand NAND4 (N1412, N1401, N909, N1379, N662);
not NOT1 (N1413, N1410);
nand NAND4 (N1414, N1408, N372, N1403, N909);
nor NOR4 (N1415, N1414, N134, N85, N724);
or OR4 (N1416, N1405, N608, N553, N1406);
xor XOR2 (N1417, N1210, N941);
not NOT1 (N1418, N1409);
nor NOR4 (N1419, N1415, N468, N153, N1356);
or OR2 (N1420, N1416, N233);
and AND4 (N1421, N1413, N249, N456, N904);
buf BUF1 (N1422, N1418);
and AND3 (N1423, N1422, N529, N380);
buf BUF1 (N1424, N1411);
or OR4 (N1425, N1412, N1187, N807, N362);
and AND2 (N1426, N1423, N1179);
not NOT1 (N1427, N1421);
not NOT1 (N1428, N1387);
and AND3 (N1429, N1428, N1166, N241);
nor NOR3 (N1430, N1420, N548, N664);
or OR2 (N1431, N1417, N872);
and AND4 (N1432, N1430, N819, N1, N359);
and AND3 (N1433, N1424, N902, N1336);
and AND2 (N1434, N1426, N194);
xor XOR2 (N1435, N1429, N732);
nand NAND2 (N1436, N1419, N736);
xor XOR2 (N1437, N1427, N55);
buf BUF1 (N1438, N1436);
nand NAND3 (N1439, N1438, N1139, N1034);
and AND2 (N1440, N1435, N14);
not NOT1 (N1441, N1373);
and AND2 (N1442, N1425, N285);
and AND3 (N1443, N1441, N534, N268);
and AND2 (N1444, N1437, N484);
and AND3 (N1445, N1432, N68, N399);
buf BUF1 (N1446, N1440);
nand NAND3 (N1447, N1431, N1396, N606);
not NOT1 (N1448, N1433);
nand NAND4 (N1449, N1442, N547, N911, N259);
xor XOR2 (N1450, N1447, N50);
nor NOR2 (N1451, N1445, N1198);
xor XOR2 (N1452, N1450, N697);
not NOT1 (N1453, N1399);
not NOT1 (N1454, N1452);
and AND3 (N1455, N1448, N349, N57);
or OR3 (N1456, N1443, N1082, N1034);
nand NAND4 (N1457, N1444, N1429, N631, N1092);
buf BUF1 (N1458, N1449);
not NOT1 (N1459, N1457);
nor NOR4 (N1460, N1434, N263, N912, N190);
nand NAND3 (N1461, N1460, N890, N19);
buf BUF1 (N1462, N1458);
buf BUF1 (N1463, N1462);
nor NOR3 (N1464, N1454, N14, N1192);
nor NOR4 (N1465, N1461, N521, N1384, N1286);
buf BUF1 (N1466, N1464);
nor NOR2 (N1467, N1451, N490);
or OR4 (N1468, N1466, N116, N85, N721);
and AND3 (N1469, N1463, N1342, N188);
or OR4 (N1470, N1446, N87, N1250, N1311);
nand NAND4 (N1471, N1470, N277, N907, N1405);
and AND4 (N1472, N1468, N1379, N129, N723);
and AND3 (N1473, N1439, N921, N233);
not NOT1 (N1474, N1453);
or OR3 (N1475, N1472, N762, N583);
xor XOR2 (N1476, N1475, N1076);
buf BUF1 (N1477, N1465);
buf BUF1 (N1478, N1467);
or OR2 (N1479, N1478, N1477);
xor XOR2 (N1480, N65, N1285);
nor NOR2 (N1481, N1459, N982);
xor XOR2 (N1482, N1456, N950);
buf BUF1 (N1483, N1482);
and AND3 (N1484, N1474, N1468, N13);
not NOT1 (N1485, N1471);
not NOT1 (N1486, N1483);
nand NAND3 (N1487, N1484, N397, N342);
and AND4 (N1488, N1469, N133, N32, N1397);
and AND4 (N1489, N1481, N757, N971, N448);
xor XOR2 (N1490, N1488, N917);
not NOT1 (N1491, N1455);
and AND2 (N1492, N1479, N962);
buf BUF1 (N1493, N1476);
buf BUF1 (N1494, N1493);
and AND3 (N1495, N1487, N695, N406);
or OR4 (N1496, N1473, N296, N1053, N54);
buf BUF1 (N1497, N1480);
xor XOR2 (N1498, N1496, N363);
nor NOR3 (N1499, N1495, N999, N1180);
buf BUF1 (N1500, N1489);
buf BUF1 (N1501, N1498);
buf BUF1 (N1502, N1492);
nand NAND3 (N1503, N1501, N1354, N372);
nand NAND4 (N1504, N1494, N952, N1131, N87);
and AND2 (N1505, N1486, N1354);
xor XOR2 (N1506, N1503, N716);
xor XOR2 (N1507, N1490, N1077);
buf BUF1 (N1508, N1502);
buf BUF1 (N1509, N1508);
not NOT1 (N1510, N1499);
or OR3 (N1511, N1491, N714, N1428);
and AND3 (N1512, N1509, N415, N773);
nor NOR4 (N1513, N1505, N187, N376, N243);
nand NAND4 (N1514, N1511, N506, N759, N162);
not NOT1 (N1515, N1500);
or OR3 (N1516, N1510, N747, N1302);
and AND4 (N1517, N1512, N642, N668, N166);
buf BUF1 (N1518, N1514);
nor NOR2 (N1519, N1515, N172);
nand NAND4 (N1520, N1513, N1029, N235, N498);
or OR2 (N1521, N1519, N966);
or OR2 (N1522, N1520, N103);
not NOT1 (N1523, N1516);
and AND3 (N1524, N1522, N1012, N279);
buf BUF1 (N1525, N1517);
not NOT1 (N1526, N1521);
buf BUF1 (N1527, N1485);
and AND2 (N1528, N1525, N598);
not NOT1 (N1529, N1497);
buf BUF1 (N1530, N1527);
xor XOR2 (N1531, N1504, N488);
xor XOR2 (N1532, N1524, N666);
not NOT1 (N1533, N1531);
and AND2 (N1534, N1529, N767);
nand NAND4 (N1535, N1533, N239, N493, N498);
nand NAND2 (N1536, N1528, N745);
buf BUF1 (N1537, N1530);
or OR3 (N1538, N1536, N700, N250);
buf BUF1 (N1539, N1518);
not NOT1 (N1540, N1523);
nor NOR2 (N1541, N1538, N628);
xor XOR2 (N1542, N1506, N714);
nand NAND2 (N1543, N1537, N1429);
not NOT1 (N1544, N1542);
xor XOR2 (N1545, N1507, N1260);
nor NOR2 (N1546, N1535, N947);
or OR3 (N1547, N1543, N68, N1323);
or OR3 (N1548, N1539, N1075, N1185);
xor XOR2 (N1549, N1548, N1);
buf BUF1 (N1550, N1532);
buf BUF1 (N1551, N1544);
xor XOR2 (N1552, N1549, N262);
or OR4 (N1553, N1547, N70, N363, N314);
nand NAND3 (N1554, N1546, N1506, N86);
xor XOR2 (N1555, N1551, N1077);
or OR2 (N1556, N1553, N1065);
nor NOR2 (N1557, N1556, N514);
not NOT1 (N1558, N1526);
or OR2 (N1559, N1540, N965);
and AND4 (N1560, N1550, N1340, N1123, N122);
and AND2 (N1561, N1534, N1242);
not NOT1 (N1562, N1554);
xor XOR2 (N1563, N1560, N1048);
or OR3 (N1564, N1561, N320, N476);
not NOT1 (N1565, N1555);
buf BUF1 (N1566, N1558);
buf BUF1 (N1567, N1565);
nor NOR4 (N1568, N1566, N1392, N372, N267);
nor NOR4 (N1569, N1562, N371, N380, N1515);
not NOT1 (N1570, N1564);
nor NOR2 (N1571, N1570, N1325);
buf BUF1 (N1572, N1557);
and AND3 (N1573, N1541, N592, N630);
nand NAND2 (N1574, N1545, N1510);
not NOT1 (N1575, N1574);
or OR2 (N1576, N1569, N697);
xor XOR2 (N1577, N1568, N1258);
nand NAND3 (N1578, N1571, N981, N734);
or OR4 (N1579, N1577, N1330, N1477, N114);
nor NOR3 (N1580, N1573, N1321, N779);
not NOT1 (N1581, N1575);
nor NOR3 (N1582, N1579, N1100, N892);
not NOT1 (N1583, N1580);
buf BUF1 (N1584, N1581);
xor XOR2 (N1585, N1578, N569);
nand NAND4 (N1586, N1567, N665, N1360, N875);
xor XOR2 (N1587, N1552, N120);
or OR2 (N1588, N1563, N177);
or OR2 (N1589, N1583, N635);
and AND3 (N1590, N1582, N1526, N1250);
xor XOR2 (N1591, N1584, N511);
nor NOR2 (N1592, N1591, N910);
buf BUF1 (N1593, N1586);
nand NAND3 (N1594, N1589, N104, N1473);
nor NOR4 (N1595, N1572, N532, N640, N1173);
xor XOR2 (N1596, N1588, N154);
buf BUF1 (N1597, N1587);
and AND2 (N1598, N1593, N704);
or OR3 (N1599, N1594, N1253, N80);
xor XOR2 (N1600, N1559, N1507);
and AND4 (N1601, N1592, N633, N727, N1108);
nor NOR4 (N1602, N1597, N1179, N1025, N559);
xor XOR2 (N1603, N1599, N1535);
and AND2 (N1604, N1590, N708);
nand NAND3 (N1605, N1598, N562, N31);
nand NAND2 (N1606, N1601, N720);
xor XOR2 (N1607, N1604, N1363);
nor NOR4 (N1608, N1605, N276, N721, N679);
nor NOR3 (N1609, N1595, N337, N498);
and AND2 (N1610, N1609, N943);
and AND4 (N1611, N1576, N943, N1568, N511);
buf BUF1 (N1612, N1606);
or OR2 (N1613, N1612, N815);
or OR3 (N1614, N1603, N99, N995);
and AND3 (N1615, N1608, N171, N1528);
not NOT1 (N1616, N1614);
buf BUF1 (N1617, N1611);
and AND3 (N1618, N1607, N1372, N679);
nand NAND3 (N1619, N1602, N575, N491);
or OR4 (N1620, N1615, N98, N195, N1427);
endmodule