// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N2997,N3010,N3012,N3005,N3004,N3013,N3008,N3009,N3007,N3015;

nand NAND3 (N16, N6, N14, N4);
xor XOR2 (N17, N13, N8);
or OR2 (N18, N15, N17);
nor NOR4 (N19, N17, N8, N8, N13);
and AND2 (N20, N7, N16);
not NOT1 (N21, N12);
nor NOR3 (N22, N11, N5, N9);
xor XOR2 (N23, N8, N21);
buf BUF1 (N24, N12);
buf BUF1 (N25, N20);
buf BUF1 (N26, N22);
xor XOR2 (N27, N1, N21);
or OR4 (N28, N16, N16, N10, N26);
and AND3 (N29, N15, N3, N21);
nand NAND2 (N30, N13, N28);
nor NOR4 (N31, N13, N17, N4, N30);
nor NOR3 (N32, N7, N17, N25);
nand NAND3 (N33, N28, N5, N12);
not NOT1 (N34, N22);
nand NAND3 (N35, N27, N5, N23);
xor XOR2 (N36, N4, N34);
xor XOR2 (N37, N15, N35);
nand NAND4 (N38, N16, N4, N22, N36);
nor NOR3 (N39, N6, N2, N35);
buf BUF1 (N40, N31);
xor XOR2 (N41, N29, N21);
not NOT1 (N42, N24);
not NOT1 (N43, N42);
and AND4 (N44, N41, N18, N32, N38);
nand NAND2 (N45, N18, N11);
xor XOR2 (N46, N6, N14);
buf BUF1 (N47, N20);
nor NOR3 (N48, N40, N3, N22);
nand NAND3 (N49, N47, N18, N22);
not NOT1 (N50, N48);
buf BUF1 (N51, N49);
not NOT1 (N52, N39);
and AND2 (N53, N44, N35);
nor NOR2 (N54, N51, N24);
not NOT1 (N55, N54);
and AND4 (N56, N33, N20, N54, N10);
not NOT1 (N57, N52);
xor XOR2 (N58, N19, N24);
not NOT1 (N59, N37);
nor NOR3 (N60, N46, N24, N12);
nand NAND3 (N61, N50, N27, N45);
nand NAND4 (N62, N18, N40, N4, N23);
and AND2 (N63, N53, N28);
nand NAND3 (N64, N63, N29, N51);
and AND2 (N65, N43, N20);
buf BUF1 (N66, N65);
not NOT1 (N67, N58);
and AND4 (N68, N55, N26, N34, N45);
buf BUF1 (N69, N66);
or OR3 (N70, N68, N21, N58);
nand NAND3 (N71, N61, N24, N24);
and AND3 (N72, N57, N46, N2);
nand NAND3 (N73, N56, N8, N69);
or OR2 (N74, N30, N71);
nand NAND4 (N75, N49, N55, N12, N20);
and AND2 (N76, N72, N18);
or OR3 (N77, N59, N72, N71);
nor NOR2 (N78, N74, N21);
buf BUF1 (N79, N78);
nor NOR4 (N80, N60, N32, N79, N21);
nor NOR2 (N81, N19, N5);
buf BUF1 (N82, N62);
not NOT1 (N83, N67);
not NOT1 (N84, N70);
xor XOR2 (N85, N82, N72);
xor XOR2 (N86, N85, N27);
or OR4 (N87, N77, N72, N85, N13);
and AND2 (N88, N76, N52);
and AND4 (N89, N64, N29, N21, N33);
and AND3 (N90, N81, N50, N12);
nor NOR4 (N91, N87, N58, N28, N19);
nor NOR3 (N92, N90, N23, N75);
not NOT1 (N93, N81);
nand NAND3 (N94, N73, N32, N25);
or OR4 (N95, N86, N53, N30, N65);
nor NOR4 (N96, N88, N65, N70, N43);
nor NOR3 (N97, N96, N94, N89);
xor XOR2 (N98, N9, N46);
nor NOR2 (N99, N31, N14);
nand NAND3 (N100, N99, N80, N26);
or OR4 (N101, N24, N100, N17, N20);
and AND2 (N102, N37, N15);
buf BUF1 (N103, N91);
not NOT1 (N104, N98);
and AND3 (N105, N93, N79, N53);
or OR4 (N106, N83, N3, N41, N37);
and AND2 (N107, N103, N89);
or OR4 (N108, N104, N59, N58, N16);
nor NOR4 (N109, N84, N27, N104, N1);
buf BUF1 (N110, N95);
or OR3 (N111, N110, N8, N57);
xor XOR2 (N112, N92, N106);
xor XOR2 (N113, N47, N16);
nor NOR4 (N114, N111, N67, N40, N53);
xor XOR2 (N115, N108, N21);
or OR2 (N116, N112, N1);
xor XOR2 (N117, N101, N42);
or OR3 (N118, N113, N94, N100);
nor NOR3 (N119, N118, N23, N79);
buf BUF1 (N120, N97);
nand NAND4 (N121, N119, N11, N78, N45);
xor XOR2 (N122, N115, N7);
or OR3 (N123, N117, N67, N55);
nand NAND2 (N124, N107, N90);
not NOT1 (N125, N116);
buf BUF1 (N126, N125);
buf BUF1 (N127, N123);
and AND3 (N128, N124, N75, N103);
not NOT1 (N129, N126);
or OR2 (N130, N109, N117);
xor XOR2 (N131, N128, N125);
and AND4 (N132, N130, N1, N44, N57);
xor XOR2 (N133, N105, N14);
or OR3 (N134, N121, N73, N29);
or OR2 (N135, N129, N61);
nor NOR4 (N136, N132, N124, N75, N19);
and AND4 (N137, N135, N125, N66, N76);
or OR2 (N138, N102, N10);
nand NAND2 (N139, N114, N15);
nand NAND3 (N140, N131, N82, N97);
nor NOR4 (N141, N139, N127, N80, N14);
not NOT1 (N142, N12);
nand NAND3 (N143, N140, N14, N85);
and AND3 (N144, N136, N23, N7);
or OR2 (N145, N122, N17);
xor XOR2 (N146, N120, N76);
and AND3 (N147, N144, N93, N27);
not NOT1 (N148, N142);
buf BUF1 (N149, N133);
xor XOR2 (N150, N146, N127);
buf BUF1 (N151, N141);
and AND3 (N152, N145, N115, N105);
nand NAND2 (N153, N152, N150);
buf BUF1 (N154, N153);
not NOT1 (N155, N120);
not NOT1 (N156, N155);
xor XOR2 (N157, N148, N126);
and AND4 (N158, N137, N23, N33, N99);
and AND2 (N159, N138, N74);
or OR2 (N160, N147, N48);
or OR2 (N161, N143, N63);
nor NOR2 (N162, N134, N148);
nand NAND4 (N163, N160, N149, N38, N93);
not NOT1 (N164, N143);
and AND3 (N165, N151, N35, N76);
not NOT1 (N166, N163);
xor XOR2 (N167, N157, N89);
and AND3 (N168, N162, N55, N105);
xor XOR2 (N169, N165, N167);
or OR4 (N170, N107, N115, N63, N124);
xor XOR2 (N171, N159, N31);
nand NAND3 (N172, N156, N133, N47);
buf BUF1 (N173, N154);
buf BUF1 (N174, N170);
buf BUF1 (N175, N169);
nand NAND4 (N176, N166, N25, N172, N78);
or OR4 (N177, N92, N54, N119, N2);
and AND4 (N178, N158, N175, N25, N175);
and AND4 (N179, N91, N84, N105, N2);
and AND3 (N180, N174, N81, N107);
not NOT1 (N181, N173);
or OR4 (N182, N181, N175, N178, N95);
and AND3 (N183, N154, N148, N11);
not NOT1 (N184, N183);
buf BUF1 (N185, N182);
not NOT1 (N186, N171);
nor NOR4 (N187, N176, N151, N128, N51);
and AND3 (N188, N184, N139, N44);
not NOT1 (N189, N187);
and AND3 (N190, N188, N43, N17);
buf BUF1 (N191, N186);
not NOT1 (N192, N189);
nor NOR2 (N193, N180, N95);
not NOT1 (N194, N161);
xor XOR2 (N195, N164, N41);
or OR2 (N196, N185, N35);
nor NOR4 (N197, N191, N32, N179, N12);
nor NOR3 (N198, N42, N195, N147);
nor NOR2 (N199, N58, N6);
and AND3 (N200, N190, N179, N184);
xor XOR2 (N201, N200, N70);
buf BUF1 (N202, N198);
and AND3 (N203, N199, N51, N160);
buf BUF1 (N204, N201);
or OR3 (N205, N203, N4, N27);
nor NOR3 (N206, N192, N63, N161);
buf BUF1 (N207, N197);
buf BUF1 (N208, N177);
nor NOR3 (N209, N206, N93, N85);
not NOT1 (N210, N207);
nand NAND4 (N211, N204, N92, N110, N69);
not NOT1 (N212, N194);
xor XOR2 (N213, N168, N148);
or OR2 (N214, N205, N158);
nor NOR2 (N215, N212, N55);
and AND3 (N216, N214, N126, N85);
xor XOR2 (N217, N202, N21);
not NOT1 (N218, N216);
and AND2 (N219, N211, N188);
nor NOR3 (N220, N208, N118, N9);
nor NOR2 (N221, N193, N204);
or OR3 (N222, N210, N13, N139);
xor XOR2 (N223, N196, N11);
and AND3 (N224, N219, N15, N89);
buf BUF1 (N225, N220);
buf BUF1 (N226, N221);
and AND3 (N227, N225, N69, N217);
xor XOR2 (N228, N179, N183);
nor NOR2 (N229, N227, N89);
or OR3 (N230, N224, N31, N107);
not NOT1 (N231, N228);
nor NOR4 (N232, N226, N178, N202, N187);
and AND2 (N233, N222, N62);
buf BUF1 (N234, N215);
and AND4 (N235, N231, N65, N10, N127);
buf BUF1 (N236, N209);
xor XOR2 (N237, N218, N191);
not NOT1 (N238, N234);
nor NOR4 (N239, N233, N48, N5, N217);
nor NOR3 (N240, N238, N163, N12);
nand NAND2 (N241, N237, N99);
buf BUF1 (N242, N229);
xor XOR2 (N243, N242, N202);
and AND4 (N244, N243, N15, N47, N59);
nand NAND3 (N245, N230, N149, N211);
and AND2 (N246, N235, N140);
xor XOR2 (N247, N239, N245);
nand NAND3 (N248, N16, N93, N163);
xor XOR2 (N249, N232, N169);
and AND3 (N250, N247, N69, N78);
or OR4 (N251, N250, N94, N76, N66);
xor XOR2 (N252, N240, N199);
buf BUF1 (N253, N252);
not NOT1 (N254, N246);
nor NOR4 (N255, N236, N157, N16, N12);
not NOT1 (N256, N251);
nand NAND3 (N257, N254, N57, N1);
xor XOR2 (N258, N241, N236);
nor NOR4 (N259, N249, N3, N31, N216);
buf BUF1 (N260, N257);
and AND4 (N261, N244, N224, N113, N189);
not NOT1 (N262, N259);
nor NOR3 (N263, N253, N22, N9);
nand NAND3 (N264, N255, N209, N43);
nand NAND3 (N265, N260, N232, N201);
nor NOR4 (N266, N213, N182, N136, N178);
not NOT1 (N267, N266);
or OR4 (N268, N265, N206, N12, N161);
xor XOR2 (N269, N256, N250);
buf BUF1 (N270, N263);
and AND3 (N271, N223, N258, N184);
nor NOR4 (N272, N4, N13, N36, N245);
buf BUF1 (N273, N272);
xor XOR2 (N274, N273, N20);
nor NOR4 (N275, N267, N204, N234, N50);
nand NAND3 (N276, N268, N118, N167);
or OR3 (N277, N274, N166, N116);
not NOT1 (N278, N271);
buf BUF1 (N279, N270);
nor NOR2 (N280, N275, N18);
or OR4 (N281, N277, N263, N165, N182);
buf BUF1 (N282, N262);
and AND3 (N283, N269, N32, N101);
or OR3 (N284, N279, N66, N78);
nor NOR2 (N285, N261, N172);
xor XOR2 (N286, N264, N100);
xor XOR2 (N287, N281, N77);
and AND4 (N288, N280, N186, N16, N150);
nand NAND2 (N289, N284, N176);
buf BUF1 (N290, N282);
or OR3 (N291, N283, N197, N201);
or OR4 (N292, N285, N30, N168, N29);
nor NOR3 (N293, N248, N233, N145);
or OR3 (N294, N278, N200, N141);
nand NAND2 (N295, N290, N176);
xor XOR2 (N296, N288, N214);
buf BUF1 (N297, N295);
or OR3 (N298, N286, N157, N70);
nor NOR2 (N299, N293, N9);
or OR2 (N300, N289, N236);
not NOT1 (N301, N276);
and AND2 (N302, N298, N83);
nand NAND3 (N303, N300, N218, N104);
and AND4 (N304, N296, N293, N300, N226);
xor XOR2 (N305, N304, N1);
or OR4 (N306, N297, N252, N295, N84);
xor XOR2 (N307, N294, N159);
buf BUF1 (N308, N292);
nor NOR3 (N309, N299, N166, N221);
nor NOR2 (N310, N307, N233);
xor XOR2 (N311, N303, N282);
or OR4 (N312, N309, N250, N303, N8);
not NOT1 (N313, N311);
or OR2 (N314, N302, N276);
nor NOR4 (N315, N306, N27, N135, N172);
and AND4 (N316, N305, N274, N101, N234);
buf BUF1 (N317, N291);
not NOT1 (N318, N287);
nor NOR4 (N319, N310, N117, N205, N268);
nand NAND3 (N320, N301, N307, N183);
and AND3 (N321, N314, N157, N210);
not NOT1 (N322, N308);
and AND2 (N323, N319, N254);
buf BUF1 (N324, N320);
buf BUF1 (N325, N318);
nor NOR3 (N326, N313, N132, N114);
buf BUF1 (N327, N316);
and AND2 (N328, N322, N200);
xor XOR2 (N329, N312, N121);
buf BUF1 (N330, N329);
xor XOR2 (N331, N323, N237);
xor XOR2 (N332, N324, N71);
nand NAND3 (N333, N317, N188, N61);
or OR3 (N334, N325, N177, N313);
and AND3 (N335, N315, N208, N210);
nor NOR2 (N336, N335, N112);
not NOT1 (N337, N321);
nand NAND2 (N338, N333, N109);
xor XOR2 (N339, N331, N323);
or OR3 (N340, N328, N79, N127);
xor XOR2 (N341, N338, N77);
or OR4 (N342, N334, N5, N124, N119);
or OR4 (N343, N340, N6, N261, N277);
xor XOR2 (N344, N330, N188);
xor XOR2 (N345, N341, N69);
xor XOR2 (N346, N343, N217);
xor XOR2 (N347, N345, N343);
nor NOR4 (N348, N332, N149, N144, N201);
and AND2 (N349, N337, N246);
and AND2 (N350, N336, N282);
and AND2 (N351, N339, N249);
not NOT1 (N352, N347);
xor XOR2 (N353, N350, N178);
and AND4 (N354, N346, N185, N236, N220);
buf BUF1 (N355, N351);
xor XOR2 (N356, N355, N16);
or OR4 (N357, N326, N64, N116, N66);
not NOT1 (N358, N352);
xor XOR2 (N359, N358, N72);
xor XOR2 (N360, N348, N18);
nor NOR4 (N361, N327, N90, N115, N30);
nand NAND3 (N362, N353, N187, N4);
not NOT1 (N363, N357);
nand NAND2 (N364, N360, N50);
or OR2 (N365, N359, N250);
xor XOR2 (N366, N342, N202);
or OR2 (N367, N363, N297);
buf BUF1 (N368, N356);
or OR3 (N369, N354, N101, N303);
or OR4 (N370, N349, N170, N200, N52);
not NOT1 (N371, N366);
buf BUF1 (N372, N361);
xor XOR2 (N373, N362, N239);
buf BUF1 (N374, N344);
not NOT1 (N375, N373);
buf BUF1 (N376, N370);
xor XOR2 (N377, N369, N75);
buf BUF1 (N378, N364);
xor XOR2 (N379, N378, N278);
nand NAND4 (N380, N376, N228, N212, N144);
not NOT1 (N381, N372);
nor NOR2 (N382, N367, N300);
and AND3 (N383, N375, N249, N36);
nand NAND2 (N384, N382, N301);
nand NAND4 (N385, N379, N211, N161, N107);
xor XOR2 (N386, N368, N246);
nor NOR4 (N387, N377, N256, N370, N280);
nor NOR4 (N388, N381, N152, N264, N32);
not NOT1 (N389, N380);
or OR2 (N390, N386, N34);
and AND4 (N391, N389, N265, N241, N105);
xor XOR2 (N392, N374, N163);
not NOT1 (N393, N384);
not NOT1 (N394, N365);
nor NOR4 (N395, N385, N110, N255, N40);
xor XOR2 (N396, N388, N176);
or OR3 (N397, N395, N272, N365);
not NOT1 (N398, N391);
and AND4 (N399, N396, N333, N241, N332);
or OR2 (N400, N393, N7);
buf BUF1 (N401, N383);
nand NAND3 (N402, N387, N128, N327);
and AND3 (N403, N390, N3, N295);
buf BUF1 (N404, N394);
xor XOR2 (N405, N399, N129);
xor XOR2 (N406, N392, N12);
and AND4 (N407, N371, N107, N109, N223);
or OR4 (N408, N407, N297, N329, N258);
buf BUF1 (N409, N400);
nor NOR3 (N410, N403, N273, N342);
and AND4 (N411, N408, N279, N235, N401);
xor XOR2 (N412, N156, N52);
nor NOR4 (N413, N410, N127, N370, N265);
nand NAND3 (N414, N411, N79, N252);
not NOT1 (N415, N398);
nand NAND2 (N416, N414, N25);
buf BUF1 (N417, N413);
and AND2 (N418, N409, N172);
or OR4 (N419, N415, N134, N86, N109);
nand NAND3 (N420, N406, N27, N214);
nand NAND4 (N421, N412, N335, N375, N226);
nor NOR4 (N422, N405, N417, N262, N303);
nor NOR4 (N423, N83, N343, N80, N187);
nand NAND2 (N424, N418, N180);
or OR2 (N425, N423, N6);
xor XOR2 (N426, N419, N417);
xor XOR2 (N427, N424, N15);
or OR4 (N428, N425, N180, N403, N6);
nand NAND4 (N429, N397, N92, N150, N65);
xor XOR2 (N430, N402, N211);
nand NAND4 (N431, N429, N129, N380, N51);
xor XOR2 (N432, N427, N372);
nand NAND3 (N433, N422, N142, N9);
not NOT1 (N434, N431);
or OR2 (N435, N421, N166);
or OR4 (N436, N430, N295, N28, N101);
or OR2 (N437, N426, N59);
nor NOR2 (N438, N436, N52);
not NOT1 (N439, N428);
or OR4 (N440, N439, N338, N290, N298);
nand NAND2 (N441, N433, N286);
buf BUF1 (N442, N434);
xor XOR2 (N443, N404, N434);
buf BUF1 (N444, N416);
not NOT1 (N445, N441);
nor NOR3 (N446, N442, N13, N138);
and AND2 (N447, N440, N61);
buf BUF1 (N448, N447);
xor XOR2 (N449, N420, N351);
buf BUF1 (N450, N435);
buf BUF1 (N451, N449);
not NOT1 (N452, N432);
not NOT1 (N453, N450);
xor XOR2 (N454, N444, N445);
nand NAND3 (N455, N432, N135, N326);
nand NAND2 (N456, N454, N329);
and AND3 (N457, N452, N381, N210);
not NOT1 (N458, N438);
nor NOR4 (N459, N437, N145, N241, N420);
xor XOR2 (N460, N446, N409);
nand NAND4 (N461, N443, N130, N163, N94);
xor XOR2 (N462, N448, N321);
buf BUF1 (N463, N458);
and AND2 (N464, N460, N458);
xor XOR2 (N465, N455, N214);
and AND2 (N466, N451, N402);
xor XOR2 (N467, N466, N415);
or OR2 (N468, N462, N447);
and AND4 (N469, N459, N70, N391, N468);
nor NOR4 (N470, N290, N197, N432, N210);
nor NOR4 (N471, N467, N152, N194, N447);
buf BUF1 (N472, N471);
and AND3 (N473, N464, N106, N215);
or OR4 (N474, N456, N317, N126, N411);
and AND4 (N475, N473, N240, N400, N403);
not NOT1 (N476, N469);
nand NAND3 (N477, N461, N191, N434);
xor XOR2 (N478, N457, N453);
and AND2 (N479, N285, N85);
nand NAND2 (N480, N470, N278);
xor XOR2 (N481, N472, N102);
nand NAND3 (N482, N481, N315, N97);
and AND3 (N483, N463, N372, N159);
buf BUF1 (N484, N477);
not NOT1 (N485, N465);
and AND4 (N486, N474, N345, N49, N470);
and AND2 (N487, N485, N300);
and AND2 (N488, N476, N123);
buf BUF1 (N489, N484);
not NOT1 (N490, N475);
nor NOR3 (N491, N489, N267, N1);
nor NOR3 (N492, N491, N389, N55);
or OR3 (N493, N479, N42, N313);
or OR3 (N494, N488, N82, N40);
nand NAND3 (N495, N493, N73, N361);
not NOT1 (N496, N482);
or OR3 (N497, N483, N35, N465);
or OR2 (N498, N492, N107);
xor XOR2 (N499, N498, N433);
buf BUF1 (N500, N495);
buf BUF1 (N501, N478);
and AND2 (N502, N480, N95);
buf BUF1 (N503, N486);
xor XOR2 (N504, N503, N456);
and AND3 (N505, N502, N301, N122);
not NOT1 (N506, N499);
nor NOR2 (N507, N501, N433);
and AND2 (N508, N504, N315);
xor XOR2 (N509, N500, N388);
nor NOR4 (N510, N494, N357, N387, N123);
xor XOR2 (N511, N490, N457);
or OR2 (N512, N509, N34);
and AND4 (N513, N496, N33, N415, N25);
nor NOR3 (N514, N506, N343, N84);
nor NOR2 (N515, N514, N194);
or OR4 (N516, N515, N330, N55, N401);
nor NOR2 (N517, N516, N271);
nor NOR3 (N518, N510, N513, N24);
and AND2 (N519, N186, N369);
nand NAND2 (N520, N519, N423);
xor XOR2 (N521, N517, N299);
and AND4 (N522, N512, N328, N104, N342);
buf BUF1 (N523, N508);
and AND4 (N524, N487, N35, N132, N183);
nor NOR4 (N525, N524, N266, N143, N7);
and AND3 (N526, N525, N221, N358);
nand NAND2 (N527, N523, N457);
buf BUF1 (N528, N507);
or OR2 (N529, N497, N342);
buf BUF1 (N530, N518);
nor NOR3 (N531, N529, N279, N273);
nor NOR2 (N532, N522, N324);
buf BUF1 (N533, N505);
xor XOR2 (N534, N527, N54);
nand NAND4 (N535, N511, N88, N365, N289);
and AND3 (N536, N526, N277, N1);
nand NAND3 (N537, N520, N454, N244);
or OR2 (N538, N536, N471);
buf BUF1 (N539, N534);
or OR4 (N540, N521, N477, N362, N394);
buf BUF1 (N541, N535);
nand NAND3 (N542, N538, N106, N248);
buf BUF1 (N543, N528);
xor XOR2 (N544, N530, N314);
or OR3 (N545, N544, N469, N446);
xor XOR2 (N546, N543, N409);
or OR3 (N547, N537, N441, N29);
not NOT1 (N548, N539);
nor NOR3 (N549, N547, N258, N395);
or OR2 (N550, N546, N85);
or OR2 (N551, N533, N312);
buf BUF1 (N552, N549);
nor NOR4 (N553, N531, N209, N465, N65);
and AND4 (N554, N532, N119, N192, N251);
and AND3 (N555, N541, N91, N341);
xor XOR2 (N556, N551, N137);
nor NOR4 (N557, N555, N135, N100, N555);
xor XOR2 (N558, N550, N508);
xor XOR2 (N559, N548, N62);
nor NOR3 (N560, N545, N308, N394);
or OR2 (N561, N540, N354);
nand NAND2 (N562, N554, N263);
or OR2 (N563, N560, N206);
xor XOR2 (N564, N562, N38);
xor XOR2 (N565, N556, N229);
buf BUF1 (N566, N561);
or OR4 (N567, N557, N26, N107, N172);
not NOT1 (N568, N559);
or OR4 (N569, N553, N180, N219, N53);
or OR3 (N570, N569, N21, N511);
xor XOR2 (N571, N566, N497);
and AND3 (N572, N563, N518, N422);
nand NAND4 (N573, N558, N369, N372, N161);
nand NAND2 (N574, N542, N544);
nor NOR4 (N575, N574, N316, N452, N104);
or OR2 (N576, N552, N566);
xor XOR2 (N577, N575, N63);
nand NAND3 (N578, N576, N489, N186);
not NOT1 (N579, N570);
and AND3 (N580, N571, N305, N21);
xor XOR2 (N581, N579, N279);
not NOT1 (N582, N580);
or OR3 (N583, N578, N327, N449);
xor XOR2 (N584, N565, N296);
buf BUF1 (N585, N564);
or OR3 (N586, N582, N40, N258);
xor XOR2 (N587, N584, N541);
not NOT1 (N588, N572);
and AND3 (N589, N567, N9, N549);
not NOT1 (N590, N573);
xor XOR2 (N591, N585, N72);
buf BUF1 (N592, N588);
nand NAND3 (N593, N577, N489, N35);
or OR2 (N594, N591, N93);
nand NAND4 (N595, N587, N150, N202, N311);
buf BUF1 (N596, N586);
xor XOR2 (N597, N581, N356);
buf BUF1 (N598, N592);
buf BUF1 (N599, N583);
buf BUF1 (N600, N589);
nand NAND4 (N601, N599, N104, N320, N9);
not NOT1 (N602, N595);
nand NAND4 (N603, N596, N213, N267, N364);
and AND2 (N604, N602, N400);
or OR4 (N605, N568, N380, N206, N361);
buf BUF1 (N606, N590);
xor XOR2 (N607, N597, N175);
nand NAND4 (N608, N604, N515, N341, N96);
nand NAND3 (N609, N598, N460, N235);
nor NOR3 (N610, N593, N16, N359);
and AND4 (N611, N606, N384, N204, N594);
xor XOR2 (N612, N328, N356);
buf BUF1 (N613, N612);
and AND2 (N614, N613, N466);
or OR3 (N615, N605, N4, N290);
buf BUF1 (N616, N615);
xor XOR2 (N617, N601, N523);
not NOT1 (N618, N616);
and AND2 (N619, N610, N494);
xor XOR2 (N620, N608, N167);
and AND4 (N621, N607, N178, N594, N217);
nor NOR2 (N622, N617, N241);
xor XOR2 (N623, N609, N36);
nor NOR4 (N624, N611, N188, N246, N85);
and AND3 (N625, N618, N40, N52);
nor NOR3 (N626, N619, N36, N441);
or OR3 (N627, N621, N506, N573);
and AND2 (N628, N622, N311);
xor XOR2 (N629, N600, N417);
or OR3 (N630, N614, N296, N576);
nor NOR2 (N631, N629, N549);
nor NOR4 (N632, N620, N372, N305, N474);
xor XOR2 (N633, N625, N307);
nor NOR2 (N634, N627, N501);
and AND2 (N635, N626, N79);
nor NOR2 (N636, N635, N80);
buf BUF1 (N637, N630);
nand NAND3 (N638, N637, N515, N299);
xor XOR2 (N639, N603, N555);
or OR4 (N640, N638, N348, N67, N141);
buf BUF1 (N641, N640);
and AND3 (N642, N639, N181, N125);
or OR4 (N643, N623, N484, N287, N375);
nor NOR3 (N644, N628, N274, N454);
and AND4 (N645, N631, N597, N225, N638);
nand NAND4 (N646, N644, N258, N176, N420);
or OR3 (N647, N641, N376, N413);
xor XOR2 (N648, N632, N488);
xor XOR2 (N649, N643, N537);
not NOT1 (N650, N648);
nand NAND4 (N651, N649, N416, N305, N225);
or OR3 (N652, N642, N462, N172);
or OR2 (N653, N647, N353);
and AND4 (N654, N645, N342, N297, N7);
nand NAND3 (N655, N652, N276, N343);
and AND3 (N656, N634, N109, N398);
or OR3 (N657, N653, N485, N515);
xor XOR2 (N658, N651, N127);
not NOT1 (N659, N646);
nor NOR4 (N660, N658, N508, N19, N230);
and AND2 (N661, N656, N605);
xor XOR2 (N662, N657, N311);
nand NAND2 (N663, N650, N348);
xor XOR2 (N664, N655, N107);
buf BUF1 (N665, N654);
xor XOR2 (N666, N636, N519);
xor XOR2 (N667, N664, N443);
xor XOR2 (N668, N663, N81);
nand NAND3 (N669, N633, N301, N393);
buf BUF1 (N670, N659);
or OR2 (N671, N661, N318);
nor NOR2 (N672, N671, N370);
xor XOR2 (N673, N669, N471);
and AND2 (N674, N667, N305);
buf BUF1 (N675, N668);
not NOT1 (N676, N660);
nand NAND2 (N677, N666, N529);
buf BUF1 (N678, N674);
and AND2 (N679, N675, N54);
not NOT1 (N680, N676);
xor XOR2 (N681, N665, N108);
and AND3 (N682, N672, N226, N181);
or OR4 (N683, N677, N661, N419, N373);
buf BUF1 (N684, N681);
buf BUF1 (N685, N624);
nor NOR3 (N686, N680, N153, N312);
or OR2 (N687, N684, N549);
xor XOR2 (N688, N685, N479);
buf BUF1 (N689, N678);
nor NOR2 (N690, N673, N410);
or OR4 (N691, N689, N368, N225, N552);
and AND4 (N692, N683, N450, N84, N486);
buf BUF1 (N693, N670);
nand NAND2 (N694, N679, N481);
and AND4 (N695, N693, N582, N491, N271);
and AND4 (N696, N682, N79, N131, N531);
nand NAND3 (N697, N695, N190, N144);
and AND2 (N698, N696, N272);
or OR3 (N699, N697, N316, N666);
nor NOR3 (N700, N690, N428, N389);
buf BUF1 (N701, N699);
nand NAND4 (N702, N687, N355, N652, N87);
nand NAND3 (N703, N688, N392, N201);
nand NAND4 (N704, N702, N456, N236, N299);
nor NOR2 (N705, N703, N448);
not NOT1 (N706, N705);
xor XOR2 (N707, N698, N590);
nor NOR3 (N708, N694, N135, N351);
and AND4 (N709, N701, N137, N597, N666);
or OR3 (N710, N686, N294, N560);
xor XOR2 (N711, N691, N244);
not NOT1 (N712, N711);
and AND3 (N713, N704, N55, N581);
xor XOR2 (N714, N710, N299);
or OR3 (N715, N700, N73, N82);
nor NOR3 (N716, N707, N532, N42);
nor NOR4 (N717, N714, N652, N657, N397);
and AND3 (N718, N713, N450, N275);
nand NAND4 (N719, N716, N100, N191, N86);
not NOT1 (N720, N709);
or OR4 (N721, N715, N388, N95, N468);
nor NOR4 (N722, N712, N298, N502, N451);
or OR2 (N723, N718, N627);
and AND4 (N724, N723, N338, N103, N508);
buf BUF1 (N725, N692);
buf BUF1 (N726, N725);
xor XOR2 (N727, N720, N584);
and AND2 (N728, N722, N450);
and AND2 (N729, N724, N142);
not NOT1 (N730, N717);
nor NOR2 (N731, N662, N522);
nand NAND3 (N732, N731, N248, N343);
buf BUF1 (N733, N728);
nor NOR2 (N734, N733, N389);
nor NOR3 (N735, N719, N614, N547);
xor XOR2 (N736, N735, N589);
nor NOR4 (N737, N727, N222, N27, N574);
xor XOR2 (N738, N729, N458);
and AND2 (N739, N736, N432);
nor NOR3 (N740, N739, N328, N340);
nand NAND2 (N741, N732, N389);
not NOT1 (N742, N726);
nand NAND3 (N743, N740, N596, N269);
nor NOR4 (N744, N721, N390, N384, N196);
nand NAND4 (N745, N708, N459, N550, N286);
nor NOR2 (N746, N738, N611);
xor XOR2 (N747, N730, N149);
or OR4 (N748, N746, N331, N387, N195);
nand NAND2 (N749, N745, N211);
nor NOR2 (N750, N748, N196);
nor NOR3 (N751, N743, N229, N569);
not NOT1 (N752, N749);
or OR4 (N753, N747, N205, N141, N103);
nor NOR4 (N754, N737, N358, N37, N679);
nor NOR3 (N755, N741, N2, N707);
xor XOR2 (N756, N751, N662);
nand NAND4 (N757, N753, N706, N271, N587);
nand NAND3 (N758, N202, N747, N529);
and AND3 (N759, N744, N259, N360);
nor NOR3 (N760, N754, N44, N249);
xor XOR2 (N761, N752, N103);
nand NAND3 (N762, N757, N124, N178);
and AND4 (N763, N750, N440, N193, N754);
nor NOR3 (N764, N758, N200, N502);
or OR2 (N765, N764, N534);
not NOT1 (N766, N759);
buf BUF1 (N767, N755);
nor NOR3 (N768, N734, N356, N725);
nor NOR3 (N769, N760, N488, N217);
buf BUF1 (N770, N756);
xor XOR2 (N771, N763, N574);
not NOT1 (N772, N762);
and AND4 (N773, N765, N113, N421, N91);
xor XOR2 (N774, N773, N452);
xor XOR2 (N775, N770, N327);
xor XOR2 (N776, N774, N153);
not NOT1 (N777, N771);
nor NOR3 (N778, N772, N673, N511);
nor NOR2 (N779, N778, N294);
nor NOR2 (N780, N777, N554);
xor XOR2 (N781, N768, N412);
xor XOR2 (N782, N775, N248);
xor XOR2 (N783, N776, N140);
buf BUF1 (N784, N780);
or OR2 (N785, N781, N127);
xor XOR2 (N786, N761, N509);
and AND2 (N787, N742, N567);
and AND3 (N788, N785, N572, N5);
and AND3 (N789, N783, N726, N380);
xor XOR2 (N790, N767, N177);
not NOT1 (N791, N787);
nor NOR2 (N792, N790, N777);
and AND4 (N793, N782, N601, N40, N737);
buf BUF1 (N794, N793);
not NOT1 (N795, N769);
or OR4 (N796, N791, N322, N525, N274);
and AND3 (N797, N794, N540, N47);
nand NAND4 (N798, N795, N631, N325, N231);
xor XOR2 (N799, N784, N143);
xor XOR2 (N800, N796, N645);
and AND2 (N801, N797, N350);
nor NOR4 (N802, N766, N609, N423, N643);
not NOT1 (N803, N800);
nand NAND3 (N804, N803, N775, N755);
nor NOR3 (N805, N802, N59, N162);
or OR3 (N806, N804, N362, N293);
not NOT1 (N807, N799);
buf BUF1 (N808, N805);
and AND3 (N809, N806, N425, N131);
nand NAND3 (N810, N789, N739, N610);
buf BUF1 (N811, N792);
or OR3 (N812, N779, N703, N87);
nand NAND4 (N813, N798, N480, N483, N216);
xor XOR2 (N814, N808, N506);
xor XOR2 (N815, N811, N785);
xor XOR2 (N816, N814, N150);
not NOT1 (N817, N812);
and AND3 (N818, N801, N536, N133);
buf BUF1 (N819, N818);
nand NAND2 (N820, N807, N398);
and AND2 (N821, N813, N336);
xor XOR2 (N822, N786, N714);
nand NAND4 (N823, N816, N122, N91, N645);
and AND3 (N824, N810, N508, N364);
nor NOR4 (N825, N823, N294, N809, N252);
and AND4 (N826, N304, N443, N482, N602);
not NOT1 (N827, N826);
xor XOR2 (N828, N825, N578);
buf BUF1 (N829, N817);
or OR4 (N830, N827, N69, N92, N107);
nand NAND4 (N831, N788, N569, N426, N679);
and AND4 (N832, N815, N292, N705, N168);
not NOT1 (N833, N824);
xor XOR2 (N834, N833, N619);
not NOT1 (N835, N831);
not NOT1 (N836, N821);
not NOT1 (N837, N832);
and AND2 (N838, N836, N3);
xor XOR2 (N839, N834, N657);
and AND2 (N840, N838, N90);
nand NAND4 (N841, N829, N665, N89, N232);
or OR2 (N842, N819, N462);
buf BUF1 (N843, N839);
buf BUF1 (N844, N828);
or OR3 (N845, N837, N604, N143);
or OR2 (N846, N845, N515);
nor NOR4 (N847, N820, N599, N404, N698);
xor XOR2 (N848, N843, N133);
buf BUF1 (N849, N846);
nor NOR2 (N850, N844, N576);
xor XOR2 (N851, N849, N71);
nand NAND3 (N852, N840, N63, N197);
not NOT1 (N853, N830);
nor NOR3 (N854, N822, N290, N367);
xor XOR2 (N855, N841, N396);
xor XOR2 (N856, N850, N523);
not NOT1 (N857, N853);
nor NOR4 (N858, N856, N147, N140, N39);
nor NOR2 (N859, N847, N288);
not NOT1 (N860, N842);
not NOT1 (N861, N848);
nor NOR4 (N862, N860, N495, N633, N185);
xor XOR2 (N863, N855, N521);
or OR3 (N864, N835, N654, N533);
not NOT1 (N865, N851);
and AND3 (N866, N859, N779, N262);
and AND2 (N867, N865, N570);
or OR4 (N868, N862, N240, N414, N506);
or OR2 (N869, N858, N632);
not NOT1 (N870, N868);
buf BUF1 (N871, N861);
nor NOR3 (N872, N857, N568, N165);
buf BUF1 (N873, N863);
or OR4 (N874, N867, N864, N678, N107);
or OR3 (N875, N806, N39, N25);
nor NOR3 (N876, N852, N837, N666);
xor XOR2 (N877, N869, N495);
and AND2 (N878, N872, N9);
xor XOR2 (N879, N875, N830);
buf BUF1 (N880, N871);
nand NAND2 (N881, N854, N652);
nand NAND4 (N882, N881, N127, N309, N390);
xor XOR2 (N883, N870, N158);
nor NOR2 (N884, N866, N445);
and AND4 (N885, N880, N241, N71, N148);
buf BUF1 (N886, N884);
or OR2 (N887, N879, N78);
or OR2 (N888, N887, N185);
nand NAND3 (N889, N878, N80, N183);
buf BUF1 (N890, N873);
nand NAND3 (N891, N883, N520, N675);
or OR3 (N892, N890, N219, N751);
nand NAND4 (N893, N882, N66, N286, N823);
not NOT1 (N894, N891);
nand NAND3 (N895, N876, N220, N86);
buf BUF1 (N896, N886);
or OR2 (N897, N893, N273);
or OR2 (N898, N874, N567);
nor NOR4 (N899, N896, N529, N679, N220);
nand NAND3 (N900, N885, N586, N136);
nor NOR3 (N901, N895, N517, N212);
nand NAND3 (N902, N888, N549, N173);
and AND3 (N903, N902, N229, N104);
or OR4 (N904, N897, N728, N215, N843);
buf BUF1 (N905, N901);
buf BUF1 (N906, N894);
or OR4 (N907, N904, N276, N850, N787);
and AND2 (N908, N907, N840);
nor NOR2 (N909, N899, N367);
nand NAND2 (N910, N909, N220);
nand NAND3 (N911, N892, N15, N666);
not NOT1 (N912, N911);
and AND3 (N913, N889, N469, N434);
and AND2 (N914, N898, N627);
or OR3 (N915, N912, N654, N96);
not NOT1 (N916, N913);
nand NAND4 (N917, N914, N115, N102, N475);
not NOT1 (N918, N905);
or OR2 (N919, N900, N326);
buf BUF1 (N920, N906);
buf BUF1 (N921, N920);
nor NOR2 (N922, N919, N668);
buf BUF1 (N923, N877);
and AND4 (N924, N923, N395, N470, N202);
xor XOR2 (N925, N916, N667);
or OR4 (N926, N924, N600, N147, N265);
not NOT1 (N927, N918);
buf BUF1 (N928, N903);
buf BUF1 (N929, N921);
not NOT1 (N930, N929);
nor NOR4 (N931, N922, N21, N781, N685);
not NOT1 (N932, N930);
nand NAND3 (N933, N910, N671, N5);
not NOT1 (N934, N915);
and AND4 (N935, N908, N669, N153, N548);
not NOT1 (N936, N917);
nor NOR4 (N937, N933, N640, N890, N544);
and AND3 (N938, N935, N215, N289);
and AND2 (N939, N927, N895);
or OR4 (N940, N928, N375, N935, N444);
and AND4 (N941, N939, N168, N96, N146);
not NOT1 (N942, N937);
buf BUF1 (N943, N932);
nand NAND4 (N944, N925, N875, N752, N465);
buf BUF1 (N945, N926);
nand NAND3 (N946, N945, N741, N694);
not NOT1 (N947, N944);
buf BUF1 (N948, N938);
nand NAND4 (N949, N931, N301, N242, N453);
and AND4 (N950, N947, N515, N367, N103);
buf BUF1 (N951, N950);
and AND4 (N952, N951, N712, N203, N900);
not NOT1 (N953, N934);
not NOT1 (N954, N941);
and AND2 (N955, N942, N481);
xor XOR2 (N956, N940, N558);
xor XOR2 (N957, N943, N612);
not NOT1 (N958, N953);
or OR2 (N959, N956, N515);
nor NOR4 (N960, N949, N683, N411, N197);
and AND4 (N961, N958, N600, N404, N156);
not NOT1 (N962, N959);
not NOT1 (N963, N960);
nor NOR3 (N964, N952, N189, N103);
not NOT1 (N965, N957);
and AND2 (N966, N954, N232);
xor XOR2 (N967, N946, N672);
nor NOR4 (N968, N965, N814, N252, N21);
and AND2 (N969, N967, N950);
nand NAND2 (N970, N968, N189);
buf BUF1 (N971, N936);
not NOT1 (N972, N971);
nor NOR4 (N973, N963, N243, N780, N539);
buf BUF1 (N974, N969);
or OR3 (N975, N962, N845, N679);
nand NAND4 (N976, N975, N418, N464, N258);
buf BUF1 (N977, N955);
xor XOR2 (N978, N961, N698);
or OR2 (N979, N978, N475);
nand NAND4 (N980, N973, N370, N165, N105);
not NOT1 (N981, N972);
or OR4 (N982, N980, N129, N731, N776);
buf BUF1 (N983, N977);
nand NAND3 (N984, N970, N594, N927);
buf BUF1 (N985, N979);
not NOT1 (N986, N981);
nand NAND2 (N987, N986, N230);
not NOT1 (N988, N964);
nor NOR2 (N989, N985, N526);
nand NAND4 (N990, N987, N510, N464, N894);
nand NAND2 (N991, N974, N672);
nor NOR4 (N992, N990, N696, N308, N376);
xor XOR2 (N993, N984, N78);
nor NOR2 (N994, N991, N972);
and AND2 (N995, N948, N606);
or OR4 (N996, N992, N618, N471, N915);
or OR2 (N997, N994, N751);
nor NOR2 (N998, N993, N742);
or OR3 (N999, N982, N36, N477);
and AND4 (N1000, N995, N412, N214, N466);
xor XOR2 (N1001, N976, N167);
nand NAND3 (N1002, N996, N422, N24);
nor NOR3 (N1003, N1002, N987, N915);
nand NAND2 (N1004, N999, N328);
or OR4 (N1005, N998, N648, N260, N330);
buf BUF1 (N1006, N997);
not NOT1 (N1007, N966);
nor NOR3 (N1008, N1004, N345, N505);
and AND3 (N1009, N1001, N587, N275);
nand NAND3 (N1010, N1006, N702, N179);
nor NOR4 (N1011, N1007, N453, N624, N733);
or OR4 (N1012, N1008, N715, N838, N916);
xor XOR2 (N1013, N1009, N320);
buf BUF1 (N1014, N983);
buf BUF1 (N1015, N1012);
or OR2 (N1016, N1015, N185);
nor NOR2 (N1017, N1005, N362);
buf BUF1 (N1018, N1013);
and AND3 (N1019, N1000, N872, N272);
or OR4 (N1020, N1011, N744, N793, N169);
and AND3 (N1021, N1018, N489, N928);
and AND3 (N1022, N1017, N192, N512);
xor XOR2 (N1023, N1003, N739);
nor NOR4 (N1024, N1022, N313, N461, N507);
and AND3 (N1025, N1020, N692, N125);
or OR2 (N1026, N1019, N358);
and AND4 (N1027, N1016, N248, N1011, N584);
nor NOR2 (N1028, N1010, N1015);
nor NOR2 (N1029, N1027, N884);
nor NOR2 (N1030, N1025, N714);
nor NOR2 (N1031, N1024, N974);
and AND3 (N1032, N1031, N709, N596);
xor XOR2 (N1033, N1021, N287);
or OR3 (N1034, N989, N407, N453);
and AND4 (N1035, N1026, N221, N703, N641);
xor XOR2 (N1036, N1035, N63);
xor XOR2 (N1037, N988, N89);
nand NAND3 (N1038, N1032, N921, N593);
xor XOR2 (N1039, N1029, N104);
xor XOR2 (N1040, N1034, N986);
nand NAND4 (N1041, N1040, N561, N467, N813);
and AND3 (N1042, N1014, N125, N862);
not NOT1 (N1043, N1028);
and AND2 (N1044, N1033, N441);
nand NAND3 (N1045, N1036, N18, N521);
nand NAND2 (N1046, N1023, N518);
not NOT1 (N1047, N1042);
not NOT1 (N1048, N1038);
nand NAND4 (N1049, N1046, N600, N2, N812);
nand NAND4 (N1050, N1041, N41, N441, N483);
not NOT1 (N1051, N1045);
nor NOR3 (N1052, N1037, N139, N246);
or OR4 (N1053, N1049, N408, N843, N28);
buf BUF1 (N1054, N1050);
not NOT1 (N1055, N1052);
nor NOR2 (N1056, N1051, N574);
nand NAND3 (N1057, N1056, N348, N637);
xor XOR2 (N1058, N1054, N869);
or OR3 (N1059, N1044, N861, N989);
or OR4 (N1060, N1048, N106, N908, N451);
xor XOR2 (N1061, N1057, N581);
nand NAND4 (N1062, N1039, N1034, N233, N850);
xor XOR2 (N1063, N1060, N84);
xor XOR2 (N1064, N1053, N725);
nand NAND4 (N1065, N1061, N830, N337, N714);
nand NAND4 (N1066, N1065, N106, N142, N471);
or OR3 (N1067, N1055, N844, N716);
not NOT1 (N1068, N1062);
buf BUF1 (N1069, N1063);
and AND4 (N1070, N1067, N883, N866, N651);
xor XOR2 (N1071, N1047, N326);
nor NOR4 (N1072, N1070, N634, N44, N370);
and AND4 (N1073, N1059, N190, N887, N599);
nand NAND2 (N1074, N1043, N1019);
or OR3 (N1075, N1074, N419, N324);
not NOT1 (N1076, N1064);
buf BUF1 (N1077, N1075);
nand NAND4 (N1078, N1073, N711, N883, N313);
not NOT1 (N1079, N1069);
and AND2 (N1080, N1071, N253);
nor NOR3 (N1081, N1080, N7, N111);
buf BUF1 (N1082, N1030);
or OR4 (N1083, N1079, N465, N198, N800);
nor NOR2 (N1084, N1066, N365);
and AND4 (N1085, N1068, N32, N306, N993);
not NOT1 (N1086, N1081);
or OR4 (N1087, N1082, N909, N538, N704);
not NOT1 (N1088, N1084);
nand NAND3 (N1089, N1072, N75, N147);
nor NOR2 (N1090, N1083, N273);
buf BUF1 (N1091, N1090);
nand NAND2 (N1092, N1087, N588);
buf BUF1 (N1093, N1088);
not NOT1 (N1094, N1093);
not NOT1 (N1095, N1085);
nand NAND2 (N1096, N1092, N192);
nor NOR3 (N1097, N1096, N917, N644);
nand NAND3 (N1098, N1078, N470, N897);
and AND3 (N1099, N1095, N421, N635);
nand NAND2 (N1100, N1089, N527);
or OR4 (N1101, N1097, N665, N962, N218);
or OR2 (N1102, N1101, N576);
nor NOR2 (N1103, N1102, N132);
buf BUF1 (N1104, N1091);
nand NAND2 (N1105, N1058, N37);
or OR4 (N1106, N1103, N211, N125, N234);
buf BUF1 (N1107, N1086);
nor NOR4 (N1108, N1099, N636, N105, N93);
nand NAND2 (N1109, N1098, N736);
xor XOR2 (N1110, N1108, N19);
nand NAND2 (N1111, N1077, N779);
nand NAND2 (N1112, N1100, N604);
buf BUF1 (N1113, N1076);
nor NOR3 (N1114, N1113, N277, N401);
buf BUF1 (N1115, N1109);
and AND3 (N1116, N1104, N242, N328);
xor XOR2 (N1117, N1106, N838);
not NOT1 (N1118, N1112);
and AND3 (N1119, N1111, N765, N47);
not NOT1 (N1120, N1105);
xor XOR2 (N1121, N1115, N473);
not NOT1 (N1122, N1119);
or OR2 (N1123, N1116, N638);
buf BUF1 (N1124, N1094);
and AND2 (N1125, N1124, N555);
nor NOR3 (N1126, N1123, N858, N119);
xor XOR2 (N1127, N1126, N192);
nor NOR4 (N1128, N1118, N981, N881, N361);
or OR3 (N1129, N1107, N1004, N1106);
not NOT1 (N1130, N1122);
buf BUF1 (N1131, N1125);
or OR3 (N1132, N1114, N614, N767);
not NOT1 (N1133, N1117);
buf BUF1 (N1134, N1110);
not NOT1 (N1135, N1120);
and AND2 (N1136, N1134, N521);
and AND2 (N1137, N1133, N1090);
not NOT1 (N1138, N1129);
buf BUF1 (N1139, N1135);
nor NOR2 (N1140, N1127, N58);
buf BUF1 (N1141, N1132);
and AND4 (N1142, N1140, N717, N326, N940);
and AND4 (N1143, N1131, N244, N77, N929);
xor XOR2 (N1144, N1130, N867);
and AND3 (N1145, N1141, N618, N207);
and AND4 (N1146, N1121, N606, N1060, N205);
nor NOR4 (N1147, N1139, N909, N228, N167);
nand NAND3 (N1148, N1143, N442, N481);
and AND2 (N1149, N1136, N681);
and AND4 (N1150, N1149, N923, N579, N594);
and AND2 (N1151, N1138, N581);
xor XOR2 (N1152, N1142, N243);
buf BUF1 (N1153, N1148);
or OR2 (N1154, N1153, N671);
buf BUF1 (N1155, N1150);
or OR2 (N1156, N1154, N435);
nor NOR4 (N1157, N1152, N411, N484, N910);
nand NAND2 (N1158, N1156, N617);
nor NOR4 (N1159, N1145, N193, N323, N997);
nor NOR3 (N1160, N1137, N1101, N80);
or OR2 (N1161, N1159, N962);
or OR4 (N1162, N1161, N731, N589, N944);
xor XOR2 (N1163, N1160, N588);
nor NOR2 (N1164, N1157, N24);
nor NOR2 (N1165, N1162, N1034);
and AND4 (N1166, N1164, N954, N91, N21);
nor NOR3 (N1167, N1155, N89, N949);
and AND4 (N1168, N1147, N908, N989, N844);
nor NOR3 (N1169, N1151, N352, N868);
nor NOR3 (N1170, N1128, N602, N369);
xor XOR2 (N1171, N1146, N724);
not NOT1 (N1172, N1158);
nand NAND4 (N1173, N1144, N130, N304, N524);
nand NAND2 (N1174, N1163, N380);
not NOT1 (N1175, N1171);
or OR4 (N1176, N1175, N1077, N727, N836);
not NOT1 (N1177, N1174);
buf BUF1 (N1178, N1165);
and AND4 (N1179, N1168, N548, N679, N845);
or OR2 (N1180, N1167, N1066);
buf BUF1 (N1181, N1178);
buf BUF1 (N1182, N1166);
buf BUF1 (N1183, N1170);
buf BUF1 (N1184, N1180);
not NOT1 (N1185, N1179);
buf BUF1 (N1186, N1173);
not NOT1 (N1187, N1169);
xor XOR2 (N1188, N1172, N158);
nor NOR2 (N1189, N1176, N780);
buf BUF1 (N1190, N1183);
not NOT1 (N1191, N1185);
nor NOR3 (N1192, N1189, N297, N569);
or OR4 (N1193, N1181, N966, N1146, N783);
nand NAND2 (N1194, N1188, N963);
not NOT1 (N1195, N1177);
not NOT1 (N1196, N1186);
buf BUF1 (N1197, N1196);
nand NAND4 (N1198, N1184, N1007, N269, N1087);
xor XOR2 (N1199, N1187, N770);
not NOT1 (N1200, N1199);
and AND4 (N1201, N1200, N1141, N528, N632);
nand NAND2 (N1202, N1192, N543);
nor NOR2 (N1203, N1190, N651);
nor NOR2 (N1204, N1182, N708);
nand NAND3 (N1205, N1204, N384, N1054);
and AND4 (N1206, N1195, N184, N904, N1);
not NOT1 (N1207, N1201);
nand NAND2 (N1208, N1197, N565);
or OR2 (N1209, N1191, N359);
buf BUF1 (N1210, N1207);
buf BUF1 (N1211, N1208);
and AND2 (N1212, N1198, N1143);
buf BUF1 (N1213, N1194);
and AND3 (N1214, N1210, N1213, N361);
nand NAND2 (N1215, N537, N321);
and AND4 (N1216, N1214, N1039, N1019, N1086);
nor NOR2 (N1217, N1212, N957);
not NOT1 (N1218, N1215);
not NOT1 (N1219, N1218);
xor XOR2 (N1220, N1216, N1024);
and AND2 (N1221, N1203, N303);
nand NAND2 (N1222, N1206, N995);
xor XOR2 (N1223, N1217, N874);
xor XOR2 (N1224, N1220, N272);
buf BUF1 (N1225, N1224);
not NOT1 (N1226, N1222);
or OR3 (N1227, N1202, N752, N644);
nand NAND2 (N1228, N1226, N298);
or OR2 (N1229, N1223, N1170);
xor XOR2 (N1230, N1193, N341);
buf BUF1 (N1231, N1205);
or OR4 (N1232, N1231, N668, N317, N557);
not NOT1 (N1233, N1228);
nand NAND4 (N1234, N1232, N1211, N1181, N869);
nand NAND2 (N1235, N1229, N1060);
not NOT1 (N1236, N901);
or OR4 (N1237, N1236, N844, N557, N275);
nand NAND2 (N1238, N1227, N166);
not NOT1 (N1239, N1225);
not NOT1 (N1240, N1221);
nor NOR4 (N1241, N1235, N72, N554, N394);
and AND2 (N1242, N1237, N141);
nand NAND2 (N1243, N1233, N524);
not NOT1 (N1244, N1234);
and AND2 (N1245, N1209, N498);
not NOT1 (N1246, N1241);
or OR4 (N1247, N1240, N65, N437, N90);
and AND4 (N1248, N1247, N626, N1068, N932);
nand NAND2 (N1249, N1239, N460);
not NOT1 (N1250, N1219);
and AND4 (N1251, N1250, N208, N472, N837);
nand NAND3 (N1252, N1251, N1132, N839);
not NOT1 (N1253, N1244);
nor NOR2 (N1254, N1242, N532);
nand NAND4 (N1255, N1248, N1183, N638, N387);
not NOT1 (N1256, N1254);
xor XOR2 (N1257, N1245, N1197);
xor XOR2 (N1258, N1253, N787);
nand NAND3 (N1259, N1257, N84, N708);
not NOT1 (N1260, N1246);
buf BUF1 (N1261, N1238);
and AND2 (N1262, N1258, N619);
xor XOR2 (N1263, N1252, N938);
not NOT1 (N1264, N1256);
xor XOR2 (N1265, N1255, N624);
or OR2 (N1266, N1230, N739);
and AND3 (N1267, N1260, N1138, N994);
buf BUF1 (N1268, N1262);
nand NAND3 (N1269, N1263, N278, N823);
and AND3 (N1270, N1267, N660, N140);
buf BUF1 (N1271, N1264);
or OR4 (N1272, N1269, N673, N49, N657);
xor XOR2 (N1273, N1259, N700);
and AND4 (N1274, N1243, N1111, N208, N116);
not NOT1 (N1275, N1268);
nand NAND2 (N1276, N1249, N401);
buf BUF1 (N1277, N1274);
nor NOR2 (N1278, N1271, N1033);
and AND2 (N1279, N1266, N611);
xor XOR2 (N1280, N1278, N466);
and AND4 (N1281, N1273, N932, N64, N955);
buf BUF1 (N1282, N1275);
not NOT1 (N1283, N1279);
buf BUF1 (N1284, N1272);
nor NOR3 (N1285, N1277, N1025, N671);
xor XOR2 (N1286, N1281, N654);
or OR2 (N1287, N1285, N777);
or OR4 (N1288, N1283, N1090, N589, N595);
not NOT1 (N1289, N1280);
xor XOR2 (N1290, N1284, N954);
buf BUF1 (N1291, N1265);
xor XOR2 (N1292, N1286, N1132);
not NOT1 (N1293, N1288);
not NOT1 (N1294, N1287);
nor NOR3 (N1295, N1289, N1141, N110);
nand NAND2 (N1296, N1276, N600);
nor NOR3 (N1297, N1296, N1194, N305);
nor NOR4 (N1298, N1290, N800, N1292, N1044);
xor XOR2 (N1299, N914, N412);
or OR4 (N1300, N1270, N474, N535, N183);
xor XOR2 (N1301, N1293, N952);
or OR4 (N1302, N1282, N275, N1184, N413);
xor XOR2 (N1303, N1302, N923);
and AND2 (N1304, N1297, N50);
nand NAND3 (N1305, N1303, N1129, N936);
nand NAND4 (N1306, N1305, N40, N1148, N1253);
nand NAND4 (N1307, N1298, N692, N401, N622);
nor NOR3 (N1308, N1306, N471, N1049);
nand NAND2 (N1309, N1304, N837);
nor NOR2 (N1310, N1309, N198);
or OR2 (N1311, N1307, N1307);
and AND4 (N1312, N1261, N63, N776, N1256);
or OR2 (N1313, N1312, N1194);
xor XOR2 (N1314, N1294, N252);
nor NOR2 (N1315, N1314, N545);
xor XOR2 (N1316, N1300, N1159);
nand NAND4 (N1317, N1301, N941, N1037, N174);
not NOT1 (N1318, N1291);
and AND2 (N1319, N1308, N1071);
nor NOR3 (N1320, N1295, N780, N1102);
nor NOR4 (N1321, N1320, N693, N194, N725);
or OR2 (N1322, N1313, N1247);
xor XOR2 (N1323, N1316, N767);
nor NOR4 (N1324, N1310, N335, N1273, N735);
buf BUF1 (N1325, N1323);
xor XOR2 (N1326, N1311, N131);
buf BUF1 (N1327, N1324);
and AND4 (N1328, N1322, N1109, N821, N328);
and AND4 (N1329, N1319, N982, N929, N587);
and AND3 (N1330, N1318, N1263, N1041);
and AND2 (N1331, N1328, N545);
nand NAND3 (N1332, N1315, N1014, N220);
not NOT1 (N1333, N1327);
and AND3 (N1334, N1321, N1140, N5);
buf BUF1 (N1335, N1332);
nor NOR3 (N1336, N1326, N1307, N187);
xor XOR2 (N1337, N1335, N737);
buf BUF1 (N1338, N1325);
nor NOR3 (N1339, N1331, N928, N558);
and AND4 (N1340, N1336, N780, N267, N717);
nor NOR2 (N1341, N1333, N367);
not NOT1 (N1342, N1337);
and AND2 (N1343, N1338, N463);
buf BUF1 (N1344, N1342);
buf BUF1 (N1345, N1344);
nand NAND2 (N1346, N1341, N346);
or OR3 (N1347, N1346, N528, N3);
or OR3 (N1348, N1343, N566, N800);
or OR2 (N1349, N1334, N652);
xor XOR2 (N1350, N1349, N126);
nand NAND2 (N1351, N1299, N386);
and AND3 (N1352, N1347, N343, N1113);
nand NAND2 (N1353, N1350, N55);
and AND4 (N1354, N1353, N345, N83, N707);
buf BUF1 (N1355, N1329);
and AND4 (N1356, N1317, N1156, N1011, N479);
buf BUF1 (N1357, N1339);
and AND4 (N1358, N1354, N967, N568, N925);
xor XOR2 (N1359, N1358, N1307);
or OR4 (N1360, N1359, N844, N299, N683);
nand NAND4 (N1361, N1356, N922, N1230, N900);
buf BUF1 (N1362, N1361);
nand NAND4 (N1363, N1348, N727, N818, N1188);
nand NAND4 (N1364, N1330, N969, N549, N560);
buf BUF1 (N1365, N1352);
or OR4 (N1366, N1364, N589, N1279, N487);
xor XOR2 (N1367, N1360, N257);
and AND4 (N1368, N1351, N714, N438, N867);
nor NOR4 (N1369, N1366, N453, N510, N1316);
xor XOR2 (N1370, N1367, N1344);
buf BUF1 (N1371, N1370);
not NOT1 (N1372, N1355);
not NOT1 (N1373, N1357);
or OR3 (N1374, N1363, N307, N44);
not NOT1 (N1375, N1345);
not NOT1 (N1376, N1371);
nand NAND2 (N1377, N1373, N1207);
and AND2 (N1378, N1362, N787);
nor NOR4 (N1379, N1375, N1118, N1098, N730);
buf BUF1 (N1380, N1340);
nor NOR3 (N1381, N1380, N414, N549);
nor NOR4 (N1382, N1372, N797, N1304, N1210);
or OR3 (N1383, N1378, N52, N1099);
nand NAND2 (N1384, N1383, N1035);
or OR3 (N1385, N1379, N1364, N650);
xor XOR2 (N1386, N1368, N270);
or OR4 (N1387, N1374, N1260, N679, N1014);
xor XOR2 (N1388, N1369, N335);
and AND4 (N1389, N1384, N493, N41, N1099);
buf BUF1 (N1390, N1385);
not NOT1 (N1391, N1377);
or OR2 (N1392, N1390, N17);
not NOT1 (N1393, N1391);
nand NAND4 (N1394, N1388, N217, N1185, N644);
xor XOR2 (N1395, N1382, N368);
buf BUF1 (N1396, N1386);
nor NOR3 (N1397, N1393, N539, N408);
buf BUF1 (N1398, N1389);
or OR3 (N1399, N1387, N1366, N1168);
and AND4 (N1400, N1399, N938, N573, N611);
buf BUF1 (N1401, N1400);
and AND3 (N1402, N1365, N1127, N315);
and AND3 (N1403, N1394, N1063, N902);
nand NAND3 (N1404, N1376, N293, N328);
and AND4 (N1405, N1395, N712, N1297, N821);
nor NOR4 (N1406, N1402, N911, N1401, N869);
nand NAND3 (N1407, N891, N850, N1169);
xor XOR2 (N1408, N1396, N210);
nand NAND2 (N1409, N1405, N466);
xor XOR2 (N1410, N1404, N649);
not NOT1 (N1411, N1410);
xor XOR2 (N1412, N1408, N1352);
buf BUF1 (N1413, N1406);
xor XOR2 (N1414, N1413, N60);
buf BUF1 (N1415, N1407);
or OR4 (N1416, N1397, N1007, N778, N344);
buf BUF1 (N1417, N1414);
xor XOR2 (N1418, N1381, N1063);
nor NOR4 (N1419, N1411, N640, N75, N718);
and AND2 (N1420, N1416, N870);
and AND2 (N1421, N1419, N431);
or OR3 (N1422, N1418, N809, N755);
xor XOR2 (N1423, N1403, N7);
and AND4 (N1424, N1412, N617, N949, N687);
and AND2 (N1425, N1398, N1);
nor NOR3 (N1426, N1421, N550, N427);
xor XOR2 (N1427, N1424, N1061);
nand NAND2 (N1428, N1427, N1033);
buf BUF1 (N1429, N1428);
or OR3 (N1430, N1409, N413, N920);
and AND4 (N1431, N1425, N1302, N44, N431);
or OR4 (N1432, N1431, N683, N1146, N424);
xor XOR2 (N1433, N1417, N965);
nor NOR3 (N1434, N1426, N1083, N1090);
nor NOR3 (N1435, N1430, N175, N1240);
buf BUF1 (N1436, N1423);
nor NOR3 (N1437, N1432, N126, N1412);
buf BUF1 (N1438, N1420);
nand NAND3 (N1439, N1435, N479, N152);
nand NAND3 (N1440, N1429, N461, N674);
nand NAND2 (N1441, N1436, N85);
or OR4 (N1442, N1415, N308, N532, N484);
buf BUF1 (N1443, N1422);
nor NOR3 (N1444, N1440, N9, N1317);
or OR3 (N1445, N1434, N867, N82);
xor XOR2 (N1446, N1445, N174);
buf BUF1 (N1447, N1444);
buf BUF1 (N1448, N1447);
nor NOR3 (N1449, N1442, N170, N191);
or OR3 (N1450, N1392, N1105, N905);
not NOT1 (N1451, N1446);
nor NOR2 (N1452, N1433, N1223);
not NOT1 (N1453, N1438);
and AND2 (N1454, N1452, N824);
nor NOR4 (N1455, N1437, N62, N972, N854);
or OR2 (N1456, N1441, N1060);
nor NOR2 (N1457, N1439, N1246);
xor XOR2 (N1458, N1455, N458);
not NOT1 (N1459, N1456);
and AND2 (N1460, N1448, N361);
buf BUF1 (N1461, N1457);
not NOT1 (N1462, N1458);
nor NOR2 (N1463, N1453, N479);
xor XOR2 (N1464, N1449, N1167);
buf BUF1 (N1465, N1464);
nand NAND2 (N1466, N1443, N371);
buf BUF1 (N1467, N1454);
not NOT1 (N1468, N1459);
not NOT1 (N1469, N1461);
xor XOR2 (N1470, N1450, N988);
not NOT1 (N1471, N1470);
xor XOR2 (N1472, N1467, N946);
xor XOR2 (N1473, N1471, N433);
or OR2 (N1474, N1466, N460);
buf BUF1 (N1475, N1462);
buf BUF1 (N1476, N1474);
buf BUF1 (N1477, N1468);
not NOT1 (N1478, N1460);
or OR2 (N1479, N1478, N801);
or OR3 (N1480, N1451, N983, N349);
nand NAND4 (N1481, N1472, N65, N933, N15);
or OR2 (N1482, N1463, N142);
not NOT1 (N1483, N1482);
or OR3 (N1484, N1475, N179, N1209);
not NOT1 (N1485, N1469);
nor NOR4 (N1486, N1465, N1, N188, N901);
and AND2 (N1487, N1481, N1127);
and AND2 (N1488, N1476, N1390);
or OR2 (N1489, N1485, N383);
nor NOR4 (N1490, N1489, N483, N1157, N807);
and AND3 (N1491, N1486, N630, N1111);
or OR2 (N1492, N1473, N1002);
nand NAND2 (N1493, N1483, N658);
buf BUF1 (N1494, N1488);
xor XOR2 (N1495, N1477, N1203);
nor NOR3 (N1496, N1480, N552, N1456);
not NOT1 (N1497, N1484);
not NOT1 (N1498, N1479);
and AND2 (N1499, N1498, N175);
not NOT1 (N1500, N1496);
and AND3 (N1501, N1493, N303, N1446);
or OR4 (N1502, N1500, N1468, N388, N618);
xor XOR2 (N1503, N1499, N267);
nand NAND3 (N1504, N1490, N1131, N138);
nand NAND2 (N1505, N1502, N10);
xor XOR2 (N1506, N1505, N1212);
nand NAND4 (N1507, N1497, N650, N325, N358);
buf BUF1 (N1508, N1491);
not NOT1 (N1509, N1494);
or OR3 (N1510, N1487, N1272, N565);
nor NOR2 (N1511, N1501, N1344);
xor XOR2 (N1512, N1507, N970);
xor XOR2 (N1513, N1506, N138);
or OR3 (N1514, N1495, N469, N317);
buf BUF1 (N1515, N1513);
nor NOR2 (N1516, N1492, N291);
buf BUF1 (N1517, N1511);
or OR4 (N1518, N1503, N1128, N174, N873);
and AND4 (N1519, N1516, N1262, N746, N1329);
nand NAND3 (N1520, N1512, N1006, N8);
nor NOR3 (N1521, N1518, N1135, N225);
nor NOR4 (N1522, N1514, N913, N457, N569);
xor XOR2 (N1523, N1519, N1223);
not NOT1 (N1524, N1520);
and AND4 (N1525, N1510, N1366, N1298, N998);
not NOT1 (N1526, N1508);
nor NOR4 (N1527, N1524, N1100, N296, N1435);
and AND3 (N1528, N1527, N819, N14);
nor NOR2 (N1529, N1528, N868);
nor NOR2 (N1530, N1517, N337);
buf BUF1 (N1531, N1529);
nand NAND4 (N1532, N1531, N913, N500, N1513);
and AND4 (N1533, N1521, N1371, N671, N1289);
or OR3 (N1534, N1515, N1207, N1266);
nand NAND4 (N1535, N1533, N1024, N337, N139);
not NOT1 (N1536, N1532);
not NOT1 (N1537, N1535);
buf BUF1 (N1538, N1536);
not NOT1 (N1539, N1523);
and AND4 (N1540, N1534, N36, N509, N639);
and AND4 (N1541, N1504, N620, N1324, N1390);
or OR4 (N1542, N1537, N266, N312, N763);
buf BUF1 (N1543, N1538);
xor XOR2 (N1544, N1543, N539);
not NOT1 (N1545, N1526);
and AND2 (N1546, N1522, N1123);
or OR4 (N1547, N1539, N719, N1342, N322);
nand NAND4 (N1548, N1525, N1520, N414, N1312);
or OR2 (N1549, N1547, N1292);
or OR2 (N1550, N1549, N502);
nor NOR4 (N1551, N1550, N50, N618, N1492);
nor NOR2 (N1552, N1541, N1052);
not NOT1 (N1553, N1509);
xor XOR2 (N1554, N1530, N1173);
not NOT1 (N1555, N1554);
buf BUF1 (N1556, N1548);
or OR4 (N1557, N1555, N536, N110, N1448);
nand NAND3 (N1558, N1544, N162, N630);
xor XOR2 (N1559, N1556, N363);
not NOT1 (N1560, N1546);
nand NAND3 (N1561, N1542, N383, N1273);
not NOT1 (N1562, N1560);
nor NOR2 (N1563, N1540, N1401);
nand NAND3 (N1564, N1559, N950, N116);
xor XOR2 (N1565, N1551, N1109);
and AND4 (N1566, N1564, N784, N31, N1238);
or OR4 (N1567, N1565, N1077, N564, N54);
nand NAND4 (N1568, N1567, N910, N1549, N330);
nor NOR3 (N1569, N1545, N1195, N318);
nor NOR4 (N1570, N1569, N402, N622, N1534);
buf BUF1 (N1571, N1552);
not NOT1 (N1572, N1558);
xor XOR2 (N1573, N1570, N1550);
and AND4 (N1574, N1572, N149, N583, N1439);
nand NAND2 (N1575, N1553, N654);
buf BUF1 (N1576, N1574);
nor NOR4 (N1577, N1571, N625, N1247, N1061);
or OR2 (N1578, N1563, N1165);
nor NOR4 (N1579, N1562, N435, N1134, N796);
or OR4 (N1580, N1568, N1185, N1477, N554);
or OR3 (N1581, N1561, N10, N564);
not NOT1 (N1582, N1579);
xor XOR2 (N1583, N1566, N313);
buf BUF1 (N1584, N1582);
not NOT1 (N1585, N1584);
xor XOR2 (N1586, N1577, N1455);
or OR3 (N1587, N1573, N508, N796);
or OR4 (N1588, N1581, N1382, N900, N1308);
and AND2 (N1589, N1583, N1284);
buf BUF1 (N1590, N1588);
and AND3 (N1591, N1576, N1380, N1173);
xor XOR2 (N1592, N1590, N813);
or OR4 (N1593, N1587, N31, N482, N968);
buf BUF1 (N1594, N1591);
nand NAND3 (N1595, N1557, N983, N429);
and AND2 (N1596, N1595, N704);
not NOT1 (N1597, N1592);
nor NOR3 (N1598, N1578, N817, N690);
not NOT1 (N1599, N1598);
or OR4 (N1600, N1580, N317, N264, N1498);
not NOT1 (N1601, N1600);
not NOT1 (N1602, N1586);
and AND2 (N1603, N1593, N1494);
or OR2 (N1604, N1597, N481);
xor XOR2 (N1605, N1604, N733);
nand NAND2 (N1606, N1575, N41);
or OR4 (N1607, N1603, N884, N1446, N775);
or OR3 (N1608, N1594, N550, N85);
xor XOR2 (N1609, N1601, N1427);
not NOT1 (N1610, N1589);
and AND3 (N1611, N1605, N757, N71);
xor XOR2 (N1612, N1606, N114);
nor NOR3 (N1613, N1602, N1395, N667);
nand NAND3 (N1614, N1610, N645, N1042);
not NOT1 (N1615, N1609);
nor NOR2 (N1616, N1599, N1270);
nand NAND3 (N1617, N1614, N660, N940);
nand NAND4 (N1618, N1596, N124, N1081, N516);
not NOT1 (N1619, N1615);
nor NOR2 (N1620, N1616, N1164);
or OR4 (N1621, N1618, N107, N413, N273);
not NOT1 (N1622, N1607);
nand NAND2 (N1623, N1585, N575);
nand NAND3 (N1624, N1612, N1615, N893);
and AND4 (N1625, N1617, N1380, N1574, N758);
nand NAND2 (N1626, N1624, N1153);
buf BUF1 (N1627, N1621);
xor XOR2 (N1628, N1625, N290);
or OR3 (N1629, N1613, N1582, N1512);
nor NOR2 (N1630, N1619, N55);
or OR3 (N1631, N1611, N1374, N693);
or OR3 (N1632, N1626, N156, N1000);
or OR2 (N1633, N1620, N496);
nor NOR3 (N1634, N1623, N297, N246);
not NOT1 (N1635, N1632);
nor NOR3 (N1636, N1622, N59, N742);
buf BUF1 (N1637, N1634);
buf BUF1 (N1638, N1608);
nand NAND3 (N1639, N1627, N352, N1619);
nand NAND2 (N1640, N1636, N394);
nor NOR2 (N1641, N1637, N1014);
nor NOR2 (N1642, N1630, N1587);
buf BUF1 (N1643, N1638);
or OR4 (N1644, N1643, N717, N1069, N26);
or OR4 (N1645, N1628, N349, N415, N1550);
and AND4 (N1646, N1640, N357, N157, N841);
nor NOR3 (N1647, N1633, N1600, N447);
buf BUF1 (N1648, N1647);
not NOT1 (N1649, N1629);
nand NAND3 (N1650, N1648, N1630, N645);
nor NOR2 (N1651, N1646, N1112);
not NOT1 (N1652, N1641);
xor XOR2 (N1653, N1652, N677);
xor XOR2 (N1654, N1639, N606);
nand NAND4 (N1655, N1642, N941, N1321, N449);
or OR2 (N1656, N1651, N1651);
xor XOR2 (N1657, N1645, N710);
or OR4 (N1658, N1653, N116, N1442, N237);
buf BUF1 (N1659, N1650);
xor XOR2 (N1660, N1657, N1280);
nor NOR2 (N1661, N1635, N1298);
xor XOR2 (N1662, N1644, N976);
and AND2 (N1663, N1662, N1071);
buf BUF1 (N1664, N1649);
xor XOR2 (N1665, N1661, N1259);
xor XOR2 (N1666, N1659, N1473);
or OR2 (N1667, N1664, N843);
or OR3 (N1668, N1667, N162, N817);
xor XOR2 (N1669, N1654, N594);
and AND3 (N1670, N1631, N1378, N379);
not NOT1 (N1671, N1660);
xor XOR2 (N1672, N1656, N769);
and AND2 (N1673, N1665, N1159);
xor XOR2 (N1674, N1673, N1339);
xor XOR2 (N1675, N1663, N6);
and AND2 (N1676, N1658, N506);
buf BUF1 (N1677, N1669);
and AND3 (N1678, N1666, N352, N1654);
and AND4 (N1679, N1675, N1568, N1393, N379);
not NOT1 (N1680, N1655);
or OR4 (N1681, N1674, N801, N952, N424);
and AND2 (N1682, N1676, N707);
or OR4 (N1683, N1671, N776, N122, N1612);
nor NOR3 (N1684, N1681, N1614, N1322);
buf BUF1 (N1685, N1668);
or OR2 (N1686, N1680, N1566);
xor XOR2 (N1687, N1686, N354);
xor XOR2 (N1688, N1685, N458);
xor XOR2 (N1689, N1672, N456);
xor XOR2 (N1690, N1670, N552);
nand NAND3 (N1691, N1684, N1534, N1580);
nand NAND3 (N1692, N1691, N1167, N1397);
or OR4 (N1693, N1690, N52, N1166, N502);
not NOT1 (N1694, N1679);
nor NOR4 (N1695, N1682, N809, N1388, N924);
and AND3 (N1696, N1693, N308, N197);
not NOT1 (N1697, N1694);
xor XOR2 (N1698, N1678, N302);
xor XOR2 (N1699, N1696, N405);
buf BUF1 (N1700, N1698);
buf BUF1 (N1701, N1688);
not NOT1 (N1702, N1677);
nand NAND2 (N1703, N1687, N1067);
not NOT1 (N1704, N1703);
buf BUF1 (N1705, N1692);
xor XOR2 (N1706, N1689, N1410);
buf BUF1 (N1707, N1706);
not NOT1 (N1708, N1683);
or OR3 (N1709, N1702, N97, N1697);
or OR3 (N1710, N680, N1508, N908);
nand NAND3 (N1711, N1708, N856, N738);
xor XOR2 (N1712, N1701, N755);
nor NOR2 (N1713, N1704, N1444);
nor NOR3 (N1714, N1713, N1022, N602);
nand NAND2 (N1715, N1710, N15);
not NOT1 (N1716, N1695);
not NOT1 (N1717, N1711);
buf BUF1 (N1718, N1715);
not NOT1 (N1719, N1705);
not NOT1 (N1720, N1707);
nor NOR3 (N1721, N1712, N158, N799);
nand NAND3 (N1722, N1719, N167, N1125);
not NOT1 (N1723, N1721);
not NOT1 (N1724, N1717);
buf BUF1 (N1725, N1720);
xor XOR2 (N1726, N1725, N1258);
not NOT1 (N1727, N1723);
not NOT1 (N1728, N1709);
buf BUF1 (N1729, N1727);
nor NOR3 (N1730, N1724, N518, N106);
buf BUF1 (N1731, N1699);
not NOT1 (N1732, N1726);
or OR3 (N1733, N1730, N888, N503);
nor NOR3 (N1734, N1716, N158, N619);
and AND3 (N1735, N1732, N1066, N618);
nor NOR4 (N1736, N1729, N1335, N202, N860);
buf BUF1 (N1737, N1728);
or OR4 (N1738, N1735, N1170, N1614, N924);
buf BUF1 (N1739, N1718);
buf BUF1 (N1740, N1734);
buf BUF1 (N1741, N1731);
xor XOR2 (N1742, N1733, N1326);
nor NOR2 (N1743, N1737, N54);
buf BUF1 (N1744, N1739);
buf BUF1 (N1745, N1743);
and AND2 (N1746, N1714, N1319);
nor NOR3 (N1747, N1700, N1220, N780);
buf BUF1 (N1748, N1742);
xor XOR2 (N1749, N1747, N368);
buf BUF1 (N1750, N1741);
nor NOR2 (N1751, N1746, N94);
not NOT1 (N1752, N1722);
nor NOR2 (N1753, N1748, N398);
buf BUF1 (N1754, N1738);
nand NAND3 (N1755, N1754, N230, N716);
not NOT1 (N1756, N1753);
not NOT1 (N1757, N1744);
not NOT1 (N1758, N1749);
buf BUF1 (N1759, N1745);
or OR3 (N1760, N1740, N1380, N979);
nor NOR4 (N1761, N1757, N1496, N1284, N1377);
xor XOR2 (N1762, N1760, N511);
not NOT1 (N1763, N1761);
and AND3 (N1764, N1763, N1634, N862);
xor XOR2 (N1765, N1759, N681);
nor NOR2 (N1766, N1758, N1717);
xor XOR2 (N1767, N1755, N468);
nor NOR3 (N1768, N1762, N1665, N519);
buf BUF1 (N1769, N1756);
nand NAND3 (N1770, N1769, N1456, N503);
nand NAND3 (N1771, N1764, N633, N857);
xor XOR2 (N1772, N1766, N936);
xor XOR2 (N1773, N1736, N1652);
nand NAND3 (N1774, N1751, N938, N1649);
buf BUF1 (N1775, N1768);
nand NAND3 (N1776, N1774, N380, N935);
and AND4 (N1777, N1773, N1499, N1747, N933);
xor XOR2 (N1778, N1750, N321);
not NOT1 (N1779, N1772);
and AND4 (N1780, N1777, N1746, N1223, N1366);
or OR4 (N1781, N1778, N737, N1431, N1414);
xor XOR2 (N1782, N1770, N391);
not NOT1 (N1783, N1765);
or OR2 (N1784, N1781, N673);
and AND3 (N1785, N1783, N1587, N464);
xor XOR2 (N1786, N1785, N390);
nand NAND4 (N1787, N1775, N1265, N361, N566);
nand NAND3 (N1788, N1767, N299, N319);
nand NAND3 (N1789, N1788, N1745, N1439);
buf BUF1 (N1790, N1786);
not NOT1 (N1791, N1790);
buf BUF1 (N1792, N1752);
and AND4 (N1793, N1779, N1215, N1382, N916);
buf BUF1 (N1794, N1771);
not NOT1 (N1795, N1789);
or OR2 (N1796, N1795, N355);
xor XOR2 (N1797, N1776, N899);
and AND3 (N1798, N1793, N855, N1703);
nand NAND3 (N1799, N1782, N15, N207);
xor XOR2 (N1800, N1798, N1124);
or OR4 (N1801, N1794, N696, N750, N356);
or OR4 (N1802, N1791, N1413, N1649, N1737);
nand NAND4 (N1803, N1787, N923, N390, N590);
not NOT1 (N1804, N1796);
and AND2 (N1805, N1803, N1801);
or OR2 (N1806, N1395, N1584);
nor NOR3 (N1807, N1792, N1379, N1396);
buf BUF1 (N1808, N1802);
or OR2 (N1809, N1807, N289);
nor NOR3 (N1810, N1780, N1486, N890);
nor NOR4 (N1811, N1806, N449, N1582, N153);
or OR2 (N1812, N1811, N1602);
xor XOR2 (N1813, N1799, N1282);
xor XOR2 (N1814, N1813, N365);
or OR2 (N1815, N1804, N361);
not NOT1 (N1816, N1805);
nand NAND4 (N1817, N1812, N1342, N732, N1353);
nand NAND3 (N1818, N1797, N959, N1497);
nor NOR4 (N1819, N1800, N168, N920, N270);
or OR2 (N1820, N1818, N1743);
not NOT1 (N1821, N1815);
or OR4 (N1822, N1821, N1816, N824, N1779);
nor NOR2 (N1823, N1627, N52);
xor XOR2 (N1824, N1810, N1693);
and AND4 (N1825, N1814, N1539, N1005, N669);
buf BUF1 (N1826, N1824);
and AND2 (N1827, N1822, N557);
and AND3 (N1828, N1825, N1756, N83);
nor NOR4 (N1829, N1808, N836, N1745, N62);
or OR4 (N1830, N1817, N455, N1785, N208);
not NOT1 (N1831, N1826);
or OR4 (N1832, N1828, N25, N471, N1037);
or OR2 (N1833, N1819, N158);
or OR4 (N1834, N1829, N19, N791, N1796);
nor NOR4 (N1835, N1830, N507, N1159, N1639);
buf BUF1 (N1836, N1834);
and AND2 (N1837, N1820, N1242);
and AND2 (N1838, N1836, N689);
nor NOR2 (N1839, N1823, N923);
not NOT1 (N1840, N1827);
not NOT1 (N1841, N1839);
or OR3 (N1842, N1835, N1829, N1838);
and AND4 (N1843, N710, N681, N303, N1772);
and AND4 (N1844, N1784, N839, N482, N47);
or OR2 (N1845, N1843, N1316);
nor NOR2 (N1846, N1837, N493);
nor NOR3 (N1847, N1840, N1459, N223);
xor XOR2 (N1848, N1831, N1024);
nand NAND4 (N1849, N1833, N104, N1165, N879);
xor XOR2 (N1850, N1842, N760);
nand NAND4 (N1851, N1844, N370, N100, N564);
not NOT1 (N1852, N1850);
not NOT1 (N1853, N1852);
not NOT1 (N1854, N1845);
or OR2 (N1855, N1847, N393);
nor NOR4 (N1856, N1841, N810, N733, N1217);
xor XOR2 (N1857, N1849, N1406);
buf BUF1 (N1858, N1853);
buf BUF1 (N1859, N1832);
nor NOR4 (N1860, N1848, N1418, N115, N135);
xor XOR2 (N1861, N1856, N94);
not NOT1 (N1862, N1860);
buf BUF1 (N1863, N1859);
nor NOR4 (N1864, N1854, N516, N41, N490);
and AND4 (N1865, N1858, N940, N710, N1711);
nand NAND4 (N1866, N1865, N1724, N1007, N1783);
nand NAND4 (N1867, N1846, N606, N55, N1633);
not NOT1 (N1868, N1867);
xor XOR2 (N1869, N1863, N423);
buf BUF1 (N1870, N1861);
not NOT1 (N1871, N1809);
and AND3 (N1872, N1851, N173, N1076);
or OR3 (N1873, N1866, N759, N1458);
nor NOR2 (N1874, N1871, N1513);
nor NOR2 (N1875, N1864, N1228);
or OR4 (N1876, N1870, N1219, N834, N606);
and AND2 (N1877, N1862, N597);
or OR2 (N1878, N1855, N116);
nor NOR2 (N1879, N1873, N414);
nand NAND2 (N1880, N1857, N1607);
nand NAND3 (N1881, N1877, N87, N582);
buf BUF1 (N1882, N1878);
not NOT1 (N1883, N1879);
not NOT1 (N1884, N1868);
or OR2 (N1885, N1869, N1742);
and AND4 (N1886, N1884, N544, N791, N1226);
and AND2 (N1887, N1880, N1853);
or OR2 (N1888, N1874, N53);
not NOT1 (N1889, N1885);
xor XOR2 (N1890, N1881, N106);
xor XOR2 (N1891, N1876, N1379);
xor XOR2 (N1892, N1875, N599);
nand NAND3 (N1893, N1889, N801, N1640);
nor NOR2 (N1894, N1888, N1137);
xor XOR2 (N1895, N1890, N1243);
and AND3 (N1896, N1894, N80, N1142);
or OR2 (N1897, N1887, N177);
not NOT1 (N1898, N1897);
xor XOR2 (N1899, N1882, N1849);
nor NOR4 (N1900, N1883, N609, N1678, N1805);
nand NAND2 (N1901, N1899, N484);
nor NOR2 (N1902, N1898, N801);
nor NOR2 (N1903, N1901, N1695);
nand NAND4 (N1904, N1895, N590, N1597, N239);
and AND4 (N1905, N1903, N1233, N472, N1396);
not NOT1 (N1906, N1872);
and AND3 (N1907, N1891, N1143, N343);
not NOT1 (N1908, N1896);
xor XOR2 (N1909, N1886, N1828);
not NOT1 (N1910, N1904);
xor XOR2 (N1911, N1909, N298);
nand NAND2 (N1912, N1893, N1168);
buf BUF1 (N1913, N1908);
buf BUF1 (N1914, N1902);
and AND3 (N1915, N1892, N535, N396);
nand NAND4 (N1916, N1906, N17, N1668, N1824);
and AND4 (N1917, N1907, N1096, N1504, N557);
nand NAND4 (N1918, N1905, N1056, N1067, N1311);
buf BUF1 (N1919, N1910);
nand NAND2 (N1920, N1914, N1018);
not NOT1 (N1921, N1913);
buf BUF1 (N1922, N1921);
or OR4 (N1923, N1915, N1177, N504, N1482);
or OR4 (N1924, N1917, N1817, N582, N679);
and AND2 (N1925, N1916, N1845);
or OR4 (N1926, N1920, N1853, N108, N869);
xor XOR2 (N1927, N1918, N712);
nor NOR3 (N1928, N1911, N1793, N1558);
or OR4 (N1929, N1928, N234, N613, N1102);
not NOT1 (N1930, N1929);
nor NOR2 (N1931, N1919, N90);
xor XOR2 (N1932, N1922, N829);
or OR2 (N1933, N1925, N1140);
not NOT1 (N1934, N1933);
or OR2 (N1935, N1912, N1294);
nand NAND4 (N1936, N1900, N388, N881, N1245);
nor NOR3 (N1937, N1923, N1514, N452);
nor NOR2 (N1938, N1935, N1765);
buf BUF1 (N1939, N1926);
xor XOR2 (N1940, N1931, N1343);
buf BUF1 (N1941, N1939);
xor XOR2 (N1942, N1936, N1885);
nor NOR2 (N1943, N1937, N389);
and AND4 (N1944, N1940, N645, N1586, N1197);
nor NOR3 (N1945, N1924, N991, N753);
nor NOR3 (N1946, N1934, N386, N1148);
nor NOR2 (N1947, N1942, N1740);
not NOT1 (N1948, N1938);
buf BUF1 (N1949, N1946);
xor XOR2 (N1950, N1944, N1210);
xor XOR2 (N1951, N1927, N1169);
buf BUF1 (N1952, N1930);
nand NAND2 (N1953, N1943, N1109);
and AND3 (N1954, N1949, N108, N723);
not NOT1 (N1955, N1954);
not NOT1 (N1956, N1953);
or OR3 (N1957, N1950, N1761, N762);
nor NOR2 (N1958, N1951, N1308);
not NOT1 (N1959, N1945);
not NOT1 (N1960, N1932);
nand NAND4 (N1961, N1958, N1831, N1351, N1614);
nor NOR4 (N1962, N1957, N699, N991, N1009);
or OR3 (N1963, N1960, N107, N1221);
xor XOR2 (N1964, N1947, N1307);
xor XOR2 (N1965, N1955, N1617);
xor XOR2 (N1966, N1952, N339);
or OR4 (N1967, N1948, N1607, N1849, N1563);
buf BUF1 (N1968, N1962);
and AND3 (N1969, N1966, N829, N954);
xor XOR2 (N1970, N1963, N1948);
xor XOR2 (N1971, N1969, N625);
not NOT1 (N1972, N1970);
nor NOR4 (N1973, N1961, N1819, N252, N309);
buf BUF1 (N1974, N1973);
xor XOR2 (N1975, N1964, N1161);
xor XOR2 (N1976, N1974, N701);
not NOT1 (N1977, N1968);
and AND3 (N1978, N1975, N1397, N1570);
buf BUF1 (N1979, N1965);
not NOT1 (N1980, N1972);
or OR3 (N1981, N1941, N1954, N891);
not NOT1 (N1982, N1978);
and AND2 (N1983, N1980, N179);
nor NOR2 (N1984, N1979, N470);
xor XOR2 (N1985, N1967, N414);
and AND2 (N1986, N1985, N968);
and AND4 (N1987, N1983, N297, N1319, N535);
nor NOR3 (N1988, N1976, N200, N272);
or OR2 (N1989, N1982, N416);
or OR3 (N1990, N1986, N916, N508);
nand NAND3 (N1991, N1990, N424, N1375);
or OR4 (N1992, N1981, N1424, N1166, N1795);
nor NOR2 (N1993, N1977, N243);
xor XOR2 (N1994, N1984, N1302);
nor NOR2 (N1995, N1994, N1970);
and AND4 (N1996, N1956, N1840, N1247, N1919);
nor NOR4 (N1997, N1995, N170, N785, N1797);
buf BUF1 (N1998, N1959);
or OR3 (N1999, N1993, N429, N192);
xor XOR2 (N2000, N1971, N193);
not NOT1 (N2001, N1991);
buf BUF1 (N2002, N1989);
nand NAND4 (N2003, N1992, N1022, N1052, N1837);
not NOT1 (N2004, N2001);
xor XOR2 (N2005, N2002, N449);
buf BUF1 (N2006, N1988);
buf BUF1 (N2007, N2003);
and AND3 (N2008, N2007, N686, N1785);
xor XOR2 (N2009, N2005, N1126);
and AND4 (N2010, N1987, N28, N1189, N1129);
nor NOR3 (N2011, N2000, N1076, N128);
nor NOR2 (N2012, N2008, N56);
xor XOR2 (N2013, N1996, N626);
or OR2 (N2014, N1998, N1471);
nor NOR4 (N2015, N2011, N1810, N137, N241);
nand NAND4 (N2016, N2012, N649, N1090, N1871);
nor NOR4 (N2017, N1997, N83, N668, N187);
xor XOR2 (N2018, N2016, N296);
nor NOR2 (N2019, N2018, N1595);
or OR2 (N2020, N2004, N990);
nand NAND4 (N2021, N2013, N429, N772, N1085);
nor NOR2 (N2022, N2017, N1155);
and AND4 (N2023, N2022, N1919, N1911, N778);
nor NOR4 (N2024, N2019, N739, N444, N1923);
nor NOR3 (N2025, N2014, N1092, N177);
not NOT1 (N2026, N2010);
xor XOR2 (N2027, N2009, N1793);
xor XOR2 (N2028, N2023, N636);
or OR2 (N2029, N2025, N650);
or OR4 (N2030, N2028, N383, N1150, N1509);
not NOT1 (N2031, N2029);
or OR2 (N2032, N2021, N1612);
or OR3 (N2033, N2024, N2003, N556);
nand NAND4 (N2034, N2026, N1295, N1118, N1250);
buf BUF1 (N2035, N2032);
or OR4 (N2036, N2031, N1222, N35, N29);
nor NOR4 (N2037, N2027, N326, N1988, N1785);
xor XOR2 (N2038, N2015, N1887);
xor XOR2 (N2039, N2037, N1753);
and AND3 (N2040, N1999, N1442, N1952);
and AND3 (N2041, N2006, N1210, N1580);
nor NOR2 (N2042, N2035, N1725);
or OR2 (N2043, N2020, N1204);
xor XOR2 (N2044, N2030, N625);
and AND3 (N2045, N2042, N1233, N1798);
xor XOR2 (N2046, N2040, N1366);
nand NAND4 (N2047, N2044, N1183, N838, N317);
nand NAND2 (N2048, N2045, N1111);
and AND3 (N2049, N2047, N1569, N1738);
buf BUF1 (N2050, N2039);
or OR2 (N2051, N2046, N1930);
nor NOR4 (N2052, N2043, N358, N136, N473);
xor XOR2 (N2053, N2050, N401);
nand NAND2 (N2054, N2051, N570);
xor XOR2 (N2055, N2033, N1693);
buf BUF1 (N2056, N2049);
or OR3 (N2057, N2034, N1940, N348);
xor XOR2 (N2058, N2054, N911);
not NOT1 (N2059, N2048);
and AND2 (N2060, N2053, N194);
xor XOR2 (N2061, N2041, N179);
buf BUF1 (N2062, N2059);
not NOT1 (N2063, N2055);
nand NAND3 (N2064, N2058, N1380, N1916);
not NOT1 (N2065, N2052);
nand NAND4 (N2066, N2063, N140, N621, N1616);
or OR2 (N2067, N2065, N677);
nor NOR3 (N2068, N2038, N521, N1874);
not NOT1 (N2069, N2068);
nand NAND4 (N2070, N2057, N740, N1652, N717);
xor XOR2 (N2071, N2070, N65);
xor XOR2 (N2072, N2069, N1425);
buf BUF1 (N2073, N2062);
buf BUF1 (N2074, N2073);
not NOT1 (N2075, N2056);
nor NOR4 (N2076, N2071, N1654, N1764, N1010);
xor XOR2 (N2077, N2064, N1951);
not NOT1 (N2078, N2076);
or OR3 (N2079, N2060, N1484, N973);
and AND3 (N2080, N2079, N112, N788);
not NOT1 (N2081, N2066);
not NOT1 (N2082, N2072);
nand NAND3 (N2083, N2074, N1636, N1329);
xor XOR2 (N2084, N2067, N219);
xor XOR2 (N2085, N2082, N1463);
nor NOR3 (N2086, N2077, N2042, N799);
and AND4 (N2087, N2061, N648, N902, N1473);
nand NAND2 (N2088, N2087, N410);
nor NOR2 (N2089, N2078, N270);
and AND3 (N2090, N2075, N524, N1544);
buf BUF1 (N2091, N2089);
and AND4 (N2092, N2081, N738, N1426, N1955);
nor NOR4 (N2093, N2090, N160, N377, N2009);
nand NAND2 (N2094, N2093, N1773);
buf BUF1 (N2095, N2088);
or OR4 (N2096, N2036, N1106, N452, N363);
buf BUF1 (N2097, N2080);
nand NAND4 (N2098, N2094, N993, N496, N1173);
or OR3 (N2099, N2096, N1105, N37);
not NOT1 (N2100, N2085);
nand NAND3 (N2101, N2092, N1325, N1791);
not NOT1 (N2102, N2091);
nor NOR3 (N2103, N2097, N989, N345);
nor NOR3 (N2104, N2098, N1232, N289);
buf BUF1 (N2105, N2099);
nor NOR2 (N2106, N2095, N1347);
not NOT1 (N2107, N2102);
or OR2 (N2108, N2106, N471);
and AND4 (N2109, N2108, N1555, N1805, N2000);
or OR2 (N2110, N2105, N1599);
and AND3 (N2111, N2084, N326, N2060);
buf BUF1 (N2112, N2111);
not NOT1 (N2113, N2100);
buf BUF1 (N2114, N2110);
xor XOR2 (N2115, N2086, N755);
and AND4 (N2116, N2115, N724, N803, N1532);
nor NOR4 (N2117, N2104, N658, N1122, N919);
xor XOR2 (N2118, N2112, N1906);
not NOT1 (N2119, N2118);
buf BUF1 (N2120, N2117);
nor NOR3 (N2121, N2113, N1594, N1788);
xor XOR2 (N2122, N2120, N752);
not NOT1 (N2123, N2101);
buf BUF1 (N2124, N2103);
and AND3 (N2125, N2124, N927, N1602);
nand NAND2 (N2126, N2107, N1318);
or OR3 (N2127, N2083, N1529, N1369);
not NOT1 (N2128, N2125);
nor NOR2 (N2129, N2114, N374);
xor XOR2 (N2130, N2119, N2050);
buf BUF1 (N2131, N2123);
buf BUF1 (N2132, N2131);
nor NOR3 (N2133, N2122, N1450, N1418);
not NOT1 (N2134, N2128);
not NOT1 (N2135, N2126);
or OR3 (N2136, N2130, N210, N1920);
nor NOR2 (N2137, N2127, N658);
xor XOR2 (N2138, N2109, N1592);
and AND2 (N2139, N2136, N906);
nand NAND4 (N2140, N2134, N1660, N1819, N1876);
nor NOR2 (N2141, N2137, N634);
nor NOR3 (N2142, N2140, N693, N862);
and AND4 (N2143, N2141, N1300, N1686, N1421);
xor XOR2 (N2144, N2143, N450);
nand NAND4 (N2145, N2116, N2133, N1211, N906);
not NOT1 (N2146, N1811);
buf BUF1 (N2147, N2144);
or OR3 (N2148, N2135, N1549, N452);
nand NAND3 (N2149, N2138, N981, N2138);
nand NAND4 (N2150, N2148, N1613, N856, N1189);
or OR2 (N2151, N2146, N1836);
xor XOR2 (N2152, N2145, N1230);
or OR4 (N2153, N2139, N1846, N2062, N728);
nor NOR3 (N2154, N2129, N29, N1966);
and AND3 (N2155, N2151, N1632, N1301);
not NOT1 (N2156, N2121);
nand NAND3 (N2157, N2156, N1310, N1020);
xor XOR2 (N2158, N2154, N424);
nor NOR3 (N2159, N2158, N610, N203);
xor XOR2 (N2160, N2142, N1785);
buf BUF1 (N2161, N2155);
buf BUF1 (N2162, N2152);
and AND3 (N2163, N2162, N574, N419);
and AND2 (N2164, N2153, N1308);
buf BUF1 (N2165, N2161);
nor NOR2 (N2166, N2164, N2033);
nand NAND4 (N2167, N2157, N1199, N611, N347);
and AND3 (N2168, N2166, N551, N1175);
nor NOR4 (N2169, N2159, N1524, N401, N575);
and AND4 (N2170, N2165, N612, N624, N729);
buf BUF1 (N2171, N2150);
nand NAND2 (N2172, N2171, N567);
nand NAND2 (N2173, N2167, N641);
buf BUF1 (N2174, N2149);
or OR3 (N2175, N2132, N575, N1045);
xor XOR2 (N2176, N2172, N1076);
or OR4 (N2177, N2169, N1671, N1513, N241);
buf BUF1 (N2178, N2170);
not NOT1 (N2179, N2177);
nand NAND3 (N2180, N2160, N1547, N106);
nand NAND2 (N2181, N2180, N729);
not NOT1 (N2182, N2175);
not NOT1 (N2183, N2179);
or OR4 (N2184, N2176, N2136, N661, N1135);
not NOT1 (N2185, N2178);
nand NAND4 (N2186, N2181, N2130, N1877, N679);
not NOT1 (N2187, N2147);
and AND2 (N2188, N2163, N485);
or OR4 (N2189, N2168, N1610, N246, N1540);
buf BUF1 (N2190, N2187);
and AND2 (N2191, N2183, N1203);
xor XOR2 (N2192, N2188, N2030);
or OR2 (N2193, N2190, N1276);
buf BUF1 (N2194, N2192);
nand NAND4 (N2195, N2184, N330, N2005, N982);
not NOT1 (N2196, N2194);
or OR2 (N2197, N2185, N583);
nor NOR2 (N2198, N2195, N1442);
buf BUF1 (N2199, N2182);
or OR4 (N2200, N2198, N1927, N1205, N2104);
buf BUF1 (N2201, N2191);
not NOT1 (N2202, N2174);
xor XOR2 (N2203, N2201, N1417);
buf BUF1 (N2204, N2203);
nand NAND3 (N2205, N2173, N2038, N973);
xor XOR2 (N2206, N2186, N667);
buf BUF1 (N2207, N2206);
and AND3 (N2208, N2207, N1571, N2108);
nand NAND3 (N2209, N2205, N216, N333);
buf BUF1 (N2210, N2199);
nand NAND4 (N2211, N2209, N405, N291, N882);
xor XOR2 (N2212, N2193, N1391);
and AND3 (N2213, N2189, N2187, N954);
or OR2 (N2214, N2212, N162);
or OR4 (N2215, N2214, N371, N1799, N1378);
and AND4 (N2216, N2213, N428, N1494, N2210);
xor XOR2 (N2217, N1673, N2049);
or OR2 (N2218, N2216, N807);
buf BUF1 (N2219, N2197);
nor NOR3 (N2220, N2218, N1316, N600);
xor XOR2 (N2221, N2204, N759);
buf BUF1 (N2222, N2221);
not NOT1 (N2223, N2220);
nor NOR2 (N2224, N2200, N1535);
and AND3 (N2225, N2224, N2000, N1897);
xor XOR2 (N2226, N2215, N711);
not NOT1 (N2227, N2208);
nor NOR2 (N2228, N2223, N2212);
not NOT1 (N2229, N2226);
nor NOR2 (N2230, N2229, N2074);
xor XOR2 (N2231, N2222, N1674);
or OR3 (N2232, N2219, N1597, N1224);
or OR3 (N2233, N2217, N880, N2140);
not NOT1 (N2234, N2227);
nand NAND2 (N2235, N2234, N754);
or OR2 (N2236, N2228, N417);
or OR4 (N2237, N2233, N277, N1960, N684);
not NOT1 (N2238, N2237);
not NOT1 (N2239, N2225);
or OR2 (N2240, N2230, N764);
nand NAND4 (N2241, N2240, N224, N2159, N448);
or OR3 (N2242, N2236, N1064, N274);
or OR2 (N2243, N2241, N1533);
and AND3 (N2244, N2235, N212, N747);
and AND4 (N2245, N2202, N1160, N248, N2184);
buf BUF1 (N2246, N2211);
xor XOR2 (N2247, N2232, N694);
nand NAND4 (N2248, N2243, N500, N361, N599);
or OR3 (N2249, N2248, N2246, N1128);
xor XOR2 (N2250, N2129, N625);
nor NOR2 (N2251, N2245, N1084);
buf BUF1 (N2252, N2244);
nand NAND3 (N2253, N2238, N1770, N2200);
nor NOR4 (N2254, N2252, N856, N1500, N322);
nand NAND2 (N2255, N2247, N1680);
nand NAND2 (N2256, N2242, N1217);
buf BUF1 (N2257, N2253);
xor XOR2 (N2258, N2255, N1531);
xor XOR2 (N2259, N2231, N811);
or OR2 (N2260, N2250, N286);
nand NAND3 (N2261, N2259, N485, N358);
or OR3 (N2262, N2254, N1653, N432);
nand NAND4 (N2263, N2251, N302, N897, N208);
or OR2 (N2264, N2260, N1866);
buf BUF1 (N2265, N2239);
not NOT1 (N2266, N2265);
nand NAND3 (N2267, N2249, N401, N356);
buf BUF1 (N2268, N2262);
xor XOR2 (N2269, N2264, N46);
not NOT1 (N2270, N2256);
buf BUF1 (N2271, N2196);
nand NAND3 (N2272, N2268, N1413, N378);
buf BUF1 (N2273, N2258);
nor NOR4 (N2274, N2263, N2041, N1469, N1129);
or OR4 (N2275, N2269, N245, N1732, N1199);
and AND3 (N2276, N2267, N199, N1460);
not NOT1 (N2277, N2272);
buf BUF1 (N2278, N2261);
xor XOR2 (N2279, N2276, N751);
or OR2 (N2280, N2275, N1566);
nand NAND4 (N2281, N2271, N756, N2017, N330);
nand NAND4 (N2282, N2270, N1994, N276, N348);
xor XOR2 (N2283, N2278, N1764);
nand NAND2 (N2284, N2279, N2206);
not NOT1 (N2285, N2282);
xor XOR2 (N2286, N2280, N2076);
not NOT1 (N2287, N2286);
not NOT1 (N2288, N2273);
nor NOR3 (N2289, N2285, N2122, N2048);
not NOT1 (N2290, N2274);
or OR2 (N2291, N2283, N732);
not NOT1 (N2292, N2277);
xor XOR2 (N2293, N2288, N909);
and AND2 (N2294, N2266, N888);
nor NOR2 (N2295, N2294, N479);
buf BUF1 (N2296, N2291);
buf BUF1 (N2297, N2295);
not NOT1 (N2298, N2287);
nor NOR3 (N2299, N2292, N589, N1458);
xor XOR2 (N2300, N2296, N1933);
xor XOR2 (N2301, N2284, N2188);
xor XOR2 (N2302, N2297, N1749);
and AND3 (N2303, N2289, N1971, N852);
not NOT1 (N2304, N2301);
xor XOR2 (N2305, N2290, N1562);
nand NAND3 (N2306, N2299, N61, N1961);
nand NAND2 (N2307, N2303, N1793);
or OR4 (N2308, N2298, N1309, N1182, N2116);
and AND4 (N2309, N2281, N2026, N606, N1461);
buf BUF1 (N2310, N2306);
xor XOR2 (N2311, N2304, N387);
xor XOR2 (N2312, N2300, N1735);
nor NOR4 (N2313, N2307, N1032, N1257, N1372);
or OR4 (N2314, N2310, N1772, N1515, N691);
buf BUF1 (N2315, N2312);
nand NAND2 (N2316, N2314, N1414);
nand NAND4 (N2317, N2311, N1107, N835, N1892);
and AND3 (N2318, N2305, N506, N782);
and AND2 (N2319, N2316, N1507);
not NOT1 (N2320, N2319);
nand NAND4 (N2321, N2315, N1222, N153, N2130);
nor NOR2 (N2322, N2320, N1744);
nor NOR4 (N2323, N2317, N1063, N1236, N1170);
or OR4 (N2324, N2321, N370, N937, N1034);
or OR4 (N2325, N2322, N788, N438, N578);
nor NOR4 (N2326, N2308, N1985, N883, N1877);
buf BUF1 (N2327, N2325);
nor NOR3 (N2328, N2257, N112, N484);
nor NOR4 (N2329, N2326, N1475, N2326, N1134);
nor NOR2 (N2330, N2293, N933);
or OR2 (N2331, N2309, N98);
not NOT1 (N2332, N2324);
or OR2 (N2333, N2318, N2161);
xor XOR2 (N2334, N2327, N889);
and AND2 (N2335, N2329, N1069);
buf BUF1 (N2336, N2328);
and AND3 (N2337, N2332, N1806, N694);
not NOT1 (N2338, N2336);
or OR4 (N2339, N2335, N85, N2153, N2005);
xor XOR2 (N2340, N2333, N1786);
xor XOR2 (N2341, N2313, N166);
buf BUF1 (N2342, N2334);
and AND3 (N2343, N2340, N1525, N1416);
xor XOR2 (N2344, N2339, N956);
buf BUF1 (N2345, N2330);
not NOT1 (N2346, N2338);
not NOT1 (N2347, N2337);
nor NOR2 (N2348, N2342, N2241);
not NOT1 (N2349, N2331);
or OR2 (N2350, N2323, N1980);
nor NOR2 (N2351, N2345, N1872);
and AND4 (N2352, N2350, N1426, N1223, N776);
xor XOR2 (N2353, N2347, N1281);
nor NOR3 (N2354, N2349, N1927, N2079);
buf BUF1 (N2355, N2346);
or OR3 (N2356, N2302, N2223, N1013);
or OR4 (N2357, N2341, N1278, N810, N1775);
nor NOR4 (N2358, N2356, N1065, N626, N2036);
and AND2 (N2359, N2343, N1093);
not NOT1 (N2360, N2354);
nand NAND2 (N2361, N2344, N2306);
buf BUF1 (N2362, N2353);
nand NAND4 (N2363, N2358, N2092, N370, N1664);
and AND4 (N2364, N2361, N1388, N481, N2033);
or OR2 (N2365, N2357, N549);
and AND3 (N2366, N2348, N2092, N879);
or OR4 (N2367, N2366, N1599, N917, N263);
and AND2 (N2368, N2360, N489);
nand NAND4 (N2369, N2352, N982, N1407, N770);
nor NOR4 (N2370, N2362, N350, N441, N665);
xor XOR2 (N2371, N2370, N846);
and AND3 (N2372, N2369, N22, N1256);
or OR2 (N2373, N2363, N1650);
buf BUF1 (N2374, N2359);
buf BUF1 (N2375, N2364);
or OR3 (N2376, N2373, N833, N2088);
xor XOR2 (N2377, N2374, N2038);
or OR4 (N2378, N2372, N1067, N2096, N1836);
nand NAND4 (N2379, N2351, N683, N1099, N1476);
xor XOR2 (N2380, N2376, N727);
buf BUF1 (N2381, N2365);
and AND3 (N2382, N2378, N2101, N563);
xor XOR2 (N2383, N2377, N1755);
and AND2 (N2384, N2382, N211);
and AND2 (N2385, N2384, N1305);
nor NOR3 (N2386, N2355, N2053, N1664);
nor NOR2 (N2387, N2381, N2253);
xor XOR2 (N2388, N2371, N1110);
nor NOR2 (N2389, N2380, N36);
and AND4 (N2390, N2383, N903, N152, N2387);
buf BUF1 (N2391, N1279);
xor XOR2 (N2392, N2391, N167);
and AND2 (N2393, N2367, N1691);
nor NOR2 (N2394, N2390, N220);
nor NOR3 (N2395, N2386, N1370, N2296);
xor XOR2 (N2396, N2385, N2075);
or OR3 (N2397, N2389, N485, N702);
not NOT1 (N2398, N2375);
or OR4 (N2399, N2379, N207, N12, N2194);
nand NAND4 (N2400, N2395, N699, N957, N393);
or OR2 (N2401, N2399, N958);
nor NOR2 (N2402, N2396, N282);
buf BUF1 (N2403, N2402);
not NOT1 (N2404, N2368);
nand NAND4 (N2405, N2403, N985, N1346, N2316);
nor NOR2 (N2406, N2392, N326);
buf BUF1 (N2407, N2400);
xor XOR2 (N2408, N2393, N337);
nand NAND4 (N2409, N2388, N50, N2256, N1588);
nor NOR4 (N2410, N2404, N2229, N522, N2327);
or OR3 (N2411, N2398, N2355, N1979);
not NOT1 (N2412, N2397);
not NOT1 (N2413, N2394);
not NOT1 (N2414, N2409);
and AND2 (N2415, N2401, N1627);
buf BUF1 (N2416, N2413);
buf BUF1 (N2417, N2407);
and AND2 (N2418, N2410, N193);
nand NAND4 (N2419, N2416, N2358, N1152, N231);
nor NOR2 (N2420, N2414, N1675);
and AND4 (N2421, N2412, N1102, N487, N931);
nand NAND3 (N2422, N2417, N2266, N1847);
xor XOR2 (N2423, N2418, N1785);
nor NOR4 (N2424, N2415, N1289, N1712, N1553);
nor NOR4 (N2425, N2424, N1979, N493, N784);
xor XOR2 (N2426, N2425, N81);
and AND4 (N2427, N2421, N1501, N2224, N153);
buf BUF1 (N2428, N2419);
or OR4 (N2429, N2405, N2327, N1183, N402);
and AND4 (N2430, N2422, N1238, N444, N174);
nand NAND2 (N2431, N2408, N1090);
buf BUF1 (N2432, N2428);
or OR2 (N2433, N2423, N2187);
not NOT1 (N2434, N2420);
not NOT1 (N2435, N2429);
not NOT1 (N2436, N2435);
nor NOR4 (N2437, N2436, N2182, N236, N1028);
nand NAND2 (N2438, N2432, N1548);
not NOT1 (N2439, N2438);
buf BUF1 (N2440, N2434);
nand NAND2 (N2441, N2406, N545);
and AND4 (N2442, N2427, N2110, N823, N471);
buf BUF1 (N2443, N2440);
nand NAND3 (N2444, N2411, N1838, N1891);
buf BUF1 (N2445, N2430);
and AND4 (N2446, N2426, N125, N231, N1636);
nand NAND2 (N2447, N2442, N1398);
nor NOR3 (N2448, N2446, N2271, N193);
nand NAND3 (N2449, N2433, N2407, N267);
xor XOR2 (N2450, N2449, N49);
xor XOR2 (N2451, N2448, N2217);
nand NAND4 (N2452, N2444, N1934, N473, N1181);
xor XOR2 (N2453, N2452, N433);
and AND3 (N2454, N2441, N1159, N301);
xor XOR2 (N2455, N2451, N1170);
buf BUF1 (N2456, N2443);
or OR3 (N2457, N2454, N744, N655);
xor XOR2 (N2458, N2453, N992);
buf BUF1 (N2459, N2458);
not NOT1 (N2460, N2457);
not NOT1 (N2461, N2460);
or OR4 (N2462, N2455, N1192, N2098, N1933);
xor XOR2 (N2463, N2447, N1476);
buf BUF1 (N2464, N2445);
buf BUF1 (N2465, N2456);
and AND3 (N2466, N2439, N128, N48);
nor NOR3 (N2467, N2466, N726, N340);
nand NAND3 (N2468, N2462, N1336, N825);
and AND3 (N2469, N2465, N1953, N376);
xor XOR2 (N2470, N2467, N553);
or OR4 (N2471, N2464, N845, N1720, N2180);
and AND3 (N2472, N2471, N1357, N1840);
nor NOR4 (N2473, N2461, N2436, N904, N2259);
buf BUF1 (N2474, N2469);
nor NOR2 (N2475, N2431, N1914);
nor NOR3 (N2476, N2437, N1181, N1370);
nand NAND3 (N2477, N2468, N400, N2003);
or OR2 (N2478, N2474, N1638);
xor XOR2 (N2479, N2473, N1764);
buf BUF1 (N2480, N2478);
nand NAND3 (N2481, N2477, N827, N2463);
xor XOR2 (N2482, N2352, N737);
nor NOR2 (N2483, N2472, N2046);
nor NOR2 (N2484, N2475, N2114);
xor XOR2 (N2485, N2459, N1545);
buf BUF1 (N2486, N2484);
or OR3 (N2487, N2450, N2355, N1397);
or OR2 (N2488, N2480, N1218);
xor XOR2 (N2489, N2487, N547);
buf BUF1 (N2490, N2483);
or OR4 (N2491, N2481, N1221, N19, N50);
nand NAND2 (N2492, N2489, N1994);
xor XOR2 (N2493, N2479, N2274);
nand NAND2 (N2494, N2482, N1790);
xor XOR2 (N2495, N2490, N1582);
nand NAND2 (N2496, N2476, N1774);
and AND2 (N2497, N2470, N2100);
not NOT1 (N2498, N2491);
nor NOR3 (N2499, N2495, N1848, N281);
xor XOR2 (N2500, N2496, N849);
and AND4 (N2501, N2498, N1026, N1115, N2478);
and AND2 (N2502, N2493, N1447);
or OR2 (N2503, N2500, N1999);
buf BUF1 (N2504, N2501);
not NOT1 (N2505, N2494);
not NOT1 (N2506, N2503);
and AND4 (N2507, N2497, N2229, N1766, N1382);
nand NAND3 (N2508, N2502, N1140, N2357);
xor XOR2 (N2509, N2485, N1969);
nor NOR4 (N2510, N2499, N2334, N1865, N2294);
or OR4 (N2511, N2488, N1958, N1140, N1094);
nand NAND4 (N2512, N2492, N17, N2478, N153);
nor NOR3 (N2513, N2506, N2131, N1220);
xor XOR2 (N2514, N2504, N737);
nor NOR2 (N2515, N2509, N219);
or OR3 (N2516, N2515, N612, N339);
xor XOR2 (N2517, N2505, N700);
nor NOR3 (N2518, N2510, N875, N356);
xor XOR2 (N2519, N2514, N629);
or OR3 (N2520, N2508, N1275, N552);
or OR2 (N2521, N2486, N2352);
buf BUF1 (N2522, N2521);
nor NOR2 (N2523, N2518, N729);
nand NAND4 (N2524, N2522, N232, N1266, N184);
not NOT1 (N2525, N2512);
not NOT1 (N2526, N2524);
buf BUF1 (N2527, N2525);
buf BUF1 (N2528, N2520);
nor NOR3 (N2529, N2527, N700, N1527);
xor XOR2 (N2530, N2513, N2526);
nand NAND4 (N2531, N422, N26, N1446, N1113);
and AND4 (N2532, N2523, N1620, N1561, N1110);
xor XOR2 (N2533, N2532, N876);
not NOT1 (N2534, N2517);
and AND2 (N2535, N2534, N1251);
nor NOR2 (N2536, N2530, N2039);
nand NAND4 (N2537, N2511, N379, N166, N544);
not NOT1 (N2538, N2535);
and AND4 (N2539, N2529, N1726, N2155, N1204);
xor XOR2 (N2540, N2538, N2406);
nor NOR3 (N2541, N2516, N168, N303);
xor XOR2 (N2542, N2507, N1228);
xor XOR2 (N2543, N2536, N1782);
nor NOR4 (N2544, N2540, N2181, N2373, N2024);
nand NAND3 (N2545, N2519, N1853, N1050);
and AND2 (N2546, N2543, N2267);
xor XOR2 (N2547, N2546, N242);
nor NOR2 (N2548, N2544, N609);
nor NOR3 (N2549, N2528, N655, N288);
and AND3 (N2550, N2531, N797, N71);
buf BUF1 (N2551, N2545);
nand NAND3 (N2552, N2539, N2266, N211);
not NOT1 (N2553, N2547);
xor XOR2 (N2554, N2537, N1824);
and AND4 (N2555, N2533, N1041, N974, N1247);
xor XOR2 (N2556, N2549, N2168);
and AND2 (N2557, N2555, N2232);
xor XOR2 (N2558, N2548, N1157);
or OR3 (N2559, N2552, N2004, N1138);
nor NOR3 (N2560, N2542, N942, N1819);
not NOT1 (N2561, N2558);
nor NOR2 (N2562, N2541, N2190);
nand NAND3 (N2563, N2553, N2, N1633);
not NOT1 (N2564, N2551);
nand NAND4 (N2565, N2562, N797, N1185, N2133);
or OR3 (N2566, N2559, N2243, N2360);
or OR3 (N2567, N2557, N1430, N421);
nand NAND3 (N2568, N2556, N1371, N203);
not NOT1 (N2569, N2568);
nand NAND3 (N2570, N2566, N2428, N1264);
nand NAND2 (N2571, N2567, N1181);
xor XOR2 (N2572, N2563, N195);
and AND4 (N2573, N2572, N237, N333, N2206);
nand NAND3 (N2574, N2561, N2139, N1012);
xor XOR2 (N2575, N2564, N2522);
or OR4 (N2576, N2550, N1528, N677, N491);
buf BUF1 (N2577, N2571);
xor XOR2 (N2578, N2575, N2033);
and AND2 (N2579, N2577, N649);
not NOT1 (N2580, N2560);
buf BUF1 (N2581, N2565);
nor NOR4 (N2582, N2579, N2562, N2103, N614);
or OR3 (N2583, N2554, N1952, N1352);
buf BUF1 (N2584, N2582);
nor NOR2 (N2585, N2569, N2415);
and AND3 (N2586, N2574, N2417, N1391);
and AND3 (N2587, N2570, N107, N755);
and AND3 (N2588, N2573, N759, N1828);
nor NOR4 (N2589, N2586, N1654, N1119, N1593);
xor XOR2 (N2590, N2587, N2204);
and AND4 (N2591, N2585, N1188, N1508, N1315);
and AND2 (N2592, N2578, N89);
buf BUF1 (N2593, N2584);
xor XOR2 (N2594, N2590, N2013);
nor NOR3 (N2595, N2592, N2384, N2201);
and AND2 (N2596, N2580, N2018);
not NOT1 (N2597, N2594);
and AND3 (N2598, N2581, N1491, N352);
buf BUF1 (N2599, N2597);
nor NOR2 (N2600, N2591, N1021);
not NOT1 (N2601, N2599);
or OR3 (N2602, N2596, N2507, N493);
nor NOR2 (N2603, N2600, N2531);
nand NAND4 (N2604, N2595, N97, N2118, N2051);
xor XOR2 (N2605, N2598, N2092);
nand NAND3 (N2606, N2604, N1509, N101);
not NOT1 (N2607, N2576);
nand NAND3 (N2608, N2593, N67, N1839);
and AND2 (N2609, N2588, N955);
nor NOR2 (N2610, N2603, N609);
buf BUF1 (N2611, N2589);
not NOT1 (N2612, N2583);
or OR3 (N2613, N2602, N1639, N1960);
or OR3 (N2614, N2613, N205, N2311);
buf BUF1 (N2615, N2611);
nor NOR4 (N2616, N2614, N1451, N285, N1809);
nor NOR2 (N2617, N2601, N2436);
buf BUF1 (N2618, N2605);
buf BUF1 (N2619, N2618);
buf BUF1 (N2620, N2609);
buf BUF1 (N2621, N2617);
buf BUF1 (N2622, N2612);
buf BUF1 (N2623, N2621);
and AND4 (N2624, N2616, N1627, N709, N501);
buf BUF1 (N2625, N2606);
and AND2 (N2626, N2624, N2450);
and AND2 (N2627, N2620, N987);
nor NOR4 (N2628, N2615, N2563, N670, N424);
nor NOR2 (N2629, N2627, N1154);
nand NAND4 (N2630, N2625, N1596, N465, N2543);
buf BUF1 (N2631, N2610);
nor NOR2 (N2632, N2628, N2629);
or OR2 (N2633, N612, N2220);
nand NAND4 (N2634, N2630, N205, N783, N765);
buf BUF1 (N2635, N2619);
not NOT1 (N2636, N2622);
or OR2 (N2637, N2636, N799);
nand NAND4 (N2638, N2634, N51, N1492, N748);
or OR4 (N2639, N2631, N64, N1803, N1184);
or OR2 (N2640, N2632, N947);
and AND4 (N2641, N2607, N1797, N562, N499);
buf BUF1 (N2642, N2640);
nor NOR2 (N2643, N2642, N1427);
nor NOR4 (N2644, N2643, N341, N1002, N1856);
buf BUF1 (N2645, N2635);
and AND2 (N2646, N2644, N1935);
nor NOR3 (N2647, N2639, N941, N2170);
buf BUF1 (N2648, N2608);
nand NAND4 (N2649, N2623, N2032, N1, N296);
not NOT1 (N2650, N2638);
nor NOR3 (N2651, N2646, N1583, N1438);
buf BUF1 (N2652, N2641);
nor NOR4 (N2653, N2637, N1138, N779, N1932);
xor XOR2 (N2654, N2650, N702);
buf BUF1 (N2655, N2654);
and AND2 (N2656, N2649, N1689);
xor XOR2 (N2657, N2653, N600);
xor XOR2 (N2658, N2647, N315);
nor NOR3 (N2659, N2651, N1108, N926);
not NOT1 (N2660, N2657);
or OR4 (N2661, N2659, N818, N1575, N311);
xor XOR2 (N2662, N2660, N611);
nor NOR4 (N2663, N2626, N757, N1664, N484);
xor XOR2 (N2664, N2652, N1520);
nand NAND3 (N2665, N2645, N552, N589);
nor NOR4 (N2666, N2633, N2526, N1497, N1355);
not NOT1 (N2667, N2661);
and AND4 (N2668, N2663, N2572, N932, N1939);
or OR4 (N2669, N2648, N1108, N877, N89);
and AND4 (N2670, N2664, N2342, N1326, N994);
nor NOR2 (N2671, N2662, N1451);
xor XOR2 (N2672, N2658, N1174);
nor NOR3 (N2673, N2655, N1702, N875);
and AND2 (N2674, N2670, N2131);
nand NAND2 (N2675, N2673, N2300);
nor NOR3 (N2676, N2667, N1247, N1899);
nand NAND2 (N2677, N2656, N64);
xor XOR2 (N2678, N2676, N1204);
xor XOR2 (N2679, N2678, N2441);
and AND4 (N2680, N2668, N1392, N2640, N1804);
and AND2 (N2681, N2665, N1682);
nand NAND4 (N2682, N2681, N858, N904, N2562);
nor NOR4 (N2683, N2671, N1542, N2339, N1950);
or OR3 (N2684, N2674, N2395, N180);
not NOT1 (N2685, N2684);
or OR3 (N2686, N2679, N2142, N2244);
not NOT1 (N2687, N2675);
not NOT1 (N2688, N2682);
xor XOR2 (N2689, N2669, N1967);
nand NAND3 (N2690, N2677, N1407, N1954);
nand NAND2 (N2691, N2688, N760);
nor NOR4 (N2692, N2691, N1437, N489, N824);
or OR4 (N2693, N2683, N352, N2550, N2182);
or OR2 (N2694, N2680, N506);
nand NAND2 (N2695, N2685, N1794);
not NOT1 (N2696, N2689);
nor NOR2 (N2697, N2672, N2246);
xor XOR2 (N2698, N2690, N1588);
xor XOR2 (N2699, N2696, N2170);
nand NAND4 (N2700, N2693, N880, N2568, N1550);
nor NOR2 (N2701, N2700, N599);
buf BUF1 (N2702, N2692);
and AND3 (N2703, N2697, N1266, N2456);
buf BUF1 (N2704, N2687);
or OR3 (N2705, N2698, N1295, N1515);
or OR4 (N2706, N2702, N1609, N2109, N1277);
nand NAND4 (N2707, N2695, N2451, N2594, N688);
xor XOR2 (N2708, N2694, N701);
nor NOR2 (N2709, N2705, N2384);
xor XOR2 (N2710, N2706, N2618);
buf BUF1 (N2711, N2666);
buf BUF1 (N2712, N2704);
buf BUF1 (N2713, N2712);
and AND3 (N2714, N2699, N2033, N410);
not NOT1 (N2715, N2709);
xor XOR2 (N2716, N2703, N2412);
or OR4 (N2717, N2716, N424, N1370, N133);
and AND2 (N2718, N2711, N182);
and AND2 (N2719, N2717, N389);
nand NAND2 (N2720, N2710, N496);
buf BUF1 (N2721, N2714);
nor NOR2 (N2722, N2701, N1954);
not NOT1 (N2723, N2708);
and AND2 (N2724, N2713, N1768);
and AND4 (N2725, N2686, N356, N243, N19);
buf BUF1 (N2726, N2718);
nand NAND3 (N2727, N2726, N1024, N2469);
buf BUF1 (N2728, N2720);
not NOT1 (N2729, N2715);
not NOT1 (N2730, N2728);
and AND3 (N2731, N2719, N2464, N1680);
or OR2 (N2732, N2729, N2051);
nand NAND3 (N2733, N2724, N2145, N1887);
nor NOR2 (N2734, N2731, N1687);
nand NAND3 (N2735, N2725, N2493, N458);
nor NOR4 (N2736, N2732, N38, N229, N2266);
and AND3 (N2737, N2736, N91, N1646);
nand NAND2 (N2738, N2730, N2570);
buf BUF1 (N2739, N2707);
nand NAND4 (N2740, N2727, N549, N2165, N2007);
buf BUF1 (N2741, N2734);
and AND3 (N2742, N2721, N1289, N2596);
buf BUF1 (N2743, N2742);
buf BUF1 (N2744, N2740);
not NOT1 (N2745, N2739);
nand NAND2 (N2746, N2745, N2212);
xor XOR2 (N2747, N2744, N1013);
not NOT1 (N2748, N2722);
buf BUF1 (N2749, N2738);
buf BUF1 (N2750, N2741);
nor NOR4 (N2751, N2733, N1830, N724, N993);
not NOT1 (N2752, N2747);
nor NOR4 (N2753, N2723, N1748, N857, N1087);
nand NAND4 (N2754, N2735, N1721, N1909, N704);
buf BUF1 (N2755, N2748);
buf BUF1 (N2756, N2750);
xor XOR2 (N2757, N2751, N2636);
buf BUF1 (N2758, N2754);
xor XOR2 (N2759, N2758, N1311);
and AND3 (N2760, N2755, N779, N2197);
and AND4 (N2761, N2752, N2745, N301, N246);
nand NAND3 (N2762, N2743, N429, N1808);
xor XOR2 (N2763, N2762, N297);
nor NOR4 (N2764, N2753, N1584, N2259, N52);
buf BUF1 (N2765, N2763);
xor XOR2 (N2766, N2737, N1361);
nand NAND3 (N2767, N2761, N2061, N651);
xor XOR2 (N2768, N2746, N313);
buf BUF1 (N2769, N2765);
nand NAND3 (N2770, N2767, N2223, N2575);
or OR3 (N2771, N2766, N187, N2091);
and AND3 (N2772, N2768, N1860, N1212);
buf BUF1 (N2773, N2759);
xor XOR2 (N2774, N2757, N2420);
not NOT1 (N2775, N2772);
buf BUF1 (N2776, N2770);
nor NOR4 (N2777, N2773, N662, N1677, N2750);
buf BUF1 (N2778, N2777);
nor NOR3 (N2779, N2769, N512, N2144);
nand NAND4 (N2780, N2779, N2139, N24, N1597);
or OR3 (N2781, N2774, N738, N1991);
or OR3 (N2782, N2776, N1778, N2355);
and AND2 (N2783, N2749, N971);
and AND3 (N2784, N2764, N2047, N634);
or OR4 (N2785, N2756, N584, N1738, N2377);
or OR4 (N2786, N2782, N620, N337, N1799);
not NOT1 (N2787, N2783);
buf BUF1 (N2788, N2775);
buf BUF1 (N2789, N2786);
nor NOR3 (N2790, N2788, N1156, N1618);
and AND2 (N2791, N2785, N27);
buf BUF1 (N2792, N2790);
xor XOR2 (N2793, N2781, N1723);
and AND4 (N2794, N2784, N1176, N836, N2192);
not NOT1 (N2795, N2771);
nand NAND4 (N2796, N2787, N252, N733, N1843);
or OR4 (N2797, N2789, N688, N2535, N2445);
nor NOR3 (N2798, N2794, N2062, N2193);
or OR4 (N2799, N2796, N325, N936, N1107);
or OR2 (N2800, N2780, N2363);
nor NOR4 (N2801, N2793, N230, N1289, N2270);
nor NOR3 (N2802, N2800, N2534, N1115);
or OR3 (N2803, N2798, N1776, N1925);
nor NOR4 (N2804, N2801, N974, N549, N2005);
not NOT1 (N2805, N2795);
nor NOR3 (N2806, N2799, N2516, N1775);
buf BUF1 (N2807, N2797);
not NOT1 (N2808, N2807);
nand NAND2 (N2809, N2778, N2229);
not NOT1 (N2810, N2760);
buf BUF1 (N2811, N2808);
not NOT1 (N2812, N2809);
not NOT1 (N2813, N2792);
or OR3 (N2814, N2805, N1827, N2151);
nor NOR3 (N2815, N2802, N2524, N446);
and AND2 (N2816, N2803, N2077);
nand NAND2 (N2817, N2811, N529);
nor NOR2 (N2818, N2813, N2364);
nor NOR2 (N2819, N2804, N1066);
nand NAND4 (N2820, N2817, N1722, N347, N239);
nor NOR3 (N2821, N2812, N1057, N1530);
or OR3 (N2822, N2806, N1985, N1512);
xor XOR2 (N2823, N2816, N81);
nand NAND3 (N2824, N2821, N2065, N566);
nand NAND4 (N2825, N2810, N76, N510, N290);
buf BUF1 (N2826, N2814);
nor NOR3 (N2827, N2826, N498, N2351);
nor NOR3 (N2828, N2825, N1960, N2652);
or OR2 (N2829, N2820, N1757);
nor NOR2 (N2830, N2828, N437);
or OR2 (N2831, N2815, N2610);
not NOT1 (N2832, N2819);
and AND2 (N2833, N2831, N2672);
and AND4 (N2834, N2830, N2181, N1366, N2579);
not NOT1 (N2835, N2832);
and AND4 (N2836, N2833, N2773, N2525, N1991);
and AND2 (N2837, N2823, N1089);
nor NOR3 (N2838, N2824, N1192, N1726);
not NOT1 (N2839, N2834);
buf BUF1 (N2840, N2791);
or OR2 (N2841, N2836, N2297);
nand NAND3 (N2842, N2827, N1253, N982);
or OR2 (N2843, N2818, N1375);
nand NAND4 (N2844, N2839, N2654, N2721, N1227);
nand NAND4 (N2845, N2840, N289, N2733, N34);
xor XOR2 (N2846, N2845, N2695);
or OR3 (N2847, N2837, N1732, N1322);
nor NOR2 (N2848, N2835, N1629);
or OR3 (N2849, N2838, N1314, N460);
not NOT1 (N2850, N2842);
nand NAND3 (N2851, N2844, N1810, N342);
not NOT1 (N2852, N2829);
not NOT1 (N2853, N2846);
nand NAND2 (N2854, N2853, N2768);
nor NOR3 (N2855, N2848, N2775, N1497);
not NOT1 (N2856, N2822);
not NOT1 (N2857, N2856);
or OR4 (N2858, N2849, N540, N705, N907);
or OR2 (N2859, N2850, N1049);
nand NAND2 (N2860, N2852, N2716);
and AND3 (N2861, N2854, N692, N254);
nor NOR4 (N2862, N2847, N1635, N539, N1055);
buf BUF1 (N2863, N2862);
nor NOR3 (N2864, N2858, N1313, N929);
or OR2 (N2865, N2841, N778);
not NOT1 (N2866, N2863);
nand NAND4 (N2867, N2855, N902, N356, N442);
nand NAND3 (N2868, N2851, N1289, N1260);
and AND3 (N2869, N2843, N796, N1733);
buf BUF1 (N2870, N2859);
nand NAND4 (N2871, N2870, N928, N1845, N948);
xor XOR2 (N2872, N2871, N2569);
and AND3 (N2873, N2864, N551, N867);
nand NAND4 (N2874, N2867, N157, N165, N2770);
nor NOR3 (N2875, N2872, N1624, N2535);
or OR4 (N2876, N2874, N1763, N87, N2713);
or OR3 (N2877, N2861, N2642, N1607);
xor XOR2 (N2878, N2877, N147);
buf BUF1 (N2879, N2869);
not NOT1 (N2880, N2873);
or OR2 (N2881, N2865, N496);
and AND2 (N2882, N2868, N767);
or OR3 (N2883, N2857, N609, N65);
not NOT1 (N2884, N2866);
and AND3 (N2885, N2876, N645, N654);
not NOT1 (N2886, N2885);
nand NAND2 (N2887, N2881, N1957);
not NOT1 (N2888, N2882);
xor XOR2 (N2889, N2875, N2364);
or OR3 (N2890, N2879, N2212, N1751);
or OR3 (N2891, N2878, N1004, N2433);
and AND3 (N2892, N2883, N605, N1270);
buf BUF1 (N2893, N2888);
and AND2 (N2894, N2891, N854);
and AND3 (N2895, N2889, N1469, N2711);
nor NOR3 (N2896, N2892, N2086, N232);
nor NOR4 (N2897, N2884, N2092, N1641, N1587);
xor XOR2 (N2898, N2887, N1276);
and AND4 (N2899, N2893, N2349, N1100, N2717);
and AND3 (N2900, N2899, N917, N2372);
nand NAND3 (N2901, N2860, N776, N738);
and AND2 (N2902, N2886, N350);
buf BUF1 (N2903, N2897);
or OR3 (N2904, N2895, N2036, N2362);
or OR3 (N2905, N2898, N1122, N484);
xor XOR2 (N2906, N2903, N351);
buf BUF1 (N2907, N2894);
nor NOR3 (N2908, N2880, N852, N931);
xor XOR2 (N2909, N2890, N2519);
and AND3 (N2910, N2907, N1247, N2727);
nand NAND4 (N2911, N2902, N928, N2865, N2698);
nor NOR2 (N2912, N2909, N2763);
nor NOR4 (N2913, N2910, N1684, N1228, N1060);
nor NOR2 (N2914, N2896, N202);
not NOT1 (N2915, N2908);
xor XOR2 (N2916, N2913, N1717);
xor XOR2 (N2917, N2916, N767);
not NOT1 (N2918, N2901);
nor NOR2 (N2919, N2900, N2702);
buf BUF1 (N2920, N2914);
and AND4 (N2921, N2905, N1236, N32, N717);
or OR2 (N2922, N2904, N645);
xor XOR2 (N2923, N2911, N2249);
and AND4 (N2924, N2923, N2042, N2069, N2619);
xor XOR2 (N2925, N2920, N1511);
nor NOR2 (N2926, N2924, N2310);
nor NOR3 (N2927, N2918, N2820, N2510);
and AND2 (N2928, N2919, N1229);
nand NAND4 (N2929, N2927, N2858, N199, N556);
or OR3 (N2930, N2906, N2882, N881);
and AND2 (N2931, N2912, N1171);
not NOT1 (N2932, N2928);
not NOT1 (N2933, N2929);
nand NAND2 (N2934, N2921, N1834);
not NOT1 (N2935, N2926);
buf BUF1 (N2936, N2932);
and AND2 (N2937, N2933, N2157);
buf BUF1 (N2938, N2936);
and AND3 (N2939, N2938, N2090, N2626);
nor NOR3 (N2940, N2934, N25, N2086);
xor XOR2 (N2941, N2935, N1602);
nor NOR4 (N2942, N2917, N349, N606, N1793);
xor XOR2 (N2943, N2922, N130);
or OR4 (N2944, N2942, N888, N893, N1414);
nand NAND3 (N2945, N2941, N1061, N746);
buf BUF1 (N2946, N2944);
xor XOR2 (N2947, N2946, N1892);
nor NOR2 (N2948, N2937, N2041);
and AND2 (N2949, N2939, N944);
nor NOR4 (N2950, N2925, N1549, N2684, N2406);
not NOT1 (N2951, N2948);
or OR4 (N2952, N2930, N1017, N2909, N428);
buf BUF1 (N2953, N2940);
nand NAND4 (N2954, N2943, N652, N2638, N81);
nand NAND3 (N2955, N2954, N2691, N2922);
buf BUF1 (N2956, N2915);
or OR4 (N2957, N2955, N1872, N2799, N2521);
and AND4 (N2958, N2957, N2874, N1944, N972);
and AND3 (N2959, N2945, N2301, N1107);
not NOT1 (N2960, N2959);
not NOT1 (N2961, N2952);
nand NAND4 (N2962, N2953, N1444, N1617, N2790);
not NOT1 (N2963, N2931);
nor NOR4 (N2964, N2961, N275, N2092, N760);
nand NAND3 (N2965, N2964, N652, N2654);
not NOT1 (N2966, N2960);
xor XOR2 (N2967, N2949, N566);
buf BUF1 (N2968, N2958);
nand NAND4 (N2969, N2967, N513, N650, N277);
xor XOR2 (N2970, N2966, N1253);
or OR4 (N2971, N2951, N2582, N550, N235);
buf BUF1 (N2972, N2950);
nand NAND2 (N2973, N2956, N484);
buf BUF1 (N2974, N2973);
xor XOR2 (N2975, N2971, N2375);
or OR3 (N2976, N2972, N814, N1986);
and AND2 (N2977, N2974, N1335);
and AND4 (N2978, N2970, N1089, N1249, N1994);
not NOT1 (N2979, N2975);
xor XOR2 (N2980, N2947, N1016);
xor XOR2 (N2981, N2963, N930);
not NOT1 (N2982, N2978);
buf BUF1 (N2983, N2969);
not NOT1 (N2984, N2977);
or OR2 (N2985, N2976, N2833);
or OR3 (N2986, N2965, N2585, N1551);
and AND2 (N2987, N2980, N1443);
not NOT1 (N2988, N2968);
nor NOR3 (N2989, N2962, N1372, N113);
xor XOR2 (N2990, N2989, N2648);
or OR4 (N2991, N2986, N2601, N1498, N1918);
xor XOR2 (N2992, N2981, N188);
nor NOR4 (N2993, N2987, N37, N1548, N360);
xor XOR2 (N2994, N2979, N1576);
and AND2 (N2995, N2994, N1885);
buf BUF1 (N2996, N2995);
xor XOR2 (N2997, N2996, N2301);
buf BUF1 (N2998, N2993);
xor XOR2 (N2999, N2983, N2086);
xor XOR2 (N3000, N2985, N1405);
not NOT1 (N3001, N2999);
buf BUF1 (N3002, N2982);
and AND3 (N3003, N2990, N2461, N2618);
nor NOR2 (N3004, N3003, N1474);
nand NAND4 (N3005, N2991, N1384, N2200, N2850);
not NOT1 (N3006, N2998);
nand NAND2 (N3007, N3002, N2160);
not NOT1 (N3008, N2992);
nand NAND3 (N3009, N3001, N892, N465);
not NOT1 (N3010, N3000);
nand NAND2 (N3011, N2988, N998);
nand NAND3 (N3012, N3011, N1707, N710);
and AND3 (N3013, N2984, N883, N2009);
not NOT1 (N3014, N3006);
buf BUF1 (N3015, N3014);
endmodule