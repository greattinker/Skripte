// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N716,N719,N668,N711,N708,N710,N717,N701,N713,N720;

and AND2 (N21, N11, N3);
or OR3 (N22, N21, N10, N3);
and AND4 (N23, N18, N3, N8, N6);
xor XOR2 (N24, N15, N22);
nand NAND4 (N25, N4, N2, N9, N10);
nand NAND2 (N26, N25, N25);
nand NAND4 (N27, N26, N15, N25, N5);
or OR4 (N28, N23, N18, N27, N26);
xor XOR2 (N29, N8, N19);
not NOT1 (N30, N6);
and AND2 (N31, N24, N21);
or OR3 (N32, N26, N22, N12);
xor XOR2 (N33, N24, N4);
buf BUF1 (N34, N21);
or OR3 (N35, N18, N4, N32);
or OR2 (N36, N14, N2);
buf BUF1 (N37, N31);
or OR2 (N38, N1, N29);
nor NOR2 (N39, N29, N33);
and AND2 (N40, N15, N30);
and AND4 (N41, N35, N29, N24, N37);
buf BUF1 (N42, N19);
nor NOR3 (N43, N38, N16, N35);
buf BUF1 (N44, N13);
nand NAND2 (N45, N15, N20);
nand NAND3 (N46, N40, N10, N13);
xor XOR2 (N47, N28, N16);
buf BUF1 (N48, N46);
and AND2 (N49, N44, N18);
buf BUF1 (N50, N45);
or OR3 (N51, N34, N3, N22);
and AND4 (N52, N48, N11, N17, N2);
not NOT1 (N53, N50);
nand NAND3 (N54, N49, N10, N32);
or OR3 (N55, N54, N21, N51);
and AND4 (N56, N49, N29, N12, N38);
not NOT1 (N57, N55);
or OR2 (N58, N56, N46);
nand NAND2 (N59, N39, N34);
nor NOR2 (N60, N57, N24);
not NOT1 (N61, N47);
not NOT1 (N62, N41);
buf BUF1 (N63, N59);
nand NAND2 (N64, N58, N41);
nand NAND4 (N65, N52, N50, N1, N1);
buf BUF1 (N66, N62);
nand NAND2 (N67, N60, N24);
xor XOR2 (N68, N36, N31);
and AND2 (N69, N64, N59);
not NOT1 (N70, N61);
or OR2 (N71, N43, N12);
nor NOR2 (N72, N65, N59);
buf BUF1 (N73, N42);
and AND3 (N74, N71, N49, N24);
xor XOR2 (N75, N67, N56);
nand NAND2 (N76, N66, N37);
or OR2 (N77, N73, N62);
xor XOR2 (N78, N53, N46);
nor NOR2 (N79, N77, N52);
buf BUF1 (N80, N74);
nor NOR2 (N81, N79, N14);
buf BUF1 (N82, N80);
xor XOR2 (N83, N63, N49);
and AND2 (N84, N70, N2);
nand NAND3 (N85, N68, N55, N19);
nor NOR2 (N86, N69, N79);
xor XOR2 (N87, N83, N26);
and AND3 (N88, N87, N84, N66);
nand NAND2 (N89, N46, N42);
nand NAND2 (N90, N88, N61);
nand NAND3 (N91, N90, N13, N20);
xor XOR2 (N92, N91, N51);
or OR2 (N93, N89, N25);
nand NAND4 (N94, N86, N39, N28, N80);
buf BUF1 (N95, N72);
xor XOR2 (N96, N95, N8);
buf BUF1 (N97, N85);
and AND2 (N98, N78, N24);
not NOT1 (N99, N75);
nor NOR4 (N100, N92, N66, N6, N14);
nor NOR2 (N101, N81, N94);
buf BUF1 (N102, N75);
xor XOR2 (N103, N96, N45);
and AND2 (N104, N103, N51);
not NOT1 (N105, N100);
nand NAND3 (N106, N97, N30, N67);
and AND3 (N107, N102, N88, N17);
buf BUF1 (N108, N93);
nand NAND4 (N109, N101, N62, N14, N14);
nand NAND2 (N110, N108, N74);
not NOT1 (N111, N105);
nor NOR3 (N112, N111, N53, N95);
nor NOR4 (N113, N106, N59, N56, N79);
or OR2 (N114, N82, N37);
and AND4 (N115, N99, N36, N84, N29);
nand NAND4 (N116, N115, N31, N84, N4);
buf BUF1 (N117, N107);
not NOT1 (N118, N76);
not NOT1 (N119, N109);
and AND2 (N120, N98, N117);
buf BUF1 (N121, N25);
nand NAND2 (N122, N110, N9);
and AND2 (N123, N114, N31);
xor XOR2 (N124, N120, N61);
and AND4 (N125, N123, N51, N41, N64);
not NOT1 (N126, N119);
nand NAND4 (N127, N113, N31, N82, N76);
or OR4 (N128, N116, N70, N5, N70);
not NOT1 (N129, N112);
or OR4 (N130, N126, N88, N14, N81);
not NOT1 (N131, N130);
buf BUF1 (N132, N129);
not NOT1 (N133, N122);
buf BUF1 (N134, N125);
nor NOR3 (N135, N121, N128, N90);
xor XOR2 (N136, N103, N83);
and AND3 (N137, N104, N111, N112);
and AND4 (N138, N135, N137, N78, N81);
not NOT1 (N139, N67);
buf BUF1 (N140, N132);
not NOT1 (N141, N131);
or OR4 (N142, N127, N1, N68, N114);
nand NAND2 (N143, N133, N40);
not NOT1 (N144, N140);
buf BUF1 (N145, N124);
buf BUF1 (N146, N142);
or OR2 (N147, N134, N138);
xor XOR2 (N148, N19, N86);
buf BUF1 (N149, N141);
xor XOR2 (N150, N148, N42);
buf BUF1 (N151, N139);
nand NAND3 (N152, N136, N8, N56);
nor NOR3 (N153, N150, N145, N65);
and AND2 (N154, N17, N108);
and AND4 (N155, N149, N137, N50, N64);
not NOT1 (N156, N144);
and AND3 (N157, N151, N116, N59);
or OR3 (N158, N147, N79, N8);
nand NAND3 (N159, N156, N29, N19);
nor NOR3 (N160, N154, N8, N63);
or OR4 (N161, N118, N46, N59, N104);
not NOT1 (N162, N160);
nor NOR4 (N163, N143, N62, N135, N42);
or OR4 (N164, N162, N5, N147, N162);
buf BUF1 (N165, N163);
nor NOR3 (N166, N157, N32, N22);
and AND2 (N167, N164, N75);
not NOT1 (N168, N146);
nor NOR3 (N169, N161, N140, N161);
and AND3 (N170, N155, N27, N134);
and AND2 (N171, N169, N133);
xor XOR2 (N172, N153, N63);
buf BUF1 (N173, N152);
or OR3 (N174, N171, N6, N93);
or OR3 (N175, N172, N113, N149);
xor XOR2 (N176, N166, N46);
or OR2 (N177, N175, N45);
and AND3 (N178, N159, N127, N63);
nor NOR3 (N179, N176, N118, N170);
nor NOR2 (N180, N28, N133);
nand NAND2 (N181, N165, N120);
xor XOR2 (N182, N173, N110);
not NOT1 (N183, N174);
buf BUF1 (N184, N178);
nand NAND2 (N185, N158, N129);
nand NAND2 (N186, N177, N62);
buf BUF1 (N187, N184);
or OR2 (N188, N179, N137);
nor NOR3 (N189, N180, N76, N110);
not NOT1 (N190, N187);
and AND2 (N191, N186, N164);
xor XOR2 (N192, N168, N27);
buf BUF1 (N193, N183);
xor XOR2 (N194, N182, N80);
xor XOR2 (N195, N188, N194);
buf BUF1 (N196, N106);
nand NAND4 (N197, N193, N159, N177, N176);
or OR4 (N198, N196, N28, N11, N153);
xor XOR2 (N199, N190, N4);
and AND2 (N200, N199, N179);
and AND2 (N201, N191, N4);
buf BUF1 (N202, N192);
nor NOR2 (N203, N181, N25);
nor NOR2 (N204, N200, N60);
or OR2 (N205, N202, N192);
buf BUF1 (N206, N195);
and AND4 (N207, N206, N15, N144, N130);
buf BUF1 (N208, N197);
buf BUF1 (N209, N167);
and AND2 (N210, N203, N59);
buf BUF1 (N211, N204);
or OR2 (N212, N185, N204);
nor NOR2 (N213, N201, N77);
and AND2 (N214, N198, N113);
and AND3 (N215, N207, N45, N83);
nor NOR3 (N216, N214, N201, N173);
nor NOR4 (N217, N215, N202, N164, N53);
nor NOR4 (N218, N189, N172, N97, N194);
buf BUF1 (N219, N218);
buf BUF1 (N220, N205);
buf BUF1 (N221, N210);
not NOT1 (N222, N217);
or OR4 (N223, N208, N166, N160, N197);
xor XOR2 (N224, N223, N180);
buf BUF1 (N225, N220);
nor NOR2 (N226, N221, N135);
buf BUF1 (N227, N216);
buf BUF1 (N228, N219);
and AND3 (N229, N224, N210, N153);
nor NOR2 (N230, N209, N24);
buf BUF1 (N231, N211);
or OR2 (N232, N227, N77);
nand NAND2 (N233, N226, N144);
buf BUF1 (N234, N213);
nand NAND3 (N235, N225, N96, N54);
or OR4 (N236, N235, N48, N128, N8);
nand NAND4 (N237, N222, N141, N81, N197);
nor NOR4 (N238, N230, N141, N98, N208);
and AND3 (N239, N231, N188, N115);
buf BUF1 (N240, N212);
and AND2 (N241, N239, N101);
not NOT1 (N242, N229);
and AND4 (N243, N242, N124, N224, N206);
or OR4 (N244, N234, N41, N72, N47);
xor XOR2 (N245, N244, N51);
buf BUF1 (N246, N243);
nor NOR2 (N247, N240, N29);
nor NOR2 (N248, N247, N138);
buf BUF1 (N249, N238);
and AND3 (N250, N236, N15, N163);
not NOT1 (N251, N241);
and AND4 (N252, N246, N5, N166, N37);
nor NOR3 (N253, N233, N165, N181);
nor NOR4 (N254, N237, N149, N84, N194);
or OR2 (N255, N228, N20);
not NOT1 (N256, N232);
or OR3 (N257, N252, N29, N229);
not NOT1 (N258, N254);
buf BUF1 (N259, N245);
not NOT1 (N260, N256);
nor NOR3 (N261, N257, N208, N22);
nor NOR4 (N262, N253, N135, N202, N58);
not NOT1 (N263, N251);
nor NOR2 (N264, N250, N189);
and AND4 (N265, N249, N30, N175, N61);
not NOT1 (N266, N263);
nand NAND2 (N267, N259, N253);
or OR4 (N268, N264, N51, N128, N205);
buf BUF1 (N269, N265);
not NOT1 (N270, N267);
or OR2 (N271, N255, N224);
nor NOR4 (N272, N269, N176, N247, N131);
not NOT1 (N273, N271);
or OR3 (N274, N273, N227, N187);
nor NOR4 (N275, N260, N151, N39, N37);
nor NOR2 (N276, N268, N6);
and AND2 (N277, N248, N11);
or OR4 (N278, N272, N231, N213, N232);
or OR2 (N279, N262, N242);
not NOT1 (N280, N275);
buf BUF1 (N281, N279);
not NOT1 (N282, N266);
nor NOR4 (N283, N274, N139, N27, N143);
nand NAND2 (N284, N278, N154);
and AND4 (N285, N277, N146, N5, N256);
buf BUF1 (N286, N280);
nor NOR2 (N287, N270, N53);
and AND2 (N288, N287, N171);
and AND3 (N289, N258, N238, N59);
nor NOR3 (N290, N285, N113, N155);
not NOT1 (N291, N289);
nand NAND4 (N292, N281, N195, N154, N23);
buf BUF1 (N293, N261);
nand NAND2 (N294, N282, N86);
and AND3 (N295, N291, N42, N272);
and AND2 (N296, N292, N140);
not NOT1 (N297, N288);
xor XOR2 (N298, N286, N162);
buf BUF1 (N299, N295);
nor NOR3 (N300, N299, N134, N190);
nand NAND4 (N301, N283, N74, N256, N273);
or OR4 (N302, N294, N46, N126, N167);
nor NOR4 (N303, N284, N105, N150, N296);
buf BUF1 (N304, N114);
or OR2 (N305, N297, N89);
buf BUF1 (N306, N293);
nand NAND3 (N307, N304, N44, N99);
xor XOR2 (N308, N300, N128);
or OR4 (N309, N276, N61, N278, N227);
xor XOR2 (N310, N305, N14);
not NOT1 (N311, N306);
buf BUF1 (N312, N311);
nand NAND4 (N313, N302, N53, N121, N21);
or OR4 (N314, N308, N217, N42, N229);
xor XOR2 (N315, N309, N152);
not NOT1 (N316, N310);
nor NOR4 (N317, N303, N29, N73, N210);
buf BUF1 (N318, N301);
and AND3 (N319, N315, N221, N287);
buf BUF1 (N320, N314);
buf BUF1 (N321, N290);
and AND3 (N322, N319, N1, N146);
buf BUF1 (N323, N320);
and AND3 (N324, N312, N25, N289);
xor XOR2 (N325, N316, N208);
or OR2 (N326, N298, N41);
and AND4 (N327, N307, N82, N232, N140);
and AND2 (N328, N326, N207);
nor NOR2 (N329, N328, N24);
or OR3 (N330, N325, N15, N211);
nand NAND2 (N331, N330, N1);
xor XOR2 (N332, N331, N292);
or OR2 (N333, N332, N131);
or OR4 (N334, N317, N84, N300, N163);
not NOT1 (N335, N323);
xor XOR2 (N336, N318, N84);
not NOT1 (N337, N322);
nor NOR2 (N338, N335, N288);
not NOT1 (N339, N327);
buf BUF1 (N340, N313);
buf BUF1 (N341, N340);
nor NOR4 (N342, N341, N62, N287, N75);
and AND3 (N343, N337, N174, N125);
nor NOR3 (N344, N324, N220, N299);
buf BUF1 (N345, N338);
buf BUF1 (N346, N336);
buf BUF1 (N347, N334);
buf BUF1 (N348, N345);
nor NOR4 (N349, N339, N92, N332, N12);
or OR4 (N350, N342, N219, N109, N153);
or OR2 (N351, N333, N233);
xor XOR2 (N352, N348, N18);
and AND2 (N353, N349, N44);
buf BUF1 (N354, N343);
xor XOR2 (N355, N353, N40);
or OR2 (N356, N329, N14);
and AND3 (N357, N321, N343, N83);
or OR4 (N358, N356, N287, N289, N237);
not NOT1 (N359, N344);
xor XOR2 (N360, N354, N308);
xor XOR2 (N361, N346, N173);
and AND4 (N362, N359, N26, N63, N23);
not NOT1 (N363, N362);
and AND4 (N364, N363, N350, N132, N74);
and AND3 (N365, N198, N128, N78);
nor NOR4 (N366, N351, N307, N193, N161);
buf BUF1 (N367, N364);
and AND4 (N368, N365, N351, N233, N225);
or OR3 (N369, N367, N221, N2);
not NOT1 (N370, N368);
nand NAND4 (N371, N347, N23, N171, N345);
nor NOR2 (N372, N360, N175);
xor XOR2 (N373, N357, N166);
not NOT1 (N374, N366);
buf BUF1 (N375, N373);
buf BUF1 (N376, N352);
or OR3 (N377, N370, N155, N38);
nand NAND4 (N378, N371, N89, N177, N353);
nand NAND2 (N379, N376, N294);
and AND3 (N380, N358, N75, N16);
nor NOR4 (N381, N378, N213, N246, N342);
or OR2 (N382, N372, N66);
nor NOR3 (N383, N381, N78, N22);
xor XOR2 (N384, N355, N113);
nand NAND4 (N385, N380, N331, N270, N129);
or OR4 (N386, N369, N273, N75, N324);
nand NAND4 (N387, N385, N239, N368, N328);
nor NOR4 (N388, N386, N15, N225, N67);
nor NOR2 (N389, N361, N72);
and AND4 (N390, N382, N165, N313, N350);
nor NOR4 (N391, N377, N101, N199, N126);
not NOT1 (N392, N379);
xor XOR2 (N393, N383, N27);
nand NAND3 (N394, N388, N260, N300);
nand NAND3 (N395, N389, N25, N107);
not NOT1 (N396, N387);
and AND3 (N397, N392, N393, N28);
not NOT1 (N398, N100);
not NOT1 (N399, N395);
or OR4 (N400, N394, N297, N157, N4);
xor XOR2 (N401, N390, N75);
and AND2 (N402, N399, N85);
nand NAND4 (N403, N401, N197, N379, N51);
or OR2 (N404, N375, N21);
buf BUF1 (N405, N398);
xor XOR2 (N406, N402, N78);
buf BUF1 (N407, N400);
xor XOR2 (N408, N406, N290);
nand NAND2 (N409, N407, N132);
nand NAND4 (N410, N391, N207, N83, N136);
or OR2 (N411, N408, N157);
not NOT1 (N412, N411);
xor XOR2 (N413, N410, N302);
xor XOR2 (N414, N396, N368);
not NOT1 (N415, N384);
and AND2 (N416, N415, N10);
or OR2 (N417, N414, N157);
xor XOR2 (N418, N413, N264);
xor XOR2 (N419, N397, N255);
nand NAND4 (N420, N403, N249, N130, N184);
xor XOR2 (N421, N412, N121);
nand NAND3 (N422, N421, N138, N413);
buf BUF1 (N423, N418);
nand NAND3 (N424, N419, N79, N353);
nor NOR3 (N425, N404, N202, N31);
xor XOR2 (N426, N405, N94);
and AND4 (N427, N417, N93, N2, N347);
xor XOR2 (N428, N374, N96);
nor NOR2 (N429, N423, N213);
or OR4 (N430, N429, N358, N38, N212);
nand NAND2 (N431, N416, N392);
or OR3 (N432, N427, N45, N335);
and AND2 (N433, N430, N281);
not NOT1 (N434, N422);
or OR2 (N435, N433, N44);
nor NOR2 (N436, N425, N333);
and AND4 (N437, N434, N417, N185, N381);
xor XOR2 (N438, N409, N229);
buf BUF1 (N439, N424);
or OR3 (N440, N435, N325, N341);
nor NOR3 (N441, N428, N66, N221);
xor XOR2 (N442, N420, N78);
nor NOR3 (N443, N439, N128, N389);
or OR2 (N444, N431, N1);
or OR4 (N445, N437, N429, N122, N328);
or OR3 (N446, N438, N84, N241);
nor NOR2 (N447, N443, N383);
or OR3 (N448, N441, N433, N349);
or OR3 (N449, N432, N231, N132);
not NOT1 (N450, N436);
not NOT1 (N451, N446);
nor NOR4 (N452, N426, N25, N247, N120);
not NOT1 (N453, N452);
buf BUF1 (N454, N442);
or OR2 (N455, N454, N204);
buf BUF1 (N456, N447);
nand NAND2 (N457, N456, N110);
and AND3 (N458, N451, N178, N106);
and AND2 (N459, N453, N135);
not NOT1 (N460, N449);
nor NOR4 (N461, N440, N430, N2, N42);
buf BUF1 (N462, N458);
nand NAND2 (N463, N457, N306);
not NOT1 (N464, N460);
or OR4 (N465, N450, N102, N30, N295);
not NOT1 (N466, N464);
and AND4 (N467, N444, N103, N177, N446);
xor XOR2 (N468, N459, N431);
nand NAND4 (N469, N465, N200, N97, N366);
and AND2 (N470, N445, N325);
not NOT1 (N471, N466);
not NOT1 (N472, N462);
nor NOR2 (N473, N461, N97);
buf BUF1 (N474, N467);
buf BUF1 (N475, N472);
or OR3 (N476, N468, N157, N455);
and AND3 (N477, N367, N353, N91);
xor XOR2 (N478, N470, N289);
buf BUF1 (N479, N478);
xor XOR2 (N480, N475, N335);
xor XOR2 (N481, N480, N427);
nor NOR4 (N482, N474, N188, N460, N152);
not NOT1 (N483, N479);
not NOT1 (N484, N481);
xor XOR2 (N485, N476, N347);
or OR2 (N486, N483, N11);
xor XOR2 (N487, N477, N58);
not NOT1 (N488, N473);
nor NOR3 (N489, N448, N194, N147);
nand NAND2 (N490, N469, N100);
buf BUF1 (N491, N490);
buf BUF1 (N492, N487);
nor NOR3 (N493, N471, N297, N139);
nand NAND3 (N494, N485, N99, N31);
not NOT1 (N495, N493);
buf BUF1 (N496, N491);
buf BUF1 (N497, N482);
not NOT1 (N498, N497);
xor XOR2 (N499, N486, N116);
xor XOR2 (N500, N489, N225);
nor NOR2 (N501, N495, N69);
and AND2 (N502, N488, N466);
nor NOR2 (N503, N499, N386);
buf BUF1 (N504, N502);
not NOT1 (N505, N494);
buf BUF1 (N506, N492);
and AND4 (N507, N501, N159, N201, N8);
buf BUF1 (N508, N506);
nand NAND3 (N509, N503, N423, N351);
or OR4 (N510, N507, N210, N308, N489);
not NOT1 (N511, N463);
not NOT1 (N512, N510);
or OR4 (N513, N484, N433, N412, N34);
not NOT1 (N514, N498);
nor NOR4 (N515, N496, N283, N351, N452);
not NOT1 (N516, N509);
buf BUF1 (N517, N515);
nor NOR4 (N518, N511, N91, N24, N20);
nor NOR3 (N519, N514, N437, N205);
nand NAND2 (N520, N508, N305);
nor NOR4 (N521, N504, N119, N232, N453);
or OR3 (N522, N517, N366, N457);
nor NOR4 (N523, N519, N200, N145, N516);
buf BUF1 (N524, N221);
and AND2 (N525, N505, N1);
nand NAND3 (N526, N525, N110, N166);
buf BUF1 (N527, N520);
xor XOR2 (N528, N524, N523);
or OR3 (N529, N302, N128, N303);
nand NAND3 (N530, N528, N190, N251);
nand NAND2 (N531, N513, N175);
and AND4 (N532, N500, N470, N473, N510);
or OR3 (N533, N522, N195, N424);
and AND4 (N534, N521, N444, N141, N170);
nor NOR4 (N535, N527, N420, N157, N299);
buf BUF1 (N536, N518);
nor NOR3 (N537, N533, N390, N497);
or OR3 (N538, N537, N411, N288);
buf BUF1 (N539, N534);
and AND2 (N540, N529, N358);
xor XOR2 (N541, N526, N240);
nor NOR4 (N542, N541, N204, N103, N498);
or OR4 (N543, N535, N459, N200, N113);
nor NOR4 (N544, N539, N304, N308, N530);
nor NOR2 (N545, N512, N454);
and AND2 (N546, N195, N99);
nor NOR2 (N547, N545, N125);
nand NAND3 (N548, N542, N395, N174);
nor NOR4 (N549, N532, N106, N122, N271);
xor XOR2 (N550, N543, N13);
and AND2 (N551, N531, N536);
nand NAND4 (N552, N93, N70, N111, N371);
not NOT1 (N553, N551);
not NOT1 (N554, N546);
or OR2 (N555, N549, N367);
not NOT1 (N556, N548);
xor XOR2 (N557, N540, N280);
and AND2 (N558, N556, N423);
buf BUF1 (N559, N544);
not NOT1 (N560, N552);
xor XOR2 (N561, N557, N127);
nand NAND4 (N562, N550, N101, N524, N167);
nand NAND4 (N563, N559, N341, N77, N94);
xor XOR2 (N564, N555, N55);
and AND2 (N565, N560, N143);
xor XOR2 (N566, N563, N142);
xor XOR2 (N567, N561, N467);
xor XOR2 (N568, N538, N501);
or OR3 (N569, N562, N222, N480);
or OR3 (N570, N564, N215, N526);
buf BUF1 (N571, N567);
xor XOR2 (N572, N553, N59);
xor XOR2 (N573, N565, N278);
not NOT1 (N574, N566);
or OR3 (N575, N571, N423, N264);
or OR3 (N576, N572, N55, N383);
nand NAND4 (N577, N573, N511, N43, N348);
or OR4 (N578, N570, N67, N329, N559);
and AND4 (N579, N576, N572, N252, N4);
not NOT1 (N580, N568);
nor NOR4 (N581, N554, N89, N73, N13);
nand NAND3 (N582, N580, N438, N157);
and AND2 (N583, N575, N26);
not NOT1 (N584, N574);
nand NAND2 (N585, N582, N189);
and AND4 (N586, N569, N169, N248, N481);
nor NOR2 (N587, N577, N22);
buf BUF1 (N588, N585);
not NOT1 (N589, N547);
buf BUF1 (N590, N586);
not NOT1 (N591, N583);
buf BUF1 (N592, N581);
nand NAND2 (N593, N558, N57);
and AND4 (N594, N590, N282, N373, N507);
nand NAND2 (N595, N588, N493);
not NOT1 (N596, N592);
not NOT1 (N597, N593);
nor NOR4 (N598, N584, N44, N304, N248);
not NOT1 (N599, N587);
or OR4 (N600, N598, N488, N50, N66);
not NOT1 (N601, N591);
not NOT1 (N602, N589);
buf BUF1 (N603, N600);
or OR3 (N604, N579, N584, N114);
and AND2 (N605, N595, N187);
buf BUF1 (N606, N597);
and AND2 (N607, N601, N374);
nand NAND4 (N608, N604, N172, N334, N343);
not NOT1 (N609, N594);
buf BUF1 (N610, N608);
not NOT1 (N611, N606);
not NOT1 (N612, N610);
xor XOR2 (N613, N611, N33);
and AND2 (N614, N612, N398);
nor NOR3 (N615, N578, N87, N244);
and AND2 (N616, N615, N350);
or OR4 (N617, N613, N608, N84, N608);
nand NAND2 (N618, N603, N192);
not NOT1 (N619, N616);
or OR4 (N620, N614, N302, N470, N221);
xor XOR2 (N621, N596, N392);
not NOT1 (N622, N617);
and AND2 (N623, N599, N175);
not NOT1 (N624, N605);
not NOT1 (N625, N609);
or OR4 (N626, N625, N430, N541, N498);
not NOT1 (N627, N620);
xor XOR2 (N628, N627, N302);
not NOT1 (N629, N618);
nand NAND4 (N630, N602, N296, N398, N11);
nor NOR4 (N631, N621, N9, N588, N612);
xor XOR2 (N632, N629, N369);
or OR3 (N633, N619, N326, N446);
not NOT1 (N634, N631);
or OR3 (N635, N633, N302, N368);
nand NAND3 (N636, N624, N399, N30);
xor XOR2 (N637, N634, N106);
nor NOR2 (N638, N630, N127);
or OR2 (N639, N635, N393);
nand NAND3 (N640, N607, N55, N285);
or OR3 (N641, N637, N181, N73);
buf BUF1 (N642, N622);
not NOT1 (N643, N640);
nand NAND2 (N644, N643, N86);
nor NOR3 (N645, N644, N611, N341);
or OR4 (N646, N642, N42, N384, N635);
not NOT1 (N647, N646);
xor XOR2 (N648, N641, N503);
and AND2 (N649, N623, N262);
not NOT1 (N650, N636);
buf BUF1 (N651, N648);
buf BUF1 (N652, N651);
nor NOR4 (N653, N649, N62, N620, N320);
not NOT1 (N654, N639);
nor NOR4 (N655, N654, N113, N272, N634);
xor XOR2 (N656, N632, N539);
buf BUF1 (N657, N650);
buf BUF1 (N658, N652);
not NOT1 (N659, N656);
or OR4 (N660, N647, N363, N5, N494);
nand NAND4 (N661, N655, N387, N42, N396);
xor XOR2 (N662, N657, N400);
nand NAND4 (N663, N645, N167, N334, N548);
nand NAND3 (N664, N662, N58, N150);
nor NOR4 (N665, N658, N439, N32, N206);
not NOT1 (N666, N626);
and AND2 (N667, N628, N244);
nand NAND2 (N668, N663, N542);
and AND2 (N669, N667, N197);
xor XOR2 (N670, N659, N216);
nor NOR3 (N671, N666, N161, N383);
xor XOR2 (N672, N671, N546);
and AND4 (N673, N672, N277, N275, N11);
nor NOR4 (N674, N670, N223, N583, N48);
xor XOR2 (N675, N674, N146);
nor NOR3 (N676, N665, N372, N262);
nor NOR4 (N677, N676, N597, N334, N464);
nor NOR3 (N678, N669, N151, N473);
or OR4 (N679, N660, N407, N405, N390);
nand NAND3 (N680, N673, N452, N87);
or OR4 (N681, N661, N658, N409, N493);
not NOT1 (N682, N679);
nor NOR2 (N683, N653, N194);
or OR4 (N684, N678, N527, N228, N86);
nand NAND4 (N685, N683, N224, N562, N400);
or OR3 (N686, N638, N606, N356);
nand NAND4 (N687, N684, N492, N343, N585);
buf BUF1 (N688, N677);
not NOT1 (N689, N664);
or OR3 (N690, N680, N396, N289);
nor NOR3 (N691, N675, N612, N214);
buf BUF1 (N692, N687);
xor XOR2 (N693, N685, N676);
nor NOR4 (N694, N682, N205, N600, N12);
nand NAND3 (N695, N692, N111, N499);
xor XOR2 (N696, N690, N516);
xor XOR2 (N697, N695, N457);
nor NOR3 (N698, N694, N472, N271);
nand NAND2 (N699, N693, N270);
or OR3 (N700, N697, N348, N40);
or OR4 (N701, N681, N320, N572, N128);
and AND3 (N702, N698, N559, N457);
xor XOR2 (N703, N688, N150);
nor NOR3 (N704, N700, N652, N516);
and AND3 (N705, N691, N225, N648);
not NOT1 (N706, N703);
and AND2 (N707, N689, N406);
nand NAND4 (N708, N704, N667, N535, N42);
nor NOR3 (N709, N707, N33, N444);
nor NOR4 (N710, N702, N386, N634, N92);
xor XOR2 (N711, N706, N359);
xor XOR2 (N712, N709, N106);
or OR2 (N713, N712, N475);
buf BUF1 (N714, N696);
nand NAND3 (N715, N714, N588, N160);
xor XOR2 (N716, N715, N219);
buf BUF1 (N717, N699);
or OR3 (N718, N686, N322, N202);
not NOT1 (N719, N705);
xor XOR2 (N720, N718, N339);
endmodule