// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N1618,N1614,N1613,N1617,N1622,N1620,N1599,N1615,N1621,N1623;

or OR4 (N24, N4, N19, N7, N17);
nand NAND4 (N25, N13, N22, N19, N7);
not NOT1 (N26, N25);
nand NAND3 (N27, N8, N1, N20);
buf BUF1 (N28, N6);
nor NOR3 (N29, N9, N15, N4);
nor NOR2 (N30, N4, N15);
not NOT1 (N31, N17);
not NOT1 (N32, N24);
nor NOR3 (N33, N12, N12, N18);
not NOT1 (N34, N6);
nor NOR2 (N35, N1, N2);
and AND3 (N36, N33, N17, N9);
or OR4 (N37, N32, N1, N1, N15);
buf BUF1 (N38, N34);
xor XOR2 (N39, N35, N30);
or OR4 (N40, N29, N26, N10, N37);
or OR2 (N41, N20, N13);
xor XOR2 (N42, N25, N39);
xor XOR2 (N43, N2, N14);
or OR4 (N44, N12, N9, N36, N6);
buf BUF1 (N45, N8);
buf BUF1 (N46, N45);
nand NAND4 (N47, N41, N5, N43, N39);
xor XOR2 (N48, N1, N33);
nand NAND2 (N49, N31, N29);
nand NAND3 (N50, N42, N1, N32);
xor XOR2 (N51, N47, N8);
nand NAND4 (N52, N27, N48, N42, N7);
or OR3 (N53, N10, N20, N36);
xor XOR2 (N54, N50, N51);
nand NAND2 (N55, N35, N1);
nor NOR3 (N56, N52, N53, N25);
not NOT1 (N57, N55);
or OR3 (N58, N23, N13, N32);
not NOT1 (N59, N58);
not NOT1 (N60, N54);
nor NOR4 (N61, N59, N17, N42, N21);
or OR4 (N62, N49, N38, N27, N12);
and AND3 (N63, N40, N48, N8);
not NOT1 (N64, N28);
or OR3 (N65, N41, N40, N63);
xor XOR2 (N66, N27, N47);
not NOT1 (N67, N64);
and AND2 (N68, N62, N23);
nand NAND3 (N69, N66, N48, N57);
xor XOR2 (N70, N61, N12);
or OR4 (N71, N54, N50, N48, N5);
not NOT1 (N72, N71);
not NOT1 (N73, N67);
buf BUF1 (N74, N65);
xor XOR2 (N75, N73, N22);
and AND4 (N76, N70, N59, N24, N27);
not NOT1 (N77, N68);
or OR2 (N78, N60, N48);
buf BUF1 (N79, N78);
buf BUF1 (N80, N79);
nand NAND4 (N81, N46, N71, N2, N4);
not NOT1 (N82, N74);
nor NOR4 (N83, N72, N5, N8, N11);
not NOT1 (N84, N81);
and AND3 (N85, N56, N70, N12);
nor NOR2 (N86, N82, N42);
nor NOR4 (N87, N69, N37, N44, N43);
nand NAND3 (N88, N76, N70, N4);
buf BUF1 (N89, N72);
or OR2 (N90, N75, N30);
or OR3 (N91, N80, N56, N47);
buf BUF1 (N92, N87);
xor XOR2 (N93, N92, N50);
nand NAND2 (N94, N89, N2);
xor XOR2 (N95, N93, N91);
xor XOR2 (N96, N33, N27);
and AND4 (N97, N77, N94, N35, N77);
nand NAND3 (N98, N77, N60, N2);
and AND3 (N99, N83, N91, N81);
nor NOR2 (N100, N97, N71);
not NOT1 (N101, N85);
or OR4 (N102, N86, N57, N42, N60);
and AND3 (N103, N88, N50, N20);
buf BUF1 (N104, N102);
buf BUF1 (N105, N95);
buf BUF1 (N106, N100);
nand NAND2 (N107, N84, N84);
nand NAND4 (N108, N104, N18, N17, N51);
buf BUF1 (N109, N108);
nor NOR3 (N110, N90, N11, N26);
or OR3 (N111, N107, N71, N54);
nand NAND3 (N112, N98, N80, N53);
not NOT1 (N113, N103);
and AND2 (N114, N106, N79);
and AND4 (N115, N101, N74, N104, N26);
or OR2 (N116, N109, N50);
not NOT1 (N117, N110);
buf BUF1 (N118, N114);
xor XOR2 (N119, N116, N62);
nand NAND3 (N120, N99, N56, N52);
not NOT1 (N121, N120);
xor XOR2 (N122, N96, N100);
buf BUF1 (N123, N121);
nand NAND3 (N124, N123, N74, N110);
and AND3 (N125, N117, N21, N9);
nand NAND2 (N126, N113, N23);
nand NAND2 (N127, N119, N103);
nand NAND4 (N128, N122, N22, N118, N120);
nor NOR4 (N129, N35, N35, N1, N66);
nand NAND3 (N130, N112, N71, N20);
xor XOR2 (N131, N128, N23);
nor NOR2 (N132, N126, N57);
and AND2 (N133, N132, N42);
buf BUF1 (N134, N105);
nor NOR3 (N135, N127, N67, N80);
not NOT1 (N136, N130);
buf BUF1 (N137, N136);
nand NAND4 (N138, N134, N113, N117, N39);
xor XOR2 (N139, N129, N104);
not NOT1 (N140, N133);
nand NAND3 (N141, N139, N140, N84);
xor XOR2 (N142, N119, N137);
buf BUF1 (N143, N127);
nor NOR2 (N144, N138, N15);
nor NOR3 (N145, N141, N137, N109);
or OR2 (N146, N144, N16);
or OR2 (N147, N146, N40);
nor NOR2 (N148, N115, N109);
or OR4 (N149, N143, N65, N60, N123);
not NOT1 (N150, N142);
buf BUF1 (N151, N111);
and AND3 (N152, N149, N81, N95);
not NOT1 (N153, N125);
nand NAND4 (N154, N131, N53, N59, N35);
and AND3 (N155, N153, N65, N3);
or OR3 (N156, N151, N64, N3);
or OR4 (N157, N156, N7, N2, N40);
nor NOR2 (N158, N148, N35);
xor XOR2 (N159, N152, N77);
xor XOR2 (N160, N157, N97);
not NOT1 (N161, N145);
xor XOR2 (N162, N161, N19);
not NOT1 (N163, N150);
and AND3 (N164, N154, N60, N121);
nand NAND4 (N165, N164, N105, N98, N33);
buf BUF1 (N166, N124);
xor XOR2 (N167, N159, N110);
xor XOR2 (N168, N167, N51);
and AND2 (N169, N166, N133);
xor XOR2 (N170, N158, N113);
xor XOR2 (N171, N147, N142);
and AND2 (N172, N170, N145);
nand NAND2 (N173, N172, N104);
buf BUF1 (N174, N169);
nor NOR4 (N175, N165, N126, N11, N107);
and AND4 (N176, N162, N135, N42, N109);
or OR3 (N177, N152, N125, N148);
or OR4 (N178, N168, N107, N163, N76);
or OR2 (N179, N97, N157);
buf BUF1 (N180, N174);
xor XOR2 (N181, N177, N94);
buf BUF1 (N182, N180);
not NOT1 (N183, N155);
xor XOR2 (N184, N182, N17);
buf BUF1 (N185, N173);
not NOT1 (N186, N179);
or OR2 (N187, N185, N112);
xor XOR2 (N188, N187, N111);
nor NOR3 (N189, N160, N32, N101);
buf BUF1 (N190, N188);
and AND3 (N191, N171, N122, N110);
nand NAND2 (N192, N178, N173);
xor XOR2 (N193, N184, N128);
not NOT1 (N194, N176);
or OR2 (N195, N192, N44);
not NOT1 (N196, N194);
and AND4 (N197, N193, N34, N122, N38);
and AND2 (N198, N186, N194);
nor NOR3 (N199, N191, N155, N100);
nor NOR3 (N200, N181, N157, N14);
xor XOR2 (N201, N175, N38);
buf BUF1 (N202, N201);
xor XOR2 (N203, N199, N35);
and AND4 (N204, N195, N92, N14, N15);
or OR4 (N205, N190, N99, N52, N112);
nand NAND3 (N206, N189, N60, N39);
buf BUF1 (N207, N204);
buf BUF1 (N208, N205);
xor XOR2 (N209, N197, N172);
nand NAND3 (N210, N207, N68, N48);
or OR4 (N211, N183, N199, N153, N70);
or OR4 (N212, N208, N92, N201, N83);
or OR3 (N213, N202, N69, N201);
or OR4 (N214, N209, N35, N119, N183);
or OR2 (N215, N206, N8);
or OR2 (N216, N200, N75);
xor XOR2 (N217, N196, N63);
buf BUF1 (N218, N214);
nor NOR4 (N219, N217, N121, N170, N46);
nor NOR2 (N220, N203, N196);
or OR3 (N221, N212, N219, N176);
and AND3 (N222, N67, N80, N45);
nand NAND2 (N223, N220, N181);
not NOT1 (N224, N216);
nor NOR4 (N225, N221, N61, N110, N207);
and AND4 (N226, N213, N42, N93, N70);
or OR4 (N227, N211, N78, N39, N214);
not NOT1 (N228, N218);
nor NOR4 (N229, N227, N198, N61, N140);
buf BUF1 (N230, N70);
xor XOR2 (N231, N229, N2);
xor XOR2 (N232, N230, N71);
xor XOR2 (N233, N222, N93);
or OR2 (N234, N215, N138);
xor XOR2 (N235, N234, N197);
xor XOR2 (N236, N232, N78);
buf BUF1 (N237, N224);
xor XOR2 (N238, N237, N199);
not NOT1 (N239, N235);
nand NAND2 (N240, N231, N63);
buf BUF1 (N241, N240);
and AND4 (N242, N226, N92, N7, N49);
buf BUF1 (N243, N233);
and AND4 (N244, N228, N8, N77, N240);
nor NOR3 (N245, N244, N40, N92);
not NOT1 (N246, N243);
not NOT1 (N247, N223);
or OR3 (N248, N247, N31, N196);
or OR4 (N249, N248, N25, N156, N153);
buf BUF1 (N250, N245);
buf BUF1 (N251, N249);
nand NAND3 (N252, N239, N115, N46);
xor XOR2 (N253, N210, N37);
nor NOR3 (N254, N251, N166, N73);
not NOT1 (N255, N242);
or OR4 (N256, N246, N185, N92, N207);
or OR3 (N257, N241, N163, N45);
not NOT1 (N258, N254);
nand NAND4 (N259, N253, N32, N207, N217);
and AND2 (N260, N236, N94);
or OR4 (N261, N252, N208, N195, N17);
not NOT1 (N262, N238);
xor XOR2 (N263, N261, N135);
xor XOR2 (N264, N258, N15);
xor XOR2 (N265, N250, N71);
and AND3 (N266, N256, N117, N177);
nand NAND2 (N267, N255, N221);
buf BUF1 (N268, N265);
nor NOR3 (N269, N225, N197, N173);
buf BUF1 (N270, N269);
nand NAND4 (N271, N270, N236, N158, N170);
xor XOR2 (N272, N268, N23);
nand NAND2 (N273, N260, N234);
not NOT1 (N274, N259);
nand NAND4 (N275, N257, N147, N272, N219);
buf BUF1 (N276, N40);
nand NAND2 (N277, N264, N120);
not NOT1 (N278, N263);
nor NOR4 (N279, N277, N99, N191, N56);
xor XOR2 (N280, N275, N176);
nor NOR2 (N281, N274, N84);
or OR2 (N282, N276, N163);
nand NAND3 (N283, N281, N216, N20);
nor NOR3 (N284, N262, N127, N249);
not NOT1 (N285, N266);
nor NOR2 (N286, N284, N48);
not NOT1 (N287, N283);
nor NOR2 (N288, N278, N67);
or OR4 (N289, N273, N163, N168, N211);
nand NAND2 (N290, N288, N157);
and AND2 (N291, N287, N39);
not NOT1 (N292, N271);
nor NOR2 (N293, N282, N235);
or OR2 (N294, N267, N55);
xor XOR2 (N295, N280, N49);
or OR4 (N296, N285, N133, N207, N174);
not NOT1 (N297, N293);
and AND2 (N298, N279, N88);
not NOT1 (N299, N290);
xor XOR2 (N300, N299, N70);
not NOT1 (N301, N291);
and AND3 (N302, N296, N257, N255);
and AND4 (N303, N294, N58, N176, N209);
xor XOR2 (N304, N297, N169);
and AND2 (N305, N304, N45);
nand NAND3 (N306, N300, N194, N22);
or OR2 (N307, N295, N49);
buf BUF1 (N308, N292);
or OR3 (N309, N306, N294, N111);
not NOT1 (N310, N302);
and AND3 (N311, N303, N93, N297);
or OR3 (N312, N310, N130, N66);
nand NAND3 (N313, N301, N158, N62);
xor XOR2 (N314, N289, N246);
nand NAND4 (N315, N313, N226, N226, N219);
buf BUF1 (N316, N309);
or OR3 (N317, N305, N264, N299);
not NOT1 (N318, N312);
nor NOR2 (N319, N307, N213);
buf BUF1 (N320, N311);
or OR2 (N321, N317, N289);
or OR4 (N322, N321, N178, N22, N80);
not NOT1 (N323, N315);
not NOT1 (N324, N318);
or OR3 (N325, N322, N20, N319);
nor NOR2 (N326, N287, N50);
buf BUF1 (N327, N323);
not NOT1 (N328, N326);
and AND4 (N329, N316, N151, N299, N94);
buf BUF1 (N330, N298);
nand NAND2 (N331, N330, N111);
buf BUF1 (N332, N328);
nand NAND3 (N333, N308, N20, N17);
buf BUF1 (N334, N332);
nand NAND2 (N335, N320, N135);
nor NOR4 (N336, N334, N67, N267, N124);
nor NOR4 (N337, N327, N73, N136, N243);
buf BUF1 (N338, N335);
or OR3 (N339, N314, N281, N331);
or OR2 (N340, N16, N171);
not NOT1 (N341, N340);
nand NAND4 (N342, N324, N102, N73, N242);
nor NOR4 (N343, N342, N142, N167, N252);
and AND2 (N344, N338, N79);
nor NOR4 (N345, N344, N309, N74, N184);
and AND3 (N346, N329, N137, N231);
not NOT1 (N347, N346);
or OR3 (N348, N343, N12, N3);
nand NAND3 (N349, N325, N203, N273);
xor XOR2 (N350, N348, N277);
nor NOR3 (N351, N337, N88, N252);
xor XOR2 (N352, N339, N125);
or OR4 (N353, N352, N209, N348, N256);
nor NOR3 (N354, N353, N321, N286);
xor XOR2 (N355, N134, N132);
nor NOR3 (N356, N336, N51, N277);
xor XOR2 (N357, N355, N269);
xor XOR2 (N358, N349, N247);
not NOT1 (N359, N350);
not NOT1 (N360, N347);
nand NAND4 (N361, N358, N301, N235, N257);
nand NAND2 (N362, N359, N207);
nand NAND4 (N363, N351, N293, N309, N77);
nor NOR4 (N364, N361, N237, N321, N110);
not NOT1 (N365, N333);
or OR2 (N366, N360, N346);
or OR4 (N367, N341, N216, N245, N60);
buf BUF1 (N368, N365);
or OR4 (N369, N364, N121, N359, N247);
nor NOR3 (N370, N366, N171, N93);
xor XOR2 (N371, N370, N12);
xor XOR2 (N372, N357, N186);
xor XOR2 (N373, N371, N197);
buf BUF1 (N374, N373);
and AND3 (N375, N356, N31, N8);
and AND2 (N376, N354, N234);
nand NAND3 (N377, N376, N182, N6);
or OR2 (N378, N374, N59);
or OR3 (N379, N363, N285, N150);
nor NOR4 (N380, N362, N163, N126, N116);
and AND3 (N381, N380, N83, N12);
nand NAND2 (N382, N381, N167);
not NOT1 (N383, N369);
or OR4 (N384, N375, N279, N136, N89);
nor NOR4 (N385, N367, N15, N253, N322);
and AND4 (N386, N382, N93, N268, N289);
buf BUF1 (N387, N345);
or OR3 (N388, N386, N345, N108);
or OR2 (N389, N372, N377);
or OR4 (N390, N68, N139, N74, N75);
not NOT1 (N391, N379);
buf BUF1 (N392, N389);
or OR3 (N393, N368, N37, N91);
buf BUF1 (N394, N384);
buf BUF1 (N395, N387);
xor XOR2 (N396, N391, N229);
nor NOR3 (N397, N396, N252, N265);
not NOT1 (N398, N392);
buf BUF1 (N399, N378);
or OR2 (N400, N395, N135);
xor XOR2 (N401, N383, N256);
and AND3 (N402, N397, N106, N51);
buf BUF1 (N403, N402);
not NOT1 (N404, N403);
not NOT1 (N405, N390);
nor NOR2 (N406, N399, N146);
nor NOR4 (N407, N388, N188, N302, N165);
and AND4 (N408, N393, N306, N21, N192);
xor XOR2 (N409, N405, N143);
nor NOR4 (N410, N385, N183, N120, N59);
nor NOR4 (N411, N398, N203, N344, N144);
nand NAND3 (N412, N410, N242, N125);
and AND2 (N413, N404, N178);
or OR3 (N414, N413, N212, N64);
not NOT1 (N415, N411);
xor XOR2 (N416, N401, N205);
buf BUF1 (N417, N394);
nor NOR4 (N418, N400, N339, N309, N403);
and AND3 (N419, N416, N2, N251);
buf BUF1 (N420, N409);
or OR4 (N421, N412, N182, N420, N376);
and AND2 (N422, N162, N228);
buf BUF1 (N423, N406);
buf BUF1 (N424, N408);
nor NOR2 (N425, N418, N254);
xor XOR2 (N426, N415, N425);
nand NAND3 (N427, N120, N75, N232);
and AND4 (N428, N423, N382, N323, N358);
nor NOR4 (N429, N427, N218, N362, N386);
not NOT1 (N430, N426);
nand NAND4 (N431, N417, N377, N389, N274);
nand NAND4 (N432, N421, N3, N386, N399);
nor NOR2 (N433, N422, N323);
or OR3 (N434, N407, N22, N317);
buf BUF1 (N435, N430);
or OR4 (N436, N432, N364, N141, N173);
or OR3 (N437, N419, N152, N408);
xor XOR2 (N438, N414, N153);
nand NAND3 (N439, N424, N122, N143);
xor XOR2 (N440, N434, N312);
nor NOR4 (N441, N439, N103, N40, N181);
buf BUF1 (N442, N438);
not NOT1 (N443, N440);
buf BUF1 (N444, N431);
and AND3 (N445, N436, N57, N238);
or OR3 (N446, N442, N183, N274);
and AND2 (N447, N446, N260);
nor NOR4 (N448, N433, N52, N4, N40);
or OR2 (N449, N447, N327);
nand NAND3 (N450, N445, N191, N210);
nand NAND2 (N451, N444, N429);
nand NAND4 (N452, N436, N427, N418, N396);
nand NAND4 (N453, N450, N310, N338, N86);
or OR4 (N454, N437, N70, N443, N119);
xor XOR2 (N455, N35, N137);
and AND2 (N456, N452, N59);
xor XOR2 (N457, N451, N284);
and AND2 (N458, N456, N149);
buf BUF1 (N459, N458);
xor XOR2 (N460, N428, N394);
xor XOR2 (N461, N454, N426);
and AND2 (N462, N453, N187);
nor NOR3 (N463, N462, N87, N179);
not NOT1 (N464, N455);
xor XOR2 (N465, N441, N221);
not NOT1 (N466, N457);
or OR2 (N467, N463, N161);
and AND4 (N468, N461, N35, N402, N118);
nor NOR3 (N469, N464, N294, N459);
nor NOR4 (N470, N413, N39, N323, N265);
nand NAND3 (N471, N469, N422, N148);
not NOT1 (N472, N449);
or OR3 (N473, N466, N10, N161);
and AND2 (N474, N460, N380);
not NOT1 (N475, N468);
buf BUF1 (N476, N470);
nand NAND2 (N477, N476, N275);
buf BUF1 (N478, N465);
nor NOR2 (N479, N473, N289);
nor NOR4 (N480, N475, N289, N437, N87);
nor NOR3 (N481, N467, N364, N446);
not NOT1 (N482, N471);
or OR2 (N483, N477, N467);
nor NOR2 (N484, N481, N251);
and AND4 (N485, N480, N331, N95, N271);
nand NAND2 (N486, N484, N452);
and AND2 (N487, N483, N417);
nor NOR3 (N488, N486, N94, N102);
and AND3 (N489, N435, N124, N63);
nor NOR2 (N490, N448, N345);
and AND3 (N491, N485, N18, N11);
buf BUF1 (N492, N479);
nand NAND3 (N493, N482, N492, N173);
buf BUF1 (N494, N156);
and AND2 (N495, N491, N217);
nor NOR2 (N496, N490, N384);
xor XOR2 (N497, N496, N277);
nand NAND3 (N498, N474, N93, N407);
xor XOR2 (N499, N472, N22);
or OR3 (N500, N495, N342, N435);
nor NOR2 (N501, N493, N456);
or OR4 (N502, N501, N239, N443, N338);
buf BUF1 (N503, N500);
and AND2 (N504, N488, N195);
nor NOR3 (N505, N494, N313, N104);
xor XOR2 (N506, N487, N230);
buf BUF1 (N507, N505);
xor XOR2 (N508, N506, N435);
xor XOR2 (N509, N508, N41);
not NOT1 (N510, N507);
xor XOR2 (N511, N509, N265);
or OR2 (N512, N489, N330);
xor XOR2 (N513, N497, N125);
and AND3 (N514, N511, N236, N266);
nand NAND4 (N515, N478, N56, N440, N182);
buf BUF1 (N516, N498);
and AND4 (N517, N504, N267, N340, N511);
buf BUF1 (N518, N516);
nor NOR2 (N519, N518, N58);
nand NAND4 (N520, N502, N375, N471, N508);
nand NAND3 (N521, N513, N240, N128);
buf BUF1 (N522, N499);
xor XOR2 (N523, N514, N431);
xor XOR2 (N524, N517, N347);
xor XOR2 (N525, N519, N242);
and AND3 (N526, N525, N242, N44);
or OR4 (N527, N524, N241, N501, N317);
not NOT1 (N528, N527);
nand NAND4 (N529, N523, N123, N482, N335);
or OR4 (N530, N512, N146, N27, N298);
or OR3 (N531, N521, N453, N263);
xor XOR2 (N532, N531, N159);
nand NAND2 (N533, N532, N175);
not NOT1 (N534, N533);
nor NOR2 (N535, N526, N477);
and AND4 (N536, N528, N207, N38, N243);
nand NAND2 (N537, N520, N49);
nand NAND4 (N538, N529, N74, N316, N341);
and AND2 (N539, N503, N443);
buf BUF1 (N540, N538);
xor XOR2 (N541, N515, N445);
buf BUF1 (N542, N530);
and AND2 (N543, N542, N354);
buf BUF1 (N544, N537);
nor NOR2 (N545, N543, N227);
buf BUF1 (N546, N534);
xor XOR2 (N547, N540, N252);
not NOT1 (N548, N539);
not NOT1 (N549, N510);
nor NOR3 (N550, N541, N235, N221);
nand NAND2 (N551, N535, N524);
nor NOR4 (N552, N546, N18, N390, N262);
nor NOR4 (N553, N522, N187, N233, N412);
not NOT1 (N554, N544);
not NOT1 (N555, N551);
xor XOR2 (N556, N555, N273);
not NOT1 (N557, N556);
nand NAND4 (N558, N547, N92, N28, N480);
xor XOR2 (N559, N548, N420);
xor XOR2 (N560, N558, N80);
nor NOR4 (N561, N552, N89, N167, N429);
and AND2 (N562, N557, N533);
nand NAND3 (N563, N554, N510, N5);
or OR2 (N564, N549, N34);
or OR4 (N565, N536, N92, N512, N452);
buf BUF1 (N566, N564);
buf BUF1 (N567, N562);
xor XOR2 (N568, N559, N185);
or OR3 (N569, N568, N377, N163);
and AND4 (N570, N545, N546, N5, N198);
or OR4 (N571, N570, N151, N293, N90);
not NOT1 (N572, N563);
nand NAND3 (N573, N569, N169, N287);
nor NOR2 (N574, N553, N431);
and AND2 (N575, N560, N246);
nand NAND3 (N576, N573, N170, N268);
or OR4 (N577, N574, N515, N255, N171);
buf BUF1 (N578, N572);
nor NOR4 (N579, N577, N156, N322, N224);
nand NAND3 (N580, N579, N158, N186);
nor NOR4 (N581, N578, N495, N201, N11);
buf BUF1 (N582, N567);
not NOT1 (N583, N566);
buf BUF1 (N584, N550);
nor NOR3 (N585, N580, N167, N152);
xor XOR2 (N586, N581, N554);
and AND2 (N587, N586, N62);
or OR3 (N588, N587, N218, N425);
and AND2 (N589, N575, N308);
nand NAND2 (N590, N583, N39);
xor XOR2 (N591, N589, N362);
nor NOR3 (N592, N582, N327, N548);
nor NOR2 (N593, N571, N224);
buf BUF1 (N594, N588);
nor NOR4 (N595, N565, N9, N539, N496);
xor XOR2 (N596, N590, N347);
or OR3 (N597, N585, N274, N362);
buf BUF1 (N598, N592);
buf BUF1 (N599, N598);
and AND2 (N600, N591, N557);
and AND2 (N601, N584, N360);
not NOT1 (N602, N597);
nor NOR2 (N603, N601, N195);
xor XOR2 (N604, N602, N157);
not NOT1 (N605, N600);
or OR4 (N606, N561, N274, N25, N495);
or OR4 (N607, N603, N244, N111, N251);
and AND2 (N608, N595, N549);
not NOT1 (N609, N606);
not NOT1 (N610, N608);
not NOT1 (N611, N609);
xor XOR2 (N612, N605, N570);
not NOT1 (N613, N607);
not NOT1 (N614, N596);
buf BUF1 (N615, N611);
nand NAND4 (N616, N612, N548, N375, N335);
or OR3 (N617, N576, N340, N174);
buf BUF1 (N618, N593);
nor NOR4 (N619, N616, N166, N242, N415);
buf BUF1 (N620, N614);
nor NOR3 (N621, N610, N484, N422);
or OR2 (N622, N620, N612);
xor XOR2 (N623, N599, N347);
buf BUF1 (N624, N618);
nor NOR3 (N625, N613, N506, N219);
nor NOR3 (N626, N594, N305, N92);
buf BUF1 (N627, N624);
buf BUF1 (N628, N619);
and AND3 (N629, N625, N54, N518);
or OR4 (N630, N627, N622, N274, N199);
or OR2 (N631, N550, N549);
xor XOR2 (N632, N628, N186);
nor NOR4 (N633, N626, N605, N247, N471);
nand NAND3 (N634, N617, N337, N202);
nand NAND3 (N635, N634, N274, N366);
xor XOR2 (N636, N630, N211);
xor XOR2 (N637, N621, N77);
and AND4 (N638, N632, N79, N253, N540);
buf BUF1 (N639, N638);
buf BUF1 (N640, N639);
xor XOR2 (N641, N635, N572);
nand NAND3 (N642, N629, N369, N636);
xor XOR2 (N643, N33, N4);
buf BUF1 (N644, N643);
xor XOR2 (N645, N623, N101);
buf BUF1 (N646, N633);
nand NAND2 (N647, N645, N324);
not NOT1 (N648, N637);
nor NOR4 (N649, N648, N494, N179, N420);
nor NOR3 (N650, N646, N178, N227);
and AND4 (N651, N642, N636, N523, N383);
not NOT1 (N652, N650);
nand NAND3 (N653, N649, N169, N171);
not NOT1 (N654, N644);
and AND2 (N655, N651, N557);
buf BUF1 (N656, N653);
and AND3 (N657, N647, N295, N240);
or OR2 (N658, N640, N58);
nor NOR3 (N659, N656, N175, N454);
buf BUF1 (N660, N659);
buf BUF1 (N661, N657);
xor XOR2 (N662, N654, N586);
not NOT1 (N663, N615);
nor NOR4 (N664, N655, N346, N467, N527);
buf BUF1 (N665, N664);
nand NAND3 (N666, N652, N583, N177);
or OR4 (N667, N631, N605, N309, N554);
or OR4 (N668, N663, N439, N642, N22);
not NOT1 (N669, N604);
nor NOR3 (N670, N666, N622, N112);
xor XOR2 (N671, N661, N505);
not NOT1 (N672, N660);
buf BUF1 (N673, N641);
or OR2 (N674, N672, N142);
nand NAND4 (N675, N662, N136, N199, N203);
nand NAND2 (N676, N667, N378);
buf BUF1 (N677, N670);
nor NOR3 (N678, N674, N204, N159);
and AND4 (N679, N675, N382, N68, N436);
not NOT1 (N680, N665);
buf BUF1 (N681, N679);
buf BUF1 (N682, N678);
xor XOR2 (N683, N671, N281);
and AND3 (N684, N680, N184, N313);
and AND3 (N685, N681, N588, N240);
not NOT1 (N686, N683);
xor XOR2 (N687, N658, N91);
or OR3 (N688, N673, N508, N91);
or OR3 (N689, N669, N233, N171);
xor XOR2 (N690, N676, N44);
or OR3 (N691, N688, N405, N5);
or OR3 (N692, N682, N413, N330);
xor XOR2 (N693, N687, N7);
xor XOR2 (N694, N668, N437);
nor NOR2 (N695, N691, N668);
not NOT1 (N696, N695);
or OR3 (N697, N689, N10, N610);
or OR4 (N698, N693, N238, N341, N149);
and AND3 (N699, N698, N304, N251);
or OR4 (N700, N690, N653, N544, N425);
nand NAND2 (N701, N686, N253);
buf BUF1 (N702, N685);
and AND4 (N703, N700, N302, N136, N302);
or OR4 (N704, N696, N91, N344, N567);
and AND4 (N705, N677, N48, N583, N256);
xor XOR2 (N706, N702, N85);
nor NOR3 (N707, N705, N306, N492);
not NOT1 (N708, N703);
or OR4 (N709, N692, N667, N442, N268);
xor XOR2 (N710, N708, N155);
not NOT1 (N711, N684);
nor NOR2 (N712, N701, N119);
nor NOR2 (N713, N697, N665);
or OR2 (N714, N707, N117);
and AND3 (N715, N714, N232, N288);
and AND4 (N716, N711, N690, N285, N17);
and AND3 (N717, N704, N655, N294);
xor XOR2 (N718, N715, N615);
or OR3 (N719, N706, N283, N390);
buf BUF1 (N720, N717);
xor XOR2 (N721, N716, N305);
not NOT1 (N722, N719);
nor NOR2 (N723, N710, N9);
buf BUF1 (N724, N720);
or OR3 (N725, N709, N722, N570);
buf BUF1 (N726, N452);
or OR4 (N727, N725, N555, N422, N596);
and AND2 (N728, N694, N589);
or OR4 (N729, N713, N714, N577, N159);
nand NAND4 (N730, N727, N329, N327, N233);
nor NOR3 (N731, N718, N471, N155);
and AND2 (N732, N724, N220);
or OR2 (N733, N726, N566);
and AND2 (N734, N732, N319);
xor XOR2 (N735, N734, N542);
or OR4 (N736, N735, N454, N631, N14);
and AND2 (N737, N733, N174);
not NOT1 (N738, N699);
xor XOR2 (N739, N712, N663);
not NOT1 (N740, N721);
nor NOR4 (N741, N739, N161, N465, N341);
not NOT1 (N742, N728);
buf BUF1 (N743, N731);
and AND2 (N744, N736, N414);
buf BUF1 (N745, N730);
not NOT1 (N746, N745);
nand NAND4 (N747, N723, N288, N27, N500);
buf BUF1 (N748, N743);
buf BUF1 (N749, N744);
xor XOR2 (N750, N742, N180);
buf BUF1 (N751, N741);
and AND4 (N752, N750, N556, N306, N33);
xor XOR2 (N753, N752, N658);
and AND2 (N754, N749, N45);
buf BUF1 (N755, N747);
and AND4 (N756, N737, N453, N197, N278);
not NOT1 (N757, N738);
nand NAND4 (N758, N754, N741, N560, N562);
not NOT1 (N759, N757);
and AND3 (N760, N755, N708, N240);
nor NOR3 (N761, N760, N253, N542);
nor NOR3 (N762, N761, N116, N362);
and AND3 (N763, N762, N252, N527);
xor XOR2 (N764, N753, N71);
and AND4 (N765, N758, N267, N265, N254);
nor NOR2 (N766, N740, N285);
not NOT1 (N767, N759);
buf BUF1 (N768, N751);
or OR2 (N769, N767, N565);
not NOT1 (N770, N763);
nor NOR2 (N771, N765, N734);
buf BUF1 (N772, N768);
xor XOR2 (N773, N746, N221);
buf BUF1 (N774, N764);
and AND3 (N775, N771, N512, N739);
not NOT1 (N776, N748);
and AND2 (N777, N774, N708);
or OR3 (N778, N772, N462, N396);
xor XOR2 (N779, N775, N456);
buf BUF1 (N780, N756);
and AND2 (N781, N776, N667);
xor XOR2 (N782, N779, N1);
xor XOR2 (N783, N729, N33);
nor NOR3 (N784, N780, N248, N320);
and AND4 (N785, N773, N257, N463, N388);
or OR4 (N786, N777, N461, N471, N202);
or OR4 (N787, N770, N13, N26, N558);
xor XOR2 (N788, N783, N251);
nand NAND3 (N789, N786, N66, N165);
xor XOR2 (N790, N781, N345);
and AND3 (N791, N789, N293, N225);
nor NOR3 (N792, N785, N571, N395);
and AND2 (N793, N778, N729);
and AND3 (N794, N782, N737, N191);
xor XOR2 (N795, N791, N197);
and AND3 (N796, N793, N160, N132);
xor XOR2 (N797, N787, N201);
nor NOR4 (N798, N795, N739, N112, N373);
or OR2 (N799, N790, N129);
and AND3 (N800, N788, N283, N647);
buf BUF1 (N801, N792);
nor NOR2 (N802, N769, N28);
buf BUF1 (N803, N798);
nand NAND3 (N804, N802, N710, N564);
nand NAND2 (N805, N799, N361);
buf BUF1 (N806, N784);
not NOT1 (N807, N794);
xor XOR2 (N808, N805, N8);
xor XOR2 (N809, N797, N597);
nand NAND4 (N810, N806, N29, N192, N699);
nand NAND2 (N811, N803, N175);
nor NOR4 (N812, N801, N682, N154, N628);
not NOT1 (N813, N766);
nor NOR4 (N814, N813, N447, N304, N803);
nand NAND4 (N815, N809, N101, N460, N683);
and AND2 (N816, N807, N775);
or OR3 (N817, N810, N409, N205);
or OR2 (N818, N811, N474);
nand NAND4 (N819, N808, N673, N345, N574);
and AND4 (N820, N812, N768, N511, N30);
not NOT1 (N821, N814);
nor NOR4 (N822, N800, N694, N201, N63);
not NOT1 (N823, N796);
not NOT1 (N824, N818);
nor NOR3 (N825, N804, N797, N535);
nand NAND4 (N826, N824, N312, N75, N427);
or OR3 (N827, N823, N738, N415);
not NOT1 (N828, N820);
xor XOR2 (N829, N827, N371);
xor XOR2 (N830, N828, N321);
nand NAND3 (N831, N829, N674, N388);
buf BUF1 (N832, N819);
nor NOR2 (N833, N822, N463);
buf BUF1 (N834, N833);
not NOT1 (N835, N826);
buf BUF1 (N836, N830);
buf BUF1 (N837, N816);
nand NAND4 (N838, N821, N395, N482, N566);
buf BUF1 (N839, N835);
xor XOR2 (N840, N836, N322);
nor NOR4 (N841, N834, N237, N473, N125);
xor XOR2 (N842, N840, N640);
not NOT1 (N843, N842);
nand NAND2 (N844, N838, N18);
xor XOR2 (N845, N831, N721);
and AND3 (N846, N844, N763, N807);
and AND2 (N847, N815, N670);
and AND2 (N848, N841, N727);
not NOT1 (N849, N825);
buf BUF1 (N850, N849);
buf BUF1 (N851, N837);
nand NAND2 (N852, N845, N187);
xor XOR2 (N853, N846, N352);
not NOT1 (N854, N843);
xor XOR2 (N855, N851, N83);
nor NOR4 (N856, N847, N854, N799, N852);
and AND4 (N857, N404, N359, N146, N750);
not NOT1 (N858, N84);
and AND2 (N859, N853, N498);
and AND3 (N860, N858, N727, N10);
nor NOR3 (N861, N857, N767, N488);
not NOT1 (N862, N861);
buf BUF1 (N863, N817);
xor XOR2 (N864, N860, N592);
buf BUF1 (N865, N856);
nand NAND3 (N866, N865, N176, N133);
buf BUF1 (N867, N866);
xor XOR2 (N868, N867, N126);
nor NOR3 (N869, N862, N53, N450);
xor XOR2 (N870, N869, N637);
or OR3 (N871, N839, N549, N316);
nand NAND4 (N872, N859, N864, N42, N505);
and AND4 (N873, N233, N844, N343, N33);
nor NOR3 (N874, N870, N63, N411);
not NOT1 (N875, N872);
and AND4 (N876, N855, N102, N565, N174);
nor NOR2 (N877, N875, N745);
nand NAND2 (N878, N848, N770);
buf BUF1 (N879, N871);
not NOT1 (N880, N874);
buf BUF1 (N881, N863);
nand NAND2 (N882, N832, N699);
or OR3 (N883, N879, N563, N367);
buf BUF1 (N884, N882);
not NOT1 (N885, N876);
not NOT1 (N886, N877);
nand NAND3 (N887, N886, N164, N613);
and AND3 (N888, N868, N92, N371);
and AND3 (N889, N873, N154, N63);
buf BUF1 (N890, N883);
buf BUF1 (N891, N884);
nor NOR3 (N892, N850, N204, N704);
or OR2 (N893, N880, N363);
and AND4 (N894, N891, N315, N143, N316);
and AND2 (N895, N890, N655);
not NOT1 (N896, N887);
nand NAND2 (N897, N894, N224);
xor XOR2 (N898, N895, N859);
or OR4 (N899, N889, N303, N3, N626);
nand NAND2 (N900, N896, N648);
nand NAND4 (N901, N892, N716, N803, N377);
xor XOR2 (N902, N881, N404);
and AND3 (N903, N900, N362, N291);
nor NOR4 (N904, N878, N712, N547, N177);
or OR3 (N905, N885, N848, N825);
nor NOR3 (N906, N903, N458, N657);
nand NAND3 (N907, N906, N118, N759);
nand NAND4 (N908, N893, N820, N47, N782);
not NOT1 (N909, N901);
or OR2 (N910, N902, N219);
buf BUF1 (N911, N898);
and AND4 (N912, N911, N590, N354, N618);
not NOT1 (N913, N905);
buf BUF1 (N914, N907);
and AND3 (N915, N888, N238, N240);
and AND3 (N916, N899, N236, N15);
or OR3 (N917, N897, N511, N383);
not NOT1 (N918, N917);
buf BUF1 (N919, N914);
nand NAND3 (N920, N908, N640, N489);
and AND4 (N921, N920, N305, N15, N415);
not NOT1 (N922, N919);
buf BUF1 (N923, N912);
nand NAND2 (N924, N909, N873);
and AND3 (N925, N924, N97, N145);
buf BUF1 (N926, N925);
buf BUF1 (N927, N923);
buf BUF1 (N928, N913);
xor XOR2 (N929, N927, N574);
or OR4 (N930, N922, N518, N248, N925);
or OR4 (N931, N926, N783, N314, N293);
not NOT1 (N932, N910);
and AND4 (N933, N931, N851, N432, N387);
or OR2 (N934, N916, N101);
nor NOR4 (N935, N929, N442, N812, N661);
nand NAND3 (N936, N933, N127, N269);
xor XOR2 (N937, N918, N415);
not NOT1 (N938, N932);
or OR4 (N939, N938, N198, N81, N891);
nor NOR2 (N940, N936, N85);
not NOT1 (N941, N928);
nor NOR3 (N942, N915, N211, N275);
nor NOR3 (N943, N941, N293, N196);
buf BUF1 (N944, N942);
not NOT1 (N945, N935);
nor NOR2 (N946, N945, N477);
not NOT1 (N947, N921);
and AND2 (N948, N904, N676);
or OR4 (N949, N947, N318, N934, N876);
nand NAND3 (N950, N324, N255, N485);
and AND2 (N951, N943, N835);
or OR3 (N952, N949, N685, N487);
nand NAND3 (N953, N951, N128, N27);
nand NAND2 (N954, N939, N217);
nor NOR2 (N955, N944, N672);
buf BUF1 (N956, N955);
xor XOR2 (N957, N940, N29);
xor XOR2 (N958, N950, N316);
or OR4 (N959, N958, N769, N594, N441);
nor NOR3 (N960, N930, N724, N753);
nand NAND2 (N961, N956, N602);
nand NAND2 (N962, N953, N277);
or OR3 (N963, N957, N626, N402);
nor NOR3 (N964, N960, N270, N216);
or OR4 (N965, N964, N612, N735, N936);
xor XOR2 (N966, N962, N835);
and AND4 (N967, N965, N654, N200, N165);
xor XOR2 (N968, N959, N834);
not NOT1 (N969, N954);
nand NAND3 (N970, N952, N6, N289);
or OR3 (N971, N963, N395, N101);
nand NAND3 (N972, N946, N627, N701);
nand NAND2 (N973, N968, N901);
buf BUF1 (N974, N970);
and AND3 (N975, N974, N197, N854);
xor XOR2 (N976, N966, N434);
xor XOR2 (N977, N967, N86);
nand NAND3 (N978, N976, N893, N221);
or OR3 (N979, N971, N85, N68);
xor XOR2 (N980, N937, N529);
not NOT1 (N981, N969);
nand NAND2 (N982, N972, N694);
and AND2 (N983, N948, N254);
not NOT1 (N984, N961);
or OR2 (N985, N975, N792);
nand NAND2 (N986, N981, N174);
buf BUF1 (N987, N984);
or OR3 (N988, N977, N838, N164);
or OR3 (N989, N986, N549, N739);
nor NOR3 (N990, N983, N810, N986);
nor NOR2 (N991, N988, N286);
or OR4 (N992, N973, N325, N399, N837);
nor NOR4 (N993, N978, N878, N711, N762);
or OR2 (N994, N987, N308);
xor XOR2 (N995, N980, N410);
nand NAND3 (N996, N991, N757, N793);
xor XOR2 (N997, N985, N397);
not NOT1 (N998, N982);
nand NAND3 (N999, N993, N1, N433);
buf BUF1 (N1000, N992);
nor NOR4 (N1001, N997, N436, N988, N609);
buf BUF1 (N1002, N995);
not NOT1 (N1003, N1002);
nand NAND2 (N1004, N979, N693);
not NOT1 (N1005, N994);
not NOT1 (N1006, N1005);
xor XOR2 (N1007, N998, N620);
nor NOR4 (N1008, N1000, N689, N647, N508);
buf BUF1 (N1009, N1007);
buf BUF1 (N1010, N1009);
and AND3 (N1011, N996, N822, N956);
buf BUF1 (N1012, N1003);
xor XOR2 (N1013, N1001, N413);
nor NOR4 (N1014, N1012, N297, N444, N980);
nor NOR3 (N1015, N1013, N411, N177);
or OR4 (N1016, N1011, N340, N604, N974);
xor XOR2 (N1017, N1010, N729);
nand NAND2 (N1018, N1004, N505);
not NOT1 (N1019, N1015);
and AND3 (N1020, N1018, N118, N672);
xor XOR2 (N1021, N1008, N414);
nor NOR3 (N1022, N1014, N992, N167);
xor XOR2 (N1023, N1016, N653);
xor XOR2 (N1024, N1019, N674);
or OR3 (N1025, N999, N545, N635);
xor XOR2 (N1026, N1023, N1020);
and AND4 (N1027, N424, N30, N221, N195);
nor NOR3 (N1028, N990, N877, N198);
not NOT1 (N1029, N1022);
nand NAND4 (N1030, N1026, N610, N717, N683);
or OR3 (N1031, N1017, N534, N111);
and AND2 (N1032, N1031, N601);
xor XOR2 (N1033, N989, N1000);
nand NAND3 (N1034, N1030, N279, N778);
buf BUF1 (N1035, N1021);
nor NOR2 (N1036, N1034, N206);
nor NOR2 (N1037, N1028, N424);
not NOT1 (N1038, N1036);
buf BUF1 (N1039, N1032);
nor NOR3 (N1040, N1024, N160, N316);
and AND4 (N1041, N1027, N1039, N133, N127);
buf BUF1 (N1042, N56);
not NOT1 (N1043, N1029);
nor NOR2 (N1044, N1037, N963);
and AND3 (N1045, N1040, N977, N973);
or OR4 (N1046, N1045, N115, N751, N672);
buf BUF1 (N1047, N1041);
nor NOR2 (N1048, N1046, N541);
or OR4 (N1049, N1042, N787, N71, N567);
nor NOR4 (N1050, N1044, N289, N466, N377);
and AND3 (N1051, N1047, N1005, N615);
nand NAND4 (N1052, N1006, N923, N315, N916);
nand NAND4 (N1053, N1050, N868, N798, N103);
not NOT1 (N1054, N1052);
not NOT1 (N1055, N1033);
and AND2 (N1056, N1035, N669);
or OR3 (N1057, N1051, N561, N991);
nor NOR2 (N1058, N1057, N702);
nor NOR2 (N1059, N1054, N102);
not NOT1 (N1060, N1059);
and AND3 (N1061, N1043, N769, N814);
nor NOR3 (N1062, N1056, N242, N870);
nor NOR4 (N1063, N1025, N316, N605, N279);
nor NOR4 (N1064, N1038, N341, N461, N76);
nor NOR3 (N1065, N1058, N322, N21);
and AND4 (N1066, N1049, N139, N411, N295);
xor XOR2 (N1067, N1065, N272);
nand NAND3 (N1068, N1067, N129, N318);
buf BUF1 (N1069, N1061);
not NOT1 (N1070, N1069);
or OR4 (N1071, N1063, N699, N114, N767);
xor XOR2 (N1072, N1068, N846);
buf BUF1 (N1073, N1072);
and AND4 (N1074, N1055, N346, N980, N910);
xor XOR2 (N1075, N1070, N566);
nand NAND4 (N1076, N1048, N608, N288, N79);
and AND2 (N1077, N1053, N30);
nand NAND2 (N1078, N1074, N207);
or OR4 (N1079, N1073, N713, N961, N1016);
xor XOR2 (N1080, N1071, N141);
buf BUF1 (N1081, N1066);
xor XOR2 (N1082, N1078, N758);
or OR2 (N1083, N1082, N546);
xor XOR2 (N1084, N1077, N822);
or OR3 (N1085, N1075, N126, N191);
xor XOR2 (N1086, N1079, N637);
buf BUF1 (N1087, N1076);
and AND3 (N1088, N1084, N707, N706);
nor NOR4 (N1089, N1062, N884, N654, N765);
and AND4 (N1090, N1089, N379, N984, N457);
not NOT1 (N1091, N1085);
nand NAND2 (N1092, N1083, N829);
nor NOR4 (N1093, N1081, N471, N535, N1032);
nand NAND4 (N1094, N1091, N1068, N413, N787);
nor NOR4 (N1095, N1064, N101, N745, N321);
xor XOR2 (N1096, N1088, N344);
nor NOR4 (N1097, N1094, N605, N881, N825);
nor NOR4 (N1098, N1092, N344, N1058, N827);
buf BUF1 (N1099, N1096);
xor XOR2 (N1100, N1098, N681);
nand NAND3 (N1101, N1090, N1076, N475);
nand NAND3 (N1102, N1060, N516, N885);
or OR3 (N1103, N1101, N536, N730);
buf BUF1 (N1104, N1087);
nand NAND2 (N1105, N1102, N657);
not NOT1 (N1106, N1103);
nor NOR3 (N1107, N1099, N545, N936);
nand NAND2 (N1108, N1097, N160);
nand NAND4 (N1109, N1080, N1012, N789, N897);
or OR3 (N1110, N1093, N528, N885);
and AND3 (N1111, N1106, N909, N904);
or OR2 (N1112, N1109, N298);
or OR3 (N1113, N1110, N935, N139);
or OR2 (N1114, N1113, N43);
and AND4 (N1115, N1111, N601, N586, N504);
and AND3 (N1116, N1115, N551, N100);
and AND4 (N1117, N1104, N1058, N657, N395);
or OR3 (N1118, N1105, N1031, N770);
xor XOR2 (N1119, N1114, N958);
not NOT1 (N1120, N1117);
nand NAND3 (N1121, N1095, N200, N82);
nand NAND4 (N1122, N1120, N464, N388, N348);
nor NOR4 (N1123, N1118, N313, N164, N502);
and AND2 (N1124, N1086, N224);
nor NOR4 (N1125, N1119, N498, N40, N797);
and AND2 (N1126, N1107, N592);
buf BUF1 (N1127, N1124);
or OR4 (N1128, N1125, N731, N365, N265);
not NOT1 (N1129, N1116);
not NOT1 (N1130, N1126);
and AND4 (N1131, N1128, N401, N766, N1082);
or OR4 (N1132, N1100, N162, N1100, N811);
xor XOR2 (N1133, N1129, N286);
xor XOR2 (N1134, N1131, N735);
xor XOR2 (N1135, N1123, N157);
buf BUF1 (N1136, N1135);
and AND3 (N1137, N1133, N155, N659);
nor NOR4 (N1138, N1136, N557, N502, N576);
nand NAND2 (N1139, N1137, N838);
nand NAND4 (N1140, N1108, N470, N811, N841);
buf BUF1 (N1141, N1127);
xor XOR2 (N1142, N1112, N479);
not NOT1 (N1143, N1141);
xor XOR2 (N1144, N1134, N253);
not NOT1 (N1145, N1132);
and AND2 (N1146, N1144, N627);
and AND2 (N1147, N1139, N392);
xor XOR2 (N1148, N1140, N892);
and AND4 (N1149, N1145, N272, N575, N343);
xor XOR2 (N1150, N1148, N954);
or OR2 (N1151, N1138, N614);
not NOT1 (N1152, N1143);
nand NAND4 (N1153, N1121, N166, N792, N190);
or OR4 (N1154, N1130, N37, N819, N202);
nand NAND2 (N1155, N1142, N32);
nand NAND4 (N1156, N1122, N781, N22, N348);
xor XOR2 (N1157, N1153, N85);
nand NAND4 (N1158, N1154, N790, N472, N152);
xor XOR2 (N1159, N1158, N1043);
not NOT1 (N1160, N1156);
nand NAND3 (N1161, N1146, N769, N317);
buf BUF1 (N1162, N1149);
nand NAND2 (N1163, N1159, N606);
xor XOR2 (N1164, N1147, N539);
and AND3 (N1165, N1157, N15, N307);
or OR4 (N1166, N1160, N964, N113, N355);
or OR4 (N1167, N1150, N282, N292, N740);
buf BUF1 (N1168, N1155);
xor XOR2 (N1169, N1152, N180);
nand NAND2 (N1170, N1162, N1047);
buf BUF1 (N1171, N1170);
or OR3 (N1172, N1169, N195, N392);
buf BUF1 (N1173, N1163);
or OR2 (N1174, N1161, N755);
or OR2 (N1175, N1174, N595);
nor NOR2 (N1176, N1165, N702);
xor XOR2 (N1177, N1164, N907);
buf BUF1 (N1178, N1171);
or OR4 (N1179, N1172, N1082, N647, N1069);
and AND4 (N1180, N1177, N380, N1100, N759);
buf BUF1 (N1181, N1180);
buf BUF1 (N1182, N1151);
or OR3 (N1183, N1167, N323, N954);
xor XOR2 (N1184, N1182, N81);
and AND3 (N1185, N1168, N141, N793);
xor XOR2 (N1186, N1183, N2);
and AND2 (N1187, N1175, N1135);
buf BUF1 (N1188, N1184);
nand NAND3 (N1189, N1173, N562, N127);
nor NOR2 (N1190, N1188, N125);
not NOT1 (N1191, N1185);
not NOT1 (N1192, N1187);
xor XOR2 (N1193, N1181, N1189);
buf BUF1 (N1194, N334);
not NOT1 (N1195, N1179);
or OR2 (N1196, N1191, N1093);
nand NAND4 (N1197, N1186, N218, N1187, N1077);
nand NAND3 (N1198, N1196, N591, N575);
and AND4 (N1199, N1178, N395, N356, N563);
not NOT1 (N1200, N1194);
buf BUF1 (N1201, N1200);
or OR2 (N1202, N1195, N493);
nor NOR2 (N1203, N1201, N306);
xor XOR2 (N1204, N1176, N529);
buf BUF1 (N1205, N1199);
and AND3 (N1206, N1202, N376, N1030);
and AND3 (N1207, N1192, N1012, N787);
and AND3 (N1208, N1193, N916, N735);
or OR3 (N1209, N1206, N1050, N389);
nand NAND4 (N1210, N1204, N481, N241, N1050);
nor NOR2 (N1211, N1197, N206);
nor NOR3 (N1212, N1205, N271, N920);
and AND4 (N1213, N1211, N81, N678, N19);
or OR4 (N1214, N1166, N62, N761, N898);
or OR2 (N1215, N1212, N1178);
and AND4 (N1216, N1207, N964, N307, N1037);
or OR3 (N1217, N1216, N519, N1132);
or OR2 (N1218, N1217, N549);
nand NAND4 (N1219, N1215, N843, N163, N217);
and AND3 (N1220, N1209, N565, N354);
nor NOR2 (N1221, N1220, N661);
not NOT1 (N1222, N1214);
or OR4 (N1223, N1219, N661, N902, N1155);
not NOT1 (N1224, N1210);
and AND3 (N1225, N1203, N764, N1124);
not NOT1 (N1226, N1225);
nor NOR4 (N1227, N1223, N214, N158, N568);
not NOT1 (N1228, N1221);
buf BUF1 (N1229, N1228);
buf BUF1 (N1230, N1190);
xor XOR2 (N1231, N1227, N1099);
nor NOR3 (N1232, N1226, N145, N440);
not NOT1 (N1233, N1224);
nor NOR4 (N1234, N1233, N337, N915, N1062);
xor XOR2 (N1235, N1213, N1044);
or OR3 (N1236, N1235, N398, N615);
not NOT1 (N1237, N1231);
nand NAND2 (N1238, N1237, N1098);
nand NAND4 (N1239, N1198, N719, N10, N420);
nor NOR4 (N1240, N1232, N176, N683, N1171);
not NOT1 (N1241, N1239);
xor XOR2 (N1242, N1234, N441);
and AND4 (N1243, N1238, N240, N199, N571);
nand NAND4 (N1244, N1230, N1207, N844, N620);
and AND2 (N1245, N1208, N1163);
or OR4 (N1246, N1218, N646, N599, N800);
nand NAND3 (N1247, N1243, N874, N457);
not NOT1 (N1248, N1244);
and AND2 (N1249, N1222, N268);
nor NOR4 (N1250, N1240, N1244, N1009, N144);
not NOT1 (N1251, N1248);
not NOT1 (N1252, N1249);
or OR2 (N1253, N1246, N772);
buf BUF1 (N1254, N1236);
nor NOR3 (N1255, N1252, N33, N814);
not NOT1 (N1256, N1242);
nand NAND2 (N1257, N1241, N420);
buf BUF1 (N1258, N1229);
and AND3 (N1259, N1251, N753, N330);
or OR4 (N1260, N1255, N509, N299, N1199);
nand NAND2 (N1261, N1253, N856);
xor XOR2 (N1262, N1245, N1148);
not NOT1 (N1263, N1262);
buf BUF1 (N1264, N1261);
buf BUF1 (N1265, N1259);
not NOT1 (N1266, N1263);
and AND4 (N1267, N1260, N1027, N1000, N1068);
buf BUF1 (N1268, N1247);
or OR2 (N1269, N1250, N535);
buf BUF1 (N1270, N1256);
nand NAND3 (N1271, N1267, N618, N305);
or OR2 (N1272, N1266, N808);
and AND3 (N1273, N1258, N202, N1112);
and AND2 (N1274, N1272, N1241);
nor NOR4 (N1275, N1274, N86, N1216, N800);
nor NOR3 (N1276, N1254, N391, N296);
nor NOR3 (N1277, N1275, N703, N431);
not NOT1 (N1278, N1271);
or OR3 (N1279, N1269, N1125, N1131);
xor XOR2 (N1280, N1264, N1185);
or OR4 (N1281, N1265, N576, N573, N904);
or OR4 (N1282, N1268, N175, N988, N348);
not NOT1 (N1283, N1280);
nand NAND2 (N1284, N1273, N946);
buf BUF1 (N1285, N1276);
and AND4 (N1286, N1279, N406, N757, N538);
xor XOR2 (N1287, N1284, N1003);
nand NAND2 (N1288, N1283, N610);
xor XOR2 (N1289, N1282, N28);
nor NOR2 (N1290, N1270, N1102);
or OR4 (N1291, N1288, N952, N762, N609);
nand NAND3 (N1292, N1257, N193, N857);
and AND2 (N1293, N1291, N828);
xor XOR2 (N1294, N1278, N919);
nor NOR4 (N1295, N1293, N238, N982, N504);
and AND4 (N1296, N1287, N387, N350, N350);
nor NOR4 (N1297, N1281, N1265, N303, N136);
nand NAND3 (N1298, N1286, N125, N793);
and AND3 (N1299, N1290, N754, N242);
buf BUF1 (N1300, N1295);
buf BUF1 (N1301, N1300);
and AND4 (N1302, N1296, N686, N1105, N861);
nand NAND4 (N1303, N1302, N39, N432, N610);
nand NAND4 (N1304, N1298, N1092, N961, N351);
nor NOR2 (N1305, N1285, N775);
not NOT1 (N1306, N1294);
nor NOR2 (N1307, N1299, N379);
xor XOR2 (N1308, N1277, N42);
nand NAND2 (N1309, N1297, N1015);
nor NOR2 (N1310, N1309, N912);
nor NOR2 (N1311, N1308, N715);
buf BUF1 (N1312, N1292);
and AND4 (N1313, N1304, N785, N256, N564);
xor XOR2 (N1314, N1305, N367);
or OR4 (N1315, N1289, N238, N639, N487);
nor NOR3 (N1316, N1315, N770, N1015);
or OR4 (N1317, N1306, N324, N679, N910);
or OR4 (N1318, N1310, N508, N103, N1083);
and AND4 (N1319, N1303, N394, N191, N298);
not NOT1 (N1320, N1317);
buf BUF1 (N1321, N1311);
nand NAND4 (N1322, N1318, N544, N444, N208);
not NOT1 (N1323, N1319);
nor NOR4 (N1324, N1322, N227, N973, N580);
and AND2 (N1325, N1323, N1230);
nand NAND4 (N1326, N1316, N480, N997, N92);
not NOT1 (N1327, N1312);
and AND2 (N1328, N1325, N772);
and AND3 (N1329, N1327, N1026, N576);
and AND4 (N1330, N1307, N717, N386, N806);
nor NOR4 (N1331, N1301, N925, N602, N512);
not NOT1 (N1332, N1328);
xor XOR2 (N1333, N1320, N1247);
and AND2 (N1334, N1313, N1210);
buf BUF1 (N1335, N1324);
and AND4 (N1336, N1314, N1089, N1274, N478);
or OR4 (N1337, N1333, N388, N545, N605);
nand NAND4 (N1338, N1332, N108, N1201, N160);
nor NOR4 (N1339, N1329, N1049, N282, N207);
not NOT1 (N1340, N1331);
buf BUF1 (N1341, N1339);
not NOT1 (N1342, N1330);
nor NOR4 (N1343, N1321, N1265, N472, N527);
xor XOR2 (N1344, N1342, N1128);
and AND2 (N1345, N1338, N952);
not NOT1 (N1346, N1336);
and AND3 (N1347, N1340, N19, N202);
or OR2 (N1348, N1345, N500);
or OR2 (N1349, N1343, N408);
xor XOR2 (N1350, N1347, N627);
not NOT1 (N1351, N1326);
and AND3 (N1352, N1334, N780, N531);
nand NAND3 (N1353, N1350, N1098, N344);
nand NAND2 (N1354, N1349, N1303);
not NOT1 (N1355, N1352);
xor XOR2 (N1356, N1337, N603);
not NOT1 (N1357, N1356);
nand NAND3 (N1358, N1335, N1200, N333);
not NOT1 (N1359, N1357);
and AND3 (N1360, N1351, N212, N30);
xor XOR2 (N1361, N1346, N223);
or OR2 (N1362, N1353, N1087);
and AND4 (N1363, N1361, N1208, N540, N598);
and AND4 (N1364, N1344, N979, N1177, N585);
xor XOR2 (N1365, N1363, N805);
or OR3 (N1366, N1341, N1003, N1258);
or OR2 (N1367, N1355, N1086);
buf BUF1 (N1368, N1367);
nand NAND3 (N1369, N1354, N1246, N710);
xor XOR2 (N1370, N1364, N531);
not NOT1 (N1371, N1365);
nand NAND2 (N1372, N1362, N1173);
nand NAND4 (N1373, N1358, N244, N175, N616);
buf BUF1 (N1374, N1348);
and AND2 (N1375, N1360, N425);
not NOT1 (N1376, N1370);
or OR4 (N1377, N1371, N1149, N354, N429);
buf BUF1 (N1378, N1376);
and AND3 (N1379, N1378, N1308, N581);
buf BUF1 (N1380, N1366);
not NOT1 (N1381, N1374);
xor XOR2 (N1382, N1379, N667);
and AND3 (N1383, N1380, N1243, N1363);
xor XOR2 (N1384, N1383, N428);
or OR2 (N1385, N1369, N1347);
and AND4 (N1386, N1382, N1101, N758, N800);
nand NAND4 (N1387, N1381, N1044, N623, N1228);
nor NOR4 (N1388, N1377, N1256, N194, N1336);
nand NAND4 (N1389, N1386, N79, N284, N137);
not NOT1 (N1390, N1368);
buf BUF1 (N1391, N1387);
buf BUF1 (N1392, N1390);
xor XOR2 (N1393, N1388, N1186);
buf BUF1 (N1394, N1373);
or OR3 (N1395, N1394, N314, N149);
not NOT1 (N1396, N1372);
and AND4 (N1397, N1393, N160, N885, N875);
and AND4 (N1398, N1385, N575, N282, N1150);
and AND3 (N1399, N1359, N884, N1126);
buf BUF1 (N1400, N1391);
xor XOR2 (N1401, N1389, N44);
buf BUF1 (N1402, N1398);
nand NAND3 (N1403, N1395, N498, N450);
or OR4 (N1404, N1401, N823, N1389, N1304);
xor XOR2 (N1405, N1399, N377);
xor XOR2 (N1406, N1400, N40);
nand NAND4 (N1407, N1397, N1036, N296, N90);
buf BUF1 (N1408, N1375);
or OR3 (N1409, N1407, N159, N333);
and AND3 (N1410, N1402, N900, N1056);
nand NAND2 (N1411, N1409, N73);
xor XOR2 (N1412, N1396, N390);
or OR3 (N1413, N1410, N1368, N1410);
or OR2 (N1414, N1411, N796);
nand NAND3 (N1415, N1408, N68, N675);
nand NAND3 (N1416, N1412, N1153, N642);
xor XOR2 (N1417, N1405, N994);
xor XOR2 (N1418, N1406, N495);
and AND2 (N1419, N1418, N1023);
not NOT1 (N1420, N1403);
and AND4 (N1421, N1415, N994, N365, N1358);
nor NOR3 (N1422, N1416, N1012, N766);
xor XOR2 (N1423, N1392, N973);
not NOT1 (N1424, N1417);
nor NOR3 (N1425, N1422, N805, N839);
nor NOR2 (N1426, N1424, N384);
nor NOR4 (N1427, N1384, N280, N1398, N553);
xor XOR2 (N1428, N1423, N1206);
buf BUF1 (N1429, N1427);
or OR4 (N1430, N1428, N1138, N188, N840);
buf BUF1 (N1431, N1413);
xor XOR2 (N1432, N1430, N1404);
nand NAND2 (N1433, N112, N312);
and AND2 (N1434, N1419, N500);
not NOT1 (N1435, N1429);
nand NAND3 (N1436, N1433, N894, N1327);
buf BUF1 (N1437, N1421);
nand NAND3 (N1438, N1414, N1057, N433);
or OR3 (N1439, N1434, N914, N562);
nor NOR4 (N1440, N1437, N569, N657, N1267);
nor NOR3 (N1441, N1438, N69, N595);
buf BUF1 (N1442, N1441);
buf BUF1 (N1443, N1435);
xor XOR2 (N1444, N1432, N1228);
xor XOR2 (N1445, N1431, N788);
not NOT1 (N1446, N1436);
xor XOR2 (N1447, N1444, N417);
nor NOR4 (N1448, N1426, N203, N208, N1140);
nand NAND3 (N1449, N1448, N81, N246);
nand NAND3 (N1450, N1445, N627, N824);
nor NOR4 (N1451, N1450, N1090, N635, N1345);
or OR2 (N1452, N1440, N1182);
nand NAND3 (N1453, N1449, N683, N1313);
and AND3 (N1454, N1447, N547, N973);
nand NAND4 (N1455, N1451, N452, N1349, N1320);
buf BUF1 (N1456, N1443);
and AND2 (N1457, N1456, N1005);
nand NAND2 (N1458, N1453, N977);
not NOT1 (N1459, N1442);
not NOT1 (N1460, N1455);
nor NOR2 (N1461, N1446, N523);
nand NAND2 (N1462, N1457, N640);
and AND4 (N1463, N1460, N689, N496, N1223);
buf BUF1 (N1464, N1420);
buf BUF1 (N1465, N1458);
nand NAND2 (N1466, N1425, N1182);
or OR4 (N1467, N1465, N716, N45, N1229);
or OR2 (N1468, N1461, N337);
nor NOR3 (N1469, N1462, N1186, N1466);
or OR4 (N1470, N1255, N832, N970, N259);
nand NAND3 (N1471, N1464, N720, N316);
buf BUF1 (N1472, N1463);
nand NAND3 (N1473, N1471, N924, N165);
not NOT1 (N1474, N1459);
xor XOR2 (N1475, N1452, N372);
not NOT1 (N1476, N1468);
nand NAND4 (N1477, N1473, N1198, N935, N172);
buf BUF1 (N1478, N1476);
xor XOR2 (N1479, N1469, N51);
nor NOR2 (N1480, N1470, N1015);
buf BUF1 (N1481, N1472);
and AND2 (N1482, N1480, N62);
not NOT1 (N1483, N1475);
xor XOR2 (N1484, N1483, N727);
and AND3 (N1485, N1467, N272, N945);
and AND2 (N1486, N1477, N1166);
not NOT1 (N1487, N1478);
nor NOR4 (N1488, N1486, N1444, N1333, N856);
and AND4 (N1489, N1488, N799, N1247, N212);
buf BUF1 (N1490, N1481);
nand NAND4 (N1491, N1479, N1296, N935, N940);
not NOT1 (N1492, N1474);
and AND3 (N1493, N1485, N1397, N1449);
buf BUF1 (N1494, N1487);
buf BUF1 (N1495, N1454);
buf BUF1 (N1496, N1491);
nor NOR4 (N1497, N1489, N418, N660, N419);
and AND2 (N1498, N1492, N25);
nor NOR3 (N1499, N1484, N748, N1424);
xor XOR2 (N1500, N1494, N350);
and AND3 (N1501, N1500, N917, N1267);
not NOT1 (N1502, N1499);
buf BUF1 (N1503, N1495);
not NOT1 (N1504, N1493);
xor XOR2 (N1505, N1504, N751);
nor NOR4 (N1506, N1496, N579, N456, N286);
nor NOR3 (N1507, N1505, N967, N156);
buf BUF1 (N1508, N1507);
not NOT1 (N1509, N1501);
or OR4 (N1510, N1439, N1001, N3, N188);
buf BUF1 (N1511, N1509);
nor NOR3 (N1512, N1497, N90, N1006);
nand NAND2 (N1513, N1508, N1492);
or OR3 (N1514, N1510, N1233, N190);
and AND3 (N1515, N1498, N1467, N941);
buf BUF1 (N1516, N1482);
xor XOR2 (N1517, N1511, N972);
xor XOR2 (N1518, N1503, N177);
xor XOR2 (N1519, N1502, N1065);
buf BUF1 (N1520, N1519);
xor XOR2 (N1521, N1514, N322);
not NOT1 (N1522, N1490);
nand NAND3 (N1523, N1515, N217, N675);
nor NOR4 (N1524, N1522, N863, N822, N737);
nor NOR2 (N1525, N1521, N24);
or OR3 (N1526, N1517, N93, N579);
or OR3 (N1527, N1516, N861, N1261);
nor NOR4 (N1528, N1512, N710, N960, N1449);
not NOT1 (N1529, N1518);
nand NAND2 (N1530, N1529, N612);
nand NAND4 (N1531, N1525, N1022, N709, N545);
or OR3 (N1532, N1524, N794, N1084);
nand NAND2 (N1533, N1513, N917);
buf BUF1 (N1534, N1528);
not NOT1 (N1535, N1533);
or OR4 (N1536, N1532, N769, N654, N420);
and AND2 (N1537, N1530, N317);
not NOT1 (N1538, N1526);
nor NOR3 (N1539, N1523, N305, N398);
nor NOR3 (N1540, N1538, N479, N491);
not NOT1 (N1541, N1537);
or OR4 (N1542, N1527, N20, N1085, N203);
and AND4 (N1543, N1535, N648, N850, N736);
xor XOR2 (N1544, N1543, N34);
buf BUF1 (N1545, N1531);
xor XOR2 (N1546, N1541, N358);
xor XOR2 (N1547, N1542, N907);
not NOT1 (N1548, N1520);
nand NAND3 (N1549, N1540, N1245, N321);
nand NAND4 (N1550, N1536, N1062, N577, N1200);
not NOT1 (N1551, N1539);
and AND4 (N1552, N1506, N32, N1439, N1338);
not NOT1 (N1553, N1549);
not NOT1 (N1554, N1553);
and AND4 (N1555, N1551, N934, N387, N1291);
nand NAND2 (N1556, N1546, N677);
xor XOR2 (N1557, N1547, N1179);
xor XOR2 (N1558, N1557, N513);
nor NOR4 (N1559, N1554, N978, N776, N471);
or OR2 (N1560, N1555, N504);
nor NOR3 (N1561, N1558, N252, N233);
nor NOR2 (N1562, N1552, N637);
nor NOR2 (N1563, N1562, N433);
nand NAND4 (N1564, N1560, N192, N891, N487);
nand NAND2 (N1565, N1544, N1091);
and AND3 (N1566, N1545, N486, N1424);
not NOT1 (N1567, N1534);
or OR2 (N1568, N1565, N406);
or OR2 (N1569, N1568, N202);
xor XOR2 (N1570, N1564, N46);
not NOT1 (N1571, N1569);
or OR2 (N1572, N1559, N321);
or OR3 (N1573, N1571, N160, N1536);
nand NAND3 (N1574, N1556, N358, N467);
xor XOR2 (N1575, N1548, N372);
not NOT1 (N1576, N1550);
nand NAND2 (N1577, N1561, N20);
buf BUF1 (N1578, N1570);
xor XOR2 (N1579, N1566, N508);
buf BUF1 (N1580, N1575);
nand NAND4 (N1581, N1574, N730, N197, N527);
not NOT1 (N1582, N1581);
not NOT1 (N1583, N1580);
xor XOR2 (N1584, N1576, N1000);
nand NAND3 (N1585, N1578, N884, N797);
buf BUF1 (N1586, N1577);
or OR2 (N1587, N1563, N83);
nand NAND3 (N1588, N1572, N634, N290);
nor NOR3 (N1589, N1586, N240, N1495);
or OR3 (N1590, N1582, N1351, N1420);
nor NOR2 (N1591, N1583, N768);
nand NAND3 (N1592, N1589, N1491, N481);
or OR4 (N1593, N1591, N572, N601, N1272);
nor NOR3 (N1594, N1587, N728, N440);
xor XOR2 (N1595, N1584, N604);
not NOT1 (N1596, N1588);
xor XOR2 (N1597, N1593, N186);
nor NOR4 (N1598, N1579, N601, N821, N39);
or OR2 (N1599, N1594, N1102);
or OR2 (N1600, N1595, N1470);
xor XOR2 (N1601, N1567, N1086);
nor NOR2 (N1602, N1573, N168);
buf BUF1 (N1603, N1601);
buf BUF1 (N1604, N1585);
nor NOR2 (N1605, N1596, N1537);
xor XOR2 (N1606, N1598, N275);
or OR3 (N1607, N1602, N739, N1300);
and AND2 (N1608, N1604, N1230);
or OR4 (N1609, N1605, N1072, N408, N1290);
not NOT1 (N1610, N1608);
nand NAND4 (N1611, N1592, N1232, N678, N305);
or OR3 (N1612, N1606, N43, N145);
or OR4 (N1613, N1603, N475, N1032, N766);
nand NAND2 (N1614, N1609, N361);
nor NOR3 (N1615, N1612, N892, N1287);
and AND2 (N1616, N1600, N1560);
or OR2 (N1617, N1611, N1337);
and AND3 (N1618, N1590, N1211, N311);
buf BUF1 (N1619, N1597);
nor NOR3 (N1620, N1607, N18, N1588);
and AND2 (N1621, N1616, N1259);
nor NOR4 (N1622, N1619, N568, N289, N493);
or OR3 (N1623, N1610, N1603, N1021);
endmodule