// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N299,N302,N296,N276,N308,N304,N307,N305,N309,N310;

buf BUF1 (N11, N1);
or OR4 (N12, N1, N11, N6, N5);
nor NOR4 (N13, N10, N12, N9, N8);
and AND3 (N14, N5, N9, N11);
or OR3 (N15, N2, N6, N2);
buf BUF1 (N16, N12);
buf BUF1 (N17, N2);
or OR4 (N18, N1, N2, N14, N9);
or OR3 (N19, N16, N9, N11);
nand NAND3 (N20, N14, N9, N14);
nor NOR2 (N21, N12, N13);
nor NOR3 (N22, N14, N11, N20);
and AND4 (N23, N22, N20, N19, N20);
not NOT1 (N24, N22);
nor NOR4 (N25, N5, N9, N4, N21);
nand NAND4 (N26, N19, N16, N6, N13);
nor NOR2 (N27, N24, N20);
xor XOR2 (N28, N15, N20);
not NOT1 (N29, N8);
or OR4 (N30, N22, N24, N19, N21);
xor XOR2 (N31, N28, N27);
buf BUF1 (N32, N20);
buf BUF1 (N33, N32);
buf BUF1 (N34, N19);
nor NOR4 (N35, N26, N27, N8, N23);
or OR3 (N36, N25, N33, N9);
nor NOR2 (N37, N21, N5);
and AND2 (N38, N23, N23);
buf BUF1 (N39, N18);
xor XOR2 (N40, N34, N5);
nand NAND2 (N41, N37, N15);
or OR3 (N42, N40, N28, N33);
buf BUF1 (N43, N30);
nor NOR2 (N44, N31, N35);
not NOT1 (N45, N27);
not NOT1 (N46, N39);
nand NAND2 (N47, N46, N40);
nor NOR3 (N48, N42, N9, N29);
nor NOR3 (N49, N21, N21, N3);
nand NAND4 (N50, N49, N5, N10, N24);
not NOT1 (N51, N17);
not NOT1 (N52, N50);
xor XOR2 (N53, N38, N3);
xor XOR2 (N54, N45, N11);
and AND3 (N55, N47, N22, N31);
or OR3 (N56, N43, N54, N47);
xor XOR2 (N57, N22, N34);
or OR3 (N58, N48, N24, N38);
xor XOR2 (N59, N44, N14);
nand NAND4 (N60, N51, N5, N9, N7);
xor XOR2 (N61, N53, N2);
not NOT1 (N62, N61);
or OR4 (N63, N55, N10, N53, N42);
not NOT1 (N64, N58);
and AND4 (N65, N63, N56, N33, N17);
or OR2 (N66, N13, N26);
nor NOR2 (N67, N66, N41);
buf BUF1 (N68, N29);
buf BUF1 (N69, N52);
buf BUF1 (N70, N64);
nor NOR4 (N71, N65, N34, N14, N40);
or OR2 (N72, N59, N41);
and AND2 (N73, N62, N40);
and AND3 (N74, N60, N52, N40);
nor NOR2 (N75, N36, N20);
not NOT1 (N76, N75);
not NOT1 (N77, N70);
nand NAND3 (N78, N69, N66, N60);
and AND2 (N79, N67, N14);
buf BUF1 (N80, N79);
xor XOR2 (N81, N80, N50);
xor XOR2 (N82, N78, N14);
and AND3 (N83, N76, N42, N72);
or OR4 (N84, N81, N71, N30, N47);
not NOT1 (N85, N47);
nor NOR2 (N86, N24, N38);
or OR4 (N87, N74, N11, N16, N54);
nor NOR3 (N88, N83, N22, N86);
and AND2 (N89, N81, N73);
or OR2 (N90, N41, N43);
buf BUF1 (N91, N85);
and AND4 (N92, N57, N86, N77, N72);
and AND2 (N93, N46, N20);
and AND3 (N94, N88, N15, N59);
nand NAND3 (N95, N82, N62, N34);
buf BUF1 (N96, N87);
nand NAND2 (N97, N95, N42);
nor NOR4 (N98, N93, N22, N46, N29);
nand NAND2 (N99, N98, N32);
nor NOR4 (N100, N96, N60, N91, N91);
nand NAND2 (N101, N82, N89);
not NOT1 (N102, N57);
buf BUF1 (N103, N97);
and AND3 (N104, N103, N89, N18);
buf BUF1 (N105, N68);
or OR4 (N106, N84, N73, N44, N15);
nand NAND2 (N107, N105, N14);
and AND3 (N108, N106, N96, N59);
or OR4 (N109, N92, N47, N84, N60);
buf BUF1 (N110, N100);
or OR4 (N111, N108, N56, N99, N29);
or OR2 (N112, N54, N19);
nand NAND4 (N113, N109, N98, N91, N42);
xor XOR2 (N114, N107, N52);
and AND3 (N115, N113, N16, N23);
nor NOR4 (N116, N104, N87, N111, N43);
and AND2 (N117, N28, N75);
nand NAND3 (N118, N94, N82, N78);
xor XOR2 (N119, N118, N114);
nor NOR2 (N120, N104, N38);
nor NOR3 (N121, N120, N29, N34);
nor NOR2 (N122, N115, N116);
xor XOR2 (N123, N2, N60);
not NOT1 (N124, N110);
buf BUF1 (N125, N90);
nand NAND4 (N126, N122, N117, N95, N31);
nand NAND2 (N127, N5, N12);
or OR3 (N128, N123, N46, N81);
nand NAND3 (N129, N112, N18, N120);
nor NOR4 (N130, N102, N15, N80, N18);
or OR2 (N131, N126, N23);
nor NOR3 (N132, N129, N68, N72);
xor XOR2 (N133, N101, N123);
not NOT1 (N134, N128);
xor XOR2 (N135, N133, N61);
nor NOR4 (N136, N130, N42, N75, N9);
not NOT1 (N137, N124);
xor XOR2 (N138, N132, N8);
or OR3 (N139, N125, N21, N92);
xor XOR2 (N140, N137, N126);
or OR2 (N141, N131, N11);
nor NOR3 (N142, N140, N53, N133);
or OR3 (N143, N127, N41, N116);
not NOT1 (N144, N143);
nor NOR4 (N145, N141, N94, N66, N27);
and AND3 (N146, N136, N36, N94);
or OR2 (N147, N119, N128);
xor XOR2 (N148, N147, N45);
nand NAND2 (N149, N148, N51);
xor XOR2 (N150, N121, N148);
nor NOR3 (N151, N138, N36, N8);
and AND4 (N152, N149, N82, N83, N76);
not NOT1 (N153, N135);
nand NAND3 (N154, N152, N46, N42);
xor XOR2 (N155, N145, N95);
not NOT1 (N156, N139);
and AND2 (N157, N153, N116);
buf BUF1 (N158, N142);
not NOT1 (N159, N150);
buf BUF1 (N160, N144);
and AND3 (N161, N160, N54, N156);
nand NAND3 (N162, N119, N62, N85);
buf BUF1 (N163, N151);
not NOT1 (N164, N155);
or OR4 (N165, N154, N136, N28, N124);
nor NOR4 (N166, N157, N133, N50, N109);
nand NAND4 (N167, N146, N87, N87, N116);
xor XOR2 (N168, N158, N129);
nor NOR3 (N169, N159, N97, N19);
buf BUF1 (N170, N134);
not NOT1 (N171, N164);
nand NAND2 (N172, N165, N82);
or OR2 (N173, N161, N123);
and AND3 (N174, N163, N84, N61);
not NOT1 (N175, N171);
or OR3 (N176, N170, N61, N64);
nand NAND4 (N177, N174, N102, N105, N26);
or OR2 (N178, N177, N174);
or OR4 (N179, N166, N173, N171, N95);
xor XOR2 (N180, N171, N141);
buf BUF1 (N181, N180);
buf BUF1 (N182, N176);
buf BUF1 (N183, N182);
xor XOR2 (N184, N168, N44);
nor NOR2 (N185, N183, N183);
xor XOR2 (N186, N172, N143);
xor XOR2 (N187, N169, N133);
buf BUF1 (N188, N167);
not NOT1 (N189, N188);
xor XOR2 (N190, N186, N23);
xor XOR2 (N191, N190, N13);
nand NAND2 (N192, N189, N59);
not NOT1 (N193, N181);
not NOT1 (N194, N179);
nand NAND3 (N195, N192, N19, N115);
xor XOR2 (N196, N162, N113);
not NOT1 (N197, N187);
not NOT1 (N198, N191);
buf BUF1 (N199, N196);
buf BUF1 (N200, N197);
not NOT1 (N201, N194);
nand NAND3 (N202, N178, N82, N95);
buf BUF1 (N203, N199);
and AND4 (N204, N195, N68, N202, N55);
nand NAND4 (N205, N103, N122, N11, N146);
nand NAND2 (N206, N198, N191);
nand NAND2 (N207, N184, N156);
and AND4 (N208, N205, N143, N112, N74);
buf BUF1 (N209, N204);
nand NAND3 (N210, N200, N78, N22);
xor XOR2 (N211, N209, N110);
and AND3 (N212, N185, N191, N54);
not NOT1 (N213, N193);
xor XOR2 (N214, N213, N146);
nor NOR3 (N215, N210, N74, N166);
nand NAND4 (N216, N214, N121, N152, N143);
buf BUF1 (N217, N212);
nor NOR4 (N218, N208, N38, N118, N97);
or OR2 (N219, N206, N10);
and AND3 (N220, N219, N196, N34);
or OR3 (N221, N216, N36, N65);
nor NOR4 (N222, N175, N60, N187, N95);
and AND4 (N223, N201, N4, N26, N121);
xor XOR2 (N224, N207, N81);
and AND2 (N225, N217, N151);
nand NAND4 (N226, N225, N199, N80, N81);
xor XOR2 (N227, N221, N182);
xor XOR2 (N228, N224, N96);
not NOT1 (N229, N227);
not NOT1 (N230, N218);
not NOT1 (N231, N223);
nor NOR4 (N232, N215, N182, N8, N52);
not NOT1 (N233, N230);
xor XOR2 (N234, N233, N107);
xor XOR2 (N235, N211, N65);
and AND2 (N236, N231, N123);
and AND2 (N237, N226, N125);
not NOT1 (N238, N235);
xor XOR2 (N239, N234, N38);
and AND3 (N240, N220, N113, N173);
buf BUF1 (N241, N203);
nor NOR2 (N242, N237, N135);
and AND3 (N243, N241, N186, N24);
and AND4 (N244, N240, N126, N152, N83);
buf BUF1 (N245, N236);
nand NAND3 (N246, N222, N114, N236);
xor XOR2 (N247, N246, N92);
and AND3 (N248, N242, N174, N43);
buf BUF1 (N249, N232);
and AND4 (N250, N238, N1, N174, N188);
or OR2 (N251, N244, N203);
nand NAND3 (N252, N251, N185, N114);
nor NOR2 (N253, N248, N60);
and AND4 (N254, N253, N88, N146, N17);
nor NOR3 (N255, N229, N167, N181);
nor NOR4 (N256, N249, N195, N154, N65);
nor NOR2 (N257, N239, N38);
nand NAND3 (N258, N252, N106, N25);
and AND3 (N259, N245, N178, N66);
and AND4 (N260, N254, N29, N181, N34);
xor XOR2 (N261, N243, N81);
xor XOR2 (N262, N250, N43);
nor NOR3 (N263, N256, N235, N20);
or OR4 (N264, N228, N162, N30, N218);
nor NOR2 (N265, N260, N181);
nor NOR3 (N266, N261, N33, N20);
nand NAND3 (N267, N255, N198, N243);
xor XOR2 (N268, N259, N66);
buf BUF1 (N269, N268);
and AND3 (N270, N265, N6, N139);
not NOT1 (N271, N262);
or OR4 (N272, N267, N33, N237, N224);
nand NAND3 (N273, N270, N139, N268);
or OR2 (N274, N271, N168);
nor NOR3 (N275, N264, N127, N98);
nand NAND4 (N276, N247, N238, N139, N114);
or OR3 (N277, N269, N64, N111);
buf BUF1 (N278, N257);
nor NOR3 (N279, N266, N274, N267);
buf BUF1 (N280, N231);
and AND2 (N281, N277, N137);
nor NOR2 (N282, N281, N65);
buf BUF1 (N283, N258);
nor NOR4 (N284, N272, N283, N223, N79);
or OR3 (N285, N77, N96, N70);
buf BUF1 (N286, N263);
nand NAND4 (N287, N273, N101, N228, N285);
xor XOR2 (N288, N271, N31);
nor NOR4 (N289, N278, N97, N202, N8);
and AND4 (N290, N289, N183, N151, N244);
or OR3 (N291, N279, N184, N201);
not NOT1 (N292, N280);
not NOT1 (N293, N287);
nand NAND4 (N294, N293, N201, N210, N46);
nand NAND3 (N295, N290, N175, N168);
and AND4 (N296, N286, N131, N111, N222);
nand NAND4 (N297, N292, N220, N88, N180);
and AND3 (N298, N284, N222, N68);
or OR3 (N299, N288, N251, N34);
and AND4 (N300, N282, N40, N62, N28);
buf BUF1 (N301, N295);
xor XOR2 (N302, N300, N132);
buf BUF1 (N303, N294);
not NOT1 (N304, N303);
buf BUF1 (N305, N275);
or OR4 (N306, N297, N91, N108, N249);
nand NAND3 (N307, N291, N37, N54);
buf BUF1 (N308, N301);
nand NAND4 (N309, N306, N298, N110, N242);
xor XOR2 (N310, N67, N145);
endmodule