// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N16009,N16018,N15999,N16023,N16021,N16012,N16017,N16022,N16016,N16024;

nor NOR4 (N25, N1, N9, N21, N13);
buf BUF1 (N26, N8);
nand NAND2 (N27, N4, N11);
and AND2 (N28, N5, N3);
not NOT1 (N29, N4);
and AND3 (N30, N28, N14, N15);
buf BUF1 (N31, N6);
buf BUF1 (N32, N25);
buf BUF1 (N33, N3);
and AND4 (N34, N23, N20, N29, N8);
nand NAND2 (N35, N22, N5);
nand NAND2 (N36, N2, N33);
or OR2 (N37, N29, N19);
not NOT1 (N38, N37);
nor NOR3 (N39, N27, N18, N30);
xor XOR2 (N40, N17, N12);
not NOT1 (N41, N22);
nand NAND4 (N42, N38, N4, N37, N33);
nand NAND2 (N43, N42, N2);
xor XOR2 (N44, N32, N41);
buf BUF1 (N45, N41);
xor XOR2 (N46, N36, N40);
xor XOR2 (N47, N46, N44);
not NOT1 (N48, N19);
and AND4 (N49, N45, N43, N27, N11);
or OR3 (N50, N11, N35, N16);
or OR4 (N51, N33, N15, N7, N23);
nor NOR2 (N52, N6, N16);
and AND4 (N53, N31, N48, N4, N48);
nand NAND4 (N54, N24, N48, N37, N28);
not NOT1 (N55, N47);
not NOT1 (N56, N51);
xor XOR2 (N57, N39, N39);
not NOT1 (N58, N50);
nand NAND3 (N59, N58, N50, N1);
nand NAND4 (N60, N54, N57, N39, N58);
or OR2 (N61, N25, N50);
buf BUF1 (N62, N26);
or OR2 (N63, N56, N45);
buf BUF1 (N64, N49);
nand NAND4 (N65, N55, N44, N17, N20);
nand NAND3 (N66, N60, N36, N15);
nand NAND2 (N67, N63, N9);
buf BUF1 (N68, N66);
xor XOR2 (N69, N61, N43);
not NOT1 (N70, N69);
xor XOR2 (N71, N68, N52);
or OR2 (N72, N68, N45);
and AND3 (N73, N34, N34, N6);
and AND3 (N74, N73, N32, N18);
and AND3 (N75, N53, N60, N21);
not NOT1 (N76, N75);
and AND4 (N77, N64, N42, N4, N34);
or OR2 (N78, N59, N74);
buf BUF1 (N79, N32);
nand NAND2 (N80, N70, N34);
nor NOR3 (N81, N78, N35, N54);
and AND2 (N82, N67, N43);
nor NOR4 (N83, N62, N49, N38, N6);
or OR3 (N84, N79, N69, N82);
or OR2 (N85, N55, N77);
and AND4 (N86, N63, N32, N73, N19);
nor NOR4 (N87, N83, N3, N9, N56);
or OR4 (N88, N65, N33, N33, N26);
or OR3 (N89, N71, N21, N82);
nor NOR4 (N90, N89, N86, N18, N39);
not NOT1 (N91, N76);
and AND3 (N92, N62, N64, N22);
buf BUF1 (N93, N84);
nor NOR4 (N94, N90, N23, N5, N59);
not NOT1 (N95, N81);
nand NAND4 (N96, N92, N65, N77, N49);
nor NOR4 (N97, N91, N73, N34, N84);
buf BUF1 (N98, N94);
buf BUF1 (N99, N85);
or OR3 (N100, N72, N75, N88);
nor NOR4 (N101, N30, N2, N45, N68);
nand NAND4 (N102, N93, N37, N9, N58);
or OR4 (N103, N97, N56, N22, N52);
xor XOR2 (N104, N87, N4);
buf BUF1 (N105, N101);
nand NAND4 (N106, N95, N24, N95, N2);
nor NOR4 (N107, N100, N100, N53, N26);
buf BUF1 (N108, N104);
nand NAND4 (N109, N99, N85, N17, N60);
buf BUF1 (N110, N108);
nand NAND2 (N111, N96, N14);
nand NAND3 (N112, N106, N44, N92);
nor NOR4 (N113, N98, N96, N86, N112);
nand NAND2 (N114, N5, N99);
not NOT1 (N115, N111);
xor XOR2 (N116, N105, N113);
nor NOR2 (N117, N56, N65);
not NOT1 (N118, N114);
and AND4 (N119, N103, N31, N33, N104);
buf BUF1 (N120, N110);
xor XOR2 (N121, N115, N65);
not NOT1 (N122, N120);
nor NOR3 (N123, N117, N66, N107);
and AND2 (N124, N80, N40);
nand NAND3 (N125, N84, N59, N78);
and AND4 (N126, N125, N47, N6, N119);
buf BUF1 (N127, N81);
nand NAND2 (N128, N116, N73);
buf BUF1 (N129, N124);
buf BUF1 (N130, N102);
or OR3 (N131, N123, N32, N23);
xor XOR2 (N132, N122, N86);
nand NAND2 (N133, N127, N69);
and AND2 (N134, N128, N78);
xor XOR2 (N135, N130, N81);
nor NOR4 (N136, N118, N102, N72, N15);
nor NOR2 (N137, N136, N121);
xor XOR2 (N138, N34, N61);
buf BUF1 (N139, N137);
not NOT1 (N140, N132);
nand NAND2 (N141, N135, N98);
and AND3 (N142, N140, N132, N114);
not NOT1 (N143, N126);
nor NOR2 (N144, N141, N20);
or OR4 (N145, N129, N66, N39, N40);
buf BUF1 (N146, N109);
nor NOR2 (N147, N134, N57);
buf BUF1 (N148, N143);
xor XOR2 (N149, N131, N112);
buf BUF1 (N150, N139);
or OR2 (N151, N138, N3);
xor XOR2 (N152, N145, N48);
and AND3 (N153, N152, N128, N111);
nand NAND2 (N154, N150, N64);
nand NAND4 (N155, N149, N146, N88, N68);
not NOT1 (N156, N44);
buf BUF1 (N157, N154);
nor NOR3 (N158, N157, N92, N12);
xor XOR2 (N159, N156, N9);
nand NAND3 (N160, N151, N11, N149);
nand NAND2 (N161, N155, N36);
nor NOR4 (N162, N153, N32, N35, N84);
or OR2 (N163, N133, N4);
buf BUF1 (N164, N144);
buf BUF1 (N165, N142);
not NOT1 (N166, N165);
xor XOR2 (N167, N159, N120);
and AND4 (N168, N163, N93, N75, N129);
or OR2 (N169, N147, N68);
not NOT1 (N170, N167);
and AND4 (N171, N169, N146, N60, N58);
not NOT1 (N172, N162);
nor NOR3 (N173, N170, N95, N98);
not NOT1 (N174, N160);
not NOT1 (N175, N164);
or OR3 (N176, N168, N59, N18);
or OR3 (N177, N158, N161, N24);
xor XOR2 (N178, N4, N14);
not NOT1 (N179, N172);
buf BUF1 (N180, N179);
or OR4 (N181, N173, N38, N34, N158);
and AND4 (N182, N177, N35, N133, N86);
nor NOR3 (N183, N176, N103, N142);
buf BUF1 (N184, N171);
not NOT1 (N185, N181);
xor XOR2 (N186, N178, N157);
nand NAND4 (N187, N166, N105, N26, N171);
not NOT1 (N188, N186);
buf BUF1 (N189, N180);
buf BUF1 (N190, N182);
nor NOR3 (N191, N190, N151, N55);
nand NAND3 (N192, N148, N85, N29);
nor NOR3 (N193, N191, N55, N119);
buf BUF1 (N194, N185);
not NOT1 (N195, N193);
nor NOR3 (N196, N184, N15, N174);
nor NOR4 (N197, N177, N40, N76, N120);
nand NAND3 (N198, N188, N79, N50);
buf BUF1 (N199, N189);
or OR3 (N200, N183, N34, N27);
not NOT1 (N201, N199);
buf BUF1 (N202, N187);
nor NOR4 (N203, N197, N25, N73, N30);
and AND2 (N204, N196, N179);
not NOT1 (N205, N175);
not NOT1 (N206, N201);
nand NAND4 (N207, N195, N35, N47, N48);
xor XOR2 (N208, N198, N8);
xor XOR2 (N209, N205, N69);
and AND2 (N210, N207, N20);
and AND4 (N211, N194, N136, N80, N8);
and AND2 (N212, N204, N10);
nor NOR3 (N213, N210, N154, N139);
xor XOR2 (N214, N208, N46);
nor NOR2 (N215, N214, N115);
and AND2 (N216, N211, N198);
or OR3 (N217, N216, N119, N192);
xor XOR2 (N218, N206, N40);
nand NAND3 (N219, N149, N167, N49);
and AND4 (N220, N212, N36, N169, N47);
nand NAND4 (N221, N213, N15, N117, N79);
and AND3 (N222, N221, N220, N213);
nand NAND3 (N223, N35, N33, N189);
and AND4 (N224, N223, N128, N38, N61);
and AND4 (N225, N202, N59, N141, N7);
buf BUF1 (N226, N200);
and AND2 (N227, N217, N190);
xor XOR2 (N228, N209, N56);
nor NOR4 (N229, N224, N162, N48, N138);
xor XOR2 (N230, N228, N143);
nand NAND3 (N231, N219, N102, N212);
nor NOR4 (N232, N227, N171, N195, N177);
and AND2 (N233, N230, N72);
nor NOR3 (N234, N203, N137, N55);
buf BUF1 (N235, N215);
nand NAND3 (N236, N226, N180, N215);
buf BUF1 (N237, N231);
not NOT1 (N238, N222);
nor NOR2 (N239, N236, N89);
buf BUF1 (N240, N234);
buf BUF1 (N241, N239);
nor NOR3 (N242, N229, N114, N169);
or OR4 (N243, N218, N165, N64, N66);
nand NAND2 (N244, N237, N53);
not NOT1 (N245, N243);
nand NAND3 (N246, N225, N29, N220);
or OR2 (N247, N232, N43);
xor XOR2 (N248, N246, N7);
xor XOR2 (N249, N247, N29);
nor NOR2 (N250, N245, N21);
nor NOR3 (N251, N235, N118, N6);
xor XOR2 (N252, N248, N148);
nand NAND4 (N253, N241, N93, N16, N186);
or OR2 (N254, N242, N249);
not NOT1 (N255, N158);
and AND3 (N256, N250, N51, N172);
nor NOR2 (N257, N244, N56);
xor XOR2 (N258, N240, N114);
nor NOR3 (N259, N251, N207, N53);
nor NOR4 (N260, N254, N54, N126, N236);
nor NOR4 (N261, N257, N214, N216, N247);
nor NOR4 (N262, N233, N142, N208, N214);
buf BUF1 (N263, N238);
buf BUF1 (N264, N253);
nand NAND4 (N265, N262, N11, N160, N65);
xor XOR2 (N266, N260, N262);
nor NOR3 (N267, N263, N137, N92);
xor XOR2 (N268, N256, N16);
not NOT1 (N269, N267);
not NOT1 (N270, N269);
nand NAND3 (N271, N268, N32, N119);
buf BUF1 (N272, N264);
or OR3 (N273, N261, N140, N114);
not NOT1 (N274, N265);
xor XOR2 (N275, N271, N230);
and AND4 (N276, N270, N122, N166, N268);
xor XOR2 (N277, N258, N148);
not NOT1 (N278, N252);
xor XOR2 (N279, N272, N227);
or OR3 (N280, N273, N207, N276);
xor XOR2 (N281, N70, N238);
nand NAND4 (N282, N274, N47, N74, N43);
and AND3 (N283, N255, N99, N159);
or OR2 (N284, N266, N117);
buf BUF1 (N285, N283);
not NOT1 (N286, N282);
xor XOR2 (N287, N281, N250);
nand NAND4 (N288, N280, N121, N153, N110);
not NOT1 (N289, N288);
and AND2 (N290, N287, N131);
and AND4 (N291, N279, N66, N222, N52);
xor XOR2 (N292, N285, N124);
and AND4 (N293, N291, N272, N42, N266);
nor NOR3 (N294, N286, N26, N252);
and AND2 (N295, N293, N245);
or OR2 (N296, N295, N144);
nand NAND2 (N297, N259, N182);
buf BUF1 (N298, N294);
nand NAND2 (N299, N289, N222);
xor XOR2 (N300, N297, N214);
nor NOR2 (N301, N277, N264);
not NOT1 (N302, N290);
not NOT1 (N303, N299);
nor NOR4 (N304, N301, N186, N211, N233);
nand NAND4 (N305, N298, N196, N32, N251);
and AND4 (N306, N303, N244, N236, N46);
nand NAND3 (N307, N305, N101, N107);
nand NAND3 (N308, N304, N70, N217);
nand NAND4 (N309, N306, N9, N263, N172);
not NOT1 (N310, N296);
nand NAND2 (N311, N275, N259);
nor NOR2 (N312, N310, N38);
xor XOR2 (N313, N302, N131);
not NOT1 (N314, N308);
nand NAND3 (N315, N312, N99, N210);
nor NOR4 (N316, N313, N268, N286, N153);
nor NOR4 (N317, N292, N40, N230, N246);
or OR2 (N318, N316, N151);
not NOT1 (N319, N300);
buf BUF1 (N320, N284);
nor NOR2 (N321, N319, N26);
and AND4 (N322, N315, N253, N207, N115);
not NOT1 (N323, N314);
nand NAND3 (N324, N322, N146, N184);
nor NOR4 (N325, N320, N84, N222, N299);
nor NOR2 (N326, N278, N269);
xor XOR2 (N327, N321, N67);
nor NOR4 (N328, N326, N236, N88, N233);
nor NOR3 (N329, N324, N178, N127);
nand NAND2 (N330, N327, N138);
and AND3 (N331, N318, N87, N279);
buf BUF1 (N332, N323);
nor NOR2 (N333, N331, N97);
nor NOR2 (N334, N307, N72);
nor NOR3 (N335, N328, N82, N51);
nand NAND3 (N336, N333, N94, N184);
xor XOR2 (N337, N309, N61);
nand NAND4 (N338, N330, N181, N135, N120);
buf BUF1 (N339, N334);
xor XOR2 (N340, N311, N158);
not NOT1 (N341, N337);
buf BUF1 (N342, N340);
xor XOR2 (N343, N338, N129);
not NOT1 (N344, N335);
nand NAND3 (N345, N317, N174, N60);
or OR4 (N346, N341, N246, N282, N185);
not NOT1 (N347, N339);
not NOT1 (N348, N329);
xor XOR2 (N349, N332, N91);
xor XOR2 (N350, N336, N72);
xor XOR2 (N351, N346, N78);
xor XOR2 (N352, N343, N14);
nor NOR4 (N353, N348, N120, N312, N229);
or OR2 (N354, N347, N5);
buf BUF1 (N355, N349);
or OR3 (N356, N345, N180, N198);
xor XOR2 (N357, N344, N310);
or OR4 (N358, N355, N268, N328, N283);
nand NAND4 (N359, N350, N77, N149, N59);
xor XOR2 (N360, N358, N284);
xor XOR2 (N361, N356, N1);
buf BUF1 (N362, N361);
nand NAND2 (N363, N354, N114);
not NOT1 (N364, N352);
nor NOR3 (N365, N360, N105, N257);
xor XOR2 (N366, N363, N136);
buf BUF1 (N367, N365);
and AND4 (N368, N359, N1, N265, N29);
or OR4 (N369, N368, N50, N245, N217);
not NOT1 (N370, N367);
nor NOR4 (N371, N369, N250, N338, N295);
nor NOR4 (N372, N362, N252, N34, N90);
and AND3 (N373, N371, N11, N22);
xor XOR2 (N374, N373, N183);
not NOT1 (N375, N357);
and AND3 (N376, N366, N87, N248);
buf BUF1 (N377, N375);
nand NAND3 (N378, N374, N63, N280);
nor NOR2 (N379, N342, N357);
nand NAND3 (N380, N351, N177, N247);
not NOT1 (N381, N325);
and AND4 (N382, N379, N196, N108, N380);
or OR4 (N383, N239, N179, N195, N106);
nor NOR4 (N384, N370, N295, N368, N275);
or OR3 (N385, N372, N126, N257);
buf BUF1 (N386, N381);
nand NAND2 (N387, N383, N281);
or OR2 (N388, N382, N105);
nor NOR2 (N389, N387, N199);
buf BUF1 (N390, N364);
and AND4 (N391, N386, N91, N272, N342);
or OR2 (N392, N391, N354);
nand NAND2 (N393, N378, N133);
and AND3 (N394, N393, N165, N343);
nand NAND3 (N395, N388, N237, N17);
buf BUF1 (N396, N377);
buf BUF1 (N397, N385);
buf BUF1 (N398, N392);
buf BUF1 (N399, N384);
xor XOR2 (N400, N399, N239);
nand NAND2 (N401, N394, N240);
or OR4 (N402, N376, N29, N1, N182);
or OR3 (N403, N398, N181, N312);
nand NAND3 (N404, N395, N314, N32);
nor NOR2 (N405, N404, N288);
nand NAND3 (N406, N390, N326, N329);
and AND4 (N407, N396, N371, N353, N227);
nand NAND3 (N408, N265, N351, N24);
not NOT1 (N409, N397);
or OR3 (N410, N406, N281, N64);
buf BUF1 (N411, N389);
nor NOR2 (N412, N405, N188);
not NOT1 (N413, N412);
not NOT1 (N414, N403);
nand NAND3 (N415, N414, N214, N137);
or OR3 (N416, N409, N147, N110);
or OR4 (N417, N416, N120, N281, N161);
xor XOR2 (N418, N413, N55);
buf BUF1 (N419, N410);
nand NAND4 (N420, N411, N395, N134, N88);
not NOT1 (N421, N420);
nor NOR2 (N422, N400, N311);
or OR2 (N423, N401, N410);
buf BUF1 (N424, N417);
and AND4 (N425, N408, N285, N183, N199);
nor NOR3 (N426, N424, N225, N289);
xor XOR2 (N427, N418, N397);
buf BUF1 (N428, N402);
or OR4 (N429, N415, N80, N236, N224);
nand NAND2 (N430, N429, N158);
buf BUF1 (N431, N427);
or OR3 (N432, N426, N23, N199);
and AND3 (N433, N407, N50, N326);
not NOT1 (N434, N422);
and AND2 (N435, N430, N253);
not NOT1 (N436, N425);
and AND3 (N437, N423, N211, N159);
not NOT1 (N438, N431);
or OR3 (N439, N434, N100, N422);
or OR4 (N440, N419, N22, N280, N353);
nand NAND3 (N441, N438, N98, N124);
xor XOR2 (N442, N421, N175);
and AND2 (N443, N432, N388);
or OR3 (N444, N437, N21, N410);
not NOT1 (N445, N440);
buf BUF1 (N446, N428);
and AND2 (N447, N444, N31);
not NOT1 (N448, N445);
and AND2 (N449, N436, N168);
nor NOR3 (N450, N448, N293, N274);
and AND2 (N451, N435, N183);
nand NAND2 (N452, N441, N339);
xor XOR2 (N453, N446, N132);
nand NAND2 (N454, N442, N371);
or OR3 (N455, N452, N131, N139);
nand NAND3 (N456, N455, N306, N360);
xor XOR2 (N457, N439, N27);
not NOT1 (N458, N451);
nand NAND3 (N459, N456, N354, N30);
nand NAND4 (N460, N449, N41, N162, N165);
and AND2 (N461, N453, N185);
not NOT1 (N462, N454);
not NOT1 (N463, N460);
and AND3 (N464, N433, N357, N367);
xor XOR2 (N465, N464, N436);
and AND2 (N466, N459, N376);
nor NOR3 (N467, N465, N359, N433);
not NOT1 (N468, N458);
or OR4 (N469, N466, N159, N194, N340);
nor NOR3 (N470, N468, N123, N406);
or OR2 (N471, N470, N31);
xor XOR2 (N472, N469, N417);
xor XOR2 (N473, N447, N271);
buf BUF1 (N474, N467);
xor XOR2 (N475, N461, N401);
or OR2 (N476, N462, N308);
nand NAND3 (N477, N474, N401, N407);
and AND3 (N478, N473, N246, N16);
xor XOR2 (N479, N475, N319);
xor XOR2 (N480, N463, N58);
buf BUF1 (N481, N477);
buf BUF1 (N482, N476);
nor NOR2 (N483, N480, N311);
and AND4 (N484, N472, N482, N277, N230);
xor XOR2 (N485, N390, N348);
or OR2 (N486, N457, N319);
nand NAND3 (N487, N486, N340, N70);
xor XOR2 (N488, N487, N130);
nand NAND3 (N489, N471, N218, N333);
nor NOR3 (N490, N479, N236, N104);
buf BUF1 (N491, N478);
not NOT1 (N492, N443);
nand NAND2 (N493, N450, N425);
nand NAND2 (N494, N491, N212);
xor XOR2 (N495, N492, N219);
xor XOR2 (N496, N489, N376);
nor NOR2 (N497, N495, N170);
xor XOR2 (N498, N483, N270);
xor XOR2 (N499, N488, N159);
and AND2 (N500, N499, N375);
not NOT1 (N501, N494);
and AND3 (N502, N481, N95, N70);
or OR4 (N503, N493, N419, N128, N25);
xor XOR2 (N504, N485, N105);
not NOT1 (N505, N500);
and AND3 (N506, N498, N34, N472);
xor XOR2 (N507, N497, N187);
and AND4 (N508, N507, N144, N182, N316);
not NOT1 (N509, N501);
nand NAND4 (N510, N496, N168, N103, N476);
buf BUF1 (N511, N508);
and AND3 (N512, N510, N174, N505);
nand NAND3 (N513, N473, N31, N25);
or OR3 (N514, N504, N126, N20);
not NOT1 (N515, N506);
or OR2 (N516, N513, N106);
not NOT1 (N517, N515);
and AND2 (N518, N503, N308);
and AND3 (N519, N490, N61, N352);
xor XOR2 (N520, N516, N197);
xor XOR2 (N521, N520, N208);
nand NAND3 (N522, N511, N472, N452);
or OR2 (N523, N519, N482);
nand NAND2 (N524, N517, N482);
nand NAND4 (N525, N509, N394, N169, N518);
xor XOR2 (N526, N29, N435);
and AND2 (N527, N525, N203);
or OR4 (N528, N523, N111, N201, N519);
or OR3 (N529, N514, N279, N8);
nand NAND3 (N530, N526, N393, N269);
buf BUF1 (N531, N502);
nor NOR3 (N532, N484, N463, N137);
not NOT1 (N533, N524);
xor XOR2 (N534, N521, N182);
not NOT1 (N535, N534);
and AND3 (N536, N512, N285, N508);
nor NOR3 (N537, N528, N267, N5);
or OR4 (N538, N537, N3, N504, N140);
xor XOR2 (N539, N530, N378);
buf BUF1 (N540, N539);
buf BUF1 (N541, N540);
not NOT1 (N542, N529);
nand NAND2 (N543, N535, N442);
nor NOR2 (N544, N527, N481);
and AND2 (N545, N532, N6);
xor XOR2 (N546, N522, N428);
not NOT1 (N547, N542);
nor NOR4 (N548, N544, N21, N246, N80);
and AND3 (N549, N533, N103, N183);
nor NOR2 (N550, N531, N269);
or OR2 (N551, N545, N68);
xor XOR2 (N552, N546, N157);
nand NAND2 (N553, N538, N153);
and AND4 (N554, N547, N221, N67, N168);
nand NAND2 (N555, N552, N97);
and AND2 (N556, N541, N312);
nand NAND4 (N557, N550, N274, N521, N128);
nand NAND4 (N558, N543, N521, N315, N295);
xor XOR2 (N559, N554, N340);
nand NAND4 (N560, N556, N498, N23, N214);
nand NAND3 (N561, N548, N466, N437);
or OR2 (N562, N555, N297);
not NOT1 (N563, N559);
buf BUF1 (N564, N558);
or OR2 (N565, N564, N378);
nand NAND2 (N566, N551, N69);
nand NAND2 (N567, N557, N65);
and AND4 (N568, N565, N382, N558, N550);
or OR4 (N569, N561, N452, N393, N303);
nor NOR2 (N570, N563, N249);
or OR3 (N571, N570, N532, N181);
nand NAND2 (N572, N567, N498);
not NOT1 (N573, N536);
nor NOR3 (N574, N571, N340, N207);
buf BUF1 (N575, N569);
nand NAND4 (N576, N572, N268, N422, N7);
nor NOR4 (N577, N553, N124, N37, N359);
nand NAND3 (N578, N575, N37, N284);
buf BUF1 (N579, N562);
nand NAND3 (N580, N568, N286, N220);
xor XOR2 (N581, N566, N13);
nor NOR2 (N582, N580, N129);
not NOT1 (N583, N579);
or OR3 (N584, N577, N99, N516);
buf BUF1 (N585, N576);
or OR2 (N586, N560, N410);
and AND2 (N587, N581, N243);
buf BUF1 (N588, N583);
or OR3 (N589, N585, N218, N220);
xor XOR2 (N590, N584, N437);
xor XOR2 (N591, N573, N396);
and AND4 (N592, N578, N573, N401, N96);
nor NOR3 (N593, N574, N371, N287);
or OR2 (N594, N593, N433);
or OR2 (N595, N582, N489);
buf BUF1 (N596, N589);
or OR4 (N597, N596, N305, N569, N288);
xor XOR2 (N598, N594, N143);
xor XOR2 (N599, N590, N250);
or OR4 (N600, N592, N287, N325, N218);
xor XOR2 (N601, N595, N298);
xor XOR2 (N602, N591, N591);
xor XOR2 (N603, N601, N391);
xor XOR2 (N604, N588, N487);
and AND4 (N605, N598, N534, N362, N563);
and AND2 (N606, N605, N11);
nand NAND4 (N607, N587, N376, N160, N332);
not NOT1 (N608, N549);
not NOT1 (N609, N602);
buf BUF1 (N610, N608);
xor XOR2 (N611, N600, N600);
and AND4 (N612, N604, N333, N216, N160);
or OR2 (N613, N599, N514);
or OR4 (N614, N597, N84, N288, N562);
xor XOR2 (N615, N607, N282);
nand NAND3 (N616, N615, N174, N263);
nand NAND2 (N617, N586, N210);
buf BUF1 (N618, N614);
nor NOR3 (N619, N617, N479, N125);
xor XOR2 (N620, N613, N439);
or OR2 (N621, N609, N127);
nand NAND2 (N622, N619, N446);
nand NAND4 (N623, N621, N494, N7, N139);
not NOT1 (N624, N618);
not NOT1 (N625, N611);
nor NOR3 (N626, N616, N87, N170);
and AND3 (N627, N606, N95, N577);
xor XOR2 (N628, N623, N256);
and AND4 (N629, N627, N42, N578, N596);
nor NOR2 (N630, N610, N35);
nor NOR3 (N631, N622, N78, N145);
nor NOR2 (N632, N628, N489);
xor XOR2 (N633, N612, N500);
nor NOR4 (N634, N625, N356, N469, N325);
not NOT1 (N635, N634);
nor NOR3 (N636, N624, N234, N561);
or OR3 (N637, N629, N275, N99);
and AND2 (N638, N637, N326);
nand NAND2 (N639, N620, N268);
not NOT1 (N640, N631);
nor NOR4 (N641, N638, N210, N290, N355);
or OR2 (N642, N640, N484);
nand NAND2 (N643, N636, N206);
buf BUF1 (N644, N626);
or OR2 (N645, N630, N122);
buf BUF1 (N646, N603);
buf BUF1 (N647, N633);
nor NOR4 (N648, N641, N103, N421, N359);
nor NOR4 (N649, N635, N612, N647, N555);
buf BUF1 (N650, N537);
xor XOR2 (N651, N650, N617);
buf BUF1 (N652, N649);
nor NOR3 (N653, N643, N450, N112);
xor XOR2 (N654, N651, N336);
nand NAND4 (N655, N652, N4, N326, N146);
nand NAND2 (N656, N645, N622);
nand NAND3 (N657, N648, N526, N111);
nor NOR4 (N658, N657, N152, N153, N290);
or OR3 (N659, N658, N61, N42);
xor XOR2 (N660, N655, N451);
not NOT1 (N661, N639);
nor NOR2 (N662, N660, N541);
xor XOR2 (N663, N644, N397);
nor NOR2 (N664, N653, N434);
nand NAND2 (N665, N659, N189);
buf BUF1 (N666, N665);
or OR4 (N667, N663, N496, N382, N644);
and AND4 (N668, N667, N393, N23, N514);
buf BUF1 (N669, N646);
nand NAND3 (N670, N669, N120, N213);
and AND4 (N671, N661, N205, N631, N72);
not NOT1 (N672, N656);
nor NOR2 (N673, N670, N222);
and AND4 (N674, N642, N375, N10, N389);
or OR3 (N675, N666, N59, N468);
nand NAND2 (N676, N671, N655);
nor NOR3 (N677, N654, N453, N525);
nor NOR4 (N678, N672, N380, N624, N594);
buf BUF1 (N679, N668);
nand NAND2 (N680, N676, N509);
not NOT1 (N681, N664);
or OR4 (N682, N674, N104, N242, N240);
nor NOR3 (N683, N662, N377, N555);
nand NAND3 (N684, N675, N226, N11);
nor NOR2 (N685, N632, N535);
not NOT1 (N686, N677);
xor XOR2 (N687, N673, N413);
or OR4 (N688, N679, N104, N455, N7);
nand NAND3 (N689, N683, N408, N95);
and AND4 (N690, N680, N73, N658, N139);
buf BUF1 (N691, N689);
xor XOR2 (N692, N682, N184);
not NOT1 (N693, N684);
nand NAND3 (N694, N688, N45, N6);
xor XOR2 (N695, N694, N403);
nor NOR4 (N696, N690, N75, N88, N542);
nand NAND4 (N697, N687, N324, N420, N481);
and AND4 (N698, N691, N338, N13, N277);
nand NAND3 (N699, N686, N374, N105);
nor NOR4 (N700, N695, N92, N146, N274);
or OR4 (N701, N700, N414, N275, N475);
buf BUF1 (N702, N685);
and AND3 (N703, N696, N255, N235);
nor NOR4 (N704, N703, N313, N404, N262);
not NOT1 (N705, N697);
or OR2 (N706, N678, N251);
nand NAND2 (N707, N698, N205);
not NOT1 (N708, N704);
not NOT1 (N709, N701);
xor XOR2 (N710, N709, N493);
nand NAND4 (N711, N699, N151, N43, N607);
or OR2 (N712, N693, N298);
and AND2 (N713, N702, N80);
xor XOR2 (N714, N711, N347);
or OR3 (N715, N710, N230, N140);
and AND4 (N716, N713, N666, N639, N562);
buf BUF1 (N717, N714);
not NOT1 (N718, N681);
or OR3 (N719, N706, N446, N556);
xor XOR2 (N720, N708, N495);
buf BUF1 (N721, N707);
xor XOR2 (N722, N721, N51);
or OR4 (N723, N705, N548, N254, N301);
not NOT1 (N724, N720);
nand NAND3 (N725, N717, N76, N508);
buf BUF1 (N726, N715);
or OR2 (N727, N723, N638);
and AND4 (N728, N716, N476, N489, N265);
nor NOR2 (N729, N724, N64);
or OR2 (N730, N728, N284);
buf BUF1 (N731, N719);
xor XOR2 (N732, N730, N169);
not NOT1 (N733, N725);
or OR2 (N734, N729, N183);
xor XOR2 (N735, N722, N73);
xor XOR2 (N736, N727, N614);
nand NAND3 (N737, N735, N310, N182);
and AND3 (N738, N736, N150, N677);
nor NOR4 (N739, N737, N470, N111, N274);
and AND3 (N740, N731, N205, N482);
not NOT1 (N741, N738);
or OR2 (N742, N739, N342);
or OR2 (N743, N734, N120);
or OR2 (N744, N740, N598);
not NOT1 (N745, N742);
buf BUF1 (N746, N745);
xor XOR2 (N747, N692, N45);
or OR4 (N748, N712, N143, N400, N68);
nor NOR4 (N749, N718, N726, N683, N403);
or OR3 (N750, N450, N666, N697);
buf BUF1 (N751, N747);
and AND2 (N752, N733, N443);
nand NAND3 (N753, N750, N414, N85);
nand NAND2 (N754, N748, N593);
buf BUF1 (N755, N743);
and AND3 (N756, N744, N609, N176);
or OR3 (N757, N756, N62, N519);
or OR4 (N758, N755, N435, N241, N588);
or OR4 (N759, N749, N180, N263, N554);
or OR4 (N760, N741, N136, N394, N185);
xor XOR2 (N761, N760, N558);
xor XOR2 (N762, N757, N580);
nand NAND4 (N763, N759, N338, N160, N198);
nand NAND4 (N764, N746, N434, N713, N674);
xor XOR2 (N765, N763, N89);
buf BUF1 (N766, N761);
or OR2 (N767, N765, N757);
buf BUF1 (N768, N753);
or OR3 (N769, N732, N236, N270);
or OR2 (N770, N767, N386);
and AND3 (N771, N766, N265, N635);
buf BUF1 (N772, N752);
not NOT1 (N773, N771);
and AND3 (N774, N773, N464, N673);
or OR4 (N775, N754, N297, N457, N363);
or OR3 (N776, N762, N34, N349);
buf BUF1 (N777, N751);
buf BUF1 (N778, N768);
nor NOR2 (N779, N775, N649);
nand NAND2 (N780, N758, N662);
and AND3 (N781, N770, N331, N399);
or OR4 (N782, N781, N749, N121, N3);
buf BUF1 (N783, N779);
xor XOR2 (N784, N772, N682);
nand NAND3 (N785, N774, N413, N481);
nand NAND2 (N786, N764, N77);
buf BUF1 (N787, N785);
buf BUF1 (N788, N778);
xor XOR2 (N789, N788, N646);
not NOT1 (N790, N777);
and AND2 (N791, N790, N102);
nand NAND4 (N792, N784, N655, N658, N564);
nand NAND3 (N793, N782, N362, N106);
not NOT1 (N794, N791);
nand NAND3 (N795, N786, N241, N124);
nor NOR2 (N796, N787, N680);
not NOT1 (N797, N783);
or OR3 (N798, N793, N304, N211);
buf BUF1 (N799, N798);
not NOT1 (N800, N797);
nor NOR4 (N801, N794, N275, N720, N508);
not NOT1 (N802, N796);
xor XOR2 (N803, N792, N512);
not NOT1 (N804, N802);
or OR2 (N805, N804, N164);
or OR4 (N806, N776, N223, N716, N496);
or OR2 (N807, N803, N55);
or OR3 (N808, N789, N745, N302);
xor XOR2 (N809, N808, N465);
or OR2 (N810, N807, N544);
and AND2 (N811, N805, N195);
and AND4 (N812, N795, N689, N32, N134);
nand NAND4 (N813, N799, N136, N138, N107);
xor XOR2 (N814, N806, N344);
not NOT1 (N815, N810);
xor XOR2 (N816, N809, N486);
not NOT1 (N817, N811);
xor XOR2 (N818, N814, N764);
nand NAND3 (N819, N801, N527, N118);
not NOT1 (N820, N800);
not NOT1 (N821, N818);
not NOT1 (N822, N812);
nand NAND3 (N823, N769, N266, N725);
xor XOR2 (N824, N822, N630);
nor NOR2 (N825, N816, N242);
or OR3 (N826, N815, N348, N309);
nand NAND3 (N827, N826, N764, N224);
nor NOR3 (N828, N817, N691, N734);
nor NOR3 (N829, N813, N380, N484);
not NOT1 (N830, N821);
and AND4 (N831, N828, N704, N446, N521);
and AND2 (N832, N825, N455);
and AND4 (N833, N832, N730, N288, N76);
or OR2 (N834, N829, N212);
and AND3 (N835, N827, N423, N229);
not NOT1 (N836, N834);
buf BUF1 (N837, N836);
or OR2 (N838, N830, N258);
and AND4 (N839, N819, N830, N101, N767);
nor NOR4 (N840, N833, N112, N51, N734);
buf BUF1 (N841, N820);
and AND2 (N842, N841, N440);
or OR4 (N843, N780, N172, N419, N159);
xor XOR2 (N844, N835, N196);
not NOT1 (N845, N839);
nand NAND2 (N846, N823, N395);
nor NOR2 (N847, N842, N713);
xor XOR2 (N848, N845, N771);
nand NAND2 (N849, N824, N809);
nor NOR4 (N850, N847, N606, N596, N294);
or OR4 (N851, N846, N225, N286, N300);
not NOT1 (N852, N849);
xor XOR2 (N853, N848, N384);
nand NAND2 (N854, N853, N629);
not NOT1 (N855, N840);
and AND3 (N856, N843, N93, N39);
nand NAND2 (N857, N851, N73);
and AND3 (N858, N854, N144, N470);
xor XOR2 (N859, N855, N210);
and AND3 (N860, N858, N431, N263);
nand NAND3 (N861, N838, N423, N749);
and AND4 (N862, N856, N796, N843, N519);
or OR4 (N863, N861, N56, N620, N317);
xor XOR2 (N864, N850, N525);
not NOT1 (N865, N844);
xor XOR2 (N866, N831, N773);
and AND4 (N867, N863, N631, N825, N692);
xor XOR2 (N868, N837, N142);
or OR4 (N869, N852, N150, N346, N47);
and AND3 (N870, N864, N706, N513);
and AND4 (N871, N866, N181, N2, N211);
buf BUF1 (N872, N865);
not NOT1 (N873, N862);
nor NOR3 (N874, N867, N535, N591);
not NOT1 (N875, N872);
and AND2 (N876, N874, N808);
or OR4 (N877, N873, N330, N778, N5);
nand NAND2 (N878, N876, N598);
not NOT1 (N879, N878);
nand NAND4 (N880, N875, N378, N3, N627);
not NOT1 (N881, N880);
buf BUF1 (N882, N868);
buf BUF1 (N883, N869);
buf BUF1 (N884, N881);
buf BUF1 (N885, N857);
nor NOR4 (N886, N870, N791, N75, N15);
xor XOR2 (N887, N860, N709);
or OR3 (N888, N883, N367, N519);
or OR4 (N889, N882, N343, N815, N354);
not NOT1 (N890, N885);
and AND4 (N891, N890, N410, N574, N297);
not NOT1 (N892, N891);
or OR4 (N893, N886, N151, N677, N218);
nor NOR4 (N894, N887, N233, N577, N4);
nor NOR2 (N895, N859, N412);
xor XOR2 (N896, N888, N652);
buf BUF1 (N897, N896);
or OR2 (N898, N894, N438);
not NOT1 (N899, N897);
nand NAND3 (N900, N895, N478, N173);
nand NAND4 (N901, N893, N11, N128, N379);
not NOT1 (N902, N900);
not NOT1 (N903, N871);
or OR4 (N904, N892, N884, N535, N671);
and AND2 (N905, N459, N776);
and AND2 (N906, N877, N903);
or OR2 (N907, N435, N442);
buf BUF1 (N908, N901);
and AND3 (N909, N904, N567, N149);
not NOT1 (N910, N909);
and AND3 (N911, N907, N381, N638);
nor NOR2 (N912, N898, N45);
and AND2 (N913, N912, N168);
nor NOR4 (N914, N908, N604, N480, N905);
not NOT1 (N915, N223);
nor NOR4 (N916, N889, N631, N32, N399);
and AND2 (N917, N913, N114);
nor NOR2 (N918, N917, N5);
or OR2 (N919, N914, N324);
or OR3 (N920, N910, N884, N467);
buf BUF1 (N921, N916);
or OR2 (N922, N921, N653);
or OR3 (N923, N902, N267, N176);
nand NAND3 (N924, N922, N431, N110);
and AND2 (N925, N923, N763);
and AND4 (N926, N911, N646, N401, N191);
not NOT1 (N927, N924);
not NOT1 (N928, N925);
and AND2 (N929, N920, N105);
nor NOR3 (N930, N929, N335, N70);
and AND3 (N931, N927, N194, N166);
or OR2 (N932, N915, N378);
and AND3 (N933, N926, N630, N649);
nor NOR2 (N934, N931, N912);
buf BUF1 (N935, N906);
nor NOR3 (N936, N919, N771, N297);
buf BUF1 (N937, N935);
or OR3 (N938, N879, N214, N324);
or OR4 (N939, N899, N232, N329, N468);
not NOT1 (N940, N932);
nor NOR2 (N941, N936, N612);
not NOT1 (N942, N937);
nor NOR4 (N943, N934, N124, N941, N882);
nor NOR2 (N944, N355, N710);
and AND2 (N945, N928, N383);
xor XOR2 (N946, N939, N777);
xor XOR2 (N947, N945, N114);
and AND3 (N948, N940, N930, N833);
and AND3 (N949, N112, N315, N706);
and AND3 (N950, N948, N703, N832);
xor XOR2 (N951, N946, N936);
nor NOR4 (N952, N951, N402, N99, N805);
nand NAND2 (N953, N949, N598);
xor XOR2 (N954, N953, N866);
or OR2 (N955, N950, N206);
buf BUF1 (N956, N918);
and AND3 (N957, N954, N164, N928);
nand NAND2 (N958, N947, N555);
or OR4 (N959, N955, N915, N400, N3);
or OR4 (N960, N944, N774, N348, N950);
and AND3 (N961, N942, N773, N109);
nor NOR4 (N962, N957, N189, N542, N926);
nand NAND2 (N963, N943, N12);
and AND2 (N964, N960, N433);
nor NOR2 (N965, N964, N911);
and AND2 (N966, N959, N490);
nor NOR4 (N967, N962, N578, N720, N200);
nor NOR4 (N968, N933, N253, N717, N261);
or OR4 (N969, N938, N332, N13, N148);
nor NOR2 (N970, N963, N965);
nand NAND4 (N971, N694, N189, N613, N698);
nor NOR3 (N972, N967, N382, N527);
xor XOR2 (N973, N956, N482);
not NOT1 (N974, N961);
not NOT1 (N975, N952);
xor XOR2 (N976, N974, N224);
buf BUF1 (N977, N971);
buf BUF1 (N978, N966);
nand NAND2 (N979, N968, N212);
not NOT1 (N980, N976);
and AND3 (N981, N977, N479, N8);
and AND3 (N982, N979, N819, N606);
nand NAND4 (N983, N975, N679, N172, N25);
buf BUF1 (N984, N970);
nand NAND4 (N985, N972, N659, N248, N458);
xor XOR2 (N986, N983, N312);
or OR3 (N987, N973, N311, N555);
buf BUF1 (N988, N982);
or OR3 (N989, N978, N309, N484);
or OR3 (N990, N988, N943, N498);
or OR3 (N991, N985, N626, N870);
nor NOR2 (N992, N991, N568);
and AND2 (N993, N969, N207);
or OR3 (N994, N980, N421, N809);
nand NAND2 (N995, N958, N743);
nor NOR2 (N996, N990, N737);
nor NOR4 (N997, N986, N792, N43, N492);
nor NOR4 (N998, N984, N283, N787, N891);
xor XOR2 (N999, N996, N981);
nand NAND3 (N1000, N242, N231, N746);
not NOT1 (N1001, N992);
not NOT1 (N1002, N995);
or OR3 (N1003, N1000, N753, N678);
xor XOR2 (N1004, N999, N869);
xor XOR2 (N1005, N1002, N571);
xor XOR2 (N1006, N1003, N300);
not NOT1 (N1007, N987);
or OR4 (N1008, N998, N93, N920, N288);
not NOT1 (N1009, N994);
or OR2 (N1010, N1008, N813);
nand NAND3 (N1011, N1007, N94, N858);
or OR3 (N1012, N1010, N18, N3);
buf BUF1 (N1013, N1006);
or OR2 (N1014, N1009, N372);
buf BUF1 (N1015, N997);
buf BUF1 (N1016, N989);
nor NOR4 (N1017, N1016, N86, N41, N76);
or OR2 (N1018, N1017, N448);
and AND2 (N1019, N1015, N13);
and AND2 (N1020, N1004, N599);
or OR4 (N1021, N1014, N18, N621, N766);
nand NAND3 (N1022, N1021, N51, N595);
xor XOR2 (N1023, N1011, N307);
or OR2 (N1024, N993, N771);
or OR2 (N1025, N1012, N728);
nor NOR4 (N1026, N1019, N352, N609, N285);
and AND2 (N1027, N1001, N941);
xor XOR2 (N1028, N1005, N549);
buf BUF1 (N1029, N1020);
buf BUF1 (N1030, N1026);
nand NAND3 (N1031, N1023, N963, N325);
xor XOR2 (N1032, N1022, N913);
buf BUF1 (N1033, N1013);
and AND3 (N1034, N1024, N817, N1005);
not NOT1 (N1035, N1025);
not NOT1 (N1036, N1033);
nor NOR3 (N1037, N1034, N365, N751);
and AND2 (N1038, N1036, N874);
nor NOR4 (N1039, N1038, N714, N194, N778);
and AND2 (N1040, N1031, N484);
or OR2 (N1041, N1030, N854);
or OR2 (N1042, N1018, N1002);
buf BUF1 (N1043, N1035);
nand NAND3 (N1044, N1028, N687, N338);
buf BUF1 (N1045, N1040);
xor XOR2 (N1046, N1041, N457);
and AND2 (N1047, N1043, N235);
and AND3 (N1048, N1039, N483, N1022);
buf BUF1 (N1049, N1027);
buf BUF1 (N1050, N1044);
and AND4 (N1051, N1045, N732, N827, N1022);
nand NAND3 (N1052, N1047, N92, N893);
not NOT1 (N1053, N1029);
not NOT1 (N1054, N1053);
nand NAND4 (N1055, N1051, N126, N983, N690);
and AND4 (N1056, N1032, N526, N953, N440);
nand NAND4 (N1057, N1048, N336, N39, N721);
or OR3 (N1058, N1037, N419, N564);
nor NOR2 (N1059, N1058, N311);
or OR3 (N1060, N1056, N1, N928);
nand NAND2 (N1061, N1054, N193);
nor NOR3 (N1062, N1042, N618, N999);
nor NOR3 (N1063, N1055, N506, N902);
not NOT1 (N1064, N1062);
not NOT1 (N1065, N1049);
or OR3 (N1066, N1061, N940, N835);
and AND2 (N1067, N1050, N534);
buf BUF1 (N1068, N1060);
xor XOR2 (N1069, N1063, N63);
not NOT1 (N1070, N1068);
not NOT1 (N1071, N1070);
buf BUF1 (N1072, N1065);
nor NOR2 (N1073, N1069, N434);
buf BUF1 (N1074, N1072);
and AND3 (N1075, N1073, N922, N565);
xor XOR2 (N1076, N1052, N6);
not NOT1 (N1077, N1074);
nand NAND3 (N1078, N1075, N858, N973);
nand NAND4 (N1079, N1057, N523, N852, N722);
not NOT1 (N1080, N1046);
nor NOR4 (N1081, N1059, N1066, N843, N380);
not NOT1 (N1082, N758);
not NOT1 (N1083, N1081);
or OR4 (N1084, N1082, N338, N921, N177);
xor XOR2 (N1085, N1064, N468);
xor XOR2 (N1086, N1078, N140);
or OR2 (N1087, N1086, N121);
nand NAND4 (N1088, N1080, N287, N574, N406);
or OR3 (N1089, N1085, N709, N491);
nand NAND4 (N1090, N1067, N69, N625, N407);
xor XOR2 (N1091, N1090, N559);
buf BUF1 (N1092, N1088);
and AND3 (N1093, N1087, N89, N584);
not NOT1 (N1094, N1084);
and AND3 (N1095, N1079, N300, N164);
nand NAND3 (N1096, N1092, N362, N1056);
buf BUF1 (N1097, N1076);
or OR2 (N1098, N1096, N266);
not NOT1 (N1099, N1094);
nand NAND3 (N1100, N1098, N910, N727);
not NOT1 (N1101, N1083);
not NOT1 (N1102, N1099);
not NOT1 (N1103, N1091);
or OR4 (N1104, N1093, N355, N768, N215);
nand NAND2 (N1105, N1071, N824);
and AND4 (N1106, N1089, N701, N118, N1039);
nand NAND2 (N1107, N1104, N551);
nand NAND4 (N1108, N1095, N893, N827, N689);
buf BUF1 (N1109, N1102);
or OR2 (N1110, N1103, N5);
not NOT1 (N1111, N1097);
nor NOR2 (N1112, N1106, N656);
nor NOR2 (N1113, N1110, N1097);
xor XOR2 (N1114, N1107, N957);
buf BUF1 (N1115, N1111);
nand NAND3 (N1116, N1101, N379, N324);
nand NAND3 (N1117, N1115, N894, N543);
nand NAND4 (N1118, N1113, N355, N850, N481);
nor NOR4 (N1119, N1108, N226, N696, N19);
nand NAND3 (N1120, N1105, N771, N447);
not NOT1 (N1121, N1077);
nor NOR3 (N1122, N1120, N966, N49);
nand NAND2 (N1123, N1116, N1035);
nand NAND3 (N1124, N1114, N495, N558);
not NOT1 (N1125, N1100);
or OR2 (N1126, N1121, N634);
nor NOR4 (N1127, N1119, N160, N155, N993);
nand NAND4 (N1128, N1126, N312, N495, N1040);
and AND2 (N1129, N1109, N168);
nor NOR3 (N1130, N1112, N659, N1112);
nor NOR3 (N1131, N1117, N53, N986);
xor XOR2 (N1132, N1122, N640);
or OR2 (N1133, N1118, N81);
nor NOR4 (N1134, N1127, N863, N252, N713);
or OR4 (N1135, N1123, N88, N13, N755);
xor XOR2 (N1136, N1131, N613);
and AND4 (N1137, N1136, N244, N179, N656);
not NOT1 (N1138, N1130);
or OR2 (N1139, N1129, N740);
nand NAND2 (N1140, N1132, N30);
buf BUF1 (N1141, N1134);
and AND4 (N1142, N1138, N893, N601, N868);
not NOT1 (N1143, N1135);
and AND4 (N1144, N1140, N1019, N135, N1107);
nor NOR2 (N1145, N1144, N830);
nor NOR2 (N1146, N1128, N742);
xor XOR2 (N1147, N1124, N50);
not NOT1 (N1148, N1143);
not NOT1 (N1149, N1146);
buf BUF1 (N1150, N1148);
not NOT1 (N1151, N1149);
and AND3 (N1152, N1150, N720, N511);
xor XOR2 (N1153, N1125, N316);
nand NAND3 (N1154, N1133, N23, N1123);
or OR2 (N1155, N1147, N852);
or OR4 (N1156, N1141, N105, N937, N506);
nand NAND3 (N1157, N1145, N226, N684);
nor NOR4 (N1158, N1152, N1095, N1089, N309);
nand NAND4 (N1159, N1137, N327, N278, N390);
or OR3 (N1160, N1154, N812, N97);
not NOT1 (N1161, N1160);
not NOT1 (N1162, N1158);
not NOT1 (N1163, N1162);
nand NAND3 (N1164, N1153, N514, N274);
and AND3 (N1165, N1161, N994, N315);
xor XOR2 (N1166, N1159, N24);
not NOT1 (N1167, N1156);
nand NAND4 (N1168, N1142, N331, N368, N796);
or OR4 (N1169, N1163, N38, N407, N170);
xor XOR2 (N1170, N1167, N626);
buf BUF1 (N1171, N1166);
or OR3 (N1172, N1171, N172, N515);
or OR4 (N1173, N1139, N1108, N427, N119);
nor NOR4 (N1174, N1169, N510, N1158, N352);
and AND3 (N1175, N1155, N687, N261);
and AND3 (N1176, N1165, N580, N887);
and AND4 (N1177, N1172, N712, N530, N25);
nand NAND3 (N1178, N1168, N161, N781);
and AND2 (N1179, N1178, N383);
xor XOR2 (N1180, N1151, N1068);
nor NOR4 (N1181, N1164, N263, N556, N1180);
nor NOR4 (N1182, N45, N356, N881, N197);
and AND3 (N1183, N1157, N367, N122);
or OR3 (N1184, N1176, N206, N727);
and AND4 (N1185, N1170, N1181, N913, N905);
nand NAND4 (N1186, N16, N931, N86, N513);
buf BUF1 (N1187, N1179);
nand NAND3 (N1188, N1174, N59, N455);
not NOT1 (N1189, N1185);
not NOT1 (N1190, N1182);
or OR4 (N1191, N1189, N380, N513, N848);
nand NAND2 (N1192, N1184, N432);
buf BUF1 (N1193, N1175);
nor NOR3 (N1194, N1193, N539, N434);
xor XOR2 (N1195, N1186, N227);
nand NAND2 (N1196, N1190, N680);
xor XOR2 (N1197, N1191, N1088);
nand NAND3 (N1198, N1197, N401, N393);
not NOT1 (N1199, N1196);
xor XOR2 (N1200, N1192, N1102);
nor NOR3 (N1201, N1195, N826, N103);
and AND4 (N1202, N1187, N948, N413, N810);
nor NOR2 (N1203, N1201, N14);
nor NOR3 (N1204, N1203, N695, N944);
and AND3 (N1205, N1177, N248, N591);
buf BUF1 (N1206, N1173);
and AND2 (N1207, N1188, N330);
or OR4 (N1208, N1198, N1002, N951, N880);
nor NOR2 (N1209, N1205, N154);
nor NOR2 (N1210, N1207, N1196);
nor NOR3 (N1211, N1209, N704, N258);
or OR3 (N1212, N1204, N397, N316);
or OR2 (N1213, N1211, N914);
nor NOR3 (N1214, N1208, N640, N639);
or OR4 (N1215, N1183, N32, N982, N1203);
buf BUF1 (N1216, N1213);
not NOT1 (N1217, N1214);
and AND4 (N1218, N1199, N974, N544, N962);
or OR4 (N1219, N1194, N1209, N840, N1082);
nand NAND3 (N1220, N1216, N548, N940);
buf BUF1 (N1221, N1217);
and AND3 (N1222, N1212, N743, N816);
and AND2 (N1223, N1210, N259);
not NOT1 (N1224, N1215);
not NOT1 (N1225, N1223);
xor XOR2 (N1226, N1202, N1060);
and AND4 (N1227, N1221, N65, N214, N42);
not NOT1 (N1228, N1219);
xor XOR2 (N1229, N1227, N1171);
or OR2 (N1230, N1229, N971);
nor NOR4 (N1231, N1226, N1211, N1011, N1225);
and AND3 (N1232, N346, N494, N1037);
not NOT1 (N1233, N1200);
nand NAND2 (N1234, N1230, N1156);
nand NAND2 (N1235, N1233, N104);
not NOT1 (N1236, N1218);
nand NAND3 (N1237, N1232, N465, N274);
nand NAND3 (N1238, N1234, N659, N551);
nand NAND4 (N1239, N1237, N768, N925, N221);
and AND3 (N1240, N1224, N948, N909);
xor XOR2 (N1241, N1238, N1118);
nor NOR2 (N1242, N1220, N529);
xor XOR2 (N1243, N1236, N952);
or OR4 (N1244, N1206, N457, N1048, N901);
buf BUF1 (N1245, N1222);
nand NAND3 (N1246, N1239, N489, N542);
and AND3 (N1247, N1246, N510, N436);
or OR2 (N1248, N1228, N929);
and AND2 (N1249, N1247, N157);
nor NOR4 (N1250, N1241, N1123, N384, N441);
not NOT1 (N1251, N1242);
and AND2 (N1252, N1248, N150);
buf BUF1 (N1253, N1240);
buf BUF1 (N1254, N1231);
xor XOR2 (N1255, N1243, N41);
and AND2 (N1256, N1251, N1247);
nor NOR3 (N1257, N1255, N468, N603);
buf BUF1 (N1258, N1250);
buf BUF1 (N1259, N1257);
not NOT1 (N1260, N1245);
not NOT1 (N1261, N1244);
buf BUF1 (N1262, N1260);
buf BUF1 (N1263, N1253);
and AND3 (N1264, N1235, N1152, N357);
not NOT1 (N1265, N1264);
and AND4 (N1266, N1262, N1151, N438, N536);
nand NAND3 (N1267, N1261, N467, N535);
nor NOR4 (N1268, N1266, N338, N580, N529);
buf BUF1 (N1269, N1254);
xor XOR2 (N1270, N1269, N133);
and AND2 (N1271, N1268, N177);
xor XOR2 (N1272, N1270, N1040);
not NOT1 (N1273, N1265);
or OR2 (N1274, N1271, N387);
buf BUF1 (N1275, N1274);
and AND2 (N1276, N1252, N66);
nor NOR4 (N1277, N1263, N18, N885, N276);
buf BUF1 (N1278, N1276);
or OR3 (N1279, N1277, N62, N184);
nand NAND3 (N1280, N1259, N1211, N1059);
nor NOR2 (N1281, N1273, N763);
nor NOR2 (N1282, N1279, N939);
xor XOR2 (N1283, N1267, N613);
nor NOR3 (N1284, N1249, N721, N847);
not NOT1 (N1285, N1278);
nand NAND2 (N1286, N1283, N1276);
buf BUF1 (N1287, N1284);
not NOT1 (N1288, N1256);
nor NOR3 (N1289, N1286, N583, N29);
or OR4 (N1290, N1289, N821, N74, N464);
nor NOR4 (N1291, N1288, N464, N280, N407);
not NOT1 (N1292, N1285);
nor NOR2 (N1293, N1272, N1250);
xor XOR2 (N1294, N1287, N261);
buf BUF1 (N1295, N1293);
nor NOR4 (N1296, N1295, N574, N458, N1154);
nor NOR3 (N1297, N1296, N167, N615);
or OR4 (N1298, N1291, N421, N499, N614);
xor XOR2 (N1299, N1298, N896);
xor XOR2 (N1300, N1280, N987);
xor XOR2 (N1301, N1297, N144);
nor NOR4 (N1302, N1292, N57, N967, N926);
nor NOR4 (N1303, N1281, N1191, N909, N132);
xor XOR2 (N1304, N1294, N461);
not NOT1 (N1305, N1275);
not NOT1 (N1306, N1304);
nand NAND3 (N1307, N1300, N901, N426);
nor NOR2 (N1308, N1303, N1251);
xor XOR2 (N1309, N1306, N786);
nor NOR4 (N1310, N1308, N869, N395, N343);
not NOT1 (N1311, N1307);
nor NOR4 (N1312, N1311, N917, N1274, N1055);
or OR2 (N1313, N1310, N804);
and AND4 (N1314, N1258, N298, N224, N175);
not NOT1 (N1315, N1282);
not NOT1 (N1316, N1314);
buf BUF1 (N1317, N1312);
not NOT1 (N1318, N1317);
and AND4 (N1319, N1316, N786, N350, N506);
buf BUF1 (N1320, N1290);
xor XOR2 (N1321, N1313, N1063);
not NOT1 (N1322, N1320);
buf BUF1 (N1323, N1315);
nand NAND4 (N1324, N1299, N1041, N619, N1200);
buf BUF1 (N1325, N1319);
xor XOR2 (N1326, N1324, N211);
and AND4 (N1327, N1309, N700, N442, N535);
not NOT1 (N1328, N1302);
nor NOR4 (N1329, N1326, N1245, N474, N1074);
nand NAND2 (N1330, N1318, N838);
nor NOR4 (N1331, N1323, N32, N983, N845);
buf BUF1 (N1332, N1325);
buf BUF1 (N1333, N1327);
buf BUF1 (N1334, N1329);
buf BUF1 (N1335, N1332);
xor XOR2 (N1336, N1333, N804);
xor XOR2 (N1337, N1328, N129);
not NOT1 (N1338, N1337);
or OR3 (N1339, N1336, N1328, N274);
or OR3 (N1340, N1331, N712, N1091);
or OR3 (N1341, N1338, N121, N949);
and AND2 (N1342, N1334, N414);
xor XOR2 (N1343, N1330, N1012);
nor NOR3 (N1344, N1343, N63, N35);
nand NAND2 (N1345, N1340, N759);
buf BUF1 (N1346, N1345);
nor NOR2 (N1347, N1346, N189);
not NOT1 (N1348, N1335);
or OR4 (N1349, N1348, N520, N425, N364);
nand NAND2 (N1350, N1339, N700);
xor XOR2 (N1351, N1349, N1103);
not NOT1 (N1352, N1351);
buf BUF1 (N1353, N1342);
or OR3 (N1354, N1341, N393, N95);
nor NOR3 (N1355, N1347, N1265, N636);
and AND4 (N1356, N1352, N341, N498, N1021);
xor XOR2 (N1357, N1355, N1205);
buf BUF1 (N1358, N1350);
not NOT1 (N1359, N1344);
or OR4 (N1360, N1357, N593, N992, N525);
xor XOR2 (N1361, N1360, N1174);
not NOT1 (N1362, N1356);
and AND4 (N1363, N1322, N273, N456, N1092);
xor XOR2 (N1364, N1321, N614);
buf BUF1 (N1365, N1358);
and AND3 (N1366, N1301, N1025, N127);
buf BUF1 (N1367, N1363);
not NOT1 (N1368, N1364);
nand NAND4 (N1369, N1362, N1032, N1104, N783);
nand NAND4 (N1370, N1365, N17, N570, N1211);
nand NAND3 (N1371, N1305, N947, N427);
nor NOR2 (N1372, N1367, N686);
or OR2 (N1373, N1359, N540);
nor NOR4 (N1374, N1371, N171, N1227, N1372);
not NOT1 (N1375, N521);
buf BUF1 (N1376, N1370);
or OR3 (N1377, N1368, N760, N756);
and AND3 (N1378, N1373, N123, N364);
xor XOR2 (N1379, N1366, N1360);
not NOT1 (N1380, N1375);
not NOT1 (N1381, N1380);
buf BUF1 (N1382, N1376);
and AND2 (N1383, N1374, N329);
or OR3 (N1384, N1354, N827, N296);
buf BUF1 (N1385, N1377);
xor XOR2 (N1386, N1378, N828);
nor NOR2 (N1387, N1369, N1103);
not NOT1 (N1388, N1382);
xor XOR2 (N1389, N1384, N457);
xor XOR2 (N1390, N1389, N1144);
or OR4 (N1391, N1381, N554, N636, N683);
not NOT1 (N1392, N1385);
and AND2 (N1393, N1388, N674);
or OR2 (N1394, N1391, N199);
or OR3 (N1395, N1379, N570, N82);
not NOT1 (N1396, N1392);
or OR3 (N1397, N1353, N917, N349);
nor NOR2 (N1398, N1393, N494);
nor NOR2 (N1399, N1386, N1303);
nand NAND2 (N1400, N1398, N430);
nor NOR2 (N1401, N1387, N1003);
not NOT1 (N1402, N1401);
xor XOR2 (N1403, N1361, N635);
buf BUF1 (N1404, N1399);
nand NAND2 (N1405, N1397, N1026);
or OR3 (N1406, N1400, N595, N811);
and AND3 (N1407, N1403, N967, N967);
buf BUF1 (N1408, N1394);
xor XOR2 (N1409, N1383, N1255);
and AND3 (N1410, N1409, N645, N1042);
not NOT1 (N1411, N1405);
and AND2 (N1412, N1390, N119);
not NOT1 (N1413, N1412);
nor NOR2 (N1414, N1396, N477);
not NOT1 (N1415, N1408);
nand NAND3 (N1416, N1404, N301, N812);
buf BUF1 (N1417, N1406);
buf BUF1 (N1418, N1416);
xor XOR2 (N1419, N1407, N801);
and AND3 (N1420, N1418, N1381, N824);
buf BUF1 (N1421, N1395);
buf BUF1 (N1422, N1414);
and AND2 (N1423, N1413, N898);
xor XOR2 (N1424, N1410, N42);
or OR2 (N1425, N1424, N1108);
and AND4 (N1426, N1422, N587, N479, N786);
and AND4 (N1427, N1423, N365, N1151, N313);
buf BUF1 (N1428, N1411);
nand NAND2 (N1429, N1421, N815);
buf BUF1 (N1430, N1425);
and AND4 (N1431, N1430, N1310, N447, N904);
xor XOR2 (N1432, N1415, N681);
buf BUF1 (N1433, N1432);
not NOT1 (N1434, N1420);
nor NOR2 (N1435, N1431, N470);
or OR2 (N1436, N1429, N909);
not NOT1 (N1437, N1428);
xor XOR2 (N1438, N1436, N596);
xor XOR2 (N1439, N1427, N588);
and AND4 (N1440, N1438, N1232, N242, N168);
buf BUF1 (N1441, N1440);
buf BUF1 (N1442, N1433);
xor XOR2 (N1443, N1417, N645);
buf BUF1 (N1444, N1443);
not NOT1 (N1445, N1426);
not NOT1 (N1446, N1434);
and AND4 (N1447, N1419, N841, N559, N1165);
nand NAND4 (N1448, N1437, N1358, N1309, N747);
and AND3 (N1449, N1439, N701, N385);
nor NOR3 (N1450, N1445, N578, N815);
buf BUF1 (N1451, N1446);
buf BUF1 (N1452, N1441);
nor NOR2 (N1453, N1452, N1424);
buf BUF1 (N1454, N1450);
and AND3 (N1455, N1448, N731, N998);
not NOT1 (N1456, N1435);
xor XOR2 (N1457, N1444, N154);
buf BUF1 (N1458, N1455);
and AND4 (N1459, N1442, N729, N491, N630);
xor XOR2 (N1460, N1457, N288);
not NOT1 (N1461, N1402);
nor NOR3 (N1462, N1461, N501, N800);
not NOT1 (N1463, N1460);
nand NAND4 (N1464, N1451, N55, N1319, N1362);
nand NAND3 (N1465, N1462, N520, N872);
not NOT1 (N1466, N1456);
xor XOR2 (N1467, N1463, N365);
buf BUF1 (N1468, N1453);
or OR2 (N1469, N1459, N1316);
nor NOR4 (N1470, N1454, N913, N1193, N1399);
not NOT1 (N1471, N1465);
and AND3 (N1472, N1447, N893, N278);
buf BUF1 (N1473, N1468);
or OR4 (N1474, N1466, N1319, N166, N1255);
not NOT1 (N1475, N1470);
nor NOR4 (N1476, N1449, N1140, N550, N1463);
xor XOR2 (N1477, N1473, N444);
and AND3 (N1478, N1467, N63, N791);
buf BUF1 (N1479, N1469);
not NOT1 (N1480, N1476);
or OR2 (N1481, N1458, N1477);
buf BUF1 (N1482, N1071);
xor XOR2 (N1483, N1479, N309);
not NOT1 (N1484, N1474);
not NOT1 (N1485, N1483);
buf BUF1 (N1486, N1482);
and AND4 (N1487, N1480, N616, N944, N918);
nand NAND4 (N1488, N1478, N219, N46, N65);
nor NOR2 (N1489, N1472, N325);
buf BUF1 (N1490, N1471);
not NOT1 (N1491, N1484);
or OR2 (N1492, N1481, N556);
buf BUF1 (N1493, N1491);
or OR2 (N1494, N1492, N645);
xor XOR2 (N1495, N1490, N562);
xor XOR2 (N1496, N1485, N84);
and AND3 (N1497, N1494, N479, N428);
not NOT1 (N1498, N1464);
not NOT1 (N1499, N1497);
nor NOR4 (N1500, N1496, N63, N561, N385);
buf BUF1 (N1501, N1495);
nand NAND3 (N1502, N1475, N651, N187);
buf BUF1 (N1503, N1500);
not NOT1 (N1504, N1498);
xor XOR2 (N1505, N1487, N1006);
buf BUF1 (N1506, N1488);
nand NAND4 (N1507, N1505, N1456, N288, N501);
not NOT1 (N1508, N1486);
and AND3 (N1509, N1506, N470, N1355);
nand NAND4 (N1510, N1489, N1397, N497, N936);
nor NOR2 (N1511, N1499, N533);
and AND4 (N1512, N1504, N1486, N818, N358);
xor XOR2 (N1513, N1502, N257);
buf BUF1 (N1514, N1503);
and AND3 (N1515, N1514, N135, N730);
buf BUF1 (N1516, N1510);
nand NAND4 (N1517, N1516, N1257, N1468, N1228);
nor NOR4 (N1518, N1513, N296, N1489, N971);
or OR3 (N1519, N1508, N689, N163);
or OR2 (N1520, N1512, N622);
nand NAND3 (N1521, N1515, N809, N800);
and AND3 (N1522, N1518, N154, N177);
nand NAND3 (N1523, N1493, N976, N3);
not NOT1 (N1524, N1520);
and AND2 (N1525, N1521, N1262);
and AND2 (N1526, N1501, N103);
or OR4 (N1527, N1526, N60, N1034, N1028);
not NOT1 (N1528, N1524);
and AND4 (N1529, N1527, N877, N379, N590);
or OR4 (N1530, N1525, N1170, N1072, N1052);
and AND4 (N1531, N1519, N743, N1526, N1375);
nand NAND2 (N1532, N1530, N1218);
and AND2 (N1533, N1528, N1062);
and AND3 (N1534, N1532, N785, N1306);
nor NOR3 (N1535, N1522, N243, N1100);
nor NOR2 (N1536, N1511, N103);
not NOT1 (N1537, N1523);
or OR3 (N1538, N1534, N345, N624);
or OR3 (N1539, N1507, N366, N1334);
not NOT1 (N1540, N1529);
buf BUF1 (N1541, N1538);
nand NAND3 (N1542, N1539, N1038, N88);
nor NOR2 (N1543, N1540, N1305);
nand NAND2 (N1544, N1543, N1118);
and AND4 (N1545, N1544, N524, N711, N213);
nand NAND4 (N1546, N1517, N1452, N1335, N1334);
or OR3 (N1547, N1542, N602, N203);
not NOT1 (N1548, N1541);
not NOT1 (N1549, N1535);
nor NOR4 (N1550, N1533, N1428, N842, N845);
nor NOR3 (N1551, N1537, N390, N1);
and AND4 (N1552, N1546, N714, N843, N1339);
nor NOR2 (N1553, N1545, N497);
nand NAND2 (N1554, N1552, N587);
xor XOR2 (N1555, N1550, N937);
nor NOR4 (N1556, N1548, N518, N1187, N855);
nand NAND2 (N1557, N1555, N667);
nand NAND4 (N1558, N1557, N594, N1289, N572);
or OR3 (N1559, N1558, N1508, N323);
xor XOR2 (N1560, N1554, N679);
xor XOR2 (N1561, N1556, N305);
nand NAND4 (N1562, N1559, N116, N954, N296);
xor XOR2 (N1563, N1547, N162);
nor NOR4 (N1564, N1562, N338, N910, N1416);
xor XOR2 (N1565, N1563, N1181);
or OR3 (N1566, N1560, N959, N453);
nor NOR2 (N1567, N1565, N983);
nand NAND3 (N1568, N1561, N286, N1071);
or OR2 (N1569, N1551, N1004);
nor NOR4 (N1570, N1567, N237, N468, N477);
not NOT1 (N1571, N1570);
buf BUF1 (N1572, N1571);
buf BUF1 (N1573, N1572);
buf BUF1 (N1574, N1549);
xor XOR2 (N1575, N1573, N1572);
nand NAND2 (N1576, N1564, N933);
nand NAND2 (N1577, N1574, N930);
xor XOR2 (N1578, N1531, N266);
and AND4 (N1579, N1569, N838, N1370, N613);
or OR3 (N1580, N1576, N1140, N813);
or OR2 (N1581, N1575, N410);
and AND3 (N1582, N1578, N136, N944);
and AND3 (N1583, N1568, N714, N169);
buf BUF1 (N1584, N1553);
not NOT1 (N1585, N1583);
nor NOR4 (N1586, N1581, N818, N782, N550);
buf BUF1 (N1587, N1579);
or OR3 (N1588, N1580, N609, N620);
not NOT1 (N1589, N1577);
nand NAND4 (N1590, N1589, N655, N615, N540);
not NOT1 (N1591, N1584);
xor XOR2 (N1592, N1586, N1186);
buf BUF1 (N1593, N1588);
not NOT1 (N1594, N1591);
nand NAND2 (N1595, N1536, N831);
not NOT1 (N1596, N1594);
nor NOR4 (N1597, N1592, N237, N432, N1114);
or OR3 (N1598, N1509, N1130, N833);
nand NAND2 (N1599, N1585, N151);
nand NAND2 (N1600, N1590, N1218);
or OR2 (N1601, N1595, N35);
not NOT1 (N1602, N1598);
or OR2 (N1603, N1593, N932);
or OR4 (N1604, N1587, N1325, N1147, N1558);
buf BUF1 (N1605, N1597);
nor NOR4 (N1606, N1599, N230, N308, N1348);
buf BUF1 (N1607, N1596);
or OR4 (N1608, N1603, N386, N642, N477);
nor NOR2 (N1609, N1602, N915);
xor XOR2 (N1610, N1608, N1090);
not NOT1 (N1611, N1609);
or OR4 (N1612, N1566, N378, N685, N1473);
nand NAND2 (N1613, N1605, N1019);
and AND2 (N1614, N1582, N134);
nor NOR2 (N1615, N1600, N1531);
not NOT1 (N1616, N1613);
and AND2 (N1617, N1601, N775);
and AND2 (N1618, N1604, N1204);
xor XOR2 (N1619, N1614, N281);
nand NAND2 (N1620, N1611, N1147);
xor XOR2 (N1621, N1620, N179);
or OR3 (N1622, N1607, N869, N904);
nand NAND3 (N1623, N1612, N525, N1456);
buf BUF1 (N1624, N1618);
buf BUF1 (N1625, N1617);
buf BUF1 (N1626, N1610);
not NOT1 (N1627, N1624);
xor XOR2 (N1628, N1625, N1091);
buf BUF1 (N1629, N1616);
buf BUF1 (N1630, N1615);
nor NOR3 (N1631, N1623, N191, N768);
or OR4 (N1632, N1627, N510, N1006, N30);
xor XOR2 (N1633, N1632, N441);
xor XOR2 (N1634, N1630, N815);
xor XOR2 (N1635, N1621, N1066);
xor XOR2 (N1636, N1628, N1044);
and AND4 (N1637, N1619, N1067, N1015, N588);
buf BUF1 (N1638, N1633);
buf BUF1 (N1639, N1606);
or OR4 (N1640, N1635, N775, N303, N304);
not NOT1 (N1641, N1637);
or OR4 (N1642, N1634, N841, N1163, N1313);
not NOT1 (N1643, N1640);
or OR4 (N1644, N1639, N1469, N680, N1216);
and AND3 (N1645, N1626, N331, N1357);
xor XOR2 (N1646, N1644, N446);
xor XOR2 (N1647, N1646, N1603);
nand NAND3 (N1648, N1642, N877, N559);
not NOT1 (N1649, N1631);
nor NOR4 (N1650, N1641, N78, N1084, N408);
not NOT1 (N1651, N1622);
or OR2 (N1652, N1649, N949);
nand NAND3 (N1653, N1648, N577, N85);
not NOT1 (N1654, N1636);
or OR2 (N1655, N1654, N539);
nand NAND2 (N1656, N1629, N1485);
xor XOR2 (N1657, N1652, N1115);
xor XOR2 (N1658, N1647, N778);
buf BUF1 (N1659, N1638);
buf BUF1 (N1660, N1656);
or OR4 (N1661, N1643, N1346, N347, N765);
not NOT1 (N1662, N1645);
and AND3 (N1663, N1659, N1265, N217);
or OR2 (N1664, N1653, N755);
xor XOR2 (N1665, N1655, N336);
xor XOR2 (N1666, N1658, N964);
and AND4 (N1667, N1665, N1445, N1046, N779);
xor XOR2 (N1668, N1660, N1337);
not NOT1 (N1669, N1663);
or OR3 (N1670, N1666, N72, N300);
not NOT1 (N1671, N1667);
xor XOR2 (N1672, N1669, N1545);
nand NAND4 (N1673, N1661, N963, N716, N654);
nand NAND4 (N1674, N1650, N381, N1425, N735);
and AND3 (N1675, N1672, N979, N1253);
xor XOR2 (N1676, N1662, N90);
nor NOR3 (N1677, N1670, N651, N213);
not NOT1 (N1678, N1651);
or OR4 (N1679, N1657, N377, N94, N1420);
nor NOR2 (N1680, N1676, N990);
not NOT1 (N1681, N1668);
nor NOR4 (N1682, N1674, N386, N1249, N1457);
nand NAND4 (N1683, N1679, N1128, N1422, N854);
nand NAND4 (N1684, N1677, N616, N378, N868);
nor NOR2 (N1685, N1682, N824);
xor XOR2 (N1686, N1681, N704);
not NOT1 (N1687, N1686);
nor NOR4 (N1688, N1675, N64, N557, N833);
xor XOR2 (N1689, N1680, N56);
and AND2 (N1690, N1689, N1266);
and AND3 (N1691, N1688, N554, N258);
or OR2 (N1692, N1690, N1153);
nor NOR3 (N1693, N1683, N239, N1107);
nor NOR3 (N1694, N1692, N1535, N565);
or OR3 (N1695, N1685, N317, N690);
or OR3 (N1696, N1671, N885, N1464);
buf BUF1 (N1697, N1664);
or OR2 (N1698, N1694, N1677);
xor XOR2 (N1699, N1678, N245);
and AND2 (N1700, N1693, N550);
nor NOR2 (N1701, N1684, N755);
or OR2 (N1702, N1701, N976);
or OR3 (N1703, N1699, N171, N862);
and AND2 (N1704, N1698, N348);
xor XOR2 (N1705, N1702, N1114);
nand NAND3 (N1706, N1673, N128, N997);
not NOT1 (N1707, N1696);
nand NAND3 (N1708, N1691, N1704, N1548);
xor XOR2 (N1709, N1613, N1068);
or OR2 (N1710, N1709, N559);
nand NAND3 (N1711, N1687, N1147, N1314);
xor XOR2 (N1712, N1705, N1256);
buf BUF1 (N1713, N1697);
xor XOR2 (N1714, N1713, N782);
nand NAND3 (N1715, N1695, N1186, N1378);
buf BUF1 (N1716, N1700);
xor XOR2 (N1717, N1712, N878);
nand NAND3 (N1718, N1706, N1007, N1563);
or OR4 (N1719, N1718, N133, N851, N550);
or OR2 (N1720, N1717, N1388);
not NOT1 (N1721, N1719);
nand NAND3 (N1722, N1720, N914, N1110);
not NOT1 (N1723, N1716);
nor NOR3 (N1724, N1723, N1299, N543);
nand NAND2 (N1725, N1724, N347);
nor NOR4 (N1726, N1710, N411, N1110, N1576);
not NOT1 (N1727, N1707);
and AND3 (N1728, N1722, N972, N1083);
nand NAND4 (N1729, N1725, N1552, N653, N46);
buf BUF1 (N1730, N1715);
buf BUF1 (N1731, N1730);
buf BUF1 (N1732, N1726);
buf BUF1 (N1733, N1708);
and AND2 (N1734, N1729, N1227);
and AND3 (N1735, N1727, N783, N1378);
buf BUF1 (N1736, N1703);
and AND3 (N1737, N1714, N114, N1509);
nand NAND4 (N1738, N1731, N1088, N1695, N675);
and AND2 (N1739, N1728, N111);
nor NOR2 (N1740, N1734, N734);
nand NAND2 (N1741, N1740, N1468);
or OR3 (N1742, N1735, N1650, N1328);
nor NOR2 (N1743, N1739, N1395);
nand NAND2 (N1744, N1743, N256);
nor NOR3 (N1745, N1732, N919, N1495);
and AND3 (N1746, N1744, N459, N1545);
or OR3 (N1747, N1738, N765, N587);
nor NOR4 (N1748, N1741, N805, N1606, N1174);
xor XOR2 (N1749, N1748, N123);
buf BUF1 (N1750, N1746);
nor NOR2 (N1751, N1737, N337);
or OR2 (N1752, N1721, N1308);
xor XOR2 (N1753, N1750, N1287);
nand NAND3 (N1754, N1711, N1520, N1421);
and AND2 (N1755, N1736, N239);
buf BUF1 (N1756, N1747);
buf BUF1 (N1757, N1749);
or OR4 (N1758, N1745, N809, N892, N1385);
buf BUF1 (N1759, N1751);
nor NOR3 (N1760, N1752, N1095, N980);
or OR2 (N1761, N1754, N42);
buf BUF1 (N1762, N1733);
not NOT1 (N1763, N1762);
and AND4 (N1764, N1756, N191, N1756, N96);
not NOT1 (N1765, N1763);
nand NAND4 (N1766, N1758, N962, N604, N1580);
nor NOR2 (N1767, N1760, N886);
or OR2 (N1768, N1753, N1581);
not NOT1 (N1769, N1761);
nor NOR2 (N1770, N1769, N1158);
and AND3 (N1771, N1767, N1375, N1345);
nor NOR4 (N1772, N1759, N555, N290, N635);
or OR4 (N1773, N1772, N1238, N1537, N698);
nand NAND4 (N1774, N1771, N664, N5, N1230);
not NOT1 (N1775, N1773);
buf BUF1 (N1776, N1770);
and AND3 (N1777, N1764, N741, N609);
nand NAND3 (N1778, N1768, N696, N891);
and AND2 (N1779, N1776, N178);
nor NOR3 (N1780, N1765, N1742, N363);
nand NAND2 (N1781, N30, N508);
and AND2 (N1782, N1781, N1156);
not NOT1 (N1783, N1779);
buf BUF1 (N1784, N1757);
not NOT1 (N1785, N1777);
buf BUF1 (N1786, N1774);
xor XOR2 (N1787, N1785, N1000);
nand NAND3 (N1788, N1755, N42, N1328);
nand NAND4 (N1789, N1766, N30, N1058, N1220);
and AND3 (N1790, N1775, N681, N596);
and AND3 (N1791, N1787, N1710, N170);
buf BUF1 (N1792, N1783);
and AND3 (N1793, N1789, N1175, N1590);
nor NOR3 (N1794, N1790, N398, N958);
not NOT1 (N1795, N1780);
and AND3 (N1796, N1788, N1564, N653);
and AND3 (N1797, N1792, N1009, N1157);
nand NAND2 (N1798, N1795, N494);
not NOT1 (N1799, N1784);
not NOT1 (N1800, N1793);
xor XOR2 (N1801, N1797, N259);
nand NAND4 (N1802, N1778, N1794, N299, N702);
nand NAND4 (N1803, N867, N1316, N994, N336);
or OR3 (N1804, N1791, N642, N1105);
and AND4 (N1805, N1804, N22, N1742, N112);
buf BUF1 (N1806, N1800);
and AND3 (N1807, N1806, N521, N376);
not NOT1 (N1808, N1801);
not NOT1 (N1809, N1796);
xor XOR2 (N1810, N1805, N242);
not NOT1 (N1811, N1782);
or OR4 (N1812, N1786, N445, N1139, N569);
not NOT1 (N1813, N1807);
or OR3 (N1814, N1802, N4, N1201);
and AND2 (N1815, N1798, N119);
nand NAND4 (N1816, N1803, N1096, N1259, N110);
buf BUF1 (N1817, N1799);
buf BUF1 (N1818, N1812);
and AND2 (N1819, N1814, N464);
nand NAND2 (N1820, N1817, N586);
and AND4 (N1821, N1815, N90, N602, N528);
xor XOR2 (N1822, N1816, N485);
or OR2 (N1823, N1808, N995);
not NOT1 (N1824, N1813);
nor NOR4 (N1825, N1819, N319, N146, N1360);
or OR2 (N1826, N1825, N293);
xor XOR2 (N1827, N1809, N1385);
nor NOR4 (N1828, N1818, N1620, N1435, N1131);
nor NOR4 (N1829, N1826, N1802, N1736, N358);
xor XOR2 (N1830, N1827, N1213);
nand NAND2 (N1831, N1823, N689);
nor NOR4 (N1832, N1829, N809, N684, N621);
nand NAND3 (N1833, N1824, N1053, N699);
xor XOR2 (N1834, N1831, N1434);
or OR3 (N1835, N1830, N496, N1437);
nand NAND4 (N1836, N1828, N1008, N326, N100);
nor NOR4 (N1837, N1820, N1708, N1637, N819);
or OR4 (N1838, N1822, N910, N1073, N571);
nand NAND3 (N1839, N1838, N416, N888);
xor XOR2 (N1840, N1837, N727);
xor XOR2 (N1841, N1832, N1290);
or OR2 (N1842, N1834, N193);
and AND4 (N1843, N1836, N1330, N229, N997);
and AND2 (N1844, N1841, N1100);
buf BUF1 (N1845, N1840);
xor XOR2 (N1846, N1844, N1619);
or OR3 (N1847, N1842, N830, N1538);
and AND3 (N1848, N1811, N1836, N347);
and AND3 (N1849, N1821, N114, N742);
or OR4 (N1850, N1810, N834, N955, N686);
nor NOR4 (N1851, N1849, N717, N1366, N623);
buf BUF1 (N1852, N1850);
xor XOR2 (N1853, N1848, N259);
nand NAND3 (N1854, N1846, N278, N1331);
nand NAND4 (N1855, N1843, N305, N1323, N1058);
or OR2 (N1856, N1847, N1364);
xor XOR2 (N1857, N1833, N143);
not NOT1 (N1858, N1852);
not NOT1 (N1859, N1845);
not NOT1 (N1860, N1853);
or OR3 (N1861, N1859, N943, N862);
nor NOR3 (N1862, N1857, N1519, N1116);
xor XOR2 (N1863, N1839, N1455);
or OR3 (N1864, N1863, N608, N1861);
buf BUF1 (N1865, N416);
xor XOR2 (N1866, N1865, N514);
nor NOR2 (N1867, N1862, N75);
not NOT1 (N1868, N1835);
or OR4 (N1869, N1868, N636, N77, N1760);
not NOT1 (N1870, N1856);
buf BUF1 (N1871, N1855);
not NOT1 (N1872, N1870);
and AND2 (N1873, N1864, N959);
nor NOR2 (N1874, N1858, N1003);
buf BUF1 (N1875, N1866);
buf BUF1 (N1876, N1873);
nor NOR3 (N1877, N1860, N717, N1055);
nor NOR3 (N1878, N1869, N91, N1660);
xor XOR2 (N1879, N1867, N573);
and AND2 (N1880, N1872, N159);
buf BUF1 (N1881, N1876);
and AND3 (N1882, N1878, N1110, N1146);
xor XOR2 (N1883, N1879, N1029);
nor NOR3 (N1884, N1854, N14, N923);
and AND3 (N1885, N1877, N800, N524);
and AND4 (N1886, N1882, N1186, N1057, N659);
not NOT1 (N1887, N1880);
or OR3 (N1888, N1887, N1591, N1472);
not NOT1 (N1889, N1883);
buf BUF1 (N1890, N1851);
nor NOR4 (N1891, N1886, N1582, N559, N503);
nand NAND3 (N1892, N1874, N282, N39);
or OR2 (N1893, N1888, N339);
xor XOR2 (N1894, N1884, N1730);
xor XOR2 (N1895, N1875, N371);
nor NOR3 (N1896, N1892, N1745, N1741);
xor XOR2 (N1897, N1894, N72);
and AND4 (N1898, N1890, N1879, N255, N1430);
nor NOR4 (N1899, N1898, N1774, N573, N1888);
nand NAND2 (N1900, N1895, N1847);
buf BUF1 (N1901, N1897);
not NOT1 (N1902, N1900);
and AND2 (N1903, N1871, N84);
xor XOR2 (N1904, N1889, N653);
buf BUF1 (N1905, N1891);
or OR4 (N1906, N1902, N1833, N12, N557);
nand NAND3 (N1907, N1896, N620, N1062);
xor XOR2 (N1908, N1885, N119);
xor XOR2 (N1909, N1907, N716);
xor XOR2 (N1910, N1903, N515);
xor XOR2 (N1911, N1893, N266);
and AND3 (N1912, N1906, N1518, N1660);
xor XOR2 (N1913, N1908, N768);
and AND4 (N1914, N1910, N1324, N420, N558);
not NOT1 (N1915, N1881);
nor NOR3 (N1916, N1912, N214, N924);
not NOT1 (N1917, N1905);
buf BUF1 (N1918, N1911);
nor NOR2 (N1919, N1917, N636);
and AND4 (N1920, N1914, N1424, N1499, N702);
nor NOR2 (N1921, N1916, N1817);
or OR3 (N1922, N1919, N24, N645);
not NOT1 (N1923, N1899);
xor XOR2 (N1924, N1909, N1505);
buf BUF1 (N1925, N1921);
xor XOR2 (N1926, N1920, N214);
and AND3 (N1927, N1918, N489, N799);
xor XOR2 (N1928, N1922, N1392);
buf BUF1 (N1929, N1901);
nor NOR2 (N1930, N1923, N1783);
buf BUF1 (N1931, N1913);
or OR3 (N1932, N1915, N1173, N1876);
nor NOR2 (N1933, N1925, N1640);
or OR2 (N1934, N1927, N1375);
not NOT1 (N1935, N1932);
or OR4 (N1936, N1930, N369, N1649, N1844);
xor XOR2 (N1937, N1904, N1223);
not NOT1 (N1938, N1924);
nand NAND3 (N1939, N1934, N1921, N1080);
or OR4 (N1940, N1928, N1213, N405, N1868);
xor XOR2 (N1941, N1937, N1001);
not NOT1 (N1942, N1929);
nand NAND3 (N1943, N1926, N257, N1925);
nand NAND4 (N1944, N1938, N316, N870, N1581);
buf BUF1 (N1945, N1933);
and AND4 (N1946, N1945, N328, N1285, N1198);
nor NOR2 (N1947, N1941, N1449);
xor XOR2 (N1948, N1947, N1929);
nand NAND3 (N1949, N1942, N1470, N1932);
xor XOR2 (N1950, N1946, N449);
or OR2 (N1951, N1950, N1647);
buf BUF1 (N1952, N1944);
nor NOR2 (N1953, N1949, N141);
nor NOR3 (N1954, N1948, N122, N154);
buf BUF1 (N1955, N1951);
and AND4 (N1956, N1955, N520, N1055, N1818);
xor XOR2 (N1957, N1954, N1436);
nor NOR4 (N1958, N1952, N1400, N1051, N850);
buf BUF1 (N1959, N1931);
or OR2 (N1960, N1957, N970);
nor NOR2 (N1961, N1953, N1236);
buf BUF1 (N1962, N1939);
or OR3 (N1963, N1962, N505, N253);
nor NOR2 (N1964, N1940, N1387);
nor NOR4 (N1965, N1956, N1867, N1677, N1417);
xor XOR2 (N1966, N1964, N1355);
nor NOR4 (N1967, N1965, N1531, N1263, N652);
or OR2 (N1968, N1958, N295);
or OR2 (N1969, N1960, N846);
nor NOR3 (N1970, N1943, N492, N1726);
nor NOR3 (N1971, N1963, N529, N165);
and AND4 (N1972, N1970, N1161, N1051, N1177);
not NOT1 (N1973, N1969);
not NOT1 (N1974, N1973);
not NOT1 (N1975, N1966);
nand NAND4 (N1976, N1972, N1893, N1701, N72);
and AND2 (N1977, N1961, N1482);
and AND4 (N1978, N1936, N375, N1361, N332);
not NOT1 (N1979, N1977);
buf BUF1 (N1980, N1959);
xor XOR2 (N1981, N1975, N1082);
nor NOR2 (N1982, N1979, N766);
nand NAND4 (N1983, N1980, N535, N336, N954);
xor XOR2 (N1984, N1981, N1972);
nor NOR3 (N1985, N1967, N557, N234);
and AND4 (N1986, N1935, N1180, N58, N942);
xor XOR2 (N1987, N1978, N788);
nor NOR3 (N1988, N1984, N409, N1887);
or OR2 (N1989, N1986, N384);
buf BUF1 (N1990, N1988);
and AND4 (N1991, N1971, N1113, N770, N79);
not NOT1 (N1992, N1989);
buf BUF1 (N1993, N1987);
and AND4 (N1994, N1990, N755, N416, N1025);
nand NAND4 (N1995, N1993, N1935, N365, N1898);
xor XOR2 (N1996, N1983, N1300);
or OR2 (N1997, N1994, N612);
nand NAND4 (N1998, N1991, N1327, N908, N1016);
not NOT1 (N1999, N1998);
nand NAND2 (N2000, N1974, N237);
xor XOR2 (N2001, N1985, N167);
nand NAND2 (N2002, N1982, N1650);
and AND3 (N2003, N2002, N1306, N1794);
or OR3 (N2004, N1968, N1671, N738);
nand NAND4 (N2005, N1997, N1431, N1443, N839);
not NOT1 (N2006, N2000);
xor XOR2 (N2007, N1992, N51);
xor XOR2 (N2008, N1995, N1447);
nor NOR2 (N2009, N2007, N230);
not NOT1 (N2010, N2001);
or OR2 (N2011, N1999, N1975);
nor NOR3 (N2012, N2003, N841, N356);
or OR3 (N2013, N1996, N1784, N1735);
or OR2 (N2014, N2012, N1290);
nand NAND3 (N2015, N2009, N1603, N129);
buf BUF1 (N2016, N2013);
nor NOR4 (N2017, N2004, N1752, N823, N1442);
nor NOR2 (N2018, N2010, N1817);
xor XOR2 (N2019, N2011, N18);
nand NAND4 (N2020, N2018, N138, N1680, N1625);
or OR3 (N2021, N2014, N922, N642);
nand NAND4 (N2022, N2019, N824, N254, N1089);
buf BUF1 (N2023, N2016);
xor XOR2 (N2024, N2020, N589);
or OR2 (N2025, N2023, N1314);
nand NAND4 (N2026, N2006, N401, N157, N1723);
xor XOR2 (N2027, N2022, N782);
or OR3 (N2028, N2027, N1805, N126);
nand NAND4 (N2029, N2025, N429, N951, N929);
or OR4 (N2030, N2008, N261, N408, N208);
buf BUF1 (N2031, N2017);
not NOT1 (N2032, N2029);
or OR4 (N2033, N2024, N61, N1330, N1607);
buf BUF1 (N2034, N2032);
and AND4 (N2035, N2033, N547, N1706, N687);
nor NOR3 (N2036, N2030, N1209, N338);
or OR4 (N2037, N2036, N1577, N1299, N1676);
buf BUF1 (N2038, N2005);
not NOT1 (N2039, N2037);
or OR3 (N2040, N2038, N558, N261);
and AND3 (N2041, N2021, N1810, N1152);
xor XOR2 (N2042, N2035, N258);
xor XOR2 (N2043, N2042, N612);
or OR2 (N2044, N2040, N994);
nor NOR3 (N2045, N2039, N1168, N1216);
nor NOR2 (N2046, N2015, N1471);
or OR4 (N2047, N1976, N616, N287, N925);
nand NAND3 (N2048, N2028, N615, N784);
nor NOR4 (N2049, N2026, N1755, N375, N1094);
buf BUF1 (N2050, N2046);
or OR3 (N2051, N2043, N2046, N1152);
not NOT1 (N2052, N2041);
or OR3 (N2053, N2050, N1420, N1105);
nand NAND3 (N2054, N2051, N796, N160);
nand NAND3 (N2055, N2054, N207, N758);
or OR4 (N2056, N2052, N841, N877, N1068);
not NOT1 (N2057, N2047);
or OR4 (N2058, N2045, N116, N2018, N342);
buf BUF1 (N2059, N2055);
not NOT1 (N2060, N2056);
nand NAND3 (N2061, N2057, N274, N665);
nand NAND4 (N2062, N2053, N1324, N1582, N1654);
xor XOR2 (N2063, N2060, N593);
xor XOR2 (N2064, N2061, N759);
not NOT1 (N2065, N2064);
buf BUF1 (N2066, N2049);
nand NAND2 (N2067, N2031, N1393);
or OR4 (N2068, N2044, N908, N22, N751);
nor NOR2 (N2069, N2066, N136);
and AND3 (N2070, N2067, N451, N927);
and AND4 (N2071, N2058, N4, N1595, N1387);
and AND2 (N2072, N2034, N701);
xor XOR2 (N2073, N2065, N1848);
not NOT1 (N2074, N2059);
xor XOR2 (N2075, N2048, N1903);
not NOT1 (N2076, N2075);
xor XOR2 (N2077, N2063, N1679);
and AND2 (N2078, N2073, N900);
buf BUF1 (N2079, N2072);
nor NOR2 (N2080, N2077, N729);
xor XOR2 (N2081, N2069, N1836);
buf BUF1 (N2082, N2062);
nand NAND3 (N2083, N2081, N1827, N1674);
nor NOR4 (N2084, N2074, N651, N1439, N1381);
nor NOR2 (N2085, N2071, N156);
not NOT1 (N2086, N2085);
and AND2 (N2087, N2082, N247);
nand NAND2 (N2088, N2078, N359);
buf BUF1 (N2089, N2083);
xor XOR2 (N2090, N2088, N138);
nor NOR3 (N2091, N2079, N87, N1358);
not NOT1 (N2092, N2076);
nor NOR2 (N2093, N2092, N1104);
xor XOR2 (N2094, N2080, N332);
xor XOR2 (N2095, N2068, N1030);
not NOT1 (N2096, N2089);
nor NOR3 (N2097, N2084, N1227, N2021);
or OR4 (N2098, N2097, N576, N1130, N1566);
nand NAND4 (N2099, N2091, N1419, N696, N1416);
not NOT1 (N2100, N2099);
not NOT1 (N2101, N2096);
nand NAND2 (N2102, N2098, N76);
and AND3 (N2103, N2087, N842, N88);
nand NAND2 (N2104, N2095, N947);
buf BUF1 (N2105, N2094);
nand NAND2 (N2106, N2093, N1979);
xor XOR2 (N2107, N2103, N452);
or OR3 (N2108, N2101, N2028, N250);
and AND4 (N2109, N2107, N1203, N681, N1587);
not NOT1 (N2110, N2070);
and AND2 (N2111, N2086, N1618);
nor NOR4 (N2112, N2110, N881, N1096, N1491);
nor NOR2 (N2113, N2104, N1924);
or OR4 (N2114, N2100, N748, N1415, N1454);
nor NOR4 (N2115, N2108, N165, N1821, N1158);
not NOT1 (N2116, N2102);
and AND3 (N2117, N2116, N1039, N1485);
or OR3 (N2118, N2114, N1082, N711);
nand NAND2 (N2119, N2090, N590);
buf BUF1 (N2120, N2115);
and AND2 (N2121, N2118, N170);
nor NOR3 (N2122, N2117, N219, N1372);
or OR4 (N2123, N2122, N1381, N1345, N838);
or OR3 (N2124, N2119, N682, N1000);
nor NOR2 (N2125, N2109, N719);
nand NAND2 (N2126, N2111, N1400);
or OR3 (N2127, N2121, N53, N2106);
and AND2 (N2128, N646, N903);
nand NAND2 (N2129, N2124, N502);
or OR4 (N2130, N2113, N1965, N664, N892);
nand NAND4 (N2131, N2128, N1217, N729, N2016);
nand NAND3 (N2132, N2131, N2063, N449);
nand NAND3 (N2133, N2130, N1320, N1191);
not NOT1 (N2134, N2132);
nor NOR2 (N2135, N2120, N1716);
or OR2 (N2136, N2105, N1848);
xor XOR2 (N2137, N2127, N1577);
xor XOR2 (N2138, N2136, N2095);
nand NAND2 (N2139, N2135, N322);
buf BUF1 (N2140, N2126);
xor XOR2 (N2141, N2123, N1516);
nor NOR2 (N2142, N2133, N1106);
buf BUF1 (N2143, N2129);
nand NAND4 (N2144, N2141, N300, N1106, N1303);
not NOT1 (N2145, N2137);
nor NOR4 (N2146, N2144, N1167, N1321, N1828);
buf BUF1 (N2147, N2139);
not NOT1 (N2148, N2125);
not NOT1 (N2149, N2140);
nand NAND2 (N2150, N2138, N1327);
or OR2 (N2151, N2145, N1544);
not NOT1 (N2152, N2149);
and AND2 (N2153, N2148, N2014);
not NOT1 (N2154, N2146);
and AND2 (N2155, N2142, N1815);
not NOT1 (N2156, N2143);
or OR4 (N2157, N2154, N1246, N493, N57);
or OR2 (N2158, N2152, N1940);
buf BUF1 (N2159, N2155);
buf BUF1 (N2160, N2156);
buf BUF1 (N2161, N2151);
nand NAND3 (N2162, N2157, N636, N366);
not NOT1 (N2163, N2112);
or OR2 (N2164, N2158, N1205);
buf BUF1 (N2165, N2161);
not NOT1 (N2166, N2160);
buf BUF1 (N2167, N2150);
xor XOR2 (N2168, N2159, N1382);
not NOT1 (N2169, N2162);
and AND2 (N2170, N2168, N1777);
nor NOR4 (N2171, N2165, N1463, N1683, N1388);
and AND4 (N2172, N2153, N1062, N1040, N1490);
buf BUF1 (N2173, N2164);
or OR3 (N2174, N2163, N1628, N20);
nand NAND3 (N2175, N2172, N572, N916);
nor NOR4 (N2176, N2166, N778, N895, N6);
nand NAND2 (N2177, N2169, N892);
and AND2 (N2178, N2167, N481);
or OR4 (N2179, N2175, N1226, N712, N1223);
xor XOR2 (N2180, N2178, N1727);
and AND3 (N2181, N2174, N891, N1360);
xor XOR2 (N2182, N2134, N699);
or OR3 (N2183, N2177, N867, N302);
or OR4 (N2184, N2181, N668, N604, N359);
xor XOR2 (N2185, N2180, N1376);
nor NOR2 (N2186, N2185, N433);
and AND4 (N2187, N2186, N1357, N1813, N1301);
or OR4 (N2188, N2147, N1148, N410, N1421);
or OR4 (N2189, N2184, N1604, N1952, N840);
and AND3 (N2190, N2187, N1179, N1174);
not NOT1 (N2191, N2170);
and AND4 (N2192, N2173, N1758, N1383, N1809);
not NOT1 (N2193, N2176);
or OR4 (N2194, N2192, N744, N376, N1567);
buf BUF1 (N2195, N2183);
and AND2 (N2196, N2191, N66);
buf BUF1 (N2197, N2171);
and AND2 (N2198, N2195, N838);
buf BUF1 (N2199, N2193);
nand NAND4 (N2200, N2179, N1608, N527, N1289);
buf BUF1 (N2201, N2197);
or OR3 (N2202, N2188, N662, N2063);
not NOT1 (N2203, N2189);
nor NOR4 (N2204, N2196, N2144, N255, N979);
and AND3 (N2205, N2182, N491, N1309);
buf BUF1 (N2206, N2198);
nor NOR2 (N2207, N2199, N132);
nor NOR2 (N2208, N2190, N1458);
xor XOR2 (N2209, N2203, N1088);
not NOT1 (N2210, N2201);
or OR3 (N2211, N2210, N234, N1612);
or OR2 (N2212, N2204, N25);
buf BUF1 (N2213, N2200);
nand NAND4 (N2214, N2202, N574, N283, N1872);
buf BUF1 (N2215, N2214);
nor NOR2 (N2216, N2215, N966);
xor XOR2 (N2217, N2205, N716);
buf BUF1 (N2218, N2194);
not NOT1 (N2219, N2207);
nor NOR3 (N2220, N2216, N918, N2218);
nand NAND3 (N2221, N1336, N1851, N1881);
xor XOR2 (N2222, N2213, N1433);
xor XOR2 (N2223, N2208, N2186);
nor NOR3 (N2224, N2212, N94, N1365);
nor NOR2 (N2225, N2209, N177);
not NOT1 (N2226, N2223);
not NOT1 (N2227, N2226);
or OR3 (N2228, N2219, N1003, N1710);
nor NOR3 (N2229, N2221, N2076, N120);
not NOT1 (N2230, N2227);
buf BUF1 (N2231, N2217);
nand NAND3 (N2232, N2211, N2176, N120);
nand NAND3 (N2233, N2230, N1632, N1016);
not NOT1 (N2234, N2222);
and AND4 (N2235, N2233, N371, N1931, N621);
xor XOR2 (N2236, N2229, N1502);
not NOT1 (N2237, N2220);
buf BUF1 (N2238, N2234);
buf BUF1 (N2239, N2236);
or OR4 (N2240, N2225, N1326, N1606, N1665);
or OR4 (N2241, N2239, N418, N1164, N907);
buf BUF1 (N2242, N2228);
buf BUF1 (N2243, N2206);
buf BUF1 (N2244, N2231);
nor NOR2 (N2245, N2237, N497);
nand NAND3 (N2246, N2235, N395, N1990);
not NOT1 (N2247, N2246);
buf BUF1 (N2248, N2247);
nand NAND3 (N2249, N2232, N2241, N300);
buf BUF1 (N2250, N1940);
nor NOR3 (N2251, N2243, N412, N1546);
or OR2 (N2252, N2240, N207);
and AND3 (N2253, N2245, N209, N2025);
not NOT1 (N2254, N2253);
not NOT1 (N2255, N2252);
not NOT1 (N2256, N2255);
and AND4 (N2257, N2248, N1142, N1911, N1790);
xor XOR2 (N2258, N2224, N435);
xor XOR2 (N2259, N2251, N226);
nor NOR2 (N2260, N2259, N63);
and AND2 (N2261, N2244, N581);
nor NOR4 (N2262, N2238, N1753, N208, N1850);
xor XOR2 (N2263, N2249, N2056);
nand NAND3 (N2264, N2250, N1585, N686);
or OR2 (N2265, N2264, N828);
nand NAND2 (N2266, N2262, N2254);
or OR2 (N2267, N405, N1342);
and AND3 (N2268, N2263, N1716, N241);
buf BUF1 (N2269, N2242);
nor NOR4 (N2270, N2266, N2141, N1003, N607);
and AND4 (N2271, N2261, N1694, N2075, N292);
nand NAND4 (N2272, N2267, N1976, N1929, N288);
nor NOR2 (N2273, N2260, N1429);
xor XOR2 (N2274, N2258, N72);
or OR4 (N2275, N2271, N1604, N1901, N457);
nand NAND3 (N2276, N2265, N2048, N1648);
or OR2 (N2277, N2269, N1242);
not NOT1 (N2278, N2274);
and AND3 (N2279, N2273, N1463, N1732);
nor NOR2 (N2280, N2276, N2120);
not NOT1 (N2281, N2280);
xor XOR2 (N2282, N2270, N381);
buf BUF1 (N2283, N2281);
buf BUF1 (N2284, N2268);
and AND2 (N2285, N2282, N1216);
not NOT1 (N2286, N2285);
nand NAND3 (N2287, N2277, N922, N1104);
or OR4 (N2288, N2287, N1647, N367, N641);
xor XOR2 (N2289, N2283, N632);
nand NAND2 (N2290, N2284, N491);
not NOT1 (N2291, N2289);
nand NAND3 (N2292, N2290, N447, N479);
buf BUF1 (N2293, N2256);
nand NAND2 (N2294, N2257, N1582);
xor XOR2 (N2295, N2293, N2010);
or OR2 (N2296, N2278, N1042);
not NOT1 (N2297, N2296);
not NOT1 (N2298, N2279);
and AND3 (N2299, N2295, N341, N662);
nand NAND2 (N2300, N2275, N590);
and AND2 (N2301, N2298, N1122);
nand NAND2 (N2302, N2291, N2203);
buf BUF1 (N2303, N2302);
or OR2 (N2304, N2288, N789);
nor NOR3 (N2305, N2297, N1086, N1298);
buf BUF1 (N2306, N2286);
buf BUF1 (N2307, N2292);
not NOT1 (N2308, N2307);
xor XOR2 (N2309, N2301, N1926);
or OR2 (N2310, N2308, N1433);
buf BUF1 (N2311, N2306);
not NOT1 (N2312, N2303);
and AND2 (N2313, N2272, N1233);
or OR4 (N2314, N2313, N1247, N1572, N1603);
and AND4 (N2315, N2305, N1252, N1542, N1967);
or OR2 (N2316, N2299, N832);
xor XOR2 (N2317, N2316, N706);
or OR2 (N2318, N2311, N1770);
nor NOR4 (N2319, N2314, N2232, N1513, N2161);
xor XOR2 (N2320, N2312, N28);
not NOT1 (N2321, N2320);
and AND4 (N2322, N2300, N655, N170, N1135);
and AND4 (N2323, N2321, N840, N1100, N782);
or OR3 (N2324, N2323, N1773, N444);
nand NAND2 (N2325, N2322, N2093);
and AND4 (N2326, N2309, N1509, N427, N1284);
buf BUF1 (N2327, N2325);
not NOT1 (N2328, N2317);
and AND2 (N2329, N2310, N143);
and AND4 (N2330, N2327, N771, N2313, N1836);
nand NAND3 (N2331, N2330, N824, N2179);
nor NOR2 (N2332, N2326, N1346);
and AND2 (N2333, N2319, N1974);
and AND4 (N2334, N2332, N215, N804, N964);
not NOT1 (N2335, N2333);
nand NAND2 (N2336, N2315, N818);
nor NOR4 (N2337, N2331, N824, N1175, N634);
buf BUF1 (N2338, N2318);
and AND3 (N2339, N2337, N1704, N1750);
xor XOR2 (N2340, N2334, N366);
or OR3 (N2341, N2329, N237, N2113);
buf BUF1 (N2342, N2340);
and AND2 (N2343, N2336, N981);
nand NAND4 (N2344, N2343, N2181, N285, N2160);
or OR2 (N2345, N2324, N1995);
xor XOR2 (N2346, N2339, N2189);
not NOT1 (N2347, N2345);
or OR3 (N2348, N2344, N1131, N1225);
or OR3 (N2349, N2338, N342, N1455);
or OR2 (N2350, N2348, N1410);
buf BUF1 (N2351, N2328);
not NOT1 (N2352, N2349);
and AND4 (N2353, N2335, N675, N1235, N2078);
nand NAND4 (N2354, N2352, N184, N386, N1848);
and AND2 (N2355, N2341, N1786);
not NOT1 (N2356, N2354);
nor NOR4 (N2357, N2304, N2076, N2337, N1922);
or OR3 (N2358, N2350, N1557, N361);
nand NAND4 (N2359, N2347, N2048, N1551, N157);
or OR4 (N2360, N2359, N774, N795, N595);
nor NOR2 (N2361, N2358, N1933);
and AND3 (N2362, N2355, N1035, N1086);
nand NAND4 (N2363, N2294, N1710, N2243, N1703);
buf BUF1 (N2364, N2361);
or OR2 (N2365, N2360, N1854);
nand NAND2 (N2366, N2357, N1493);
and AND2 (N2367, N2362, N750);
xor XOR2 (N2368, N2342, N1852);
nand NAND2 (N2369, N2367, N2310);
xor XOR2 (N2370, N2366, N479);
buf BUF1 (N2371, N2363);
xor XOR2 (N2372, N2371, N38);
xor XOR2 (N2373, N2370, N1850);
xor XOR2 (N2374, N2346, N1166);
nand NAND3 (N2375, N2356, N1233, N256);
nand NAND3 (N2376, N2374, N2211, N2154);
nor NOR4 (N2377, N2376, N1832, N947, N412);
or OR2 (N2378, N2375, N1831);
or OR2 (N2379, N2377, N537);
buf BUF1 (N2380, N2351);
or OR3 (N2381, N2372, N210, N2101);
buf BUF1 (N2382, N2364);
not NOT1 (N2383, N2373);
not NOT1 (N2384, N2383);
and AND3 (N2385, N2384, N797, N237);
xor XOR2 (N2386, N2385, N1198);
buf BUF1 (N2387, N2369);
and AND3 (N2388, N2368, N2088, N884);
buf BUF1 (N2389, N2380);
nand NAND4 (N2390, N2378, N1305, N10, N1730);
nand NAND3 (N2391, N2386, N806, N2356);
and AND3 (N2392, N2381, N334, N502);
nor NOR3 (N2393, N2353, N633, N277);
not NOT1 (N2394, N2390);
xor XOR2 (N2395, N2392, N1139);
xor XOR2 (N2396, N2391, N888);
buf BUF1 (N2397, N2394);
nor NOR4 (N2398, N2387, N1917, N222, N951);
or OR3 (N2399, N2379, N716, N137);
buf BUF1 (N2400, N2388);
xor XOR2 (N2401, N2382, N992);
nand NAND3 (N2402, N2396, N15, N849);
or OR2 (N2403, N2401, N2350);
xor XOR2 (N2404, N2389, N1352);
or OR4 (N2405, N2398, N1217, N1963, N1600);
and AND3 (N2406, N2403, N584, N1629);
nand NAND2 (N2407, N2395, N891);
buf BUF1 (N2408, N2405);
buf BUF1 (N2409, N2397);
and AND4 (N2410, N2407, N100, N1578, N1100);
buf BUF1 (N2411, N2409);
not NOT1 (N2412, N2399);
or OR2 (N2413, N2406, N681);
nand NAND4 (N2414, N2393, N2119, N1442, N101);
not NOT1 (N2415, N2413);
nor NOR2 (N2416, N2365, N732);
nand NAND3 (N2417, N2402, N1528, N542);
nor NOR4 (N2418, N2414, N234, N1737, N1029);
not NOT1 (N2419, N2400);
buf BUF1 (N2420, N2412);
nand NAND4 (N2421, N2408, N2045, N311, N867);
and AND4 (N2422, N2411, N802, N864, N1563);
not NOT1 (N2423, N2418);
not NOT1 (N2424, N2423);
nand NAND3 (N2425, N2417, N581, N1609);
and AND4 (N2426, N2404, N1261, N1048, N1964);
buf BUF1 (N2427, N2422);
buf BUF1 (N2428, N2421);
buf BUF1 (N2429, N2420);
and AND4 (N2430, N2419, N371, N1727, N1447);
not NOT1 (N2431, N2426);
or OR3 (N2432, N2415, N1, N2243);
xor XOR2 (N2433, N2429, N611);
xor XOR2 (N2434, N2416, N2292);
buf BUF1 (N2435, N2431);
buf BUF1 (N2436, N2427);
nand NAND2 (N2437, N2435, N503);
nand NAND3 (N2438, N2433, N665, N151);
not NOT1 (N2439, N2410);
buf BUF1 (N2440, N2438);
buf BUF1 (N2441, N2437);
not NOT1 (N2442, N2425);
nand NAND2 (N2443, N2441, N601);
nand NAND4 (N2444, N2428, N956, N544, N372);
nor NOR3 (N2445, N2439, N1246, N757);
not NOT1 (N2446, N2443);
nand NAND2 (N2447, N2424, N1912);
xor XOR2 (N2448, N2447, N1426);
not NOT1 (N2449, N2444);
and AND2 (N2450, N2430, N1439);
and AND2 (N2451, N2434, N1965);
or OR2 (N2452, N2446, N335);
nand NAND3 (N2453, N2442, N630, N972);
nand NAND4 (N2454, N2440, N2151, N475, N858);
buf BUF1 (N2455, N2436);
and AND3 (N2456, N2455, N778, N1134);
buf BUF1 (N2457, N2432);
xor XOR2 (N2458, N2448, N1451);
or OR2 (N2459, N2453, N2037);
xor XOR2 (N2460, N2457, N179);
or OR3 (N2461, N2454, N43, N532);
not NOT1 (N2462, N2449);
nand NAND2 (N2463, N2451, N728);
or OR4 (N2464, N2458, N1602, N86, N17);
nor NOR3 (N2465, N2459, N1175, N1370);
xor XOR2 (N2466, N2452, N155);
or OR3 (N2467, N2464, N1211, N1522);
or OR2 (N2468, N2467, N729);
nor NOR4 (N2469, N2463, N225, N1948, N1671);
not NOT1 (N2470, N2466);
buf BUF1 (N2471, N2456);
not NOT1 (N2472, N2460);
or OR2 (N2473, N2461, N321);
nor NOR4 (N2474, N2472, N1610, N1188, N1251);
and AND2 (N2475, N2471, N2113);
and AND3 (N2476, N2469, N2263, N1712);
buf BUF1 (N2477, N2445);
or OR2 (N2478, N2476, N2205);
nand NAND2 (N2479, N2474, N131);
not NOT1 (N2480, N2465);
xor XOR2 (N2481, N2468, N2361);
buf BUF1 (N2482, N2450);
xor XOR2 (N2483, N2478, N188);
or OR3 (N2484, N2483, N157, N348);
or OR2 (N2485, N2480, N2189);
nand NAND4 (N2486, N2462, N828, N351, N2476);
not NOT1 (N2487, N2475);
or OR2 (N2488, N2485, N2140);
buf BUF1 (N2489, N2477);
nor NOR4 (N2490, N2489, N353, N1693, N1641);
or OR4 (N2491, N2479, N1073, N699, N804);
nor NOR4 (N2492, N2491, N1024, N693, N1512);
and AND2 (N2493, N2484, N195);
xor XOR2 (N2494, N2470, N590);
xor XOR2 (N2495, N2482, N2062);
not NOT1 (N2496, N2490);
nor NOR4 (N2497, N2494, N2163, N1526, N842);
not NOT1 (N2498, N2492);
nand NAND4 (N2499, N2498, N506, N436, N1902);
and AND4 (N2500, N2495, N1101, N1982, N898);
nand NAND3 (N2501, N2487, N69, N230);
and AND4 (N2502, N2488, N756, N750, N2178);
xor XOR2 (N2503, N2473, N1062);
nor NOR4 (N2504, N2486, N1018, N48, N2401);
and AND3 (N2505, N2504, N2307, N1787);
and AND3 (N2506, N2497, N966, N2195);
not NOT1 (N2507, N2505);
buf BUF1 (N2508, N2493);
and AND3 (N2509, N2503, N1370, N1703);
or OR3 (N2510, N2501, N2211, N269);
or OR3 (N2511, N2507, N1237, N2306);
and AND4 (N2512, N2508, N1279, N853, N561);
buf BUF1 (N2513, N2511);
or OR2 (N2514, N2506, N1255);
buf BUF1 (N2515, N2502);
buf BUF1 (N2516, N2481);
nor NOR3 (N2517, N2500, N2472, N1745);
buf BUF1 (N2518, N2516);
and AND2 (N2519, N2499, N1734);
and AND4 (N2520, N2512, N1136, N1324, N1424);
xor XOR2 (N2521, N2513, N1672);
nand NAND3 (N2522, N2514, N699, N2460);
nand NAND2 (N2523, N2509, N942);
xor XOR2 (N2524, N2519, N2218);
or OR4 (N2525, N2522, N2225, N2099, N805);
nand NAND4 (N2526, N2515, N1479, N1409, N432);
nand NAND3 (N2527, N2510, N2225, N1301);
and AND3 (N2528, N2525, N146, N602);
and AND3 (N2529, N2527, N261, N1876);
buf BUF1 (N2530, N2529);
xor XOR2 (N2531, N2521, N941);
or OR2 (N2532, N2518, N1705);
and AND4 (N2533, N2530, N1544, N2177, N1992);
buf BUF1 (N2534, N2496);
and AND3 (N2535, N2531, N2485, N693);
xor XOR2 (N2536, N2532, N2255);
xor XOR2 (N2537, N2517, N1919);
not NOT1 (N2538, N2528);
not NOT1 (N2539, N2535);
and AND3 (N2540, N2534, N386, N2164);
nand NAND4 (N2541, N2524, N1183, N2479, N1944);
or OR3 (N2542, N2523, N1151, N911);
buf BUF1 (N2543, N2526);
nor NOR4 (N2544, N2536, N1120, N1342, N964);
or OR3 (N2545, N2538, N1248, N1599);
nor NOR4 (N2546, N2541, N1824, N1081, N367);
not NOT1 (N2547, N2520);
nor NOR2 (N2548, N2537, N718);
nand NAND2 (N2549, N2539, N541);
buf BUF1 (N2550, N2549);
or OR3 (N2551, N2547, N837, N2143);
nor NOR3 (N2552, N2548, N2242, N1058);
not NOT1 (N2553, N2543);
and AND2 (N2554, N2550, N2392);
buf BUF1 (N2555, N2551);
nand NAND2 (N2556, N2554, N2438);
buf BUF1 (N2557, N2552);
or OR2 (N2558, N2546, N317);
xor XOR2 (N2559, N2557, N2124);
nor NOR3 (N2560, N2556, N1526, N1388);
or OR4 (N2561, N2555, N1360, N107, N447);
and AND4 (N2562, N2544, N2246, N1149, N2478);
nor NOR3 (N2563, N2560, N982, N609);
nand NAND3 (N2564, N2540, N1914, N37);
nand NAND3 (N2565, N2561, N824, N1054);
nor NOR3 (N2566, N2533, N2241, N2021);
buf BUF1 (N2567, N2566);
and AND2 (N2568, N2564, N2441);
nor NOR3 (N2569, N2558, N234, N300);
nor NOR4 (N2570, N2563, N170, N1640, N901);
nand NAND4 (N2571, N2559, N712, N74, N1406);
not NOT1 (N2572, N2545);
xor XOR2 (N2573, N2562, N1328);
not NOT1 (N2574, N2565);
xor XOR2 (N2575, N2569, N968);
xor XOR2 (N2576, N2575, N2448);
and AND4 (N2577, N2576, N2108, N1936, N748);
and AND3 (N2578, N2567, N405, N1550);
not NOT1 (N2579, N2542);
nand NAND2 (N2580, N2577, N2239);
buf BUF1 (N2581, N2568);
buf BUF1 (N2582, N2580);
nor NOR2 (N2583, N2579, N816);
nor NOR4 (N2584, N2581, N1202, N782, N1913);
and AND3 (N2585, N2584, N430, N1081);
nor NOR3 (N2586, N2570, N413, N2382);
xor XOR2 (N2587, N2574, N908);
xor XOR2 (N2588, N2586, N583);
xor XOR2 (N2589, N2582, N1329);
xor XOR2 (N2590, N2578, N523);
buf BUF1 (N2591, N2589);
xor XOR2 (N2592, N2571, N2550);
or OR2 (N2593, N2592, N136);
nor NOR3 (N2594, N2583, N2493, N655);
or OR3 (N2595, N2572, N1320, N979);
nor NOR4 (N2596, N2594, N2017, N779, N1815);
xor XOR2 (N2597, N2596, N557);
nand NAND3 (N2598, N2587, N1462, N2480);
xor XOR2 (N2599, N2595, N646);
or OR3 (N2600, N2599, N1285, N1680);
nor NOR2 (N2601, N2590, N2337);
xor XOR2 (N2602, N2588, N55);
nand NAND4 (N2603, N2602, N48, N1821, N2031);
xor XOR2 (N2604, N2591, N2337);
and AND3 (N2605, N2601, N2184, N606);
xor XOR2 (N2606, N2605, N2027);
xor XOR2 (N2607, N2593, N2294);
not NOT1 (N2608, N2604);
not NOT1 (N2609, N2603);
or OR3 (N2610, N2607, N2099, N1453);
nor NOR4 (N2611, N2573, N1252, N1487, N1998);
nand NAND3 (N2612, N2610, N1077, N1565);
nand NAND3 (N2613, N2600, N2160, N2088);
and AND4 (N2614, N2606, N2191, N270, N930);
not NOT1 (N2615, N2553);
and AND4 (N2616, N2614, N1517, N10, N1986);
not NOT1 (N2617, N2585);
not NOT1 (N2618, N2615);
xor XOR2 (N2619, N2617, N1950);
and AND2 (N2620, N2597, N320);
buf BUF1 (N2621, N2620);
and AND3 (N2622, N2612, N1690, N16);
and AND4 (N2623, N2619, N2395, N1462, N1137);
xor XOR2 (N2624, N2618, N168);
xor XOR2 (N2625, N2624, N1565);
nand NAND2 (N2626, N2611, N2360);
nand NAND3 (N2627, N2598, N1297, N2614);
nor NOR3 (N2628, N2622, N1943, N279);
xor XOR2 (N2629, N2621, N2347);
xor XOR2 (N2630, N2609, N422);
buf BUF1 (N2631, N2628);
buf BUF1 (N2632, N2625);
nor NOR3 (N2633, N2608, N107, N2143);
or OR3 (N2634, N2633, N2340, N35);
nor NOR2 (N2635, N2626, N1183);
xor XOR2 (N2636, N2630, N597);
nor NOR2 (N2637, N2636, N341);
and AND3 (N2638, N2637, N2042, N1465);
buf BUF1 (N2639, N2616);
not NOT1 (N2640, N2627);
xor XOR2 (N2641, N2640, N2288);
nor NOR2 (N2642, N2629, N1522);
nor NOR3 (N2643, N2623, N896, N1376);
not NOT1 (N2644, N2643);
xor XOR2 (N2645, N2631, N1949);
buf BUF1 (N2646, N2642);
nand NAND2 (N2647, N2639, N2467);
buf BUF1 (N2648, N2647);
buf BUF1 (N2649, N2641);
xor XOR2 (N2650, N2649, N772);
or OR3 (N2651, N2632, N968, N1302);
nand NAND3 (N2652, N2645, N666, N1017);
or OR4 (N2653, N2635, N148, N2329, N1963);
nor NOR3 (N2654, N2650, N203, N1824);
buf BUF1 (N2655, N2654);
not NOT1 (N2656, N2638);
buf BUF1 (N2657, N2644);
nand NAND2 (N2658, N2646, N1222);
buf BUF1 (N2659, N2651);
or OR4 (N2660, N2648, N185, N2020, N418);
xor XOR2 (N2661, N2656, N1040);
and AND4 (N2662, N2659, N800, N2225, N396);
xor XOR2 (N2663, N2634, N1710);
not NOT1 (N2664, N2658);
buf BUF1 (N2665, N2653);
nor NOR4 (N2666, N2613, N1302, N2291, N1056);
xor XOR2 (N2667, N2664, N1203);
xor XOR2 (N2668, N2667, N195);
or OR4 (N2669, N2661, N2169, N2445, N1001);
xor XOR2 (N2670, N2655, N96);
not NOT1 (N2671, N2669);
nand NAND4 (N2672, N2668, N662, N543, N2488);
nor NOR2 (N2673, N2666, N1450);
buf BUF1 (N2674, N2670);
not NOT1 (N2675, N2652);
xor XOR2 (N2676, N2673, N233);
xor XOR2 (N2677, N2675, N1011);
nor NOR3 (N2678, N2660, N2663, N2020);
nand NAND4 (N2679, N2660, N513, N828, N1686);
not NOT1 (N2680, N2678);
or OR3 (N2681, N2677, N1237, N2604);
nand NAND4 (N2682, N2674, N1875, N2447, N682);
nand NAND3 (N2683, N2676, N561, N1450);
xor XOR2 (N2684, N2681, N87);
nor NOR2 (N2685, N2680, N1888);
nor NOR2 (N2686, N2684, N61);
and AND4 (N2687, N2682, N1817, N2464, N2085);
and AND3 (N2688, N2679, N1419, N1006);
buf BUF1 (N2689, N2683);
or OR4 (N2690, N2686, N975, N305, N1477);
and AND3 (N2691, N2689, N1422, N1404);
nand NAND3 (N2692, N2662, N1947, N142);
xor XOR2 (N2693, N2688, N1398);
xor XOR2 (N2694, N2693, N2026);
buf BUF1 (N2695, N2657);
nand NAND2 (N2696, N2665, N77);
and AND2 (N2697, N2671, N143);
nor NOR4 (N2698, N2690, N662, N1454, N1741);
xor XOR2 (N2699, N2692, N2182);
xor XOR2 (N2700, N2699, N2103);
buf BUF1 (N2701, N2698);
buf BUF1 (N2702, N2695);
buf BUF1 (N2703, N2696);
buf BUF1 (N2704, N2672);
not NOT1 (N2705, N2687);
nand NAND2 (N2706, N2691, N2691);
xor XOR2 (N2707, N2697, N2351);
or OR2 (N2708, N2707, N2470);
nand NAND3 (N2709, N2694, N2544, N1567);
buf BUF1 (N2710, N2702);
or OR2 (N2711, N2705, N1296);
or OR2 (N2712, N2701, N560);
nand NAND3 (N2713, N2710, N1662, N2544);
xor XOR2 (N2714, N2706, N2494);
buf BUF1 (N2715, N2700);
xor XOR2 (N2716, N2714, N2177);
not NOT1 (N2717, N2685);
buf BUF1 (N2718, N2709);
nand NAND3 (N2719, N2713, N2155, N773);
nor NOR4 (N2720, N2716, N885, N2291, N1199);
not NOT1 (N2721, N2720);
buf BUF1 (N2722, N2715);
not NOT1 (N2723, N2704);
and AND2 (N2724, N2722, N1743);
buf BUF1 (N2725, N2712);
nor NOR3 (N2726, N2723, N1986, N973);
nand NAND3 (N2727, N2725, N1296, N1014);
buf BUF1 (N2728, N2721);
xor XOR2 (N2729, N2718, N1763);
nand NAND3 (N2730, N2703, N484, N1664);
xor XOR2 (N2731, N2711, N1641);
or OR3 (N2732, N2708, N1671, N1063);
or OR3 (N2733, N2729, N2051, N1066);
nand NAND2 (N2734, N2717, N1696);
and AND3 (N2735, N2728, N2334, N95);
nor NOR2 (N2736, N2735, N283);
or OR2 (N2737, N2733, N1423);
buf BUF1 (N2738, N2736);
not NOT1 (N2739, N2727);
or OR4 (N2740, N2724, N1524, N1656, N77);
nand NAND3 (N2741, N2732, N138, N687);
not NOT1 (N2742, N2739);
not NOT1 (N2743, N2742);
nand NAND4 (N2744, N2741, N1, N2585, N1351);
nor NOR2 (N2745, N2738, N1835);
or OR2 (N2746, N2726, N1174);
xor XOR2 (N2747, N2737, N2073);
nand NAND3 (N2748, N2731, N11, N806);
or OR3 (N2749, N2740, N87, N450);
or OR4 (N2750, N2745, N2452, N517, N583);
nor NOR3 (N2751, N2734, N763, N1680);
nor NOR2 (N2752, N2749, N353);
buf BUF1 (N2753, N2730);
buf BUF1 (N2754, N2746);
nand NAND2 (N2755, N2719, N2595);
and AND2 (N2756, N2748, N1686);
nand NAND4 (N2757, N2750, N1108, N1256, N686);
or OR2 (N2758, N2744, N87);
not NOT1 (N2759, N2757);
nor NOR2 (N2760, N2759, N2375);
nor NOR3 (N2761, N2760, N1752, N2003);
or OR4 (N2762, N2743, N2095, N2042, N1961);
and AND3 (N2763, N2761, N63, N435);
nand NAND2 (N2764, N2754, N1881);
xor XOR2 (N2765, N2752, N2052);
nor NOR2 (N2766, N2753, N907);
or OR2 (N2767, N2764, N1203);
or OR3 (N2768, N2763, N2283, N87);
or OR4 (N2769, N2768, N2346, N862, N762);
xor XOR2 (N2770, N2758, N2720);
nand NAND3 (N2771, N2751, N2384, N1215);
nor NOR2 (N2772, N2769, N841);
not NOT1 (N2773, N2747);
not NOT1 (N2774, N2762);
buf BUF1 (N2775, N2765);
nor NOR2 (N2776, N2767, N242);
not NOT1 (N2777, N2772);
xor XOR2 (N2778, N2776, N637);
nor NOR4 (N2779, N2756, N2398, N1611, N1872);
buf BUF1 (N2780, N2766);
nor NOR2 (N2781, N2777, N603);
xor XOR2 (N2782, N2755, N2054);
nand NAND2 (N2783, N2782, N637);
nand NAND2 (N2784, N2781, N453);
buf BUF1 (N2785, N2771);
and AND4 (N2786, N2780, N2585, N2032, N2500);
buf BUF1 (N2787, N2785);
xor XOR2 (N2788, N2770, N1725);
not NOT1 (N2789, N2787);
buf BUF1 (N2790, N2778);
and AND3 (N2791, N2789, N2505, N1099);
xor XOR2 (N2792, N2779, N1943);
nand NAND4 (N2793, N2792, N196, N2087, N593);
not NOT1 (N2794, N2784);
not NOT1 (N2795, N2794);
and AND2 (N2796, N2791, N1287);
xor XOR2 (N2797, N2790, N1931);
not NOT1 (N2798, N2783);
nand NAND4 (N2799, N2775, N1238, N1952, N241);
buf BUF1 (N2800, N2788);
nor NOR3 (N2801, N2796, N451, N1397);
and AND2 (N2802, N2786, N360);
nand NAND2 (N2803, N2793, N1062);
xor XOR2 (N2804, N2799, N784);
buf BUF1 (N2805, N2803);
buf BUF1 (N2806, N2797);
nand NAND2 (N2807, N2773, N462);
or OR2 (N2808, N2805, N1486);
and AND4 (N2809, N2774, N691, N1595, N2786);
nor NOR2 (N2810, N2804, N849);
nor NOR2 (N2811, N2801, N2567);
not NOT1 (N2812, N2807);
nand NAND3 (N2813, N2802, N1194, N806);
or OR3 (N2814, N2806, N2556, N539);
not NOT1 (N2815, N2811);
nand NAND2 (N2816, N2808, N697);
nor NOR2 (N2817, N2798, N554);
xor XOR2 (N2818, N2795, N1167);
not NOT1 (N2819, N2818);
nand NAND3 (N2820, N2816, N2335, N595);
buf BUF1 (N2821, N2820);
nor NOR2 (N2822, N2809, N179);
nor NOR3 (N2823, N2813, N980, N324);
nand NAND4 (N2824, N2819, N1775, N230, N2214);
buf BUF1 (N2825, N2822);
xor XOR2 (N2826, N2812, N51);
or OR4 (N2827, N2810, N1022, N1897, N253);
or OR4 (N2828, N2824, N355, N902, N1797);
nand NAND4 (N2829, N2815, N2257, N2347, N2204);
and AND2 (N2830, N2828, N1691);
xor XOR2 (N2831, N2817, N388);
not NOT1 (N2832, N2826);
nand NAND4 (N2833, N2832, N1292, N1656, N2370);
buf BUF1 (N2834, N2831);
buf BUF1 (N2835, N2825);
xor XOR2 (N2836, N2821, N1199);
nor NOR3 (N2837, N2800, N605, N727);
not NOT1 (N2838, N2829);
nor NOR2 (N2839, N2836, N2371);
buf BUF1 (N2840, N2835);
not NOT1 (N2841, N2837);
xor XOR2 (N2842, N2841, N106);
not NOT1 (N2843, N2842);
xor XOR2 (N2844, N2827, N1310);
buf BUF1 (N2845, N2838);
nor NOR3 (N2846, N2833, N1382, N908);
and AND3 (N2847, N2823, N2641, N293);
and AND4 (N2848, N2830, N2645, N1126, N1104);
nor NOR2 (N2849, N2845, N2699);
or OR4 (N2850, N2849, N2420, N2263, N1575);
nor NOR3 (N2851, N2846, N1463, N1587);
xor XOR2 (N2852, N2834, N1262);
or OR3 (N2853, N2850, N179, N1153);
buf BUF1 (N2854, N2814);
nor NOR4 (N2855, N2839, N1259, N1264, N1770);
nor NOR3 (N2856, N2843, N1376, N2442);
not NOT1 (N2857, N2855);
nor NOR3 (N2858, N2844, N601, N903);
xor XOR2 (N2859, N2853, N2086);
or OR4 (N2860, N2856, N1188, N2759, N246);
and AND3 (N2861, N2860, N1013, N366);
or OR4 (N2862, N2858, N2612, N564, N2206);
not NOT1 (N2863, N2848);
nand NAND2 (N2864, N2857, N2295);
not NOT1 (N2865, N2847);
buf BUF1 (N2866, N2859);
and AND2 (N2867, N2864, N1784);
xor XOR2 (N2868, N2865, N1277);
not NOT1 (N2869, N2866);
and AND4 (N2870, N2840, N2736, N744, N1812);
buf BUF1 (N2871, N2868);
xor XOR2 (N2872, N2854, N1296);
nor NOR4 (N2873, N2870, N2199, N314, N310);
nor NOR2 (N2874, N2873, N1001);
or OR2 (N2875, N2869, N31);
or OR4 (N2876, N2872, N1533, N2367, N2486);
buf BUF1 (N2877, N2863);
and AND3 (N2878, N2876, N2818, N2207);
not NOT1 (N2879, N2875);
not NOT1 (N2880, N2879);
or OR2 (N2881, N2877, N2561);
nand NAND3 (N2882, N2867, N790, N821);
not NOT1 (N2883, N2871);
or OR3 (N2884, N2861, N992, N1002);
buf BUF1 (N2885, N2851);
nor NOR4 (N2886, N2874, N767, N2128, N2027);
nand NAND4 (N2887, N2885, N934, N853, N1456);
or OR3 (N2888, N2862, N1922, N755);
nor NOR4 (N2889, N2882, N345, N1673, N1680);
nand NAND4 (N2890, N2886, N2275, N1888, N1366);
or OR2 (N2891, N2887, N2274);
buf BUF1 (N2892, N2881);
nand NAND4 (N2893, N2892, N1681, N1834, N273);
nor NOR2 (N2894, N2893, N947);
not NOT1 (N2895, N2884);
nor NOR4 (N2896, N2891, N2701, N900, N1282);
or OR4 (N2897, N2852, N941, N2516, N1117);
xor XOR2 (N2898, N2888, N2335);
xor XOR2 (N2899, N2878, N2888);
nor NOR2 (N2900, N2890, N2739);
and AND4 (N2901, N2900, N2856, N438, N1261);
or OR4 (N2902, N2880, N1920, N1154, N1672);
and AND3 (N2903, N2894, N536, N1831);
nor NOR2 (N2904, N2898, N414);
and AND2 (N2905, N2895, N1958);
not NOT1 (N2906, N2897);
xor XOR2 (N2907, N2896, N1703);
xor XOR2 (N2908, N2883, N8);
and AND2 (N2909, N2905, N1600);
xor XOR2 (N2910, N2901, N1417);
nand NAND4 (N2911, N2910, N955, N1810, N1601);
nor NOR4 (N2912, N2906, N1101, N1341, N1756);
nand NAND4 (N2913, N2899, N1591, N479, N2662);
not NOT1 (N2914, N2904);
and AND4 (N2915, N2889, N262, N2726, N1708);
xor XOR2 (N2916, N2912, N2778);
or OR2 (N2917, N2916, N2008);
buf BUF1 (N2918, N2908);
nor NOR2 (N2919, N2914, N272);
xor XOR2 (N2920, N2907, N1585);
or OR3 (N2921, N2911, N1214, N244);
nor NOR4 (N2922, N2915, N1150, N2803, N1436);
buf BUF1 (N2923, N2917);
buf BUF1 (N2924, N2903);
and AND3 (N2925, N2902, N1617, N1311);
buf BUF1 (N2926, N2919);
nand NAND2 (N2927, N2924, N1122);
buf BUF1 (N2928, N2925);
xor XOR2 (N2929, N2926, N2219);
and AND4 (N2930, N2921, N2164, N730, N2196);
buf BUF1 (N2931, N2928);
or OR4 (N2932, N2930, N1796, N2616, N514);
nand NAND2 (N2933, N2923, N1409);
not NOT1 (N2934, N2929);
buf BUF1 (N2935, N2933);
nor NOR3 (N2936, N2918, N2790, N2605);
or OR2 (N2937, N2931, N2465);
not NOT1 (N2938, N2934);
and AND2 (N2939, N2932, N2248);
not NOT1 (N2940, N2922);
and AND3 (N2941, N2927, N45, N1403);
buf BUF1 (N2942, N2936);
and AND4 (N2943, N2935, N2482, N1091, N495);
not NOT1 (N2944, N2942);
and AND3 (N2945, N2943, N1251, N1750);
buf BUF1 (N2946, N2939);
xor XOR2 (N2947, N2945, N2117);
buf BUF1 (N2948, N2940);
not NOT1 (N2949, N2938);
buf BUF1 (N2950, N2909);
and AND2 (N2951, N2950, N818);
not NOT1 (N2952, N2937);
or OR3 (N2953, N2944, N477, N1235);
xor XOR2 (N2954, N2948, N1663);
xor XOR2 (N2955, N2947, N2246);
nor NOR4 (N2956, N2953, N1050, N2491, N1022);
not NOT1 (N2957, N2954);
nand NAND3 (N2958, N2913, N520, N2777);
nor NOR4 (N2959, N2952, N1097, N925, N2727);
nor NOR4 (N2960, N2949, N232, N1094, N1975);
and AND3 (N2961, N2951, N1063, N2461);
xor XOR2 (N2962, N2957, N1926);
nor NOR3 (N2963, N2946, N1867, N2759);
nor NOR3 (N2964, N2956, N58, N47);
or OR4 (N2965, N2941, N1547, N980, N2929);
buf BUF1 (N2966, N2960);
nand NAND2 (N2967, N2961, N1153);
buf BUF1 (N2968, N2963);
nand NAND2 (N2969, N2959, N1275);
or OR4 (N2970, N2969, N1915, N1699, N1549);
not NOT1 (N2971, N2968);
nand NAND4 (N2972, N2958, N1089, N2111, N1662);
nand NAND3 (N2973, N2967, N2342, N1835);
or OR4 (N2974, N2972, N2551, N1212, N1254);
not NOT1 (N2975, N2955);
not NOT1 (N2976, N2970);
and AND4 (N2977, N2920, N2847, N211, N1036);
nor NOR4 (N2978, N2966, N1958, N1764, N2613);
or OR3 (N2979, N2965, N2693, N476);
and AND4 (N2980, N2975, N694, N1767, N2559);
nand NAND4 (N2981, N2979, N2290, N2159, N13);
xor XOR2 (N2982, N2974, N522);
not NOT1 (N2983, N2973);
nor NOR4 (N2984, N2962, N2701, N2208, N2668);
xor XOR2 (N2985, N2981, N1771);
not NOT1 (N2986, N2985);
not NOT1 (N2987, N2980);
or OR2 (N2988, N2978, N2546);
not NOT1 (N2989, N2984);
or OR2 (N2990, N2986, N2464);
buf BUF1 (N2991, N2989);
or OR4 (N2992, N2990, N1976, N1905, N1251);
buf BUF1 (N2993, N2976);
buf BUF1 (N2994, N2987);
buf BUF1 (N2995, N2983);
nand NAND4 (N2996, N2992, N1452, N147, N2708);
and AND4 (N2997, N2994, N2490, N1251, N2551);
xor XOR2 (N2998, N2977, N1111);
xor XOR2 (N2999, N2982, N1174);
buf BUF1 (N3000, N2997);
or OR4 (N3001, N2964, N130, N993, N2747);
nor NOR2 (N3002, N2995, N542);
nand NAND2 (N3003, N2971, N582);
xor XOR2 (N3004, N2999, N2066);
not NOT1 (N3005, N3000);
buf BUF1 (N3006, N3001);
nor NOR3 (N3007, N3002, N2000, N1954);
not NOT1 (N3008, N2998);
or OR4 (N3009, N3003, N2129, N662, N2803);
not NOT1 (N3010, N3006);
xor XOR2 (N3011, N3009, N2515);
not NOT1 (N3012, N2996);
and AND3 (N3013, N3012, N549, N2548);
not NOT1 (N3014, N2991);
nor NOR4 (N3015, N3010, N919, N1122, N1400);
buf BUF1 (N3016, N3014);
not NOT1 (N3017, N3015);
nor NOR2 (N3018, N2988, N277);
nor NOR2 (N3019, N3005, N1351);
nor NOR3 (N3020, N3019, N2213, N2206);
not NOT1 (N3021, N3007);
or OR3 (N3022, N3021, N1093, N197);
xor XOR2 (N3023, N3018, N2087);
or OR2 (N3024, N3020, N1625);
and AND3 (N3025, N2993, N2127, N374);
nand NAND3 (N3026, N3023, N1828, N893);
nor NOR3 (N3027, N3008, N2856, N170);
buf BUF1 (N3028, N3026);
xor XOR2 (N3029, N3004, N804);
nor NOR2 (N3030, N3025, N471);
or OR2 (N3031, N3016, N1613);
buf BUF1 (N3032, N3011);
and AND4 (N3033, N3022, N1144, N2763, N822);
xor XOR2 (N3034, N3031, N1259);
or OR3 (N3035, N3013, N2089, N1404);
xor XOR2 (N3036, N3027, N1005);
xor XOR2 (N3037, N3028, N2750);
buf BUF1 (N3038, N3024);
and AND2 (N3039, N3034, N105);
or OR3 (N3040, N3017, N2204, N2190);
nor NOR3 (N3041, N3036, N577, N906);
not NOT1 (N3042, N3038);
buf BUF1 (N3043, N3040);
xor XOR2 (N3044, N3032, N983);
not NOT1 (N3045, N3039);
nor NOR3 (N3046, N3029, N1020, N2972);
not NOT1 (N3047, N3044);
or OR3 (N3048, N3041, N158, N2207);
nand NAND2 (N3049, N3048, N513);
not NOT1 (N3050, N3030);
nand NAND4 (N3051, N3033, N2614, N925, N1437);
not NOT1 (N3052, N3046);
not NOT1 (N3053, N3037);
xor XOR2 (N3054, N3045, N2005);
not NOT1 (N3055, N3054);
or OR4 (N3056, N3052, N591, N2695, N1140);
nand NAND4 (N3057, N3035, N574, N987, N1103);
not NOT1 (N3058, N3051);
xor XOR2 (N3059, N3042, N760);
xor XOR2 (N3060, N3043, N856);
xor XOR2 (N3061, N3060, N591);
xor XOR2 (N3062, N3049, N2784);
nand NAND2 (N3063, N3047, N231);
buf BUF1 (N3064, N3062);
and AND2 (N3065, N3058, N3056);
or OR4 (N3066, N2909, N911, N2139, N1630);
and AND4 (N3067, N3050, N1197, N779, N2249);
not NOT1 (N3068, N3067);
not NOT1 (N3069, N3068);
nor NOR4 (N3070, N3065, N2983, N2282, N736);
and AND3 (N3071, N3061, N1671, N3027);
and AND2 (N3072, N3064, N2877);
nor NOR2 (N3073, N3055, N2478);
xor XOR2 (N3074, N3072, N785);
nand NAND3 (N3075, N3070, N1142, N2254);
xor XOR2 (N3076, N3063, N2067);
and AND3 (N3077, N3073, N2420, N2513);
not NOT1 (N3078, N3076);
xor XOR2 (N3079, N3074, N2512);
not NOT1 (N3080, N3066);
or OR3 (N3081, N3075, N2965, N2370);
xor XOR2 (N3082, N3059, N1970);
and AND3 (N3083, N3077, N2568, N880);
xor XOR2 (N3084, N3080, N1981);
and AND3 (N3085, N3069, N1446, N1812);
buf BUF1 (N3086, N3084);
buf BUF1 (N3087, N3057);
buf BUF1 (N3088, N3085);
xor XOR2 (N3089, N3071, N1493);
or OR4 (N3090, N3078, N3003, N2382, N602);
not NOT1 (N3091, N3087);
nor NOR2 (N3092, N3091, N1915);
or OR3 (N3093, N3081, N2667, N731);
nor NOR3 (N3094, N3088, N2953, N1254);
and AND2 (N3095, N3082, N2438);
and AND4 (N3096, N3095, N1639, N1952, N2117);
or OR4 (N3097, N3083, N461, N561, N1313);
or OR3 (N3098, N3053, N1003, N138);
nand NAND4 (N3099, N3090, N1915, N2289, N1556);
or OR3 (N3100, N3099, N2257, N120);
not NOT1 (N3101, N3094);
xor XOR2 (N3102, N3079, N1191);
nand NAND4 (N3103, N3102, N2804, N2681, N2154);
and AND3 (N3104, N3101, N701, N1054);
nand NAND3 (N3105, N3104, N3059, N1804);
nand NAND2 (N3106, N3105, N537);
nand NAND4 (N3107, N3098, N750, N220, N2094);
xor XOR2 (N3108, N3092, N1563);
or OR4 (N3109, N3093, N1029, N2079, N1751);
nor NOR4 (N3110, N3096, N246, N681, N2495);
nand NAND3 (N3111, N3109, N523, N734);
nand NAND3 (N3112, N3111, N353, N2030);
not NOT1 (N3113, N3089);
xor XOR2 (N3114, N3100, N561);
not NOT1 (N3115, N3097);
xor XOR2 (N3116, N3113, N36);
xor XOR2 (N3117, N3112, N3011);
xor XOR2 (N3118, N3107, N679);
not NOT1 (N3119, N3117);
nand NAND3 (N3120, N3106, N2136, N2759);
nand NAND2 (N3121, N3115, N178);
not NOT1 (N3122, N3108);
buf BUF1 (N3123, N3122);
nor NOR4 (N3124, N3119, N210, N675, N2513);
buf BUF1 (N3125, N3110);
or OR4 (N3126, N3114, N2862, N2689, N755);
and AND2 (N3127, N3124, N2261);
nor NOR2 (N3128, N3123, N941);
not NOT1 (N3129, N3125);
not NOT1 (N3130, N3126);
buf BUF1 (N3131, N3116);
not NOT1 (N3132, N3128);
nor NOR2 (N3133, N3120, N936);
nand NAND3 (N3134, N3132, N1314, N1347);
xor XOR2 (N3135, N3103, N2560);
xor XOR2 (N3136, N3121, N2204);
nand NAND4 (N3137, N3133, N1754, N1718, N489);
nor NOR3 (N3138, N3131, N253, N1667);
not NOT1 (N3139, N3136);
buf BUF1 (N3140, N3127);
nor NOR4 (N3141, N3140, N839, N1720, N2194);
nand NAND2 (N3142, N3138, N1960);
or OR4 (N3143, N3086, N2894, N1937, N131);
not NOT1 (N3144, N3137);
and AND2 (N3145, N3141, N1593);
nand NAND2 (N3146, N3143, N2698);
or OR3 (N3147, N3139, N614, N1010);
not NOT1 (N3148, N3118);
buf BUF1 (N3149, N3142);
or OR2 (N3150, N3130, N2046);
or OR2 (N3151, N3149, N2013);
buf BUF1 (N3152, N3135);
buf BUF1 (N3153, N3148);
nand NAND2 (N3154, N3147, N2916);
and AND4 (N3155, N3129, N1214, N1570, N3147);
buf BUF1 (N3156, N3145);
buf BUF1 (N3157, N3152);
and AND4 (N3158, N3154, N144, N2657, N1503);
or OR2 (N3159, N3146, N2350);
nand NAND3 (N3160, N3159, N1628, N1935);
nor NOR2 (N3161, N3144, N3054);
not NOT1 (N3162, N3151);
or OR2 (N3163, N3134, N871);
and AND3 (N3164, N3155, N477, N1817);
buf BUF1 (N3165, N3161);
xor XOR2 (N3166, N3164, N496);
or OR2 (N3167, N3157, N2043);
nor NOR3 (N3168, N3162, N2926, N2616);
not NOT1 (N3169, N3153);
xor XOR2 (N3170, N3163, N965);
or OR3 (N3171, N3165, N383, N2303);
or OR4 (N3172, N3167, N1433, N3027, N1948);
nor NOR4 (N3173, N3171, N1708, N2669, N706);
and AND4 (N3174, N3158, N1578, N164, N1375);
xor XOR2 (N3175, N3168, N329);
not NOT1 (N3176, N3160);
not NOT1 (N3177, N3172);
not NOT1 (N3178, N3170);
nand NAND3 (N3179, N3156, N2881, N715);
xor XOR2 (N3180, N3169, N2372);
nor NOR2 (N3181, N3174, N954);
xor XOR2 (N3182, N3178, N1456);
buf BUF1 (N3183, N3176);
and AND4 (N3184, N3166, N2940, N2168, N2122);
or OR3 (N3185, N3180, N3043, N205);
nor NOR4 (N3186, N3175, N1337, N1111, N1417);
or OR2 (N3187, N3179, N515);
not NOT1 (N3188, N3173);
or OR2 (N3189, N3183, N2150);
or OR3 (N3190, N3188, N3167, N339);
buf BUF1 (N3191, N3187);
nand NAND4 (N3192, N3177, N418, N2131, N491);
nor NOR3 (N3193, N3186, N518, N1936);
not NOT1 (N3194, N3185);
nor NOR3 (N3195, N3192, N214, N2718);
or OR4 (N3196, N3182, N2738, N349, N932);
xor XOR2 (N3197, N3189, N1025);
nand NAND3 (N3198, N3191, N1088, N1813);
buf BUF1 (N3199, N3196);
and AND3 (N3200, N3195, N2957, N1754);
buf BUF1 (N3201, N3190);
nand NAND2 (N3202, N3198, N30);
nor NOR2 (N3203, N3184, N767);
or OR2 (N3204, N3201, N1800);
buf BUF1 (N3205, N3181);
xor XOR2 (N3206, N3197, N219);
buf BUF1 (N3207, N3199);
not NOT1 (N3208, N3207);
nor NOR2 (N3209, N3150, N1722);
not NOT1 (N3210, N3202);
nor NOR4 (N3211, N3210, N1399, N2225, N702);
buf BUF1 (N3212, N3206);
and AND4 (N3213, N3193, N2736, N1409, N244);
nand NAND2 (N3214, N3213, N1997);
xor XOR2 (N3215, N3194, N1139);
nor NOR4 (N3216, N3203, N2888, N2972, N671);
nor NOR3 (N3217, N3214, N3180, N1711);
or OR3 (N3218, N3216, N716, N26);
nand NAND4 (N3219, N3205, N2069, N871, N505);
nand NAND3 (N3220, N3218, N2099, N391);
nand NAND4 (N3221, N3204, N1277, N2993, N1804);
or OR2 (N3222, N3208, N2774);
nand NAND3 (N3223, N3211, N1060, N2088);
and AND3 (N3224, N3223, N2236, N3189);
or OR2 (N3225, N3220, N2512);
or OR2 (N3226, N3212, N1710);
and AND3 (N3227, N3226, N2356, N252);
nor NOR2 (N3228, N3221, N1534);
and AND3 (N3229, N3219, N2578, N2372);
nor NOR2 (N3230, N3222, N784);
or OR3 (N3231, N3200, N996, N315);
nor NOR2 (N3232, N3230, N3227);
xor XOR2 (N3233, N695, N1146);
xor XOR2 (N3234, N3228, N2639);
nor NOR2 (N3235, N3217, N1959);
or OR3 (N3236, N3215, N326, N581);
or OR3 (N3237, N3233, N1908, N385);
not NOT1 (N3238, N3236);
buf BUF1 (N3239, N3225);
nand NAND2 (N3240, N3234, N211);
nor NOR4 (N3241, N3239, N3015, N320, N773);
nand NAND3 (N3242, N3241, N2878, N1224);
buf BUF1 (N3243, N3237);
nor NOR4 (N3244, N3243, N792, N1654, N999);
and AND3 (N3245, N3229, N1698, N3179);
xor XOR2 (N3246, N3232, N2425);
buf BUF1 (N3247, N3238);
xor XOR2 (N3248, N3242, N1952);
not NOT1 (N3249, N3235);
or OR3 (N3250, N3240, N1234, N822);
nand NAND2 (N3251, N3249, N1834);
nand NAND2 (N3252, N3251, N173);
and AND3 (N3253, N3246, N2707, N3171);
nand NAND2 (N3254, N3245, N1420);
buf BUF1 (N3255, N3254);
and AND2 (N3256, N3209, N1031);
and AND3 (N3257, N3224, N2673, N1695);
not NOT1 (N3258, N3253);
nor NOR2 (N3259, N3257, N2395);
nor NOR4 (N3260, N3252, N801, N787, N1436);
buf BUF1 (N3261, N3255);
buf BUF1 (N3262, N3260);
or OR4 (N3263, N3231, N2399, N1576, N786);
buf BUF1 (N3264, N3256);
xor XOR2 (N3265, N3244, N3058);
buf BUF1 (N3266, N3247);
and AND3 (N3267, N3262, N373, N1739);
not NOT1 (N3268, N3266);
xor XOR2 (N3269, N3248, N1771);
xor XOR2 (N3270, N3264, N1836);
and AND2 (N3271, N3258, N502);
nor NOR2 (N3272, N3267, N2682);
not NOT1 (N3273, N3268);
xor XOR2 (N3274, N3263, N1052);
xor XOR2 (N3275, N3270, N2751);
and AND3 (N3276, N3261, N519, N622);
nor NOR2 (N3277, N3273, N2786);
nand NAND3 (N3278, N3250, N492, N2194);
buf BUF1 (N3279, N3277);
buf BUF1 (N3280, N3278);
nand NAND4 (N3281, N3271, N3275, N1020, N897);
not NOT1 (N3282, N2826);
xor XOR2 (N3283, N3276, N822);
and AND2 (N3284, N3265, N1131);
nor NOR4 (N3285, N3259, N829, N455, N366);
or OR4 (N3286, N3285, N2371, N425, N20);
not NOT1 (N3287, N3269);
and AND3 (N3288, N3282, N1124, N3192);
and AND4 (N3289, N3280, N2541, N2747, N3044);
buf BUF1 (N3290, N3272);
buf BUF1 (N3291, N3279);
nand NAND2 (N3292, N3289, N2580);
nor NOR4 (N3293, N3287, N2348, N714, N1079);
nor NOR3 (N3294, N3286, N3185, N3108);
or OR2 (N3295, N3292, N2867);
nor NOR4 (N3296, N3274, N1727, N817, N191);
buf BUF1 (N3297, N3288);
buf BUF1 (N3298, N3283);
and AND4 (N3299, N3295, N755, N2454, N3243);
buf BUF1 (N3300, N3293);
or OR2 (N3301, N3294, N2970);
or OR2 (N3302, N3298, N877);
and AND4 (N3303, N3291, N3004, N2979, N1417);
nand NAND3 (N3304, N3281, N938, N296);
buf BUF1 (N3305, N3301);
and AND2 (N3306, N3300, N1229);
xor XOR2 (N3307, N3304, N3001);
buf BUF1 (N3308, N3306);
nor NOR3 (N3309, N3299, N1649, N606);
xor XOR2 (N3310, N3290, N1812);
not NOT1 (N3311, N3296);
xor XOR2 (N3312, N3305, N1645);
nand NAND3 (N3313, N3284, N916, N672);
xor XOR2 (N3314, N3302, N261);
or OR4 (N3315, N3314, N1328, N1891, N1915);
or OR2 (N3316, N3310, N2528);
not NOT1 (N3317, N3313);
or OR2 (N3318, N3315, N2053);
buf BUF1 (N3319, N3307);
and AND3 (N3320, N3317, N3163, N909);
buf BUF1 (N3321, N3311);
and AND3 (N3322, N3309, N1835, N3154);
xor XOR2 (N3323, N3312, N1232);
or OR3 (N3324, N3297, N237, N804);
or OR4 (N3325, N3322, N1275, N934, N1528);
nor NOR4 (N3326, N3325, N611, N739, N287);
not NOT1 (N3327, N3316);
not NOT1 (N3328, N3327);
buf BUF1 (N3329, N3321);
buf BUF1 (N3330, N3303);
or OR3 (N3331, N3308, N515, N578);
xor XOR2 (N3332, N3318, N541);
nor NOR2 (N3333, N3323, N2863);
xor XOR2 (N3334, N3330, N1273);
or OR3 (N3335, N3329, N2286, N2508);
buf BUF1 (N3336, N3319);
or OR3 (N3337, N3326, N3259, N1906);
and AND2 (N3338, N3324, N1091);
buf BUF1 (N3339, N3320);
xor XOR2 (N3340, N3334, N2842);
nand NAND2 (N3341, N3337, N797);
or OR4 (N3342, N3336, N2854, N3339, N1970);
nor NOR2 (N3343, N492, N1707);
nand NAND3 (N3344, N3343, N1874, N1417);
xor XOR2 (N3345, N3328, N2404);
and AND2 (N3346, N3342, N957);
nand NAND3 (N3347, N3341, N677, N2454);
xor XOR2 (N3348, N3346, N2698);
not NOT1 (N3349, N3344);
buf BUF1 (N3350, N3340);
or OR3 (N3351, N3350, N483, N1486);
or OR4 (N3352, N3345, N18, N2685, N2341);
xor XOR2 (N3353, N3332, N2357);
nand NAND3 (N3354, N3353, N3094, N2010);
nor NOR3 (N3355, N3354, N616, N2812);
xor XOR2 (N3356, N3347, N3240);
or OR3 (N3357, N3356, N1179, N2663);
nor NOR2 (N3358, N3351, N76);
not NOT1 (N3359, N3338);
not NOT1 (N3360, N3357);
and AND3 (N3361, N3352, N2219, N1162);
xor XOR2 (N3362, N3349, N3208);
or OR3 (N3363, N3333, N1015, N2346);
and AND2 (N3364, N3359, N856);
and AND2 (N3365, N3348, N1607);
nand NAND2 (N3366, N3360, N2753);
xor XOR2 (N3367, N3363, N207);
xor XOR2 (N3368, N3362, N2556);
nor NOR4 (N3369, N3361, N2072, N3190, N2677);
nor NOR3 (N3370, N3355, N2970, N72);
nor NOR2 (N3371, N3367, N504);
nor NOR3 (N3372, N3366, N175, N510);
or OR3 (N3373, N3371, N1928, N3036);
not NOT1 (N3374, N3368);
xor XOR2 (N3375, N3364, N1031);
and AND4 (N3376, N3370, N2130, N2729, N3026);
nor NOR4 (N3377, N3335, N2441, N1592, N3060);
nand NAND2 (N3378, N3365, N1087);
or OR4 (N3379, N3372, N3217, N397, N2870);
or OR3 (N3380, N3331, N1034, N2153);
and AND4 (N3381, N3378, N2800, N134, N2248);
xor XOR2 (N3382, N3373, N2554);
not NOT1 (N3383, N3375);
nand NAND4 (N3384, N3377, N2542, N202, N3300);
xor XOR2 (N3385, N3381, N892);
xor XOR2 (N3386, N3380, N2446);
xor XOR2 (N3387, N3379, N3173);
buf BUF1 (N3388, N3383);
nor NOR3 (N3389, N3374, N2694, N2252);
nor NOR2 (N3390, N3388, N1943);
nand NAND4 (N3391, N3390, N2342, N883, N2443);
nand NAND4 (N3392, N3385, N2282, N1092, N558);
nor NOR3 (N3393, N3376, N391, N2833);
or OR3 (N3394, N3389, N510, N1226);
nor NOR3 (N3395, N3392, N1924, N3087);
nand NAND2 (N3396, N3384, N1045);
nor NOR2 (N3397, N3358, N763);
not NOT1 (N3398, N3382);
nor NOR3 (N3399, N3391, N917, N310);
or OR2 (N3400, N3393, N2645);
nor NOR4 (N3401, N3386, N2008, N1291, N1183);
and AND2 (N3402, N3401, N3190);
nor NOR3 (N3403, N3398, N1058, N994);
nor NOR4 (N3404, N3387, N2783, N3365, N206);
or OR4 (N3405, N3403, N3302, N2326, N949);
xor XOR2 (N3406, N3399, N1678);
xor XOR2 (N3407, N3400, N886);
or OR4 (N3408, N3395, N3334, N550, N16);
nand NAND4 (N3409, N3397, N482, N2727, N2081);
or OR3 (N3410, N3404, N618, N1455);
and AND4 (N3411, N3402, N271, N975, N757);
buf BUF1 (N3412, N3411);
not NOT1 (N3413, N3394);
or OR3 (N3414, N3408, N867, N538);
and AND2 (N3415, N3414, N781);
nor NOR4 (N3416, N3407, N1862, N2973, N1645);
buf BUF1 (N3417, N3405);
nand NAND4 (N3418, N3412, N1217, N2556, N2470);
xor XOR2 (N3419, N3396, N3412);
xor XOR2 (N3420, N3417, N1561);
or OR4 (N3421, N3418, N2819, N1263, N3279);
xor XOR2 (N3422, N3406, N2734);
nand NAND2 (N3423, N3416, N1075);
xor XOR2 (N3424, N3420, N1287);
buf BUF1 (N3425, N3424);
nand NAND3 (N3426, N3421, N2586, N1447);
or OR2 (N3427, N3422, N2718);
or OR3 (N3428, N3369, N1786, N2573);
or OR2 (N3429, N3410, N1526);
buf BUF1 (N3430, N3426);
or OR2 (N3431, N3413, N673);
or OR2 (N3432, N3425, N1639);
buf BUF1 (N3433, N3427);
nor NOR3 (N3434, N3429, N119, N158);
not NOT1 (N3435, N3419);
or OR3 (N3436, N3409, N2124, N713);
not NOT1 (N3437, N3432);
xor XOR2 (N3438, N3423, N1955);
and AND4 (N3439, N3415, N3346, N2087, N2232);
or OR3 (N3440, N3430, N179, N1155);
or OR4 (N3441, N3438, N1054, N3268, N3138);
nor NOR4 (N3442, N3436, N1688, N2297, N663);
nor NOR2 (N3443, N3435, N1805);
xor XOR2 (N3444, N3441, N810);
buf BUF1 (N3445, N3442);
not NOT1 (N3446, N3437);
nand NAND3 (N3447, N3443, N2689, N609);
not NOT1 (N3448, N3447);
nor NOR4 (N3449, N3431, N2834, N124, N3109);
nand NAND3 (N3450, N3439, N3288, N1038);
nand NAND2 (N3451, N3446, N3417);
buf BUF1 (N3452, N3428);
nor NOR2 (N3453, N3448, N2684);
buf BUF1 (N3454, N3444);
xor XOR2 (N3455, N3452, N1695);
xor XOR2 (N3456, N3440, N1964);
nor NOR2 (N3457, N3450, N537);
nand NAND3 (N3458, N3453, N288, N196);
buf BUF1 (N3459, N3445);
nand NAND4 (N3460, N3455, N2020, N2584, N521);
nor NOR3 (N3461, N3451, N1714, N2084);
nand NAND4 (N3462, N3454, N1386, N1339, N312);
buf BUF1 (N3463, N3456);
and AND4 (N3464, N3460, N2872, N899, N906);
nand NAND3 (N3465, N3459, N2950, N2074);
nor NOR3 (N3466, N3449, N1316, N279);
or OR3 (N3467, N3462, N1395, N2405);
or OR4 (N3468, N3464, N1773, N630, N2238);
and AND4 (N3469, N3465, N1494, N3295, N1366);
xor XOR2 (N3470, N3457, N514);
or OR2 (N3471, N3434, N1991);
xor XOR2 (N3472, N3466, N2704);
and AND3 (N3473, N3463, N3194, N3258);
buf BUF1 (N3474, N3469);
or OR2 (N3475, N3473, N144);
nor NOR4 (N3476, N3467, N94, N60, N1653);
and AND2 (N3477, N3475, N1116);
or OR4 (N3478, N3468, N2078, N2144, N3361);
and AND3 (N3479, N3433, N3141, N2179);
buf BUF1 (N3480, N3458);
and AND2 (N3481, N3471, N2597);
nor NOR4 (N3482, N3472, N2384, N1307, N2612);
and AND3 (N3483, N3480, N3258, N1765);
nand NAND4 (N3484, N3478, N3299, N3014, N524);
nor NOR4 (N3485, N3479, N1321, N2940, N1603);
and AND2 (N3486, N3470, N2211);
buf BUF1 (N3487, N3483);
buf BUF1 (N3488, N3482);
or OR2 (N3489, N3477, N2493);
or OR4 (N3490, N3485, N1071, N2318, N936);
and AND4 (N3491, N3461, N2358, N1485, N1858);
and AND2 (N3492, N3491, N409);
nand NAND4 (N3493, N3474, N2959, N618, N2926);
not NOT1 (N3494, N3489);
or OR4 (N3495, N3494, N3041, N2852, N1678);
not NOT1 (N3496, N3493);
and AND3 (N3497, N3481, N712, N113);
and AND3 (N3498, N3488, N2088, N1423);
and AND2 (N3499, N3476, N985);
nand NAND3 (N3500, N3497, N3413, N918);
buf BUF1 (N3501, N3495);
xor XOR2 (N3502, N3490, N3162);
and AND3 (N3503, N3492, N509, N1420);
nor NOR3 (N3504, N3503, N1900, N2717);
and AND4 (N3505, N3499, N1045, N275, N2308);
or OR4 (N3506, N3504, N1273, N2141, N450);
and AND4 (N3507, N3498, N2987, N308, N2656);
xor XOR2 (N3508, N3486, N1134);
buf BUF1 (N3509, N3508);
not NOT1 (N3510, N3484);
nor NOR2 (N3511, N3496, N1527);
not NOT1 (N3512, N3511);
and AND2 (N3513, N3509, N2668);
xor XOR2 (N3514, N3512, N238);
or OR3 (N3515, N3510, N2193, N2366);
not NOT1 (N3516, N3514);
and AND3 (N3517, N3500, N2628, N1916);
nand NAND4 (N3518, N3517, N1510, N1421, N735);
and AND2 (N3519, N3501, N406);
nand NAND2 (N3520, N3502, N3341);
xor XOR2 (N3521, N3516, N3462);
or OR3 (N3522, N3519, N854, N3017);
not NOT1 (N3523, N3513);
or OR4 (N3524, N3506, N1475, N861, N2444);
and AND4 (N3525, N3518, N2489, N947, N1241);
xor XOR2 (N3526, N3505, N3479);
and AND2 (N3527, N3524, N2095);
xor XOR2 (N3528, N3515, N863);
xor XOR2 (N3529, N3523, N2254);
and AND2 (N3530, N3527, N2434);
buf BUF1 (N3531, N3529);
buf BUF1 (N3532, N3530);
buf BUF1 (N3533, N3528);
or OR2 (N3534, N3522, N511);
buf BUF1 (N3535, N3532);
and AND3 (N3536, N3525, N2999, N3234);
nor NOR4 (N3537, N3536, N639, N3383, N3216);
nand NAND4 (N3538, N3520, N176, N1030, N3533);
or OR2 (N3539, N1575, N2808);
nor NOR3 (N3540, N3531, N3153, N1910);
nand NAND2 (N3541, N3535, N2155);
and AND3 (N3542, N3507, N729, N3023);
not NOT1 (N3543, N3542);
or OR2 (N3544, N3487, N1580);
nand NAND3 (N3545, N3540, N2081, N2653);
and AND3 (N3546, N3543, N3029, N592);
nor NOR2 (N3547, N3544, N1799);
buf BUF1 (N3548, N3521);
not NOT1 (N3549, N3547);
and AND4 (N3550, N3537, N3094, N1687, N2241);
nand NAND4 (N3551, N3526, N96, N88, N1743);
xor XOR2 (N3552, N3534, N330);
nand NAND2 (N3553, N3538, N3278);
buf BUF1 (N3554, N3553);
xor XOR2 (N3555, N3545, N1320);
buf BUF1 (N3556, N3554);
nand NAND2 (N3557, N3551, N433);
or OR2 (N3558, N3555, N243);
or OR3 (N3559, N3552, N1991, N3096);
or OR4 (N3560, N3559, N3538, N879, N985);
and AND3 (N3561, N3549, N1410, N2043);
and AND3 (N3562, N3541, N3095, N1335);
or OR3 (N3563, N3539, N2304, N3418);
buf BUF1 (N3564, N3561);
nand NAND2 (N3565, N3546, N3452);
or OR3 (N3566, N3564, N170, N2543);
nand NAND3 (N3567, N3550, N2111, N738);
not NOT1 (N3568, N3558);
nand NAND4 (N3569, N3562, N377, N2385, N1129);
xor XOR2 (N3570, N3556, N2782);
nand NAND4 (N3571, N3565, N1092, N2392, N1466);
not NOT1 (N3572, N3571);
nand NAND3 (N3573, N3557, N2435, N3221);
not NOT1 (N3574, N3567);
nor NOR3 (N3575, N3566, N2153, N2309);
not NOT1 (N3576, N3563);
or OR4 (N3577, N3574, N1910, N1716, N2542);
xor XOR2 (N3578, N3573, N354);
buf BUF1 (N3579, N3548);
buf BUF1 (N3580, N3576);
nand NAND2 (N3581, N3579, N2823);
xor XOR2 (N3582, N3568, N2648);
not NOT1 (N3583, N3578);
nand NAND3 (N3584, N3575, N2970, N1089);
nor NOR3 (N3585, N3580, N2990, N1668);
not NOT1 (N3586, N3584);
nor NOR3 (N3587, N3581, N1761, N1632);
nand NAND4 (N3588, N3570, N1948, N2442, N2433);
xor XOR2 (N3589, N3585, N1725);
nand NAND2 (N3590, N3583, N2611);
xor XOR2 (N3591, N3586, N3187);
not NOT1 (N3592, N3560);
or OR4 (N3593, N3592, N571, N2023, N3144);
nand NAND4 (N3594, N3590, N3032, N341, N2049);
nand NAND4 (N3595, N3588, N388, N3407, N1982);
nor NOR3 (N3596, N3589, N1821, N624);
nor NOR2 (N3597, N3595, N2496);
xor XOR2 (N3598, N3594, N1644);
buf BUF1 (N3599, N3569);
xor XOR2 (N3600, N3572, N261);
buf BUF1 (N3601, N3597);
buf BUF1 (N3602, N3582);
nand NAND3 (N3603, N3602, N958, N1102);
and AND3 (N3604, N3591, N1402, N921);
or OR3 (N3605, N3600, N3136, N2090);
and AND4 (N3606, N3577, N1988, N395, N3119);
buf BUF1 (N3607, N3599);
nor NOR2 (N3608, N3603, N622);
or OR3 (N3609, N3607, N3097, N2554);
not NOT1 (N3610, N3601);
or OR2 (N3611, N3609, N3223);
not NOT1 (N3612, N3596);
buf BUF1 (N3613, N3610);
nor NOR4 (N3614, N3612, N1949, N31, N3452);
and AND3 (N3615, N3587, N2278, N1183);
nor NOR4 (N3616, N3611, N2469, N639, N1112);
and AND2 (N3617, N3593, N1304);
xor XOR2 (N3618, N3617, N1291);
nor NOR4 (N3619, N3618, N1696, N1858, N654);
not NOT1 (N3620, N3614);
xor XOR2 (N3621, N3616, N2568);
buf BUF1 (N3622, N3605);
or OR3 (N3623, N3621, N482, N1739);
and AND2 (N3624, N3604, N149);
nand NAND4 (N3625, N3613, N1058, N381, N18);
not NOT1 (N3626, N3624);
nor NOR2 (N3627, N3615, N1139);
xor XOR2 (N3628, N3619, N1049);
and AND3 (N3629, N3622, N1991, N454);
nor NOR4 (N3630, N3606, N739, N1694, N1456);
not NOT1 (N3631, N3620);
xor XOR2 (N3632, N3631, N2097);
nand NAND4 (N3633, N3632, N2000, N258, N336);
nor NOR3 (N3634, N3633, N1647, N163);
xor XOR2 (N3635, N3626, N342);
nand NAND2 (N3636, N3608, N148);
and AND3 (N3637, N3628, N1584, N1928);
or OR2 (N3638, N3627, N1858);
and AND4 (N3639, N3636, N3160, N2553, N2675);
buf BUF1 (N3640, N3635);
buf BUF1 (N3641, N3637);
not NOT1 (N3642, N3623);
or OR4 (N3643, N3639, N267, N161, N2651);
not NOT1 (N3644, N3630);
not NOT1 (N3645, N3642);
nand NAND3 (N3646, N3598, N1868, N3563);
nand NAND2 (N3647, N3638, N1937);
and AND2 (N3648, N3641, N2411);
not NOT1 (N3649, N3640);
nand NAND3 (N3650, N3646, N2486, N366);
nand NAND3 (N3651, N3629, N2826, N3634);
not NOT1 (N3652, N956);
nand NAND2 (N3653, N3643, N2337);
and AND4 (N3654, N3649, N865, N572, N2894);
not NOT1 (N3655, N3645);
nand NAND4 (N3656, N3647, N1185, N337, N1129);
nand NAND2 (N3657, N3625, N1970);
or OR2 (N3658, N3655, N3330);
xor XOR2 (N3659, N3653, N2272);
nand NAND4 (N3660, N3658, N3358, N2171, N905);
xor XOR2 (N3661, N3651, N3649);
buf BUF1 (N3662, N3656);
or OR4 (N3663, N3648, N1790, N368, N485);
xor XOR2 (N3664, N3663, N3586);
nor NOR3 (N3665, N3660, N3657, N601);
nand NAND4 (N3666, N2381, N384, N2171, N2561);
nand NAND4 (N3667, N3662, N1243, N1443, N970);
and AND4 (N3668, N3650, N3173, N2978, N3474);
and AND2 (N3669, N3652, N3477);
nor NOR3 (N3670, N3661, N634, N2408);
xor XOR2 (N3671, N3659, N2403);
and AND2 (N3672, N3666, N3459);
and AND2 (N3673, N3669, N1253);
or OR4 (N3674, N3673, N3523, N2101, N3213);
or OR3 (N3675, N3672, N2051, N1168);
and AND2 (N3676, N3644, N2324);
buf BUF1 (N3677, N3676);
buf BUF1 (N3678, N3671);
xor XOR2 (N3679, N3654, N2466);
not NOT1 (N3680, N3674);
nor NOR2 (N3681, N3667, N215);
xor XOR2 (N3682, N3679, N2141);
nor NOR2 (N3683, N3677, N1685);
not NOT1 (N3684, N3665);
and AND4 (N3685, N3683, N608, N2129, N684);
or OR3 (N3686, N3685, N868, N1921);
xor XOR2 (N3687, N3670, N1135);
nand NAND2 (N3688, N3664, N288);
nand NAND2 (N3689, N3686, N2970);
xor XOR2 (N3690, N3684, N12);
not NOT1 (N3691, N3678);
nand NAND4 (N3692, N3690, N792, N2322, N153);
buf BUF1 (N3693, N3681);
and AND2 (N3694, N3687, N3293);
not NOT1 (N3695, N3691);
not NOT1 (N3696, N3680);
buf BUF1 (N3697, N3693);
or OR3 (N3698, N3695, N3508, N3190);
not NOT1 (N3699, N3675);
nand NAND4 (N3700, N3692, N3694, N3441, N1966);
buf BUF1 (N3701, N2787);
nor NOR3 (N3702, N3696, N237, N133);
nand NAND4 (N3703, N3698, N1828, N2374, N3041);
or OR4 (N3704, N3689, N2828, N735, N1603);
not NOT1 (N3705, N3697);
not NOT1 (N3706, N3704);
nor NOR3 (N3707, N3703, N270, N2592);
not NOT1 (N3708, N3706);
xor XOR2 (N3709, N3702, N3265);
and AND2 (N3710, N3705, N826);
xor XOR2 (N3711, N3707, N1318);
nor NOR3 (N3712, N3700, N2074, N43);
and AND2 (N3713, N3688, N160);
buf BUF1 (N3714, N3709);
nand NAND3 (N3715, N3714, N3396, N2070);
and AND4 (N3716, N3711, N2907, N3459, N1017);
not NOT1 (N3717, N3699);
nor NOR4 (N3718, N3708, N616, N1275, N2512);
nand NAND2 (N3719, N3712, N700);
buf BUF1 (N3720, N3719);
nor NOR3 (N3721, N3668, N1592, N1667);
not NOT1 (N3722, N3710);
nor NOR3 (N3723, N3715, N3524, N1035);
and AND3 (N3724, N3723, N851, N2686);
or OR2 (N3725, N3713, N102);
buf BUF1 (N3726, N3721);
xor XOR2 (N3727, N3726, N2842);
nor NOR3 (N3728, N3716, N2106, N1596);
or OR4 (N3729, N3727, N3617, N2092, N3598);
and AND4 (N3730, N3725, N989, N1347, N345);
nor NOR4 (N3731, N3729, N2614, N2361, N2921);
nand NAND3 (N3732, N3717, N957, N845);
buf BUF1 (N3733, N3701);
xor XOR2 (N3734, N3722, N688);
or OR3 (N3735, N3720, N1313, N1172);
buf BUF1 (N3736, N3735);
and AND3 (N3737, N3731, N383, N1981);
buf BUF1 (N3738, N3718);
xor XOR2 (N3739, N3728, N595);
or OR3 (N3740, N3736, N1471, N278);
buf BUF1 (N3741, N3682);
and AND3 (N3742, N3734, N1006, N3409);
nor NOR3 (N3743, N3740, N1581, N520);
nand NAND2 (N3744, N3738, N2287);
buf BUF1 (N3745, N3741);
xor XOR2 (N3746, N3730, N3062);
nand NAND2 (N3747, N3746, N480);
nor NOR4 (N3748, N3744, N1816, N3619, N1014);
nor NOR4 (N3749, N3745, N1007, N3427, N3201);
and AND2 (N3750, N3748, N1541);
and AND4 (N3751, N3750, N1177, N1241, N1189);
and AND2 (N3752, N3737, N1100);
not NOT1 (N3753, N3749);
not NOT1 (N3754, N3742);
buf BUF1 (N3755, N3753);
or OR4 (N3756, N3724, N881, N2506, N2394);
or OR2 (N3757, N3756, N1881);
buf BUF1 (N3758, N3732);
not NOT1 (N3759, N3757);
nor NOR4 (N3760, N3758, N215, N2972, N3480);
and AND3 (N3761, N3751, N2285, N2883);
and AND4 (N3762, N3760, N239, N2566, N1458);
not NOT1 (N3763, N3761);
nor NOR3 (N3764, N3762, N3371, N1200);
and AND3 (N3765, N3754, N2524, N1184);
or OR2 (N3766, N3759, N353);
not NOT1 (N3767, N3747);
xor XOR2 (N3768, N3739, N35);
nand NAND3 (N3769, N3767, N3432, N952);
buf BUF1 (N3770, N3764);
nand NAND3 (N3771, N3765, N1513, N3130);
not NOT1 (N3772, N3743);
nor NOR2 (N3773, N3771, N1493);
xor XOR2 (N3774, N3768, N376);
and AND3 (N3775, N3766, N1479, N1609);
nor NOR3 (N3776, N3733, N1046, N2173);
nand NAND2 (N3777, N3763, N1141);
and AND3 (N3778, N3774, N1997, N2186);
xor XOR2 (N3779, N3770, N1274);
not NOT1 (N3780, N3779);
not NOT1 (N3781, N3752);
not NOT1 (N3782, N3776);
buf BUF1 (N3783, N3775);
nor NOR3 (N3784, N3777, N81, N488);
nor NOR2 (N3785, N3784, N176);
nand NAND4 (N3786, N3785, N1597, N700, N1398);
not NOT1 (N3787, N3769);
xor XOR2 (N3788, N3772, N388);
or OR2 (N3789, N3778, N2905);
buf BUF1 (N3790, N3782);
and AND3 (N3791, N3781, N796, N1448);
or OR2 (N3792, N3790, N2864);
and AND4 (N3793, N3792, N3358, N3211, N2519);
nor NOR2 (N3794, N3793, N2981);
nand NAND4 (N3795, N3786, N2248, N1384, N1594);
nand NAND4 (N3796, N3780, N3674, N3009, N2552);
or OR2 (N3797, N3773, N3741);
nand NAND3 (N3798, N3789, N3667, N1176);
nand NAND3 (N3799, N3755, N3593, N447);
xor XOR2 (N3800, N3797, N2910);
not NOT1 (N3801, N3787);
nand NAND3 (N3802, N3796, N3051, N2125);
nor NOR4 (N3803, N3791, N2342, N649, N126);
and AND3 (N3804, N3788, N3625, N2810);
nand NAND4 (N3805, N3804, N3383, N2687, N360);
and AND4 (N3806, N3794, N177, N2243, N1868);
nor NOR3 (N3807, N3803, N1536, N876);
and AND3 (N3808, N3783, N322, N2804);
and AND3 (N3809, N3805, N979, N914);
or OR2 (N3810, N3800, N2014);
not NOT1 (N3811, N3799);
or OR4 (N3812, N3806, N1727, N1739, N1407);
and AND2 (N3813, N3809, N2980);
xor XOR2 (N3814, N3798, N2988);
and AND3 (N3815, N3795, N200, N568);
nor NOR4 (N3816, N3807, N501, N1106, N1072);
or OR2 (N3817, N3814, N3658);
or OR2 (N3818, N3808, N1354);
nor NOR2 (N3819, N3802, N3126);
and AND4 (N3820, N3812, N1638, N1341, N700);
and AND2 (N3821, N3818, N2921);
nand NAND4 (N3822, N3817, N3172, N1458, N2645);
not NOT1 (N3823, N3816);
and AND4 (N3824, N3811, N225, N765, N1326);
nand NAND2 (N3825, N3823, N3580);
or OR2 (N3826, N3820, N2772);
buf BUF1 (N3827, N3826);
nor NOR4 (N3828, N3810, N3777, N1513, N491);
or OR3 (N3829, N3828, N89, N1795);
nand NAND2 (N3830, N3819, N1435);
xor XOR2 (N3831, N3801, N2720);
nand NAND4 (N3832, N3821, N774, N1221, N1686);
not NOT1 (N3833, N3830);
nand NAND4 (N3834, N3813, N1539, N2387, N200);
buf BUF1 (N3835, N3827);
or OR2 (N3836, N3831, N1336);
nand NAND3 (N3837, N3824, N1413, N1020);
nand NAND3 (N3838, N3829, N556, N1525);
and AND2 (N3839, N3833, N507);
nand NAND2 (N3840, N3832, N3306);
buf BUF1 (N3841, N3836);
and AND2 (N3842, N3841, N64);
buf BUF1 (N3843, N3837);
xor XOR2 (N3844, N3835, N1127);
and AND4 (N3845, N3843, N500, N3252, N626);
xor XOR2 (N3846, N3822, N3759);
and AND3 (N3847, N3840, N2980, N2621);
nor NOR4 (N3848, N3845, N3153, N147, N938);
not NOT1 (N3849, N3842);
nor NOR4 (N3850, N3849, N3247, N1504, N2035);
buf BUF1 (N3851, N3839);
nor NOR2 (N3852, N3825, N1690);
not NOT1 (N3853, N3852);
nor NOR4 (N3854, N3844, N2335, N1664, N3779);
nor NOR3 (N3855, N3847, N1246, N99);
xor XOR2 (N3856, N3854, N91);
xor XOR2 (N3857, N3838, N1985);
xor XOR2 (N3858, N3848, N3566);
and AND4 (N3859, N3858, N240, N2639, N1248);
not NOT1 (N3860, N3846);
nand NAND2 (N3861, N3857, N2192);
nor NOR2 (N3862, N3861, N3585);
xor XOR2 (N3863, N3853, N3181);
or OR3 (N3864, N3860, N2317, N1148);
nor NOR3 (N3865, N3863, N277, N1153);
nand NAND4 (N3866, N3865, N1649, N2489, N2044);
xor XOR2 (N3867, N3834, N3815);
and AND4 (N3868, N1842, N1937, N3334, N1176);
or OR4 (N3869, N3856, N996, N369, N828);
nand NAND3 (N3870, N3855, N1778, N1762);
nor NOR2 (N3871, N3862, N947);
not NOT1 (N3872, N3871);
or OR3 (N3873, N3859, N365, N184);
nor NOR4 (N3874, N3868, N3817, N2125, N3437);
or OR3 (N3875, N3864, N1336, N84);
not NOT1 (N3876, N3874);
or OR3 (N3877, N3869, N2702, N2462);
buf BUF1 (N3878, N3866);
buf BUF1 (N3879, N3851);
or OR3 (N3880, N3876, N3106, N2198);
and AND3 (N3881, N3873, N2413, N869);
nor NOR3 (N3882, N3867, N702, N1769);
and AND3 (N3883, N3878, N1992, N982);
xor XOR2 (N3884, N3870, N1832);
nand NAND2 (N3885, N3879, N1125);
or OR4 (N3886, N3883, N2071, N461, N1230);
nand NAND4 (N3887, N3886, N1966, N2934, N1500);
nor NOR2 (N3888, N3875, N106);
nand NAND4 (N3889, N3872, N1542, N1062, N734);
xor XOR2 (N3890, N3880, N2004);
xor XOR2 (N3891, N3887, N1591);
buf BUF1 (N3892, N3888);
nor NOR2 (N3893, N3885, N770);
or OR2 (N3894, N3882, N3083);
buf BUF1 (N3895, N3884);
xor XOR2 (N3896, N3877, N708);
xor XOR2 (N3897, N3891, N2793);
or OR3 (N3898, N3881, N3681, N3530);
not NOT1 (N3899, N3898);
not NOT1 (N3900, N3897);
not NOT1 (N3901, N3890);
nor NOR4 (N3902, N3900, N570, N2766, N383);
or OR2 (N3903, N3893, N607);
buf BUF1 (N3904, N3899);
and AND2 (N3905, N3892, N2802);
nand NAND3 (N3906, N3905, N843, N868);
nand NAND2 (N3907, N3901, N2586);
and AND4 (N3908, N3903, N2843, N2901, N3441);
nor NOR4 (N3909, N3850, N540, N2488, N2269);
nand NAND4 (N3910, N3906, N1294, N2580, N2005);
buf BUF1 (N3911, N3904);
or OR4 (N3912, N3894, N1229, N2562, N3796);
xor XOR2 (N3913, N3912, N2603);
nand NAND3 (N3914, N3902, N991, N2253);
xor XOR2 (N3915, N3907, N243);
and AND3 (N3916, N3908, N2871, N1049);
xor XOR2 (N3917, N3916, N1153);
nand NAND2 (N3918, N3889, N1162);
not NOT1 (N3919, N3895);
buf BUF1 (N3920, N3910);
nor NOR2 (N3921, N3909, N3843);
nand NAND2 (N3922, N3915, N1009);
xor XOR2 (N3923, N3914, N1452);
buf BUF1 (N3924, N3919);
nor NOR2 (N3925, N3924, N3878);
nor NOR2 (N3926, N3917, N1481);
nand NAND2 (N3927, N3926, N3470);
nor NOR3 (N3928, N3927, N3192, N619);
nor NOR4 (N3929, N3913, N2864, N2297, N442);
buf BUF1 (N3930, N3923);
buf BUF1 (N3931, N3930);
not NOT1 (N3932, N3925);
nor NOR2 (N3933, N3896, N358);
nor NOR2 (N3934, N3911, N2642);
nor NOR4 (N3935, N3931, N2899, N2211, N938);
and AND3 (N3936, N3932, N2555, N3433);
nand NAND4 (N3937, N3929, N3386, N46, N767);
nand NAND3 (N3938, N3921, N3011, N2999);
not NOT1 (N3939, N3935);
buf BUF1 (N3940, N3920);
not NOT1 (N3941, N3928);
nor NOR3 (N3942, N3937, N3179, N754);
nor NOR4 (N3943, N3942, N3243, N3536, N3807);
and AND2 (N3944, N3936, N787);
not NOT1 (N3945, N3939);
and AND3 (N3946, N3918, N1696, N2840);
buf BUF1 (N3947, N3946);
or OR3 (N3948, N3933, N2377, N2741);
not NOT1 (N3949, N3943);
or OR2 (N3950, N3934, N3362);
or OR4 (N3951, N3940, N2182, N3121, N2454);
nor NOR4 (N3952, N3951, N906, N2459, N2312);
buf BUF1 (N3953, N3941);
buf BUF1 (N3954, N3922);
buf BUF1 (N3955, N3938);
nand NAND4 (N3956, N3944, N46, N3733, N2309);
buf BUF1 (N3957, N3953);
nand NAND4 (N3958, N3957, N2384, N1085, N2737);
or OR2 (N3959, N3947, N604);
and AND3 (N3960, N3945, N985, N3614);
buf BUF1 (N3961, N3960);
buf BUF1 (N3962, N3958);
not NOT1 (N3963, N3962);
not NOT1 (N3964, N3948);
nor NOR4 (N3965, N3949, N2012, N100, N2596);
and AND2 (N3966, N3950, N1650);
not NOT1 (N3967, N3954);
buf BUF1 (N3968, N3965);
nor NOR4 (N3969, N3966, N3747, N2027, N2782);
nand NAND3 (N3970, N3961, N2461, N3930);
nand NAND2 (N3971, N3959, N1575);
and AND3 (N3972, N3964, N3952, N360);
not NOT1 (N3973, N2697);
nand NAND4 (N3974, N3968, N3329, N2498, N2130);
nand NAND3 (N3975, N3956, N1808, N2853);
not NOT1 (N3976, N3974);
nand NAND2 (N3977, N3972, N230);
or OR2 (N3978, N3973, N2987);
not NOT1 (N3979, N3976);
nand NAND4 (N3980, N3967, N2694, N994, N522);
not NOT1 (N3981, N3971);
nand NAND2 (N3982, N3978, N2816);
not NOT1 (N3983, N3980);
xor XOR2 (N3984, N3977, N2874);
nand NAND4 (N3985, N3963, N3350, N223, N3437);
nor NOR3 (N3986, N3969, N2283, N1930);
nor NOR4 (N3987, N3975, N475, N3024, N1249);
and AND4 (N3988, N3982, N2161, N777, N2856);
nor NOR3 (N3989, N3984, N1265, N2174);
nor NOR2 (N3990, N3970, N2010);
xor XOR2 (N3991, N3988, N2148);
nand NAND4 (N3992, N3979, N2516, N637, N224);
and AND2 (N3993, N3992, N645);
buf BUF1 (N3994, N3985);
nand NAND4 (N3995, N3987, N3913, N2897, N2763);
nor NOR2 (N3996, N3991, N1431);
nor NOR4 (N3997, N3995, N1676, N669, N1873);
nand NAND2 (N3998, N3981, N1754);
buf BUF1 (N3999, N3990);
buf BUF1 (N4000, N3989);
buf BUF1 (N4001, N3993);
xor XOR2 (N4002, N3986, N777);
or OR3 (N4003, N4001, N3940, N867);
nand NAND2 (N4004, N3955, N3964);
buf BUF1 (N4005, N3983);
buf BUF1 (N4006, N3998);
or OR2 (N4007, N3996, N864);
and AND4 (N4008, N4004, N877, N675, N906);
xor XOR2 (N4009, N3999, N1743);
or OR3 (N4010, N4007, N2951, N3551);
buf BUF1 (N4011, N3997);
buf BUF1 (N4012, N4008);
nor NOR4 (N4013, N4011, N1052, N2136, N2449);
or OR4 (N4014, N4013, N25, N3261, N2365);
and AND3 (N4015, N4002, N3360, N154);
xor XOR2 (N4016, N3994, N1329);
xor XOR2 (N4017, N4010, N3826);
buf BUF1 (N4018, N4017);
not NOT1 (N4019, N4015);
nor NOR2 (N4020, N4005, N1778);
or OR2 (N4021, N4009, N1104);
buf BUF1 (N4022, N4018);
or OR2 (N4023, N4014, N310);
and AND4 (N4024, N4023, N133, N893, N362);
nand NAND4 (N4025, N4016, N1293, N2371, N957);
and AND4 (N4026, N4000, N249, N837, N550);
buf BUF1 (N4027, N4006);
and AND2 (N4028, N4020, N1178);
nor NOR3 (N4029, N4003, N856, N36);
nor NOR2 (N4030, N4012, N3005);
nand NAND2 (N4031, N4028, N993);
or OR3 (N4032, N4027, N3385, N1356);
buf BUF1 (N4033, N4022);
or OR3 (N4034, N4025, N3173, N1194);
xor XOR2 (N4035, N4019, N3208);
and AND2 (N4036, N4024, N180);
nand NAND3 (N4037, N4032, N3936, N646);
xor XOR2 (N4038, N4034, N1092);
and AND3 (N4039, N4037, N302, N3629);
nor NOR4 (N4040, N4026, N2899, N1567, N3304);
not NOT1 (N4041, N4033);
buf BUF1 (N4042, N4040);
and AND4 (N4043, N4031, N3165, N3001, N3103);
nand NAND3 (N4044, N4035, N1449, N3927);
and AND4 (N4045, N4021, N1767, N485, N2571);
and AND2 (N4046, N4043, N1656);
and AND4 (N4047, N4045, N1495, N3393, N1127);
buf BUF1 (N4048, N4029);
buf BUF1 (N4049, N4041);
buf BUF1 (N4050, N4046);
buf BUF1 (N4051, N4036);
nand NAND4 (N4052, N4039, N858, N2282, N717);
or OR2 (N4053, N4051, N2360);
xor XOR2 (N4054, N4042, N3511);
nand NAND4 (N4055, N4053, N1761, N2406, N1326);
or OR2 (N4056, N4047, N2772);
nand NAND2 (N4057, N4044, N1347);
nand NAND4 (N4058, N4038, N1711, N3122, N130);
or OR4 (N4059, N4030, N1255, N2301, N2714);
nand NAND2 (N4060, N4048, N470);
not NOT1 (N4061, N4049);
nor NOR4 (N4062, N4057, N2901, N2361, N3932);
not NOT1 (N4063, N4061);
nor NOR2 (N4064, N4058, N3454);
or OR4 (N4065, N4056, N2912, N2626, N454);
not NOT1 (N4066, N4062);
buf BUF1 (N4067, N4063);
and AND4 (N4068, N4065, N1761, N2716, N1546);
and AND4 (N4069, N4067, N1256, N2896, N2925);
not NOT1 (N4070, N4069);
buf BUF1 (N4071, N4050);
and AND4 (N4072, N4059, N3820, N3534, N2696);
or OR3 (N4073, N4068, N2112, N18);
and AND3 (N4074, N4072, N1716, N3244);
xor XOR2 (N4075, N4074, N2328);
xor XOR2 (N4076, N4066, N1766);
xor XOR2 (N4077, N4064, N2871);
nand NAND4 (N4078, N4076, N4038, N1410, N159);
nand NAND2 (N4079, N4052, N3545);
nor NOR2 (N4080, N4077, N2081);
or OR3 (N4081, N4075, N3711, N2887);
and AND3 (N4082, N4080, N964, N3558);
nand NAND2 (N4083, N4071, N2841);
buf BUF1 (N4084, N4082);
and AND4 (N4085, N4073, N2715, N506, N1885);
nor NOR4 (N4086, N4054, N1571, N494, N1039);
and AND4 (N4087, N4079, N2596, N282, N3852);
xor XOR2 (N4088, N4060, N3476);
nor NOR2 (N4089, N4087, N2881);
and AND3 (N4090, N4085, N662, N589);
xor XOR2 (N4091, N4090, N2497);
xor XOR2 (N4092, N4091, N1992);
or OR3 (N4093, N4092, N430, N2466);
xor XOR2 (N4094, N4055, N265);
nor NOR4 (N4095, N4089, N747, N1210, N3195);
buf BUF1 (N4096, N4093);
not NOT1 (N4097, N4096);
nand NAND3 (N4098, N4084, N1414, N365);
or OR2 (N4099, N4098, N1564);
and AND2 (N4100, N4095, N3605);
and AND3 (N4101, N4081, N2927, N2053);
and AND2 (N4102, N4083, N1928);
not NOT1 (N4103, N4088);
or OR3 (N4104, N4102, N3912, N1064);
not NOT1 (N4105, N4099);
xor XOR2 (N4106, N4070, N3966);
nor NOR3 (N4107, N4097, N935, N1701);
not NOT1 (N4108, N4104);
and AND2 (N4109, N4086, N124);
buf BUF1 (N4110, N4094);
nand NAND2 (N4111, N4105, N2593);
or OR3 (N4112, N4110, N1003, N794);
buf BUF1 (N4113, N4106);
buf BUF1 (N4114, N4113);
xor XOR2 (N4115, N4078, N1086);
nand NAND2 (N4116, N4111, N2532);
xor XOR2 (N4117, N4112, N3394);
and AND3 (N4118, N4107, N4064, N1050);
not NOT1 (N4119, N4117);
buf BUF1 (N4120, N4118);
not NOT1 (N4121, N4109);
nand NAND2 (N4122, N4121, N3057);
and AND4 (N4123, N4114, N714, N3336, N4119);
and AND4 (N4124, N927, N2251, N3437, N788);
not NOT1 (N4125, N4101);
nor NOR2 (N4126, N4115, N3978);
and AND3 (N4127, N4122, N919, N1268);
xor XOR2 (N4128, N4103, N3939);
nand NAND3 (N4129, N4100, N1637, N3414);
xor XOR2 (N4130, N4125, N3061);
and AND4 (N4131, N4120, N618, N1922, N2165);
buf BUF1 (N4132, N4130);
buf BUF1 (N4133, N4132);
not NOT1 (N4134, N4133);
or OR4 (N4135, N4124, N3600, N1259, N368);
nand NAND4 (N4136, N4135, N2036, N1524, N688);
or OR3 (N4137, N4129, N3270, N2849);
buf BUF1 (N4138, N4126);
and AND3 (N4139, N4116, N1759, N2715);
not NOT1 (N4140, N4123);
not NOT1 (N4141, N4140);
nor NOR3 (N4142, N4134, N93, N3010);
nor NOR2 (N4143, N4139, N2658);
nand NAND3 (N4144, N4108, N2292, N1182);
not NOT1 (N4145, N4136);
nand NAND2 (N4146, N4144, N3091);
and AND4 (N4147, N4146, N3185, N1191, N2048);
and AND2 (N4148, N4141, N1875);
buf BUF1 (N4149, N4128);
not NOT1 (N4150, N4145);
nor NOR3 (N4151, N4143, N3299, N1362);
and AND2 (N4152, N4148, N1999);
and AND3 (N4153, N4152, N768, N1586);
or OR3 (N4154, N4137, N1314, N2828);
nor NOR4 (N4155, N4151, N2369, N3252, N2000);
xor XOR2 (N4156, N4127, N2448);
and AND2 (N4157, N4131, N1432);
xor XOR2 (N4158, N4157, N2826);
nand NAND3 (N4159, N4153, N4081, N582);
nand NAND2 (N4160, N4147, N2554);
nor NOR4 (N4161, N4138, N408, N2786, N2043);
and AND4 (N4162, N4150, N4003, N1792, N686);
nand NAND3 (N4163, N4149, N2624, N913);
nor NOR2 (N4164, N4162, N3714);
and AND4 (N4165, N4159, N2372, N483, N2675);
not NOT1 (N4166, N4142);
not NOT1 (N4167, N4165);
xor XOR2 (N4168, N4166, N2316);
nor NOR4 (N4169, N4160, N3864, N1343, N7);
or OR3 (N4170, N4168, N2081, N522);
or OR2 (N4171, N4167, N75);
nand NAND3 (N4172, N4161, N411, N2307);
and AND3 (N4173, N4158, N1926, N369);
buf BUF1 (N4174, N4170);
nand NAND4 (N4175, N4156, N2888, N174, N4007);
buf BUF1 (N4176, N4173);
not NOT1 (N4177, N4164);
buf BUF1 (N4178, N4175);
not NOT1 (N4179, N4155);
or OR3 (N4180, N4176, N3648, N2569);
nand NAND4 (N4181, N4179, N1136, N2735, N412);
or OR3 (N4182, N4174, N3527, N1960);
nor NOR3 (N4183, N4169, N485, N1761);
nand NAND2 (N4184, N4180, N1235);
buf BUF1 (N4185, N4172);
not NOT1 (N4186, N4185);
nand NAND3 (N4187, N4171, N2048, N1772);
xor XOR2 (N4188, N4181, N1408);
and AND4 (N4189, N4183, N3383, N2515, N907);
xor XOR2 (N4190, N4163, N3384);
nand NAND3 (N4191, N4188, N2830, N3861);
nand NAND4 (N4192, N4190, N1778, N2834, N3177);
and AND2 (N4193, N4177, N2778);
nor NOR3 (N4194, N4178, N1295, N1156);
nor NOR3 (N4195, N4192, N831, N571);
and AND4 (N4196, N4194, N3928, N1435, N724);
xor XOR2 (N4197, N4191, N662);
or OR4 (N4198, N4186, N398, N3126, N663);
not NOT1 (N4199, N4198);
and AND3 (N4200, N4154, N3796, N360);
not NOT1 (N4201, N4193);
not NOT1 (N4202, N4184);
xor XOR2 (N4203, N4187, N3919);
and AND4 (N4204, N4197, N2698, N384, N4133);
buf BUF1 (N4205, N4182);
or OR3 (N4206, N4203, N1633, N3466);
xor XOR2 (N4207, N4206, N1244);
or OR3 (N4208, N4195, N801, N2715);
xor XOR2 (N4209, N4207, N4026);
xor XOR2 (N4210, N4205, N926);
not NOT1 (N4211, N4210);
buf BUF1 (N4212, N4211);
xor XOR2 (N4213, N4189, N3789);
xor XOR2 (N4214, N4204, N3097);
or OR4 (N4215, N4212, N3919, N692, N2041);
nand NAND4 (N4216, N4214, N2073, N630, N2263);
not NOT1 (N4217, N4213);
and AND2 (N4218, N4216, N2397);
and AND4 (N4219, N4199, N2233, N3147, N3676);
nor NOR2 (N4220, N4209, N1141);
not NOT1 (N4221, N4202);
not NOT1 (N4222, N4218);
xor XOR2 (N4223, N4215, N1939);
nor NOR3 (N4224, N4208, N2870, N3474);
nand NAND3 (N4225, N4196, N1957, N2472);
or OR3 (N4226, N4200, N1138, N3546);
nor NOR3 (N4227, N4224, N715, N554);
buf BUF1 (N4228, N4219);
nand NAND3 (N4229, N4220, N1700, N188);
not NOT1 (N4230, N4221);
xor XOR2 (N4231, N4229, N1687);
or OR4 (N4232, N4222, N2255, N2173, N329);
buf BUF1 (N4233, N4217);
nand NAND3 (N4234, N4232, N833, N1060);
not NOT1 (N4235, N4225);
nand NAND2 (N4236, N4228, N1650);
and AND2 (N4237, N4201, N579);
xor XOR2 (N4238, N4233, N2920);
and AND3 (N4239, N4226, N1323, N2050);
or OR2 (N4240, N4234, N3305);
and AND2 (N4241, N4223, N3443);
buf BUF1 (N4242, N4230);
buf BUF1 (N4243, N4242);
or OR4 (N4244, N4243, N951, N4221, N73);
nand NAND4 (N4245, N4241, N2463, N4074, N2434);
xor XOR2 (N4246, N4238, N865);
buf BUF1 (N4247, N4235);
and AND4 (N4248, N4236, N1228, N204, N4178);
and AND3 (N4249, N4231, N2049, N2475);
nand NAND2 (N4250, N4237, N3394);
and AND2 (N4251, N4239, N1615);
buf BUF1 (N4252, N4251);
nor NOR4 (N4253, N4227, N2660, N491, N202);
nor NOR4 (N4254, N4246, N504, N1627, N1096);
or OR2 (N4255, N4245, N2050);
not NOT1 (N4256, N4248);
and AND3 (N4257, N4252, N1676, N579);
buf BUF1 (N4258, N4249);
xor XOR2 (N4259, N4255, N1774);
buf BUF1 (N4260, N4244);
nor NOR3 (N4261, N4240, N4248, N1784);
not NOT1 (N4262, N4260);
xor XOR2 (N4263, N4257, N3450);
or OR4 (N4264, N4258, N911, N712, N3141);
xor XOR2 (N4265, N4263, N3777);
not NOT1 (N4266, N4259);
or OR2 (N4267, N4250, N1237);
xor XOR2 (N4268, N4262, N1482);
not NOT1 (N4269, N4264);
buf BUF1 (N4270, N4254);
and AND3 (N4271, N4270, N2576, N3830);
buf BUF1 (N4272, N4265);
or OR4 (N4273, N4271, N1086, N2137, N1438);
not NOT1 (N4274, N4272);
xor XOR2 (N4275, N4247, N3926);
xor XOR2 (N4276, N4275, N2845);
and AND2 (N4277, N4256, N1062);
buf BUF1 (N4278, N4276);
nand NAND2 (N4279, N4274, N3872);
nand NAND3 (N4280, N4269, N450, N3967);
or OR3 (N4281, N4261, N4261, N2810);
buf BUF1 (N4282, N4273);
buf BUF1 (N4283, N4281);
nand NAND2 (N4284, N4278, N3884);
nor NOR4 (N4285, N4279, N3256, N1028, N1296);
buf BUF1 (N4286, N4280);
xor XOR2 (N4287, N4284, N241);
buf BUF1 (N4288, N4268);
xor XOR2 (N4289, N4286, N1663);
xor XOR2 (N4290, N4282, N1774);
buf BUF1 (N4291, N4289);
xor XOR2 (N4292, N4253, N410);
or OR4 (N4293, N4288, N3974, N2934, N3719);
not NOT1 (N4294, N4293);
or OR3 (N4295, N4291, N1036, N145);
nand NAND4 (N4296, N4294, N890, N1920, N596);
not NOT1 (N4297, N4292);
not NOT1 (N4298, N4295);
or OR4 (N4299, N4287, N1465, N1875, N1013);
xor XOR2 (N4300, N4266, N2056);
xor XOR2 (N4301, N4300, N2167);
xor XOR2 (N4302, N4299, N2818);
nor NOR4 (N4303, N4297, N3910, N1841, N400);
or OR3 (N4304, N4290, N3302, N3232);
not NOT1 (N4305, N4304);
not NOT1 (N4306, N4285);
buf BUF1 (N4307, N4283);
nand NAND3 (N4308, N4302, N4059, N4120);
and AND4 (N4309, N4303, N4294, N2131, N824);
nand NAND4 (N4310, N4298, N2054, N1486, N527);
xor XOR2 (N4311, N4296, N4005);
not NOT1 (N4312, N4308);
nor NOR4 (N4313, N4305, N2843, N427, N2778);
nand NAND4 (N4314, N4310, N2210, N1650, N4184);
xor XOR2 (N4315, N4277, N2755);
not NOT1 (N4316, N4311);
nand NAND2 (N4317, N4301, N3295);
not NOT1 (N4318, N4306);
and AND3 (N4319, N4318, N168, N642);
and AND2 (N4320, N4317, N3352);
nand NAND2 (N4321, N4320, N1126);
xor XOR2 (N4322, N4309, N261);
or OR4 (N4323, N4322, N3202, N2217, N3836);
buf BUF1 (N4324, N4321);
buf BUF1 (N4325, N4319);
nand NAND4 (N4326, N4316, N1306, N4260, N1943);
and AND3 (N4327, N4307, N3628, N1177);
nor NOR3 (N4328, N4314, N2826, N3117);
and AND2 (N4329, N4312, N3773);
xor XOR2 (N4330, N4267, N4107);
buf BUF1 (N4331, N4330);
nor NOR4 (N4332, N4315, N767, N1769, N1819);
not NOT1 (N4333, N4326);
nand NAND3 (N4334, N4329, N2782, N800);
or OR3 (N4335, N4331, N3685, N3785);
nand NAND3 (N4336, N4313, N3594, N3836);
not NOT1 (N4337, N4336);
and AND2 (N4338, N4327, N2523);
nor NOR2 (N4339, N4335, N978);
or OR2 (N4340, N4339, N1900);
nor NOR3 (N4341, N4333, N4317, N329);
buf BUF1 (N4342, N4328);
not NOT1 (N4343, N4338);
buf BUF1 (N4344, N4324);
or OR2 (N4345, N4342, N4007);
and AND3 (N4346, N4345, N367, N3937);
and AND4 (N4347, N4341, N2100, N103, N2026);
nand NAND3 (N4348, N4347, N866, N2327);
nand NAND4 (N4349, N4334, N2553, N3937, N1043);
xor XOR2 (N4350, N4323, N474);
nand NAND2 (N4351, N4343, N3792);
not NOT1 (N4352, N4346);
nor NOR3 (N4353, N4350, N2774, N4043);
nor NOR2 (N4354, N4344, N3497);
nor NOR2 (N4355, N4353, N1716);
xor XOR2 (N4356, N4340, N2060);
or OR2 (N4357, N4325, N1043);
nand NAND4 (N4358, N4337, N2223, N414, N584);
or OR4 (N4359, N4354, N1147, N4174, N1032);
nor NOR4 (N4360, N4348, N3904, N2104, N4122);
and AND4 (N4361, N4349, N3532, N925, N2296);
buf BUF1 (N4362, N4360);
or OR2 (N4363, N4352, N775);
nor NOR4 (N4364, N4359, N228, N514, N3075);
or OR2 (N4365, N4357, N2388);
xor XOR2 (N4366, N4362, N900);
buf BUF1 (N4367, N4356);
nand NAND2 (N4368, N4364, N3875);
or OR2 (N4369, N4367, N1014);
xor XOR2 (N4370, N4369, N3330);
and AND4 (N4371, N4332, N3733, N909, N3804);
and AND2 (N4372, N4370, N2165);
nor NOR3 (N4373, N4355, N1162, N2487);
nor NOR3 (N4374, N4361, N3347, N1934);
and AND3 (N4375, N4365, N370, N3974);
xor XOR2 (N4376, N4368, N3536);
xor XOR2 (N4377, N4375, N3682);
buf BUF1 (N4378, N4376);
xor XOR2 (N4379, N4373, N2572);
nor NOR2 (N4380, N4372, N2425);
not NOT1 (N4381, N4363);
and AND3 (N4382, N4351, N2430, N1786);
nand NAND4 (N4383, N4380, N3316, N4200, N3252);
xor XOR2 (N4384, N4378, N689);
xor XOR2 (N4385, N4383, N698);
buf BUF1 (N4386, N4379);
nor NOR2 (N4387, N4366, N217);
xor XOR2 (N4388, N4381, N3837);
nand NAND4 (N4389, N4377, N2252, N1242, N1893);
buf BUF1 (N4390, N4387);
not NOT1 (N4391, N4374);
not NOT1 (N4392, N4386);
not NOT1 (N4393, N4358);
nor NOR3 (N4394, N4371, N2994, N2378);
or OR3 (N4395, N4392, N4120, N1723);
or OR4 (N4396, N4391, N3653, N364, N3263);
and AND3 (N4397, N4385, N1687, N2424);
or OR2 (N4398, N4390, N4129);
xor XOR2 (N4399, N4384, N2557);
not NOT1 (N4400, N4396);
nand NAND4 (N4401, N4399, N2164, N3619, N710);
and AND4 (N4402, N4397, N1808, N185, N1346);
not NOT1 (N4403, N4395);
buf BUF1 (N4404, N4402);
xor XOR2 (N4405, N4389, N2596);
not NOT1 (N4406, N4398);
not NOT1 (N4407, N4400);
nor NOR3 (N4408, N4406, N2229, N2455);
not NOT1 (N4409, N4393);
and AND3 (N4410, N4404, N1726, N3521);
buf BUF1 (N4411, N4394);
not NOT1 (N4412, N4409);
xor XOR2 (N4413, N4403, N2618);
xor XOR2 (N4414, N4413, N2781);
nand NAND4 (N4415, N4382, N2350, N3081, N1906);
not NOT1 (N4416, N4401);
and AND2 (N4417, N4388, N1850);
or OR4 (N4418, N4411, N1230, N4007, N3798);
or OR3 (N4419, N4412, N3424, N2978);
not NOT1 (N4420, N4405);
nand NAND3 (N4421, N4408, N1295, N3170);
nand NAND2 (N4422, N4407, N795);
nand NAND2 (N4423, N4415, N4040);
xor XOR2 (N4424, N4410, N1099);
nor NOR2 (N4425, N4422, N268);
nor NOR4 (N4426, N4423, N1522, N1797, N4073);
and AND2 (N4427, N4419, N3012);
nand NAND2 (N4428, N4424, N140);
and AND3 (N4429, N4414, N4258, N3025);
and AND2 (N4430, N4426, N3174);
not NOT1 (N4431, N4421);
buf BUF1 (N4432, N4431);
and AND3 (N4433, N4429, N1408, N3978);
xor XOR2 (N4434, N4418, N3982);
or OR4 (N4435, N4428, N2199, N4371, N1049);
nor NOR2 (N4436, N4420, N3924);
buf BUF1 (N4437, N4435);
nor NOR4 (N4438, N4430, N3520, N1479, N492);
nand NAND3 (N4439, N4416, N2461, N3833);
nor NOR3 (N4440, N4425, N1574, N1202);
nor NOR2 (N4441, N4434, N2753);
buf BUF1 (N4442, N4432);
or OR2 (N4443, N4441, N2820);
buf BUF1 (N4444, N4439);
or OR3 (N4445, N4438, N4248, N1089);
and AND3 (N4446, N4427, N2008, N2740);
and AND2 (N4447, N4442, N4163);
or OR2 (N4448, N4433, N1651);
buf BUF1 (N4449, N4448);
and AND2 (N4450, N4449, N4397);
xor XOR2 (N4451, N4444, N3928);
or OR2 (N4452, N4451, N1500);
buf BUF1 (N4453, N4436);
not NOT1 (N4454, N4450);
not NOT1 (N4455, N4445);
and AND4 (N4456, N4452, N2009, N4357, N929);
nand NAND3 (N4457, N4417, N2982, N2125);
nand NAND2 (N4458, N4440, N2112);
buf BUF1 (N4459, N4453);
nand NAND3 (N4460, N4437, N4015, N3192);
not NOT1 (N4461, N4457);
buf BUF1 (N4462, N4461);
xor XOR2 (N4463, N4459, N1543);
not NOT1 (N4464, N4455);
not NOT1 (N4465, N4443);
nand NAND4 (N4466, N4464, N3073, N1565, N244);
nand NAND3 (N4467, N4456, N1830, N3764);
and AND3 (N4468, N4447, N4067, N2651);
not NOT1 (N4469, N4468);
and AND2 (N4470, N4460, N1863);
nand NAND4 (N4471, N4458, N3768, N3371, N1121);
or OR4 (N4472, N4469, N3945, N2374, N3946);
nor NOR4 (N4473, N4446, N992, N431, N3279);
and AND3 (N4474, N4467, N2222, N66);
or OR4 (N4475, N4470, N2214, N34, N2520);
and AND4 (N4476, N4474, N875, N240, N1356);
or OR3 (N4477, N4462, N3864, N385);
nand NAND4 (N4478, N4472, N992, N3270, N784);
nor NOR4 (N4479, N4465, N2424, N747, N323);
not NOT1 (N4480, N4473);
nand NAND2 (N4481, N4480, N4423);
buf BUF1 (N4482, N4454);
buf BUF1 (N4483, N4475);
buf BUF1 (N4484, N4483);
nor NOR2 (N4485, N4466, N3756);
buf BUF1 (N4486, N4482);
xor XOR2 (N4487, N4486, N1156);
and AND3 (N4488, N4484, N1214, N2352);
or OR4 (N4489, N4479, N331, N1112, N4454);
nand NAND4 (N4490, N4487, N147, N4390, N2473);
buf BUF1 (N4491, N4489);
buf BUF1 (N4492, N4476);
or OR2 (N4493, N4490, N1135);
xor XOR2 (N4494, N4481, N2739);
or OR3 (N4495, N4471, N2908, N2360);
and AND3 (N4496, N4477, N2647, N3615);
not NOT1 (N4497, N4485);
nand NAND2 (N4498, N4478, N2001);
nor NOR3 (N4499, N4463, N4471, N1843);
not NOT1 (N4500, N4493);
or OR2 (N4501, N4497, N3884);
nor NOR4 (N4502, N4495, N3983, N3792, N541);
xor XOR2 (N4503, N4500, N3855);
nand NAND2 (N4504, N4492, N1815);
buf BUF1 (N4505, N4491);
nor NOR3 (N4506, N4494, N912, N326);
buf BUF1 (N4507, N4488);
and AND3 (N4508, N4502, N4397, N2633);
or OR2 (N4509, N4503, N3685);
nand NAND3 (N4510, N4509, N3742, N1467);
nor NOR4 (N4511, N4501, N2154, N3205, N1842);
and AND3 (N4512, N4499, N1105, N366);
buf BUF1 (N4513, N4508);
buf BUF1 (N4514, N4505);
xor XOR2 (N4515, N4510, N2749);
not NOT1 (N4516, N4514);
nand NAND4 (N4517, N4515, N2787, N2874, N4222);
or OR3 (N4518, N4512, N2307, N2223);
buf BUF1 (N4519, N4516);
nand NAND4 (N4520, N4496, N2477, N2415, N3247);
not NOT1 (N4521, N4507);
buf BUF1 (N4522, N4506);
nand NAND2 (N4523, N4518, N24);
nand NAND3 (N4524, N4504, N4252, N3928);
and AND3 (N4525, N4511, N3254, N993);
buf BUF1 (N4526, N4521);
xor XOR2 (N4527, N4525, N1178);
and AND2 (N4528, N4527, N2831);
nor NOR4 (N4529, N4526, N2970, N3295, N4471);
and AND3 (N4530, N4522, N1220, N142);
nor NOR2 (N4531, N4523, N2666);
and AND4 (N4532, N4498, N1617, N2872, N339);
buf BUF1 (N4533, N4528);
nor NOR4 (N4534, N4524, N3066, N799, N1459);
nand NAND3 (N4535, N4520, N4119, N532);
or OR4 (N4536, N4517, N210, N95, N2982);
xor XOR2 (N4537, N4513, N2438);
or OR2 (N4538, N4531, N4065);
buf BUF1 (N4539, N4532);
nor NOR2 (N4540, N4519, N1929);
buf BUF1 (N4541, N4535);
not NOT1 (N4542, N4529);
not NOT1 (N4543, N4541);
xor XOR2 (N4544, N4530, N1853);
and AND3 (N4545, N4533, N1320, N2814);
not NOT1 (N4546, N4538);
not NOT1 (N4547, N4546);
buf BUF1 (N4548, N4545);
not NOT1 (N4549, N4539);
nor NOR4 (N4550, N4537, N2884, N3909, N2971);
nor NOR3 (N4551, N4549, N4118, N1018);
or OR4 (N4552, N4540, N2908, N2637, N3552);
xor XOR2 (N4553, N4544, N353);
nor NOR4 (N4554, N4547, N3324, N2829, N1809);
and AND4 (N4555, N4543, N1059, N656, N311);
or OR2 (N4556, N4555, N557);
and AND2 (N4557, N4553, N829);
xor XOR2 (N4558, N4554, N4546);
xor XOR2 (N4559, N4551, N2158);
nor NOR4 (N4560, N4550, N2987, N2118, N3405);
buf BUF1 (N4561, N4536);
xor XOR2 (N4562, N4558, N3202);
nand NAND2 (N4563, N4548, N1840);
buf BUF1 (N4564, N4557);
and AND3 (N4565, N4560, N90, N1894);
xor XOR2 (N4566, N4562, N2126);
buf BUF1 (N4567, N4542);
nand NAND3 (N4568, N4552, N412, N3701);
and AND2 (N4569, N4567, N561);
xor XOR2 (N4570, N4534, N2721);
xor XOR2 (N4571, N4559, N699);
and AND4 (N4572, N4565, N1699, N3533, N3798);
not NOT1 (N4573, N4568);
or OR2 (N4574, N4556, N3108);
nand NAND4 (N4575, N4572, N1527, N1177, N221);
and AND3 (N4576, N4575, N3928, N178);
xor XOR2 (N4577, N4563, N4389);
or OR4 (N4578, N4561, N2617, N3983, N2028);
nand NAND3 (N4579, N4571, N3751, N2630);
or OR4 (N4580, N4574, N3293, N4056, N3200);
and AND4 (N4581, N4566, N169, N2830, N1900);
or OR3 (N4582, N4581, N4242, N3452);
not NOT1 (N4583, N4570);
buf BUF1 (N4584, N4580);
nor NOR2 (N4585, N4584, N2411);
nand NAND4 (N4586, N4585, N603, N899, N1063);
and AND3 (N4587, N4564, N3376, N4365);
and AND4 (N4588, N4582, N2586, N380, N327);
and AND4 (N4589, N4583, N3590, N4297, N3480);
nor NOR2 (N4590, N4577, N2964);
nor NOR4 (N4591, N4588, N3860, N2909, N3564);
not NOT1 (N4592, N4590);
xor XOR2 (N4593, N4579, N3831);
and AND4 (N4594, N4573, N4138, N1199, N2526);
xor XOR2 (N4595, N4589, N2197);
or OR4 (N4596, N4576, N2757, N3135, N1062);
not NOT1 (N4597, N4569);
or OR2 (N4598, N4593, N2679);
buf BUF1 (N4599, N4594);
or OR2 (N4600, N4599, N198);
buf BUF1 (N4601, N4595);
nand NAND4 (N4602, N4597, N2036, N89, N3419);
nor NOR2 (N4603, N4602, N895);
buf BUF1 (N4604, N4578);
and AND4 (N4605, N4596, N3841, N4149, N4462);
and AND4 (N4606, N4600, N34, N1031, N2711);
xor XOR2 (N4607, N4587, N1083);
or OR2 (N4608, N4603, N2472);
nand NAND3 (N4609, N4605, N407, N1574);
nand NAND2 (N4610, N4598, N3932);
buf BUF1 (N4611, N4609);
or OR3 (N4612, N4586, N286, N1928);
not NOT1 (N4613, N4607);
nand NAND4 (N4614, N4612, N3527, N4333, N3853);
and AND2 (N4615, N4608, N4339);
buf BUF1 (N4616, N4601);
or OR4 (N4617, N4616, N2832, N3884, N3496);
nor NOR2 (N4618, N4613, N1668);
nor NOR3 (N4619, N4615, N2062, N1544);
nand NAND2 (N4620, N4618, N1704);
not NOT1 (N4621, N4604);
buf BUF1 (N4622, N4617);
not NOT1 (N4623, N4620);
nor NOR3 (N4624, N4614, N239, N2226);
nand NAND2 (N4625, N4622, N1183);
and AND2 (N4626, N4611, N1843);
buf BUF1 (N4627, N4619);
and AND3 (N4628, N4591, N4431, N367);
nor NOR3 (N4629, N4626, N987, N3760);
or OR4 (N4630, N4628, N3037, N4167, N576);
xor XOR2 (N4631, N4625, N3080);
nor NOR3 (N4632, N4627, N2679, N1897);
or OR3 (N4633, N4631, N960, N572);
and AND4 (N4634, N4633, N3662, N2139, N649);
not NOT1 (N4635, N4606);
or OR3 (N4636, N4624, N2924, N2704);
nand NAND4 (N4637, N4621, N4365, N2528, N361);
and AND4 (N4638, N4634, N2447, N1549, N2946);
xor XOR2 (N4639, N4636, N3997);
buf BUF1 (N4640, N4592);
not NOT1 (N4641, N4637);
nand NAND3 (N4642, N4630, N946, N1005);
nand NAND2 (N4643, N4639, N2347);
buf BUF1 (N4644, N4642);
and AND2 (N4645, N4638, N2009);
nor NOR3 (N4646, N4635, N550, N2275);
not NOT1 (N4647, N4629);
buf BUF1 (N4648, N4640);
and AND4 (N4649, N4646, N3379, N3214, N3949);
nand NAND4 (N4650, N4632, N2637, N1833, N3300);
nor NOR4 (N4651, N4649, N1112, N2824, N1220);
nand NAND2 (N4652, N4643, N1932);
buf BUF1 (N4653, N4647);
buf BUF1 (N4654, N4650);
xor XOR2 (N4655, N4645, N3904);
nand NAND2 (N4656, N4652, N935);
xor XOR2 (N4657, N4655, N1346);
or OR2 (N4658, N4657, N3985);
nand NAND3 (N4659, N4658, N2877, N1701);
or OR3 (N4660, N4659, N1078, N3202);
not NOT1 (N4661, N4660);
nor NOR2 (N4662, N4661, N256);
nand NAND4 (N4663, N4644, N2365, N4189, N671);
xor XOR2 (N4664, N4610, N2597);
nor NOR2 (N4665, N4654, N4302);
nor NOR2 (N4666, N4651, N4208);
xor XOR2 (N4667, N4663, N4523);
nand NAND2 (N4668, N4667, N2606);
not NOT1 (N4669, N4653);
and AND3 (N4670, N4669, N532, N3372);
buf BUF1 (N4671, N4664);
or OR3 (N4672, N4670, N529, N2463);
and AND2 (N4673, N4671, N356);
or OR4 (N4674, N4656, N1145, N2135, N2781);
buf BUF1 (N4675, N4665);
nand NAND2 (N4676, N4672, N3125);
not NOT1 (N4677, N4641);
buf BUF1 (N4678, N4674);
or OR3 (N4679, N4677, N1276, N2082);
nand NAND3 (N4680, N4668, N4037, N3102);
xor XOR2 (N4681, N4623, N4355);
xor XOR2 (N4682, N4681, N1198);
buf BUF1 (N4683, N4680);
xor XOR2 (N4684, N4666, N4457);
or OR2 (N4685, N4662, N6);
nor NOR2 (N4686, N4679, N3817);
nor NOR2 (N4687, N4683, N4359);
and AND2 (N4688, N4687, N2638);
buf BUF1 (N4689, N4686);
xor XOR2 (N4690, N4688, N1527);
buf BUF1 (N4691, N4673);
nor NOR2 (N4692, N4682, N1579);
or OR2 (N4693, N4648, N1427);
not NOT1 (N4694, N4693);
buf BUF1 (N4695, N4692);
and AND3 (N4696, N4690, N4555, N2843);
xor XOR2 (N4697, N4678, N797);
or OR2 (N4698, N4689, N1480);
xor XOR2 (N4699, N4695, N2341);
or OR3 (N4700, N4696, N2974, N18);
not NOT1 (N4701, N4700);
nand NAND3 (N4702, N4699, N919, N1316);
buf BUF1 (N4703, N4702);
or OR3 (N4704, N4694, N2968, N2146);
not NOT1 (N4705, N4701);
or OR4 (N4706, N4684, N2839, N1301, N1135);
or OR4 (N4707, N4706, N2221, N409, N2326);
not NOT1 (N4708, N4703);
nor NOR4 (N4709, N4685, N555, N1964, N1579);
or OR3 (N4710, N4698, N1716, N96);
or OR4 (N4711, N4707, N4373, N12, N386);
nand NAND3 (N4712, N4675, N3047, N276);
not NOT1 (N4713, N4712);
or OR3 (N4714, N4676, N4682, N1989);
buf BUF1 (N4715, N4711);
nand NAND2 (N4716, N4709, N1599);
nand NAND4 (N4717, N4697, N2346, N2708, N192);
nand NAND4 (N4718, N4691, N508, N1668, N345);
and AND3 (N4719, N4705, N3008, N2629);
and AND4 (N4720, N4719, N2731, N4673, N1332);
buf BUF1 (N4721, N4718);
xor XOR2 (N4722, N4704, N1388);
xor XOR2 (N4723, N4708, N4363);
nand NAND2 (N4724, N4716, N625);
nand NAND4 (N4725, N4721, N4611, N576, N3350);
nor NOR3 (N4726, N4724, N3389, N2226);
nor NOR2 (N4727, N4715, N2064);
or OR4 (N4728, N4710, N3438, N3532, N497);
nor NOR3 (N4729, N4717, N3022, N3632);
not NOT1 (N4730, N4722);
buf BUF1 (N4731, N4720);
or OR3 (N4732, N4725, N2346, N4180);
nand NAND4 (N4733, N4729, N1662, N4128, N379);
or OR3 (N4734, N4726, N1224, N1009);
or OR3 (N4735, N4732, N1950, N280);
and AND2 (N4736, N4714, N3825);
or OR4 (N4737, N4728, N1284, N3681, N3008);
nor NOR2 (N4738, N4730, N511);
nor NOR2 (N4739, N4733, N3901);
and AND2 (N4740, N4735, N3140);
not NOT1 (N4741, N4727);
nor NOR3 (N4742, N4738, N67, N1548);
and AND4 (N4743, N4713, N4393, N3590, N4577);
not NOT1 (N4744, N4739);
nor NOR4 (N4745, N4741, N3285, N309, N1954);
xor XOR2 (N4746, N4744, N264);
nand NAND2 (N4747, N4731, N4297);
nor NOR3 (N4748, N4742, N2931, N4276);
or OR4 (N4749, N4734, N3065, N4077, N2122);
xor XOR2 (N4750, N4745, N473);
or OR2 (N4751, N4723, N209);
or OR2 (N4752, N4746, N1114);
not NOT1 (N4753, N4740);
or OR4 (N4754, N4736, N4512, N189, N768);
buf BUF1 (N4755, N4743);
and AND2 (N4756, N4747, N1514);
nand NAND3 (N4757, N4756, N1073, N4065);
or OR4 (N4758, N4750, N1161, N4528, N1830);
not NOT1 (N4759, N4748);
xor XOR2 (N4760, N4755, N3002);
nor NOR4 (N4761, N4753, N3227, N3367, N3403);
not NOT1 (N4762, N4752);
buf BUF1 (N4763, N4762);
and AND3 (N4764, N4737, N4744, N2384);
not NOT1 (N4765, N4751);
not NOT1 (N4766, N4761);
or OR4 (N4767, N4766, N2718, N2641, N211);
and AND3 (N4768, N4767, N4473, N39);
buf BUF1 (N4769, N4763);
or OR4 (N4770, N4769, N3771, N4684, N4396);
nand NAND4 (N4771, N4770, N1649, N3473, N3997);
buf BUF1 (N4772, N4758);
or OR2 (N4773, N4760, N1143);
buf BUF1 (N4774, N4772);
nor NOR3 (N4775, N4754, N664, N2293);
nand NAND4 (N4776, N4749, N4699, N3031, N191);
not NOT1 (N4777, N4765);
buf BUF1 (N4778, N4768);
xor XOR2 (N4779, N4777, N3765);
xor XOR2 (N4780, N4776, N3188);
or OR3 (N4781, N4780, N4212, N4551);
or OR4 (N4782, N4764, N1179, N4670, N3702);
xor XOR2 (N4783, N4779, N1650);
buf BUF1 (N4784, N4782);
and AND3 (N4785, N4778, N2932, N3867);
and AND4 (N4786, N4773, N2342, N2560, N3072);
buf BUF1 (N4787, N4786);
buf BUF1 (N4788, N4775);
and AND3 (N4789, N4783, N391, N682);
or OR4 (N4790, N4789, N1769, N1856, N3553);
nand NAND3 (N4791, N4790, N1180, N4065);
or OR2 (N4792, N4788, N4653);
or OR3 (N4793, N4759, N4105, N726);
not NOT1 (N4794, N4774);
not NOT1 (N4795, N4791);
not NOT1 (N4796, N4781);
not NOT1 (N4797, N4792);
nand NAND2 (N4798, N4771, N885);
nor NOR2 (N4799, N4757, N2053);
not NOT1 (N4800, N4795);
and AND3 (N4801, N4796, N1275, N3411);
nor NOR4 (N4802, N4784, N714, N4267, N805);
nand NAND2 (N4803, N4794, N1812);
nand NAND3 (N4804, N4800, N2857, N1834);
nand NAND2 (N4805, N4797, N1801);
or OR4 (N4806, N4802, N1559, N1338, N4567);
nor NOR4 (N4807, N4801, N2289, N1818, N1364);
xor XOR2 (N4808, N4798, N735);
buf BUF1 (N4809, N4793);
or OR4 (N4810, N4803, N2361, N425, N1342);
or OR4 (N4811, N4806, N1593, N4361, N4040);
xor XOR2 (N4812, N4810, N1859);
or OR4 (N4813, N4787, N1395, N4238, N1155);
buf BUF1 (N4814, N4805);
and AND2 (N4815, N4813, N3585);
nor NOR3 (N4816, N4814, N1828, N4057);
xor XOR2 (N4817, N4807, N2415);
not NOT1 (N4818, N4815);
and AND4 (N4819, N4812, N1077, N4678, N1669);
nand NAND4 (N4820, N4809, N1289, N2649, N4106);
nand NAND3 (N4821, N4785, N3390, N1965);
nor NOR4 (N4822, N4820, N1734, N3109, N626);
or OR2 (N4823, N4816, N2041);
xor XOR2 (N4824, N4818, N1993);
nor NOR3 (N4825, N4822, N2579, N1560);
nand NAND3 (N4826, N4811, N1266, N3928);
or OR4 (N4827, N4808, N1702, N729, N3308);
and AND2 (N4828, N4799, N2635);
or OR4 (N4829, N4804, N364, N1907, N598);
not NOT1 (N4830, N4819);
nor NOR3 (N4831, N4817, N2537, N3819);
not NOT1 (N4832, N4826);
not NOT1 (N4833, N4821);
buf BUF1 (N4834, N4833);
not NOT1 (N4835, N4832);
not NOT1 (N4836, N4825);
buf BUF1 (N4837, N4834);
xor XOR2 (N4838, N4837, N1330);
xor XOR2 (N4839, N4828, N2099);
nor NOR4 (N4840, N4830, N750, N3348, N445);
and AND4 (N4841, N4836, N2434, N4820, N4104);
buf BUF1 (N4842, N4831);
xor XOR2 (N4843, N4839, N624);
buf BUF1 (N4844, N4842);
xor XOR2 (N4845, N4840, N2835);
nor NOR2 (N4846, N4844, N1408);
buf BUF1 (N4847, N4827);
xor XOR2 (N4848, N4846, N2853);
nand NAND3 (N4849, N4843, N1340, N2309);
xor XOR2 (N4850, N4841, N4196);
or OR2 (N4851, N4824, N4062);
xor XOR2 (N4852, N4838, N4277);
not NOT1 (N4853, N4852);
xor XOR2 (N4854, N4848, N2307);
buf BUF1 (N4855, N4829);
nor NOR3 (N4856, N4855, N3526, N4787);
and AND3 (N4857, N4823, N146, N892);
nor NOR4 (N4858, N4851, N1469, N1948, N762);
or OR3 (N4859, N4847, N2808, N2627);
buf BUF1 (N4860, N4850);
not NOT1 (N4861, N4854);
nor NOR2 (N4862, N4835, N77);
buf BUF1 (N4863, N4861);
or OR2 (N4864, N4845, N172);
and AND4 (N4865, N4862, N2310, N3901, N1858);
nand NAND3 (N4866, N4849, N765, N3017);
xor XOR2 (N4867, N4866, N3710);
xor XOR2 (N4868, N4867, N112);
nor NOR3 (N4869, N4856, N1106, N3683);
and AND4 (N4870, N4858, N130, N3327, N3900);
xor XOR2 (N4871, N4869, N880);
not NOT1 (N4872, N4871);
or OR3 (N4873, N4865, N1527, N3910);
and AND3 (N4874, N4860, N4399, N4328);
nor NOR3 (N4875, N4872, N4417, N3422);
nand NAND4 (N4876, N4857, N3183, N3552, N1729);
not NOT1 (N4877, N4863);
xor XOR2 (N4878, N4859, N3702);
buf BUF1 (N4879, N4877);
xor XOR2 (N4880, N4864, N3068);
nor NOR4 (N4881, N4874, N4238, N3294, N2380);
nand NAND2 (N4882, N4870, N1728);
buf BUF1 (N4883, N4882);
buf BUF1 (N4884, N4873);
xor XOR2 (N4885, N4875, N4042);
buf BUF1 (N4886, N4884);
xor XOR2 (N4887, N4853, N1646);
and AND4 (N4888, N4881, N3208, N3428, N1939);
xor XOR2 (N4889, N4879, N3602);
nand NAND4 (N4890, N4880, N4764, N1467, N3625);
and AND3 (N4891, N4876, N1075, N1777);
and AND2 (N4892, N4883, N3826);
and AND3 (N4893, N4891, N3488, N4762);
not NOT1 (N4894, N4888);
and AND4 (N4895, N4878, N4120, N2879, N1348);
xor XOR2 (N4896, N4890, N17);
or OR4 (N4897, N4896, N2227, N2601, N2131);
and AND4 (N4898, N4893, N980, N1549, N3333);
nand NAND4 (N4899, N4885, N1644, N1300, N3007);
nand NAND3 (N4900, N4868, N1348, N613);
not NOT1 (N4901, N4887);
and AND3 (N4902, N4889, N2842, N578);
xor XOR2 (N4903, N4894, N1109);
not NOT1 (N4904, N4903);
not NOT1 (N4905, N4899);
not NOT1 (N4906, N4892);
and AND4 (N4907, N4904, N426, N737, N811);
not NOT1 (N4908, N4902);
xor XOR2 (N4909, N4907, N4491);
buf BUF1 (N4910, N4906);
nor NOR4 (N4911, N4900, N2085, N1480, N279);
not NOT1 (N4912, N4897);
xor XOR2 (N4913, N4912, N1381);
and AND3 (N4914, N4908, N4411, N2731);
nand NAND3 (N4915, N4913, N301, N4910);
not NOT1 (N4916, N524);
or OR4 (N4917, N4895, N451, N3020, N312);
or OR4 (N4918, N4886, N1635, N3848, N1179);
not NOT1 (N4919, N4911);
and AND2 (N4920, N4915, N2501);
buf BUF1 (N4921, N4909);
nor NOR2 (N4922, N4905, N1755);
nand NAND3 (N4923, N4898, N3801, N2431);
nor NOR3 (N4924, N4921, N4455, N2564);
and AND4 (N4925, N4923, N4708, N1935, N4915);
nand NAND2 (N4926, N4924, N2319);
and AND2 (N4927, N4916, N3299);
and AND2 (N4928, N4926, N4865);
and AND2 (N4929, N4901, N1001);
nand NAND3 (N4930, N4925, N391, N1751);
not NOT1 (N4931, N4920);
or OR2 (N4932, N4918, N4068);
and AND4 (N4933, N4928, N1294, N650, N1000);
xor XOR2 (N4934, N4927, N533);
nor NOR2 (N4935, N4932, N699);
nor NOR2 (N4936, N4934, N3245);
not NOT1 (N4937, N4931);
nand NAND4 (N4938, N4935, N2702, N2232, N204);
nand NAND3 (N4939, N4938, N451, N2397);
or OR3 (N4940, N4914, N3845, N3084);
nand NAND2 (N4941, N4919, N2577);
or OR2 (N4942, N4937, N1449);
and AND2 (N4943, N4939, N3769);
buf BUF1 (N4944, N4942);
nand NAND2 (N4945, N4943, N112);
or OR3 (N4946, N4936, N2502, N3621);
nor NOR2 (N4947, N4929, N2538);
xor XOR2 (N4948, N4945, N1810);
and AND4 (N4949, N4946, N83, N1718, N3130);
nor NOR4 (N4950, N4930, N4067, N753, N4756);
and AND4 (N4951, N4944, N3873, N1307, N125);
nand NAND2 (N4952, N4947, N888);
not NOT1 (N4953, N4948);
nand NAND2 (N4954, N4953, N3199);
nand NAND2 (N4955, N4951, N1410);
nand NAND4 (N4956, N4922, N965, N3459, N3442);
or OR2 (N4957, N4933, N2384);
nand NAND2 (N4958, N4955, N1811);
xor XOR2 (N4959, N4954, N4695);
xor XOR2 (N4960, N4959, N4957);
xor XOR2 (N4961, N926, N2167);
not NOT1 (N4962, N4949);
buf BUF1 (N4963, N4941);
not NOT1 (N4964, N4950);
not NOT1 (N4965, N4952);
nor NOR3 (N4966, N4964, N4399, N842);
and AND2 (N4967, N4940, N2046);
and AND4 (N4968, N4967, N1365, N4323, N1157);
nor NOR2 (N4969, N4966, N4769);
nand NAND2 (N4970, N4958, N653);
or OR3 (N4971, N4961, N2428, N3559);
not NOT1 (N4972, N4970);
xor XOR2 (N4973, N4956, N4509);
nand NAND2 (N4974, N4917, N2708);
or OR4 (N4975, N4968, N3256, N1554, N2816);
buf BUF1 (N4976, N4960);
nor NOR2 (N4977, N4963, N570);
and AND3 (N4978, N4977, N3017, N2927);
and AND4 (N4979, N4962, N4967, N2525, N3282);
xor XOR2 (N4980, N4974, N1773);
not NOT1 (N4981, N4979);
xor XOR2 (N4982, N4975, N1836);
not NOT1 (N4983, N4981);
not NOT1 (N4984, N4980);
and AND2 (N4985, N4965, N2868);
and AND2 (N4986, N4983, N1892);
or OR2 (N4987, N4971, N898);
buf BUF1 (N4988, N4985);
xor XOR2 (N4989, N4973, N154);
nand NAND2 (N4990, N4987, N641);
xor XOR2 (N4991, N4990, N971);
and AND2 (N4992, N4976, N2928);
xor XOR2 (N4993, N4991, N4607);
nand NAND3 (N4994, N4969, N1006, N1753);
nand NAND2 (N4995, N4978, N4439);
or OR2 (N4996, N4988, N4850);
nand NAND2 (N4997, N4992, N3443);
and AND3 (N4998, N4996, N725, N3210);
nor NOR4 (N4999, N4972, N511, N1074, N1031);
buf BUF1 (N5000, N4989);
xor XOR2 (N5001, N4999, N1848);
xor XOR2 (N5002, N5001, N1422);
and AND3 (N5003, N4994, N829, N1516);
nor NOR2 (N5004, N5000, N2925);
nand NAND2 (N5005, N5002, N3585);
not NOT1 (N5006, N4993);
not NOT1 (N5007, N5003);
not NOT1 (N5008, N5006);
not NOT1 (N5009, N4984);
nand NAND3 (N5010, N4982, N2786, N3722);
buf BUF1 (N5011, N5005);
xor XOR2 (N5012, N5010, N1200);
buf BUF1 (N5013, N5007);
nor NOR2 (N5014, N4995, N3080);
xor XOR2 (N5015, N4997, N2904);
nor NOR3 (N5016, N4998, N229, N576);
or OR2 (N5017, N5009, N318);
or OR2 (N5018, N5004, N3267);
nand NAND4 (N5019, N5018, N1782, N707, N4582);
nor NOR4 (N5020, N5016, N1536, N1798, N3794);
nor NOR3 (N5021, N4986, N4139, N74);
not NOT1 (N5022, N5012);
buf BUF1 (N5023, N5015);
nor NOR2 (N5024, N5014, N4447);
not NOT1 (N5025, N5022);
xor XOR2 (N5026, N5023, N4131);
or OR4 (N5027, N5021, N3728, N1324, N3247);
nand NAND4 (N5028, N5013, N3056, N1857, N4974);
buf BUF1 (N5029, N5025);
nand NAND3 (N5030, N5017, N1407, N4224);
buf BUF1 (N5031, N5024);
or OR2 (N5032, N5029, N2795);
not NOT1 (N5033, N5031);
or OR4 (N5034, N5028, N4765, N4032, N4952);
buf BUF1 (N5035, N5032);
xor XOR2 (N5036, N5020, N3789);
buf BUF1 (N5037, N5019);
and AND2 (N5038, N5035, N1977);
nor NOR4 (N5039, N5026, N4719, N1643, N1340);
nor NOR2 (N5040, N5036, N104);
xor XOR2 (N5041, N5008, N3355);
and AND4 (N5042, N5040, N2844, N522, N2586);
nor NOR2 (N5043, N5039, N3913);
nor NOR2 (N5044, N5042, N137);
nor NOR2 (N5045, N5041, N3905);
xor XOR2 (N5046, N5027, N4640);
xor XOR2 (N5047, N5043, N3579);
and AND2 (N5048, N5033, N3217);
or OR4 (N5049, N5046, N664, N1265, N3335);
or OR2 (N5050, N5011, N1584);
nor NOR4 (N5051, N5049, N1818, N3324, N1241);
nand NAND4 (N5052, N5051, N3032, N1527, N1700);
buf BUF1 (N5053, N5044);
not NOT1 (N5054, N5045);
or OR3 (N5055, N5047, N4289, N3171);
and AND2 (N5056, N5052, N598);
not NOT1 (N5057, N5030);
and AND4 (N5058, N5057, N3931, N374, N4506);
nand NAND3 (N5059, N5037, N3367, N2836);
and AND2 (N5060, N5050, N4641);
nor NOR3 (N5061, N5048, N2390, N295);
nand NAND3 (N5062, N5038, N3621, N4565);
or OR2 (N5063, N5058, N4350);
and AND2 (N5064, N5053, N2190);
nor NOR4 (N5065, N5034, N1006, N2684, N4138);
not NOT1 (N5066, N5064);
buf BUF1 (N5067, N5059);
or OR2 (N5068, N5065, N2679);
not NOT1 (N5069, N5054);
and AND4 (N5070, N5068, N2606, N1209, N2124);
buf BUF1 (N5071, N5062);
xor XOR2 (N5072, N5060, N2128);
and AND4 (N5073, N5069, N3119, N875, N3132);
nor NOR2 (N5074, N5056, N1475);
xor XOR2 (N5075, N5063, N4442);
nand NAND4 (N5076, N5066, N1767, N75, N1246);
buf BUF1 (N5077, N5072);
nand NAND2 (N5078, N5075, N188);
not NOT1 (N5079, N5055);
nor NOR3 (N5080, N5073, N3076, N4589);
or OR4 (N5081, N5078, N1935, N1962, N2251);
nand NAND3 (N5082, N5081, N4292, N3773);
and AND4 (N5083, N5067, N172, N4253, N1567);
nand NAND2 (N5084, N5077, N4581);
nand NAND4 (N5085, N5076, N1521, N4209, N4278);
nand NAND3 (N5086, N5061, N1830, N728);
xor XOR2 (N5087, N5084, N3530);
buf BUF1 (N5088, N5071);
xor XOR2 (N5089, N5088, N3970);
buf BUF1 (N5090, N5083);
and AND4 (N5091, N5080, N2464, N3278, N2462);
nor NOR3 (N5092, N5079, N456, N460);
xor XOR2 (N5093, N5082, N2119);
buf BUF1 (N5094, N5091);
nor NOR3 (N5095, N5086, N3536, N4847);
nor NOR4 (N5096, N5089, N4101, N4527, N2226);
nand NAND3 (N5097, N5070, N2743, N4361);
or OR3 (N5098, N5097, N1903, N507);
xor XOR2 (N5099, N5093, N3499);
nor NOR4 (N5100, N5087, N2770, N3916, N4591);
and AND2 (N5101, N5094, N2897);
xor XOR2 (N5102, N5101, N1352);
nor NOR3 (N5103, N5095, N906, N4242);
xor XOR2 (N5104, N5074, N196);
not NOT1 (N5105, N5104);
and AND4 (N5106, N5099, N3150, N1552, N4709);
not NOT1 (N5107, N5096);
or OR3 (N5108, N5090, N753, N345);
or OR2 (N5109, N5105, N4868);
and AND2 (N5110, N5098, N635);
not NOT1 (N5111, N5103);
nand NAND2 (N5112, N5102, N3066);
or OR3 (N5113, N5085, N1335, N1765);
and AND3 (N5114, N5109, N3863, N2961);
xor XOR2 (N5115, N5112, N662);
nor NOR2 (N5116, N5110, N250);
nor NOR4 (N5117, N5108, N749, N1167, N3203);
buf BUF1 (N5118, N5107);
xor XOR2 (N5119, N5100, N266);
not NOT1 (N5120, N5106);
xor XOR2 (N5121, N5092, N1845);
nor NOR4 (N5122, N5115, N1026, N4673, N3856);
nand NAND3 (N5123, N5117, N4081, N878);
and AND2 (N5124, N5118, N2835);
buf BUF1 (N5125, N5124);
and AND3 (N5126, N5119, N3643, N2114);
xor XOR2 (N5127, N5122, N2532);
not NOT1 (N5128, N5113);
not NOT1 (N5129, N5111);
nor NOR4 (N5130, N5116, N960, N1026, N2500);
and AND3 (N5131, N5128, N1725, N2777);
and AND2 (N5132, N5114, N2543);
and AND4 (N5133, N5130, N976, N3984, N3378);
buf BUF1 (N5134, N5127);
and AND4 (N5135, N5120, N2630, N2394, N852);
and AND3 (N5136, N5125, N289, N2415);
xor XOR2 (N5137, N5133, N5078);
not NOT1 (N5138, N5132);
nand NAND4 (N5139, N5138, N747, N4473, N363);
nand NAND2 (N5140, N5123, N3340);
not NOT1 (N5141, N5139);
nand NAND3 (N5142, N5129, N2673, N4339);
not NOT1 (N5143, N5131);
xor XOR2 (N5144, N5136, N1845);
not NOT1 (N5145, N5134);
nand NAND3 (N5146, N5141, N2234, N1778);
nand NAND3 (N5147, N5145, N2945, N880);
nor NOR4 (N5148, N5146, N1915, N3290, N1868);
buf BUF1 (N5149, N5140);
xor XOR2 (N5150, N5126, N4969);
buf BUF1 (N5151, N5149);
and AND3 (N5152, N5142, N2443, N4130);
nor NOR4 (N5153, N5151, N582, N550, N3342);
nor NOR2 (N5154, N5152, N4039);
xor XOR2 (N5155, N5135, N3168);
or OR4 (N5156, N5121, N1609, N1572, N4018);
buf BUF1 (N5157, N5150);
not NOT1 (N5158, N5154);
xor XOR2 (N5159, N5155, N4267);
xor XOR2 (N5160, N5137, N841);
not NOT1 (N5161, N5159);
nor NOR2 (N5162, N5147, N1816);
nor NOR4 (N5163, N5153, N1827, N1892, N4104);
xor XOR2 (N5164, N5160, N5);
or OR2 (N5165, N5156, N2060);
and AND4 (N5166, N5165, N5062, N1697, N515);
or OR2 (N5167, N5148, N894);
and AND4 (N5168, N5166, N4784, N600, N1021);
or OR3 (N5169, N5158, N3053, N1359);
xor XOR2 (N5170, N5162, N460);
xor XOR2 (N5171, N5157, N681);
not NOT1 (N5172, N5163);
not NOT1 (N5173, N5169);
buf BUF1 (N5174, N5161);
nand NAND2 (N5175, N5171, N4555);
buf BUF1 (N5176, N5164);
or OR2 (N5177, N5175, N1580);
not NOT1 (N5178, N5170);
or OR4 (N5179, N5168, N2759, N1724, N41);
or OR3 (N5180, N5172, N3529, N1963);
xor XOR2 (N5181, N5167, N3345);
buf BUF1 (N5182, N5178);
not NOT1 (N5183, N5143);
nand NAND4 (N5184, N5182, N4702, N1189, N4527);
and AND4 (N5185, N5184, N1870, N2094, N571);
not NOT1 (N5186, N5180);
or OR2 (N5187, N5185, N2413);
or OR3 (N5188, N5177, N3940, N2605);
and AND4 (N5189, N5183, N3205, N4278, N2355);
xor XOR2 (N5190, N5189, N3715);
nand NAND4 (N5191, N5144, N967, N4574, N3316);
xor XOR2 (N5192, N5181, N4952);
xor XOR2 (N5193, N5176, N2814);
or OR4 (N5194, N5173, N1348, N3251, N3989);
or OR3 (N5195, N5193, N3708, N4870);
nand NAND2 (N5196, N5192, N1351);
nor NOR2 (N5197, N5191, N537);
or OR4 (N5198, N5194, N3267, N2532, N673);
and AND4 (N5199, N5174, N3073, N4143, N2823);
or OR2 (N5200, N5179, N4759);
not NOT1 (N5201, N5198);
xor XOR2 (N5202, N5186, N2652);
buf BUF1 (N5203, N5199);
buf BUF1 (N5204, N5196);
nor NOR2 (N5205, N5200, N1203);
buf BUF1 (N5206, N5190);
xor XOR2 (N5207, N5195, N2039);
nand NAND2 (N5208, N5202, N1172);
xor XOR2 (N5209, N5207, N3294);
or OR3 (N5210, N5188, N3384, N40);
nand NAND3 (N5211, N5201, N1084, N4639);
or OR3 (N5212, N5187, N2701, N2474);
buf BUF1 (N5213, N5212);
buf BUF1 (N5214, N5211);
not NOT1 (N5215, N5209);
not NOT1 (N5216, N5208);
and AND2 (N5217, N5206, N1348);
xor XOR2 (N5218, N5216, N2659);
xor XOR2 (N5219, N5203, N3390);
and AND2 (N5220, N5214, N289);
and AND3 (N5221, N5220, N1046, N5165);
buf BUF1 (N5222, N5205);
and AND3 (N5223, N5219, N1098, N2476);
nor NOR2 (N5224, N5218, N4865);
not NOT1 (N5225, N5204);
nand NAND3 (N5226, N5221, N582, N3326);
not NOT1 (N5227, N5224);
xor XOR2 (N5228, N5217, N4936);
or OR3 (N5229, N5210, N1955, N4095);
not NOT1 (N5230, N5213);
nand NAND2 (N5231, N5227, N265);
or OR3 (N5232, N5223, N2357, N1954);
nand NAND4 (N5233, N5215, N4958, N4989, N2586);
not NOT1 (N5234, N5233);
xor XOR2 (N5235, N5231, N4288);
nor NOR3 (N5236, N5197, N1075, N382);
nor NOR4 (N5237, N5225, N912, N5055, N1491);
or OR2 (N5238, N5222, N3591);
xor XOR2 (N5239, N5232, N768);
and AND2 (N5240, N5228, N4408);
not NOT1 (N5241, N5230);
buf BUF1 (N5242, N5241);
and AND2 (N5243, N5239, N3560);
nor NOR2 (N5244, N5240, N2890);
or OR4 (N5245, N5237, N721, N3221, N4460);
nand NAND3 (N5246, N5226, N1194, N33);
nor NOR2 (N5247, N5229, N3669);
nand NAND3 (N5248, N5238, N691, N622);
xor XOR2 (N5249, N5234, N3210);
nor NOR4 (N5250, N5242, N986, N5068, N1302);
and AND3 (N5251, N5245, N4594, N2902);
buf BUF1 (N5252, N5243);
buf BUF1 (N5253, N5248);
nand NAND2 (N5254, N5246, N4373);
xor XOR2 (N5255, N5254, N2198);
not NOT1 (N5256, N5236);
nor NOR4 (N5257, N5255, N3564, N2025, N1437);
nor NOR2 (N5258, N5253, N268);
not NOT1 (N5259, N5257);
or OR3 (N5260, N5249, N492, N1253);
nand NAND2 (N5261, N5252, N417);
not NOT1 (N5262, N5258);
nor NOR3 (N5263, N5262, N3142, N3874);
nand NAND4 (N5264, N5250, N1499, N4276, N4173);
xor XOR2 (N5265, N5235, N1265);
not NOT1 (N5266, N5264);
not NOT1 (N5267, N5265);
nor NOR4 (N5268, N5263, N3754, N4948, N1803);
and AND3 (N5269, N5251, N2267, N2308);
or OR4 (N5270, N5244, N739, N246, N1378);
and AND4 (N5271, N5266, N2494, N5041, N922);
not NOT1 (N5272, N5260);
xor XOR2 (N5273, N5271, N1515);
or OR4 (N5274, N5272, N4446, N862, N2081);
xor XOR2 (N5275, N5261, N3213);
nor NOR3 (N5276, N5267, N1449, N1299);
and AND4 (N5277, N5268, N5216, N4355, N5067);
or OR4 (N5278, N5247, N4851, N3349, N4857);
or OR2 (N5279, N5275, N1458);
or OR3 (N5280, N5279, N3416, N1007);
xor XOR2 (N5281, N5256, N3426);
xor XOR2 (N5282, N5277, N192);
xor XOR2 (N5283, N5280, N1478);
and AND4 (N5284, N5273, N3095, N1672, N4012);
buf BUF1 (N5285, N5270);
not NOT1 (N5286, N5274);
nand NAND4 (N5287, N5278, N5031, N617, N4666);
xor XOR2 (N5288, N5286, N4973);
xor XOR2 (N5289, N5281, N511);
and AND3 (N5290, N5276, N4797, N546);
nand NAND2 (N5291, N5284, N1999);
nor NOR2 (N5292, N5259, N184);
or OR3 (N5293, N5282, N3158, N4354);
xor XOR2 (N5294, N5283, N1809);
and AND2 (N5295, N5292, N1932);
nor NOR3 (N5296, N5287, N4132, N3684);
buf BUF1 (N5297, N5296);
and AND4 (N5298, N5291, N3783, N4085, N614);
not NOT1 (N5299, N5298);
xor XOR2 (N5300, N5299, N2678);
nor NOR3 (N5301, N5288, N4468, N3106);
or OR3 (N5302, N5290, N1910, N1708);
or OR2 (N5303, N5285, N3429);
xor XOR2 (N5304, N5303, N1858);
or OR4 (N5305, N5289, N734, N2899, N1828);
and AND3 (N5306, N5300, N2175, N4228);
and AND3 (N5307, N5297, N233, N3075);
and AND2 (N5308, N5269, N3469);
xor XOR2 (N5309, N5301, N3795);
nor NOR2 (N5310, N5309, N1475);
nand NAND3 (N5311, N5295, N177, N3133);
or OR2 (N5312, N5307, N2642);
xor XOR2 (N5313, N5293, N2556);
and AND4 (N5314, N5311, N735, N683, N2147);
nand NAND3 (N5315, N5310, N3412, N356);
nor NOR4 (N5316, N5315, N1746, N1251, N2006);
buf BUF1 (N5317, N5312);
nand NAND2 (N5318, N5306, N4148);
buf BUF1 (N5319, N5314);
xor XOR2 (N5320, N5318, N4230);
not NOT1 (N5321, N5316);
not NOT1 (N5322, N5319);
buf BUF1 (N5323, N5321);
or OR4 (N5324, N5322, N637, N960, N39);
or OR4 (N5325, N5320, N3750, N649, N3748);
nor NOR4 (N5326, N5308, N3825, N2931, N3428);
and AND2 (N5327, N5324, N5114);
nand NAND2 (N5328, N5304, N5168);
xor XOR2 (N5329, N5323, N1175);
nand NAND3 (N5330, N5328, N4533, N4886);
and AND2 (N5331, N5329, N2631);
xor XOR2 (N5332, N5317, N4657);
nor NOR3 (N5333, N5294, N1036, N4475);
nor NOR2 (N5334, N5326, N1649);
not NOT1 (N5335, N5302);
nand NAND4 (N5336, N5305, N1415, N881, N3315);
nor NOR2 (N5337, N5332, N710);
and AND4 (N5338, N5335, N2421, N5129, N4616);
buf BUF1 (N5339, N5336);
buf BUF1 (N5340, N5339);
nor NOR4 (N5341, N5337, N2649, N1687, N2900);
not NOT1 (N5342, N5325);
nand NAND4 (N5343, N5313, N442, N4079, N5287);
not NOT1 (N5344, N5338);
and AND4 (N5345, N5333, N1459, N761, N3809);
not NOT1 (N5346, N5342);
buf BUF1 (N5347, N5346);
buf BUF1 (N5348, N5334);
or OR3 (N5349, N5344, N1104, N2934);
or OR4 (N5350, N5327, N4413, N1392, N1535);
buf BUF1 (N5351, N5331);
and AND4 (N5352, N5340, N4488, N5056, N2176);
xor XOR2 (N5353, N5352, N3089);
xor XOR2 (N5354, N5349, N3547);
buf BUF1 (N5355, N5343);
not NOT1 (N5356, N5350);
buf BUF1 (N5357, N5353);
and AND2 (N5358, N5357, N3060);
buf BUF1 (N5359, N5348);
or OR3 (N5360, N5341, N3825, N3567);
and AND2 (N5361, N5358, N880);
or OR3 (N5362, N5355, N3501, N350);
nor NOR3 (N5363, N5360, N1658, N4892);
nor NOR4 (N5364, N5351, N72, N1321, N1056);
nor NOR3 (N5365, N5330, N607, N2444);
buf BUF1 (N5366, N5347);
and AND3 (N5367, N5361, N1196, N4488);
or OR4 (N5368, N5345, N2483, N2623, N4792);
nor NOR3 (N5369, N5364, N4957, N987);
buf BUF1 (N5370, N5354);
and AND4 (N5371, N5366, N913, N209, N2539);
not NOT1 (N5372, N5368);
or OR3 (N5373, N5370, N1341, N1543);
and AND3 (N5374, N5369, N4384, N3183);
nor NOR3 (N5375, N5367, N1449, N3099);
or OR4 (N5376, N5371, N441, N3990, N2500);
not NOT1 (N5377, N5375);
not NOT1 (N5378, N5359);
or OR4 (N5379, N5372, N1616, N2235, N1561);
and AND2 (N5380, N5377, N3939);
buf BUF1 (N5381, N5379);
not NOT1 (N5382, N5376);
not NOT1 (N5383, N5365);
and AND4 (N5384, N5382, N98, N4919, N586);
nand NAND4 (N5385, N5378, N4407, N1048, N5032);
and AND2 (N5386, N5362, N3607);
xor XOR2 (N5387, N5380, N3026);
xor XOR2 (N5388, N5373, N4886);
not NOT1 (N5389, N5385);
buf BUF1 (N5390, N5388);
or OR2 (N5391, N5387, N458);
nand NAND3 (N5392, N5390, N2319, N2215);
nand NAND4 (N5393, N5381, N2807, N3729, N448);
buf BUF1 (N5394, N5374);
nor NOR2 (N5395, N5383, N1787);
nand NAND4 (N5396, N5395, N1186, N1527, N3660);
xor XOR2 (N5397, N5391, N3596);
or OR3 (N5398, N5356, N4126, N2515);
xor XOR2 (N5399, N5363, N2914);
or OR4 (N5400, N5393, N5110, N4877, N2967);
not NOT1 (N5401, N5386);
or OR3 (N5402, N5384, N2778, N1361);
xor XOR2 (N5403, N5389, N2965);
not NOT1 (N5404, N5399);
buf BUF1 (N5405, N5398);
not NOT1 (N5406, N5392);
xor XOR2 (N5407, N5403, N1862);
buf BUF1 (N5408, N5397);
nand NAND2 (N5409, N5400, N2695);
not NOT1 (N5410, N5402);
not NOT1 (N5411, N5394);
nor NOR2 (N5412, N5408, N5330);
nor NOR3 (N5413, N5404, N746, N1725);
not NOT1 (N5414, N5401);
nand NAND4 (N5415, N5405, N3606, N482, N2478);
nor NOR4 (N5416, N5414, N2249, N2732, N1295);
buf BUF1 (N5417, N5407);
buf BUF1 (N5418, N5410);
and AND4 (N5419, N5411, N28, N920, N4573);
buf BUF1 (N5420, N5396);
nor NOR4 (N5421, N5418, N3549, N4538, N4208);
nor NOR3 (N5422, N5413, N3796, N677);
nand NAND2 (N5423, N5420, N2045);
buf BUF1 (N5424, N5422);
and AND3 (N5425, N5409, N4982, N1975);
nand NAND3 (N5426, N5421, N2807, N2733);
or OR4 (N5427, N5412, N2284, N4092, N3896);
or OR4 (N5428, N5427, N779, N173, N1149);
buf BUF1 (N5429, N5416);
xor XOR2 (N5430, N5424, N2831);
not NOT1 (N5431, N5419);
xor XOR2 (N5432, N5428, N3989);
buf BUF1 (N5433, N5406);
or OR3 (N5434, N5423, N4220, N1500);
nor NOR2 (N5435, N5430, N1022);
nand NAND3 (N5436, N5434, N2125, N4787);
buf BUF1 (N5437, N5436);
buf BUF1 (N5438, N5425);
buf BUF1 (N5439, N5438);
xor XOR2 (N5440, N5437, N3798);
nand NAND3 (N5441, N5431, N287, N4441);
buf BUF1 (N5442, N5415);
not NOT1 (N5443, N5426);
and AND2 (N5444, N5441, N2309);
and AND4 (N5445, N5417, N1072, N1743, N4684);
xor XOR2 (N5446, N5440, N2982);
nor NOR4 (N5447, N5439, N171, N1019, N1445);
xor XOR2 (N5448, N5443, N3279);
not NOT1 (N5449, N5446);
or OR3 (N5450, N5449, N5176, N496);
buf BUF1 (N5451, N5429);
and AND2 (N5452, N5442, N218);
xor XOR2 (N5453, N5435, N1773);
and AND2 (N5454, N5445, N2944);
xor XOR2 (N5455, N5432, N2445);
nand NAND3 (N5456, N5455, N3401, N3004);
buf BUF1 (N5457, N5451);
or OR4 (N5458, N5456, N458, N5187, N752);
xor XOR2 (N5459, N5452, N2660);
nor NOR3 (N5460, N5459, N3946, N1581);
buf BUF1 (N5461, N5457);
nand NAND4 (N5462, N5448, N2393, N5388, N849);
and AND3 (N5463, N5454, N2170, N4527);
nor NOR2 (N5464, N5450, N4992);
and AND3 (N5465, N5458, N1728, N250);
and AND3 (N5466, N5462, N1117, N528);
buf BUF1 (N5467, N5465);
nor NOR2 (N5468, N5466, N1291);
or OR2 (N5469, N5433, N4008);
nand NAND2 (N5470, N5453, N1184);
nand NAND4 (N5471, N5463, N3989, N2372, N3512);
xor XOR2 (N5472, N5460, N1148);
xor XOR2 (N5473, N5470, N2143);
nor NOR4 (N5474, N5469, N120, N1178, N4717);
or OR2 (N5475, N5447, N2713);
or OR4 (N5476, N5468, N4467, N2123, N1730);
not NOT1 (N5477, N5472);
or OR3 (N5478, N5444, N1986, N5052);
and AND4 (N5479, N5478, N263, N2969, N5125);
not NOT1 (N5480, N5471);
xor XOR2 (N5481, N5477, N1110);
not NOT1 (N5482, N5461);
xor XOR2 (N5483, N5464, N2154);
and AND3 (N5484, N5476, N3333, N1774);
xor XOR2 (N5485, N5482, N4671);
xor XOR2 (N5486, N5484, N1653);
or OR2 (N5487, N5474, N1304);
and AND3 (N5488, N5485, N1844, N4035);
nor NOR3 (N5489, N5475, N1501, N4844);
nand NAND4 (N5490, N5486, N4501, N2969, N682);
not NOT1 (N5491, N5479);
nand NAND3 (N5492, N5490, N4211, N337);
not NOT1 (N5493, N5467);
not NOT1 (N5494, N5483);
not NOT1 (N5495, N5492);
and AND4 (N5496, N5481, N473, N2846, N5074);
xor XOR2 (N5497, N5493, N4777);
buf BUF1 (N5498, N5489);
nand NAND3 (N5499, N5497, N4094, N346);
or OR3 (N5500, N5487, N4005, N422);
xor XOR2 (N5501, N5494, N76);
buf BUF1 (N5502, N5473);
not NOT1 (N5503, N5480);
xor XOR2 (N5504, N5496, N5259);
buf BUF1 (N5505, N5502);
and AND4 (N5506, N5505, N2174, N5176, N1349);
buf BUF1 (N5507, N5491);
buf BUF1 (N5508, N5504);
not NOT1 (N5509, N5507);
xor XOR2 (N5510, N5499, N1958);
nor NOR3 (N5511, N5501, N379, N5373);
or OR3 (N5512, N5503, N614, N5158);
nand NAND3 (N5513, N5506, N240, N3216);
buf BUF1 (N5514, N5510);
and AND4 (N5515, N5500, N27, N4791, N3385);
or OR3 (N5516, N5508, N2503, N4391);
xor XOR2 (N5517, N5488, N1315);
and AND3 (N5518, N5509, N1517, N2304);
and AND4 (N5519, N5513, N2928, N5467, N4351);
buf BUF1 (N5520, N5515);
and AND2 (N5521, N5518, N4911);
not NOT1 (N5522, N5521);
nand NAND2 (N5523, N5512, N2938);
nand NAND2 (N5524, N5522, N4633);
and AND2 (N5525, N5524, N652);
xor XOR2 (N5526, N5495, N4145);
not NOT1 (N5527, N5526);
buf BUF1 (N5528, N5519);
buf BUF1 (N5529, N5525);
buf BUF1 (N5530, N5520);
buf BUF1 (N5531, N5529);
nand NAND2 (N5532, N5523, N4455);
nor NOR2 (N5533, N5511, N3911);
and AND2 (N5534, N5531, N813);
not NOT1 (N5535, N5517);
and AND3 (N5536, N5514, N1779, N4769);
nor NOR2 (N5537, N5516, N1113);
nor NOR3 (N5538, N5537, N584, N1253);
buf BUF1 (N5539, N5528);
nor NOR3 (N5540, N5534, N4815, N2858);
not NOT1 (N5541, N5538);
buf BUF1 (N5542, N5539);
or OR3 (N5543, N5542, N2048, N4768);
nand NAND3 (N5544, N5541, N2572, N3323);
or OR2 (N5545, N5527, N5202);
and AND2 (N5546, N5536, N545);
or OR2 (N5547, N5543, N84);
and AND4 (N5548, N5535, N2208, N1776, N783);
and AND3 (N5549, N5548, N3265, N2809);
or OR4 (N5550, N5532, N3234, N4083, N4090);
and AND2 (N5551, N5549, N2716);
nor NOR3 (N5552, N5540, N955, N4898);
not NOT1 (N5553, N5552);
nand NAND4 (N5554, N5550, N2904, N4309, N309);
or OR4 (N5555, N5547, N255, N2997, N3410);
nand NAND2 (N5556, N5498, N1445);
or OR3 (N5557, N5553, N2939, N2239);
nor NOR2 (N5558, N5556, N1536);
not NOT1 (N5559, N5533);
nand NAND3 (N5560, N5559, N3998, N2003);
nand NAND3 (N5561, N5545, N4912, N2597);
not NOT1 (N5562, N5554);
and AND2 (N5563, N5561, N2868);
nor NOR3 (N5564, N5558, N559, N2152);
or OR3 (N5565, N5560, N27, N811);
or OR4 (N5566, N5557, N1563, N5216, N4629);
nand NAND3 (N5567, N5566, N1239, N4322);
not NOT1 (N5568, N5551);
nor NOR3 (N5569, N5562, N885, N2547);
not NOT1 (N5570, N5544);
and AND3 (N5571, N5567, N1794, N29);
nand NAND2 (N5572, N5571, N3962);
and AND3 (N5573, N5563, N4726, N3507);
buf BUF1 (N5574, N5564);
nor NOR3 (N5575, N5568, N3243, N1136);
and AND3 (N5576, N5570, N5382, N1921);
or OR2 (N5577, N5569, N2593);
not NOT1 (N5578, N5573);
nor NOR3 (N5579, N5578, N5223, N4342);
xor XOR2 (N5580, N5574, N3840);
nor NOR3 (N5581, N5565, N1324, N4441);
nand NAND4 (N5582, N5575, N1226, N3602, N217);
nand NAND3 (N5583, N5581, N636, N4610);
nand NAND2 (N5584, N5572, N3536);
nand NAND2 (N5585, N5530, N4075);
buf BUF1 (N5586, N5579);
not NOT1 (N5587, N5577);
and AND2 (N5588, N5586, N639);
and AND2 (N5589, N5582, N4086);
or OR2 (N5590, N5546, N1447);
xor XOR2 (N5591, N5555, N4237);
and AND4 (N5592, N5587, N1028, N2587, N4119);
nand NAND2 (N5593, N5588, N4376);
and AND2 (N5594, N5589, N523);
xor XOR2 (N5595, N5576, N1994);
buf BUF1 (N5596, N5583);
buf BUF1 (N5597, N5595);
xor XOR2 (N5598, N5596, N3731);
buf BUF1 (N5599, N5593);
nor NOR3 (N5600, N5580, N3967, N3159);
xor XOR2 (N5601, N5598, N2819);
buf BUF1 (N5602, N5585);
and AND2 (N5603, N5597, N44);
not NOT1 (N5604, N5600);
and AND3 (N5605, N5601, N5292, N519);
or OR3 (N5606, N5584, N3894, N2855);
buf BUF1 (N5607, N5599);
or OR4 (N5608, N5603, N5191, N3618, N4982);
nand NAND4 (N5609, N5608, N4995, N1410, N3280);
nand NAND4 (N5610, N5590, N720, N3438, N97);
or OR2 (N5611, N5592, N2055);
not NOT1 (N5612, N5610);
nor NOR2 (N5613, N5611, N4336);
not NOT1 (N5614, N5609);
buf BUF1 (N5615, N5594);
or OR4 (N5616, N5614, N2970, N3947, N2031);
and AND4 (N5617, N5607, N5287, N524, N76);
nor NOR4 (N5618, N5604, N353, N4233, N5484);
not NOT1 (N5619, N5612);
not NOT1 (N5620, N5605);
or OR3 (N5621, N5615, N3660, N1241);
and AND4 (N5622, N5621, N2365, N5075, N909);
and AND4 (N5623, N5619, N779, N171, N2948);
nor NOR4 (N5624, N5618, N5516, N455, N1582);
buf BUF1 (N5625, N5602);
nor NOR3 (N5626, N5624, N4659, N3803);
nor NOR4 (N5627, N5606, N5178, N2491, N1548);
and AND4 (N5628, N5626, N5542, N2749, N891);
buf BUF1 (N5629, N5628);
buf BUF1 (N5630, N5591);
or OR4 (N5631, N5613, N5575, N5116, N4578);
buf BUF1 (N5632, N5623);
nor NOR2 (N5633, N5631, N5182);
or OR2 (N5634, N5627, N904);
and AND3 (N5635, N5616, N4321, N3368);
or OR4 (N5636, N5622, N1320, N4343, N1830);
nor NOR4 (N5637, N5625, N1662, N2117, N3073);
or OR3 (N5638, N5635, N178, N3272);
not NOT1 (N5639, N5629);
nor NOR4 (N5640, N5617, N613, N1786, N3630);
xor XOR2 (N5641, N5632, N1919);
buf BUF1 (N5642, N5630);
nand NAND2 (N5643, N5636, N3318);
and AND3 (N5644, N5637, N3163, N4208);
nand NAND4 (N5645, N5639, N4872, N1832, N5528);
nand NAND2 (N5646, N5640, N846);
and AND2 (N5647, N5634, N3242);
not NOT1 (N5648, N5641);
buf BUF1 (N5649, N5647);
xor XOR2 (N5650, N5648, N5165);
nand NAND2 (N5651, N5643, N3890);
and AND2 (N5652, N5646, N1152);
nand NAND2 (N5653, N5620, N1347);
not NOT1 (N5654, N5653);
nor NOR3 (N5655, N5650, N5398, N5247);
or OR3 (N5656, N5652, N3668, N4888);
buf BUF1 (N5657, N5654);
nand NAND2 (N5658, N5642, N1066);
nor NOR3 (N5659, N5656, N2862, N2013);
not NOT1 (N5660, N5655);
nor NOR4 (N5661, N5633, N54, N4542, N2004);
and AND4 (N5662, N5658, N1580, N777, N4316);
nor NOR2 (N5663, N5638, N2704);
and AND3 (N5664, N5645, N537, N1151);
or OR4 (N5665, N5651, N4613, N5594, N288);
not NOT1 (N5666, N5662);
buf BUF1 (N5667, N5665);
xor XOR2 (N5668, N5667, N1133);
or OR2 (N5669, N5649, N3479);
and AND4 (N5670, N5666, N5414, N3626, N2005);
and AND2 (N5671, N5644, N3103);
and AND2 (N5672, N5661, N4578);
xor XOR2 (N5673, N5669, N4865);
buf BUF1 (N5674, N5663);
not NOT1 (N5675, N5674);
buf BUF1 (N5676, N5657);
buf BUF1 (N5677, N5670);
buf BUF1 (N5678, N5671);
nor NOR3 (N5679, N5675, N2869, N2730);
nand NAND4 (N5680, N5678, N4833, N4860, N5382);
and AND2 (N5681, N5680, N4720);
xor XOR2 (N5682, N5681, N4361);
buf BUF1 (N5683, N5676);
nand NAND2 (N5684, N5668, N1754);
nand NAND4 (N5685, N5683, N4989, N3416, N1145);
not NOT1 (N5686, N5682);
and AND2 (N5687, N5685, N4358);
and AND4 (N5688, N5684, N5113, N2926, N135);
and AND4 (N5689, N5688, N1952, N2816, N1179);
buf BUF1 (N5690, N5687);
not NOT1 (N5691, N5664);
buf BUF1 (N5692, N5691);
nand NAND3 (N5693, N5677, N4471, N5623);
and AND4 (N5694, N5693, N364, N17, N1983);
buf BUF1 (N5695, N5659);
buf BUF1 (N5696, N5679);
nor NOR3 (N5697, N5694, N4371, N1744);
nand NAND2 (N5698, N5673, N4438);
not NOT1 (N5699, N5686);
or OR2 (N5700, N5692, N432);
xor XOR2 (N5701, N5700, N742);
xor XOR2 (N5702, N5660, N3625);
not NOT1 (N5703, N5689);
nand NAND2 (N5704, N5701, N82);
xor XOR2 (N5705, N5704, N1155);
nand NAND4 (N5706, N5696, N4082, N4991, N4841);
xor XOR2 (N5707, N5695, N1355);
and AND2 (N5708, N5702, N4410);
not NOT1 (N5709, N5706);
and AND3 (N5710, N5697, N1513, N1824);
nor NOR4 (N5711, N5705, N5480, N756, N1841);
nor NOR3 (N5712, N5709, N404, N225);
buf BUF1 (N5713, N5703);
nor NOR4 (N5714, N5712, N1498, N139, N5301);
buf BUF1 (N5715, N5708);
nor NOR3 (N5716, N5699, N1318, N247);
and AND3 (N5717, N5710, N3068, N4445);
buf BUF1 (N5718, N5672);
not NOT1 (N5719, N5711);
nor NOR4 (N5720, N5714, N519, N4793, N5380);
nand NAND4 (N5721, N5698, N2322, N1997, N203);
and AND4 (N5722, N5716, N1690, N2469, N4112);
and AND3 (N5723, N5713, N3931, N1634);
nor NOR4 (N5724, N5718, N811, N4560, N2407);
not NOT1 (N5725, N5690);
or OR3 (N5726, N5725, N4613, N4044);
or OR2 (N5727, N5717, N148);
not NOT1 (N5728, N5721);
nand NAND4 (N5729, N5719, N1556, N4194, N4337);
buf BUF1 (N5730, N5724);
nor NOR2 (N5731, N5723, N1479);
not NOT1 (N5732, N5726);
or OR2 (N5733, N5728, N2777);
or OR3 (N5734, N5730, N4335, N4045);
xor XOR2 (N5735, N5715, N5504);
xor XOR2 (N5736, N5727, N119);
or OR3 (N5737, N5732, N2856, N368);
or OR2 (N5738, N5733, N1052);
nand NAND4 (N5739, N5722, N3924, N974, N2602);
nand NAND4 (N5740, N5720, N3140, N4587, N3812);
buf BUF1 (N5741, N5734);
or OR4 (N5742, N5736, N5137, N1228, N3381);
buf BUF1 (N5743, N5729);
not NOT1 (N5744, N5735);
or OR2 (N5745, N5707, N4891);
nor NOR3 (N5746, N5731, N188, N213);
nor NOR3 (N5747, N5740, N4957, N293);
buf BUF1 (N5748, N5739);
or OR4 (N5749, N5744, N2809, N3757, N4888);
nor NOR2 (N5750, N5738, N1527);
nand NAND2 (N5751, N5741, N4729);
buf BUF1 (N5752, N5750);
nor NOR3 (N5753, N5743, N1309, N2786);
xor XOR2 (N5754, N5747, N1375);
nor NOR2 (N5755, N5752, N1954);
nor NOR3 (N5756, N5753, N2764, N5063);
nor NOR2 (N5757, N5749, N792);
not NOT1 (N5758, N5748);
not NOT1 (N5759, N5737);
nand NAND2 (N5760, N5745, N2857);
xor XOR2 (N5761, N5742, N1650);
nand NAND2 (N5762, N5760, N3588);
xor XOR2 (N5763, N5762, N4973);
xor XOR2 (N5764, N5754, N2486);
and AND2 (N5765, N5761, N3142);
or OR3 (N5766, N5755, N3735, N2937);
nand NAND3 (N5767, N5758, N2360, N5668);
not NOT1 (N5768, N5756);
or OR4 (N5769, N5768, N1551, N2421, N1490);
buf BUF1 (N5770, N5751);
and AND3 (N5771, N5764, N988, N84);
xor XOR2 (N5772, N5771, N1479);
xor XOR2 (N5773, N5769, N344);
or OR3 (N5774, N5773, N5699, N206);
or OR3 (N5775, N5767, N2325, N1929);
nand NAND4 (N5776, N5765, N2421, N5608, N4815);
xor XOR2 (N5777, N5757, N4457);
buf BUF1 (N5778, N5763);
buf BUF1 (N5779, N5776);
nor NOR2 (N5780, N5746, N4285);
nor NOR3 (N5781, N5780, N4618, N2235);
or OR2 (N5782, N5777, N5454);
or OR4 (N5783, N5778, N3543, N987, N3335);
nor NOR4 (N5784, N5759, N1305, N4553, N4108);
nand NAND3 (N5785, N5781, N2039, N5242);
and AND3 (N5786, N5782, N4109, N1410);
not NOT1 (N5787, N5786);
and AND3 (N5788, N5779, N3954, N1835);
nor NOR2 (N5789, N5775, N5176);
nand NAND4 (N5790, N5772, N1308, N3876, N3442);
xor XOR2 (N5791, N5770, N5053);
buf BUF1 (N5792, N5774);
not NOT1 (N5793, N5766);
buf BUF1 (N5794, N5784);
or OR4 (N5795, N5793, N377, N2707, N862);
nand NAND3 (N5796, N5788, N5585, N710);
xor XOR2 (N5797, N5792, N3178);
buf BUF1 (N5798, N5789);
xor XOR2 (N5799, N5790, N3810);
not NOT1 (N5800, N5799);
buf BUF1 (N5801, N5785);
nand NAND4 (N5802, N5801, N3142, N1014, N5457);
nand NAND2 (N5803, N5796, N5748);
or OR3 (N5804, N5795, N297, N1893);
buf BUF1 (N5805, N5800);
and AND4 (N5806, N5794, N5484, N1462, N2937);
not NOT1 (N5807, N5806);
xor XOR2 (N5808, N5802, N4319);
not NOT1 (N5809, N5783);
not NOT1 (N5810, N5805);
xor XOR2 (N5811, N5798, N4805);
or OR3 (N5812, N5791, N2647, N1790);
or OR3 (N5813, N5804, N1634, N5425);
not NOT1 (N5814, N5809);
nor NOR2 (N5815, N5787, N197);
or OR2 (N5816, N5797, N2223);
or OR2 (N5817, N5810, N5076);
and AND4 (N5818, N5807, N5406, N674, N3733);
xor XOR2 (N5819, N5811, N4861);
or OR3 (N5820, N5808, N3118, N5291);
or OR2 (N5821, N5818, N1764);
not NOT1 (N5822, N5813);
buf BUF1 (N5823, N5817);
and AND3 (N5824, N5819, N2439, N1847);
and AND2 (N5825, N5823, N2430);
buf BUF1 (N5826, N5822);
or OR3 (N5827, N5825, N5698, N746);
buf BUF1 (N5828, N5812);
nor NOR4 (N5829, N5803, N3676, N5503, N3551);
nor NOR3 (N5830, N5816, N3723, N4283);
xor XOR2 (N5831, N5828, N4539);
not NOT1 (N5832, N5815);
or OR4 (N5833, N5821, N3812, N4249, N4513);
or OR2 (N5834, N5829, N1748);
and AND2 (N5835, N5834, N2533);
buf BUF1 (N5836, N5831);
not NOT1 (N5837, N5833);
or OR2 (N5838, N5824, N1880);
or OR4 (N5839, N5820, N2079, N5691, N2515);
or OR4 (N5840, N5814, N2575, N3131, N1355);
not NOT1 (N5841, N5837);
xor XOR2 (N5842, N5838, N3352);
nand NAND2 (N5843, N5836, N1445);
nor NOR4 (N5844, N5840, N1521, N1288, N1377);
and AND2 (N5845, N5841, N5324);
buf BUF1 (N5846, N5826);
nand NAND2 (N5847, N5839, N1019);
buf BUF1 (N5848, N5843);
nand NAND4 (N5849, N5848, N3106, N2333, N3231);
not NOT1 (N5850, N5846);
buf BUF1 (N5851, N5827);
not NOT1 (N5852, N5850);
not NOT1 (N5853, N5851);
or OR2 (N5854, N5835, N4599);
buf BUF1 (N5855, N5845);
buf BUF1 (N5856, N5844);
not NOT1 (N5857, N5853);
buf BUF1 (N5858, N5832);
or OR3 (N5859, N5847, N4559, N2643);
xor XOR2 (N5860, N5854, N3433);
and AND2 (N5861, N5856, N259);
and AND4 (N5862, N5842, N540, N529, N3141);
and AND3 (N5863, N5857, N4375, N3136);
xor XOR2 (N5864, N5855, N5582);
nor NOR4 (N5865, N5864, N125, N2105, N3919);
or OR3 (N5866, N5859, N3563, N630);
buf BUF1 (N5867, N5862);
nand NAND4 (N5868, N5860, N432, N2702, N627);
and AND2 (N5869, N5830, N548);
or OR2 (N5870, N5866, N3161);
nand NAND3 (N5871, N5852, N4007, N2630);
xor XOR2 (N5872, N5858, N4131);
nand NAND4 (N5873, N5849, N5829, N2504, N1615);
not NOT1 (N5874, N5865);
xor XOR2 (N5875, N5863, N4579);
nand NAND3 (N5876, N5873, N3180, N1873);
nor NOR2 (N5877, N5867, N631);
buf BUF1 (N5878, N5877);
nand NAND4 (N5879, N5871, N741, N1433, N452);
or OR2 (N5880, N5868, N3903);
or OR2 (N5881, N5872, N1811);
xor XOR2 (N5882, N5880, N1148);
and AND2 (N5883, N5878, N2201);
or OR4 (N5884, N5861, N4433, N1182, N95);
and AND2 (N5885, N5884, N3483);
not NOT1 (N5886, N5883);
nor NOR3 (N5887, N5881, N2568, N3348);
xor XOR2 (N5888, N5887, N4154);
xor XOR2 (N5889, N5876, N285);
buf BUF1 (N5890, N5870);
not NOT1 (N5891, N5889);
nor NOR3 (N5892, N5891, N1590, N1758);
xor XOR2 (N5893, N5875, N4220);
not NOT1 (N5894, N5882);
xor XOR2 (N5895, N5886, N4657);
buf BUF1 (N5896, N5890);
and AND2 (N5897, N5888, N3431);
and AND2 (N5898, N5885, N4699);
xor XOR2 (N5899, N5879, N2608);
xor XOR2 (N5900, N5892, N1661);
not NOT1 (N5901, N5894);
buf BUF1 (N5902, N5900);
nor NOR2 (N5903, N5869, N3931);
not NOT1 (N5904, N5895);
xor XOR2 (N5905, N5898, N4276);
xor XOR2 (N5906, N5899, N3834);
not NOT1 (N5907, N5901);
nand NAND3 (N5908, N5905, N2118, N4907);
nand NAND3 (N5909, N5897, N1055, N1531);
buf BUF1 (N5910, N5874);
xor XOR2 (N5911, N5903, N1276);
nor NOR2 (N5912, N5908, N4259);
xor XOR2 (N5913, N5909, N1683);
and AND4 (N5914, N5912, N3520, N4476, N5467);
or OR4 (N5915, N5904, N2917, N5531, N570);
nand NAND2 (N5916, N5914, N5372);
nand NAND3 (N5917, N5916, N785, N846);
nand NAND2 (N5918, N5907, N3288);
nor NOR4 (N5919, N5913, N1916, N5486, N2469);
xor XOR2 (N5920, N5910, N5734);
and AND3 (N5921, N5917, N5484, N172);
buf BUF1 (N5922, N5915);
and AND2 (N5923, N5922, N5395);
or OR3 (N5924, N5893, N1721, N4526);
and AND3 (N5925, N5919, N3564, N3404);
not NOT1 (N5926, N5920);
nand NAND2 (N5927, N5923, N3070);
or OR3 (N5928, N5927, N4849, N4131);
not NOT1 (N5929, N5896);
xor XOR2 (N5930, N5906, N5630);
nand NAND4 (N5931, N5902, N938, N4457, N5004);
nand NAND3 (N5932, N5930, N5605, N3364);
nand NAND4 (N5933, N5931, N1802, N2090, N3873);
nor NOR3 (N5934, N5929, N2217, N870);
or OR4 (N5935, N5911, N4669, N935, N3987);
and AND4 (N5936, N5918, N3149, N2039, N4731);
or OR2 (N5937, N5926, N5318);
nor NOR3 (N5938, N5932, N3359, N5804);
xor XOR2 (N5939, N5935, N4839);
xor XOR2 (N5940, N5937, N4777);
xor XOR2 (N5941, N5936, N1244);
nand NAND3 (N5942, N5938, N2303, N3898);
and AND2 (N5943, N5941, N5889);
not NOT1 (N5944, N5924);
or OR2 (N5945, N5925, N4491);
buf BUF1 (N5946, N5942);
not NOT1 (N5947, N5944);
nand NAND2 (N5948, N5933, N3269);
xor XOR2 (N5949, N5921, N3044);
and AND3 (N5950, N5939, N4564, N4088);
buf BUF1 (N5951, N5928);
not NOT1 (N5952, N5943);
and AND3 (N5953, N5952, N3499, N4989);
or OR2 (N5954, N5950, N5139);
and AND3 (N5955, N5946, N4259, N5363);
not NOT1 (N5956, N5934);
xor XOR2 (N5957, N5956, N2956);
nor NOR4 (N5958, N5953, N2016, N505, N3506);
nand NAND3 (N5959, N5951, N276, N4357);
nor NOR4 (N5960, N5940, N3108, N4019, N923);
and AND4 (N5961, N5948, N44, N3556, N3724);
nand NAND4 (N5962, N5959, N3913, N3927, N2212);
nand NAND3 (N5963, N5961, N4100, N548);
and AND3 (N5964, N5960, N3651, N2327);
nand NAND2 (N5965, N5947, N1705);
not NOT1 (N5966, N5965);
xor XOR2 (N5967, N5955, N4262);
or OR2 (N5968, N5967, N4635);
buf BUF1 (N5969, N5954);
nor NOR3 (N5970, N5966, N4721, N5652);
nand NAND4 (N5971, N5949, N4060, N2760, N5805);
not NOT1 (N5972, N5962);
nor NOR2 (N5973, N5945, N3482);
not NOT1 (N5974, N5972);
nor NOR3 (N5975, N5957, N5722, N5718);
not NOT1 (N5976, N5958);
nand NAND4 (N5977, N5973, N2263, N440, N5100);
nand NAND4 (N5978, N5974, N5258, N339, N3285);
nand NAND3 (N5979, N5976, N3875, N1876);
and AND4 (N5980, N5970, N3906, N131, N5951);
nand NAND4 (N5981, N5980, N2127, N3663, N3737);
buf BUF1 (N5982, N5981);
not NOT1 (N5983, N5971);
nand NAND4 (N5984, N5963, N4151, N1715, N5865);
not NOT1 (N5985, N5983);
and AND3 (N5986, N5975, N2600, N794);
xor XOR2 (N5987, N5982, N4040);
buf BUF1 (N5988, N5968);
not NOT1 (N5989, N5964);
and AND2 (N5990, N5984, N2788);
xor XOR2 (N5991, N5989, N1460);
not NOT1 (N5992, N5977);
nor NOR4 (N5993, N5986, N4522, N363, N4417);
nand NAND3 (N5994, N5992, N2632, N471);
nor NOR3 (N5995, N5969, N5602, N3269);
buf BUF1 (N5996, N5994);
and AND3 (N5997, N5987, N2964, N1651);
or OR4 (N5998, N5985, N5648, N5096, N3356);
nor NOR4 (N5999, N5991, N858, N5871, N3651);
xor XOR2 (N6000, N5988, N410);
xor XOR2 (N6001, N5997, N4102);
xor XOR2 (N6002, N5998, N4297);
not NOT1 (N6003, N5990);
nand NAND4 (N6004, N5993, N743, N4249, N3706);
not NOT1 (N6005, N5979);
buf BUF1 (N6006, N6005);
xor XOR2 (N6007, N6004, N2483);
not NOT1 (N6008, N6002);
nor NOR2 (N6009, N5995, N5938);
nand NAND2 (N6010, N6007, N5776);
nor NOR3 (N6011, N6006, N4504, N1056);
or OR2 (N6012, N6008, N5067);
nand NAND4 (N6013, N6003, N19, N1721, N3204);
nor NOR2 (N6014, N5999, N3869);
not NOT1 (N6015, N5996);
not NOT1 (N6016, N6012);
or OR4 (N6017, N6010, N2920, N3272, N2808);
not NOT1 (N6018, N6017);
and AND2 (N6019, N6009, N4411);
nor NOR2 (N6020, N6016, N2800);
nand NAND3 (N6021, N6011, N4369, N802);
xor XOR2 (N6022, N6021, N3584);
xor XOR2 (N6023, N6018, N4808);
or OR3 (N6024, N6023, N3613, N3861);
nand NAND4 (N6025, N6020, N196, N2150, N255);
nand NAND4 (N6026, N6000, N5816, N20, N2517);
xor XOR2 (N6027, N6022, N7);
xor XOR2 (N6028, N5978, N1409);
buf BUF1 (N6029, N6024);
not NOT1 (N6030, N6028);
xor XOR2 (N6031, N6014, N44);
buf BUF1 (N6032, N6026);
or OR3 (N6033, N6030, N667, N475);
nand NAND4 (N6034, N6025, N407, N3374, N4357);
xor XOR2 (N6035, N6034, N4090);
nand NAND3 (N6036, N6019, N2874, N460);
and AND4 (N6037, N6001, N1863, N5185, N3979);
or OR3 (N6038, N6035, N4459, N5492);
nor NOR3 (N6039, N6037, N1791, N1375);
or OR3 (N6040, N6027, N4899, N3617);
and AND2 (N6041, N6040, N4947);
and AND4 (N6042, N6038, N5699, N4990, N2207);
buf BUF1 (N6043, N6041);
xor XOR2 (N6044, N6042, N3681);
not NOT1 (N6045, N6013);
xor XOR2 (N6046, N6033, N3995);
not NOT1 (N6047, N6045);
or OR3 (N6048, N6015, N329, N1155);
or OR2 (N6049, N6029, N4522);
or OR4 (N6050, N6046, N111, N2823, N877);
nand NAND3 (N6051, N6036, N4456, N668);
nor NOR2 (N6052, N6050, N660);
not NOT1 (N6053, N6049);
nor NOR4 (N6054, N6051, N2694, N1064, N5957);
buf BUF1 (N6055, N6044);
not NOT1 (N6056, N6043);
or OR3 (N6057, N6054, N2322, N5438);
buf BUF1 (N6058, N6047);
or OR4 (N6059, N6032, N4544, N1179, N1563);
not NOT1 (N6060, N6059);
xor XOR2 (N6061, N6052, N1794);
or OR4 (N6062, N6056, N1884, N3650, N5318);
buf BUF1 (N6063, N6061);
buf BUF1 (N6064, N6060);
buf BUF1 (N6065, N6055);
or OR2 (N6066, N6062, N4018);
not NOT1 (N6067, N6031);
and AND3 (N6068, N6065, N131, N3791);
nand NAND2 (N6069, N6039, N1543);
nand NAND3 (N6070, N6067, N85, N1993);
nand NAND2 (N6071, N6053, N185);
xor XOR2 (N6072, N6066, N2936);
nor NOR2 (N6073, N6063, N4706);
nand NAND4 (N6074, N6073, N6015, N1012, N1908);
not NOT1 (N6075, N6070);
nand NAND2 (N6076, N6071, N5954);
xor XOR2 (N6077, N6048, N2197);
nor NOR2 (N6078, N6077, N5116);
and AND2 (N6079, N6078, N382);
buf BUF1 (N6080, N6058);
buf BUF1 (N6081, N6076);
not NOT1 (N6082, N6079);
nand NAND2 (N6083, N6080, N120);
and AND3 (N6084, N6081, N3767, N5559);
and AND4 (N6085, N6064, N296, N3907, N124);
or OR3 (N6086, N6085, N1228, N4393);
nand NAND3 (N6087, N6069, N2429, N5316);
or OR3 (N6088, N6075, N2124, N1824);
buf BUF1 (N6089, N6068);
not NOT1 (N6090, N6086);
buf BUF1 (N6091, N6088);
and AND2 (N6092, N6089, N3133);
not NOT1 (N6093, N6083);
not NOT1 (N6094, N6084);
or OR2 (N6095, N6091, N926);
nor NOR4 (N6096, N6092, N3534, N2216, N3980);
buf BUF1 (N6097, N6087);
or OR3 (N6098, N6057, N4612, N4902);
xor XOR2 (N6099, N6074, N1938);
nor NOR2 (N6100, N6093, N3846);
buf BUF1 (N6101, N6094);
xor XOR2 (N6102, N6072, N1207);
nand NAND2 (N6103, N6097, N5570);
or OR2 (N6104, N6100, N2771);
xor XOR2 (N6105, N6103, N142);
nand NAND3 (N6106, N6098, N3692, N1809);
and AND2 (N6107, N6101, N1763);
nand NAND3 (N6108, N6106, N2614, N5332);
nor NOR4 (N6109, N6099, N651, N2336, N5260);
buf BUF1 (N6110, N6090);
nor NOR4 (N6111, N6107, N4840, N6085, N3640);
or OR2 (N6112, N6082, N5869);
xor XOR2 (N6113, N6108, N1806);
not NOT1 (N6114, N6111);
and AND4 (N6115, N6105, N3824, N3997, N203);
not NOT1 (N6116, N6104);
buf BUF1 (N6117, N6112);
or OR4 (N6118, N6110, N351, N437, N754);
not NOT1 (N6119, N6117);
or OR2 (N6120, N6102, N2484);
nand NAND4 (N6121, N6095, N3172, N3835, N3350);
or OR3 (N6122, N6121, N3648, N917);
nor NOR2 (N6123, N6119, N3051);
buf BUF1 (N6124, N6122);
buf BUF1 (N6125, N6116);
nor NOR3 (N6126, N6114, N1583, N4252);
or OR3 (N6127, N6124, N1775, N4264);
xor XOR2 (N6128, N6113, N394);
buf BUF1 (N6129, N6128);
or OR3 (N6130, N6126, N3325, N4580);
or OR3 (N6131, N6096, N1697, N4663);
xor XOR2 (N6132, N6115, N890);
not NOT1 (N6133, N6125);
or OR2 (N6134, N6131, N4154);
and AND2 (N6135, N6127, N5337);
xor XOR2 (N6136, N6135, N5544);
not NOT1 (N6137, N6118);
not NOT1 (N6138, N6123);
nand NAND2 (N6139, N6132, N2225);
buf BUF1 (N6140, N6139);
not NOT1 (N6141, N6137);
and AND4 (N6142, N6109, N3453, N413, N2322);
and AND2 (N6143, N6138, N1357);
nor NOR2 (N6144, N6142, N1867);
and AND3 (N6145, N6130, N4485, N784);
not NOT1 (N6146, N6133);
xor XOR2 (N6147, N6145, N1109);
nor NOR4 (N6148, N6129, N2466, N411, N2066);
and AND2 (N6149, N6147, N1241);
buf BUF1 (N6150, N6149);
not NOT1 (N6151, N6140);
nor NOR4 (N6152, N6141, N6010, N1277, N4438);
not NOT1 (N6153, N6136);
buf BUF1 (N6154, N6143);
xor XOR2 (N6155, N6144, N3210);
nor NOR4 (N6156, N6146, N3727, N279, N4594);
buf BUF1 (N6157, N6155);
xor XOR2 (N6158, N6120, N3721);
or OR3 (N6159, N6151, N1806, N326);
nand NAND4 (N6160, N6134, N5742, N1919, N1794);
not NOT1 (N6161, N6156);
buf BUF1 (N6162, N6159);
or OR3 (N6163, N6150, N2283, N479);
nor NOR2 (N6164, N6148, N3626);
nand NAND2 (N6165, N6160, N5732);
xor XOR2 (N6166, N6157, N546);
nor NOR3 (N6167, N6158, N4952, N3014);
nor NOR3 (N6168, N6154, N513, N2816);
buf BUF1 (N6169, N6166);
buf BUF1 (N6170, N6162);
nor NOR4 (N6171, N6161, N3071, N3061, N4333);
nand NAND3 (N6172, N6164, N3451, N5890);
nor NOR3 (N6173, N6172, N5713, N4936);
and AND4 (N6174, N6165, N1397, N5352, N214);
not NOT1 (N6175, N6153);
or OR4 (N6176, N6173, N1970, N4699, N4625);
and AND2 (N6177, N6167, N4524);
buf BUF1 (N6178, N6171);
buf BUF1 (N6179, N6169);
nand NAND3 (N6180, N6152, N5639, N5622);
nor NOR4 (N6181, N6180, N3389, N3288, N196);
nand NAND4 (N6182, N6181, N3484, N5616, N2581);
buf BUF1 (N6183, N6175);
nand NAND4 (N6184, N6163, N5391, N3191, N5170);
nand NAND4 (N6185, N6176, N1432, N4047, N4481);
or OR2 (N6186, N6182, N4196);
and AND4 (N6187, N6178, N3384, N757, N2176);
not NOT1 (N6188, N6177);
or OR2 (N6189, N6187, N891);
buf BUF1 (N6190, N6185);
not NOT1 (N6191, N6179);
not NOT1 (N6192, N6170);
xor XOR2 (N6193, N6188, N3617);
nor NOR2 (N6194, N6174, N45);
or OR4 (N6195, N6184, N1484, N4439, N5329);
or OR2 (N6196, N6183, N1199);
buf BUF1 (N6197, N6194);
buf BUF1 (N6198, N6168);
nand NAND2 (N6199, N6192, N5615);
xor XOR2 (N6200, N6195, N1121);
nor NOR3 (N6201, N6186, N4795, N612);
nand NAND4 (N6202, N6193, N112, N3486, N4898);
xor XOR2 (N6203, N6191, N4986);
nor NOR2 (N6204, N6198, N2275);
nand NAND2 (N6205, N6189, N3279);
and AND4 (N6206, N6204, N1917, N3653, N2999);
or OR2 (N6207, N6190, N3435);
buf BUF1 (N6208, N6205);
nor NOR4 (N6209, N6207, N4744, N3713, N5889);
buf BUF1 (N6210, N6197);
and AND2 (N6211, N6200, N5061);
xor XOR2 (N6212, N6199, N2040);
nand NAND2 (N6213, N6196, N715);
xor XOR2 (N6214, N6203, N5626);
buf BUF1 (N6215, N6214);
not NOT1 (N6216, N6215);
or OR2 (N6217, N6206, N1363);
and AND3 (N6218, N6217, N182, N5246);
nor NOR2 (N6219, N6216, N3408);
buf BUF1 (N6220, N6202);
nor NOR4 (N6221, N6220, N86, N195, N2048);
and AND2 (N6222, N6208, N1567);
and AND3 (N6223, N6221, N4947, N1564);
nand NAND4 (N6224, N6222, N5804, N3137, N2706);
xor XOR2 (N6225, N6210, N5569);
nor NOR3 (N6226, N6211, N3751, N5489);
or OR3 (N6227, N6225, N2328, N3321);
or OR3 (N6228, N6227, N3247, N6086);
buf BUF1 (N6229, N6223);
not NOT1 (N6230, N6228);
nand NAND4 (N6231, N6230, N5676, N3860, N4002);
or OR2 (N6232, N6229, N5159);
not NOT1 (N6233, N6212);
and AND4 (N6234, N6218, N2472, N3743, N3389);
or OR4 (N6235, N6231, N1747, N1360, N6030);
and AND2 (N6236, N6201, N4501);
nand NAND3 (N6237, N6236, N176, N818);
nor NOR2 (N6238, N6235, N5621);
buf BUF1 (N6239, N6224);
and AND2 (N6240, N6234, N3647);
buf BUF1 (N6241, N6213);
buf BUF1 (N6242, N6233);
xor XOR2 (N6243, N6219, N46);
xor XOR2 (N6244, N6242, N6007);
nor NOR2 (N6245, N6239, N2273);
nand NAND2 (N6246, N6226, N1030);
nand NAND2 (N6247, N6246, N3707);
nand NAND2 (N6248, N6241, N5492);
nand NAND3 (N6249, N6232, N4092, N1292);
or OR2 (N6250, N6248, N5387);
not NOT1 (N6251, N6247);
nand NAND3 (N6252, N6238, N380, N2980);
or OR3 (N6253, N6251, N126, N3594);
or OR3 (N6254, N6209, N3155, N3733);
buf BUF1 (N6255, N6244);
nor NOR4 (N6256, N6243, N1885, N4981, N3647);
or OR3 (N6257, N6245, N673, N4218);
xor XOR2 (N6258, N6249, N3443);
buf BUF1 (N6259, N6257);
buf BUF1 (N6260, N6253);
or OR3 (N6261, N6240, N145, N5551);
xor XOR2 (N6262, N6259, N130);
or OR4 (N6263, N6258, N2806, N4896, N5184);
and AND3 (N6264, N6250, N100, N1334);
or OR4 (N6265, N6255, N1143, N853, N3728);
nand NAND4 (N6266, N6263, N3020, N5081, N2304);
or OR4 (N6267, N6265, N4571, N1220, N2182);
and AND4 (N6268, N6260, N3648, N2347, N5083);
nor NOR2 (N6269, N6261, N3672);
or OR2 (N6270, N6254, N4991);
nor NOR3 (N6271, N6268, N4188, N6053);
not NOT1 (N6272, N6262);
nand NAND4 (N6273, N6252, N5673, N4157, N2025);
and AND3 (N6274, N6273, N5093, N1510);
and AND3 (N6275, N6270, N884, N2865);
xor XOR2 (N6276, N6256, N4639);
xor XOR2 (N6277, N6237, N5339);
xor XOR2 (N6278, N6264, N5932);
nand NAND4 (N6279, N6277, N4706, N3232, N2034);
buf BUF1 (N6280, N6272);
xor XOR2 (N6281, N6266, N4028);
and AND2 (N6282, N6274, N3123);
xor XOR2 (N6283, N6281, N3671);
or OR2 (N6284, N6271, N737);
nand NAND4 (N6285, N6267, N820, N4686, N1263);
nor NOR4 (N6286, N6269, N4998, N1850, N6137);
not NOT1 (N6287, N6280);
xor XOR2 (N6288, N6285, N780);
or OR4 (N6289, N6283, N2312, N2169, N1759);
not NOT1 (N6290, N6282);
not NOT1 (N6291, N6288);
or OR3 (N6292, N6284, N2286, N1807);
xor XOR2 (N6293, N6290, N2522);
nor NOR2 (N6294, N6279, N1099);
and AND4 (N6295, N6293, N414, N3034, N3288);
nor NOR3 (N6296, N6287, N4351, N2307);
and AND4 (N6297, N6276, N1508, N1070, N2772);
buf BUF1 (N6298, N6289);
nor NOR3 (N6299, N6292, N4448, N837);
and AND2 (N6300, N6296, N2460);
or OR4 (N6301, N6295, N6156, N237, N3361);
nand NAND4 (N6302, N6301, N1777, N407, N79);
not NOT1 (N6303, N6286);
or OR2 (N6304, N6302, N3556);
or OR2 (N6305, N6303, N571);
not NOT1 (N6306, N6298);
not NOT1 (N6307, N6305);
or OR4 (N6308, N6304, N4064, N1540, N2933);
or OR2 (N6309, N6299, N1624);
nor NOR4 (N6310, N6306, N2976, N4718, N2890);
xor XOR2 (N6311, N6307, N1550);
nand NAND2 (N6312, N6310, N1055);
nand NAND3 (N6313, N6278, N573, N2066);
nor NOR3 (N6314, N6312, N1845, N307);
xor XOR2 (N6315, N6294, N6145);
or OR4 (N6316, N6275, N2684, N5781, N4032);
nor NOR2 (N6317, N6316, N524);
nand NAND2 (N6318, N6315, N2758);
buf BUF1 (N6319, N6313);
xor XOR2 (N6320, N6297, N2168);
nand NAND3 (N6321, N6320, N4263, N469);
buf BUF1 (N6322, N6311);
nand NAND2 (N6323, N6318, N5747);
or OR4 (N6324, N6291, N2315, N4796, N2423);
buf BUF1 (N6325, N6324);
not NOT1 (N6326, N6309);
not NOT1 (N6327, N6317);
nand NAND2 (N6328, N6327, N1937);
xor XOR2 (N6329, N6322, N920);
xor XOR2 (N6330, N6319, N2611);
and AND4 (N6331, N6328, N3660, N4281, N3343);
and AND4 (N6332, N6321, N2554, N2684, N5892);
buf BUF1 (N6333, N6331);
or OR3 (N6334, N6332, N5777, N2316);
nand NAND2 (N6335, N6326, N3451);
buf BUF1 (N6336, N6334);
nor NOR4 (N6337, N6323, N771, N3553, N386);
nand NAND2 (N6338, N6335, N1229);
not NOT1 (N6339, N6300);
and AND4 (N6340, N6337, N4312, N4179, N2538);
and AND2 (N6341, N6338, N4698);
and AND2 (N6342, N6341, N3599);
not NOT1 (N6343, N6340);
not NOT1 (N6344, N6330);
nor NOR4 (N6345, N6314, N2343, N3379, N2819);
buf BUF1 (N6346, N6329);
and AND4 (N6347, N6336, N1695, N2168, N3572);
or OR3 (N6348, N6347, N5435, N793);
buf BUF1 (N6349, N6308);
or OR3 (N6350, N6339, N3341, N6043);
not NOT1 (N6351, N6344);
or OR2 (N6352, N6348, N3347);
xor XOR2 (N6353, N6343, N4844);
nand NAND2 (N6354, N6350, N2365);
and AND3 (N6355, N6333, N6198, N1194);
buf BUF1 (N6356, N6352);
or OR3 (N6357, N6354, N1581, N1528);
not NOT1 (N6358, N6345);
not NOT1 (N6359, N6349);
and AND3 (N6360, N6342, N983, N6325);
xor XOR2 (N6361, N4851, N458);
not NOT1 (N6362, N6356);
nand NAND3 (N6363, N6351, N2852, N3749);
nand NAND2 (N6364, N6358, N6115);
or OR4 (N6365, N6362, N130, N5178, N3068);
or OR3 (N6366, N6357, N3210, N1533);
nor NOR2 (N6367, N6355, N3735);
nor NOR3 (N6368, N6361, N334, N3877);
nor NOR2 (N6369, N6363, N495);
not NOT1 (N6370, N6353);
nand NAND2 (N6371, N6368, N5496);
nand NAND2 (N6372, N6346, N4711);
buf BUF1 (N6373, N6369);
not NOT1 (N6374, N6373);
xor XOR2 (N6375, N6372, N5283);
not NOT1 (N6376, N6370);
or OR4 (N6377, N6367, N2689, N4919, N5603);
not NOT1 (N6378, N6377);
buf BUF1 (N6379, N6374);
and AND4 (N6380, N6371, N1399, N4262, N660);
xor XOR2 (N6381, N6360, N1911);
not NOT1 (N6382, N6366);
or OR4 (N6383, N6359, N168, N5827, N3326);
buf BUF1 (N6384, N6379);
xor XOR2 (N6385, N6381, N2439);
nor NOR4 (N6386, N6365, N2996, N1403, N1286);
buf BUF1 (N6387, N6382);
and AND4 (N6388, N6385, N4462, N2041, N2926);
buf BUF1 (N6389, N6378);
nor NOR2 (N6390, N6388, N2927);
nor NOR2 (N6391, N6384, N2003);
buf BUF1 (N6392, N6376);
buf BUF1 (N6393, N6389);
buf BUF1 (N6394, N6392);
nor NOR4 (N6395, N6393, N2831, N4575, N4285);
xor XOR2 (N6396, N6364, N465);
not NOT1 (N6397, N6394);
xor XOR2 (N6398, N6395, N445);
and AND3 (N6399, N6387, N4393, N2580);
and AND4 (N6400, N6383, N4770, N2199, N1665);
and AND3 (N6401, N6380, N823, N748);
and AND4 (N6402, N6390, N3176, N2426, N1030);
nor NOR3 (N6403, N6391, N3701, N1844);
nor NOR4 (N6404, N6402, N2691, N2460, N2614);
not NOT1 (N6405, N6397);
xor XOR2 (N6406, N6405, N4477);
nor NOR3 (N6407, N6399, N350, N733);
nor NOR4 (N6408, N6400, N4085, N174, N1547);
xor XOR2 (N6409, N6407, N4791);
or OR2 (N6410, N6401, N2409);
buf BUF1 (N6411, N6410);
nor NOR2 (N6412, N6406, N1603);
nor NOR4 (N6413, N6404, N2679, N3582, N4114);
nor NOR4 (N6414, N6408, N2779, N5646, N5520);
nand NAND4 (N6415, N6396, N2627, N6310, N1332);
nand NAND3 (N6416, N6386, N5406, N3879);
nor NOR4 (N6417, N6411, N2931, N2450, N1188);
nor NOR2 (N6418, N6409, N426);
not NOT1 (N6419, N6375);
or OR2 (N6420, N6416, N3590);
xor XOR2 (N6421, N6403, N2934);
xor XOR2 (N6422, N6420, N1636);
xor XOR2 (N6423, N6412, N4824);
or OR2 (N6424, N6418, N4844);
and AND3 (N6425, N6423, N5096, N5203);
or OR4 (N6426, N6421, N4935, N2179, N3839);
nor NOR4 (N6427, N6424, N4340, N3989, N1733);
and AND4 (N6428, N6417, N4146, N2651, N6025);
or OR2 (N6429, N6413, N1296);
and AND2 (N6430, N6414, N3283);
nand NAND4 (N6431, N6422, N713, N2232, N2622);
buf BUF1 (N6432, N6425);
or OR4 (N6433, N6398, N5971, N1346, N4005);
nor NOR3 (N6434, N6430, N3605, N2226);
nor NOR2 (N6435, N6415, N440);
not NOT1 (N6436, N6419);
buf BUF1 (N6437, N6428);
not NOT1 (N6438, N6435);
and AND2 (N6439, N6436, N3630);
xor XOR2 (N6440, N6429, N2787);
not NOT1 (N6441, N6431);
and AND2 (N6442, N6437, N3532);
nand NAND2 (N6443, N6433, N1236);
nand NAND3 (N6444, N6439, N3670, N2711);
nor NOR4 (N6445, N6438, N1172, N216, N678);
not NOT1 (N6446, N6426);
or OR2 (N6447, N6434, N1433);
buf BUF1 (N6448, N6427);
xor XOR2 (N6449, N6448, N5217);
nor NOR4 (N6450, N6440, N80, N3822, N1390);
or OR2 (N6451, N6443, N483);
and AND4 (N6452, N6449, N5925, N5371, N5569);
xor XOR2 (N6453, N6442, N1078);
xor XOR2 (N6454, N6441, N6422);
not NOT1 (N6455, N6432);
buf BUF1 (N6456, N6444);
not NOT1 (N6457, N6447);
not NOT1 (N6458, N6457);
nand NAND3 (N6459, N6445, N1524, N1701);
or OR3 (N6460, N6454, N3612, N4951);
or OR3 (N6461, N6451, N2445, N1743);
not NOT1 (N6462, N6453);
xor XOR2 (N6463, N6452, N3638);
or OR4 (N6464, N6450, N2765, N2856, N3209);
nor NOR2 (N6465, N6455, N1259);
and AND4 (N6466, N6458, N1950, N5625, N733);
or OR2 (N6467, N6461, N3237);
and AND3 (N6468, N6462, N5050, N3612);
and AND3 (N6469, N6456, N619, N5295);
nand NAND2 (N6470, N6468, N860);
or OR4 (N6471, N6470, N1690, N5340, N4864);
xor XOR2 (N6472, N6464, N5901);
nor NOR4 (N6473, N6471, N5274, N4112, N3535);
or OR3 (N6474, N6459, N87, N1131);
not NOT1 (N6475, N6469);
or OR3 (N6476, N6474, N4426, N127);
not NOT1 (N6477, N6465);
nor NOR2 (N6478, N6473, N6346);
nand NAND3 (N6479, N6460, N2292, N2809);
not NOT1 (N6480, N6472);
and AND3 (N6481, N6476, N1147, N4542);
nand NAND2 (N6482, N6481, N1220);
nor NOR2 (N6483, N6479, N4521);
not NOT1 (N6484, N6480);
and AND3 (N6485, N6483, N1025, N930);
and AND2 (N6486, N6482, N4849);
and AND3 (N6487, N6478, N1899, N4716);
or OR2 (N6488, N6446, N1301);
and AND3 (N6489, N6466, N6383, N5687);
and AND3 (N6490, N6486, N6470, N4229);
nand NAND2 (N6491, N6490, N601);
or OR2 (N6492, N6477, N6317);
or OR3 (N6493, N6485, N2834, N3548);
buf BUF1 (N6494, N6493);
buf BUF1 (N6495, N6494);
xor XOR2 (N6496, N6475, N6328);
nor NOR3 (N6497, N6487, N4493, N2377);
buf BUF1 (N6498, N6497);
buf BUF1 (N6499, N6463);
nand NAND4 (N6500, N6492, N105, N485, N90);
buf BUF1 (N6501, N6500);
and AND2 (N6502, N6484, N251);
or OR2 (N6503, N6489, N6203);
xor XOR2 (N6504, N6496, N4363);
nor NOR4 (N6505, N6488, N5034, N6018, N4526);
or OR4 (N6506, N6503, N630, N1035, N5037);
buf BUF1 (N6507, N6498);
xor XOR2 (N6508, N6467, N2285);
or OR4 (N6509, N6506, N1282, N4937, N4887);
xor XOR2 (N6510, N6509, N6063);
buf BUF1 (N6511, N6505);
not NOT1 (N6512, N6502);
buf BUF1 (N6513, N6499);
nand NAND4 (N6514, N6510, N1939, N5070, N4827);
or OR4 (N6515, N6511, N2610, N1400, N3257);
buf BUF1 (N6516, N6515);
or OR3 (N6517, N6507, N6444, N5415);
buf BUF1 (N6518, N6514);
nand NAND3 (N6519, N6512, N2613, N2257);
and AND4 (N6520, N6501, N2230, N2274, N2661);
and AND4 (N6521, N6516, N4141, N4521, N2721);
or OR2 (N6522, N6521, N5412);
and AND3 (N6523, N6508, N2117, N3166);
buf BUF1 (N6524, N6491);
buf BUF1 (N6525, N6523);
buf BUF1 (N6526, N6525);
nor NOR3 (N6527, N6522, N139, N6461);
nand NAND4 (N6528, N6504, N5202, N3352, N2238);
nor NOR2 (N6529, N6520, N2542);
or OR2 (N6530, N6524, N4445);
or OR2 (N6531, N6517, N1433);
buf BUF1 (N6532, N6518);
not NOT1 (N6533, N6519);
and AND3 (N6534, N6530, N5613, N1656);
nand NAND3 (N6535, N6526, N6526, N1329);
nand NAND3 (N6536, N6529, N3049, N5399);
and AND2 (N6537, N6535, N6385);
nand NAND4 (N6538, N6495, N5160, N2391, N1108);
buf BUF1 (N6539, N6528);
xor XOR2 (N6540, N6537, N3757);
not NOT1 (N6541, N6533);
or OR2 (N6542, N6541, N3422);
buf BUF1 (N6543, N6539);
or OR2 (N6544, N6534, N1912);
not NOT1 (N6545, N6543);
nand NAND3 (N6546, N6513, N1786, N3912);
and AND4 (N6547, N6540, N5050, N2858, N668);
and AND3 (N6548, N6531, N5477, N2591);
not NOT1 (N6549, N6527);
or OR3 (N6550, N6546, N407, N5710);
xor XOR2 (N6551, N6550, N4366);
nor NOR3 (N6552, N6547, N2460, N373);
xor XOR2 (N6553, N6551, N2362);
not NOT1 (N6554, N6549);
buf BUF1 (N6555, N6536);
and AND4 (N6556, N6545, N5785, N6265, N815);
buf BUF1 (N6557, N6555);
not NOT1 (N6558, N6542);
or OR2 (N6559, N6558, N4349);
not NOT1 (N6560, N6548);
and AND4 (N6561, N6544, N1981, N3499, N5573);
and AND3 (N6562, N6553, N880, N3211);
or OR3 (N6563, N6554, N782, N1853);
or OR4 (N6564, N6552, N4426, N4572, N208);
not NOT1 (N6565, N6538);
not NOT1 (N6566, N6557);
buf BUF1 (N6567, N6563);
and AND3 (N6568, N6556, N1881, N589);
nor NOR3 (N6569, N6562, N6232, N1246);
xor XOR2 (N6570, N6566, N4651);
or OR4 (N6571, N6567, N1020, N5403, N3547);
or OR4 (N6572, N6569, N3145, N2765, N387);
buf BUF1 (N6573, N6560);
nand NAND3 (N6574, N6565, N3739, N95);
or OR3 (N6575, N6568, N2346, N3849);
not NOT1 (N6576, N6571);
nand NAND3 (N6577, N6564, N2041, N4905);
buf BUF1 (N6578, N6575);
and AND4 (N6579, N6577, N1196, N1910, N679);
or OR3 (N6580, N6578, N6208, N4970);
buf BUF1 (N6581, N6574);
nor NOR2 (N6582, N6580, N611);
or OR4 (N6583, N6532, N2628, N3850, N6388);
xor XOR2 (N6584, N6576, N4081);
and AND3 (N6585, N6583, N4533, N43);
nand NAND3 (N6586, N6585, N6330, N5076);
and AND4 (N6587, N6584, N916, N3832, N1339);
or OR3 (N6588, N6586, N1402, N2452);
or OR2 (N6589, N6570, N39);
nand NAND4 (N6590, N6582, N1326, N5266, N4048);
xor XOR2 (N6591, N6573, N3404);
or OR2 (N6592, N6589, N1296);
nor NOR3 (N6593, N6579, N1953, N4015);
not NOT1 (N6594, N6581);
xor XOR2 (N6595, N6561, N5856);
buf BUF1 (N6596, N6593);
and AND3 (N6597, N6572, N1723, N5422);
and AND3 (N6598, N6591, N4963, N6160);
nand NAND4 (N6599, N6596, N2501, N4854, N5761);
nor NOR4 (N6600, N6592, N972, N5818, N3244);
and AND2 (N6601, N6599, N1958);
and AND3 (N6602, N6598, N1961, N511);
nor NOR3 (N6603, N6595, N1864, N6075);
buf BUF1 (N6604, N6603);
buf BUF1 (N6605, N6597);
nand NAND2 (N6606, N6587, N5537);
nor NOR3 (N6607, N6605, N2778, N4661);
and AND4 (N6608, N6604, N2303, N3931, N129);
xor XOR2 (N6609, N6559, N5504);
buf BUF1 (N6610, N6606);
and AND3 (N6611, N6601, N6175, N3675);
not NOT1 (N6612, N6610);
nand NAND2 (N6613, N6612, N2364);
or OR2 (N6614, N6613, N4419);
and AND3 (N6615, N6609, N2386, N4561);
buf BUF1 (N6616, N6600);
buf BUF1 (N6617, N6614);
not NOT1 (N6618, N6617);
xor XOR2 (N6619, N6611, N3565);
and AND4 (N6620, N6608, N6024, N6434, N551);
not NOT1 (N6621, N6594);
nand NAND3 (N6622, N6588, N5429, N4975);
nand NAND2 (N6623, N6619, N5663);
and AND2 (N6624, N6623, N4224);
nor NOR4 (N6625, N6620, N1405, N2712, N1065);
nor NOR2 (N6626, N6607, N6121);
xor XOR2 (N6627, N6625, N3381);
not NOT1 (N6628, N6624);
or OR2 (N6629, N6622, N853);
nand NAND2 (N6630, N6628, N6097);
nand NAND2 (N6631, N6626, N1127);
nand NAND3 (N6632, N6621, N418, N708);
nand NAND4 (N6633, N6615, N2862, N2640, N3524);
nor NOR4 (N6634, N6631, N3799, N5527, N4101);
and AND3 (N6635, N6633, N4593, N6349);
not NOT1 (N6636, N6590);
not NOT1 (N6637, N6629);
buf BUF1 (N6638, N6636);
nand NAND3 (N6639, N6637, N955, N5025);
or OR2 (N6640, N6630, N5851);
nand NAND4 (N6641, N6635, N2609, N2681, N4071);
xor XOR2 (N6642, N6638, N2193);
xor XOR2 (N6643, N6618, N1087);
and AND2 (N6644, N6627, N2806);
nor NOR3 (N6645, N6640, N480, N634);
buf BUF1 (N6646, N6602);
buf BUF1 (N6647, N6645);
buf BUF1 (N6648, N6632);
and AND2 (N6649, N6641, N4175);
nor NOR2 (N6650, N6642, N473);
nand NAND2 (N6651, N6650, N1693);
not NOT1 (N6652, N6646);
nand NAND2 (N6653, N6649, N896);
buf BUF1 (N6654, N6653);
buf BUF1 (N6655, N6644);
xor XOR2 (N6656, N6643, N468);
not NOT1 (N6657, N6651);
or OR3 (N6658, N6657, N2615, N1795);
nand NAND3 (N6659, N6655, N3716, N778);
xor XOR2 (N6660, N6639, N5400);
nand NAND3 (N6661, N6659, N2537, N6009);
or OR3 (N6662, N6647, N817, N2491);
nor NOR4 (N6663, N6661, N5896, N1537, N1406);
buf BUF1 (N6664, N6662);
not NOT1 (N6665, N6654);
not NOT1 (N6666, N6634);
buf BUF1 (N6667, N6658);
nor NOR4 (N6668, N6652, N2620, N6239, N3890);
nand NAND2 (N6669, N6648, N56);
xor XOR2 (N6670, N6664, N6159);
nor NOR2 (N6671, N6666, N556);
nor NOR3 (N6672, N6663, N3957, N6477);
nand NAND3 (N6673, N6616, N2942, N2482);
and AND3 (N6674, N6671, N4784, N3793);
not NOT1 (N6675, N6674);
not NOT1 (N6676, N6660);
and AND2 (N6677, N6668, N935);
or OR3 (N6678, N6672, N6355, N5477);
nor NOR4 (N6679, N6665, N5633, N5079, N1935);
buf BUF1 (N6680, N6669);
xor XOR2 (N6681, N6673, N3943);
nor NOR4 (N6682, N6670, N3532, N893, N1546);
not NOT1 (N6683, N6675);
xor XOR2 (N6684, N6678, N3401);
not NOT1 (N6685, N6679);
buf BUF1 (N6686, N6685);
and AND3 (N6687, N6680, N572, N5088);
xor XOR2 (N6688, N6677, N1311);
nor NOR2 (N6689, N6667, N2413);
buf BUF1 (N6690, N6676);
nor NOR4 (N6691, N6688, N6393, N2278, N5610);
not NOT1 (N6692, N6681);
xor XOR2 (N6693, N6691, N3808);
not NOT1 (N6694, N6656);
buf BUF1 (N6695, N6687);
nand NAND4 (N6696, N6686, N4653, N1297, N4539);
nor NOR4 (N6697, N6692, N3929, N2020, N4143);
or OR4 (N6698, N6684, N2707, N4845, N5648);
nand NAND3 (N6699, N6682, N644, N2291);
buf BUF1 (N6700, N6683);
nor NOR3 (N6701, N6697, N414, N3955);
or OR4 (N6702, N6690, N1932, N4913, N4006);
and AND4 (N6703, N6701, N1074, N358, N794);
and AND3 (N6704, N6693, N3686, N5688);
and AND2 (N6705, N6700, N3944);
nor NOR2 (N6706, N6694, N4688);
buf BUF1 (N6707, N6698);
or OR4 (N6708, N6702, N5451, N6627, N159);
nand NAND4 (N6709, N6705, N5953, N626, N4931);
not NOT1 (N6710, N6704);
nand NAND4 (N6711, N6710, N697, N4358, N1992);
and AND4 (N6712, N6711, N3965, N4864, N4020);
buf BUF1 (N6713, N6703);
buf BUF1 (N6714, N6696);
xor XOR2 (N6715, N6689, N3186);
nand NAND2 (N6716, N6715, N762);
nor NOR3 (N6717, N6714, N1036, N103);
or OR3 (N6718, N6713, N2264, N1043);
and AND2 (N6719, N6706, N2612);
xor XOR2 (N6720, N6719, N4316);
xor XOR2 (N6721, N6708, N1304);
or OR4 (N6722, N6699, N4452, N6678, N638);
not NOT1 (N6723, N6720);
buf BUF1 (N6724, N6721);
xor XOR2 (N6725, N6712, N1019);
nand NAND4 (N6726, N6695, N5181, N6616, N5708);
not NOT1 (N6727, N6709);
buf BUF1 (N6728, N6717);
nor NOR2 (N6729, N6718, N355);
or OR4 (N6730, N6725, N2005, N594, N548);
and AND3 (N6731, N6723, N1208, N872);
buf BUF1 (N6732, N6716);
nor NOR2 (N6733, N6724, N115);
xor XOR2 (N6734, N6731, N2905);
xor XOR2 (N6735, N6722, N4868);
xor XOR2 (N6736, N6730, N5878);
nand NAND3 (N6737, N6729, N3394, N5928);
buf BUF1 (N6738, N6736);
not NOT1 (N6739, N6728);
not NOT1 (N6740, N6727);
buf BUF1 (N6741, N6733);
nor NOR2 (N6742, N6707, N4959);
nand NAND2 (N6743, N6737, N2175);
not NOT1 (N6744, N6739);
not NOT1 (N6745, N6726);
nor NOR4 (N6746, N6732, N5908, N4231, N1518);
not NOT1 (N6747, N6742);
not NOT1 (N6748, N6747);
and AND3 (N6749, N6738, N4424, N5675);
nand NAND4 (N6750, N6744, N2603, N2319, N4073);
and AND4 (N6751, N6748, N5143, N6164, N2211);
nor NOR4 (N6752, N6746, N6153, N220, N370);
buf BUF1 (N6753, N6743);
buf BUF1 (N6754, N6735);
and AND2 (N6755, N6750, N6121);
buf BUF1 (N6756, N6753);
not NOT1 (N6757, N6754);
nor NOR4 (N6758, N6757, N4270, N3735, N2142);
buf BUF1 (N6759, N6745);
or OR3 (N6760, N6758, N1444, N279);
not NOT1 (N6761, N6740);
nand NAND4 (N6762, N6749, N4594, N3100, N559);
nor NOR2 (N6763, N6755, N4988);
xor XOR2 (N6764, N6763, N2655);
nor NOR4 (N6765, N6751, N3712, N3159, N1209);
buf BUF1 (N6766, N6760);
buf BUF1 (N6767, N6766);
or OR4 (N6768, N6762, N5139, N5163, N5018);
buf BUF1 (N6769, N6752);
and AND2 (N6770, N6764, N5888);
xor XOR2 (N6771, N6765, N5737);
and AND3 (N6772, N6756, N3901, N3691);
not NOT1 (N6773, N6759);
nor NOR3 (N6774, N6769, N5935, N2034);
or OR3 (N6775, N6767, N5378, N3635);
nand NAND2 (N6776, N6741, N1399);
nand NAND3 (N6777, N6774, N5644, N1839);
xor XOR2 (N6778, N6775, N6318);
not NOT1 (N6779, N6771);
nor NOR4 (N6780, N6779, N362, N5765, N3541);
or OR3 (N6781, N6777, N3978, N4053);
nor NOR2 (N6782, N6780, N3803);
and AND2 (N6783, N6768, N6370);
xor XOR2 (N6784, N6734, N6425);
and AND4 (N6785, N6781, N4690, N6489, N1537);
or OR4 (N6786, N6761, N3278, N5815, N1597);
xor XOR2 (N6787, N6776, N5307);
xor XOR2 (N6788, N6770, N6340);
and AND2 (N6789, N6772, N1258);
not NOT1 (N6790, N6783);
not NOT1 (N6791, N6787);
nand NAND3 (N6792, N6789, N3140, N2285);
not NOT1 (N6793, N6785);
nor NOR4 (N6794, N6786, N1892, N4352, N2141);
buf BUF1 (N6795, N6784);
nand NAND4 (N6796, N6795, N4947, N6264, N3377);
nor NOR3 (N6797, N6792, N772, N1565);
or OR3 (N6798, N6778, N90, N3298);
nor NOR2 (N6799, N6797, N6648);
buf BUF1 (N6800, N6790);
not NOT1 (N6801, N6800);
and AND2 (N6802, N6793, N272);
buf BUF1 (N6803, N6802);
not NOT1 (N6804, N6791);
xor XOR2 (N6805, N6804, N4957);
and AND2 (N6806, N6794, N3411);
or OR3 (N6807, N6798, N1130, N6095);
nand NAND3 (N6808, N6799, N2836, N5235);
buf BUF1 (N6809, N6801);
or OR4 (N6810, N6809, N6806, N5190, N5351);
buf BUF1 (N6811, N5620);
nor NOR3 (N6812, N6796, N3815, N2867);
not NOT1 (N6813, N6808);
or OR4 (N6814, N6788, N995, N37, N1322);
xor XOR2 (N6815, N6810, N2515);
buf BUF1 (N6816, N6814);
and AND3 (N6817, N6815, N3616, N2123);
xor XOR2 (N6818, N6816, N3994);
buf BUF1 (N6819, N6773);
nand NAND2 (N6820, N6819, N1548);
and AND3 (N6821, N6817, N4602, N2982);
not NOT1 (N6822, N6807);
nand NAND4 (N6823, N6803, N2737, N1091, N145);
not NOT1 (N6824, N6820);
xor XOR2 (N6825, N6812, N3906);
not NOT1 (N6826, N6811);
and AND3 (N6827, N6822, N4003, N3057);
or OR2 (N6828, N6782, N1567);
and AND3 (N6829, N6828, N6009, N4066);
xor XOR2 (N6830, N6823, N4247);
not NOT1 (N6831, N6827);
and AND3 (N6832, N6831, N1154, N3282);
nand NAND4 (N6833, N6832, N4573, N5851, N945);
nor NOR2 (N6834, N6813, N1324);
or OR3 (N6835, N6821, N3240, N6640);
nand NAND3 (N6836, N6835, N627, N1058);
nor NOR3 (N6837, N6824, N2842, N3867);
not NOT1 (N6838, N6805);
nor NOR4 (N6839, N6836, N3550, N2917, N3779);
and AND2 (N6840, N6826, N491);
or OR2 (N6841, N6825, N1864);
nor NOR4 (N6842, N6840, N6196, N5542, N5664);
not NOT1 (N6843, N6834);
buf BUF1 (N6844, N6843);
xor XOR2 (N6845, N6829, N5777);
not NOT1 (N6846, N6845);
or OR2 (N6847, N6833, N5314);
buf BUF1 (N6848, N6830);
nor NOR3 (N6849, N6818, N2320, N726);
not NOT1 (N6850, N6837);
buf BUF1 (N6851, N6842);
xor XOR2 (N6852, N6850, N2619);
xor XOR2 (N6853, N6846, N1382);
nand NAND2 (N6854, N6847, N511);
xor XOR2 (N6855, N6839, N2061);
buf BUF1 (N6856, N6852);
not NOT1 (N6857, N6854);
or OR2 (N6858, N6841, N5461);
and AND3 (N6859, N6855, N214, N4609);
not NOT1 (N6860, N6856);
xor XOR2 (N6861, N6860, N345);
and AND4 (N6862, N6851, N3827, N3569, N6289);
and AND3 (N6863, N6853, N4374, N3694);
xor XOR2 (N6864, N6848, N6046);
buf BUF1 (N6865, N6864);
and AND2 (N6866, N6849, N4338);
buf BUF1 (N6867, N6858);
nor NOR2 (N6868, N6859, N1208);
nand NAND2 (N6869, N6866, N5425);
or OR4 (N6870, N6844, N6251, N288, N6160);
nor NOR3 (N6871, N6838, N4192, N4943);
or OR2 (N6872, N6857, N2260);
xor XOR2 (N6873, N6870, N1300);
xor XOR2 (N6874, N6867, N1777);
and AND4 (N6875, N6861, N4099, N4275, N2855);
xor XOR2 (N6876, N6873, N1972);
not NOT1 (N6877, N6862);
buf BUF1 (N6878, N6869);
nor NOR3 (N6879, N6878, N968, N4416);
and AND2 (N6880, N6874, N2573);
xor XOR2 (N6881, N6880, N2171);
or OR4 (N6882, N6875, N5371, N4448, N432);
or OR3 (N6883, N6882, N145, N281);
and AND2 (N6884, N6883, N4057);
nand NAND2 (N6885, N6868, N539);
nand NAND2 (N6886, N6885, N3681);
or OR3 (N6887, N6881, N2886, N2310);
xor XOR2 (N6888, N6872, N5311);
and AND4 (N6889, N6884, N5421, N200, N6766);
nand NAND3 (N6890, N6879, N603, N5878);
nor NOR2 (N6891, N6877, N4225);
buf BUF1 (N6892, N6891);
nor NOR2 (N6893, N6886, N74);
not NOT1 (N6894, N6888);
not NOT1 (N6895, N6876);
buf BUF1 (N6896, N6890);
not NOT1 (N6897, N6889);
buf BUF1 (N6898, N6893);
buf BUF1 (N6899, N6865);
or OR2 (N6900, N6898, N1961);
nand NAND2 (N6901, N6900, N2837);
or OR4 (N6902, N6871, N5818, N6138, N754);
or OR4 (N6903, N6899, N4789, N1105, N1789);
xor XOR2 (N6904, N6897, N4178);
xor XOR2 (N6905, N6896, N1253);
and AND2 (N6906, N6904, N860);
buf BUF1 (N6907, N6892);
and AND3 (N6908, N6863, N6486, N1405);
buf BUF1 (N6909, N6908);
nor NOR2 (N6910, N6887, N6316);
nand NAND2 (N6911, N6902, N6084);
and AND3 (N6912, N6894, N3437, N5353);
and AND4 (N6913, N6901, N6339, N6462, N4378);
not NOT1 (N6914, N6909);
buf BUF1 (N6915, N6913);
xor XOR2 (N6916, N6906, N3041);
nand NAND2 (N6917, N6915, N1485);
nand NAND2 (N6918, N6912, N5018);
xor XOR2 (N6919, N6905, N4706);
xor XOR2 (N6920, N6916, N958);
nor NOR2 (N6921, N6907, N717);
or OR2 (N6922, N6911, N2853);
not NOT1 (N6923, N6914);
nor NOR2 (N6924, N6910, N879);
or OR2 (N6925, N6903, N6773);
xor XOR2 (N6926, N6919, N6230);
nand NAND2 (N6927, N6895, N784);
buf BUF1 (N6928, N6922);
and AND3 (N6929, N6926, N642, N5936);
nor NOR2 (N6930, N6918, N6107);
nand NAND3 (N6931, N6923, N6106, N3212);
buf BUF1 (N6932, N6931);
and AND3 (N6933, N6924, N6220, N6694);
nand NAND3 (N6934, N6917, N5955, N399);
not NOT1 (N6935, N6934);
and AND3 (N6936, N6927, N1387, N5253);
buf BUF1 (N6937, N6925);
or OR4 (N6938, N6920, N159, N1004, N5383);
buf BUF1 (N6939, N6928);
nand NAND4 (N6940, N6935, N1754, N5467, N4094);
not NOT1 (N6941, N6933);
nor NOR2 (N6942, N6941, N1958);
buf BUF1 (N6943, N6930);
nor NOR2 (N6944, N6938, N5613);
not NOT1 (N6945, N6921);
buf BUF1 (N6946, N6942);
buf BUF1 (N6947, N6943);
buf BUF1 (N6948, N6937);
and AND2 (N6949, N6945, N1486);
or OR2 (N6950, N6947, N4060);
or OR3 (N6951, N6936, N3665, N850);
buf BUF1 (N6952, N6951);
xor XOR2 (N6953, N6952, N5195);
not NOT1 (N6954, N6939);
and AND3 (N6955, N6932, N3275, N525);
nor NOR2 (N6956, N6940, N1360);
xor XOR2 (N6957, N6948, N259);
nand NAND2 (N6958, N6955, N3797);
nor NOR3 (N6959, N6958, N4994, N1373);
nand NAND3 (N6960, N6957, N1478, N2306);
or OR2 (N6961, N6953, N5999);
buf BUF1 (N6962, N6956);
not NOT1 (N6963, N6946);
and AND3 (N6964, N6961, N2605, N6677);
not NOT1 (N6965, N6929);
not NOT1 (N6966, N6959);
nor NOR3 (N6967, N6966, N5386, N4841);
or OR3 (N6968, N6944, N2795, N5428);
buf BUF1 (N6969, N6962);
nand NAND3 (N6970, N6967, N2974, N6154);
not NOT1 (N6971, N6968);
buf BUF1 (N6972, N6963);
nor NOR4 (N6973, N6969, N2204, N5150, N3834);
nor NOR2 (N6974, N6950, N1114);
or OR4 (N6975, N6970, N4975, N6876, N4995);
or OR4 (N6976, N6971, N3670, N2138, N2902);
and AND4 (N6977, N6949, N3985, N6747, N3078);
not NOT1 (N6978, N6965);
xor XOR2 (N6979, N6954, N3203);
nor NOR2 (N6980, N6978, N51);
xor XOR2 (N6981, N6974, N5262);
nand NAND4 (N6982, N6981, N195, N4079, N6418);
xor XOR2 (N6983, N6977, N6931);
not NOT1 (N6984, N6982);
buf BUF1 (N6985, N6973);
or OR4 (N6986, N6964, N5496, N4898, N2140);
or OR4 (N6987, N6976, N1449, N4190, N1893);
nor NOR3 (N6988, N6979, N6377, N2469);
or OR3 (N6989, N6972, N6520, N1779);
nand NAND4 (N6990, N6988, N3757, N6612, N3842);
not NOT1 (N6991, N6985);
nor NOR4 (N6992, N6984, N2948, N5410, N592);
or OR3 (N6993, N6975, N307, N4022);
xor XOR2 (N6994, N6992, N852);
and AND4 (N6995, N6987, N6100, N6113, N4283);
nand NAND2 (N6996, N6986, N2810);
not NOT1 (N6997, N6994);
and AND3 (N6998, N6990, N2673, N4431);
and AND3 (N6999, N6993, N839, N3698);
nor NOR4 (N7000, N6960, N6332, N1369, N5836);
and AND2 (N7001, N6980, N1323);
nand NAND3 (N7002, N6999, N98, N1430);
nor NOR4 (N7003, N6995, N1664, N5986, N3665);
nand NAND4 (N7004, N7001, N6381, N3905, N6721);
and AND4 (N7005, N6996, N1895, N5856, N2635);
nor NOR3 (N7006, N6998, N660, N6335);
or OR4 (N7007, N7005, N4899, N694, N2231);
not NOT1 (N7008, N7006);
nand NAND3 (N7009, N6989, N2595, N6551);
or OR3 (N7010, N6991, N6922, N714);
nand NAND2 (N7011, N7007, N173);
buf BUF1 (N7012, N7008);
not NOT1 (N7013, N7010);
not NOT1 (N7014, N7009);
xor XOR2 (N7015, N6983, N1904);
not NOT1 (N7016, N7000);
not NOT1 (N7017, N7012);
buf BUF1 (N7018, N7014);
nor NOR4 (N7019, N7013, N3889, N4079, N1637);
nand NAND3 (N7020, N6997, N6406, N1704);
nand NAND4 (N7021, N7004, N3924, N955, N3761);
or OR3 (N7022, N7011, N6472, N4206);
not NOT1 (N7023, N7015);
and AND4 (N7024, N7016, N3248, N4978, N3302);
nand NAND2 (N7025, N7024, N1516);
xor XOR2 (N7026, N7019, N3435);
or OR3 (N7027, N7022, N928, N4501);
or OR4 (N7028, N7025, N6369, N4598, N3766);
and AND4 (N7029, N7028, N537, N6620, N1194);
buf BUF1 (N7030, N7021);
nand NAND3 (N7031, N7020, N6018, N4329);
nand NAND4 (N7032, N7026, N5387, N4073, N3070);
nand NAND2 (N7033, N7018, N6404);
not NOT1 (N7034, N7002);
nand NAND4 (N7035, N7031, N3049, N1578, N1994);
nor NOR3 (N7036, N7029, N5936, N4336);
buf BUF1 (N7037, N7032);
or OR4 (N7038, N7033, N4208, N1727, N2442);
and AND2 (N7039, N7036, N395);
nand NAND2 (N7040, N7035, N2883);
not NOT1 (N7041, N7023);
nor NOR4 (N7042, N7034, N4726, N6847, N1851);
nand NAND4 (N7043, N7040, N3589, N2454, N3745);
nand NAND3 (N7044, N7039, N1423, N4171);
not NOT1 (N7045, N7030);
xor XOR2 (N7046, N7044, N5830);
not NOT1 (N7047, N7038);
buf BUF1 (N7048, N7047);
or OR2 (N7049, N7017, N717);
or OR2 (N7050, N7042, N1019);
xor XOR2 (N7051, N7043, N261);
buf BUF1 (N7052, N7037);
or OR3 (N7053, N7051, N2165, N1406);
xor XOR2 (N7054, N7053, N5935);
not NOT1 (N7055, N7027);
nor NOR4 (N7056, N7052, N888, N191, N800);
xor XOR2 (N7057, N7048, N4615);
nand NAND2 (N7058, N7057, N308);
or OR2 (N7059, N7003, N6287);
and AND3 (N7060, N7049, N6304, N1093);
and AND4 (N7061, N7050, N1209, N2961, N6030);
nor NOR3 (N7062, N7056, N1278, N1322);
nor NOR3 (N7063, N7046, N1665, N4311);
xor XOR2 (N7064, N7060, N6225);
nor NOR4 (N7065, N7061, N1529, N2119, N1116);
xor XOR2 (N7066, N7054, N402);
nor NOR2 (N7067, N7055, N2314);
nor NOR4 (N7068, N7065, N4023, N5324, N2428);
and AND3 (N7069, N7045, N4807, N341);
not NOT1 (N7070, N7064);
buf BUF1 (N7071, N7062);
buf BUF1 (N7072, N7068);
and AND3 (N7073, N7041, N6340, N1226);
nand NAND2 (N7074, N7067, N5302);
or OR4 (N7075, N7074, N1985, N6940, N6438);
and AND3 (N7076, N7058, N2744, N1729);
or OR2 (N7077, N7075, N4378);
nor NOR3 (N7078, N7063, N3767, N2650);
not NOT1 (N7079, N7077);
and AND4 (N7080, N7071, N62, N1078, N2456);
nor NOR3 (N7081, N7066, N4901, N5989);
nor NOR2 (N7082, N7059, N4110);
or OR2 (N7083, N7072, N4779);
nand NAND4 (N7084, N7082, N3654, N3255, N3211);
buf BUF1 (N7085, N7079);
buf BUF1 (N7086, N7081);
nand NAND3 (N7087, N7070, N59, N5800);
nor NOR3 (N7088, N7069, N2521, N4168);
nand NAND3 (N7089, N7086, N3410, N674);
xor XOR2 (N7090, N7078, N5043);
not NOT1 (N7091, N7083);
not NOT1 (N7092, N7085);
xor XOR2 (N7093, N7084, N3520);
nor NOR4 (N7094, N7093, N662, N134, N1193);
or OR2 (N7095, N7080, N6947);
not NOT1 (N7096, N7089);
not NOT1 (N7097, N7088);
xor XOR2 (N7098, N7095, N1622);
buf BUF1 (N7099, N7073);
and AND3 (N7100, N7087, N390, N2631);
xor XOR2 (N7101, N7097, N1167);
nor NOR3 (N7102, N7099, N2865, N5939);
not NOT1 (N7103, N7098);
nand NAND2 (N7104, N7100, N755);
not NOT1 (N7105, N7104);
buf BUF1 (N7106, N7091);
or OR4 (N7107, N7101, N3244, N4653, N1775);
nor NOR4 (N7108, N7090, N5561, N1294, N5396);
nor NOR2 (N7109, N7076, N4782);
buf BUF1 (N7110, N7092);
nand NAND4 (N7111, N7110, N4464, N2263, N881);
buf BUF1 (N7112, N7106);
not NOT1 (N7113, N7103);
or OR2 (N7114, N7105, N6154);
or OR4 (N7115, N7096, N4185, N4190, N3591);
and AND2 (N7116, N7094, N1483);
buf BUF1 (N7117, N7102);
buf BUF1 (N7118, N7115);
or OR3 (N7119, N7116, N2090, N6144);
nand NAND3 (N7120, N7118, N302, N3172);
or OR2 (N7121, N7112, N3639);
nor NOR2 (N7122, N7119, N4655);
or OR4 (N7123, N7108, N6362, N2911, N4695);
and AND2 (N7124, N7114, N1686);
not NOT1 (N7125, N7109);
nand NAND2 (N7126, N7123, N3508);
or OR3 (N7127, N7122, N1562, N2213);
not NOT1 (N7128, N7113);
buf BUF1 (N7129, N7120);
or OR4 (N7130, N7128, N1094, N606, N1170);
and AND2 (N7131, N7111, N4507);
nand NAND3 (N7132, N7125, N2249, N3400);
xor XOR2 (N7133, N7131, N2678);
xor XOR2 (N7134, N7117, N4788);
and AND2 (N7135, N7121, N4710);
or OR2 (N7136, N7133, N571);
nand NAND4 (N7137, N7132, N3188, N6484, N5080);
not NOT1 (N7138, N7107);
buf BUF1 (N7139, N7129);
or OR4 (N7140, N7139, N3725, N165, N6680);
or OR4 (N7141, N7136, N6154, N6363, N6033);
nor NOR3 (N7142, N7138, N3804, N5439);
buf BUF1 (N7143, N7127);
or OR2 (N7144, N7140, N4760);
nor NOR2 (N7145, N7141, N2217);
buf BUF1 (N7146, N7145);
xor XOR2 (N7147, N7134, N1216);
buf BUF1 (N7148, N7124);
buf BUF1 (N7149, N7130);
and AND3 (N7150, N7143, N2375, N7129);
or OR4 (N7151, N7146, N2942, N5105, N1441);
xor XOR2 (N7152, N7147, N4937);
not NOT1 (N7153, N7126);
not NOT1 (N7154, N7150);
not NOT1 (N7155, N7144);
not NOT1 (N7156, N7151);
xor XOR2 (N7157, N7135, N2311);
buf BUF1 (N7158, N7157);
nor NOR4 (N7159, N7155, N6564, N1114, N144);
xor XOR2 (N7160, N7137, N3310);
or OR3 (N7161, N7160, N880, N4517);
and AND4 (N7162, N7148, N354, N1019, N5491);
buf BUF1 (N7163, N7162);
buf BUF1 (N7164, N7142);
or OR2 (N7165, N7156, N4407);
xor XOR2 (N7166, N7159, N4660);
or OR4 (N7167, N7154, N2756, N4669, N5538);
nand NAND2 (N7168, N7158, N2332);
buf BUF1 (N7169, N7167);
or OR4 (N7170, N7166, N1138, N5512, N4229);
xor XOR2 (N7171, N7163, N825);
xor XOR2 (N7172, N7165, N6327);
and AND4 (N7173, N7152, N6300, N4437, N3097);
or OR2 (N7174, N7149, N268);
or OR3 (N7175, N7161, N582, N5336);
buf BUF1 (N7176, N7164);
buf BUF1 (N7177, N7173);
nand NAND3 (N7178, N7174, N6050, N6373);
xor XOR2 (N7179, N7178, N6999);
and AND4 (N7180, N7179, N3075, N3983, N3113);
and AND4 (N7181, N7180, N4690, N406, N454);
xor XOR2 (N7182, N7172, N6384);
xor XOR2 (N7183, N7182, N4181);
not NOT1 (N7184, N7177);
xor XOR2 (N7185, N7181, N1569);
not NOT1 (N7186, N7169);
nand NAND2 (N7187, N7176, N5477);
not NOT1 (N7188, N7175);
nand NAND4 (N7189, N7183, N4510, N4398, N4168);
nor NOR2 (N7190, N7188, N5218);
not NOT1 (N7191, N7184);
nor NOR3 (N7192, N7171, N4072, N3597);
not NOT1 (N7193, N7187);
and AND2 (N7194, N7186, N1236);
nand NAND3 (N7195, N7190, N397, N2567);
buf BUF1 (N7196, N7193);
nand NAND4 (N7197, N7192, N3080, N2151, N5981);
nor NOR2 (N7198, N7197, N2050);
buf BUF1 (N7199, N7198);
buf BUF1 (N7200, N7191);
or OR4 (N7201, N7194, N3846, N2467, N2809);
not NOT1 (N7202, N7153);
xor XOR2 (N7203, N7200, N3968);
buf BUF1 (N7204, N7185);
not NOT1 (N7205, N7195);
not NOT1 (N7206, N7168);
or OR3 (N7207, N7196, N1993, N6324);
or OR2 (N7208, N7206, N2073);
buf BUF1 (N7209, N7189);
and AND4 (N7210, N7203, N4702, N5585, N4109);
buf BUF1 (N7211, N7199);
nor NOR2 (N7212, N7201, N6665);
nor NOR3 (N7213, N7208, N3804, N7171);
nand NAND2 (N7214, N7212, N943);
and AND3 (N7215, N7211, N1779, N1021);
xor XOR2 (N7216, N7207, N998);
nor NOR2 (N7217, N7214, N3160);
xor XOR2 (N7218, N7202, N5166);
and AND2 (N7219, N7218, N4521);
and AND3 (N7220, N7209, N4114, N1297);
not NOT1 (N7221, N7217);
not NOT1 (N7222, N7219);
and AND3 (N7223, N7204, N5022, N1645);
nor NOR2 (N7224, N7216, N4783);
nand NAND3 (N7225, N7215, N5959, N2218);
nor NOR4 (N7226, N7223, N7075, N6323, N3952);
xor XOR2 (N7227, N7222, N5804);
not NOT1 (N7228, N7221);
xor XOR2 (N7229, N7205, N4804);
buf BUF1 (N7230, N7224);
and AND2 (N7231, N7228, N4786);
and AND3 (N7232, N7229, N959, N645);
and AND2 (N7233, N7220, N4526);
or OR4 (N7234, N7230, N6481, N3602, N3108);
or OR3 (N7235, N7225, N5095, N3898);
nor NOR3 (N7236, N7231, N4793, N3582);
and AND3 (N7237, N7232, N6336, N3168);
nor NOR3 (N7238, N7235, N715, N2084);
and AND4 (N7239, N7238, N2627, N3573, N5107);
nor NOR3 (N7240, N7213, N4605, N914);
nand NAND4 (N7241, N7239, N429, N2150, N263);
or OR2 (N7242, N7241, N5817);
nor NOR2 (N7243, N7210, N6842);
nor NOR3 (N7244, N7233, N6878, N2353);
nand NAND4 (N7245, N7242, N5629, N810, N6938);
not NOT1 (N7246, N7243);
not NOT1 (N7247, N7227);
not NOT1 (N7248, N7234);
nor NOR4 (N7249, N7240, N2586, N334, N5821);
nor NOR3 (N7250, N7245, N2874, N820);
nor NOR2 (N7251, N7244, N1839);
not NOT1 (N7252, N7226);
not NOT1 (N7253, N7237);
nor NOR4 (N7254, N7170, N1992, N2505, N4448);
xor XOR2 (N7255, N7254, N4982);
xor XOR2 (N7256, N7253, N2496);
nand NAND2 (N7257, N7255, N5560);
buf BUF1 (N7258, N7252);
xor XOR2 (N7259, N7248, N870);
buf BUF1 (N7260, N7258);
not NOT1 (N7261, N7249);
and AND4 (N7262, N7261, N6578, N4629, N7244);
nor NOR2 (N7263, N7259, N6378);
nand NAND2 (N7264, N7263, N5546);
xor XOR2 (N7265, N7264, N6607);
not NOT1 (N7266, N7250);
nor NOR3 (N7267, N7251, N5037, N5813);
xor XOR2 (N7268, N7256, N4915);
and AND2 (N7269, N7260, N3312);
nand NAND3 (N7270, N7262, N4138, N3887);
xor XOR2 (N7271, N7269, N382);
buf BUF1 (N7272, N7265);
nor NOR3 (N7273, N7268, N58, N3739);
buf BUF1 (N7274, N7271);
or OR3 (N7275, N7274, N2949, N3443);
buf BUF1 (N7276, N7247);
nor NOR2 (N7277, N7272, N6294);
and AND4 (N7278, N7276, N93, N3609, N2672);
or OR2 (N7279, N7267, N184);
nor NOR2 (N7280, N7279, N4451);
and AND4 (N7281, N7275, N4379, N358, N1901);
and AND4 (N7282, N7246, N2254, N674, N3361);
and AND3 (N7283, N7270, N6499, N4418);
nor NOR4 (N7284, N7266, N4510, N603, N4366);
xor XOR2 (N7285, N7280, N288);
not NOT1 (N7286, N7282);
not NOT1 (N7287, N7283);
or OR4 (N7288, N7286, N7027, N5914, N4931);
nand NAND3 (N7289, N7236, N4236, N3865);
and AND4 (N7290, N7288, N477, N4464, N106);
buf BUF1 (N7291, N7284);
nor NOR4 (N7292, N7290, N4307, N6299, N4135);
not NOT1 (N7293, N7281);
nand NAND2 (N7294, N7277, N4136);
nor NOR3 (N7295, N7289, N6693, N3572);
not NOT1 (N7296, N7294);
not NOT1 (N7297, N7273);
or OR3 (N7298, N7278, N5815, N6444);
buf BUF1 (N7299, N7297);
or OR4 (N7300, N7293, N2635, N3396, N85);
or OR4 (N7301, N7285, N5528, N1891, N5134);
xor XOR2 (N7302, N7295, N6214);
xor XOR2 (N7303, N7302, N4943);
not NOT1 (N7304, N7287);
or OR4 (N7305, N7291, N7033, N3667, N2291);
not NOT1 (N7306, N7301);
buf BUF1 (N7307, N7292);
not NOT1 (N7308, N7307);
nor NOR2 (N7309, N7296, N2821);
nand NAND3 (N7310, N7299, N1940, N3562);
not NOT1 (N7311, N7304);
nor NOR3 (N7312, N7308, N7153, N5155);
buf BUF1 (N7313, N7300);
nand NAND2 (N7314, N7312, N5493);
buf BUF1 (N7315, N7314);
nand NAND4 (N7316, N7303, N391, N6603, N2344);
buf BUF1 (N7317, N7298);
and AND2 (N7318, N7313, N2287);
nor NOR4 (N7319, N7306, N5711, N2384, N2697);
nand NAND3 (N7320, N7315, N2432, N6549);
xor XOR2 (N7321, N7317, N6926);
xor XOR2 (N7322, N7318, N1211);
nand NAND2 (N7323, N7309, N6199);
buf BUF1 (N7324, N7311);
not NOT1 (N7325, N7316);
or OR2 (N7326, N7323, N3319);
nand NAND3 (N7327, N7257, N181, N7036);
or OR2 (N7328, N7305, N2982);
or OR4 (N7329, N7322, N131, N3130, N5681);
nand NAND2 (N7330, N7327, N5479);
nand NAND3 (N7331, N7319, N3264, N1708);
and AND2 (N7332, N7330, N4347);
not NOT1 (N7333, N7325);
xor XOR2 (N7334, N7326, N1914);
nand NAND2 (N7335, N7332, N6521);
buf BUF1 (N7336, N7328);
not NOT1 (N7337, N7335);
buf BUF1 (N7338, N7321);
or OR4 (N7339, N7336, N2466, N6113, N791);
or OR4 (N7340, N7337, N4868, N4559, N3019);
or OR3 (N7341, N7334, N3332, N5766);
buf BUF1 (N7342, N7333);
nand NAND3 (N7343, N7329, N6887, N6237);
nor NOR4 (N7344, N7338, N2936, N1032, N6370);
and AND2 (N7345, N7340, N2926);
buf BUF1 (N7346, N7341);
xor XOR2 (N7347, N7343, N4710);
and AND2 (N7348, N7345, N4016);
nor NOR3 (N7349, N7346, N2389, N5080);
or OR3 (N7350, N7339, N3534, N2643);
or OR2 (N7351, N7342, N3849);
buf BUF1 (N7352, N7349);
and AND2 (N7353, N7310, N1461);
nand NAND3 (N7354, N7352, N7175, N3708);
buf BUF1 (N7355, N7331);
not NOT1 (N7356, N7344);
xor XOR2 (N7357, N7353, N370);
nor NOR4 (N7358, N7356, N1251, N2026, N2213);
or OR2 (N7359, N7351, N684);
nor NOR4 (N7360, N7320, N4348, N1907, N3841);
nand NAND2 (N7361, N7354, N6549);
buf BUF1 (N7362, N7358);
nor NOR2 (N7363, N7357, N4538);
buf BUF1 (N7364, N7348);
not NOT1 (N7365, N7360);
nor NOR4 (N7366, N7359, N4308, N3802, N6921);
not NOT1 (N7367, N7361);
xor XOR2 (N7368, N7367, N430);
or OR2 (N7369, N7366, N5948);
and AND4 (N7370, N7350, N6937, N2802, N4913);
and AND3 (N7371, N7362, N3942, N2610);
nor NOR2 (N7372, N7371, N4266);
buf BUF1 (N7373, N7355);
nand NAND4 (N7374, N7363, N2403, N1833, N2019);
nor NOR3 (N7375, N7373, N3127, N881);
xor XOR2 (N7376, N7375, N2672);
xor XOR2 (N7377, N7364, N2572);
nor NOR3 (N7378, N7374, N2484, N5103);
buf BUF1 (N7379, N7369);
nand NAND4 (N7380, N7378, N4645, N6056, N4884);
nor NOR2 (N7381, N7347, N5123);
not NOT1 (N7382, N7365);
and AND3 (N7383, N7368, N7349, N1555);
or OR4 (N7384, N7324, N1722, N2003, N2445);
xor XOR2 (N7385, N7380, N7101);
nand NAND4 (N7386, N7376, N2878, N43, N783);
and AND4 (N7387, N7382, N852, N4131, N6749);
buf BUF1 (N7388, N7370);
buf BUF1 (N7389, N7383);
nor NOR4 (N7390, N7381, N2755, N4359, N4931);
not NOT1 (N7391, N7379);
not NOT1 (N7392, N7387);
not NOT1 (N7393, N7388);
nand NAND4 (N7394, N7385, N6109, N4819, N1400);
buf BUF1 (N7395, N7384);
buf BUF1 (N7396, N7389);
nand NAND3 (N7397, N7391, N3247, N6236);
nand NAND2 (N7398, N7395, N5247);
xor XOR2 (N7399, N7390, N670);
nor NOR3 (N7400, N7399, N4847, N2200);
not NOT1 (N7401, N7396);
or OR3 (N7402, N7372, N1116, N7032);
not NOT1 (N7403, N7392);
buf BUF1 (N7404, N7403);
and AND2 (N7405, N7398, N257);
nor NOR3 (N7406, N7394, N721, N5884);
xor XOR2 (N7407, N7405, N7066);
xor XOR2 (N7408, N7407, N1990);
not NOT1 (N7409, N7401);
or OR4 (N7410, N7402, N6075, N6873, N6704);
nand NAND4 (N7411, N7409, N6950, N6554, N3557);
or OR2 (N7412, N7377, N3007);
xor XOR2 (N7413, N7408, N6328);
buf BUF1 (N7414, N7386);
not NOT1 (N7415, N7393);
buf BUF1 (N7416, N7406);
nand NAND2 (N7417, N7410, N5218);
xor XOR2 (N7418, N7400, N3127);
xor XOR2 (N7419, N7416, N1216);
and AND3 (N7420, N7411, N2856, N3669);
and AND2 (N7421, N7397, N4884);
nand NAND4 (N7422, N7420, N405, N6154, N3275);
and AND3 (N7423, N7417, N3407, N2425);
not NOT1 (N7424, N7422);
not NOT1 (N7425, N7418);
buf BUF1 (N7426, N7419);
nor NOR2 (N7427, N7415, N5407);
or OR2 (N7428, N7427, N1275);
and AND2 (N7429, N7412, N3034);
buf BUF1 (N7430, N7404);
and AND4 (N7431, N7413, N3459, N2567, N640);
nor NOR4 (N7432, N7425, N2278, N6074, N5448);
and AND4 (N7433, N7424, N5681, N636, N6062);
or OR2 (N7434, N7414, N1009);
buf BUF1 (N7435, N7432);
or OR2 (N7436, N7431, N1807);
and AND3 (N7437, N7421, N3265, N3853);
and AND2 (N7438, N7428, N2043);
not NOT1 (N7439, N7438);
xor XOR2 (N7440, N7423, N2939);
nand NAND4 (N7441, N7429, N4301, N292, N6844);
nor NOR2 (N7442, N7430, N2100);
nand NAND3 (N7443, N7435, N5502, N2969);
and AND4 (N7444, N7434, N707, N800, N1744);
nor NOR2 (N7445, N7436, N4265);
and AND4 (N7446, N7445, N4428, N4691, N5008);
not NOT1 (N7447, N7437);
buf BUF1 (N7448, N7439);
or OR2 (N7449, N7433, N7344);
nor NOR4 (N7450, N7440, N2857, N3814, N5540);
or OR3 (N7451, N7442, N7283, N424);
xor XOR2 (N7452, N7446, N2811);
nand NAND4 (N7453, N7441, N2149, N5832, N2169);
and AND3 (N7454, N7450, N4595, N6073);
nand NAND3 (N7455, N7451, N3914, N1496);
and AND3 (N7456, N7426, N3483, N5130);
and AND2 (N7457, N7449, N4502);
xor XOR2 (N7458, N7443, N2441);
not NOT1 (N7459, N7455);
nand NAND3 (N7460, N7454, N4943, N6218);
buf BUF1 (N7461, N7456);
nor NOR2 (N7462, N7460, N5756);
buf BUF1 (N7463, N7452);
or OR3 (N7464, N7447, N6816, N3460);
nor NOR3 (N7465, N7463, N6828, N1396);
nand NAND2 (N7466, N7457, N5325);
buf BUF1 (N7467, N7462);
not NOT1 (N7468, N7461);
nor NOR4 (N7469, N7466, N1283, N3910, N151);
nand NAND4 (N7470, N7453, N463, N2471, N1066);
not NOT1 (N7471, N7444);
nand NAND3 (N7472, N7469, N1036, N579);
buf BUF1 (N7473, N7470);
and AND4 (N7474, N7468, N2629, N7316, N5146);
and AND2 (N7475, N7473, N6264);
not NOT1 (N7476, N7465);
not NOT1 (N7477, N7472);
or OR2 (N7478, N7467, N874);
not NOT1 (N7479, N7448);
not NOT1 (N7480, N7479);
xor XOR2 (N7481, N7459, N4851);
buf BUF1 (N7482, N7478);
or OR3 (N7483, N7471, N6385, N6730);
and AND4 (N7484, N7482, N4759, N4438, N3419);
xor XOR2 (N7485, N7464, N6100);
nor NOR3 (N7486, N7485, N2943, N3683);
not NOT1 (N7487, N7458);
xor XOR2 (N7488, N7475, N5693);
and AND2 (N7489, N7474, N2118);
not NOT1 (N7490, N7480);
xor XOR2 (N7491, N7477, N331);
not NOT1 (N7492, N7490);
or OR4 (N7493, N7492, N5701, N1502, N5854);
xor XOR2 (N7494, N7481, N5244);
not NOT1 (N7495, N7486);
or OR2 (N7496, N7493, N1761);
or OR3 (N7497, N7483, N1850, N4567);
xor XOR2 (N7498, N7488, N7319);
nor NOR2 (N7499, N7495, N1218);
or OR4 (N7500, N7489, N3396, N3628, N6816);
buf BUF1 (N7501, N7491);
nand NAND2 (N7502, N7494, N7091);
and AND2 (N7503, N7487, N3968);
nor NOR3 (N7504, N7496, N5066, N4077);
or OR2 (N7505, N7498, N599);
not NOT1 (N7506, N7497);
not NOT1 (N7507, N7502);
buf BUF1 (N7508, N7505);
buf BUF1 (N7509, N7508);
not NOT1 (N7510, N7484);
xor XOR2 (N7511, N7509, N3952);
not NOT1 (N7512, N7511);
or OR2 (N7513, N7501, N5539);
nor NOR2 (N7514, N7504, N5254);
and AND3 (N7515, N7507, N4356, N4174);
and AND4 (N7516, N7510, N7196, N1036, N2122);
or OR2 (N7517, N7513, N3592);
nand NAND2 (N7518, N7499, N538);
not NOT1 (N7519, N7518);
xor XOR2 (N7520, N7476, N1864);
nor NOR3 (N7521, N7515, N5800, N2504);
nor NOR3 (N7522, N7512, N3054, N4065);
nand NAND2 (N7523, N7506, N2342);
nor NOR4 (N7524, N7521, N625, N6811, N4244);
xor XOR2 (N7525, N7523, N1085);
nor NOR3 (N7526, N7519, N4159, N1365);
or OR2 (N7527, N7503, N6053);
nand NAND3 (N7528, N7524, N2503, N6355);
buf BUF1 (N7529, N7526);
nand NAND2 (N7530, N7516, N666);
xor XOR2 (N7531, N7529, N233);
not NOT1 (N7532, N7522);
and AND4 (N7533, N7500, N6033, N5249, N4725);
buf BUF1 (N7534, N7517);
and AND2 (N7535, N7531, N2742);
not NOT1 (N7536, N7530);
nand NAND2 (N7537, N7525, N6426);
nand NAND2 (N7538, N7527, N3297);
xor XOR2 (N7539, N7536, N6988);
nand NAND2 (N7540, N7520, N4404);
nor NOR2 (N7541, N7535, N4356);
not NOT1 (N7542, N7538);
nor NOR2 (N7543, N7537, N293);
xor XOR2 (N7544, N7532, N4831);
buf BUF1 (N7545, N7528);
xor XOR2 (N7546, N7541, N6981);
buf BUF1 (N7547, N7544);
not NOT1 (N7548, N7545);
nand NAND4 (N7549, N7546, N188, N5248, N4690);
not NOT1 (N7550, N7534);
buf BUF1 (N7551, N7548);
xor XOR2 (N7552, N7543, N547);
or OR3 (N7553, N7550, N2385, N3996);
and AND4 (N7554, N7547, N4020, N4401, N5245);
not NOT1 (N7555, N7514);
xor XOR2 (N7556, N7553, N6747);
nand NAND3 (N7557, N7540, N5277, N5912);
not NOT1 (N7558, N7549);
nand NAND3 (N7559, N7533, N5910, N5130);
and AND3 (N7560, N7557, N2358, N5995);
nand NAND3 (N7561, N7551, N5993, N4831);
and AND3 (N7562, N7556, N4426, N804);
nand NAND2 (N7563, N7552, N4333);
or OR2 (N7564, N7559, N2417);
nor NOR4 (N7565, N7558, N6731, N2387, N6892);
nor NOR3 (N7566, N7560, N5406, N2277);
buf BUF1 (N7567, N7539);
or OR3 (N7568, N7564, N7438, N2578);
xor XOR2 (N7569, N7554, N3723);
nor NOR3 (N7570, N7567, N130, N3791);
not NOT1 (N7571, N7566);
and AND2 (N7572, N7569, N1229);
and AND4 (N7573, N7572, N6618, N2812, N2920);
or OR2 (N7574, N7565, N2727);
xor XOR2 (N7575, N7568, N4388);
nand NAND3 (N7576, N7574, N913, N222);
and AND3 (N7577, N7576, N3413, N4676);
nor NOR2 (N7578, N7573, N1407);
nand NAND2 (N7579, N7563, N6223);
and AND4 (N7580, N7579, N5409, N5978, N225);
or OR4 (N7581, N7561, N1070, N933, N4214);
xor XOR2 (N7582, N7575, N6894);
nand NAND3 (N7583, N7581, N2987, N1965);
xor XOR2 (N7584, N7578, N4788);
or OR3 (N7585, N7562, N2456, N1489);
nand NAND3 (N7586, N7582, N1354, N2893);
nor NOR3 (N7587, N7577, N180, N4315);
and AND3 (N7588, N7584, N622, N4259);
or OR2 (N7589, N7587, N2943);
buf BUF1 (N7590, N7585);
xor XOR2 (N7591, N7580, N5239);
not NOT1 (N7592, N7591);
nor NOR3 (N7593, N7570, N3142, N2079);
nor NOR4 (N7594, N7590, N492, N6356, N4467);
xor XOR2 (N7595, N7555, N2414);
nand NAND4 (N7596, N7586, N2356, N490, N5734);
xor XOR2 (N7597, N7592, N1398);
buf BUF1 (N7598, N7542);
nand NAND2 (N7599, N7588, N287);
buf BUF1 (N7600, N7595);
nor NOR4 (N7601, N7598, N1843, N4403, N6179);
xor XOR2 (N7602, N7571, N2850);
xor XOR2 (N7603, N7596, N5750);
nor NOR3 (N7604, N7602, N5591, N1638);
nand NAND3 (N7605, N7593, N4792, N3839);
or OR3 (N7606, N7603, N3309, N755);
xor XOR2 (N7607, N7597, N1808);
not NOT1 (N7608, N7599);
and AND3 (N7609, N7608, N5231, N5858);
or OR4 (N7610, N7594, N4102, N6840, N1945);
nand NAND2 (N7611, N7601, N6768);
not NOT1 (N7612, N7610);
not NOT1 (N7613, N7600);
and AND2 (N7614, N7589, N4774);
nor NOR4 (N7615, N7604, N4602, N2737, N6195);
and AND2 (N7616, N7609, N3424);
nand NAND4 (N7617, N7616, N6332, N1714, N7034);
xor XOR2 (N7618, N7617, N2319);
buf BUF1 (N7619, N7605);
nand NAND2 (N7620, N7614, N1408);
buf BUF1 (N7621, N7612);
buf BUF1 (N7622, N7615);
and AND2 (N7623, N7613, N162);
nand NAND4 (N7624, N7619, N6858, N7502, N1975);
not NOT1 (N7625, N7620);
nand NAND2 (N7626, N7618, N5309);
nor NOR2 (N7627, N7607, N192);
and AND4 (N7628, N7624, N5, N3617, N196);
not NOT1 (N7629, N7583);
not NOT1 (N7630, N7621);
buf BUF1 (N7631, N7627);
nor NOR4 (N7632, N7628, N4991, N1375, N623);
nor NOR3 (N7633, N7625, N3858, N6154);
buf BUF1 (N7634, N7633);
nor NOR2 (N7635, N7629, N6041);
xor XOR2 (N7636, N7611, N5637);
or OR4 (N7637, N7631, N5419, N4624, N3606);
or OR3 (N7638, N7636, N1844, N2060);
buf BUF1 (N7639, N7632);
nand NAND2 (N7640, N7635, N1345);
nor NOR2 (N7641, N7638, N503);
buf BUF1 (N7642, N7640);
buf BUF1 (N7643, N7637);
xor XOR2 (N7644, N7643, N6713);
not NOT1 (N7645, N7642);
xor XOR2 (N7646, N7622, N293);
xor XOR2 (N7647, N7639, N1629);
xor XOR2 (N7648, N7646, N1236);
buf BUF1 (N7649, N7644);
and AND3 (N7650, N7634, N3603, N3927);
nor NOR4 (N7651, N7645, N7085, N4247, N994);
buf BUF1 (N7652, N7651);
xor XOR2 (N7653, N7649, N6443);
not NOT1 (N7654, N7650);
nor NOR2 (N7655, N7653, N5680);
nor NOR3 (N7656, N7626, N2891, N7213);
nor NOR4 (N7657, N7656, N7256, N2789, N5792);
xor XOR2 (N7658, N7648, N3483);
or OR4 (N7659, N7606, N1672, N3788, N6885);
nand NAND4 (N7660, N7657, N4117, N7124, N6967);
xor XOR2 (N7661, N7654, N2931);
nor NOR4 (N7662, N7623, N2541, N5753, N3448);
or OR2 (N7663, N7658, N7356);
buf BUF1 (N7664, N7661);
buf BUF1 (N7665, N7647);
buf BUF1 (N7666, N7630);
nand NAND2 (N7667, N7655, N2181);
nand NAND4 (N7668, N7665, N3114, N4847, N7413);
buf BUF1 (N7669, N7641);
or OR4 (N7670, N7668, N1543, N2647, N6806);
or OR2 (N7671, N7666, N5492);
or OR3 (N7672, N7660, N5564, N5378);
xor XOR2 (N7673, N7670, N19);
nor NOR3 (N7674, N7662, N3317, N6030);
or OR4 (N7675, N7672, N3492, N5705, N1011);
not NOT1 (N7676, N7659);
or OR3 (N7677, N7667, N569, N923);
xor XOR2 (N7678, N7671, N7103);
and AND4 (N7679, N7652, N3522, N3086, N2602);
buf BUF1 (N7680, N7676);
and AND3 (N7681, N7675, N6109, N5354);
nor NOR3 (N7682, N7680, N7124, N6531);
xor XOR2 (N7683, N7682, N4899);
and AND4 (N7684, N7683, N7619, N5639, N4817);
xor XOR2 (N7685, N7684, N3666);
not NOT1 (N7686, N7677);
nor NOR4 (N7687, N7686, N1565, N5646, N3478);
or OR3 (N7688, N7664, N3332, N2013);
nand NAND3 (N7689, N7673, N5375, N1430);
buf BUF1 (N7690, N7688);
and AND4 (N7691, N7663, N2014, N2078, N1301);
xor XOR2 (N7692, N7674, N6856);
xor XOR2 (N7693, N7678, N3802);
nand NAND3 (N7694, N7669, N6503, N1168);
nor NOR4 (N7695, N7681, N5480, N6949, N3112);
nand NAND4 (N7696, N7690, N235, N496, N5615);
buf BUF1 (N7697, N7685);
nand NAND2 (N7698, N7687, N7636);
buf BUF1 (N7699, N7693);
not NOT1 (N7700, N7689);
xor XOR2 (N7701, N7699, N3183);
not NOT1 (N7702, N7696);
nor NOR2 (N7703, N7698, N2160);
nand NAND3 (N7704, N7691, N7068, N7050);
nor NOR3 (N7705, N7704, N3622, N555);
nand NAND2 (N7706, N7702, N6941);
xor XOR2 (N7707, N7700, N5490);
or OR4 (N7708, N7706, N189, N190, N3423);
nand NAND4 (N7709, N7707, N3343, N2582, N5741);
and AND3 (N7710, N7692, N4851, N3378);
or OR4 (N7711, N7679, N6299, N2065, N6106);
buf BUF1 (N7712, N7695);
buf BUF1 (N7713, N7694);
xor XOR2 (N7714, N7701, N4474);
buf BUF1 (N7715, N7708);
xor XOR2 (N7716, N7705, N1385);
nor NOR3 (N7717, N7710, N4585, N1761);
nand NAND4 (N7718, N7712, N1430, N1492, N7394);
not NOT1 (N7719, N7709);
buf BUF1 (N7720, N7697);
nor NOR3 (N7721, N7718, N4384, N860);
and AND3 (N7722, N7719, N6704, N4670);
nand NAND3 (N7723, N7715, N3270, N3506);
not NOT1 (N7724, N7723);
buf BUF1 (N7725, N7722);
or OR2 (N7726, N7724, N4235);
buf BUF1 (N7727, N7720);
nand NAND3 (N7728, N7721, N6785, N2327);
and AND2 (N7729, N7727, N5725);
buf BUF1 (N7730, N7729);
not NOT1 (N7731, N7730);
xor XOR2 (N7732, N7728, N5265);
or OR3 (N7733, N7703, N6647, N6848);
xor XOR2 (N7734, N7713, N4807);
nand NAND4 (N7735, N7734, N2932, N1307, N6001);
not NOT1 (N7736, N7717);
xor XOR2 (N7737, N7732, N6710);
not NOT1 (N7738, N7725);
buf BUF1 (N7739, N7737);
not NOT1 (N7740, N7739);
buf BUF1 (N7741, N7711);
nor NOR3 (N7742, N7716, N3600, N2227);
or OR3 (N7743, N7740, N3723, N1464);
nand NAND4 (N7744, N7731, N5229, N2851, N1977);
and AND4 (N7745, N7743, N2429, N2077, N428);
or OR3 (N7746, N7714, N6759, N2159);
xor XOR2 (N7747, N7738, N2227);
nor NOR4 (N7748, N7744, N6801, N2177, N4831);
nor NOR3 (N7749, N7745, N6681, N2904);
or OR2 (N7750, N7746, N4974);
nand NAND3 (N7751, N7750, N3520, N1882);
nor NOR3 (N7752, N7733, N7137, N2640);
nand NAND4 (N7753, N7752, N5313, N3284, N6185);
buf BUF1 (N7754, N7741);
nand NAND3 (N7755, N7748, N4998, N4002);
buf BUF1 (N7756, N7755);
not NOT1 (N7757, N7747);
xor XOR2 (N7758, N7753, N7612);
buf BUF1 (N7759, N7758);
buf BUF1 (N7760, N7754);
or OR4 (N7761, N7751, N6572, N3085, N2288);
or OR4 (N7762, N7756, N81, N5104, N7024);
xor XOR2 (N7763, N7757, N6873);
not NOT1 (N7764, N7762);
nor NOR2 (N7765, N7749, N578);
buf BUF1 (N7766, N7736);
or OR2 (N7767, N7761, N3528);
buf BUF1 (N7768, N7735);
xor XOR2 (N7769, N7766, N5218);
nor NOR2 (N7770, N7765, N4445);
and AND3 (N7771, N7742, N32, N2211);
xor XOR2 (N7772, N7770, N924);
or OR4 (N7773, N7768, N4956, N164, N4496);
nand NAND4 (N7774, N7767, N2685, N5279, N2113);
or OR3 (N7775, N7763, N3611, N4442);
nand NAND4 (N7776, N7760, N2446, N408, N4642);
buf BUF1 (N7777, N7771);
nor NOR4 (N7778, N7777, N7262, N5978, N6641);
xor XOR2 (N7779, N7775, N5409);
xor XOR2 (N7780, N7776, N2757);
not NOT1 (N7781, N7772);
buf BUF1 (N7782, N7780);
not NOT1 (N7783, N7764);
and AND4 (N7784, N7783, N2385, N1032, N2039);
nor NOR3 (N7785, N7779, N4159, N6228);
nand NAND3 (N7786, N7782, N1128, N6157);
or OR2 (N7787, N7781, N684);
nor NOR3 (N7788, N7773, N341, N1270);
buf BUF1 (N7789, N7787);
nand NAND2 (N7790, N7784, N4883);
nor NOR3 (N7791, N7769, N6221, N5815);
xor XOR2 (N7792, N7789, N5553);
buf BUF1 (N7793, N7774);
nor NOR4 (N7794, N7785, N5843, N4822, N6296);
not NOT1 (N7795, N7726);
xor XOR2 (N7796, N7794, N366);
buf BUF1 (N7797, N7791);
not NOT1 (N7798, N7790);
not NOT1 (N7799, N7793);
not NOT1 (N7800, N7759);
nor NOR2 (N7801, N7786, N4639);
nand NAND4 (N7802, N7792, N3515, N4555, N4047);
or OR4 (N7803, N7801, N6538, N5248, N1245);
buf BUF1 (N7804, N7802);
xor XOR2 (N7805, N7795, N6535);
and AND2 (N7806, N7778, N1566);
not NOT1 (N7807, N7805);
or OR3 (N7808, N7788, N4519, N4143);
nor NOR3 (N7809, N7807, N3744, N3851);
xor XOR2 (N7810, N7806, N5477);
and AND4 (N7811, N7809, N5952, N7562, N1257);
and AND2 (N7812, N7808, N5505);
nor NOR3 (N7813, N7797, N4208, N7087);
not NOT1 (N7814, N7810);
not NOT1 (N7815, N7811);
nor NOR4 (N7816, N7796, N3871, N3853, N2481);
xor XOR2 (N7817, N7814, N359);
not NOT1 (N7818, N7813);
nor NOR2 (N7819, N7803, N1811);
xor XOR2 (N7820, N7818, N2010);
nor NOR4 (N7821, N7820, N5893, N2610, N3902);
and AND4 (N7822, N7815, N1614, N5933, N5369);
or OR2 (N7823, N7819, N1070);
and AND4 (N7824, N7798, N5708, N2870, N5085);
nand NAND2 (N7825, N7821, N1489);
not NOT1 (N7826, N7823);
nor NOR3 (N7827, N7817, N1242, N5777);
nand NAND4 (N7828, N7824, N2535, N4209, N1429);
nand NAND2 (N7829, N7822, N7508);
nand NAND2 (N7830, N7804, N4986);
and AND4 (N7831, N7828, N5308, N3383, N4176);
nand NAND4 (N7832, N7830, N7078, N2393, N5197);
or OR2 (N7833, N7812, N5556);
not NOT1 (N7834, N7799);
or OR3 (N7835, N7827, N3932, N5508);
nor NOR3 (N7836, N7832, N1460, N6424);
buf BUF1 (N7837, N7835);
buf BUF1 (N7838, N7800);
buf BUF1 (N7839, N7837);
and AND2 (N7840, N7834, N6860);
not NOT1 (N7841, N7825);
nor NOR2 (N7842, N7841, N4440);
not NOT1 (N7843, N7826);
nand NAND3 (N7844, N7836, N2099, N7150);
nor NOR2 (N7845, N7833, N1474);
nand NAND3 (N7846, N7844, N3642, N1685);
and AND3 (N7847, N7831, N3625, N5330);
or OR2 (N7848, N7845, N4141);
nand NAND3 (N7849, N7846, N5121, N560);
buf BUF1 (N7850, N7816);
nand NAND2 (N7851, N7839, N2751);
or OR2 (N7852, N7848, N7559);
or OR3 (N7853, N7850, N2983, N5927);
nor NOR4 (N7854, N7842, N7563, N959, N3829);
not NOT1 (N7855, N7847);
not NOT1 (N7856, N7843);
nand NAND3 (N7857, N7851, N7660, N6943);
buf BUF1 (N7858, N7840);
xor XOR2 (N7859, N7853, N2921);
nand NAND3 (N7860, N7856, N144, N2912);
nand NAND3 (N7861, N7829, N1341, N2936);
and AND3 (N7862, N7838, N3896, N6982);
and AND3 (N7863, N7854, N6079, N4174);
buf BUF1 (N7864, N7859);
and AND2 (N7865, N7852, N2984);
or OR4 (N7866, N7857, N2692, N1293, N4179);
xor XOR2 (N7867, N7864, N2074);
xor XOR2 (N7868, N7860, N6179);
xor XOR2 (N7869, N7849, N6987);
and AND4 (N7870, N7867, N3863, N7327, N6608);
xor XOR2 (N7871, N7870, N5187);
xor XOR2 (N7872, N7863, N6492);
nor NOR4 (N7873, N7869, N1347, N2734, N555);
nor NOR4 (N7874, N7871, N1117, N5342, N3143);
nand NAND3 (N7875, N7868, N2432, N4024);
buf BUF1 (N7876, N7855);
nand NAND2 (N7877, N7874, N7416);
not NOT1 (N7878, N7865);
not NOT1 (N7879, N7876);
not NOT1 (N7880, N7879);
nand NAND4 (N7881, N7858, N1897, N7656, N140);
nand NAND3 (N7882, N7861, N1066, N3544);
not NOT1 (N7883, N7877);
not NOT1 (N7884, N7878);
nand NAND3 (N7885, N7873, N4448, N3674);
not NOT1 (N7886, N7883);
buf BUF1 (N7887, N7880);
not NOT1 (N7888, N7885);
nor NOR3 (N7889, N7884, N506, N234);
nor NOR4 (N7890, N7887, N4665, N6821, N1089);
nand NAND3 (N7891, N7862, N2067, N564);
not NOT1 (N7892, N7890);
buf BUF1 (N7893, N7882);
buf BUF1 (N7894, N7866);
xor XOR2 (N7895, N7888, N180);
not NOT1 (N7896, N7875);
nor NOR4 (N7897, N7872, N120, N3169, N7819);
buf BUF1 (N7898, N7889);
xor XOR2 (N7899, N7893, N2403);
buf BUF1 (N7900, N7898);
nand NAND3 (N7901, N7899, N2819, N7112);
buf BUF1 (N7902, N7901);
nor NOR3 (N7903, N7881, N4665, N2600);
nand NAND4 (N7904, N7903, N6962, N4542, N5476);
xor XOR2 (N7905, N7902, N2779);
or OR4 (N7906, N7892, N6658, N6194, N3718);
not NOT1 (N7907, N7905);
or OR4 (N7908, N7886, N4140, N356, N6709);
and AND3 (N7909, N7904, N7824, N6992);
xor XOR2 (N7910, N7894, N2659);
not NOT1 (N7911, N7900);
or OR3 (N7912, N7910, N2076, N7374);
nor NOR4 (N7913, N7908, N3017, N4048, N5763);
and AND2 (N7914, N7897, N5126);
and AND4 (N7915, N7896, N1193, N1516, N7880);
or OR3 (N7916, N7913, N7337, N1971);
xor XOR2 (N7917, N7907, N3385);
or OR3 (N7918, N7895, N3798, N1765);
or OR4 (N7919, N7906, N1684, N6973, N4054);
buf BUF1 (N7920, N7914);
or OR3 (N7921, N7916, N3474, N5304);
buf BUF1 (N7922, N7918);
nand NAND3 (N7923, N7909, N2695, N5774);
nor NOR4 (N7924, N7921, N5227, N708, N3924);
nor NOR4 (N7925, N7919, N1099, N1720, N7022);
or OR4 (N7926, N7925, N777, N6141, N7403);
xor XOR2 (N7927, N7923, N1091);
nand NAND4 (N7928, N7891, N505, N2029, N5271);
and AND2 (N7929, N7912, N5086);
nor NOR2 (N7930, N7928, N2137);
nand NAND4 (N7931, N7922, N5200, N5200, N4088);
buf BUF1 (N7932, N7924);
nand NAND2 (N7933, N7927, N3485);
not NOT1 (N7934, N7917);
nand NAND3 (N7935, N7929, N233, N2049);
buf BUF1 (N7936, N7911);
buf BUF1 (N7937, N7926);
not NOT1 (N7938, N7932);
buf BUF1 (N7939, N7937);
not NOT1 (N7940, N7915);
not NOT1 (N7941, N7936);
buf BUF1 (N7942, N7920);
not NOT1 (N7943, N7939);
and AND4 (N7944, N7941, N3998, N7414, N3974);
and AND2 (N7945, N7944, N3495);
and AND4 (N7946, N7935, N2815, N4355, N4068);
xor XOR2 (N7947, N7931, N3905);
nand NAND2 (N7948, N7933, N6342);
and AND4 (N7949, N7943, N1616, N7104, N5185);
nand NAND2 (N7950, N7948, N6029);
not NOT1 (N7951, N7940);
nor NOR4 (N7952, N7946, N5417, N5264, N1991);
nand NAND3 (N7953, N7938, N1706, N5515);
not NOT1 (N7954, N7951);
not NOT1 (N7955, N7949);
not NOT1 (N7956, N7950);
buf BUF1 (N7957, N7947);
xor XOR2 (N7958, N7945, N5953);
not NOT1 (N7959, N7957);
nand NAND2 (N7960, N7953, N7948);
and AND4 (N7961, N7959, N3020, N7246, N697);
buf BUF1 (N7962, N7961);
buf BUF1 (N7963, N7956);
or OR3 (N7964, N7960, N4773, N4222);
or OR4 (N7965, N7962, N4436, N4220, N4876);
nor NOR4 (N7966, N7964, N4517, N3588, N7581);
and AND4 (N7967, N7958, N3935, N7181, N7471);
nand NAND4 (N7968, N7966, N4688, N6123, N6391);
not NOT1 (N7969, N7967);
nor NOR3 (N7970, N7968, N4281, N4610);
xor XOR2 (N7971, N7963, N3872);
nor NOR2 (N7972, N7955, N3880);
and AND3 (N7973, N7965, N3137, N6732);
not NOT1 (N7974, N7973);
not NOT1 (N7975, N7972);
nand NAND2 (N7976, N7952, N4958);
buf BUF1 (N7977, N7975);
nand NAND3 (N7978, N7930, N2483, N3338);
not NOT1 (N7979, N7934);
xor XOR2 (N7980, N7971, N3754);
xor XOR2 (N7981, N7954, N1182);
and AND4 (N7982, N7979, N1257, N4714, N2646);
not NOT1 (N7983, N7970);
or OR4 (N7984, N7982, N247, N5123, N3818);
or OR3 (N7985, N7978, N1494, N1322);
and AND4 (N7986, N7969, N2028, N1636, N2155);
not NOT1 (N7987, N7977);
and AND2 (N7988, N7981, N5925);
xor XOR2 (N7989, N7942, N3967);
nand NAND2 (N7990, N7974, N3616);
xor XOR2 (N7991, N7986, N2492);
or OR2 (N7992, N7980, N935);
and AND4 (N7993, N7991, N4068, N1532, N3239);
buf BUF1 (N7994, N7983);
nand NAND2 (N7995, N7990, N728);
not NOT1 (N7996, N7994);
nor NOR3 (N7997, N7976, N5715, N4369);
xor XOR2 (N7998, N7997, N5697);
or OR4 (N7999, N7998, N4752, N1380, N7341);
nand NAND4 (N8000, N7987, N3747, N7829, N6183);
or OR3 (N8001, N7995, N1748, N6469);
xor XOR2 (N8002, N8000, N2477);
nand NAND2 (N8003, N8001, N1320);
xor XOR2 (N8004, N7984, N6358);
nand NAND3 (N8005, N7989, N476, N4918);
buf BUF1 (N8006, N8004);
buf BUF1 (N8007, N7996);
nor NOR3 (N8008, N8006, N5183, N1257);
buf BUF1 (N8009, N8003);
xor XOR2 (N8010, N7992, N315);
not NOT1 (N8011, N7985);
not NOT1 (N8012, N8011);
xor XOR2 (N8013, N8007, N2818);
nor NOR4 (N8014, N8008, N137, N302, N3126);
and AND3 (N8015, N8005, N3589, N164);
buf BUF1 (N8016, N8009);
buf BUF1 (N8017, N7993);
not NOT1 (N8018, N8010);
and AND3 (N8019, N8013, N3032, N1443);
not NOT1 (N8020, N8015);
nor NOR4 (N8021, N8002, N1849, N2232, N3859);
xor XOR2 (N8022, N8017, N3852);
xor XOR2 (N8023, N8014, N3895);
or OR2 (N8024, N8022, N177);
or OR2 (N8025, N8020, N1740);
or OR2 (N8026, N8024, N1674);
and AND4 (N8027, N8012, N5166, N5512, N5205);
nor NOR3 (N8028, N8019, N4, N1216);
and AND3 (N8029, N7988, N767, N7173);
nor NOR2 (N8030, N8023, N5209);
nand NAND3 (N8031, N8018, N612, N5195);
or OR3 (N8032, N8031, N92, N3808);
or OR2 (N8033, N8030, N5536);
not NOT1 (N8034, N8033);
or OR4 (N8035, N8029, N7959, N7180, N3761);
not NOT1 (N8036, N8025);
or OR4 (N8037, N8028, N3996, N3426, N2900);
or OR4 (N8038, N8034, N4096, N5700, N7949);
xor XOR2 (N8039, N8035, N3582);
not NOT1 (N8040, N8021);
and AND4 (N8041, N8026, N7943, N2799, N2138);
nand NAND2 (N8042, N8039, N1980);
buf BUF1 (N8043, N8042);
nor NOR3 (N8044, N8037, N7288, N2081);
and AND4 (N8045, N8040, N5025, N6955, N1932);
not NOT1 (N8046, N8036);
nor NOR4 (N8047, N8043, N4351, N5573, N2353);
nand NAND4 (N8048, N8047, N6628, N7138, N6711);
or OR2 (N8049, N8027, N1129);
buf BUF1 (N8050, N8046);
xor XOR2 (N8051, N8048, N5825);
not NOT1 (N8052, N8041);
nor NOR2 (N8053, N8016, N2939);
or OR2 (N8054, N8053, N7365);
xor XOR2 (N8055, N8051, N2304);
and AND2 (N8056, N8032, N1444);
nand NAND2 (N8057, N8049, N3048);
buf BUF1 (N8058, N8057);
or OR2 (N8059, N8050, N6494);
xor XOR2 (N8060, N8059, N184);
nand NAND4 (N8061, N8054, N4045, N5635, N2336);
nand NAND3 (N8062, N8055, N6086, N6390);
and AND2 (N8063, N8052, N4830);
not NOT1 (N8064, N8060);
not NOT1 (N8065, N8056);
or OR4 (N8066, N8064, N4550, N3665, N1355);
nor NOR3 (N8067, N8065, N3513, N1293);
and AND4 (N8068, N8038, N266, N4819, N2446);
not NOT1 (N8069, N8068);
not NOT1 (N8070, N8067);
and AND4 (N8071, N8061, N4403, N4383, N4263);
not NOT1 (N8072, N8069);
or OR2 (N8073, N8045, N1885);
nor NOR3 (N8074, N8073, N7454, N1535);
or OR3 (N8075, N8062, N294, N7703);
xor XOR2 (N8076, N8072, N1746);
or OR4 (N8077, N7999, N7134, N1433, N5085);
nand NAND3 (N8078, N8063, N5257, N344);
nor NOR3 (N8079, N8076, N4957, N4352);
nand NAND4 (N8080, N8074, N7363, N4114, N5242);
buf BUF1 (N8081, N8078);
nor NOR3 (N8082, N8044, N1793, N5013);
buf BUF1 (N8083, N8077);
or OR4 (N8084, N8079, N3946, N2036, N7975);
xor XOR2 (N8085, N8075, N5544);
and AND3 (N8086, N8058, N6989, N1758);
or OR2 (N8087, N8082, N3738);
or OR2 (N8088, N8071, N6049);
nand NAND2 (N8089, N8084, N5042);
not NOT1 (N8090, N8081);
nand NAND4 (N8091, N8070, N5824, N7107, N6298);
not NOT1 (N8092, N8086);
buf BUF1 (N8093, N8090);
nand NAND3 (N8094, N8088, N2557, N3687);
or OR3 (N8095, N8066, N1817, N6073);
xor XOR2 (N8096, N8089, N7784);
or OR2 (N8097, N8091, N7123);
or OR3 (N8098, N8094, N7346, N6881);
and AND3 (N8099, N8087, N843, N4027);
nand NAND2 (N8100, N8080, N4851);
buf BUF1 (N8101, N8096);
buf BUF1 (N8102, N8100);
xor XOR2 (N8103, N8095, N2062);
or OR2 (N8104, N8097, N7999);
nor NOR2 (N8105, N8098, N2059);
nand NAND3 (N8106, N8105, N74, N4687);
nor NOR4 (N8107, N8103, N2240, N7907, N5914);
and AND4 (N8108, N8092, N845, N1028, N3391);
not NOT1 (N8109, N8108);
nor NOR3 (N8110, N8109, N7555, N4733);
nand NAND3 (N8111, N8110, N2606, N6349);
xor XOR2 (N8112, N8099, N2432);
or OR2 (N8113, N8102, N3994);
buf BUF1 (N8114, N8113);
nor NOR2 (N8115, N8112, N5964);
nor NOR4 (N8116, N8114, N5644, N1354, N2272);
nor NOR2 (N8117, N8115, N7615);
nor NOR3 (N8118, N8116, N4563, N5938);
nor NOR2 (N8119, N8104, N6284);
nor NOR2 (N8120, N8117, N162);
and AND4 (N8121, N8083, N2785, N863, N4704);
and AND2 (N8122, N8121, N3553);
and AND4 (N8123, N8107, N6931, N2175, N1847);
nand NAND2 (N8124, N8122, N2778);
xor XOR2 (N8125, N8093, N2742);
xor XOR2 (N8126, N8119, N7013);
or OR3 (N8127, N8126, N1496, N1461);
nand NAND3 (N8128, N8123, N1799, N1463);
nor NOR2 (N8129, N8128, N7817);
and AND3 (N8130, N8101, N3500, N7146);
xor XOR2 (N8131, N8124, N5998);
buf BUF1 (N8132, N8106);
nor NOR2 (N8133, N8120, N3365);
or OR2 (N8134, N8130, N6835);
not NOT1 (N8135, N8129);
xor XOR2 (N8136, N8118, N6845);
xor XOR2 (N8137, N8085, N6974);
not NOT1 (N8138, N8127);
xor XOR2 (N8139, N8133, N4839);
buf BUF1 (N8140, N8134);
nor NOR4 (N8141, N8132, N5268, N7336, N1955);
and AND2 (N8142, N8139, N7166);
or OR2 (N8143, N8136, N6227);
or OR3 (N8144, N8137, N7138, N362);
not NOT1 (N8145, N8143);
and AND2 (N8146, N8141, N3077);
not NOT1 (N8147, N8111);
xor XOR2 (N8148, N8147, N68);
or OR4 (N8149, N8146, N5757, N6420, N969);
not NOT1 (N8150, N8145);
nor NOR3 (N8151, N8131, N4079, N2977);
not NOT1 (N8152, N8135);
not NOT1 (N8153, N8140);
nand NAND4 (N8154, N8151, N4130, N4148, N3771);
or OR3 (N8155, N8138, N2726, N4939);
not NOT1 (N8156, N8148);
and AND2 (N8157, N8152, N2963);
or OR3 (N8158, N8142, N7995, N1719);
buf BUF1 (N8159, N8157);
or OR2 (N8160, N8144, N6302);
xor XOR2 (N8161, N8158, N7199);
nand NAND4 (N8162, N8156, N4575, N3847, N4118);
xor XOR2 (N8163, N8149, N7576);
nand NAND4 (N8164, N8162, N3862, N3301, N5175);
and AND3 (N8165, N8155, N7606, N3315);
and AND3 (N8166, N8165, N7642, N698);
nor NOR2 (N8167, N8159, N186);
nand NAND2 (N8168, N8153, N5678);
or OR2 (N8169, N8150, N6238);
not NOT1 (N8170, N8166);
or OR4 (N8171, N8163, N154, N6024, N4382);
buf BUF1 (N8172, N8125);
xor XOR2 (N8173, N8171, N2240);
xor XOR2 (N8174, N8172, N3911);
not NOT1 (N8175, N8164);
buf BUF1 (N8176, N8160);
or OR2 (N8177, N8170, N3311);
xor XOR2 (N8178, N8174, N4162);
nand NAND4 (N8179, N8176, N7465, N5133, N2856);
xor XOR2 (N8180, N8179, N4585);
not NOT1 (N8181, N8175);
not NOT1 (N8182, N8178);
nand NAND2 (N8183, N8161, N1448);
or OR4 (N8184, N8168, N925, N507, N4908);
and AND3 (N8185, N8169, N6550, N1036);
or OR4 (N8186, N8173, N3321, N3961, N333);
or OR3 (N8187, N8182, N406, N1199);
and AND4 (N8188, N8154, N6794, N4510, N112);
nor NOR4 (N8189, N8186, N8009, N7698, N7882);
or OR2 (N8190, N8187, N4986);
nor NOR3 (N8191, N8190, N281, N4426);
nand NAND4 (N8192, N8177, N1778, N333, N3026);
nor NOR3 (N8193, N8183, N5829, N3173);
buf BUF1 (N8194, N8180);
or OR2 (N8195, N8184, N1283);
nor NOR4 (N8196, N8167, N7383, N300, N6696);
not NOT1 (N8197, N8189);
nor NOR3 (N8198, N8193, N4344, N414);
not NOT1 (N8199, N8196);
nand NAND4 (N8200, N8198, N2964, N5371, N360);
and AND2 (N8201, N8191, N4740);
xor XOR2 (N8202, N8197, N6355);
xor XOR2 (N8203, N8199, N5027);
and AND4 (N8204, N8188, N7219, N6952, N2666);
and AND4 (N8205, N8203, N3824, N2, N5002);
nand NAND4 (N8206, N8201, N405, N3155, N2052);
not NOT1 (N8207, N8181);
and AND2 (N8208, N8207, N7981);
nand NAND4 (N8209, N8185, N4068, N6316, N548);
or OR2 (N8210, N8192, N3873);
buf BUF1 (N8211, N8202);
xor XOR2 (N8212, N8200, N6757);
nor NOR2 (N8213, N8209, N6256);
not NOT1 (N8214, N8206);
or OR3 (N8215, N8205, N4627, N6405);
nor NOR4 (N8216, N8195, N5543, N7857, N4929);
buf BUF1 (N8217, N8213);
nand NAND2 (N8218, N8215, N7029);
nor NOR3 (N8219, N8217, N3200, N5685);
xor XOR2 (N8220, N8218, N4998);
and AND4 (N8221, N8204, N6085, N6715, N2856);
nor NOR3 (N8222, N8210, N3342, N2274);
and AND2 (N8223, N8216, N5141);
buf BUF1 (N8224, N8219);
not NOT1 (N8225, N8211);
buf BUF1 (N8226, N8225);
nor NOR2 (N8227, N8221, N2831);
and AND2 (N8228, N8224, N7256);
not NOT1 (N8229, N8223);
not NOT1 (N8230, N8226);
or OR4 (N8231, N8228, N6444, N6180, N7159);
and AND2 (N8232, N8214, N4070);
or OR4 (N8233, N8231, N2859, N5000, N864);
nor NOR3 (N8234, N8227, N3763, N8106);
buf BUF1 (N8235, N8234);
and AND2 (N8236, N8208, N5210);
xor XOR2 (N8237, N8220, N7251);
xor XOR2 (N8238, N8194, N6439);
and AND2 (N8239, N8229, N6245);
buf BUF1 (N8240, N8232);
not NOT1 (N8241, N8236);
or OR3 (N8242, N8233, N8070, N1254);
and AND3 (N8243, N8238, N5100, N7671);
xor XOR2 (N8244, N8239, N239);
not NOT1 (N8245, N8240);
nand NAND3 (N8246, N8242, N5202, N4339);
buf BUF1 (N8247, N8246);
buf BUF1 (N8248, N8245);
not NOT1 (N8249, N8212);
nor NOR3 (N8250, N8230, N7871, N4469);
nand NAND3 (N8251, N8243, N7298, N83);
xor XOR2 (N8252, N8250, N4028);
xor XOR2 (N8253, N8249, N1215);
buf BUF1 (N8254, N8235);
xor XOR2 (N8255, N8244, N4159);
or OR3 (N8256, N8251, N982, N5155);
buf BUF1 (N8257, N8237);
and AND2 (N8258, N8254, N439);
buf BUF1 (N8259, N8258);
nand NAND4 (N8260, N8241, N2304, N7926, N7490);
or OR2 (N8261, N8222, N524);
and AND2 (N8262, N8247, N7096);
nand NAND4 (N8263, N8260, N3457, N92, N4365);
nand NAND4 (N8264, N8255, N1242, N3628, N5441);
nand NAND2 (N8265, N8259, N8047);
and AND3 (N8266, N8257, N6350, N5838);
or OR3 (N8267, N8264, N7204, N729);
or OR3 (N8268, N8256, N6198, N1779);
nand NAND3 (N8269, N8267, N6241, N6886);
not NOT1 (N8270, N8266);
nor NOR3 (N8271, N8269, N4766, N916);
xor XOR2 (N8272, N8252, N271);
or OR2 (N8273, N8272, N5001);
not NOT1 (N8274, N8268);
nor NOR3 (N8275, N8253, N5776, N2486);
not NOT1 (N8276, N8275);
nor NOR4 (N8277, N8276, N3437, N3321, N3412);
buf BUF1 (N8278, N8271);
nor NOR2 (N8279, N8261, N2067);
or OR3 (N8280, N8262, N1690, N5544);
buf BUF1 (N8281, N8280);
not NOT1 (N8282, N8274);
nand NAND3 (N8283, N8279, N3259, N1527);
nor NOR3 (N8284, N8248, N2754, N5327);
and AND3 (N8285, N8270, N3459, N4640);
not NOT1 (N8286, N8281);
buf BUF1 (N8287, N8285);
not NOT1 (N8288, N8265);
not NOT1 (N8289, N8263);
and AND3 (N8290, N8277, N4874, N8273);
nand NAND3 (N8291, N5072, N1688, N3432);
xor XOR2 (N8292, N8286, N5218);
nor NOR4 (N8293, N8278, N995, N8168, N3367);
and AND2 (N8294, N8290, N3410);
nor NOR3 (N8295, N8293, N7502, N2036);
or OR2 (N8296, N8292, N7353);
or OR3 (N8297, N8294, N2906, N2185);
not NOT1 (N8298, N8284);
buf BUF1 (N8299, N8297);
not NOT1 (N8300, N8291);
nor NOR2 (N8301, N8287, N7256);
buf BUF1 (N8302, N8299);
nand NAND4 (N8303, N8301, N2932, N4422, N2414);
and AND3 (N8304, N8283, N3577, N1280);
xor XOR2 (N8305, N8303, N2172);
nor NOR4 (N8306, N8298, N7501, N6808, N5284);
nor NOR3 (N8307, N8296, N4009, N5626);
or OR4 (N8308, N8295, N3766, N3552, N3795);
xor XOR2 (N8309, N8306, N5694);
nor NOR4 (N8310, N8308, N5875, N2635, N7259);
nor NOR3 (N8311, N8302, N3747, N6671);
nand NAND3 (N8312, N8288, N2477, N6877);
nor NOR3 (N8313, N8305, N1115, N1390);
xor XOR2 (N8314, N8304, N6959);
xor XOR2 (N8315, N8309, N2937);
buf BUF1 (N8316, N8282);
not NOT1 (N8317, N8307);
nor NOR3 (N8318, N8300, N8115, N2762);
and AND2 (N8319, N8315, N3566);
not NOT1 (N8320, N8311);
xor XOR2 (N8321, N8317, N6823);
or OR2 (N8322, N8319, N4857);
xor XOR2 (N8323, N8310, N4695);
buf BUF1 (N8324, N8314);
not NOT1 (N8325, N8320);
or OR2 (N8326, N8322, N6489);
buf BUF1 (N8327, N8312);
or OR4 (N8328, N8316, N4918, N1282, N2465);
and AND3 (N8329, N8328, N3880, N5218);
not NOT1 (N8330, N8321);
nand NAND4 (N8331, N8324, N5444, N1012, N8036);
and AND2 (N8332, N8327, N2786);
xor XOR2 (N8333, N8331, N6777);
nand NAND3 (N8334, N8330, N7905, N1111);
and AND3 (N8335, N8289, N5499, N101);
buf BUF1 (N8336, N8326);
nand NAND3 (N8337, N8333, N4939, N191);
not NOT1 (N8338, N8325);
and AND2 (N8339, N8329, N5540);
or OR3 (N8340, N8332, N4934, N4474);
buf BUF1 (N8341, N8336);
and AND2 (N8342, N8337, N1292);
not NOT1 (N8343, N8339);
nor NOR4 (N8344, N8340, N4362, N4331, N1172);
nor NOR2 (N8345, N8343, N6112);
buf BUF1 (N8346, N8335);
not NOT1 (N8347, N8341);
buf BUF1 (N8348, N8338);
nand NAND3 (N8349, N8334, N706, N24);
nand NAND2 (N8350, N8342, N1707);
nor NOR4 (N8351, N8323, N3121, N3459, N2212);
nand NAND3 (N8352, N8345, N307, N2998);
buf BUF1 (N8353, N8318);
not NOT1 (N8354, N8352);
not NOT1 (N8355, N8346);
buf BUF1 (N8356, N8353);
nor NOR2 (N8357, N8351, N468);
nor NOR2 (N8358, N8313, N7608);
and AND4 (N8359, N8357, N2405, N7272, N2116);
buf BUF1 (N8360, N8355);
xor XOR2 (N8361, N8359, N3325);
or OR2 (N8362, N8350, N1285);
nand NAND4 (N8363, N8360, N2594, N4826, N2961);
nor NOR3 (N8364, N8361, N4935, N5622);
nand NAND2 (N8365, N8362, N1040);
and AND3 (N8366, N8354, N5850, N3534);
not NOT1 (N8367, N8344);
nor NOR2 (N8368, N8363, N6802);
xor XOR2 (N8369, N8368, N4717);
buf BUF1 (N8370, N8356);
buf BUF1 (N8371, N8358);
not NOT1 (N8372, N8364);
nor NOR3 (N8373, N8366, N5392, N6715);
nor NOR4 (N8374, N8347, N1825, N5504, N1110);
or OR3 (N8375, N8348, N6434, N8008);
and AND4 (N8376, N8371, N220, N6819, N6979);
xor XOR2 (N8377, N8372, N3412);
buf BUF1 (N8378, N8367);
not NOT1 (N8379, N8375);
buf BUF1 (N8380, N8379);
xor XOR2 (N8381, N8374, N1369);
not NOT1 (N8382, N8380);
nand NAND2 (N8383, N8377, N3961);
buf BUF1 (N8384, N8349);
and AND4 (N8385, N8383, N2176, N6303, N7357);
buf BUF1 (N8386, N8378);
nand NAND2 (N8387, N8381, N116);
not NOT1 (N8388, N8373);
or OR3 (N8389, N8369, N85, N2407);
nor NOR2 (N8390, N8386, N456);
nand NAND2 (N8391, N8387, N960);
not NOT1 (N8392, N8382);
nand NAND2 (N8393, N8388, N7218);
nand NAND2 (N8394, N8393, N7740);
buf BUF1 (N8395, N8391);
or OR4 (N8396, N8365, N3920, N1902, N1206);
or OR2 (N8397, N8384, N2007);
not NOT1 (N8398, N8390);
nand NAND2 (N8399, N8370, N4604);
and AND4 (N8400, N8389, N1664, N959, N7127);
nor NOR2 (N8401, N8395, N1483);
and AND3 (N8402, N8399, N5573, N808);
nor NOR2 (N8403, N8397, N5418);
nor NOR4 (N8404, N8385, N5182, N181, N4579);
nand NAND3 (N8405, N8401, N5394, N5553);
and AND3 (N8406, N8396, N623, N7570);
nand NAND3 (N8407, N8403, N1010, N4089);
or OR2 (N8408, N8407, N5023);
not NOT1 (N8409, N8406);
xor XOR2 (N8410, N8404, N8162);
buf BUF1 (N8411, N8400);
and AND2 (N8412, N8398, N4106);
buf BUF1 (N8413, N8410);
and AND4 (N8414, N8413, N3127, N2251, N6414);
nand NAND2 (N8415, N8405, N1789);
buf BUF1 (N8416, N8412);
and AND3 (N8417, N8376, N6877, N1925);
or OR2 (N8418, N8408, N2356);
xor XOR2 (N8419, N8402, N2829);
xor XOR2 (N8420, N8417, N4292);
or OR4 (N8421, N8419, N3035, N8054, N5429);
nor NOR2 (N8422, N8421, N4017);
nor NOR3 (N8423, N8394, N1097, N3968);
xor XOR2 (N8424, N8409, N1200);
or OR4 (N8425, N8420, N6653, N3464, N4803);
not NOT1 (N8426, N8414);
and AND4 (N8427, N8392, N6936, N8267, N4304);
nand NAND2 (N8428, N8415, N5907);
nor NOR3 (N8429, N8422, N1642, N7165);
and AND4 (N8430, N8418, N7160, N5176, N1833);
xor XOR2 (N8431, N8428, N1507);
and AND4 (N8432, N8430, N3305, N1588, N5767);
nand NAND2 (N8433, N8432, N7217);
nand NAND4 (N8434, N8429, N4442, N3407, N4554);
and AND3 (N8435, N8431, N7063, N7927);
xor XOR2 (N8436, N8416, N7209);
nor NOR2 (N8437, N8427, N3753);
buf BUF1 (N8438, N8425);
and AND4 (N8439, N8411, N2132, N5400, N5087);
buf BUF1 (N8440, N8439);
and AND4 (N8441, N8435, N3865, N7275, N7852);
xor XOR2 (N8442, N8441, N3004);
buf BUF1 (N8443, N8423);
buf BUF1 (N8444, N8442);
buf BUF1 (N8445, N8434);
or OR4 (N8446, N8433, N610, N5425, N4837);
nand NAND3 (N8447, N8436, N6606, N412);
or OR2 (N8448, N8440, N1937);
xor XOR2 (N8449, N8443, N4017);
or OR4 (N8450, N8448, N998, N5779, N6239);
nand NAND2 (N8451, N8426, N540);
buf BUF1 (N8452, N8447);
xor XOR2 (N8453, N8424, N6767);
nand NAND3 (N8454, N8444, N3742, N2709);
xor XOR2 (N8455, N8446, N2095);
xor XOR2 (N8456, N8453, N4694);
not NOT1 (N8457, N8445);
buf BUF1 (N8458, N8456);
and AND3 (N8459, N8438, N595, N2857);
nor NOR4 (N8460, N8459, N2281, N7434, N5776);
or OR3 (N8461, N8452, N8079, N960);
or OR3 (N8462, N8437, N4797, N6693);
nor NOR4 (N8463, N8454, N2236, N4164, N4613);
xor XOR2 (N8464, N8463, N705);
nand NAND3 (N8465, N8449, N4579, N1528);
buf BUF1 (N8466, N8465);
or OR4 (N8467, N8461, N4332, N8133, N5751);
or OR4 (N8468, N8450, N2188, N4131, N7926);
nand NAND4 (N8469, N8462, N8062, N1121, N4647);
xor XOR2 (N8470, N8460, N4213);
or OR4 (N8471, N8451, N6010, N7633, N4178);
nor NOR4 (N8472, N8469, N917, N1793, N1134);
or OR4 (N8473, N8458, N6120, N7774, N7086);
and AND4 (N8474, N8468, N5088, N4816, N4076);
and AND3 (N8475, N8470, N2294, N2547);
buf BUF1 (N8476, N8475);
and AND3 (N8477, N8464, N6264, N5427);
and AND4 (N8478, N8467, N5531, N3769, N6199);
or OR4 (N8479, N8466, N4003, N6014, N5706);
nand NAND3 (N8480, N8476, N4865, N1235);
not NOT1 (N8481, N8473);
nor NOR4 (N8482, N8480, N5242, N2682, N3548);
buf BUF1 (N8483, N8471);
nand NAND3 (N8484, N8482, N5107, N748);
nand NAND4 (N8485, N8472, N1934, N8034, N1947);
nand NAND2 (N8486, N8477, N3885);
nor NOR2 (N8487, N8455, N3846);
xor XOR2 (N8488, N8457, N3468);
buf BUF1 (N8489, N8485);
buf BUF1 (N8490, N8486);
or OR2 (N8491, N8479, N3756);
and AND3 (N8492, N8490, N4939, N34);
nand NAND3 (N8493, N8478, N80, N2195);
not NOT1 (N8494, N8493);
nor NOR3 (N8495, N8491, N7164, N1440);
buf BUF1 (N8496, N8484);
and AND3 (N8497, N8487, N4689, N2915);
buf BUF1 (N8498, N8483);
buf BUF1 (N8499, N8495);
nand NAND4 (N8500, N8492, N6233, N8018, N6126);
xor XOR2 (N8501, N8497, N1793);
nand NAND4 (N8502, N8481, N6727, N5939, N3090);
and AND3 (N8503, N8501, N7861, N3498);
buf BUF1 (N8504, N8494);
buf BUF1 (N8505, N8503);
nor NOR3 (N8506, N8499, N8030, N5117);
and AND2 (N8507, N8474, N7293);
or OR4 (N8508, N8498, N2228, N7496, N1376);
nor NOR2 (N8509, N8506, N7413);
or OR2 (N8510, N8489, N2765);
not NOT1 (N8511, N8510);
nand NAND2 (N8512, N8509, N1730);
buf BUF1 (N8513, N8488);
and AND2 (N8514, N8511, N2482);
not NOT1 (N8515, N8514);
xor XOR2 (N8516, N8504, N8459);
buf BUF1 (N8517, N8507);
xor XOR2 (N8518, N8515, N2029);
or OR4 (N8519, N8496, N6537, N3013, N7935);
and AND3 (N8520, N8512, N3312, N8282);
buf BUF1 (N8521, N8517);
nand NAND3 (N8522, N8519, N3311, N5548);
and AND3 (N8523, N8513, N3498, N4575);
and AND4 (N8524, N8522, N8153, N1624, N3845);
not NOT1 (N8525, N8500);
nor NOR4 (N8526, N8524, N5002, N7663, N3232);
not NOT1 (N8527, N8502);
buf BUF1 (N8528, N8516);
and AND4 (N8529, N8520, N6072, N1108, N1356);
nor NOR4 (N8530, N8505, N2336, N7550, N2182);
buf BUF1 (N8531, N8526);
xor XOR2 (N8532, N8531, N3704);
nand NAND2 (N8533, N8528, N2530);
xor XOR2 (N8534, N8527, N648);
nor NOR2 (N8535, N8532, N3443);
nand NAND4 (N8536, N8535, N4586, N3406, N4306);
buf BUF1 (N8537, N8534);
and AND3 (N8538, N8533, N7757, N2005);
nor NOR4 (N8539, N8537, N3895, N7709, N1026);
or OR2 (N8540, N8529, N4706);
nor NOR4 (N8541, N8540, N3247, N7167, N6311);
and AND3 (N8542, N8508, N7763, N3920);
or OR2 (N8543, N8521, N794);
or OR3 (N8544, N8523, N1103, N2999);
xor XOR2 (N8545, N8543, N7667);
or OR2 (N8546, N8545, N1929);
or OR4 (N8547, N8536, N3772, N3987, N6849);
not NOT1 (N8548, N8546);
and AND4 (N8549, N8518, N6420, N3951, N3543);
or OR3 (N8550, N8547, N627, N5200);
nand NAND2 (N8551, N8548, N4112);
nor NOR4 (N8552, N8549, N4456, N4351, N4410);
and AND4 (N8553, N8541, N3023, N8241, N1787);
nand NAND4 (N8554, N8538, N1791, N7523, N1549);
xor XOR2 (N8555, N8550, N535);
nand NAND3 (N8556, N8551, N3791, N4596);
xor XOR2 (N8557, N8544, N8058);
xor XOR2 (N8558, N8555, N76);
or OR2 (N8559, N8554, N5967);
nor NOR4 (N8560, N8552, N2745, N4199, N7834);
and AND2 (N8561, N8542, N1860);
xor XOR2 (N8562, N8559, N4608);
or OR2 (N8563, N8557, N599);
not NOT1 (N8564, N8553);
buf BUF1 (N8565, N8561);
nor NOR2 (N8566, N8558, N6299);
buf BUF1 (N8567, N8539);
and AND2 (N8568, N8564, N3184);
buf BUF1 (N8569, N8562);
buf BUF1 (N8570, N8560);
and AND2 (N8571, N8569, N420);
nand NAND2 (N8572, N8567, N3081);
nand NAND3 (N8573, N8566, N2228, N56);
nand NAND3 (N8574, N8525, N1394, N5393);
or OR3 (N8575, N8574, N7667, N6110);
nor NOR3 (N8576, N8572, N3834, N6299);
xor XOR2 (N8577, N8565, N478);
and AND2 (N8578, N8530, N2100);
or OR4 (N8579, N8576, N814, N1184, N6298);
not NOT1 (N8580, N8563);
not NOT1 (N8581, N8570);
or OR4 (N8582, N8577, N6974, N5902, N5909);
and AND3 (N8583, N8556, N5428, N5085);
xor XOR2 (N8584, N8575, N5468);
not NOT1 (N8585, N8573);
or OR4 (N8586, N8571, N3566, N3008, N5958);
and AND4 (N8587, N8582, N4951, N8207, N4295);
not NOT1 (N8588, N8568);
buf BUF1 (N8589, N8588);
nor NOR3 (N8590, N8586, N6917, N730);
nor NOR3 (N8591, N8590, N914, N4723);
not NOT1 (N8592, N8589);
xor XOR2 (N8593, N8580, N3755);
or OR4 (N8594, N8593, N5563, N1643, N6346);
buf BUF1 (N8595, N8584);
xor XOR2 (N8596, N8594, N7015);
or OR3 (N8597, N8591, N753, N7188);
nor NOR2 (N8598, N8596, N2226);
not NOT1 (N8599, N8578);
xor XOR2 (N8600, N8595, N3734);
xor XOR2 (N8601, N8583, N2239);
nand NAND2 (N8602, N8579, N2302);
xor XOR2 (N8603, N8602, N8447);
buf BUF1 (N8604, N8592);
xor XOR2 (N8605, N8603, N865);
and AND2 (N8606, N8599, N6673);
nand NAND2 (N8607, N8604, N4428);
and AND4 (N8608, N8601, N1802, N3526, N8020);
or OR2 (N8609, N8606, N363);
nand NAND4 (N8610, N8608, N355, N1606, N3617);
xor XOR2 (N8611, N8605, N314);
not NOT1 (N8612, N8607);
buf BUF1 (N8613, N8581);
buf BUF1 (N8614, N8610);
nand NAND3 (N8615, N8614, N1987, N3787);
not NOT1 (N8616, N8597);
buf BUF1 (N8617, N8615);
buf BUF1 (N8618, N8600);
or OR4 (N8619, N8587, N3836, N725, N6558);
or OR3 (N8620, N8618, N7293, N6153);
nor NOR2 (N8621, N8585, N6407);
xor XOR2 (N8622, N8621, N5235);
not NOT1 (N8623, N8617);
not NOT1 (N8624, N8623);
buf BUF1 (N8625, N8624);
and AND3 (N8626, N8613, N7241, N597);
nor NOR3 (N8627, N8609, N2676, N5668);
nor NOR3 (N8628, N8619, N3815, N6728);
nand NAND3 (N8629, N8628, N7317, N8486);
and AND3 (N8630, N8612, N6655, N5945);
and AND4 (N8631, N8622, N448, N890, N1957);
buf BUF1 (N8632, N8620);
buf BUF1 (N8633, N8598);
and AND2 (N8634, N8627, N5447);
nor NOR4 (N8635, N8611, N3516, N215, N1360);
or OR4 (N8636, N8616, N919, N5342, N5360);
buf BUF1 (N8637, N8635);
buf BUF1 (N8638, N8625);
nor NOR2 (N8639, N8634, N4076);
or OR4 (N8640, N8638, N2358, N1509, N1481);
not NOT1 (N8641, N8639);
not NOT1 (N8642, N8629);
nand NAND4 (N8643, N8626, N4319, N813, N1173);
and AND3 (N8644, N8636, N6343, N96);
nand NAND4 (N8645, N8644, N5832, N4891, N5523);
nor NOR4 (N8646, N8637, N241, N2151, N1571);
or OR3 (N8647, N8646, N7398, N888);
and AND2 (N8648, N8647, N1736);
xor XOR2 (N8649, N8642, N422);
and AND2 (N8650, N8632, N8584);
xor XOR2 (N8651, N8630, N665);
or OR3 (N8652, N8645, N6537, N7524);
nand NAND4 (N8653, N8641, N5431, N8373, N5272);
xor XOR2 (N8654, N8643, N492);
nand NAND2 (N8655, N8652, N6736);
or OR2 (N8656, N8631, N1625);
or OR2 (N8657, N8654, N3445);
nand NAND3 (N8658, N8633, N3300, N1304);
xor XOR2 (N8659, N8648, N5952);
buf BUF1 (N8660, N8657);
or OR3 (N8661, N8658, N4321, N2754);
buf BUF1 (N8662, N8650);
and AND4 (N8663, N8651, N5700, N4863, N3784);
and AND4 (N8664, N8659, N3182, N7645, N186);
xor XOR2 (N8665, N8656, N6047);
or OR4 (N8666, N8661, N5399, N3219, N6538);
not NOT1 (N8667, N8655);
or OR4 (N8668, N8663, N3167, N5122, N7165);
or OR3 (N8669, N8664, N4425, N2942);
nand NAND2 (N8670, N8669, N7649);
and AND4 (N8671, N8670, N8507, N2213, N3964);
buf BUF1 (N8672, N8660);
not NOT1 (N8673, N8662);
xor XOR2 (N8674, N8668, N8428);
buf BUF1 (N8675, N8674);
and AND2 (N8676, N8675, N4199);
or OR3 (N8677, N8671, N2400, N2404);
not NOT1 (N8678, N8649);
nor NOR4 (N8679, N8653, N444, N5362, N4805);
and AND3 (N8680, N8666, N2526, N7901);
or OR2 (N8681, N8673, N6008);
xor XOR2 (N8682, N8679, N5384);
and AND4 (N8683, N8678, N6200, N7132, N6006);
or OR4 (N8684, N8676, N6120, N6828, N167);
not NOT1 (N8685, N8681);
xor XOR2 (N8686, N8665, N3310);
nor NOR4 (N8687, N8684, N2672, N3620, N4853);
nand NAND2 (N8688, N8640, N6936);
nand NAND3 (N8689, N8682, N6712, N7262);
xor XOR2 (N8690, N8687, N4833);
and AND4 (N8691, N8686, N8238, N4096, N7422);
nor NOR2 (N8692, N8690, N3964);
nand NAND3 (N8693, N8688, N5831, N6485);
xor XOR2 (N8694, N8693, N5043);
buf BUF1 (N8695, N8672);
buf BUF1 (N8696, N8685);
xor XOR2 (N8697, N8696, N5276);
xor XOR2 (N8698, N8680, N7365);
nor NOR2 (N8699, N8695, N4141);
nor NOR3 (N8700, N8699, N3036, N7264);
not NOT1 (N8701, N8694);
nand NAND2 (N8702, N8683, N6523);
nand NAND3 (N8703, N8667, N7857, N5647);
nand NAND2 (N8704, N8700, N2374);
buf BUF1 (N8705, N8692);
xor XOR2 (N8706, N8677, N6566);
not NOT1 (N8707, N8702);
nor NOR4 (N8708, N8697, N2098, N6387, N4060);
or OR2 (N8709, N8706, N3786);
xor XOR2 (N8710, N8698, N1069);
or OR3 (N8711, N8691, N2696, N7419);
and AND2 (N8712, N8689, N5876);
and AND2 (N8713, N8711, N105);
xor XOR2 (N8714, N8704, N6917);
and AND3 (N8715, N8705, N5595, N3623);
nand NAND2 (N8716, N8712, N5949);
nand NAND3 (N8717, N8707, N6212, N6564);
not NOT1 (N8718, N8715);
or OR4 (N8719, N8710, N212, N243, N5788);
buf BUF1 (N8720, N8716);
xor XOR2 (N8721, N8714, N1846);
or OR4 (N8722, N8709, N370, N7080, N2941);
and AND3 (N8723, N8719, N6165, N4288);
buf BUF1 (N8724, N8708);
xor XOR2 (N8725, N8722, N7248);
nand NAND4 (N8726, N8713, N4478, N3167, N5696);
nand NAND3 (N8727, N8724, N7251, N5477);
or OR3 (N8728, N8717, N6454, N863);
xor XOR2 (N8729, N8721, N4739);
buf BUF1 (N8730, N8723);
nand NAND2 (N8731, N8730, N1493);
not NOT1 (N8732, N8718);
and AND3 (N8733, N8727, N5224, N3803);
or OR2 (N8734, N8732, N4740);
buf BUF1 (N8735, N8729);
and AND2 (N8736, N8701, N8310);
and AND2 (N8737, N8734, N7685);
xor XOR2 (N8738, N8703, N5776);
not NOT1 (N8739, N8731);
nor NOR2 (N8740, N8739, N1851);
and AND3 (N8741, N8733, N321, N8295);
xor XOR2 (N8742, N8728, N3840);
and AND3 (N8743, N8742, N428, N1178);
xor XOR2 (N8744, N8720, N2110);
nand NAND2 (N8745, N8735, N7179);
buf BUF1 (N8746, N8725);
xor XOR2 (N8747, N8741, N8602);
not NOT1 (N8748, N8745);
buf BUF1 (N8749, N8740);
nor NOR2 (N8750, N8726, N1206);
or OR4 (N8751, N8738, N238, N4474, N6771);
nand NAND2 (N8752, N8750, N2767);
buf BUF1 (N8753, N8752);
buf BUF1 (N8754, N8746);
nor NOR3 (N8755, N8749, N4079, N6467);
xor XOR2 (N8756, N8753, N945);
xor XOR2 (N8757, N8747, N7790);
nor NOR4 (N8758, N8744, N8198, N3734, N2060);
not NOT1 (N8759, N8748);
buf BUF1 (N8760, N8756);
nand NAND4 (N8761, N8759, N3664, N6481, N795);
xor XOR2 (N8762, N8736, N3519);
or OR2 (N8763, N8761, N3573);
buf BUF1 (N8764, N8737);
buf BUF1 (N8765, N8743);
nor NOR4 (N8766, N8754, N7780, N3081, N7401);
buf BUF1 (N8767, N8766);
buf BUF1 (N8768, N8755);
nor NOR2 (N8769, N8758, N2714);
xor XOR2 (N8770, N8765, N4115);
not NOT1 (N8771, N8757);
and AND3 (N8772, N8769, N3604, N1523);
buf BUF1 (N8773, N8763);
and AND3 (N8774, N8767, N1577, N5418);
and AND2 (N8775, N8770, N8197);
not NOT1 (N8776, N8772);
or OR2 (N8777, N8764, N6167);
xor XOR2 (N8778, N8776, N1160);
nand NAND3 (N8779, N8774, N895, N6705);
xor XOR2 (N8780, N8778, N3283);
nand NAND4 (N8781, N8760, N7038, N8315, N6313);
nor NOR4 (N8782, N8773, N4795, N8241, N2910);
not NOT1 (N8783, N8771);
xor XOR2 (N8784, N8782, N6095);
not NOT1 (N8785, N8751);
nor NOR4 (N8786, N8779, N1725, N6202, N5569);
and AND4 (N8787, N8783, N3955, N7663, N6897);
and AND4 (N8788, N8777, N2892, N5939, N5067);
buf BUF1 (N8789, N8762);
nor NOR3 (N8790, N8768, N8307, N5132);
and AND2 (N8791, N8784, N5939);
and AND2 (N8792, N8790, N195);
and AND3 (N8793, N8785, N1719, N8166);
nand NAND4 (N8794, N8786, N952, N7191, N3348);
and AND4 (N8795, N8793, N5645, N1952, N2625);
nor NOR3 (N8796, N8781, N8462, N1838);
and AND4 (N8797, N8775, N725, N7695, N8047);
and AND2 (N8798, N8789, N275);
xor XOR2 (N8799, N8798, N1710);
nor NOR3 (N8800, N8795, N1461, N8214);
nor NOR4 (N8801, N8800, N96, N7456, N2745);
not NOT1 (N8802, N8788);
xor XOR2 (N8803, N8801, N1758);
nor NOR4 (N8804, N8792, N7603, N7233, N4446);
nor NOR4 (N8805, N8787, N4218, N383, N3915);
xor XOR2 (N8806, N8791, N2597);
buf BUF1 (N8807, N8804);
and AND4 (N8808, N8797, N5492, N4902, N6138);
not NOT1 (N8809, N8780);
buf BUF1 (N8810, N8808);
buf BUF1 (N8811, N8803);
nor NOR3 (N8812, N8794, N8368, N3054);
buf BUF1 (N8813, N8812);
nor NOR4 (N8814, N8813, N4996, N4051, N4208);
buf BUF1 (N8815, N8814);
nand NAND3 (N8816, N8807, N4412, N5972);
or OR3 (N8817, N8815, N5255, N8430);
xor XOR2 (N8818, N8796, N413);
nor NOR3 (N8819, N8806, N5457, N6712);
xor XOR2 (N8820, N8810, N6837);
not NOT1 (N8821, N8820);
or OR4 (N8822, N8821, N266, N3706, N3781);
not NOT1 (N8823, N8817);
nor NOR2 (N8824, N8818, N7484);
and AND4 (N8825, N8802, N2575, N7572, N2666);
nand NAND2 (N8826, N8809, N6711);
and AND4 (N8827, N8822, N6138, N8227, N2636);
not NOT1 (N8828, N8823);
and AND3 (N8829, N8826, N4000, N1266);
xor XOR2 (N8830, N8824, N905);
or OR4 (N8831, N8829, N8518, N7207, N7832);
or OR4 (N8832, N8828, N1547, N4916, N1737);
not NOT1 (N8833, N8832);
nor NOR3 (N8834, N8799, N1886, N4191);
or OR4 (N8835, N8805, N1884, N884, N6985);
not NOT1 (N8836, N8833);
or OR4 (N8837, N8834, N6857, N5357, N7438);
and AND3 (N8838, N8819, N2773, N7304);
nor NOR4 (N8839, N8835, N4647, N7625, N2556);
not NOT1 (N8840, N8816);
buf BUF1 (N8841, N8838);
buf BUF1 (N8842, N8830);
xor XOR2 (N8843, N8836, N7556);
not NOT1 (N8844, N8841);
nor NOR3 (N8845, N8840, N8819, N1287);
xor XOR2 (N8846, N8827, N690);
or OR4 (N8847, N8825, N6513, N1070, N5929);
xor XOR2 (N8848, N8837, N5195);
xor XOR2 (N8849, N8811, N6210);
not NOT1 (N8850, N8846);
nor NOR2 (N8851, N8849, N6848);
not NOT1 (N8852, N8850);
and AND2 (N8853, N8851, N3811);
xor XOR2 (N8854, N8842, N542);
and AND3 (N8855, N8848, N403, N2950);
buf BUF1 (N8856, N8839);
or OR2 (N8857, N8856, N5413);
nand NAND2 (N8858, N8844, N6479);
not NOT1 (N8859, N8852);
xor XOR2 (N8860, N8853, N52);
or OR3 (N8861, N8847, N6253, N2626);
and AND2 (N8862, N8843, N2772);
and AND3 (N8863, N8831, N337, N1334);
and AND2 (N8864, N8855, N7124);
or OR3 (N8865, N8860, N8100, N723);
nor NOR4 (N8866, N8863, N268, N5207, N8692);
nand NAND3 (N8867, N8857, N779, N8591);
not NOT1 (N8868, N8859);
nor NOR4 (N8869, N8854, N472, N2283, N2557);
and AND2 (N8870, N8869, N3187);
nor NOR2 (N8871, N8868, N4097);
xor XOR2 (N8872, N8864, N4975);
not NOT1 (N8873, N8862);
and AND2 (N8874, N8873, N4337);
nand NAND2 (N8875, N8870, N143);
nand NAND3 (N8876, N8866, N2129, N3462);
nand NAND2 (N8877, N8876, N1229);
nand NAND4 (N8878, N8871, N1651, N846, N1847);
buf BUF1 (N8879, N8858);
xor XOR2 (N8880, N8861, N5388);
or OR2 (N8881, N8867, N6672);
not NOT1 (N8882, N8845);
not NOT1 (N8883, N8872);
xor XOR2 (N8884, N8874, N2736);
nand NAND2 (N8885, N8883, N7660);
nand NAND3 (N8886, N8875, N1700, N869);
xor XOR2 (N8887, N8880, N6698);
not NOT1 (N8888, N8882);
not NOT1 (N8889, N8878);
xor XOR2 (N8890, N8877, N6127);
xor XOR2 (N8891, N8889, N7227);
or OR3 (N8892, N8886, N779, N7248);
or OR3 (N8893, N8885, N4722, N4757);
nand NAND4 (N8894, N8893, N1716, N3634, N2923);
nor NOR4 (N8895, N8865, N1233, N7396, N5562);
not NOT1 (N8896, N8895);
not NOT1 (N8897, N8891);
not NOT1 (N8898, N8887);
and AND4 (N8899, N8890, N239, N4318, N1967);
and AND2 (N8900, N8897, N6363);
and AND4 (N8901, N8879, N2956, N3290, N3094);
and AND4 (N8902, N8898, N5971, N1195, N5841);
nand NAND2 (N8903, N8902, N1293);
buf BUF1 (N8904, N8884);
buf BUF1 (N8905, N8881);
nor NOR3 (N8906, N8892, N7840, N5642);
nand NAND3 (N8907, N8894, N2322, N6028);
not NOT1 (N8908, N8896);
or OR2 (N8909, N8907, N3949);
or OR3 (N8910, N8909, N8403, N7508);
nor NOR3 (N8911, N8906, N6440, N1474);
or OR2 (N8912, N8903, N6814);
nand NAND2 (N8913, N8911, N7322);
not NOT1 (N8914, N8908);
or OR2 (N8915, N8913, N7690);
or OR3 (N8916, N8904, N8105, N2822);
or OR2 (N8917, N8888, N1184);
nor NOR4 (N8918, N8917, N6663, N2737, N5393);
xor XOR2 (N8919, N8910, N885);
nor NOR3 (N8920, N8918, N8650, N7450);
nor NOR3 (N8921, N8915, N89, N6617);
and AND4 (N8922, N8914, N5625, N2310, N8265);
not NOT1 (N8923, N8912);
and AND4 (N8924, N8900, N3380, N6793, N5349);
and AND2 (N8925, N8919, N1507);
xor XOR2 (N8926, N8924, N5227);
nor NOR4 (N8927, N8905, N8827, N800, N2842);
not NOT1 (N8928, N8916);
xor XOR2 (N8929, N8920, N7601);
xor XOR2 (N8930, N8923, N3951);
nand NAND4 (N8931, N8927, N809, N7510, N969);
or OR3 (N8932, N8928, N4372, N7821);
buf BUF1 (N8933, N8925);
not NOT1 (N8934, N8932);
and AND2 (N8935, N8922, N6168);
nand NAND3 (N8936, N8929, N3053, N1909);
not NOT1 (N8937, N8921);
or OR3 (N8938, N8926, N5822, N7634);
not NOT1 (N8939, N8901);
and AND3 (N8940, N8934, N8635, N6580);
nand NAND4 (N8941, N8935, N1653, N6280, N5158);
and AND4 (N8942, N8938, N2490, N6358, N4216);
xor XOR2 (N8943, N8936, N756);
nor NOR3 (N8944, N8939, N5078, N475);
not NOT1 (N8945, N8944);
nor NOR3 (N8946, N8933, N5386, N2602);
not NOT1 (N8947, N8899);
and AND4 (N8948, N8930, N216, N1485, N5790);
nand NAND2 (N8949, N8947, N3416);
and AND4 (N8950, N8931, N8307, N6962, N8427);
not NOT1 (N8951, N8943);
not NOT1 (N8952, N8940);
nor NOR2 (N8953, N8948, N7916);
and AND2 (N8954, N8942, N3226);
buf BUF1 (N8955, N8950);
and AND3 (N8956, N8937, N3409, N1658);
xor XOR2 (N8957, N8956, N3713);
or OR4 (N8958, N8949, N7834, N6856, N1212);
buf BUF1 (N8959, N8954);
not NOT1 (N8960, N8945);
or OR3 (N8961, N8957, N89, N3024);
or OR2 (N8962, N8959, N8413);
xor XOR2 (N8963, N8958, N7014);
nor NOR2 (N8964, N8953, N3276);
or OR2 (N8965, N8951, N8516);
not NOT1 (N8966, N8961);
xor XOR2 (N8967, N8960, N1050);
not NOT1 (N8968, N8955);
xor XOR2 (N8969, N8964, N2862);
nand NAND2 (N8970, N8941, N303);
nor NOR4 (N8971, N8952, N559, N1825, N4129);
nand NAND2 (N8972, N8963, N1207);
or OR3 (N8973, N8972, N2766, N2314);
or OR2 (N8974, N8970, N4503);
buf BUF1 (N8975, N8968);
xor XOR2 (N8976, N8974, N4754);
or OR3 (N8977, N8965, N8771, N231);
nand NAND3 (N8978, N8967, N591, N6);
buf BUF1 (N8979, N8962);
xor XOR2 (N8980, N8969, N6655);
not NOT1 (N8981, N8971);
nand NAND3 (N8982, N8975, N3895, N7156);
and AND3 (N8983, N8966, N7902, N551);
buf BUF1 (N8984, N8980);
buf BUF1 (N8985, N8982);
and AND2 (N8986, N8977, N973);
buf BUF1 (N8987, N8976);
or OR3 (N8988, N8973, N7438, N370);
buf BUF1 (N8989, N8988);
or OR3 (N8990, N8983, N365, N6700);
nand NAND3 (N8991, N8986, N5735, N5650);
xor XOR2 (N8992, N8985, N2806);
nand NAND4 (N8993, N8987, N6122, N8235, N6834);
nor NOR4 (N8994, N8946, N3029, N632, N8663);
xor XOR2 (N8995, N8989, N4759);
or OR4 (N8996, N8994, N4330, N5806, N566);
nor NOR3 (N8997, N8991, N6395, N128);
xor XOR2 (N8998, N8996, N1801);
or OR3 (N8999, N8978, N4266, N2929);
buf BUF1 (N9000, N8981);
buf BUF1 (N9001, N8990);
or OR3 (N9002, N8993, N5338, N6067);
nand NAND4 (N9003, N8992, N5788, N5911, N4846);
nand NAND3 (N9004, N8998, N8370, N154);
nor NOR2 (N9005, N9004, N4188);
xor XOR2 (N9006, N8979, N3299);
buf BUF1 (N9007, N9006);
and AND4 (N9008, N9005, N59, N1096, N7958);
not NOT1 (N9009, N8995);
nor NOR2 (N9010, N9008, N3155);
and AND2 (N9011, N8999, N8095);
nand NAND4 (N9012, N9010, N7828, N1326, N4910);
not NOT1 (N9013, N9009);
or OR2 (N9014, N9011, N8729);
or OR4 (N9015, N9012, N4061, N1368, N4294);
and AND4 (N9016, N9001, N4255, N7801, N4288);
xor XOR2 (N9017, N9013, N4548);
xor XOR2 (N9018, N9015, N4836);
buf BUF1 (N9019, N9002);
buf BUF1 (N9020, N9003);
and AND4 (N9021, N9020, N2005, N2332, N256);
nor NOR3 (N9022, N8984, N2683, N8249);
not NOT1 (N9023, N9022);
and AND3 (N9024, N9021, N440, N728);
not NOT1 (N9025, N9023);
and AND4 (N9026, N8997, N1467, N5431, N2312);
or OR4 (N9027, N9014, N4591, N2430, N4808);
nor NOR3 (N9028, N9025, N298, N1669);
and AND4 (N9029, N9007, N3220, N7269, N6698);
nor NOR3 (N9030, N9000, N7396, N6024);
nand NAND2 (N9031, N9016, N3910);
nor NOR2 (N9032, N9030, N8758);
not NOT1 (N9033, N9029);
and AND2 (N9034, N9017, N367);
and AND3 (N9035, N9018, N1446, N1212);
or OR4 (N9036, N9027, N5340, N6865, N3599);
xor XOR2 (N9037, N9035, N1528);
and AND4 (N9038, N9032, N7081, N3807, N5832);
and AND4 (N9039, N9034, N2302, N3055, N8656);
and AND4 (N9040, N9037, N8915, N7402, N8251);
nor NOR2 (N9041, N9031, N5308);
xor XOR2 (N9042, N9019, N5038);
not NOT1 (N9043, N9040);
nor NOR2 (N9044, N9038, N2901);
and AND4 (N9045, N9024, N1533, N4325, N8754);
not NOT1 (N9046, N9039);
or OR3 (N9047, N9036, N6995, N8353);
not NOT1 (N9048, N9047);
xor XOR2 (N9049, N9041, N5048);
xor XOR2 (N9050, N9045, N3547);
nand NAND2 (N9051, N9049, N7968);
buf BUF1 (N9052, N9033);
nand NAND2 (N9053, N9042, N8013);
and AND4 (N9054, N9043, N7444, N8012, N5709);
not NOT1 (N9055, N9028);
buf BUF1 (N9056, N9044);
not NOT1 (N9057, N9048);
nand NAND3 (N9058, N9026, N7095, N5446);
or OR4 (N9059, N9055, N1480, N2120, N2405);
and AND3 (N9060, N9054, N4766, N17);
or OR3 (N9061, N9060, N4648, N1687);
nand NAND4 (N9062, N9050, N3288, N5092, N3320);
and AND4 (N9063, N9051, N3447, N7639, N4863);
xor XOR2 (N9064, N9046, N8706);
nand NAND2 (N9065, N9064, N1093);
nand NAND4 (N9066, N9063, N6237, N5563, N5665);
buf BUF1 (N9067, N9058);
xor XOR2 (N9068, N9059, N3494);
or OR4 (N9069, N9062, N8594, N7264, N667);
buf BUF1 (N9070, N9069);
or OR3 (N9071, N9066, N1890, N6291);
not NOT1 (N9072, N9067);
and AND2 (N9073, N9072, N635);
nor NOR3 (N9074, N9073, N3337, N5146);
not NOT1 (N9075, N9053);
xor XOR2 (N9076, N9074, N4927);
and AND3 (N9077, N9070, N880, N8586);
nor NOR3 (N9078, N9056, N2605, N7405);
nor NOR4 (N9079, N9061, N448, N3032, N6083);
nor NOR4 (N9080, N9079, N4801, N8804, N5812);
nand NAND2 (N9081, N9077, N4852);
buf BUF1 (N9082, N9071);
nor NOR4 (N9083, N9065, N1324, N2934, N8565);
or OR3 (N9084, N9078, N3599, N5752);
buf BUF1 (N9085, N9084);
or OR3 (N9086, N9085, N2845, N654);
and AND4 (N9087, N9057, N1600, N7405, N7002);
not NOT1 (N9088, N9081);
nand NAND4 (N9089, N9076, N5655, N8771, N8052);
and AND2 (N9090, N9086, N7102);
xor XOR2 (N9091, N9075, N8338);
and AND3 (N9092, N9082, N5290, N1899);
or OR2 (N9093, N9092, N7271);
xor XOR2 (N9094, N9091, N8507);
xor XOR2 (N9095, N9093, N5092);
or OR3 (N9096, N9068, N6386, N6466);
nand NAND2 (N9097, N9083, N8737);
xor XOR2 (N9098, N9088, N2144);
and AND3 (N9099, N9097, N2168, N3807);
and AND3 (N9100, N9094, N1357, N8490);
nand NAND2 (N9101, N9087, N3629);
nand NAND3 (N9102, N9098, N3204, N7946);
nand NAND3 (N9103, N9089, N9028, N689);
xor XOR2 (N9104, N9096, N9058);
and AND2 (N9105, N9099, N1371);
xor XOR2 (N9106, N9103, N2833);
and AND4 (N9107, N9105, N4347, N3306, N4613);
and AND4 (N9108, N9080, N2390, N8914, N8746);
buf BUF1 (N9109, N9102);
and AND4 (N9110, N9108, N1865, N1586, N3472);
nand NAND4 (N9111, N9052, N3728, N4692, N5349);
and AND4 (N9112, N9100, N3267, N8182, N8717);
buf BUF1 (N9113, N9106);
xor XOR2 (N9114, N9109, N7428);
buf BUF1 (N9115, N9112);
or OR4 (N9116, N9090, N6474, N451, N9039);
not NOT1 (N9117, N9107);
nand NAND4 (N9118, N9113, N1808, N3040, N3631);
nor NOR2 (N9119, N9101, N411);
or OR2 (N9120, N9104, N349);
and AND2 (N9121, N9116, N645);
nor NOR2 (N9122, N9118, N8276);
not NOT1 (N9123, N9119);
not NOT1 (N9124, N9115);
xor XOR2 (N9125, N9117, N3318);
nand NAND3 (N9126, N9095, N2806, N7440);
not NOT1 (N9127, N9114);
nor NOR2 (N9128, N9111, N4724);
and AND2 (N9129, N9121, N6015);
nor NOR2 (N9130, N9126, N2939);
xor XOR2 (N9131, N9124, N5556);
and AND2 (N9132, N9128, N7122);
and AND2 (N9133, N9130, N3200);
and AND2 (N9134, N9131, N8654);
nor NOR2 (N9135, N9122, N238);
xor XOR2 (N9136, N9132, N8847);
buf BUF1 (N9137, N9125);
xor XOR2 (N9138, N9134, N1827);
nor NOR2 (N9139, N9129, N3431);
or OR2 (N9140, N9133, N1277);
not NOT1 (N9141, N9120);
xor XOR2 (N9142, N9127, N2812);
xor XOR2 (N9143, N9135, N5163);
xor XOR2 (N9144, N9140, N5657);
xor XOR2 (N9145, N9123, N6552);
and AND3 (N9146, N9141, N7387, N6263);
or OR4 (N9147, N9143, N6157, N340, N6171);
nand NAND3 (N9148, N9142, N8597, N5897);
xor XOR2 (N9149, N9148, N5797);
or OR4 (N9150, N9136, N2650, N5314, N693);
buf BUF1 (N9151, N9137);
not NOT1 (N9152, N9151);
nand NAND3 (N9153, N9145, N9036, N8579);
buf BUF1 (N9154, N9152);
nand NAND3 (N9155, N9144, N5833, N8392);
nand NAND3 (N9156, N9154, N4847, N1787);
xor XOR2 (N9157, N9138, N4682);
xor XOR2 (N9158, N9155, N6404);
buf BUF1 (N9159, N9153);
nor NOR2 (N9160, N9156, N4619);
xor XOR2 (N9161, N9149, N6157);
buf BUF1 (N9162, N9157);
buf BUF1 (N9163, N9158);
nand NAND2 (N9164, N9147, N2765);
nor NOR4 (N9165, N9164, N4992, N7103, N8116);
not NOT1 (N9166, N9139);
buf BUF1 (N9167, N9160);
xor XOR2 (N9168, N9161, N2049);
nand NAND4 (N9169, N9168, N515, N2318, N417);
nor NOR3 (N9170, N9162, N4763, N2446);
or OR2 (N9171, N9163, N7215);
not NOT1 (N9172, N9170);
nor NOR2 (N9173, N9146, N7951);
nand NAND4 (N9174, N9159, N8636, N1545, N8905);
nor NOR2 (N9175, N9169, N7862);
buf BUF1 (N9176, N9150);
xor XOR2 (N9177, N9176, N3697);
nand NAND4 (N9178, N9165, N8964, N6607, N784);
nor NOR4 (N9179, N9175, N6996, N7247, N5906);
not NOT1 (N9180, N9171);
not NOT1 (N9181, N9166);
not NOT1 (N9182, N9173);
xor XOR2 (N9183, N9182, N625);
or OR4 (N9184, N9180, N2754, N7560, N6291);
nand NAND2 (N9185, N9172, N2446);
and AND2 (N9186, N9184, N2043);
and AND3 (N9187, N9178, N7844, N2373);
buf BUF1 (N9188, N9187);
not NOT1 (N9189, N9110);
or OR2 (N9190, N9181, N1997);
buf BUF1 (N9191, N9183);
nand NAND4 (N9192, N9167, N3076, N6726, N3084);
nand NAND3 (N9193, N9188, N6930, N8309);
or OR2 (N9194, N9190, N4743);
not NOT1 (N9195, N9191);
xor XOR2 (N9196, N9185, N7831);
buf BUF1 (N9197, N9196);
not NOT1 (N9198, N9179);
nand NAND3 (N9199, N9174, N3185, N7190);
and AND2 (N9200, N9186, N4669);
xor XOR2 (N9201, N9197, N110);
and AND2 (N9202, N9193, N7588);
or OR2 (N9203, N9195, N829);
nor NOR2 (N9204, N9189, N4511);
nor NOR4 (N9205, N9198, N207, N5491, N5791);
nor NOR3 (N9206, N9204, N599, N3366);
nand NAND2 (N9207, N9177, N5199);
or OR3 (N9208, N9207, N4078, N6207);
nand NAND4 (N9209, N9192, N90, N4241, N3606);
and AND4 (N9210, N9200, N276, N2134, N2003);
or OR2 (N9211, N9205, N4938);
buf BUF1 (N9212, N9208);
nand NAND2 (N9213, N9202, N5580);
xor XOR2 (N9214, N9199, N8895);
and AND2 (N9215, N9213, N2970);
nor NOR3 (N9216, N9203, N2050, N9063);
or OR2 (N9217, N9201, N8375);
xor XOR2 (N9218, N9211, N5302);
nand NAND3 (N9219, N9209, N7098, N329);
buf BUF1 (N9220, N9212);
or OR3 (N9221, N9215, N604, N4770);
xor XOR2 (N9222, N9219, N5648);
and AND2 (N9223, N9218, N6213);
nor NOR3 (N9224, N9194, N8178, N4021);
buf BUF1 (N9225, N9221);
and AND2 (N9226, N9214, N2471);
and AND2 (N9227, N9216, N4109);
and AND2 (N9228, N9224, N4705);
and AND3 (N9229, N9210, N8522, N5756);
nand NAND2 (N9230, N9223, N921);
xor XOR2 (N9231, N9206, N3370);
nor NOR2 (N9232, N9217, N7302);
and AND3 (N9233, N9228, N8765, N5220);
nand NAND3 (N9234, N9233, N2818, N4457);
or OR4 (N9235, N9222, N2490, N9101, N2126);
not NOT1 (N9236, N9232);
not NOT1 (N9237, N9231);
nand NAND4 (N9238, N9236, N8106, N6252, N63);
and AND2 (N9239, N9235, N4498);
and AND3 (N9240, N9239, N312, N2064);
xor XOR2 (N9241, N9225, N7437);
or OR3 (N9242, N9226, N5650, N3452);
buf BUF1 (N9243, N9227);
not NOT1 (N9244, N9243);
buf BUF1 (N9245, N9229);
or OR2 (N9246, N9220, N5437);
nor NOR2 (N9247, N9246, N2154);
and AND3 (N9248, N9238, N1984, N8514);
nand NAND4 (N9249, N9241, N6363, N7045, N6653);
not NOT1 (N9250, N9234);
and AND2 (N9251, N9249, N4847);
xor XOR2 (N9252, N9247, N4227);
and AND4 (N9253, N9252, N1270, N5733, N6076);
nor NOR2 (N9254, N9248, N8950);
xor XOR2 (N9255, N9250, N7284);
buf BUF1 (N9256, N9253);
nand NAND3 (N9257, N9255, N1841, N483);
or OR4 (N9258, N9237, N8292, N9184, N6474);
nand NAND2 (N9259, N9242, N6100);
nor NOR2 (N9260, N9256, N6911);
buf BUF1 (N9261, N9245);
xor XOR2 (N9262, N9240, N441);
nand NAND4 (N9263, N9257, N3066, N3506, N8243);
nor NOR4 (N9264, N9254, N4336, N5345, N39);
or OR3 (N9265, N9260, N3701, N8440);
nor NOR2 (N9266, N9259, N1956);
nand NAND2 (N9267, N9265, N7839);
and AND3 (N9268, N9263, N7768, N7320);
nand NAND3 (N9269, N9264, N2080, N1122);
not NOT1 (N9270, N9251);
xor XOR2 (N9271, N9262, N4191);
nand NAND2 (N9272, N9267, N6886);
xor XOR2 (N9273, N9271, N5927);
not NOT1 (N9274, N9230);
nor NOR2 (N9275, N9244, N4328);
xor XOR2 (N9276, N9275, N2547);
buf BUF1 (N9277, N9258);
nand NAND2 (N9278, N9277, N2252);
xor XOR2 (N9279, N9266, N5917);
or OR4 (N9280, N9272, N7168, N3791, N5948);
buf BUF1 (N9281, N9278);
nor NOR3 (N9282, N9261, N656, N7312);
buf BUF1 (N9283, N9274);
and AND4 (N9284, N9283, N6408, N6345, N6091);
or OR3 (N9285, N9279, N3885, N1671);
nor NOR3 (N9286, N9273, N7205, N6230);
not NOT1 (N9287, N9268);
xor XOR2 (N9288, N9285, N7916);
not NOT1 (N9289, N9287);
or OR4 (N9290, N9281, N2298, N1598, N126);
and AND2 (N9291, N9282, N6862);
buf BUF1 (N9292, N9270);
and AND4 (N9293, N9292, N3440, N805, N8286);
or OR3 (N9294, N9276, N1245, N204);
xor XOR2 (N9295, N9291, N4241);
not NOT1 (N9296, N9295);
nor NOR3 (N9297, N9296, N6181, N117);
nand NAND3 (N9298, N9280, N4806, N4500);
nand NAND4 (N9299, N9290, N8297, N2490, N2730);
not NOT1 (N9300, N9293);
not NOT1 (N9301, N9288);
and AND4 (N9302, N9300, N4002, N3680, N1991);
nand NAND4 (N9303, N9298, N6479, N7960, N1336);
nand NAND2 (N9304, N9269, N5095);
buf BUF1 (N9305, N9303);
and AND4 (N9306, N9284, N1348, N7420, N7261);
buf BUF1 (N9307, N9294);
not NOT1 (N9308, N9286);
xor XOR2 (N9309, N9302, N7927);
xor XOR2 (N9310, N9289, N4344);
buf BUF1 (N9311, N9309);
xor XOR2 (N9312, N9299, N8845);
buf BUF1 (N9313, N9307);
nand NAND2 (N9314, N9313, N8514);
nor NOR3 (N9315, N9305, N1373, N6304);
or OR3 (N9316, N9297, N3889, N2587);
buf BUF1 (N9317, N9301);
nand NAND2 (N9318, N9304, N8290);
buf BUF1 (N9319, N9318);
not NOT1 (N9320, N9314);
buf BUF1 (N9321, N9317);
xor XOR2 (N9322, N9316, N358);
xor XOR2 (N9323, N9320, N2542);
xor XOR2 (N9324, N9315, N3752);
and AND2 (N9325, N9323, N6728);
buf BUF1 (N9326, N9324);
buf BUF1 (N9327, N9319);
and AND4 (N9328, N9311, N9167, N7834, N7924);
and AND4 (N9329, N9322, N3765, N5463, N2274);
buf BUF1 (N9330, N9325);
nor NOR3 (N9331, N9330, N7416, N2249);
or OR3 (N9332, N9312, N1458, N6562);
and AND3 (N9333, N9306, N4837, N6595);
or OR2 (N9334, N9332, N6954);
or OR2 (N9335, N9329, N5723);
nand NAND2 (N9336, N9335, N409);
buf BUF1 (N9337, N9333);
not NOT1 (N9338, N9337);
nor NOR3 (N9339, N9310, N1733, N3464);
buf BUF1 (N9340, N9326);
or OR2 (N9341, N9308, N7504);
nand NAND3 (N9342, N9321, N6493, N7801);
buf BUF1 (N9343, N9339);
and AND3 (N9344, N9343, N5593, N4604);
not NOT1 (N9345, N9342);
xor XOR2 (N9346, N9344, N2458);
not NOT1 (N9347, N9336);
nand NAND2 (N9348, N9347, N5627);
buf BUF1 (N9349, N9331);
buf BUF1 (N9350, N9348);
not NOT1 (N9351, N9328);
xor XOR2 (N9352, N9341, N5803);
buf BUF1 (N9353, N9340);
xor XOR2 (N9354, N9327, N8595);
not NOT1 (N9355, N9334);
nand NAND4 (N9356, N9352, N7913, N4599, N1330);
or OR2 (N9357, N9345, N105);
and AND3 (N9358, N9353, N4283, N3416);
nand NAND4 (N9359, N9355, N6481, N7690, N141);
nand NAND4 (N9360, N9359, N8426, N6228, N7106);
or OR3 (N9361, N9354, N3874, N1203);
or OR3 (N9362, N9356, N1798, N3125);
nand NAND3 (N9363, N9349, N1702, N2122);
and AND3 (N9364, N9361, N5815, N2388);
or OR2 (N9365, N9350, N2997);
buf BUF1 (N9366, N9346);
and AND3 (N9367, N9363, N2038, N2464);
buf BUF1 (N9368, N9364);
and AND2 (N9369, N9366, N6498);
or OR3 (N9370, N9358, N2997, N4696);
or OR4 (N9371, N9351, N8269, N7106, N6496);
or OR2 (N9372, N9370, N223);
buf BUF1 (N9373, N9367);
nand NAND4 (N9374, N9373, N5820, N4804, N5293);
nand NAND3 (N9375, N9374, N1991, N4247);
not NOT1 (N9376, N9360);
xor XOR2 (N9377, N9338, N2898);
nand NAND3 (N9378, N9377, N2048, N6520);
nand NAND3 (N9379, N9375, N9123, N8502);
and AND4 (N9380, N9378, N1457, N6754, N8325);
not NOT1 (N9381, N9371);
not NOT1 (N9382, N9380);
or OR4 (N9383, N9357, N8859, N4643, N8801);
not NOT1 (N9384, N9379);
nor NOR3 (N9385, N9376, N1766, N7054);
xor XOR2 (N9386, N9369, N7070);
xor XOR2 (N9387, N9362, N146);
and AND4 (N9388, N9382, N5999, N1277, N7205);
not NOT1 (N9389, N9388);
buf BUF1 (N9390, N9387);
not NOT1 (N9391, N9386);
xor XOR2 (N9392, N9383, N75);
or OR3 (N9393, N9384, N2001, N7864);
buf BUF1 (N9394, N9393);
xor XOR2 (N9395, N9381, N6058);
or OR4 (N9396, N9365, N7183, N6983, N2943);
or OR3 (N9397, N9368, N950, N1795);
xor XOR2 (N9398, N9397, N4225);
nor NOR4 (N9399, N9389, N2552, N4966, N3384);
xor XOR2 (N9400, N9372, N3925);
nand NAND2 (N9401, N9400, N5375);
not NOT1 (N9402, N9401);
buf BUF1 (N9403, N9385);
nor NOR2 (N9404, N9403, N5907);
nor NOR2 (N9405, N9396, N3089);
or OR2 (N9406, N9404, N805);
or OR4 (N9407, N9392, N1856, N256, N1949);
not NOT1 (N9408, N9399);
xor XOR2 (N9409, N9394, N357);
nor NOR4 (N9410, N9407, N9381, N2552, N4250);
nand NAND3 (N9411, N9405, N3801, N22);
and AND3 (N9412, N9410, N1075, N8893);
and AND4 (N9413, N9409, N5263, N6470, N936);
xor XOR2 (N9414, N9390, N8696);
and AND4 (N9415, N9406, N472, N7979, N4052);
xor XOR2 (N9416, N9391, N289);
xor XOR2 (N9417, N9415, N7135);
buf BUF1 (N9418, N9413);
not NOT1 (N9419, N9418);
or OR2 (N9420, N9419, N2404);
and AND4 (N9421, N9420, N5720, N3226, N5108);
not NOT1 (N9422, N9395);
nand NAND4 (N9423, N9421, N564, N1988, N604);
xor XOR2 (N9424, N9414, N4361);
and AND2 (N9425, N9423, N6453);
or OR4 (N9426, N9424, N5046, N9265, N8288);
nand NAND3 (N9427, N9422, N860, N7929);
and AND3 (N9428, N9408, N6898, N387);
xor XOR2 (N9429, N9425, N1790);
and AND2 (N9430, N9398, N4809);
nand NAND3 (N9431, N9429, N8453, N6168);
and AND3 (N9432, N9411, N3070, N7176);
nor NOR2 (N9433, N9402, N2394);
buf BUF1 (N9434, N9412);
nor NOR3 (N9435, N9432, N1233, N3377);
or OR2 (N9436, N9416, N1278);
buf BUF1 (N9437, N9427);
xor XOR2 (N9438, N9430, N9076);
nand NAND2 (N9439, N9435, N6256);
xor XOR2 (N9440, N9434, N8547);
and AND3 (N9441, N9426, N4664, N2651);
nor NOR2 (N9442, N9433, N5092);
not NOT1 (N9443, N9441);
xor XOR2 (N9444, N9428, N6726);
or OR2 (N9445, N9439, N5202);
xor XOR2 (N9446, N9442, N936);
or OR4 (N9447, N9443, N6562, N2183, N2901);
nor NOR3 (N9448, N9431, N8328, N7916);
buf BUF1 (N9449, N9436);
not NOT1 (N9450, N9449);
buf BUF1 (N9451, N9437);
buf BUF1 (N9452, N9447);
xor XOR2 (N9453, N9438, N3127);
buf BUF1 (N9454, N9448);
nor NOR3 (N9455, N9440, N8205, N1155);
not NOT1 (N9456, N9417);
or OR3 (N9457, N9446, N534, N7485);
not NOT1 (N9458, N9454);
nor NOR3 (N9459, N9458, N2584, N4328);
buf BUF1 (N9460, N9450);
nor NOR2 (N9461, N9453, N5221);
nand NAND3 (N9462, N9444, N7305, N2463);
not NOT1 (N9463, N9462);
buf BUF1 (N9464, N9445);
and AND3 (N9465, N9457, N676, N2739);
buf BUF1 (N9466, N9456);
buf BUF1 (N9467, N9459);
xor XOR2 (N9468, N9461, N7825);
nand NAND4 (N9469, N9460, N8926, N2800, N3715);
nor NOR4 (N9470, N9467, N9441, N6980, N2377);
nand NAND3 (N9471, N9452, N1380, N8098);
or OR4 (N9472, N9465, N7929, N5170, N5651);
not NOT1 (N9473, N9468);
xor XOR2 (N9474, N9472, N6985);
nor NOR2 (N9475, N9451, N886);
buf BUF1 (N9476, N9463);
xor XOR2 (N9477, N9455, N3938);
or OR4 (N9478, N9473, N5430, N3991, N3903);
xor XOR2 (N9479, N9475, N8163);
not NOT1 (N9480, N9476);
or OR2 (N9481, N9470, N4348);
buf BUF1 (N9482, N9464);
nand NAND2 (N9483, N9471, N7256);
or OR2 (N9484, N9482, N6540);
nor NOR2 (N9485, N9478, N5408);
nor NOR2 (N9486, N9474, N6734);
or OR2 (N9487, N9481, N5944);
not NOT1 (N9488, N9469);
nand NAND4 (N9489, N9477, N4455, N3088, N1378);
nand NAND3 (N9490, N9480, N407, N6165);
and AND3 (N9491, N9487, N4643, N5887);
nand NAND3 (N9492, N9488, N6302, N765);
or OR2 (N9493, N9489, N4850);
not NOT1 (N9494, N9466);
xor XOR2 (N9495, N9483, N2609);
buf BUF1 (N9496, N9490);
nand NAND2 (N9497, N9493, N8195);
nor NOR3 (N9498, N9479, N8121, N7099);
nand NAND3 (N9499, N9491, N9397, N4943);
nor NOR4 (N9500, N9496, N895, N3275, N8250);
and AND2 (N9501, N9499, N7330);
and AND2 (N9502, N9497, N6963);
not NOT1 (N9503, N9492);
not NOT1 (N9504, N9502);
nor NOR2 (N9505, N9486, N2618);
xor XOR2 (N9506, N9500, N7272);
xor XOR2 (N9507, N9484, N9306);
nor NOR3 (N9508, N9485, N4002, N8824);
not NOT1 (N9509, N9505);
xor XOR2 (N9510, N9494, N8623);
xor XOR2 (N9511, N9508, N7019);
or OR3 (N9512, N9506, N6954, N6476);
nand NAND2 (N9513, N9509, N8846);
buf BUF1 (N9514, N9501);
nand NAND2 (N9515, N9507, N5233);
xor XOR2 (N9516, N9498, N3009);
or OR4 (N9517, N9516, N8075, N6646, N9229);
not NOT1 (N9518, N9495);
nor NOR3 (N9519, N9515, N6720, N8005);
not NOT1 (N9520, N9511);
xor XOR2 (N9521, N9503, N33);
nor NOR2 (N9522, N9520, N5786);
buf BUF1 (N9523, N9521);
buf BUF1 (N9524, N9512);
buf BUF1 (N9525, N9522);
or OR4 (N9526, N9504, N9279, N2008, N7390);
nand NAND3 (N9527, N9525, N2758, N4661);
buf BUF1 (N9528, N9517);
not NOT1 (N9529, N9524);
nand NAND3 (N9530, N9518, N8635, N8901);
and AND3 (N9531, N9523, N1858, N5503);
buf BUF1 (N9532, N9513);
nand NAND4 (N9533, N9529, N5048, N5325, N2498);
nor NOR4 (N9534, N9533, N5, N1552, N2511);
not NOT1 (N9535, N9527);
xor XOR2 (N9536, N9534, N3891);
buf BUF1 (N9537, N9530);
and AND2 (N9538, N9519, N2517);
not NOT1 (N9539, N9538);
or OR3 (N9540, N9539, N5146, N6013);
nor NOR2 (N9541, N9540, N3885);
nor NOR3 (N9542, N9541, N943, N9213);
buf BUF1 (N9543, N9537);
xor XOR2 (N9544, N9542, N1795);
xor XOR2 (N9545, N9532, N1933);
buf BUF1 (N9546, N9510);
xor XOR2 (N9547, N9535, N4496);
xor XOR2 (N9548, N9544, N2478);
buf BUF1 (N9549, N9536);
nand NAND3 (N9550, N9543, N3669, N8724);
nor NOR3 (N9551, N9546, N8131, N173);
nor NOR2 (N9552, N9549, N2442);
buf BUF1 (N9553, N9514);
nand NAND3 (N9554, N9553, N4978, N4939);
nor NOR2 (N9555, N9548, N7415);
nand NAND3 (N9556, N9545, N113, N6175);
nor NOR4 (N9557, N9552, N4845, N9204, N8602);
not NOT1 (N9558, N9531);
xor XOR2 (N9559, N9551, N2077);
xor XOR2 (N9560, N9547, N5976);
not NOT1 (N9561, N9560);
xor XOR2 (N9562, N9556, N6067);
and AND4 (N9563, N9559, N2554, N6084, N7646);
or OR3 (N9564, N9557, N2486, N118);
nor NOR4 (N9565, N9526, N5333, N543, N674);
or OR2 (N9566, N9565, N1206);
or OR3 (N9567, N9564, N7902, N9408);
or OR4 (N9568, N9528, N4527, N7077, N7880);
buf BUF1 (N9569, N9568);
not NOT1 (N9570, N9561);
or OR3 (N9571, N9554, N469, N3840);
or OR4 (N9572, N9563, N2771, N7947, N6093);
or OR3 (N9573, N9558, N1628, N6313);
and AND2 (N9574, N9572, N6208);
nand NAND4 (N9575, N9555, N9151, N1262, N2391);
or OR4 (N9576, N9566, N8907, N8428, N8410);
xor XOR2 (N9577, N9550, N8335);
or OR4 (N9578, N9576, N2186, N5635, N2354);
and AND3 (N9579, N9567, N1795, N2711);
xor XOR2 (N9580, N9573, N3079);
or OR2 (N9581, N9570, N1573);
and AND4 (N9582, N9574, N3850, N9399, N9579);
not NOT1 (N9583, N8051);
nor NOR4 (N9584, N9582, N2090, N8201, N2553);
xor XOR2 (N9585, N9571, N729);
xor XOR2 (N9586, N9584, N6038);
buf BUF1 (N9587, N9562);
nand NAND3 (N9588, N9580, N5829, N6170);
nand NAND3 (N9589, N9587, N3666, N3200);
nor NOR4 (N9590, N9569, N6415, N1903, N6096);
buf BUF1 (N9591, N9577);
nor NOR2 (N9592, N9581, N7574);
and AND4 (N9593, N9585, N6894, N4933, N7038);
buf BUF1 (N9594, N9583);
nand NAND2 (N9595, N9578, N4205);
not NOT1 (N9596, N9595);
and AND3 (N9597, N9586, N3902, N4998);
not NOT1 (N9598, N9575);
and AND3 (N9599, N9593, N3698, N4606);
buf BUF1 (N9600, N9599);
xor XOR2 (N9601, N9600, N3019);
buf BUF1 (N9602, N9588);
nor NOR4 (N9603, N9597, N6040, N8474, N3876);
buf BUF1 (N9604, N9602);
nand NAND2 (N9605, N9598, N915);
and AND3 (N9606, N9605, N9446, N1789);
xor XOR2 (N9607, N9591, N6721);
buf BUF1 (N9608, N9596);
or OR2 (N9609, N9603, N8320);
or OR2 (N9610, N9609, N7124);
nor NOR3 (N9611, N9592, N8586, N8356);
not NOT1 (N9612, N9607);
nor NOR3 (N9613, N9611, N4339, N8994);
nand NAND3 (N9614, N9590, N1376, N4914);
nor NOR3 (N9615, N9613, N2836, N8445);
nor NOR2 (N9616, N9601, N8610);
buf BUF1 (N9617, N9610);
buf BUF1 (N9618, N9612);
nor NOR2 (N9619, N9606, N8068);
or OR4 (N9620, N9616, N175, N916, N5998);
xor XOR2 (N9621, N9617, N1513);
nor NOR3 (N9622, N9614, N1667, N5601);
buf BUF1 (N9623, N9620);
nand NAND3 (N9624, N9589, N8988, N7824);
nand NAND3 (N9625, N9604, N9356, N7711);
xor XOR2 (N9626, N9623, N3697);
buf BUF1 (N9627, N9608);
and AND4 (N9628, N9624, N1422, N6913, N8446);
and AND3 (N9629, N9627, N2677, N1037);
or OR3 (N9630, N9594, N3299, N5124);
nor NOR2 (N9631, N9621, N6447);
nand NAND3 (N9632, N9622, N9589, N2841);
and AND3 (N9633, N9618, N4914, N6646);
buf BUF1 (N9634, N9630);
and AND3 (N9635, N9631, N569, N4950);
and AND2 (N9636, N9625, N4097);
nor NOR4 (N9637, N9636, N5790, N3458, N4257);
and AND4 (N9638, N9619, N5991, N3486, N2058);
not NOT1 (N9639, N9629);
buf BUF1 (N9640, N9638);
nand NAND2 (N9641, N9632, N135);
nor NOR2 (N9642, N9639, N3139);
nor NOR2 (N9643, N9641, N1700);
buf BUF1 (N9644, N9637);
nand NAND4 (N9645, N9640, N4280, N4626, N3016);
buf BUF1 (N9646, N9634);
not NOT1 (N9647, N9646);
and AND3 (N9648, N9647, N4034, N2399);
and AND3 (N9649, N9642, N7402, N5325);
and AND2 (N9650, N9645, N1269);
and AND3 (N9651, N9626, N4458, N7645);
and AND2 (N9652, N9650, N7815);
buf BUF1 (N9653, N9643);
not NOT1 (N9654, N9644);
xor XOR2 (N9655, N9653, N6538);
not NOT1 (N9656, N9651);
nand NAND3 (N9657, N9633, N6651, N5411);
nor NOR3 (N9658, N9652, N8805, N4598);
or OR2 (N9659, N9649, N6377);
nand NAND3 (N9660, N9657, N6057, N8112);
nor NOR2 (N9661, N9655, N7274);
and AND2 (N9662, N9648, N8581);
xor XOR2 (N9663, N9661, N9095);
or OR3 (N9664, N9635, N329, N6481);
buf BUF1 (N9665, N9658);
buf BUF1 (N9666, N9664);
nor NOR3 (N9667, N9628, N8423, N445);
and AND4 (N9668, N9666, N6818, N2373, N8443);
not NOT1 (N9669, N9656);
and AND2 (N9670, N9654, N6996);
and AND2 (N9671, N9669, N3866);
nor NOR3 (N9672, N9662, N5581, N5478);
nor NOR3 (N9673, N9663, N6393, N8904);
buf BUF1 (N9674, N9660);
nand NAND3 (N9675, N9674, N4612, N8387);
nand NAND3 (N9676, N9675, N4493, N5216);
buf BUF1 (N9677, N9671);
or OR4 (N9678, N9659, N3718, N9664, N8415);
or OR4 (N9679, N9667, N4617, N2961, N3462);
xor XOR2 (N9680, N9665, N2126);
not NOT1 (N9681, N9676);
nand NAND3 (N9682, N9668, N6896, N84);
buf BUF1 (N9683, N9678);
xor XOR2 (N9684, N9683, N1125);
nand NAND2 (N9685, N9670, N9069);
not NOT1 (N9686, N9680);
buf BUF1 (N9687, N9681);
buf BUF1 (N9688, N9615);
not NOT1 (N9689, N9672);
buf BUF1 (N9690, N9684);
or OR2 (N9691, N9673, N6585);
nand NAND4 (N9692, N9682, N4746, N8610, N9103);
or OR3 (N9693, N9687, N9288, N8582);
buf BUF1 (N9694, N9689);
or OR2 (N9695, N9686, N6079);
or OR3 (N9696, N9693, N1248, N7704);
nor NOR3 (N9697, N9695, N6155, N5750);
buf BUF1 (N9698, N9677);
buf BUF1 (N9699, N9692);
nor NOR2 (N9700, N9679, N2352);
and AND3 (N9701, N9696, N7074, N9659);
not NOT1 (N9702, N9697);
nor NOR3 (N9703, N9691, N6383, N4452);
not NOT1 (N9704, N9703);
buf BUF1 (N9705, N9702);
nand NAND3 (N9706, N9699, N1773, N7388);
or OR2 (N9707, N9688, N8951);
nand NAND3 (N9708, N9690, N3468, N3615);
not NOT1 (N9709, N9705);
buf BUF1 (N9710, N9698);
not NOT1 (N9711, N9706);
or OR2 (N9712, N9711, N8721);
xor XOR2 (N9713, N9710, N2065);
and AND2 (N9714, N9685, N5223);
or OR2 (N9715, N9708, N5688);
not NOT1 (N9716, N9694);
nand NAND3 (N9717, N9715, N348, N4297);
xor XOR2 (N9718, N9700, N8519);
nor NOR4 (N9719, N9716, N2560, N6325, N9103);
xor XOR2 (N9720, N9719, N2350);
nor NOR4 (N9721, N9714, N1661, N1167, N344);
xor XOR2 (N9722, N9707, N379);
and AND2 (N9723, N9718, N668);
nor NOR4 (N9724, N9709, N5360, N4740, N2893);
buf BUF1 (N9725, N9720);
nor NOR2 (N9726, N9725, N4829);
and AND4 (N9727, N9701, N7097, N3391, N5987);
buf BUF1 (N9728, N9727);
not NOT1 (N9729, N9713);
xor XOR2 (N9730, N9726, N5700);
not NOT1 (N9731, N9728);
and AND2 (N9732, N9729, N2016);
buf BUF1 (N9733, N9712);
nor NOR2 (N9734, N9724, N666);
xor XOR2 (N9735, N9704, N5833);
not NOT1 (N9736, N9735);
not NOT1 (N9737, N9733);
nand NAND4 (N9738, N9721, N4166, N1184, N6082);
or OR2 (N9739, N9737, N8269);
nand NAND3 (N9740, N9731, N9019, N4725);
xor XOR2 (N9741, N9717, N621);
or OR2 (N9742, N9738, N1993);
buf BUF1 (N9743, N9723);
buf BUF1 (N9744, N9732);
nand NAND2 (N9745, N9743, N8674);
nor NOR3 (N9746, N9740, N9154, N2346);
and AND3 (N9747, N9736, N4753, N8944);
not NOT1 (N9748, N9742);
or OR2 (N9749, N9730, N6318);
buf BUF1 (N9750, N9748);
xor XOR2 (N9751, N9741, N5194);
nor NOR2 (N9752, N9745, N4412);
buf BUF1 (N9753, N9722);
or OR3 (N9754, N9747, N3397, N4461);
and AND2 (N9755, N9734, N9027);
or OR2 (N9756, N9749, N2591);
not NOT1 (N9757, N9739);
buf BUF1 (N9758, N9744);
buf BUF1 (N9759, N9756);
or OR2 (N9760, N9751, N6698);
and AND4 (N9761, N9757, N882, N4390, N2201);
or OR4 (N9762, N9759, N6794, N8538, N8159);
and AND3 (N9763, N9752, N6814, N2586);
and AND4 (N9764, N9750, N6166, N4592, N8282);
and AND4 (N9765, N9754, N5809, N5367, N542);
or OR3 (N9766, N9761, N5811, N3982);
and AND2 (N9767, N9753, N1185);
nor NOR3 (N9768, N9760, N5770, N2936);
and AND4 (N9769, N9764, N5669, N9341, N6486);
xor XOR2 (N9770, N9768, N9538);
buf BUF1 (N9771, N9769);
nand NAND4 (N9772, N9746, N8683, N8378, N5172);
nand NAND2 (N9773, N9772, N2879);
and AND2 (N9774, N9765, N5527);
buf BUF1 (N9775, N9766);
nor NOR4 (N9776, N9755, N8202, N9009, N8677);
or OR3 (N9777, N9758, N7081, N5496);
xor XOR2 (N9778, N9775, N7162);
or OR4 (N9779, N9774, N5948, N9510, N5116);
buf BUF1 (N9780, N9779);
buf BUF1 (N9781, N9773);
nor NOR2 (N9782, N9763, N9036);
or OR4 (N9783, N9780, N4029, N9196, N690);
nor NOR3 (N9784, N9767, N1644, N2082);
and AND3 (N9785, N9777, N1732, N8024);
or OR3 (N9786, N9762, N705, N5428);
nor NOR2 (N9787, N9770, N7917);
and AND2 (N9788, N9782, N1989);
nor NOR2 (N9789, N9788, N1996);
nand NAND3 (N9790, N9787, N4236, N7326);
and AND3 (N9791, N9785, N3534, N4596);
xor XOR2 (N9792, N9778, N5780);
not NOT1 (N9793, N9781);
and AND2 (N9794, N9791, N2804);
nor NOR2 (N9795, N9789, N9646);
and AND3 (N9796, N9786, N5431, N3866);
or OR3 (N9797, N9783, N3262, N7160);
xor XOR2 (N9798, N9796, N9559);
and AND3 (N9799, N9793, N1764, N7683);
and AND2 (N9800, N9799, N4858);
or OR3 (N9801, N9794, N5987, N8532);
not NOT1 (N9802, N9784);
or OR2 (N9803, N9795, N8106);
nand NAND2 (N9804, N9803, N8775);
or OR3 (N9805, N9801, N6325, N3530);
nand NAND2 (N9806, N9790, N2689);
not NOT1 (N9807, N9806);
nor NOR3 (N9808, N9771, N1249, N8363);
and AND4 (N9809, N9808, N5715, N7939, N6995);
or OR4 (N9810, N9809, N4510, N7466, N9763);
nor NOR3 (N9811, N9776, N5455, N4153);
not NOT1 (N9812, N9802);
xor XOR2 (N9813, N9810, N5223);
nor NOR3 (N9814, N9797, N4445, N9193);
nand NAND2 (N9815, N9798, N1079);
and AND2 (N9816, N9807, N9719);
and AND4 (N9817, N9812, N8467, N2649, N2644);
nor NOR3 (N9818, N9814, N8118, N1795);
nor NOR3 (N9819, N9818, N1181, N8652);
and AND3 (N9820, N9813, N6973, N8803);
nor NOR4 (N9821, N9817, N6452, N5714, N5768);
or OR4 (N9822, N9819, N8116, N4620, N532);
xor XOR2 (N9823, N9821, N8979);
not NOT1 (N9824, N9823);
not NOT1 (N9825, N9792);
or OR2 (N9826, N9804, N2643);
and AND4 (N9827, N9805, N4706, N950, N172);
and AND2 (N9828, N9800, N9790);
nand NAND3 (N9829, N9827, N9491, N7138);
nor NOR2 (N9830, N9815, N3834);
nor NOR3 (N9831, N9829, N1691, N5364);
nand NAND2 (N9832, N9811, N1442);
nand NAND4 (N9833, N9831, N5616, N8527, N6679);
nand NAND4 (N9834, N9825, N7164, N2042, N2415);
not NOT1 (N9835, N9826);
and AND2 (N9836, N9828, N1545);
not NOT1 (N9837, N9835);
not NOT1 (N9838, N9830);
xor XOR2 (N9839, N9838, N5931);
and AND3 (N9840, N9839, N4087, N152);
not NOT1 (N9841, N9836);
buf BUF1 (N9842, N9822);
and AND4 (N9843, N9840, N2868, N2737, N7993);
nand NAND3 (N9844, N9824, N9078, N1207);
xor XOR2 (N9845, N9833, N9146);
buf BUF1 (N9846, N9820);
xor XOR2 (N9847, N9834, N2518);
and AND4 (N9848, N9832, N2417, N8203, N404);
and AND4 (N9849, N9842, N6084, N2817, N7748);
or OR3 (N9850, N9847, N3553, N5024);
and AND4 (N9851, N9841, N7918, N2733, N5430);
nand NAND4 (N9852, N9843, N1039, N3387, N1853);
xor XOR2 (N9853, N9850, N7722);
not NOT1 (N9854, N9853);
xor XOR2 (N9855, N9844, N6037);
or OR4 (N9856, N9845, N504, N3286, N1183);
nor NOR3 (N9857, N9837, N3393, N9579);
not NOT1 (N9858, N9848);
nand NAND4 (N9859, N9816, N1013, N9447, N5164);
or OR2 (N9860, N9855, N7029);
xor XOR2 (N9861, N9854, N8379);
nand NAND4 (N9862, N9857, N9410, N5935, N1066);
nor NOR2 (N9863, N9849, N4285);
and AND2 (N9864, N9861, N1585);
or OR2 (N9865, N9863, N8805);
nand NAND2 (N9866, N9852, N9393);
nand NAND3 (N9867, N9860, N8226, N2201);
and AND3 (N9868, N9851, N2580, N5412);
nand NAND4 (N9869, N9859, N493, N6027, N7332);
or OR4 (N9870, N9867, N1693, N4187, N7830);
or OR4 (N9871, N9870, N343, N3393, N3193);
or OR2 (N9872, N9856, N2045);
and AND2 (N9873, N9868, N3450);
not NOT1 (N9874, N9865);
xor XOR2 (N9875, N9872, N1657);
nor NOR3 (N9876, N9874, N6666, N9413);
buf BUF1 (N9877, N9873);
not NOT1 (N9878, N9875);
nor NOR2 (N9879, N9864, N313);
nand NAND4 (N9880, N9862, N909, N4540, N1571);
nor NOR3 (N9881, N9866, N1327, N7086);
or OR3 (N9882, N9881, N5887, N6322);
or OR2 (N9883, N9846, N6997);
nand NAND2 (N9884, N9869, N2441);
not NOT1 (N9885, N9883);
nor NOR4 (N9886, N9878, N9805, N3007, N8887);
nand NAND2 (N9887, N9858, N9400);
not NOT1 (N9888, N9886);
nand NAND2 (N9889, N9882, N6221);
xor XOR2 (N9890, N9888, N8859);
or OR4 (N9891, N9879, N5908, N6226, N6692);
xor XOR2 (N9892, N9877, N9439);
buf BUF1 (N9893, N9890);
not NOT1 (N9894, N9876);
and AND4 (N9895, N9893, N6669, N2504, N7003);
nor NOR2 (N9896, N9880, N5743);
buf BUF1 (N9897, N9891);
xor XOR2 (N9898, N9887, N2883);
or OR4 (N9899, N9898, N636, N1829, N7249);
or OR3 (N9900, N9894, N9831, N4191);
nor NOR3 (N9901, N9899, N1543, N2403);
nor NOR3 (N9902, N9892, N1411, N5193);
nand NAND3 (N9903, N9885, N7030, N1653);
nand NAND3 (N9904, N9889, N8057, N4133);
buf BUF1 (N9905, N9897);
not NOT1 (N9906, N9903);
or OR4 (N9907, N9900, N6005, N2716, N3918);
nand NAND2 (N9908, N9871, N3685);
buf BUF1 (N9909, N9905);
xor XOR2 (N9910, N9906, N6498);
xor XOR2 (N9911, N9895, N2523);
xor XOR2 (N9912, N9907, N2872);
xor XOR2 (N9913, N9912, N5534);
nand NAND3 (N9914, N9901, N2102, N6467);
nor NOR3 (N9915, N9909, N6003, N6330);
not NOT1 (N9916, N9910);
nor NOR3 (N9917, N9884, N7258, N728);
not NOT1 (N9918, N9908);
nor NOR2 (N9919, N9918, N7111);
nor NOR4 (N9920, N9916, N2662, N7008, N4301);
buf BUF1 (N9921, N9919);
nor NOR4 (N9922, N9917, N848, N3482, N3790);
buf BUF1 (N9923, N9904);
nor NOR2 (N9924, N9920, N7241);
nor NOR2 (N9925, N9902, N7304);
or OR3 (N9926, N9923, N5315, N1772);
buf BUF1 (N9927, N9926);
or OR2 (N9928, N9927, N3372);
xor XOR2 (N9929, N9924, N293);
nor NOR3 (N9930, N9928, N4606, N2239);
buf BUF1 (N9931, N9929);
xor XOR2 (N9932, N9914, N2323);
buf BUF1 (N9933, N9911);
buf BUF1 (N9934, N9922);
buf BUF1 (N9935, N9921);
not NOT1 (N9936, N9915);
or OR2 (N9937, N9935, N1280);
nor NOR2 (N9938, N9936, N6345);
and AND2 (N9939, N9934, N1979);
nand NAND4 (N9940, N9937, N7187, N6324, N7883);
and AND4 (N9941, N9938, N1557, N5830, N2831);
buf BUF1 (N9942, N9930);
buf BUF1 (N9943, N9913);
nor NOR2 (N9944, N9943, N5278);
and AND3 (N9945, N9933, N8527, N5384);
and AND3 (N9946, N9932, N5926, N5142);
or OR4 (N9947, N9896, N6610, N61, N4642);
and AND2 (N9948, N9946, N8317);
nand NAND2 (N9949, N9940, N2807);
xor XOR2 (N9950, N9947, N9488);
and AND2 (N9951, N9925, N8363);
not NOT1 (N9952, N9945);
buf BUF1 (N9953, N9942);
xor XOR2 (N9954, N9948, N11);
nand NAND4 (N9955, N9931, N8218, N4468, N5557);
and AND3 (N9956, N9951, N6386, N3170);
nor NOR2 (N9957, N9941, N5610);
xor XOR2 (N9958, N9949, N3475);
and AND3 (N9959, N9953, N6495, N2510);
or OR4 (N9960, N9939, N2361, N2416, N3704);
nand NAND2 (N9961, N9959, N3431);
xor XOR2 (N9962, N9944, N9109);
not NOT1 (N9963, N9961);
nand NAND4 (N9964, N9952, N4048, N5876, N9098);
and AND4 (N9965, N9962, N2237, N2825, N7378);
and AND3 (N9966, N9958, N218, N2875);
and AND2 (N9967, N9963, N8752);
nor NOR2 (N9968, N9950, N4979);
and AND4 (N9969, N9968, N6686, N3438, N4810);
xor XOR2 (N9970, N9957, N8708);
buf BUF1 (N9971, N9965);
nand NAND4 (N9972, N9955, N9661, N6234, N2776);
nand NAND3 (N9973, N9967, N7658, N4495);
and AND4 (N9974, N9956, N8970, N1574, N6869);
buf BUF1 (N9975, N9964);
or OR4 (N9976, N9960, N5731, N510, N5980);
nor NOR3 (N9977, N9969, N5599, N9831);
nor NOR4 (N9978, N9972, N1723, N617, N190);
buf BUF1 (N9979, N9971);
buf BUF1 (N9980, N9978);
or OR2 (N9981, N9966, N7555);
nor NOR3 (N9982, N9974, N6263, N7910);
or OR4 (N9983, N9979, N2059, N1224, N2304);
nand NAND4 (N9984, N9973, N3209, N3326, N4793);
or OR3 (N9985, N9977, N9358, N6207);
xor XOR2 (N9986, N9984, N2390);
xor XOR2 (N9987, N9986, N2818);
not NOT1 (N9988, N9954);
nor NOR4 (N9989, N9981, N4569, N5042, N9304);
xor XOR2 (N9990, N9980, N3356);
or OR3 (N9991, N9987, N1394, N3071);
nand NAND2 (N9992, N9983, N2313);
nor NOR3 (N9993, N9975, N98, N9698);
buf BUF1 (N9994, N9992);
nand NAND3 (N9995, N9985, N2145, N2410);
and AND4 (N9996, N9988, N8860, N2141, N7125);
not NOT1 (N9997, N9993);
or OR2 (N9998, N9991, N8983);
xor XOR2 (N9999, N9997, N6344);
nor NOR2 (N10000, N9998, N4859);
nor NOR2 (N10001, N9976, N919);
nand NAND3 (N10002, N9996, N303, N1177);
xor XOR2 (N10003, N9994, N1767);
not NOT1 (N10004, N9970);
or OR2 (N10005, N10003, N1519);
nand NAND2 (N10006, N10000, N4020);
nor NOR2 (N10007, N9999, N270);
and AND2 (N10008, N10006, N7974);
or OR4 (N10009, N10008, N8301, N1349, N8414);
xor XOR2 (N10010, N10004, N4154);
nand NAND3 (N10011, N10009, N6558, N9529);
xor XOR2 (N10012, N10005, N9938);
buf BUF1 (N10013, N10012);
buf BUF1 (N10014, N10013);
not NOT1 (N10015, N10014);
or OR4 (N10016, N9995, N8508, N3678, N7565);
and AND4 (N10017, N9990, N407, N3846, N3398);
buf BUF1 (N10018, N9989);
not NOT1 (N10019, N10015);
xor XOR2 (N10020, N10001, N8930);
buf BUF1 (N10021, N10019);
buf BUF1 (N10022, N10016);
and AND4 (N10023, N10020, N3272, N4320, N5552);
xor XOR2 (N10024, N10002, N3041);
nand NAND4 (N10025, N10022, N6383, N1375, N3083);
xor XOR2 (N10026, N10024, N9644);
nand NAND2 (N10027, N10011, N3234);
nand NAND3 (N10028, N10027, N9158, N9454);
buf BUF1 (N10029, N10026);
not NOT1 (N10030, N10028);
xor XOR2 (N10031, N10018, N25);
or OR2 (N10032, N10029, N7042);
and AND3 (N10033, N9982, N5769, N7860);
buf BUF1 (N10034, N10017);
buf BUF1 (N10035, N10025);
or OR2 (N10036, N10033, N1262);
nor NOR4 (N10037, N10035, N6091, N4185, N6523);
buf BUF1 (N10038, N10037);
buf BUF1 (N10039, N10032);
nor NOR4 (N10040, N10038, N8277, N542, N1104);
not NOT1 (N10041, N10039);
nor NOR2 (N10042, N10010, N2316);
or OR3 (N10043, N10042, N4229, N1460);
and AND4 (N10044, N10031, N1838, N5385, N2533);
or OR2 (N10045, N10036, N5020);
and AND2 (N10046, N10023, N1104);
xor XOR2 (N10047, N10021, N3585);
nand NAND3 (N10048, N10045, N8405, N6615);
nor NOR2 (N10049, N10007, N3533);
nor NOR3 (N10050, N10046, N1100, N2249);
and AND4 (N10051, N10049, N326, N1627, N4691);
not NOT1 (N10052, N10034);
buf BUF1 (N10053, N10043);
or OR3 (N10054, N10047, N8571, N1920);
or OR3 (N10055, N10050, N1470, N3500);
and AND4 (N10056, N10055, N7918, N1195, N7183);
and AND3 (N10057, N10056, N2053, N1563);
nor NOR4 (N10058, N10044, N3484, N7771, N4535);
or OR4 (N10059, N10053, N3435, N5864, N4550);
buf BUF1 (N10060, N10041);
and AND2 (N10061, N10057, N4233);
nor NOR4 (N10062, N10061, N7326, N4285, N4147);
nand NAND3 (N10063, N10059, N1689, N5439);
not NOT1 (N10064, N10030);
nor NOR3 (N10065, N10052, N7306, N230);
buf BUF1 (N10066, N10040);
or OR2 (N10067, N10060, N7738);
not NOT1 (N10068, N10048);
nor NOR2 (N10069, N10062, N7176);
nand NAND4 (N10070, N10067, N6987, N6803, N763);
xor XOR2 (N10071, N10058, N7298);
xor XOR2 (N10072, N10070, N3590);
nand NAND2 (N10073, N10051, N86);
xor XOR2 (N10074, N10064, N8546);
nand NAND4 (N10075, N10065, N5300, N3728, N1155);
nand NAND2 (N10076, N10066, N6019);
nor NOR2 (N10077, N10073, N7844);
and AND4 (N10078, N10074, N1382, N854, N1792);
nor NOR3 (N10079, N10063, N9032, N607);
xor XOR2 (N10080, N10054, N6766);
buf BUF1 (N10081, N10075);
and AND2 (N10082, N10068, N1892);
nand NAND4 (N10083, N10071, N2362, N2875, N10065);
not NOT1 (N10084, N10080);
nand NAND4 (N10085, N10069, N8194, N9117, N2129);
xor XOR2 (N10086, N10084, N447);
nor NOR3 (N10087, N10076, N4105, N3331);
xor XOR2 (N10088, N10085, N114);
or OR4 (N10089, N10077, N1173, N7205, N5736);
not NOT1 (N10090, N10072);
not NOT1 (N10091, N10090);
buf BUF1 (N10092, N10089);
not NOT1 (N10093, N10088);
not NOT1 (N10094, N10091);
xor XOR2 (N10095, N10079, N5321);
xor XOR2 (N10096, N10078, N5082);
buf BUF1 (N10097, N10094);
xor XOR2 (N10098, N10086, N1646);
xor XOR2 (N10099, N10082, N5154);
nor NOR3 (N10100, N10098, N1862, N8391);
and AND2 (N10101, N10100, N7093);
nor NOR3 (N10102, N10092, N3058, N5407);
nor NOR2 (N10103, N10095, N9000);
or OR2 (N10104, N10103, N8744);
buf BUF1 (N10105, N10096);
nand NAND2 (N10106, N10104, N938);
or OR4 (N10107, N10093, N3854, N2442, N10011);
and AND4 (N10108, N10102, N2965, N3989, N4371);
and AND2 (N10109, N10108, N6961);
nor NOR4 (N10110, N10081, N9076, N4862, N5831);
buf BUF1 (N10111, N10099);
buf BUF1 (N10112, N10111);
nand NAND4 (N10113, N10110, N3823, N5626, N1551);
buf BUF1 (N10114, N10087);
or OR3 (N10115, N10113, N5098, N1150);
nor NOR4 (N10116, N10115, N1960, N526, N436);
not NOT1 (N10117, N10112);
not NOT1 (N10118, N10083);
or OR3 (N10119, N10107, N6106, N6507);
nor NOR3 (N10120, N10105, N5194, N7624);
nor NOR2 (N10121, N10119, N7617);
not NOT1 (N10122, N10101);
or OR3 (N10123, N10120, N7666, N9194);
or OR3 (N10124, N10121, N7906, N5179);
and AND3 (N10125, N10123, N2593, N665);
not NOT1 (N10126, N10117);
not NOT1 (N10127, N10114);
xor XOR2 (N10128, N10109, N1884);
nor NOR4 (N10129, N10124, N2011, N4806, N615);
and AND3 (N10130, N10126, N2364, N9729);
nor NOR4 (N10131, N10125, N8293, N7429, N6451);
or OR2 (N10132, N10131, N3149);
nor NOR4 (N10133, N10128, N1, N3478, N9312);
nor NOR3 (N10134, N10118, N4491, N7478);
nor NOR4 (N10135, N10129, N2290, N9473, N7490);
and AND3 (N10136, N10132, N1631, N7963);
nand NAND2 (N10137, N10122, N3812);
buf BUF1 (N10138, N10135);
or OR2 (N10139, N10130, N7491);
xor XOR2 (N10140, N10138, N2016);
nand NAND3 (N10141, N10097, N4206, N6032);
and AND3 (N10142, N10106, N5741, N1605);
nand NAND3 (N10143, N10134, N4550, N379);
not NOT1 (N10144, N10139);
buf BUF1 (N10145, N10144);
buf BUF1 (N10146, N10141);
nor NOR2 (N10147, N10146, N2837);
nor NOR2 (N10148, N10116, N629);
buf BUF1 (N10149, N10148);
or OR3 (N10150, N10145, N1338, N5679);
or OR3 (N10151, N10127, N1559, N5676);
or OR3 (N10152, N10140, N3151, N1999);
or OR2 (N10153, N10151, N1356);
buf BUF1 (N10154, N10147);
nand NAND3 (N10155, N10153, N752, N4260);
and AND4 (N10156, N10155, N944, N9934, N1123);
or OR4 (N10157, N10137, N3713, N3834, N4266);
not NOT1 (N10158, N10152);
nor NOR2 (N10159, N10136, N2816);
buf BUF1 (N10160, N10133);
nor NOR3 (N10161, N10150, N3713, N7960);
nor NOR2 (N10162, N10158, N1208);
xor XOR2 (N10163, N10143, N3664);
buf BUF1 (N10164, N10161);
xor XOR2 (N10165, N10142, N9470);
xor XOR2 (N10166, N10149, N8538);
and AND2 (N10167, N10163, N5715);
xor XOR2 (N10168, N10160, N3140);
not NOT1 (N10169, N10166);
or OR3 (N10170, N10156, N9297, N4390);
nor NOR2 (N10171, N10170, N5303);
or OR4 (N10172, N10167, N9399, N5826, N1628);
or OR3 (N10173, N10169, N1210, N8173);
xor XOR2 (N10174, N10168, N1928);
nand NAND3 (N10175, N10154, N8798, N8436);
not NOT1 (N10176, N10174);
and AND3 (N10177, N10173, N6304, N5474);
xor XOR2 (N10178, N10176, N7370);
xor XOR2 (N10179, N10159, N4025);
nor NOR2 (N10180, N10178, N7602);
nand NAND2 (N10181, N10175, N5921);
or OR4 (N10182, N10177, N3768, N9088, N4070);
nor NOR3 (N10183, N10162, N9102, N3033);
buf BUF1 (N10184, N10157);
buf BUF1 (N10185, N10171);
nor NOR4 (N10186, N10164, N7240, N4265, N360);
buf BUF1 (N10187, N10181);
nand NAND4 (N10188, N10187, N9866, N9943, N6951);
not NOT1 (N10189, N10188);
not NOT1 (N10190, N10180);
nand NAND2 (N10191, N10183, N200);
xor XOR2 (N10192, N10165, N4654);
xor XOR2 (N10193, N10185, N8799);
and AND4 (N10194, N10179, N464, N7084, N7470);
xor XOR2 (N10195, N10190, N3316);
nor NOR4 (N10196, N10194, N351, N1057, N377);
or OR3 (N10197, N10195, N6533, N1623);
and AND4 (N10198, N10197, N2405, N7518, N6680);
xor XOR2 (N10199, N10193, N2722);
buf BUF1 (N10200, N10191);
buf BUF1 (N10201, N10198);
not NOT1 (N10202, N10199);
buf BUF1 (N10203, N10196);
nand NAND4 (N10204, N10192, N1316, N8215, N4831);
buf BUF1 (N10205, N10201);
nand NAND3 (N10206, N10204, N4382, N4802);
and AND2 (N10207, N10203, N3504);
nand NAND3 (N10208, N10172, N4265, N271);
and AND2 (N10209, N10182, N9731);
not NOT1 (N10210, N10207);
and AND4 (N10211, N10200, N8056, N5469, N9490);
buf BUF1 (N10212, N10184);
nand NAND2 (N10213, N10205, N6986);
not NOT1 (N10214, N10212);
and AND4 (N10215, N10186, N7445, N8384, N8467);
and AND4 (N10216, N10189, N9064, N3080, N8043);
not NOT1 (N10217, N10209);
buf BUF1 (N10218, N10213);
nand NAND4 (N10219, N10218, N4554, N3098, N8692);
buf BUF1 (N10220, N10215);
nor NOR4 (N10221, N10202, N118, N6055, N9291);
and AND3 (N10222, N10211, N1327, N9543);
nand NAND3 (N10223, N10216, N3462, N3495);
not NOT1 (N10224, N10222);
and AND4 (N10225, N10210, N5208, N6184, N4133);
buf BUF1 (N10226, N10224);
xor XOR2 (N10227, N10223, N4734);
buf BUF1 (N10228, N10226);
xor XOR2 (N10229, N10219, N2783);
xor XOR2 (N10230, N10227, N7216);
or OR3 (N10231, N10229, N4741, N10039);
nor NOR3 (N10232, N10221, N4105, N851);
not NOT1 (N10233, N10214);
and AND4 (N10234, N10233, N1297, N9645, N3078);
nand NAND4 (N10235, N10208, N5021, N5237, N6108);
buf BUF1 (N10236, N10232);
xor XOR2 (N10237, N10235, N5811);
nand NAND2 (N10238, N10237, N3601);
not NOT1 (N10239, N10206);
and AND2 (N10240, N10220, N4247);
and AND2 (N10241, N10239, N6033);
not NOT1 (N10242, N10225);
not NOT1 (N10243, N10230);
nand NAND2 (N10244, N10241, N8707);
xor XOR2 (N10245, N10234, N7644);
nand NAND3 (N10246, N10243, N469, N7656);
buf BUF1 (N10247, N10236);
xor XOR2 (N10248, N10244, N5588);
not NOT1 (N10249, N10228);
and AND4 (N10250, N10240, N6211, N3382, N7651);
xor XOR2 (N10251, N10245, N8459);
not NOT1 (N10252, N10246);
and AND2 (N10253, N10247, N7994);
nand NAND2 (N10254, N10231, N1430);
or OR4 (N10255, N10251, N1501, N10036, N2378);
buf BUF1 (N10256, N10250);
nor NOR4 (N10257, N10249, N3500, N6865, N3386);
nor NOR4 (N10258, N10253, N235, N6955, N8441);
and AND3 (N10259, N10238, N3798, N5519);
and AND4 (N10260, N10256, N8361, N6246, N9407);
or OR4 (N10261, N10259, N4761, N4570, N3981);
nor NOR3 (N10262, N10255, N1163, N130);
nor NOR4 (N10263, N10262, N5808, N3913, N3395);
or OR4 (N10264, N10261, N9885, N5935, N9259);
and AND3 (N10265, N10217, N2311, N3964);
or OR4 (N10266, N10265, N3654, N824, N6923);
and AND3 (N10267, N10254, N4745, N6711);
nor NOR3 (N10268, N10260, N405, N5893);
and AND4 (N10269, N10257, N7991, N8035, N5798);
not NOT1 (N10270, N10263);
buf BUF1 (N10271, N10264);
nand NAND3 (N10272, N10269, N4886, N4497);
xor XOR2 (N10273, N10270, N4377);
or OR3 (N10274, N10242, N2221, N274);
not NOT1 (N10275, N10274);
nand NAND2 (N10276, N10272, N6505);
xor XOR2 (N10277, N10267, N2758);
or OR4 (N10278, N10276, N293, N3569, N983);
or OR2 (N10279, N10278, N6840);
buf BUF1 (N10280, N10277);
or OR3 (N10281, N10271, N2537, N1323);
xor XOR2 (N10282, N10266, N1396);
and AND3 (N10283, N10275, N1602, N828);
xor XOR2 (N10284, N10268, N161);
and AND3 (N10285, N10284, N8259, N5220);
nor NOR2 (N10286, N10258, N5380);
or OR2 (N10287, N10281, N7468);
nand NAND3 (N10288, N10282, N98, N140);
and AND3 (N10289, N10252, N4540, N8456);
nand NAND2 (N10290, N10273, N7570);
and AND3 (N10291, N10283, N4094, N8118);
buf BUF1 (N10292, N10290);
or OR4 (N10293, N10288, N10176, N3462, N8961);
xor XOR2 (N10294, N10279, N9494);
buf BUF1 (N10295, N10287);
nor NOR4 (N10296, N10280, N8899, N2419, N6448);
buf BUF1 (N10297, N10295);
and AND4 (N10298, N10296, N852, N912, N3192);
and AND3 (N10299, N10291, N480, N5316);
nor NOR3 (N10300, N10248, N3118, N8058);
buf BUF1 (N10301, N10294);
and AND4 (N10302, N10299, N1441, N8090, N6834);
not NOT1 (N10303, N10300);
or OR4 (N10304, N10303, N6116, N6394, N4983);
xor XOR2 (N10305, N10304, N2709);
and AND4 (N10306, N10293, N6919, N4149, N10248);
xor XOR2 (N10307, N10305, N4166);
not NOT1 (N10308, N10285);
xor XOR2 (N10309, N10289, N4699);
or OR3 (N10310, N10302, N5404, N5357);
xor XOR2 (N10311, N10298, N3559);
nand NAND3 (N10312, N10301, N8877, N5503);
or OR4 (N10313, N10297, N9611, N9572, N890);
or OR2 (N10314, N10313, N4969);
xor XOR2 (N10315, N10310, N8611);
nand NAND3 (N10316, N10292, N8451, N8292);
and AND3 (N10317, N10308, N7068, N7673);
or OR2 (N10318, N10311, N5364);
not NOT1 (N10319, N10317);
xor XOR2 (N10320, N10316, N926);
xor XOR2 (N10321, N10320, N8375);
nor NOR3 (N10322, N10312, N2335, N3061);
xor XOR2 (N10323, N10286, N7185);
not NOT1 (N10324, N10314);
nor NOR3 (N10325, N10307, N4212, N3222);
nor NOR4 (N10326, N10324, N1736, N7101, N3538);
xor XOR2 (N10327, N10315, N8110);
and AND2 (N10328, N10325, N3178);
buf BUF1 (N10329, N10321);
nand NAND4 (N10330, N10326, N1995, N2641, N1479);
nand NAND2 (N10331, N10327, N470);
buf BUF1 (N10332, N10306);
buf BUF1 (N10333, N10323);
or OR3 (N10334, N10309, N4479, N3165);
buf BUF1 (N10335, N10318);
and AND3 (N10336, N10328, N8464, N5451);
nand NAND2 (N10337, N10331, N6000);
and AND4 (N10338, N10330, N3005, N7035, N8272);
and AND3 (N10339, N10322, N4080, N4478);
nand NAND3 (N10340, N10334, N8622, N8208);
or OR2 (N10341, N10338, N6111);
nor NOR4 (N10342, N10339, N3417, N2467, N433);
or OR2 (N10343, N10336, N352);
and AND4 (N10344, N10319, N542, N6457, N2730);
not NOT1 (N10345, N10344);
xor XOR2 (N10346, N10329, N2840);
buf BUF1 (N10347, N10335);
nand NAND2 (N10348, N10345, N4945);
nor NOR4 (N10349, N10333, N3765, N1837, N8833);
nor NOR3 (N10350, N10349, N1976, N7285);
and AND3 (N10351, N10332, N9520, N8783);
not NOT1 (N10352, N10346);
nor NOR2 (N10353, N10343, N5000);
nand NAND2 (N10354, N10350, N7912);
nor NOR4 (N10355, N10353, N9443, N6571, N697);
buf BUF1 (N10356, N10341);
nor NOR4 (N10357, N10342, N5952, N3862, N3787);
or OR3 (N10358, N10351, N9445, N9350);
and AND2 (N10359, N10348, N9014);
or OR2 (N10360, N10354, N978);
buf BUF1 (N10361, N10355);
xor XOR2 (N10362, N10358, N3222);
or OR3 (N10363, N10359, N9771, N889);
not NOT1 (N10364, N10352);
not NOT1 (N10365, N10364);
not NOT1 (N10366, N10356);
and AND2 (N10367, N10340, N543);
or OR2 (N10368, N10347, N3418);
buf BUF1 (N10369, N10366);
nand NAND3 (N10370, N10368, N8834, N4629);
xor XOR2 (N10371, N10362, N9933);
xor XOR2 (N10372, N10365, N9564);
nand NAND3 (N10373, N10372, N8790, N5982);
nor NOR2 (N10374, N10371, N188);
buf BUF1 (N10375, N10363);
and AND3 (N10376, N10367, N4972, N8543);
and AND4 (N10377, N10357, N4426, N9682, N487);
buf BUF1 (N10378, N10337);
xor XOR2 (N10379, N10378, N9599);
not NOT1 (N10380, N10379);
xor XOR2 (N10381, N10361, N1555);
nand NAND4 (N10382, N10377, N320, N4745, N8152);
xor XOR2 (N10383, N10382, N3092);
xor XOR2 (N10384, N10376, N3131);
buf BUF1 (N10385, N10373);
and AND3 (N10386, N10370, N6844, N487);
nand NAND4 (N10387, N10383, N1571, N2151, N2928);
nor NOR3 (N10388, N10387, N6595, N6920);
and AND3 (N10389, N10380, N3245, N2462);
xor XOR2 (N10390, N10386, N3393);
xor XOR2 (N10391, N10384, N2329);
xor XOR2 (N10392, N10389, N703);
not NOT1 (N10393, N10360);
nand NAND3 (N10394, N10369, N9204, N5690);
not NOT1 (N10395, N10381);
and AND2 (N10396, N10393, N1377);
not NOT1 (N10397, N10394);
nand NAND2 (N10398, N10390, N7142);
buf BUF1 (N10399, N10395);
buf BUF1 (N10400, N10374);
buf BUF1 (N10401, N10400);
and AND4 (N10402, N10375, N4646, N9756, N3209);
and AND3 (N10403, N10401, N1125, N8796);
xor XOR2 (N10404, N10398, N6888);
xor XOR2 (N10405, N10392, N5701);
buf BUF1 (N10406, N10385);
nand NAND4 (N10407, N10391, N3123, N6797, N8008);
nor NOR3 (N10408, N10407, N8980, N710);
not NOT1 (N10409, N10396);
not NOT1 (N10410, N10405);
nand NAND3 (N10411, N10409, N9238, N4674);
nand NAND2 (N10412, N10408, N347);
nor NOR4 (N10413, N10388, N1168, N773, N6156);
xor XOR2 (N10414, N10399, N10254);
nor NOR4 (N10415, N10406, N6057, N834, N7744);
and AND3 (N10416, N10397, N4465, N1346);
and AND3 (N10417, N10416, N424, N6937);
xor XOR2 (N10418, N10417, N2894);
buf BUF1 (N10419, N10414);
and AND3 (N10420, N10404, N3995, N1224);
or OR2 (N10421, N10420, N762);
and AND2 (N10422, N10402, N6446);
not NOT1 (N10423, N10419);
buf BUF1 (N10424, N10413);
nand NAND2 (N10425, N10411, N278);
xor XOR2 (N10426, N10412, N683);
xor XOR2 (N10427, N10410, N6636);
not NOT1 (N10428, N10424);
buf BUF1 (N10429, N10426);
buf BUF1 (N10430, N10403);
or OR3 (N10431, N10415, N7672, N2994);
buf BUF1 (N10432, N10428);
not NOT1 (N10433, N10430);
buf BUF1 (N10434, N10427);
nor NOR2 (N10435, N10425, N8069);
nand NAND4 (N10436, N10422, N2127, N3963, N5431);
not NOT1 (N10437, N10432);
or OR2 (N10438, N10431, N7448);
or OR3 (N10439, N10418, N2585, N1128);
nor NOR4 (N10440, N10439, N3909, N5321, N10341);
or OR4 (N10441, N10433, N3059, N1996, N2848);
buf BUF1 (N10442, N10437);
nand NAND3 (N10443, N10421, N8883, N4247);
xor XOR2 (N10444, N10440, N634);
nand NAND3 (N10445, N10436, N6310, N4105);
and AND4 (N10446, N10434, N2304, N9905, N7371);
xor XOR2 (N10447, N10446, N4935);
nand NAND3 (N10448, N10441, N1374, N3058);
nor NOR4 (N10449, N10444, N5598, N3191, N8548);
not NOT1 (N10450, N10449);
nor NOR4 (N10451, N10438, N1081, N8480, N7860);
and AND3 (N10452, N10442, N6651, N6504);
xor XOR2 (N10453, N10450, N106);
and AND4 (N10454, N10429, N3595, N4130, N4083);
xor XOR2 (N10455, N10423, N4165);
and AND4 (N10456, N10452, N6438, N10117, N2227);
and AND3 (N10457, N10451, N2274, N9335);
buf BUF1 (N10458, N10455);
buf BUF1 (N10459, N10453);
buf BUF1 (N10460, N10457);
buf BUF1 (N10461, N10447);
xor XOR2 (N10462, N10460, N3691);
nor NOR4 (N10463, N10443, N599, N9053, N7057);
not NOT1 (N10464, N10445);
not NOT1 (N10465, N10458);
nor NOR2 (N10466, N10464, N5461);
not NOT1 (N10467, N10456);
and AND4 (N10468, N10461, N1235, N9879, N4578);
nand NAND4 (N10469, N10454, N3259, N5928, N3393);
buf BUF1 (N10470, N10448);
nor NOR3 (N10471, N10465, N1242, N5219);
xor XOR2 (N10472, N10468, N8323);
and AND3 (N10473, N10472, N8415, N9436);
nor NOR2 (N10474, N10466, N3028);
and AND3 (N10475, N10467, N7747, N8497);
or OR3 (N10476, N10462, N10388, N5881);
nand NAND4 (N10477, N10473, N1627, N4399, N2362);
buf BUF1 (N10478, N10471);
buf BUF1 (N10479, N10435);
nor NOR2 (N10480, N10479, N5582);
xor XOR2 (N10481, N10469, N4255);
nor NOR3 (N10482, N10477, N4561, N5285);
not NOT1 (N10483, N10482);
not NOT1 (N10484, N10481);
not NOT1 (N10485, N10478);
or OR3 (N10486, N10484, N1970, N4440);
xor XOR2 (N10487, N10474, N8483);
xor XOR2 (N10488, N10476, N7870);
or OR4 (N10489, N10459, N6084, N3118, N1585);
nor NOR4 (N10490, N10485, N1229, N6795, N3592);
nand NAND4 (N10491, N10475, N8726, N622, N9962);
buf BUF1 (N10492, N10463);
or OR3 (N10493, N10492, N241, N6290);
xor XOR2 (N10494, N10486, N10330);
nand NAND3 (N10495, N10493, N6638, N912);
nor NOR4 (N10496, N10490, N1823, N3554, N7182);
not NOT1 (N10497, N10470);
or OR4 (N10498, N10483, N6504, N7313, N5791);
nand NAND4 (N10499, N10488, N3292, N2591, N7799);
nand NAND3 (N10500, N10494, N6283, N6136);
nand NAND4 (N10501, N10495, N1494, N8849, N5804);
nand NAND3 (N10502, N10496, N1005, N1502);
xor XOR2 (N10503, N10489, N4990);
nand NAND2 (N10504, N10500, N323);
nor NOR4 (N10505, N10480, N6201, N3690, N7388);
not NOT1 (N10506, N10498);
not NOT1 (N10507, N10499);
not NOT1 (N10508, N10504);
and AND2 (N10509, N10487, N10233);
nand NAND2 (N10510, N10505, N2446);
and AND2 (N10511, N10501, N9825);
buf BUF1 (N10512, N10491);
and AND3 (N10513, N10503, N1036, N9009);
xor XOR2 (N10514, N10507, N2164);
or OR2 (N10515, N10514, N7875);
or OR2 (N10516, N10506, N1748);
buf BUF1 (N10517, N10512);
not NOT1 (N10518, N10516);
and AND3 (N10519, N10502, N5395, N2430);
or OR4 (N10520, N10508, N3273, N9956, N4609);
not NOT1 (N10521, N10520);
or OR4 (N10522, N10521, N1893, N10196, N9928);
nor NOR3 (N10523, N10517, N9875, N3136);
buf BUF1 (N10524, N10523);
not NOT1 (N10525, N10497);
and AND3 (N10526, N10513, N697, N4877);
not NOT1 (N10527, N10515);
nand NAND3 (N10528, N10525, N6619, N6665);
nand NAND3 (N10529, N10528, N5020, N7599);
buf BUF1 (N10530, N10519);
nand NAND4 (N10531, N10524, N2698, N5134, N7817);
xor XOR2 (N10532, N10531, N3777);
nor NOR2 (N10533, N10526, N1892);
xor XOR2 (N10534, N10510, N9294);
nor NOR2 (N10535, N10518, N4385);
xor XOR2 (N10536, N10529, N9430);
nor NOR2 (N10537, N10527, N6290);
nor NOR3 (N10538, N10537, N3517, N3475);
not NOT1 (N10539, N10522);
and AND2 (N10540, N10534, N307);
not NOT1 (N10541, N10536);
buf BUF1 (N10542, N10509);
buf BUF1 (N10543, N10535);
buf BUF1 (N10544, N10533);
xor XOR2 (N10545, N10511, N8536);
buf BUF1 (N10546, N10538);
nor NOR3 (N10547, N10541, N8474, N6608);
or OR3 (N10548, N10540, N6465, N178);
nor NOR3 (N10549, N10545, N7661, N2851);
nand NAND4 (N10550, N10547, N3676, N9318, N5682);
nand NAND3 (N10551, N10542, N9255, N7896);
nor NOR4 (N10552, N10543, N5728, N7079, N7544);
xor XOR2 (N10553, N10530, N359);
and AND2 (N10554, N10548, N8810);
nand NAND3 (N10555, N10552, N7376, N6176);
nand NAND2 (N10556, N10546, N5016);
or OR2 (N10557, N10551, N1053);
and AND2 (N10558, N10532, N6811);
not NOT1 (N10559, N10556);
nand NAND2 (N10560, N10549, N5941);
and AND4 (N10561, N10560, N5879, N8773, N7454);
and AND2 (N10562, N10554, N2380);
nor NOR4 (N10563, N10558, N10264, N1179, N324);
not NOT1 (N10564, N10539);
nor NOR4 (N10565, N10555, N4105, N76, N7388);
and AND3 (N10566, N10550, N6000, N6103);
not NOT1 (N10567, N10566);
xor XOR2 (N10568, N10553, N2861);
and AND4 (N10569, N10559, N1906, N6333, N72);
buf BUF1 (N10570, N10568);
buf BUF1 (N10571, N10565);
not NOT1 (N10572, N10567);
and AND4 (N10573, N10562, N816, N2779, N1770);
not NOT1 (N10574, N10569);
nand NAND4 (N10575, N10557, N3656, N3050, N8294);
nor NOR2 (N10576, N10564, N9459);
nand NAND2 (N10577, N10573, N7835);
not NOT1 (N10578, N10561);
xor XOR2 (N10579, N10572, N1137);
or OR2 (N10580, N10563, N5615);
nand NAND2 (N10581, N10580, N6615);
xor XOR2 (N10582, N10544, N5940);
and AND2 (N10583, N10578, N1122);
buf BUF1 (N10584, N10577);
xor XOR2 (N10585, N10571, N8724);
or OR4 (N10586, N10582, N6122, N4770, N4551);
xor XOR2 (N10587, N10570, N7964);
and AND2 (N10588, N10583, N551);
or OR3 (N10589, N10574, N8321, N2452);
xor XOR2 (N10590, N10576, N3222);
nor NOR3 (N10591, N10586, N4390, N4371);
not NOT1 (N10592, N10590);
buf BUF1 (N10593, N10585);
nand NAND2 (N10594, N10589, N3237);
or OR4 (N10595, N10581, N1087, N9658, N6284);
or OR3 (N10596, N10593, N6775, N929);
or OR2 (N10597, N10594, N5651);
not NOT1 (N10598, N10575);
nor NOR3 (N10599, N10588, N6322, N316);
buf BUF1 (N10600, N10598);
nand NAND2 (N10601, N10595, N5134);
buf BUF1 (N10602, N10579);
buf BUF1 (N10603, N10584);
and AND4 (N10604, N10602, N6036, N6147, N4585);
buf BUF1 (N10605, N10597);
nor NOR4 (N10606, N10592, N2756, N1398, N4302);
not NOT1 (N10607, N10599);
buf BUF1 (N10608, N10600);
not NOT1 (N10609, N10591);
nand NAND3 (N10610, N10601, N7446, N5316);
nand NAND3 (N10611, N10604, N9223, N704);
not NOT1 (N10612, N10609);
nor NOR3 (N10613, N10603, N2924, N2452);
nand NAND4 (N10614, N10596, N1151, N3125, N3072);
and AND3 (N10615, N10612, N9787, N8108);
nor NOR4 (N10616, N10587, N10360, N5914, N8412);
not NOT1 (N10617, N10610);
xor XOR2 (N10618, N10607, N3489);
and AND4 (N10619, N10614, N8238, N7821, N3671);
xor XOR2 (N10620, N10617, N2249);
nand NAND3 (N10621, N10615, N5938, N6281);
not NOT1 (N10622, N10613);
nand NAND2 (N10623, N10606, N8459);
xor XOR2 (N10624, N10605, N10436);
nor NOR3 (N10625, N10622, N2875, N3727);
xor XOR2 (N10626, N10619, N7615);
nand NAND3 (N10627, N10618, N9829, N3756);
nor NOR4 (N10628, N10627, N6066, N4347, N8025);
nand NAND4 (N10629, N10611, N4465, N7140, N10400);
xor XOR2 (N10630, N10624, N8231);
and AND3 (N10631, N10630, N4592, N798);
not NOT1 (N10632, N10631);
nand NAND4 (N10633, N10616, N7648, N6939, N7125);
nor NOR2 (N10634, N10620, N4657);
or OR3 (N10635, N10628, N1849, N939);
not NOT1 (N10636, N10633);
nand NAND4 (N10637, N10634, N8557, N7832, N8539);
buf BUF1 (N10638, N10626);
not NOT1 (N10639, N10635);
nor NOR3 (N10640, N10638, N4517, N9402);
not NOT1 (N10641, N10640);
xor XOR2 (N10642, N10637, N2309);
buf BUF1 (N10643, N10636);
nand NAND4 (N10644, N10642, N2597, N3701, N4592);
not NOT1 (N10645, N10608);
not NOT1 (N10646, N10629);
xor XOR2 (N10647, N10644, N7532);
not NOT1 (N10648, N10632);
not NOT1 (N10649, N10648);
not NOT1 (N10650, N10621);
not NOT1 (N10651, N10641);
not NOT1 (N10652, N10646);
and AND4 (N10653, N10639, N7970, N9489, N9011);
nor NOR3 (N10654, N10649, N1079, N5985);
buf BUF1 (N10655, N10647);
or OR2 (N10656, N10643, N2709);
xor XOR2 (N10657, N10656, N3270);
and AND2 (N10658, N10625, N2085);
not NOT1 (N10659, N10651);
buf BUF1 (N10660, N10659);
not NOT1 (N10661, N10650);
or OR3 (N10662, N10645, N6197, N8446);
or OR3 (N10663, N10652, N9526, N20);
and AND3 (N10664, N10623, N3079, N8509);
or OR4 (N10665, N10661, N7928, N6517, N9717);
nand NAND4 (N10666, N10658, N7932, N7859, N4957);
nand NAND3 (N10667, N10662, N490, N523);
buf BUF1 (N10668, N10657);
buf BUF1 (N10669, N10663);
not NOT1 (N10670, N10665);
or OR3 (N10671, N10668, N1679, N5017);
and AND2 (N10672, N10660, N7205);
nor NOR2 (N10673, N10655, N9218);
or OR3 (N10674, N10670, N3961, N8423);
and AND3 (N10675, N10666, N1176, N10113);
and AND3 (N10676, N10654, N2391, N6587);
or OR3 (N10677, N10669, N1937, N3785);
not NOT1 (N10678, N10672);
or OR2 (N10679, N10653, N7236);
nand NAND4 (N10680, N10664, N3099, N9239, N4876);
not NOT1 (N10681, N10674);
xor XOR2 (N10682, N10675, N392);
xor XOR2 (N10683, N10667, N7965);
xor XOR2 (N10684, N10676, N2338);
nand NAND2 (N10685, N10673, N10371);
nand NAND4 (N10686, N10671, N2020, N4052, N8666);
or OR2 (N10687, N10680, N5487);
or OR3 (N10688, N10678, N9852, N3093);
xor XOR2 (N10689, N10688, N526);
not NOT1 (N10690, N10686);
buf BUF1 (N10691, N10679);
not NOT1 (N10692, N10691);
xor XOR2 (N10693, N10690, N7349);
not NOT1 (N10694, N10687);
nor NOR4 (N10695, N10689, N5275, N3761, N3267);
and AND4 (N10696, N10693, N5674, N9098, N1878);
xor XOR2 (N10697, N10692, N5358);
nand NAND4 (N10698, N10682, N7629, N176, N8668);
nand NAND3 (N10699, N10681, N3434, N9329);
not NOT1 (N10700, N10696);
and AND2 (N10701, N10684, N3213);
nand NAND4 (N10702, N10700, N69, N6661, N3580);
or OR4 (N10703, N10699, N8547, N9575, N8323);
not NOT1 (N10704, N10697);
nand NAND3 (N10705, N10703, N2391, N5651);
not NOT1 (N10706, N10695);
xor XOR2 (N10707, N10677, N5429);
not NOT1 (N10708, N10706);
and AND3 (N10709, N10685, N6786, N3996);
not NOT1 (N10710, N10683);
not NOT1 (N10711, N10694);
nor NOR4 (N10712, N10704, N3481, N7702, N9071);
buf BUF1 (N10713, N10710);
xor XOR2 (N10714, N10712, N3796);
not NOT1 (N10715, N10701);
not NOT1 (N10716, N10698);
and AND2 (N10717, N10709, N8070);
nor NOR2 (N10718, N10702, N9757);
or OR3 (N10719, N10713, N8134, N4502);
or OR3 (N10720, N10717, N10445, N3518);
or OR3 (N10721, N10715, N4363, N256);
xor XOR2 (N10722, N10714, N8317);
not NOT1 (N10723, N10711);
or OR3 (N10724, N10718, N7776, N6452);
nor NOR3 (N10725, N10724, N7623, N1162);
and AND2 (N10726, N10716, N2590);
not NOT1 (N10727, N10719);
xor XOR2 (N10728, N10720, N938);
not NOT1 (N10729, N10726);
nor NOR3 (N10730, N10729, N9798, N4182);
buf BUF1 (N10731, N10723);
xor XOR2 (N10732, N10731, N6286);
or OR4 (N10733, N10728, N9223, N77, N448);
buf BUF1 (N10734, N10733);
nand NAND2 (N10735, N10722, N4849);
and AND2 (N10736, N10705, N9703);
xor XOR2 (N10737, N10734, N9723);
not NOT1 (N10738, N10727);
and AND4 (N10739, N10708, N7828, N4761, N2607);
buf BUF1 (N10740, N10736);
nand NAND2 (N10741, N10732, N9097);
xor XOR2 (N10742, N10725, N7089);
buf BUF1 (N10743, N10737);
or OR2 (N10744, N10741, N8983);
not NOT1 (N10745, N10739);
or OR4 (N10746, N10738, N8731, N4388, N1574);
nor NOR3 (N10747, N10743, N4711, N5938);
and AND4 (N10748, N10747, N9893, N5132, N10404);
buf BUF1 (N10749, N10707);
or OR2 (N10750, N10740, N5557);
nand NAND2 (N10751, N10721, N7434);
xor XOR2 (N10752, N10748, N8214);
buf BUF1 (N10753, N10752);
nand NAND2 (N10754, N10750, N2454);
xor XOR2 (N10755, N10749, N8762);
buf BUF1 (N10756, N10745);
buf BUF1 (N10757, N10755);
or OR4 (N10758, N10735, N5317, N6433, N8194);
and AND3 (N10759, N10756, N6755, N8038);
and AND4 (N10760, N10754, N8083, N10010, N5491);
xor XOR2 (N10761, N10757, N10673);
buf BUF1 (N10762, N10730);
xor XOR2 (N10763, N10761, N542);
not NOT1 (N10764, N10763);
nor NOR2 (N10765, N10759, N2248);
or OR3 (N10766, N10751, N7971, N2757);
nor NOR3 (N10767, N10760, N5281, N9965);
nand NAND3 (N10768, N10753, N6897, N4202);
buf BUF1 (N10769, N10766);
buf BUF1 (N10770, N10758);
nand NAND3 (N10771, N10764, N8433, N5192);
or OR4 (N10772, N10771, N8650, N7208, N5555);
or OR2 (N10773, N10772, N7187);
buf BUF1 (N10774, N10765);
and AND4 (N10775, N10770, N3563, N8411, N6549);
nor NOR2 (N10776, N10767, N9298);
or OR3 (N10777, N10773, N8284, N8226);
nand NAND3 (N10778, N10762, N9272, N10688);
buf BUF1 (N10779, N10744);
buf BUF1 (N10780, N10775);
and AND3 (N10781, N10742, N8603, N395);
or OR3 (N10782, N10746, N7823, N1125);
nand NAND3 (N10783, N10768, N6354, N6083);
xor XOR2 (N10784, N10779, N10653);
buf BUF1 (N10785, N10782);
nand NAND4 (N10786, N10774, N7235, N2366, N2520);
nand NAND3 (N10787, N10769, N5392, N4061);
buf BUF1 (N10788, N10777);
or OR2 (N10789, N10784, N7705);
xor XOR2 (N10790, N10786, N3705);
or OR4 (N10791, N10776, N2114, N7865, N7357);
not NOT1 (N10792, N10787);
and AND2 (N10793, N10790, N812);
nand NAND2 (N10794, N10791, N4006);
and AND2 (N10795, N10788, N8094);
xor XOR2 (N10796, N10794, N1187);
not NOT1 (N10797, N10785);
or OR4 (N10798, N10796, N9522, N3294, N5820);
and AND3 (N10799, N10780, N1736, N1576);
or OR4 (N10800, N10793, N10392, N475, N61);
not NOT1 (N10801, N10778);
buf BUF1 (N10802, N10801);
or OR4 (N10803, N10799, N6699, N2303, N10182);
nor NOR4 (N10804, N10792, N6065, N1258, N8817);
nand NAND2 (N10805, N10795, N8679);
or OR2 (N10806, N10800, N3959);
buf BUF1 (N10807, N10789);
or OR4 (N10808, N10781, N2310, N4353, N10211);
xor XOR2 (N10809, N10803, N8780);
not NOT1 (N10810, N10807);
nor NOR2 (N10811, N10809, N5588);
buf BUF1 (N10812, N10802);
nand NAND3 (N10813, N10797, N3485, N7693);
not NOT1 (N10814, N10798);
nand NAND2 (N10815, N10811, N2664);
and AND3 (N10816, N10783, N1317, N3955);
xor XOR2 (N10817, N10813, N9709);
or OR2 (N10818, N10814, N127);
and AND3 (N10819, N10810, N1572, N2669);
buf BUF1 (N10820, N10808);
nor NOR3 (N10821, N10817, N4528, N176);
nor NOR4 (N10822, N10812, N2747, N3039, N4156);
or OR4 (N10823, N10804, N153, N1211, N2674);
and AND4 (N10824, N10821, N3781, N2948, N7453);
nand NAND3 (N10825, N10815, N4385, N2294);
not NOT1 (N10826, N10825);
or OR4 (N10827, N10820, N9496, N5355, N2150);
nand NAND4 (N10828, N10823, N5485, N10263, N4788);
nand NAND4 (N10829, N10827, N8073, N2205, N5302);
xor XOR2 (N10830, N10828, N7876);
or OR2 (N10831, N10816, N6330);
nand NAND3 (N10832, N10818, N1195, N6265);
and AND4 (N10833, N10806, N1807, N477, N1960);
nor NOR4 (N10834, N10822, N1105, N2990, N9156);
not NOT1 (N10835, N10830);
xor XOR2 (N10836, N10805, N1883);
and AND3 (N10837, N10832, N2426, N7306);
or OR3 (N10838, N10829, N8755, N7878);
nand NAND2 (N10839, N10819, N875);
and AND2 (N10840, N10838, N6015);
not NOT1 (N10841, N10833);
or OR4 (N10842, N10840, N7305, N6738, N277);
nand NAND2 (N10843, N10835, N10384);
not NOT1 (N10844, N10843);
nand NAND2 (N10845, N10826, N9713);
nand NAND4 (N10846, N10841, N7591, N4278, N2123);
or OR3 (N10847, N10842, N5803, N3896);
nand NAND4 (N10848, N10831, N3867, N1483, N7042);
and AND3 (N10849, N10844, N4393, N7375);
nand NAND2 (N10850, N10837, N3977);
nor NOR4 (N10851, N10847, N1069, N1494, N2364);
or OR2 (N10852, N10845, N3130);
and AND4 (N10853, N10846, N7403, N5999, N1278);
nor NOR2 (N10854, N10836, N6084);
or OR4 (N10855, N10824, N5367, N2382, N798);
or OR4 (N10856, N10850, N7687, N6003, N9223);
nand NAND3 (N10857, N10849, N9876, N888);
buf BUF1 (N10858, N10854);
xor XOR2 (N10859, N10855, N7121);
not NOT1 (N10860, N10853);
xor XOR2 (N10861, N10839, N9028);
nor NOR4 (N10862, N10834, N4095, N7706, N5569);
nor NOR3 (N10863, N10856, N3595, N7196);
not NOT1 (N10864, N10861);
nand NAND3 (N10865, N10859, N2446, N1933);
and AND4 (N10866, N10864, N31, N5433, N5038);
nand NAND4 (N10867, N10852, N976, N7618, N1088);
nor NOR4 (N10868, N10860, N3580, N8275, N3563);
nor NOR2 (N10869, N10863, N2191);
xor XOR2 (N10870, N10862, N1120);
or OR2 (N10871, N10848, N869);
nand NAND2 (N10872, N10870, N8330);
xor XOR2 (N10873, N10866, N6282);
and AND4 (N10874, N10851, N5588, N4464, N771);
xor XOR2 (N10875, N10872, N3492);
not NOT1 (N10876, N10875);
and AND2 (N10877, N10874, N2820);
and AND3 (N10878, N10876, N1556, N5407);
buf BUF1 (N10879, N10873);
xor XOR2 (N10880, N10858, N1977);
buf BUF1 (N10881, N10878);
or OR3 (N10882, N10867, N8195, N5236);
nand NAND2 (N10883, N10857, N4981);
nand NAND3 (N10884, N10869, N697, N8492);
not NOT1 (N10885, N10880);
nand NAND2 (N10886, N10881, N4564);
nand NAND4 (N10887, N10883, N9258, N5169, N7208);
nand NAND4 (N10888, N10868, N10285, N1465, N1079);
buf BUF1 (N10889, N10886);
not NOT1 (N10890, N10882);
not NOT1 (N10891, N10890);
xor XOR2 (N10892, N10888, N7752);
xor XOR2 (N10893, N10871, N6914);
not NOT1 (N10894, N10887);
xor XOR2 (N10895, N10893, N389);
xor XOR2 (N10896, N10889, N4807);
nor NOR2 (N10897, N10895, N1926);
and AND2 (N10898, N10896, N4274);
not NOT1 (N10899, N10865);
xor XOR2 (N10900, N10899, N8306);
and AND4 (N10901, N10900, N6828, N3188, N3064);
and AND3 (N10902, N10898, N4807, N7438);
and AND4 (N10903, N10891, N9244, N6934, N10276);
nand NAND4 (N10904, N10894, N7225, N5156, N6540);
and AND2 (N10905, N10877, N428);
buf BUF1 (N10906, N10902);
xor XOR2 (N10907, N10892, N7869);
buf BUF1 (N10908, N10901);
buf BUF1 (N10909, N10897);
or OR4 (N10910, N10905, N10872, N3327, N6751);
or OR2 (N10911, N10910, N486);
buf BUF1 (N10912, N10908);
nand NAND2 (N10913, N10911, N1347);
nand NAND3 (N10914, N10912, N3943, N14);
or OR3 (N10915, N10906, N7144, N5333);
nor NOR2 (N10916, N10884, N7695);
not NOT1 (N10917, N10915);
nand NAND2 (N10918, N10909, N4941);
nand NAND4 (N10919, N10907, N2571, N1290, N10066);
not NOT1 (N10920, N10916);
not NOT1 (N10921, N10918);
nor NOR3 (N10922, N10919, N944, N9185);
nor NOR3 (N10923, N10921, N10370, N8276);
and AND2 (N10924, N10923, N1054);
xor XOR2 (N10925, N10914, N10309);
nand NAND4 (N10926, N10917, N7691, N1952, N9619);
buf BUF1 (N10927, N10879);
not NOT1 (N10928, N10920);
buf BUF1 (N10929, N10904);
or OR2 (N10930, N10913, N7780);
not NOT1 (N10931, N10924);
buf BUF1 (N10932, N10927);
nand NAND3 (N10933, N10931, N9026, N49);
and AND4 (N10934, N10925, N5959, N9028, N10091);
or OR4 (N10935, N10928, N1742, N4235, N7995);
buf BUF1 (N10936, N10922);
and AND3 (N10937, N10932, N4481, N5393);
xor XOR2 (N10938, N10926, N2826);
nor NOR3 (N10939, N10930, N3136, N3570);
or OR2 (N10940, N10885, N4885);
not NOT1 (N10941, N10936);
nor NOR3 (N10942, N10903, N2019, N7614);
and AND3 (N10943, N10934, N556, N3951);
and AND3 (N10944, N10937, N8962, N3700);
xor XOR2 (N10945, N10935, N731);
nor NOR2 (N10946, N10941, N834);
nand NAND2 (N10947, N10946, N6546);
nand NAND3 (N10948, N10942, N26, N8695);
and AND4 (N10949, N10947, N3226, N4932, N2670);
and AND4 (N10950, N10945, N8291, N8134, N10444);
or OR3 (N10951, N10950, N8248, N10136);
not NOT1 (N10952, N10944);
and AND4 (N10953, N10939, N10929, N631, N1315);
xor XOR2 (N10954, N824, N563);
xor XOR2 (N10955, N10938, N2327);
or OR4 (N10956, N10933, N5429, N621, N1713);
not NOT1 (N10957, N10953);
nand NAND2 (N10958, N10957, N10856);
or OR4 (N10959, N10954, N2901, N10110, N542);
nand NAND3 (N10960, N10959, N8086, N7701);
xor XOR2 (N10961, N10956, N1719);
or OR3 (N10962, N10955, N7422, N1985);
xor XOR2 (N10963, N10962, N492);
xor XOR2 (N10964, N10958, N9140);
and AND4 (N10965, N10964, N1573, N3154, N2979);
buf BUF1 (N10966, N10961);
not NOT1 (N10967, N10943);
or OR4 (N10968, N10963, N8042, N1625, N10580);
xor XOR2 (N10969, N10940, N8916);
nor NOR4 (N10970, N10966, N10267, N5713, N1223);
xor XOR2 (N10971, N10967, N7346);
nand NAND3 (N10972, N10968, N10761, N5498);
and AND3 (N10973, N10952, N10918, N9157);
buf BUF1 (N10974, N10973);
not NOT1 (N10975, N10948);
buf BUF1 (N10976, N10949);
nand NAND3 (N10977, N10970, N2679, N2902);
and AND2 (N10978, N10972, N2505);
xor XOR2 (N10979, N10976, N6322);
not NOT1 (N10980, N10977);
and AND2 (N10981, N10980, N9538);
not NOT1 (N10982, N10981);
buf BUF1 (N10983, N10982);
and AND2 (N10984, N10983, N2724);
buf BUF1 (N10985, N10971);
buf BUF1 (N10986, N10985);
not NOT1 (N10987, N10978);
buf BUF1 (N10988, N10974);
not NOT1 (N10989, N10969);
nand NAND4 (N10990, N10987, N7402, N542, N8833);
or OR4 (N10991, N10988, N1725, N1393, N6525);
buf BUF1 (N10992, N10951);
nor NOR4 (N10993, N10984, N9114, N4122, N5281);
nor NOR2 (N10994, N10975, N4691);
nor NOR3 (N10995, N10993, N8854, N5126);
buf BUF1 (N10996, N10986);
nor NOR2 (N10997, N10994, N6105);
nor NOR3 (N10998, N10996, N208, N544);
xor XOR2 (N10999, N10995, N417);
not NOT1 (N11000, N10997);
nor NOR3 (N11001, N10992, N10511, N4946);
or OR3 (N11002, N10960, N3848, N6413);
xor XOR2 (N11003, N11002, N4977);
and AND4 (N11004, N10990, N907, N4500, N2207);
or OR3 (N11005, N10999, N7240, N6551);
nor NOR4 (N11006, N11001, N1853, N825, N6136);
xor XOR2 (N11007, N10991, N3907);
nand NAND2 (N11008, N11006, N9761);
and AND3 (N11009, N11005, N8253, N248);
nand NAND4 (N11010, N10979, N5218, N3659, N10578);
not NOT1 (N11011, N11010);
xor XOR2 (N11012, N10989, N3539);
xor XOR2 (N11013, N11012, N2407);
not NOT1 (N11014, N11011);
not NOT1 (N11015, N11007);
and AND3 (N11016, N11000, N3923, N2785);
nor NOR3 (N11017, N11015, N7122, N2434);
not NOT1 (N11018, N11013);
not NOT1 (N11019, N11004);
nor NOR3 (N11020, N10965, N10398, N9067);
or OR2 (N11021, N10998, N2295);
and AND3 (N11022, N11019, N9494, N9134);
xor XOR2 (N11023, N11022, N9186);
xor XOR2 (N11024, N11008, N6192);
xor XOR2 (N11025, N11020, N10960);
xor XOR2 (N11026, N11009, N3815);
and AND2 (N11027, N11016, N7939);
nand NAND4 (N11028, N11026, N1262, N6294, N9507);
or OR4 (N11029, N11018, N1231, N5613, N2169);
or OR3 (N11030, N11025, N2838, N10101);
and AND4 (N11031, N11014, N2693, N2390, N10119);
xor XOR2 (N11032, N11024, N9916);
or OR3 (N11033, N11021, N9171, N10471);
nand NAND2 (N11034, N11029, N6731);
or OR4 (N11035, N11017, N6143, N5143, N3977);
not NOT1 (N11036, N11035);
nor NOR3 (N11037, N11023, N2650, N984);
or OR2 (N11038, N11028, N8388);
nor NOR3 (N11039, N11033, N8011, N5657);
nor NOR2 (N11040, N11032, N816);
or OR3 (N11041, N11036, N6679, N2767);
nor NOR2 (N11042, N11034, N7627);
nand NAND2 (N11043, N11042, N1591);
nor NOR2 (N11044, N11038, N9228);
or OR4 (N11045, N11044, N924, N6759, N10875);
xor XOR2 (N11046, N11003, N8575);
buf BUF1 (N11047, N11031);
nor NOR4 (N11048, N11045, N3050, N7337, N3666);
buf BUF1 (N11049, N11043);
or OR3 (N11050, N11040, N4001, N10302);
nand NAND3 (N11051, N11030, N7712, N8222);
buf BUF1 (N11052, N11039);
nand NAND2 (N11053, N11046, N9845);
buf BUF1 (N11054, N11047);
or OR3 (N11055, N11054, N9379, N1095);
buf BUF1 (N11056, N11051);
not NOT1 (N11057, N11027);
and AND4 (N11058, N11041, N434, N8866, N9548);
not NOT1 (N11059, N11058);
nor NOR4 (N11060, N11059, N7127, N6599, N131);
and AND2 (N11061, N11048, N8825);
xor XOR2 (N11062, N11056, N385);
and AND2 (N11063, N11061, N4922);
nand NAND3 (N11064, N11050, N2372, N2922);
nor NOR3 (N11065, N11037, N3739, N3524);
buf BUF1 (N11066, N11062);
nand NAND2 (N11067, N11060, N9848);
and AND4 (N11068, N11057, N9355, N8729, N2393);
and AND4 (N11069, N11064, N6470, N7293, N2837);
buf BUF1 (N11070, N11063);
not NOT1 (N11071, N11053);
nand NAND4 (N11072, N11071, N7082, N10513, N10350);
and AND4 (N11073, N11052, N68, N4227, N3685);
buf BUF1 (N11074, N11067);
or OR4 (N11075, N11074, N2821, N4274, N9202);
or OR4 (N11076, N11066, N6623, N8116, N8731);
buf BUF1 (N11077, N11072);
nand NAND4 (N11078, N11055, N4776, N6256, N3333);
and AND3 (N11079, N11075, N10582, N8113);
xor XOR2 (N11080, N11077, N3094);
nor NOR4 (N11081, N11073, N153, N2690, N4054);
buf BUF1 (N11082, N11080);
nand NAND4 (N11083, N11068, N5866, N7877, N2996);
nor NOR2 (N11084, N11079, N8242);
nand NAND3 (N11085, N11076, N3013, N5152);
buf BUF1 (N11086, N11070);
xor XOR2 (N11087, N11085, N6812);
not NOT1 (N11088, N11086);
nor NOR3 (N11089, N11083, N7095, N10584);
not NOT1 (N11090, N11049);
nand NAND3 (N11091, N11089, N3416, N2801);
nand NAND2 (N11092, N11088, N2538);
buf BUF1 (N11093, N11082);
buf BUF1 (N11094, N11087);
nand NAND3 (N11095, N11065, N10171, N10764);
nand NAND2 (N11096, N11090, N4308);
xor XOR2 (N11097, N11081, N7071);
or OR4 (N11098, N11095, N26, N1027, N5940);
nand NAND4 (N11099, N11097, N9465, N9844, N2762);
xor XOR2 (N11100, N11069, N8618);
not NOT1 (N11101, N11093);
and AND4 (N11102, N11096, N6376, N5142, N5521);
or OR3 (N11103, N11101, N8194, N5553);
not NOT1 (N11104, N11100);
not NOT1 (N11105, N11102);
or OR2 (N11106, N11078, N1368);
not NOT1 (N11107, N11106);
and AND2 (N11108, N11104, N7541);
not NOT1 (N11109, N11103);
nor NOR3 (N11110, N11094, N3660, N4213);
buf BUF1 (N11111, N11107);
nand NAND3 (N11112, N11092, N8694, N9938);
xor XOR2 (N11113, N11105, N9166);
not NOT1 (N11114, N11084);
or OR3 (N11115, N11098, N5515, N6979);
nor NOR2 (N11116, N11108, N6857);
nand NAND4 (N11117, N11115, N2173, N2439, N2560);
or OR4 (N11118, N11113, N10776, N8842, N1136);
buf BUF1 (N11119, N11117);
not NOT1 (N11120, N11114);
not NOT1 (N11121, N11091);
not NOT1 (N11122, N11112);
nor NOR2 (N11123, N11116, N8015);
nor NOR3 (N11124, N11120, N3087, N9269);
buf BUF1 (N11125, N11119);
not NOT1 (N11126, N11099);
not NOT1 (N11127, N11126);
buf BUF1 (N11128, N11124);
or OR2 (N11129, N11121, N5032);
or OR2 (N11130, N11128, N5761);
nor NOR3 (N11131, N11111, N6530, N9375);
or OR3 (N11132, N11125, N5460, N6124);
xor XOR2 (N11133, N11131, N10537);
and AND4 (N11134, N11129, N6009, N1994, N2071);
not NOT1 (N11135, N11122);
not NOT1 (N11136, N11118);
nand NAND3 (N11137, N11136, N6925, N1939);
xor XOR2 (N11138, N11110, N5918);
nor NOR2 (N11139, N11127, N5596);
or OR2 (N11140, N11139, N2268);
nor NOR2 (N11141, N11134, N3828);
nor NOR4 (N11142, N11133, N3187, N745, N8772);
nand NAND2 (N11143, N11140, N8601);
buf BUF1 (N11144, N11143);
buf BUF1 (N11145, N11141);
xor XOR2 (N11146, N11145, N8007);
or OR3 (N11147, N11142, N11065, N3485);
not NOT1 (N11148, N11135);
or OR2 (N11149, N11137, N2816);
buf BUF1 (N11150, N11147);
buf BUF1 (N11151, N11148);
buf BUF1 (N11152, N11138);
or OR2 (N11153, N11151, N1501);
nor NOR4 (N11154, N11132, N2782, N2024, N157);
nor NOR3 (N11155, N11154, N7526, N6094);
xor XOR2 (N11156, N11123, N1885);
nor NOR4 (N11157, N11152, N8310, N2995, N4297);
nor NOR2 (N11158, N11109, N8056);
or OR2 (N11159, N11146, N6203);
or OR2 (N11160, N11157, N204);
nand NAND2 (N11161, N11160, N3798);
buf BUF1 (N11162, N11161);
xor XOR2 (N11163, N11159, N1459);
or OR2 (N11164, N11130, N4782);
nand NAND4 (N11165, N11163, N9707, N9867, N4510);
nor NOR3 (N11166, N11144, N8019, N4298);
xor XOR2 (N11167, N11162, N3038);
nor NOR3 (N11168, N11150, N1169, N8979);
buf BUF1 (N11169, N11149);
xor XOR2 (N11170, N11167, N1964);
not NOT1 (N11171, N11156);
or OR2 (N11172, N11165, N5624);
nand NAND4 (N11173, N11155, N10841, N7291, N3192);
nand NAND4 (N11174, N11169, N1623, N1339, N378);
buf BUF1 (N11175, N11170);
buf BUF1 (N11176, N11168);
and AND4 (N11177, N11158, N420, N6654, N7888);
not NOT1 (N11178, N11177);
nand NAND3 (N11179, N11172, N10490, N8628);
nor NOR4 (N11180, N11179, N7690, N6474, N2182);
xor XOR2 (N11181, N11175, N8360);
or OR2 (N11182, N11164, N4233);
nor NOR4 (N11183, N11181, N8476, N5394, N11059);
not NOT1 (N11184, N11166);
not NOT1 (N11185, N11173);
xor XOR2 (N11186, N11182, N2557);
not NOT1 (N11187, N11178);
buf BUF1 (N11188, N11186);
buf BUF1 (N11189, N11176);
or OR2 (N11190, N11183, N7891);
not NOT1 (N11191, N11187);
xor XOR2 (N11192, N11185, N7161);
or OR3 (N11193, N11171, N5401, N1602);
and AND3 (N11194, N11174, N6180, N3530);
not NOT1 (N11195, N11194);
or OR4 (N11196, N11188, N5570, N10014, N7205);
or OR4 (N11197, N11193, N5104, N4591, N2104);
and AND3 (N11198, N11196, N9568, N1382);
not NOT1 (N11199, N11153);
nand NAND4 (N11200, N11195, N9546, N534, N815);
buf BUF1 (N11201, N11198);
nor NOR2 (N11202, N11190, N2472);
not NOT1 (N11203, N11199);
buf BUF1 (N11204, N11189);
not NOT1 (N11205, N11200);
or OR3 (N11206, N11201, N9265, N6776);
not NOT1 (N11207, N11191);
xor XOR2 (N11208, N11197, N5071);
nand NAND4 (N11209, N11184, N7951, N7367, N3226);
and AND4 (N11210, N11202, N8454, N8719, N9239);
xor XOR2 (N11211, N11192, N11042);
nand NAND3 (N11212, N11211, N757, N3699);
buf BUF1 (N11213, N11204);
xor XOR2 (N11214, N11180, N2944);
not NOT1 (N11215, N11208);
xor XOR2 (N11216, N11207, N2903);
nand NAND4 (N11217, N11210, N9476, N9480, N1969);
xor XOR2 (N11218, N11212, N10039);
not NOT1 (N11219, N11217);
or OR2 (N11220, N11203, N11203);
and AND3 (N11221, N11215, N10618, N1874);
or OR2 (N11222, N11216, N7125);
or OR2 (N11223, N11219, N11100);
not NOT1 (N11224, N11209);
not NOT1 (N11225, N11206);
nand NAND4 (N11226, N11214, N5767, N870, N2102);
and AND4 (N11227, N11213, N2181, N6688, N8554);
not NOT1 (N11228, N11225);
xor XOR2 (N11229, N11223, N1861);
buf BUF1 (N11230, N11224);
not NOT1 (N11231, N11226);
xor XOR2 (N11232, N11228, N2560);
nand NAND4 (N11233, N11221, N9267, N6196, N9616);
nor NOR2 (N11234, N11231, N6450);
nand NAND2 (N11235, N11205, N1594);
xor XOR2 (N11236, N11222, N3958);
nor NOR3 (N11237, N11233, N3954, N10651);
not NOT1 (N11238, N11235);
nand NAND3 (N11239, N11227, N10278, N3380);
buf BUF1 (N11240, N11237);
nand NAND4 (N11241, N11240, N7612, N4707, N8482);
not NOT1 (N11242, N11234);
not NOT1 (N11243, N11241);
buf BUF1 (N11244, N11230);
nand NAND2 (N11245, N11243, N4717);
and AND3 (N11246, N11238, N2753, N6133);
or OR3 (N11247, N11239, N10490, N3180);
nand NAND4 (N11248, N11232, N397, N1249, N4168);
xor XOR2 (N11249, N11248, N3472);
xor XOR2 (N11250, N11247, N9261);
and AND3 (N11251, N11249, N10677, N1990);
nor NOR4 (N11252, N11242, N5993, N11012, N8253);
and AND3 (N11253, N11218, N1960, N409);
or OR2 (N11254, N11252, N2228);
xor XOR2 (N11255, N11245, N4993);
nand NAND3 (N11256, N11250, N1016, N7485);
buf BUF1 (N11257, N11246);
xor XOR2 (N11258, N11244, N8618);
xor XOR2 (N11259, N11236, N9800);
or OR3 (N11260, N11256, N25, N4207);
nand NAND3 (N11261, N11258, N9710, N7621);
and AND2 (N11262, N11253, N4008);
buf BUF1 (N11263, N11229);
nand NAND4 (N11264, N11261, N8976, N3957, N3559);
buf BUF1 (N11265, N11263);
nand NAND3 (N11266, N11265, N1881, N4538);
nor NOR2 (N11267, N11257, N7422);
xor XOR2 (N11268, N11251, N6629);
nor NOR3 (N11269, N11260, N4265, N9980);
not NOT1 (N11270, N11254);
or OR4 (N11271, N11269, N10215, N7631, N2384);
and AND3 (N11272, N11268, N1763, N1609);
nand NAND3 (N11273, N11271, N1987, N6052);
or OR4 (N11274, N11267, N1516, N6739, N1599);
and AND4 (N11275, N11264, N1064, N3262, N6758);
and AND4 (N11276, N11262, N9168, N3529, N1549);
xor XOR2 (N11277, N11273, N4098);
buf BUF1 (N11278, N11275);
buf BUF1 (N11279, N11266);
nand NAND3 (N11280, N11274, N10513, N7839);
nor NOR3 (N11281, N11259, N8252, N3699);
nor NOR3 (N11282, N11278, N3129, N7117);
buf BUF1 (N11283, N11270);
nor NOR4 (N11284, N11255, N9740, N2315, N2234);
buf BUF1 (N11285, N11282);
xor XOR2 (N11286, N11272, N10163);
buf BUF1 (N11287, N11280);
buf BUF1 (N11288, N11279);
buf BUF1 (N11289, N11284);
not NOT1 (N11290, N11283);
nand NAND3 (N11291, N11288, N409, N3315);
xor XOR2 (N11292, N11291, N3592);
xor XOR2 (N11293, N11290, N1092);
buf BUF1 (N11294, N11286);
and AND2 (N11295, N11276, N8870);
not NOT1 (N11296, N11285);
not NOT1 (N11297, N11287);
or OR3 (N11298, N11293, N3441, N8126);
xor XOR2 (N11299, N11292, N11237);
not NOT1 (N11300, N11295);
buf BUF1 (N11301, N11294);
nor NOR4 (N11302, N11299, N11008, N6586, N8090);
nor NOR2 (N11303, N11220, N1101);
nand NAND4 (N11304, N11277, N378, N10761, N7764);
and AND2 (N11305, N11298, N7718);
not NOT1 (N11306, N11305);
not NOT1 (N11307, N11281);
buf BUF1 (N11308, N11303);
not NOT1 (N11309, N11306);
nor NOR4 (N11310, N11289, N7482, N542, N3869);
nand NAND3 (N11311, N11308, N3338, N10475);
and AND2 (N11312, N11311, N10314);
not NOT1 (N11313, N11297);
and AND4 (N11314, N11307, N4478, N1246, N7839);
not NOT1 (N11315, N11304);
buf BUF1 (N11316, N11309);
buf BUF1 (N11317, N11313);
xor XOR2 (N11318, N11316, N1097);
xor XOR2 (N11319, N11300, N9829);
xor XOR2 (N11320, N11319, N2996);
or OR4 (N11321, N11302, N8118, N3953, N6232);
and AND3 (N11322, N11315, N7325, N743);
or OR3 (N11323, N11318, N806, N6769);
not NOT1 (N11324, N11320);
xor XOR2 (N11325, N11323, N4025);
or OR3 (N11326, N11324, N1837, N1154);
nor NOR2 (N11327, N11325, N3723);
nand NAND4 (N11328, N11326, N10663, N1462, N10129);
nand NAND2 (N11329, N11317, N2697);
nor NOR2 (N11330, N11314, N1034);
and AND2 (N11331, N11296, N1735);
and AND4 (N11332, N11330, N6123, N9012, N5669);
xor XOR2 (N11333, N11327, N11280);
and AND4 (N11334, N11312, N7305, N11002, N6345);
xor XOR2 (N11335, N11332, N8377);
xor XOR2 (N11336, N11335, N1622);
and AND4 (N11337, N11336, N712, N7314, N3167);
not NOT1 (N11338, N11331);
not NOT1 (N11339, N11329);
or OR3 (N11340, N11338, N10425, N8657);
xor XOR2 (N11341, N11337, N10748);
buf BUF1 (N11342, N11333);
buf BUF1 (N11343, N11341);
and AND4 (N11344, N11328, N6548, N9133, N9722);
or OR4 (N11345, N11343, N1724, N7698, N7759);
xor XOR2 (N11346, N11334, N7781);
or OR3 (N11347, N11346, N6953, N1346);
nand NAND2 (N11348, N11344, N3076);
or OR3 (N11349, N11310, N5906, N4034);
nand NAND4 (N11350, N11322, N7739, N4160, N5960);
nand NAND3 (N11351, N11350, N3365, N6653);
not NOT1 (N11352, N11301);
and AND2 (N11353, N11351, N3462);
nor NOR3 (N11354, N11339, N6648, N4202);
nand NAND2 (N11355, N11347, N10270);
not NOT1 (N11356, N11355);
xor XOR2 (N11357, N11353, N7180);
and AND3 (N11358, N11345, N7594, N520);
not NOT1 (N11359, N11352);
or OR4 (N11360, N11340, N3778, N2325, N6941);
nand NAND2 (N11361, N11342, N116);
or OR4 (N11362, N11358, N6459, N7298, N2649);
buf BUF1 (N11363, N11349);
or OR2 (N11364, N11321, N6506);
xor XOR2 (N11365, N11362, N7330);
nand NAND3 (N11366, N11365, N10867, N2537);
not NOT1 (N11367, N11354);
buf BUF1 (N11368, N11367);
buf BUF1 (N11369, N11360);
not NOT1 (N11370, N11368);
and AND2 (N11371, N11370, N7915);
not NOT1 (N11372, N11357);
not NOT1 (N11373, N11363);
xor XOR2 (N11374, N11356, N3675);
buf BUF1 (N11375, N11348);
and AND2 (N11376, N11371, N3612);
xor XOR2 (N11377, N11359, N5368);
not NOT1 (N11378, N11374);
nor NOR3 (N11379, N11378, N7003, N10208);
xor XOR2 (N11380, N11369, N9972);
buf BUF1 (N11381, N11376);
buf BUF1 (N11382, N11372);
buf BUF1 (N11383, N11379);
not NOT1 (N11384, N11383);
nor NOR4 (N11385, N11373, N8440, N9145, N586);
and AND3 (N11386, N11366, N3333, N2474);
nor NOR3 (N11387, N11385, N2666, N9829);
or OR4 (N11388, N11375, N1749, N1585, N5882);
nand NAND3 (N11389, N11380, N735, N10663);
xor XOR2 (N11390, N11389, N251);
nor NOR4 (N11391, N11386, N843, N10061, N8769);
buf BUF1 (N11392, N11388);
or OR2 (N11393, N11377, N9923);
buf BUF1 (N11394, N11361);
and AND2 (N11395, N11387, N3572);
not NOT1 (N11396, N11384);
or OR2 (N11397, N11364, N3583);
buf BUF1 (N11398, N11382);
xor XOR2 (N11399, N11396, N4383);
and AND3 (N11400, N11394, N4311, N10152);
and AND4 (N11401, N11381, N6679, N11378, N8268);
not NOT1 (N11402, N11398);
xor XOR2 (N11403, N11391, N2718);
and AND3 (N11404, N11401, N2387, N2228);
and AND3 (N11405, N11402, N5197, N5263);
nand NAND3 (N11406, N11390, N203, N10547);
xor XOR2 (N11407, N11397, N3601);
nand NAND2 (N11408, N11405, N7998);
xor XOR2 (N11409, N11395, N1731);
nand NAND4 (N11410, N11400, N4618, N3069, N13);
or OR3 (N11411, N11399, N6980, N5049);
and AND4 (N11412, N11393, N10614, N6550, N2401);
or OR2 (N11413, N11408, N9528);
nand NAND2 (N11414, N11412, N785);
xor XOR2 (N11415, N11406, N10589);
nor NOR4 (N11416, N11392, N448, N1611, N10492);
xor XOR2 (N11417, N11410, N928);
or OR3 (N11418, N11416, N4071, N515);
not NOT1 (N11419, N11413);
or OR4 (N11420, N11418, N802, N585, N11298);
not NOT1 (N11421, N11417);
and AND4 (N11422, N11419, N5492, N3182, N2066);
or OR4 (N11423, N11420, N5524, N4378, N2470);
and AND4 (N11424, N11415, N5204, N5815, N6);
nor NOR3 (N11425, N11421, N283, N2474);
xor XOR2 (N11426, N11424, N1953);
xor XOR2 (N11427, N11409, N5168);
or OR4 (N11428, N11407, N6905, N6447, N8755);
xor XOR2 (N11429, N11428, N8320);
not NOT1 (N11430, N11422);
buf BUF1 (N11431, N11426);
and AND2 (N11432, N11414, N2763);
and AND3 (N11433, N11430, N8308, N7010);
nand NAND4 (N11434, N11403, N1295, N11110, N11054);
or OR4 (N11435, N11433, N8643, N9001, N3542);
xor XOR2 (N11436, N11411, N2371);
xor XOR2 (N11437, N11434, N9935);
xor XOR2 (N11438, N11432, N4069);
not NOT1 (N11439, N11435);
nor NOR2 (N11440, N11427, N7452);
or OR3 (N11441, N11436, N10468, N5159);
nor NOR4 (N11442, N11425, N631, N3972, N5416);
xor XOR2 (N11443, N11429, N3458);
not NOT1 (N11444, N11438);
and AND4 (N11445, N11442, N3626, N10897, N9850);
and AND4 (N11446, N11431, N6299, N10430, N3630);
buf BUF1 (N11447, N11404);
and AND4 (N11448, N11447, N10055, N5495, N11043);
or OR2 (N11449, N11445, N5066);
or OR3 (N11450, N11449, N6974, N7957);
and AND4 (N11451, N11446, N10337, N3402, N7856);
not NOT1 (N11452, N11444);
or OR2 (N11453, N11423, N4163);
and AND3 (N11454, N11451, N199, N8577);
nand NAND3 (N11455, N11437, N8790, N4919);
xor XOR2 (N11456, N11440, N5221);
nor NOR3 (N11457, N11453, N85, N1844);
or OR2 (N11458, N11443, N5590);
not NOT1 (N11459, N11458);
and AND4 (N11460, N11448, N4047, N8120, N1196);
nand NAND2 (N11461, N11452, N8618);
xor XOR2 (N11462, N11459, N2670);
or OR3 (N11463, N11461, N544, N153);
and AND2 (N11464, N11454, N6062);
not NOT1 (N11465, N11456);
nand NAND3 (N11466, N11441, N758, N9693);
not NOT1 (N11467, N11457);
nand NAND2 (N11468, N11439, N11453);
nand NAND3 (N11469, N11460, N2757, N4264);
buf BUF1 (N11470, N11455);
and AND4 (N11471, N11450, N8433, N8458, N3544);
nand NAND3 (N11472, N11465, N3820, N7498);
not NOT1 (N11473, N11468);
xor XOR2 (N11474, N11473, N5206);
buf BUF1 (N11475, N11463);
xor XOR2 (N11476, N11474, N2307);
nand NAND3 (N11477, N11472, N2589, N8632);
nor NOR2 (N11478, N11477, N4990);
nor NOR3 (N11479, N11478, N724, N294);
and AND2 (N11480, N11479, N9369);
nor NOR4 (N11481, N11469, N6705, N1905, N1829);
not NOT1 (N11482, N11480);
nand NAND2 (N11483, N11470, N9300);
nor NOR4 (N11484, N11464, N3322, N5829, N4560);
not NOT1 (N11485, N11462);
buf BUF1 (N11486, N11476);
nor NOR4 (N11487, N11481, N2471, N1082, N10783);
xor XOR2 (N11488, N11485, N10327);
or OR2 (N11489, N11471, N10466);
and AND3 (N11490, N11482, N8276, N1961);
not NOT1 (N11491, N11488);
nor NOR3 (N11492, N11484, N5793, N750);
buf BUF1 (N11493, N11491);
nor NOR4 (N11494, N11466, N10632, N10812, N8541);
buf BUF1 (N11495, N11489);
xor XOR2 (N11496, N11494, N6042);
nor NOR4 (N11497, N11495, N10804, N7687, N3389);
nand NAND3 (N11498, N11483, N7831, N5720);
nor NOR2 (N11499, N11467, N9858);
nand NAND3 (N11500, N11496, N3899, N1647);
nand NAND2 (N11501, N11497, N4033);
not NOT1 (N11502, N11475);
not NOT1 (N11503, N11498);
and AND3 (N11504, N11486, N3860, N748);
nor NOR2 (N11505, N11500, N11484);
not NOT1 (N11506, N11499);
and AND4 (N11507, N11505, N3938, N6560, N1732);
buf BUF1 (N11508, N11507);
or OR2 (N11509, N11504, N9919);
xor XOR2 (N11510, N11506, N5411);
buf BUF1 (N11511, N11502);
not NOT1 (N11512, N11492);
and AND4 (N11513, N11510, N10036, N7057, N3361);
nand NAND3 (N11514, N11509, N9580, N2386);
nand NAND4 (N11515, N11508, N2223, N8718, N8448);
or OR3 (N11516, N11487, N8893, N637);
and AND4 (N11517, N11515, N4235, N6943, N7769);
xor XOR2 (N11518, N11512, N8969);
not NOT1 (N11519, N11514);
xor XOR2 (N11520, N11490, N7148);
not NOT1 (N11521, N11493);
nand NAND2 (N11522, N11516, N1324);
or OR2 (N11523, N11521, N6587);
nor NOR4 (N11524, N11519, N7134, N470, N178);
and AND3 (N11525, N11503, N7763, N10377);
and AND4 (N11526, N11522, N8331, N7041, N4871);
nand NAND3 (N11527, N11525, N595, N4324);
not NOT1 (N11528, N11527);
nor NOR3 (N11529, N11513, N1827, N1374);
or OR4 (N11530, N11517, N6733, N10433, N8400);
and AND2 (N11531, N11529, N4147);
xor XOR2 (N11532, N11501, N3652);
or OR3 (N11533, N11511, N2741, N6393);
not NOT1 (N11534, N11528);
and AND4 (N11535, N11533, N7136, N6062, N9092);
buf BUF1 (N11536, N11524);
not NOT1 (N11537, N11531);
nor NOR3 (N11538, N11526, N7447, N5727);
or OR4 (N11539, N11535, N10378, N10650, N957);
xor XOR2 (N11540, N11538, N7755);
and AND4 (N11541, N11539, N7708, N10011, N7905);
or OR4 (N11542, N11541, N9510, N10614, N9065);
or OR2 (N11543, N11520, N9583);
not NOT1 (N11544, N11543);
or OR4 (N11545, N11523, N1230, N9496, N7869);
and AND4 (N11546, N11532, N8808, N108, N3149);
and AND3 (N11547, N11544, N10165, N3984);
not NOT1 (N11548, N11547);
nor NOR2 (N11549, N11537, N4680);
and AND2 (N11550, N11540, N2929);
or OR3 (N11551, N11518, N2503, N7871);
not NOT1 (N11552, N11545);
buf BUF1 (N11553, N11546);
xor XOR2 (N11554, N11551, N1099);
not NOT1 (N11555, N11549);
nand NAND2 (N11556, N11554, N8337);
nor NOR4 (N11557, N11550, N10558, N5973, N11544);
xor XOR2 (N11558, N11555, N9090);
not NOT1 (N11559, N11557);
nand NAND2 (N11560, N11559, N4288);
nand NAND3 (N11561, N11556, N2914, N8872);
buf BUF1 (N11562, N11548);
not NOT1 (N11563, N11562);
nor NOR3 (N11564, N11553, N8026, N3964);
nand NAND4 (N11565, N11542, N10994, N6129, N7501);
buf BUF1 (N11566, N11534);
not NOT1 (N11567, N11536);
nand NAND4 (N11568, N11566, N3844, N3260, N6226);
buf BUF1 (N11569, N11567);
xor XOR2 (N11570, N11563, N824);
xor XOR2 (N11571, N11558, N4002);
nor NOR2 (N11572, N11565, N11);
buf BUF1 (N11573, N11564);
nand NAND2 (N11574, N11561, N3357);
or OR3 (N11575, N11570, N8060, N10674);
nand NAND3 (N11576, N11530, N5588, N7012);
nand NAND3 (N11577, N11552, N6571, N7940);
buf BUF1 (N11578, N11569);
nand NAND2 (N11579, N11568, N9325);
and AND2 (N11580, N11576, N3465);
or OR2 (N11581, N11580, N3078);
and AND2 (N11582, N11574, N2470);
buf BUF1 (N11583, N11577);
and AND2 (N11584, N11583, N1504);
buf BUF1 (N11585, N11578);
buf BUF1 (N11586, N11582);
nor NOR4 (N11587, N11575, N7999, N10123, N5093);
or OR4 (N11588, N11585, N3541, N4852, N4035);
xor XOR2 (N11589, N11571, N33);
xor XOR2 (N11590, N11560, N10107);
xor XOR2 (N11591, N11579, N9273);
or OR2 (N11592, N11587, N10891);
nor NOR4 (N11593, N11589, N7841, N2494, N7219);
not NOT1 (N11594, N11592);
nor NOR3 (N11595, N11572, N2788, N3487);
and AND3 (N11596, N11591, N3934, N843);
nand NAND4 (N11597, N11594, N1558, N5436, N7648);
not NOT1 (N11598, N11573);
or OR3 (N11599, N11586, N9404, N3617);
xor XOR2 (N11600, N11598, N7320);
or OR4 (N11601, N11596, N6178, N11305, N9235);
not NOT1 (N11602, N11581);
xor XOR2 (N11603, N11601, N2932);
buf BUF1 (N11604, N11593);
buf BUF1 (N11605, N11597);
xor XOR2 (N11606, N11604, N3830);
nor NOR2 (N11607, N11590, N8822);
xor XOR2 (N11608, N11603, N7902);
nor NOR3 (N11609, N11602, N8440, N6066);
nand NAND3 (N11610, N11599, N2693, N10771);
or OR3 (N11611, N11605, N2120, N1859);
buf BUF1 (N11612, N11584);
not NOT1 (N11613, N11606);
not NOT1 (N11614, N11588);
nand NAND4 (N11615, N11614, N3043, N2479, N6640);
xor XOR2 (N11616, N11611, N4841);
nand NAND2 (N11617, N11615, N5586);
nor NOR3 (N11618, N11612, N6972, N10744);
nand NAND2 (N11619, N11617, N10620);
or OR2 (N11620, N11608, N1234);
nand NAND3 (N11621, N11595, N4840, N7908);
and AND3 (N11622, N11620, N6149, N1517);
nor NOR4 (N11623, N11613, N6157, N4362, N5676);
xor XOR2 (N11624, N11623, N76);
and AND3 (N11625, N11621, N8023, N4294);
not NOT1 (N11626, N11624);
and AND2 (N11627, N11619, N11229);
xor XOR2 (N11628, N11600, N10329);
or OR2 (N11629, N11616, N5705);
and AND2 (N11630, N11618, N8911);
nor NOR2 (N11631, N11610, N7509);
and AND2 (N11632, N11629, N3702);
buf BUF1 (N11633, N11632);
and AND2 (N11634, N11633, N1605);
and AND2 (N11635, N11630, N10254);
and AND4 (N11636, N11634, N8745, N3129, N10209);
and AND3 (N11637, N11636, N11429, N235);
nand NAND4 (N11638, N11622, N8535, N1416, N9247);
nor NOR2 (N11639, N11625, N9941);
xor XOR2 (N11640, N11639, N5518);
buf BUF1 (N11641, N11637);
and AND4 (N11642, N11609, N10874, N3500, N10609);
nor NOR3 (N11643, N11607, N9668, N5113);
nand NAND2 (N11644, N11635, N8200);
and AND4 (N11645, N11628, N8781, N7038, N3029);
nand NAND3 (N11646, N11641, N4235, N11248);
or OR2 (N11647, N11645, N8357);
and AND3 (N11648, N11640, N4259, N4778);
xor XOR2 (N11649, N11642, N6777);
nor NOR4 (N11650, N11647, N6581, N7562, N3535);
buf BUF1 (N11651, N11627);
nor NOR4 (N11652, N11649, N633, N1437, N600);
not NOT1 (N11653, N11638);
buf BUF1 (N11654, N11643);
buf BUF1 (N11655, N11644);
xor XOR2 (N11656, N11654, N6309);
xor XOR2 (N11657, N11652, N3855);
or OR2 (N11658, N11656, N3689);
and AND2 (N11659, N11653, N7626);
buf BUF1 (N11660, N11650);
xor XOR2 (N11661, N11659, N10240);
nand NAND2 (N11662, N11651, N8162);
or OR3 (N11663, N11648, N656, N1317);
not NOT1 (N11664, N11660);
nor NOR2 (N11665, N11663, N3232);
not NOT1 (N11666, N11658);
and AND3 (N11667, N11664, N2941, N2367);
or OR4 (N11668, N11626, N3931, N5003, N8649);
xor XOR2 (N11669, N11667, N9690);
buf BUF1 (N11670, N11661);
buf BUF1 (N11671, N11670);
not NOT1 (N11672, N11662);
or OR4 (N11673, N11665, N6222, N5342, N1507);
or OR4 (N11674, N11646, N10614, N8535, N7161);
and AND4 (N11675, N11672, N9066, N7841, N1490);
and AND3 (N11676, N11668, N3974, N2506);
and AND4 (N11677, N11674, N8045, N8443, N7937);
not NOT1 (N11678, N11631);
not NOT1 (N11679, N11676);
buf BUF1 (N11680, N11657);
nand NAND3 (N11681, N11669, N10848, N6424);
buf BUF1 (N11682, N11677);
xor XOR2 (N11683, N11655, N9206);
nand NAND3 (N11684, N11666, N7726, N257);
not NOT1 (N11685, N11675);
nor NOR2 (N11686, N11685, N10387);
xor XOR2 (N11687, N11681, N8638);
xor XOR2 (N11688, N11678, N10891);
or OR3 (N11689, N11673, N2810, N4269);
buf BUF1 (N11690, N11683);
buf BUF1 (N11691, N11690);
buf BUF1 (N11692, N11680);
or OR4 (N11693, N11692, N9351, N7640, N8491);
or OR3 (N11694, N11691, N4756, N5015);
nand NAND3 (N11695, N11686, N1384, N10641);
nand NAND3 (N11696, N11693, N10689, N3225);
or OR4 (N11697, N11671, N1921, N8648, N6416);
nand NAND2 (N11698, N11689, N6487);
or OR3 (N11699, N11687, N10841, N7462);
nand NAND4 (N11700, N11698, N3164, N1019, N10215);
xor XOR2 (N11701, N11684, N10853);
nor NOR2 (N11702, N11688, N967);
xor XOR2 (N11703, N11700, N8386);
and AND4 (N11704, N11695, N4779, N1289, N4297);
or OR4 (N11705, N11702, N1809, N5027, N5630);
buf BUF1 (N11706, N11705);
nor NOR3 (N11707, N11694, N4661, N5645);
xor XOR2 (N11708, N11679, N3);
nor NOR4 (N11709, N11703, N5462, N2165, N3026);
nand NAND4 (N11710, N11682, N3440, N10399, N7890);
and AND3 (N11711, N11696, N9801, N9027);
nor NOR2 (N11712, N11699, N8732);
nand NAND4 (N11713, N11709, N8430, N8787, N10984);
or OR2 (N11714, N11710, N3815);
nand NAND3 (N11715, N11712, N780, N7161);
or OR4 (N11716, N11706, N11348, N1341, N5871);
and AND2 (N11717, N11714, N1725);
xor XOR2 (N11718, N11715, N982);
not NOT1 (N11719, N11697);
not NOT1 (N11720, N11704);
buf BUF1 (N11721, N11701);
not NOT1 (N11722, N11713);
and AND3 (N11723, N11721, N56, N1598);
buf BUF1 (N11724, N11717);
buf BUF1 (N11725, N11722);
buf BUF1 (N11726, N11711);
xor XOR2 (N11727, N11725, N2792);
not NOT1 (N11728, N11727);
buf BUF1 (N11729, N11707);
not NOT1 (N11730, N11719);
nor NOR4 (N11731, N11720, N10396, N6151, N3005);
nor NOR2 (N11732, N11716, N4759);
and AND2 (N11733, N11723, N6773);
and AND2 (N11734, N11724, N3071);
nor NOR3 (N11735, N11729, N3028, N11679);
and AND3 (N11736, N11734, N3007, N6218);
not NOT1 (N11737, N11726);
nand NAND4 (N11738, N11730, N781, N66, N6336);
not NOT1 (N11739, N11738);
and AND2 (N11740, N11732, N1268);
nor NOR4 (N11741, N11736, N9716, N9512, N8857);
nand NAND2 (N11742, N11708, N2319);
nor NOR4 (N11743, N11739, N1284, N2527, N368);
buf BUF1 (N11744, N11742);
buf BUF1 (N11745, N11728);
or OR4 (N11746, N11741, N7053, N7400, N7092);
nand NAND2 (N11747, N11743, N2952);
nand NAND2 (N11748, N11731, N5731);
nand NAND2 (N11749, N11735, N4692);
or OR4 (N11750, N11737, N1695, N9358, N10367);
not NOT1 (N11751, N11744);
nor NOR3 (N11752, N11748, N244, N7);
nor NOR3 (N11753, N11752, N11092, N10389);
nor NOR2 (N11754, N11753, N8254);
and AND4 (N11755, N11718, N1679, N361, N7755);
and AND3 (N11756, N11733, N1165, N9777);
not NOT1 (N11757, N11755);
xor XOR2 (N11758, N11745, N2596);
or OR2 (N11759, N11740, N9405);
xor XOR2 (N11760, N11757, N8363);
and AND2 (N11761, N11746, N3993);
nor NOR4 (N11762, N11761, N8475, N7486, N11230);
nand NAND4 (N11763, N11749, N4938, N5142, N6128);
xor XOR2 (N11764, N11751, N10505);
nor NOR2 (N11765, N11754, N3952);
or OR4 (N11766, N11747, N2580, N9880, N7506);
buf BUF1 (N11767, N11763);
nor NOR2 (N11768, N11767, N3727);
xor XOR2 (N11769, N11768, N7399);
buf BUF1 (N11770, N11756);
nor NOR2 (N11771, N11770, N10180);
or OR3 (N11772, N11764, N8381, N6392);
nand NAND4 (N11773, N11750, N3348, N3448, N8758);
xor XOR2 (N11774, N11773, N4736);
nand NAND4 (N11775, N11762, N1255, N1967, N2472);
or OR3 (N11776, N11769, N3842, N7490);
not NOT1 (N11777, N11766);
or OR4 (N11778, N11775, N11457, N5970, N7658);
nand NAND3 (N11779, N11777, N1879, N6682);
or OR4 (N11780, N11776, N4034, N5501, N6921);
xor XOR2 (N11781, N11774, N2156);
nor NOR2 (N11782, N11781, N10459);
and AND3 (N11783, N11780, N3706, N8941);
and AND3 (N11784, N11779, N6807, N903);
nand NAND4 (N11785, N11772, N9541, N2617, N2278);
and AND2 (N11786, N11778, N3003);
nor NOR4 (N11787, N11765, N11730, N595, N967);
and AND2 (N11788, N11787, N11420);
not NOT1 (N11789, N11760);
xor XOR2 (N11790, N11789, N8967);
nand NAND2 (N11791, N11782, N7481);
nand NAND3 (N11792, N11786, N8675, N10630);
buf BUF1 (N11793, N11785);
or OR2 (N11794, N11758, N1463);
nand NAND2 (N11795, N11794, N5106);
not NOT1 (N11796, N11783);
or OR3 (N11797, N11793, N63, N6691);
xor XOR2 (N11798, N11784, N1872);
nor NOR3 (N11799, N11791, N8862, N6170);
nor NOR2 (N11800, N11795, N2714);
not NOT1 (N11801, N11792);
xor XOR2 (N11802, N11799, N6445);
buf BUF1 (N11803, N11797);
not NOT1 (N11804, N11803);
xor XOR2 (N11805, N11801, N5959);
and AND4 (N11806, N11805, N8973, N8705, N5213);
not NOT1 (N11807, N11802);
not NOT1 (N11808, N11800);
or OR2 (N11809, N11759, N2210);
not NOT1 (N11810, N11807);
nor NOR2 (N11811, N11790, N1410);
or OR3 (N11812, N11788, N9813, N5106);
buf BUF1 (N11813, N11798);
nand NAND3 (N11814, N11804, N9006, N11127);
xor XOR2 (N11815, N11812, N11806);
xor XOR2 (N11816, N578, N1387);
and AND4 (N11817, N11796, N1054, N5408, N9619);
or OR3 (N11818, N11811, N6003, N9042);
and AND4 (N11819, N11818, N3727, N3117, N6570);
nor NOR3 (N11820, N11815, N6006, N10378);
or OR4 (N11821, N11813, N7935, N534, N9130);
and AND3 (N11822, N11771, N2641, N826);
xor XOR2 (N11823, N11808, N4022);
buf BUF1 (N11824, N11816);
buf BUF1 (N11825, N11810);
and AND4 (N11826, N11823, N5030, N3341, N5713);
not NOT1 (N11827, N11824);
xor XOR2 (N11828, N11820, N6375);
buf BUF1 (N11829, N11822);
nor NOR3 (N11830, N11826, N2845, N6772);
buf BUF1 (N11831, N11827);
xor XOR2 (N11832, N11828, N9710);
or OR2 (N11833, N11825, N1951);
not NOT1 (N11834, N11832);
and AND3 (N11835, N11809, N1354, N6672);
buf BUF1 (N11836, N11831);
and AND3 (N11837, N11819, N8492, N2567);
and AND2 (N11838, N11835, N7620);
or OR3 (N11839, N11821, N5198, N10341);
nand NAND2 (N11840, N11833, N6413);
nand NAND4 (N11841, N11814, N8824, N2773, N9036);
xor XOR2 (N11842, N11841, N2008);
xor XOR2 (N11843, N11817, N8691);
or OR4 (N11844, N11838, N981, N9614, N10223);
not NOT1 (N11845, N11830);
not NOT1 (N11846, N11843);
and AND3 (N11847, N11834, N8567, N8507);
not NOT1 (N11848, N11837);
and AND2 (N11849, N11829, N3483);
and AND3 (N11850, N11836, N6969, N4099);
or OR3 (N11851, N11840, N480, N6889);
not NOT1 (N11852, N11851);
xor XOR2 (N11853, N11849, N7999);
xor XOR2 (N11854, N11850, N10585);
or OR3 (N11855, N11844, N5377, N11538);
nor NOR4 (N11856, N11852, N9380, N11220, N9938);
or OR2 (N11857, N11845, N8172);
xor XOR2 (N11858, N11839, N5014);
nor NOR4 (N11859, N11853, N4994, N10417, N1892);
and AND2 (N11860, N11855, N8336);
nand NAND4 (N11861, N11848, N1593, N7777, N7487);
nor NOR4 (N11862, N11861, N4148, N331, N8330);
nand NAND4 (N11863, N11857, N5277, N2258, N1051);
buf BUF1 (N11864, N11847);
not NOT1 (N11865, N11846);
nand NAND4 (N11866, N11858, N2159, N8162, N6675);
xor XOR2 (N11867, N11865, N7498);
not NOT1 (N11868, N11864);
nor NOR2 (N11869, N11867, N5595);
nand NAND2 (N11870, N11868, N1089);
or OR4 (N11871, N11862, N4753, N6485, N3281);
nand NAND3 (N11872, N11870, N5638, N2203);
buf BUF1 (N11873, N11869);
or OR3 (N11874, N11842, N5212, N8040);
xor XOR2 (N11875, N11873, N5034);
and AND4 (N11876, N11856, N1946, N6760, N382);
or OR4 (N11877, N11863, N8159, N2572, N8906);
or OR3 (N11878, N11859, N9666, N1824);
or OR2 (N11879, N11854, N3481);
not NOT1 (N11880, N11875);
nand NAND3 (N11881, N11880, N3289, N680);
buf BUF1 (N11882, N11872);
xor XOR2 (N11883, N11878, N3204);
and AND3 (N11884, N11877, N7235, N3959);
xor XOR2 (N11885, N11860, N5191);
or OR3 (N11886, N11883, N9342, N2909);
not NOT1 (N11887, N11876);
xor XOR2 (N11888, N11871, N7915);
not NOT1 (N11889, N11881);
nor NOR4 (N11890, N11879, N2729, N1097, N4441);
or OR3 (N11891, N11874, N10623, N1556);
nor NOR2 (N11892, N11891, N1923);
nor NOR2 (N11893, N11890, N11291);
nor NOR3 (N11894, N11882, N1916, N1006);
not NOT1 (N11895, N11884);
not NOT1 (N11896, N11866);
or OR4 (N11897, N11885, N1382, N8241, N3078);
or OR4 (N11898, N11892, N2271, N7120, N2658);
nor NOR3 (N11899, N11898, N11561, N9162);
nor NOR3 (N11900, N11893, N8649, N8939);
nand NAND3 (N11901, N11894, N167, N2018);
not NOT1 (N11902, N11897);
or OR3 (N11903, N11895, N1804, N4568);
xor XOR2 (N11904, N11889, N11040);
xor XOR2 (N11905, N11888, N6224);
xor XOR2 (N11906, N11902, N260);
or OR3 (N11907, N11904, N6988, N1945);
xor XOR2 (N11908, N11906, N3714);
or OR2 (N11909, N11908, N4141);
and AND3 (N11910, N11905, N2757, N10967);
xor XOR2 (N11911, N11903, N9449);
xor XOR2 (N11912, N11900, N7470);
buf BUF1 (N11913, N11896);
nor NOR4 (N11914, N11912, N3056, N10414, N6560);
or OR4 (N11915, N11886, N2683, N2392, N2561);
and AND3 (N11916, N11911, N6966, N4162);
buf BUF1 (N11917, N11910);
xor XOR2 (N11918, N11909, N3273);
or OR2 (N11919, N11918, N550);
not NOT1 (N11920, N11917);
not NOT1 (N11921, N11913);
not NOT1 (N11922, N11921);
not NOT1 (N11923, N11922);
not NOT1 (N11924, N11901);
xor XOR2 (N11925, N11899, N7883);
buf BUF1 (N11926, N11915);
not NOT1 (N11927, N11920);
not NOT1 (N11928, N11907);
or OR3 (N11929, N11926, N5496, N7372);
or OR2 (N11930, N11919, N5638);
xor XOR2 (N11931, N11887, N9532);
and AND4 (N11932, N11916, N6510, N4024, N621);
not NOT1 (N11933, N11932);
or OR3 (N11934, N11914, N7617, N763);
nor NOR4 (N11935, N11925, N7404, N3771, N9098);
nor NOR2 (N11936, N11931, N5656);
and AND4 (N11937, N11935, N5840, N10665, N4826);
and AND4 (N11938, N11936, N9113, N11528, N9724);
buf BUF1 (N11939, N11929);
nand NAND4 (N11940, N11933, N4402, N4712, N7306);
nand NAND2 (N11941, N11928, N4194);
buf BUF1 (N11942, N11934);
nand NAND2 (N11943, N11939, N6507);
nor NOR4 (N11944, N11941, N4499, N11708, N5355);
xor XOR2 (N11945, N11943, N8106);
not NOT1 (N11946, N11927);
and AND2 (N11947, N11945, N2348);
nor NOR2 (N11948, N11923, N81);
and AND3 (N11949, N11938, N602, N3590);
nor NOR3 (N11950, N11924, N11232, N7738);
and AND2 (N11951, N11947, N6042);
xor XOR2 (N11952, N11930, N10278);
nand NAND2 (N11953, N11950, N5340);
buf BUF1 (N11954, N11937);
xor XOR2 (N11955, N11940, N751);
not NOT1 (N11956, N11944);
and AND3 (N11957, N11952, N8671, N1845);
buf BUF1 (N11958, N11951);
and AND2 (N11959, N11953, N8195);
nor NOR2 (N11960, N11946, N2012);
nor NOR4 (N11961, N11960, N3661, N2338, N10019);
not NOT1 (N11962, N11948);
nand NAND2 (N11963, N11956, N3591);
nor NOR2 (N11964, N11954, N7447);
buf BUF1 (N11965, N11955);
nand NAND3 (N11966, N11961, N7467, N4942);
or OR3 (N11967, N11963, N9054, N107);
xor XOR2 (N11968, N11966, N10781);
buf BUF1 (N11969, N11968);
not NOT1 (N11970, N11965);
not NOT1 (N11971, N11957);
and AND3 (N11972, N11969, N11905, N11097);
nand NAND3 (N11973, N11970, N3706, N10483);
buf BUF1 (N11974, N11971);
not NOT1 (N11975, N11949);
nand NAND4 (N11976, N11959, N4607, N8068, N9145);
and AND4 (N11977, N11976, N6075, N7356, N788);
and AND4 (N11978, N11973, N7457, N5441, N6991);
nor NOR4 (N11979, N11964, N3516, N9670, N7935);
and AND4 (N11980, N11979, N1263, N7970, N2840);
not NOT1 (N11981, N11974);
and AND2 (N11982, N11977, N1398);
not NOT1 (N11983, N11942);
and AND3 (N11984, N11972, N8866, N10071);
nand NAND3 (N11985, N11984, N9578, N6412);
and AND4 (N11986, N11958, N10793, N797, N7900);
or OR4 (N11987, N11986, N10041, N9595, N7091);
nor NOR3 (N11988, N11978, N9255, N9629);
not NOT1 (N11989, N11985);
or OR4 (N11990, N11980, N5949, N5653, N3745);
or OR4 (N11991, N11981, N9531, N1499, N2277);
or OR2 (N11992, N11967, N1445);
nand NAND4 (N11993, N11962, N8119, N3827, N11150);
and AND4 (N11994, N11990, N6814, N8987, N11451);
nand NAND3 (N11995, N11989, N7433, N4678);
buf BUF1 (N11996, N11983);
and AND3 (N11997, N11992, N1414, N5671);
buf BUF1 (N11998, N11996);
xor XOR2 (N11999, N11994, N8048);
nor NOR4 (N12000, N11991, N6315, N10308, N2804);
or OR3 (N12001, N11975, N3906, N7822);
not NOT1 (N12002, N11999);
xor XOR2 (N12003, N11995, N4496);
not NOT1 (N12004, N11998);
or OR3 (N12005, N11993, N1257, N2983);
xor XOR2 (N12006, N12000, N8889);
nand NAND4 (N12007, N11982, N5486, N7013, N2017);
not NOT1 (N12008, N12002);
or OR2 (N12009, N12008, N5840);
nand NAND4 (N12010, N12003, N3518, N2035, N8772);
not NOT1 (N12011, N12005);
and AND2 (N12012, N11988, N8222);
nand NAND3 (N12013, N12007, N6850, N6687);
nand NAND2 (N12014, N12006, N3879);
nor NOR3 (N12015, N12001, N4345, N11311);
or OR2 (N12016, N12012, N2766);
nor NOR3 (N12017, N12013, N8810, N9886);
or OR4 (N12018, N12004, N3511, N6463, N4006);
buf BUF1 (N12019, N12009);
nand NAND3 (N12020, N11987, N6418, N4002);
nor NOR4 (N12021, N12019, N3871, N4625, N1319);
nor NOR4 (N12022, N12021, N2625, N3955, N1878);
xor XOR2 (N12023, N12010, N4609);
nor NOR2 (N12024, N11997, N1686);
nand NAND4 (N12025, N12023, N695, N5658, N3156);
buf BUF1 (N12026, N12015);
buf BUF1 (N12027, N12022);
nor NOR2 (N12028, N12016, N3232);
not NOT1 (N12029, N12011);
not NOT1 (N12030, N12025);
nand NAND3 (N12031, N12014, N5238, N10359);
or OR3 (N12032, N12030, N4511, N1089);
xor XOR2 (N12033, N12028, N5816);
xor XOR2 (N12034, N12018, N5516);
xor XOR2 (N12035, N12024, N6352);
xor XOR2 (N12036, N12020, N9707);
and AND4 (N12037, N12035, N4106, N11935, N7408);
nand NAND3 (N12038, N12026, N5037, N4397);
not NOT1 (N12039, N12027);
and AND2 (N12040, N12033, N8302);
nor NOR2 (N12041, N12017, N4781);
or OR3 (N12042, N12039, N10050, N945);
and AND2 (N12043, N12038, N5793);
xor XOR2 (N12044, N12029, N769);
xor XOR2 (N12045, N12036, N9631);
nor NOR2 (N12046, N12034, N1433);
xor XOR2 (N12047, N12041, N1843);
and AND2 (N12048, N12032, N6903);
xor XOR2 (N12049, N12043, N5555);
xor XOR2 (N12050, N12047, N8876);
buf BUF1 (N12051, N12045);
not NOT1 (N12052, N12040);
nor NOR4 (N12053, N12049, N9942, N1837, N11756);
nand NAND3 (N12054, N12051, N11930, N10019);
nor NOR4 (N12055, N12037, N2982, N5807, N6527);
and AND3 (N12056, N12050, N4475, N11420);
or OR2 (N12057, N12048, N148);
xor XOR2 (N12058, N12042, N1240);
not NOT1 (N12059, N12058);
nor NOR2 (N12060, N12054, N10659);
buf BUF1 (N12061, N12052);
or OR3 (N12062, N12060, N5364, N9094);
not NOT1 (N12063, N12056);
buf BUF1 (N12064, N12046);
or OR2 (N12065, N12057, N2902);
xor XOR2 (N12066, N12064, N8868);
buf BUF1 (N12067, N12053);
and AND2 (N12068, N12055, N2197);
nor NOR3 (N12069, N12044, N1638, N1319);
nand NAND4 (N12070, N12061, N1301, N9994, N8524);
nand NAND4 (N12071, N12068, N6535, N8573, N8220);
xor XOR2 (N12072, N12065, N8172);
and AND3 (N12073, N12071, N3776, N738);
and AND4 (N12074, N12069, N4494, N2617, N10175);
not NOT1 (N12075, N12059);
nand NAND3 (N12076, N12070, N4553, N11022);
xor XOR2 (N12077, N12031, N8900);
nand NAND3 (N12078, N12063, N5949, N4020);
and AND3 (N12079, N12072, N11234, N3780);
nand NAND4 (N12080, N12066, N6143, N10764, N8913);
nor NOR3 (N12081, N12067, N3785, N10161);
nand NAND2 (N12082, N12079, N9629);
xor XOR2 (N12083, N12078, N1405);
not NOT1 (N12084, N12077);
not NOT1 (N12085, N12083);
xor XOR2 (N12086, N12075, N3682);
or OR2 (N12087, N12074, N9564);
and AND4 (N12088, N12082, N6664, N830, N563);
nand NAND2 (N12089, N12086, N10529);
buf BUF1 (N12090, N12084);
nor NOR4 (N12091, N12073, N5316, N4400, N6434);
or OR3 (N12092, N12089, N11892, N4014);
not NOT1 (N12093, N12080);
nor NOR2 (N12094, N12088, N6364);
not NOT1 (N12095, N12076);
and AND3 (N12096, N12094, N5274, N3766);
not NOT1 (N12097, N12087);
nor NOR4 (N12098, N12081, N8887, N1399, N6888);
or OR4 (N12099, N12092, N11193, N3186, N9011);
not NOT1 (N12100, N12062);
xor XOR2 (N12101, N12098, N7368);
xor XOR2 (N12102, N12099, N219);
xor XOR2 (N12103, N12093, N8785);
and AND2 (N12104, N12091, N2429);
nor NOR3 (N12105, N12103, N8995, N1197);
nor NOR2 (N12106, N12102, N268);
xor XOR2 (N12107, N12105, N7801);
nand NAND4 (N12108, N12096, N10973, N3491, N11544);
nand NAND4 (N12109, N12095, N9261, N6337, N6776);
xor XOR2 (N12110, N12107, N850);
nor NOR3 (N12111, N12085, N6978, N9683);
and AND4 (N12112, N12104, N10893, N3258, N11295);
and AND4 (N12113, N12101, N4926, N5180, N9285);
xor XOR2 (N12114, N12100, N10250);
nor NOR3 (N12115, N12109, N727, N54);
and AND2 (N12116, N12090, N2668);
or OR3 (N12117, N12110, N3717, N3278);
nand NAND3 (N12118, N12114, N11063, N5946);
not NOT1 (N12119, N12116);
nand NAND2 (N12120, N12118, N7597);
or OR3 (N12121, N12115, N8132, N6809);
buf BUF1 (N12122, N12097);
and AND3 (N12123, N12121, N5858, N5932);
and AND4 (N12124, N12106, N8604, N1851, N11696);
xor XOR2 (N12125, N12117, N6787);
buf BUF1 (N12126, N12124);
buf BUF1 (N12127, N12111);
buf BUF1 (N12128, N12112);
buf BUF1 (N12129, N12119);
xor XOR2 (N12130, N12113, N9781);
or OR3 (N12131, N12122, N3559, N1533);
and AND2 (N12132, N12108, N1192);
xor XOR2 (N12133, N12129, N7346);
xor XOR2 (N12134, N12127, N8793);
not NOT1 (N12135, N12125);
nand NAND2 (N12136, N12123, N3870);
buf BUF1 (N12137, N12133);
nand NAND3 (N12138, N12131, N7660, N2581);
or OR4 (N12139, N12128, N3379, N649, N6482);
nor NOR2 (N12140, N12136, N2283);
not NOT1 (N12141, N12126);
or OR4 (N12142, N12135, N770, N5787, N2764);
and AND2 (N12143, N12130, N10002);
not NOT1 (N12144, N12141);
nand NAND4 (N12145, N12132, N6509, N11218, N668);
xor XOR2 (N12146, N12145, N9616);
nand NAND3 (N12147, N12137, N12037, N5890);
not NOT1 (N12148, N12139);
not NOT1 (N12149, N12134);
and AND4 (N12150, N12143, N9869, N2463, N3706);
xor XOR2 (N12151, N12148, N10827);
nor NOR4 (N12152, N12142, N10188, N1006, N9631);
not NOT1 (N12153, N12149);
or OR4 (N12154, N12140, N2138, N4144, N5673);
not NOT1 (N12155, N12120);
and AND4 (N12156, N12155, N6292, N532, N9453);
nor NOR2 (N12157, N12154, N3243);
xor XOR2 (N12158, N12151, N4965);
xor XOR2 (N12159, N12138, N11851);
or OR4 (N12160, N12144, N9173, N11676, N7265);
xor XOR2 (N12161, N12160, N2356);
not NOT1 (N12162, N12147);
xor XOR2 (N12163, N12152, N11);
nand NAND4 (N12164, N12162, N4770, N4746, N8374);
buf BUF1 (N12165, N12158);
or OR4 (N12166, N12165, N6339, N4298, N2174);
xor XOR2 (N12167, N12166, N10623);
nor NOR3 (N12168, N12150, N2674, N5391);
or OR4 (N12169, N12156, N11835, N9850, N11494);
xor XOR2 (N12170, N12164, N2022);
nand NAND2 (N12171, N12157, N6845);
or OR4 (N12172, N12169, N1872, N10045, N10389);
buf BUF1 (N12173, N12159);
and AND4 (N12174, N12168, N4367, N2147, N9707);
or OR3 (N12175, N12173, N6628, N1312);
buf BUF1 (N12176, N12163);
nor NOR2 (N12177, N12171, N7108);
or OR3 (N12178, N12146, N4395, N4452);
nand NAND2 (N12179, N12178, N823);
nand NAND3 (N12180, N12177, N5713, N3231);
xor XOR2 (N12181, N12167, N10413);
xor XOR2 (N12182, N12174, N11008);
or OR2 (N12183, N12176, N7227);
nor NOR3 (N12184, N12183, N714, N10246);
buf BUF1 (N12185, N12179);
nand NAND4 (N12186, N12161, N9992, N5800, N11341);
nor NOR4 (N12187, N12181, N5852, N2578, N12139);
not NOT1 (N12188, N12180);
buf BUF1 (N12189, N12187);
buf BUF1 (N12190, N12185);
and AND3 (N12191, N12188, N3334, N5438);
buf BUF1 (N12192, N12191);
nor NOR4 (N12193, N12170, N8516, N2, N117);
nand NAND4 (N12194, N12192, N10948, N635, N8623);
not NOT1 (N12195, N12186);
or OR4 (N12196, N12195, N674, N2152, N9156);
not NOT1 (N12197, N12196);
not NOT1 (N12198, N12193);
xor XOR2 (N12199, N12172, N1518);
xor XOR2 (N12200, N12197, N9050);
or OR3 (N12201, N12184, N5949, N4719);
nor NOR4 (N12202, N12182, N11086, N5635, N2505);
nor NOR4 (N12203, N12194, N2379, N10000, N1059);
xor XOR2 (N12204, N12199, N11428);
and AND3 (N12205, N12175, N10154, N6829);
buf BUF1 (N12206, N12198);
and AND2 (N12207, N12201, N9434);
not NOT1 (N12208, N12200);
not NOT1 (N12209, N12204);
not NOT1 (N12210, N12203);
buf BUF1 (N12211, N12208);
buf BUF1 (N12212, N12207);
nor NOR4 (N12213, N12202, N3047, N2975, N3548);
xor XOR2 (N12214, N12205, N8331);
buf BUF1 (N12215, N12210);
and AND2 (N12216, N12213, N6904);
buf BUF1 (N12217, N12215);
not NOT1 (N12218, N12153);
xor XOR2 (N12219, N12216, N807);
buf BUF1 (N12220, N12211);
or OR2 (N12221, N12219, N7937);
xor XOR2 (N12222, N12206, N1712);
xor XOR2 (N12223, N12221, N4783);
nor NOR2 (N12224, N12217, N9346);
buf BUF1 (N12225, N12224);
nor NOR4 (N12226, N12189, N5809, N9508, N2458);
not NOT1 (N12227, N12223);
nand NAND4 (N12228, N12218, N1283, N10327, N7035);
nor NOR3 (N12229, N12190, N9818, N4085);
or OR4 (N12230, N12229, N6423, N9213, N5299);
xor XOR2 (N12231, N12220, N6099);
xor XOR2 (N12232, N12225, N9691);
and AND3 (N12233, N12222, N6692, N5376);
and AND3 (N12234, N12232, N8357, N9681);
and AND2 (N12235, N12234, N9271);
nand NAND4 (N12236, N12212, N11032, N3231, N5102);
nand NAND3 (N12237, N12228, N164, N9528);
not NOT1 (N12238, N12235);
nor NOR4 (N12239, N12209, N3897, N9147, N3796);
xor XOR2 (N12240, N12214, N5546);
or OR2 (N12241, N12231, N8184);
buf BUF1 (N12242, N12230);
or OR3 (N12243, N12241, N8455, N8881);
and AND3 (N12244, N12227, N976, N2860);
or OR4 (N12245, N12243, N3099, N4054, N7612);
xor XOR2 (N12246, N12237, N10403);
or OR2 (N12247, N12238, N11728);
nand NAND3 (N12248, N12240, N9066, N8454);
nand NAND3 (N12249, N12246, N1802, N10523);
not NOT1 (N12250, N12242);
nand NAND4 (N12251, N12249, N8440, N10972, N7043);
not NOT1 (N12252, N12233);
nor NOR3 (N12253, N12226, N1045, N10782);
or OR3 (N12254, N12239, N6556, N9483);
or OR4 (N12255, N12252, N4293, N1604, N6940);
nor NOR3 (N12256, N12254, N12145, N1003);
xor XOR2 (N12257, N12244, N7168);
nand NAND4 (N12258, N12255, N5681, N3448, N6868);
not NOT1 (N12259, N12256);
and AND3 (N12260, N12257, N6286, N4015);
nor NOR4 (N12261, N12260, N4099, N7408, N2833);
nand NAND3 (N12262, N12247, N6541, N5425);
and AND2 (N12263, N12259, N4291);
and AND3 (N12264, N12258, N473, N10972);
nor NOR3 (N12265, N12261, N9800, N6916);
not NOT1 (N12266, N12236);
and AND4 (N12267, N12251, N2508, N2501, N3853);
xor XOR2 (N12268, N12263, N7441);
or OR4 (N12269, N12248, N9774, N4323, N2845);
buf BUF1 (N12270, N12264);
buf BUF1 (N12271, N12253);
nor NOR3 (N12272, N12271, N11782, N11519);
xor XOR2 (N12273, N12266, N12131);
nor NOR4 (N12274, N12267, N1750, N8734, N1185);
and AND4 (N12275, N12262, N5314, N5096, N9412);
buf BUF1 (N12276, N12270);
and AND3 (N12277, N12272, N3697, N1376);
nor NOR4 (N12278, N12274, N1529, N6998, N8863);
nor NOR2 (N12279, N12268, N7210);
nand NAND3 (N12280, N12245, N9112, N1323);
or OR2 (N12281, N12277, N5595);
nand NAND3 (N12282, N12265, N6995, N3838);
or OR2 (N12283, N12282, N3417);
nand NAND4 (N12284, N12279, N11980, N2307, N11368);
nor NOR2 (N12285, N12281, N7379);
not NOT1 (N12286, N12250);
nor NOR2 (N12287, N12284, N5700);
nor NOR4 (N12288, N12283, N6082, N2037, N11967);
not NOT1 (N12289, N12278);
and AND4 (N12290, N12273, N1845, N2720, N1855);
and AND3 (N12291, N12287, N2219, N2982);
nor NOR2 (N12292, N12269, N8320);
or OR2 (N12293, N12290, N7932);
nand NAND2 (N12294, N12285, N2674);
nand NAND2 (N12295, N12286, N10229);
nand NAND3 (N12296, N12292, N6088, N3381);
buf BUF1 (N12297, N12296);
and AND2 (N12298, N12289, N4914);
nand NAND2 (N12299, N12295, N3905);
xor XOR2 (N12300, N12297, N1821);
and AND4 (N12301, N12298, N7145, N6825, N2686);
and AND4 (N12302, N12299, N4263, N4844, N3067);
nand NAND2 (N12303, N12276, N11178);
and AND3 (N12304, N12288, N10775, N3594);
or OR4 (N12305, N12291, N6989, N9294, N1740);
and AND4 (N12306, N12294, N3767, N7020, N6727);
not NOT1 (N12307, N12305);
buf BUF1 (N12308, N12304);
nand NAND4 (N12309, N12308, N8425, N9175, N3680);
not NOT1 (N12310, N12303);
nor NOR4 (N12311, N12306, N11407, N1385, N7954);
xor XOR2 (N12312, N12311, N8583);
nand NAND3 (N12313, N12300, N1064, N1073);
or OR4 (N12314, N12312, N7846, N3215, N4702);
and AND2 (N12315, N12275, N11745);
xor XOR2 (N12316, N12314, N3580);
nor NOR4 (N12317, N12307, N4253, N404, N2806);
or OR2 (N12318, N12316, N2977);
or OR2 (N12319, N12317, N6292);
xor XOR2 (N12320, N12310, N563);
or OR3 (N12321, N12318, N4539, N10803);
not NOT1 (N12322, N12280);
nand NAND3 (N12323, N12301, N5337, N2196);
or OR4 (N12324, N12302, N2617, N5992, N10032);
not NOT1 (N12325, N12293);
or OR4 (N12326, N12313, N7326, N5886, N6658);
buf BUF1 (N12327, N12322);
not NOT1 (N12328, N12320);
nor NOR2 (N12329, N12324, N3920);
not NOT1 (N12330, N12326);
or OR3 (N12331, N12323, N1430, N354);
xor XOR2 (N12332, N12329, N7896);
nand NAND3 (N12333, N12325, N6218, N11464);
or OR3 (N12334, N12328, N10003, N7359);
buf BUF1 (N12335, N12319);
or OR4 (N12336, N12327, N7346, N347, N3560);
buf BUF1 (N12337, N12331);
buf BUF1 (N12338, N12315);
nand NAND3 (N12339, N12337, N11710, N10634);
nand NAND4 (N12340, N12330, N7000, N9680, N3695);
buf BUF1 (N12341, N12338);
xor XOR2 (N12342, N12341, N3994);
and AND3 (N12343, N12339, N3701, N6306);
nand NAND4 (N12344, N12321, N1764, N6232, N10652);
xor XOR2 (N12345, N12332, N6553);
not NOT1 (N12346, N12340);
buf BUF1 (N12347, N12342);
buf BUF1 (N12348, N12336);
buf BUF1 (N12349, N12334);
or OR4 (N12350, N12349, N4349, N4927, N3304);
nor NOR3 (N12351, N12309, N5386, N5434);
not NOT1 (N12352, N12333);
not NOT1 (N12353, N12345);
or OR3 (N12354, N12352, N919, N11760);
nor NOR3 (N12355, N12350, N2221, N8466);
and AND3 (N12356, N12348, N701, N10445);
and AND2 (N12357, N12335, N740);
xor XOR2 (N12358, N12353, N10943);
and AND3 (N12359, N12356, N6320, N10619);
buf BUF1 (N12360, N12354);
xor XOR2 (N12361, N12347, N467);
not NOT1 (N12362, N12360);
xor XOR2 (N12363, N12358, N8067);
not NOT1 (N12364, N12361);
nand NAND3 (N12365, N12362, N7673, N11656);
or OR2 (N12366, N12344, N1234);
nand NAND4 (N12367, N12365, N11655, N5594, N5581);
xor XOR2 (N12368, N12346, N7108);
or OR4 (N12369, N12368, N8639, N6564, N7277);
buf BUF1 (N12370, N12355);
nor NOR4 (N12371, N12367, N7752, N9323, N10081);
nand NAND3 (N12372, N12363, N8096, N7157);
nand NAND2 (N12373, N12351, N2371);
or OR3 (N12374, N12364, N8003, N2843);
nand NAND2 (N12375, N12359, N1722);
buf BUF1 (N12376, N12374);
nand NAND4 (N12377, N12366, N4944, N10795, N9889);
nand NAND3 (N12378, N12372, N1007, N4276);
not NOT1 (N12379, N12373);
or OR4 (N12380, N12357, N2336, N7396, N8301);
buf BUF1 (N12381, N12377);
nand NAND3 (N12382, N12370, N6667, N4536);
xor XOR2 (N12383, N12379, N7108);
not NOT1 (N12384, N12371);
nand NAND4 (N12385, N12380, N8253, N4051, N374);
buf BUF1 (N12386, N12384);
and AND2 (N12387, N12343, N10602);
not NOT1 (N12388, N12387);
nor NOR4 (N12389, N12375, N1165, N6618, N1895);
nand NAND4 (N12390, N12383, N1281, N4677, N1350);
buf BUF1 (N12391, N12369);
not NOT1 (N12392, N12385);
not NOT1 (N12393, N12388);
buf BUF1 (N12394, N12392);
and AND4 (N12395, N12390, N4654, N9264, N650);
xor XOR2 (N12396, N12386, N11584);
and AND3 (N12397, N12394, N2651, N11237);
and AND3 (N12398, N12378, N8074, N11095);
or OR3 (N12399, N12396, N12356, N3856);
nand NAND4 (N12400, N12393, N2863, N244, N7441);
xor XOR2 (N12401, N12389, N3720);
and AND2 (N12402, N12395, N10267);
nand NAND2 (N12403, N12397, N7839);
xor XOR2 (N12404, N12391, N10805);
nand NAND2 (N12405, N12402, N8483);
nor NOR4 (N12406, N12400, N11977, N7358, N6486);
nand NAND3 (N12407, N12398, N3701, N6355);
xor XOR2 (N12408, N12401, N3722);
and AND4 (N12409, N12405, N1648, N7546, N1582);
nand NAND2 (N12410, N12403, N11916);
not NOT1 (N12411, N12410);
buf BUF1 (N12412, N12407);
nand NAND2 (N12413, N12411, N10098);
nor NOR3 (N12414, N12382, N7839, N2406);
or OR3 (N12415, N12413, N527, N1711);
nor NOR3 (N12416, N12412, N8460, N439);
or OR2 (N12417, N12408, N8303);
and AND3 (N12418, N12409, N5911, N8882);
and AND3 (N12419, N12414, N9575, N4717);
nand NAND3 (N12420, N12404, N3258, N1794);
nor NOR2 (N12421, N12381, N8632);
and AND4 (N12422, N12416, N5602, N7570, N11161);
nand NAND2 (N12423, N12419, N7307);
or OR4 (N12424, N12420, N12030, N4836, N9241);
buf BUF1 (N12425, N12423);
nor NOR3 (N12426, N12422, N7477, N316);
nand NAND3 (N12427, N12417, N928, N229);
not NOT1 (N12428, N12421);
buf BUF1 (N12429, N12376);
buf BUF1 (N12430, N12415);
nor NOR2 (N12431, N12399, N3615);
buf BUF1 (N12432, N12431);
and AND2 (N12433, N12425, N12421);
and AND4 (N12434, N12429, N3956, N4312, N10310);
xor XOR2 (N12435, N12406, N9356);
buf BUF1 (N12436, N12432);
buf BUF1 (N12437, N12424);
nand NAND2 (N12438, N12437, N11855);
and AND2 (N12439, N12433, N5927);
nand NAND4 (N12440, N12436, N11571, N5046, N1596);
or OR4 (N12441, N12426, N3228, N2990, N10851);
and AND2 (N12442, N12430, N7115);
nand NAND2 (N12443, N12442, N5713);
xor XOR2 (N12444, N12434, N1039);
buf BUF1 (N12445, N12441);
nor NOR2 (N12446, N12418, N2245);
not NOT1 (N12447, N12440);
or OR2 (N12448, N12447, N8000);
buf BUF1 (N12449, N12444);
nand NAND2 (N12450, N12428, N5998);
or OR4 (N12451, N12446, N574, N349, N1104);
or OR3 (N12452, N12448, N8962, N816);
nor NOR3 (N12453, N12450, N1937, N6219);
nor NOR2 (N12454, N12445, N9373);
buf BUF1 (N12455, N12435);
xor XOR2 (N12456, N12438, N3910);
nor NOR4 (N12457, N12427, N5782, N9576, N1100);
not NOT1 (N12458, N12449);
nand NAND2 (N12459, N12457, N8180);
nand NAND3 (N12460, N12439, N11507, N4070);
buf BUF1 (N12461, N12458);
nor NOR4 (N12462, N12452, N10809, N11443, N3832);
nor NOR4 (N12463, N12443, N9265, N3661, N5420);
xor XOR2 (N12464, N12451, N12205);
not NOT1 (N12465, N12461);
buf BUF1 (N12466, N12464);
not NOT1 (N12467, N12463);
nand NAND4 (N12468, N12462, N9947, N5143, N2032);
nand NAND3 (N12469, N12454, N8733, N7357);
buf BUF1 (N12470, N12466);
nand NAND2 (N12471, N12455, N12142);
xor XOR2 (N12472, N12471, N9969);
buf BUF1 (N12473, N12460);
not NOT1 (N12474, N12470);
xor XOR2 (N12475, N12469, N1155);
and AND4 (N12476, N12467, N498, N10759, N9653);
or OR4 (N12477, N12465, N3139, N6400, N9941);
and AND3 (N12478, N12475, N5375, N3640);
nand NAND2 (N12479, N12473, N2091);
nor NOR2 (N12480, N12479, N2865);
xor XOR2 (N12481, N12456, N8118);
not NOT1 (N12482, N12481);
and AND2 (N12483, N12472, N9225);
nor NOR3 (N12484, N12478, N11440, N7136);
nand NAND3 (N12485, N12482, N1754, N1905);
and AND2 (N12486, N12459, N2274);
nor NOR4 (N12487, N12486, N3370, N4854, N9719);
xor XOR2 (N12488, N12468, N6831);
or OR2 (N12489, N12485, N6665);
buf BUF1 (N12490, N12453);
xor XOR2 (N12491, N12480, N10991);
or OR4 (N12492, N12477, N6808, N1524, N6720);
nor NOR2 (N12493, N12489, N11101);
not NOT1 (N12494, N12487);
or OR4 (N12495, N12474, N4169, N6940, N1881);
buf BUF1 (N12496, N12476);
and AND2 (N12497, N12483, N7050);
nor NOR3 (N12498, N12490, N7539, N2979);
not NOT1 (N12499, N12496);
nand NAND3 (N12500, N12498, N4712, N4017);
nor NOR4 (N12501, N12484, N5531, N5723, N11058);
not NOT1 (N12502, N12488);
buf BUF1 (N12503, N12497);
nor NOR3 (N12504, N12501, N6175, N3440);
and AND2 (N12505, N12504, N3150);
nand NAND2 (N12506, N12502, N2101);
and AND2 (N12507, N12493, N1755);
nor NOR3 (N12508, N12506, N11768, N2937);
and AND2 (N12509, N12494, N639);
or OR2 (N12510, N12492, N10207);
nand NAND3 (N12511, N12503, N9983, N11855);
nor NOR4 (N12512, N12508, N4431, N56, N8043);
or OR4 (N12513, N12495, N8466, N4420, N7599);
nor NOR2 (N12514, N12505, N1592);
not NOT1 (N12515, N12509);
nand NAND2 (N12516, N12491, N783);
not NOT1 (N12517, N12499);
buf BUF1 (N12518, N12512);
buf BUF1 (N12519, N12518);
not NOT1 (N12520, N12511);
buf BUF1 (N12521, N12500);
and AND4 (N12522, N12516, N9539, N12333, N2113);
nor NOR3 (N12523, N12510, N7409, N2197);
buf BUF1 (N12524, N12513);
nand NAND2 (N12525, N12521, N5105);
nor NOR2 (N12526, N12523, N12151);
and AND4 (N12527, N12520, N9273, N549, N1260);
nand NAND2 (N12528, N12515, N9276);
or OR4 (N12529, N12517, N3968, N8015, N904);
and AND4 (N12530, N12519, N4230, N7721, N627);
nor NOR3 (N12531, N12530, N10475, N1185);
or OR2 (N12532, N12526, N11703);
and AND3 (N12533, N12524, N3287, N5317);
or OR2 (N12534, N12529, N11819);
and AND2 (N12535, N12525, N2822);
not NOT1 (N12536, N12533);
not NOT1 (N12537, N12532);
not NOT1 (N12538, N12537);
xor XOR2 (N12539, N12522, N5698);
not NOT1 (N12540, N12531);
nor NOR2 (N12541, N12536, N10377);
not NOT1 (N12542, N12541);
buf BUF1 (N12543, N12539);
buf BUF1 (N12544, N12543);
buf BUF1 (N12545, N12528);
or OR3 (N12546, N12544, N10183, N7725);
and AND4 (N12547, N12514, N4852, N3334, N10940);
buf BUF1 (N12548, N12546);
xor XOR2 (N12549, N12534, N9600);
buf BUF1 (N12550, N12527);
not NOT1 (N12551, N12550);
nand NAND2 (N12552, N12551, N4505);
nand NAND3 (N12553, N12538, N10913, N2088);
xor XOR2 (N12554, N12540, N10758);
and AND3 (N12555, N12553, N4772, N7150);
nor NOR4 (N12556, N12552, N3033, N1382, N3823);
and AND4 (N12557, N12549, N10296, N8459, N1462);
xor XOR2 (N12558, N12557, N3939);
nand NAND3 (N12559, N12545, N10051, N7690);
xor XOR2 (N12560, N12554, N10803);
nor NOR2 (N12561, N12560, N6573);
or OR4 (N12562, N12547, N1458, N1714, N2462);
and AND2 (N12563, N12558, N1358);
not NOT1 (N12564, N12556);
buf BUF1 (N12565, N12563);
not NOT1 (N12566, N12555);
xor XOR2 (N12567, N12548, N10601);
xor XOR2 (N12568, N12535, N2320);
xor XOR2 (N12569, N12562, N598);
and AND4 (N12570, N12507, N4111, N8032, N7764);
not NOT1 (N12571, N12559);
not NOT1 (N12572, N12571);
not NOT1 (N12573, N12567);
and AND2 (N12574, N12564, N1858);
and AND3 (N12575, N12574, N6217, N6697);
and AND4 (N12576, N12572, N7154, N6349, N5808);
not NOT1 (N12577, N12568);
nor NOR2 (N12578, N12577, N3236);
xor XOR2 (N12579, N12578, N451);
or OR4 (N12580, N12575, N8115, N12139, N5248);
or OR4 (N12581, N12566, N4189, N7722, N11259);
or OR2 (N12582, N12581, N3164);
nand NAND2 (N12583, N12565, N900);
buf BUF1 (N12584, N12561);
not NOT1 (N12585, N12570);
not NOT1 (N12586, N12583);
or OR4 (N12587, N12580, N9302, N2468, N2191);
buf BUF1 (N12588, N12579);
not NOT1 (N12589, N12585);
buf BUF1 (N12590, N12573);
nor NOR2 (N12591, N12586, N5305);
nand NAND3 (N12592, N12587, N4434, N5521);
not NOT1 (N12593, N12569);
buf BUF1 (N12594, N12590);
and AND3 (N12595, N12591, N8341, N451);
nor NOR2 (N12596, N12589, N9295);
nand NAND4 (N12597, N12592, N4619, N4871, N9258);
and AND4 (N12598, N12582, N10191, N7292, N7713);
xor XOR2 (N12599, N12598, N6637);
nor NOR4 (N12600, N12588, N6379, N11859, N841);
buf BUF1 (N12601, N12542);
nand NAND2 (N12602, N12597, N10695);
or OR4 (N12603, N12584, N11177, N3474, N10345);
or OR2 (N12604, N12600, N9282);
and AND3 (N12605, N12593, N6590, N9190);
nor NOR3 (N12606, N12599, N7010, N9374);
xor XOR2 (N12607, N12602, N11968);
not NOT1 (N12608, N12607);
buf BUF1 (N12609, N12605);
and AND2 (N12610, N12594, N3062);
nor NOR2 (N12611, N12595, N3032);
xor XOR2 (N12612, N12596, N8443);
nand NAND3 (N12613, N12609, N1173, N6033);
xor XOR2 (N12614, N12603, N11680);
nand NAND4 (N12615, N12601, N1024, N11096, N6417);
and AND2 (N12616, N12613, N10185);
not NOT1 (N12617, N12606);
not NOT1 (N12618, N12608);
nand NAND4 (N12619, N12611, N7955, N3423, N12301);
buf BUF1 (N12620, N12610);
not NOT1 (N12621, N12615);
and AND2 (N12622, N12620, N7920);
xor XOR2 (N12623, N12619, N3616);
and AND3 (N12624, N12618, N11551, N9116);
buf BUF1 (N12625, N12624);
xor XOR2 (N12626, N12621, N2692);
and AND2 (N12627, N12604, N2937);
or OR2 (N12628, N12616, N8479);
buf BUF1 (N12629, N12576);
buf BUF1 (N12630, N12629);
buf BUF1 (N12631, N12630);
nor NOR2 (N12632, N12612, N89);
and AND4 (N12633, N12625, N6289, N2169, N1710);
nand NAND3 (N12634, N12622, N2108, N3064);
or OR4 (N12635, N12623, N859, N614, N10864);
nor NOR2 (N12636, N12635, N1984);
not NOT1 (N12637, N12626);
xor XOR2 (N12638, N12614, N1794);
and AND2 (N12639, N12634, N3331);
nor NOR2 (N12640, N12637, N2003);
nand NAND4 (N12641, N12631, N11379, N6171, N8473);
xor XOR2 (N12642, N12641, N6425);
xor XOR2 (N12643, N12638, N2019);
xor XOR2 (N12644, N12636, N9248);
nor NOR2 (N12645, N12617, N4332);
xor XOR2 (N12646, N12627, N10379);
xor XOR2 (N12647, N12645, N2723);
xor XOR2 (N12648, N12628, N12326);
or OR2 (N12649, N12647, N832);
nor NOR2 (N12650, N12643, N2872);
not NOT1 (N12651, N12648);
not NOT1 (N12652, N12639);
nand NAND3 (N12653, N12652, N5038, N9345);
not NOT1 (N12654, N12649);
or OR3 (N12655, N12651, N6446, N9563);
buf BUF1 (N12656, N12640);
nand NAND4 (N12657, N12646, N10751, N8287, N9382);
buf BUF1 (N12658, N12655);
nand NAND2 (N12659, N12658, N5828);
or OR4 (N12660, N12650, N3569, N4350, N9728);
nor NOR4 (N12661, N12656, N11562, N4372, N11841);
nor NOR4 (N12662, N12653, N5191, N3734, N1933);
xor XOR2 (N12663, N12632, N4334);
and AND2 (N12664, N12644, N2864);
buf BUF1 (N12665, N12642);
not NOT1 (N12666, N12659);
buf BUF1 (N12667, N12666);
buf BUF1 (N12668, N12663);
nand NAND2 (N12669, N12664, N11246);
and AND2 (N12670, N12669, N7643);
buf BUF1 (N12671, N12654);
buf BUF1 (N12672, N12633);
xor XOR2 (N12673, N12662, N11113);
nand NAND2 (N12674, N12671, N5984);
buf BUF1 (N12675, N12672);
not NOT1 (N12676, N12660);
or OR2 (N12677, N12661, N7149);
and AND4 (N12678, N12674, N3902, N5004, N3558);
buf BUF1 (N12679, N12657);
or OR2 (N12680, N12676, N4711);
nand NAND3 (N12681, N12673, N11065, N1835);
and AND2 (N12682, N12668, N6674);
or OR4 (N12683, N12670, N395, N11248, N6257);
buf BUF1 (N12684, N12667);
nand NAND3 (N12685, N12680, N12295, N1900);
buf BUF1 (N12686, N12684);
not NOT1 (N12687, N12679);
buf BUF1 (N12688, N12678);
not NOT1 (N12689, N12681);
buf BUF1 (N12690, N12677);
buf BUF1 (N12691, N12683);
nand NAND2 (N12692, N12687, N12586);
nor NOR2 (N12693, N12665, N12539);
xor XOR2 (N12694, N12693, N4339);
and AND2 (N12695, N12689, N12083);
not NOT1 (N12696, N12686);
xor XOR2 (N12697, N12695, N10177);
buf BUF1 (N12698, N12696);
nand NAND2 (N12699, N12692, N10223);
xor XOR2 (N12700, N12694, N1642);
nor NOR4 (N12701, N12691, N10789, N5142, N10072);
nor NOR2 (N12702, N12700, N11503);
not NOT1 (N12703, N12688);
nor NOR4 (N12704, N12690, N12693, N8431, N351);
buf BUF1 (N12705, N12682);
nand NAND3 (N12706, N12699, N12243, N2291);
nand NAND2 (N12707, N12698, N2106);
not NOT1 (N12708, N12702);
xor XOR2 (N12709, N12708, N8949);
or OR4 (N12710, N12705, N469, N11765, N4229);
not NOT1 (N12711, N12707);
nand NAND3 (N12712, N12710, N7486, N3304);
not NOT1 (N12713, N12703);
not NOT1 (N12714, N12709);
and AND4 (N12715, N12675, N12316, N2507, N3899);
xor XOR2 (N12716, N12712, N7500);
xor XOR2 (N12717, N12685, N8394);
or OR3 (N12718, N12714, N5050, N7231);
buf BUF1 (N12719, N12701);
buf BUF1 (N12720, N12713);
buf BUF1 (N12721, N12711);
or OR2 (N12722, N12704, N2336);
nor NOR4 (N12723, N12697, N3463, N10046, N750);
nor NOR4 (N12724, N12717, N4518, N180, N11294);
buf BUF1 (N12725, N12722);
nor NOR2 (N12726, N12716, N1356);
and AND4 (N12727, N12721, N4043, N2806, N2561);
and AND2 (N12728, N12723, N9423);
not NOT1 (N12729, N12724);
xor XOR2 (N12730, N12715, N5972);
buf BUF1 (N12731, N12728);
and AND2 (N12732, N12729, N2164);
and AND3 (N12733, N12720, N11277, N5855);
buf BUF1 (N12734, N12733);
or OR4 (N12735, N12706, N1123, N1852, N8346);
nand NAND4 (N12736, N12735, N7436, N3567, N4914);
and AND2 (N12737, N12732, N11488);
or OR2 (N12738, N12734, N12405);
not NOT1 (N12739, N12727);
nand NAND4 (N12740, N12738, N4401, N4984, N12427);
nand NAND2 (N12741, N12718, N5760);
nand NAND4 (N12742, N12719, N7331, N7172, N959);
nand NAND2 (N12743, N12739, N298);
nand NAND4 (N12744, N12742, N11103, N465, N3004);
nand NAND2 (N12745, N12744, N2371);
and AND4 (N12746, N12737, N7846, N3737, N12542);
not NOT1 (N12747, N12730);
or OR2 (N12748, N12740, N7063);
nand NAND2 (N12749, N12741, N8355);
and AND3 (N12750, N12731, N691, N8599);
and AND2 (N12751, N12726, N12154);
xor XOR2 (N12752, N12746, N168);
or OR2 (N12753, N12743, N7838);
nand NAND3 (N12754, N12752, N11887, N1136);
xor XOR2 (N12755, N12747, N9185);
nand NAND2 (N12756, N12754, N10187);
xor XOR2 (N12757, N12750, N4211);
nor NOR2 (N12758, N12745, N12705);
not NOT1 (N12759, N12749);
xor XOR2 (N12760, N12753, N2054);
xor XOR2 (N12761, N12736, N10919);
xor XOR2 (N12762, N12760, N5743);
and AND4 (N12763, N12762, N9841, N12737, N12399);
buf BUF1 (N12764, N12751);
nor NOR2 (N12765, N12763, N10424);
or OR3 (N12766, N12756, N10282, N7297);
buf BUF1 (N12767, N12755);
nand NAND2 (N12768, N12765, N9155);
not NOT1 (N12769, N12761);
and AND2 (N12770, N12748, N9289);
or OR3 (N12771, N12757, N5970, N12597);
nand NAND2 (N12772, N12764, N5043);
not NOT1 (N12773, N12758);
xor XOR2 (N12774, N12770, N5248);
nor NOR2 (N12775, N12759, N7941);
nor NOR3 (N12776, N12725, N8077, N3558);
nor NOR3 (N12777, N12776, N7185, N5095);
nor NOR2 (N12778, N12767, N7763);
buf BUF1 (N12779, N12778);
nand NAND2 (N12780, N12771, N11864);
xor XOR2 (N12781, N12774, N11732);
xor XOR2 (N12782, N12777, N2920);
not NOT1 (N12783, N12775);
not NOT1 (N12784, N12782);
or OR2 (N12785, N12766, N6203);
xor XOR2 (N12786, N12768, N1348);
buf BUF1 (N12787, N12773);
nor NOR4 (N12788, N12785, N1292, N8429, N3389);
buf BUF1 (N12789, N12772);
nand NAND2 (N12790, N12783, N3394);
not NOT1 (N12791, N12788);
or OR3 (N12792, N12790, N4944, N8321);
xor XOR2 (N12793, N12780, N3181);
nand NAND4 (N12794, N12791, N3187, N3548, N6164);
or OR3 (N12795, N12784, N2984, N4394);
nand NAND4 (N12796, N12781, N560, N2752, N1401);
xor XOR2 (N12797, N12792, N2512);
not NOT1 (N12798, N12795);
or OR4 (N12799, N12793, N559, N5917, N12433);
not NOT1 (N12800, N12786);
nand NAND3 (N12801, N12799, N10895, N232);
nor NOR4 (N12802, N12798, N10294, N12431, N813);
nand NAND3 (N12803, N12797, N3854, N3215);
not NOT1 (N12804, N12779);
nand NAND2 (N12805, N12804, N4175);
buf BUF1 (N12806, N12803);
not NOT1 (N12807, N12789);
xor XOR2 (N12808, N12794, N11699);
not NOT1 (N12809, N12808);
xor XOR2 (N12810, N12809, N7266);
xor XOR2 (N12811, N12787, N1635);
xor XOR2 (N12812, N12811, N2823);
nand NAND2 (N12813, N12805, N9592);
xor XOR2 (N12814, N12796, N970);
or OR2 (N12815, N12806, N2379);
not NOT1 (N12816, N12812);
xor XOR2 (N12817, N12800, N12622);
nor NOR4 (N12818, N12813, N1815, N9685, N257);
and AND2 (N12819, N12817, N8351);
and AND2 (N12820, N12819, N1888);
xor XOR2 (N12821, N12807, N12456);
and AND2 (N12822, N12821, N10603);
or OR3 (N12823, N12802, N10416, N7963);
buf BUF1 (N12824, N12818);
not NOT1 (N12825, N12824);
not NOT1 (N12826, N12822);
or OR4 (N12827, N12769, N10034, N7638, N2756);
or OR3 (N12828, N12825, N12666, N10115);
and AND4 (N12829, N12828, N4548, N1877, N10567);
buf BUF1 (N12830, N12801);
xor XOR2 (N12831, N12823, N5343);
not NOT1 (N12832, N12815);
and AND2 (N12833, N12826, N12621);
nand NAND2 (N12834, N12832, N10565);
nand NAND4 (N12835, N12829, N10070, N2495, N4102);
not NOT1 (N12836, N12816);
nor NOR4 (N12837, N12827, N10885, N8902, N4361);
nand NAND3 (N12838, N12836, N5116, N2017);
xor XOR2 (N12839, N12835, N553);
nor NOR2 (N12840, N12833, N4106);
buf BUF1 (N12841, N12840);
or OR3 (N12842, N12810, N484, N11396);
and AND3 (N12843, N12837, N12148, N2694);
buf BUF1 (N12844, N12838);
buf BUF1 (N12845, N12842);
and AND2 (N12846, N12845, N10975);
nor NOR4 (N12847, N12834, N6755, N12239, N10628);
buf BUF1 (N12848, N12820);
not NOT1 (N12849, N12843);
nor NOR2 (N12850, N12839, N5347);
nor NOR4 (N12851, N12850, N9794, N8073, N1155);
buf BUF1 (N12852, N12814);
and AND2 (N12853, N12849, N3284);
not NOT1 (N12854, N12846);
xor XOR2 (N12855, N12851, N9437);
xor XOR2 (N12856, N12841, N2349);
xor XOR2 (N12857, N12830, N3717);
xor XOR2 (N12858, N12854, N9838);
xor XOR2 (N12859, N12852, N5046);
nor NOR3 (N12860, N12848, N10106, N11619);
or OR3 (N12861, N12831, N7234, N3131);
nand NAND4 (N12862, N12856, N176, N5858, N5727);
buf BUF1 (N12863, N12861);
buf BUF1 (N12864, N12858);
nand NAND4 (N12865, N12857, N2627, N3524, N8605);
or OR4 (N12866, N12865, N5101, N9540, N37);
xor XOR2 (N12867, N12844, N10741);
nand NAND3 (N12868, N12847, N574, N8160);
xor XOR2 (N12869, N12853, N12719);
not NOT1 (N12870, N12855);
or OR3 (N12871, N12859, N2437, N818);
buf BUF1 (N12872, N12862);
nor NOR3 (N12873, N12868, N11408, N5223);
and AND3 (N12874, N12867, N7802, N4633);
xor XOR2 (N12875, N12872, N10732);
and AND3 (N12876, N12874, N4113, N6868);
buf BUF1 (N12877, N12876);
and AND2 (N12878, N12860, N4650);
nand NAND4 (N12879, N12873, N10029, N12302, N658);
nand NAND4 (N12880, N12869, N516, N4290, N5515);
nand NAND4 (N12881, N12866, N9929, N4486, N12370);
nand NAND4 (N12882, N12875, N1578, N8984, N807);
buf BUF1 (N12883, N12880);
or OR4 (N12884, N12864, N4421, N5011, N4831);
or OR2 (N12885, N12870, N3475);
nor NOR4 (N12886, N12882, N1916, N6105, N2251);
nor NOR2 (N12887, N12878, N3198);
buf BUF1 (N12888, N12887);
nand NAND3 (N12889, N12883, N6988, N9191);
or OR3 (N12890, N12879, N8255, N1848);
nor NOR2 (N12891, N12877, N12448);
not NOT1 (N12892, N12889);
or OR3 (N12893, N12863, N5911, N10583);
not NOT1 (N12894, N12881);
nand NAND3 (N12895, N12871, N8065, N9256);
buf BUF1 (N12896, N12886);
xor XOR2 (N12897, N12892, N5978);
or OR2 (N12898, N12897, N6177);
and AND4 (N12899, N12893, N2824, N6941, N8920);
not NOT1 (N12900, N12896);
nand NAND4 (N12901, N12894, N9339, N10148, N2087);
buf BUF1 (N12902, N12885);
and AND3 (N12903, N12888, N428, N12015);
buf BUF1 (N12904, N12903);
and AND2 (N12905, N12898, N4996);
nand NAND2 (N12906, N12904, N4246);
nand NAND3 (N12907, N12895, N12127, N1176);
nand NAND4 (N12908, N12902, N1697, N12300, N8973);
xor XOR2 (N12909, N12899, N649);
not NOT1 (N12910, N12890);
and AND2 (N12911, N12910, N3442);
not NOT1 (N12912, N12906);
and AND2 (N12913, N12912, N4075);
xor XOR2 (N12914, N12901, N7659);
not NOT1 (N12915, N12884);
nand NAND2 (N12916, N12913, N4048);
xor XOR2 (N12917, N12905, N9605);
nor NOR2 (N12918, N12907, N7845);
xor XOR2 (N12919, N12900, N10030);
and AND3 (N12920, N12919, N9428, N7810);
nand NAND3 (N12921, N12918, N11644, N12191);
nor NOR2 (N12922, N12914, N6723);
xor XOR2 (N12923, N12915, N3126);
buf BUF1 (N12924, N12916);
and AND3 (N12925, N12921, N10981, N1483);
not NOT1 (N12926, N12924);
nand NAND3 (N12927, N12891, N6545, N5882);
nor NOR4 (N12928, N12925, N11890, N4023, N5160);
or OR4 (N12929, N12922, N2427, N2024, N4312);
xor XOR2 (N12930, N12909, N4227);
xor XOR2 (N12931, N12929, N2585);
xor XOR2 (N12932, N12931, N597);
buf BUF1 (N12933, N12927);
and AND3 (N12934, N12911, N9636, N1730);
nand NAND3 (N12935, N12908, N434, N6023);
nor NOR2 (N12936, N12923, N7548);
not NOT1 (N12937, N12932);
nor NOR4 (N12938, N12934, N1695, N2388, N996);
or OR4 (N12939, N12937, N9134, N8510, N2216);
not NOT1 (N12940, N12933);
xor XOR2 (N12941, N12930, N4808);
not NOT1 (N12942, N12928);
and AND2 (N12943, N12939, N5809);
xor XOR2 (N12944, N12917, N11638);
nor NOR2 (N12945, N12926, N1889);
nor NOR2 (N12946, N12942, N11280);
and AND4 (N12947, N12936, N2428, N1957, N7844);
or OR2 (N12948, N12920, N3970);
xor XOR2 (N12949, N12938, N12647);
xor XOR2 (N12950, N12947, N9589);
nor NOR2 (N12951, N12935, N82);
not NOT1 (N12952, N12941);
nand NAND3 (N12953, N12945, N7460, N2804);
nor NOR4 (N12954, N12948, N7342, N2661, N5242);
or OR2 (N12955, N12944, N3886);
not NOT1 (N12956, N12950);
or OR3 (N12957, N12953, N7281, N7535);
xor XOR2 (N12958, N12946, N12436);
buf BUF1 (N12959, N12955);
not NOT1 (N12960, N12952);
or OR4 (N12961, N12951, N2831, N10481, N4607);
not NOT1 (N12962, N12949);
not NOT1 (N12963, N12958);
not NOT1 (N12964, N12956);
or OR2 (N12965, N12954, N4743);
nor NOR4 (N12966, N12962, N12574, N392, N11478);
buf BUF1 (N12967, N12963);
xor XOR2 (N12968, N12943, N4734);
xor XOR2 (N12969, N12957, N11279);
not NOT1 (N12970, N12968);
buf BUF1 (N12971, N12961);
buf BUF1 (N12972, N12970);
nor NOR4 (N12973, N12967, N8614, N11260, N4111);
and AND3 (N12974, N12969, N10836, N2117);
and AND3 (N12975, N12966, N10232, N5925);
xor XOR2 (N12976, N12972, N7);
and AND3 (N12977, N12974, N12616, N3138);
xor XOR2 (N12978, N12959, N6827);
or OR3 (N12979, N12960, N3515, N149);
nor NOR2 (N12980, N12973, N2394);
buf BUF1 (N12981, N12978);
nor NOR2 (N12982, N12971, N5760);
buf BUF1 (N12983, N12965);
or OR2 (N12984, N12979, N1422);
xor XOR2 (N12985, N12983, N1424);
buf BUF1 (N12986, N12982);
nand NAND4 (N12987, N12986, N10003, N11135, N10856);
not NOT1 (N12988, N12940);
nor NOR2 (N12989, N12975, N2204);
and AND3 (N12990, N12989, N8902, N10723);
xor XOR2 (N12991, N12990, N4491);
and AND4 (N12992, N12981, N866, N11606, N10896);
nand NAND3 (N12993, N12985, N3930, N6692);
not NOT1 (N12994, N12988);
nor NOR4 (N12995, N12992, N8342, N12619, N246);
xor XOR2 (N12996, N12993, N3165);
xor XOR2 (N12997, N12995, N3613);
xor XOR2 (N12998, N12980, N9916);
and AND4 (N12999, N12991, N5847, N3207, N1258);
nor NOR2 (N13000, N12996, N133);
nor NOR3 (N13001, N12997, N3401, N8544);
not NOT1 (N13002, N12987);
or OR3 (N13003, N12984, N3379, N3927);
nor NOR4 (N13004, N12998, N11518, N6065, N3865);
buf BUF1 (N13005, N12999);
xor XOR2 (N13006, N13005, N4539);
buf BUF1 (N13007, N12964);
nand NAND4 (N13008, N12994, N8872, N23, N8461);
xor XOR2 (N13009, N13006, N11221);
or OR4 (N13010, N13009, N3813, N5773, N9652);
xor XOR2 (N13011, N13002, N7919);
xor XOR2 (N13012, N13004, N2371);
or OR4 (N13013, N13003, N263, N11001, N1785);
and AND3 (N13014, N13011, N1177, N10492);
nand NAND4 (N13015, N13014, N2806, N4909, N5531);
nand NAND2 (N13016, N13010, N8462);
or OR3 (N13017, N13000, N618, N173);
or OR4 (N13018, N12977, N11557, N8138, N2925);
nor NOR4 (N13019, N13012, N2484, N361, N2418);
or OR3 (N13020, N13018, N5805, N9475);
xor XOR2 (N13021, N13015, N8336);
xor XOR2 (N13022, N12976, N7393);
nand NAND4 (N13023, N13007, N8573, N3768, N4653);
xor XOR2 (N13024, N13020, N10033);
xor XOR2 (N13025, N13022, N842);
nor NOR4 (N13026, N13025, N8673, N12483, N4310);
xor XOR2 (N13027, N13021, N5546);
or OR3 (N13028, N13023, N6993, N4482);
xor XOR2 (N13029, N13028, N2589);
xor XOR2 (N13030, N13013, N10447);
xor XOR2 (N13031, N13024, N12162);
or OR3 (N13032, N13017, N6483, N12109);
and AND2 (N13033, N13001, N9465);
and AND4 (N13034, N13008, N8119, N9995, N11371);
xor XOR2 (N13035, N13016, N12603);
nor NOR4 (N13036, N13031, N5611, N599, N2718);
nor NOR2 (N13037, N13033, N6226);
and AND4 (N13038, N13030, N8008, N3964, N2444);
and AND4 (N13039, N13029, N5435, N1421, N7316);
not NOT1 (N13040, N13037);
nor NOR4 (N13041, N13039, N3085, N465, N6742);
nand NAND4 (N13042, N13026, N8879, N11456, N8208);
xor XOR2 (N13043, N13038, N4062);
nand NAND2 (N13044, N13043, N5820);
xor XOR2 (N13045, N13032, N12805);
nor NOR3 (N13046, N13036, N1450, N5642);
or OR2 (N13047, N13034, N201);
nor NOR4 (N13048, N13042, N7117, N317, N7116);
buf BUF1 (N13049, N13046);
nand NAND2 (N13050, N13048, N5634);
buf BUF1 (N13051, N13040);
buf BUF1 (N13052, N13027);
and AND3 (N13053, N13019, N3290, N2573);
buf BUF1 (N13054, N13047);
nor NOR3 (N13055, N13035, N1729, N7759);
and AND3 (N13056, N13050, N7726, N6114);
buf BUF1 (N13057, N13049);
or OR2 (N13058, N13041, N7370);
or OR3 (N13059, N13053, N7518, N2274);
nor NOR3 (N13060, N13058, N11832, N12787);
or OR4 (N13061, N13052, N153, N6335, N6206);
or OR2 (N13062, N13057, N7674);
or OR2 (N13063, N13054, N12247);
nand NAND3 (N13064, N13060, N5433, N4037);
and AND4 (N13065, N13051, N4844, N3719, N494);
not NOT1 (N13066, N13064);
and AND2 (N13067, N13045, N8040);
xor XOR2 (N13068, N13067, N4098);
and AND3 (N13069, N13066, N7726, N8856);
nor NOR4 (N13070, N13056, N9270, N9156, N3610);
not NOT1 (N13071, N13062);
nor NOR3 (N13072, N13071, N9527, N8558);
not NOT1 (N13073, N13068);
nand NAND2 (N13074, N13059, N5379);
buf BUF1 (N13075, N13072);
or OR2 (N13076, N13061, N11484);
xor XOR2 (N13077, N13073, N1776);
and AND3 (N13078, N13063, N4901, N10381);
or OR2 (N13079, N13074, N8368);
not NOT1 (N13080, N13076);
nand NAND3 (N13081, N13065, N10281, N12795);
nand NAND2 (N13082, N13055, N2736);
not NOT1 (N13083, N13080);
or OR2 (N13084, N13070, N3190);
or OR2 (N13085, N13082, N8143);
not NOT1 (N13086, N13069);
not NOT1 (N13087, N13086);
not NOT1 (N13088, N13077);
not NOT1 (N13089, N13044);
or OR2 (N13090, N13083, N6128);
not NOT1 (N13091, N13088);
or OR2 (N13092, N13090, N4431);
xor XOR2 (N13093, N13091, N12257);
nand NAND3 (N13094, N13078, N4399, N10149);
nand NAND3 (N13095, N13075, N2642, N10983);
xor XOR2 (N13096, N13089, N2086);
xor XOR2 (N13097, N13079, N11171);
and AND4 (N13098, N13097, N11939, N6510, N8666);
buf BUF1 (N13099, N13096);
buf BUF1 (N13100, N13087);
not NOT1 (N13101, N13084);
nor NOR2 (N13102, N13095, N4106);
not NOT1 (N13103, N13081);
buf BUF1 (N13104, N13085);
nor NOR3 (N13105, N13094, N3045, N4838);
or OR4 (N13106, N13099, N1506, N8658, N10932);
xor XOR2 (N13107, N13092, N4007);
or OR3 (N13108, N13106, N5617, N280);
nor NOR3 (N13109, N13108, N8388, N2659);
xor XOR2 (N13110, N13101, N11393);
nand NAND2 (N13111, N13109, N4899);
nand NAND4 (N13112, N13110, N10925, N9040, N4651);
not NOT1 (N13113, N13102);
buf BUF1 (N13114, N13105);
nand NAND2 (N13115, N13113, N5778);
or OR3 (N13116, N13107, N2456, N4113);
and AND4 (N13117, N13115, N5980, N8376, N6329);
and AND4 (N13118, N13100, N9041, N2150, N40);
xor XOR2 (N13119, N13114, N3838);
xor XOR2 (N13120, N13112, N2314);
nor NOR3 (N13121, N13116, N7673, N2535);
and AND4 (N13122, N13118, N2435, N5117, N6430);
not NOT1 (N13123, N13122);
or OR2 (N13124, N13123, N10424);
or OR4 (N13125, N13111, N1061, N11509, N4114);
buf BUF1 (N13126, N13098);
nand NAND4 (N13127, N13119, N10878, N8289, N1387);
and AND3 (N13128, N13117, N188, N6271);
nand NAND2 (N13129, N13121, N1279);
nor NOR3 (N13130, N13120, N6886, N11717);
nor NOR2 (N13131, N13127, N2010);
not NOT1 (N13132, N13130);
not NOT1 (N13133, N13104);
and AND3 (N13134, N13133, N7952, N1073);
xor XOR2 (N13135, N13093, N12864);
or OR2 (N13136, N13128, N7291);
and AND3 (N13137, N13125, N1118, N6267);
nor NOR3 (N13138, N13103, N4720, N5851);
nand NAND4 (N13139, N13129, N2000, N6302, N5982);
and AND3 (N13140, N13124, N694, N4154);
buf BUF1 (N13141, N13131);
nand NAND2 (N13142, N13138, N11689);
not NOT1 (N13143, N13141);
or OR2 (N13144, N13142, N6609);
buf BUF1 (N13145, N13139);
xor XOR2 (N13146, N13126, N11209);
or OR4 (N13147, N13146, N7079, N13082, N2894);
not NOT1 (N13148, N13145);
not NOT1 (N13149, N13144);
nand NAND4 (N13150, N13137, N1056, N4985, N9825);
buf BUF1 (N13151, N13148);
buf BUF1 (N13152, N13150);
nor NOR2 (N13153, N13152, N13047);
and AND3 (N13154, N13135, N12634, N12020);
not NOT1 (N13155, N13140);
nand NAND2 (N13156, N13134, N9512);
and AND4 (N13157, N13154, N3554, N12814, N3400);
or OR3 (N13158, N13136, N3650, N6874);
buf BUF1 (N13159, N13151);
or OR3 (N13160, N13159, N12098, N2206);
buf BUF1 (N13161, N13147);
and AND3 (N13162, N13161, N3313, N998);
or OR3 (N13163, N13132, N657, N2562);
and AND4 (N13164, N13160, N1698, N1585, N1214);
and AND3 (N13165, N13149, N10996, N4538);
buf BUF1 (N13166, N13156);
or OR2 (N13167, N13143, N418);
and AND3 (N13168, N13165, N12847, N2233);
or OR2 (N13169, N13158, N3097);
not NOT1 (N13170, N13169);
or OR3 (N13171, N13162, N7473, N1857);
buf BUF1 (N13172, N13164);
not NOT1 (N13173, N13166);
or OR3 (N13174, N13155, N3678, N7327);
and AND2 (N13175, N13163, N4348);
nor NOR3 (N13176, N13171, N5428, N6873);
nor NOR2 (N13177, N13168, N10803);
buf BUF1 (N13178, N13176);
not NOT1 (N13179, N13177);
xor XOR2 (N13180, N13174, N12133);
and AND3 (N13181, N13157, N8302, N12453);
nand NAND3 (N13182, N13179, N2812, N8036);
xor XOR2 (N13183, N13172, N4420);
nand NAND3 (N13184, N13153, N8439, N12330);
nand NAND4 (N13185, N13181, N6594, N3128, N11070);
xor XOR2 (N13186, N13170, N10114);
buf BUF1 (N13187, N13178);
not NOT1 (N13188, N13180);
and AND2 (N13189, N13167, N4597);
xor XOR2 (N13190, N13183, N655);
xor XOR2 (N13191, N13184, N11784);
not NOT1 (N13192, N13189);
and AND2 (N13193, N13187, N5091);
buf BUF1 (N13194, N13173);
nor NOR3 (N13195, N13185, N9290, N5074);
xor XOR2 (N13196, N13195, N7205);
xor XOR2 (N13197, N13194, N4967);
nand NAND2 (N13198, N13193, N11635);
buf BUF1 (N13199, N13197);
nor NOR2 (N13200, N13198, N91);
or OR4 (N13201, N13186, N9071, N7280, N2368);
nand NAND3 (N13202, N13191, N790, N2831);
xor XOR2 (N13203, N13192, N11529);
not NOT1 (N13204, N13203);
and AND3 (N13205, N13204, N5812, N2500);
and AND3 (N13206, N13175, N1866, N13162);
xor XOR2 (N13207, N13200, N2529);
or OR2 (N13208, N13201, N3489);
xor XOR2 (N13209, N13199, N6252);
or OR2 (N13210, N13205, N380);
not NOT1 (N13211, N13210);
buf BUF1 (N13212, N13188);
xor XOR2 (N13213, N13190, N3687);
or OR2 (N13214, N13196, N4371);
not NOT1 (N13215, N13214);
and AND4 (N13216, N13211, N7822, N7859, N7426);
not NOT1 (N13217, N13202);
and AND2 (N13218, N13208, N2605);
xor XOR2 (N13219, N13207, N1661);
nand NAND3 (N13220, N13216, N9665, N924);
buf BUF1 (N13221, N13220);
not NOT1 (N13222, N13218);
nor NOR2 (N13223, N13217, N3564);
nor NOR4 (N13224, N13213, N11110, N526, N12935);
nand NAND3 (N13225, N13206, N2773, N5894);
and AND2 (N13226, N13219, N7157);
buf BUF1 (N13227, N13222);
or OR3 (N13228, N13226, N12583, N8038);
not NOT1 (N13229, N13224);
or OR4 (N13230, N13209, N6908, N2518, N4770);
buf BUF1 (N13231, N13215);
nand NAND3 (N13232, N13212, N5436, N3525);
nor NOR3 (N13233, N13229, N10633, N109);
nor NOR2 (N13234, N13225, N3976);
not NOT1 (N13235, N13230);
nor NOR2 (N13236, N13182, N11986);
nand NAND3 (N13237, N13233, N12119, N9297);
not NOT1 (N13238, N13223);
xor XOR2 (N13239, N13221, N1173);
and AND2 (N13240, N13235, N3089);
and AND3 (N13241, N13237, N11170, N1069);
buf BUF1 (N13242, N13234);
nor NOR3 (N13243, N13232, N6286, N1703);
xor XOR2 (N13244, N13231, N12946);
nor NOR2 (N13245, N13239, N13036);
and AND2 (N13246, N13227, N7292);
buf BUF1 (N13247, N13228);
buf BUF1 (N13248, N13245);
not NOT1 (N13249, N13244);
nand NAND4 (N13250, N13249, N6235, N843, N427);
or OR4 (N13251, N13248, N1835, N7811, N12009);
and AND2 (N13252, N13243, N5182);
or OR2 (N13253, N13251, N8933);
and AND3 (N13254, N13236, N9644, N1836);
and AND2 (N13255, N13254, N9571);
xor XOR2 (N13256, N13255, N9552);
nand NAND3 (N13257, N13246, N7174, N5683);
or OR4 (N13258, N13250, N2562, N967, N135);
nor NOR2 (N13259, N13258, N9376);
or OR3 (N13260, N13253, N564, N8427);
nand NAND3 (N13261, N13240, N4077, N4161);
not NOT1 (N13262, N13261);
or OR4 (N13263, N13262, N7879, N453, N3673);
not NOT1 (N13264, N13259);
nor NOR3 (N13265, N13263, N10809, N12678);
nor NOR3 (N13266, N13264, N11671, N9436);
nand NAND2 (N13267, N13257, N9949);
buf BUF1 (N13268, N13266);
not NOT1 (N13269, N13260);
and AND3 (N13270, N13265, N1053, N6945);
or OR3 (N13271, N13238, N2142, N13187);
or OR2 (N13272, N13268, N11103);
and AND2 (N13273, N13247, N7638);
not NOT1 (N13274, N13270);
nor NOR4 (N13275, N13269, N206, N7932, N13081);
and AND3 (N13276, N13274, N13138, N5819);
xor XOR2 (N13277, N13256, N6622);
and AND3 (N13278, N13271, N6158, N12574);
xor XOR2 (N13279, N13252, N8544);
buf BUF1 (N13280, N13241);
nor NOR4 (N13281, N13280, N5332, N6418, N3534);
xor XOR2 (N13282, N13242, N2147);
buf BUF1 (N13283, N13276);
nand NAND2 (N13284, N13277, N4201);
nand NAND4 (N13285, N13275, N929, N4428, N12036);
xor XOR2 (N13286, N13267, N3483);
and AND4 (N13287, N13279, N11402, N3557, N12795);
or OR3 (N13288, N13281, N7020, N13256);
buf BUF1 (N13289, N13288);
not NOT1 (N13290, N13272);
not NOT1 (N13291, N13284);
nand NAND2 (N13292, N13290, N3018);
xor XOR2 (N13293, N13285, N5874);
buf BUF1 (N13294, N13292);
nor NOR2 (N13295, N13293, N13148);
and AND4 (N13296, N13291, N10439, N7719, N12571);
nor NOR4 (N13297, N13287, N2546, N4298, N12246);
and AND3 (N13298, N13295, N4800, N13086);
or OR4 (N13299, N13297, N12919, N2815, N4769);
nand NAND4 (N13300, N13286, N6996, N2487, N1882);
not NOT1 (N13301, N13283);
xor XOR2 (N13302, N13296, N10708);
or OR3 (N13303, N13282, N8201, N6577);
buf BUF1 (N13304, N13302);
not NOT1 (N13305, N13299);
buf BUF1 (N13306, N13305);
nand NAND3 (N13307, N13273, N4741, N1589);
not NOT1 (N13308, N13306);
not NOT1 (N13309, N13301);
xor XOR2 (N13310, N13278, N2547);
nor NOR4 (N13311, N13289, N1661, N2341, N9279);
not NOT1 (N13312, N13304);
nand NAND2 (N13313, N13294, N3728);
buf BUF1 (N13314, N13303);
buf BUF1 (N13315, N13314);
xor XOR2 (N13316, N13313, N11665);
nand NAND3 (N13317, N13312, N10848, N4709);
and AND3 (N13318, N13311, N10112, N4043);
and AND4 (N13319, N13298, N13072, N7832, N7922);
and AND2 (N13320, N13319, N5191);
or OR4 (N13321, N13315, N7104, N3802, N8770);
buf BUF1 (N13322, N13309);
and AND3 (N13323, N13320, N9141, N1340);
or OR4 (N13324, N13310, N4773, N12588, N782);
xor XOR2 (N13325, N13324, N4174);
not NOT1 (N13326, N13322);
or OR2 (N13327, N13321, N11537);
nor NOR4 (N13328, N13318, N4418, N178, N354);
nand NAND4 (N13329, N13308, N1514, N2449, N10236);
and AND2 (N13330, N13323, N3918);
nand NAND2 (N13331, N13330, N40);
buf BUF1 (N13332, N13300);
buf BUF1 (N13333, N13328);
not NOT1 (N13334, N13331);
buf BUF1 (N13335, N13333);
xor XOR2 (N13336, N13332, N1725);
buf BUF1 (N13337, N13327);
not NOT1 (N13338, N13326);
nand NAND4 (N13339, N13335, N9144, N3321, N1492);
buf BUF1 (N13340, N13329);
or OR2 (N13341, N13337, N3136);
and AND4 (N13342, N13316, N1603, N4839, N1987);
nand NAND2 (N13343, N13342, N638);
nor NOR3 (N13344, N13339, N7567, N1716);
nor NOR2 (N13345, N13341, N1243);
buf BUF1 (N13346, N13334);
xor XOR2 (N13347, N13340, N3282);
and AND2 (N13348, N13307, N13177);
and AND2 (N13349, N13343, N2936);
buf BUF1 (N13350, N13338);
buf BUF1 (N13351, N13350);
not NOT1 (N13352, N13345);
or OR2 (N13353, N13351, N2842);
or OR2 (N13354, N13336, N9085);
nor NOR2 (N13355, N13354, N2055);
not NOT1 (N13356, N13352);
nor NOR3 (N13357, N13353, N12835, N10323);
not NOT1 (N13358, N13325);
xor XOR2 (N13359, N13317, N2960);
or OR2 (N13360, N13347, N9745);
nor NOR4 (N13361, N13344, N3216, N7134, N9441);
not NOT1 (N13362, N13355);
buf BUF1 (N13363, N13349);
or OR3 (N13364, N13363, N5732, N8172);
xor XOR2 (N13365, N13348, N12675);
and AND4 (N13366, N13356, N9262, N3931, N2714);
nand NAND4 (N13367, N13361, N7617, N6853, N12762);
xor XOR2 (N13368, N13365, N13254);
not NOT1 (N13369, N13358);
and AND3 (N13370, N13346, N12914, N8843);
nor NOR4 (N13371, N13366, N12702, N1656, N12142);
xor XOR2 (N13372, N13357, N8984);
xor XOR2 (N13373, N13368, N7191);
xor XOR2 (N13374, N13373, N3940);
or OR4 (N13375, N13360, N2595, N2206, N932);
nand NAND2 (N13376, N13367, N2286);
buf BUF1 (N13377, N13364);
nor NOR4 (N13378, N13359, N9263, N9724, N11704);
nand NAND3 (N13379, N13370, N6408, N8725);
nand NAND4 (N13380, N13375, N13228, N9828, N2892);
xor XOR2 (N13381, N13379, N1023);
not NOT1 (N13382, N13377);
not NOT1 (N13383, N13380);
nor NOR3 (N13384, N13374, N8975, N4920);
nor NOR2 (N13385, N13378, N2504);
and AND4 (N13386, N13383, N7646, N2806, N7641);
nor NOR4 (N13387, N13369, N7575, N11009, N12194);
and AND2 (N13388, N13381, N5557);
nand NAND2 (N13389, N13372, N4842);
nor NOR2 (N13390, N13386, N10722);
buf BUF1 (N13391, N13387);
nor NOR2 (N13392, N13376, N5365);
and AND3 (N13393, N13385, N11110, N6465);
or OR4 (N13394, N13388, N2249, N11048, N681);
nor NOR4 (N13395, N13382, N4864, N8731, N4701);
xor XOR2 (N13396, N13384, N12277);
and AND4 (N13397, N13392, N6817, N1541, N1434);
not NOT1 (N13398, N13390);
or OR4 (N13399, N13391, N7771, N4057, N12437);
xor XOR2 (N13400, N13389, N8149);
not NOT1 (N13401, N13396);
not NOT1 (N13402, N13400);
not NOT1 (N13403, N13398);
xor XOR2 (N13404, N13393, N4475);
nor NOR3 (N13405, N13404, N10906, N7809);
and AND4 (N13406, N13397, N11634, N12661, N4581);
nor NOR4 (N13407, N13403, N13243, N4574, N12038);
buf BUF1 (N13408, N13406);
and AND4 (N13409, N13401, N11464, N7962, N3125);
nand NAND2 (N13410, N13395, N7370);
not NOT1 (N13411, N13402);
not NOT1 (N13412, N13405);
and AND2 (N13413, N13371, N911);
nor NOR4 (N13414, N13411, N996, N779, N11609);
buf BUF1 (N13415, N13399);
not NOT1 (N13416, N13415);
or OR2 (N13417, N13408, N544);
not NOT1 (N13418, N13417);
nor NOR4 (N13419, N13409, N8505, N5645, N2784);
xor XOR2 (N13420, N13394, N1121);
buf BUF1 (N13421, N13407);
or OR4 (N13422, N13420, N899, N9729, N8752);
xor XOR2 (N13423, N13416, N9431);
not NOT1 (N13424, N13419);
nand NAND4 (N13425, N13412, N4876, N2044, N7857);
and AND4 (N13426, N13423, N6196, N8868, N7630);
buf BUF1 (N13427, N13425);
nor NOR3 (N13428, N13414, N2724, N6121);
not NOT1 (N13429, N13426);
nor NOR3 (N13430, N13428, N758, N586);
nand NAND4 (N13431, N13422, N5371, N1359, N12872);
xor XOR2 (N13432, N13429, N12534);
and AND4 (N13433, N13421, N10596, N3129, N9073);
or OR3 (N13434, N13413, N7028, N3631);
and AND3 (N13435, N13430, N9229, N8394);
buf BUF1 (N13436, N13410);
xor XOR2 (N13437, N13418, N8562);
buf BUF1 (N13438, N13432);
nor NOR2 (N13439, N13424, N12319);
xor XOR2 (N13440, N13436, N6432);
or OR3 (N13441, N13433, N12704, N3994);
xor XOR2 (N13442, N13362, N311);
or OR4 (N13443, N13431, N5216, N12666, N9608);
or OR4 (N13444, N13437, N11096, N6463, N6577);
nor NOR4 (N13445, N13439, N1588, N9068, N357);
and AND3 (N13446, N13445, N3474, N5569);
and AND3 (N13447, N13444, N9930, N614);
nand NAND4 (N13448, N13434, N2978, N8773, N6752);
and AND4 (N13449, N13441, N2812, N12659, N3067);
and AND2 (N13450, N13435, N2002);
xor XOR2 (N13451, N13447, N8671);
not NOT1 (N13452, N13450);
buf BUF1 (N13453, N13449);
or OR4 (N13454, N13446, N12896, N13406, N12587);
nand NAND3 (N13455, N13453, N10039, N13374);
nand NAND3 (N13456, N13448, N1326, N10289);
nand NAND2 (N13457, N13455, N555);
buf BUF1 (N13458, N13456);
nand NAND2 (N13459, N13438, N9702);
not NOT1 (N13460, N13440);
buf BUF1 (N13461, N13457);
not NOT1 (N13462, N13460);
nand NAND3 (N13463, N13459, N2399, N464);
xor XOR2 (N13464, N13451, N12543);
nor NOR3 (N13465, N13463, N10139, N3504);
or OR2 (N13466, N13462, N13131);
or OR3 (N13467, N13466, N10733, N7203);
buf BUF1 (N13468, N13454);
nand NAND2 (N13469, N13467, N4887);
buf BUF1 (N13470, N13461);
and AND4 (N13471, N13427, N12324, N2271, N8963);
xor XOR2 (N13472, N13470, N5071);
or OR2 (N13473, N13468, N12253);
nor NOR3 (N13474, N13473, N12572, N3542);
nor NOR4 (N13475, N13443, N2553, N1122, N9755);
nor NOR4 (N13476, N13465, N5689, N11845, N423);
not NOT1 (N13477, N13452);
and AND2 (N13478, N13458, N1642);
or OR3 (N13479, N13471, N7025, N4637);
xor XOR2 (N13480, N13475, N4514);
xor XOR2 (N13481, N13476, N7838);
not NOT1 (N13482, N13469);
nor NOR4 (N13483, N13481, N9836, N4397, N3683);
nor NOR4 (N13484, N13477, N11123, N1526, N13222);
buf BUF1 (N13485, N13483);
buf BUF1 (N13486, N13484);
nor NOR3 (N13487, N13482, N5582, N12825);
nand NAND3 (N13488, N13485, N12921, N5919);
xor XOR2 (N13489, N13442, N8852);
and AND3 (N13490, N13486, N8332, N10881);
buf BUF1 (N13491, N13464);
nand NAND4 (N13492, N13487, N9603, N6320, N9715);
xor XOR2 (N13493, N13492, N649);
nand NAND4 (N13494, N13491, N6418, N9616, N5719);
nor NOR3 (N13495, N13494, N9417, N10513);
xor XOR2 (N13496, N13495, N12405);
nand NAND2 (N13497, N13496, N12784);
and AND4 (N13498, N13488, N8855, N1437, N11666);
xor XOR2 (N13499, N13493, N5590);
nor NOR3 (N13500, N13480, N6099, N2630);
buf BUF1 (N13501, N13500);
or OR3 (N13502, N13489, N3400, N10895);
nor NOR3 (N13503, N13498, N201, N8972);
nand NAND3 (N13504, N13503, N2162, N5191);
xor XOR2 (N13505, N13490, N7613);
or OR3 (N13506, N13479, N1166, N2649);
nand NAND2 (N13507, N13497, N6949);
xor XOR2 (N13508, N13507, N588);
buf BUF1 (N13509, N13505);
or OR2 (N13510, N13472, N5010);
xor XOR2 (N13511, N13506, N7237);
nand NAND3 (N13512, N13478, N7588, N6837);
nand NAND3 (N13513, N13511, N8737, N1470);
not NOT1 (N13514, N13512);
nor NOR2 (N13515, N13509, N11707);
nand NAND4 (N13516, N13474, N3314, N792, N10641);
and AND2 (N13517, N13499, N3483);
nand NAND2 (N13518, N13514, N1297);
not NOT1 (N13519, N13502);
nand NAND3 (N13520, N13515, N205, N142);
and AND2 (N13521, N13520, N3692);
or OR4 (N13522, N13519, N12572, N5078, N10871);
nand NAND4 (N13523, N13508, N11575, N5051, N11309);
or OR4 (N13524, N13516, N9614, N784, N10579);
or OR4 (N13525, N13524, N958, N12406, N909);
not NOT1 (N13526, N13523);
or OR2 (N13527, N13517, N6213);
buf BUF1 (N13528, N13501);
buf BUF1 (N13529, N13527);
xor XOR2 (N13530, N13525, N640);
nor NOR2 (N13531, N13504, N10769);
not NOT1 (N13532, N13518);
nor NOR3 (N13533, N13513, N1141, N4440);
and AND2 (N13534, N13522, N2537);
and AND3 (N13535, N13526, N1621, N7996);
buf BUF1 (N13536, N13530);
xor XOR2 (N13537, N13521, N2194);
or OR3 (N13538, N13532, N6682, N2972);
or OR4 (N13539, N13531, N11577, N11973, N6180);
and AND3 (N13540, N13529, N4008, N9277);
buf BUF1 (N13541, N13534);
buf BUF1 (N13542, N13540);
xor XOR2 (N13543, N13533, N2084);
or OR3 (N13544, N13510, N13091, N4835);
nand NAND2 (N13545, N13536, N954);
or OR2 (N13546, N13545, N7647);
xor XOR2 (N13547, N13538, N10693);
and AND2 (N13548, N13537, N12691);
buf BUF1 (N13549, N13535);
or OR2 (N13550, N13546, N1981);
and AND3 (N13551, N13548, N2003, N8636);
not NOT1 (N13552, N13544);
or OR4 (N13553, N13539, N3825, N12101, N3560);
and AND2 (N13554, N13528, N10371);
nor NOR4 (N13555, N13551, N6635, N3574, N1499);
and AND4 (N13556, N13555, N10749, N11986, N9171);
nor NOR4 (N13557, N13547, N2051, N10107, N4101);
xor XOR2 (N13558, N13553, N1217);
or OR2 (N13559, N13556, N1995);
not NOT1 (N13560, N13550);
buf BUF1 (N13561, N13557);
buf BUF1 (N13562, N13552);
buf BUF1 (N13563, N13541);
xor XOR2 (N13564, N13558, N12937);
nand NAND4 (N13565, N13560, N7693, N3742, N3055);
buf BUF1 (N13566, N13565);
nor NOR3 (N13567, N13563, N5958, N9442);
or OR2 (N13568, N13549, N11043);
nor NOR2 (N13569, N13561, N7993);
or OR2 (N13570, N13566, N12312);
not NOT1 (N13571, N13543);
nor NOR3 (N13572, N13571, N6134, N13340);
nand NAND4 (N13573, N13569, N9220, N4197, N8507);
or OR2 (N13574, N13564, N2239);
nand NAND3 (N13575, N13554, N132, N7509);
and AND4 (N13576, N13559, N4074, N9994, N3210);
buf BUF1 (N13577, N13567);
not NOT1 (N13578, N13542);
buf BUF1 (N13579, N13574);
or OR4 (N13580, N13572, N10258, N12175, N4333);
xor XOR2 (N13581, N13579, N1460);
not NOT1 (N13582, N13578);
xor XOR2 (N13583, N13575, N12017);
not NOT1 (N13584, N13577);
not NOT1 (N13585, N13573);
nand NAND4 (N13586, N13584, N8529, N2030, N6226);
and AND4 (N13587, N13581, N6636, N1212, N586);
not NOT1 (N13588, N13568);
nor NOR4 (N13589, N13583, N10283, N5779, N10371);
nor NOR3 (N13590, N13570, N7171, N3312);
and AND3 (N13591, N13586, N10058, N6425);
nand NAND4 (N13592, N13587, N5156, N8082, N5023);
xor XOR2 (N13593, N13576, N11240);
xor XOR2 (N13594, N13585, N3557);
nor NOR4 (N13595, N13594, N12777, N12815, N2635);
not NOT1 (N13596, N13588);
not NOT1 (N13597, N13592);
nand NAND4 (N13598, N13596, N10155, N8373, N11096);
xor XOR2 (N13599, N13580, N4526);
not NOT1 (N13600, N13598);
xor XOR2 (N13601, N13582, N10718);
xor XOR2 (N13602, N13600, N12447);
buf BUF1 (N13603, N13593);
nor NOR3 (N13604, N13595, N13159, N6440);
nand NAND3 (N13605, N13603, N7303, N2869);
not NOT1 (N13606, N13562);
not NOT1 (N13607, N13604);
xor XOR2 (N13608, N13591, N6872);
nor NOR4 (N13609, N13608, N12588, N11999, N197);
and AND4 (N13610, N13601, N5824, N7477, N1395);
xor XOR2 (N13611, N13606, N11368);
and AND2 (N13612, N13599, N7790);
and AND3 (N13613, N13589, N7190, N13339);
and AND3 (N13614, N13613, N12129, N8263);
nand NAND2 (N13615, N13612, N2708);
and AND4 (N13616, N13602, N408, N3851, N4075);
or OR3 (N13617, N13615, N1798, N2508);
and AND3 (N13618, N13607, N7022, N11467);
nand NAND4 (N13619, N13616, N9645, N6204, N5266);
nor NOR3 (N13620, N13617, N5647, N791);
nand NAND2 (N13621, N13610, N9180);
and AND4 (N13622, N13609, N2853, N12435, N11815);
not NOT1 (N13623, N13597);
buf BUF1 (N13624, N13622);
or OR3 (N13625, N13623, N4635, N12332);
xor XOR2 (N13626, N13605, N2361);
xor XOR2 (N13627, N13626, N10059);
and AND4 (N13628, N13627, N10045, N3891, N9363);
buf BUF1 (N13629, N13618);
or OR4 (N13630, N13624, N12391, N11994, N7217);
not NOT1 (N13631, N13614);
xor XOR2 (N13632, N13621, N9603);
and AND4 (N13633, N13629, N5377, N5306, N13163);
or OR3 (N13634, N13625, N6334, N12484);
nand NAND2 (N13635, N13620, N902);
xor XOR2 (N13636, N13611, N11034);
buf BUF1 (N13637, N13633);
nand NAND3 (N13638, N13636, N9351, N629);
nor NOR4 (N13639, N13632, N10326, N9836, N353);
and AND2 (N13640, N13630, N788);
xor XOR2 (N13641, N13590, N9646);
nor NOR3 (N13642, N13641, N12658, N7378);
or OR4 (N13643, N13634, N2946, N2952, N7649);
or OR3 (N13644, N13635, N11298, N3580);
or OR2 (N13645, N13619, N11414);
nand NAND3 (N13646, N13645, N12974, N11058);
not NOT1 (N13647, N13639);
buf BUF1 (N13648, N13647);
or OR4 (N13649, N13638, N216, N5472, N8033);
xor XOR2 (N13650, N13628, N12486);
and AND2 (N13651, N13637, N10064);
nand NAND3 (N13652, N13646, N5518, N1936);
xor XOR2 (N13653, N13652, N10671);
or OR3 (N13654, N13650, N6676, N655);
buf BUF1 (N13655, N13642);
and AND4 (N13656, N13651, N11968, N7264, N4144);
xor XOR2 (N13657, N13648, N1551);
not NOT1 (N13658, N13643);
nand NAND3 (N13659, N13631, N9778, N4557);
not NOT1 (N13660, N13649);
and AND4 (N13661, N13656, N3024, N8156, N10223);
not NOT1 (N13662, N13659);
buf BUF1 (N13663, N13654);
buf BUF1 (N13664, N13640);
nand NAND4 (N13665, N13653, N3395, N5779, N9421);
xor XOR2 (N13666, N13665, N4470);
nand NAND3 (N13667, N13663, N11123, N9996);
and AND2 (N13668, N13661, N2877);
not NOT1 (N13669, N13655);
not NOT1 (N13670, N13662);
xor XOR2 (N13671, N13670, N8221);
buf BUF1 (N13672, N13668);
xor XOR2 (N13673, N13664, N3820);
nand NAND2 (N13674, N13658, N7657);
nand NAND2 (N13675, N13673, N11262);
buf BUF1 (N13676, N13657);
or OR4 (N13677, N13672, N2592, N6049, N2591);
not NOT1 (N13678, N13677);
buf BUF1 (N13679, N13667);
nand NAND2 (N13680, N13660, N5866);
buf BUF1 (N13681, N13675);
buf BUF1 (N13682, N13644);
nor NOR2 (N13683, N13682, N11169);
nor NOR3 (N13684, N13669, N8915, N5031);
and AND2 (N13685, N13666, N12995);
xor XOR2 (N13686, N13680, N3702);
and AND4 (N13687, N13678, N8049, N11315, N446);
and AND4 (N13688, N13684, N7721, N13261, N5493);
or OR2 (N13689, N13679, N6538);
and AND3 (N13690, N13671, N5012, N12743);
xor XOR2 (N13691, N13685, N4127);
not NOT1 (N13692, N13686);
nor NOR4 (N13693, N13674, N5292, N7392, N12725);
nor NOR4 (N13694, N13692, N12393, N2386, N10824);
xor XOR2 (N13695, N13689, N8604);
nor NOR4 (N13696, N13695, N8153, N4856, N5283);
nor NOR2 (N13697, N13687, N10894);
nand NAND2 (N13698, N13681, N7226);
and AND3 (N13699, N13690, N4751, N1954);
or OR4 (N13700, N13697, N736, N9016, N3643);
nor NOR4 (N13701, N13676, N5709, N811, N8586);
or OR3 (N13702, N13700, N13313, N451);
nand NAND3 (N13703, N13693, N10294, N5326);
not NOT1 (N13704, N13701);
buf BUF1 (N13705, N13704);
nor NOR2 (N13706, N13683, N11720);
not NOT1 (N13707, N13698);
and AND4 (N13708, N13688, N7906, N8708, N2286);
and AND4 (N13709, N13705, N2754, N2510, N788);
xor XOR2 (N13710, N13699, N10431);
and AND3 (N13711, N13706, N1508, N3523);
not NOT1 (N13712, N13710);
nor NOR2 (N13713, N13709, N7648);
buf BUF1 (N13714, N13708);
and AND3 (N13715, N13713, N9714, N606);
and AND4 (N13716, N13696, N11764, N9923, N7938);
not NOT1 (N13717, N13711);
nor NOR4 (N13718, N13707, N9736, N1422, N8984);
nor NOR2 (N13719, N13703, N7972);
and AND2 (N13720, N13714, N11287);
xor XOR2 (N13721, N13720, N2113);
or OR4 (N13722, N13716, N4172, N12213, N5514);
nand NAND2 (N13723, N13702, N6060);
nand NAND4 (N13724, N13694, N2678, N806, N5691);
and AND4 (N13725, N13721, N11897, N7164, N7141);
nand NAND2 (N13726, N13718, N13715);
xor XOR2 (N13727, N9398, N7685);
nand NAND3 (N13728, N13722, N5070, N3280);
not NOT1 (N13729, N13724);
and AND3 (N13730, N13728, N8089, N4042);
nand NAND3 (N13731, N13691, N2661, N13259);
nor NOR2 (N13732, N13712, N1761);
or OR2 (N13733, N13732, N944);
or OR3 (N13734, N13725, N7420, N2554);
buf BUF1 (N13735, N13730);
buf BUF1 (N13736, N13734);
or OR4 (N13737, N13733, N7837, N6096, N3006);
xor XOR2 (N13738, N13726, N13722);
buf BUF1 (N13739, N13727);
nand NAND4 (N13740, N13737, N1385, N1815, N7014);
xor XOR2 (N13741, N13736, N1778);
and AND3 (N13742, N13738, N9362, N12147);
nand NAND3 (N13743, N13731, N86, N1216);
xor XOR2 (N13744, N13741, N10722);
and AND4 (N13745, N13740, N5244, N2239, N4835);
not NOT1 (N13746, N13742);
nor NOR2 (N13747, N13746, N1635);
and AND2 (N13748, N13717, N12014);
nor NOR4 (N13749, N13729, N4212, N849, N4147);
xor XOR2 (N13750, N13743, N2485);
or OR4 (N13751, N13749, N2160, N4499, N1699);
or OR4 (N13752, N13739, N3783, N10143, N5391);
xor XOR2 (N13753, N13747, N2192);
nor NOR2 (N13754, N13751, N2094);
xor XOR2 (N13755, N13753, N11381);
and AND3 (N13756, N13754, N10866, N5083);
or OR3 (N13757, N13719, N6643, N8642);
nor NOR2 (N13758, N13744, N804);
buf BUF1 (N13759, N13752);
buf BUF1 (N13760, N13758);
not NOT1 (N13761, N13756);
buf BUF1 (N13762, N13760);
nand NAND4 (N13763, N13757, N7399, N6892, N5099);
not NOT1 (N13764, N13750);
buf BUF1 (N13765, N13748);
and AND2 (N13766, N13723, N7130);
not NOT1 (N13767, N13745);
not NOT1 (N13768, N13766);
not NOT1 (N13769, N13735);
nor NOR2 (N13770, N13767, N9621);
and AND2 (N13771, N13761, N7430);
or OR4 (N13772, N13759, N6506, N1586, N5052);
or OR4 (N13773, N13764, N1928, N1408, N5889);
or OR4 (N13774, N13762, N4218, N10070, N7927);
xor XOR2 (N13775, N13772, N1597);
nor NOR4 (N13776, N13768, N4223, N9517, N6799);
not NOT1 (N13777, N13769);
nand NAND2 (N13778, N13774, N11873);
nor NOR4 (N13779, N13773, N10874, N7200, N6768);
and AND3 (N13780, N13779, N9507, N7399);
xor XOR2 (N13781, N13771, N12033);
nor NOR3 (N13782, N13780, N7045, N1427);
nand NAND4 (N13783, N13763, N6701, N3057, N762);
xor XOR2 (N13784, N13765, N7470);
or OR4 (N13785, N13777, N8685, N11494, N10314);
or OR3 (N13786, N13785, N13454, N13417);
or OR4 (N13787, N13778, N9404, N629, N12242);
and AND3 (N13788, N13787, N2310, N12316);
nand NAND2 (N13789, N13770, N651);
xor XOR2 (N13790, N13784, N6445);
nand NAND4 (N13791, N13789, N13506, N3052, N13334);
nand NAND4 (N13792, N13775, N5461, N7433, N1658);
nand NAND2 (N13793, N13776, N9532);
not NOT1 (N13794, N13788);
or OR2 (N13795, N13791, N8882);
and AND3 (N13796, N13793, N3259, N9151);
nor NOR3 (N13797, N13792, N8749, N544);
buf BUF1 (N13798, N13783);
and AND3 (N13799, N13795, N2432, N12779);
or OR3 (N13800, N13755, N6755, N5883);
nor NOR2 (N13801, N13799, N7341);
buf BUF1 (N13802, N13801);
nand NAND4 (N13803, N13781, N2613, N1055, N5713);
and AND3 (N13804, N13798, N4304, N3644);
nor NOR4 (N13805, N13802, N3622, N7057, N12903);
and AND2 (N13806, N13794, N6045);
and AND3 (N13807, N13782, N9395, N6889);
nand NAND4 (N13808, N13786, N7475, N10778, N10883);
xor XOR2 (N13809, N13808, N5984);
xor XOR2 (N13810, N13797, N10984);
xor XOR2 (N13811, N13809, N1147);
nand NAND2 (N13812, N13804, N3425);
buf BUF1 (N13813, N13806);
not NOT1 (N13814, N13811);
nor NOR3 (N13815, N13796, N7373, N6056);
nor NOR3 (N13816, N13805, N10792, N12578);
and AND4 (N13817, N13800, N597, N11458, N1114);
not NOT1 (N13818, N13790);
or OR4 (N13819, N13817, N2368, N7735, N2044);
and AND4 (N13820, N13810, N7529, N13666, N11876);
nand NAND3 (N13821, N13814, N7404, N939);
nor NOR3 (N13822, N13819, N5111, N5914);
not NOT1 (N13823, N13821);
buf BUF1 (N13824, N13807);
nand NAND3 (N13825, N13803, N3336, N1074);
nor NOR3 (N13826, N13815, N4467, N13657);
nand NAND2 (N13827, N13820, N1715);
and AND3 (N13828, N13822, N3193, N442);
not NOT1 (N13829, N13826);
or OR2 (N13830, N13818, N3926);
and AND2 (N13831, N13812, N7351);
nand NAND3 (N13832, N13828, N13617, N4245);
buf BUF1 (N13833, N13816);
xor XOR2 (N13834, N13830, N4155);
nand NAND2 (N13835, N13824, N5389);
nor NOR4 (N13836, N13834, N8952, N846, N13796);
and AND3 (N13837, N13831, N1268, N1925);
xor XOR2 (N13838, N13835, N8855);
nor NOR2 (N13839, N13813, N2551);
nor NOR4 (N13840, N13823, N8390, N1189, N12482);
xor XOR2 (N13841, N13837, N12901);
not NOT1 (N13842, N13839);
nand NAND4 (N13843, N13840, N5701, N6791, N10663);
nor NOR3 (N13844, N13833, N6932, N10279);
nand NAND2 (N13845, N13829, N13532);
xor XOR2 (N13846, N13825, N9833);
or OR3 (N13847, N13838, N4276, N5705);
and AND4 (N13848, N13847, N5128, N3833, N10956);
or OR2 (N13849, N13827, N9137);
not NOT1 (N13850, N13832);
not NOT1 (N13851, N13850);
not NOT1 (N13852, N13845);
nand NAND4 (N13853, N13848, N5849, N1983, N9058);
nor NOR4 (N13854, N13851, N2328, N10071, N5235);
buf BUF1 (N13855, N13842);
xor XOR2 (N13856, N13854, N6275);
and AND4 (N13857, N13841, N8122, N9734, N4968);
xor XOR2 (N13858, N13855, N10538);
and AND3 (N13859, N13852, N11100, N6082);
xor XOR2 (N13860, N13856, N9844);
and AND3 (N13861, N13836, N5641, N4446);
nand NAND4 (N13862, N13843, N945, N5350, N10999);
not NOT1 (N13863, N13844);
or OR3 (N13864, N13860, N212, N13455);
buf BUF1 (N13865, N13861);
or OR3 (N13866, N13849, N2209, N6771);
nor NOR4 (N13867, N13859, N5605, N3879, N1532);
nand NAND3 (N13868, N13857, N7590, N6390);
and AND4 (N13869, N13846, N7743, N9494, N2821);
or OR2 (N13870, N13858, N4671);
not NOT1 (N13871, N13869);
nor NOR3 (N13872, N13865, N10672, N8132);
and AND4 (N13873, N13870, N13774, N3521, N10562);
buf BUF1 (N13874, N13867);
and AND4 (N13875, N13874, N6280, N6708, N13577);
xor XOR2 (N13876, N13864, N1568);
nand NAND2 (N13877, N13876, N8623);
not NOT1 (N13878, N13875);
xor XOR2 (N13879, N13863, N12608);
nor NOR3 (N13880, N13866, N1417, N9434);
not NOT1 (N13881, N13873);
or OR4 (N13882, N13853, N9938, N8440, N9742);
nand NAND4 (N13883, N13871, N3664, N1908, N8417);
or OR4 (N13884, N13882, N2378, N6701, N13464);
not NOT1 (N13885, N13881);
nand NAND4 (N13886, N13862, N8039, N3928, N13301);
not NOT1 (N13887, N13885);
xor XOR2 (N13888, N13883, N13317);
and AND4 (N13889, N13872, N18, N5840, N263);
nand NAND4 (N13890, N13877, N2564, N2720, N3143);
nor NOR3 (N13891, N13890, N98, N2514);
or OR3 (N13892, N13868, N8890, N513);
or OR2 (N13893, N13889, N12947);
or OR3 (N13894, N13880, N9955, N3471);
and AND4 (N13895, N13894, N5029, N8627, N9837);
buf BUF1 (N13896, N13878);
buf BUF1 (N13897, N13884);
and AND4 (N13898, N13886, N13427, N1840, N2617);
or OR4 (N13899, N13895, N9657, N9568, N3793);
xor XOR2 (N13900, N13879, N3170);
not NOT1 (N13901, N13898);
and AND3 (N13902, N13893, N3635, N1567);
nand NAND4 (N13903, N13892, N6957, N5844, N4617);
nor NOR3 (N13904, N13903, N1055, N8020);
buf BUF1 (N13905, N13888);
or OR3 (N13906, N13902, N4201, N4462);
nand NAND4 (N13907, N13900, N8889, N7608, N8);
buf BUF1 (N13908, N13905);
not NOT1 (N13909, N13904);
xor XOR2 (N13910, N13909, N9489);
and AND3 (N13911, N13896, N13842, N13406);
nand NAND2 (N13912, N13910, N12938);
xor XOR2 (N13913, N13899, N11776);
and AND3 (N13914, N13887, N7698, N1444);
nor NOR4 (N13915, N13913, N11512, N10476, N5441);
nor NOR3 (N13916, N13915, N10804, N4535);
buf BUF1 (N13917, N13912);
nand NAND2 (N13918, N13907, N877);
buf BUF1 (N13919, N13891);
and AND3 (N13920, N13897, N5931, N3633);
xor XOR2 (N13921, N13919, N10235);
nor NOR2 (N13922, N13917, N2846);
nor NOR3 (N13923, N13920, N12796, N8708);
nor NOR4 (N13924, N13916, N4722, N7329, N8409);
and AND3 (N13925, N13923, N1204, N4835);
nor NOR4 (N13926, N13922, N3971, N5499, N5952);
and AND2 (N13927, N13901, N9959);
and AND4 (N13928, N13906, N7585, N12449, N11927);
or OR3 (N13929, N13928, N12578, N7170);
or OR2 (N13930, N13924, N2599);
or OR4 (N13931, N13911, N9439, N8192, N6134);
and AND4 (N13932, N13931, N6083, N6292, N3761);
xor XOR2 (N13933, N13918, N10344);
nor NOR3 (N13934, N13926, N1089, N4654);
not NOT1 (N13935, N13930);
xor XOR2 (N13936, N13934, N6827);
nand NAND2 (N13937, N13927, N8166);
and AND4 (N13938, N13935, N1309, N156, N3155);
buf BUF1 (N13939, N13932);
and AND3 (N13940, N13925, N744, N7720);
and AND2 (N13941, N13929, N3959);
and AND2 (N13942, N13908, N9693);
nor NOR4 (N13943, N13936, N635, N4328, N4634);
not NOT1 (N13944, N13938);
nand NAND2 (N13945, N13943, N6231);
buf BUF1 (N13946, N13941);
not NOT1 (N13947, N13933);
xor XOR2 (N13948, N13940, N13018);
xor XOR2 (N13949, N13946, N8311);
not NOT1 (N13950, N13942);
and AND2 (N13951, N13939, N8060);
buf BUF1 (N13952, N13937);
or OR3 (N13953, N13914, N7419, N2999);
buf BUF1 (N13954, N13921);
xor XOR2 (N13955, N13950, N8227);
xor XOR2 (N13956, N13953, N13177);
xor XOR2 (N13957, N13945, N13943);
xor XOR2 (N13958, N13957, N13786);
buf BUF1 (N13959, N13952);
or OR2 (N13960, N13944, N3749);
nand NAND4 (N13961, N13955, N1144, N5194, N7096);
xor XOR2 (N13962, N13959, N3432);
nand NAND2 (N13963, N13948, N10696);
buf BUF1 (N13964, N13960);
buf BUF1 (N13965, N13951);
nand NAND4 (N13966, N13964, N8293, N1004, N5901);
xor XOR2 (N13967, N13956, N6174);
nor NOR3 (N13968, N13954, N8830, N6764);
and AND2 (N13969, N13963, N6486);
xor XOR2 (N13970, N13968, N11221);
nor NOR3 (N13971, N13966, N9617, N9211);
or OR2 (N13972, N13949, N13545);
buf BUF1 (N13973, N13969);
or OR4 (N13974, N13965, N3140, N13117, N10217);
buf BUF1 (N13975, N13971);
nand NAND2 (N13976, N13973, N13246);
or OR4 (N13977, N13975, N6437, N12599, N5791);
not NOT1 (N13978, N13967);
xor XOR2 (N13979, N13972, N12148);
buf BUF1 (N13980, N13977);
not NOT1 (N13981, N13962);
and AND4 (N13982, N13961, N3637, N9523, N8206);
buf BUF1 (N13983, N13958);
and AND2 (N13984, N13979, N1117);
not NOT1 (N13985, N13974);
buf BUF1 (N13986, N13978);
buf BUF1 (N13987, N13986);
not NOT1 (N13988, N13976);
nand NAND2 (N13989, N13984, N12046);
and AND2 (N13990, N13947, N1189);
nand NAND2 (N13991, N13988, N1085);
nor NOR3 (N13992, N13983, N1829, N13306);
and AND3 (N13993, N13981, N6134, N1208);
xor XOR2 (N13994, N13990, N3064);
xor XOR2 (N13995, N13985, N13476);
not NOT1 (N13996, N13995);
or OR3 (N13997, N13980, N9185, N12506);
and AND4 (N13998, N13994, N12456, N11601, N5700);
not NOT1 (N13999, N13998);
or OR3 (N14000, N13992, N8905, N1214);
not NOT1 (N14001, N13996);
xor XOR2 (N14002, N13991, N6766);
nor NOR2 (N14003, N13993, N2735);
not NOT1 (N14004, N13987);
xor XOR2 (N14005, N13999, N8999);
xor XOR2 (N14006, N13997, N8848);
and AND3 (N14007, N14002, N4354, N13189);
xor XOR2 (N14008, N14000, N577);
and AND2 (N14009, N14007, N8553);
not NOT1 (N14010, N13989);
buf BUF1 (N14011, N14001);
buf BUF1 (N14012, N13982);
buf BUF1 (N14013, N14011);
nand NAND4 (N14014, N14013, N10320, N12609, N9450);
xor XOR2 (N14015, N14003, N1378);
xor XOR2 (N14016, N14014, N7417);
not NOT1 (N14017, N14008);
not NOT1 (N14018, N13970);
nand NAND2 (N14019, N14005, N11620);
and AND3 (N14020, N14010, N11955, N9827);
not NOT1 (N14021, N14020);
nand NAND3 (N14022, N14016, N2645, N13903);
buf BUF1 (N14023, N14006);
or OR4 (N14024, N14015, N3765, N12620, N10636);
not NOT1 (N14025, N14004);
not NOT1 (N14026, N14017);
xor XOR2 (N14027, N14019, N13686);
and AND2 (N14028, N14018, N2443);
or OR3 (N14029, N14025, N2214, N7147);
nor NOR3 (N14030, N14009, N12327, N3113);
and AND2 (N14031, N14029, N10757);
xor XOR2 (N14032, N14022, N11340);
buf BUF1 (N14033, N14030);
not NOT1 (N14034, N14012);
and AND4 (N14035, N14034, N7786, N4348, N55);
nand NAND2 (N14036, N14026, N2374);
nor NOR4 (N14037, N14027, N13253, N11116, N4765);
nand NAND3 (N14038, N14031, N10934, N8359);
buf BUF1 (N14039, N14023);
buf BUF1 (N14040, N14021);
buf BUF1 (N14041, N14033);
or OR2 (N14042, N14038, N2716);
xor XOR2 (N14043, N14032, N13591);
and AND3 (N14044, N14035, N5790, N1855);
and AND3 (N14045, N14037, N9966, N7107);
nand NAND2 (N14046, N14044, N3419);
or OR4 (N14047, N14042, N10991, N7951, N7644);
not NOT1 (N14048, N14043);
xor XOR2 (N14049, N14036, N9868);
not NOT1 (N14050, N14049);
nand NAND3 (N14051, N14050, N6121, N6749);
nor NOR4 (N14052, N14041, N1643, N1566, N2093);
not NOT1 (N14053, N14048);
nand NAND3 (N14054, N14028, N9408, N6908);
not NOT1 (N14055, N14046);
nand NAND2 (N14056, N14054, N10737);
xor XOR2 (N14057, N14047, N12976);
buf BUF1 (N14058, N14039);
or OR4 (N14059, N14057, N6326, N10480, N5427);
nand NAND3 (N14060, N14024, N5692, N432);
nand NAND2 (N14061, N14045, N3857);
xor XOR2 (N14062, N14061, N12681);
buf BUF1 (N14063, N14055);
xor XOR2 (N14064, N14040, N1462);
buf BUF1 (N14065, N14059);
xor XOR2 (N14066, N14058, N6062);
nand NAND4 (N14067, N14060, N11861, N5168, N6807);
or OR4 (N14068, N14065, N3768, N4621, N4129);
or OR4 (N14069, N14067, N12489, N5467, N3584);
nor NOR4 (N14070, N14052, N2638, N13764, N9218);
xor XOR2 (N14071, N14053, N3363);
and AND2 (N14072, N14056, N4034);
nor NOR4 (N14073, N14071, N10126, N5807, N4854);
nor NOR4 (N14074, N14066, N8547, N6342, N4488);
or OR4 (N14075, N14070, N4074, N11407, N8355);
nor NOR2 (N14076, N14051, N1938);
xor XOR2 (N14077, N14076, N2948);
buf BUF1 (N14078, N14064);
and AND3 (N14079, N14069, N5210, N3299);
nand NAND3 (N14080, N14079, N3986, N9350);
buf BUF1 (N14081, N14072);
xor XOR2 (N14082, N14073, N10854);
xor XOR2 (N14083, N14063, N10557);
xor XOR2 (N14084, N14082, N11058);
xor XOR2 (N14085, N14084, N4689);
and AND2 (N14086, N14083, N2980);
buf BUF1 (N14087, N14062);
and AND2 (N14088, N14077, N8883);
nand NAND4 (N14089, N14068, N5386, N13715, N12612);
not NOT1 (N14090, N14085);
or OR2 (N14091, N14090, N2234);
nand NAND2 (N14092, N14086, N4059);
buf BUF1 (N14093, N14092);
nor NOR2 (N14094, N14080, N8243);
or OR3 (N14095, N14081, N1476, N2204);
and AND3 (N14096, N14094, N6845, N11890);
and AND3 (N14097, N14078, N10098, N4228);
not NOT1 (N14098, N14075);
nor NOR2 (N14099, N14097, N11659);
and AND3 (N14100, N14095, N9595, N8983);
nand NAND3 (N14101, N14089, N9223, N4942);
nor NOR4 (N14102, N14093, N5556, N13878, N7441);
buf BUF1 (N14103, N14098);
xor XOR2 (N14104, N14099, N9273);
nand NAND3 (N14105, N14088, N10943, N12090);
nor NOR3 (N14106, N14103, N8415, N10302);
not NOT1 (N14107, N14106);
nand NAND3 (N14108, N14101, N6248, N5535);
or OR2 (N14109, N14107, N10405);
buf BUF1 (N14110, N14091);
nor NOR2 (N14111, N14074, N11394);
not NOT1 (N14112, N14102);
nor NOR3 (N14113, N14111, N12368, N30);
buf BUF1 (N14114, N14087);
not NOT1 (N14115, N14100);
xor XOR2 (N14116, N14113, N8921);
buf BUF1 (N14117, N14096);
and AND4 (N14118, N14105, N5749, N108, N4448);
not NOT1 (N14119, N14109);
not NOT1 (N14120, N14118);
xor XOR2 (N14121, N14120, N9345);
nor NOR4 (N14122, N14121, N11384, N9255, N9847);
buf BUF1 (N14123, N14104);
and AND2 (N14124, N14119, N811);
or OR3 (N14125, N14117, N13225, N1060);
or OR2 (N14126, N14114, N981);
nand NAND4 (N14127, N14123, N2298, N10817, N13370);
or OR2 (N14128, N14110, N10420);
buf BUF1 (N14129, N14125);
nand NAND4 (N14130, N14112, N2156, N8988, N5024);
nor NOR4 (N14131, N14122, N8017, N11485, N10596);
buf BUF1 (N14132, N14116);
nor NOR2 (N14133, N14128, N7366);
not NOT1 (N14134, N14115);
and AND4 (N14135, N14132, N5326, N2215, N6768);
buf BUF1 (N14136, N14134);
or OR2 (N14137, N14133, N13711);
nor NOR2 (N14138, N14130, N5106);
nor NOR4 (N14139, N14136, N7906, N11888, N13463);
nand NAND2 (N14140, N14124, N5236);
buf BUF1 (N14141, N14135);
buf BUF1 (N14142, N14126);
buf BUF1 (N14143, N14142);
buf BUF1 (N14144, N14129);
nand NAND2 (N14145, N14144, N12584);
not NOT1 (N14146, N14108);
xor XOR2 (N14147, N14145, N10677);
nand NAND4 (N14148, N14141, N2990, N260, N8948);
xor XOR2 (N14149, N14146, N1142);
and AND2 (N14150, N14143, N3523);
buf BUF1 (N14151, N14127);
xor XOR2 (N14152, N14131, N4839);
or OR3 (N14153, N14148, N9889, N7217);
xor XOR2 (N14154, N14151, N1649);
xor XOR2 (N14155, N14150, N723);
not NOT1 (N14156, N14137);
xor XOR2 (N14157, N14140, N804);
or OR2 (N14158, N14154, N6907);
or OR3 (N14159, N14158, N10737, N10015);
buf BUF1 (N14160, N14139);
buf BUF1 (N14161, N14147);
buf BUF1 (N14162, N14159);
nor NOR3 (N14163, N14153, N4337, N10661);
and AND3 (N14164, N14149, N12931, N2238);
or OR4 (N14165, N14162, N9100, N347, N10147);
and AND2 (N14166, N14156, N1607);
and AND4 (N14167, N14165, N2413, N3546, N5578);
nand NAND2 (N14168, N14152, N4214);
buf BUF1 (N14169, N14138);
and AND3 (N14170, N14168, N10028, N6310);
nor NOR3 (N14171, N14157, N4316, N2416);
and AND4 (N14172, N14166, N10830, N13183, N1231);
not NOT1 (N14173, N14171);
or OR3 (N14174, N14172, N894, N3635);
nor NOR2 (N14175, N14160, N3037);
and AND3 (N14176, N14163, N13502, N6832);
and AND4 (N14177, N14173, N1767, N8672, N13570);
nor NOR2 (N14178, N14175, N548);
xor XOR2 (N14179, N14167, N13912);
and AND3 (N14180, N14155, N6323, N4210);
xor XOR2 (N14181, N14164, N11335);
buf BUF1 (N14182, N14176);
buf BUF1 (N14183, N14170);
buf BUF1 (N14184, N14183);
xor XOR2 (N14185, N14174, N90);
buf BUF1 (N14186, N14185);
or OR3 (N14187, N14178, N9389, N8030);
and AND4 (N14188, N14177, N148, N6295, N1259);
nand NAND4 (N14189, N14182, N6807, N6751, N7666);
buf BUF1 (N14190, N14186);
and AND3 (N14191, N14188, N7785, N13649);
and AND2 (N14192, N14169, N2835);
buf BUF1 (N14193, N14161);
nand NAND3 (N14194, N14180, N931, N11871);
not NOT1 (N14195, N14190);
buf BUF1 (N14196, N14189);
nand NAND3 (N14197, N14179, N8618, N5121);
xor XOR2 (N14198, N14187, N13058);
and AND4 (N14199, N14184, N8437, N6468, N8922);
nor NOR2 (N14200, N14199, N10780);
nor NOR2 (N14201, N14191, N7424);
nor NOR3 (N14202, N14194, N2440, N13988);
xor XOR2 (N14203, N14192, N2089);
and AND3 (N14204, N14201, N7493, N3117);
not NOT1 (N14205, N14195);
and AND2 (N14206, N14197, N13413);
xor XOR2 (N14207, N14198, N1397);
or OR3 (N14208, N14204, N13906, N5736);
nor NOR2 (N14209, N14206, N6647);
nand NAND3 (N14210, N14205, N2672, N898);
and AND3 (N14211, N14193, N13982, N13819);
nand NAND2 (N14212, N14203, N14193);
xor XOR2 (N14213, N14208, N7408);
nor NOR2 (N14214, N14181, N8925);
or OR2 (N14215, N14196, N4159);
nand NAND4 (N14216, N14200, N13139, N8279, N9714);
not NOT1 (N14217, N14213);
not NOT1 (N14218, N14212);
or OR4 (N14219, N14218, N9088, N2855, N2818);
or OR3 (N14220, N14207, N7259, N7273);
xor XOR2 (N14221, N14210, N1367);
nand NAND2 (N14222, N14220, N1196);
or OR2 (N14223, N14214, N9516);
not NOT1 (N14224, N14221);
xor XOR2 (N14225, N14215, N6040);
nor NOR3 (N14226, N14223, N11807, N9435);
not NOT1 (N14227, N14209);
xor XOR2 (N14228, N14222, N7120);
xor XOR2 (N14229, N14219, N1824);
nand NAND2 (N14230, N14202, N5884);
nand NAND3 (N14231, N14227, N3793, N9624);
buf BUF1 (N14232, N14226);
xor XOR2 (N14233, N14232, N778);
not NOT1 (N14234, N14231);
nand NAND2 (N14235, N14229, N2611);
or OR2 (N14236, N14225, N6724);
nor NOR4 (N14237, N14230, N4353, N9476, N3565);
nor NOR2 (N14238, N14234, N11731);
or OR4 (N14239, N14228, N13287, N6600, N12192);
and AND4 (N14240, N14216, N8783, N8707, N10338);
and AND3 (N14241, N14238, N2240, N4091);
xor XOR2 (N14242, N14211, N4131);
not NOT1 (N14243, N14224);
and AND4 (N14244, N14236, N3590, N131, N9109);
and AND2 (N14245, N14244, N7350);
not NOT1 (N14246, N14241);
nor NOR4 (N14247, N14239, N11984, N12927, N2341);
nor NOR3 (N14248, N14242, N14148, N3920);
and AND3 (N14249, N14243, N3682, N4107);
nor NOR4 (N14250, N14235, N5842, N5764, N8881);
nor NOR4 (N14251, N14250, N11952, N13147, N13178);
or OR3 (N14252, N14233, N3927, N10465);
buf BUF1 (N14253, N14247);
and AND2 (N14254, N14248, N13478);
buf BUF1 (N14255, N14237);
not NOT1 (N14256, N14217);
buf BUF1 (N14257, N14255);
not NOT1 (N14258, N14252);
buf BUF1 (N14259, N14249);
and AND2 (N14260, N14246, N9642);
or OR3 (N14261, N14259, N10769, N12388);
buf BUF1 (N14262, N14240);
xor XOR2 (N14263, N14262, N7157);
xor XOR2 (N14264, N14256, N7475);
and AND4 (N14265, N14264, N13043, N4201, N2709);
or OR4 (N14266, N14265, N2707, N10401, N5430);
and AND3 (N14267, N14245, N7600, N5666);
and AND3 (N14268, N14251, N646, N427);
buf BUF1 (N14269, N14253);
or OR3 (N14270, N14263, N1300, N11053);
and AND2 (N14271, N14268, N10947);
nor NOR3 (N14272, N14258, N4867, N11138);
nor NOR2 (N14273, N14271, N7490);
and AND2 (N14274, N14272, N10361);
not NOT1 (N14275, N14254);
not NOT1 (N14276, N14275);
or OR4 (N14277, N14274, N2590, N5333, N12692);
or OR4 (N14278, N14269, N11708, N11886, N12087);
nor NOR4 (N14279, N14267, N14048, N9077, N12853);
and AND2 (N14280, N14273, N2506);
buf BUF1 (N14281, N14279);
xor XOR2 (N14282, N14276, N887);
and AND3 (N14283, N14257, N637, N2674);
buf BUF1 (N14284, N14260);
buf BUF1 (N14285, N14282);
buf BUF1 (N14286, N14280);
and AND3 (N14287, N14284, N6585, N9442);
or OR2 (N14288, N14285, N3255);
or OR2 (N14289, N14286, N4986);
buf BUF1 (N14290, N14261);
nor NOR4 (N14291, N14289, N3416, N1845, N11004);
or OR3 (N14292, N14277, N5008, N11351);
or OR4 (N14293, N14288, N13492, N880, N2581);
xor XOR2 (N14294, N14291, N8888);
and AND4 (N14295, N14290, N6226, N1627, N8188);
not NOT1 (N14296, N14281);
nand NAND4 (N14297, N14278, N5400, N3834, N1555);
xor XOR2 (N14298, N14297, N11599);
and AND2 (N14299, N14292, N9554);
nor NOR3 (N14300, N14283, N7361, N10345);
or OR2 (N14301, N14299, N7412);
not NOT1 (N14302, N14295);
nand NAND3 (N14303, N14302, N2902, N7118);
nor NOR4 (N14304, N14293, N7152, N8605, N13119);
xor XOR2 (N14305, N14296, N9392);
nor NOR3 (N14306, N14287, N7861, N923);
not NOT1 (N14307, N14306);
nand NAND4 (N14308, N14303, N10399, N360, N12656);
nand NAND4 (N14309, N14266, N6337, N9838, N7651);
xor XOR2 (N14310, N14298, N9133);
buf BUF1 (N14311, N14301);
xor XOR2 (N14312, N14304, N5553);
buf BUF1 (N14313, N14305);
nor NOR2 (N14314, N14307, N2903);
and AND3 (N14315, N14309, N6781, N5561);
or OR3 (N14316, N14294, N13017, N813);
buf BUF1 (N14317, N14310);
nor NOR2 (N14318, N14270, N4167);
xor XOR2 (N14319, N14308, N10671);
not NOT1 (N14320, N14311);
nor NOR4 (N14321, N14317, N2739, N7582, N14231);
xor XOR2 (N14322, N14300, N3805);
buf BUF1 (N14323, N14319);
nand NAND2 (N14324, N14323, N9416);
or OR2 (N14325, N14321, N1164);
or OR3 (N14326, N14313, N5078, N4600);
buf BUF1 (N14327, N14320);
and AND4 (N14328, N14324, N1444, N7665, N3993);
or OR3 (N14329, N14312, N9309, N2543);
and AND4 (N14330, N14315, N6116, N266, N2171);
not NOT1 (N14331, N14328);
or OR3 (N14332, N14329, N11970, N5551);
xor XOR2 (N14333, N14316, N722);
xor XOR2 (N14334, N14322, N10991);
nand NAND2 (N14335, N14333, N6394);
not NOT1 (N14336, N14335);
or OR4 (N14337, N14332, N5472, N3765, N3644);
buf BUF1 (N14338, N14325);
nor NOR2 (N14339, N14338, N6121);
and AND2 (N14340, N14330, N544);
buf BUF1 (N14341, N14340);
or OR3 (N14342, N14334, N9852, N1284);
nand NAND2 (N14343, N14341, N2794);
xor XOR2 (N14344, N14337, N14024);
and AND4 (N14345, N14343, N4001, N2774, N5378);
nand NAND2 (N14346, N14331, N9839);
and AND3 (N14347, N14344, N11710, N1685);
xor XOR2 (N14348, N14347, N4896);
not NOT1 (N14349, N14327);
nand NAND3 (N14350, N14345, N13026, N1858);
nand NAND3 (N14351, N14318, N13012, N6591);
not NOT1 (N14352, N14348);
xor XOR2 (N14353, N14349, N4808);
buf BUF1 (N14354, N14314);
or OR4 (N14355, N14342, N7233, N829, N2730);
buf BUF1 (N14356, N14355);
nor NOR4 (N14357, N14353, N2860, N3628, N13006);
xor XOR2 (N14358, N14351, N2292);
nand NAND4 (N14359, N14354, N5522, N13552, N12885);
not NOT1 (N14360, N14336);
or OR4 (N14361, N14356, N9722, N13458, N4721);
or OR4 (N14362, N14326, N9630, N1378, N13045);
buf BUF1 (N14363, N14339);
buf BUF1 (N14364, N14346);
nand NAND3 (N14365, N14352, N5183, N10881);
xor XOR2 (N14366, N14359, N6443);
xor XOR2 (N14367, N14358, N11058);
xor XOR2 (N14368, N14350, N11370);
or OR3 (N14369, N14361, N4888, N11265);
xor XOR2 (N14370, N14357, N6511);
not NOT1 (N14371, N14370);
not NOT1 (N14372, N14365);
xor XOR2 (N14373, N14362, N9714);
or OR3 (N14374, N14364, N10220, N5452);
and AND4 (N14375, N14371, N8405, N1783, N6102);
xor XOR2 (N14376, N14363, N5764);
or OR2 (N14377, N14372, N9791);
not NOT1 (N14378, N14360);
not NOT1 (N14379, N14367);
xor XOR2 (N14380, N14366, N11916);
not NOT1 (N14381, N14380);
or OR4 (N14382, N14377, N6832, N13018, N10894);
nand NAND3 (N14383, N14379, N4520, N10718);
and AND4 (N14384, N14378, N184, N4222, N3015);
nand NAND4 (N14385, N14382, N7120, N13008, N6482);
not NOT1 (N14386, N14384);
and AND4 (N14387, N14369, N2620, N7197, N278);
and AND3 (N14388, N14386, N4355, N6525);
nor NOR4 (N14389, N14383, N923, N14009, N9516);
xor XOR2 (N14390, N14368, N4201);
not NOT1 (N14391, N14390);
or OR2 (N14392, N14385, N5821);
xor XOR2 (N14393, N14392, N5814);
nor NOR2 (N14394, N14381, N7207);
nor NOR2 (N14395, N14374, N6876);
and AND2 (N14396, N14389, N2690);
xor XOR2 (N14397, N14376, N266);
buf BUF1 (N14398, N14395);
not NOT1 (N14399, N14398);
buf BUF1 (N14400, N14394);
buf BUF1 (N14401, N14400);
or OR2 (N14402, N14401, N13630);
and AND2 (N14403, N14387, N8436);
or OR4 (N14404, N14393, N3054, N8227, N11982);
not NOT1 (N14405, N14388);
buf BUF1 (N14406, N14373);
nand NAND2 (N14407, N14404, N9526);
or OR4 (N14408, N14375, N14314, N9965, N12593);
not NOT1 (N14409, N14405);
and AND4 (N14410, N14402, N1611, N8131, N14256);
or OR4 (N14411, N14408, N9336, N10611, N683);
or OR2 (N14412, N14391, N14181);
xor XOR2 (N14413, N14396, N727);
xor XOR2 (N14414, N14411, N8546);
not NOT1 (N14415, N14407);
and AND2 (N14416, N14399, N10082);
or OR2 (N14417, N14410, N4559);
nor NOR4 (N14418, N14413, N6057, N5588, N584);
and AND4 (N14419, N14403, N10882, N8976, N9928);
nand NAND3 (N14420, N14418, N2061, N1463);
nand NAND3 (N14421, N14420, N11858, N5570);
nand NAND2 (N14422, N14421, N7565);
nand NAND3 (N14423, N14412, N8998, N10388);
xor XOR2 (N14424, N14406, N818);
xor XOR2 (N14425, N14414, N2356);
not NOT1 (N14426, N14425);
xor XOR2 (N14427, N14415, N10975);
not NOT1 (N14428, N14417);
not NOT1 (N14429, N14416);
or OR2 (N14430, N14422, N8344);
not NOT1 (N14431, N14423);
xor XOR2 (N14432, N14426, N12667);
nor NOR3 (N14433, N14419, N13468, N3826);
xor XOR2 (N14434, N14427, N1187);
buf BUF1 (N14435, N14409);
and AND2 (N14436, N14430, N2375);
or OR3 (N14437, N14434, N10482, N9760);
nor NOR4 (N14438, N14424, N8631, N8494, N2306);
and AND3 (N14439, N14432, N10644, N3153);
and AND4 (N14440, N14437, N653, N3835, N13505);
nand NAND2 (N14441, N14397, N2725);
nand NAND4 (N14442, N14431, N7426, N2342, N4386);
nor NOR2 (N14443, N14435, N11306);
nand NAND4 (N14444, N14442, N14381, N8236, N14378);
nand NAND4 (N14445, N14438, N6784, N14443, N8572);
nand NAND4 (N14446, N345, N9413, N2212, N5161);
nor NOR2 (N14447, N14439, N8580);
xor XOR2 (N14448, N14446, N5275);
or OR4 (N14449, N14436, N8949, N7688, N10542);
or OR3 (N14450, N14441, N4243, N6494);
xor XOR2 (N14451, N14440, N13383);
nor NOR2 (N14452, N14450, N5732);
nand NAND3 (N14453, N14448, N1146, N4980);
and AND3 (N14454, N14428, N10982, N2975);
not NOT1 (N14455, N14445);
and AND4 (N14456, N14454, N4019, N3014, N3855);
and AND4 (N14457, N14433, N6729, N12963, N646);
nand NAND2 (N14458, N14452, N5703);
and AND3 (N14459, N14451, N10900, N13446);
xor XOR2 (N14460, N14459, N10140);
and AND4 (N14461, N14460, N757, N9453, N10879);
or OR3 (N14462, N14447, N621, N6291);
not NOT1 (N14463, N14462);
buf BUF1 (N14464, N14429);
and AND4 (N14465, N14461, N3543, N806, N1280);
xor XOR2 (N14466, N14463, N12761);
xor XOR2 (N14467, N14453, N1807);
nor NOR3 (N14468, N14455, N5956, N14410);
buf BUF1 (N14469, N14465);
nor NOR2 (N14470, N14467, N7715);
not NOT1 (N14471, N14470);
not NOT1 (N14472, N14449);
and AND2 (N14473, N14464, N7677);
buf BUF1 (N14474, N14466);
not NOT1 (N14475, N14457);
buf BUF1 (N14476, N14471);
xor XOR2 (N14477, N14456, N5165);
nor NOR3 (N14478, N14475, N5890, N13135);
not NOT1 (N14479, N14444);
not NOT1 (N14480, N14472);
nand NAND2 (N14481, N14468, N9446);
buf BUF1 (N14482, N14479);
or OR4 (N14483, N14482, N7621, N7607, N1187);
nor NOR2 (N14484, N14473, N6129);
nor NOR4 (N14485, N14458, N13365, N6804, N4034);
or OR2 (N14486, N14485, N13035);
xor XOR2 (N14487, N14476, N11817);
nand NAND3 (N14488, N14487, N3699, N9102);
not NOT1 (N14489, N14483);
and AND2 (N14490, N14489, N3592);
nor NOR3 (N14491, N14486, N3967, N5093);
and AND3 (N14492, N14474, N9860, N5143);
or OR3 (N14493, N14491, N7058, N2448);
or OR3 (N14494, N14484, N7490, N12086);
nor NOR4 (N14495, N14490, N3770, N11543, N11695);
or OR2 (N14496, N14478, N5092);
nor NOR3 (N14497, N14492, N13111, N11078);
or OR3 (N14498, N14494, N7712, N3887);
nand NAND3 (N14499, N14496, N5288, N1950);
not NOT1 (N14500, N14469);
nand NAND2 (N14501, N14495, N11771);
not NOT1 (N14502, N14493);
buf BUF1 (N14503, N14488);
not NOT1 (N14504, N14481);
nor NOR3 (N14505, N14504, N11716, N130);
buf BUF1 (N14506, N14480);
xor XOR2 (N14507, N14497, N8212);
or OR3 (N14508, N14477, N4337, N7863);
and AND2 (N14509, N14506, N822);
not NOT1 (N14510, N14505);
or OR4 (N14511, N14502, N14286, N11822, N5001);
and AND3 (N14512, N14507, N5498, N7377);
xor XOR2 (N14513, N14510, N12674);
not NOT1 (N14514, N14500);
buf BUF1 (N14515, N14503);
or OR3 (N14516, N14509, N10456, N12267);
or OR2 (N14517, N14508, N4808);
xor XOR2 (N14518, N14511, N11823);
nand NAND2 (N14519, N14499, N3855);
or OR4 (N14520, N14515, N180, N11683, N9743);
nor NOR4 (N14521, N14516, N6898, N10134, N9410);
nor NOR4 (N14522, N14498, N12717, N8478, N3224);
and AND4 (N14523, N14522, N2862, N1245, N3510);
buf BUF1 (N14524, N14517);
xor XOR2 (N14525, N14513, N9452);
nand NAND4 (N14526, N14525, N12447, N2825, N12604);
nor NOR3 (N14527, N14518, N5697, N7007);
and AND3 (N14528, N14527, N11604, N12286);
buf BUF1 (N14529, N14526);
buf BUF1 (N14530, N14523);
nand NAND3 (N14531, N14528, N7895, N2930);
buf BUF1 (N14532, N14521);
not NOT1 (N14533, N14532);
or OR4 (N14534, N14519, N12180, N11749, N431);
not NOT1 (N14535, N14529);
nor NOR4 (N14536, N14533, N6698, N5706, N2907);
nor NOR2 (N14537, N14530, N4596);
or OR2 (N14538, N14520, N11703);
nand NAND4 (N14539, N14538, N5167, N6471, N4678);
nand NAND4 (N14540, N14537, N13753, N1641, N11856);
or OR3 (N14541, N14524, N5667, N8483);
nand NAND4 (N14542, N14512, N7081, N2825, N781);
and AND4 (N14543, N14501, N3152, N6955, N3582);
or OR4 (N14544, N14542, N715, N5369, N2309);
not NOT1 (N14545, N14531);
buf BUF1 (N14546, N14534);
and AND4 (N14547, N14545, N2659, N2136, N8339);
and AND2 (N14548, N14535, N13543);
not NOT1 (N14549, N14547);
nand NAND4 (N14550, N14539, N6303, N2225, N1049);
nor NOR4 (N14551, N14549, N10553, N12627, N22);
buf BUF1 (N14552, N14541);
xor XOR2 (N14553, N14551, N4823);
nor NOR4 (N14554, N14552, N14467, N8570, N1724);
xor XOR2 (N14555, N14550, N6449);
nor NOR3 (N14556, N14548, N7547, N14478);
not NOT1 (N14557, N14546);
nand NAND2 (N14558, N14553, N9515);
or OR3 (N14559, N14557, N7613, N1945);
xor XOR2 (N14560, N14540, N6537);
nand NAND2 (N14561, N14544, N8580);
not NOT1 (N14562, N14559);
not NOT1 (N14563, N14561);
not NOT1 (N14564, N14555);
or OR2 (N14565, N14560, N3066);
nand NAND4 (N14566, N14563, N10178, N12592, N9476);
nor NOR4 (N14567, N14566, N12889, N1406, N9459);
and AND2 (N14568, N14565, N3074);
nand NAND3 (N14569, N14514, N13460, N11031);
or OR3 (N14570, N14558, N3778, N3314);
xor XOR2 (N14571, N14536, N9327);
or OR4 (N14572, N14569, N12464, N4513, N6818);
xor XOR2 (N14573, N14568, N529);
buf BUF1 (N14574, N14554);
nor NOR4 (N14575, N14573, N12820, N10033, N6461);
buf BUF1 (N14576, N14562);
nand NAND2 (N14577, N14576, N733);
not NOT1 (N14578, N14577);
nor NOR2 (N14579, N14564, N10253);
or OR2 (N14580, N14572, N1961);
or OR3 (N14581, N14543, N4773, N10294);
xor XOR2 (N14582, N14571, N10579);
xor XOR2 (N14583, N14578, N7876);
not NOT1 (N14584, N14575);
and AND3 (N14585, N14579, N12035, N5254);
xor XOR2 (N14586, N14556, N3917);
nand NAND4 (N14587, N14582, N9509, N4768, N10784);
not NOT1 (N14588, N14584);
xor XOR2 (N14589, N14567, N5637);
and AND3 (N14590, N14583, N3016, N5018);
or OR2 (N14591, N14581, N13523);
or OR4 (N14592, N14570, N2523, N402, N3242);
and AND2 (N14593, N14588, N5978);
nor NOR4 (N14594, N14593, N8708, N5258, N1029);
or OR2 (N14595, N14585, N13928);
nor NOR4 (N14596, N14590, N1686, N12711, N4131);
and AND3 (N14597, N14594, N1605, N1368);
buf BUF1 (N14598, N14574);
not NOT1 (N14599, N14591);
buf BUF1 (N14600, N14598);
not NOT1 (N14601, N14597);
buf BUF1 (N14602, N14600);
and AND3 (N14603, N14602, N11240, N12098);
or OR2 (N14604, N14589, N3167);
nor NOR2 (N14605, N14580, N13556);
or OR4 (N14606, N14604, N11978, N7183, N9204);
xor XOR2 (N14607, N14599, N13363);
and AND4 (N14608, N14605, N9279, N7118, N9247);
nand NAND3 (N14609, N14601, N1333, N11285);
not NOT1 (N14610, N14587);
not NOT1 (N14611, N14603);
nand NAND3 (N14612, N14606, N8624, N7939);
nand NAND4 (N14613, N14595, N1091, N14001, N2615);
nor NOR3 (N14614, N14612, N14364, N1751);
buf BUF1 (N14615, N14614);
or OR4 (N14616, N14609, N3397, N7261, N10834);
buf BUF1 (N14617, N14613);
or OR4 (N14618, N14586, N14210, N4898, N1419);
nand NAND3 (N14619, N14616, N9406, N283);
or OR2 (N14620, N14611, N11232);
and AND2 (N14621, N14617, N6007);
and AND4 (N14622, N14620, N4591, N9852, N7225);
nand NAND3 (N14623, N14622, N6341, N14164);
and AND2 (N14624, N14610, N6785);
or OR3 (N14625, N14621, N5095, N14239);
buf BUF1 (N14626, N14596);
nand NAND4 (N14627, N14592, N12523, N9287, N2804);
not NOT1 (N14628, N14607);
nor NOR2 (N14629, N14608, N8613);
nor NOR2 (N14630, N14627, N9103);
buf BUF1 (N14631, N14624);
nor NOR3 (N14632, N14623, N4402, N10624);
and AND2 (N14633, N14630, N10406);
not NOT1 (N14634, N14628);
xor XOR2 (N14635, N14634, N2869);
or OR4 (N14636, N14615, N12157, N4348, N11127);
nand NAND4 (N14637, N14625, N10511, N13035, N10457);
buf BUF1 (N14638, N14635);
nor NOR2 (N14639, N14638, N7404);
nor NOR3 (N14640, N14636, N14637, N11667);
nor NOR3 (N14641, N14146, N13282, N5012);
not NOT1 (N14642, N14618);
xor XOR2 (N14643, N14641, N10268);
nor NOR2 (N14644, N14619, N8615);
nand NAND4 (N14645, N14629, N4900, N6942, N7130);
and AND2 (N14646, N14645, N771);
xor XOR2 (N14647, N14644, N7891);
nand NAND3 (N14648, N14646, N8833, N13148);
or OR3 (N14649, N14631, N8571, N12262);
nor NOR4 (N14650, N14649, N6916, N11760, N12974);
or OR2 (N14651, N14632, N12644);
nand NAND4 (N14652, N14643, N9819, N13446, N7448);
nand NAND3 (N14653, N14651, N5876, N2941);
nor NOR4 (N14654, N14640, N5830, N10806, N11851);
or OR2 (N14655, N14647, N2992);
and AND4 (N14656, N14626, N14574, N2504, N13124);
or OR3 (N14657, N14639, N10869, N6435);
nand NAND4 (N14658, N14657, N148, N1740, N9007);
and AND3 (N14659, N14654, N3179, N7702);
nor NOR4 (N14660, N14656, N11447, N5538, N7676);
not NOT1 (N14661, N14652);
not NOT1 (N14662, N14661);
buf BUF1 (N14663, N14659);
not NOT1 (N14664, N14662);
and AND4 (N14665, N14648, N9498, N14352, N14135);
buf BUF1 (N14666, N14665);
nor NOR2 (N14667, N14633, N4268);
and AND4 (N14668, N14642, N2456, N8183, N4935);
and AND2 (N14669, N14663, N9651);
xor XOR2 (N14670, N14666, N4206);
xor XOR2 (N14671, N14668, N9229);
or OR3 (N14672, N14655, N1879, N10347);
and AND4 (N14673, N14667, N8879, N8525, N2793);
or OR2 (N14674, N14664, N1939);
xor XOR2 (N14675, N14660, N2806);
xor XOR2 (N14676, N14669, N2827);
nor NOR4 (N14677, N14674, N2077, N6618, N4425);
nor NOR4 (N14678, N14677, N12509, N3825, N13524);
and AND2 (N14679, N14653, N3203);
nor NOR4 (N14680, N14676, N6133, N10374, N1363);
nor NOR4 (N14681, N14678, N4561, N5351, N11235);
nand NAND3 (N14682, N14675, N5528, N13720);
and AND3 (N14683, N14671, N2519, N13313);
not NOT1 (N14684, N14658);
buf BUF1 (N14685, N14673);
buf BUF1 (N14686, N14682);
nor NOR3 (N14687, N14670, N12940, N5691);
or OR3 (N14688, N14672, N9873, N5276);
nor NOR2 (N14689, N14685, N10555);
xor XOR2 (N14690, N14687, N13207);
or OR2 (N14691, N14684, N13501);
and AND3 (N14692, N14680, N4443, N5796);
not NOT1 (N14693, N14692);
and AND4 (N14694, N14686, N4650, N14015, N11325);
nand NAND3 (N14695, N14679, N13391, N1089);
xor XOR2 (N14696, N14691, N6113);
and AND2 (N14697, N14683, N13494);
or OR4 (N14698, N14689, N4386, N6600, N10564);
nand NAND2 (N14699, N14697, N10502);
xor XOR2 (N14700, N14694, N13151);
or OR2 (N14701, N14693, N12030);
and AND4 (N14702, N14701, N10391, N14449, N9137);
buf BUF1 (N14703, N14699);
and AND3 (N14704, N14681, N13581, N5711);
and AND3 (N14705, N14690, N11938, N6942);
not NOT1 (N14706, N14704);
nor NOR3 (N14707, N14705, N9053, N10601);
xor XOR2 (N14708, N14698, N2061);
nor NOR4 (N14709, N14688, N6914, N11242, N9826);
nand NAND3 (N14710, N14703, N12909, N9536);
and AND3 (N14711, N14707, N14097, N4036);
xor XOR2 (N14712, N14696, N2597);
or OR4 (N14713, N14706, N11876, N7116, N2539);
not NOT1 (N14714, N14700);
nor NOR3 (N14715, N14702, N10460, N12968);
nor NOR2 (N14716, N14715, N2071);
and AND3 (N14717, N14695, N10533, N206);
buf BUF1 (N14718, N14712);
and AND2 (N14719, N14713, N1300);
nor NOR4 (N14720, N14714, N9868, N7663, N287);
nor NOR3 (N14721, N14716, N6077, N10232);
nand NAND3 (N14722, N14719, N161, N7171);
and AND2 (N14723, N14718, N12496);
nand NAND3 (N14724, N14650, N7077, N2441);
or OR3 (N14725, N14709, N114, N6309);
or OR3 (N14726, N14722, N769, N2219);
buf BUF1 (N14727, N14711);
xor XOR2 (N14728, N14721, N12328);
buf BUF1 (N14729, N14726);
and AND2 (N14730, N14717, N1919);
xor XOR2 (N14731, N14729, N14555);
or OR3 (N14732, N14731, N8824, N14248);
buf BUF1 (N14733, N14732);
not NOT1 (N14734, N14730);
buf BUF1 (N14735, N14723);
or OR2 (N14736, N14724, N2980);
and AND3 (N14737, N14725, N1006, N12237);
not NOT1 (N14738, N14734);
buf BUF1 (N14739, N14710);
xor XOR2 (N14740, N14727, N1028);
not NOT1 (N14741, N14739);
xor XOR2 (N14742, N14738, N12369);
nand NAND2 (N14743, N14728, N4544);
not NOT1 (N14744, N14708);
or OR4 (N14745, N14733, N11566, N6191, N9235);
xor XOR2 (N14746, N14736, N6887);
xor XOR2 (N14747, N14735, N2231);
or OR2 (N14748, N14740, N233);
buf BUF1 (N14749, N14743);
nand NAND3 (N14750, N14747, N8191, N6692);
nor NOR2 (N14751, N14744, N12643);
buf BUF1 (N14752, N14745);
nand NAND3 (N14753, N14742, N12348, N2548);
nand NAND4 (N14754, N14746, N8972, N11761, N12998);
nor NOR3 (N14755, N14751, N1938, N13765);
or OR3 (N14756, N14720, N12207, N7664);
and AND2 (N14757, N14741, N13627);
not NOT1 (N14758, N14757);
buf BUF1 (N14759, N14756);
or OR2 (N14760, N14750, N14495);
or OR2 (N14761, N14748, N6840);
buf BUF1 (N14762, N14758);
and AND2 (N14763, N14737, N1261);
nand NAND2 (N14764, N14760, N2503);
or OR3 (N14765, N14761, N12402, N474);
and AND3 (N14766, N14763, N7376, N10200);
buf BUF1 (N14767, N14765);
xor XOR2 (N14768, N14752, N9663);
and AND2 (N14769, N14754, N5069);
xor XOR2 (N14770, N14755, N11556);
nand NAND4 (N14771, N14762, N1912, N5812, N163);
xor XOR2 (N14772, N14770, N13920);
or OR3 (N14773, N14767, N2742, N11856);
and AND4 (N14774, N14749, N4608, N3204, N10766);
buf BUF1 (N14775, N14769);
and AND3 (N14776, N14753, N7625, N11804);
nand NAND2 (N14777, N14776, N8320);
and AND4 (N14778, N14766, N8935, N12224, N7588);
buf BUF1 (N14779, N14772);
nor NOR4 (N14780, N14775, N12603, N5871, N5957);
or OR3 (N14781, N14764, N12103, N4978);
or OR2 (N14782, N14779, N483);
not NOT1 (N14783, N14777);
nor NOR2 (N14784, N14781, N11070);
not NOT1 (N14785, N14774);
nor NOR3 (N14786, N14771, N7447, N13101);
nor NOR4 (N14787, N14773, N14040, N6714, N11219);
and AND4 (N14788, N14787, N4207, N10364, N7113);
nand NAND4 (N14789, N14780, N4939, N12949, N13508);
or OR3 (N14790, N14782, N8199, N9035);
nand NAND3 (N14791, N14768, N3004, N7263);
nand NAND3 (N14792, N14790, N12373, N9455);
buf BUF1 (N14793, N14788);
buf BUF1 (N14794, N14786);
and AND2 (N14795, N14759, N11376);
nor NOR4 (N14796, N14783, N2229, N12060, N9617);
buf BUF1 (N14797, N14792);
and AND4 (N14798, N14784, N14763, N8560, N10418);
nand NAND3 (N14799, N14778, N10585, N12552);
nand NAND4 (N14800, N14799, N9768, N5151, N313);
nand NAND3 (N14801, N14789, N5393, N3642);
nand NAND4 (N14802, N14796, N12925, N6946, N14203);
or OR4 (N14803, N14801, N3361, N13506, N684);
nor NOR2 (N14804, N14795, N7325);
buf BUF1 (N14805, N14800);
xor XOR2 (N14806, N14805, N7359);
nor NOR3 (N14807, N14794, N11639, N10013);
buf BUF1 (N14808, N14791);
buf BUF1 (N14809, N14798);
xor XOR2 (N14810, N14793, N14673);
nor NOR2 (N14811, N14803, N2100);
nor NOR4 (N14812, N14811, N7494, N5451, N5696);
and AND4 (N14813, N14809, N13602, N7160, N76);
nand NAND4 (N14814, N14810, N10459, N11904, N1200);
xor XOR2 (N14815, N14813, N8304);
nand NAND3 (N14816, N14807, N6820, N4264);
not NOT1 (N14817, N14815);
buf BUF1 (N14818, N14802);
nand NAND2 (N14819, N14797, N168);
not NOT1 (N14820, N14812);
not NOT1 (N14821, N14808);
xor XOR2 (N14822, N14821, N10749);
nand NAND4 (N14823, N14814, N13953, N731, N9952);
buf BUF1 (N14824, N14823);
buf BUF1 (N14825, N14824);
nor NOR4 (N14826, N14785, N3816, N12332, N12801);
not NOT1 (N14827, N14826);
and AND4 (N14828, N14818, N5157, N5819, N12193);
nand NAND4 (N14829, N14822, N795, N10249, N14438);
and AND2 (N14830, N14804, N690);
xor XOR2 (N14831, N14820, N1809);
and AND4 (N14832, N14819, N640, N13991, N2047);
buf BUF1 (N14833, N14817);
and AND2 (N14834, N14831, N11192);
nor NOR3 (N14835, N14832, N8766, N10232);
buf BUF1 (N14836, N14806);
or OR4 (N14837, N14834, N12750, N105, N8444);
or OR2 (N14838, N14829, N3915);
buf BUF1 (N14839, N14830);
nand NAND3 (N14840, N14835, N10027, N9627);
buf BUF1 (N14841, N14825);
not NOT1 (N14842, N14841);
buf BUF1 (N14843, N14837);
xor XOR2 (N14844, N14840, N7645);
and AND4 (N14845, N14827, N1516, N13149, N5282);
nand NAND2 (N14846, N14836, N14474);
xor XOR2 (N14847, N14838, N13675);
and AND2 (N14848, N14828, N13856);
nor NOR2 (N14849, N14846, N5785);
not NOT1 (N14850, N14847);
and AND4 (N14851, N14833, N2580, N13544, N11236);
nor NOR4 (N14852, N14839, N2749, N13220, N2278);
nand NAND4 (N14853, N14851, N6656, N8920, N10564);
buf BUF1 (N14854, N14842);
buf BUF1 (N14855, N14852);
and AND3 (N14856, N14849, N6059, N7532);
not NOT1 (N14857, N14853);
xor XOR2 (N14858, N14845, N6062);
nor NOR2 (N14859, N14857, N14405);
or OR3 (N14860, N14816, N12193, N6310);
nor NOR4 (N14861, N14848, N157, N7133, N13531);
nor NOR2 (N14862, N14855, N3815);
xor XOR2 (N14863, N14856, N5549);
xor XOR2 (N14864, N14861, N14512);
and AND3 (N14865, N14858, N946, N3283);
xor XOR2 (N14866, N14862, N9187);
and AND2 (N14867, N14859, N53);
nand NAND4 (N14868, N14844, N2468, N12423, N9784);
not NOT1 (N14869, N14867);
and AND2 (N14870, N14860, N5825);
nand NAND2 (N14871, N14864, N8103);
not NOT1 (N14872, N14854);
nand NAND2 (N14873, N14863, N9413);
not NOT1 (N14874, N14843);
or OR4 (N14875, N14874, N10166, N6578, N2548);
not NOT1 (N14876, N14875);
or OR3 (N14877, N14873, N6028, N14110);
or OR3 (N14878, N14877, N2649, N4879);
nor NOR2 (N14879, N14876, N10637);
xor XOR2 (N14880, N14865, N1676);
nand NAND3 (N14881, N14850, N14593, N1966);
nand NAND2 (N14882, N14869, N6025);
nand NAND2 (N14883, N14870, N11494);
nor NOR3 (N14884, N14879, N6118, N14648);
xor XOR2 (N14885, N14884, N10483);
xor XOR2 (N14886, N14872, N6896);
or OR4 (N14887, N14881, N8093, N14406, N10418);
or OR2 (N14888, N14883, N10057);
xor XOR2 (N14889, N14887, N9053);
xor XOR2 (N14890, N14880, N10512);
nand NAND4 (N14891, N14871, N12916, N14725, N1946);
or OR2 (N14892, N14868, N11430);
or OR3 (N14893, N14892, N389, N256);
not NOT1 (N14894, N14882);
nand NAND2 (N14895, N14886, N10331);
xor XOR2 (N14896, N14893, N6592);
and AND3 (N14897, N14889, N1114, N4722);
nor NOR3 (N14898, N14895, N4664, N5201);
or OR4 (N14899, N14866, N6943, N6262, N9650);
buf BUF1 (N14900, N14894);
not NOT1 (N14901, N14878);
nand NAND4 (N14902, N14899, N9867, N1864, N3304);
or OR3 (N14903, N14891, N489, N13666);
buf BUF1 (N14904, N14890);
and AND4 (N14905, N14898, N3500, N5914, N7160);
xor XOR2 (N14906, N14888, N14728);
not NOT1 (N14907, N14896);
nand NAND2 (N14908, N14904, N7893);
xor XOR2 (N14909, N14901, N4083);
nor NOR2 (N14910, N14900, N8108);
and AND3 (N14911, N14907, N8510, N13845);
xor XOR2 (N14912, N14906, N3357);
nor NOR3 (N14913, N14885, N8184, N630);
nand NAND3 (N14914, N14912, N1580, N14706);
and AND3 (N14915, N14908, N3984, N2);
or OR3 (N14916, N14913, N11475, N3526);
nand NAND3 (N14917, N14909, N8451, N1934);
nand NAND2 (N14918, N14917, N14164);
or OR4 (N14919, N14918, N3979, N12195, N14694);
and AND4 (N14920, N14914, N14485, N14383, N11193);
nor NOR4 (N14921, N14902, N5121, N12372, N1813);
or OR3 (N14922, N14905, N12582, N9878);
nand NAND4 (N14923, N14921, N13897, N4995, N2009);
and AND4 (N14924, N14920, N9825, N3826, N8016);
nor NOR4 (N14925, N14915, N10165, N11041, N7663);
nand NAND4 (N14926, N14910, N5775, N14119, N2956);
nor NOR3 (N14927, N14923, N7817, N14570);
not NOT1 (N14928, N14903);
nor NOR3 (N14929, N14922, N2220, N9272);
or OR3 (N14930, N14897, N8819, N1094);
nor NOR4 (N14931, N14919, N8177, N14444, N6498);
nor NOR4 (N14932, N14931, N9105, N7943, N995);
not NOT1 (N14933, N14924);
xor XOR2 (N14934, N14930, N9842);
nand NAND4 (N14935, N14926, N2831, N12550, N8369);
xor XOR2 (N14936, N14911, N10614);
not NOT1 (N14937, N14932);
xor XOR2 (N14938, N14937, N13546);
not NOT1 (N14939, N14935);
and AND3 (N14940, N14939, N12304, N3861);
and AND4 (N14941, N14936, N1990, N5129, N7654);
not NOT1 (N14942, N14916);
or OR2 (N14943, N14929, N14513);
nor NOR4 (N14944, N14927, N1192, N14419, N9310);
and AND3 (N14945, N14942, N4047, N13772);
nor NOR2 (N14946, N14938, N13359);
nor NOR2 (N14947, N14946, N342);
or OR4 (N14948, N14944, N3197, N13520, N3877);
or OR4 (N14949, N14928, N14587, N1142, N3733);
xor XOR2 (N14950, N14934, N960);
and AND2 (N14951, N14925, N8575);
not NOT1 (N14952, N14949);
or OR3 (N14953, N14950, N10615, N14797);
nor NOR2 (N14954, N14948, N14030);
and AND4 (N14955, N14951, N576, N4305, N12237);
buf BUF1 (N14956, N14943);
and AND4 (N14957, N14947, N1734, N2735, N4810);
or OR4 (N14958, N14957, N3116, N8765, N13052);
and AND3 (N14959, N14945, N11163, N14288);
xor XOR2 (N14960, N14953, N9185);
nor NOR3 (N14961, N14952, N12203, N12384);
xor XOR2 (N14962, N14955, N12337);
not NOT1 (N14963, N14956);
and AND3 (N14964, N14954, N5351, N6381);
or OR2 (N14965, N14958, N2418);
nor NOR4 (N14966, N14959, N8658, N510, N1830);
not NOT1 (N14967, N14933);
nor NOR4 (N14968, N14962, N11526, N12364, N9033);
not NOT1 (N14969, N14966);
nand NAND4 (N14970, N14968, N14204, N12917, N12731);
nor NOR2 (N14971, N14963, N3716);
not NOT1 (N14972, N14969);
or OR3 (N14973, N14967, N9141, N7500);
not NOT1 (N14974, N14941);
buf BUF1 (N14975, N14965);
nand NAND4 (N14976, N14971, N256, N13179, N5482);
xor XOR2 (N14977, N14974, N11920);
or OR4 (N14978, N14970, N9244, N14807, N14738);
not NOT1 (N14979, N14964);
nand NAND2 (N14980, N14973, N12825);
and AND4 (N14981, N14960, N7631, N6596, N7982);
or OR2 (N14982, N14972, N12814);
buf BUF1 (N14983, N14961);
buf BUF1 (N14984, N14981);
xor XOR2 (N14985, N14980, N1938);
nand NAND4 (N14986, N14983, N2381, N11609, N7961);
nand NAND3 (N14987, N14979, N4832, N11592);
nand NAND3 (N14988, N14986, N3377, N6211);
or OR4 (N14989, N14978, N14641, N1652, N2898);
nor NOR3 (N14990, N14940, N6117, N11778);
not NOT1 (N14991, N14977);
or OR4 (N14992, N14989, N14112, N12973, N13235);
buf BUF1 (N14993, N14976);
or OR4 (N14994, N14993, N2953, N5593, N10456);
or OR3 (N14995, N14990, N9277, N13601);
nand NAND3 (N14996, N14984, N8593, N14779);
or OR2 (N14997, N14994, N6978);
nand NAND2 (N14998, N14995, N1852);
not NOT1 (N14999, N14982);
xor XOR2 (N15000, N14992, N11126);
or OR3 (N15001, N14998, N5189, N2973);
buf BUF1 (N15002, N14985);
buf BUF1 (N15003, N14975);
buf BUF1 (N15004, N14997);
nor NOR3 (N15005, N15002, N11659, N3945);
and AND2 (N15006, N14991, N9855);
and AND4 (N15007, N14996, N3379, N8590, N3401);
nor NOR4 (N15008, N15001, N4353, N4633, N9452);
buf BUF1 (N15009, N15003);
nand NAND4 (N15010, N15008, N3532, N4504, N4023);
or OR3 (N15011, N15000, N14767, N7611);
buf BUF1 (N15012, N14999);
xor XOR2 (N15013, N15006, N4952);
or OR2 (N15014, N15012, N8963);
or OR4 (N15015, N15004, N10271, N12995, N5718);
and AND3 (N15016, N15011, N12131, N2634);
nor NOR4 (N15017, N15013, N13808, N11913, N12515);
or OR4 (N15018, N15009, N11697, N14148, N765);
and AND4 (N15019, N15015, N4126, N10596, N5367);
or OR4 (N15020, N15017, N3049, N1267, N857);
xor XOR2 (N15021, N15010, N2259);
buf BUF1 (N15022, N15018);
and AND4 (N15023, N15007, N10397, N596, N11261);
nand NAND3 (N15024, N15023, N8794, N9166);
or OR4 (N15025, N15021, N2679, N8689, N8871);
nor NOR2 (N15026, N15014, N3690);
buf BUF1 (N15027, N15020);
xor XOR2 (N15028, N15022, N7755);
or OR4 (N15029, N15027, N11228, N2716, N2208);
nor NOR4 (N15030, N15016, N6425, N698, N10031);
buf BUF1 (N15031, N15024);
nor NOR4 (N15032, N15025, N2809, N13595, N8560);
nor NOR2 (N15033, N15030, N6853);
not NOT1 (N15034, N15005);
nor NOR4 (N15035, N15033, N14532, N4609, N1466);
xor XOR2 (N15036, N15026, N5050);
not NOT1 (N15037, N15035);
nand NAND2 (N15038, N14988, N10398);
and AND3 (N15039, N15031, N13064, N4472);
nor NOR3 (N15040, N15029, N9213, N7966);
not NOT1 (N15041, N15036);
or OR3 (N15042, N15041, N1075, N5923);
and AND4 (N15043, N15019, N13663, N10389, N6368);
and AND2 (N15044, N15038, N6108);
and AND4 (N15045, N14987, N1962, N1077, N1667);
nand NAND4 (N15046, N15042, N13924, N12833, N11240);
xor XOR2 (N15047, N15039, N11332);
and AND2 (N15048, N15034, N2932);
xor XOR2 (N15049, N15032, N13070);
xor XOR2 (N15050, N15046, N4202);
xor XOR2 (N15051, N15040, N14936);
nand NAND2 (N15052, N15048, N11922);
xor XOR2 (N15053, N15047, N11804);
not NOT1 (N15054, N15049);
nor NOR4 (N15055, N15052, N6976, N896, N993);
xor XOR2 (N15056, N15043, N7112);
or OR3 (N15057, N15055, N564, N4383);
nor NOR3 (N15058, N15051, N14687, N10614);
or OR2 (N15059, N15028, N10130);
not NOT1 (N15060, N15053);
nand NAND2 (N15061, N15054, N3530);
or OR2 (N15062, N15037, N6601);
nor NOR2 (N15063, N15056, N27);
buf BUF1 (N15064, N15059);
nor NOR4 (N15065, N15058, N202, N471, N12931);
and AND2 (N15066, N15060, N4295);
nand NAND3 (N15067, N15065, N10349, N1987);
nor NOR3 (N15068, N15057, N14417, N14921);
and AND2 (N15069, N15067, N13782);
nor NOR2 (N15070, N15068, N15041);
and AND3 (N15071, N15044, N3043, N11522);
or OR2 (N15072, N15071, N4739);
buf BUF1 (N15073, N15070);
nand NAND4 (N15074, N15061, N7472, N3410, N8732);
and AND2 (N15075, N15050, N14257);
nand NAND4 (N15076, N15066, N12944, N2672, N553);
and AND2 (N15077, N15076, N7132);
buf BUF1 (N15078, N15069);
or OR4 (N15079, N15077, N6769, N10714, N8834);
or OR3 (N15080, N15063, N14399, N7910);
nand NAND3 (N15081, N15075, N13464, N1503);
nand NAND3 (N15082, N15080, N13167, N1047);
nand NAND4 (N15083, N15074, N1901, N294, N1478);
and AND2 (N15084, N15072, N1263);
and AND4 (N15085, N15073, N3964, N11003, N11566);
not NOT1 (N15086, N15085);
or OR3 (N15087, N15081, N7160, N8309);
nand NAND3 (N15088, N15086, N2379, N1132);
xor XOR2 (N15089, N15062, N11730);
or OR3 (N15090, N15089, N6289, N5853);
xor XOR2 (N15091, N15088, N12295);
nor NOR2 (N15092, N15078, N4644);
nor NOR3 (N15093, N15083, N10771, N7676);
and AND2 (N15094, N15093, N2532);
and AND3 (N15095, N15064, N9587, N3467);
or OR2 (N15096, N15087, N4363);
nor NOR3 (N15097, N15084, N1991, N9314);
or OR2 (N15098, N15096, N8126);
not NOT1 (N15099, N15045);
and AND3 (N15100, N15097, N9544, N13544);
xor XOR2 (N15101, N15099, N1269);
and AND4 (N15102, N15095, N7073, N8598, N7115);
and AND2 (N15103, N15102, N14767);
nand NAND4 (N15104, N15079, N10895, N6566, N13577);
nand NAND4 (N15105, N15092, N965, N9278, N7250);
nor NOR3 (N15106, N15104, N9249, N1853);
or OR3 (N15107, N15098, N9112, N5966);
and AND4 (N15108, N15105, N289, N13032, N6363);
buf BUF1 (N15109, N15082);
and AND4 (N15110, N15103, N8874, N1593, N13913);
buf BUF1 (N15111, N15110);
not NOT1 (N15112, N15109);
not NOT1 (N15113, N15106);
not NOT1 (N15114, N15101);
and AND4 (N15115, N15112, N7524, N1953, N5209);
buf BUF1 (N15116, N15113);
nor NOR2 (N15117, N15111, N12926);
buf BUF1 (N15118, N15094);
not NOT1 (N15119, N15108);
nor NOR4 (N15120, N15090, N5748, N13507, N4298);
buf BUF1 (N15121, N15091);
xor XOR2 (N15122, N15114, N8675);
buf BUF1 (N15123, N15119);
nand NAND4 (N15124, N15116, N13215, N6384, N1480);
and AND2 (N15125, N15122, N527);
nor NOR4 (N15126, N15107, N10666, N13000, N7898);
buf BUF1 (N15127, N15123);
buf BUF1 (N15128, N15118);
nor NOR3 (N15129, N15115, N11578, N12380);
not NOT1 (N15130, N15128);
or OR4 (N15131, N15125, N10968, N1932, N13920);
nor NOR3 (N15132, N15126, N8595, N12629);
nor NOR4 (N15133, N15121, N9126, N3370, N14920);
nand NAND4 (N15134, N15133, N3012, N6347, N5728);
xor XOR2 (N15135, N15132, N2175);
xor XOR2 (N15136, N15134, N1639);
nor NOR3 (N15137, N15117, N6850, N2649);
xor XOR2 (N15138, N15131, N3714);
not NOT1 (N15139, N15120);
xor XOR2 (N15140, N15100, N10573);
nand NAND3 (N15141, N15127, N6610, N13083);
buf BUF1 (N15142, N15129);
xor XOR2 (N15143, N15139, N12990);
or OR2 (N15144, N15137, N12894);
or OR4 (N15145, N15130, N14602, N6706, N4887);
nand NAND4 (N15146, N15124, N2887, N1042, N3129);
not NOT1 (N15147, N15141);
not NOT1 (N15148, N15140);
nor NOR4 (N15149, N15142, N11422, N5263, N4975);
and AND4 (N15150, N15143, N12816, N5528, N7520);
or OR3 (N15151, N15138, N13627, N1105);
xor XOR2 (N15152, N15135, N11859);
or OR4 (N15153, N15136, N2180, N14418, N4594);
nand NAND3 (N15154, N15144, N12088, N2111);
buf BUF1 (N15155, N15150);
and AND4 (N15156, N15152, N10686, N14172, N12154);
or OR3 (N15157, N15148, N145, N14882);
nand NAND2 (N15158, N15149, N1109);
buf BUF1 (N15159, N15147);
and AND4 (N15160, N15158, N12676, N9667, N10377);
buf BUF1 (N15161, N15151);
or OR4 (N15162, N15156, N2835, N2248, N891);
or OR4 (N15163, N15157, N13113, N1130, N87);
and AND4 (N15164, N15159, N841, N8810, N3877);
buf BUF1 (N15165, N15163);
not NOT1 (N15166, N15155);
nor NOR2 (N15167, N15153, N10239);
and AND2 (N15168, N15160, N3738);
or OR2 (N15169, N15145, N5154);
xor XOR2 (N15170, N15167, N2770);
buf BUF1 (N15171, N15164);
nor NOR3 (N15172, N15171, N15071, N12213);
buf BUF1 (N15173, N15169);
nand NAND3 (N15174, N15172, N11239, N4975);
not NOT1 (N15175, N15146);
or OR3 (N15176, N15161, N3336, N13415);
xor XOR2 (N15177, N15176, N14046);
buf BUF1 (N15178, N15174);
and AND4 (N15179, N15166, N6147, N12320, N14201);
not NOT1 (N15180, N15175);
buf BUF1 (N15181, N15178);
nand NAND3 (N15182, N15173, N3517, N14317);
or OR2 (N15183, N15182, N10152);
and AND3 (N15184, N15181, N12358, N5141);
not NOT1 (N15185, N15183);
nor NOR2 (N15186, N15154, N683);
nand NAND3 (N15187, N15165, N10543, N15012);
and AND3 (N15188, N15162, N7112, N12884);
nand NAND4 (N15189, N15188, N5330, N2842, N4549);
nor NOR4 (N15190, N15179, N12431, N2881, N12075);
nand NAND2 (N15191, N15170, N137);
buf BUF1 (N15192, N15189);
and AND2 (N15193, N15184, N12500);
and AND4 (N15194, N15193, N10550, N13605, N950);
and AND4 (N15195, N15191, N4391, N7308, N1707);
xor XOR2 (N15196, N15195, N2707);
nor NOR2 (N15197, N15177, N11468);
buf BUF1 (N15198, N15196);
xor XOR2 (N15199, N15198, N6448);
xor XOR2 (N15200, N15197, N2842);
nand NAND3 (N15201, N15190, N498, N9239);
nor NOR3 (N15202, N15168, N7747, N13316);
nor NOR3 (N15203, N15202, N14946, N87);
not NOT1 (N15204, N15200);
or OR3 (N15205, N15194, N6447, N3143);
nor NOR2 (N15206, N15201, N14576);
nor NOR3 (N15207, N15206, N920, N7940);
xor XOR2 (N15208, N15180, N5857);
nor NOR4 (N15209, N15185, N1742, N12531, N8681);
not NOT1 (N15210, N15203);
nand NAND2 (N15211, N15209, N13283);
and AND2 (N15212, N15207, N3079);
nor NOR2 (N15213, N15205, N14598);
and AND3 (N15214, N15210, N8594, N1174);
buf BUF1 (N15215, N15208);
or OR2 (N15216, N15211, N7780);
and AND3 (N15217, N15216, N12771, N3528);
nand NAND4 (N15218, N15217, N2403, N9948, N6597);
not NOT1 (N15219, N15199);
or OR3 (N15220, N15212, N4750, N241);
nor NOR3 (N15221, N15215, N394, N1217);
nor NOR4 (N15222, N15219, N8761, N4000, N1453);
or OR4 (N15223, N15221, N14531, N11768, N11577);
or OR3 (N15224, N15192, N4792, N11518);
nand NAND3 (N15225, N15218, N11938, N10378);
nor NOR2 (N15226, N15223, N7447);
nand NAND3 (N15227, N15186, N14501, N108);
buf BUF1 (N15228, N15225);
not NOT1 (N15229, N15226);
nand NAND3 (N15230, N15224, N3385, N1915);
or OR3 (N15231, N15229, N925, N7886);
nor NOR3 (N15232, N15204, N12300, N12097);
buf BUF1 (N15233, N15232);
xor XOR2 (N15234, N15228, N3267);
buf BUF1 (N15235, N15187);
nor NOR4 (N15236, N15227, N2874, N14238, N9329);
not NOT1 (N15237, N15213);
and AND3 (N15238, N15220, N7693, N2877);
and AND3 (N15239, N15233, N10455, N9086);
and AND4 (N15240, N15239, N9406, N11466, N8777);
nand NAND2 (N15241, N15214, N8701);
nand NAND3 (N15242, N15234, N10479, N11003);
and AND2 (N15243, N15222, N13475);
nor NOR3 (N15244, N15236, N8574, N10133);
and AND4 (N15245, N15238, N1232, N5599, N12139);
nor NOR2 (N15246, N15244, N2819);
xor XOR2 (N15247, N15243, N7341);
nor NOR3 (N15248, N15231, N3712, N7071);
xor XOR2 (N15249, N15241, N14311);
not NOT1 (N15250, N15237);
xor XOR2 (N15251, N15250, N13990);
not NOT1 (N15252, N15230);
nor NOR3 (N15253, N15251, N7149, N1265);
buf BUF1 (N15254, N15252);
nor NOR4 (N15255, N15246, N4626, N3372, N8828);
nand NAND4 (N15256, N15242, N5230, N6578, N1375);
nand NAND3 (N15257, N15254, N4762, N2211);
not NOT1 (N15258, N15255);
and AND2 (N15259, N15256, N1658);
nand NAND4 (N15260, N15258, N2696, N15046, N2450);
and AND2 (N15261, N15248, N13046);
nand NAND2 (N15262, N15249, N11392);
nor NOR4 (N15263, N15261, N11585, N7481, N2322);
buf BUF1 (N15264, N15253);
nand NAND4 (N15265, N15260, N13519, N4365, N11577);
and AND2 (N15266, N15245, N11112);
and AND3 (N15267, N15263, N1585, N3300);
or OR2 (N15268, N15267, N3642);
and AND3 (N15269, N15259, N11140, N7711);
not NOT1 (N15270, N15257);
and AND2 (N15271, N15240, N4850);
or OR4 (N15272, N15269, N11139, N4464, N495);
nor NOR4 (N15273, N15272, N12639, N14728, N5833);
and AND4 (N15274, N15271, N4776, N6795, N1260);
buf BUF1 (N15275, N15268);
not NOT1 (N15276, N15265);
or OR4 (N15277, N15262, N7107, N15008, N14386);
and AND3 (N15278, N15274, N14980, N3833);
buf BUF1 (N15279, N15275);
nor NOR4 (N15280, N15278, N7203, N13241, N11770);
or OR4 (N15281, N15276, N8407, N12386, N10059);
buf BUF1 (N15282, N15277);
or OR2 (N15283, N15279, N3656);
nand NAND3 (N15284, N15283, N14273, N11048);
buf BUF1 (N15285, N15264);
or OR4 (N15286, N15282, N4537, N10833, N14800);
and AND2 (N15287, N15266, N14419);
or OR2 (N15288, N15270, N13473);
nor NOR3 (N15289, N15247, N14200, N8867);
not NOT1 (N15290, N15273);
not NOT1 (N15291, N15287);
not NOT1 (N15292, N15290);
nor NOR2 (N15293, N15285, N11805);
nor NOR3 (N15294, N15293, N4925, N13639);
nand NAND4 (N15295, N15281, N4849, N13187, N14212);
or OR3 (N15296, N15288, N8031, N12797);
nor NOR2 (N15297, N15286, N2179);
buf BUF1 (N15298, N15297);
not NOT1 (N15299, N15295);
not NOT1 (N15300, N15296);
xor XOR2 (N15301, N15298, N2876);
nor NOR2 (N15302, N15294, N9210);
buf BUF1 (N15303, N15289);
nand NAND3 (N15304, N15291, N2345, N4776);
xor XOR2 (N15305, N15280, N4900);
buf BUF1 (N15306, N15305);
nand NAND4 (N15307, N15301, N6240, N4074, N10941);
nand NAND3 (N15308, N15300, N5494, N1726);
xor XOR2 (N15309, N15304, N6268);
nor NOR3 (N15310, N15284, N8002, N1047);
or OR2 (N15311, N15235, N7176);
nand NAND4 (N15312, N15311, N14807, N5616, N6748);
not NOT1 (N15313, N15303);
nand NAND4 (N15314, N15312, N10170, N3248, N15253);
nor NOR4 (N15315, N15308, N2458, N11574, N13886);
not NOT1 (N15316, N15292);
or OR2 (N15317, N15315, N1099);
not NOT1 (N15318, N15309);
buf BUF1 (N15319, N15318);
nand NAND3 (N15320, N15313, N13899, N1340);
nor NOR4 (N15321, N15302, N4282, N214, N9857);
or OR3 (N15322, N15317, N14044, N1005);
and AND2 (N15323, N15320, N7981);
or OR4 (N15324, N15299, N1934, N4581, N7832);
xor XOR2 (N15325, N15322, N8793);
nand NAND3 (N15326, N15325, N2164, N2629);
nand NAND3 (N15327, N15310, N11059, N4387);
xor XOR2 (N15328, N15307, N7834);
not NOT1 (N15329, N15323);
nand NAND3 (N15330, N15314, N3858, N5039);
or OR4 (N15331, N15316, N3311, N3723, N7920);
or OR2 (N15332, N15321, N13201);
not NOT1 (N15333, N15324);
buf BUF1 (N15334, N15326);
nand NAND2 (N15335, N15328, N10146);
nor NOR3 (N15336, N15332, N13086, N9190);
and AND2 (N15337, N15336, N7632);
buf BUF1 (N15338, N15337);
or OR2 (N15339, N15327, N6275);
or OR4 (N15340, N15306, N14018, N8360, N8250);
nor NOR3 (N15341, N15331, N2015, N7837);
not NOT1 (N15342, N15339);
or OR3 (N15343, N15334, N1222, N10525);
not NOT1 (N15344, N15330);
and AND3 (N15345, N15341, N5447, N12463);
buf BUF1 (N15346, N15319);
nand NAND3 (N15347, N15346, N12533, N6042);
xor XOR2 (N15348, N15333, N5468);
or OR4 (N15349, N15338, N6546, N6715, N1674);
nand NAND4 (N15350, N15348, N2722, N10201, N4538);
nor NOR2 (N15351, N15342, N6452);
not NOT1 (N15352, N15347);
nor NOR2 (N15353, N15340, N4717);
not NOT1 (N15354, N15349);
buf BUF1 (N15355, N15329);
and AND3 (N15356, N15335, N3829, N4333);
nand NAND2 (N15357, N15355, N8939);
nor NOR4 (N15358, N15352, N6410, N14040, N4012);
not NOT1 (N15359, N15357);
or OR4 (N15360, N15345, N3052, N6244, N12475);
not NOT1 (N15361, N15360);
or OR3 (N15362, N15344, N11613, N11918);
xor XOR2 (N15363, N15356, N11298);
xor XOR2 (N15364, N15343, N2366);
or OR3 (N15365, N15350, N2350, N1433);
nand NAND4 (N15366, N15358, N12709, N9287, N424);
not NOT1 (N15367, N15353);
nand NAND2 (N15368, N15364, N3149);
not NOT1 (N15369, N15351);
and AND4 (N15370, N15367, N8535, N10576, N11016);
or OR3 (N15371, N15361, N7925, N9009);
and AND2 (N15372, N15370, N12573);
and AND3 (N15373, N15359, N1385, N1213);
and AND3 (N15374, N15354, N4201, N7642);
xor XOR2 (N15375, N15372, N601);
buf BUF1 (N15376, N15363);
nand NAND3 (N15377, N15366, N9899, N3437);
and AND4 (N15378, N15375, N12979, N9624, N4886);
not NOT1 (N15379, N15362);
and AND3 (N15380, N15368, N3169, N7254);
buf BUF1 (N15381, N15371);
and AND4 (N15382, N15369, N11687, N13479, N2828);
xor XOR2 (N15383, N15373, N11319);
nor NOR3 (N15384, N15379, N9278, N7982);
nor NOR4 (N15385, N15377, N12024, N5673, N11704);
nor NOR3 (N15386, N15385, N7826, N4915);
not NOT1 (N15387, N15384);
buf BUF1 (N15388, N15365);
nand NAND4 (N15389, N15382, N4036, N665, N11553);
not NOT1 (N15390, N15388);
buf BUF1 (N15391, N15390);
nor NOR3 (N15392, N15383, N1353, N2191);
nand NAND3 (N15393, N15389, N9174, N12839);
not NOT1 (N15394, N15386);
not NOT1 (N15395, N15393);
and AND2 (N15396, N15378, N2881);
and AND3 (N15397, N15392, N12741, N5376);
nand NAND2 (N15398, N15380, N12507);
or OR3 (N15399, N15374, N12430, N3079);
buf BUF1 (N15400, N15399);
or OR4 (N15401, N15398, N5483, N15048, N1305);
nand NAND3 (N15402, N15394, N2758, N1165);
or OR2 (N15403, N15397, N14817);
and AND2 (N15404, N15395, N2322);
buf BUF1 (N15405, N15402);
not NOT1 (N15406, N15404);
buf BUF1 (N15407, N15406);
not NOT1 (N15408, N15387);
nor NOR3 (N15409, N15401, N11491, N4068);
xor XOR2 (N15410, N15408, N6307);
not NOT1 (N15411, N15400);
xor XOR2 (N15412, N15405, N3826);
nor NOR4 (N15413, N15376, N4610, N911, N4034);
nor NOR4 (N15414, N15412, N3904, N4620, N5129);
not NOT1 (N15415, N15413);
nor NOR2 (N15416, N15415, N2624);
nand NAND3 (N15417, N15416, N12415, N3513);
nor NOR3 (N15418, N15410, N6848, N4146);
buf BUF1 (N15419, N15381);
nand NAND3 (N15420, N15419, N1371, N2507);
or OR4 (N15421, N15407, N15153, N11087, N8866);
buf BUF1 (N15422, N15403);
not NOT1 (N15423, N15418);
nor NOR3 (N15424, N15422, N9033, N13870);
or OR4 (N15425, N15424, N7252, N3610, N320);
and AND3 (N15426, N15414, N9156, N14778);
and AND2 (N15427, N15409, N3148);
not NOT1 (N15428, N15391);
or OR3 (N15429, N15396, N2284, N9873);
nor NOR2 (N15430, N15428, N14751);
xor XOR2 (N15431, N15421, N5723);
not NOT1 (N15432, N15425);
not NOT1 (N15433, N15411);
not NOT1 (N15434, N15420);
or OR2 (N15435, N15431, N13940);
buf BUF1 (N15436, N15430);
not NOT1 (N15437, N15426);
buf BUF1 (N15438, N15434);
nand NAND2 (N15439, N15438, N14627);
xor XOR2 (N15440, N15436, N9181);
not NOT1 (N15441, N15429);
nand NAND4 (N15442, N15423, N13665, N9135, N7037);
buf BUF1 (N15443, N15417);
nand NAND4 (N15444, N15441, N14623, N614, N13532);
buf BUF1 (N15445, N15432);
buf BUF1 (N15446, N15445);
xor XOR2 (N15447, N15427, N1801);
not NOT1 (N15448, N15440);
not NOT1 (N15449, N15437);
and AND2 (N15450, N15447, N3304);
and AND4 (N15451, N15443, N13067, N9219, N5239);
xor XOR2 (N15452, N15439, N5608);
nor NOR3 (N15453, N15450, N1058, N2411);
nor NOR2 (N15454, N15452, N12704);
not NOT1 (N15455, N15435);
nor NOR4 (N15456, N15448, N7611, N12665, N9213);
nand NAND2 (N15457, N15456, N5089);
or OR4 (N15458, N15457, N5226, N6849, N4173);
and AND4 (N15459, N15433, N3437, N13299, N5019);
or OR2 (N15460, N15446, N6713);
or OR3 (N15461, N15460, N10052, N5202);
buf BUF1 (N15462, N15458);
and AND4 (N15463, N15454, N3897, N8595, N5755);
buf BUF1 (N15464, N15451);
not NOT1 (N15465, N15461);
and AND2 (N15466, N15455, N3628);
nor NOR2 (N15467, N15465, N2674);
nand NAND4 (N15468, N15466, N14193, N3184, N10859);
buf BUF1 (N15469, N15453);
or OR2 (N15470, N15442, N9641);
not NOT1 (N15471, N15464);
or OR4 (N15472, N15459, N301, N11375, N10983);
nor NOR3 (N15473, N15468, N73, N14593);
nand NAND3 (N15474, N15473, N10059, N2283);
and AND4 (N15475, N15474, N14249, N7397, N4973);
buf BUF1 (N15476, N15469);
nand NAND4 (N15477, N15472, N1028, N6995, N15153);
nand NAND3 (N15478, N15477, N941, N13417);
and AND4 (N15479, N15462, N14673, N9046, N901);
not NOT1 (N15480, N15444);
xor XOR2 (N15481, N15480, N1976);
not NOT1 (N15482, N15475);
nand NAND2 (N15483, N15463, N11252);
and AND2 (N15484, N15478, N7629);
not NOT1 (N15485, N15476);
xor XOR2 (N15486, N15483, N13273);
buf BUF1 (N15487, N15481);
or OR4 (N15488, N15449, N10178, N716, N10561);
buf BUF1 (N15489, N15467);
buf BUF1 (N15490, N15487);
not NOT1 (N15491, N15489);
nor NOR2 (N15492, N15485, N12384);
nor NOR2 (N15493, N15471, N13613);
buf BUF1 (N15494, N15479);
and AND4 (N15495, N15491, N2365, N4976, N3174);
xor XOR2 (N15496, N15488, N4044);
and AND2 (N15497, N15496, N12251);
buf BUF1 (N15498, N15490);
not NOT1 (N15499, N15495);
and AND2 (N15500, N15493, N15485);
nand NAND2 (N15501, N15484, N8300);
nor NOR4 (N15502, N15486, N2942, N10554, N1656);
or OR4 (N15503, N15499, N15362, N9556, N1073);
or OR3 (N15504, N15502, N10781, N11056);
nor NOR3 (N15505, N15482, N13962, N12639);
nor NOR4 (N15506, N15505, N15448, N5872, N5671);
xor XOR2 (N15507, N15492, N3999);
and AND3 (N15508, N15498, N15244, N4628);
xor XOR2 (N15509, N15504, N11799);
or OR2 (N15510, N15501, N6609);
and AND3 (N15511, N15494, N15033, N1475);
buf BUF1 (N15512, N15503);
not NOT1 (N15513, N15507);
and AND3 (N15514, N15511, N6370, N13628);
nand NAND4 (N15515, N15508, N8391, N11249, N7572);
nand NAND2 (N15516, N15512, N12228);
or OR4 (N15517, N15497, N14453, N1150, N12442);
nand NAND2 (N15518, N15470, N5566);
buf BUF1 (N15519, N15500);
buf BUF1 (N15520, N15513);
or OR2 (N15521, N15506, N13098);
nor NOR4 (N15522, N15519, N3115, N11749, N10525);
or OR2 (N15523, N15520, N11980);
or OR4 (N15524, N15517, N9008, N10092, N11672);
and AND3 (N15525, N15522, N5265, N23);
nor NOR4 (N15526, N15525, N7917, N7567, N2106);
or OR2 (N15527, N15518, N2953);
nand NAND2 (N15528, N15514, N11990);
nor NOR2 (N15529, N15524, N4148);
nand NAND4 (N15530, N15526, N7287, N12394, N12932);
nand NAND3 (N15531, N15523, N10712, N15415);
not NOT1 (N15532, N15515);
xor XOR2 (N15533, N15528, N5089);
xor XOR2 (N15534, N15521, N6710);
or OR2 (N15535, N15510, N6114);
xor XOR2 (N15536, N15527, N940);
nor NOR3 (N15537, N15509, N3459, N5374);
nand NAND4 (N15538, N15529, N9779, N9032, N6107);
and AND4 (N15539, N15530, N5702, N15348, N10035);
and AND2 (N15540, N15538, N15390);
xor XOR2 (N15541, N15535, N8684);
or OR4 (N15542, N15532, N3672, N14775, N11221);
nor NOR4 (N15543, N15539, N10329, N14477, N522);
not NOT1 (N15544, N15543);
and AND3 (N15545, N15544, N10211, N10070);
and AND4 (N15546, N15516, N4351, N7980, N141);
buf BUF1 (N15547, N15537);
nand NAND2 (N15548, N15540, N7172);
and AND4 (N15549, N15531, N13183, N69, N12123);
xor XOR2 (N15550, N15541, N3648);
not NOT1 (N15551, N15545);
and AND3 (N15552, N15536, N1652, N1323);
xor XOR2 (N15553, N15534, N1846);
nor NOR4 (N15554, N15553, N913, N5990, N4463);
nand NAND2 (N15555, N15550, N309);
not NOT1 (N15556, N15549);
or OR3 (N15557, N15547, N11658, N12013);
xor XOR2 (N15558, N15548, N10325);
buf BUF1 (N15559, N15557);
nor NOR2 (N15560, N15542, N12046);
xor XOR2 (N15561, N15556, N4336);
or OR2 (N15562, N15561, N8742);
and AND4 (N15563, N15533, N12152, N5140, N12337);
and AND3 (N15564, N15562, N7294, N8336);
nor NOR3 (N15565, N15552, N7177, N9516);
buf BUF1 (N15566, N15555);
or OR2 (N15567, N15558, N387);
not NOT1 (N15568, N15565);
xor XOR2 (N15569, N15567, N15300);
not NOT1 (N15570, N15560);
and AND3 (N15571, N15568, N1545, N9805);
not NOT1 (N15572, N15566);
xor XOR2 (N15573, N15564, N812);
not NOT1 (N15574, N15571);
or OR4 (N15575, N15570, N12246, N8156, N10253);
and AND2 (N15576, N15554, N1368);
buf BUF1 (N15577, N15575);
nor NOR4 (N15578, N15572, N7344, N3908, N11676);
or OR4 (N15579, N15551, N14216, N12947, N5439);
not NOT1 (N15580, N15579);
not NOT1 (N15581, N15574);
buf BUF1 (N15582, N15573);
nand NAND2 (N15583, N15563, N3568);
buf BUF1 (N15584, N15580);
or OR3 (N15585, N15581, N10992, N13048);
nor NOR2 (N15586, N15582, N6556);
and AND3 (N15587, N15584, N1535, N9450);
buf BUF1 (N15588, N15576);
nor NOR3 (N15589, N15578, N10804, N15169);
nor NOR2 (N15590, N15587, N12730);
or OR2 (N15591, N15586, N14914);
or OR2 (N15592, N15559, N12442);
buf BUF1 (N15593, N15577);
buf BUF1 (N15594, N15583);
and AND4 (N15595, N15594, N12896, N785, N8910);
buf BUF1 (N15596, N15590);
or OR4 (N15597, N15589, N10177, N9512, N10193);
or OR4 (N15598, N15592, N6305, N10077, N6777);
nand NAND3 (N15599, N15593, N4391, N3090);
or OR2 (N15600, N15546, N9830);
and AND2 (N15601, N15588, N12758);
buf BUF1 (N15602, N15569);
or OR2 (N15603, N15598, N7016);
and AND2 (N15604, N15600, N12313);
and AND3 (N15605, N15595, N3023, N12892);
buf BUF1 (N15606, N15599);
and AND3 (N15607, N15591, N7329, N1945);
nand NAND2 (N15608, N15604, N6286);
or OR3 (N15609, N15596, N12347, N14175);
nor NOR3 (N15610, N15606, N13059, N8065);
buf BUF1 (N15611, N15602);
nor NOR2 (N15612, N15611, N14642);
buf BUF1 (N15613, N15603);
buf BUF1 (N15614, N15597);
or OR4 (N15615, N15610, N9475, N5810, N12655);
and AND3 (N15616, N15608, N10828, N6574);
not NOT1 (N15617, N15585);
nand NAND4 (N15618, N15616, N10942, N1662, N10803);
not NOT1 (N15619, N15612);
buf BUF1 (N15620, N15601);
nand NAND2 (N15621, N15618, N11808);
not NOT1 (N15622, N15614);
nor NOR2 (N15623, N15620, N3723);
nand NAND4 (N15624, N15622, N3843, N4417, N14574);
and AND4 (N15625, N15607, N12868, N11950, N9528);
or OR2 (N15626, N15613, N2326);
nor NOR4 (N15627, N15615, N10291, N4574, N13012);
nor NOR4 (N15628, N15605, N1396, N11523, N2787);
xor XOR2 (N15629, N15625, N9812);
xor XOR2 (N15630, N15619, N13427);
nor NOR3 (N15631, N15627, N13457, N6644);
nand NAND3 (N15632, N15628, N3443, N1431);
nand NAND4 (N15633, N15623, N228, N8680, N15558);
nor NOR2 (N15634, N15632, N3258);
nand NAND2 (N15635, N15626, N4818);
not NOT1 (N15636, N15634);
and AND2 (N15637, N15630, N4474);
nor NOR3 (N15638, N15609, N1777, N15116);
nand NAND4 (N15639, N15617, N5594, N13810, N10661);
and AND3 (N15640, N15635, N3988, N12872);
nand NAND4 (N15641, N15637, N12313, N10930, N8235);
not NOT1 (N15642, N15624);
not NOT1 (N15643, N15641);
and AND2 (N15644, N15643, N5200);
nor NOR4 (N15645, N15640, N5861, N6310, N2647);
xor XOR2 (N15646, N15644, N6233);
or OR2 (N15647, N15639, N1828);
nand NAND4 (N15648, N15636, N9653, N12010, N9855);
xor XOR2 (N15649, N15629, N7665);
buf BUF1 (N15650, N15633);
not NOT1 (N15651, N15649);
and AND4 (N15652, N15645, N4072, N6886, N10225);
xor XOR2 (N15653, N15651, N648);
nand NAND2 (N15654, N15652, N8131);
xor XOR2 (N15655, N15638, N13491);
nand NAND3 (N15656, N15655, N6724, N5988);
buf BUF1 (N15657, N15648);
xor XOR2 (N15658, N15654, N7770);
buf BUF1 (N15659, N15642);
xor XOR2 (N15660, N15647, N13480);
xor XOR2 (N15661, N15653, N1687);
or OR4 (N15662, N15659, N8421, N4335, N3314);
buf BUF1 (N15663, N15660);
not NOT1 (N15664, N15621);
and AND4 (N15665, N15664, N509, N7857, N6174);
nand NAND4 (N15666, N15662, N5703, N2838, N13899);
not NOT1 (N15667, N15663);
or OR2 (N15668, N15667, N2905);
nand NAND3 (N15669, N15661, N13276, N7278);
nor NOR2 (N15670, N15668, N1170);
and AND3 (N15671, N15646, N12261, N2784);
and AND4 (N15672, N15631, N3852, N15292, N4266);
xor XOR2 (N15673, N15658, N13534);
nor NOR3 (N15674, N15665, N2959, N15461);
and AND3 (N15675, N15672, N13519, N14679);
or OR4 (N15676, N15673, N2615, N2286, N5659);
buf BUF1 (N15677, N15676);
not NOT1 (N15678, N15656);
or OR3 (N15679, N15666, N1769, N11784);
not NOT1 (N15680, N15678);
nor NOR3 (N15681, N15650, N13540, N11706);
nor NOR2 (N15682, N15657, N9283);
buf BUF1 (N15683, N15675);
not NOT1 (N15684, N15671);
not NOT1 (N15685, N15677);
not NOT1 (N15686, N15679);
and AND3 (N15687, N15686, N845, N14684);
xor XOR2 (N15688, N15682, N195);
nand NAND4 (N15689, N15688, N1211, N1696, N747);
buf BUF1 (N15690, N15674);
nor NOR2 (N15691, N15687, N9143);
not NOT1 (N15692, N15680);
buf BUF1 (N15693, N15685);
nand NAND4 (N15694, N15684, N213, N12344, N6490);
nand NAND2 (N15695, N15683, N3297);
not NOT1 (N15696, N15669);
not NOT1 (N15697, N15693);
nand NAND3 (N15698, N15697, N4577, N3888);
xor XOR2 (N15699, N15681, N2965);
not NOT1 (N15700, N15689);
xor XOR2 (N15701, N15692, N10370);
xor XOR2 (N15702, N15701, N11628);
nand NAND2 (N15703, N15699, N11672);
nor NOR3 (N15704, N15690, N10109, N713);
nor NOR3 (N15705, N15704, N7079, N12003);
not NOT1 (N15706, N15696);
xor XOR2 (N15707, N15698, N9336);
not NOT1 (N15708, N15694);
and AND2 (N15709, N15708, N14911);
nor NOR4 (N15710, N15709, N14573, N3168, N8007);
nor NOR4 (N15711, N15707, N8260, N13344, N5196);
not NOT1 (N15712, N15711);
nand NAND3 (N15713, N15706, N7785, N14781);
not NOT1 (N15714, N15703);
not NOT1 (N15715, N15695);
not NOT1 (N15716, N15691);
buf BUF1 (N15717, N15670);
buf BUF1 (N15718, N15713);
not NOT1 (N15719, N15718);
nand NAND4 (N15720, N15717, N15655, N12300, N3523);
nand NAND2 (N15721, N15705, N3209);
and AND4 (N15722, N15714, N11445, N14028, N14926);
nand NAND3 (N15723, N15712, N4894, N958);
and AND4 (N15724, N15719, N10077, N13643, N3722);
nand NAND2 (N15725, N15716, N13419);
buf BUF1 (N15726, N15700);
xor XOR2 (N15727, N15723, N3885);
nand NAND4 (N15728, N15721, N6515, N8343, N8182);
not NOT1 (N15729, N15710);
nand NAND3 (N15730, N15727, N15340, N4183);
nor NOR4 (N15731, N15729, N4773, N11350, N3336);
and AND2 (N15732, N15702, N4402);
xor XOR2 (N15733, N15720, N1317);
xor XOR2 (N15734, N15728, N15015);
nor NOR4 (N15735, N15733, N13638, N4228, N1706);
buf BUF1 (N15736, N15726);
and AND3 (N15737, N15736, N13572, N2886);
nand NAND4 (N15738, N15732, N10837, N11982, N3307);
or OR2 (N15739, N15715, N6794);
xor XOR2 (N15740, N15725, N6406);
xor XOR2 (N15741, N15731, N13429);
buf BUF1 (N15742, N15722);
not NOT1 (N15743, N15739);
buf BUF1 (N15744, N15734);
nor NOR4 (N15745, N15742, N7401, N12326, N12891);
nand NAND4 (N15746, N15745, N12867, N7726, N4181);
nor NOR4 (N15747, N15737, N13881, N13363, N8500);
not NOT1 (N15748, N15746);
xor XOR2 (N15749, N15730, N1591);
not NOT1 (N15750, N15748);
not NOT1 (N15751, N15740);
buf BUF1 (N15752, N15735);
buf BUF1 (N15753, N15743);
or OR3 (N15754, N15738, N7837, N4886);
buf BUF1 (N15755, N15747);
buf BUF1 (N15756, N15724);
or OR4 (N15757, N15749, N13664, N9921, N12018);
nand NAND2 (N15758, N15752, N14041);
not NOT1 (N15759, N15750);
nor NOR3 (N15760, N15755, N8330, N5506);
and AND4 (N15761, N15760, N3868, N7208, N2463);
buf BUF1 (N15762, N15756);
nand NAND2 (N15763, N15753, N3155);
not NOT1 (N15764, N15744);
not NOT1 (N15765, N15751);
buf BUF1 (N15766, N15754);
and AND2 (N15767, N15766, N13261);
buf BUF1 (N15768, N15767);
not NOT1 (N15769, N15762);
and AND3 (N15770, N15763, N7238, N7300);
buf BUF1 (N15771, N15759);
or OR3 (N15772, N15768, N12372, N11592);
nand NAND3 (N15773, N15757, N4550, N7273);
buf BUF1 (N15774, N15769);
not NOT1 (N15775, N15774);
not NOT1 (N15776, N15758);
nor NOR4 (N15777, N15772, N2433, N13234, N7629);
and AND2 (N15778, N15775, N11697);
not NOT1 (N15779, N15776);
not NOT1 (N15780, N15770);
not NOT1 (N15781, N15778);
nor NOR4 (N15782, N15765, N5917, N13311, N7455);
not NOT1 (N15783, N15761);
xor XOR2 (N15784, N15771, N8491);
nor NOR4 (N15785, N15781, N2436, N14229, N2584);
not NOT1 (N15786, N15783);
nand NAND3 (N15787, N15773, N14972, N4921);
or OR2 (N15788, N15780, N8533);
or OR4 (N15789, N15787, N4410, N5801, N8737);
and AND4 (N15790, N15764, N1621, N5852, N10523);
nor NOR4 (N15791, N15785, N6387, N3011, N15299);
or OR3 (N15792, N15790, N6789, N9782);
not NOT1 (N15793, N15786);
buf BUF1 (N15794, N15791);
not NOT1 (N15795, N15792);
nand NAND2 (N15796, N15793, N13329);
or OR3 (N15797, N15796, N2910, N3975);
and AND3 (N15798, N15794, N9711, N10702);
not NOT1 (N15799, N15741);
nand NAND3 (N15800, N15798, N8253, N11156);
not NOT1 (N15801, N15788);
nor NOR4 (N15802, N15801, N6954, N4682, N6174);
not NOT1 (N15803, N15789);
nor NOR4 (N15804, N15800, N15176, N14549, N8564);
or OR3 (N15805, N15782, N2166, N5331);
nand NAND2 (N15806, N15784, N15762);
xor XOR2 (N15807, N15799, N6238);
not NOT1 (N15808, N15804);
buf BUF1 (N15809, N15803);
or OR3 (N15810, N15777, N3835, N1010);
buf BUF1 (N15811, N15805);
nand NAND2 (N15812, N15802, N11191);
xor XOR2 (N15813, N15812, N11853);
xor XOR2 (N15814, N15811, N1287);
xor XOR2 (N15815, N15809, N15173);
not NOT1 (N15816, N15815);
or OR4 (N15817, N15795, N2887, N9015, N6376);
and AND2 (N15818, N15817, N8544);
buf BUF1 (N15819, N15797);
xor XOR2 (N15820, N15813, N7131);
xor XOR2 (N15821, N15810, N1808);
xor XOR2 (N15822, N15820, N1791);
and AND3 (N15823, N15807, N11140, N5978);
not NOT1 (N15824, N15806);
buf BUF1 (N15825, N15779);
or OR3 (N15826, N15823, N9562, N7420);
nor NOR4 (N15827, N15826, N4572, N10965, N974);
nor NOR2 (N15828, N15818, N3324);
and AND2 (N15829, N15822, N9626);
nand NAND4 (N15830, N15824, N11244, N7486, N2852);
or OR4 (N15831, N15816, N12499, N8571, N8118);
xor XOR2 (N15832, N15830, N9256);
or OR3 (N15833, N15828, N11326, N15781);
nor NOR3 (N15834, N15829, N11144, N6475);
and AND4 (N15835, N15821, N5502, N13753, N3869);
and AND2 (N15836, N15827, N6547);
or OR4 (N15837, N15833, N7416, N10441, N5509);
nand NAND3 (N15838, N15836, N1937, N281);
xor XOR2 (N15839, N15819, N15075);
buf BUF1 (N15840, N15825);
xor XOR2 (N15841, N15808, N8444);
xor XOR2 (N15842, N15835, N1720);
buf BUF1 (N15843, N15834);
buf BUF1 (N15844, N15842);
xor XOR2 (N15845, N15841, N8526);
nor NOR2 (N15846, N15838, N14907);
and AND3 (N15847, N15846, N6871, N11589);
not NOT1 (N15848, N15814);
xor XOR2 (N15849, N15847, N4300);
xor XOR2 (N15850, N15844, N11472);
and AND3 (N15851, N15849, N8408, N4590);
not NOT1 (N15852, N15839);
buf BUF1 (N15853, N15843);
buf BUF1 (N15854, N15831);
not NOT1 (N15855, N15854);
nor NOR2 (N15856, N15851, N9832);
and AND2 (N15857, N15850, N15570);
and AND3 (N15858, N15832, N4247, N8360);
or OR2 (N15859, N15856, N313);
nand NAND2 (N15860, N15852, N8558);
nand NAND2 (N15861, N15840, N3808);
buf BUF1 (N15862, N15859);
and AND2 (N15863, N15857, N9540);
buf BUF1 (N15864, N15853);
nor NOR2 (N15865, N15864, N3514);
or OR4 (N15866, N15848, N833, N3467, N12242);
and AND3 (N15867, N15866, N7357, N4989);
not NOT1 (N15868, N15867);
nor NOR3 (N15869, N15860, N11970, N14318);
xor XOR2 (N15870, N15855, N8584);
nand NAND3 (N15871, N15845, N13505, N1938);
nor NOR2 (N15872, N15863, N9651);
not NOT1 (N15873, N15861);
nor NOR3 (N15874, N15873, N9142, N6364);
not NOT1 (N15875, N15858);
or OR2 (N15876, N15875, N9165);
nor NOR4 (N15877, N15874, N224, N8756, N2840);
xor XOR2 (N15878, N15870, N1419);
not NOT1 (N15879, N15837);
buf BUF1 (N15880, N15876);
nand NAND3 (N15881, N15878, N13783, N11066);
nand NAND2 (N15882, N15865, N3076);
and AND3 (N15883, N15882, N7088, N14729);
buf BUF1 (N15884, N15871);
xor XOR2 (N15885, N15881, N8723);
nor NOR3 (N15886, N15869, N6992, N9186);
buf BUF1 (N15887, N15862);
and AND2 (N15888, N15887, N10032);
not NOT1 (N15889, N15879);
xor XOR2 (N15890, N15880, N3495);
xor XOR2 (N15891, N15886, N12389);
not NOT1 (N15892, N15877);
or OR4 (N15893, N15885, N176, N6847, N1133);
nand NAND2 (N15894, N15883, N5706);
buf BUF1 (N15895, N15889);
or OR3 (N15896, N15868, N2208, N13090);
nor NOR2 (N15897, N15894, N14919);
nand NAND4 (N15898, N15892, N6199, N2769, N6805);
not NOT1 (N15899, N15888);
buf BUF1 (N15900, N15891);
or OR3 (N15901, N15898, N7145, N8285);
xor XOR2 (N15902, N15890, N2999);
nor NOR3 (N15903, N15895, N6421, N6280);
or OR3 (N15904, N15897, N14396, N10485);
nand NAND4 (N15905, N15904, N7775, N15720, N8166);
xor XOR2 (N15906, N15902, N10154);
buf BUF1 (N15907, N15896);
buf BUF1 (N15908, N15893);
not NOT1 (N15909, N15872);
nor NOR3 (N15910, N15901, N12371, N2697);
buf BUF1 (N15911, N15910);
xor XOR2 (N15912, N15899, N1882);
xor XOR2 (N15913, N15900, N11290);
buf BUF1 (N15914, N15911);
nand NAND2 (N15915, N15913, N4092);
and AND2 (N15916, N15915, N12814);
buf BUF1 (N15917, N15912);
and AND4 (N15918, N15908, N2245, N9148, N4051);
and AND4 (N15919, N15884, N13417, N10562, N11349);
nand NAND4 (N15920, N15905, N5804, N11071, N13199);
nor NOR2 (N15921, N15917, N4665);
nor NOR4 (N15922, N15914, N10989, N11397, N9984);
nor NOR3 (N15923, N15906, N15429, N12901);
nand NAND2 (N15924, N15919, N1971);
or OR4 (N15925, N15903, N10962, N8990, N2014);
xor XOR2 (N15926, N15924, N7250);
xor XOR2 (N15927, N15909, N829);
nor NOR3 (N15928, N15907, N824, N7660);
nand NAND3 (N15929, N15922, N2346, N10939);
or OR2 (N15930, N15927, N322);
xor XOR2 (N15931, N15925, N13626);
not NOT1 (N15932, N15930);
nand NAND2 (N15933, N15928, N2067);
buf BUF1 (N15934, N15932);
or OR3 (N15935, N15916, N13094, N15573);
not NOT1 (N15936, N15923);
or OR3 (N15937, N15918, N2343, N15082);
or OR3 (N15938, N15931, N9297, N15396);
xor XOR2 (N15939, N15920, N13223);
not NOT1 (N15940, N15933);
buf BUF1 (N15941, N15934);
nor NOR4 (N15942, N15940, N4964, N5254, N11771);
xor XOR2 (N15943, N15929, N11322);
nor NOR4 (N15944, N15939, N5606, N669, N2728);
or OR3 (N15945, N15935, N5295, N14813);
not NOT1 (N15946, N15944);
and AND4 (N15947, N15941, N6205, N8684, N2006);
and AND2 (N15948, N15946, N15613);
not NOT1 (N15949, N15948);
not NOT1 (N15950, N15936);
and AND4 (N15951, N15950, N860, N12408, N5815);
xor XOR2 (N15952, N15943, N14829);
and AND3 (N15953, N15942, N2482, N12777);
or OR2 (N15954, N15937, N14879);
buf BUF1 (N15955, N15945);
and AND3 (N15956, N15954, N7647, N2390);
and AND2 (N15957, N15951, N246);
not NOT1 (N15958, N15921);
not NOT1 (N15959, N15938);
or OR3 (N15960, N15956, N11960, N5800);
nand NAND3 (N15961, N15952, N2917, N13008);
not NOT1 (N15962, N15961);
buf BUF1 (N15963, N15949);
or OR2 (N15964, N15953, N4638);
buf BUF1 (N15965, N15962);
nand NAND2 (N15966, N15963, N9197);
buf BUF1 (N15967, N15955);
and AND2 (N15968, N15958, N2723);
buf BUF1 (N15969, N15957);
buf BUF1 (N15970, N15964);
nand NAND4 (N15971, N15947, N12575, N11910, N15653);
or OR3 (N15972, N15970, N7583, N4730);
and AND3 (N15973, N15967, N11793, N6460);
buf BUF1 (N15974, N15968);
not NOT1 (N15975, N15974);
nor NOR2 (N15976, N15975, N6519);
nor NOR3 (N15977, N15965, N10642, N14580);
and AND4 (N15978, N15926, N14144, N12418, N5065);
or OR4 (N15979, N15978, N409, N225, N14556);
or OR3 (N15980, N15966, N15950, N6379);
nand NAND3 (N15981, N15979, N2605, N11248);
nand NAND2 (N15982, N15976, N3006);
or OR4 (N15983, N15981, N11930, N4308, N14128);
buf BUF1 (N15984, N15971);
nand NAND3 (N15985, N15982, N2521, N15096);
nand NAND4 (N15986, N15985, N10684, N6065, N11173);
or OR4 (N15987, N15983, N9572, N15186, N11637);
not NOT1 (N15988, N15959);
not NOT1 (N15989, N15984);
not NOT1 (N15990, N15969);
xor XOR2 (N15991, N15986, N10509);
nand NAND4 (N15992, N15987, N10535, N3153, N2096);
or OR2 (N15993, N15989, N13646);
nand NAND4 (N15994, N15993, N15899, N7014, N14912);
not NOT1 (N15995, N15994);
nor NOR2 (N15996, N15995, N8589);
nor NOR2 (N15997, N15972, N1597);
nor NOR3 (N15998, N15992, N11234, N638);
and AND3 (N15999, N15998, N7878, N13301);
nand NAND2 (N16000, N15960, N12174);
buf BUF1 (N16001, N16000);
nand NAND3 (N16002, N15988, N8896, N8919);
nor NOR4 (N16003, N15990, N15949, N7267, N5727);
or OR4 (N16004, N15977, N14297, N3422, N2800);
or OR3 (N16005, N16003, N1999, N7966);
buf BUF1 (N16006, N15973);
or OR3 (N16007, N15996, N12861, N6712);
buf BUF1 (N16008, N16006);
and AND2 (N16009, N15991, N10269);
xor XOR2 (N16010, N16004, N11067);
nor NOR2 (N16011, N16002, N13153);
not NOT1 (N16012, N16008);
nand NAND4 (N16013, N16001, N11744, N5615, N1869);
xor XOR2 (N16014, N16010, N11247);
or OR4 (N16015, N16007, N9564, N296, N2905);
nor NOR2 (N16016, N16014, N10818);
nor NOR2 (N16017, N16013, N5478);
nand NAND4 (N16018, N15997, N8077, N7686, N8364);
and AND2 (N16019, N16005, N6182);
and AND3 (N16020, N15980, N673, N3791);
not NOT1 (N16021, N16019);
nand NAND3 (N16022, N16020, N11989, N14019);
not NOT1 (N16023, N16011);
and AND2 (N16024, N16015, N111);
endmodule