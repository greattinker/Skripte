// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N403,N408,N413,N411,N414,N407,N410,N406,N412,N416;

xor XOR2 (N17, N8, N1);
nand NAND3 (N18, N10, N1, N12);
and AND2 (N19, N17, N3);
not NOT1 (N20, N4);
xor XOR2 (N21, N3, N19);
buf BUF1 (N22, N12);
not NOT1 (N23, N3);
and AND3 (N24, N18, N17, N4);
xor XOR2 (N25, N24, N10);
or OR2 (N26, N25, N16);
not NOT1 (N27, N9);
not NOT1 (N28, N21);
nand NAND2 (N29, N11, N12);
or OR4 (N30, N14, N12, N20, N1);
and AND4 (N31, N6, N14, N14, N28);
buf BUF1 (N32, N29);
not NOT1 (N33, N21);
and AND2 (N34, N18, N29);
or OR4 (N35, N3, N3, N14, N9);
not NOT1 (N36, N26);
nand NAND2 (N37, N34, N31);
not NOT1 (N38, N34);
not NOT1 (N39, N22);
nor NOR4 (N40, N37, N26, N37, N35);
or OR2 (N41, N11, N6);
or OR3 (N42, N30, N29, N38);
xor XOR2 (N43, N6, N30);
nor NOR2 (N44, N23, N30);
nand NAND2 (N45, N36, N5);
buf BUF1 (N46, N40);
not NOT1 (N47, N33);
nand NAND4 (N48, N39, N30, N24, N8);
xor XOR2 (N49, N48, N28);
and AND3 (N50, N47, N20, N1);
and AND4 (N51, N45, N30, N10, N16);
or OR2 (N52, N27, N3);
xor XOR2 (N53, N49, N48);
xor XOR2 (N54, N32, N45);
buf BUF1 (N55, N54);
not NOT1 (N56, N53);
or OR2 (N57, N56, N41);
xor XOR2 (N58, N50, N11);
or OR4 (N59, N32, N54, N15, N15);
xor XOR2 (N60, N59, N46);
buf BUF1 (N61, N38);
and AND3 (N62, N57, N40, N47);
or OR2 (N63, N42, N37);
and AND3 (N64, N44, N47, N17);
and AND4 (N65, N64, N26, N61, N55);
not NOT1 (N66, N63);
or OR2 (N67, N35, N5);
or OR4 (N68, N31, N16, N20, N5);
buf BUF1 (N69, N66);
and AND4 (N70, N52, N16, N61, N7);
not NOT1 (N71, N65);
or OR3 (N72, N71, N24, N20);
not NOT1 (N73, N72);
nor NOR3 (N74, N70, N4, N55);
buf BUF1 (N75, N69);
and AND3 (N76, N51, N19, N35);
buf BUF1 (N77, N75);
or OR3 (N78, N62, N46, N49);
and AND3 (N79, N43, N41, N24);
xor XOR2 (N80, N79, N44);
not NOT1 (N81, N78);
and AND2 (N82, N60, N48);
nand NAND3 (N83, N76, N49, N82);
not NOT1 (N84, N26);
nor NOR2 (N85, N68, N8);
xor XOR2 (N86, N80, N15);
not NOT1 (N87, N67);
buf BUF1 (N88, N86);
xor XOR2 (N89, N58, N31);
and AND4 (N90, N74, N41, N60, N7);
xor XOR2 (N91, N90, N14);
nand NAND3 (N92, N83, N68, N80);
nand NAND3 (N93, N81, N54, N78);
buf BUF1 (N94, N73);
and AND3 (N95, N89, N31, N3);
nand NAND2 (N96, N84, N12);
not NOT1 (N97, N88);
or OR3 (N98, N77, N11, N67);
or OR2 (N99, N87, N75);
buf BUF1 (N100, N96);
not NOT1 (N101, N98);
and AND3 (N102, N97, N32, N12);
nand NAND2 (N103, N94, N63);
or OR3 (N104, N101, N90, N17);
not NOT1 (N105, N103);
nor NOR4 (N106, N102, N47, N82, N57);
or OR3 (N107, N93, N44, N105);
buf BUF1 (N108, N99);
or OR3 (N109, N23, N82, N57);
not NOT1 (N110, N106);
xor XOR2 (N111, N104, N74);
nor NOR3 (N112, N107, N76, N31);
nor NOR3 (N113, N92, N17, N47);
nand NAND3 (N114, N95, N88, N78);
nor NOR4 (N115, N85, N22, N85, N75);
nor NOR3 (N116, N109, N64, N69);
not NOT1 (N117, N115);
nor NOR2 (N118, N117, N83);
and AND4 (N119, N100, N56, N100, N3);
nor NOR4 (N120, N118, N49, N75, N34);
xor XOR2 (N121, N91, N62);
xor XOR2 (N122, N113, N53);
and AND4 (N123, N108, N39, N105, N121);
and AND4 (N124, N23, N98, N116, N55);
or OR2 (N125, N15, N20);
nand NAND3 (N126, N112, N82, N37);
not NOT1 (N127, N110);
nor NOR3 (N128, N122, N120, N119);
buf BUF1 (N129, N53);
xor XOR2 (N130, N37, N129);
nand NAND2 (N131, N19, N112);
buf BUF1 (N132, N114);
xor XOR2 (N133, N126, N83);
not NOT1 (N134, N128);
nand NAND4 (N135, N134, N129, N101, N106);
not NOT1 (N136, N123);
xor XOR2 (N137, N131, N16);
nand NAND2 (N138, N125, N17);
nand NAND2 (N139, N111, N87);
not NOT1 (N140, N127);
xor XOR2 (N141, N130, N21);
nand NAND2 (N142, N136, N57);
and AND3 (N143, N139, N101, N33);
xor XOR2 (N144, N133, N98);
not NOT1 (N145, N132);
nor NOR4 (N146, N141, N72, N136, N145);
or OR4 (N147, N11, N102, N72, N26);
nand NAND3 (N148, N144, N125, N120);
buf BUF1 (N149, N137);
and AND4 (N150, N142, N113, N39, N22);
and AND2 (N151, N135, N4);
buf BUF1 (N152, N138);
buf BUF1 (N153, N146);
buf BUF1 (N154, N151);
and AND3 (N155, N154, N101, N96);
buf BUF1 (N156, N148);
xor XOR2 (N157, N156, N81);
xor XOR2 (N158, N140, N134);
nand NAND4 (N159, N153, N96, N123, N57);
xor XOR2 (N160, N157, N81);
or OR2 (N161, N159, N118);
and AND3 (N162, N147, N128, N41);
or OR4 (N163, N152, N126, N26, N114);
not NOT1 (N164, N124);
nand NAND3 (N165, N155, N119, N98);
xor XOR2 (N166, N149, N36);
nor NOR3 (N167, N161, N88, N138);
xor XOR2 (N168, N166, N1);
xor XOR2 (N169, N143, N33);
nand NAND2 (N170, N164, N141);
nand NAND2 (N171, N167, N121);
buf BUF1 (N172, N170);
not NOT1 (N173, N171);
nand NAND3 (N174, N158, N5, N52);
and AND3 (N175, N168, N132, N27);
xor XOR2 (N176, N165, N127);
nand NAND2 (N177, N169, N23);
nor NOR3 (N178, N176, N167, N113);
nand NAND4 (N179, N172, N31, N54, N31);
and AND2 (N180, N175, N57);
not NOT1 (N181, N163);
not NOT1 (N182, N150);
and AND4 (N183, N179, N30, N54, N171);
not NOT1 (N184, N160);
and AND3 (N185, N177, N184, N18);
and AND3 (N186, N126, N173, N70);
nor NOR3 (N187, N146, N59, N34);
nand NAND3 (N188, N185, N2, N7);
nand NAND2 (N189, N180, N88);
xor XOR2 (N190, N174, N92);
and AND3 (N191, N178, N149, N110);
not NOT1 (N192, N191);
not NOT1 (N193, N192);
buf BUF1 (N194, N188);
or OR2 (N195, N183, N44);
and AND3 (N196, N182, N18, N97);
nand NAND4 (N197, N186, N147, N19, N48);
nand NAND2 (N198, N195, N54);
nand NAND4 (N199, N197, N116, N63, N162);
not NOT1 (N200, N67);
not NOT1 (N201, N200);
xor XOR2 (N202, N181, N84);
and AND4 (N203, N199, N42, N197, N43);
nand NAND4 (N204, N190, N88, N100, N98);
nor NOR3 (N205, N196, N182, N174);
buf BUF1 (N206, N203);
or OR2 (N207, N205, N123);
buf BUF1 (N208, N202);
nor NOR4 (N209, N208, N103, N184, N69);
nand NAND3 (N210, N209, N174, N178);
nand NAND4 (N211, N187, N207, N15, N128);
buf BUF1 (N212, N141);
nor NOR3 (N213, N193, N163, N44);
nor NOR3 (N214, N206, N16, N180);
nor NOR4 (N215, N201, N134, N18, N214);
buf BUF1 (N216, N74);
and AND3 (N217, N215, N209, N28);
and AND3 (N218, N216, N216, N129);
xor XOR2 (N219, N218, N189);
buf BUF1 (N220, N188);
nand NAND4 (N221, N212, N168, N113, N142);
buf BUF1 (N222, N198);
and AND2 (N223, N213, N204);
nor NOR2 (N224, N110, N2);
nor NOR3 (N225, N224, N68, N151);
buf BUF1 (N226, N222);
not NOT1 (N227, N220);
buf BUF1 (N228, N225);
xor XOR2 (N229, N227, N21);
and AND2 (N230, N211, N194);
or OR4 (N231, N81, N136, N74, N118);
or OR3 (N232, N226, N133, N152);
xor XOR2 (N233, N229, N79);
xor XOR2 (N234, N217, N104);
buf BUF1 (N235, N234);
and AND2 (N236, N230, N148);
buf BUF1 (N237, N233);
and AND2 (N238, N223, N45);
nor NOR4 (N239, N238, N126, N90, N179);
not NOT1 (N240, N236);
not NOT1 (N241, N239);
or OR2 (N242, N221, N170);
xor XOR2 (N243, N235, N53);
and AND2 (N244, N240, N19);
or OR4 (N245, N232, N91, N19, N207);
nor NOR4 (N246, N243, N87, N178, N55);
not NOT1 (N247, N228);
and AND2 (N248, N219, N41);
nand NAND4 (N249, N245, N33, N194, N160);
nor NOR3 (N250, N231, N9, N117);
buf BUF1 (N251, N250);
nand NAND4 (N252, N210, N133, N9, N249);
buf BUF1 (N253, N56);
nand NAND2 (N254, N247, N55);
xor XOR2 (N255, N241, N124);
buf BUF1 (N256, N251);
not NOT1 (N257, N255);
not NOT1 (N258, N252);
buf BUF1 (N259, N237);
or OR3 (N260, N259, N182, N35);
or OR4 (N261, N248, N180, N134, N259);
and AND4 (N262, N254, N187, N72, N239);
buf BUF1 (N263, N260);
and AND3 (N264, N244, N257, N34);
or OR3 (N265, N165, N98, N150);
nor NOR4 (N266, N263, N81, N54, N221);
and AND2 (N267, N256, N80);
buf BUF1 (N268, N261);
and AND3 (N269, N265, N72, N201);
xor XOR2 (N270, N258, N89);
and AND2 (N271, N270, N227);
xor XOR2 (N272, N269, N115);
xor XOR2 (N273, N246, N256);
or OR2 (N274, N273, N124);
buf BUF1 (N275, N264);
nand NAND4 (N276, N267, N242, N232, N208);
xor XOR2 (N277, N257, N29);
or OR4 (N278, N253, N16, N261, N217);
nor NOR4 (N279, N268, N221, N274, N234);
and AND2 (N280, N243, N118);
not NOT1 (N281, N272);
nor NOR4 (N282, N266, N272, N184, N17);
buf BUF1 (N283, N275);
nor NOR2 (N284, N279, N95);
buf BUF1 (N285, N262);
buf BUF1 (N286, N277);
nor NOR3 (N287, N285, N21, N87);
not NOT1 (N288, N287);
xor XOR2 (N289, N271, N245);
buf BUF1 (N290, N288);
nand NAND4 (N291, N290, N150, N1, N84);
nor NOR4 (N292, N283, N119, N98, N161);
not NOT1 (N293, N286);
nand NAND4 (N294, N289, N107, N90, N141);
and AND2 (N295, N276, N219);
nor NOR2 (N296, N281, N277);
buf BUF1 (N297, N280);
nand NAND3 (N298, N294, N135, N47);
buf BUF1 (N299, N296);
xor XOR2 (N300, N299, N249);
buf BUF1 (N301, N298);
buf BUF1 (N302, N300);
buf BUF1 (N303, N282);
not NOT1 (N304, N297);
xor XOR2 (N305, N304, N57);
nand NAND2 (N306, N305, N134);
and AND4 (N307, N295, N197, N19, N185);
and AND3 (N308, N302, N252, N191);
buf BUF1 (N309, N307);
or OR3 (N310, N284, N283, N146);
nor NOR2 (N311, N310, N182);
xor XOR2 (N312, N306, N120);
nor NOR3 (N313, N311, N157, N88);
or OR3 (N314, N291, N258, N250);
xor XOR2 (N315, N312, N63);
nand NAND2 (N316, N309, N73);
xor XOR2 (N317, N316, N162);
buf BUF1 (N318, N308);
nand NAND3 (N319, N301, N157, N194);
not NOT1 (N320, N318);
buf BUF1 (N321, N319);
xor XOR2 (N322, N320, N252);
and AND4 (N323, N293, N175, N153, N265);
and AND2 (N324, N292, N250);
not NOT1 (N325, N315);
nor NOR4 (N326, N317, N257, N238, N277);
not NOT1 (N327, N303);
not NOT1 (N328, N326);
or OR3 (N329, N328, N37, N33);
buf BUF1 (N330, N313);
buf BUF1 (N331, N278);
and AND2 (N332, N324, N220);
nor NOR4 (N333, N323, N280, N233, N187);
xor XOR2 (N334, N314, N317);
buf BUF1 (N335, N330);
buf BUF1 (N336, N322);
xor XOR2 (N337, N335, N135);
nor NOR2 (N338, N327, N232);
buf BUF1 (N339, N336);
buf BUF1 (N340, N333);
nand NAND4 (N341, N340, N160, N241, N128);
or OR4 (N342, N321, N175, N31, N195);
xor XOR2 (N343, N339, N245);
or OR2 (N344, N329, N130);
nand NAND3 (N345, N337, N146, N192);
xor XOR2 (N346, N342, N238);
xor XOR2 (N347, N343, N343);
or OR4 (N348, N325, N200, N28, N284);
and AND2 (N349, N348, N100);
xor XOR2 (N350, N334, N205);
nand NAND3 (N351, N350, N44, N55);
not NOT1 (N352, N345);
nor NOR3 (N353, N341, N181, N241);
or OR2 (N354, N352, N277);
nand NAND4 (N355, N331, N101, N110, N176);
nand NAND4 (N356, N355, N166, N129, N28);
buf BUF1 (N357, N349);
nand NAND4 (N358, N351, N110, N169, N160);
nor NOR2 (N359, N357, N68);
or OR3 (N360, N356, N121, N13);
xor XOR2 (N361, N344, N78);
nand NAND3 (N362, N332, N40, N66);
or OR3 (N363, N338, N210, N193);
buf BUF1 (N364, N354);
not NOT1 (N365, N362);
buf BUF1 (N366, N363);
or OR2 (N367, N353, N230);
and AND4 (N368, N347, N136, N131, N132);
and AND2 (N369, N361, N275);
buf BUF1 (N370, N358);
buf BUF1 (N371, N364);
not NOT1 (N372, N365);
nand NAND4 (N373, N372, N26, N314, N11);
not NOT1 (N374, N359);
not NOT1 (N375, N346);
and AND4 (N376, N373, N216, N191, N125);
and AND4 (N377, N360, N207, N45, N132);
not NOT1 (N378, N370);
and AND4 (N379, N369, N163, N172, N204);
buf BUF1 (N380, N367);
nor NOR3 (N381, N376, N137, N246);
nand NAND4 (N382, N368, N372, N244, N252);
nor NOR4 (N383, N382, N380, N79, N242);
xor XOR2 (N384, N152, N4);
nand NAND2 (N385, N384, N282);
not NOT1 (N386, N383);
xor XOR2 (N387, N378, N338);
nand NAND2 (N388, N377, N342);
not NOT1 (N389, N374);
not NOT1 (N390, N379);
buf BUF1 (N391, N366);
nand NAND4 (N392, N381, N26, N127, N224);
buf BUF1 (N393, N390);
and AND4 (N394, N387, N119, N14, N219);
nand NAND4 (N395, N391, N188, N28, N183);
and AND2 (N396, N385, N59);
not NOT1 (N397, N389);
nand NAND4 (N398, N375, N106, N109, N302);
not NOT1 (N399, N392);
xor XOR2 (N400, N395, N251);
nor NOR3 (N401, N394, N260, N373);
or OR4 (N402, N397, N170, N315, N118);
buf BUF1 (N403, N398);
or OR3 (N404, N393, N25, N24);
or OR3 (N405, N371, N118, N187);
buf BUF1 (N406, N388);
or OR3 (N407, N401, N3, N400);
nor NOR3 (N408, N286, N288, N73);
or OR3 (N409, N399, N398, N286);
and AND3 (N410, N402, N47, N80);
xor XOR2 (N411, N404, N27);
buf BUF1 (N412, N386);
xor XOR2 (N413, N409, N228);
and AND4 (N414, N396, N160, N66, N325);
not NOT1 (N415, N405);
nand NAND3 (N416, N415, N214, N256);
endmodule