// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N511,N513,N501,N505,N506,N496,N507,N482,N512,N514;

nor NOR4 (N15, N13, N8, N8, N1);
nand NAND4 (N16, N11, N14, N6, N11);
not NOT1 (N17, N9);
xor XOR2 (N18, N3, N10);
not NOT1 (N19, N11);
not NOT1 (N20, N6);
xor XOR2 (N21, N6, N2);
buf BUF1 (N22, N15);
buf BUF1 (N23, N13);
nor NOR3 (N24, N10, N7, N5);
buf BUF1 (N25, N16);
not NOT1 (N26, N7);
or OR4 (N27, N18, N5, N18, N25);
nor NOR3 (N28, N19, N6, N13);
or OR3 (N29, N3, N12, N9);
buf BUF1 (N30, N28);
not NOT1 (N31, N20);
not NOT1 (N32, N23);
nor NOR3 (N33, N31, N4, N1);
or OR3 (N34, N27, N25, N26);
and AND4 (N35, N21, N32, N12, N22);
xor XOR2 (N36, N1, N18);
nor NOR3 (N37, N24, N4, N11);
nand NAND3 (N38, N7, N23, N10);
nor NOR2 (N39, N30, N10);
not NOT1 (N40, N35);
buf BUF1 (N41, N35);
nand NAND2 (N42, N34, N36);
nand NAND3 (N43, N6, N14, N33);
xor XOR2 (N44, N36, N39);
or OR4 (N45, N7, N14, N24, N1);
or OR3 (N46, N41, N4, N31);
nor NOR2 (N47, N42, N5);
buf BUF1 (N48, N43);
or OR4 (N49, N44, N46, N20, N19);
xor XOR2 (N50, N37, N38);
or OR4 (N51, N17, N41, N10, N35);
nor NOR2 (N52, N4, N37);
not NOT1 (N53, N27);
and AND3 (N54, N47, N51, N5);
buf BUF1 (N55, N37);
not NOT1 (N56, N29);
and AND3 (N57, N54, N21, N17);
buf BUF1 (N58, N40);
xor XOR2 (N59, N48, N16);
or OR2 (N60, N53, N59);
not NOT1 (N61, N31);
or OR4 (N62, N55, N23, N3, N40);
nor NOR3 (N63, N52, N62, N33);
buf BUF1 (N64, N21);
or OR2 (N65, N61, N55);
or OR4 (N66, N64, N32, N5, N62);
nor NOR2 (N67, N58, N23);
buf BUF1 (N68, N56);
not NOT1 (N69, N63);
nand NAND4 (N70, N49, N32, N42, N45);
nor NOR4 (N71, N7, N11, N68, N8);
nor NOR2 (N72, N25, N50);
or OR4 (N73, N48, N37, N17, N8);
nor NOR2 (N74, N57, N60);
xor XOR2 (N75, N30, N54);
buf BUF1 (N76, N65);
buf BUF1 (N77, N66);
nand NAND2 (N78, N74, N72);
or OR3 (N79, N42, N74, N15);
xor XOR2 (N80, N73, N61);
buf BUF1 (N81, N80);
xor XOR2 (N82, N77, N24);
or OR2 (N83, N67, N62);
nand NAND3 (N84, N79, N75, N80);
not NOT1 (N85, N51);
nor NOR4 (N86, N83, N51, N40, N14);
xor XOR2 (N87, N85, N23);
nor NOR3 (N88, N86, N80, N47);
and AND4 (N89, N81, N68, N79, N8);
xor XOR2 (N90, N70, N44);
nor NOR2 (N91, N76, N13);
and AND2 (N92, N90, N39);
nor NOR4 (N93, N78, N47, N59, N77);
buf BUF1 (N94, N89);
nand NAND2 (N95, N82, N85);
buf BUF1 (N96, N92);
or OR4 (N97, N84, N76, N82, N6);
nor NOR4 (N98, N96, N70, N41, N25);
buf BUF1 (N99, N71);
nor NOR4 (N100, N87, N94, N23, N29);
nand NAND4 (N101, N47, N83, N44, N24);
nor NOR4 (N102, N101, N88, N66, N35);
and AND3 (N103, N26, N73, N12);
xor XOR2 (N104, N102, N67);
xor XOR2 (N105, N93, N68);
buf BUF1 (N106, N105);
nand NAND4 (N107, N99, N61, N11, N105);
buf BUF1 (N108, N103);
buf BUF1 (N109, N69);
xor XOR2 (N110, N106, N42);
or OR2 (N111, N107, N26);
nor NOR3 (N112, N95, N20, N92);
nor NOR2 (N113, N112, N22);
and AND3 (N114, N111, N54, N81);
nor NOR2 (N115, N110, N83);
not NOT1 (N116, N91);
xor XOR2 (N117, N114, N61);
xor XOR2 (N118, N109, N13);
nand NAND2 (N119, N104, N82);
xor XOR2 (N120, N118, N52);
or OR3 (N121, N97, N15, N52);
buf BUF1 (N122, N120);
nor NOR3 (N123, N115, N76, N36);
nor NOR4 (N124, N108, N12, N39, N20);
nand NAND4 (N125, N100, N48, N71, N2);
xor XOR2 (N126, N119, N63);
nand NAND4 (N127, N121, N62, N58, N79);
not NOT1 (N128, N123);
or OR2 (N129, N125, N72);
or OR2 (N130, N117, N10);
nor NOR2 (N131, N124, N37);
and AND3 (N132, N116, N22, N131);
not NOT1 (N133, N86);
xor XOR2 (N134, N133, N74);
nor NOR3 (N135, N132, N96, N86);
or OR2 (N136, N135, N105);
nor NOR2 (N137, N127, N67);
or OR4 (N138, N113, N65, N11, N98);
nand NAND3 (N139, N13, N10, N105);
or OR3 (N140, N129, N52, N108);
xor XOR2 (N141, N139, N68);
nor NOR4 (N142, N140, N137, N100, N85);
xor XOR2 (N143, N55, N113);
or OR3 (N144, N142, N23, N105);
nand NAND4 (N145, N141, N3, N74, N55);
nor NOR4 (N146, N134, N30, N87, N78);
xor XOR2 (N147, N122, N30);
not NOT1 (N148, N144);
xor XOR2 (N149, N126, N68);
xor XOR2 (N150, N145, N56);
nand NAND2 (N151, N128, N150);
buf BUF1 (N152, N121);
nand NAND2 (N153, N151, N3);
nor NOR4 (N154, N153, N3, N149, N93);
not NOT1 (N155, N79);
or OR2 (N156, N152, N41);
buf BUF1 (N157, N154);
nor NOR3 (N158, N156, N43, N104);
buf BUF1 (N159, N157);
nand NAND2 (N160, N147, N91);
nand NAND3 (N161, N136, N61, N64);
nor NOR4 (N162, N160, N110, N113, N29);
xor XOR2 (N163, N146, N66);
and AND2 (N164, N130, N72);
or OR4 (N165, N148, N30, N86, N10);
not NOT1 (N166, N155);
nand NAND4 (N167, N161, N36, N145, N85);
buf BUF1 (N168, N158);
not NOT1 (N169, N167);
xor XOR2 (N170, N138, N74);
nor NOR4 (N171, N168, N43, N95, N127);
buf BUF1 (N172, N162);
xor XOR2 (N173, N169, N165);
or OR3 (N174, N114, N141, N5);
and AND4 (N175, N172, N37, N161, N118);
buf BUF1 (N176, N170);
or OR4 (N177, N173, N144, N144, N90);
buf BUF1 (N178, N159);
and AND3 (N179, N175, N20, N133);
buf BUF1 (N180, N178);
and AND3 (N181, N143, N143, N178);
and AND2 (N182, N171, N151);
nor NOR4 (N183, N164, N120, N130, N121);
nor NOR2 (N184, N163, N24);
or OR3 (N185, N177, N114, N62);
buf BUF1 (N186, N179);
or OR3 (N187, N185, N16, N56);
or OR2 (N188, N182, N110);
or OR2 (N189, N188, N143);
or OR3 (N190, N174, N129, N156);
buf BUF1 (N191, N184);
xor XOR2 (N192, N186, N79);
buf BUF1 (N193, N166);
and AND3 (N194, N181, N40, N62);
and AND4 (N195, N191, N190, N59, N117);
not NOT1 (N196, N36);
nand NAND2 (N197, N195, N86);
xor XOR2 (N198, N180, N42);
and AND4 (N199, N198, N143, N178, N195);
xor XOR2 (N200, N187, N82);
xor XOR2 (N201, N192, N21);
buf BUF1 (N202, N193);
xor XOR2 (N203, N176, N12);
not NOT1 (N204, N202);
and AND3 (N205, N201, N163, N173);
or OR2 (N206, N203, N167);
and AND2 (N207, N196, N158);
xor XOR2 (N208, N189, N89);
buf BUF1 (N209, N205);
or OR3 (N210, N207, N23, N43);
and AND2 (N211, N199, N10);
buf BUF1 (N212, N208);
buf BUF1 (N213, N204);
xor XOR2 (N214, N194, N54);
and AND3 (N215, N211, N42, N96);
or OR4 (N216, N214, N16, N125, N148);
xor XOR2 (N217, N206, N67);
and AND3 (N218, N197, N98, N78);
and AND3 (N219, N209, N145, N23);
buf BUF1 (N220, N183);
xor XOR2 (N221, N213, N171);
and AND2 (N222, N217, N57);
buf BUF1 (N223, N218);
nand NAND4 (N224, N215, N171, N26, N44);
nand NAND3 (N225, N222, N142, N129);
not NOT1 (N226, N212);
buf BUF1 (N227, N216);
and AND4 (N228, N226, N5, N80, N213);
xor XOR2 (N229, N200, N184);
and AND4 (N230, N221, N190, N121, N178);
xor XOR2 (N231, N225, N11);
not NOT1 (N232, N228);
or OR4 (N233, N230, N221, N193, N97);
nand NAND2 (N234, N220, N28);
nand NAND2 (N235, N223, N66);
or OR2 (N236, N232, N142);
buf BUF1 (N237, N233);
xor XOR2 (N238, N236, N200);
not NOT1 (N239, N235);
buf BUF1 (N240, N237);
nor NOR4 (N241, N224, N192, N122, N97);
not NOT1 (N242, N240);
nand NAND4 (N243, N242, N10, N82, N215);
and AND2 (N244, N229, N88);
not NOT1 (N245, N244);
xor XOR2 (N246, N219, N128);
and AND4 (N247, N234, N31, N101, N89);
nor NOR2 (N248, N231, N170);
xor XOR2 (N249, N227, N246);
xor XOR2 (N250, N18, N26);
nand NAND4 (N251, N250, N68, N60, N7);
nor NOR4 (N252, N238, N151, N205, N96);
buf BUF1 (N253, N245);
not NOT1 (N254, N210);
or OR3 (N255, N249, N96, N139);
buf BUF1 (N256, N239);
and AND3 (N257, N251, N104, N216);
nor NOR3 (N258, N256, N181, N198);
not NOT1 (N259, N253);
xor XOR2 (N260, N257, N101);
nand NAND2 (N261, N252, N151);
or OR2 (N262, N243, N51);
not NOT1 (N263, N241);
buf BUF1 (N264, N260);
buf BUF1 (N265, N258);
not NOT1 (N266, N261);
xor XOR2 (N267, N254, N93);
nand NAND2 (N268, N248, N142);
nor NOR2 (N269, N255, N262);
not NOT1 (N270, N252);
not NOT1 (N271, N264);
not NOT1 (N272, N268);
and AND3 (N273, N247, N272, N197);
buf BUF1 (N274, N22);
buf BUF1 (N275, N267);
buf BUF1 (N276, N269);
nor NOR4 (N277, N265, N93, N189, N19);
nand NAND2 (N278, N271, N132);
xor XOR2 (N279, N278, N56);
and AND3 (N280, N259, N267, N118);
not NOT1 (N281, N270);
not NOT1 (N282, N266);
buf BUF1 (N283, N263);
or OR4 (N284, N277, N141, N90, N126);
or OR3 (N285, N283, N76, N139);
and AND4 (N286, N273, N144, N185, N260);
or OR4 (N287, N285, N80, N169, N67);
not NOT1 (N288, N284);
and AND3 (N289, N281, N130, N124);
buf BUF1 (N290, N276);
xor XOR2 (N291, N287, N196);
and AND4 (N292, N289, N138, N52, N160);
xor XOR2 (N293, N286, N85);
nand NAND2 (N294, N293, N259);
nor NOR3 (N295, N274, N49, N151);
buf BUF1 (N296, N275);
buf BUF1 (N297, N292);
buf BUF1 (N298, N295);
not NOT1 (N299, N294);
buf BUF1 (N300, N298);
xor XOR2 (N301, N300, N153);
buf BUF1 (N302, N296);
buf BUF1 (N303, N288);
or OR2 (N304, N279, N23);
nand NAND3 (N305, N304, N257, N292);
nor NOR3 (N306, N297, N91, N137);
xor XOR2 (N307, N306, N286);
nand NAND3 (N308, N299, N268, N24);
xor XOR2 (N309, N308, N237);
and AND2 (N310, N309, N38);
nor NOR4 (N311, N303, N21, N78, N261);
nand NAND3 (N312, N290, N269, N131);
and AND4 (N313, N311, N168, N47, N65);
not NOT1 (N314, N307);
buf BUF1 (N315, N280);
nor NOR3 (N316, N305, N290, N66);
and AND3 (N317, N301, N40, N199);
nand NAND4 (N318, N315, N194, N234, N267);
nand NAND4 (N319, N310, N314, N274, N141);
or OR3 (N320, N179, N143, N82);
buf BUF1 (N321, N312);
and AND3 (N322, N319, N77, N170);
nand NAND2 (N323, N318, N186);
xor XOR2 (N324, N320, N24);
xor XOR2 (N325, N291, N81);
nand NAND2 (N326, N313, N234);
buf BUF1 (N327, N322);
buf BUF1 (N328, N323);
not NOT1 (N329, N316);
or OR4 (N330, N321, N57, N186, N266);
not NOT1 (N331, N282);
and AND4 (N332, N328, N206, N302, N230);
nand NAND2 (N333, N315, N323);
not NOT1 (N334, N325);
buf BUF1 (N335, N333);
and AND2 (N336, N329, N6);
nand NAND4 (N337, N332, N243, N240, N251);
buf BUF1 (N338, N336);
nand NAND4 (N339, N326, N70, N331, N154);
nor NOR3 (N340, N55, N59, N233);
buf BUF1 (N341, N339);
buf BUF1 (N342, N337);
xor XOR2 (N343, N338, N152);
or OR4 (N344, N340, N234, N26, N212);
and AND2 (N345, N330, N175);
or OR4 (N346, N343, N131, N242, N245);
or OR2 (N347, N335, N10);
nand NAND4 (N348, N345, N222, N229, N4);
or OR3 (N349, N334, N330, N150);
and AND2 (N350, N344, N143);
buf BUF1 (N351, N350);
xor XOR2 (N352, N348, N232);
xor XOR2 (N353, N347, N260);
or OR3 (N354, N317, N168, N239);
nand NAND4 (N355, N346, N74, N190, N5);
nand NAND4 (N356, N349, N79, N234, N298);
not NOT1 (N357, N327);
xor XOR2 (N358, N351, N146);
nand NAND2 (N359, N354, N174);
xor XOR2 (N360, N356, N71);
xor XOR2 (N361, N324, N323);
nand NAND3 (N362, N341, N76, N91);
and AND4 (N363, N359, N213, N220, N337);
nor NOR3 (N364, N353, N115, N324);
xor XOR2 (N365, N361, N244);
not NOT1 (N366, N362);
buf BUF1 (N367, N358);
nor NOR4 (N368, N365, N21, N253, N141);
and AND4 (N369, N342, N313, N146, N277);
and AND3 (N370, N364, N23, N108);
buf BUF1 (N371, N370);
not NOT1 (N372, N360);
nand NAND2 (N373, N372, N298);
nor NOR3 (N374, N357, N76, N133);
or OR2 (N375, N366, N2);
buf BUF1 (N376, N352);
or OR3 (N377, N374, N271, N110);
buf BUF1 (N378, N375);
nor NOR3 (N379, N378, N213, N144);
xor XOR2 (N380, N367, N261);
nor NOR2 (N381, N355, N17);
or OR4 (N382, N373, N239, N144, N118);
nor NOR2 (N383, N369, N46);
or OR3 (N384, N381, N107, N19);
and AND4 (N385, N368, N366, N292, N131);
nor NOR2 (N386, N384, N50);
nor NOR4 (N387, N382, N23, N17, N265);
not NOT1 (N388, N383);
or OR3 (N389, N387, N145, N218);
buf BUF1 (N390, N386);
nand NAND2 (N391, N371, N179);
and AND4 (N392, N377, N96, N200, N230);
or OR4 (N393, N363, N285, N336, N364);
or OR3 (N394, N385, N49, N288);
not NOT1 (N395, N391);
buf BUF1 (N396, N389);
nor NOR4 (N397, N388, N25, N216, N391);
not NOT1 (N398, N376);
not NOT1 (N399, N395);
nand NAND3 (N400, N394, N163, N115);
xor XOR2 (N401, N380, N297);
not NOT1 (N402, N392);
nor NOR3 (N403, N400, N217, N69);
nand NAND4 (N404, N396, N330, N151, N113);
and AND3 (N405, N390, N353, N392);
buf BUF1 (N406, N405);
buf BUF1 (N407, N402);
buf BUF1 (N408, N379);
not NOT1 (N409, N397);
nand NAND2 (N410, N401, N393);
nand NAND3 (N411, N398, N278, N300);
xor XOR2 (N412, N331, N11);
xor XOR2 (N413, N404, N150);
xor XOR2 (N414, N411, N222);
nor NOR3 (N415, N412, N362, N194);
not NOT1 (N416, N407);
nor NOR4 (N417, N414, N332, N248, N175);
nor NOR4 (N418, N409, N218, N297, N19);
not NOT1 (N419, N418);
xor XOR2 (N420, N419, N162);
buf BUF1 (N421, N399);
or OR4 (N422, N420, N227, N24, N124);
nor NOR3 (N423, N410, N187, N328);
nor NOR3 (N424, N416, N337, N291);
and AND4 (N425, N422, N344, N406, N391);
or OR2 (N426, N90, N346);
nor NOR3 (N427, N423, N425, N157);
buf BUF1 (N428, N342);
or OR3 (N429, N426, N143, N206);
nor NOR3 (N430, N429, N171, N411);
or OR4 (N431, N403, N212, N85, N278);
nand NAND2 (N432, N431, N380);
buf BUF1 (N433, N427);
and AND2 (N434, N433, N426);
nand NAND3 (N435, N434, N293, N292);
buf BUF1 (N436, N435);
nor NOR2 (N437, N408, N400);
or OR4 (N438, N421, N130, N431, N383);
buf BUF1 (N439, N437);
nor NOR4 (N440, N439, N133, N347, N393);
or OR4 (N441, N413, N94, N207, N322);
not NOT1 (N442, N441);
or OR4 (N443, N428, N106, N21, N346);
nor NOR4 (N444, N436, N265, N134, N96);
buf BUF1 (N445, N444);
and AND4 (N446, N443, N383, N334, N213);
xor XOR2 (N447, N424, N399);
nand NAND4 (N448, N432, N433, N135, N103);
buf BUF1 (N449, N446);
xor XOR2 (N450, N417, N366);
not NOT1 (N451, N445);
buf BUF1 (N452, N430);
nor NOR2 (N453, N451, N238);
xor XOR2 (N454, N449, N111);
not NOT1 (N455, N452);
buf BUF1 (N456, N455);
nor NOR4 (N457, N415, N6, N356, N214);
xor XOR2 (N458, N447, N199);
not NOT1 (N459, N438);
and AND2 (N460, N456, N263);
and AND4 (N461, N454, N220, N260, N243);
nand NAND4 (N462, N457, N306, N88, N69);
xor XOR2 (N463, N458, N215);
xor XOR2 (N464, N459, N198);
nand NAND2 (N465, N464, N329);
buf BUF1 (N466, N440);
nand NAND3 (N467, N466, N291, N168);
not NOT1 (N468, N467);
not NOT1 (N469, N468);
not NOT1 (N470, N460);
nor NOR4 (N471, N448, N358, N178, N11);
or OR3 (N472, N470, N361, N295);
or OR3 (N473, N442, N171, N95);
buf BUF1 (N474, N465);
and AND4 (N475, N453, N51, N200, N244);
buf BUF1 (N476, N472);
and AND3 (N477, N475, N120, N251);
nand NAND2 (N478, N477, N88);
not NOT1 (N479, N471);
xor XOR2 (N480, N462, N244);
and AND3 (N481, N478, N193, N348);
nor NOR3 (N482, N473, N314, N195);
buf BUF1 (N483, N463);
and AND4 (N484, N476, N413, N341, N355);
nor NOR2 (N485, N483, N14);
or OR3 (N486, N479, N295, N434);
nand NAND3 (N487, N461, N412, N322);
not NOT1 (N488, N474);
or OR3 (N489, N488, N63, N345);
xor XOR2 (N490, N450, N34);
or OR4 (N491, N481, N447, N462, N140);
nand NAND3 (N492, N489, N366, N47);
buf BUF1 (N493, N491);
xor XOR2 (N494, N484, N41);
buf BUF1 (N495, N480);
or OR3 (N496, N490, N463, N132);
not NOT1 (N497, N495);
xor XOR2 (N498, N486, N464);
buf BUF1 (N499, N497);
xor XOR2 (N500, N485, N329);
nand NAND2 (N501, N492, N346);
buf BUF1 (N502, N493);
nor NOR3 (N503, N498, N260, N350);
buf BUF1 (N504, N500);
xor XOR2 (N505, N504, N16);
nor NOR3 (N506, N502, N103, N173);
nand NAND4 (N507, N494, N100, N287, N112);
xor XOR2 (N508, N499, N368);
and AND4 (N509, N508, N282, N100, N107);
nor NOR3 (N510, N503, N82, N408);
nand NAND3 (N511, N510, N391, N475);
nor NOR2 (N512, N487, N215);
xor XOR2 (N513, N469, N462);
not NOT1 (N514, N509);
endmodule