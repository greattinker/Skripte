// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N712,N703,N713,N714,N716,N707,N717,N711,N676,N718;

nand NAND3 (N19, N11, N14, N6);
and AND4 (N20, N17, N14, N17, N6);
buf BUF1 (N21, N15);
buf BUF1 (N22, N12);
nor NOR2 (N23, N11, N2);
xor XOR2 (N24, N11, N18);
buf BUF1 (N25, N20);
and AND4 (N26, N14, N13, N22, N3);
nand NAND2 (N27, N8, N4);
and AND4 (N28, N8, N5, N23, N6);
xor XOR2 (N29, N3, N17);
not NOT1 (N30, N17);
or OR2 (N31, N7, N10);
nor NOR3 (N32, N25, N18, N12);
nor NOR3 (N33, N30, N19, N20);
nor NOR2 (N34, N32, N10);
buf BUF1 (N35, N16);
and AND4 (N36, N27, N10, N3, N30);
nand NAND4 (N37, N21, N36, N18, N13);
not NOT1 (N38, N22);
or OR3 (N39, N33, N32, N2);
nor NOR2 (N40, N39, N7);
not NOT1 (N41, N34);
nor NOR4 (N42, N24, N24, N32, N35);
or OR4 (N43, N4, N16, N40, N25);
or OR4 (N44, N37, N4, N43, N5);
xor XOR2 (N45, N4, N26);
buf BUF1 (N46, N36);
buf BUF1 (N47, N20);
and AND4 (N48, N41, N9, N47, N22);
or OR4 (N49, N3, N35, N41, N14);
not NOT1 (N50, N31);
nor NOR2 (N51, N46, N25);
and AND3 (N52, N45, N24, N15);
or OR4 (N53, N51, N26, N34, N50);
nand NAND4 (N54, N42, N11, N37, N15);
xor XOR2 (N55, N43, N6);
or OR4 (N56, N52, N43, N9, N50);
nor NOR4 (N57, N53, N24, N10, N48);
or OR3 (N58, N36, N46, N57);
nor NOR2 (N59, N47, N27);
nor NOR2 (N60, N59, N57);
xor XOR2 (N61, N56, N6);
nand NAND4 (N62, N55, N41, N15, N3);
and AND4 (N63, N60, N19, N38, N46);
not NOT1 (N64, N58);
nand NAND3 (N65, N44, N1, N58);
nand NAND2 (N66, N39, N62);
buf BUF1 (N67, N59);
xor XOR2 (N68, N65, N31);
nand NAND2 (N69, N68, N53);
buf BUF1 (N70, N49);
nor NOR3 (N71, N54, N7, N17);
buf BUF1 (N72, N70);
not NOT1 (N73, N71);
nand NAND3 (N74, N69, N7, N48);
not NOT1 (N75, N67);
nor NOR2 (N76, N75, N71);
and AND3 (N77, N66, N55, N22);
xor XOR2 (N78, N74, N56);
xor XOR2 (N79, N28, N25);
and AND4 (N80, N79, N14, N56, N46);
xor XOR2 (N81, N73, N72);
not NOT1 (N82, N13);
buf BUF1 (N83, N81);
or OR4 (N84, N82, N78, N10, N23);
nand NAND3 (N85, N65, N21, N18);
buf BUF1 (N86, N64);
and AND4 (N87, N83, N53, N12, N70);
and AND3 (N88, N61, N51, N43);
or OR4 (N89, N84, N78, N78, N76);
xor XOR2 (N90, N7, N48);
and AND2 (N91, N89, N5);
nor NOR4 (N92, N85, N80, N50, N4);
xor XOR2 (N93, N2, N79);
buf BUF1 (N94, N91);
buf BUF1 (N95, N63);
buf BUF1 (N96, N86);
nand NAND2 (N97, N94, N44);
xor XOR2 (N98, N87, N88);
or OR4 (N99, N28, N98, N45, N26);
nor NOR2 (N100, N95, N5);
buf BUF1 (N101, N59);
nand NAND3 (N102, N100, N79, N17);
xor XOR2 (N103, N99, N92);
or OR2 (N104, N79, N22);
nor NOR4 (N105, N90, N37, N94, N39);
nor NOR2 (N106, N105, N61);
and AND2 (N107, N102, N105);
xor XOR2 (N108, N93, N22);
nand NAND4 (N109, N97, N58, N62, N10);
and AND4 (N110, N107, N90, N100, N23);
nor NOR4 (N111, N101, N31, N67, N14);
nand NAND2 (N112, N110, N34);
xor XOR2 (N113, N112, N104);
nor NOR3 (N114, N103, N79, N13);
not NOT1 (N115, N8);
buf BUF1 (N116, N114);
and AND3 (N117, N96, N37, N13);
xor XOR2 (N118, N106, N6);
nor NOR2 (N119, N111, N84);
xor XOR2 (N120, N119, N102);
not NOT1 (N121, N117);
buf BUF1 (N122, N77);
not NOT1 (N123, N113);
not NOT1 (N124, N122);
or OR2 (N125, N120, N35);
nand NAND3 (N126, N124, N85, N47);
buf BUF1 (N127, N109);
nand NAND3 (N128, N118, N9, N44);
xor XOR2 (N129, N29, N23);
xor XOR2 (N130, N128, N76);
buf BUF1 (N131, N123);
or OR3 (N132, N121, N124, N21);
or OR3 (N133, N127, N65, N28);
nand NAND3 (N134, N126, N80, N2);
nor NOR2 (N135, N125, N61);
nor NOR4 (N136, N115, N56, N94, N123);
not NOT1 (N137, N135);
or OR2 (N138, N130, N84);
nand NAND3 (N139, N138, N38, N122);
not NOT1 (N140, N133);
nor NOR3 (N141, N134, N83, N140);
or OR4 (N142, N36, N103, N124, N12);
and AND3 (N143, N131, N62, N106);
nor NOR4 (N144, N129, N62, N69, N32);
nor NOR4 (N145, N132, N76, N108, N13);
buf BUF1 (N146, N85);
nand NAND4 (N147, N143, N129, N58, N6);
xor XOR2 (N148, N139, N145);
buf BUF1 (N149, N72);
and AND2 (N150, N142, N37);
xor XOR2 (N151, N137, N125);
nand NAND2 (N152, N149, N116);
nand NAND2 (N153, N70, N120);
buf BUF1 (N154, N151);
nor NOR4 (N155, N141, N13, N59, N153);
nor NOR3 (N156, N132, N79, N28);
not NOT1 (N157, N144);
nor NOR2 (N158, N156, N3);
nand NAND4 (N159, N155, N139, N107, N144);
or OR2 (N160, N148, N59);
and AND4 (N161, N146, N100, N38, N130);
buf BUF1 (N162, N158);
nor NOR2 (N163, N136, N46);
not NOT1 (N164, N160);
or OR3 (N165, N147, N160, N15);
not NOT1 (N166, N165);
xor XOR2 (N167, N162, N155);
nor NOR4 (N168, N157, N128, N167, N85);
buf BUF1 (N169, N47);
nor NOR2 (N170, N164, N52);
and AND4 (N171, N163, N154, N54, N24);
nor NOR2 (N172, N27, N9);
not NOT1 (N173, N169);
xor XOR2 (N174, N171, N49);
and AND3 (N175, N152, N37, N134);
nand NAND4 (N176, N150, N168, N146, N45);
nor NOR3 (N177, N2, N48, N127);
or OR2 (N178, N176, N104);
nand NAND3 (N179, N175, N20, N131);
and AND2 (N180, N174, N30);
and AND3 (N181, N172, N17, N53);
and AND2 (N182, N170, N121);
or OR4 (N183, N182, N20, N113, N135);
nand NAND4 (N184, N173, N158, N39, N132);
and AND3 (N185, N159, N10, N113);
nor NOR2 (N186, N185, N62);
and AND4 (N187, N183, N103, N125, N50);
buf BUF1 (N188, N166);
xor XOR2 (N189, N186, N28);
nor NOR3 (N190, N179, N124, N9);
nor NOR4 (N191, N181, N56, N125, N129);
or OR3 (N192, N180, N114, N40);
or OR4 (N193, N178, N85, N187, N93);
xor XOR2 (N194, N6, N93);
nand NAND4 (N195, N188, N14, N134, N31);
xor XOR2 (N196, N191, N45);
or OR4 (N197, N177, N143, N64, N85);
xor XOR2 (N198, N195, N97);
xor XOR2 (N199, N189, N61);
nand NAND2 (N200, N194, N167);
xor XOR2 (N201, N192, N130);
nor NOR2 (N202, N190, N125);
and AND3 (N203, N193, N94, N75);
not NOT1 (N204, N200);
not NOT1 (N205, N204);
nor NOR3 (N206, N199, N153, N16);
buf BUF1 (N207, N198);
nand NAND3 (N208, N205, N95, N33);
and AND3 (N209, N161, N4, N150);
nor NOR3 (N210, N184, N137, N152);
nor NOR3 (N211, N203, N207, N68);
xor XOR2 (N212, N92, N7);
nand NAND2 (N213, N209, N212);
not NOT1 (N214, N15);
xor XOR2 (N215, N213, N33);
nand NAND2 (N216, N206, N180);
and AND2 (N217, N196, N38);
not NOT1 (N218, N217);
not NOT1 (N219, N211);
xor XOR2 (N220, N218, N29);
xor XOR2 (N221, N219, N126);
xor XOR2 (N222, N214, N194);
nor NOR2 (N223, N197, N20);
and AND2 (N224, N215, N26);
nand NAND2 (N225, N224, N49);
or OR4 (N226, N210, N146, N82, N184);
nor NOR3 (N227, N201, N3, N49);
nand NAND3 (N228, N227, N47, N35);
nand NAND3 (N229, N216, N38, N89);
xor XOR2 (N230, N226, N158);
and AND2 (N231, N208, N206);
buf BUF1 (N232, N222);
buf BUF1 (N233, N221);
nand NAND4 (N234, N232, N218, N81, N77);
xor XOR2 (N235, N231, N228);
nand NAND2 (N236, N185, N127);
nor NOR4 (N237, N235, N68, N10, N156);
buf BUF1 (N238, N230);
xor XOR2 (N239, N223, N164);
not NOT1 (N240, N225);
and AND2 (N241, N237, N232);
and AND4 (N242, N239, N35, N69, N38);
xor XOR2 (N243, N229, N107);
xor XOR2 (N244, N243, N22);
buf BUF1 (N245, N238);
nand NAND3 (N246, N244, N3, N15);
nor NOR4 (N247, N240, N95, N21, N154);
nand NAND2 (N248, N202, N6);
nand NAND2 (N249, N233, N76);
or OR2 (N250, N234, N203);
nor NOR4 (N251, N236, N9, N25, N127);
or OR4 (N252, N247, N31, N89, N247);
buf BUF1 (N253, N248);
xor XOR2 (N254, N249, N76);
not NOT1 (N255, N252);
not NOT1 (N256, N254);
xor XOR2 (N257, N245, N241);
or OR2 (N258, N182, N99);
nand NAND4 (N259, N242, N190, N105, N176);
nand NAND3 (N260, N220, N226, N157);
nor NOR2 (N261, N250, N137);
xor XOR2 (N262, N258, N110);
or OR4 (N263, N257, N167, N123, N221);
not NOT1 (N264, N261);
xor XOR2 (N265, N251, N214);
nor NOR4 (N266, N253, N124, N244, N111);
or OR2 (N267, N266, N234);
buf BUF1 (N268, N264);
and AND4 (N269, N263, N35, N151, N213);
and AND4 (N270, N255, N184, N141, N33);
nand NAND3 (N271, N256, N61, N233);
nand NAND2 (N272, N268, N49);
and AND3 (N273, N269, N84, N191);
nand NAND2 (N274, N259, N30);
and AND2 (N275, N246, N69);
or OR2 (N276, N267, N54);
buf BUF1 (N277, N271);
nor NOR3 (N278, N270, N229, N225);
xor XOR2 (N279, N260, N223);
nor NOR2 (N280, N273, N272);
not NOT1 (N281, N129);
not NOT1 (N282, N262);
nor NOR2 (N283, N278, N104);
or OR3 (N284, N280, N147, N17);
not NOT1 (N285, N275);
not NOT1 (N286, N285);
buf BUF1 (N287, N282);
or OR4 (N288, N274, N234, N202, N37);
nand NAND3 (N289, N288, N233, N197);
xor XOR2 (N290, N281, N232);
and AND2 (N291, N283, N287);
buf BUF1 (N292, N248);
and AND2 (N293, N289, N198);
buf BUF1 (N294, N293);
buf BUF1 (N295, N276);
or OR2 (N296, N279, N143);
nor NOR4 (N297, N295, N205, N143, N197);
buf BUF1 (N298, N294);
not NOT1 (N299, N265);
buf BUF1 (N300, N297);
nand NAND4 (N301, N296, N293, N141, N232);
or OR4 (N302, N290, N61, N144, N69);
and AND3 (N303, N302, N30, N137);
and AND4 (N304, N301, N94, N92, N266);
buf BUF1 (N305, N292);
xor XOR2 (N306, N277, N152);
or OR2 (N307, N299, N100);
not NOT1 (N308, N300);
not NOT1 (N309, N284);
xor XOR2 (N310, N308, N225);
and AND4 (N311, N309, N91, N296, N62);
xor XOR2 (N312, N298, N252);
nor NOR3 (N313, N291, N119, N307);
xor XOR2 (N314, N136, N20);
or OR4 (N315, N286, N76, N156, N75);
buf BUF1 (N316, N311);
nand NAND2 (N317, N303, N45);
xor XOR2 (N318, N305, N311);
xor XOR2 (N319, N314, N3);
nand NAND2 (N320, N313, N194);
nor NOR3 (N321, N316, N48, N219);
not NOT1 (N322, N312);
or OR3 (N323, N320, N33, N212);
xor XOR2 (N324, N321, N40);
or OR2 (N325, N324, N282);
and AND4 (N326, N310, N320, N129, N80);
and AND3 (N327, N304, N281, N29);
xor XOR2 (N328, N323, N27);
xor XOR2 (N329, N328, N320);
and AND2 (N330, N322, N152);
xor XOR2 (N331, N330, N157);
not NOT1 (N332, N317);
and AND2 (N333, N331, N47);
not NOT1 (N334, N319);
xor XOR2 (N335, N325, N162);
nand NAND2 (N336, N327, N44);
nor NOR3 (N337, N332, N321, N133);
xor XOR2 (N338, N337, N46);
not NOT1 (N339, N336);
nor NOR4 (N340, N338, N220, N133, N267);
and AND4 (N341, N340, N203, N27, N245);
buf BUF1 (N342, N306);
and AND3 (N343, N335, N58, N1);
nor NOR3 (N344, N342, N156, N226);
and AND3 (N345, N333, N123, N231);
nor NOR4 (N346, N326, N147, N237, N48);
or OR4 (N347, N329, N233, N260, N93);
not NOT1 (N348, N341);
not NOT1 (N349, N344);
and AND3 (N350, N315, N285, N224);
nand NAND2 (N351, N346, N163);
nand NAND3 (N352, N351, N66, N152);
nor NOR2 (N353, N347, N340);
nor NOR3 (N354, N339, N5, N39);
buf BUF1 (N355, N354);
and AND4 (N356, N355, N333, N72, N111);
xor XOR2 (N357, N345, N142);
buf BUF1 (N358, N356);
and AND3 (N359, N343, N123, N343);
buf BUF1 (N360, N318);
buf BUF1 (N361, N358);
buf BUF1 (N362, N350);
and AND4 (N363, N359, N131, N275, N52);
not NOT1 (N364, N349);
xor XOR2 (N365, N334, N360);
xor XOR2 (N366, N59, N252);
nor NOR2 (N367, N353, N360);
or OR3 (N368, N348, N80, N217);
and AND4 (N369, N368, N68, N356, N294);
or OR2 (N370, N366, N114);
nor NOR4 (N371, N370, N50, N164, N13);
nor NOR3 (N372, N367, N97, N343);
or OR3 (N373, N363, N259, N264);
nor NOR4 (N374, N373, N74, N29, N115);
xor XOR2 (N375, N361, N151);
nor NOR4 (N376, N374, N50, N374, N221);
buf BUF1 (N377, N369);
xor XOR2 (N378, N364, N332);
buf BUF1 (N379, N378);
nor NOR4 (N380, N379, N181, N187, N89);
buf BUF1 (N381, N365);
nand NAND3 (N382, N381, N155, N107);
nand NAND4 (N383, N357, N376, N304, N337);
and AND4 (N384, N12, N201, N92, N162);
not NOT1 (N385, N375);
not NOT1 (N386, N382);
nand NAND4 (N387, N362, N120, N352, N336);
nor NOR4 (N388, N257, N387, N378, N380);
xor XOR2 (N389, N298, N365);
and AND3 (N390, N382, N282, N370);
nor NOR2 (N391, N388, N44);
and AND3 (N392, N384, N51, N106);
xor XOR2 (N393, N372, N316);
not NOT1 (N394, N393);
buf BUF1 (N395, N394);
nand NAND4 (N396, N392, N203, N108, N252);
or OR2 (N397, N371, N316);
nor NOR3 (N398, N377, N281, N355);
xor XOR2 (N399, N391, N160);
or OR2 (N400, N399, N353);
or OR2 (N401, N396, N32);
nand NAND3 (N402, N385, N311, N124);
nand NAND2 (N403, N386, N119);
nand NAND3 (N404, N401, N289, N238);
not NOT1 (N405, N404);
xor XOR2 (N406, N397, N375);
buf BUF1 (N407, N398);
and AND4 (N408, N405, N248, N356, N396);
nand NAND3 (N409, N408, N379, N239);
nor NOR2 (N410, N400, N261);
or OR2 (N411, N395, N282);
not NOT1 (N412, N403);
nand NAND2 (N413, N383, N332);
nand NAND4 (N414, N389, N240, N300, N77);
buf BUF1 (N415, N409);
not NOT1 (N416, N415);
xor XOR2 (N417, N411, N81);
buf BUF1 (N418, N417);
and AND3 (N419, N402, N192, N415);
not NOT1 (N420, N414);
or OR4 (N421, N410, N401, N132, N182);
xor XOR2 (N422, N406, N270);
not NOT1 (N423, N418);
nand NAND2 (N424, N413, N25);
xor XOR2 (N425, N421, N277);
or OR3 (N426, N419, N107, N89);
and AND3 (N427, N420, N151, N203);
nor NOR4 (N428, N412, N38, N95, N149);
not NOT1 (N429, N390);
buf BUF1 (N430, N423);
not NOT1 (N431, N426);
nor NOR4 (N432, N422, N151, N70, N154);
xor XOR2 (N433, N424, N334);
nand NAND3 (N434, N425, N295, N252);
and AND3 (N435, N416, N132, N318);
xor XOR2 (N436, N434, N282);
xor XOR2 (N437, N432, N111);
not NOT1 (N438, N428);
not NOT1 (N439, N433);
or OR3 (N440, N437, N192, N378);
not NOT1 (N441, N407);
or OR3 (N442, N441, N175, N276);
nand NAND3 (N443, N430, N175, N260);
and AND2 (N444, N442, N110);
or OR3 (N445, N429, N131, N414);
nor NOR4 (N446, N444, N402, N234, N83);
buf BUF1 (N447, N436);
buf BUF1 (N448, N440);
nand NAND4 (N449, N447, N282, N287, N74);
buf BUF1 (N450, N435);
nand NAND3 (N451, N431, N132, N183);
buf BUF1 (N452, N448);
and AND2 (N453, N443, N355);
and AND4 (N454, N446, N210, N248, N153);
and AND4 (N455, N452, N332, N376, N347);
not NOT1 (N456, N451);
or OR4 (N457, N438, N456, N311, N257);
not NOT1 (N458, N43);
or OR3 (N459, N439, N258, N318);
nor NOR4 (N460, N459, N206, N333, N157);
xor XOR2 (N461, N454, N411);
not NOT1 (N462, N455);
nand NAND4 (N463, N450, N85, N437, N291);
not NOT1 (N464, N462);
buf BUF1 (N465, N445);
xor XOR2 (N466, N427, N155);
and AND2 (N467, N457, N84);
and AND4 (N468, N465, N418, N180, N83);
or OR2 (N469, N466, N53);
xor XOR2 (N470, N460, N86);
nor NOR4 (N471, N449, N400, N447, N384);
buf BUF1 (N472, N470);
nand NAND2 (N473, N472, N26);
buf BUF1 (N474, N468);
xor XOR2 (N475, N453, N227);
nor NOR4 (N476, N467, N465, N227, N171);
or OR4 (N477, N464, N293, N404, N140);
nor NOR2 (N478, N471, N47);
or OR2 (N479, N463, N471);
nor NOR4 (N480, N476, N291, N201, N56);
not NOT1 (N481, N473);
and AND4 (N482, N477, N145, N58, N90);
nor NOR2 (N483, N475, N63);
xor XOR2 (N484, N480, N4);
nand NAND3 (N485, N461, N482, N179);
xor XOR2 (N486, N405, N307);
not NOT1 (N487, N486);
xor XOR2 (N488, N487, N219);
or OR4 (N489, N479, N448, N53, N261);
buf BUF1 (N490, N481);
or OR2 (N491, N469, N306);
xor XOR2 (N492, N474, N451);
nand NAND3 (N493, N491, N201, N484);
and AND2 (N494, N292, N368);
not NOT1 (N495, N478);
nand NAND2 (N496, N494, N298);
nor NOR2 (N497, N458, N149);
and AND2 (N498, N485, N353);
buf BUF1 (N499, N497);
nor NOR4 (N500, N496, N403, N170, N350);
not NOT1 (N501, N488);
buf BUF1 (N502, N501);
nor NOR4 (N503, N483, N109, N376, N489);
buf BUF1 (N504, N97);
nor NOR4 (N505, N504, N491, N240, N169);
buf BUF1 (N506, N505);
buf BUF1 (N507, N498);
xor XOR2 (N508, N503, N247);
and AND2 (N509, N507, N404);
nand NAND3 (N510, N502, N244, N224);
xor XOR2 (N511, N495, N267);
nand NAND4 (N512, N493, N160, N463, N95);
xor XOR2 (N513, N512, N359);
not NOT1 (N514, N509);
nand NAND2 (N515, N490, N140);
xor XOR2 (N516, N500, N464);
nor NOR3 (N517, N514, N19, N124);
nor NOR2 (N518, N517, N46);
or OR4 (N519, N499, N72, N128, N259);
nand NAND3 (N520, N515, N36, N156);
and AND4 (N521, N519, N201, N497, N287);
not NOT1 (N522, N506);
xor XOR2 (N523, N513, N141);
not NOT1 (N524, N520);
and AND4 (N525, N523, N7, N181, N373);
not NOT1 (N526, N522);
xor XOR2 (N527, N526, N258);
xor XOR2 (N528, N524, N423);
buf BUF1 (N529, N521);
buf BUF1 (N530, N528);
nor NOR3 (N531, N510, N283, N263);
nor NOR2 (N532, N531, N441);
xor XOR2 (N533, N518, N161);
xor XOR2 (N534, N529, N399);
not NOT1 (N535, N492);
buf BUF1 (N536, N508);
xor XOR2 (N537, N511, N192);
not NOT1 (N538, N536);
or OR2 (N539, N533, N117);
and AND4 (N540, N530, N534, N81, N460);
or OR2 (N541, N105, N428);
nand NAND3 (N542, N525, N201, N344);
xor XOR2 (N543, N532, N229);
nor NOR4 (N544, N516, N243, N237, N425);
nand NAND3 (N545, N539, N381, N331);
nand NAND4 (N546, N545, N243, N162, N167);
xor XOR2 (N547, N537, N315);
buf BUF1 (N548, N538);
or OR4 (N549, N544, N259, N431, N442);
not NOT1 (N550, N542);
buf BUF1 (N551, N540);
nand NAND4 (N552, N549, N183, N199, N216);
or OR4 (N553, N547, N230, N175, N57);
nand NAND2 (N554, N548, N475);
nor NOR3 (N555, N546, N201, N89);
buf BUF1 (N556, N552);
nor NOR2 (N557, N535, N105);
not NOT1 (N558, N541);
and AND3 (N559, N551, N270, N400);
and AND3 (N560, N553, N117, N442);
not NOT1 (N561, N558);
buf BUF1 (N562, N557);
or OR4 (N563, N556, N40, N503, N369);
xor XOR2 (N564, N560, N105);
buf BUF1 (N565, N543);
xor XOR2 (N566, N561, N255);
nor NOR2 (N567, N565, N320);
not NOT1 (N568, N527);
nand NAND2 (N569, N564, N30);
or OR3 (N570, N559, N152, N248);
buf BUF1 (N571, N554);
xor XOR2 (N572, N569, N167);
and AND3 (N573, N563, N334, N536);
or OR3 (N574, N572, N448, N322);
nor NOR2 (N575, N568, N416);
not NOT1 (N576, N575);
buf BUF1 (N577, N567);
buf BUF1 (N578, N573);
xor XOR2 (N579, N576, N539);
xor XOR2 (N580, N577, N392);
buf BUF1 (N581, N562);
nor NOR2 (N582, N580, N247);
xor XOR2 (N583, N579, N528);
not NOT1 (N584, N582);
buf BUF1 (N585, N578);
buf BUF1 (N586, N570);
nand NAND2 (N587, N574, N503);
xor XOR2 (N588, N585, N359);
xor XOR2 (N589, N555, N366);
and AND2 (N590, N584, N111);
nand NAND4 (N591, N571, N523, N491, N90);
nor NOR3 (N592, N588, N406, N191);
and AND4 (N593, N583, N303, N229, N518);
not NOT1 (N594, N590);
xor XOR2 (N595, N581, N114);
and AND2 (N596, N586, N82);
or OR3 (N597, N594, N555, N218);
and AND4 (N598, N595, N7, N464, N295);
nor NOR2 (N599, N587, N179);
or OR4 (N600, N589, N231, N422, N393);
or OR2 (N601, N591, N221);
not NOT1 (N602, N593);
nor NOR3 (N603, N601, N222, N577);
xor XOR2 (N604, N602, N99);
or OR3 (N605, N566, N206, N119);
or OR3 (N606, N603, N602, N64);
nor NOR3 (N607, N592, N215, N412);
xor XOR2 (N608, N607, N569);
nor NOR4 (N609, N606, N124, N386, N288);
or OR2 (N610, N596, N302);
xor XOR2 (N611, N598, N344);
nand NAND4 (N612, N608, N387, N540, N175);
nand NAND2 (N613, N597, N263);
buf BUF1 (N614, N613);
buf BUF1 (N615, N604);
xor XOR2 (N616, N605, N141);
not NOT1 (N617, N616);
and AND3 (N618, N550, N596, N203);
nor NOR3 (N619, N599, N483, N458);
nand NAND2 (N620, N618, N75);
and AND3 (N621, N600, N222, N51);
nand NAND2 (N622, N609, N317);
nand NAND3 (N623, N611, N417, N79);
nand NAND3 (N624, N612, N412, N290);
not NOT1 (N625, N610);
or OR3 (N626, N622, N432, N15);
or OR4 (N627, N624, N156, N547, N594);
not NOT1 (N628, N621);
nand NAND3 (N629, N620, N459, N62);
or OR4 (N630, N629, N396, N485, N465);
or OR2 (N631, N623, N483);
xor XOR2 (N632, N614, N230);
nand NAND4 (N633, N627, N453, N625, N159);
xor XOR2 (N634, N345, N103);
xor XOR2 (N635, N626, N139);
xor XOR2 (N636, N635, N560);
and AND4 (N637, N615, N57, N154, N503);
buf BUF1 (N638, N634);
xor XOR2 (N639, N633, N357);
buf BUF1 (N640, N619);
nor NOR4 (N641, N632, N366, N602, N164);
nand NAND4 (N642, N636, N357, N195, N435);
nand NAND4 (N643, N617, N384, N363, N161);
and AND4 (N644, N640, N150, N598, N560);
or OR4 (N645, N631, N133, N32, N553);
buf BUF1 (N646, N643);
buf BUF1 (N647, N638);
and AND4 (N648, N630, N96, N249, N25);
buf BUF1 (N649, N642);
or OR2 (N650, N646, N576);
or OR4 (N651, N645, N389, N337, N158);
and AND2 (N652, N647, N644);
nor NOR2 (N653, N641, N321);
nor NOR3 (N654, N327, N114, N481);
nor NOR4 (N655, N651, N220, N589, N261);
xor XOR2 (N656, N648, N619);
buf BUF1 (N657, N639);
xor XOR2 (N658, N657, N568);
not NOT1 (N659, N650);
nand NAND2 (N660, N652, N161);
not NOT1 (N661, N628);
nor NOR2 (N662, N660, N598);
xor XOR2 (N663, N654, N24);
nand NAND4 (N664, N663, N130, N182, N189);
nor NOR4 (N665, N658, N461, N434, N627);
xor XOR2 (N666, N665, N26);
not NOT1 (N667, N656);
xor XOR2 (N668, N661, N275);
buf BUF1 (N669, N655);
buf BUF1 (N670, N666);
nand NAND2 (N671, N659, N420);
xor XOR2 (N672, N664, N249);
not NOT1 (N673, N653);
and AND2 (N674, N637, N429);
xor XOR2 (N675, N672, N501);
xor XOR2 (N676, N662, N305);
nor NOR2 (N677, N668, N260);
xor XOR2 (N678, N671, N161);
nor NOR2 (N679, N649, N604);
nor NOR4 (N680, N670, N622, N584, N287);
xor XOR2 (N681, N675, N232);
nand NAND2 (N682, N669, N153);
not NOT1 (N683, N681);
xor XOR2 (N684, N677, N311);
buf BUF1 (N685, N684);
nor NOR4 (N686, N673, N497, N150, N17);
nor NOR3 (N687, N683, N331, N298);
not NOT1 (N688, N679);
xor XOR2 (N689, N682, N54);
nand NAND2 (N690, N685, N639);
not NOT1 (N691, N678);
xor XOR2 (N692, N690, N512);
xor XOR2 (N693, N688, N90);
and AND4 (N694, N687, N631, N312, N620);
or OR3 (N695, N693, N471, N426);
and AND3 (N696, N680, N499, N207);
and AND2 (N697, N674, N537);
nand NAND3 (N698, N696, N488, N146);
nor NOR2 (N699, N689, N408);
nand NAND4 (N700, N667, N197, N615, N451);
buf BUF1 (N701, N698);
nor NOR2 (N702, N699, N138);
nor NOR4 (N703, N695, N398, N165, N154);
not NOT1 (N704, N692);
nand NAND3 (N705, N700, N522, N193);
nand NAND2 (N706, N697, N73);
not NOT1 (N707, N702);
buf BUF1 (N708, N694);
not NOT1 (N709, N701);
buf BUF1 (N710, N691);
buf BUF1 (N711, N709);
nor NOR3 (N712, N704, N591, N396);
and AND3 (N713, N708, N5, N181);
xor XOR2 (N714, N686, N472);
not NOT1 (N715, N706);
buf BUF1 (N716, N705);
nor NOR2 (N717, N715, N312);
buf BUF1 (N718, N710);
endmodule