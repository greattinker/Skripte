// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N7999,N8006,N7998,N8008,N8009,N7991,N8003,N7992,N8001,N8010;

xor XOR2 (N11, N8, N1);
and AND3 (N12, N8, N3, N7);
or OR3 (N13, N10, N7, N4);
nor NOR4 (N14, N1, N7, N4, N3);
and AND3 (N15, N11, N3, N8);
and AND4 (N16, N8, N15, N9, N4);
not NOT1 (N17, N2);
nor NOR4 (N18, N1, N3, N5, N12);
xor XOR2 (N19, N10, N13);
nand NAND2 (N20, N17, N13);
nand NAND3 (N21, N5, N18, N16);
nor NOR2 (N22, N6, N2);
xor XOR2 (N23, N13, N17);
buf BUF1 (N24, N20);
and AND2 (N25, N17, N16);
not NOT1 (N26, N2);
xor XOR2 (N27, N14, N14);
nand NAND4 (N28, N17, N6, N19, N13);
xor XOR2 (N29, N7, N11);
nor NOR2 (N30, N22, N3);
not NOT1 (N31, N29);
nor NOR3 (N32, N11, N8, N1);
buf BUF1 (N33, N24);
not NOT1 (N34, N25);
not NOT1 (N35, N34);
and AND3 (N36, N23, N6, N26);
and AND2 (N37, N36, N27);
not NOT1 (N38, N24);
and AND3 (N39, N5, N25, N18);
nor NOR2 (N40, N32, N27);
or OR2 (N41, N35, N14);
and AND2 (N42, N31, N39);
and AND4 (N43, N2, N2, N33, N9);
nor NOR2 (N44, N21, N11);
and AND4 (N45, N17, N12, N17, N5);
nor NOR4 (N46, N40, N27, N8, N22);
xor XOR2 (N47, N42, N17);
or OR3 (N48, N41, N38, N30);
buf BUF1 (N49, N41);
or OR3 (N50, N37, N46, N37);
nor NOR4 (N51, N1, N2, N15, N19);
or OR2 (N52, N15, N4);
and AND4 (N53, N50, N11, N3, N6);
and AND2 (N54, N48, N50);
nor NOR3 (N55, N47, N40, N15);
nor NOR3 (N56, N28, N16, N26);
not NOT1 (N57, N43);
xor XOR2 (N58, N57, N33);
nand NAND2 (N59, N49, N52);
buf BUF1 (N60, N29);
not NOT1 (N61, N59);
or OR4 (N62, N55, N31, N34, N16);
buf BUF1 (N63, N51);
and AND4 (N64, N62, N45, N44, N49);
xor XOR2 (N65, N33, N17);
and AND2 (N66, N64, N58);
or OR3 (N67, N63, N4, N3);
and AND2 (N68, N11, N20);
nand NAND4 (N69, N30, N1, N40, N18);
nor NOR4 (N70, N67, N49, N50, N50);
nor NOR3 (N71, N54, N69, N34);
buf BUF1 (N72, N2);
nand NAND3 (N73, N66, N1, N63);
nand NAND4 (N74, N70, N23, N16, N68);
buf BUF1 (N75, N62);
not NOT1 (N76, N65);
xor XOR2 (N77, N72, N28);
not NOT1 (N78, N76);
and AND3 (N79, N75, N56, N43);
and AND2 (N80, N35, N69);
or OR4 (N81, N80, N23, N24, N32);
xor XOR2 (N82, N74, N28);
nand NAND4 (N83, N53, N76, N26, N68);
xor XOR2 (N84, N73, N13);
nand NAND3 (N85, N81, N31, N77);
buf BUF1 (N86, N53);
or OR4 (N87, N61, N73, N69, N8);
nand NAND2 (N88, N83, N60);
not NOT1 (N89, N44);
nand NAND4 (N90, N85, N43, N38, N13);
nor NOR2 (N91, N90, N69);
nor NOR4 (N92, N86, N79, N76, N5);
nand NAND2 (N93, N91, N68);
not NOT1 (N94, N60);
buf BUF1 (N95, N92);
and AND2 (N96, N78, N52);
and AND2 (N97, N89, N23);
nand NAND4 (N98, N82, N74, N90, N75);
or OR4 (N99, N88, N32, N7, N26);
xor XOR2 (N100, N97, N92);
and AND2 (N101, N87, N6);
xor XOR2 (N102, N71, N3);
nand NAND4 (N103, N95, N78, N54, N14);
not NOT1 (N104, N103);
nand NAND2 (N105, N101, N7);
and AND4 (N106, N105, N51, N6, N3);
nand NAND2 (N107, N104, N30);
nand NAND2 (N108, N93, N52);
buf BUF1 (N109, N94);
buf BUF1 (N110, N100);
nand NAND2 (N111, N102, N69);
or OR3 (N112, N111, N65, N79);
nor NOR2 (N113, N110, N99);
nand NAND3 (N114, N71, N83, N57);
and AND4 (N115, N84, N32, N11, N78);
and AND4 (N116, N115, N72, N31, N7);
or OR4 (N117, N107, N8, N67, N69);
or OR3 (N118, N106, N8, N67);
nand NAND2 (N119, N112, N56);
nor NOR3 (N120, N98, N80, N69);
or OR4 (N121, N119, N104, N9, N20);
or OR3 (N122, N96, N77, N102);
xor XOR2 (N123, N122, N78);
nor NOR4 (N124, N120, N65, N25, N38);
nor NOR2 (N125, N124, N7);
nor NOR3 (N126, N121, N82, N78);
and AND2 (N127, N108, N13);
xor XOR2 (N128, N126, N84);
and AND2 (N129, N116, N45);
buf BUF1 (N130, N129);
nor NOR3 (N131, N114, N125, N6);
buf BUF1 (N132, N39);
xor XOR2 (N133, N113, N109);
not NOT1 (N134, N123);
nor NOR4 (N135, N123, N7, N63, N19);
nand NAND2 (N136, N128, N71);
xor XOR2 (N137, N136, N9);
and AND2 (N138, N117, N1);
buf BUF1 (N139, N133);
xor XOR2 (N140, N139, N91);
or OR4 (N141, N140, N83, N52, N23);
not NOT1 (N142, N135);
or OR3 (N143, N134, N104, N8);
or OR4 (N144, N118, N69, N128, N45);
or OR4 (N145, N130, N80, N64, N12);
xor XOR2 (N146, N132, N141);
not NOT1 (N147, N109);
xor XOR2 (N148, N127, N115);
not NOT1 (N149, N145);
nand NAND3 (N150, N146, N112, N25);
nand NAND2 (N151, N150, N147);
nand NAND2 (N152, N40, N128);
not NOT1 (N153, N143);
and AND4 (N154, N138, N107, N136, N95);
buf BUF1 (N155, N152);
nand NAND3 (N156, N153, N115, N62);
and AND2 (N157, N131, N134);
buf BUF1 (N158, N144);
buf BUF1 (N159, N151);
not NOT1 (N160, N158);
nand NAND3 (N161, N155, N50, N109);
buf BUF1 (N162, N137);
xor XOR2 (N163, N149, N153);
xor XOR2 (N164, N160, N85);
and AND3 (N165, N156, N127, N9);
xor XOR2 (N166, N142, N71);
xor XOR2 (N167, N161, N107);
not NOT1 (N168, N162);
or OR3 (N169, N168, N76, N115);
and AND3 (N170, N154, N33, N83);
and AND2 (N171, N170, N160);
and AND3 (N172, N169, N161, N48);
buf BUF1 (N173, N166);
not NOT1 (N174, N171);
and AND4 (N175, N159, N39, N144, N133);
or OR3 (N176, N172, N12, N170);
xor XOR2 (N177, N148, N81);
not NOT1 (N178, N177);
nand NAND3 (N179, N178, N28, N59);
nor NOR3 (N180, N163, N164, N1);
nand NAND4 (N181, N105, N140, N141, N179);
or OR4 (N182, N64, N174, N141, N34);
or OR3 (N183, N7, N31, N175);
xor XOR2 (N184, N98, N137);
buf BUF1 (N185, N180);
buf BUF1 (N186, N165);
and AND3 (N187, N157, N135, N180);
buf BUF1 (N188, N176);
nor NOR4 (N189, N182, N66, N130, N114);
nor NOR4 (N190, N167, N31, N161, N97);
and AND3 (N191, N184, N143, N71);
not NOT1 (N192, N173);
xor XOR2 (N193, N188, N48);
or OR3 (N194, N181, N144, N43);
not NOT1 (N195, N186);
and AND2 (N196, N183, N139);
buf BUF1 (N197, N196);
nand NAND3 (N198, N185, N124, N147);
xor XOR2 (N199, N194, N7);
nand NAND2 (N200, N189, N39);
buf BUF1 (N201, N200);
nand NAND2 (N202, N197, N106);
and AND2 (N203, N190, N165);
nor NOR3 (N204, N187, N95, N166);
buf BUF1 (N205, N204);
and AND4 (N206, N193, N58, N96, N46);
nand NAND2 (N207, N206, N38);
nand NAND4 (N208, N198, N207, N44, N40);
not NOT1 (N209, N28);
or OR4 (N210, N202, N19, N134, N201);
not NOT1 (N211, N175);
xor XOR2 (N212, N210, N150);
xor XOR2 (N213, N209, N180);
and AND2 (N214, N191, N86);
nor NOR3 (N215, N208, N141, N115);
and AND3 (N216, N212, N192, N9);
and AND3 (N217, N56, N44, N169);
nor NOR2 (N218, N199, N198);
nand NAND4 (N219, N203, N61, N113, N45);
and AND2 (N220, N217, N209);
not NOT1 (N221, N213);
not NOT1 (N222, N221);
buf BUF1 (N223, N218);
or OR4 (N224, N216, N102, N60, N74);
or OR3 (N225, N224, N119, N120);
buf BUF1 (N226, N225);
not NOT1 (N227, N226);
nand NAND4 (N228, N214, N134, N165, N1);
nor NOR3 (N229, N219, N88, N177);
and AND3 (N230, N220, N66, N89);
nand NAND3 (N231, N227, N78, N226);
and AND3 (N232, N211, N172, N10);
xor XOR2 (N233, N195, N210);
or OR2 (N234, N229, N147);
nand NAND3 (N235, N222, N61, N189);
and AND3 (N236, N205, N130, N146);
not NOT1 (N237, N236);
xor XOR2 (N238, N231, N228);
not NOT1 (N239, N116);
or OR3 (N240, N232, N109, N233);
nor NOR2 (N241, N83, N206);
nand NAND4 (N242, N241, N41, N192, N5);
nor NOR2 (N243, N223, N97);
and AND2 (N244, N239, N108);
xor XOR2 (N245, N237, N141);
or OR2 (N246, N234, N239);
xor XOR2 (N247, N235, N198);
or OR2 (N248, N245, N120);
and AND2 (N249, N240, N188);
not NOT1 (N250, N244);
and AND2 (N251, N243, N83);
nor NOR3 (N252, N249, N155, N206);
and AND4 (N253, N246, N113, N87, N204);
and AND2 (N254, N238, N6);
nor NOR2 (N255, N215, N112);
not NOT1 (N256, N254);
not NOT1 (N257, N253);
nand NAND3 (N258, N242, N17, N96);
nor NOR4 (N259, N258, N215, N245, N139);
or OR3 (N260, N250, N28, N2);
buf BUF1 (N261, N230);
buf BUF1 (N262, N251);
xor XOR2 (N263, N252, N109);
and AND2 (N264, N260, N132);
xor XOR2 (N265, N262, N94);
buf BUF1 (N266, N259);
nor NOR2 (N267, N257, N124);
or OR3 (N268, N265, N81, N161);
not NOT1 (N269, N268);
and AND2 (N270, N263, N224);
xor XOR2 (N271, N264, N21);
buf BUF1 (N272, N247);
or OR4 (N273, N267, N69, N260, N159);
nand NAND4 (N274, N270, N54, N201, N198);
nand NAND3 (N275, N256, N248, N251);
buf BUF1 (N276, N137);
not NOT1 (N277, N272);
or OR4 (N278, N269, N253, N238, N223);
nand NAND2 (N279, N275, N185);
xor XOR2 (N280, N277, N55);
nand NAND4 (N281, N266, N120, N121, N235);
or OR3 (N282, N255, N129, N139);
nand NAND4 (N283, N273, N34, N9, N135);
or OR2 (N284, N274, N192);
not NOT1 (N285, N284);
and AND4 (N286, N261, N95, N37, N106);
not NOT1 (N287, N286);
and AND3 (N288, N282, N206, N275);
and AND3 (N289, N288, N254, N229);
xor XOR2 (N290, N271, N89);
buf BUF1 (N291, N276);
buf BUF1 (N292, N283);
nor NOR2 (N293, N279, N260);
not NOT1 (N294, N291);
nand NAND3 (N295, N285, N105, N213);
xor XOR2 (N296, N293, N51);
not NOT1 (N297, N287);
nand NAND3 (N298, N296, N223, N280);
buf BUF1 (N299, N208);
not NOT1 (N300, N298);
not NOT1 (N301, N289);
and AND2 (N302, N290, N242);
not NOT1 (N303, N297);
nor NOR3 (N304, N301, N58, N59);
nand NAND4 (N305, N299, N4, N16, N13);
nor NOR3 (N306, N295, N299, N33);
and AND4 (N307, N281, N121, N241, N49);
nor NOR2 (N308, N303, N168);
buf BUF1 (N309, N307);
buf BUF1 (N310, N302);
nand NAND4 (N311, N309, N136, N79, N129);
or OR3 (N312, N292, N236, N6);
nor NOR4 (N313, N294, N181, N232, N197);
not NOT1 (N314, N312);
and AND2 (N315, N304, N160);
buf BUF1 (N316, N311);
nor NOR3 (N317, N314, N7, N216);
xor XOR2 (N318, N313, N60);
buf BUF1 (N319, N300);
not NOT1 (N320, N319);
or OR2 (N321, N305, N297);
nand NAND3 (N322, N320, N166, N34);
not NOT1 (N323, N306);
nand NAND4 (N324, N308, N277, N56, N204);
nor NOR3 (N325, N315, N119, N150);
not NOT1 (N326, N310);
and AND2 (N327, N324, N202);
and AND3 (N328, N317, N284, N28);
xor XOR2 (N329, N316, N23);
or OR2 (N330, N323, N182);
nor NOR2 (N331, N326, N234);
or OR2 (N332, N321, N238);
and AND4 (N333, N332, N60, N160, N243);
or OR4 (N334, N318, N325, N36, N196);
not NOT1 (N335, N133);
buf BUF1 (N336, N322);
nor NOR4 (N337, N336, N180, N27, N172);
not NOT1 (N338, N329);
buf BUF1 (N339, N327);
not NOT1 (N340, N333);
buf BUF1 (N341, N334);
not NOT1 (N342, N340);
buf BUF1 (N343, N328);
and AND4 (N344, N331, N46, N281, N66);
not NOT1 (N345, N342);
nand NAND4 (N346, N330, N230, N5, N60);
or OR3 (N347, N341, N313, N165);
buf BUF1 (N348, N335);
not NOT1 (N349, N346);
buf BUF1 (N350, N347);
nand NAND4 (N351, N339, N69, N248, N267);
xor XOR2 (N352, N337, N268);
and AND4 (N353, N348, N114, N206, N91);
nor NOR2 (N354, N345, N268);
and AND3 (N355, N354, N338, N114);
xor XOR2 (N356, N109, N64);
or OR2 (N357, N352, N147);
xor XOR2 (N358, N349, N275);
buf BUF1 (N359, N356);
xor XOR2 (N360, N358, N300);
xor XOR2 (N361, N355, N278);
nand NAND3 (N362, N185, N240, N165);
and AND4 (N363, N361, N79, N223, N353);
not NOT1 (N364, N162);
or OR2 (N365, N350, N36);
nor NOR4 (N366, N344, N169, N328, N363);
not NOT1 (N367, N281);
nand NAND4 (N368, N351, N15, N354, N52);
buf BUF1 (N369, N343);
not NOT1 (N370, N362);
not NOT1 (N371, N370);
nor NOR4 (N372, N369, N309, N154, N82);
xor XOR2 (N373, N364, N314);
and AND2 (N374, N371, N277);
nor NOR4 (N375, N374, N229, N349, N113);
nand NAND3 (N376, N373, N174, N247);
and AND3 (N377, N372, N326, N92);
nor NOR3 (N378, N357, N144, N181);
buf BUF1 (N379, N376);
nand NAND3 (N380, N359, N364, N266);
not NOT1 (N381, N379);
buf BUF1 (N382, N377);
xor XOR2 (N383, N366, N260);
not NOT1 (N384, N368);
not NOT1 (N385, N380);
xor XOR2 (N386, N383, N345);
not NOT1 (N387, N365);
not NOT1 (N388, N360);
buf BUF1 (N389, N378);
xor XOR2 (N390, N387, N388);
not NOT1 (N391, N50);
nand NAND4 (N392, N390, N73, N188, N124);
xor XOR2 (N393, N384, N375);
nand NAND4 (N394, N131, N78, N53, N138);
and AND4 (N395, N386, N325, N178, N227);
nor NOR3 (N396, N381, N119, N222);
xor XOR2 (N397, N395, N171);
nand NAND3 (N398, N391, N300, N218);
buf BUF1 (N399, N398);
nor NOR2 (N400, N396, N275);
and AND3 (N401, N382, N48, N52);
nor NOR2 (N402, N367, N24);
xor XOR2 (N403, N389, N267);
or OR2 (N404, N392, N74);
nand NAND3 (N405, N403, N237, N213);
buf BUF1 (N406, N400);
nand NAND2 (N407, N385, N195);
xor XOR2 (N408, N401, N334);
not NOT1 (N409, N407);
and AND2 (N410, N393, N44);
nor NOR3 (N411, N394, N62, N361);
and AND2 (N412, N406, N216);
xor XOR2 (N413, N410, N401);
buf BUF1 (N414, N404);
nor NOR2 (N415, N413, N97);
and AND3 (N416, N402, N337, N266);
or OR2 (N417, N405, N319);
xor XOR2 (N418, N408, N271);
and AND2 (N419, N416, N77);
and AND4 (N420, N411, N411, N221, N116);
xor XOR2 (N421, N420, N347);
nand NAND4 (N422, N414, N248, N373, N220);
nand NAND3 (N423, N415, N269, N289);
nor NOR4 (N424, N422, N89, N213, N359);
buf BUF1 (N425, N421);
or OR2 (N426, N424, N161);
nor NOR2 (N427, N397, N210);
and AND2 (N428, N419, N138);
not NOT1 (N429, N409);
and AND3 (N430, N427, N284, N201);
or OR3 (N431, N430, N303, N144);
nor NOR3 (N432, N425, N244, N324);
nor NOR2 (N433, N426, N181);
not NOT1 (N434, N412);
xor XOR2 (N435, N418, N237);
or OR4 (N436, N423, N384, N110, N36);
xor XOR2 (N437, N435, N8);
nand NAND2 (N438, N399, N318);
nor NOR4 (N439, N432, N436, N423, N195);
or OR4 (N440, N16, N88, N350, N39);
buf BUF1 (N441, N439);
or OR2 (N442, N434, N244);
buf BUF1 (N443, N437);
buf BUF1 (N444, N438);
and AND3 (N445, N431, N82, N185);
xor XOR2 (N446, N440, N434);
xor XOR2 (N447, N417, N28);
or OR2 (N448, N445, N400);
or OR2 (N449, N443, N317);
not NOT1 (N450, N447);
nand NAND2 (N451, N446, N319);
nor NOR4 (N452, N444, N255, N271, N15);
nand NAND2 (N453, N448, N325);
not NOT1 (N454, N452);
nand NAND4 (N455, N428, N117, N167, N370);
nand NAND4 (N456, N451, N50, N225, N262);
xor XOR2 (N457, N441, N118);
nand NAND4 (N458, N449, N71, N65, N164);
buf BUF1 (N459, N457);
buf BUF1 (N460, N454);
buf BUF1 (N461, N442);
nor NOR4 (N462, N459, N259, N430, N202);
nor NOR4 (N463, N462, N369, N321, N325);
xor XOR2 (N464, N456, N41);
not NOT1 (N465, N463);
nor NOR4 (N466, N429, N188, N303, N157);
nand NAND4 (N467, N461, N125, N184, N138);
and AND4 (N468, N450, N305, N204, N305);
xor XOR2 (N469, N458, N180);
nor NOR3 (N470, N468, N207, N313);
xor XOR2 (N471, N467, N168);
not NOT1 (N472, N470);
xor XOR2 (N473, N472, N229);
nor NOR4 (N474, N433, N168, N6, N348);
buf BUF1 (N475, N471);
nor NOR4 (N476, N465, N187, N4, N162);
nor NOR3 (N477, N473, N15, N214);
xor XOR2 (N478, N455, N19);
nor NOR3 (N479, N466, N191, N411);
buf BUF1 (N480, N475);
or OR2 (N481, N476, N266);
nand NAND3 (N482, N474, N245, N351);
nor NOR4 (N483, N479, N82, N191, N194);
and AND2 (N484, N460, N153);
not NOT1 (N485, N464);
and AND3 (N486, N453, N71, N242);
nor NOR4 (N487, N482, N350, N381, N173);
not NOT1 (N488, N483);
xor XOR2 (N489, N480, N207);
or OR2 (N490, N485, N203);
nor NOR4 (N491, N487, N374, N88, N442);
or OR2 (N492, N486, N426);
and AND2 (N493, N469, N359);
and AND2 (N494, N484, N112);
not NOT1 (N495, N491);
not NOT1 (N496, N490);
not NOT1 (N497, N494);
not NOT1 (N498, N477);
xor XOR2 (N499, N498, N393);
xor XOR2 (N500, N492, N94);
buf BUF1 (N501, N496);
xor XOR2 (N502, N478, N67);
buf BUF1 (N503, N495);
nor NOR2 (N504, N502, N87);
not NOT1 (N505, N488);
or OR2 (N506, N497, N387);
or OR4 (N507, N489, N175, N359, N41);
xor XOR2 (N508, N499, N130);
not NOT1 (N509, N506);
and AND2 (N510, N508, N274);
and AND3 (N511, N493, N300, N331);
or OR3 (N512, N500, N158, N2);
nand NAND3 (N513, N512, N199, N93);
buf BUF1 (N514, N509);
and AND2 (N515, N505, N509);
buf BUF1 (N516, N501);
and AND4 (N517, N510, N79, N4, N387);
nor NOR2 (N518, N517, N456);
not NOT1 (N519, N515);
or OR4 (N520, N481, N385, N2, N118);
and AND2 (N521, N511, N214);
nand NAND4 (N522, N516, N30, N6, N236);
nand NAND2 (N523, N522, N346);
nand NAND3 (N524, N513, N142, N412);
or OR2 (N525, N503, N188);
xor XOR2 (N526, N524, N383);
and AND4 (N527, N519, N196, N477, N318);
nand NAND2 (N528, N507, N26);
nand NAND4 (N529, N520, N353, N191, N408);
not NOT1 (N530, N518);
buf BUF1 (N531, N514);
and AND3 (N532, N525, N435, N258);
and AND2 (N533, N530, N520);
and AND3 (N534, N523, N482, N479);
nor NOR2 (N535, N534, N179);
and AND4 (N536, N533, N36, N207, N68);
and AND3 (N537, N529, N388, N65);
nand NAND3 (N538, N528, N102, N328);
buf BUF1 (N539, N538);
or OR3 (N540, N536, N463, N439);
or OR2 (N541, N540, N458);
and AND2 (N542, N541, N64);
and AND4 (N543, N531, N319, N217, N399);
and AND3 (N544, N532, N124, N41);
and AND2 (N545, N527, N310);
not NOT1 (N546, N526);
nor NOR4 (N547, N542, N467, N465, N116);
or OR4 (N548, N545, N67, N488, N166);
nor NOR3 (N549, N548, N363, N228);
or OR3 (N550, N549, N429, N448);
and AND4 (N551, N537, N476, N1, N284);
nor NOR3 (N552, N547, N228, N174);
nor NOR3 (N553, N521, N486, N150);
nor NOR4 (N554, N552, N297, N287, N445);
and AND3 (N555, N554, N44, N242);
nor NOR3 (N556, N539, N109, N523);
xor XOR2 (N557, N546, N340);
or OR2 (N558, N555, N196);
nor NOR4 (N559, N556, N336, N413, N330);
and AND2 (N560, N559, N141);
xor XOR2 (N561, N544, N494);
xor XOR2 (N562, N558, N156);
xor XOR2 (N563, N504, N17);
not NOT1 (N564, N543);
xor XOR2 (N565, N535, N294);
not NOT1 (N566, N562);
nor NOR2 (N567, N561, N544);
not NOT1 (N568, N565);
nor NOR2 (N569, N567, N197);
not NOT1 (N570, N551);
xor XOR2 (N571, N568, N176);
or OR2 (N572, N553, N531);
and AND2 (N573, N570, N269);
nor NOR3 (N574, N563, N66, N533);
and AND3 (N575, N569, N161, N230);
and AND3 (N576, N566, N249, N515);
buf BUF1 (N577, N564);
nand NAND2 (N578, N574, N522);
buf BUF1 (N579, N571);
and AND4 (N580, N577, N534, N34, N366);
xor XOR2 (N581, N580, N89);
xor XOR2 (N582, N557, N215);
and AND4 (N583, N575, N370, N440, N109);
buf BUF1 (N584, N572);
nor NOR2 (N585, N560, N230);
or OR4 (N586, N582, N565, N401, N482);
and AND4 (N587, N550, N173, N425, N296);
and AND2 (N588, N573, N388);
not NOT1 (N589, N579);
nand NAND3 (N590, N588, N416, N286);
and AND4 (N591, N583, N434, N201, N76);
nand NAND3 (N592, N581, N213, N394);
nor NOR4 (N593, N576, N451, N89, N141);
or OR3 (N594, N593, N333, N558);
or OR2 (N595, N585, N374);
not NOT1 (N596, N590);
buf BUF1 (N597, N594);
nand NAND4 (N598, N586, N323, N425, N233);
nor NOR4 (N599, N598, N583, N386, N254);
xor XOR2 (N600, N584, N337);
or OR4 (N601, N596, N304, N355, N249);
and AND3 (N602, N601, N184, N158);
nand NAND2 (N603, N595, N584);
nand NAND4 (N604, N600, N350, N417, N307);
buf BUF1 (N605, N589);
xor XOR2 (N606, N602, N388);
not NOT1 (N607, N605);
buf BUF1 (N608, N606);
buf BUF1 (N609, N587);
buf BUF1 (N610, N607);
buf BUF1 (N611, N608);
or OR2 (N612, N609, N371);
nand NAND4 (N613, N603, N358, N158, N150);
not NOT1 (N614, N592);
not NOT1 (N615, N611);
not NOT1 (N616, N615);
nor NOR2 (N617, N604, N308);
xor XOR2 (N618, N578, N164);
nor NOR3 (N619, N613, N381, N585);
or OR2 (N620, N612, N79);
nor NOR2 (N621, N617, N389);
nand NAND2 (N622, N616, N1);
or OR3 (N623, N597, N272, N333);
and AND4 (N624, N623, N599, N191, N122);
and AND2 (N625, N452, N56);
not NOT1 (N626, N620);
or OR2 (N627, N625, N262);
nor NOR4 (N628, N624, N299, N44, N368);
buf BUF1 (N629, N628);
not NOT1 (N630, N618);
buf BUF1 (N631, N619);
or OR2 (N632, N622, N129);
nor NOR2 (N633, N626, N551);
nand NAND3 (N634, N630, N464, N597);
buf BUF1 (N635, N634);
or OR4 (N636, N631, N520, N405, N336);
xor XOR2 (N637, N610, N253);
buf BUF1 (N638, N637);
not NOT1 (N639, N614);
not NOT1 (N640, N621);
nor NOR4 (N641, N633, N103, N364, N466);
xor XOR2 (N642, N632, N448);
not NOT1 (N643, N638);
buf BUF1 (N644, N642);
or OR4 (N645, N639, N586, N352, N445);
nand NAND3 (N646, N643, N492, N612);
xor XOR2 (N647, N591, N40);
not NOT1 (N648, N641);
and AND3 (N649, N648, N297, N629);
not NOT1 (N650, N405);
nor NOR4 (N651, N647, N440, N212, N351);
buf BUF1 (N652, N635);
or OR2 (N653, N645, N340);
or OR4 (N654, N640, N395, N503, N360);
not NOT1 (N655, N653);
nor NOR3 (N656, N644, N62, N529);
not NOT1 (N657, N650);
nand NAND4 (N658, N649, N126, N314, N212);
or OR3 (N659, N652, N48, N304);
and AND2 (N660, N658, N267);
nand NAND2 (N661, N656, N627);
and AND2 (N662, N63, N150);
buf BUF1 (N663, N646);
and AND2 (N664, N663, N631);
nand NAND3 (N665, N651, N402, N382);
nor NOR2 (N666, N664, N267);
nand NAND2 (N667, N654, N124);
buf BUF1 (N668, N660);
buf BUF1 (N669, N657);
xor XOR2 (N670, N661, N461);
nor NOR4 (N671, N666, N159, N520, N186);
not NOT1 (N672, N671);
nand NAND4 (N673, N670, N670, N152, N549);
or OR3 (N674, N669, N141, N85);
nand NAND2 (N675, N655, N196);
buf BUF1 (N676, N662);
not NOT1 (N677, N675);
and AND4 (N678, N659, N199, N200, N47);
nand NAND3 (N679, N668, N334, N534);
and AND2 (N680, N679, N47);
nand NAND3 (N681, N665, N31, N378);
and AND4 (N682, N667, N99, N677, N670);
buf BUF1 (N683, N655);
and AND3 (N684, N674, N413, N221);
not NOT1 (N685, N684);
nand NAND2 (N686, N636, N98);
nand NAND2 (N687, N686, N167);
nor NOR2 (N688, N676, N388);
xor XOR2 (N689, N687, N411);
xor XOR2 (N690, N683, N396);
or OR3 (N691, N678, N199, N56);
nor NOR4 (N692, N673, N227, N76, N33);
not NOT1 (N693, N682);
or OR3 (N694, N693, N33, N68);
or OR2 (N695, N688, N464);
not NOT1 (N696, N690);
nand NAND4 (N697, N691, N567, N223, N330);
and AND3 (N698, N680, N327, N240);
not NOT1 (N699, N696);
buf BUF1 (N700, N698);
buf BUF1 (N701, N692);
nand NAND4 (N702, N685, N380, N23, N521);
xor XOR2 (N703, N701, N380);
xor XOR2 (N704, N697, N330);
and AND2 (N705, N689, N544);
and AND4 (N706, N702, N423, N384, N20);
xor XOR2 (N707, N672, N274);
xor XOR2 (N708, N704, N351);
not NOT1 (N709, N707);
buf BUF1 (N710, N708);
and AND3 (N711, N703, N587, N614);
nor NOR3 (N712, N700, N453, N533);
buf BUF1 (N713, N705);
nor NOR4 (N714, N710, N647, N85, N467);
nor NOR3 (N715, N681, N610, N26);
nand NAND3 (N716, N712, N192, N421);
xor XOR2 (N717, N711, N253);
nor NOR4 (N718, N706, N96, N683, N105);
or OR2 (N719, N714, N223);
nor NOR4 (N720, N716, N426, N236, N303);
nand NAND3 (N721, N713, N450, N634);
xor XOR2 (N722, N717, N65);
and AND2 (N723, N721, N363);
not NOT1 (N724, N718);
nand NAND2 (N725, N694, N64);
buf BUF1 (N726, N725);
nor NOR4 (N727, N722, N489, N376, N605);
not NOT1 (N728, N726);
buf BUF1 (N729, N699);
nor NOR4 (N730, N695, N679, N147, N67);
nand NAND2 (N731, N720, N19);
not NOT1 (N732, N727);
and AND4 (N733, N731, N458, N634, N448);
not NOT1 (N734, N724);
xor XOR2 (N735, N729, N257);
nor NOR3 (N736, N733, N106, N20);
not NOT1 (N737, N715);
nor NOR2 (N738, N709, N331);
buf BUF1 (N739, N735);
buf BUF1 (N740, N738);
not NOT1 (N741, N737);
xor XOR2 (N742, N734, N239);
and AND2 (N743, N741, N333);
not NOT1 (N744, N723);
not NOT1 (N745, N730);
buf BUF1 (N746, N745);
nor NOR4 (N747, N742, N742, N693, N330);
not NOT1 (N748, N747);
or OR3 (N749, N732, N410, N319);
and AND2 (N750, N746, N536);
nand NAND2 (N751, N719, N213);
nor NOR2 (N752, N748, N436);
buf BUF1 (N753, N744);
not NOT1 (N754, N751);
not NOT1 (N755, N740);
or OR2 (N756, N754, N460);
nor NOR3 (N757, N736, N30, N4);
or OR4 (N758, N752, N649, N421, N652);
not NOT1 (N759, N739);
or OR2 (N760, N757, N319);
nor NOR2 (N761, N755, N398);
not NOT1 (N762, N750);
nand NAND3 (N763, N759, N392, N400);
and AND4 (N764, N763, N342, N607, N209);
nand NAND4 (N765, N756, N289, N396, N58);
not NOT1 (N766, N753);
xor XOR2 (N767, N761, N532);
or OR4 (N768, N760, N524, N521, N581);
nor NOR4 (N769, N749, N334, N602, N553);
xor XOR2 (N770, N728, N769);
or OR4 (N771, N243, N597, N614, N267);
not NOT1 (N772, N766);
or OR3 (N773, N762, N248, N249);
or OR4 (N774, N773, N419, N705, N682);
nand NAND3 (N775, N771, N314, N426);
and AND2 (N776, N765, N658);
nand NAND4 (N777, N767, N494, N130, N447);
nand NAND2 (N778, N764, N640);
nor NOR2 (N779, N775, N2);
or OR3 (N780, N774, N329, N548);
and AND2 (N781, N778, N466);
or OR2 (N782, N780, N40);
nor NOR2 (N783, N743, N585);
buf BUF1 (N784, N777);
not NOT1 (N785, N770);
buf BUF1 (N786, N785);
not NOT1 (N787, N783);
buf BUF1 (N788, N768);
nand NAND3 (N789, N788, N663, N6);
or OR2 (N790, N758, N124);
xor XOR2 (N791, N789, N658);
nor NOR3 (N792, N786, N167, N171);
nand NAND4 (N793, N792, N322, N682, N453);
buf BUF1 (N794, N779);
not NOT1 (N795, N782);
xor XOR2 (N796, N776, N339);
and AND4 (N797, N791, N33, N227, N659);
not NOT1 (N798, N790);
nor NOR3 (N799, N794, N39, N298);
and AND4 (N800, N772, N703, N309, N15);
and AND4 (N801, N787, N768, N442, N419);
nand NAND3 (N802, N793, N183, N42);
nor NOR3 (N803, N800, N734, N720);
not NOT1 (N804, N801);
or OR3 (N805, N781, N346, N400);
not NOT1 (N806, N795);
nor NOR2 (N807, N805, N739);
buf BUF1 (N808, N798);
nor NOR2 (N809, N797, N155);
not NOT1 (N810, N806);
not NOT1 (N811, N796);
xor XOR2 (N812, N809, N282);
buf BUF1 (N813, N804);
xor XOR2 (N814, N811, N597);
nor NOR4 (N815, N803, N11, N22, N258);
or OR4 (N816, N807, N28, N114, N677);
xor XOR2 (N817, N814, N633);
not NOT1 (N818, N799);
buf BUF1 (N819, N802);
and AND2 (N820, N816, N489);
buf BUF1 (N821, N819);
not NOT1 (N822, N813);
nand NAND3 (N823, N818, N637, N761);
xor XOR2 (N824, N823, N243);
and AND2 (N825, N824, N383);
xor XOR2 (N826, N784, N260);
and AND2 (N827, N817, N591);
nand NAND4 (N828, N810, N776, N124, N430);
not NOT1 (N829, N808);
nand NAND2 (N830, N812, N646);
nand NAND3 (N831, N829, N87, N296);
nand NAND2 (N832, N820, N369);
not NOT1 (N833, N826);
nand NAND4 (N834, N822, N144, N159, N728);
xor XOR2 (N835, N830, N543);
buf BUF1 (N836, N828);
not NOT1 (N837, N835);
or OR4 (N838, N836, N316, N597, N175);
not NOT1 (N839, N832);
nand NAND2 (N840, N838, N215);
nor NOR2 (N841, N825, N403);
nand NAND2 (N842, N840, N709);
xor XOR2 (N843, N821, N834);
and AND2 (N844, N577, N282);
nor NOR2 (N845, N843, N90);
nand NAND2 (N846, N845, N298);
xor XOR2 (N847, N833, N137);
and AND4 (N848, N847, N131, N32, N257);
xor XOR2 (N849, N839, N648);
nand NAND3 (N850, N844, N692, N529);
or OR2 (N851, N831, N376);
not NOT1 (N852, N848);
and AND3 (N853, N842, N8, N836);
buf BUF1 (N854, N841);
buf BUF1 (N855, N827);
xor XOR2 (N856, N837, N610);
and AND4 (N857, N854, N475, N178, N117);
and AND4 (N858, N852, N695, N835, N430);
nor NOR3 (N859, N851, N150, N88);
not NOT1 (N860, N846);
buf BUF1 (N861, N815);
nand NAND3 (N862, N858, N671, N853);
and AND2 (N863, N748, N42);
and AND4 (N864, N849, N852, N301, N714);
or OR3 (N865, N857, N505, N192);
buf BUF1 (N866, N862);
not NOT1 (N867, N856);
and AND2 (N868, N867, N640);
xor XOR2 (N869, N865, N174);
not NOT1 (N870, N869);
nand NAND2 (N871, N860, N8);
and AND4 (N872, N870, N116, N705, N730);
xor XOR2 (N873, N859, N345);
buf BUF1 (N874, N871);
xor XOR2 (N875, N874, N441);
xor XOR2 (N876, N866, N15);
and AND2 (N877, N861, N440);
nand NAND2 (N878, N872, N542);
not NOT1 (N879, N864);
not NOT1 (N880, N850);
nand NAND3 (N881, N875, N494, N263);
or OR3 (N882, N873, N654, N630);
buf BUF1 (N883, N881);
nor NOR4 (N884, N877, N439, N708, N690);
nor NOR4 (N885, N879, N847, N47, N766);
buf BUF1 (N886, N863);
not NOT1 (N887, N868);
xor XOR2 (N888, N885, N84);
and AND4 (N889, N888, N883, N850, N34);
nand NAND2 (N890, N10, N183);
buf BUF1 (N891, N890);
nor NOR2 (N892, N884, N159);
buf BUF1 (N893, N855);
nor NOR4 (N894, N889, N680, N853, N538);
not NOT1 (N895, N880);
nor NOR4 (N896, N876, N261, N219, N863);
not NOT1 (N897, N887);
nand NAND4 (N898, N893, N477, N329, N260);
and AND4 (N899, N897, N416, N4, N693);
or OR2 (N900, N891, N34);
or OR4 (N901, N882, N566, N342, N418);
or OR4 (N902, N878, N300, N250, N20);
not NOT1 (N903, N902);
nor NOR3 (N904, N899, N129, N379);
nor NOR3 (N905, N901, N760, N72);
not NOT1 (N906, N900);
buf BUF1 (N907, N894);
and AND4 (N908, N905, N895, N744, N836);
buf BUF1 (N909, N73);
nand NAND4 (N910, N903, N197, N832, N531);
not NOT1 (N911, N896);
nor NOR3 (N912, N898, N65, N733);
xor XOR2 (N913, N908, N890);
or OR4 (N914, N904, N282, N48, N905);
or OR2 (N915, N907, N119);
buf BUF1 (N916, N910);
or OR3 (N917, N911, N642, N523);
xor XOR2 (N918, N913, N175);
not NOT1 (N919, N917);
nor NOR3 (N920, N912, N249, N494);
xor XOR2 (N921, N919, N496);
or OR2 (N922, N921, N139);
nor NOR3 (N923, N909, N118, N27);
not NOT1 (N924, N914);
nand NAND4 (N925, N916, N389, N111, N784);
nor NOR4 (N926, N886, N823, N317, N2);
xor XOR2 (N927, N915, N106);
not NOT1 (N928, N920);
and AND4 (N929, N926, N255, N219, N20);
and AND3 (N930, N924, N273, N545);
nand NAND2 (N931, N923, N923);
xor XOR2 (N932, N906, N839);
xor XOR2 (N933, N932, N856);
not NOT1 (N934, N933);
and AND3 (N935, N934, N841, N718);
xor XOR2 (N936, N922, N671);
nand NAND4 (N937, N925, N335, N199, N478);
nor NOR4 (N938, N935, N585, N216, N189);
nand NAND4 (N939, N938, N875, N144, N207);
or OR4 (N940, N936, N825, N641, N262);
or OR2 (N941, N892, N37);
and AND4 (N942, N918, N20, N674, N306);
xor XOR2 (N943, N930, N5);
not NOT1 (N944, N939);
or OR4 (N945, N944, N262, N620, N726);
buf BUF1 (N946, N937);
nand NAND4 (N947, N931, N659, N130, N762);
xor XOR2 (N948, N946, N943);
nand NAND2 (N949, N438, N878);
or OR3 (N950, N945, N511, N188);
or OR4 (N951, N947, N596, N26, N663);
or OR4 (N952, N941, N829, N233, N504);
xor XOR2 (N953, N940, N224);
nor NOR2 (N954, N928, N387);
not NOT1 (N955, N927);
buf BUF1 (N956, N954);
not NOT1 (N957, N956);
nor NOR4 (N958, N950, N110, N858, N312);
not NOT1 (N959, N951);
not NOT1 (N960, N955);
buf BUF1 (N961, N949);
not NOT1 (N962, N960);
and AND3 (N963, N952, N838, N348);
and AND4 (N964, N948, N491, N471, N293);
nor NOR4 (N965, N959, N468, N683, N480);
nand NAND3 (N966, N965, N857, N572);
and AND2 (N967, N958, N427);
buf BUF1 (N968, N953);
buf BUF1 (N969, N962);
nand NAND2 (N970, N968, N537);
and AND3 (N971, N963, N155, N759);
and AND2 (N972, N961, N316);
xor XOR2 (N973, N942, N359);
buf BUF1 (N974, N969);
xor XOR2 (N975, N972, N478);
or OR2 (N976, N966, N353);
nor NOR3 (N977, N967, N138, N238);
buf BUF1 (N978, N964);
not NOT1 (N979, N971);
buf BUF1 (N980, N973);
and AND4 (N981, N970, N584, N384, N804);
not NOT1 (N982, N979);
nor NOR2 (N983, N980, N403);
xor XOR2 (N984, N978, N774);
not NOT1 (N985, N982);
nor NOR3 (N986, N981, N91, N134);
or OR3 (N987, N976, N471, N735);
not NOT1 (N988, N957);
not NOT1 (N989, N986);
buf BUF1 (N990, N977);
nand NAND2 (N991, N974, N325);
and AND2 (N992, N989, N383);
xor XOR2 (N993, N985, N361);
and AND3 (N994, N987, N277, N202);
and AND2 (N995, N975, N145);
buf BUF1 (N996, N984);
or OR4 (N997, N994, N79, N685, N369);
and AND3 (N998, N991, N622, N932);
nand NAND4 (N999, N929, N628, N444, N291);
buf BUF1 (N1000, N992);
and AND2 (N1001, N993, N209);
not NOT1 (N1002, N983);
nor NOR3 (N1003, N1000, N21, N173);
or OR3 (N1004, N988, N137, N282);
nand NAND4 (N1005, N999, N213, N788, N542);
or OR3 (N1006, N998, N114, N331);
or OR2 (N1007, N1001, N265);
buf BUF1 (N1008, N1005);
buf BUF1 (N1009, N1002);
nor NOR4 (N1010, N995, N476, N240, N761);
nor NOR4 (N1011, N1007, N64, N550, N754);
not NOT1 (N1012, N1010);
buf BUF1 (N1013, N996);
xor XOR2 (N1014, N1009, N855);
buf BUF1 (N1015, N1003);
xor XOR2 (N1016, N1014, N836);
nor NOR2 (N1017, N1011, N49);
not NOT1 (N1018, N1012);
nand NAND4 (N1019, N990, N173, N514, N50);
nor NOR2 (N1020, N1006, N506);
xor XOR2 (N1021, N1016, N847);
xor XOR2 (N1022, N1013, N709);
nor NOR2 (N1023, N1015, N385);
nand NAND2 (N1024, N1018, N538);
nand NAND2 (N1025, N1023, N416);
nand NAND3 (N1026, N997, N21, N452);
nand NAND2 (N1027, N1004, N398);
buf BUF1 (N1028, N1022);
nor NOR2 (N1029, N1027, N842);
nand NAND3 (N1030, N1026, N170, N504);
nand NAND3 (N1031, N1021, N809, N157);
and AND3 (N1032, N1025, N655, N387);
xor XOR2 (N1033, N1030, N110);
or OR3 (N1034, N1019, N609, N398);
or OR3 (N1035, N1008, N148, N320);
nor NOR2 (N1036, N1032, N339);
not NOT1 (N1037, N1033);
not NOT1 (N1038, N1024);
nor NOR3 (N1039, N1020, N963, N69);
nand NAND3 (N1040, N1017, N333, N215);
nand NAND4 (N1041, N1035, N603, N68, N105);
nor NOR2 (N1042, N1028, N279);
not NOT1 (N1043, N1029);
xor XOR2 (N1044, N1042, N406);
nand NAND4 (N1045, N1039, N277, N420, N939);
xor XOR2 (N1046, N1040, N281);
nand NAND2 (N1047, N1041, N340);
or OR2 (N1048, N1047, N1005);
buf BUF1 (N1049, N1045);
buf BUF1 (N1050, N1034);
or OR4 (N1051, N1037, N790, N722, N582);
nand NAND4 (N1052, N1044, N128, N500, N213);
xor XOR2 (N1053, N1050, N907);
buf BUF1 (N1054, N1038);
xor XOR2 (N1055, N1049, N18);
nand NAND3 (N1056, N1055, N687, N320);
buf BUF1 (N1057, N1031);
nor NOR4 (N1058, N1056, N188, N707, N419);
or OR2 (N1059, N1052, N422);
not NOT1 (N1060, N1057);
or OR3 (N1061, N1058, N558, N65);
xor XOR2 (N1062, N1054, N1035);
buf BUF1 (N1063, N1043);
or OR3 (N1064, N1036, N769, N239);
not NOT1 (N1065, N1046);
xor XOR2 (N1066, N1062, N398);
not NOT1 (N1067, N1063);
and AND4 (N1068, N1048, N387, N963, N1034);
or OR3 (N1069, N1061, N877, N900);
not NOT1 (N1070, N1051);
not NOT1 (N1071, N1067);
or OR2 (N1072, N1053, N857);
nand NAND3 (N1073, N1066, N406, N185);
nand NAND3 (N1074, N1059, N723, N38);
nand NAND2 (N1075, N1072, N516);
and AND3 (N1076, N1071, N610, N959);
or OR2 (N1077, N1064, N382);
xor XOR2 (N1078, N1074, N893);
nor NOR4 (N1079, N1077, N829, N340, N410);
and AND2 (N1080, N1075, N16);
buf BUF1 (N1081, N1060);
nand NAND4 (N1082, N1078, N668, N449, N356);
and AND4 (N1083, N1069, N101, N98, N599);
and AND3 (N1084, N1082, N828, N597);
buf BUF1 (N1085, N1068);
or OR2 (N1086, N1081, N176);
or OR3 (N1087, N1079, N572, N197);
or OR2 (N1088, N1070, N594);
xor XOR2 (N1089, N1080, N785);
xor XOR2 (N1090, N1089, N668);
nand NAND3 (N1091, N1076, N469, N512);
nor NOR2 (N1092, N1085, N837);
nor NOR2 (N1093, N1090, N101);
nand NAND4 (N1094, N1092, N913, N898, N285);
nor NOR3 (N1095, N1086, N206, N311);
and AND2 (N1096, N1073, N63);
and AND3 (N1097, N1094, N553, N871);
and AND3 (N1098, N1084, N949, N45);
nor NOR2 (N1099, N1097, N339);
xor XOR2 (N1100, N1093, N505);
nor NOR3 (N1101, N1088, N344, N948);
and AND3 (N1102, N1099, N1054, N961);
nor NOR3 (N1103, N1065, N1007, N86);
nand NAND2 (N1104, N1100, N389);
nor NOR4 (N1105, N1083, N256, N564, N118);
nand NAND4 (N1106, N1098, N871, N738, N1045);
nand NAND3 (N1107, N1106, N588, N409);
nand NAND4 (N1108, N1103, N1095, N953, N193);
and AND4 (N1109, N525, N65, N471, N1043);
buf BUF1 (N1110, N1091);
and AND4 (N1111, N1109, N755, N1037, N341);
not NOT1 (N1112, N1108);
buf BUF1 (N1113, N1111);
xor XOR2 (N1114, N1102, N921);
and AND4 (N1115, N1096, N794, N987, N335);
buf BUF1 (N1116, N1114);
not NOT1 (N1117, N1113);
and AND4 (N1118, N1087, N1106, N807, N736);
nand NAND2 (N1119, N1104, N263);
not NOT1 (N1120, N1119);
nand NAND3 (N1121, N1120, N445, N515);
and AND3 (N1122, N1116, N814, N430);
not NOT1 (N1123, N1121);
xor XOR2 (N1124, N1112, N25);
nand NAND4 (N1125, N1101, N70, N314, N994);
xor XOR2 (N1126, N1118, N806);
xor XOR2 (N1127, N1122, N857);
xor XOR2 (N1128, N1123, N228);
xor XOR2 (N1129, N1125, N1006);
and AND3 (N1130, N1124, N724, N810);
not NOT1 (N1131, N1115);
xor XOR2 (N1132, N1131, N921);
nand NAND2 (N1133, N1110, N128);
xor XOR2 (N1134, N1128, N613);
not NOT1 (N1135, N1126);
nor NOR2 (N1136, N1134, N448);
xor XOR2 (N1137, N1129, N802);
nand NAND4 (N1138, N1130, N1098, N624, N834);
nor NOR4 (N1139, N1135, N726, N214, N677);
nor NOR3 (N1140, N1132, N917, N812);
xor XOR2 (N1141, N1137, N396);
and AND3 (N1142, N1105, N603, N70);
or OR3 (N1143, N1138, N897, N90);
and AND2 (N1144, N1141, N593);
and AND4 (N1145, N1117, N483, N602, N804);
nand NAND3 (N1146, N1136, N945, N431);
or OR2 (N1147, N1127, N378);
or OR2 (N1148, N1139, N39);
and AND2 (N1149, N1143, N443);
not NOT1 (N1150, N1142);
nor NOR2 (N1151, N1147, N939);
not NOT1 (N1152, N1149);
xor XOR2 (N1153, N1148, N693);
xor XOR2 (N1154, N1144, N447);
buf BUF1 (N1155, N1145);
and AND4 (N1156, N1153, N721, N526, N512);
not NOT1 (N1157, N1154);
xor XOR2 (N1158, N1155, N495);
and AND2 (N1159, N1157, N365);
buf BUF1 (N1160, N1146);
nor NOR3 (N1161, N1156, N1039, N404);
or OR2 (N1162, N1150, N1013);
not NOT1 (N1163, N1133);
and AND3 (N1164, N1140, N767, N354);
not NOT1 (N1165, N1152);
xor XOR2 (N1166, N1161, N175);
or OR4 (N1167, N1107, N488, N981, N422);
nor NOR4 (N1168, N1166, N466, N621, N475);
xor XOR2 (N1169, N1163, N1133);
and AND4 (N1170, N1169, N668, N242, N154);
nor NOR4 (N1171, N1165, N623, N1, N747);
nand NAND2 (N1172, N1162, N216);
nor NOR2 (N1173, N1159, N998);
xor XOR2 (N1174, N1160, N178);
or OR2 (N1175, N1167, N1079);
nand NAND3 (N1176, N1164, N588, N263);
buf BUF1 (N1177, N1171);
xor XOR2 (N1178, N1170, N750);
and AND2 (N1179, N1158, N791);
nand NAND4 (N1180, N1177, N913, N183, N227);
or OR2 (N1181, N1168, N180);
and AND4 (N1182, N1172, N244, N466, N929);
xor XOR2 (N1183, N1175, N969);
xor XOR2 (N1184, N1173, N751);
buf BUF1 (N1185, N1178);
not NOT1 (N1186, N1179);
or OR2 (N1187, N1181, N463);
nor NOR4 (N1188, N1187, N137, N773, N1034);
and AND4 (N1189, N1174, N138, N431, N970);
not NOT1 (N1190, N1183);
not NOT1 (N1191, N1189);
and AND2 (N1192, N1190, N318);
nand NAND3 (N1193, N1176, N585, N1143);
nor NOR2 (N1194, N1188, N398);
buf BUF1 (N1195, N1192);
nor NOR3 (N1196, N1180, N517, N524);
and AND2 (N1197, N1184, N665);
buf BUF1 (N1198, N1194);
and AND3 (N1199, N1151, N442, N817);
buf BUF1 (N1200, N1186);
and AND2 (N1201, N1185, N839);
buf BUF1 (N1202, N1195);
not NOT1 (N1203, N1182);
and AND3 (N1204, N1201, N391, N963);
buf BUF1 (N1205, N1196);
nor NOR4 (N1206, N1202, N410, N1057, N1180);
nand NAND2 (N1207, N1206, N1102);
nand NAND2 (N1208, N1198, N471);
or OR4 (N1209, N1203, N717, N488, N675);
or OR3 (N1210, N1204, N189, N670);
not NOT1 (N1211, N1191);
nand NAND4 (N1212, N1205, N698, N994, N836);
nor NOR4 (N1213, N1208, N63, N265, N516);
nor NOR2 (N1214, N1213, N1156);
buf BUF1 (N1215, N1212);
nor NOR2 (N1216, N1214, N167);
buf BUF1 (N1217, N1199);
xor XOR2 (N1218, N1217, N978);
nand NAND4 (N1219, N1209, N1066, N992, N398);
or OR3 (N1220, N1200, N74, N732);
buf BUF1 (N1221, N1207);
nand NAND2 (N1222, N1197, N900);
buf BUF1 (N1223, N1210);
nand NAND4 (N1224, N1222, N1117, N1084, N410);
xor XOR2 (N1225, N1219, N155);
buf BUF1 (N1226, N1193);
not NOT1 (N1227, N1220);
nand NAND2 (N1228, N1224, N964);
nand NAND2 (N1229, N1227, N437);
not NOT1 (N1230, N1221);
or OR2 (N1231, N1211, N235);
and AND2 (N1232, N1215, N285);
xor XOR2 (N1233, N1231, N784);
not NOT1 (N1234, N1225);
buf BUF1 (N1235, N1233);
buf BUF1 (N1236, N1228);
and AND3 (N1237, N1232, N974, N239);
xor XOR2 (N1238, N1226, N122);
nor NOR2 (N1239, N1229, N411);
or OR3 (N1240, N1216, N1013, N54);
not NOT1 (N1241, N1237);
and AND4 (N1242, N1238, N326, N866, N374);
xor XOR2 (N1243, N1218, N881);
xor XOR2 (N1244, N1239, N850);
nand NAND2 (N1245, N1230, N396);
nor NOR4 (N1246, N1240, N1012, N306, N1088);
and AND2 (N1247, N1242, N669);
not NOT1 (N1248, N1223);
or OR4 (N1249, N1234, N180, N41, N55);
not NOT1 (N1250, N1244);
buf BUF1 (N1251, N1247);
buf BUF1 (N1252, N1246);
buf BUF1 (N1253, N1235);
nand NAND2 (N1254, N1251, N231);
nor NOR2 (N1255, N1236, N1050);
nor NOR3 (N1256, N1245, N238, N328);
or OR3 (N1257, N1241, N629, N469);
buf BUF1 (N1258, N1254);
nor NOR2 (N1259, N1249, N906);
nor NOR3 (N1260, N1259, N1228, N651);
nand NAND3 (N1261, N1248, N1041, N333);
not NOT1 (N1262, N1260);
or OR2 (N1263, N1255, N34);
or OR2 (N1264, N1256, N1117);
or OR4 (N1265, N1261, N30, N607, N223);
not NOT1 (N1266, N1262);
and AND4 (N1267, N1266, N1103, N1139, N9);
or OR3 (N1268, N1253, N830, N130);
nand NAND2 (N1269, N1252, N593);
buf BUF1 (N1270, N1263);
and AND4 (N1271, N1250, N624, N951, N1210);
not NOT1 (N1272, N1243);
xor XOR2 (N1273, N1265, N24);
not NOT1 (N1274, N1264);
nand NAND2 (N1275, N1258, N979);
buf BUF1 (N1276, N1257);
and AND3 (N1277, N1268, N1276, N1276);
or OR3 (N1278, N523, N367, N393);
xor XOR2 (N1279, N1274, N241);
and AND4 (N1280, N1269, N195, N105, N188);
xor XOR2 (N1281, N1278, N1280);
not NOT1 (N1282, N108);
buf BUF1 (N1283, N1277);
and AND4 (N1284, N1275, N1113, N1200, N1188);
xor XOR2 (N1285, N1279, N224);
xor XOR2 (N1286, N1282, N935);
buf BUF1 (N1287, N1284);
buf BUF1 (N1288, N1287);
buf BUF1 (N1289, N1272);
buf BUF1 (N1290, N1283);
and AND3 (N1291, N1286, N775, N526);
xor XOR2 (N1292, N1291, N230);
xor XOR2 (N1293, N1273, N623);
or OR3 (N1294, N1271, N1208, N984);
xor XOR2 (N1295, N1267, N443);
or OR2 (N1296, N1293, N797);
or OR3 (N1297, N1296, N442, N345);
not NOT1 (N1298, N1294);
not NOT1 (N1299, N1281);
nand NAND4 (N1300, N1288, N1206, N1019, N962);
not NOT1 (N1301, N1292);
buf BUF1 (N1302, N1300);
or OR4 (N1303, N1285, N947, N1063, N458);
not NOT1 (N1304, N1299);
or OR4 (N1305, N1290, N507, N1020, N330);
not NOT1 (N1306, N1304);
nor NOR2 (N1307, N1298, N677);
xor XOR2 (N1308, N1301, N724);
nand NAND4 (N1309, N1308, N213, N976, N799);
nand NAND3 (N1310, N1302, N801, N1186);
nor NOR4 (N1311, N1306, N202, N640, N1035);
nand NAND3 (N1312, N1297, N1049, N777);
and AND4 (N1313, N1270, N947, N1133, N928);
and AND2 (N1314, N1305, N271);
and AND4 (N1315, N1310, N1206, N1177, N253);
or OR3 (N1316, N1309, N992, N383);
or OR2 (N1317, N1311, N251);
xor XOR2 (N1318, N1312, N1113);
nor NOR4 (N1319, N1307, N601, N479, N1276);
or OR2 (N1320, N1303, N1062);
nor NOR3 (N1321, N1313, N110, N645);
not NOT1 (N1322, N1289);
xor XOR2 (N1323, N1314, N688);
buf BUF1 (N1324, N1323);
not NOT1 (N1325, N1316);
xor XOR2 (N1326, N1318, N1286);
or OR2 (N1327, N1321, N338);
or OR2 (N1328, N1322, N1117);
not NOT1 (N1329, N1320);
not NOT1 (N1330, N1325);
xor XOR2 (N1331, N1319, N865);
buf BUF1 (N1332, N1326);
not NOT1 (N1333, N1331);
and AND3 (N1334, N1295, N978, N1288);
nor NOR2 (N1335, N1333, N55);
and AND3 (N1336, N1324, N255, N1061);
not NOT1 (N1337, N1334);
buf BUF1 (N1338, N1329);
xor XOR2 (N1339, N1315, N539);
not NOT1 (N1340, N1328);
xor XOR2 (N1341, N1335, N1128);
buf BUF1 (N1342, N1337);
nor NOR2 (N1343, N1340, N144);
nand NAND3 (N1344, N1327, N82, N923);
nor NOR3 (N1345, N1338, N401, N1062);
nand NAND3 (N1346, N1345, N801, N1305);
xor XOR2 (N1347, N1343, N1221);
and AND3 (N1348, N1332, N1267, N621);
not NOT1 (N1349, N1317);
and AND4 (N1350, N1330, N1291, N1050, N374);
not NOT1 (N1351, N1339);
or OR2 (N1352, N1350, N1305);
buf BUF1 (N1353, N1347);
nor NOR4 (N1354, N1353, N1129, N1010, N1297);
not NOT1 (N1355, N1344);
and AND4 (N1356, N1354, N1329, N323, N903);
and AND3 (N1357, N1342, N265, N302);
buf BUF1 (N1358, N1349);
and AND4 (N1359, N1351, N644, N368, N1259);
buf BUF1 (N1360, N1357);
nand NAND4 (N1361, N1352, N1153, N480, N784);
nand NAND3 (N1362, N1359, N874, N705);
and AND2 (N1363, N1348, N608);
xor XOR2 (N1364, N1362, N246);
nor NOR2 (N1365, N1364, N335);
buf BUF1 (N1366, N1341);
nand NAND3 (N1367, N1366, N35, N654);
xor XOR2 (N1368, N1360, N1006);
or OR4 (N1369, N1346, N383, N613, N1360);
xor XOR2 (N1370, N1361, N843);
not NOT1 (N1371, N1336);
nand NAND2 (N1372, N1363, N271);
nand NAND4 (N1373, N1365, N611, N1103, N1127);
nor NOR2 (N1374, N1358, N763);
xor XOR2 (N1375, N1367, N696);
and AND4 (N1376, N1372, N289, N590, N1036);
not NOT1 (N1377, N1356);
or OR3 (N1378, N1376, N340, N551);
and AND3 (N1379, N1368, N604, N862);
not NOT1 (N1380, N1377);
xor XOR2 (N1381, N1374, N1115);
and AND3 (N1382, N1375, N685, N1349);
or OR2 (N1383, N1382, N197);
or OR4 (N1384, N1381, N926, N880, N854);
or OR4 (N1385, N1373, N369, N1218, N561);
xor XOR2 (N1386, N1384, N630);
or OR4 (N1387, N1369, N1095, N189, N688);
or OR2 (N1388, N1385, N263);
or OR2 (N1389, N1386, N682);
buf BUF1 (N1390, N1378);
or OR3 (N1391, N1390, N293, N1303);
and AND2 (N1392, N1388, N1390);
buf BUF1 (N1393, N1391);
xor XOR2 (N1394, N1370, N1338);
not NOT1 (N1395, N1371);
not NOT1 (N1396, N1392);
xor XOR2 (N1397, N1387, N606);
not NOT1 (N1398, N1395);
nand NAND2 (N1399, N1396, N464);
nor NOR2 (N1400, N1394, N1115);
or OR4 (N1401, N1380, N1087, N600, N822);
nor NOR4 (N1402, N1397, N464, N647, N482);
or OR2 (N1403, N1398, N668);
not NOT1 (N1404, N1383);
buf BUF1 (N1405, N1401);
nor NOR3 (N1406, N1399, N9, N916);
not NOT1 (N1407, N1402);
and AND4 (N1408, N1404, N453, N1182, N187);
or OR4 (N1409, N1406, N1009, N993, N295);
buf BUF1 (N1410, N1407);
or OR3 (N1411, N1409, N111, N24);
buf BUF1 (N1412, N1355);
buf BUF1 (N1413, N1408);
xor XOR2 (N1414, N1412, N881);
or OR2 (N1415, N1400, N33);
or OR2 (N1416, N1379, N1249);
xor XOR2 (N1417, N1413, N139);
xor XOR2 (N1418, N1411, N614);
or OR4 (N1419, N1416, N320, N630, N45);
not NOT1 (N1420, N1415);
buf BUF1 (N1421, N1403);
nor NOR3 (N1422, N1417, N729, N1037);
or OR2 (N1423, N1393, N731);
not NOT1 (N1424, N1421);
and AND4 (N1425, N1423, N911, N645, N833);
and AND3 (N1426, N1420, N418, N1414);
or OR3 (N1427, N244, N507, N92);
nand NAND4 (N1428, N1419, N1232, N214, N890);
or OR3 (N1429, N1389, N406, N1119);
and AND3 (N1430, N1426, N504, N592);
not NOT1 (N1431, N1424);
buf BUF1 (N1432, N1410);
nand NAND3 (N1433, N1431, N202, N580);
nand NAND2 (N1434, N1422, N1172);
nand NAND4 (N1435, N1428, N485, N258, N611);
or OR4 (N1436, N1418, N1207, N941, N797);
or OR4 (N1437, N1434, N1358, N1333, N459);
buf BUF1 (N1438, N1437);
xor XOR2 (N1439, N1405, N1333);
buf BUF1 (N1440, N1430);
nand NAND4 (N1441, N1433, N138, N569, N1058);
buf BUF1 (N1442, N1429);
xor XOR2 (N1443, N1435, N818);
buf BUF1 (N1444, N1432);
nand NAND4 (N1445, N1440, N251, N325, N545);
or OR3 (N1446, N1438, N1306, N144);
or OR3 (N1447, N1425, N1342, N102);
not NOT1 (N1448, N1442);
not NOT1 (N1449, N1436);
not NOT1 (N1450, N1448);
nand NAND2 (N1451, N1447, N296);
buf BUF1 (N1452, N1441);
xor XOR2 (N1453, N1445, N480);
and AND3 (N1454, N1446, N461, N798);
and AND2 (N1455, N1427, N699);
or OR2 (N1456, N1454, N1313);
xor XOR2 (N1457, N1449, N69);
buf BUF1 (N1458, N1453);
buf BUF1 (N1459, N1444);
xor XOR2 (N1460, N1452, N1446);
and AND2 (N1461, N1457, N1176);
xor XOR2 (N1462, N1451, N1313);
or OR4 (N1463, N1462, N978, N242, N1175);
buf BUF1 (N1464, N1459);
or OR3 (N1465, N1443, N906, N1128);
xor XOR2 (N1466, N1464, N411);
not NOT1 (N1467, N1439);
nand NAND3 (N1468, N1463, N3, N296);
buf BUF1 (N1469, N1458);
nor NOR4 (N1470, N1466, N1003, N1455, N299);
xor XOR2 (N1471, N502, N874);
nor NOR4 (N1472, N1469, N150, N459, N16);
xor XOR2 (N1473, N1460, N761);
xor XOR2 (N1474, N1467, N171);
or OR4 (N1475, N1472, N1399, N282, N366);
nor NOR4 (N1476, N1471, N676, N1121, N1044);
not NOT1 (N1477, N1475);
buf BUF1 (N1478, N1474);
and AND4 (N1479, N1478, N1120, N67, N454);
nor NOR2 (N1480, N1468, N909);
nor NOR4 (N1481, N1476, N248, N1185, N1044);
xor XOR2 (N1482, N1461, N52);
nand NAND3 (N1483, N1465, N109, N1432);
not NOT1 (N1484, N1470);
or OR2 (N1485, N1450, N1227);
nand NAND3 (N1486, N1482, N839, N1029);
xor XOR2 (N1487, N1456, N1028);
nor NOR3 (N1488, N1486, N707, N504);
nor NOR3 (N1489, N1479, N76, N644);
and AND4 (N1490, N1485, N909, N604, N323);
buf BUF1 (N1491, N1483);
not NOT1 (N1492, N1480);
xor XOR2 (N1493, N1491, N1403);
nor NOR3 (N1494, N1489, N46, N751);
and AND2 (N1495, N1492, N219);
buf BUF1 (N1496, N1487);
nand NAND4 (N1497, N1473, N1455, N856, N264);
buf BUF1 (N1498, N1484);
buf BUF1 (N1499, N1498);
xor XOR2 (N1500, N1493, N1383);
or OR3 (N1501, N1477, N1425, N872);
not NOT1 (N1502, N1501);
and AND2 (N1503, N1496, N1150);
or OR3 (N1504, N1494, N392, N1220);
xor XOR2 (N1505, N1500, N318);
and AND2 (N1506, N1502, N1040);
nor NOR3 (N1507, N1506, N767, N254);
nor NOR3 (N1508, N1488, N234, N1395);
xor XOR2 (N1509, N1504, N1318);
not NOT1 (N1510, N1507);
nand NAND2 (N1511, N1505, N944);
buf BUF1 (N1512, N1497);
xor XOR2 (N1513, N1499, N1474);
or OR2 (N1514, N1510, N1484);
buf BUF1 (N1515, N1512);
buf BUF1 (N1516, N1503);
nor NOR2 (N1517, N1511, N295);
buf BUF1 (N1518, N1508);
nor NOR2 (N1519, N1495, N442);
nor NOR3 (N1520, N1515, N862, N636);
xor XOR2 (N1521, N1509, N189);
nor NOR4 (N1522, N1518, N411, N1340, N1287);
not NOT1 (N1523, N1490);
nor NOR4 (N1524, N1516, N617, N1332, N1427);
nor NOR3 (N1525, N1513, N39, N775);
xor XOR2 (N1526, N1524, N368);
not NOT1 (N1527, N1519);
or OR3 (N1528, N1526, N15, N1139);
buf BUF1 (N1529, N1481);
xor XOR2 (N1530, N1527, N1229);
and AND2 (N1531, N1530, N773);
and AND2 (N1532, N1531, N3);
xor XOR2 (N1533, N1529, N707);
xor XOR2 (N1534, N1520, N434);
nor NOR4 (N1535, N1517, N185, N1258, N1278);
nor NOR4 (N1536, N1525, N82, N508, N859);
and AND2 (N1537, N1534, N530);
nor NOR2 (N1538, N1537, N1145);
xor XOR2 (N1539, N1522, N909);
buf BUF1 (N1540, N1528);
or OR2 (N1541, N1523, N288);
or OR3 (N1542, N1514, N1261, N1512);
nand NAND3 (N1543, N1521, N283, N1016);
not NOT1 (N1544, N1542);
nand NAND4 (N1545, N1544, N552, N242, N943);
nand NAND4 (N1546, N1539, N1429, N476, N1103);
not NOT1 (N1547, N1538);
buf BUF1 (N1548, N1532);
and AND2 (N1549, N1548, N209);
buf BUF1 (N1550, N1535);
and AND2 (N1551, N1543, N514);
or OR2 (N1552, N1545, N636);
nand NAND2 (N1553, N1550, N991);
or OR3 (N1554, N1549, N1202, N531);
nand NAND2 (N1555, N1536, N1418);
not NOT1 (N1556, N1540);
buf BUF1 (N1557, N1546);
xor XOR2 (N1558, N1556, N990);
or OR2 (N1559, N1533, N1388);
and AND4 (N1560, N1555, N1369, N1461, N1248);
buf BUF1 (N1561, N1547);
not NOT1 (N1562, N1553);
or OR3 (N1563, N1551, N584, N1138);
xor XOR2 (N1564, N1554, N168);
xor XOR2 (N1565, N1560, N1412);
xor XOR2 (N1566, N1565, N1041);
or OR2 (N1567, N1564, N638);
nand NAND4 (N1568, N1562, N1356, N739, N1492);
xor XOR2 (N1569, N1568, N915);
not NOT1 (N1570, N1541);
xor XOR2 (N1571, N1569, N57);
xor XOR2 (N1572, N1566, N1414);
nand NAND3 (N1573, N1561, N764, N1185);
or OR3 (N1574, N1563, N631, N1352);
nor NOR4 (N1575, N1558, N285, N1324, N1519);
xor XOR2 (N1576, N1559, N1045);
and AND4 (N1577, N1574, N40, N1185, N1265);
buf BUF1 (N1578, N1576);
or OR3 (N1579, N1557, N1236, N799);
not NOT1 (N1580, N1570);
buf BUF1 (N1581, N1580);
or OR4 (N1582, N1567, N1384, N705, N669);
buf BUF1 (N1583, N1581);
nor NOR4 (N1584, N1572, N1133, N1335, N557);
nand NAND3 (N1585, N1571, N1364, N1244);
and AND3 (N1586, N1583, N619, N775);
and AND3 (N1587, N1584, N275, N8);
nand NAND4 (N1588, N1586, N730, N1380, N1057);
xor XOR2 (N1589, N1587, N1042);
not NOT1 (N1590, N1552);
nor NOR2 (N1591, N1575, N1539);
and AND3 (N1592, N1590, N554, N1141);
and AND3 (N1593, N1589, N735, N1320);
buf BUF1 (N1594, N1579);
not NOT1 (N1595, N1588);
nor NOR4 (N1596, N1592, N638, N640, N465);
not NOT1 (N1597, N1591);
or OR2 (N1598, N1597, N599);
buf BUF1 (N1599, N1596);
nand NAND4 (N1600, N1599, N907, N187, N819);
buf BUF1 (N1601, N1585);
buf BUF1 (N1602, N1578);
and AND4 (N1603, N1602, N1365, N898, N256);
or OR4 (N1604, N1600, N322, N1406, N921);
nand NAND4 (N1605, N1595, N544, N469, N1204);
nor NOR2 (N1606, N1582, N1364);
buf BUF1 (N1607, N1593);
nand NAND3 (N1608, N1607, N1188, N1505);
and AND3 (N1609, N1594, N1378, N599);
and AND4 (N1610, N1606, N1323, N103, N134);
nor NOR2 (N1611, N1604, N265);
xor XOR2 (N1612, N1611, N1479);
nand NAND4 (N1613, N1573, N1525, N1306, N64);
and AND2 (N1614, N1612, N1427);
and AND4 (N1615, N1601, N1600, N113, N698);
and AND4 (N1616, N1605, N943, N661, N119);
xor XOR2 (N1617, N1598, N1514);
nor NOR3 (N1618, N1610, N991, N1384);
not NOT1 (N1619, N1616);
not NOT1 (N1620, N1608);
nand NAND3 (N1621, N1619, N1052, N1612);
nor NOR3 (N1622, N1617, N1345, N1606);
buf BUF1 (N1623, N1618);
buf BUF1 (N1624, N1613);
not NOT1 (N1625, N1614);
xor XOR2 (N1626, N1620, N1183);
buf BUF1 (N1627, N1625);
nand NAND4 (N1628, N1624, N1391, N919, N338);
not NOT1 (N1629, N1577);
xor XOR2 (N1630, N1626, N1301);
nor NOR4 (N1631, N1615, N572, N1306, N365);
xor XOR2 (N1632, N1628, N263);
buf BUF1 (N1633, N1632);
not NOT1 (N1634, N1630);
or OR2 (N1635, N1634, N885);
not NOT1 (N1636, N1627);
nor NOR4 (N1637, N1603, N346, N897, N92);
and AND4 (N1638, N1621, N145, N755, N516);
xor XOR2 (N1639, N1633, N855);
and AND4 (N1640, N1635, N1234, N841, N576);
xor XOR2 (N1641, N1609, N916);
and AND2 (N1642, N1636, N998);
buf BUF1 (N1643, N1623);
buf BUF1 (N1644, N1638);
not NOT1 (N1645, N1629);
buf BUF1 (N1646, N1622);
nand NAND3 (N1647, N1645, N500, N554);
or OR4 (N1648, N1643, N476, N973, N1032);
nand NAND3 (N1649, N1646, N46, N71);
not NOT1 (N1650, N1647);
buf BUF1 (N1651, N1641);
not NOT1 (N1652, N1639);
and AND2 (N1653, N1650, N1442);
or OR4 (N1654, N1642, N359, N1495, N781);
not NOT1 (N1655, N1637);
and AND4 (N1656, N1655, N236, N696, N1395);
buf BUF1 (N1657, N1651);
and AND3 (N1658, N1648, N1646, N4);
and AND4 (N1659, N1654, N778, N620, N809);
xor XOR2 (N1660, N1640, N1375);
nor NOR2 (N1661, N1658, N728);
xor XOR2 (N1662, N1652, N1340);
xor XOR2 (N1663, N1659, N555);
and AND3 (N1664, N1660, N1294, N1609);
and AND3 (N1665, N1656, N914, N707);
buf BUF1 (N1666, N1662);
nor NOR3 (N1667, N1657, N1509, N1132);
and AND4 (N1668, N1665, N163, N64, N693);
nand NAND4 (N1669, N1667, N908, N788, N179);
and AND4 (N1670, N1661, N1509, N664, N1453);
or OR2 (N1671, N1669, N55);
buf BUF1 (N1672, N1671);
and AND4 (N1673, N1653, N1576, N920, N929);
buf BUF1 (N1674, N1631);
or OR3 (N1675, N1644, N456, N374);
xor XOR2 (N1676, N1672, N1601);
nor NOR4 (N1677, N1674, N131, N516, N1389);
buf BUF1 (N1678, N1664);
xor XOR2 (N1679, N1668, N347);
nand NAND2 (N1680, N1649, N807);
buf BUF1 (N1681, N1680);
buf BUF1 (N1682, N1675);
or OR4 (N1683, N1676, N746, N999, N783);
nand NAND2 (N1684, N1678, N891);
nor NOR4 (N1685, N1683, N688, N1628, N1518);
buf BUF1 (N1686, N1681);
xor XOR2 (N1687, N1673, N1279);
not NOT1 (N1688, N1687);
xor XOR2 (N1689, N1663, N202);
xor XOR2 (N1690, N1685, N846);
nor NOR3 (N1691, N1688, N730, N257);
and AND3 (N1692, N1682, N903, N479);
buf BUF1 (N1693, N1690);
and AND4 (N1694, N1666, N576, N101, N303);
buf BUF1 (N1695, N1689);
or OR2 (N1696, N1677, N254);
nand NAND4 (N1697, N1679, N632, N292, N1468);
xor XOR2 (N1698, N1697, N735);
not NOT1 (N1699, N1686);
and AND3 (N1700, N1696, N1536, N1571);
not NOT1 (N1701, N1698);
and AND4 (N1702, N1691, N595, N1283, N794);
xor XOR2 (N1703, N1692, N1249);
nor NOR2 (N1704, N1694, N1115);
or OR3 (N1705, N1684, N838, N305);
buf BUF1 (N1706, N1704);
nor NOR4 (N1707, N1670, N441, N557, N933);
and AND3 (N1708, N1702, N768, N383);
nor NOR3 (N1709, N1705, N1030, N687);
or OR2 (N1710, N1708, N14);
or OR4 (N1711, N1700, N783, N1117, N398);
or OR4 (N1712, N1706, N63, N1639, N716);
xor XOR2 (N1713, N1693, N1532);
nand NAND4 (N1714, N1711, N1417, N1649, N1194);
xor XOR2 (N1715, N1713, N56);
or OR2 (N1716, N1707, N568);
nand NAND3 (N1717, N1703, N308, N13);
nand NAND4 (N1718, N1699, N1042, N472, N687);
nand NAND4 (N1719, N1718, N279, N1595, N1273);
buf BUF1 (N1720, N1712);
nor NOR3 (N1721, N1716, N1490, N600);
and AND3 (N1722, N1710, N637, N1007);
or OR3 (N1723, N1715, N1639, N1099);
not NOT1 (N1724, N1719);
and AND2 (N1725, N1724, N392);
not NOT1 (N1726, N1714);
nand NAND2 (N1727, N1723, N1034);
or OR3 (N1728, N1722, N1060, N853);
nand NAND3 (N1729, N1695, N129, N143);
buf BUF1 (N1730, N1729);
xor XOR2 (N1731, N1720, N1161);
nand NAND3 (N1732, N1709, N1155, N1045);
xor XOR2 (N1733, N1727, N261);
xor XOR2 (N1734, N1730, N833);
nor NOR3 (N1735, N1734, N1717, N1555);
nor NOR3 (N1736, N577, N1179, N955);
or OR3 (N1737, N1731, N1351, N547);
nand NAND4 (N1738, N1732, N445, N1712, N842);
xor XOR2 (N1739, N1726, N742);
xor XOR2 (N1740, N1737, N1468);
xor XOR2 (N1741, N1739, N1495);
xor XOR2 (N1742, N1741, N160);
or OR3 (N1743, N1742, N1563, N884);
or OR4 (N1744, N1721, N142, N1509, N1530);
buf BUF1 (N1745, N1740);
xor XOR2 (N1746, N1725, N265);
nand NAND4 (N1747, N1735, N617, N253, N1574);
nor NOR2 (N1748, N1701, N595);
nor NOR3 (N1749, N1743, N1081, N1714);
not NOT1 (N1750, N1733);
nand NAND4 (N1751, N1738, N810, N616, N733);
nor NOR2 (N1752, N1747, N1627);
and AND2 (N1753, N1745, N758);
buf BUF1 (N1754, N1744);
buf BUF1 (N1755, N1752);
buf BUF1 (N1756, N1754);
nor NOR3 (N1757, N1753, N1705, N1350);
nand NAND3 (N1758, N1757, N1045, N1318);
nand NAND2 (N1759, N1756, N1662);
not NOT1 (N1760, N1750);
and AND4 (N1761, N1748, N1112, N1745, N760);
not NOT1 (N1762, N1758);
not NOT1 (N1763, N1728);
nor NOR2 (N1764, N1736, N1231);
nand NAND4 (N1765, N1763, N160, N1175, N469);
buf BUF1 (N1766, N1751);
xor XOR2 (N1767, N1764, N82);
nand NAND2 (N1768, N1755, N934);
and AND3 (N1769, N1768, N1518, N1405);
not NOT1 (N1770, N1746);
buf BUF1 (N1771, N1767);
nor NOR4 (N1772, N1769, N1294, N1467, N1212);
not NOT1 (N1773, N1770);
or OR2 (N1774, N1773, N538);
nand NAND3 (N1775, N1771, N1489, N1284);
or OR2 (N1776, N1774, N1383);
nand NAND4 (N1777, N1749, N1423, N123, N1516);
nor NOR3 (N1778, N1777, N231, N1197);
or OR2 (N1779, N1776, N1473);
or OR3 (N1780, N1762, N2, N303);
nor NOR2 (N1781, N1775, N306);
buf BUF1 (N1782, N1772);
buf BUF1 (N1783, N1760);
xor XOR2 (N1784, N1778, N1010);
xor XOR2 (N1785, N1759, N1139);
xor XOR2 (N1786, N1785, N394);
nor NOR2 (N1787, N1783, N475);
or OR4 (N1788, N1780, N1247, N200, N683);
nand NAND3 (N1789, N1765, N582, N1127);
nor NOR2 (N1790, N1781, N1463);
and AND2 (N1791, N1786, N987);
or OR3 (N1792, N1791, N1312, N943);
nor NOR4 (N1793, N1789, N1495, N1527, N359);
nand NAND3 (N1794, N1766, N1485, N564);
not NOT1 (N1795, N1787);
nand NAND4 (N1796, N1794, N1742, N1603, N1775);
buf BUF1 (N1797, N1784);
and AND3 (N1798, N1790, N1603, N1155);
buf BUF1 (N1799, N1797);
or OR3 (N1800, N1798, N231, N1600);
or OR4 (N1801, N1795, N1432, N706, N947);
nand NAND3 (N1802, N1793, N460, N957);
nand NAND2 (N1803, N1796, N1676);
not NOT1 (N1804, N1803);
nor NOR2 (N1805, N1779, N923);
buf BUF1 (N1806, N1801);
nand NAND2 (N1807, N1788, N961);
and AND2 (N1808, N1806, N534);
nor NOR2 (N1809, N1761, N862);
and AND2 (N1810, N1792, N847);
xor XOR2 (N1811, N1810, N590);
buf BUF1 (N1812, N1799);
nor NOR4 (N1813, N1809, N1059, N1429, N794);
not NOT1 (N1814, N1811);
or OR4 (N1815, N1807, N52, N1719, N1288);
not NOT1 (N1816, N1800);
and AND2 (N1817, N1812, N989);
buf BUF1 (N1818, N1802);
not NOT1 (N1819, N1818);
or OR2 (N1820, N1805, N1153);
not NOT1 (N1821, N1808);
buf BUF1 (N1822, N1813);
not NOT1 (N1823, N1822);
xor XOR2 (N1824, N1814, N920);
buf BUF1 (N1825, N1782);
nand NAND4 (N1826, N1823, N224, N1724, N1671);
or OR2 (N1827, N1825, N502);
nor NOR2 (N1828, N1820, N1386);
not NOT1 (N1829, N1804);
and AND4 (N1830, N1826, N1828, N1536, N855);
xor XOR2 (N1831, N715, N257);
nand NAND3 (N1832, N1816, N757, N593);
not NOT1 (N1833, N1819);
xor XOR2 (N1834, N1821, N1624);
or OR4 (N1835, N1827, N99, N416, N1185);
nor NOR2 (N1836, N1832, N674);
nand NAND4 (N1837, N1835, N829, N960, N1234);
not NOT1 (N1838, N1833);
nor NOR3 (N1839, N1817, N575, N1112);
nand NAND4 (N1840, N1831, N1723, N768, N1528);
buf BUF1 (N1841, N1834);
not NOT1 (N1842, N1840);
nor NOR3 (N1843, N1836, N1727, N223);
not NOT1 (N1844, N1824);
not NOT1 (N1845, N1837);
xor XOR2 (N1846, N1842, N346);
buf BUF1 (N1847, N1838);
nor NOR3 (N1848, N1846, N847, N442);
xor XOR2 (N1849, N1815, N208);
xor XOR2 (N1850, N1829, N930);
not NOT1 (N1851, N1830);
or OR4 (N1852, N1844, N984, N847, N189);
not NOT1 (N1853, N1852);
nand NAND3 (N1854, N1845, N392, N819);
or OR2 (N1855, N1849, N889);
not NOT1 (N1856, N1855);
buf BUF1 (N1857, N1841);
nor NOR2 (N1858, N1843, N118);
not NOT1 (N1859, N1851);
and AND4 (N1860, N1859, N1279, N1622, N998);
buf BUF1 (N1861, N1858);
not NOT1 (N1862, N1861);
or OR2 (N1863, N1853, N1189);
not NOT1 (N1864, N1848);
and AND4 (N1865, N1863, N1857, N1740, N1357);
xor XOR2 (N1866, N1200, N1232);
xor XOR2 (N1867, N1862, N594);
nor NOR4 (N1868, N1867, N1675, N1649, N526);
not NOT1 (N1869, N1865);
not NOT1 (N1870, N1847);
and AND3 (N1871, N1854, N1674, N1111);
buf BUF1 (N1872, N1866);
nor NOR2 (N1873, N1839, N1698);
buf BUF1 (N1874, N1856);
nand NAND3 (N1875, N1850, N124, N431);
buf BUF1 (N1876, N1875);
nor NOR2 (N1877, N1864, N1543);
not NOT1 (N1878, N1860);
nand NAND4 (N1879, N1878, N164, N1860, N616);
and AND3 (N1880, N1869, N119, N1247);
nor NOR2 (N1881, N1879, N1157);
not NOT1 (N1882, N1873);
not NOT1 (N1883, N1881);
nor NOR2 (N1884, N1870, N1146);
and AND3 (N1885, N1880, N1243, N1876);
buf BUF1 (N1886, N1641);
and AND4 (N1887, N1868, N1131, N628, N533);
buf BUF1 (N1888, N1886);
not NOT1 (N1889, N1882);
buf BUF1 (N1890, N1888);
or OR3 (N1891, N1872, N1291, N1103);
nand NAND4 (N1892, N1874, N1822, N322, N1847);
not NOT1 (N1893, N1871);
buf BUF1 (N1894, N1890);
not NOT1 (N1895, N1893);
xor XOR2 (N1896, N1885, N1348);
and AND4 (N1897, N1877, N636, N179, N1116);
and AND2 (N1898, N1889, N1790);
buf BUF1 (N1899, N1883);
nor NOR2 (N1900, N1895, N528);
buf BUF1 (N1901, N1891);
not NOT1 (N1902, N1887);
buf BUF1 (N1903, N1901);
and AND3 (N1904, N1894, N1027, N1052);
xor XOR2 (N1905, N1903, N1029);
buf BUF1 (N1906, N1892);
xor XOR2 (N1907, N1898, N1403);
not NOT1 (N1908, N1884);
nand NAND2 (N1909, N1899, N960);
or OR4 (N1910, N1902, N1351, N234, N783);
not NOT1 (N1911, N1906);
buf BUF1 (N1912, N1911);
nand NAND2 (N1913, N1907, N1889);
nor NOR4 (N1914, N1913, N723, N671, N958);
and AND4 (N1915, N1910, N96, N1414, N580);
and AND3 (N1916, N1909, N785, N365);
xor XOR2 (N1917, N1897, N1808);
not NOT1 (N1918, N1905);
and AND3 (N1919, N1900, N1649, N1065);
not NOT1 (N1920, N1914);
nand NAND2 (N1921, N1917, N1173);
or OR2 (N1922, N1904, N293);
buf BUF1 (N1923, N1920);
not NOT1 (N1924, N1922);
or OR3 (N1925, N1916, N325, N1515);
nand NAND4 (N1926, N1925, N1274, N1226, N744);
nor NOR4 (N1927, N1912, N371, N1204, N136);
xor XOR2 (N1928, N1915, N903);
not NOT1 (N1929, N1918);
xor XOR2 (N1930, N1928, N364);
and AND3 (N1931, N1908, N1110, N903);
not NOT1 (N1932, N1930);
xor XOR2 (N1933, N1921, N1647);
buf BUF1 (N1934, N1929);
and AND4 (N1935, N1927, N1763, N403, N1369);
buf BUF1 (N1936, N1935);
buf BUF1 (N1937, N1923);
or OR2 (N1938, N1931, N1530);
nand NAND3 (N1939, N1896, N1916, N833);
xor XOR2 (N1940, N1926, N1322);
xor XOR2 (N1941, N1924, N1597);
nor NOR4 (N1942, N1940, N226, N329, N580);
xor XOR2 (N1943, N1937, N565);
not NOT1 (N1944, N1932);
nand NAND2 (N1945, N1936, N1136);
nor NOR3 (N1946, N1939, N570, N1236);
and AND2 (N1947, N1943, N743);
nand NAND3 (N1948, N1933, N376, N803);
buf BUF1 (N1949, N1919);
or OR2 (N1950, N1945, N1411);
or OR3 (N1951, N1941, N1369, N1120);
xor XOR2 (N1952, N1944, N1142);
not NOT1 (N1953, N1946);
not NOT1 (N1954, N1947);
nor NOR3 (N1955, N1942, N1463, N1114);
and AND2 (N1956, N1938, N780);
not NOT1 (N1957, N1952);
not NOT1 (N1958, N1948);
and AND2 (N1959, N1957, N1763);
nand NAND2 (N1960, N1951, N1231);
xor XOR2 (N1961, N1949, N1245);
or OR4 (N1962, N1954, N1030, N1404, N555);
and AND2 (N1963, N1950, N1630);
buf BUF1 (N1964, N1934);
xor XOR2 (N1965, N1959, N534);
xor XOR2 (N1966, N1961, N1370);
xor XOR2 (N1967, N1962, N1303);
and AND3 (N1968, N1963, N259, N711);
nor NOR3 (N1969, N1953, N582, N1201);
xor XOR2 (N1970, N1955, N1965);
or OR2 (N1971, N641, N1359);
nand NAND4 (N1972, N1969, N1741, N55, N1032);
nor NOR3 (N1973, N1968, N1462, N797);
or OR3 (N1974, N1972, N1011, N123);
not NOT1 (N1975, N1973);
not NOT1 (N1976, N1964);
xor XOR2 (N1977, N1958, N1681);
and AND3 (N1978, N1975, N697, N544);
or OR3 (N1979, N1977, N1904, N394);
or OR2 (N1980, N1978, N936);
nor NOR4 (N1981, N1970, N1800, N447, N1653);
nand NAND3 (N1982, N1974, N608, N205);
nor NOR2 (N1983, N1976, N888);
and AND3 (N1984, N1966, N399, N1292);
nand NAND3 (N1985, N1982, N1929, N838);
not NOT1 (N1986, N1960);
nand NAND4 (N1987, N1981, N492, N558, N1030);
nor NOR3 (N1988, N1987, N1598, N5);
not NOT1 (N1989, N1988);
not NOT1 (N1990, N1983);
not NOT1 (N1991, N1971);
nand NAND3 (N1992, N1986, N744, N803);
nor NOR2 (N1993, N1989, N214);
nand NAND2 (N1994, N1967, N395);
and AND2 (N1995, N1993, N1304);
xor XOR2 (N1996, N1992, N736);
or OR2 (N1997, N1980, N1912);
xor XOR2 (N1998, N1956, N618);
nand NAND3 (N1999, N1997, N1460, N986);
and AND3 (N2000, N1985, N342, N564);
and AND2 (N2001, N1984, N1821);
and AND3 (N2002, N1994, N882, N1953);
or OR4 (N2003, N2000, N346, N1688, N29);
xor XOR2 (N2004, N2002, N284);
or OR3 (N2005, N1990, N1525, N1500);
buf BUF1 (N2006, N1991);
xor XOR2 (N2007, N2004, N481);
nor NOR3 (N2008, N1995, N1184, N1371);
or OR3 (N2009, N1999, N1144, N778);
or OR3 (N2010, N1998, N487, N998);
nor NOR4 (N2011, N2006, N2001, N244, N346);
nand NAND4 (N2012, N1924, N1257, N640, N392);
and AND2 (N2013, N2003, N1127);
not NOT1 (N2014, N2008);
or OR3 (N2015, N2012, N1559, N456);
xor XOR2 (N2016, N2009, N399);
nor NOR3 (N2017, N2010, N266, N1723);
nor NOR2 (N2018, N2007, N383);
or OR4 (N2019, N2016, N1269, N756, N393);
nor NOR2 (N2020, N2013, N1312);
xor XOR2 (N2021, N2014, N1460);
buf BUF1 (N2022, N2019);
xor XOR2 (N2023, N2022, N211);
or OR4 (N2024, N2021, N1449, N1803, N1190);
not NOT1 (N2025, N1979);
or OR4 (N2026, N2023, N1421, N1739, N1879);
and AND4 (N2027, N2025, N1005, N478, N1483);
or OR2 (N2028, N2011, N1925);
nand NAND2 (N2029, N2028, N1614);
nand NAND4 (N2030, N2029, N328, N1188, N446);
nand NAND3 (N2031, N1996, N1091, N1811);
not NOT1 (N2032, N2017);
nand NAND4 (N2033, N2032, N1560, N562, N699);
and AND3 (N2034, N2024, N415, N1886);
not NOT1 (N2035, N2020);
and AND3 (N2036, N2030, N1340, N828);
nand NAND4 (N2037, N2035, N1516, N637, N374);
xor XOR2 (N2038, N2033, N19);
not NOT1 (N2039, N2036);
nand NAND2 (N2040, N2015, N637);
or OR2 (N2041, N2040, N1784);
nor NOR4 (N2042, N2026, N1022, N526, N1726);
buf BUF1 (N2043, N2005);
nand NAND4 (N2044, N2039, N1720, N1234, N67);
xor XOR2 (N2045, N2037, N64);
nor NOR2 (N2046, N2043, N626);
buf BUF1 (N2047, N2044);
not NOT1 (N2048, N2046);
xor XOR2 (N2049, N2042, N481);
nor NOR3 (N2050, N2034, N2018, N186);
or OR4 (N2051, N747, N1740, N1301, N380);
xor XOR2 (N2052, N2049, N1503);
not NOT1 (N2053, N2051);
nor NOR2 (N2054, N2050, N1555);
not NOT1 (N2055, N2031);
and AND3 (N2056, N2027, N695, N1779);
or OR4 (N2057, N2038, N1738, N1873, N403);
xor XOR2 (N2058, N2045, N2047);
nor NOR2 (N2059, N1729, N1698);
nor NOR2 (N2060, N2056, N1547);
and AND3 (N2061, N2059, N1544, N49);
xor XOR2 (N2062, N2055, N822);
and AND4 (N2063, N2062, N350, N177, N756);
nor NOR3 (N2064, N2053, N1095, N673);
nand NAND2 (N2065, N2061, N1705);
not NOT1 (N2066, N2048);
xor XOR2 (N2067, N2052, N625);
not NOT1 (N2068, N2066);
and AND3 (N2069, N2054, N135, N694);
or OR3 (N2070, N2057, N1232, N1646);
buf BUF1 (N2071, N2060);
nor NOR4 (N2072, N2065, N21, N147, N2044);
nand NAND3 (N2073, N2071, N1297, N1434);
buf BUF1 (N2074, N2069);
buf BUF1 (N2075, N2058);
nand NAND2 (N2076, N2064, N1893);
and AND3 (N2077, N2074, N1915, N1896);
not NOT1 (N2078, N2072);
or OR4 (N2079, N2068, N1670, N1540, N1124);
or OR2 (N2080, N2077, N616);
buf BUF1 (N2081, N2076);
buf BUF1 (N2082, N2080);
or OR2 (N2083, N2079, N279);
xor XOR2 (N2084, N2083, N494);
xor XOR2 (N2085, N2041, N251);
or OR2 (N2086, N2067, N1734);
nand NAND3 (N2087, N2075, N1601, N1196);
or OR2 (N2088, N2078, N2066);
and AND2 (N2089, N2088, N413);
buf BUF1 (N2090, N2086);
or OR3 (N2091, N2087, N412, N1123);
nor NOR4 (N2092, N2089, N1009, N390, N1751);
xor XOR2 (N2093, N2092, N272);
nor NOR2 (N2094, N2093, N1111);
and AND4 (N2095, N2091, N890, N1259, N1834);
and AND4 (N2096, N2082, N20, N111, N190);
nand NAND4 (N2097, N2084, N300, N941, N1312);
xor XOR2 (N2098, N2073, N1024);
xor XOR2 (N2099, N2096, N1936);
or OR2 (N2100, N2090, N785);
buf BUF1 (N2101, N2095);
buf BUF1 (N2102, N2101);
nand NAND2 (N2103, N2094, N441);
xor XOR2 (N2104, N2081, N240);
nor NOR4 (N2105, N2063, N1923, N753, N856);
nor NOR3 (N2106, N2097, N1498, N824);
not NOT1 (N2107, N2085);
xor XOR2 (N2108, N2105, N172);
not NOT1 (N2109, N2108);
buf BUF1 (N2110, N2100);
buf BUF1 (N2111, N2098);
and AND4 (N2112, N2109, N720, N233, N823);
and AND2 (N2113, N2102, N505);
nand NAND4 (N2114, N2099, N1450, N161, N1106);
nor NOR4 (N2115, N2110, N956, N1091, N1809);
and AND4 (N2116, N2114, N798, N1448, N625);
buf BUF1 (N2117, N2106);
nand NAND4 (N2118, N2107, N508, N1995, N1757);
and AND4 (N2119, N2070, N825, N544, N1246);
nor NOR2 (N2120, N2117, N204);
nor NOR3 (N2121, N2119, N1146, N1001);
and AND4 (N2122, N2118, N1173, N676, N631);
nand NAND2 (N2123, N2103, N975);
nor NOR2 (N2124, N2121, N1964);
xor XOR2 (N2125, N2116, N1697);
or OR4 (N2126, N2104, N39, N1195, N437);
xor XOR2 (N2127, N2122, N877);
buf BUF1 (N2128, N2115);
xor XOR2 (N2129, N2123, N337);
not NOT1 (N2130, N2124);
xor XOR2 (N2131, N2111, N545);
xor XOR2 (N2132, N2126, N1524);
and AND3 (N2133, N2125, N104, N938);
nand NAND4 (N2134, N2127, N926, N1317, N1449);
nand NAND4 (N2135, N2128, N11, N1585, N262);
or OR2 (N2136, N2130, N1938);
xor XOR2 (N2137, N2120, N1653);
buf BUF1 (N2138, N2137);
and AND2 (N2139, N2112, N613);
nor NOR3 (N2140, N2113, N240, N1091);
nand NAND4 (N2141, N2129, N1523, N1582, N2053);
buf BUF1 (N2142, N2133);
xor XOR2 (N2143, N2134, N885);
and AND3 (N2144, N2132, N1379, N1254);
buf BUF1 (N2145, N2136);
xor XOR2 (N2146, N2135, N1009);
xor XOR2 (N2147, N2138, N43);
nor NOR4 (N2148, N2142, N1616, N328, N658);
nor NOR4 (N2149, N2147, N56, N872, N937);
nand NAND2 (N2150, N2144, N730);
and AND3 (N2151, N2143, N1104, N1124);
nand NAND4 (N2152, N2146, N1619, N1316, N1878);
and AND4 (N2153, N2141, N1680, N1858, N938);
and AND2 (N2154, N2131, N1389);
nand NAND4 (N2155, N2148, N105, N1121, N1789);
and AND2 (N2156, N2140, N274);
or OR3 (N2157, N2154, N462, N457);
and AND4 (N2158, N2151, N1284, N1353, N603);
and AND3 (N2159, N2158, N190, N1333);
or OR2 (N2160, N2139, N305);
or OR2 (N2161, N2150, N574);
xor XOR2 (N2162, N2145, N1146);
or OR4 (N2163, N2156, N1998, N1565, N1465);
nand NAND3 (N2164, N2162, N1037, N1016);
xor XOR2 (N2165, N2152, N1798);
xor XOR2 (N2166, N2160, N336);
buf BUF1 (N2167, N2161);
nand NAND2 (N2168, N2163, N179);
and AND3 (N2169, N2164, N761, N944);
buf BUF1 (N2170, N2165);
xor XOR2 (N2171, N2168, N991);
or OR4 (N2172, N2155, N1313, N1387, N303);
buf BUF1 (N2173, N2170);
not NOT1 (N2174, N2149);
nor NOR3 (N2175, N2159, N2114, N1477);
nand NAND3 (N2176, N2172, N1380, N783);
or OR3 (N2177, N2153, N2014, N889);
nor NOR2 (N2178, N2167, N642);
nor NOR4 (N2179, N2171, N156, N570, N426);
not NOT1 (N2180, N2174);
nand NAND4 (N2181, N2177, N1410, N1402, N1207);
and AND2 (N2182, N2173, N17);
buf BUF1 (N2183, N2182);
not NOT1 (N2184, N2176);
xor XOR2 (N2185, N2180, N1407);
and AND2 (N2186, N2166, N1229);
nor NOR4 (N2187, N2185, N1783, N110, N655);
xor XOR2 (N2188, N2181, N1591);
or OR2 (N2189, N2188, N635);
buf BUF1 (N2190, N2178);
nand NAND3 (N2191, N2187, N1318, N1474);
xor XOR2 (N2192, N2157, N20);
xor XOR2 (N2193, N2183, N545);
or OR3 (N2194, N2184, N523, N2093);
not NOT1 (N2195, N2194);
buf BUF1 (N2196, N2175);
and AND3 (N2197, N2192, N1069, N1877);
nand NAND2 (N2198, N2179, N67);
nor NOR3 (N2199, N2189, N312, N861);
buf BUF1 (N2200, N2197);
not NOT1 (N2201, N2198);
or OR3 (N2202, N2196, N1952, N1463);
or OR4 (N2203, N2191, N1899, N2086, N286);
nand NAND2 (N2204, N2199, N244);
and AND3 (N2205, N2169, N1, N1406);
or OR4 (N2206, N2202, N642, N1334, N261);
or OR2 (N2207, N2203, N1860);
or OR3 (N2208, N2190, N1643, N403);
nor NOR4 (N2209, N2204, N1260, N417, N1525);
nor NOR2 (N2210, N2208, N423);
and AND2 (N2211, N2205, N1684);
nor NOR4 (N2212, N2209, N1678, N873, N598);
nand NAND3 (N2213, N2186, N1921, N1835);
and AND2 (N2214, N2195, N1174);
nand NAND3 (N2215, N2214, N1386, N648);
xor XOR2 (N2216, N2213, N689);
or OR4 (N2217, N2206, N466, N1873, N386);
and AND4 (N2218, N2210, N195, N861, N964);
nand NAND3 (N2219, N2207, N1999, N2034);
and AND2 (N2220, N2218, N932);
nand NAND2 (N2221, N2200, N1288);
buf BUF1 (N2222, N2215);
or OR2 (N2223, N2219, N660);
buf BUF1 (N2224, N2211);
xor XOR2 (N2225, N2223, N1967);
buf BUF1 (N2226, N2221);
not NOT1 (N2227, N2222);
buf BUF1 (N2228, N2216);
or OR3 (N2229, N2193, N842, N1754);
xor XOR2 (N2230, N2228, N1301);
not NOT1 (N2231, N2226);
not NOT1 (N2232, N2231);
not NOT1 (N2233, N2212);
buf BUF1 (N2234, N2225);
and AND3 (N2235, N2232, N1935, N534);
xor XOR2 (N2236, N2233, N125);
and AND3 (N2237, N2217, N1554, N1504);
nand NAND3 (N2238, N2220, N1453, N1654);
nand NAND4 (N2239, N2229, N1971, N2222, N1559);
nand NAND3 (N2240, N2234, N2078, N960);
not NOT1 (N2241, N2230);
nor NOR2 (N2242, N2236, N2126);
nand NAND2 (N2243, N2224, N62);
buf BUF1 (N2244, N2201);
nor NOR4 (N2245, N2239, N1259, N552, N2129);
or OR2 (N2246, N2241, N1311);
xor XOR2 (N2247, N2243, N2202);
nor NOR2 (N2248, N2247, N161);
or OR4 (N2249, N2242, N858, N1728, N1190);
buf BUF1 (N2250, N2235);
nor NOR2 (N2251, N2244, N1766);
not NOT1 (N2252, N2227);
nand NAND3 (N2253, N2251, N1175, N871);
buf BUF1 (N2254, N2252);
xor XOR2 (N2255, N2250, N206);
nand NAND2 (N2256, N2245, N1756);
xor XOR2 (N2257, N2249, N602);
nor NOR3 (N2258, N2240, N1540, N691);
xor XOR2 (N2259, N2258, N861);
xor XOR2 (N2260, N2246, N981);
and AND3 (N2261, N2259, N1040, N1139);
and AND3 (N2262, N2256, N1406, N178);
not NOT1 (N2263, N2262);
nor NOR2 (N2264, N2255, N1750);
xor XOR2 (N2265, N2260, N2110);
not NOT1 (N2266, N2265);
xor XOR2 (N2267, N2263, N74);
nand NAND2 (N2268, N2237, N1901);
buf BUF1 (N2269, N2254);
nor NOR3 (N2270, N2261, N782, N1065);
or OR4 (N2271, N2266, N1108, N862, N969);
and AND2 (N2272, N2248, N1698);
buf BUF1 (N2273, N2269);
and AND2 (N2274, N2257, N1322);
not NOT1 (N2275, N2264);
nor NOR2 (N2276, N2271, N1462);
nand NAND2 (N2277, N2270, N640);
nor NOR2 (N2278, N2268, N1282);
and AND2 (N2279, N2238, N613);
or OR4 (N2280, N2274, N1963, N2044, N1819);
nor NOR4 (N2281, N2267, N1249, N1472, N197);
and AND3 (N2282, N2276, N1932, N86);
nand NAND3 (N2283, N2281, N846, N850);
and AND2 (N2284, N2280, N1380);
not NOT1 (N2285, N2275);
nor NOR4 (N2286, N2278, N259, N1453, N1975);
nand NAND3 (N2287, N2284, N62, N1929);
or OR3 (N2288, N2282, N1205, N546);
not NOT1 (N2289, N2285);
and AND2 (N2290, N2277, N1561);
not NOT1 (N2291, N2253);
not NOT1 (N2292, N2279);
not NOT1 (N2293, N2291);
buf BUF1 (N2294, N2288);
or OR2 (N2295, N2283, N676);
and AND4 (N2296, N2286, N395, N993, N941);
nand NAND4 (N2297, N2273, N349, N385, N1535);
buf BUF1 (N2298, N2294);
nor NOR4 (N2299, N2287, N595, N724, N2289);
buf BUF1 (N2300, N855);
buf BUF1 (N2301, N2300);
buf BUF1 (N2302, N2295);
buf BUF1 (N2303, N2290);
nor NOR2 (N2304, N2301, N500);
and AND4 (N2305, N2292, N1696, N1813, N161);
nor NOR4 (N2306, N2302, N717, N1053, N787);
nor NOR4 (N2307, N2296, N1266, N849, N736);
nand NAND3 (N2308, N2272, N590, N1787);
not NOT1 (N2309, N2307);
buf BUF1 (N2310, N2299);
nand NAND2 (N2311, N2297, N1617);
nand NAND4 (N2312, N2306, N241, N213, N2279);
xor XOR2 (N2313, N2309, N1062);
nand NAND4 (N2314, N2303, N433, N409, N1997);
nor NOR3 (N2315, N2304, N1872, N2071);
nand NAND3 (N2316, N2298, N1737, N2016);
and AND3 (N2317, N2316, N1804, N1489);
nand NAND3 (N2318, N2315, N129, N1112);
nand NAND3 (N2319, N2312, N720, N2258);
nor NOR2 (N2320, N2308, N1304);
xor XOR2 (N2321, N2319, N602);
nand NAND3 (N2322, N2320, N375, N1220);
buf BUF1 (N2323, N2317);
nand NAND4 (N2324, N2318, N2169, N415, N1923);
xor XOR2 (N2325, N2322, N225);
nor NOR4 (N2326, N2311, N111, N1202, N1552);
nand NAND3 (N2327, N2314, N2044, N1466);
nand NAND4 (N2328, N2323, N955, N1668, N985);
buf BUF1 (N2329, N2326);
nor NOR2 (N2330, N2324, N406);
xor XOR2 (N2331, N2330, N569);
xor XOR2 (N2332, N2325, N871);
not NOT1 (N2333, N2328);
buf BUF1 (N2334, N2321);
not NOT1 (N2335, N2310);
xor XOR2 (N2336, N2331, N1737);
xor XOR2 (N2337, N2329, N1826);
and AND4 (N2338, N2327, N1606, N2240, N1605);
and AND4 (N2339, N2337, N133, N1564, N2307);
xor XOR2 (N2340, N2333, N1217);
not NOT1 (N2341, N2334);
nand NAND3 (N2342, N2336, N1225, N1808);
or OR3 (N2343, N2335, N288, N147);
xor XOR2 (N2344, N2313, N595);
buf BUF1 (N2345, N2341);
nor NOR4 (N2346, N2342, N639, N99, N2068);
buf BUF1 (N2347, N2343);
buf BUF1 (N2348, N2305);
nor NOR3 (N2349, N2332, N442, N79);
and AND2 (N2350, N2347, N200);
and AND4 (N2351, N2345, N99, N785, N1099);
or OR3 (N2352, N2344, N817, N1768);
or OR4 (N2353, N2348, N882, N611, N48);
nor NOR3 (N2354, N2349, N98, N2101);
nor NOR2 (N2355, N2338, N693);
or OR3 (N2356, N2354, N2312, N1256);
not NOT1 (N2357, N2346);
and AND4 (N2358, N2350, N2209, N1142, N2137);
not NOT1 (N2359, N2340);
and AND3 (N2360, N2359, N610, N1264);
buf BUF1 (N2361, N2356);
not NOT1 (N2362, N2361);
nand NAND3 (N2363, N2355, N1672, N609);
buf BUF1 (N2364, N2362);
and AND3 (N2365, N2293, N1493, N403);
or OR4 (N2366, N2351, N1817, N890, N1423);
and AND3 (N2367, N2357, N2350, N355);
and AND4 (N2368, N2352, N639, N1970, N281);
not NOT1 (N2369, N2358);
buf BUF1 (N2370, N2365);
or OR3 (N2371, N2367, N1226, N718);
nand NAND4 (N2372, N2371, N784, N1514, N1553);
not NOT1 (N2373, N2369);
buf BUF1 (N2374, N2363);
buf BUF1 (N2375, N2353);
nor NOR3 (N2376, N2375, N1745, N864);
buf BUF1 (N2377, N2373);
nor NOR4 (N2378, N2370, N2258, N2051, N1022);
xor XOR2 (N2379, N2374, N2235);
not NOT1 (N2380, N2339);
and AND2 (N2381, N2380, N914);
and AND4 (N2382, N2379, N1526, N989, N318);
or OR4 (N2383, N2372, N173, N1319, N2285);
xor XOR2 (N2384, N2377, N2140);
not NOT1 (N2385, N2382);
or OR3 (N2386, N2366, N1923, N1289);
nand NAND3 (N2387, N2385, N1637, N295);
nor NOR4 (N2388, N2368, N425, N512, N492);
nor NOR3 (N2389, N2383, N187, N39);
xor XOR2 (N2390, N2360, N1329);
or OR4 (N2391, N2378, N2183, N1466, N674);
buf BUF1 (N2392, N2389);
xor XOR2 (N2393, N2376, N1918);
buf BUF1 (N2394, N2391);
buf BUF1 (N2395, N2364);
or OR3 (N2396, N2393, N528, N1951);
xor XOR2 (N2397, N2381, N79);
buf BUF1 (N2398, N2395);
buf BUF1 (N2399, N2396);
buf BUF1 (N2400, N2386);
buf BUF1 (N2401, N2399);
and AND2 (N2402, N2397, N1164);
xor XOR2 (N2403, N2394, N630);
xor XOR2 (N2404, N2398, N1410);
nand NAND3 (N2405, N2387, N1149, N924);
and AND3 (N2406, N2388, N2168, N2);
nor NOR4 (N2407, N2400, N552, N600, N293);
and AND4 (N2408, N2407, N1620, N1540, N1763);
and AND3 (N2409, N2402, N866, N1252);
xor XOR2 (N2410, N2384, N1737);
and AND3 (N2411, N2392, N835, N604);
and AND4 (N2412, N2390, N199, N1149, N868);
and AND4 (N2413, N2406, N91, N2143, N1262);
buf BUF1 (N2414, N2405);
nand NAND3 (N2415, N2413, N244, N1909);
not NOT1 (N2416, N2414);
xor XOR2 (N2417, N2410, N893);
nand NAND3 (N2418, N2403, N2343, N519);
nor NOR2 (N2419, N2417, N732);
buf BUF1 (N2420, N2409);
nor NOR2 (N2421, N2411, N741);
and AND3 (N2422, N2416, N584, N2253);
and AND2 (N2423, N2420, N941);
nand NAND3 (N2424, N2404, N168, N37);
xor XOR2 (N2425, N2408, N1270);
and AND2 (N2426, N2423, N1211);
buf BUF1 (N2427, N2421);
nor NOR3 (N2428, N2422, N772, N1219);
nand NAND2 (N2429, N2427, N1980);
or OR3 (N2430, N2401, N907, N1117);
and AND3 (N2431, N2426, N2013, N1858);
not NOT1 (N2432, N2428);
xor XOR2 (N2433, N2431, N526);
xor XOR2 (N2434, N2418, N2372);
and AND4 (N2435, N2412, N840, N398, N1909);
not NOT1 (N2436, N2430);
and AND4 (N2437, N2436, N815, N78, N1601);
xor XOR2 (N2438, N2435, N129);
and AND3 (N2439, N2415, N1414, N179);
xor XOR2 (N2440, N2424, N1084);
nor NOR3 (N2441, N2419, N263, N1461);
and AND2 (N2442, N2441, N888);
nor NOR2 (N2443, N2434, N2089);
xor XOR2 (N2444, N2429, N1885);
not NOT1 (N2445, N2443);
buf BUF1 (N2446, N2442);
xor XOR2 (N2447, N2439, N1937);
not NOT1 (N2448, N2447);
nor NOR2 (N2449, N2437, N381);
xor XOR2 (N2450, N2440, N1325);
and AND4 (N2451, N2445, N632, N1606, N675);
not NOT1 (N2452, N2438);
nand NAND4 (N2453, N2444, N97, N8, N423);
xor XOR2 (N2454, N2453, N2364);
not NOT1 (N2455, N2452);
or OR3 (N2456, N2451, N1537, N1717);
xor XOR2 (N2457, N2454, N2096);
xor XOR2 (N2458, N2448, N1974);
or OR2 (N2459, N2425, N2340);
buf BUF1 (N2460, N2459);
not NOT1 (N2461, N2449);
or OR4 (N2462, N2455, N913, N1321, N794);
and AND2 (N2463, N2457, N2366);
and AND3 (N2464, N2450, N1003, N1978);
buf BUF1 (N2465, N2446);
not NOT1 (N2466, N2460);
xor XOR2 (N2467, N2461, N1648);
or OR2 (N2468, N2465, N2310);
xor XOR2 (N2469, N2432, N2060);
xor XOR2 (N2470, N2466, N120);
nor NOR3 (N2471, N2470, N1486, N1917);
nor NOR2 (N2472, N2467, N837);
nand NAND2 (N2473, N2456, N212);
not NOT1 (N2474, N2464);
and AND3 (N2475, N2469, N481, N1255);
or OR3 (N2476, N2473, N2187, N1840);
not NOT1 (N2477, N2471);
not NOT1 (N2478, N2475);
nor NOR2 (N2479, N2468, N411);
not NOT1 (N2480, N2478);
xor XOR2 (N2481, N2480, N329);
xor XOR2 (N2482, N2433, N1271);
or OR2 (N2483, N2481, N1299);
nand NAND4 (N2484, N2477, N2309, N1338, N616);
nand NAND2 (N2485, N2479, N554);
xor XOR2 (N2486, N2485, N432);
xor XOR2 (N2487, N2472, N1746);
nand NAND4 (N2488, N2483, N2071, N2291, N1431);
and AND4 (N2489, N2462, N295, N1230, N698);
nand NAND3 (N2490, N2482, N2290, N1961);
or OR4 (N2491, N2488, N1114, N2169, N14);
nand NAND3 (N2492, N2476, N1311, N2249);
nor NOR2 (N2493, N2489, N2463);
and AND3 (N2494, N2184, N1305, N2172);
buf BUF1 (N2495, N2493);
not NOT1 (N2496, N2491);
and AND2 (N2497, N2484, N424);
nand NAND2 (N2498, N2496, N582);
buf BUF1 (N2499, N2492);
xor XOR2 (N2500, N2458, N2006);
or OR3 (N2501, N2500, N1398, N426);
nor NOR2 (N2502, N2497, N63);
nand NAND4 (N2503, N2487, N2365, N1651, N2053);
buf BUF1 (N2504, N2499);
nand NAND3 (N2505, N2502, N1600, N366);
not NOT1 (N2506, N2498);
and AND2 (N2507, N2494, N1954);
not NOT1 (N2508, N2490);
nand NAND4 (N2509, N2508, N1796, N2497, N1673);
not NOT1 (N2510, N2474);
nor NOR3 (N2511, N2510, N338, N953);
nor NOR3 (N2512, N2511, N1994, N693);
xor XOR2 (N2513, N2501, N1013);
nor NOR2 (N2514, N2486, N2333);
not NOT1 (N2515, N2505);
buf BUF1 (N2516, N2513);
not NOT1 (N2517, N2503);
and AND2 (N2518, N2512, N1079);
buf BUF1 (N2519, N2504);
and AND3 (N2520, N2506, N913, N95);
nand NAND4 (N2521, N2514, N2037, N590, N870);
xor XOR2 (N2522, N2507, N2496);
xor XOR2 (N2523, N2521, N599);
xor XOR2 (N2524, N2522, N1547);
xor XOR2 (N2525, N2509, N2395);
nand NAND3 (N2526, N2517, N995, N1069);
nand NAND3 (N2527, N2526, N2305, N1336);
nor NOR4 (N2528, N2524, N649, N840, N580);
nor NOR2 (N2529, N2528, N1795);
and AND2 (N2530, N2519, N407);
nand NAND3 (N2531, N2516, N1489, N839);
nor NOR3 (N2532, N2527, N1568, N364);
nor NOR2 (N2533, N2515, N1699);
buf BUF1 (N2534, N2523);
nor NOR4 (N2535, N2525, N1217, N1880, N566);
and AND2 (N2536, N2518, N895);
nand NAND2 (N2537, N2495, N712);
buf BUF1 (N2538, N2529);
nor NOR4 (N2539, N2537, N875, N199, N1665);
not NOT1 (N2540, N2520);
not NOT1 (N2541, N2536);
buf BUF1 (N2542, N2534);
nand NAND4 (N2543, N2531, N25, N1553, N906);
nand NAND4 (N2544, N2530, N21, N2375, N1347);
xor XOR2 (N2545, N2532, N616);
nand NAND4 (N2546, N2538, N1825, N334, N85);
or OR2 (N2547, N2544, N544);
not NOT1 (N2548, N2535);
or OR4 (N2549, N2548, N1740, N2228, N1085);
and AND2 (N2550, N2546, N508);
nand NAND2 (N2551, N2540, N1469);
and AND3 (N2552, N2533, N1813, N122);
nand NAND3 (N2553, N2552, N20, N1873);
buf BUF1 (N2554, N2542);
and AND2 (N2555, N2547, N570);
nor NOR4 (N2556, N2550, N579, N942, N2083);
xor XOR2 (N2557, N2539, N365);
xor XOR2 (N2558, N2543, N393);
buf BUF1 (N2559, N2549);
or OR2 (N2560, N2558, N432);
or OR2 (N2561, N2556, N2495);
or OR2 (N2562, N2560, N2281);
and AND2 (N2563, N2545, N68);
nor NOR2 (N2564, N2541, N1460);
and AND2 (N2565, N2554, N2482);
nor NOR3 (N2566, N2564, N578, N2363);
and AND2 (N2567, N2565, N1045);
nor NOR3 (N2568, N2566, N704, N1587);
not NOT1 (N2569, N2553);
nor NOR4 (N2570, N2562, N1138, N2482, N2506);
xor XOR2 (N2571, N2555, N451);
buf BUF1 (N2572, N2569);
buf BUF1 (N2573, N2551);
and AND3 (N2574, N2557, N1100, N1326);
not NOT1 (N2575, N2571);
not NOT1 (N2576, N2563);
xor XOR2 (N2577, N2575, N966);
or OR2 (N2578, N2572, N2196);
nand NAND4 (N2579, N2567, N2000, N158, N1061);
buf BUF1 (N2580, N2573);
buf BUF1 (N2581, N2570);
xor XOR2 (N2582, N2577, N1621);
nor NOR2 (N2583, N2578, N984);
and AND3 (N2584, N2568, N205, N2195);
and AND2 (N2585, N2579, N2449);
and AND3 (N2586, N2582, N2277, N1961);
nand NAND2 (N2587, N2581, N186);
xor XOR2 (N2588, N2574, N544);
nor NOR2 (N2589, N2583, N33);
not NOT1 (N2590, N2580);
nand NAND3 (N2591, N2559, N1830, N830);
and AND2 (N2592, N2584, N2240);
not NOT1 (N2593, N2588);
xor XOR2 (N2594, N2593, N548);
not NOT1 (N2595, N2587);
buf BUF1 (N2596, N2561);
nand NAND2 (N2597, N2596, N1221);
buf BUF1 (N2598, N2595);
not NOT1 (N2599, N2598);
not NOT1 (N2600, N2591);
and AND2 (N2601, N2592, N1290);
xor XOR2 (N2602, N2594, N725);
xor XOR2 (N2603, N2602, N2120);
and AND3 (N2604, N2590, N874, N1292);
nor NOR2 (N2605, N2597, N2584);
and AND4 (N2606, N2601, N1637, N478, N784);
and AND2 (N2607, N2589, N623);
nand NAND2 (N2608, N2600, N110);
or OR4 (N2609, N2599, N1527, N1323, N268);
not NOT1 (N2610, N2608);
buf BUF1 (N2611, N2576);
or OR4 (N2612, N2610, N2244, N1936, N1496);
buf BUF1 (N2613, N2606);
and AND3 (N2614, N2585, N1023, N663);
nor NOR2 (N2615, N2613, N1027);
buf BUF1 (N2616, N2603);
xor XOR2 (N2617, N2605, N2379);
or OR2 (N2618, N2604, N4);
buf BUF1 (N2619, N2616);
buf BUF1 (N2620, N2586);
and AND2 (N2621, N2612, N2458);
or OR3 (N2622, N2609, N546, N300);
and AND4 (N2623, N2619, N1468, N1246, N2523);
not NOT1 (N2624, N2617);
buf BUF1 (N2625, N2618);
nand NAND3 (N2626, N2623, N1575, N247);
nand NAND2 (N2627, N2626, N1672);
xor XOR2 (N2628, N2607, N2608);
or OR3 (N2629, N2615, N683, N2473);
buf BUF1 (N2630, N2625);
nand NAND3 (N2631, N2627, N405, N2497);
nand NAND3 (N2632, N2628, N239, N503);
nand NAND4 (N2633, N2631, N2570, N475, N50);
buf BUF1 (N2634, N2633);
not NOT1 (N2635, N2620);
nand NAND3 (N2636, N2611, N263, N1881);
not NOT1 (N2637, N2634);
xor XOR2 (N2638, N2621, N1595);
nand NAND2 (N2639, N2624, N1866);
xor XOR2 (N2640, N2614, N169);
nor NOR4 (N2641, N2635, N1921, N1332, N537);
nand NAND3 (N2642, N2640, N2036, N685);
xor XOR2 (N2643, N2622, N1134);
and AND3 (N2644, N2632, N1087, N1001);
or OR3 (N2645, N2643, N1839, N722);
nor NOR3 (N2646, N2638, N1740, N79);
nor NOR3 (N2647, N2644, N2419, N2198);
nor NOR3 (N2648, N2637, N509, N2454);
and AND2 (N2649, N2641, N118);
nor NOR3 (N2650, N2629, N2305, N587);
not NOT1 (N2651, N2645);
or OR4 (N2652, N2646, N1546, N1568, N2514);
nand NAND3 (N2653, N2642, N804, N1492);
nand NAND3 (N2654, N2653, N1465, N2577);
buf BUF1 (N2655, N2630);
buf BUF1 (N2656, N2648);
xor XOR2 (N2657, N2647, N1051);
not NOT1 (N2658, N2651);
not NOT1 (N2659, N2658);
xor XOR2 (N2660, N2636, N676);
xor XOR2 (N2661, N2639, N1252);
xor XOR2 (N2662, N2650, N1126);
nor NOR4 (N2663, N2654, N2396, N1447, N440);
nor NOR4 (N2664, N2663, N2282, N114, N1879);
or OR2 (N2665, N2659, N2093);
xor XOR2 (N2666, N2661, N700);
nand NAND2 (N2667, N2666, N2323);
not NOT1 (N2668, N2665);
or OR2 (N2669, N2649, N2609);
buf BUF1 (N2670, N2660);
nand NAND3 (N2671, N2652, N850, N1519);
nand NAND4 (N2672, N2669, N2085, N2185, N1924);
not NOT1 (N2673, N2670);
buf BUF1 (N2674, N2667);
or OR4 (N2675, N2674, N2025, N1559, N2492);
nor NOR4 (N2676, N2662, N1992, N1625, N2414);
not NOT1 (N2677, N2657);
and AND4 (N2678, N2677, N2516, N393, N1412);
nor NOR4 (N2679, N2664, N1305, N1510, N178);
buf BUF1 (N2680, N2672);
nor NOR4 (N2681, N2655, N1380, N2391, N149);
buf BUF1 (N2682, N2679);
nor NOR3 (N2683, N2678, N1114, N1077);
nor NOR3 (N2684, N2673, N1293, N1053);
and AND4 (N2685, N2682, N1821, N959, N1353);
nand NAND3 (N2686, N2676, N1114, N765);
xor XOR2 (N2687, N2671, N596);
and AND3 (N2688, N2675, N213, N1187);
or OR4 (N2689, N2688, N555, N988, N1492);
or OR4 (N2690, N2685, N1469, N553, N2150);
xor XOR2 (N2691, N2684, N1722);
or OR4 (N2692, N2656, N1958, N226, N330);
buf BUF1 (N2693, N2686);
and AND4 (N2694, N2692, N335, N2470, N356);
nand NAND4 (N2695, N2690, N1693, N2544, N2156);
or OR2 (N2696, N2693, N738);
nor NOR4 (N2697, N2689, N1959, N802, N310);
xor XOR2 (N2698, N2683, N361);
xor XOR2 (N2699, N2695, N657);
buf BUF1 (N2700, N2699);
buf BUF1 (N2701, N2696);
buf BUF1 (N2702, N2687);
buf BUF1 (N2703, N2681);
buf BUF1 (N2704, N2697);
and AND2 (N2705, N2700, N1988);
not NOT1 (N2706, N2701);
nor NOR2 (N2707, N2706, N2177);
or OR3 (N2708, N2691, N657, N2389);
not NOT1 (N2709, N2707);
xor XOR2 (N2710, N2694, N2008);
not NOT1 (N2711, N2705);
nand NAND3 (N2712, N2708, N1061, N2650);
not NOT1 (N2713, N2709);
buf BUF1 (N2714, N2702);
nor NOR2 (N2715, N2710, N414);
xor XOR2 (N2716, N2698, N386);
and AND4 (N2717, N2704, N122, N1791, N273);
nand NAND4 (N2718, N2713, N1070, N1677, N1515);
buf BUF1 (N2719, N2712);
nand NAND4 (N2720, N2680, N1607, N274, N330);
not NOT1 (N2721, N2668);
nor NOR3 (N2722, N2721, N473, N848);
xor XOR2 (N2723, N2716, N302);
xor XOR2 (N2724, N2717, N1090);
or OR2 (N2725, N2722, N1962);
xor XOR2 (N2726, N2720, N175);
nand NAND3 (N2727, N2726, N1376, N1316);
nand NAND4 (N2728, N2723, N353, N2151, N1147);
nor NOR3 (N2729, N2718, N536, N1719);
nor NOR4 (N2730, N2715, N2461, N569, N2474);
nor NOR2 (N2731, N2725, N1899);
not NOT1 (N2732, N2729);
nand NAND3 (N2733, N2731, N154, N400);
not NOT1 (N2734, N2714);
nor NOR2 (N2735, N2727, N1435);
nor NOR3 (N2736, N2732, N1504, N2124);
nand NAND2 (N2737, N2736, N2050);
not NOT1 (N2738, N2703);
xor XOR2 (N2739, N2734, N1484);
and AND4 (N2740, N2728, N2297, N72, N650);
xor XOR2 (N2741, N2737, N1870);
buf BUF1 (N2742, N2740);
and AND2 (N2743, N2741, N761);
nand NAND4 (N2744, N2739, N1622, N1722, N1452);
or OR2 (N2745, N2742, N528);
and AND2 (N2746, N2719, N1999);
not NOT1 (N2747, N2738);
and AND4 (N2748, N2711, N2050, N816, N702);
or OR4 (N2749, N2748, N2119, N348, N1874);
buf BUF1 (N2750, N2747);
xor XOR2 (N2751, N2750, N984);
nor NOR3 (N2752, N2730, N1149, N2443);
buf BUF1 (N2753, N2751);
not NOT1 (N2754, N2744);
buf BUF1 (N2755, N2745);
nand NAND4 (N2756, N2733, N2123, N1605, N590);
xor XOR2 (N2757, N2752, N1570);
nor NOR2 (N2758, N2756, N1300);
or OR2 (N2759, N2746, N1259);
nor NOR2 (N2760, N2757, N544);
nor NOR2 (N2761, N2755, N1122);
not NOT1 (N2762, N2754);
not NOT1 (N2763, N2760);
nor NOR3 (N2764, N2759, N115, N2715);
not NOT1 (N2765, N2763);
nand NAND4 (N2766, N2749, N491, N1190, N1195);
nor NOR3 (N2767, N2758, N560, N1908);
and AND2 (N2768, N2764, N917);
xor XOR2 (N2769, N2735, N2718);
xor XOR2 (N2770, N2765, N1870);
xor XOR2 (N2771, N2761, N1352);
and AND3 (N2772, N2769, N673, N2081);
and AND3 (N2773, N2767, N1611, N915);
not NOT1 (N2774, N2753);
buf BUF1 (N2775, N2771);
buf BUF1 (N2776, N2770);
buf BUF1 (N2777, N2775);
not NOT1 (N2778, N2724);
nor NOR2 (N2779, N2777, N384);
nand NAND4 (N2780, N2743, N822, N2771, N1823);
buf BUF1 (N2781, N2772);
xor XOR2 (N2782, N2768, N1412);
xor XOR2 (N2783, N2782, N1727);
or OR3 (N2784, N2776, N1064, N180);
not NOT1 (N2785, N2784);
and AND4 (N2786, N2762, N2158, N714, N2694);
xor XOR2 (N2787, N2783, N284);
nor NOR4 (N2788, N2781, N1468, N1067, N2724);
and AND4 (N2789, N2774, N1432, N2375, N852);
buf BUF1 (N2790, N2787);
or OR2 (N2791, N2785, N86);
and AND4 (N2792, N2786, N627, N2278, N914);
buf BUF1 (N2793, N2780);
xor XOR2 (N2794, N2779, N1401);
xor XOR2 (N2795, N2773, N434);
xor XOR2 (N2796, N2793, N256);
or OR3 (N2797, N2789, N108, N63);
or OR3 (N2798, N2791, N3, N2306);
buf BUF1 (N2799, N2796);
xor XOR2 (N2800, N2766, N1238);
xor XOR2 (N2801, N2797, N1993);
and AND4 (N2802, N2800, N1841, N2325, N2093);
or OR4 (N2803, N2792, N165, N1103, N1321);
nor NOR4 (N2804, N2790, N2233, N490, N1325);
and AND3 (N2805, N2778, N1256, N1460);
or OR3 (N2806, N2804, N700, N640);
not NOT1 (N2807, N2798);
nor NOR2 (N2808, N2806, N2536);
nand NAND3 (N2809, N2805, N940, N1788);
not NOT1 (N2810, N2803);
and AND4 (N2811, N2808, N113, N2096, N1087);
or OR2 (N2812, N2807, N2803);
nand NAND2 (N2813, N2788, N1450);
buf BUF1 (N2814, N2812);
xor XOR2 (N2815, N2799, N83);
xor XOR2 (N2816, N2794, N542);
xor XOR2 (N2817, N2809, N1667);
xor XOR2 (N2818, N2815, N2811);
buf BUF1 (N2819, N1442);
buf BUF1 (N2820, N2817);
nor NOR2 (N2821, N2801, N1200);
nand NAND3 (N2822, N2813, N370, N2434);
and AND2 (N2823, N2822, N456);
nor NOR3 (N2824, N2816, N2613, N2251);
xor XOR2 (N2825, N2823, N1602);
nand NAND2 (N2826, N2825, N2072);
nand NAND2 (N2827, N2810, N2117);
or OR2 (N2828, N2814, N1501);
nor NOR3 (N2829, N2821, N1642, N1207);
nor NOR2 (N2830, N2826, N1560);
nor NOR3 (N2831, N2820, N921, N1468);
and AND4 (N2832, N2818, N669, N2295, N2136);
buf BUF1 (N2833, N2830);
nand NAND4 (N2834, N2829, N1105, N1665, N198);
xor XOR2 (N2835, N2833, N592);
not NOT1 (N2836, N2824);
xor XOR2 (N2837, N2836, N2561);
nand NAND2 (N2838, N2834, N2577);
nand NAND2 (N2839, N2837, N2381);
nor NOR2 (N2840, N2802, N1352);
and AND2 (N2841, N2835, N287);
not NOT1 (N2842, N2839);
not NOT1 (N2843, N2828);
nand NAND3 (N2844, N2842, N2813, N213);
nor NOR2 (N2845, N2831, N185);
or OR2 (N2846, N2844, N170);
and AND3 (N2847, N2819, N1177, N336);
nor NOR3 (N2848, N2840, N654, N127);
not NOT1 (N2849, N2841);
or OR2 (N2850, N2847, N104);
nor NOR2 (N2851, N2827, N2484);
xor XOR2 (N2852, N2851, N578);
and AND2 (N2853, N2838, N1282);
not NOT1 (N2854, N2795);
not NOT1 (N2855, N2845);
and AND2 (N2856, N2848, N1993);
nor NOR3 (N2857, N2855, N1664, N681);
not NOT1 (N2858, N2857);
not NOT1 (N2859, N2853);
or OR4 (N2860, N2843, N663, N1177, N2162);
buf BUF1 (N2861, N2854);
nor NOR2 (N2862, N2861, N251);
buf BUF1 (N2863, N2860);
nand NAND4 (N2864, N2856, N2011, N1703, N2541);
or OR4 (N2865, N2859, N1365, N1682, N1131);
buf BUF1 (N2866, N2852);
buf BUF1 (N2867, N2846);
or OR4 (N2868, N2849, N1407, N533, N1281);
xor XOR2 (N2869, N2858, N324);
and AND3 (N2870, N2868, N560, N2151);
nor NOR2 (N2871, N2866, N2373);
not NOT1 (N2872, N2869);
xor XOR2 (N2873, N2862, N2710);
buf BUF1 (N2874, N2865);
not NOT1 (N2875, N2872);
not NOT1 (N2876, N2873);
or OR3 (N2877, N2874, N26, N1994);
nand NAND4 (N2878, N2832, N2467, N2250, N686);
and AND4 (N2879, N2875, N403, N619, N1104);
nand NAND2 (N2880, N2863, N366);
and AND2 (N2881, N2850, N2787);
nand NAND4 (N2882, N2879, N1372, N1315, N167);
and AND2 (N2883, N2871, N1968);
nor NOR3 (N2884, N2867, N59, N1861);
and AND2 (N2885, N2864, N1894);
not NOT1 (N2886, N2885);
not NOT1 (N2887, N2876);
nand NAND4 (N2888, N2887, N1691, N2882, N899);
not NOT1 (N2889, N2695);
nand NAND2 (N2890, N2881, N953);
nand NAND3 (N2891, N2877, N502, N1739);
buf BUF1 (N2892, N2870);
xor XOR2 (N2893, N2890, N1772);
not NOT1 (N2894, N2883);
and AND4 (N2895, N2886, N2337, N1517, N559);
not NOT1 (N2896, N2893);
xor XOR2 (N2897, N2896, N1368);
and AND4 (N2898, N2880, N2106, N31, N2791);
and AND2 (N2899, N2891, N551);
nor NOR3 (N2900, N2884, N2880, N1257);
xor XOR2 (N2901, N2894, N2207);
not NOT1 (N2902, N2892);
not NOT1 (N2903, N2898);
xor XOR2 (N2904, N2899, N1633);
not NOT1 (N2905, N2897);
nor NOR3 (N2906, N2904, N287, N1237);
and AND3 (N2907, N2903, N1655, N198);
nand NAND3 (N2908, N2901, N2827, N2493);
nor NOR3 (N2909, N2905, N2448, N947);
or OR2 (N2910, N2878, N2666);
buf BUF1 (N2911, N2907);
and AND2 (N2912, N2908, N2537);
xor XOR2 (N2913, N2906, N55);
not NOT1 (N2914, N2910);
nor NOR3 (N2915, N2911, N167, N2831);
nor NOR2 (N2916, N2888, N2083);
buf BUF1 (N2917, N2895);
nor NOR2 (N2918, N2913, N2313);
nor NOR4 (N2919, N2915, N1233, N635, N406);
buf BUF1 (N2920, N2900);
and AND4 (N2921, N2920, N1477, N2345, N1065);
not NOT1 (N2922, N2912);
buf BUF1 (N2923, N2916);
and AND4 (N2924, N2914, N1843, N789, N1323);
nor NOR3 (N2925, N2923, N2241, N636);
buf BUF1 (N2926, N2902);
buf BUF1 (N2927, N2926);
xor XOR2 (N2928, N2927, N2527);
nand NAND4 (N2929, N2922, N2910, N1816, N1302);
xor XOR2 (N2930, N2929, N599);
nand NAND4 (N2931, N2917, N2378, N670, N2889);
and AND2 (N2932, N391, N823);
nor NOR2 (N2933, N2931, N2812);
nor NOR3 (N2934, N2924, N1583, N191);
xor XOR2 (N2935, N2909, N1522);
xor XOR2 (N2936, N2933, N370);
nand NAND2 (N2937, N2925, N2516);
and AND3 (N2938, N2932, N575, N2276);
and AND2 (N2939, N2935, N2058);
not NOT1 (N2940, N2936);
nand NAND4 (N2941, N2940, N2695, N1966, N507);
nand NAND2 (N2942, N2928, N2552);
nand NAND4 (N2943, N2938, N353, N2504, N1983);
xor XOR2 (N2944, N2921, N625);
not NOT1 (N2945, N2937);
and AND2 (N2946, N2934, N202);
nand NAND2 (N2947, N2943, N1671);
nor NOR3 (N2948, N2939, N1595, N255);
nand NAND3 (N2949, N2942, N2002, N2002);
xor XOR2 (N2950, N2918, N1740);
nand NAND2 (N2951, N2948, N765);
xor XOR2 (N2952, N2949, N1449);
or OR4 (N2953, N2919, N2579, N693, N1454);
nand NAND4 (N2954, N2941, N2328, N1982, N384);
or OR4 (N2955, N2954, N2690, N2444, N2777);
buf BUF1 (N2956, N2944);
not NOT1 (N2957, N2946);
xor XOR2 (N2958, N2951, N2496);
and AND2 (N2959, N2945, N2587);
and AND3 (N2960, N2955, N1604, N1881);
or OR2 (N2961, N2953, N732);
not NOT1 (N2962, N2957);
buf BUF1 (N2963, N2958);
buf BUF1 (N2964, N2952);
nor NOR2 (N2965, N2962, N2849);
and AND2 (N2966, N2963, N2635);
nor NOR3 (N2967, N2965, N119, N553);
nor NOR2 (N2968, N2956, N2879);
nor NOR4 (N2969, N2966, N1051, N694, N1604);
xor XOR2 (N2970, N2959, N1334);
nand NAND3 (N2971, N2964, N1005, N2114);
or OR2 (N2972, N2947, N1253);
buf BUF1 (N2973, N2960);
not NOT1 (N2974, N2971);
nor NOR4 (N2975, N2968, N571, N2840, N1943);
or OR4 (N2976, N2930, N1356, N1601, N2109);
or OR3 (N2977, N2961, N1963, N2926);
or OR4 (N2978, N2975, N1998, N303, N70);
buf BUF1 (N2979, N2976);
or OR2 (N2980, N2972, N1908);
xor XOR2 (N2981, N2950, N2281);
nor NOR3 (N2982, N2979, N1678, N1767);
not NOT1 (N2983, N2970);
xor XOR2 (N2984, N2981, N1789);
not NOT1 (N2985, N2967);
xor XOR2 (N2986, N2969, N2139);
nor NOR3 (N2987, N2974, N341, N2422);
xor XOR2 (N2988, N2985, N478);
nand NAND4 (N2989, N2980, N2395, N710, N1171);
not NOT1 (N2990, N2987);
or OR4 (N2991, N2982, N2941, N1877, N2083);
nor NOR3 (N2992, N2988, N149, N1761);
not NOT1 (N2993, N2989);
buf BUF1 (N2994, N2983);
nor NOR4 (N2995, N2986, N703, N531, N1553);
not NOT1 (N2996, N2973);
buf BUF1 (N2997, N2977);
buf BUF1 (N2998, N2992);
buf BUF1 (N2999, N2994);
nor NOR3 (N3000, N2999, N524, N676);
or OR2 (N3001, N3000, N2876);
and AND3 (N3002, N2984, N526, N2380);
xor XOR2 (N3003, N3001, N2282);
nand NAND2 (N3004, N2998, N2772);
buf BUF1 (N3005, N2991);
nor NOR4 (N3006, N3002, N2313, N1167, N1012);
xor XOR2 (N3007, N2978, N1220);
xor XOR2 (N3008, N2993, N532);
xor XOR2 (N3009, N2995, N1040);
not NOT1 (N3010, N2996);
not NOT1 (N3011, N3008);
nand NAND4 (N3012, N3006, N843, N1434, N526);
xor XOR2 (N3013, N2997, N1934);
xor XOR2 (N3014, N3013, N922);
nor NOR4 (N3015, N3011, N2827, N1550, N1672);
buf BUF1 (N3016, N3007);
or OR2 (N3017, N3003, N935);
nor NOR3 (N3018, N2990, N808, N2626);
and AND2 (N3019, N3018, N877);
xor XOR2 (N3020, N3019, N752);
or OR4 (N3021, N3009, N115, N741, N2325);
xor XOR2 (N3022, N3020, N574);
and AND3 (N3023, N3016, N845, N269);
or OR2 (N3024, N3012, N583);
nor NOR4 (N3025, N3015, N1976, N1320, N1368);
or OR2 (N3026, N3005, N549);
nand NAND2 (N3027, N3014, N2687);
xor XOR2 (N3028, N3004, N1827);
or OR2 (N3029, N3028, N2291);
nand NAND2 (N3030, N3017, N1638);
nor NOR4 (N3031, N3030, N48, N1402, N2732);
not NOT1 (N3032, N3031);
or OR3 (N3033, N3025, N1335, N3018);
xor XOR2 (N3034, N3027, N2917);
not NOT1 (N3035, N3021);
not NOT1 (N3036, N3032);
not NOT1 (N3037, N3023);
and AND2 (N3038, N3034, N868);
not NOT1 (N3039, N3038);
not NOT1 (N3040, N3029);
buf BUF1 (N3041, N3037);
or OR2 (N3042, N3022, N2423);
buf BUF1 (N3043, N3039);
xor XOR2 (N3044, N3035, N2751);
or OR2 (N3045, N3043, N2613);
nand NAND3 (N3046, N3040, N742, N207);
and AND4 (N3047, N3042, N2030, N17, N2314);
xor XOR2 (N3048, N3045, N2966);
and AND2 (N3049, N3041, N2336);
not NOT1 (N3050, N3047);
or OR2 (N3051, N3033, N118);
nand NAND4 (N3052, N3051, N1994, N1686, N2720);
or OR2 (N3053, N3026, N2011);
not NOT1 (N3054, N3024);
nand NAND3 (N3055, N3054, N468, N2706);
not NOT1 (N3056, N3048);
nand NAND3 (N3057, N3055, N1773, N1721);
or OR4 (N3058, N3052, N2898, N1697, N1084);
or OR4 (N3059, N3058, N1790, N942, N24);
nand NAND2 (N3060, N3036, N1671);
or OR2 (N3061, N3010, N467);
or OR2 (N3062, N3057, N1212);
buf BUF1 (N3063, N3059);
nand NAND2 (N3064, N3053, N1843);
nand NAND2 (N3065, N3064, N449);
or OR3 (N3066, N3044, N1273, N227);
nand NAND4 (N3067, N3046, N592, N876, N3060);
nand NAND3 (N3068, N154, N2033, N1691);
nand NAND3 (N3069, N3065, N594, N2255);
buf BUF1 (N3070, N3050);
not NOT1 (N3071, N3069);
nor NOR2 (N3072, N3063, N657);
nor NOR4 (N3073, N3056, N1901, N1345, N2404);
nor NOR2 (N3074, N3061, N1378);
and AND3 (N3075, N3073, N2262, N838);
and AND4 (N3076, N3071, N2907, N1705, N3);
nor NOR3 (N3077, N3076, N719, N1507);
and AND4 (N3078, N3062, N1396, N1343, N1387);
nand NAND4 (N3079, N3068, N173, N2809, N96);
nor NOR2 (N3080, N3079, N1976);
xor XOR2 (N3081, N3075, N1052);
buf BUF1 (N3082, N3077);
nor NOR4 (N3083, N3080, N811, N2720, N1422);
not NOT1 (N3084, N3081);
nor NOR3 (N3085, N3082, N3046, N1100);
nor NOR3 (N3086, N3084, N253, N2661);
or OR4 (N3087, N3085, N3042, N1328, N1090);
buf BUF1 (N3088, N3074);
nor NOR4 (N3089, N3087, N1028, N2410, N1123);
buf BUF1 (N3090, N3083);
xor XOR2 (N3091, N3090, N1329);
nand NAND4 (N3092, N3088, N1280, N235, N717);
xor XOR2 (N3093, N3067, N515);
and AND3 (N3094, N3091, N526, N1106);
nand NAND3 (N3095, N3094, N3055, N2889);
xor XOR2 (N3096, N3095, N1301);
or OR3 (N3097, N3049, N2114, N2403);
not NOT1 (N3098, N3086);
xor XOR2 (N3099, N3089, N1474);
nand NAND2 (N3100, N3070, N1661);
buf BUF1 (N3101, N3093);
xor XOR2 (N3102, N3098, N2851);
xor XOR2 (N3103, N3078, N171);
not NOT1 (N3104, N3101);
nand NAND2 (N3105, N3104, N3002);
nand NAND2 (N3106, N3100, N3099);
nand NAND3 (N3107, N2488, N754, N79);
and AND4 (N3108, N3105, N687, N63, N1310);
or OR3 (N3109, N3106, N1152, N3028);
not NOT1 (N3110, N3072);
buf BUF1 (N3111, N3107);
buf BUF1 (N3112, N3096);
nor NOR4 (N3113, N3109, N2481, N2747, N2424);
and AND2 (N3114, N3112, N2218);
nand NAND2 (N3115, N3113, N974);
buf BUF1 (N3116, N3066);
xor XOR2 (N3117, N3102, N1959);
xor XOR2 (N3118, N3097, N2361);
nor NOR4 (N3119, N3111, N2222, N2614, N305);
nand NAND4 (N3120, N3103, N607, N31, N883);
xor XOR2 (N3121, N3108, N1680);
not NOT1 (N3122, N3120);
nand NAND2 (N3123, N3122, N2917);
xor XOR2 (N3124, N3115, N1360);
xor XOR2 (N3125, N3110, N2144);
and AND3 (N3126, N3117, N2891, N1998);
or OR3 (N3127, N3121, N955, N2924);
or OR3 (N3128, N3114, N2855, N1675);
nor NOR4 (N3129, N3123, N1073, N2530, N2);
xor XOR2 (N3130, N3119, N2484);
xor XOR2 (N3131, N3127, N2586);
buf BUF1 (N3132, N3116);
nor NOR4 (N3133, N3125, N965, N2417, N161);
and AND3 (N3134, N3128, N734, N1987);
nor NOR4 (N3135, N3131, N933, N2032, N333);
not NOT1 (N3136, N3092);
xor XOR2 (N3137, N3135, N1867);
not NOT1 (N3138, N3124);
and AND2 (N3139, N3129, N2874);
or OR4 (N3140, N3138, N380, N2289, N190);
not NOT1 (N3141, N3140);
and AND3 (N3142, N3126, N652, N960);
not NOT1 (N3143, N3141);
buf BUF1 (N3144, N3132);
nor NOR4 (N3145, N3130, N1380, N1098, N2444);
buf BUF1 (N3146, N3136);
nor NOR4 (N3147, N3133, N2446, N324, N1771);
or OR4 (N3148, N3134, N2505, N208, N2055);
nand NAND4 (N3149, N3142, N1329, N3064, N3126);
nor NOR2 (N3150, N3146, N994);
xor XOR2 (N3151, N3144, N1468);
or OR3 (N3152, N3137, N1156, N762);
buf BUF1 (N3153, N3148);
xor XOR2 (N3154, N3139, N2783);
nor NOR2 (N3155, N3118, N2332);
nand NAND3 (N3156, N3149, N1910, N2802);
buf BUF1 (N3157, N3156);
not NOT1 (N3158, N3143);
not NOT1 (N3159, N3147);
or OR2 (N3160, N3158, N898);
nor NOR2 (N3161, N3160, N1499);
and AND3 (N3162, N3145, N1587, N1646);
or OR4 (N3163, N3154, N370, N2223, N2797);
nand NAND4 (N3164, N3159, N2699, N812, N3000);
nor NOR2 (N3165, N3164, N1698);
xor XOR2 (N3166, N3162, N447);
nand NAND3 (N3167, N3152, N2887, N614);
nand NAND4 (N3168, N3167, N1122, N477, N3095);
nor NOR4 (N3169, N3157, N500, N175, N2538);
buf BUF1 (N3170, N3169);
buf BUF1 (N3171, N3166);
not NOT1 (N3172, N3155);
and AND2 (N3173, N3163, N1758);
xor XOR2 (N3174, N3150, N212);
and AND3 (N3175, N3172, N2883, N907);
and AND2 (N3176, N3153, N1005);
or OR4 (N3177, N3173, N218, N911, N800);
nor NOR4 (N3178, N3174, N90, N520, N1194);
nand NAND2 (N3179, N3168, N1923);
or OR4 (N3180, N3178, N519, N2278, N2806);
buf BUF1 (N3181, N3176);
buf BUF1 (N3182, N3180);
nor NOR3 (N3183, N3170, N995, N3049);
and AND3 (N3184, N3161, N1577, N1428);
or OR4 (N3185, N3175, N3097, N2198, N378);
and AND4 (N3186, N3177, N1855, N519, N3136);
and AND3 (N3187, N3185, N2451, N2571);
xor XOR2 (N3188, N3165, N1674);
or OR4 (N3189, N3186, N1903, N2963, N2269);
buf BUF1 (N3190, N3151);
nor NOR2 (N3191, N3183, N227);
xor XOR2 (N3192, N3187, N1656);
buf BUF1 (N3193, N3179);
buf BUF1 (N3194, N3191);
or OR4 (N3195, N3193, N123, N2891, N3029);
not NOT1 (N3196, N3184);
nand NAND4 (N3197, N3171, N2732, N1201, N2191);
or OR2 (N3198, N3181, N3120);
and AND4 (N3199, N3188, N2882, N2457, N1907);
and AND3 (N3200, N3197, N1907, N2591);
or OR3 (N3201, N3192, N2490, N2409);
xor XOR2 (N3202, N3196, N1668);
and AND3 (N3203, N3190, N431, N2658);
not NOT1 (N3204, N3195);
nand NAND4 (N3205, N3182, N2546, N1861, N18);
buf BUF1 (N3206, N3205);
not NOT1 (N3207, N3199);
nand NAND2 (N3208, N3203, N1020);
not NOT1 (N3209, N3206);
and AND2 (N3210, N3189, N1298);
buf BUF1 (N3211, N3200);
not NOT1 (N3212, N3194);
buf BUF1 (N3213, N3198);
nor NOR3 (N3214, N3202, N3164, N2163);
nor NOR2 (N3215, N3213, N3185);
buf BUF1 (N3216, N3207);
nand NAND2 (N3217, N3216, N1500);
xor XOR2 (N3218, N3201, N1287);
nand NAND4 (N3219, N3215, N2247, N2180, N2504);
and AND2 (N3220, N3209, N3004);
xor XOR2 (N3221, N3214, N1401);
or OR3 (N3222, N3208, N928, N2969);
nand NAND3 (N3223, N3210, N2909, N2670);
not NOT1 (N3224, N3218);
not NOT1 (N3225, N3217);
or OR2 (N3226, N3221, N702);
nand NAND4 (N3227, N3220, N1244, N1181, N2473);
and AND2 (N3228, N3224, N2432);
buf BUF1 (N3229, N3219);
and AND4 (N3230, N3228, N1480, N1232, N93);
not NOT1 (N3231, N3211);
xor XOR2 (N3232, N3204, N289);
or OR3 (N3233, N3212, N2010, N2183);
nor NOR4 (N3234, N3223, N108, N3225, N2053);
nand NAND4 (N3235, N1295, N2249, N2126, N290);
xor XOR2 (N3236, N3233, N2795);
xor XOR2 (N3237, N3227, N2815);
xor XOR2 (N3238, N3232, N1178);
or OR2 (N3239, N3229, N2110);
not NOT1 (N3240, N3236);
and AND4 (N3241, N3235, N3169, N2077, N1950);
and AND4 (N3242, N3241, N2852, N254, N2031);
buf BUF1 (N3243, N3238);
nor NOR4 (N3244, N3242, N2872, N2154, N118);
and AND3 (N3245, N3230, N125, N3203);
not NOT1 (N3246, N3231);
xor XOR2 (N3247, N3234, N426);
nor NOR3 (N3248, N3247, N2723, N1902);
or OR3 (N3249, N3239, N2272, N1596);
and AND3 (N3250, N3226, N1371, N350);
and AND4 (N3251, N3246, N1567, N2958, N293);
nand NAND2 (N3252, N3250, N1629);
or OR3 (N3253, N3251, N1637, N2569);
or OR3 (N3254, N3249, N1944, N1041);
and AND3 (N3255, N3237, N806, N22);
not NOT1 (N3256, N3245);
and AND4 (N3257, N3243, N3074, N2518, N116);
and AND4 (N3258, N3244, N874, N506, N2960);
or OR4 (N3259, N3254, N2937, N1288, N1570);
nor NOR2 (N3260, N3257, N883);
xor XOR2 (N3261, N3222, N2022);
nor NOR4 (N3262, N3255, N2627, N889, N3205);
and AND3 (N3263, N3253, N2788, N2332);
and AND3 (N3264, N3262, N3021, N2345);
buf BUF1 (N3265, N3256);
not NOT1 (N3266, N3260);
xor XOR2 (N3267, N3248, N2237);
xor XOR2 (N3268, N3261, N2741);
not NOT1 (N3269, N3240);
nand NAND3 (N3270, N3252, N2059, N129);
nor NOR2 (N3271, N3263, N700);
nand NAND4 (N3272, N3269, N2325, N149, N2181);
nand NAND4 (N3273, N3267, N3190, N424, N3130);
xor XOR2 (N3274, N3259, N1325);
nor NOR4 (N3275, N3271, N1724, N2970, N2924);
or OR3 (N3276, N3264, N33, N3144);
and AND2 (N3277, N3274, N2942);
nor NOR3 (N3278, N3276, N3001, N1563);
nand NAND4 (N3279, N3258, N2950, N2754, N2446);
not NOT1 (N3280, N3268);
buf BUF1 (N3281, N3266);
nor NOR4 (N3282, N3272, N2730, N870, N3238);
or OR4 (N3283, N3277, N1872, N496, N2938);
or OR4 (N3284, N3281, N2903, N1396, N2751);
buf BUF1 (N3285, N3270);
and AND3 (N3286, N3282, N2143, N2027);
or OR3 (N3287, N3275, N2448, N1825);
buf BUF1 (N3288, N3284);
and AND2 (N3289, N3280, N1834);
nor NOR4 (N3290, N3278, N631, N610, N44);
xor XOR2 (N3291, N3283, N19);
buf BUF1 (N3292, N3285);
or OR2 (N3293, N3279, N578);
not NOT1 (N3294, N3273);
not NOT1 (N3295, N3291);
buf BUF1 (N3296, N3290);
not NOT1 (N3297, N3292);
xor XOR2 (N3298, N3294, N2944);
xor XOR2 (N3299, N3265, N1230);
and AND4 (N3300, N3288, N3243, N1659, N3116);
or OR3 (N3301, N3297, N2670, N1422);
nor NOR2 (N3302, N3301, N2505);
buf BUF1 (N3303, N3286);
and AND4 (N3304, N3303, N1760, N779, N2836);
buf BUF1 (N3305, N3299);
xor XOR2 (N3306, N3287, N2510);
and AND4 (N3307, N3305, N2800, N2236, N2825);
or OR3 (N3308, N3306, N2295, N1763);
nor NOR2 (N3309, N3298, N184);
or OR3 (N3310, N3295, N1712, N2518);
nand NAND2 (N3311, N3293, N58);
nor NOR2 (N3312, N3300, N989);
nand NAND3 (N3313, N3304, N2795, N2192);
xor XOR2 (N3314, N3309, N1733);
buf BUF1 (N3315, N3296);
or OR3 (N3316, N3302, N1230, N1428);
or OR2 (N3317, N3308, N2821);
or OR2 (N3318, N3307, N1850);
nand NAND4 (N3319, N3318, N3227, N147, N694);
not NOT1 (N3320, N3310);
buf BUF1 (N3321, N3317);
nand NAND4 (N3322, N3319, N2481, N1790, N400);
nand NAND4 (N3323, N3315, N2032, N3309, N954);
or OR4 (N3324, N3312, N2498, N2704, N2600);
xor XOR2 (N3325, N3322, N921);
xor XOR2 (N3326, N3314, N1308);
or OR2 (N3327, N3321, N2583);
nor NOR4 (N3328, N3324, N3130, N431, N815);
or OR2 (N3329, N3327, N2944);
buf BUF1 (N3330, N3326);
buf BUF1 (N3331, N3313);
nand NAND2 (N3332, N3316, N2849);
nor NOR3 (N3333, N3323, N2977, N1483);
nor NOR3 (N3334, N3289, N2213, N1106);
nor NOR3 (N3335, N3333, N2723, N1034);
not NOT1 (N3336, N3335);
not NOT1 (N3337, N3328);
nor NOR4 (N3338, N3330, N2911, N928, N737);
and AND4 (N3339, N3331, N2287, N1882, N2434);
nor NOR3 (N3340, N3325, N2551, N1489);
nand NAND4 (N3341, N3311, N1905, N846, N1389);
nor NOR4 (N3342, N3340, N1548, N3263, N2663);
nand NAND3 (N3343, N3332, N1006, N2010);
nand NAND2 (N3344, N3320, N2047);
not NOT1 (N3345, N3329);
nor NOR2 (N3346, N3345, N2715);
nor NOR2 (N3347, N3341, N54);
nor NOR2 (N3348, N3336, N838);
or OR4 (N3349, N3346, N3278, N3130, N1870);
nand NAND4 (N3350, N3349, N284, N3344, N640);
or OR3 (N3351, N1348, N848, N921);
nand NAND4 (N3352, N3339, N1088, N2293, N2017);
nand NAND2 (N3353, N3352, N1633);
or OR3 (N3354, N3353, N842, N68);
or OR2 (N3355, N3343, N1710);
buf BUF1 (N3356, N3355);
xor XOR2 (N3357, N3354, N274);
xor XOR2 (N3358, N3347, N2474);
nor NOR4 (N3359, N3351, N329, N2369, N886);
not NOT1 (N3360, N3342);
buf BUF1 (N3361, N3359);
buf BUF1 (N3362, N3350);
or OR2 (N3363, N3337, N851);
nand NAND2 (N3364, N3361, N1349);
not NOT1 (N3365, N3356);
nand NAND2 (N3366, N3365, N1789);
nand NAND4 (N3367, N3348, N3256, N1982, N2192);
not NOT1 (N3368, N3334);
not NOT1 (N3369, N3357);
or OR3 (N3370, N3358, N2890, N1133);
xor XOR2 (N3371, N3364, N2411);
or OR4 (N3372, N3338, N2674, N2082, N2229);
not NOT1 (N3373, N3366);
nand NAND3 (N3374, N3373, N2163, N3187);
or OR4 (N3375, N3370, N2572, N1462, N2342);
buf BUF1 (N3376, N3360);
buf BUF1 (N3377, N3368);
or OR2 (N3378, N3363, N1333);
and AND3 (N3379, N3362, N3139, N564);
and AND4 (N3380, N3378, N831, N567, N2112);
and AND2 (N3381, N3375, N464);
nor NOR2 (N3382, N3369, N353);
nand NAND2 (N3383, N3372, N1784);
xor XOR2 (N3384, N3381, N2644);
not NOT1 (N3385, N3384);
and AND4 (N3386, N3379, N2012, N2428, N406);
buf BUF1 (N3387, N3380);
nand NAND4 (N3388, N3371, N2125, N2106, N3294);
nor NOR4 (N3389, N3367, N2141, N698, N532);
buf BUF1 (N3390, N3389);
or OR4 (N3391, N3387, N3221, N3207, N2746);
or OR3 (N3392, N3377, N467, N2729);
and AND4 (N3393, N3391, N451, N1919, N1590);
xor XOR2 (N3394, N3388, N2705);
xor XOR2 (N3395, N3383, N1137);
nand NAND2 (N3396, N3392, N1094);
buf BUF1 (N3397, N3385);
nand NAND3 (N3398, N3397, N2639, N3056);
and AND4 (N3399, N3394, N770, N2988, N838);
xor XOR2 (N3400, N3393, N3395);
and AND2 (N3401, N3374, N1879);
not NOT1 (N3402, N3130);
nor NOR2 (N3403, N3382, N894);
not NOT1 (N3404, N3401);
or OR4 (N3405, N3390, N802, N1726, N957);
xor XOR2 (N3406, N3386, N440);
nor NOR3 (N3407, N3403, N2128, N1169);
buf BUF1 (N3408, N3399);
and AND3 (N3409, N3404, N3136, N201);
buf BUF1 (N3410, N3402);
or OR2 (N3411, N3405, N9);
nand NAND4 (N3412, N3396, N3196, N1071, N2092);
nand NAND3 (N3413, N3406, N93, N2306);
nand NAND2 (N3414, N3408, N297);
or OR4 (N3415, N3409, N1425, N2299, N2577);
and AND3 (N3416, N3410, N963, N1965);
buf BUF1 (N3417, N3412);
or OR4 (N3418, N3398, N2206, N864, N4);
nand NAND4 (N3419, N3407, N2306, N1531, N2703);
nor NOR3 (N3420, N3400, N1804, N722);
buf BUF1 (N3421, N3418);
nor NOR2 (N3422, N3421, N1139);
and AND4 (N3423, N3411, N2432, N1697, N3193);
or OR4 (N3424, N3417, N480, N1552, N1611);
xor XOR2 (N3425, N3420, N2420);
not NOT1 (N3426, N3425);
and AND3 (N3427, N3414, N1093, N1730);
or OR2 (N3428, N3376, N1701);
not NOT1 (N3429, N3413);
buf BUF1 (N3430, N3426);
buf BUF1 (N3431, N3427);
nand NAND3 (N3432, N3419, N409, N3266);
nand NAND4 (N3433, N3422, N3071, N1496, N3113);
nand NAND2 (N3434, N3431, N2762);
buf BUF1 (N3435, N3416);
xor XOR2 (N3436, N3423, N1868);
not NOT1 (N3437, N3433);
nand NAND3 (N3438, N3428, N1160, N1211);
or OR2 (N3439, N3429, N1098);
nand NAND2 (N3440, N3424, N1266);
and AND3 (N3441, N3430, N2845, N2414);
and AND3 (N3442, N3439, N2657, N1715);
not NOT1 (N3443, N3434);
nor NOR3 (N3444, N3432, N2931, N2458);
and AND2 (N3445, N3415, N730);
nand NAND3 (N3446, N3440, N2275, N1491);
nand NAND4 (N3447, N3444, N1423, N3284, N574);
nand NAND3 (N3448, N3447, N3270, N1610);
buf BUF1 (N3449, N3443);
or OR3 (N3450, N3445, N323, N198);
xor XOR2 (N3451, N3449, N216);
and AND4 (N3452, N3448, N1671, N1198, N1455);
or OR2 (N3453, N3450, N3177);
not NOT1 (N3454, N3438);
nor NOR2 (N3455, N3436, N984);
and AND2 (N3456, N3442, N1635);
or OR4 (N3457, N3453, N967, N486, N2657);
and AND3 (N3458, N3456, N2967, N765);
nor NOR3 (N3459, N3452, N1355, N2311);
not NOT1 (N3460, N3458);
not NOT1 (N3461, N3441);
xor XOR2 (N3462, N3437, N3201);
not NOT1 (N3463, N3461);
not NOT1 (N3464, N3455);
nand NAND3 (N3465, N3463, N853, N1397);
nor NOR3 (N3466, N3464, N3015, N2223);
not NOT1 (N3467, N3462);
buf BUF1 (N3468, N3467);
and AND2 (N3469, N3446, N61);
and AND2 (N3470, N3457, N621);
or OR3 (N3471, N3454, N439, N887);
or OR2 (N3472, N3466, N3351);
not NOT1 (N3473, N3460);
nor NOR4 (N3474, N3435, N2222, N3081, N2471);
and AND3 (N3475, N3468, N2090, N733);
xor XOR2 (N3476, N3459, N1646);
and AND4 (N3477, N3470, N2046, N367, N1144);
nand NAND2 (N3478, N3465, N22);
nor NOR2 (N3479, N3474, N1246);
or OR2 (N3480, N3473, N3153);
nor NOR4 (N3481, N3478, N1514, N729, N209);
buf BUF1 (N3482, N3476);
not NOT1 (N3483, N3481);
not NOT1 (N3484, N3483);
and AND3 (N3485, N3477, N2358, N1985);
or OR3 (N3486, N3471, N641, N681);
and AND3 (N3487, N3482, N1566, N1864);
xor XOR2 (N3488, N3475, N1893);
buf BUF1 (N3489, N3485);
nand NAND3 (N3490, N3484, N196, N3061);
nor NOR3 (N3491, N3486, N97, N602);
nand NAND3 (N3492, N3479, N2149, N1394);
or OR3 (N3493, N3489, N8, N2562);
buf BUF1 (N3494, N3490);
xor XOR2 (N3495, N3488, N935);
buf BUF1 (N3496, N3495);
nor NOR3 (N3497, N3491, N24, N787);
nor NOR3 (N3498, N3497, N257, N2988);
not NOT1 (N3499, N3492);
buf BUF1 (N3500, N3494);
nand NAND2 (N3501, N3480, N3118);
nand NAND4 (N3502, N3496, N1822, N1178, N1700);
xor XOR2 (N3503, N3501, N3256);
nor NOR3 (N3504, N3469, N355, N398);
nand NAND4 (N3505, N3500, N590, N1763, N344);
buf BUF1 (N3506, N3505);
buf BUF1 (N3507, N3487);
nor NOR2 (N3508, N3451, N2424);
and AND4 (N3509, N3502, N531, N789, N1240);
or OR4 (N3510, N3507, N1067, N2376, N1674);
nand NAND2 (N3511, N3509, N2147);
not NOT1 (N3512, N3503);
or OR4 (N3513, N3493, N3203, N2898, N2379);
buf BUF1 (N3514, N3511);
or OR2 (N3515, N3472, N3423);
xor XOR2 (N3516, N3513, N1185);
and AND4 (N3517, N3514, N2373, N2670, N329);
xor XOR2 (N3518, N3515, N70);
buf BUF1 (N3519, N3506);
and AND3 (N3520, N3519, N2700, N687);
nand NAND4 (N3521, N3498, N3513, N1669, N741);
nand NAND4 (N3522, N3518, N1159, N949, N907);
buf BUF1 (N3523, N3520);
nor NOR2 (N3524, N3521, N187);
buf BUF1 (N3525, N3524);
or OR4 (N3526, N3525, N998, N2427, N2958);
nor NOR3 (N3527, N3512, N2981, N1124);
nor NOR2 (N3528, N3526, N1289);
buf BUF1 (N3529, N3508);
and AND3 (N3530, N3510, N2909, N3360);
or OR2 (N3531, N3499, N120);
and AND3 (N3532, N3530, N501, N1086);
nor NOR2 (N3533, N3532, N109);
nand NAND2 (N3534, N3504, N427);
buf BUF1 (N3535, N3533);
or OR4 (N3536, N3535, N1043, N2446, N3297);
not NOT1 (N3537, N3536);
nor NOR3 (N3538, N3517, N2939, N3506);
and AND2 (N3539, N3522, N3220);
not NOT1 (N3540, N3528);
or OR2 (N3541, N3534, N2294);
nor NOR3 (N3542, N3529, N1689, N1894);
and AND2 (N3543, N3537, N3100);
nand NAND3 (N3544, N3540, N1088, N444);
nor NOR4 (N3545, N3543, N224, N371, N780);
nand NAND4 (N3546, N3523, N1870, N1922, N2027);
nor NOR4 (N3547, N3516, N859, N2287, N647);
not NOT1 (N3548, N3539);
nand NAND4 (N3549, N3538, N3044, N1417, N678);
not NOT1 (N3550, N3527);
nor NOR3 (N3551, N3550, N842, N3233);
not NOT1 (N3552, N3542);
buf BUF1 (N3553, N3551);
nand NAND4 (N3554, N3553, N466, N1443, N3356);
not NOT1 (N3555, N3549);
nor NOR4 (N3556, N3546, N3195, N2082, N1253);
or OR2 (N3557, N3544, N2916);
xor XOR2 (N3558, N3548, N1604);
not NOT1 (N3559, N3545);
xor XOR2 (N3560, N3554, N2658);
or OR4 (N3561, N3555, N1497, N1045, N653);
xor XOR2 (N3562, N3557, N3077);
nor NOR3 (N3563, N3560, N2739, N1358);
nand NAND4 (N3564, N3563, N2742, N113, N795);
nor NOR4 (N3565, N3561, N1812, N3053, N2952);
nor NOR2 (N3566, N3558, N3163);
not NOT1 (N3567, N3556);
xor XOR2 (N3568, N3552, N1101);
buf BUF1 (N3569, N3564);
nand NAND3 (N3570, N3547, N615, N1669);
or OR4 (N3571, N3541, N3142, N2716, N10);
nand NAND4 (N3572, N3568, N2955, N2259, N2812);
xor XOR2 (N3573, N3562, N2080);
buf BUF1 (N3574, N3566);
buf BUF1 (N3575, N3565);
or OR3 (N3576, N3531, N3216, N1228);
buf BUF1 (N3577, N3571);
buf BUF1 (N3578, N3575);
buf BUF1 (N3579, N3573);
or OR2 (N3580, N3567, N2412);
and AND3 (N3581, N3570, N1250, N2010);
nor NOR3 (N3582, N3579, N1039, N3307);
not NOT1 (N3583, N3582);
buf BUF1 (N3584, N3583);
nor NOR2 (N3585, N3578, N2164);
nor NOR4 (N3586, N3572, N624, N2794, N1382);
buf BUF1 (N3587, N3574);
nor NOR2 (N3588, N3580, N2270);
xor XOR2 (N3589, N3585, N1162);
and AND4 (N3590, N3589, N3240, N3209, N313);
buf BUF1 (N3591, N3576);
xor XOR2 (N3592, N3590, N2077);
and AND3 (N3593, N3577, N3169, N1750);
nor NOR2 (N3594, N3584, N249);
nor NOR4 (N3595, N3591, N3497, N6, N574);
buf BUF1 (N3596, N3586);
and AND2 (N3597, N3594, N1473);
nor NOR4 (N3598, N3559, N2362, N691, N888);
and AND4 (N3599, N3593, N1978, N3294, N1059);
xor XOR2 (N3600, N3596, N34);
and AND3 (N3601, N3597, N1970, N2419);
or OR2 (N3602, N3595, N2495);
and AND3 (N3603, N3588, N26, N1647);
nor NOR3 (N3604, N3602, N816, N924);
nor NOR2 (N3605, N3598, N3158);
nor NOR4 (N3606, N3569, N1734, N2509, N483);
nand NAND2 (N3607, N3600, N2838);
nor NOR4 (N3608, N3601, N966, N2656, N3338);
nand NAND3 (N3609, N3606, N1519, N2473);
nand NAND3 (N3610, N3587, N915, N3063);
nand NAND2 (N3611, N3608, N1975);
nand NAND4 (N3612, N3603, N697, N1439, N1902);
or OR4 (N3613, N3607, N650, N312, N2643);
nor NOR2 (N3614, N3592, N2337);
buf BUF1 (N3615, N3611);
xor XOR2 (N3616, N3615, N3425);
nand NAND3 (N3617, N3599, N306, N2580);
nand NAND4 (N3618, N3616, N2041, N493, N3045);
or OR3 (N3619, N3610, N3504, N624);
and AND4 (N3620, N3619, N1124, N2130, N290);
nand NAND2 (N3621, N3605, N977);
and AND2 (N3622, N3612, N709);
nand NAND4 (N3623, N3622, N3294, N1241, N3062);
nand NAND4 (N3624, N3581, N1818, N1840, N292);
nor NOR3 (N3625, N3613, N2994, N2798);
not NOT1 (N3626, N3625);
nand NAND4 (N3627, N3618, N3346, N3210, N3339);
xor XOR2 (N3628, N3614, N1416);
or OR4 (N3629, N3604, N534, N2686, N891);
xor XOR2 (N3630, N3617, N2574);
nor NOR4 (N3631, N3609, N448, N3147, N1055);
nand NAND3 (N3632, N3631, N2127, N1538);
xor XOR2 (N3633, N3624, N2036);
or OR4 (N3634, N3623, N442, N199, N1623);
and AND4 (N3635, N3630, N953, N1974, N941);
nor NOR3 (N3636, N3632, N315, N819);
buf BUF1 (N3637, N3634);
or OR4 (N3638, N3627, N1419, N2036, N599);
not NOT1 (N3639, N3626);
buf BUF1 (N3640, N3633);
or OR2 (N3641, N3637, N1759);
nor NOR3 (N3642, N3638, N3441, N2341);
and AND2 (N3643, N3636, N1122);
not NOT1 (N3644, N3642);
buf BUF1 (N3645, N3640);
buf BUF1 (N3646, N3639);
or OR4 (N3647, N3628, N2834, N2090, N714);
or OR4 (N3648, N3646, N2562, N3033, N2179);
nor NOR3 (N3649, N3621, N3500, N1884);
buf BUF1 (N3650, N3647);
nand NAND3 (N3651, N3649, N1880, N1831);
buf BUF1 (N3652, N3651);
xor XOR2 (N3653, N3648, N2763);
buf BUF1 (N3654, N3629);
or OR2 (N3655, N3641, N3092);
buf BUF1 (N3656, N3645);
not NOT1 (N3657, N3635);
not NOT1 (N3658, N3643);
and AND2 (N3659, N3653, N122);
xor XOR2 (N3660, N3652, N116);
buf BUF1 (N3661, N3620);
xor XOR2 (N3662, N3657, N933);
nand NAND3 (N3663, N3650, N2446, N536);
or OR4 (N3664, N3661, N3091, N552, N2715);
buf BUF1 (N3665, N3660);
nand NAND4 (N3666, N3655, N2338, N186, N2351);
xor XOR2 (N3667, N3665, N3520);
not NOT1 (N3668, N3656);
buf BUF1 (N3669, N3644);
nand NAND2 (N3670, N3667, N2722);
nand NAND3 (N3671, N3668, N2911, N3552);
nand NAND4 (N3672, N3654, N577, N775, N3132);
or OR2 (N3673, N3670, N1209);
and AND3 (N3674, N3658, N645, N1418);
buf BUF1 (N3675, N3669);
nor NOR4 (N3676, N3663, N129, N3020, N3477);
nor NOR4 (N3677, N3675, N2947, N3596, N1041);
or OR4 (N3678, N3677, N2006, N1479, N238);
and AND4 (N3679, N3664, N2740, N3621, N1948);
or OR3 (N3680, N3679, N1499, N2539);
and AND3 (N3681, N3680, N1976, N1569);
or OR3 (N3682, N3659, N3342, N2430);
nor NOR4 (N3683, N3676, N33, N1883, N1275);
or OR4 (N3684, N3672, N1845, N2138, N1696);
xor XOR2 (N3685, N3674, N391);
buf BUF1 (N3686, N3681);
and AND3 (N3687, N3683, N2624, N2138);
nor NOR4 (N3688, N3684, N3514, N1953, N904);
not NOT1 (N3689, N3678);
nor NOR4 (N3690, N3662, N1950, N1344, N476);
buf BUF1 (N3691, N3671);
buf BUF1 (N3692, N3666);
and AND4 (N3693, N3687, N182, N3677, N3677);
and AND3 (N3694, N3673, N1944, N1040);
or OR2 (N3695, N3688, N3056);
or OR2 (N3696, N3690, N2290);
or OR3 (N3697, N3686, N689, N328);
and AND4 (N3698, N3695, N272, N1554, N1110);
nand NAND3 (N3699, N3685, N2887, N833);
nor NOR2 (N3700, N3694, N1472);
or OR3 (N3701, N3696, N1326, N2989);
nor NOR4 (N3702, N3682, N1027, N1884, N1330);
not NOT1 (N3703, N3689);
xor XOR2 (N3704, N3703, N1304);
or OR3 (N3705, N3700, N1937, N1218);
and AND3 (N3706, N3691, N2529, N3022);
or OR2 (N3707, N3701, N2032);
not NOT1 (N3708, N3692);
and AND4 (N3709, N3697, N544, N1555, N422);
nor NOR4 (N3710, N3704, N2129, N347, N3431);
or OR4 (N3711, N3698, N2678, N3073, N1459);
buf BUF1 (N3712, N3711);
nor NOR4 (N3713, N3708, N587, N3173, N697);
nand NAND2 (N3714, N3705, N1260);
xor XOR2 (N3715, N3706, N1072);
buf BUF1 (N3716, N3715);
nand NAND2 (N3717, N3693, N3676);
nor NOR2 (N3718, N3702, N2346);
xor XOR2 (N3719, N3709, N1279);
or OR2 (N3720, N3707, N1582);
or OR2 (N3721, N3716, N1026);
nor NOR4 (N3722, N3721, N1448, N698, N3604);
buf BUF1 (N3723, N3712);
nand NAND3 (N3724, N3723, N213, N3336);
nand NAND4 (N3725, N3719, N2491, N2145, N3059);
nand NAND2 (N3726, N3718, N1890);
buf BUF1 (N3727, N3725);
xor XOR2 (N3728, N3724, N2168);
and AND2 (N3729, N3728, N769);
buf BUF1 (N3730, N3710);
buf BUF1 (N3731, N3699);
or OR4 (N3732, N3717, N2502, N673, N280);
and AND2 (N3733, N3732, N3026);
buf BUF1 (N3734, N3727);
xor XOR2 (N3735, N3720, N1299);
xor XOR2 (N3736, N3733, N974);
not NOT1 (N3737, N3736);
buf BUF1 (N3738, N3735);
and AND3 (N3739, N3729, N2576, N1559);
or OR3 (N3740, N3714, N372, N636);
nor NOR2 (N3741, N3738, N731);
buf BUF1 (N3742, N3713);
nor NOR2 (N3743, N3739, N1199);
nor NOR2 (N3744, N3740, N2288);
xor XOR2 (N3745, N3734, N822);
nand NAND2 (N3746, N3741, N3699);
and AND3 (N3747, N3746, N2400, N488);
buf BUF1 (N3748, N3731);
or OR3 (N3749, N3748, N975, N1059);
and AND2 (N3750, N3749, N1655);
nand NAND2 (N3751, N3743, N2838);
buf BUF1 (N3752, N3750);
or OR3 (N3753, N3737, N1603, N6);
not NOT1 (N3754, N3752);
and AND4 (N3755, N3751, N2257, N837, N294);
nand NAND4 (N3756, N3745, N1954, N3321, N3128);
xor XOR2 (N3757, N3742, N2801);
or OR4 (N3758, N3755, N3197, N3432, N2105);
buf BUF1 (N3759, N3730);
buf BUF1 (N3760, N3722);
nor NOR2 (N3761, N3754, N2208);
buf BUF1 (N3762, N3756);
nand NAND4 (N3763, N3759, N99, N316, N1168);
or OR2 (N3764, N3726, N1635);
or OR3 (N3765, N3744, N2967, N2302);
buf BUF1 (N3766, N3764);
buf BUF1 (N3767, N3763);
nor NOR4 (N3768, N3753, N41, N652, N1233);
not NOT1 (N3769, N3765);
nor NOR2 (N3770, N3766, N808);
or OR2 (N3771, N3761, N1170);
or OR3 (N3772, N3758, N760, N1802);
nor NOR2 (N3773, N3762, N2217);
buf BUF1 (N3774, N3768);
xor XOR2 (N3775, N3770, N3299);
and AND4 (N3776, N3773, N1520, N3244, N2280);
buf BUF1 (N3777, N3771);
not NOT1 (N3778, N3760);
and AND4 (N3779, N3769, N45, N3577, N1770);
xor XOR2 (N3780, N3777, N239);
nand NAND2 (N3781, N3780, N1263);
not NOT1 (N3782, N3767);
xor XOR2 (N3783, N3774, N3217);
nor NOR3 (N3784, N3779, N2816, N2904);
or OR3 (N3785, N3784, N1816, N3518);
nand NAND4 (N3786, N3776, N3568, N2694, N3544);
xor XOR2 (N3787, N3783, N376);
not NOT1 (N3788, N3775);
nor NOR2 (N3789, N3785, N2285);
xor XOR2 (N3790, N3787, N372);
nand NAND3 (N3791, N3782, N2333, N2527);
nand NAND3 (N3792, N3772, N1396, N3064);
nor NOR2 (N3793, N3786, N60);
buf BUF1 (N3794, N3793);
nand NAND4 (N3795, N3778, N750, N285, N429);
nor NOR3 (N3796, N3790, N20, N2349);
or OR4 (N3797, N3796, N883, N1021, N1691);
not NOT1 (N3798, N3794);
or OR2 (N3799, N3757, N1015);
or OR3 (N3800, N3792, N1607, N3760);
and AND4 (N3801, N3800, N3768, N3591, N416);
nand NAND2 (N3802, N3789, N1928);
not NOT1 (N3803, N3797);
buf BUF1 (N3804, N3803);
or OR2 (N3805, N3799, N912);
nand NAND4 (N3806, N3747, N299, N2298, N2990);
and AND3 (N3807, N3801, N559, N1718);
xor XOR2 (N3808, N3791, N3784);
xor XOR2 (N3809, N3807, N1344);
xor XOR2 (N3810, N3809, N3442);
buf BUF1 (N3811, N3808);
and AND2 (N3812, N3806, N793);
or OR4 (N3813, N3811, N1713, N891, N3572);
or OR2 (N3814, N3802, N690);
nor NOR4 (N3815, N3812, N3461, N3035, N2105);
nor NOR3 (N3816, N3805, N3716, N2917);
xor XOR2 (N3817, N3804, N683);
or OR3 (N3818, N3815, N3731, N285);
and AND2 (N3819, N3798, N1296);
not NOT1 (N3820, N3781);
nor NOR4 (N3821, N3820, N370, N3017, N337);
or OR3 (N3822, N3788, N1406, N1288);
xor XOR2 (N3823, N3816, N2186);
or OR3 (N3824, N3823, N2812, N2234);
nor NOR4 (N3825, N3817, N3211, N125, N997);
xor XOR2 (N3826, N3795, N1841);
or OR2 (N3827, N3813, N591);
xor XOR2 (N3828, N3822, N3098);
or OR2 (N3829, N3825, N136);
not NOT1 (N3830, N3824);
xor XOR2 (N3831, N3829, N2976);
nand NAND3 (N3832, N3818, N174, N2687);
and AND4 (N3833, N3819, N2543, N2954, N3777);
and AND4 (N3834, N3827, N92, N616, N2438);
nor NOR4 (N3835, N3821, N3149, N2109, N2892);
xor XOR2 (N3836, N3810, N1595);
not NOT1 (N3837, N3830);
or OR2 (N3838, N3835, N2918);
buf BUF1 (N3839, N3837);
nor NOR3 (N3840, N3833, N1362, N187);
xor XOR2 (N3841, N3828, N172);
nand NAND3 (N3842, N3840, N131, N3037);
and AND3 (N3843, N3814, N2044, N1037);
and AND3 (N3844, N3839, N67, N2618);
nor NOR2 (N3845, N3831, N2957);
and AND3 (N3846, N3845, N53, N679);
nand NAND2 (N3847, N3836, N3714);
nor NOR3 (N3848, N3842, N2523, N1964);
nor NOR4 (N3849, N3841, N3313, N1071, N1153);
xor XOR2 (N3850, N3832, N2042);
nand NAND3 (N3851, N3848, N2134, N2395);
xor XOR2 (N3852, N3847, N2075);
buf BUF1 (N3853, N3851);
nor NOR4 (N3854, N3846, N2235, N1157, N1377);
buf BUF1 (N3855, N3853);
nand NAND3 (N3856, N3849, N3386, N3496);
or OR2 (N3857, N3843, N3463);
xor XOR2 (N3858, N3850, N1346);
buf BUF1 (N3859, N3852);
xor XOR2 (N3860, N3834, N3560);
and AND4 (N3861, N3844, N3614, N3567, N3844);
xor XOR2 (N3862, N3861, N2780);
xor XOR2 (N3863, N3859, N614);
xor XOR2 (N3864, N3862, N398);
or OR2 (N3865, N3855, N520);
and AND4 (N3866, N3826, N3394, N3072, N3127);
buf BUF1 (N3867, N3866);
xor XOR2 (N3868, N3856, N3214);
nand NAND2 (N3869, N3868, N228);
and AND3 (N3870, N3865, N2147, N2952);
and AND4 (N3871, N3867, N3265, N2099, N1204);
or OR3 (N3872, N3854, N3653, N2125);
nor NOR3 (N3873, N3857, N675, N1997);
buf BUF1 (N3874, N3873);
xor XOR2 (N3875, N3860, N1445);
nand NAND2 (N3876, N3863, N2222);
or OR3 (N3877, N3869, N2445, N2985);
buf BUF1 (N3878, N3838);
buf BUF1 (N3879, N3874);
or OR2 (N3880, N3870, N2840);
nor NOR4 (N3881, N3877, N2744, N1810, N281);
nor NOR2 (N3882, N3880, N3614);
nor NOR4 (N3883, N3864, N1751, N140, N3112);
or OR2 (N3884, N3883, N592);
or OR4 (N3885, N3879, N421, N308, N1414);
or OR3 (N3886, N3876, N1494, N2338);
nand NAND2 (N3887, N3871, N3601);
not NOT1 (N3888, N3878);
and AND4 (N3889, N3884, N2289, N1248, N1482);
nand NAND2 (N3890, N3875, N3305);
buf BUF1 (N3891, N3872);
xor XOR2 (N3892, N3887, N3883);
not NOT1 (N3893, N3889);
xor XOR2 (N3894, N3888, N1955);
buf BUF1 (N3895, N3893);
xor XOR2 (N3896, N3890, N810);
nor NOR4 (N3897, N3882, N3294, N982, N839);
buf BUF1 (N3898, N3891);
not NOT1 (N3899, N3885);
not NOT1 (N3900, N3897);
or OR4 (N3901, N3881, N1041, N179, N3872);
buf BUF1 (N3902, N3900);
or OR2 (N3903, N3899, N2416);
and AND3 (N3904, N3898, N1713, N591);
or OR2 (N3905, N3894, N1780);
buf BUF1 (N3906, N3892);
or OR2 (N3907, N3901, N3621);
xor XOR2 (N3908, N3904, N2107);
not NOT1 (N3909, N3908);
nor NOR3 (N3910, N3886, N813, N2304);
nand NAND2 (N3911, N3902, N2346);
not NOT1 (N3912, N3910);
not NOT1 (N3913, N3903);
and AND3 (N3914, N3858, N3242, N3593);
nand NAND2 (N3915, N3905, N1270);
nor NOR3 (N3916, N3913, N3359, N3167);
buf BUF1 (N3917, N3906);
buf BUF1 (N3918, N3914);
not NOT1 (N3919, N3916);
xor XOR2 (N3920, N3909, N2814);
or OR2 (N3921, N3912, N941);
buf BUF1 (N3922, N3907);
and AND2 (N3923, N3895, N3872);
and AND3 (N3924, N3915, N2426, N2606);
and AND4 (N3925, N3922, N2857, N118, N2913);
not NOT1 (N3926, N3918);
buf BUF1 (N3927, N3920);
not NOT1 (N3928, N3927);
nand NAND4 (N3929, N3911, N87, N264, N1370);
buf BUF1 (N3930, N3926);
xor XOR2 (N3931, N3921, N2386);
and AND3 (N3932, N3924, N1291, N1556);
xor XOR2 (N3933, N3932, N95);
not NOT1 (N3934, N3925);
xor XOR2 (N3935, N3896, N1616);
buf BUF1 (N3936, N3930);
buf BUF1 (N3937, N3934);
nor NOR2 (N3938, N3931, N1864);
nor NOR2 (N3939, N3937, N2391);
xor XOR2 (N3940, N3919, N2565);
nor NOR3 (N3941, N3917, N422, N2805);
xor XOR2 (N3942, N3941, N3834);
nand NAND3 (N3943, N3933, N3417, N998);
nand NAND4 (N3944, N3938, N475, N3311, N3462);
nor NOR3 (N3945, N3928, N3584, N1474);
and AND3 (N3946, N3939, N3268, N2174);
or OR3 (N3947, N3942, N3854, N167);
and AND4 (N3948, N3923, N1615, N403, N1393);
and AND3 (N3949, N3935, N2801, N2270);
xor XOR2 (N3950, N3944, N72);
buf BUF1 (N3951, N3947);
nand NAND2 (N3952, N3951, N1709);
and AND4 (N3953, N3943, N3298, N2533, N242);
nor NOR3 (N3954, N3952, N2904, N1392);
buf BUF1 (N3955, N3950);
nor NOR3 (N3956, N3948, N3432, N180);
buf BUF1 (N3957, N3936);
not NOT1 (N3958, N3953);
xor XOR2 (N3959, N3954, N3790);
or OR4 (N3960, N3940, N3119, N1039, N2295);
not NOT1 (N3961, N3929);
not NOT1 (N3962, N3960);
and AND3 (N3963, N3955, N785, N119);
nor NOR4 (N3964, N3946, N3732, N1290, N755);
nor NOR4 (N3965, N3945, N158, N3938, N771);
buf BUF1 (N3966, N3962);
xor XOR2 (N3967, N3961, N556);
and AND4 (N3968, N3964, N1223, N314, N2191);
buf BUF1 (N3969, N3967);
nand NAND2 (N3970, N3957, N3346);
and AND3 (N3971, N3958, N2509, N1430);
xor XOR2 (N3972, N3970, N3528);
nand NAND4 (N3973, N3949, N2375, N3891, N1770);
nand NAND4 (N3974, N3971, N1737, N285, N3275);
or OR4 (N3975, N3963, N161, N2373, N1904);
nand NAND2 (N3976, N3959, N2311);
not NOT1 (N3977, N3956);
nand NAND4 (N3978, N3972, N3624, N2679, N2820);
or OR3 (N3979, N3969, N95, N790);
nand NAND4 (N3980, N3968, N42, N994, N275);
and AND3 (N3981, N3977, N791, N2163);
not NOT1 (N3982, N3974);
nor NOR4 (N3983, N3976, N955, N3921, N350);
buf BUF1 (N3984, N3981);
nand NAND3 (N3985, N3984, N3227, N568);
buf BUF1 (N3986, N3975);
buf BUF1 (N3987, N3985);
or OR4 (N3988, N3978, N1650, N3200, N3573);
nand NAND3 (N3989, N3966, N2856, N1307);
xor XOR2 (N3990, N3979, N3051);
or OR4 (N3991, N3983, N524, N688, N380);
or OR2 (N3992, N3990, N2228);
xor XOR2 (N3993, N3989, N1701);
xor XOR2 (N3994, N3982, N1654);
nor NOR4 (N3995, N3988, N374, N2312, N1645);
buf BUF1 (N3996, N3986);
xor XOR2 (N3997, N3992, N1252);
nor NOR2 (N3998, N3980, N3598);
and AND3 (N3999, N3991, N3988, N1480);
nand NAND2 (N4000, N3998, N1265);
not NOT1 (N4001, N3993);
not NOT1 (N4002, N3965);
buf BUF1 (N4003, N4000);
buf BUF1 (N4004, N3999);
nor NOR2 (N4005, N3973, N3276);
nor NOR3 (N4006, N3996, N253, N3873);
nor NOR4 (N4007, N4001, N1938, N2246, N871);
nand NAND4 (N4008, N4003, N2760, N2284, N4007);
nor NOR4 (N4009, N2809, N2852, N1526, N2493);
nand NAND2 (N4010, N3997, N3960);
not NOT1 (N4011, N4005);
not NOT1 (N4012, N4010);
buf BUF1 (N4013, N4002);
buf BUF1 (N4014, N3994);
or OR2 (N4015, N4006, N3828);
nand NAND3 (N4016, N4013, N2139, N3699);
or OR3 (N4017, N4008, N2788, N2691);
buf BUF1 (N4018, N3987);
or OR3 (N4019, N4012, N1609, N980);
nor NOR3 (N4020, N4004, N2255, N1557);
buf BUF1 (N4021, N4011);
nor NOR4 (N4022, N4014, N633, N1741, N248);
not NOT1 (N4023, N3995);
nand NAND3 (N4024, N4018, N777, N3387);
buf BUF1 (N4025, N4022);
not NOT1 (N4026, N4023);
or OR2 (N4027, N4016, N1621);
xor XOR2 (N4028, N4026, N2402);
and AND4 (N4029, N4009, N198, N3915, N1818);
and AND2 (N4030, N4017, N2807);
nand NAND2 (N4031, N4024, N3676);
nor NOR4 (N4032, N4030, N2037, N2756, N80);
and AND2 (N4033, N4029, N1248);
buf BUF1 (N4034, N4028);
or OR2 (N4035, N4015, N620);
not NOT1 (N4036, N4033);
buf BUF1 (N4037, N4027);
buf BUF1 (N4038, N4021);
not NOT1 (N4039, N4037);
or OR2 (N4040, N4035, N1883);
nand NAND4 (N4041, N4020, N3224, N964, N296);
xor XOR2 (N4042, N4041, N2755);
nor NOR3 (N4043, N4025, N2055, N3251);
buf BUF1 (N4044, N4042);
and AND2 (N4045, N4034, N1373);
xor XOR2 (N4046, N4040, N882);
xor XOR2 (N4047, N4032, N3250);
not NOT1 (N4048, N4046);
or OR2 (N4049, N4039, N661);
xor XOR2 (N4050, N4049, N4015);
nor NOR4 (N4051, N4047, N688, N718, N2436);
or OR2 (N4052, N4031, N1058);
xor XOR2 (N4053, N4019, N208);
buf BUF1 (N4054, N4050);
or OR4 (N4055, N4036, N1820, N1308, N3095);
nand NAND4 (N4056, N4054, N962, N2575, N806);
nand NAND3 (N4057, N4055, N3668, N1124);
nor NOR3 (N4058, N4052, N1763, N1077);
buf BUF1 (N4059, N4043);
nor NOR3 (N4060, N4056, N1369, N2969);
xor XOR2 (N4061, N4058, N3382);
not NOT1 (N4062, N4038);
nor NOR2 (N4063, N4044, N533);
not NOT1 (N4064, N4059);
nand NAND2 (N4065, N4051, N3873);
nand NAND2 (N4066, N4057, N3787);
or OR2 (N4067, N4064, N3673);
buf BUF1 (N4068, N4066);
buf BUF1 (N4069, N4062);
buf BUF1 (N4070, N4068);
or OR2 (N4071, N4067, N561);
and AND4 (N4072, N4063, N3695, N113, N198);
nand NAND3 (N4073, N4065, N3200, N3509);
buf BUF1 (N4074, N4072);
nor NOR4 (N4075, N4060, N3516, N127, N3655);
or OR2 (N4076, N4074, N4008);
xor XOR2 (N4077, N4070, N710);
and AND3 (N4078, N4071, N94, N1101);
nor NOR3 (N4079, N4076, N2444, N1196);
nand NAND4 (N4080, N4073, N2682, N3862, N2423);
not NOT1 (N4081, N4045);
nor NOR3 (N4082, N4078, N594, N130);
nor NOR4 (N4083, N4075, N1731, N2261, N2532);
nand NAND3 (N4084, N4081, N3722, N1877);
nor NOR2 (N4085, N4077, N1809);
or OR3 (N4086, N4080, N3557, N3592);
nand NAND2 (N4087, N4053, N495);
and AND4 (N4088, N4085, N3484, N23, N1229);
and AND2 (N4089, N4087, N2914);
or OR3 (N4090, N4084, N3407, N3061);
and AND3 (N4091, N4048, N2851, N2614);
xor XOR2 (N4092, N4082, N3582);
nor NOR3 (N4093, N4079, N2655, N654);
nand NAND4 (N4094, N4093, N2610, N1588, N3598);
or OR3 (N4095, N4091, N2386, N901);
nand NAND3 (N4096, N4092, N2971, N3712);
nand NAND3 (N4097, N4090, N2943, N3448);
nor NOR4 (N4098, N4097, N2835, N3126, N3801);
xor XOR2 (N4099, N4095, N2900);
nand NAND4 (N4100, N4069, N2522, N1477, N1139);
or OR2 (N4101, N4098, N3345);
not NOT1 (N4102, N4088);
and AND3 (N4103, N4094, N2886, N3234);
nand NAND4 (N4104, N4089, N3533, N3179, N1188);
and AND2 (N4105, N4104, N3403);
and AND4 (N4106, N4099, N417, N1122, N854);
or OR2 (N4107, N4061, N3179);
and AND3 (N4108, N4086, N216, N2120);
or OR3 (N4109, N4102, N696, N2723);
and AND4 (N4110, N4083, N1892, N608, N3277);
not NOT1 (N4111, N4101);
nor NOR3 (N4112, N4111, N3656, N677);
or OR2 (N4113, N4100, N3146);
buf BUF1 (N4114, N4109);
nand NAND2 (N4115, N4106, N3490);
or OR2 (N4116, N4115, N2389);
not NOT1 (N4117, N4114);
nor NOR4 (N4118, N4112, N2161, N400, N3753);
nor NOR3 (N4119, N4110, N3449, N3612);
and AND3 (N4120, N4113, N1115, N889);
buf BUF1 (N4121, N4116);
xor XOR2 (N4122, N4121, N1373);
and AND4 (N4123, N4108, N2251, N2733, N71);
nor NOR4 (N4124, N4118, N1213, N449, N2495);
nand NAND3 (N4125, N4120, N2658, N2056);
nor NOR4 (N4126, N4123, N3166, N3068, N283);
buf BUF1 (N4127, N4107);
nor NOR3 (N4128, N4096, N715, N2022);
nor NOR3 (N4129, N4126, N1501, N3109);
buf BUF1 (N4130, N4119);
buf BUF1 (N4131, N4127);
nor NOR2 (N4132, N4117, N5);
and AND3 (N4133, N4131, N2702, N2165);
xor XOR2 (N4134, N4130, N3490);
nor NOR3 (N4135, N4124, N1266, N850);
buf BUF1 (N4136, N4105);
not NOT1 (N4137, N4132);
nand NAND3 (N4138, N4136, N2583, N3148);
or OR2 (N4139, N4122, N3057);
xor XOR2 (N4140, N4135, N548);
nand NAND3 (N4141, N4133, N588, N136);
xor XOR2 (N4142, N4138, N617);
and AND3 (N4143, N4141, N1989, N3117);
buf BUF1 (N4144, N4128);
nand NAND3 (N4145, N4137, N3835, N1889);
xor XOR2 (N4146, N4103, N2568);
nand NAND3 (N4147, N4143, N3818, N1431);
buf BUF1 (N4148, N4140);
and AND3 (N4149, N4125, N933, N1315);
or OR3 (N4150, N4139, N2700, N1330);
or OR4 (N4151, N4147, N1227, N2040, N2470);
xor XOR2 (N4152, N4149, N3121);
xor XOR2 (N4153, N4129, N2366);
or OR4 (N4154, N4150, N1830, N4137, N3603);
and AND4 (N4155, N4145, N1072, N269, N2625);
or OR2 (N4156, N4142, N3589);
not NOT1 (N4157, N4154);
nor NOR2 (N4158, N4152, N1177);
nor NOR3 (N4159, N4158, N1208, N5);
nand NAND4 (N4160, N4153, N586, N1204, N820);
nor NOR2 (N4161, N4146, N1241);
and AND3 (N4162, N4161, N1388, N2507);
and AND4 (N4163, N4155, N208, N3820, N973);
nand NAND2 (N4164, N4148, N2861);
not NOT1 (N4165, N4163);
or OR4 (N4166, N4144, N1496, N2684, N2213);
xor XOR2 (N4167, N4156, N3905);
buf BUF1 (N4168, N4160);
nor NOR4 (N4169, N4151, N1172, N3057, N683);
nand NAND3 (N4170, N4167, N3118, N2122);
nor NOR2 (N4171, N4165, N890);
buf BUF1 (N4172, N4162);
buf BUF1 (N4173, N4134);
buf BUF1 (N4174, N4170);
nand NAND4 (N4175, N4174, N1583, N2992, N2174);
nor NOR2 (N4176, N4166, N1101);
nor NOR2 (N4177, N4157, N1348);
not NOT1 (N4178, N4171);
buf BUF1 (N4179, N4164);
and AND3 (N4180, N4179, N906, N3345);
nor NOR4 (N4181, N4169, N2913, N2305, N644);
and AND2 (N4182, N4168, N632);
nor NOR3 (N4183, N4176, N1606, N224);
xor XOR2 (N4184, N4172, N3851);
buf BUF1 (N4185, N4173);
nand NAND3 (N4186, N4183, N1011, N911);
or OR4 (N4187, N4175, N3072, N2768, N3825);
nor NOR3 (N4188, N4177, N3109, N2418);
nor NOR2 (N4189, N4187, N649);
xor XOR2 (N4190, N4188, N2470);
nand NAND2 (N4191, N4184, N839);
xor XOR2 (N4192, N4181, N4001);
nand NAND2 (N4193, N4159, N2008);
or OR2 (N4194, N4185, N303);
nor NOR3 (N4195, N4189, N2981, N1105);
or OR3 (N4196, N4191, N2162, N292);
and AND4 (N4197, N4178, N2349, N1958, N85);
xor XOR2 (N4198, N4192, N1199);
nand NAND3 (N4199, N4198, N4167, N200);
xor XOR2 (N4200, N4194, N546);
nor NOR2 (N4201, N4182, N3815);
buf BUF1 (N4202, N4201);
or OR4 (N4203, N4180, N862, N3672, N3712);
buf BUF1 (N4204, N4197);
not NOT1 (N4205, N4196);
nor NOR4 (N4206, N4204, N762, N3143, N297);
not NOT1 (N4207, N4203);
and AND4 (N4208, N4200, N3857, N1438, N1238);
xor XOR2 (N4209, N4207, N3458);
nand NAND2 (N4210, N4199, N3217);
buf BUF1 (N4211, N4209);
or OR3 (N4212, N4195, N3617, N982);
or OR3 (N4213, N4202, N3141, N1841);
not NOT1 (N4214, N4205);
buf BUF1 (N4215, N4212);
nand NAND3 (N4216, N4193, N1744, N2916);
buf BUF1 (N4217, N4211);
buf BUF1 (N4218, N4217);
nand NAND3 (N4219, N4218, N2258, N3625);
xor XOR2 (N4220, N4186, N3801);
nor NOR2 (N4221, N4213, N2580);
nand NAND2 (N4222, N4221, N321);
and AND3 (N4223, N4208, N363, N521);
nand NAND4 (N4224, N4206, N2075, N3250, N126);
buf BUF1 (N4225, N4190);
xor XOR2 (N4226, N4219, N1238);
buf BUF1 (N4227, N4222);
or OR2 (N4228, N4224, N3130);
nor NOR4 (N4229, N4220, N2286, N1108, N3793);
xor XOR2 (N4230, N4223, N974);
xor XOR2 (N4231, N4215, N3519);
buf BUF1 (N4232, N4225);
or OR4 (N4233, N4229, N2147, N721, N3222);
buf BUF1 (N4234, N4230);
and AND3 (N4235, N4214, N4045, N3084);
xor XOR2 (N4236, N4231, N851);
nand NAND4 (N4237, N4227, N4105, N2199, N1837);
xor XOR2 (N4238, N4216, N3886);
or OR4 (N4239, N4235, N3283, N3788, N3231);
nor NOR2 (N4240, N4233, N1475);
nand NAND4 (N4241, N4238, N2773, N3858, N1180);
nor NOR3 (N4242, N4226, N2311, N3725);
and AND4 (N4243, N4228, N1341, N1256, N855);
xor XOR2 (N4244, N4210, N1704);
nor NOR4 (N4245, N4239, N2351, N705, N579);
not NOT1 (N4246, N4242);
buf BUF1 (N4247, N4234);
nor NOR4 (N4248, N4245, N2217, N2517, N3213);
or OR3 (N4249, N4244, N1965, N3176);
buf BUF1 (N4250, N4246);
nor NOR4 (N4251, N4250, N1266, N1594, N1725);
not NOT1 (N4252, N4232);
not NOT1 (N4253, N4249);
not NOT1 (N4254, N4236);
nor NOR4 (N4255, N4251, N1403, N941, N2291);
nor NOR2 (N4256, N4254, N3553);
nand NAND3 (N4257, N4247, N3439, N2725);
xor XOR2 (N4258, N4256, N1703);
nand NAND4 (N4259, N4253, N996, N1045, N2462);
nor NOR4 (N4260, N4243, N2010, N1873, N238);
and AND4 (N4261, N4252, N2128, N1410, N3899);
not NOT1 (N4262, N4241);
or OR3 (N4263, N4262, N4126, N2705);
or OR3 (N4264, N4263, N2504, N823);
xor XOR2 (N4265, N4261, N1014);
nand NAND4 (N4266, N4248, N831, N2876, N788);
nand NAND4 (N4267, N4258, N1176, N2076, N3958);
or OR4 (N4268, N4259, N3204, N459, N470);
xor XOR2 (N4269, N4266, N2698);
nor NOR4 (N4270, N4240, N1664, N1145, N3849);
or OR2 (N4271, N4257, N2507);
not NOT1 (N4272, N4237);
nor NOR2 (N4273, N4265, N1409);
not NOT1 (N4274, N4273);
nand NAND2 (N4275, N4267, N865);
buf BUF1 (N4276, N4269);
or OR3 (N4277, N4255, N1397, N526);
nor NOR3 (N4278, N4276, N4164, N402);
or OR2 (N4279, N4264, N2620);
nor NOR3 (N4280, N4268, N2403, N970);
and AND4 (N4281, N4260, N4269, N2106, N895);
and AND3 (N4282, N4277, N2223, N1775);
not NOT1 (N4283, N4274);
and AND4 (N4284, N4275, N828, N1212, N1284);
or OR2 (N4285, N4281, N1720);
xor XOR2 (N4286, N4271, N3144);
xor XOR2 (N4287, N4279, N3137);
xor XOR2 (N4288, N4282, N1381);
nand NAND4 (N4289, N4286, N4020, N1411, N3754);
or OR3 (N4290, N4289, N3037, N1014);
nand NAND4 (N4291, N4283, N2619, N246, N738);
not NOT1 (N4292, N4288);
nor NOR3 (N4293, N4284, N3893, N3022);
nand NAND2 (N4294, N4270, N4185);
and AND4 (N4295, N4287, N3139, N67, N397);
nor NOR4 (N4296, N4294, N4073, N1764, N3688);
not NOT1 (N4297, N4293);
nand NAND4 (N4298, N4291, N3493, N418, N3718);
not NOT1 (N4299, N4296);
and AND4 (N4300, N4295, N3297, N2222, N3659);
xor XOR2 (N4301, N4298, N1342);
nor NOR3 (N4302, N4300, N165, N63);
nand NAND2 (N4303, N4297, N2171);
not NOT1 (N4304, N4280);
buf BUF1 (N4305, N4303);
buf BUF1 (N4306, N4302);
and AND4 (N4307, N4306, N3251, N1711, N3258);
and AND3 (N4308, N4307, N1312, N692);
and AND3 (N4309, N4304, N3167, N1125);
buf BUF1 (N4310, N4290);
and AND4 (N4311, N4305, N2197, N1780, N2504);
xor XOR2 (N4312, N4285, N1305);
or OR4 (N4313, N4308, N1666, N4212, N1674);
or OR4 (N4314, N4299, N578, N3630, N3111);
nor NOR3 (N4315, N4278, N3837, N3232);
xor XOR2 (N4316, N4315, N4077);
xor XOR2 (N4317, N4313, N342);
or OR2 (N4318, N4311, N480);
nand NAND4 (N4319, N4316, N2603, N4, N639);
buf BUF1 (N4320, N4318);
nand NAND4 (N4321, N4310, N3117, N3332, N2921);
not NOT1 (N4322, N4292);
xor XOR2 (N4323, N4319, N829);
buf BUF1 (N4324, N4317);
nor NOR3 (N4325, N4272, N1960, N813);
and AND2 (N4326, N4320, N2149);
not NOT1 (N4327, N4321);
or OR2 (N4328, N4327, N485);
nand NAND4 (N4329, N4301, N3882, N1542, N2678);
or OR2 (N4330, N4324, N1021);
nor NOR3 (N4331, N4314, N324, N202);
xor XOR2 (N4332, N4322, N836);
not NOT1 (N4333, N4309);
nor NOR4 (N4334, N4312, N2318, N2596, N2495);
nand NAND3 (N4335, N4325, N1582, N1918);
and AND2 (N4336, N4330, N1705);
buf BUF1 (N4337, N4333);
xor XOR2 (N4338, N4331, N582);
nor NOR2 (N4339, N4336, N3164);
nor NOR3 (N4340, N4332, N718, N2597);
or OR2 (N4341, N4335, N370);
buf BUF1 (N4342, N4339);
xor XOR2 (N4343, N4328, N3126);
or OR4 (N4344, N4323, N2708, N2745, N3995);
nor NOR2 (N4345, N4329, N56);
not NOT1 (N4346, N4344);
and AND2 (N4347, N4342, N307);
nor NOR2 (N4348, N4347, N3085);
nand NAND3 (N4349, N4346, N2943, N91);
nor NOR3 (N4350, N4345, N4330, N2485);
and AND2 (N4351, N4348, N1439);
nand NAND2 (N4352, N4338, N590);
nor NOR4 (N4353, N4343, N1410, N4056, N273);
not NOT1 (N4354, N4340);
not NOT1 (N4355, N4350);
nand NAND3 (N4356, N4337, N3737, N1212);
nand NAND3 (N4357, N4351, N1123, N2631);
xor XOR2 (N4358, N4355, N3662);
or OR2 (N4359, N4358, N1316);
and AND3 (N4360, N4326, N605, N2388);
nand NAND4 (N4361, N4360, N3981, N4121, N2199);
xor XOR2 (N4362, N4361, N2678);
xor XOR2 (N4363, N4334, N3060);
not NOT1 (N4364, N4352);
or OR4 (N4365, N4354, N3946, N84, N1652);
nor NOR3 (N4366, N4341, N234, N2299);
and AND2 (N4367, N4357, N2604);
nor NOR4 (N4368, N4353, N2768, N745, N2479);
xor XOR2 (N4369, N4364, N2112);
nor NOR2 (N4370, N4367, N137);
not NOT1 (N4371, N4369);
nand NAND4 (N4372, N4349, N2063, N972, N3606);
buf BUF1 (N4373, N4372);
not NOT1 (N4374, N4365);
or OR3 (N4375, N4374, N1684, N3467);
not NOT1 (N4376, N4363);
xor XOR2 (N4377, N4362, N3811);
or OR4 (N4378, N4368, N800, N3148, N2299);
xor XOR2 (N4379, N4366, N1399);
and AND4 (N4380, N4376, N1592, N3211, N1345);
xor XOR2 (N4381, N4379, N3433);
nor NOR2 (N4382, N4377, N1773);
nand NAND2 (N4383, N4382, N2523);
xor XOR2 (N4384, N4373, N3922);
xor XOR2 (N4385, N4381, N1342);
and AND2 (N4386, N4371, N3275);
and AND3 (N4387, N4385, N3593, N2138);
or OR2 (N4388, N4356, N441);
xor XOR2 (N4389, N4370, N1550);
not NOT1 (N4390, N4389);
and AND4 (N4391, N4380, N2308, N1159, N3997);
or OR2 (N4392, N4387, N3227);
not NOT1 (N4393, N4392);
buf BUF1 (N4394, N4375);
or OR4 (N4395, N4386, N3094, N2686, N2978);
buf BUF1 (N4396, N4395);
or OR3 (N4397, N4359, N3228, N3903);
or OR4 (N4398, N4388, N1890, N974, N2153);
nor NOR2 (N4399, N4383, N2904);
nand NAND2 (N4400, N4398, N2554);
xor XOR2 (N4401, N4400, N1749);
nand NAND3 (N4402, N4391, N2258, N2851);
and AND3 (N4403, N4399, N2039, N839);
and AND3 (N4404, N4378, N3464, N354);
or OR4 (N4405, N4403, N2829, N798, N16);
not NOT1 (N4406, N4404);
or OR2 (N4407, N4402, N1415);
not NOT1 (N4408, N4397);
not NOT1 (N4409, N4406);
nor NOR4 (N4410, N4384, N2256, N3623, N3227);
nor NOR4 (N4411, N4396, N769, N2735, N2540);
xor XOR2 (N4412, N4411, N600);
nor NOR2 (N4413, N4393, N3916);
not NOT1 (N4414, N4401);
buf BUF1 (N4415, N4407);
nand NAND3 (N4416, N4409, N225, N529);
not NOT1 (N4417, N4416);
or OR2 (N4418, N4394, N3642);
and AND3 (N4419, N4418, N2221, N3768);
not NOT1 (N4420, N4408);
not NOT1 (N4421, N4405);
buf BUF1 (N4422, N4415);
nor NOR4 (N4423, N4421, N2223, N3329, N3723);
buf BUF1 (N4424, N4423);
buf BUF1 (N4425, N4390);
xor XOR2 (N4426, N4424, N807);
not NOT1 (N4427, N4425);
not NOT1 (N4428, N4414);
or OR2 (N4429, N4410, N173);
buf BUF1 (N4430, N4428);
buf BUF1 (N4431, N4417);
nand NAND3 (N4432, N4429, N419, N122);
nor NOR3 (N4433, N4413, N2397, N3951);
nand NAND4 (N4434, N4431, N3827, N1949, N741);
nor NOR2 (N4435, N4419, N3842);
buf BUF1 (N4436, N4434);
and AND3 (N4437, N4435, N2723, N955);
or OR2 (N4438, N4412, N2980);
or OR2 (N4439, N4436, N3421);
nor NOR4 (N4440, N4430, N903, N3921, N1173);
nand NAND4 (N4441, N4427, N2532, N1386, N3323);
or OR4 (N4442, N4420, N2687, N739, N1198);
and AND4 (N4443, N4442, N3411, N648, N2194);
nor NOR4 (N4444, N4438, N2570, N1425, N419);
and AND4 (N4445, N4432, N3879, N1418, N4161);
nor NOR4 (N4446, N4433, N226, N2074, N1487);
not NOT1 (N4447, N4446);
or OR3 (N4448, N4426, N1783, N1549);
xor XOR2 (N4449, N4437, N4277);
and AND2 (N4450, N4444, N2734);
nor NOR3 (N4451, N4422, N4096, N1714);
nand NAND2 (N4452, N4443, N566);
nor NOR4 (N4453, N4449, N2014, N1462, N4404);
nand NAND3 (N4454, N4445, N3130, N901);
nor NOR2 (N4455, N4450, N1481);
xor XOR2 (N4456, N4453, N1571);
or OR4 (N4457, N4448, N2127, N4404, N2748);
nand NAND2 (N4458, N4451, N2270);
nand NAND2 (N4459, N4458, N1511);
nand NAND2 (N4460, N4459, N3419);
and AND2 (N4461, N4441, N3512);
xor XOR2 (N4462, N4454, N1662);
or OR4 (N4463, N4456, N2681, N1230, N1039);
buf BUF1 (N4464, N4439);
xor XOR2 (N4465, N4462, N2024);
not NOT1 (N4466, N4461);
or OR2 (N4467, N4464, N1025);
or OR3 (N4468, N4467, N1230, N2627);
buf BUF1 (N4469, N4440);
nor NOR2 (N4470, N4469, N3190);
xor XOR2 (N4471, N4447, N816);
xor XOR2 (N4472, N4471, N2439);
nor NOR3 (N4473, N4452, N1460, N4071);
nand NAND3 (N4474, N4457, N3572, N182);
nand NAND2 (N4475, N4472, N951);
or OR4 (N4476, N4466, N1735, N3987, N184);
nor NOR3 (N4477, N4473, N3869, N2210);
buf BUF1 (N4478, N4475);
nand NAND2 (N4479, N4476, N3874);
buf BUF1 (N4480, N4477);
or OR3 (N4481, N4478, N2238, N2400);
and AND2 (N4482, N4470, N4056);
and AND3 (N4483, N4455, N4388, N2072);
nor NOR2 (N4484, N4480, N977);
nand NAND4 (N4485, N4479, N4330, N4156, N220);
not NOT1 (N4486, N4482);
nand NAND3 (N4487, N4486, N1103, N2507);
buf BUF1 (N4488, N4481);
or OR2 (N4489, N4487, N1053);
nand NAND3 (N4490, N4483, N3519, N1574);
nand NAND3 (N4491, N4488, N4138, N1705);
nand NAND4 (N4492, N4465, N3370, N98, N1233);
and AND4 (N4493, N4485, N782, N3020, N4191);
nor NOR3 (N4494, N4474, N3461, N2999);
or OR2 (N4495, N4490, N463);
nor NOR2 (N4496, N4489, N369);
nand NAND3 (N4497, N4468, N1001, N1715);
buf BUF1 (N4498, N4493);
xor XOR2 (N4499, N4460, N2763);
not NOT1 (N4500, N4495);
or OR4 (N4501, N4463, N2310, N1633, N1303);
or OR4 (N4502, N4500, N3884, N1962, N3178);
not NOT1 (N4503, N4496);
and AND2 (N4504, N4502, N2802);
buf BUF1 (N4505, N4501);
or OR3 (N4506, N4503, N3723, N1878);
and AND4 (N4507, N4504, N4068, N2933, N618);
and AND4 (N4508, N4505, N3540, N2147, N1725);
and AND4 (N4509, N4484, N3988, N1454, N2779);
nor NOR2 (N4510, N4498, N4260);
and AND2 (N4511, N4508, N4140);
buf BUF1 (N4512, N4497);
or OR4 (N4513, N4511, N2315, N2517, N537);
buf BUF1 (N4514, N4507);
and AND2 (N4515, N4499, N4471);
xor XOR2 (N4516, N4491, N4512);
not NOT1 (N4517, N4294);
buf BUF1 (N4518, N4492);
nor NOR2 (N4519, N4506, N1644);
buf BUF1 (N4520, N4515);
or OR2 (N4521, N4520, N3190);
nor NOR2 (N4522, N4521, N4155);
not NOT1 (N4523, N4517);
nor NOR2 (N4524, N4510, N2250);
nand NAND2 (N4525, N4514, N860);
nor NOR3 (N4526, N4522, N385, N1319);
xor XOR2 (N4527, N4518, N533);
and AND4 (N4528, N4509, N824, N4096, N1919);
nor NOR4 (N4529, N4527, N4423, N1746, N149);
buf BUF1 (N4530, N4525);
nand NAND4 (N4531, N4526, N1375, N136, N3928);
nor NOR4 (N4532, N4519, N405, N1261, N550);
or OR2 (N4533, N4524, N3086);
nor NOR2 (N4534, N4494, N1738);
nand NAND4 (N4535, N4528, N1434, N416, N359);
or OR4 (N4536, N4532, N3084, N2029, N4151);
xor XOR2 (N4537, N4534, N4307);
nor NOR4 (N4538, N4516, N3086, N2002, N1583);
nand NAND4 (N4539, N4523, N3504, N1465, N4049);
xor XOR2 (N4540, N4539, N92);
nand NAND4 (N4541, N4540, N3157, N3304, N292);
nand NAND4 (N4542, N4529, N169, N1004, N33);
xor XOR2 (N4543, N4537, N2279);
nand NAND3 (N4544, N4542, N4396, N2931);
xor XOR2 (N4545, N4513, N1435);
or OR4 (N4546, N4538, N248, N2807, N3839);
nor NOR3 (N4547, N4545, N2103, N2586);
xor XOR2 (N4548, N4547, N2188);
buf BUF1 (N4549, N4541);
nand NAND3 (N4550, N4531, N2849, N2342);
and AND4 (N4551, N4536, N2673, N2083, N3174);
nand NAND4 (N4552, N4535, N1411, N1595, N37);
or OR2 (N4553, N4530, N3705);
not NOT1 (N4554, N4548);
not NOT1 (N4555, N4550);
or OR3 (N4556, N4551, N21, N3482);
xor XOR2 (N4557, N4552, N2248);
buf BUF1 (N4558, N4557);
nand NAND3 (N4559, N4533, N4244, N979);
not NOT1 (N4560, N4555);
or OR4 (N4561, N4553, N156, N742, N3834);
nand NAND2 (N4562, N4556, N1167);
nand NAND4 (N4563, N4558, N579, N502, N3445);
or OR3 (N4564, N4562, N3597, N604);
or OR2 (N4565, N4564, N4047);
nor NOR4 (N4566, N4543, N4164, N2524, N3177);
and AND2 (N4567, N4566, N700);
or OR4 (N4568, N4563, N18, N2084, N3704);
nand NAND3 (N4569, N4546, N736, N3513);
not NOT1 (N4570, N4559);
buf BUF1 (N4571, N4560);
not NOT1 (N4572, N4569);
or OR2 (N4573, N4561, N4567);
xor XOR2 (N4574, N226, N1436);
xor XOR2 (N4575, N4565, N3147);
nand NAND2 (N4576, N4554, N669);
or OR4 (N4577, N4573, N1907, N2687, N523);
xor XOR2 (N4578, N4568, N3175);
xor XOR2 (N4579, N4577, N4362);
and AND4 (N4580, N4575, N2195, N3392, N1624);
or OR3 (N4581, N4580, N1849, N3634);
or OR4 (N4582, N4579, N3914, N452, N1535);
xor XOR2 (N4583, N4544, N4335);
nand NAND3 (N4584, N4549, N1295, N1236);
or OR2 (N4585, N4578, N1931);
xor XOR2 (N4586, N4585, N2849);
or OR4 (N4587, N4582, N2631, N4240, N3902);
buf BUF1 (N4588, N4570);
or OR3 (N4589, N4571, N2755, N1719);
and AND4 (N4590, N4581, N1590, N4441, N4330);
buf BUF1 (N4591, N4587);
nor NOR4 (N4592, N4589, N1675, N524, N2022);
xor XOR2 (N4593, N4590, N3467);
not NOT1 (N4594, N4591);
buf BUF1 (N4595, N4586);
or OR4 (N4596, N4584, N1911, N1090, N1256);
nor NOR4 (N4597, N4588, N547, N233, N689);
nand NAND3 (N4598, N4572, N2989, N3255);
not NOT1 (N4599, N4574);
xor XOR2 (N4600, N4593, N4041);
and AND2 (N4601, N4598, N1103);
buf BUF1 (N4602, N4576);
buf BUF1 (N4603, N4601);
and AND4 (N4604, N4600, N2500, N1309, N3578);
not NOT1 (N4605, N4592);
nor NOR4 (N4606, N4594, N2607, N1933, N1166);
and AND3 (N4607, N4605, N4462, N2332);
not NOT1 (N4608, N4596);
buf BUF1 (N4609, N4597);
buf BUF1 (N4610, N4603);
or OR4 (N4611, N4606, N2610, N2456, N99);
not NOT1 (N4612, N4583);
or OR3 (N4613, N4595, N2113, N3019);
and AND3 (N4614, N4610, N2660, N4221);
buf BUF1 (N4615, N4604);
nand NAND3 (N4616, N4602, N204, N1334);
nand NAND2 (N4617, N4612, N2425);
or OR4 (N4618, N4607, N4129, N1123, N2064);
or OR4 (N4619, N4617, N4375, N2935, N3319);
and AND3 (N4620, N4609, N1966, N2319);
nor NOR2 (N4621, N4615, N451);
nand NAND4 (N4622, N4618, N2213, N1684, N1841);
and AND3 (N4623, N4620, N1572, N3018);
or OR3 (N4624, N4599, N2441, N3496);
and AND4 (N4625, N4621, N2754, N2034, N325);
nand NAND3 (N4626, N4624, N1318, N3589);
nand NAND2 (N4627, N4623, N3726);
or OR4 (N4628, N4625, N3677, N4601, N4476);
not NOT1 (N4629, N4628);
and AND2 (N4630, N4611, N3445);
buf BUF1 (N4631, N4616);
xor XOR2 (N4632, N4630, N2173);
or OR2 (N4633, N4613, N1237);
nand NAND4 (N4634, N4619, N2688, N4337, N2165);
buf BUF1 (N4635, N4633);
nor NOR3 (N4636, N4608, N2889, N394);
not NOT1 (N4637, N4622);
not NOT1 (N4638, N4626);
buf BUF1 (N4639, N4627);
not NOT1 (N4640, N4632);
not NOT1 (N4641, N4640);
nand NAND4 (N4642, N4614, N357, N3676, N1108);
xor XOR2 (N4643, N4631, N3617);
buf BUF1 (N4644, N4635);
xor XOR2 (N4645, N4634, N3398);
nor NOR4 (N4646, N4642, N3536, N4621, N3402);
buf BUF1 (N4647, N4629);
buf BUF1 (N4648, N4636);
nand NAND3 (N4649, N4641, N3288, N4187);
buf BUF1 (N4650, N4639);
or OR4 (N4651, N4649, N1846, N636, N4269);
or OR2 (N4652, N4651, N2349);
not NOT1 (N4653, N4650);
xor XOR2 (N4654, N4646, N2934);
nor NOR2 (N4655, N4647, N1541);
not NOT1 (N4656, N4655);
not NOT1 (N4657, N4638);
nand NAND3 (N4658, N4644, N3158, N2366);
and AND3 (N4659, N4643, N2843, N1376);
not NOT1 (N4660, N4656);
xor XOR2 (N4661, N4652, N4556);
xor XOR2 (N4662, N4658, N2868);
xor XOR2 (N4663, N4645, N3716);
not NOT1 (N4664, N4663);
nand NAND3 (N4665, N4654, N1830, N3455);
nor NOR3 (N4666, N4664, N3973, N2893);
nand NAND4 (N4667, N4665, N1525, N1058, N2808);
not NOT1 (N4668, N4667);
xor XOR2 (N4669, N4648, N2274);
and AND2 (N4670, N4653, N1002);
buf BUF1 (N4671, N4666);
nand NAND4 (N4672, N4660, N578, N4145, N4367);
nor NOR3 (N4673, N4668, N1787, N3520);
xor XOR2 (N4674, N4661, N2096);
not NOT1 (N4675, N4659);
nand NAND3 (N4676, N4673, N3411, N3239);
nor NOR4 (N4677, N4637, N1320, N813, N3274);
nand NAND2 (N4678, N4657, N3535);
buf BUF1 (N4679, N4674);
nand NAND4 (N4680, N4675, N4443, N2717, N762);
not NOT1 (N4681, N4672);
nor NOR2 (N4682, N4681, N1821);
nand NAND2 (N4683, N4662, N3066);
not NOT1 (N4684, N4679);
nor NOR3 (N4685, N4684, N97, N3438);
not NOT1 (N4686, N4683);
nor NOR3 (N4687, N4677, N2933, N1093);
xor XOR2 (N4688, N4687, N332);
buf BUF1 (N4689, N4688);
or OR4 (N4690, N4678, N2246, N3937, N1003);
and AND2 (N4691, N4690, N4148);
buf BUF1 (N4692, N4680);
nand NAND2 (N4693, N4689, N3885);
or OR3 (N4694, N4671, N1782, N967);
nand NAND4 (N4695, N4676, N1334, N2397, N56);
buf BUF1 (N4696, N4692);
not NOT1 (N4697, N4669);
buf BUF1 (N4698, N4696);
nand NAND3 (N4699, N4670, N2898, N2068);
or OR4 (N4700, N4691, N2173, N3859, N228);
buf BUF1 (N4701, N4698);
not NOT1 (N4702, N4700);
buf BUF1 (N4703, N4693);
nand NAND2 (N4704, N4695, N2657);
and AND3 (N4705, N4699, N592, N584);
and AND2 (N4706, N4705, N1099);
nor NOR4 (N4707, N4703, N1719, N70, N1002);
nor NOR3 (N4708, N4701, N2970, N1542);
xor XOR2 (N4709, N4707, N1865);
and AND4 (N4710, N4685, N72, N1360, N4521);
and AND4 (N4711, N4708, N3717, N3051, N2142);
nand NAND4 (N4712, N4710, N3468, N1098, N2783);
not NOT1 (N4713, N4704);
not NOT1 (N4714, N4712);
and AND4 (N4715, N4694, N830, N1891, N1773);
nor NOR3 (N4716, N4711, N1360, N2096);
nor NOR2 (N4717, N4706, N2876);
buf BUF1 (N4718, N4717);
nand NAND3 (N4719, N4718, N4710, N3061);
xor XOR2 (N4720, N4709, N1056);
not NOT1 (N4721, N4715);
xor XOR2 (N4722, N4713, N3491);
nor NOR3 (N4723, N4721, N4634, N441);
nand NAND4 (N4724, N4682, N1653, N4416, N1677);
not NOT1 (N4725, N4723);
and AND4 (N4726, N4719, N3058, N3708, N1285);
nand NAND3 (N4727, N4714, N3501, N30);
and AND3 (N4728, N4720, N1492, N2797);
xor XOR2 (N4729, N4724, N873);
buf BUF1 (N4730, N4697);
nand NAND3 (N4731, N4722, N357, N3486);
not NOT1 (N4732, N4729);
and AND3 (N4733, N4716, N4655, N84);
nand NAND2 (N4734, N4686, N202);
nor NOR2 (N4735, N4725, N4536);
or OR2 (N4736, N4728, N4108);
not NOT1 (N4737, N4730);
nand NAND3 (N4738, N4726, N484, N2917);
nand NAND3 (N4739, N4737, N1380, N789);
nand NAND2 (N4740, N4727, N1554);
nor NOR4 (N4741, N4738, N1770, N4697, N3561);
nand NAND4 (N4742, N4736, N4159, N1036, N2958);
or OR3 (N4743, N4732, N1237, N2842);
buf BUF1 (N4744, N4731);
xor XOR2 (N4745, N4733, N4121);
and AND3 (N4746, N4740, N114, N2741);
nor NOR2 (N4747, N4702, N3912);
or OR4 (N4748, N4747, N3537, N4737, N3974);
and AND4 (N4749, N4742, N1098, N2868, N1313);
buf BUF1 (N4750, N4734);
xor XOR2 (N4751, N4743, N1396);
xor XOR2 (N4752, N4749, N1887);
xor XOR2 (N4753, N4746, N3662);
or OR3 (N4754, N4748, N2864, N772);
buf BUF1 (N4755, N4754);
nor NOR4 (N4756, N4753, N1123, N934, N2527);
nand NAND2 (N4757, N4739, N1633);
and AND2 (N4758, N4755, N1591);
or OR2 (N4759, N4750, N3570);
nor NOR2 (N4760, N4759, N3520);
nand NAND3 (N4761, N4756, N2415, N487);
and AND3 (N4762, N4735, N462, N429);
buf BUF1 (N4763, N4741);
nor NOR4 (N4764, N4752, N1172, N2319, N40);
nor NOR3 (N4765, N4744, N789, N328);
xor XOR2 (N4766, N4762, N2340);
nor NOR2 (N4767, N4763, N2088);
xor XOR2 (N4768, N4758, N1527);
nand NAND2 (N4769, N4765, N4558);
and AND4 (N4770, N4767, N2684, N2298, N292);
nor NOR2 (N4771, N4764, N533);
buf BUF1 (N4772, N4761);
or OR3 (N4773, N4766, N1565, N2782);
buf BUF1 (N4774, N4757);
buf BUF1 (N4775, N4771);
not NOT1 (N4776, N4774);
nand NAND4 (N4777, N4773, N3664, N1183, N3531);
xor XOR2 (N4778, N4769, N3074);
xor XOR2 (N4779, N4778, N662);
nor NOR3 (N4780, N4776, N1610, N899);
and AND4 (N4781, N4760, N3960, N356, N2840);
nor NOR3 (N4782, N4745, N4117, N3090);
buf BUF1 (N4783, N4782);
or OR3 (N4784, N4772, N1032, N3632);
not NOT1 (N4785, N4781);
nor NOR2 (N4786, N4768, N3395);
nor NOR4 (N4787, N4770, N3738, N1420, N2447);
and AND3 (N4788, N4787, N3387, N3328);
not NOT1 (N4789, N4775);
not NOT1 (N4790, N4751);
and AND3 (N4791, N4779, N878, N1791);
not NOT1 (N4792, N4790);
or OR3 (N4793, N4791, N1584, N3467);
buf BUF1 (N4794, N4783);
nand NAND3 (N4795, N4777, N4607, N1159);
not NOT1 (N4796, N4794);
xor XOR2 (N4797, N4785, N3560);
buf BUF1 (N4798, N4793);
not NOT1 (N4799, N4788);
not NOT1 (N4800, N4798);
nor NOR2 (N4801, N4797, N3259);
or OR3 (N4802, N4792, N2087, N2206);
buf BUF1 (N4803, N4795);
xor XOR2 (N4804, N4799, N2998);
or OR2 (N4805, N4796, N1572);
or OR2 (N4806, N4805, N3876);
nor NOR3 (N4807, N4802, N374, N2034);
and AND4 (N4808, N4786, N364, N2870, N3479);
buf BUF1 (N4809, N4807);
and AND3 (N4810, N4808, N3905, N4674);
nand NAND4 (N4811, N4806, N3976, N1107, N1215);
xor XOR2 (N4812, N4800, N2452);
buf BUF1 (N4813, N4784);
or OR2 (N4814, N4789, N3449);
nand NAND4 (N4815, N4780, N611, N3793, N2572);
not NOT1 (N4816, N4815);
nor NOR3 (N4817, N4811, N1810, N4649);
xor XOR2 (N4818, N4809, N4616);
and AND3 (N4819, N4803, N4129, N1718);
xor XOR2 (N4820, N4818, N4779);
nand NAND3 (N4821, N4819, N964, N1123);
and AND4 (N4822, N4813, N2302, N1964, N3441);
nand NAND3 (N4823, N4817, N3757, N4428);
and AND3 (N4824, N4816, N2191, N4522);
buf BUF1 (N4825, N4801);
buf BUF1 (N4826, N4824);
buf BUF1 (N4827, N4826);
and AND2 (N4828, N4814, N1034);
nor NOR4 (N4829, N4825, N1695, N231, N3610);
xor XOR2 (N4830, N4810, N3521);
nor NOR3 (N4831, N4830, N4664, N2686);
buf BUF1 (N4832, N4827);
and AND3 (N4833, N4820, N3154, N638);
not NOT1 (N4834, N4804);
not NOT1 (N4835, N4832);
xor XOR2 (N4836, N4812, N3189);
buf BUF1 (N4837, N4834);
nor NOR3 (N4838, N4829, N568, N4778);
nand NAND2 (N4839, N4828, N531);
nor NOR2 (N4840, N4835, N3414);
buf BUF1 (N4841, N4837);
nand NAND4 (N4842, N4833, N2020, N2362, N1728);
xor XOR2 (N4843, N4823, N4379);
nor NOR4 (N4844, N4841, N3009, N3621, N4140);
and AND3 (N4845, N4843, N918, N651);
and AND4 (N4846, N4831, N4362, N4684, N2874);
and AND4 (N4847, N4844, N3588, N2133, N2705);
not NOT1 (N4848, N4839);
buf BUF1 (N4849, N4842);
and AND4 (N4850, N4821, N157, N2277, N1261);
nor NOR4 (N4851, N4850, N191, N2363, N503);
nor NOR4 (N4852, N4847, N618, N1504, N2678);
not NOT1 (N4853, N4851);
nand NAND4 (N4854, N4822, N2835, N3011, N2457);
nand NAND2 (N4855, N4846, N2769);
xor XOR2 (N4856, N4849, N3116);
not NOT1 (N4857, N4845);
nor NOR3 (N4858, N4852, N1758, N104);
nand NAND3 (N4859, N4855, N3274, N4369);
not NOT1 (N4860, N4848);
xor XOR2 (N4861, N4856, N1963);
not NOT1 (N4862, N4854);
not NOT1 (N4863, N4860);
or OR2 (N4864, N4836, N1122);
and AND2 (N4865, N4853, N274);
and AND2 (N4866, N4859, N181);
xor XOR2 (N4867, N4838, N1234);
buf BUF1 (N4868, N4858);
or OR4 (N4869, N4868, N819, N4118, N3029);
or OR4 (N4870, N4864, N570, N3669, N4565);
nor NOR2 (N4871, N4840, N698);
xor XOR2 (N4872, N4867, N1272);
and AND4 (N4873, N4865, N22, N1651, N587);
xor XOR2 (N4874, N4862, N136);
nor NOR3 (N4875, N4872, N2758, N4613);
or OR2 (N4876, N4861, N2768);
and AND3 (N4877, N4875, N4524, N2982);
buf BUF1 (N4878, N4869);
not NOT1 (N4879, N4878);
or OR3 (N4880, N4879, N564, N2649);
nand NAND2 (N4881, N4876, N2230);
and AND4 (N4882, N4857, N4512, N2661, N1069);
xor XOR2 (N4883, N4882, N2538);
not NOT1 (N4884, N4870);
nor NOR2 (N4885, N4880, N2017);
nor NOR3 (N4886, N4866, N1346, N4406);
xor XOR2 (N4887, N4873, N1149);
nor NOR3 (N4888, N4883, N140, N4712);
xor XOR2 (N4889, N4884, N499);
nand NAND2 (N4890, N4877, N4025);
or OR4 (N4891, N4881, N286, N4756, N3491);
buf BUF1 (N4892, N4891);
and AND3 (N4893, N4885, N4546, N1082);
not NOT1 (N4894, N4889);
and AND2 (N4895, N4863, N3385);
nand NAND3 (N4896, N4887, N1108, N3544);
not NOT1 (N4897, N4886);
xor XOR2 (N4898, N4874, N1759);
nand NAND2 (N4899, N4888, N2280);
or OR2 (N4900, N4892, N3794);
or OR4 (N4901, N4898, N3257, N4606, N3028);
and AND3 (N4902, N4896, N4496, N4033);
xor XOR2 (N4903, N4902, N2809);
buf BUF1 (N4904, N4903);
and AND3 (N4905, N4897, N2691, N1611);
xor XOR2 (N4906, N4901, N4212);
buf BUF1 (N4907, N4895);
xor XOR2 (N4908, N4871, N352);
xor XOR2 (N4909, N4899, N3437);
xor XOR2 (N4910, N4894, N1837);
not NOT1 (N4911, N4907);
and AND4 (N4912, N4910, N3766, N1122, N3824);
nand NAND4 (N4913, N4906, N4681, N1662, N301);
and AND2 (N4914, N4893, N194);
or OR4 (N4915, N4912, N1365, N3842, N555);
or OR4 (N4916, N4908, N4014, N1011, N2021);
not NOT1 (N4917, N4909);
buf BUF1 (N4918, N4915);
buf BUF1 (N4919, N4911);
or OR3 (N4920, N4918, N3635, N3357);
not NOT1 (N4921, N4919);
or OR3 (N4922, N4916, N905, N4031);
or OR3 (N4923, N4914, N263, N2813);
nand NAND2 (N4924, N4904, N602);
or OR4 (N4925, N4917, N4553, N4690, N1801);
buf BUF1 (N4926, N4913);
nand NAND2 (N4927, N4905, N904);
not NOT1 (N4928, N4900);
or OR3 (N4929, N4890, N1887, N879);
or OR2 (N4930, N4924, N795);
xor XOR2 (N4931, N4921, N976);
and AND2 (N4932, N4925, N3810);
nor NOR2 (N4933, N4929, N46);
not NOT1 (N4934, N4922);
xor XOR2 (N4935, N4920, N3434);
nor NOR3 (N4936, N4935, N4671, N814);
or OR3 (N4937, N4926, N1789, N185);
not NOT1 (N4938, N4937);
and AND4 (N4939, N4928, N2281, N2755, N4291);
nand NAND3 (N4940, N4936, N764, N2206);
nor NOR3 (N4941, N4940, N4917, N1899);
nor NOR3 (N4942, N4923, N3021, N881);
nand NAND4 (N4943, N4939, N2209, N1952, N4395);
and AND4 (N4944, N4933, N2173, N2543, N3805);
nand NAND4 (N4945, N4931, N461, N4539, N1119);
and AND3 (N4946, N4943, N4940, N2216);
nor NOR3 (N4947, N4942, N4658, N4228);
or OR4 (N4948, N4938, N2266, N864, N2373);
or OR2 (N4949, N4930, N1437);
or OR2 (N4950, N4947, N4574);
not NOT1 (N4951, N4944);
and AND3 (N4952, N4934, N4228, N4604);
buf BUF1 (N4953, N4941);
nor NOR3 (N4954, N4932, N2630, N3412);
xor XOR2 (N4955, N4951, N3948);
nor NOR4 (N4956, N4946, N4695, N1073, N1546);
buf BUF1 (N4957, N4953);
xor XOR2 (N4958, N4927, N1645);
nor NOR3 (N4959, N4955, N3683, N1078);
nor NOR4 (N4960, N4945, N631, N306, N110);
nand NAND3 (N4961, N4958, N2735, N317);
or OR3 (N4962, N4960, N260, N3821);
buf BUF1 (N4963, N4957);
or OR2 (N4964, N4956, N3595);
and AND3 (N4965, N4949, N3408, N1955);
not NOT1 (N4966, N4950);
or OR3 (N4967, N4959, N3177, N2836);
not NOT1 (N4968, N4964);
nand NAND3 (N4969, N4962, N1650, N1051);
buf BUF1 (N4970, N4967);
nand NAND3 (N4971, N4961, N1903, N972);
or OR3 (N4972, N4954, N3564, N3001);
not NOT1 (N4973, N4969);
xor XOR2 (N4974, N4971, N244);
buf BUF1 (N4975, N4973);
and AND2 (N4976, N4970, N4267);
xor XOR2 (N4977, N4952, N1066);
or OR2 (N4978, N4972, N2131);
not NOT1 (N4979, N4968);
nand NAND2 (N4980, N4974, N1516);
xor XOR2 (N4981, N4948, N691);
and AND3 (N4982, N4981, N2670, N2492);
or OR2 (N4983, N4966, N2120);
not NOT1 (N4984, N4975);
buf BUF1 (N4985, N4978);
and AND2 (N4986, N4982, N3187);
nand NAND3 (N4987, N4983, N1939, N3106);
not NOT1 (N4988, N4985);
buf BUF1 (N4989, N4979);
and AND4 (N4990, N4988, N2644, N3255, N4275);
and AND4 (N4991, N4980, N3669, N476, N3071);
or OR4 (N4992, N4965, N4544, N1399, N1846);
nand NAND2 (N4993, N4992, N4976);
not NOT1 (N4994, N2767);
nor NOR4 (N4995, N4987, N4777, N3553, N3164);
and AND4 (N4996, N4963, N3920, N1187, N2336);
or OR4 (N4997, N4977, N354, N3612, N4902);
nand NAND2 (N4998, N4996, N2140);
buf BUF1 (N4999, N4993);
buf BUF1 (N5000, N4999);
xor XOR2 (N5001, N4998, N2807);
buf BUF1 (N5002, N4984);
not NOT1 (N5003, N4986);
or OR2 (N5004, N4990, N2790);
nand NAND3 (N5005, N4989, N3651, N2075);
and AND4 (N5006, N5005, N1100, N4139, N49);
and AND2 (N5007, N5002, N4366);
buf BUF1 (N5008, N5007);
nor NOR3 (N5009, N4991, N3194, N4569);
nand NAND2 (N5010, N4994, N3343);
not NOT1 (N5011, N5000);
xor XOR2 (N5012, N5003, N742);
not NOT1 (N5013, N5012);
xor XOR2 (N5014, N5004, N2778);
and AND3 (N5015, N5001, N3465, N3739);
not NOT1 (N5016, N5013);
xor XOR2 (N5017, N4997, N4102);
buf BUF1 (N5018, N5015);
nand NAND2 (N5019, N5011, N2444);
xor XOR2 (N5020, N5010, N682);
not NOT1 (N5021, N5020);
nand NAND2 (N5022, N5018, N2498);
and AND4 (N5023, N5016, N4986, N4013, N4704);
xor XOR2 (N5024, N5022, N2439);
xor XOR2 (N5025, N5023, N367);
not NOT1 (N5026, N5014);
nand NAND4 (N5027, N5021, N3400, N709, N4517);
buf BUF1 (N5028, N5024);
and AND4 (N5029, N5028, N3157, N2048, N2258);
nand NAND2 (N5030, N5017, N4020);
nand NAND3 (N5031, N5009, N2288, N4012);
nand NAND4 (N5032, N5027, N2752, N2624, N4684);
xor XOR2 (N5033, N5029, N4486);
buf BUF1 (N5034, N5019);
not NOT1 (N5035, N4995);
nor NOR3 (N5036, N5006, N4658, N4437);
nand NAND4 (N5037, N5032, N3080, N3160, N2899);
buf BUF1 (N5038, N5035);
xor XOR2 (N5039, N5025, N1076);
buf BUF1 (N5040, N5034);
nand NAND3 (N5041, N5036, N1679, N3063);
or OR4 (N5042, N5037, N2815, N4421, N238);
or OR2 (N5043, N5042, N3372);
not NOT1 (N5044, N5030);
and AND3 (N5045, N5040, N2558, N2903);
or OR4 (N5046, N5045, N2682, N3989, N2995);
nand NAND4 (N5047, N5039, N4680, N4873, N3959);
nor NOR3 (N5048, N5026, N47, N4679);
nor NOR4 (N5049, N5008, N3640, N1276, N3748);
buf BUF1 (N5050, N5031);
nor NOR2 (N5051, N5049, N3574);
nand NAND3 (N5052, N5046, N2519, N2353);
xor XOR2 (N5053, N5043, N4236);
nand NAND3 (N5054, N5033, N164, N700);
nor NOR3 (N5055, N5044, N4517, N3007);
not NOT1 (N5056, N5038);
or OR4 (N5057, N5056, N4453, N331, N3829);
nor NOR2 (N5058, N5052, N1994);
buf BUF1 (N5059, N5051);
and AND2 (N5060, N5055, N4482);
or OR2 (N5061, N5047, N1487);
nand NAND2 (N5062, N5048, N4474);
nand NAND4 (N5063, N5050, N4897, N3273, N384);
xor XOR2 (N5064, N5058, N1626);
buf BUF1 (N5065, N5041);
not NOT1 (N5066, N5063);
buf BUF1 (N5067, N5059);
xor XOR2 (N5068, N5062, N4740);
not NOT1 (N5069, N5064);
buf BUF1 (N5070, N5067);
not NOT1 (N5071, N5066);
xor XOR2 (N5072, N5071, N2318);
xor XOR2 (N5073, N5053, N1392);
buf BUF1 (N5074, N5057);
not NOT1 (N5075, N5068);
not NOT1 (N5076, N5069);
xor XOR2 (N5077, N5061, N2696);
or OR3 (N5078, N5060, N1063, N4116);
nor NOR2 (N5079, N5065, N1674);
nor NOR2 (N5080, N5072, N4399);
and AND3 (N5081, N5076, N2574, N3910);
and AND3 (N5082, N5078, N3848, N1317);
and AND2 (N5083, N5079, N3033);
nand NAND3 (N5084, N5082, N3321, N1308);
xor XOR2 (N5085, N5054, N4611);
nor NOR2 (N5086, N5084, N2187);
xor XOR2 (N5087, N5080, N2252);
buf BUF1 (N5088, N5070);
nand NAND4 (N5089, N5087, N2811, N1003, N3706);
buf BUF1 (N5090, N5073);
xor XOR2 (N5091, N5075, N4298);
xor XOR2 (N5092, N5074, N2914);
nor NOR2 (N5093, N5091, N4405);
or OR3 (N5094, N5085, N1583, N2366);
and AND3 (N5095, N5089, N1609, N175);
xor XOR2 (N5096, N5083, N669);
and AND2 (N5097, N5093, N335);
nor NOR4 (N5098, N5090, N2968, N2642, N3782);
or OR2 (N5099, N5096, N3173);
and AND2 (N5100, N5098, N1018);
nor NOR4 (N5101, N5099, N2424, N922, N3733);
buf BUF1 (N5102, N5100);
or OR3 (N5103, N5077, N3182, N925);
or OR4 (N5104, N5102, N650, N5034, N1902);
not NOT1 (N5105, N5092);
buf BUF1 (N5106, N5097);
and AND4 (N5107, N5088, N4945, N4773, N3790);
not NOT1 (N5108, N5103);
xor XOR2 (N5109, N5108, N4649);
or OR3 (N5110, N5086, N2909, N4184);
or OR3 (N5111, N5095, N5110, N3800);
nand NAND4 (N5112, N1161, N2747, N681, N4476);
nand NAND4 (N5113, N5109, N864, N4361, N3898);
nor NOR3 (N5114, N5111, N1827, N180);
not NOT1 (N5115, N5105);
buf BUF1 (N5116, N5115);
buf BUF1 (N5117, N5104);
nor NOR3 (N5118, N5107, N1417, N264);
and AND2 (N5119, N5112, N211);
nand NAND2 (N5120, N5116, N1659);
nor NOR4 (N5121, N5094, N1975, N3603, N3325);
and AND4 (N5122, N5120, N1691, N3485, N2129);
buf BUF1 (N5123, N5106);
or OR3 (N5124, N5118, N377, N3888);
xor XOR2 (N5125, N5117, N1255);
buf BUF1 (N5126, N5124);
not NOT1 (N5127, N5123);
xor XOR2 (N5128, N5122, N3286);
xor XOR2 (N5129, N5127, N3842);
buf BUF1 (N5130, N5114);
buf BUF1 (N5131, N5121);
xor XOR2 (N5132, N5129, N4608);
xor XOR2 (N5133, N5126, N1849);
or OR4 (N5134, N5101, N225, N3018, N154);
xor XOR2 (N5135, N5113, N1660);
not NOT1 (N5136, N5131);
buf BUF1 (N5137, N5132);
not NOT1 (N5138, N5081);
not NOT1 (N5139, N5130);
nor NOR4 (N5140, N5125, N4333, N100, N2066);
nor NOR2 (N5141, N5134, N4839);
not NOT1 (N5142, N5135);
xor XOR2 (N5143, N5138, N2031);
nand NAND4 (N5144, N5119, N1772, N4672, N3212);
nand NAND2 (N5145, N5141, N3437);
xor XOR2 (N5146, N5128, N3416);
or OR2 (N5147, N5139, N482);
nand NAND4 (N5148, N5145, N4445, N968, N602);
nand NAND4 (N5149, N5143, N687, N2884, N2123);
nand NAND4 (N5150, N5133, N2436, N1075, N3227);
or OR4 (N5151, N5146, N1643, N4198, N1169);
buf BUF1 (N5152, N5136);
and AND3 (N5153, N5137, N2449, N2221);
nor NOR2 (N5154, N5148, N4096);
or OR3 (N5155, N5151, N520, N2728);
xor XOR2 (N5156, N5150, N2058);
xor XOR2 (N5157, N5147, N895);
nand NAND2 (N5158, N5153, N3958);
or OR2 (N5159, N5140, N3474);
nor NOR4 (N5160, N5144, N267, N1271, N2294);
not NOT1 (N5161, N5158);
xor XOR2 (N5162, N5159, N4980);
not NOT1 (N5163, N5157);
buf BUF1 (N5164, N5154);
nand NAND3 (N5165, N5164, N455, N4100);
nor NOR3 (N5166, N5160, N4205, N519);
buf BUF1 (N5167, N5155);
nand NAND3 (N5168, N5161, N927, N3360);
not NOT1 (N5169, N5167);
xor XOR2 (N5170, N5165, N1406);
not NOT1 (N5171, N5166);
nand NAND2 (N5172, N5170, N2573);
xor XOR2 (N5173, N5171, N4127);
nor NOR2 (N5174, N5142, N441);
nand NAND4 (N5175, N5173, N320, N888, N3356);
and AND4 (N5176, N5172, N3480, N451, N4022);
and AND3 (N5177, N5163, N4781, N3932);
xor XOR2 (N5178, N5149, N4600);
and AND4 (N5179, N5178, N99, N5149, N212);
nor NOR3 (N5180, N5179, N434, N1307);
nor NOR3 (N5181, N5177, N311, N518);
nand NAND2 (N5182, N5156, N1876);
xor XOR2 (N5183, N5180, N1663);
xor XOR2 (N5184, N5169, N2686);
buf BUF1 (N5185, N5176);
nand NAND4 (N5186, N5175, N712, N4434, N3970);
buf BUF1 (N5187, N5168);
not NOT1 (N5188, N5181);
nor NOR3 (N5189, N5188, N2197, N2847);
nand NAND3 (N5190, N5185, N1504, N3672);
nand NAND4 (N5191, N5182, N3799, N4510, N4627);
nor NOR3 (N5192, N5187, N835, N3383);
nand NAND2 (N5193, N5174, N2297);
and AND3 (N5194, N5190, N2624, N672);
nand NAND2 (N5195, N5184, N1172);
or OR3 (N5196, N5193, N2369, N4321);
nor NOR3 (N5197, N5194, N2304, N4107);
and AND4 (N5198, N5191, N2664, N4873, N5016);
buf BUF1 (N5199, N5197);
nand NAND3 (N5200, N5162, N5185, N4514);
nand NAND2 (N5201, N5198, N1881);
nor NOR2 (N5202, N5195, N3104);
or OR3 (N5203, N5183, N4431, N630);
nor NOR3 (N5204, N5202, N4096, N3057);
and AND2 (N5205, N5203, N859);
or OR4 (N5206, N5189, N1409, N372, N5020);
not NOT1 (N5207, N5205);
xor XOR2 (N5208, N5201, N155);
not NOT1 (N5209, N5196);
nor NOR3 (N5210, N5208, N4739, N1867);
nand NAND4 (N5211, N5199, N4961, N1607, N1915);
and AND4 (N5212, N5192, N3434, N4361, N5199);
and AND2 (N5213, N5152, N1587);
nand NAND3 (N5214, N5204, N3230, N2692);
nor NOR2 (N5215, N5200, N5125);
not NOT1 (N5216, N5213);
nor NOR2 (N5217, N5216, N4642);
xor XOR2 (N5218, N5207, N975);
nor NOR3 (N5219, N5218, N234, N5022);
xor XOR2 (N5220, N5219, N3548);
buf BUF1 (N5221, N5211);
or OR4 (N5222, N5220, N4550, N3767, N2592);
buf BUF1 (N5223, N5214);
nand NAND4 (N5224, N5222, N391, N2636, N2581);
nand NAND4 (N5225, N5221, N1638, N4659, N3903);
nor NOR2 (N5226, N5225, N2395);
or OR2 (N5227, N5212, N2301);
buf BUF1 (N5228, N5223);
not NOT1 (N5229, N5186);
nor NOR2 (N5230, N5217, N896);
or OR2 (N5231, N5229, N4238);
not NOT1 (N5232, N5215);
buf BUF1 (N5233, N5209);
not NOT1 (N5234, N5227);
nand NAND3 (N5235, N5233, N1116, N409);
nor NOR4 (N5236, N5226, N4911, N3871, N232);
and AND2 (N5237, N5234, N1101);
not NOT1 (N5238, N5231);
and AND4 (N5239, N5224, N5113, N4783, N2477);
buf BUF1 (N5240, N5230);
nor NOR4 (N5241, N5232, N937, N3661, N2167);
xor XOR2 (N5242, N5210, N1856);
nand NAND3 (N5243, N5242, N1901, N694);
and AND3 (N5244, N5237, N2196, N3778);
not NOT1 (N5245, N5243);
buf BUF1 (N5246, N5228);
nor NOR2 (N5247, N5206, N4061);
nand NAND3 (N5248, N5245, N3966, N4380);
buf BUF1 (N5249, N5241);
not NOT1 (N5250, N5238);
nor NOR2 (N5251, N5248, N4612);
or OR4 (N5252, N5247, N2419, N622, N4198);
nor NOR2 (N5253, N5251, N1255);
xor XOR2 (N5254, N5253, N421);
and AND3 (N5255, N5239, N2229, N3478);
nand NAND2 (N5256, N5236, N3078);
xor XOR2 (N5257, N5256, N1914);
nand NAND4 (N5258, N5257, N4336, N2846, N2982);
xor XOR2 (N5259, N5255, N3170);
not NOT1 (N5260, N5254);
not NOT1 (N5261, N5258);
or OR3 (N5262, N5240, N4030, N2831);
xor XOR2 (N5263, N5261, N5247);
not NOT1 (N5264, N5235);
xor XOR2 (N5265, N5262, N118);
nor NOR4 (N5266, N5246, N5152, N997, N3840);
nor NOR2 (N5267, N5244, N1078);
buf BUF1 (N5268, N5250);
not NOT1 (N5269, N5265);
and AND3 (N5270, N5263, N247, N333);
buf BUF1 (N5271, N5252);
nand NAND4 (N5272, N5260, N3599, N4633, N1190);
not NOT1 (N5273, N5268);
buf BUF1 (N5274, N5272);
nand NAND3 (N5275, N5273, N1451, N4916);
not NOT1 (N5276, N5275);
not NOT1 (N5277, N5267);
not NOT1 (N5278, N5274);
buf BUF1 (N5279, N5277);
xor XOR2 (N5280, N5278, N1627);
buf BUF1 (N5281, N5266);
nor NOR2 (N5282, N5281, N565);
xor XOR2 (N5283, N5276, N4548);
nor NOR2 (N5284, N5249, N3249);
buf BUF1 (N5285, N5284);
buf BUF1 (N5286, N5280);
xor XOR2 (N5287, N5259, N3745);
buf BUF1 (N5288, N5287);
nor NOR4 (N5289, N5264, N608, N3281, N1976);
nor NOR3 (N5290, N5285, N5192, N699);
not NOT1 (N5291, N5282);
buf BUF1 (N5292, N5279);
xor XOR2 (N5293, N5270, N1589);
buf BUF1 (N5294, N5291);
buf BUF1 (N5295, N5286);
xor XOR2 (N5296, N5292, N1976);
xor XOR2 (N5297, N5288, N3992);
xor XOR2 (N5298, N5294, N2523);
nand NAND2 (N5299, N5295, N2327);
xor XOR2 (N5300, N5296, N3981);
not NOT1 (N5301, N5290);
and AND4 (N5302, N5283, N4430, N3032, N2390);
or OR2 (N5303, N5301, N4973);
and AND3 (N5304, N5298, N3710, N1126);
or OR4 (N5305, N5297, N3135, N5134, N639);
xor XOR2 (N5306, N5289, N3408);
not NOT1 (N5307, N5302);
xor XOR2 (N5308, N5269, N1292);
nand NAND3 (N5309, N5304, N2769, N371);
buf BUF1 (N5310, N5307);
nor NOR3 (N5311, N5308, N2820, N4629);
not NOT1 (N5312, N5300);
or OR2 (N5313, N5306, N4847);
nor NOR3 (N5314, N5303, N4390, N4813);
xor XOR2 (N5315, N5314, N1603);
nand NAND3 (N5316, N5312, N3630, N404);
and AND4 (N5317, N5299, N108, N351, N4514);
buf BUF1 (N5318, N5313);
not NOT1 (N5319, N5305);
not NOT1 (N5320, N5310);
not NOT1 (N5321, N5318);
nand NAND4 (N5322, N5293, N4729, N4760, N3463);
nor NOR4 (N5323, N5317, N826, N1592, N5191);
not NOT1 (N5324, N5319);
nor NOR2 (N5325, N5320, N1744);
and AND2 (N5326, N5311, N1776);
nor NOR3 (N5327, N5271, N2718, N1695);
nor NOR2 (N5328, N5315, N903);
nand NAND3 (N5329, N5326, N4291, N3440);
nand NAND4 (N5330, N5323, N2328, N2876, N1177);
not NOT1 (N5331, N5322);
not NOT1 (N5332, N5309);
buf BUF1 (N5333, N5321);
or OR3 (N5334, N5316, N2552, N799);
and AND4 (N5335, N5331, N4144, N1876, N3644);
and AND4 (N5336, N5328, N2890, N1944, N4029);
or OR3 (N5337, N5332, N3655, N738);
and AND2 (N5338, N5335, N2502);
and AND3 (N5339, N5336, N835, N1814);
not NOT1 (N5340, N5329);
or OR4 (N5341, N5334, N2867, N166, N1406);
and AND2 (N5342, N5327, N4771);
or OR2 (N5343, N5330, N1900);
nor NOR2 (N5344, N5340, N1595);
or OR2 (N5345, N5339, N3054);
not NOT1 (N5346, N5337);
nand NAND4 (N5347, N5324, N1761, N3886, N3461);
not NOT1 (N5348, N5346);
nand NAND3 (N5349, N5345, N5296, N5317);
and AND3 (N5350, N5325, N2015, N3061);
or OR2 (N5351, N5343, N2965);
not NOT1 (N5352, N5341);
and AND3 (N5353, N5344, N895, N4005);
not NOT1 (N5354, N5350);
buf BUF1 (N5355, N5333);
or OR2 (N5356, N5338, N788);
not NOT1 (N5357, N5352);
and AND2 (N5358, N5354, N5155);
or OR3 (N5359, N5358, N5182, N3219);
nand NAND3 (N5360, N5342, N2243, N4952);
or OR4 (N5361, N5357, N958, N2270, N801);
and AND3 (N5362, N5348, N918, N3566);
xor XOR2 (N5363, N5356, N2916);
not NOT1 (N5364, N5359);
nor NOR2 (N5365, N5355, N4286);
and AND4 (N5366, N5347, N4308, N781, N1545);
nand NAND3 (N5367, N5351, N953, N2030);
nand NAND3 (N5368, N5366, N1144, N849);
buf BUF1 (N5369, N5353);
or OR4 (N5370, N5349, N2985, N4267, N772);
xor XOR2 (N5371, N5360, N4568);
not NOT1 (N5372, N5364);
or OR4 (N5373, N5368, N966, N2769, N3360);
nand NAND2 (N5374, N5370, N4872);
not NOT1 (N5375, N5372);
nor NOR3 (N5376, N5373, N4064, N1039);
nor NOR2 (N5377, N5376, N760);
xor XOR2 (N5378, N5363, N1810);
or OR3 (N5379, N5371, N3153, N3752);
xor XOR2 (N5380, N5369, N5133);
xor XOR2 (N5381, N5365, N4554);
not NOT1 (N5382, N5378);
and AND2 (N5383, N5361, N2511);
nor NOR2 (N5384, N5383, N4657);
and AND2 (N5385, N5362, N3069);
xor XOR2 (N5386, N5379, N1552);
nor NOR3 (N5387, N5385, N1189, N3588);
xor XOR2 (N5388, N5386, N474);
buf BUF1 (N5389, N5377);
xor XOR2 (N5390, N5389, N3744);
xor XOR2 (N5391, N5374, N1308);
and AND3 (N5392, N5391, N5252, N1645);
buf BUF1 (N5393, N5392);
nand NAND4 (N5394, N5384, N4508, N859, N819);
or OR4 (N5395, N5390, N3923, N4506, N2502);
and AND2 (N5396, N5380, N932);
xor XOR2 (N5397, N5394, N3799);
nand NAND3 (N5398, N5397, N1114, N1867);
xor XOR2 (N5399, N5375, N2803);
xor XOR2 (N5400, N5382, N1869);
buf BUF1 (N5401, N5399);
nor NOR3 (N5402, N5367, N1952, N2465);
and AND2 (N5403, N5402, N3419);
buf BUF1 (N5404, N5400);
buf BUF1 (N5405, N5393);
and AND3 (N5406, N5387, N75, N1733);
not NOT1 (N5407, N5401);
nor NOR4 (N5408, N5398, N4324, N1235, N3002);
and AND3 (N5409, N5407, N3911, N1208);
and AND3 (N5410, N5405, N1577, N1526);
nor NOR2 (N5411, N5388, N1297);
and AND2 (N5412, N5381, N1369);
xor XOR2 (N5413, N5395, N685);
not NOT1 (N5414, N5408);
xor XOR2 (N5415, N5411, N1267);
or OR2 (N5416, N5412, N1721);
not NOT1 (N5417, N5415);
xor XOR2 (N5418, N5410, N3836);
xor XOR2 (N5419, N5396, N232);
not NOT1 (N5420, N5413);
and AND4 (N5421, N5416, N1692, N4066, N2318);
not NOT1 (N5422, N5417);
nand NAND2 (N5423, N5420, N1102);
or OR2 (N5424, N5406, N2220);
or OR4 (N5425, N5421, N4937, N257, N1411);
not NOT1 (N5426, N5404);
or OR2 (N5427, N5423, N2395);
and AND4 (N5428, N5427, N1384, N190, N1283);
not NOT1 (N5429, N5414);
and AND2 (N5430, N5409, N5302);
nand NAND2 (N5431, N5419, N2237);
not NOT1 (N5432, N5424);
not NOT1 (N5433, N5403);
xor XOR2 (N5434, N5418, N648);
buf BUF1 (N5435, N5434);
and AND3 (N5436, N5428, N3064, N266);
and AND2 (N5437, N5422, N1855);
not NOT1 (N5438, N5432);
nand NAND2 (N5439, N5437, N1701);
or OR2 (N5440, N5438, N2647);
buf BUF1 (N5441, N5440);
and AND2 (N5442, N5425, N3163);
and AND3 (N5443, N5430, N1304, N1413);
and AND3 (N5444, N5426, N3643, N3915);
nor NOR2 (N5445, N5429, N2030);
and AND2 (N5446, N5431, N2932);
xor XOR2 (N5447, N5443, N1552);
nand NAND4 (N5448, N5441, N4264, N4187, N961);
not NOT1 (N5449, N5433);
nand NAND2 (N5450, N5447, N1255);
buf BUF1 (N5451, N5435);
not NOT1 (N5452, N5444);
not NOT1 (N5453, N5445);
and AND4 (N5454, N5439, N3847, N1902, N2275);
not NOT1 (N5455, N5452);
xor XOR2 (N5456, N5450, N5144);
buf BUF1 (N5457, N5446);
not NOT1 (N5458, N5457);
not NOT1 (N5459, N5451);
nor NOR4 (N5460, N5453, N483, N4935, N4761);
not NOT1 (N5461, N5455);
or OR3 (N5462, N5456, N600, N4847);
nand NAND2 (N5463, N5449, N854);
xor XOR2 (N5464, N5448, N3457);
xor XOR2 (N5465, N5460, N4280);
nand NAND2 (N5466, N5459, N262);
nand NAND4 (N5467, N5463, N2567, N536, N3230);
buf BUF1 (N5468, N5466);
and AND2 (N5469, N5436, N1863);
xor XOR2 (N5470, N5462, N850);
nor NOR2 (N5471, N5470, N1822);
xor XOR2 (N5472, N5465, N657);
or OR3 (N5473, N5461, N2390, N1296);
nor NOR3 (N5474, N5454, N3929, N4667);
xor XOR2 (N5475, N5472, N180);
and AND4 (N5476, N5467, N3788, N1451, N2209);
xor XOR2 (N5477, N5468, N5122);
nand NAND2 (N5478, N5473, N2685);
not NOT1 (N5479, N5458);
or OR3 (N5480, N5471, N2413, N2932);
and AND4 (N5481, N5476, N2867, N4027, N351);
nor NOR3 (N5482, N5474, N4678, N4962);
not NOT1 (N5483, N5477);
not NOT1 (N5484, N5475);
buf BUF1 (N5485, N5478);
not NOT1 (N5486, N5483);
and AND4 (N5487, N5442, N5278, N902, N739);
or OR2 (N5488, N5469, N635);
and AND4 (N5489, N5485, N4699, N1389, N5416);
nor NOR4 (N5490, N5481, N3486, N5193, N4160);
buf BUF1 (N5491, N5489);
buf BUF1 (N5492, N5487);
xor XOR2 (N5493, N5486, N5255);
and AND4 (N5494, N5484, N695, N296, N1650);
nor NOR3 (N5495, N5491, N1966, N3881);
xor XOR2 (N5496, N5495, N688);
xor XOR2 (N5497, N5479, N4585);
and AND4 (N5498, N5492, N1108, N2782, N4180);
buf BUF1 (N5499, N5464);
or OR3 (N5500, N5482, N4333, N4966);
buf BUF1 (N5501, N5490);
or OR4 (N5502, N5499, N1480, N939, N1148);
not NOT1 (N5503, N5488);
nor NOR4 (N5504, N5503, N1917, N1975, N3586);
and AND4 (N5505, N5502, N1907, N4829, N4953);
buf BUF1 (N5506, N5498);
buf BUF1 (N5507, N5500);
nor NOR2 (N5508, N5506, N1364);
xor XOR2 (N5509, N5480, N2298);
xor XOR2 (N5510, N5508, N3204);
not NOT1 (N5511, N5510);
xor XOR2 (N5512, N5496, N1593);
and AND4 (N5513, N5512, N4640, N1032, N1942);
nand NAND4 (N5514, N5507, N2363, N3967, N1894);
not NOT1 (N5515, N5501);
and AND3 (N5516, N5509, N1818, N3208);
nand NAND4 (N5517, N5504, N1178, N4634, N3160);
not NOT1 (N5518, N5513);
buf BUF1 (N5519, N5505);
nor NOR4 (N5520, N5494, N1946, N5310, N3681);
nor NOR3 (N5521, N5497, N222, N3785);
buf BUF1 (N5522, N5511);
not NOT1 (N5523, N5516);
not NOT1 (N5524, N5520);
xor XOR2 (N5525, N5517, N4758);
and AND2 (N5526, N5522, N2059);
nor NOR4 (N5527, N5519, N723, N3818, N3648);
buf BUF1 (N5528, N5526);
xor XOR2 (N5529, N5518, N4338);
xor XOR2 (N5530, N5527, N1584);
buf BUF1 (N5531, N5530);
or OR2 (N5532, N5514, N2202);
nand NAND4 (N5533, N5521, N5300, N5050, N434);
buf BUF1 (N5534, N5525);
nor NOR2 (N5535, N5533, N828);
nand NAND2 (N5536, N5532, N1632);
nand NAND3 (N5537, N5531, N503, N796);
nand NAND3 (N5538, N5536, N1378, N996);
not NOT1 (N5539, N5537);
or OR4 (N5540, N5538, N43, N4174, N3115);
buf BUF1 (N5541, N5523);
buf BUF1 (N5542, N5493);
nor NOR4 (N5543, N5541, N5506, N2762, N2523);
or OR2 (N5544, N5539, N304);
or OR3 (N5545, N5529, N5459, N3531);
or OR4 (N5546, N5540, N2450, N878, N2411);
nor NOR4 (N5547, N5542, N5290, N1877, N589);
and AND2 (N5548, N5524, N557);
and AND2 (N5549, N5543, N1205);
or OR2 (N5550, N5546, N2494);
xor XOR2 (N5551, N5545, N1041);
or OR4 (N5552, N5544, N4448, N4586, N3073);
or OR4 (N5553, N5549, N3419, N1484, N1086);
not NOT1 (N5554, N5552);
nand NAND4 (N5555, N5547, N3113, N2352, N4103);
or OR4 (N5556, N5534, N2902, N2411, N1959);
or OR3 (N5557, N5535, N142, N3048);
nand NAND2 (N5558, N5528, N1955);
and AND3 (N5559, N5556, N851, N3962);
buf BUF1 (N5560, N5554);
xor XOR2 (N5561, N5515, N1161);
xor XOR2 (N5562, N5548, N525);
or OR3 (N5563, N5562, N2438, N1424);
and AND4 (N5564, N5558, N3824, N5335, N5189);
or OR3 (N5565, N5561, N1287, N355);
nor NOR3 (N5566, N5565, N467, N1998);
nor NOR4 (N5567, N5564, N117, N3376, N4688);
buf BUF1 (N5568, N5553);
buf BUF1 (N5569, N5567);
nand NAND4 (N5570, N5560, N5271, N2600, N3388);
and AND2 (N5571, N5551, N662);
and AND3 (N5572, N5571, N4665, N3678);
or OR4 (N5573, N5559, N3145, N1699, N4120);
nand NAND3 (N5574, N5555, N4223, N386);
not NOT1 (N5575, N5573);
nand NAND3 (N5576, N5575, N2440, N4846);
xor XOR2 (N5577, N5568, N1661);
nor NOR4 (N5578, N5570, N2057, N2761, N4343);
not NOT1 (N5579, N5576);
and AND2 (N5580, N5563, N3452);
not NOT1 (N5581, N5578);
nor NOR2 (N5582, N5557, N225);
xor XOR2 (N5583, N5569, N2984);
not NOT1 (N5584, N5583);
nor NOR4 (N5585, N5584, N1450, N4419, N3067);
nor NOR4 (N5586, N5577, N3699, N4723, N1582);
or OR3 (N5587, N5580, N4648, N1662);
xor XOR2 (N5588, N5579, N4437);
xor XOR2 (N5589, N5587, N5488);
not NOT1 (N5590, N5574);
xor XOR2 (N5591, N5566, N1669);
xor XOR2 (N5592, N5550, N521);
nand NAND3 (N5593, N5581, N206, N1862);
xor XOR2 (N5594, N5582, N1909);
nand NAND2 (N5595, N5594, N4528);
or OR4 (N5596, N5595, N5445, N4944, N2851);
not NOT1 (N5597, N5592);
and AND4 (N5598, N5591, N5389, N1254, N3981);
nor NOR4 (N5599, N5586, N3249, N2551, N5505);
xor XOR2 (N5600, N5590, N1759);
nor NOR3 (N5601, N5597, N3772, N4261);
or OR3 (N5602, N5589, N505, N3151);
not NOT1 (N5603, N5572);
buf BUF1 (N5604, N5602);
nor NOR2 (N5605, N5588, N5485);
or OR2 (N5606, N5604, N5137);
or OR3 (N5607, N5599, N554, N1119);
xor XOR2 (N5608, N5603, N2029);
or OR3 (N5609, N5606, N909, N4326);
or OR4 (N5610, N5600, N5107, N5007, N1507);
nor NOR4 (N5611, N5607, N435, N941, N964);
and AND3 (N5612, N5611, N4180, N3379);
and AND2 (N5613, N5601, N1083);
or OR3 (N5614, N5608, N1111, N3842);
nor NOR3 (N5615, N5593, N2774, N1545);
or OR2 (N5616, N5612, N2165);
nand NAND3 (N5617, N5613, N1377, N4220);
nor NOR3 (N5618, N5609, N597, N2258);
buf BUF1 (N5619, N5618);
not NOT1 (N5620, N5585);
xor XOR2 (N5621, N5620, N494);
nor NOR2 (N5622, N5616, N3794);
nor NOR3 (N5623, N5605, N1440, N5589);
not NOT1 (N5624, N5614);
and AND3 (N5625, N5596, N4828, N5310);
buf BUF1 (N5626, N5625);
nand NAND2 (N5627, N5598, N1581);
buf BUF1 (N5628, N5626);
not NOT1 (N5629, N5617);
not NOT1 (N5630, N5619);
buf BUF1 (N5631, N5629);
buf BUF1 (N5632, N5610);
buf BUF1 (N5633, N5622);
buf BUF1 (N5634, N5632);
buf BUF1 (N5635, N5624);
and AND2 (N5636, N5633, N5134);
nor NOR4 (N5637, N5623, N2542, N1161, N3284);
nand NAND3 (N5638, N5628, N2140, N401);
not NOT1 (N5639, N5631);
nor NOR3 (N5640, N5621, N3593, N3187);
not NOT1 (N5641, N5635);
or OR4 (N5642, N5637, N3423, N67, N2727);
and AND2 (N5643, N5627, N1985);
buf BUF1 (N5644, N5615);
xor XOR2 (N5645, N5638, N4312);
buf BUF1 (N5646, N5645);
buf BUF1 (N5647, N5636);
not NOT1 (N5648, N5641);
or OR2 (N5649, N5644, N600);
nand NAND4 (N5650, N5639, N4692, N2795, N906);
nor NOR3 (N5651, N5642, N3913, N5329);
xor XOR2 (N5652, N5634, N4351);
or OR3 (N5653, N5630, N1718, N4417);
xor XOR2 (N5654, N5640, N842);
not NOT1 (N5655, N5643);
nor NOR3 (N5656, N5652, N2632, N5151);
xor XOR2 (N5657, N5655, N3577);
nand NAND2 (N5658, N5649, N899);
buf BUF1 (N5659, N5656);
nand NAND4 (N5660, N5654, N3274, N5556, N3484);
nor NOR2 (N5661, N5658, N4812);
nor NOR2 (N5662, N5660, N363);
nand NAND2 (N5663, N5650, N5299);
nor NOR2 (N5664, N5653, N334);
nand NAND4 (N5665, N5664, N4888, N5099, N3816);
nand NAND2 (N5666, N5647, N5209);
not NOT1 (N5667, N5646);
and AND4 (N5668, N5667, N4068, N2250, N555);
buf BUF1 (N5669, N5657);
and AND4 (N5670, N5648, N4546, N3899, N3456);
buf BUF1 (N5671, N5666);
xor XOR2 (N5672, N5665, N4587);
not NOT1 (N5673, N5663);
or OR2 (N5674, N5668, N3556);
nor NOR4 (N5675, N5662, N2040, N4831, N4369);
not NOT1 (N5676, N5651);
or OR2 (N5677, N5671, N5228);
nor NOR3 (N5678, N5673, N5080, N5204);
and AND2 (N5679, N5675, N215);
not NOT1 (N5680, N5661);
not NOT1 (N5681, N5672);
xor XOR2 (N5682, N5674, N3064);
not NOT1 (N5683, N5679);
and AND2 (N5684, N5680, N4630);
not NOT1 (N5685, N5677);
nor NOR2 (N5686, N5684, N1880);
and AND4 (N5687, N5676, N3840, N2532, N1900);
xor XOR2 (N5688, N5686, N1930);
not NOT1 (N5689, N5685);
and AND4 (N5690, N5681, N614, N2573, N771);
nor NOR4 (N5691, N5682, N3284, N3962, N3479);
nor NOR2 (N5692, N5659, N1849);
xor XOR2 (N5693, N5692, N3020);
nand NAND3 (N5694, N5688, N1548, N5505);
nor NOR4 (N5695, N5694, N1654, N2625, N4718);
xor XOR2 (N5696, N5690, N2087);
nor NOR4 (N5697, N5683, N4526, N331, N4103);
and AND3 (N5698, N5696, N5545, N853);
or OR4 (N5699, N5670, N2083, N671, N5310);
not NOT1 (N5700, N5669);
nor NOR2 (N5701, N5678, N4048);
buf BUF1 (N5702, N5699);
and AND2 (N5703, N5698, N4472);
buf BUF1 (N5704, N5697);
xor XOR2 (N5705, N5695, N2025);
xor XOR2 (N5706, N5701, N3378);
xor XOR2 (N5707, N5700, N3102);
nand NAND3 (N5708, N5707, N2157, N2993);
or OR2 (N5709, N5706, N3136);
buf BUF1 (N5710, N5702);
nand NAND2 (N5711, N5708, N1417);
and AND3 (N5712, N5704, N3715, N5596);
nor NOR3 (N5713, N5687, N889, N2245);
xor XOR2 (N5714, N5693, N5003);
nor NOR2 (N5715, N5705, N3697);
and AND3 (N5716, N5709, N2791, N1776);
buf BUF1 (N5717, N5703);
and AND3 (N5718, N5715, N2165, N2886);
not NOT1 (N5719, N5691);
or OR4 (N5720, N5719, N2859, N3391, N5154);
nor NOR2 (N5721, N5713, N5116);
or OR4 (N5722, N5716, N2478, N5315, N4803);
and AND2 (N5723, N5720, N3543);
xor XOR2 (N5724, N5689, N2230);
buf BUF1 (N5725, N5723);
xor XOR2 (N5726, N5714, N3699);
nor NOR2 (N5727, N5721, N246);
and AND3 (N5728, N5718, N3492, N3);
nand NAND3 (N5729, N5722, N633, N2115);
nand NAND3 (N5730, N5727, N4663, N552);
not NOT1 (N5731, N5712);
nor NOR4 (N5732, N5724, N5163, N76, N2051);
nor NOR2 (N5733, N5726, N5174);
nor NOR3 (N5734, N5711, N3713, N320);
nor NOR4 (N5735, N5729, N131, N4860, N4050);
nor NOR2 (N5736, N5728, N4408);
nand NAND4 (N5737, N5733, N4555, N5287, N5335);
and AND4 (N5738, N5725, N644, N5542, N246);
nor NOR4 (N5739, N5731, N2796, N2738, N942);
xor XOR2 (N5740, N5735, N1951);
not NOT1 (N5741, N5736);
or OR4 (N5742, N5710, N241, N5537, N4180);
buf BUF1 (N5743, N5738);
xor XOR2 (N5744, N5741, N1734);
buf BUF1 (N5745, N5737);
and AND2 (N5746, N5739, N2400);
or OR4 (N5747, N5745, N14, N275, N3274);
not NOT1 (N5748, N5730);
nand NAND2 (N5749, N5747, N2999);
or OR4 (N5750, N5746, N3698, N4053, N2353);
and AND3 (N5751, N5743, N1462, N5528);
nand NAND2 (N5752, N5742, N5343);
not NOT1 (N5753, N5752);
and AND2 (N5754, N5717, N4835);
or OR3 (N5755, N5744, N856, N5133);
buf BUF1 (N5756, N5734);
and AND2 (N5757, N5749, N1656);
or OR4 (N5758, N5750, N5546, N89, N2515);
and AND3 (N5759, N5756, N2961, N2953);
and AND3 (N5760, N5740, N376, N2039);
not NOT1 (N5761, N5760);
or OR4 (N5762, N5753, N4329, N158, N5118);
and AND3 (N5763, N5754, N260, N1557);
nand NAND4 (N5764, N5751, N3717, N4628, N1024);
buf BUF1 (N5765, N5757);
or OR2 (N5766, N5763, N3613);
nand NAND3 (N5767, N5732, N1191, N4694);
nor NOR4 (N5768, N5761, N2848, N3622, N1069);
nor NOR3 (N5769, N5764, N4255, N3559);
nand NAND3 (N5770, N5765, N1818, N4382);
nand NAND3 (N5771, N5769, N2281, N730);
and AND2 (N5772, N5768, N1789);
nor NOR3 (N5773, N5766, N2957, N4447);
nor NOR4 (N5774, N5771, N728, N554, N3377);
nand NAND4 (N5775, N5774, N1864, N2049, N1502);
and AND2 (N5776, N5773, N2078);
nor NOR2 (N5777, N5775, N449);
nor NOR3 (N5778, N5772, N5153, N4700);
nor NOR2 (N5779, N5755, N5269);
nor NOR4 (N5780, N5778, N320, N4724, N3381);
xor XOR2 (N5781, N5748, N4113);
nand NAND3 (N5782, N5777, N1931, N3164);
or OR2 (N5783, N5781, N1390);
nand NAND2 (N5784, N5780, N1053);
nor NOR3 (N5785, N5770, N2552, N3862);
not NOT1 (N5786, N5785);
or OR3 (N5787, N5759, N2086, N4983);
or OR3 (N5788, N5776, N3274, N2085);
nor NOR2 (N5789, N5786, N2325);
or OR2 (N5790, N5762, N122);
or OR4 (N5791, N5790, N5037, N625, N838);
nand NAND4 (N5792, N5788, N2752, N2762, N4453);
and AND3 (N5793, N5784, N2575, N2437);
and AND4 (N5794, N5767, N1364, N4629, N4846);
or OR2 (N5795, N5787, N4804);
xor XOR2 (N5796, N5782, N530);
xor XOR2 (N5797, N5792, N132);
nand NAND2 (N5798, N5791, N3493);
nor NOR2 (N5799, N5797, N4349);
or OR4 (N5800, N5779, N944, N3377, N2259);
nand NAND4 (N5801, N5789, N380, N2589, N1705);
xor XOR2 (N5802, N5795, N884);
nand NAND2 (N5803, N5800, N3937);
and AND4 (N5804, N5798, N886, N10, N5171);
and AND4 (N5805, N5783, N215, N4126, N1595);
buf BUF1 (N5806, N5758);
xor XOR2 (N5807, N5804, N3534);
xor XOR2 (N5808, N5805, N2746);
buf BUF1 (N5809, N5808);
nor NOR2 (N5810, N5794, N5396);
or OR4 (N5811, N5802, N3099, N2393, N1488);
nand NAND2 (N5812, N5803, N3775);
nand NAND4 (N5813, N5812, N5448, N1119, N2984);
xor XOR2 (N5814, N5806, N1742);
not NOT1 (N5815, N5813);
xor XOR2 (N5816, N5811, N1454);
not NOT1 (N5817, N5801);
not NOT1 (N5818, N5810);
not NOT1 (N5819, N5809);
nor NOR3 (N5820, N5814, N2296, N3806);
xor XOR2 (N5821, N5819, N4505);
or OR4 (N5822, N5799, N4357, N4118, N4013);
nor NOR3 (N5823, N5796, N1958, N343);
and AND2 (N5824, N5822, N1318);
buf BUF1 (N5825, N5793);
or OR2 (N5826, N5815, N5673);
xor XOR2 (N5827, N5816, N301);
or OR3 (N5828, N5826, N1026, N3619);
buf BUF1 (N5829, N5820);
or OR4 (N5830, N5829, N4061, N1313, N4933);
and AND3 (N5831, N5824, N2878, N84);
xor XOR2 (N5832, N5807, N2050);
or OR4 (N5833, N5821, N1125, N4786, N822);
nor NOR4 (N5834, N5831, N5181, N676, N551);
and AND2 (N5835, N5834, N4528);
not NOT1 (N5836, N5823);
nor NOR4 (N5837, N5818, N758, N750, N4057);
not NOT1 (N5838, N5833);
not NOT1 (N5839, N5827);
xor XOR2 (N5840, N5839, N4673);
nor NOR2 (N5841, N5830, N3620);
nor NOR2 (N5842, N5835, N1688);
not NOT1 (N5843, N5842);
not NOT1 (N5844, N5840);
nand NAND4 (N5845, N5843, N2098, N5421, N3229);
or OR4 (N5846, N5838, N4491, N3681, N492);
nor NOR3 (N5847, N5845, N4625, N2091);
nor NOR3 (N5848, N5832, N2048, N106);
and AND3 (N5849, N5817, N1657, N5506);
nor NOR4 (N5850, N5836, N2148, N3113, N1284);
buf BUF1 (N5851, N5837);
xor XOR2 (N5852, N5851, N4636);
not NOT1 (N5853, N5847);
or OR2 (N5854, N5848, N2957);
and AND4 (N5855, N5850, N1430, N2921, N100);
nand NAND2 (N5856, N5855, N949);
buf BUF1 (N5857, N5856);
nor NOR2 (N5858, N5857, N2488);
buf BUF1 (N5859, N5858);
nand NAND2 (N5860, N5854, N3731);
not NOT1 (N5861, N5828);
buf BUF1 (N5862, N5859);
nand NAND2 (N5863, N5846, N3082);
buf BUF1 (N5864, N5863);
nand NAND4 (N5865, N5864, N5336, N1946, N1718);
nand NAND4 (N5866, N5853, N3516, N2948, N1156);
nand NAND2 (N5867, N5841, N1343);
nand NAND2 (N5868, N5849, N1074);
nand NAND4 (N5869, N5868, N1954, N5403, N2870);
xor XOR2 (N5870, N5860, N662);
not NOT1 (N5871, N5867);
and AND4 (N5872, N5870, N2576, N3094, N1117);
nor NOR4 (N5873, N5825, N3999, N1054, N4688);
buf BUF1 (N5874, N5869);
and AND4 (N5875, N5873, N2338, N2091, N5865);
or OR2 (N5876, N5426, N1626);
or OR4 (N5877, N5871, N5322, N570, N3195);
nand NAND4 (N5878, N5861, N5527, N780, N5307);
buf BUF1 (N5879, N5862);
xor XOR2 (N5880, N5876, N596);
nand NAND3 (N5881, N5879, N4393, N4025);
or OR2 (N5882, N5878, N3020);
nand NAND2 (N5883, N5866, N5706);
xor XOR2 (N5884, N5883, N4666);
xor XOR2 (N5885, N5844, N2054);
xor XOR2 (N5886, N5881, N3772);
nand NAND2 (N5887, N5885, N2890);
nor NOR4 (N5888, N5875, N2849, N1377, N1433);
buf BUF1 (N5889, N5886);
and AND2 (N5890, N5887, N3370);
and AND3 (N5891, N5874, N2642, N3409);
and AND4 (N5892, N5890, N3828, N1392, N4565);
nor NOR3 (N5893, N5872, N2698, N5560);
xor XOR2 (N5894, N5884, N2973);
xor XOR2 (N5895, N5891, N3454);
nor NOR3 (N5896, N5882, N1443, N5453);
or OR2 (N5897, N5894, N5730);
or OR3 (N5898, N5888, N2372, N2535);
xor XOR2 (N5899, N5893, N4837);
xor XOR2 (N5900, N5898, N5077);
or OR4 (N5901, N5880, N5565, N4256, N3277);
nand NAND4 (N5902, N5877, N5873, N4402, N1365);
nor NOR4 (N5903, N5897, N603, N4221, N374);
or OR2 (N5904, N5901, N3530);
nor NOR3 (N5905, N5903, N2692, N3032);
and AND4 (N5906, N5899, N225, N3886, N1592);
and AND4 (N5907, N5892, N2583, N3550, N3125);
xor XOR2 (N5908, N5902, N299);
buf BUF1 (N5909, N5895);
buf BUF1 (N5910, N5906);
or OR2 (N5911, N5908, N1869);
or OR2 (N5912, N5905, N1238);
and AND3 (N5913, N5912, N3705, N5428);
or OR2 (N5914, N5909, N4543);
nand NAND2 (N5915, N5904, N3097);
nor NOR2 (N5916, N5915, N1435);
nand NAND2 (N5917, N5910, N1987);
and AND2 (N5918, N5900, N5741);
buf BUF1 (N5919, N5918);
and AND3 (N5920, N5916, N4794, N4270);
xor XOR2 (N5921, N5852, N211);
or OR3 (N5922, N5913, N5402, N5463);
xor XOR2 (N5923, N5911, N2716);
nand NAND2 (N5924, N5896, N5436);
not NOT1 (N5925, N5917);
or OR2 (N5926, N5907, N5305);
buf BUF1 (N5927, N5922);
nand NAND2 (N5928, N5919, N3353);
or OR3 (N5929, N5927, N1213, N4787);
not NOT1 (N5930, N5921);
buf BUF1 (N5931, N5920);
and AND2 (N5932, N5928, N5144);
nand NAND4 (N5933, N5930, N3168, N3349, N4397);
not NOT1 (N5934, N5929);
nand NAND2 (N5935, N5923, N1541);
not NOT1 (N5936, N5933);
and AND4 (N5937, N5926, N3932, N4637, N4398);
buf BUF1 (N5938, N5934);
xor XOR2 (N5939, N5935, N3023);
and AND4 (N5940, N5925, N3638, N1661, N3049);
or OR3 (N5941, N5940, N2254, N581);
nor NOR4 (N5942, N5938, N3865, N2654, N650);
or OR4 (N5943, N5939, N458, N4400, N3842);
not NOT1 (N5944, N5889);
not NOT1 (N5945, N5942);
buf BUF1 (N5946, N5944);
nand NAND2 (N5947, N5924, N4367);
and AND4 (N5948, N5941, N353, N2362, N2877);
and AND4 (N5949, N5947, N3904, N1749, N2736);
nor NOR3 (N5950, N5948, N903, N131);
nand NAND3 (N5951, N5937, N2142, N3101);
nor NOR3 (N5952, N5936, N1622, N3060);
not NOT1 (N5953, N5949);
or OR3 (N5954, N5943, N4948, N4999);
nand NAND4 (N5955, N5951, N2427, N5113, N103);
not NOT1 (N5956, N5945);
xor XOR2 (N5957, N5914, N5781);
and AND3 (N5958, N5953, N48, N1732);
nand NAND4 (N5959, N5950, N3005, N2631, N2183);
and AND2 (N5960, N5946, N2078);
and AND2 (N5961, N5960, N2616);
xor XOR2 (N5962, N5956, N1140);
and AND4 (N5963, N5962, N4395, N232, N1114);
nand NAND4 (N5964, N5931, N2602, N1320, N898);
or OR4 (N5965, N5964, N2571, N1031, N4887);
nor NOR4 (N5966, N5965, N1234, N5660, N3963);
nor NOR2 (N5967, N5959, N1039);
and AND4 (N5968, N5932, N1336, N5821, N4518);
and AND4 (N5969, N5954, N5812, N528, N5137);
nor NOR3 (N5970, N5958, N807, N4044);
nor NOR2 (N5971, N5963, N3872);
buf BUF1 (N5972, N5957);
and AND2 (N5973, N5969, N2583);
buf BUF1 (N5974, N5971);
nor NOR3 (N5975, N5966, N4724, N4054);
nand NAND3 (N5976, N5968, N1824, N3295);
nor NOR4 (N5977, N5970, N4762, N971, N2572);
and AND2 (N5978, N5961, N5328);
nor NOR3 (N5979, N5978, N3011, N4766);
nor NOR3 (N5980, N5967, N4708, N5758);
xor XOR2 (N5981, N5972, N1674);
nor NOR4 (N5982, N5976, N3781, N4080, N165);
and AND4 (N5983, N5980, N3653, N4214, N5085);
nor NOR3 (N5984, N5982, N3213, N4170);
nor NOR4 (N5985, N5974, N1402, N5323, N3853);
nor NOR4 (N5986, N5985, N2023, N2616, N4917);
xor XOR2 (N5987, N5979, N1888);
and AND2 (N5988, N5973, N296);
nor NOR2 (N5989, N5955, N1177);
buf BUF1 (N5990, N5952);
not NOT1 (N5991, N5988);
nand NAND4 (N5992, N5986, N1795, N5989, N412);
not NOT1 (N5993, N1869);
xor XOR2 (N5994, N5975, N5183);
and AND3 (N5995, N5992, N3882, N4293);
or OR2 (N5996, N5993, N4762);
or OR3 (N5997, N5996, N730, N1953);
not NOT1 (N5998, N5983);
xor XOR2 (N5999, N5997, N4696);
xor XOR2 (N6000, N5999, N3996);
not NOT1 (N6001, N5995);
and AND3 (N6002, N5984, N3714, N1966);
xor XOR2 (N6003, N6001, N260);
nand NAND3 (N6004, N5990, N5965, N2544);
or OR2 (N6005, N6002, N2628);
nor NOR4 (N6006, N5998, N2653, N1295, N4181);
nor NOR2 (N6007, N5981, N2881);
nand NAND4 (N6008, N6000, N2401, N2003, N2672);
not NOT1 (N6009, N6004);
or OR4 (N6010, N6007, N5251, N2248, N3634);
buf BUF1 (N6011, N6010);
not NOT1 (N6012, N5994);
nor NOR4 (N6013, N5977, N3833, N518, N4021);
and AND2 (N6014, N6008, N5577);
buf BUF1 (N6015, N6006);
or OR2 (N6016, N6003, N4599);
or OR2 (N6017, N5991, N3101);
or OR2 (N6018, N6013, N126);
nor NOR3 (N6019, N6005, N3354, N1792);
buf BUF1 (N6020, N6016);
nor NOR4 (N6021, N6018, N1797, N1068, N377);
not NOT1 (N6022, N6021);
buf BUF1 (N6023, N6014);
or OR3 (N6024, N6017, N2551, N4415);
buf BUF1 (N6025, N6022);
buf BUF1 (N6026, N6025);
nand NAND4 (N6027, N6019, N1713, N1642, N431);
nand NAND4 (N6028, N6012, N2586, N5109, N2017);
xor XOR2 (N6029, N6026, N527);
and AND3 (N6030, N6015, N5968, N1069);
buf BUF1 (N6031, N6030);
not NOT1 (N6032, N6029);
xor XOR2 (N6033, N6027, N5630);
buf BUF1 (N6034, N6033);
nand NAND3 (N6035, N6020, N2270, N3760);
and AND4 (N6036, N6011, N153, N4012, N2098);
and AND2 (N6037, N5987, N3937);
xor XOR2 (N6038, N6024, N287);
not NOT1 (N6039, N6034);
and AND4 (N6040, N6039, N2495, N4418, N5515);
or OR3 (N6041, N6023, N4073, N5256);
buf BUF1 (N6042, N6040);
or OR4 (N6043, N6038, N3258, N782, N2119);
buf BUF1 (N6044, N6031);
xor XOR2 (N6045, N6043, N1397);
nor NOR4 (N6046, N6041, N4348, N5798, N5167);
buf BUF1 (N6047, N6046);
not NOT1 (N6048, N6032);
and AND4 (N6049, N6045, N4219, N5490, N2878);
not NOT1 (N6050, N6049);
xor XOR2 (N6051, N6050, N4191);
xor XOR2 (N6052, N6044, N338);
or OR3 (N6053, N6009, N534, N2603);
buf BUF1 (N6054, N6048);
or OR4 (N6055, N6042, N5831, N1203, N2749);
and AND2 (N6056, N6054, N2344);
or OR4 (N6057, N6051, N5838, N3297, N3538);
not NOT1 (N6058, N6035);
nand NAND4 (N6059, N6057, N5521, N1611, N5390);
not NOT1 (N6060, N6036);
nand NAND2 (N6061, N6059, N881);
nand NAND2 (N6062, N6053, N5132);
not NOT1 (N6063, N6060);
xor XOR2 (N6064, N6047, N128);
xor XOR2 (N6065, N6056, N50);
and AND2 (N6066, N6055, N2939);
buf BUF1 (N6067, N6064);
or OR4 (N6068, N6062, N1941, N2987, N3590);
and AND4 (N6069, N6037, N4251, N1784, N2723);
and AND3 (N6070, N6066, N2038, N1261);
or OR4 (N6071, N6069, N58, N5613, N4058);
buf BUF1 (N6072, N6071);
and AND2 (N6073, N6063, N2391);
not NOT1 (N6074, N6065);
xor XOR2 (N6075, N6052, N5114);
nand NAND3 (N6076, N6070, N3415, N60);
or OR2 (N6077, N6058, N2166);
not NOT1 (N6078, N6028);
nand NAND2 (N6079, N6067, N4889);
nor NOR2 (N6080, N6061, N3616);
nand NAND4 (N6081, N6068, N3285, N3586, N4426);
or OR3 (N6082, N6073, N1537, N5558);
not NOT1 (N6083, N6072);
buf BUF1 (N6084, N6078);
or OR3 (N6085, N6083, N3712, N5663);
or OR4 (N6086, N6079, N3517, N586, N1279);
buf BUF1 (N6087, N6077);
nor NOR3 (N6088, N6086, N1675, N2057);
or OR2 (N6089, N6074, N1866);
buf BUF1 (N6090, N6080);
or OR2 (N6091, N6090, N978);
xor XOR2 (N6092, N6089, N2817);
nand NAND2 (N6093, N6076, N1083);
xor XOR2 (N6094, N6082, N5957);
not NOT1 (N6095, N6092);
not NOT1 (N6096, N6094);
nor NOR4 (N6097, N6084, N5017, N3848, N4630);
xor XOR2 (N6098, N6093, N2457);
xor XOR2 (N6099, N6087, N5799);
or OR2 (N6100, N6096, N3439);
nor NOR3 (N6101, N6081, N466, N4530);
xor XOR2 (N6102, N6091, N1392);
or OR3 (N6103, N6088, N4619, N4362);
nor NOR3 (N6104, N6097, N5864, N3699);
or OR3 (N6105, N6100, N5088, N2040);
not NOT1 (N6106, N6095);
xor XOR2 (N6107, N6099, N1034);
buf BUF1 (N6108, N6075);
xor XOR2 (N6109, N6102, N257);
buf BUF1 (N6110, N6108);
buf BUF1 (N6111, N6103);
not NOT1 (N6112, N6111);
not NOT1 (N6113, N6109);
buf BUF1 (N6114, N6105);
nand NAND4 (N6115, N6114, N5507, N4106, N4753);
and AND2 (N6116, N6115, N2300);
and AND4 (N6117, N6107, N4600, N1746, N863);
nor NOR2 (N6118, N6117, N5299);
nor NOR4 (N6119, N6085, N513, N3040, N1777);
and AND2 (N6120, N6116, N2962);
or OR4 (N6121, N6101, N3089, N3119, N677);
or OR4 (N6122, N6112, N4589, N2268, N703);
and AND4 (N6123, N6121, N3279, N68, N4657);
nor NOR3 (N6124, N6118, N1503, N5333);
nand NAND4 (N6125, N6113, N1865, N1991, N5412);
xor XOR2 (N6126, N6120, N3704);
xor XOR2 (N6127, N6126, N4120);
xor XOR2 (N6128, N6125, N4747);
nand NAND3 (N6129, N6124, N285, N3979);
xor XOR2 (N6130, N6123, N1173);
or OR4 (N6131, N6110, N5131, N3265, N3134);
nand NAND2 (N6132, N6130, N511);
and AND4 (N6133, N6131, N705, N4098, N2563);
and AND2 (N6134, N6106, N4092);
nor NOR4 (N6135, N6133, N3593, N4144, N822);
xor XOR2 (N6136, N6098, N3649);
buf BUF1 (N6137, N6127);
and AND3 (N6138, N6122, N3174, N2515);
nor NOR3 (N6139, N6132, N2771, N2269);
nor NOR3 (N6140, N6128, N4803, N2138);
xor XOR2 (N6141, N6138, N4579);
nor NOR2 (N6142, N6135, N1550);
xor XOR2 (N6143, N6119, N4113);
buf BUF1 (N6144, N6136);
and AND2 (N6145, N6142, N2934);
buf BUF1 (N6146, N6129);
nor NOR3 (N6147, N6143, N4986, N901);
and AND3 (N6148, N6104, N2826, N2221);
nand NAND4 (N6149, N6146, N2068, N464, N3754);
and AND2 (N6150, N6149, N5340);
xor XOR2 (N6151, N6140, N4250);
nand NAND4 (N6152, N6137, N1688, N5405, N1967);
or OR4 (N6153, N6150, N6139, N726, N1202);
xor XOR2 (N6154, N1149, N6151);
not NOT1 (N6155, N388);
nand NAND3 (N6156, N6134, N1162, N1970);
not NOT1 (N6157, N6152);
nor NOR2 (N6158, N6148, N2981);
not NOT1 (N6159, N6156);
and AND4 (N6160, N6159, N4977, N4299, N1213);
and AND2 (N6161, N6147, N86);
nand NAND3 (N6162, N6158, N3471, N466);
nor NOR2 (N6163, N6161, N4552);
buf BUF1 (N6164, N6163);
buf BUF1 (N6165, N6160);
or OR4 (N6166, N6145, N736, N5202, N5233);
or OR3 (N6167, N6164, N3486, N228);
nand NAND3 (N6168, N6154, N6115, N1973);
nand NAND4 (N6169, N6155, N2276, N2130, N6007);
nor NOR4 (N6170, N6153, N3992, N4260, N3498);
or OR2 (N6171, N6157, N1861);
nor NOR2 (N6172, N6162, N2771);
not NOT1 (N6173, N6165);
buf BUF1 (N6174, N6169);
and AND3 (N6175, N6170, N643, N4390);
xor XOR2 (N6176, N6166, N3265);
xor XOR2 (N6177, N6173, N1416);
xor XOR2 (N6178, N6141, N3742);
nand NAND3 (N6179, N6144, N5000, N208);
or OR2 (N6180, N6174, N594);
not NOT1 (N6181, N6180);
nor NOR4 (N6182, N6179, N1520, N2969, N3172);
or OR3 (N6183, N6178, N960, N740);
nand NAND2 (N6184, N6167, N5264);
not NOT1 (N6185, N6184);
nor NOR2 (N6186, N6185, N3534);
and AND2 (N6187, N6177, N3475);
xor XOR2 (N6188, N6168, N1372);
or OR4 (N6189, N6171, N108, N3848, N2262);
or OR3 (N6190, N6189, N4298, N2258);
nand NAND4 (N6191, N6181, N1271, N30, N4010);
not NOT1 (N6192, N6188);
buf BUF1 (N6193, N6183);
buf BUF1 (N6194, N6192);
not NOT1 (N6195, N6186);
nor NOR4 (N6196, N6176, N1698, N38, N2717);
xor XOR2 (N6197, N6195, N3428);
nor NOR2 (N6198, N6187, N316);
or OR3 (N6199, N6194, N4995, N5374);
buf BUF1 (N6200, N6197);
or OR2 (N6201, N6196, N5527);
and AND4 (N6202, N6198, N2522, N1574, N83);
nor NOR4 (N6203, N6201, N1886, N3612, N3933);
xor XOR2 (N6204, N6175, N524);
xor XOR2 (N6205, N6199, N4785);
or OR4 (N6206, N6190, N3990, N5999, N6123);
or OR4 (N6207, N6182, N532, N1222, N1731);
xor XOR2 (N6208, N6206, N1801);
nand NAND2 (N6209, N6172, N2747);
xor XOR2 (N6210, N6200, N4432);
nand NAND3 (N6211, N6202, N1950, N3795);
and AND4 (N6212, N6191, N1332, N5213, N686);
not NOT1 (N6213, N6193);
nand NAND2 (N6214, N6208, N770);
or OR4 (N6215, N6205, N6077, N3048, N962);
nor NOR3 (N6216, N6213, N3310, N675);
and AND3 (N6217, N6211, N5607, N5867);
buf BUF1 (N6218, N6203);
not NOT1 (N6219, N6204);
buf BUF1 (N6220, N6212);
buf BUF1 (N6221, N6207);
xor XOR2 (N6222, N6220, N3240);
nand NAND4 (N6223, N6219, N2035, N5942, N1572);
nor NOR2 (N6224, N6221, N448);
xor XOR2 (N6225, N6209, N4209);
nand NAND3 (N6226, N6210, N159, N4976);
buf BUF1 (N6227, N6224);
xor XOR2 (N6228, N6218, N3400);
not NOT1 (N6229, N6223);
or OR4 (N6230, N6228, N2551, N2129, N329);
not NOT1 (N6231, N6226);
and AND2 (N6232, N6227, N5632);
and AND3 (N6233, N6214, N1639, N4781);
buf BUF1 (N6234, N6232);
nor NOR4 (N6235, N6222, N2505, N2420, N4809);
nand NAND2 (N6236, N6216, N408);
not NOT1 (N6237, N6215);
nand NAND2 (N6238, N6231, N4743);
not NOT1 (N6239, N6217);
and AND4 (N6240, N6233, N3444, N5069, N3527);
nor NOR2 (N6241, N6234, N6189);
or OR2 (N6242, N6241, N941);
nor NOR3 (N6243, N6240, N1612, N2822);
nand NAND4 (N6244, N6238, N3926, N1294, N616);
nor NOR4 (N6245, N6239, N253, N550, N2892);
or OR3 (N6246, N6243, N2659, N1009);
and AND4 (N6247, N6245, N260, N1118, N4309);
nor NOR2 (N6248, N6244, N1463);
xor XOR2 (N6249, N6246, N294);
nand NAND4 (N6250, N6236, N4194, N2366, N5182);
buf BUF1 (N6251, N6229);
and AND2 (N6252, N6235, N4063);
nand NAND2 (N6253, N6242, N3603);
not NOT1 (N6254, N6251);
or OR4 (N6255, N6252, N829, N4664, N2986);
not NOT1 (N6256, N6237);
or OR4 (N6257, N6254, N1393, N2631, N3278);
and AND2 (N6258, N6247, N3057);
xor XOR2 (N6259, N6258, N3755);
or OR4 (N6260, N6259, N2336, N1628, N1445);
and AND2 (N6261, N6249, N1300);
buf BUF1 (N6262, N6225);
nor NOR3 (N6263, N6260, N4043, N5996);
xor XOR2 (N6264, N6255, N3717);
xor XOR2 (N6265, N6264, N2058);
nand NAND2 (N6266, N6257, N3381);
nor NOR3 (N6267, N6266, N4565, N4110);
or OR3 (N6268, N6230, N3309, N5789);
not NOT1 (N6269, N6263);
not NOT1 (N6270, N6269);
and AND2 (N6271, N6262, N2164);
nand NAND2 (N6272, N6248, N1074);
xor XOR2 (N6273, N6265, N1162);
or OR2 (N6274, N6270, N1825);
nor NOR4 (N6275, N6274, N2090, N2083, N5464);
not NOT1 (N6276, N6253);
nor NOR4 (N6277, N6261, N1719, N4548, N493);
nand NAND3 (N6278, N6275, N3051, N6095);
xor XOR2 (N6279, N6268, N2440);
nand NAND4 (N6280, N6279, N2975, N6223, N1832);
and AND2 (N6281, N6256, N1920);
buf BUF1 (N6282, N6281);
buf BUF1 (N6283, N6277);
buf BUF1 (N6284, N6273);
nor NOR4 (N6285, N6271, N4276, N3344, N2138);
nor NOR2 (N6286, N6272, N5771);
and AND2 (N6287, N6250, N2994);
nand NAND2 (N6288, N6280, N1394);
or OR2 (N6289, N6285, N1447);
xor XOR2 (N6290, N6267, N2715);
nand NAND4 (N6291, N6283, N5434, N1137, N2245);
not NOT1 (N6292, N6290);
nand NAND4 (N6293, N6278, N3067, N2172, N4319);
buf BUF1 (N6294, N6286);
not NOT1 (N6295, N6293);
not NOT1 (N6296, N6289);
and AND2 (N6297, N6287, N534);
or OR2 (N6298, N6276, N6142);
buf BUF1 (N6299, N6284);
buf BUF1 (N6300, N6299);
not NOT1 (N6301, N6295);
nor NOR4 (N6302, N6298, N5106, N253, N2057);
nand NAND3 (N6303, N6294, N6181, N5657);
not NOT1 (N6304, N6297);
or OR3 (N6305, N6300, N745, N1291);
or OR2 (N6306, N6304, N5288);
or OR3 (N6307, N6296, N5697, N5627);
not NOT1 (N6308, N6291);
and AND3 (N6309, N6302, N6029, N6251);
buf BUF1 (N6310, N6288);
or OR4 (N6311, N6282, N5048, N5707, N3361);
nand NAND2 (N6312, N6303, N1478);
and AND4 (N6313, N6309, N5699, N3951, N855);
buf BUF1 (N6314, N6308);
or OR4 (N6315, N6312, N3552, N2821, N269);
buf BUF1 (N6316, N6301);
nand NAND3 (N6317, N6311, N810, N5211);
nand NAND4 (N6318, N6314, N1488, N1803, N1092);
and AND3 (N6319, N6313, N475, N4719);
nor NOR4 (N6320, N6319, N4910, N4948, N2385);
xor XOR2 (N6321, N6307, N5179);
or OR2 (N6322, N6310, N5340);
buf BUF1 (N6323, N6322);
xor XOR2 (N6324, N6292, N187);
xor XOR2 (N6325, N6318, N3494);
nor NOR4 (N6326, N6325, N2257, N313, N2580);
not NOT1 (N6327, N6323);
buf BUF1 (N6328, N6305);
nand NAND3 (N6329, N6328, N5526, N1606);
buf BUF1 (N6330, N6306);
or OR4 (N6331, N6330, N4651, N2743, N3375);
and AND4 (N6332, N6321, N2238, N2705, N5161);
not NOT1 (N6333, N6332);
not NOT1 (N6334, N6316);
or OR3 (N6335, N6317, N2589, N2604);
nor NOR4 (N6336, N6320, N4302, N2519, N5232);
and AND3 (N6337, N6329, N3002, N818);
and AND2 (N6338, N6336, N351);
nand NAND3 (N6339, N6326, N314, N6244);
or OR4 (N6340, N6335, N4014, N4252, N1262);
not NOT1 (N6341, N6337);
or OR2 (N6342, N6327, N4644);
nand NAND3 (N6343, N6334, N2328, N4041);
or OR2 (N6344, N6331, N6114);
nor NOR4 (N6345, N6344, N785, N1424, N1105);
buf BUF1 (N6346, N6345);
or OR4 (N6347, N6346, N23, N3324, N637);
or OR3 (N6348, N6341, N3601, N1998);
and AND4 (N6349, N6347, N4739, N1240, N4688);
or OR4 (N6350, N6349, N3747, N3129, N3220);
nand NAND3 (N6351, N6338, N2923, N1158);
or OR4 (N6352, N6348, N2221, N2819, N2067);
buf BUF1 (N6353, N6333);
xor XOR2 (N6354, N6352, N2929);
xor XOR2 (N6355, N6339, N5053);
xor XOR2 (N6356, N6342, N5180);
nand NAND3 (N6357, N6353, N3917, N1876);
nand NAND2 (N6358, N6351, N4330);
nand NAND4 (N6359, N6324, N4042, N1942, N1323);
and AND4 (N6360, N6315, N5361, N4186, N1443);
nor NOR4 (N6361, N6343, N2812, N3376, N1079);
xor XOR2 (N6362, N6359, N5391);
buf BUF1 (N6363, N6360);
and AND2 (N6364, N6363, N4273);
and AND2 (N6365, N6358, N6057);
and AND2 (N6366, N6340, N3520);
or OR2 (N6367, N6362, N1814);
xor XOR2 (N6368, N6366, N5203);
not NOT1 (N6369, N6368);
and AND2 (N6370, N6357, N5024);
or OR2 (N6371, N6364, N3747);
or OR2 (N6372, N6369, N4354);
xor XOR2 (N6373, N6355, N908);
or OR3 (N6374, N6370, N138, N244);
and AND3 (N6375, N6367, N3541, N727);
xor XOR2 (N6376, N6354, N4692);
not NOT1 (N6377, N6374);
xor XOR2 (N6378, N6373, N893);
and AND3 (N6379, N6376, N3532, N6143);
not NOT1 (N6380, N6375);
xor XOR2 (N6381, N6371, N4456);
or OR2 (N6382, N6381, N20);
not NOT1 (N6383, N6372);
nand NAND2 (N6384, N6365, N4109);
buf BUF1 (N6385, N6380);
and AND2 (N6386, N6356, N2086);
buf BUF1 (N6387, N6379);
or OR3 (N6388, N6387, N5310, N5416);
or OR4 (N6389, N6361, N3981, N3377, N4804);
or OR2 (N6390, N6386, N6014);
and AND2 (N6391, N6377, N5379);
not NOT1 (N6392, N6384);
xor XOR2 (N6393, N6382, N2328);
or OR3 (N6394, N6383, N2086, N2515);
nand NAND2 (N6395, N6385, N5854);
nand NAND3 (N6396, N6388, N3261, N6108);
not NOT1 (N6397, N6393);
nor NOR3 (N6398, N6392, N1138, N1045);
not NOT1 (N6399, N6378);
nand NAND2 (N6400, N6389, N4690);
nand NAND3 (N6401, N6395, N5522, N5757);
xor XOR2 (N6402, N6390, N6128);
nor NOR4 (N6403, N6396, N4328, N5041, N1280);
nand NAND3 (N6404, N6350, N1316, N3282);
or OR2 (N6405, N6400, N3324);
xor XOR2 (N6406, N6394, N4095);
xor XOR2 (N6407, N6397, N3393);
nor NOR2 (N6408, N6404, N5847);
or OR2 (N6409, N6406, N4520);
or OR4 (N6410, N6391, N2617, N4817, N1632);
and AND3 (N6411, N6407, N2402, N3699);
or OR2 (N6412, N6408, N1531);
buf BUF1 (N6413, N6403);
not NOT1 (N6414, N6411);
and AND3 (N6415, N6412, N57, N1499);
nand NAND3 (N6416, N6409, N1800, N4838);
buf BUF1 (N6417, N6413);
nand NAND4 (N6418, N6417, N3625, N700, N4624);
nor NOR3 (N6419, N6418, N355, N590);
or OR3 (N6420, N6401, N5811, N4248);
buf BUF1 (N6421, N6405);
xor XOR2 (N6422, N6410, N473);
xor XOR2 (N6423, N6421, N2266);
buf BUF1 (N6424, N6399);
nor NOR3 (N6425, N6402, N4166, N4749);
not NOT1 (N6426, N6416);
nor NOR2 (N6427, N6425, N2173);
not NOT1 (N6428, N6424);
and AND4 (N6429, N6423, N5533, N3477, N1332);
not NOT1 (N6430, N6429);
or OR3 (N6431, N6398, N187, N825);
or OR2 (N6432, N6420, N1573);
not NOT1 (N6433, N6414);
nand NAND4 (N6434, N6415, N3121, N425, N3111);
buf BUF1 (N6435, N6433);
or OR4 (N6436, N6434, N4040, N4749, N4791);
buf BUF1 (N6437, N6419);
buf BUF1 (N6438, N6436);
and AND4 (N6439, N6432, N3518, N2604, N2961);
xor XOR2 (N6440, N6422, N3960);
or OR4 (N6441, N6438, N5918, N5063, N3686);
and AND3 (N6442, N6428, N6072, N6050);
buf BUF1 (N6443, N6430);
buf BUF1 (N6444, N6439);
nand NAND4 (N6445, N6441, N51, N705, N2233);
buf BUF1 (N6446, N6427);
nor NOR3 (N6447, N6437, N646, N129);
buf BUF1 (N6448, N6426);
or OR4 (N6449, N6444, N4064, N6408, N5200);
and AND2 (N6450, N6440, N4280);
and AND4 (N6451, N6442, N3424, N621, N4176);
and AND2 (N6452, N6445, N3232);
nor NOR4 (N6453, N6448, N4523, N5485, N5393);
not NOT1 (N6454, N6431);
xor XOR2 (N6455, N6454, N3500);
or OR2 (N6456, N6450, N5045);
nand NAND3 (N6457, N6455, N6429, N4794);
or OR4 (N6458, N6449, N4359, N4230, N4512);
nor NOR4 (N6459, N6451, N2061, N3356, N3391);
and AND2 (N6460, N6447, N3308);
buf BUF1 (N6461, N6457);
nor NOR4 (N6462, N6443, N2644, N2766, N5822);
not NOT1 (N6463, N6461);
nor NOR4 (N6464, N6458, N3081, N5810, N2735);
nor NOR2 (N6465, N6463, N3315);
and AND3 (N6466, N6459, N1599, N5861);
or OR2 (N6467, N6456, N4977);
not NOT1 (N6468, N6446);
buf BUF1 (N6469, N6464);
xor XOR2 (N6470, N6468, N4906);
or OR4 (N6471, N6453, N166, N4000, N599);
not NOT1 (N6472, N6469);
xor XOR2 (N6473, N6466, N5552);
or OR4 (N6474, N6460, N2875, N6083, N4318);
xor XOR2 (N6475, N6465, N5293);
and AND2 (N6476, N6467, N3307);
and AND3 (N6477, N6474, N3345, N3297);
nor NOR2 (N6478, N6462, N1053);
not NOT1 (N6479, N6470);
nand NAND3 (N6480, N6452, N1649, N3830);
not NOT1 (N6481, N6477);
not NOT1 (N6482, N6478);
and AND3 (N6483, N6475, N3548, N2847);
and AND4 (N6484, N6435, N5628, N5335, N432);
or OR2 (N6485, N6481, N4067);
and AND2 (N6486, N6483, N1560);
nand NAND2 (N6487, N6472, N5706);
not NOT1 (N6488, N6486);
not NOT1 (N6489, N6485);
nor NOR2 (N6490, N6480, N5607);
and AND4 (N6491, N6482, N4347, N1459, N3754);
and AND2 (N6492, N6476, N5105);
nand NAND2 (N6493, N6473, N4217);
not NOT1 (N6494, N6479);
or OR3 (N6495, N6484, N6437, N3392);
nor NOR2 (N6496, N6493, N1027);
not NOT1 (N6497, N6492);
and AND2 (N6498, N6495, N3978);
or OR2 (N6499, N6491, N4872);
not NOT1 (N6500, N6489);
buf BUF1 (N6501, N6490);
not NOT1 (N6502, N6500);
and AND2 (N6503, N6471, N4892);
or OR2 (N6504, N6498, N1446);
and AND4 (N6505, N6494, N965, N4013, N1591);
nor NOR3 (N6506, N6488, N4460, N384);
and AND2 (N6507, N6502, N6304);
xor XOR2 (N6508, N6503, N498);
xor XOR2 (N6509, N6508, N4505);
or OR4 (N6510, N6487, N3573, N3639, N2773);
or OR2 (N6511, N6497, N3913);
and AND4 (N6512, N6505, N2978, N568, N2001);
nor NOR2 (N6513, N6510, N3879);
not NOT1 (N6514, N6501);
nand NAND2 (N6515, N6514, N1610);
and AND3 (N6516, N6509, N6353, N422);
nand NAND2 (N6517, N6499, N4478);
nand NAND4 (N6518, N6511, N989, N2754, N456);
not NOT1 (N6519, N6504);
xor XOR2 (N6520, N6507, N5004);
not NOT1 (N6521, N6517);
or OR4 (N6522, N6513, N452, N2819, N5418);
nor NOR2 (N6523, N6496, N6293);
nor NOR2 (N6524, N6515, N6199);
nor NOR2 (N6525, N6516, N5772);
and AND2 (N6526, N6512, N4792);
nor NOR4 (N6527, N6524, N1257, N4093, N3397);
and AND4 (N6528, N6527, N3658, N7, N2842);
nor NOR4 (N6529, N6525, N5196, N5046, N653);
not NOT1 (N6530, N6522);
and AND3 (N6531, N6518, N4490, N6352);
xor XOR2 (N6532, N6506, N1193);
nand NAND4 (N6533, N6528, N6013, N5465, N3978);
nor NOR2 (N6534, N6526, N3117);
nor NOR4 (N6535, N6520, N1049, N1902, N5690);
not NOT1 (N6536, N6535);
and AND4 (N6537, N6523, N2583, N1013, N4715);
nor NOR4 (N6538, N6536, N5314, N1957, N6216);
or OR2 (N6539, N6529, N3500);
nand NAND3 (N6540, N6531, N5435, N1427);
buf BUF1 (N6541, N6533);
buf BUF1 (N6542, N6519);
and AND2 (N6543, N6540, N3959);
and AND3 (N6544, N6539, N1651, N3658);
or OR2 (N6545, N6541, N2271);
or OR4 (N6546, N6534, N5032, N2287, N2731);
and AND3 (N6547, N6521, N1187, N362);
nor NOR4 (N6548, N6546, N5971, N2390, N2157);
not NOT1 (N6549, N6542);
xor XOR2 (N6550, N6544, N415);
xor XOR2 (N6551, N6550, N667);
buf BUF1 (N6552, N6543);
and AND2 (N6553, N6549, N2959);
xor XOR2 (N6554, N6532, N2111);
xor XOR2 (N6555, N6538, N3287);
not NOT1 (N6556, N6547);
buf BUF1 (N6557, N6530);
and AND4 (N6558, N6553, N1744, N2540, N4312);
and AND4 (N6559, N6556, N3854, N5686, N5545);
and AND2 (N6560, N6552, N2713);
nand NAND4 (N6561, N6537, N6317, N3946, N1371);
buf BUF1 (N6562, N6558);
and AND2 (N6563, N6562, N2962);
buf BUF1 (N6564, N6560);
nand NAND2 (N6565, N6545, N5877);
nor NOR2 (N6566, N6559, N5674);
or OR3 (N6567, N6555, N6343, N2197);
xor XOR2 (N6568, N6551, N6006);
buf BUF1 (N6569, N6565);
not NOT1 (N6570, N6569);
buf BUF1 (N6571, N6557);
xor XOR2 (N6572, N6568, N3878);
xor XOR2 (N6573, N6567, N4216);
nand NAND4 (N6574, N6554, N6232, N3027, N6338);
buf BUF1 (N6575, N6548);
and AND3 (N6576, N6573, N1507, N3698);
and AND3 (N6577, N6570, N1907, N5760);
and AND3 (N6578, N6566, N611, N3995);
or OR2 (N6579, N6564, N4146);
buf BUF1 (N6580, N6572);
and AND4 (N6581, N6577, N2816, N566, N1414);
or OR4 (N6582, N6563, N1454, N2121, N5922);
and AND2 (N6583, N6580, N2176);
and AND2 (N6584, N6579, N2895);
and AND2 (N6585, N6584, N557);
not NOT1 (N6586, N6581);
nor NOR2 (N6587, N6578, N5648);
buf BUF1 (N6588, N6582);
xor XOR2 (N6589, N6586, N4666);
not NOT1 (N6590, N6583);
nor NOR4 (N6591, N6574, N3237, N3777, N3079);
not NOT1 (N6592, N6585);
and AND4 (N6593, N6592, N4153, N840, N4262);
nor NOR2 (N6594, N6575, N5852);
or OR3 (N6595, N6571, N2959, N1940);
or OR4 (N6596, N6591, N221, N3318, N4896);
buf BUF1 (N6597, N6587);
nand NAND2 (N6598, N6595, N6334);
buf BUF1 (N6599, N6576);
nor NOR4 (N6600, N6590, N666, N5890, N19);
buf BUF1 (N6601, N6597);
buf BUF1 (N6602, N6594);
buf BUF1 (N6603, N6601);
nand NAND4 (N6604, N6588, N5289, N4646, N365);
and AND2 (N6605, N6602, N212);
nor NOR3 (N6606, N6603, N2721, N1727);
and AND2 (N6607, N6598, N3652);
xor XOR2 (N6608, N6596, N4414);
not NOT1 (N6609, N6599);
buf BUF1 (N6610, N6607);
nor NOR2 (N6611, N6608, N5236);
nand NAND4 (N6612, N6604, N6102, N1194, N21);
or OR2 (N6613, N6589, N3170);
nand NAND2 (N6614, N6612, N2376);
or OR3 (N6615, N6609, N1487, N1372);
buf BUF1 (N6616, N6615);
not NOT1 (N6617, N6561);
xor XOR2 (N6618, N6605, N840);
nand NAND2 (N6619, N6610, N4643);
buf BUF1 (N6620, N6600);
not NOT1 (N6621, N6620);
and AND4 (N6622, N6613, N5480, N3679, N2457);
and AND4 (N6623, N6619, N2162, N1086, N4196);
nor NOR4 (N6624, N6614, N2550, N6550, N4973);
xor XOR2 (N6625, N6617, N1858);
xor XOR2 (N6626, N6593, N5258);
xor XOR2 (N6627, N6621, N2923);
not NOT1 (N6628, N6611);
nand NAND4 (N6629, N6623, N2630, N2032, N6530);
xor XOR2 (N6630, N6628, N5178);
nand NAND4 (N6631, N6606, N4134, N5755, N4577);
buf BUF1 (N6632, N6618);
not NOT1 (N6633, N6622);
buf BUF1 (N6634, N6624);
nor NOR2 (N6635, N6625, N4326);
xor XOR2 (N6636, N6630, N5422);
nand NAND2 (N6637, N6626, N2479);
and AND2 (N6638, N6635, N2962);
nand NAND4 (N6639, N6629, N5385, N631, N2572);
xor XOR2 (N6640, N6638, N315);
nand NAND4 (N6641, N6637, N5831, N1744, N1560);
nor NOR2 (N6642, N6639, N707);
xor XOR2 (N6643, N6636, N6111);
nor NOR4 (N6644, N6642, N4389, N4320, N1821);
or OR4 (N6645, N6627, N2943, N2159, N5014);
and AND3 (N6646, N6631, N1951, N2961);
buf BUF1 (N6647, N6633);
nand NAND2 (N6648, N6647, N2530);
or OR4 (N6649, N6632, N3477, N319, N2280);
not NOT1 (N6650, N6640);
xor XOR2 (N6651, N6649, N1967);
nand NAND2 (N6652, N6634, N1497);
xor XOR2 (N6653, N6651, N2227);
not NOT1 (N6654, N6646);
nor NOR4 (N6655, N6616, N5975, N3841, N2507);
nand NAND3 (N6656, N6650, N320, N3334);
xor XOR2 (N6657, N6655, N904);
buf BUF1 (N6658, N6645);
or OR2 (N6659, N6657, N1674);
or OR4 (N6660, N6653, N2553, N10, N3369);
nor NOR4 (N6661, N6659, N3553, N505, N5468);
buf BUF1 (N6662, N6658);
nand NAND2 (N6663, N6643, N5049);
nor NOR2 (N6664, N6644, N6387);
and AND3 (N6665, N6662, N1701, N1873);
nor NOR4 (N6666, N6665, N2169, N2687, N5681);
nand NAND3 (N6667, N6660, N3909, N918);
or OR2 (N6668, N6666, N1664);
buf BUF1 (N6669, N6656);
not NOT1 (N6670, N6641);
buf BUF1 (N6671, N6663);
and AND2 (N6672, N6654, N1973);
and AND4 (N6673, N6667, N6139, N2759, N2319);
nand NAND3 (N6674, N6670, N235, N5036);
or OR2 (N6675, N6671, N677);
nor NOR3 (N6676, N6675, N1463, N1429);
or OR4 (N6677, N6664, N1303, N2600, N6332);
and AND4 (N6678, N6677, N1386, N3653, N398);
or OR4 (N6679, N6669, N59, N6241, N2270);
or OR3 (N6680, N6668, N4489, N3114);
nand NAND4 (N6681, N6661, N3346, N2941, N2880);
nand NAND3 (N6682, N6652, N6338, N4614);
or OR3 (N6683, N6682, N3999, N6045);
and AND2 (N6684, N6680, N3742);
buf BUF1 (N6685, N6673);
xor XOR2 (N6686, N6684, N6376);
xor XOR2 (N6687, N6686, N4113);
buf BUF1 (N6688, N6678);
xor XOR2 (N6689, N6687, N1124);
buf BUF1 (N6690, N6672);
or OR3 (N6691, N6685, N4782, N6124);
buf BUF1 (N6692, N6688);
and AND3 (N6693, N6691, N137, N4819);
or OR3 (N6694, N6690, N1185, N4325);
or OR3 (N6695, N6683, N3068, N4166);
not NOT1 (N6696, N6693);
buf BUF1 (N6697, N6692);
or OR2 (N6698, N6681, N2708);
and AND4 (N6699, N6648, N4922, N1639, N4815);
and AND3 (N6700, N6679, N41, N5955);
xor XOR2 (N6701, N6689, N1608);
or OR3 (N6702, N6701, N6685, N5662);
xor XOR2 (N6703, N6674, N157);
and AND4 (N6704, N6698, N3613, N1403, N5523);
xor XOR2 (N6705, N6699, N3240);
not NOT1 (N6706, N6704);
nor NOR3 (N6707, N6694, N3623, N5478);
nand NAND4 (N6708, N6695, N6164, N2929, N4161);
not NOT1 (N6709, N6697);
and AND3 (N6710, N6702, N4772, N2721);
buf BUF1 (N6711, N6696);
xor XOR2 (N6712, N6676, N5618);
or OR2 (N6713, N6707, N3342);
and AND3 (N6714, N6712, N6453, N5335);
nand NAND4 (N6715, N6703, N4793, N3372, N4943);
nand NAND3 (N6716, N6708, N1704, N5928);
nor NOR3 (N6717, N6713, N6411, N4648);
not NOT1 (N6718, N6709);
buf BUF1 (N6719, N6718);
and AND2 (N6720, N6705, N1827);
and AND2 (N6721, N6719, N5331);
nor NOR4 (N6722, N6714, N4204, N5238, N1597);
not NOT1 (N6723, N6716);
xor XOR2 (N6724, N6711, N1560);
not NOT1 (N6725, N6717);
and AND3 (N6726, N6722, N2033, N3330);
and AND3 (N6727, N6715, N4816, N2881);
nor NOR3 (N6728, N6726, N5313, N6708);
or OR2 (N6729, N6720, N5598);
xor XOR2 (N6730, N6710, N3990);
and AND2 (N6731, N6700, N3430);
and AND4 (N6732, N6729, N2370, N4769, N1649);
and AND4 (N6733, N6725, N5910, N1708, N236);
nand NAND4 (N6734, N6721, N2582, N1281, N891);
buf BUF1 (N6735, N6728);
xor XOR2 (N6736, N6724, N266);
not NOT1 (N6737, N6706);
and AND3 (N6738, N6731, N6095, N5923);
and AND3 (N6739, N6737, N5739, N1376);
and AND4 (N6740, N6732, N3887, N6410, N578);
nand NAND3 (N6741, N6723, N4425, N4101);
and AND3 (N6742, N6733, N6611, N2793);
or OR2 (N6743, N6740, N4416);
buf BUF1 (N6744, N6742);
nand NAND4 (N6745, N6744, N4885, N4009, N6313);
or OR2 (N6746, N6738, N325);
or OR2 (N6747, N6735, N6234);
not NOT1 (N6748, N6741);
not NOT1 (N6749, N6734);
nand NAND2 (N6750, N6747, N2421);
not NOT1 (N6751, N6746);
nor NOR4 (N6752, N6751, N645, N2870, N4419);
not NOT1 (N6753, N6752);
or OR2 (N6754, N6750, N6717);
buf BUF1 (N6755, N6749);
nand NAND2 (N6756, N6753, N2824);
buf BUF1 (N6757, N6755);
nand NAND4 (N6758, N6743, N1480, N755, N5524);
buf BUF1 (N6759, N6757);
or OR4 (N6760, N6730, N4913, N720, N708);
not NOT1 (N6761, N6760);
or OR2 (N6762, N6736, N6323);
nor NOR3 (N6763, N6759, N2750, N2069);
not NOT1 (N6764, N6754);
or OR2 (N6765, N6748, N2452);
nand NAND4 (N6766, N6756, N3907, N1029, N2805);
nor NOR2 (N6767, N6763, N6648);
not NOT1 (N6768, N6727);
nor NOR4 (N6769, N6764, N278, N3344, N6111);
or OR4 (N6770, N6768, N3709, N4843, N5383);
and AND4 (N6771, N6739, N5994, N1198, N5276);
and AND3 (N6772, N6766, N6007, N5108);
not NOT1 (N6773, N6745);
xor XOR2 (N6774, N6762, N6655);
xor XOR2 (N6775, N6761, N6229);
not NOT1 (N6776, N6771);
buf BUF1 (N6777, N6772);
nand NAND2 (N6778, N6758, N1044);
buf BUF1 (N6779, N6776);
and AND3 (N6780, N6765, N1999, N5722);
not NOT1 (N6781, N6767);
xor XOR2 (N6782, N6781, N463);
xor XOR2 (N6783, N6782, N106);
and AND3 (N6784, N6779, N4050, N5460);
buf BUF1 (N6785, N6774);
and AND4 (N6786, N6780, N2244, N1464, N2675);
not NOT1 (N6787, N6785);
buf BUF1 (N6788, N6784);
xor XOR2 (N6789, N6787, N2545);
or OR2 (N6790, N6769, N5993);
nor NOR3 (N6791, N6786, N3098, N4684);
xor XOR2 (N6792, N6775, N2801);
or OR4 (N6793, N6778, N6430, N6059, N5232);
xor XOR2 (N6794, N6790, N5529);
xor XOR2 (N6795, N6794, N6504);
xor XOR2 (N6796, N6795, N627);
buf BUF1 (N6797, N6796);
buf BUF1 (N6798, N6792);
nand NAND4 (N6799, N6777, N280, N2833, N1229);
and AND2 (N6800, N6793, N3099);
and AND3 (N6801, N6788, N1840, N246);
xor XOR2 (N6802, N6770, N1791);
xor XOR2 (N6803, N6783, N2173);
xor XOR2 (N6804, N6797, N700);
buf BUF1 (N6805, N6800);
buf BUF1 (N6806, N6801);
nand NAND4 (N6807, N6799, N1777, N199, N1849);
xor XOR2 (N6808, N6804, N6337);
or OR3 (N6809, N6807, N6707, N4023);
and AND2 (N6810, N6806, N4172);
nor NOR2 (N6811, N6809, N4296);
buf BUF1 (N6812, N6808);
and AND4 (N6813, N6805, N4014, N618, N125);
buf BUF1 (N6814, N6811);
xor XOR2 (N6815, N6803, N110);
nor NOR4 (N6816, N6810, N4565, N1524, N3897);
nand NAND2 (N6817, N6812, N5577);
and AND4 (N6818, N6815, N4370, N6159, N6141);
not NOT1 (N6819, N6818);
nor NOR2 (N6820, N6789, N3353);
or OR4 (N6821, N6819, N6000, N4670, N5523);
xor XOR2 (N6822, N6773, N644);
and AND4 (N6823, N6798, N6159, N5641, N6066);
buf BUF1 (N6824, N6821);
buf BUF1 (N6825, N6817);
nand NAND2 (N6826, N6802, N888);
nand NAND4 (N6827, N6813, N5195, N613, N1612);
nor NOR4 (N6828, N6823, N1470, N5624, N978);
xor XOR2 (N6829, N6827, N5052);
and AND3 (N6830, N6824, N1676, N6116);
not NOT1 (N6831, N6828);
not NOT1 (N6832, N6829);
nand NAND2 (N6833, N6825, N2964);
not NOT1 (N6834, N6830);
or OR2 (N6835, N6822, N3031);
buf BUF1 (N6836, N6833);
buf BUF1 (N6837, N6834);
not NOT1 (N6838, N6831);
nor NOR3 (N6839, N6814, N3412, N1321);
or OR4 (N6840, N6832, N637, N3007, N3592);
or OR2 (N6841, N6839, N1823);
or OR3 (N6842, N6841, N6551, N4968);
xor XOR2 (N6843, N6816, N3798);
or OR3 (N6844, N6838, N1593, N2977);
not NOT1 (N6845, N6840);
buf BUF1 (N6846, N6837);
and AND4 (N6847, N6835, N6836, N3339, N738);
or OR3 (N6848, N431, N252, N5101);
buf BUF1 (N6849, N6845);
nor NOR3 (N6850, N6843, N6640, N5387);
xor XOR2 (N6851, N6846, N2712);
nor NOR4 (N6852, N6842, N6553, N4062, N1682);
or OR2 (N6853, N6820, N4112);
or OR4 (N6854, N6844, N5348, N2283, N1120);
xor XOR2 (N6855, N6850, N2391);
nand NAND4 (N6856, N6852, N4801, N5153, N5492);
or OR4 (N6857, N6856, N3779, N3308, N5071);
xor XOR2 (N6858, N6847, N5963);
and AND4 (N6859, N6858, N3821, N3198, N4980);
not NOT1 (N6860, N6855);
nand NAND4 (N6861, N6849, N5248, N5896, N6468);
nor NOR3 (N6862, N6861, N2607, N5438);
buf BUF1 (N6863, N6851);
not NOT1 (N6864, N6848);
buf BUF1 (N6865, N6826);
buf BUF1 (N6866, N6791);
nor NOR4 (N6867, N6863, N1473, N1602, N3710);
not NOT1 (N6868, N6862);
nor NOR2 (N6869, N6857, N5994);
nor NOR3 (N6870, N6859, N2047, N3828);
nand NAND4 (N6871, N6854, N2999, N4302, N5292);
nor NOR4 (N6872, N6869, N410, N2053, N1532);
xor XOR2 (N6873, N6871, N83);
nor NOR4 (N6874, N6860, N4020, N2695, N4356);
or OR4 (N6875, N6872, N3706, N4151, N2334);
nor NOR3 (N6876, N6867, N3812, N6206);
nor NOR4 (N6877, N6873, N4038, N64, N3245);
and AND4 (N6878, N6874, N976, N2112, N4121);
nand NAND2 (N6879, N6864, N3321);
or OR4 (N6880, N6876, N1567, N4743, N706);
nor NOR4 (N6881, N6878, N3720, N2889, N2921);
xor XOR2 (N6882, N6870, N4368);
xor XOR2 (N6883, N6882, N911);
buf BUF1 (N6884, N6879);
not NOT1 (N6885, N6881);
and AND3 (N6886, N6880, N2047, N144);
not NOT1 (N6887, N6868);
nor NOR2 (N6888, N6884, N2116);
buf BUF1 (N6889, N6888);
and AND2 (N6890, N6883, N3886);
xor XOR2 (N6891, N6853, N1265);
nor NOR4 (N6892, N6889, N1546, N3439, N3463);
nor NOR3 (N6893, N6892, N3483, N1177);
nor NOR4 (N6894, N6885, N6095, N6287, N390);
buf BUF1 (N6895, N6894);
nand NAND2 (N6896, N6886, N5002);
not NOT1 (N6897, N6865);
and AND3 (N6898, N6877, N347, N465);
xor XOR2 (N6899, N6875, N1784);
or OR4 (N6900, N6890, N3266, N2134, N5032);
nor NOR4 (N6901, N6866, N65, N4528, N19);
or OR3 (N6902, N6900, N4650, N5567);
not NOT1 (N6903, N6898);
and AND3 (N6904, N6899, N5988, N4061);
buf BUF1 (N6905, N6893);
nand NAND3 (N6906, N6903, N2556, N2013);
or OR3 (N6907, N6896, N3169, N5335);
and AND4 (N6908, N6901, N5423, N6463, N4272);
buf BUF1 (N6909, N6887);
xor XOR2 (N6910, N6891, N3222);
and AND3 (N6911, N6897, N313, N5956);
nand NAND3 (N6912, N6910, N2640, N2793);
xor XOR2 (N6913, N6902, N1029);
buf BUF1 (N6914, N6913);
buf BUF1 (N6915, N6911);
buf BUF1 (N6916, N6905);
not NOT1 (N6917, N6912);
nor NOR2 (N6918, N6916, N3657);
buf BUF1 (N6919, N6908);
or OR2 (N6920, N6918, N2702);
buf BUF1 (N6921, N6917);
or OR2 (N6922, N6909, N6759);
or OR4 (N6923, N6904, N5589, N2594, N3668);
nand NAND4 (N6924, N6915, N6403, N2986, N5151);
nand NAND2 (N6925, N6924, N2133);
or OR4 (N6926, N6919, N266, N1149, N6143);
buf BUF1 (N6927, N6920);
or OR4 (N6928, N6921, N971, N4114, N2517);
or OR3 (N6929, N6928, N4692, N1153);
and AND4 (N6930, N6922, N4258, N5896, N192);
not NOT1 (N6931, N6930);
nor NOR2 (N6932, N6931, N2574);
and AND4 (N6933, N6932, N5298, N1911, N4282);
nand NAND4 (N6934, N6926, N5166, N4466, N4811);
nand NAND3 (N6935, N6934, N1135, N3118);
nor NOR2 (N6936, N6914, N6340);
buf BUF1 (N6937, N6925);
xor XOR2 (N6938, N6935, N2066);
nor NOR2 (N6939, N6895, N4905);
or OR4 (N6940, N6939, N2851, N5528, N5512);
not NOT1 (N6941, N6906);
and AND2 (N6942, N6923, N5970);
or OR3 (N6943, N6941, N265, N2048);
nor NOR2 (N6944, N6907, N630);
and AND3 (N6945, N6943, N300, N3943);
and AND3 (N6946, N6937, N2883, N2328);
not NOT1 (N6947, N6933);
xor XOR2 (N6948, N6942, N832);
nand NAND4 (N6949, N6929, N4824, N4911, N4780);
not NOT1 (N6950, N6948);
nand NAND3 (N6951, N6945, N4425, N4320);
xor XOR2 (N6952, N6940, N219);
xor XOR2 (N6953, N6927, N3078);
and AND3 (N6954, N6952, N2325, N3750);
nand NAND4 (N6955, N6936, N3404, N5657, N6209);
xor XOR2 (N6956, N6954, N1661);
xor XOR2 (N6957, N6944, N3136);
and AND2 (N6958, N6951, N6426);
xor XOR2 (N6959, N6946, N1508);
or OR3 (N6960, N6956, N4440, N3437);
and AND2 (N6961, N6950, N623);
xor XOR2 (N6962, N6949, N4655);
xor XOR2 (N6963, N6961, N5523);
nand NAND3 (N6964, N6962, N5233, N191);
xor XOR2 (N6965, N6963, N4924);
or OR3 (N6966, N6953, N2038, N6777);
xor XOR2 (N6967, N6947, N4653);
nor NOR3 (N6968, N6955, N1369, N366);
or OR3 (N6969, N6968, N1754, N1929);
nor NOR3 (N6970, N6938, N5515, N1610);
buf BUF1 (N6971, N6960);
nand NAND3 (N6972, N6971, N4748, N4641);
not NOT1 (N6973, N6959);
buf BUF1 (N6974, N6967);
nor NOR2 (N6975, N6969, N6956);
nand NAND3 (N6976, N6965, N4428, N778);
buf BUF1 (N6977, N6974);
nand NAND3 (N6978, N6977, N1653, N1318);
or OR2 (N6979, N6966, N3822);
nor NOR2 (N6980, N6958, N2358);
buf BUF1 (N6981, N6979);
not NOT1 (N6982, N6980);
buf BUF1 (N6983, N6957);
or OR2 (N6984, N6970, N3106);
or OR2 (N6985, N6972, N432);
buf BUF1 (N6986, N6981);
nand NAND2 (N6987, N6986, N1696);
and AND2 (N6988, N6978, N422);
not NOT1 (N6989, N6984);
not NOT1 (N6990, N6985);
xor XOR2 (N6991, N6964, N5374);
nor NOR3 (N6992, N6991, N2638, N4827);
buf BUF1 (N6993, N6988);
buf BUF1 (N6994, N6982);
xor XOR2 (N6995, N6975, N6946);
nand NAND4 (N6996, N6973, N6730, N567, N6641);
or OR4 (N6997, N6995, N4230, N2709, N1470);
buf BUF1 (N6998, N6990);
nor NOR4 (N6999, N6996, N6347, N6297, N1265);
nand NAND4 (N7000, N6987, N1368, N3333, N2957);
xor XOR2 (N7001, N6998, N5344);
or OR3 (N7002, N6983, N189, N164);
and AND3 (N7003, N6993, N673, N6578);
and AND4 (N7004, N6994, N6838, N1367, N1241);
nor NOR3 (N7005, N7004, N318, N3386);
xor XOR2 (N7006, N7002, N1137);
and AND4 (N7007, N7005, N4791, N4264, N5776);
or OR4 (N7008, N7001, N630, N1649, N1338);
xor XOR2 (N7009, N7006, N807);
nand NAND3 (N7010, N6976, N4954, N3765);
buf BUF1 (N7011, N7010);
not NOT1 (N7012, N6989);
xor XOR2 (N7013, N7008, N6259);
xor XOR2 (N7014, N7011, N1905);
nand NAND2 (N7015, N7012, N5237);
buf BUF1 (N7016, N7003);
xor XOR2 (N7017, N7000, N5473);
not NOT1 (N7018, N6999);
and AND3 (N7019, N7014, N437, N4205);
buf BUF1 (N7020, N6997);
nand NAND3 (N7021, N6992, N2163, N3921);
nor NOR4 (N7022, N7017, N4785, N1540, N5715);
nor NOR2 (N7023, N7015, N1424);
or OR2 (N7024, N7016, N3050);
xor XOR2 (N7025, N7007, N5441);
and AND4 (N7026, N7023, N5509, N2500, N4650);
or OR4 (N7027, N7009, N6117, N3356, N6973);
nor NOR3 (N7028, N7022, N5284, N3716);
and AND4 (N7029, N7020, N6495, N1840, N6547);
buf BUF1 (N7030, N7013);
nand NAND3 (N7031, N7026, N6407, N4384);
nor NOR2 (N7032, N7019, N1889);
buf BUF1 (N7033, N7029);
nor NOR4 (N7034, N7021, N1151, N6837, N4514);
nor NOR4 (N7035, N7024, N4690, N4746, N4676);
nor NOR4 (N7036, N7018, N1587, N3285, N3676);
buf BUF1 (N7037, N7027);
not NOT1 (N7038, N7032);
buf BUF1 (N7039, N7031);
not NOT1 (N7040, N7025);
xor XOR2 (N7041, N7034, N4467);
and AND4 (N7042, N7033, N6337, N2530, N1911);
not NOT1 (N7043, N7039);
nor NOR2 (N7044, N7043, N964);
or OR3 (N7045, N7042, N2711, N748);
not NOT1 (N7046, N7035);
not NOT1 (N7047, N7044);
and AND3 (N7048, N7040, N1731, N4589);
not NOT1 (N7049, N7047);
and AND2 (N7050, N7049, N1006);
buf BUF1 (N7051, N7046);
xor XOR2 (N7052, N7030, N2714);
buf BUF1 (N7053, N7036);
nor NOR3 (N7054, N7038, N2436, N3780);
and AND4 (N7055, N7053, N4463, N2126, N3286);
nand NAND2 (N7056, N7052, N3087);
xor XOR2 (N7057, N7048, N4059);
or OR4 (N7058, N7057, N5007, N713, N4704);
buf BUF1 (N7059, N7058);
or OR4 (N7060, N7028, N666, N3831, N205);
and AND2 (N7061, N7059, N7045);
nor NOR2 (N7062, N797, N649);
buf BUF1 (N7063, N7056);
nor NOR3 (N7064, N7060, N4433, N873);
or OR4 (N7065, N7061, N4839, N5014, N2886);
nand NAND2 (N7066, N7064, N5347);
not NOT1 (N7067, N7062);
and AND4 (N7068, N7037, N6363, N1638, N5230);
and AND3 (N7069, N7067, N5043, N4268);
nor NOR4 (N7070, N7054, N6037, N4175, N980);
not NOT1 (N7071, N7066);
nand NAND3 (N7072, N7055, N3924, N5625);
or OR3 (N7073, N7041, N1733, N534);
buf BUF1 (N7074, N7050);
buf BUF1 (N7075, N7074);
or OR3 (N7076, N7072, N268, N5553);
nand NAND3 (N7077, N7075, N3105, N6304);
or OR3 (N7078, N7073, N4993, N6958);
buf BUF1 (N7079, N7076);
nor NOR4 (N7080, N7069, N6165, N5416, N3598);
xor XOR2 (N7081, N7070, N2497);
not NOT1 (N7082, N7081);
nor NOR4 (N7083, N7051, N1010, N4344, N2112);
buf BUF1 (N7084, N7068);
nand NAND4 (N7085, N7077, N2467, N5133, N1395);
or OR2 (N7086, N7071, N5827);
and AND4 (N7087, N7086, N6071, N457, N4783);
nand NAND3 (N7088, N7078, N1252, N2016);
and AND2 (N7089, N7084, N5046);
or OR3 (N7090, N7085, N1373, N3419);
nand NAND2 (N7091, N7079, N3383);
not NOT1 (N7092, N7080);
nor NOR3 (N7093, N7065, N390, N6668);
and AND4 (N7094, N7089, N5705, N127, N5086);
nor NOR3 (N7095, N7091, N3107, N5190);
xor XOR2 (N7096, N7095, N5948);
xor XOR2 (N7097, N7088, N6676);
or OR4 (N7098, N7096, N4363, N6493, N2404);
xor XOR2 (N7099, N7092, N1502);
and AND3 (N7100, N7098, N2699, N6867);
xor XOR2 (N7101, N7100, N3399);
buf BUF1 (N7102, N7082);
or OR2 (N7103, N7102, N3967);
or OR2 (N7104, N7099, N52);
buf BUF1 (N7105, N7104);
nor NOR3 (N7106, N7063, N5817, N1635);
nor NOR4 (N7107, N7083, N5514, N743, N4547);
buf BUF1 (N7108, N7107);
xor XOR2 (N7109, N7105, N3812);
or OR4 (N7110, N7108, N3414, N4708, N6701);
xor XOR2 (N7111, N7109, N895);
buf BUF1 (N7112, N7101);
and AND4 (N7113, N7097, N1701, N1529, N2434);
not NOT1 (N7114, N7087);
nor NOR4 (N7115, N7106, N3924, N3330, N2864);
nand NAND3 (N7116, N7093, N165, N6541);
nand NAND2 (N7117, N7116, N2808);
buf BUF1 (N7118, N7111);
buf BUF1 (N7119, N7103);
not NOT1 (N7120, N7110);
or OR3 (N7121, N7120, N2466, N4130);
not NOT1 (N7122, N7118);
or OR4 (N7123, N7094, N1071, N6733, N6215);
or OR3 (N7124, N7113, N3898, N4763);
not NOT1 (N7125, N7090);
and AND4 (N7126, N7122, N1559, N3741, N531);
buf BUF1 (N7127, N7117);
xor XOR2 (N7128, N7127, N352);
xor XOR2 (N7129, N7114, N5353);
not NOT1 (N7130, N7128);
or OR3 (N7131, N7130, N4205, N3519);
and AND3 (N7132, N7129, N4999, N86);
and AND2 (N7133, N7123, N114);
nand NAND2 (N7134, N7115, N2849);
not NOT1 (N7135, N7131);
not NOT1 (N7136, N7126);
not NOT1 (N7137, N7121);
not NOT1 (N7138, N7134);
buf BUF1 (N7139, N7112);
or OR2 (N7140, N7132, N4372);
not NOT1 (N7141, N7119);
or OR2 (N7142, N7136, N4463);
and AND3 (N7143, N7133, N4905, N2471);
xor XOR2 (N7144, N7140, N6385);
nor NOR4 (N7145, N7142, N4872, N6543, N5641);
buf BUF1 (N7146, N7145);
xor XOR2 (N7147, N7141, N6055);
nand NAND4 (N7148, N7143, N3749, N3041, N1670);
nor NOR4 (N7149, N7144, N2180, N7132, N6230);
buf BUF1 (N7150, N7124);
nor NOR4 (N7151, N7147, N4325, N6844, N4544);
not NOT1 (N7152, N7148);
or OR2 (N7153, N7150, N3723);
nand NAND3 (N7154, N7153, N6339, N5795);
or OR2 (N7155, N7149, N5412);
nor NOR4 (N7156, N7155, N5669, N6030, N1419);
nor NOR2 (N7157, N7156, N6200);
nor NOR4 (N7158, N7138, N3028, N266, N3385);
nor NOR3 (N7159, N7137, N3725, N7042);
not NOT1 (N7160, N7146);
nor NOR4 (N7161, N7157, N222, N5260, N1649);
xor XOR2 (N7162, N7158, N1527);
not NOT1 (N7163, N7151);
nor NOR2 (N7164, N7162, N1781);
and AND2 (N7165, N7163, N3573);
nor NOR2 (N7166, N7165, N4257);
and AND3 (N7167, N7152, N6801, N3125);
nor NOR2 (N7168, N7135, N278);
nand NAND4 (N7169, N7139, N4431, N6374, N6252);
and AND3 (N7170, N7167, N1830, N184);
nor NOR2 (N7171, N7161, N62);
not NOT1 (N7172, N7166);
xor XOR2 (N7173, N7169, N4401);
not NOT1 (N7174, N7154);
buf BUF1 (N7175, N7125);
xor XOR2 (N7176, N7173, N2673);
and AND2 (N7177, N7172, N4464);
buf BUF1 (N7178, N7164);
nor NOR4 (N7179, N7159, N2840, N4683, N2686);
nor NOR3 (N7180, N7168, N4810, N5299);
nand NAND3 (N7181, N7171, N5956, N2959);
buf BUF1 (N7182, N7170);
or OR3 (N7183, N7176, N6111, N3367);
xor XOR2 (N7184, N7160, N3454);
not NOT1 (N7185, N7184);
not NOT1 (N7186, N7179);
not NOT1 (N7187, N7181);
nor NOR2 (N7188, N7174, N5241);
nor NOR4 (N7189, N7182, N1138, N6953, N2972);
not NOT1 (N7190, N7178);
xor XOR2 (N7191, N7180, N1096);
buf BUF1 (N7192, N7188);
xor XOR2 (N7193, N7186, N5590);
buf BUF1 (N7194, N7175);
buf BUF1 (N7195, N7187);
buf BUF1 (N7196, N7189);
or OR2 (N7197, N7196, N5475);
not NOT1 (N7198, N7194);
and AND3 (N7199, N7198, N2770, N6503);
xor XOR2 (N7200, N7185, N502);
or OR3 (N7201, N7200, N3974, N6736);
xor XOR2 (N7202, N7201, N2497);
nand NAND4 (N7203, N7195, N2928, N5730, N1970);
and AND3 (N7204, N7183, N6472, N1039);
xor XOR2 (N7205, N7204, N4948);
not NOT1 (N7206, N7197);
nor NOR2 (N7207, N7202, N4898);
nor NOR4 (N7208, N7203, N6691, N3113, N6904);
xor XOR2 (N7209, N7208, N5184);
or OR4 (N7210, N7192, N6273, N2730, N416);
nor NOR2 (N7211, N7177, N6392);
and AND2 (N7212, N7210, N5610);
and AND3 (N7213, N7199, N3782, N2615);
and AND2 (N7214, N7191, N1525);
xor XOR2 (N7215, N7205, N842);
not NOT1 (N7216, N7209);
nand NAND2 (N7217, N7190, N2145);
nand NAND4 (N7218, N7214, N4576, N6438, N5053);
nand NAND3 (N7219, N7211, N3188, N3514);
nor NOR4 (N7220, N7207, N2438, N1256, N3362);
or OR2 (N7221, N7216, N1456);
nand NAND4 (N7222, N7221, N2428, N7, N2515);
buf BUF1 (N7223, N7217);
not NOT1 (N7224, N7215);
and AND3 (N7225, N7219, N680, N4724);
buf BUF1 (N7226, N7212);
or OR3 (N7227, N7213, N6184, N6822);
nor NOR2 (N7228, N7223, N573);
xor XOR2 (N7229, N7228, N2134);
not NOT1 (N7230, N7193);
nand NAND2 (N7231, N7229, N1423);
nor NOR3 (N7232, N7224, N2426, N5723);
or OR3 (N7233, N7225, N5134, N903);
or OR3 (N7234, N7220, N2829, N3526);
or OR3 (N7235, N7234, N7045, N6408);
xor XOR2 (N7236, N7233, N5941);
not NOT1 (N7237, N7222);
nand NAND4 (N7238, N7218, N792, N2725, N4131);
nor NOR4 (N7239, N7230, N6594, N3505, N4477);
xor XOR2 (N7240, N7232, N5068);
or OR2 (N7241, N7206, N6468);
or OR3 (N7242, N7241, N6553, N2340);
xor XOR2 (N7243, N7240, N403);
nor NOR4 (N7244, N7237, N7075, N2076, N5017);
buf BUF1 (N7245, N7243);
or OR4 (N7246, N7239, N5294, N83, N7075);
nand NAND2 (N7247, N7242, N6990);
xor XOR2 (N7248, N7238, N6918);
nor NOR3 (N7249, N7227, N1863, N910);
not NOT1 (N7250, N7245);
xor XOR2 (N7251, N7249, N2789);
nor NOR2 (N7252, N7247, N3154);
buf BUF1 (N7253, N7236);
nand NAND4 (N7254, N7251, N6478, N4392, N2523);
nand NAND2 (N7255, N7244, N4725);
nand NAND2 (N7256, N7252, N2476);
not NOT1 (N7257, N7256);
nand NAND3 (N7258, N7235, N2120, N3279);
buf BUF1 (N7259, N7231);
and AND4 (N7260, N7253, N1365, N4041, N6165);
or OR4 (N7261, N7260, N5489, N2000, N5132);
not NOT1 (N7262, N7261);
or OR4 (N7263, N7246, N4056, N593, N4474);
or OR2 (N7264, N7263, N5966);
or OR2 (N7265, N7257, N1948);
xor XOR2 (N7266, N7264, N2476);
buf BUF1 (N7267, N7262);
not NOT1 (N7268, N7254);
or OR4 (N7269, N7250, N2132, N2401, N3319);
nand NAND2 (N7270, N7226, N7097);
nand NAND2 (N7271, N7266, N4545);
or OR3 (N7272, N7248, N1261, N533);
not NOT1 (N7273, N7270);
or OR2 (N7274, N7255, N3463);
nand NAND4 (N7275, N7259, N4670, N869, N2007);
or OR2 (N7276, N7275, N728);
xor XOR2 (N7277, N7272, N4014);
xor XOR2 (N7278, N7267, N4170);
or OR2 (N7279, N7269, N5392);
not NOT1 (N7280, N7276);
buf BUF1 (N7281, N7271);
buf BUF1 (N7282, N7268);
xor XOR2 (N7283, N7277, N3957);
nor NOR3 (N7284, N7278, N3760, N404);
nor NOR2 (N7285, N7274, N5504);
buf BUF1 (N7286, N7279);
nand NAND4 (N7287, N7282, N5876, N168, N4156);
xor XOR2 (N7288, N7287, N5443);
or OR3 (N7289, N7281, N3783, N2749);
nand NAND2 (N7290, N7280, N2557);
and AND4 (N7291, N7286, N1015, N3361, N3011);
not NOT1 (N7292, N7285);
buf BUF1 (N7293, N7290);
not NOT1 (N7294, N7273);
nor NOR2 (N7295, N7291, N1463);
not NOT1 (N7296, N7265);
nor NOR4 (N7297, N7292, N5169, N1426, N6135);
or OR2 (N7298, N7295, N1959);
nand NAND3 (N7299, N7258, N27, N839);
not NOT1 (N7300, N7299);
not NOT1 (N7301, N7296);
nor NOR4 (N7302, N7284, N1895, N6834, N744);
and AND3 (N7303, N7283, N4285, N6079);
and AND2 (N7304, N7294, N3950);
not NOT1 (N7305, N7301);
not NOT1 (N7306, N7297);
and AND2 (N7307, N7288, N6652);
nor NOR4 (N7308, N7293, N4719, N515, N210);
or OR3 (N7309, N7300, N5439, N5358);
nand NAND4 (N7310, N7303, N4684, N3385, N3886);
and AND4 (N7311, N7289, N4939, N4106, N1535);
and AND2 (N7312, N7298, N1420);
xor XOR2 (N7313, N7309, N148);
or OR3 (N7314, N7307, N6930, N6408);
buf BUF1 (N7315, N7314);
or OR3 (N7316, N7304, N1207, N4017);
xor XOR2 (N7317, N7308, N4819);
buf BUF1 (N7318, N7302);
nand NAND2 (N7319, N7313, N3953);
nor NOR4 (N7320, N7315, N5071, N6109, N2494);
xor XOR2 (N7321, N7320, N1400);
nor NOR3 (N7322, N7319, N2975, N6736);
buf BUF1 (N7323, N7321);
nor NOR2 (N7324, N7312, N1368);
nor NOR3 (N7325, N7322, N5317, N3393);
nor NOR4 (N7326, N7325, N2637, N5213, N6142);
not NOT1 (N7327, N7324);
or OR4 (N7328, N7305, N1683, N5757, N6775);
or OR3 (N7329, N7310, N7062, N661);
xor XOR2 (N7330, N7327, N1527);
and AND2 (N7331, N7328, N7035);
and AND4 (N7332, N7323, N1654, N1307, N6003);
not NOT1 (N7333, N7330);
nand NAND4 (N7334, N7317, N5861, N5441, N4519);
nand NAND2 (N7335, N7311, N6037);
or OR4 (N7336, N7329, N1406, N3986, N609);
buf BUF1 (N7337, N7318);
nor NOR3 (N7338, N7334, N4166, N449);
xor XOR2 (N7339, N7331, N2527);
nand NAND3 (N7340, N7333, N5866, N1451);
not NOT1 (N7341, N7340);
and AND2 (N7342, N7332, N1964);
or OR4 (N7343, N7336, N6474, N6242, N1956);
buf BUF1 (N7344, N7306);
not NOT1 (N7345, N7342);
xor XOR2 (N7346, N7326, N6411);
or OR2 (N7347, N7343, N6187);
and AND4 (N7348, N7344, N5558, N1558, N2112);
nor NOR3 (N7349, N7345, N1668, N3238);
buf BUF1 (N7350, N7349);
or OR4 (N7351, N7347, N2072, N6692, N1732);
buf BUF1 (N7352, N7346);
buf BUF1 (N7353, N7348);
nor NOR2 (N7354, N7338, N537);
or OR3 (N7355, N7353, N3674, N3266);
buf BUF1 (N7356, N7337);
nor NOR4 (N7357, N7351, N498, N172, N1845);
not NOT1 (N7358, N7352);
or OR3 (N7359, N7356, N2227, N5831);
or OR2 (N7360, N7316, N1088);
or OR2 (N7361, N7357, N7252);
nand NAND2 (N7362, N7358, N2290);
and AND4 (N7363, N7355, N7258, N2569, N1748);
not NOT1 (N7364, N7361);
not NOT1 (N7365, N7364);
not NOT1 (N7366, N7339);
or OR4 (N7367, N7360, N3699, N3921, N295);
buf BUF1 (N7368, N7341);
nor NOR3 (N7369, N7367, N138, N860);
not NOT1 (N7370, N7359);
xor XOR2 (N7371, N7335, N2701);
buf BUF1 (N7372, N7369);
buf BUF1 (N7373, N7350);
nor NOR2 (N7374, N7362, N4347);
and AND2 (N7375, N7372, N1412);
and AND2 (N7376, N7365, N4096);
and AND2 (N7377, N7373, N6249);
or OR2 (N7378, N7371, N6377);
xor XOR2 (N7379, N7370, N693);
nand NAND4 (N7380, N7377, N7142, N6584, N1502);
and AND3 (N7381, N7376, N5187, N2979);
buf BUF1 (N7382, N7374);
and AND4 (N7383, N7379, N6689, N3362, N1543);
or OR2 (N7384, N7366, N6739);
and AND3 (N7385, N7378, N2043, N2628);
xor XOR2 (N7386, N7368, N6001);
nor NOR4 (N7387, N7375, N4448, N2670, N6785);
nand NAND2 (N7388, N7354, N4567);
and AND4 (N7389, N7386, N7043, N4324, N974);
nor NOR3 (N7390, N7381, N568, N3838);
xor XOR2 (N7391, N7390, N1956);
xor XOR2 (N7392, N7383, N724);
nor NOR2 (N7393, N7384, N7035);
buf BUF1 (N7394, N7382);
buf BUF1 (N7395, N7388);
and AND4 (N7396, N7394, N4776, N6502, N1868);
and AND4 (N7397, N7385, N3960, N7300, N3850);
xor XOR2 (N7398, N7396, N1185);
nor NOR3 (N7399, N7392, N4176, N6123);
not NOT1 (N7400, N7389);
or OR2 (N7401, N7395, N7073);
nand NAND3 (N7402, N7380, N7284, N1585);
nor NOR3 (N7403, N7393, N5404, N2789);
xor XOR2 (N7404, N7387, N4159);
and AND3 (N7405, N7397, N3410, N1208);
buf BUF1 (N7406, N7363);
xor XOR2 (N7407, N7401, N4425);
or OR3 (N7408, N7402, N1275, N3500);
buf BUF1 (N7409, N7405);
not NOT1 (N7410, N7406);
and AND4 (N7411, N7391, N805, N3812, N332);
and AND3 (N7412, N7400, N6978, N4320);
xor XOR2 (N7413, N7398, N5023);
or OR2 (N7414, N7413, N6265);
and AND4 (N7415, N7404, N3966, N1428, N7000);
or OR4 (N7416, N7403, N1634, N1831, N3783);
and AND3 (N7417, N7416, N4506, N2538);
not NOT1 (N7418, N7417);
buf BUF1 (N7419, N7407);
not NOT1 (N7420, N7419);
nor NOR3 (N7421, N7420, N4413, N6751);
xor XOR2 (N7422, N7408, N210);
not NOT1 (N7423, N7410);
or OR4 (N7424, N7422, N5630, N4695, N148);
or OR4 (N7425, N7421, N5945, N6986, N3904);
or OR3 (N7426, N7411, N2506, N3704);
nand NAND2 (N7427, N7412, N2466);
buf BUF1 (N7428, N7426);
and AND4 (N7429, N7418, N1607, N3391, N235);
nand NAND3 (N7430, N7424, N1528, N5038);
not NOT1 (N7431, N7428);
nand NAND2 (N7432, N7423, N1002);
nor NOR2 (N7433, N7415, N3192);
not NOT1 (N7434, N7399);
xor XOR2 (N7435, N7425, N4886);
nand NAND4 (N7436, N7429, N246, N5789, N1645);
not NOT1 (N7437, N7435);
nor NOR4 (N7438, N7430, N3365, N1929, N1038);
xor XOR2 (N7439, N7414, N2855);
not NOT1 (N7440, N7434);
or OR2 (N7441, N7438, N4148);
buf BUF1 (N7442, N7437);
and AND3 (N7443, N7436, N4275, N3514);
not NOT1 (N7444, N7432);
buf BUF1 (N7445, N7443);
or OR2 (N7446, N7433, N5820);
nor NOR4 (N7447, N7409, N5403, N4413, N6632);
buf BUF1 (N7448, N7444);
buf BUF1 (N7449, N7442);
xor XOR2 (N7450, N7448, N540);
and AND2 (N7451, N7449, N5712);
or OR3 (N7452, N7427, N1563, N254);
nand NAND3 (N7453, N7451, N6875, N2145);
buf BUF1 (N7454, N7439);
nor NOR2 (N7455, N7454, N5695);
xor XOR2 (N7456, N7447, N5696);
not NOT1 (N7457, N7446);
or OR2 (N7458, N7441, N6885);
or OR3 (N7459, N7440, N3651, N6639);
or OR3 (N7460, N7459, N7336, N7129);
buf BUF1 (N7461, N7453);
xor XOR2 (N7462, N7452, N4065);
xor XOR2 (N7463, N7460, N1060);
xor XOR2 (N7464, N7445, N3951);
nand NAND3 (N7465, N7455, N1923, N4954);
xor XOR2 (N7466, N7465, N2335);
buf BUF1 (N7467, N7462);
and AND3 (N7468, N7457, N1125, N7249);
buf BUF1 (N7469, N7461);
nand NAND4 (N7470, N7469, N3349, N2196, N1922);
xor XOR2 (N7471, N7470, N6881);
not NOT1 (N7472, N7471);
nor NOR2 (N7473, N7458, N1101);
nor NOR4 (N7474, N7456, N6608, N4902, N1711);
buf BUF1 (N7475, N7473);
or OR4 (N7476, N7466, N5220, N3412, N5429);
xor XOR2 (N7477, N7474, N2540);
nor NOR4 (N7478, N7467, N2343, N6900, N5698);
or OR3 (N7479, N7475, N2520, N1375);
nor NOR4 (N7480, N7431, N3440, N617, N3482);
nor NOR3 (N7481, N7477, N7044, N3616);
or OR2 (N7482, N7472, N1596);
and AND3 (N7483, N7463, N552, N6871);
not NOT1 (N7484, N7450);
buf BUF1 (N7485, N7484);
not NOT1 (N7486, N7468);
buf BUF1 (N7487, N7480);
and AND2 (N7488, N7476, N3137);
and AND2 (N7489, N7479, N1238);
buf BUF1 (N7490, N7485);
and AND4 (N7491, N7464, N5540, N5665, N2654);
or OR4 (N7492, N7489, N3205, N3396, N1368);
and AND4 (N7493, N7488, N6459, N7389, N3048);
nor NOR2 (N7494, N7493, N6730);
or OR3 (N7495, N7478, N4170, N4758);
and AND3 (N7496, N7483, N6390, N2995);
and AND2 (N7497, N7494, N5967);
buf BUF1 (N7498, N7492);
or OR3 (N7499, N7486, N6996, N7495);
nor NOR3 (N7500, N7268, N762, N904);
not NOT1 (N7501, N7497);
and AND4 (N7502, N7496, N914, N3328, N1091);
xor XOR2 (N7503, N7482, N1562);
or OR3 (N7504, N7490, N6613, N1340);
buf BUF1 (N7505, N7502);
and AND2 (N7506, N7491, N3533);
or OR3 (N7507, N7505, N1708, N1895);
buf BUF1 (N7508, N7498);
not NOT1 (N7509, N7500);
buf BUF1 (N7510, N7506);
and AND3 (N7511, N7503, N1522, N4812);
nand NAND2 (N7512, N7499, N6671);
or OR2 (N7513, N7507, N1784);
nand NAND2 (N7514, N7481, N934);
nor NOR2 (N7515, N7508, N3355);
xor XOR2 (N7516, N7504, N1431);
buf BUF1 (N7517, N7511);
nor NOR2 (N7518, N7509, N6522);
and AND2 (N7519, N7512, N5008);
and AND4 (N7520, N7516, N6928, N740, N6843);
and AND3 (N7521, N7519, N4178, N1529);
xor XOR2 (N7522, N7517, N2439);
xor XOR2 (N7523, N7514, N3346);
xor XOR2 (N7524, N7523, N3948);
and AND3 (N7525, N7520, N13, N6999);
nor NOR4 (N7526, N7524, N819, N6885, N7351);
nand NAND2 (N7527, N7515, N3788);
xor XOR2 (N7528, N7518, N4950);
or OR4 (N7529, N7525, N2783, N6147, N5036);
and AND3 (N7530, N7522, N33, N37);
nor NOR3 (N7531, N7526, N973, N5335);
not NOT1 (N7532, N7531);
nand NAND4 (N7533, N7529, N1429, N4696, N7279);
not NOT1 (N7534, N7501);
buf BUF1 (N7535, N7510);
xor XOR2 (N7536, N7487, N7385);
and AND2 (N7537, N7535, N880);
nor NOR3 (N7538, N7534, N3787, N2463);
or OR2 (N7539, N7528, N2324);
nand NAND2 (N7540, N7527, N5861);
nor NOR4 (N7541, N7532, N3101, N1858, N5181);
buf BUF1 (N7542, N7537);
nand NAND4 (N7543, N7542, N6232, N963, N1575);
and AND3 (N7544, N7530, N6842, N660);
xor XOR2 (N7545, N7536, N4854);
nor NOR3 (N7546, N7540, N3332, N7444);
xor XOR2 (N7547, N7546, N7467);
nand NAND4 (N7548, N7543, N1912, N854, N4361);
xor XOR2 (N7549, N7539, N7286);
and AND2 (N7550, N7549, N7000);
or OR3 (N7551, N7521, N967, N4823);
xor XOR2 (N7552, N7513, N110);
buf BUF1 (N7553, N7533);
xor XOR2 (N7554, N7538, N7080);
and AND2 (N7555, N7541, N3457);
nor NOR3 (N7556, N7548, N3619, N2581);
nand NAND4 (N7557, N7547, N4285, N1311, N713);
and AND4 (N7558, N7545, N349, N1705, N2501);
and AND2 (N7559, N7558, N6899);
nor NOR2 (N7560, N7559, N4781);
and AND4 (N7561, N7553, N3933, N858, N5825);
nor NOR2 (N7562, N7561, N1482);
xor XOR2 (N7563, N7562, N907);
buf BUF1 (N7564, N7556);
nor NOR2 (N7565, N7551, N4989);
nand NAND4 (N7566, N7554, N2953, N4434, N5771);
or OR4 (N7567, N7550, N5307, N742, N1034);
buf BUF1 (N7568, N7564);
nor NOR2 (N7569, N7567, N1902);
not NOT1 (N7570, N7544);
xor XOR2 (N7571, N7557, N5961);
xor XOR2 (N7572, N7552, N6993);
and AND3 (N7573, N7566, N7355, N4404);
or OR3 (N7574, N7569, N7332, N6565);
nor NOR2 (N7575, N7563, N3574);
and AND3 (N7576, N7555, N5109, N113);
xor XOR2 (N7577, N7565, N5853);
or OR4 (N7578, N7560, N5404, N787, N1718);
nand NAND2 (N7579, N7577, N5989);
nor NOR4 (N7580, N7570, N7032, N2714, N5110);
nor NOR3 (N7581, N7568, N2633, N1850);
buf BUF1 (N7582, N7575);
nor NOR2 (N7583, N7578, N3691);
and AND4 (N7584, N7583, N6056, N3617, N1988);
not NOT1 (N7585, N7574);
or OR2 (N7586, N7580, N102);
xor XOR2 (N7587, N7572, N1860);
and AND2 (N7588, N7571, N2541);
not NOT1 (N7589, N7588);
not NOT1 (N7590, N7581);
nand NAND4 (N7591, N7584, N2790, N2820, N3680);
xor XOR2 (N7592, N7590, N2387);
nor NOR4 (N7593, N7576, N3643, N4343, N7387);
xor XOR2 (N7594, N7582, N4445);
nand NAND4 (N7595, N7593, N1874, N5675, N2206);
or OR4 (N7596, N7573, N4188, N1398, N1895);
or OR4 (N7597, N7587, N2074, N1887, N29);
or OR4 (N7598, N7591, N298, N5063, N2616);
buf BUF1 (N7599, N7589);
or OR3 (N7600, N7598, N1567, N5027);
nor NOR3 (N7601, N7585, N1051, N162);
nor NOR2 (N7602, N7596, N750);
nand NAND4 (N7603, N7600, N3880, N4319, N3359);
nand NAND3 (N7604, N7595, N1079, N2766);
and AND4 (N7605, N7586, N5638, N6315, N7385);
or OR4 (N7606, N7597, N5688, N2759, N4398);
nand NAND2 (N7607, N7601, N1418);
xor XOR2 (N7608, N7599, N4484);
buf BUF1 (N7609, N7592);
not NOT1 (N7610, N7603);
nand NAND2 (N7611, N7606, N6887);
nor NOR3 (N7612, N7604, N3708, N2269);
or OR2 (N7613, N7611, N2281);
or OR2 (N7614, N7613, N3910);
buf BUF1 (N7615, N7612);
or OR4 (N7616, N7607, N4213, N4698, N2322);
nor NOR3 (N7617, N7605, N2000, N5745);
not NOT1 (N7618, N7594);
xor XOR2 (N7619, N7615, N5886);
and AND4 (N7620, N7602, N629, N2769, N3035);
or OR2 (N7621, N7620, N474);
or OR3 (N7622, N7618, N6620, N742);
or OR4 (N7623, N7621, N2102, N2226, N1806);
xor XOR2 (N7624, N7614, N893);
and AND3 (N7625, N7616, N1319, N7537);
nor NOR4 (N7626, N7617, N2429, N1650, N1151);
xor XOR2 (N7627, N7623, N6625);
not NOT1 (N7628, N7610);
xor XOR2 (N7629, N7624, N3020);
nor NOR3 (N7630, N7622, N3919, N7404);
not NOT1 (N7631, N7627);
xor XOR2 (N7632, N7619, N5762);
buf BUF1 (N7633, N7625);
buf BUF1 (N7634, N7628);
or OR3 (N7635, N7629, N3432, N7345);
not NOT1 (N7636, N7632);
buf BUF1 (N7637, N7634);
or OR2 (N7638, N7636, N1941);
nor NOR3 (N7639, N7638, N1798, N725);
buf BUF1 (N7640, N7630);
nor NOR2 (N7641, N7579, N6351);
buf BUF1 (N7642, N7609);
buf BUF1 (N7643, N7640);
not NOT1 (N7644, N7608);
nor NOR2 (N7645, N7631, N77);
not NOT1 (N7646, N7633);
not NOT1 (N7647, N7626);
nand NAND3 (N7648, N7635, N899, N856);
buf BUF1 (N7649, N7641);
or OR2 (N7650, N7643, N2854);
xor XOR2 (N7651, N7649, N4819);
and AND3 (N7652, N7646, N6782, N4190);
xor XOR2 (N7653, N7642, N936);
or OR4 (N7654, N7652, N235, N489, N6390);
or OR3 (N7655, N7648, N4663, N3109);
nand NAND2 (N7656, N7654, N597);
nor NOR4 (N7657, N7645, N1034, N1414, N6711);
nor NOR4 (N7658, N7644, N3192, N3299, N5401);
and AND2 (N7659, N7658, N2682);
or OR3 (N7660, N7647, N7491, N6441);
not NOT1 (N7661, N7659);
xor XOR2 (N7662, N7657, N2330);
not NOT1 (N7663, N7656);
buf BUF1 (N7664, N7650);
not NOT1 (N7665, N7664);
or OR2 (N7666, N7660, N147);
buf BUF1 (N7667, N7666);
or OR2 (N7668, N7639, N7299);
xor XOR2 (N7669, N7665, N2064);
or OR3 (N7670, N7651, N6873, N6983);
nand NAND3 (N7671, N7661, N4667, N3853);
nand NAND3 (N7672, N7671, N2051, N4170);
or OR3 (N7673, N7670, N4177, N2793);
not NOT1 (N7674, N7672);
nand NAND3 (N7675, N7655, N5596, N1995);
xor XOR2 (N7676, N7667, N1327);
nand NAND4 (N7677, N7674, N3986, N5415, N5528);
nor NOR2 (N7678, N7669, N5384);
or OR3 (N7679, N7662, N87, N2570);
and AND3 (N7680, N7668, N4718, N5984);
buf BUF1 (N7681, N7677);
buf BUF1 (N7682, N7663);
nor NOR3 (N7683, N7680, N2205, N1955);
not NOT1 (N7684, N7683);
not NOT1 (N7685, N7637);
buf BUF1 (N7686, N7685);
xor XOR2 (N7687, N7653, N4307);
xor XOR2 (N7688, N7676, N4363);
and AND3 (N7689, N7684, N688, N3257);
nand NAND3 (N7690, N7689, N4776, N4558);
nor NOR3 (N7691, N7682, N7468, N2662);
not NOT1 (N7692, N7681);
buf BUF1 (N7693, N7686);
not NOT1 (N7694, N7690);
buf BUF1 (N7695, N7687);
xor XOR2 (N7696, N7693, N6936);
buf BUF1 (N7697, N7678);
nand NAND3 (N7698, N7696, N3240, N551);
nor NOR3 (N7699, N7688, N1876, N1028);
xor XOR2 (N7700, N7697, N1045);
nor NOR4 (N7701, N7699, N6179, N1182, N2514);
and AND4 (N7702, N7679, N6932, N5712, N5290);
xor XOR2 (N7703, N7675, N7501);
not NOT1 (N7704, N7695);
or OR2 (N7705, N7701, N47);
nand NAND2 (N7706, N7692, N4977);
nor NOR3 (N7707, N7700, N6160, N355);
buf BUF1 (N7708, N7706);
or OR4 (N7709, N7708, N1598, N4942, N5652);
nor NOR2 (N7710, N7702, N7342);
xor XOR2 (N7711, N7703, N6190);
nand NAND2 (N7712, N7707, N973);
nand NAND3 (N7713, N7691, N4110, N1672);
and AND4 (N7714, N7713, N175, N5389, N834);
not NOT1 (N7715, N7704);
not NOT1 (N7716, N7709);
buf BUF1 (N7717, N7711);
nor NOR2 (N7718, N7717, N662);
and AND4 (N7719, N7710, N5688, N2031, N4001);
and AND4 (N7720, N7719, N2777, N5271, N640);
nand NAND3 (N7721, N7712, N5663, N624);
or OR2 (N7722, N7694, N6667);
not NOT1 (N7723, N7715);
and AND4 (N7724, N7718, N4505, N1886, N2871);
or OR3 (N7725, N7720, N4579, N339);
nand NAND3 (N7726, N7705, N5047, N924);
nor NOR2 (N7727, N7716, N2140);
and AND4 (N7728, N7698, N3921, N4291, N4440);
or OR4 (N7729, N7721, N3200, N2185, N4066);
or OR3 (N7730, N7725, N6025, N1227);
nor NOR3 (N7731, N7729, N4088, N543);
xor XOR2 (N7732, N7728, N6404);
and AND4 (N7733, N7722, N229, N3122, N2877);
nand NAND4 (N7734, N7733, N3081, N6421, N4638);
nor NOR2 (N7735, N7731, N6437);
not NOT1 (N7736, N7673);
nand NAND2 (N7737, N7734, N650);
xor XOR2 (N7738, N7714, N385);
xor XOR2 (N7739, N7723, N1430);
nand NAND2 (N7740, N7735, N2022);
not NOT1 (N7741, N7739);
xor XOR2 (N7742, N7738, N4156);
buf BUF1 (N7743, N7730);
buf BUF1 (N7744, N7727);
or OR4 (N7745, N7732, N2032, N4240, N6227);
xor XOR2 (N7746, N7744, N55);
or OR2 (N7747, N7745, N140);
xor XOR2 (N7748, N7736, N264);
buf BUF1 (N7749, N7740);
xor XOR2 (N7750, N7748, N1543);
or OR2 (N7751, N7741, N5180);
xor XOR2 (N7752, N7726, N2055);
buf BUF1 (N7753, N7751);
and AND2 (N7754, N7749, N69);
and AND3 (N7755, N7742, N845, N2957);
not NOT1 (N7756, N7746);
nand NAND4 (N7757, N7747, N3910, N2789, N955);
nor NOR4 (N7758, N7756, N4542, N6772, N2699);
not NOT1 (N7759, N7757);
buf BUF1 (N7760, N7754);
buf BUF1 (N7761, N7737);
nor NOR3 (N7762, N7724, N6695, N343);
and AND2 (N7763, N7743, N562);
not NOT1 (N7764, N7759);
or OR3 (N7765, N7755, N1697, N7369);
xor XOR2 (N7766, N7763, N4531);
not NOT1 (N7767, N7761);
and AND3 (N7768, N7750, N2356, N644);
buf BUF1 (N7769, N7765);
buf BUF1 (N7770, N7766);
buf BUF1 (N7771, N7767);
or OR3 (N7772, N7753, N525, N2968);
not NOT1 (N7773, N7771);
or OR3 (N7774, N7773, N2692, N4582);
nand NAND4 (N7775, N7769, N2082, N1159, N7344);
nand NAND4 (N7776, N7774, N7157, N2056, N5818);
not NOT1 (N7777, N7758);
or OR3 (N7778, N7777, N6800, N4593);
nor NOR2 (N7779, N7776, N5791);
not NOT1 (N7780, N7762);
not NOT1 (N7781, N7760);
nor NOR2 (N7782, N7764, N3996);
or OR3 (N7783, N7768, N6404, N727);
nor NOR3 (N7784, N7775, N2443, N4600);
nand NAND3 (N7785, N7783, N6655, N6958);
buf BUF1 (N7786, N7784);
buf BUF1 (N7787, N7752);
xor XOR2 (N7788, N7770, N2033);
nand NAND3 (N7789, N7786, N7257, N1190);
nand NAND4 (N7790, N7789, N7611, N2825, N4425);
and AND2 (N7791, N7778, N7266);
xor XOR2 (N7792, N7787, N6179);
nor NOR4 (N7793, N7788, N5744, N6736, N5897);
and AND4 (N7794, N7781, N1943, N4455, N3353);
not NOT1 (N7795, N7772);
nor NOR2 (N7796, N7785, N7068);
not NOT1 (N7797, N7795);
xor XOR2 (N7798, N7782, N3802);
nand NAND2 (N7799, N7796, N1300);
buf BUF1 (N7800, N7794);
not NOT1 (N7801, N7780);
buf BUF1 (N7802, N7793);
not NOT1 (N7803, N7779);
nand NAND4 (N7804, N7802, N5005, N2730, N5472);
not NOT1 (N7805, N7791);
and AND2 (N7806, N7798, N6329);
not NOT1 (N7807, N7800);
not NOT1 (N7808, N7790);
nand NAND4 (N7809, N7808, N6801, N7547, N1378);
or OR4 (N7810, N7801, N7395, N4796, N5623);
buf BUF1 (N7811, N7799);
or OR4 (N7812, N7797, N3999, N1898, N1211);
nand NAND2 (N7813, N7812, N1909);
and AND4 (N7814, N7807, N4836, N6169, N7665);
nor NOR4 (N7815, N7810, N3967, N3203, N4966);
or OR4 (N7816, N7813, N3867, N6565, N424);
and AND3 (N7817, N7803, N5637, N722);
and AND4 (N7818, N7805, N3628, N1459, N5267);
nor NOR3 (N7819, N7817, N48, N2320);
and AND4 (N7820, N7818, N7118, N3424, N2414);
xor XOR2 (N7821, N7814, N7012);
xor XOR2 (N7822, N7815, N6743);
buf BUF1 (N7823, N7804);
not NOT1 (N7824, N7819);
not NOT1 (N7825, N7822);
not NOT1 (N7826, N7811);
not NOT1 (N7827, N7792);
xor XOR2 (N7828, N7821, N400);
not NOT1 (N7829, N7825);
not NOT1 (N7830, N7828);
not NOT1 (N7831, N7806);
xor XOR2 (N7832, N7824, N7232);
nor NOR2 (N7833, N7829, N6895);
xor XOR2 (N7834, N7833, N6752);
and AND4 (N7835, N7834, N2260, N4316, N5830);
not NOT1 (N7836, N7809);
and AND2 (N7837, N7820, N5288);
or OR2 (N7838, N7830, N7538);
and AND3 (N7839, N7831, N6969, N1260);
or OR4 (N7840, N7832, N6002, N5066, N6737);
buf BUF1 (N7841, N7836);
or OR2 (N7842, N7840, N4923);
buf BUF1 (N7843, N7823);
buf BUF1 (N7844, N7816);
nand NAND3 (N7845, N7827, N4589, N946);
or OR3 (N7846, N7835, N4244, N3011);
or OR3 (N7847, N7841, N2205, N2202);
nor NOR2 (N7848, N7842, N5462);
buf BUF1 (N7849, N7848);
not NOT1 (N7850, N7839);
xor XOR2 (N7851, N7847, N4584);
not NOT1 (N7852, N7849);
xor XOR2 (N7853, N7843, N2133);
not NOT1 (N7854, N7852);
xor XOR2 (N7855, N7853, N1633);
xor XOR2 (N7856, N7855, N7319);
nor NOR4 (N7857, N7850, N2128, N2476, N6217);
not NOT1 (N7858, N7838);
xor XOR2 (N7859, N7854, N5815);
not NOT1 (N7860, N7857);
nor NOR2 (N7861, N7859, N308);
nand NAND4 (N7862, N7856, N5567, N4298, N55);
nand NAND4 (N7863, N7851, N5981, N2430, N7372);
xor XOR2 (N7864, N7837, N1765);
buf BUF1 (N7865, N7862);
and AND4 (N7866, N7861, N5432, N756, N6529);
not NOT1 (N7867, N7846);
nor NOR4 (N7868, N7860, N2120, N7725, N1208);
nor NOR3 (N7869, N7844, N2133, N7290);
nand NAND3 (N7870, N7864, N5686, N935);
not NOT1 (N7871, N7826);
buf BUF1 (N7872, N7868);
not NOT1 (N7873, N7871);
xor XOR2 (N7874, N7873, N4790);
or OR4 (N7875, N7867, N949, N2208, N7253);
nor NOR3 (N7876, N7845, N6981, N2135);
nand NAND3 (N7877, N7876, N71, N5250);
or OR3 (N7878, N7863, N4906, N2179);
not NOT1 (N7879, N7872);
nor NOR4 (N7880, N7879, N4592, N6155, N7450);
xor XOR2 (N7881, N7869, N7273);
nor NOR3 (N7882, N7858, N1338, N387);
buf BUF1 (N7883, N7877);
buf BUF1 (N7884, N7881);
and AND4 (N7885, N7884, N7685, N1999, N7471);
or OR4 (N7886, N7882, N6480, N1356, N7481);
xor XOR2 (N7887, N7874, N4850);
nand NAND3 (N7888, N7885, N306, N5932);
or OR4 (N7889, N7866, N3295, N3780, N7605);
not NOT1 (N7890, N7887);
buf BUF1 (N7891, N7888);
xor XOR2 (N7892, N7875, N3872);
not NOT1 (N7893, N7892);
not NOT1 (N7894, N7880);
not NOT1 (N7895, N7865);
and AND2 (N7896, N7895, N5317);
not NOT1 (N7897, N7870);
or OR2 (N7898, N7883, N3165);
or OR3 (N7899, N7893, N3828, N7315);
xor XOR2 (N7900, N7898, N4191);
nand NAND3 (N7901, N7890, N7794, N3010);
or OR4 (N7902, N7878, N3935, N3325, N6997);
nor NOR4 (N7903, N7899, N604, N2559, N7492);
not NOT1 (N7904, N7901);
xor XOR2 (N7905, N7886, N3339);
buf BUF1 (N7906, N7903);
xor XOR2 (N7907, N7905, N5218);
nand NAND4 (N7908, N7894, N103, N7541, N2989);
or OR3 (N7909, N7891, N3643, N7448);
nand NAND2 (N7910, N7904, N7192);
or OR4 (N7911, N7902, N7402, N5886, N4353);
and AND4 (N7912, N7897, N7250, N10, N1193);
and AND3 (N7913, N7911, N3325, N4597);
xor XOR2 (N7914, N7900, N7427);
buf BUF1 (N7915, N7914);
and AND3 (N7916, N7906, N4837, N7471);
and AND4 (N7917, N7913, N2875, N2789, N2494);
or OR2 (N7918, N7896, N5525);
or OR2 (N7919, N7910, N4783);
nor NOR3 (N7920, N7915, N7884, N7092);
nor NOR2 (N7921, N7920, N5494);
or OR4 (N7922, N7912, N3450, N1055, N3255);
xor XOR2 (N7923, N7918, N866);
and AND3 (N7924, N7909, N5345, N6525);
nand NAND4 (N7925, N7922, N3349, N5222, N5701);
buf BUF1 (N7926, N7916);
nand NAND4 (N7927, N7925, N6264, N2071, N2634);
not NOT1 (N7928, N7924);
buf BUF1 (N7929, N7907);
xor XOR2 (N7930, N7921, N5411);
nand NAND4 (N7931, N7926, N6777, N7510, N802);
not NOT1 (N7932, N7919);
not NOT1 (N7933, N7917);
or OR3 (N7934, N7932, N75, N4847);
not NOT1 (N7935, N7931);
nor NOR4 (N7936, N7933, N3222, N6666, N5841);
xor XOR2 (N7937, N7929, N5523);
buf BUF1 (N7938, N7927);
or OR4 (N7939, N7923, N2929, N1985, N1045);
xor XOR2 (N7940, N7934, N5556);
nor NOR4 (N7941, N7928, N4113, N7033, N5156);
nand NAND3 (N7942, N7939, N1946, N5294);
nor NOR3 (N7943, N7940, N2079, N7707);
xor XOR2 (N7944, N7936, N257);
buf BUF1 (N7945, N7889);
buf BUF1 (N7946, N7908);
or OR3 (N7947, N7945, N903, N558);
buf BUF1 (N7948, N7937);
not NOT1 (N7949, N7946);
nor NOR2 (N7950, N7944, N4765);
buf BUF1 (N7951, N7950);
xor XOR2 (N7952, N7951, N4424);
buf BUF1 (N7953, N7949);
nor NOR3 (N7954, N7935, N5029, N7612);
or OR2 (N7955, N7954, N7888);
xor XOR2 (N7956, N7942, N7424);
nor NOR2 (N7957, N7941, N326);
nor NOR2 (N7958, N7943, N323);
or OR3 (N7959, N7953, N5478, N2556);
or OR2 (N7960, N7947, N3402);
xor XOR2 (N7961, N7952, N2963);
xor XOR2 (N7962, N7960, N4535);
buf BUF1 (N7963, N7955);
xor XOR2 (N7964, N7962, N5481);
buf BUF1 (N7965, N7957);
not NOT1 (N7966, N7964);
buf BUF1 (N7967, N7938);
nand NAND2 (N7968, N7961, N6829);
buf BUF1 (N7969, N7967);
nor NOR2 (N7970, N7959, N6160);
xor XOR2 (N7971, N7969, N7273);
and AND2 (N7972, N7958, N7772);
xor XOR2 (N7973, N7963, N6265);
or OR4 (N7974, N7966, N1675, N2754, N2369);
xor XOR2 (N7975, N7968, N6639);
nor NOR3 (N7976, N7956, N3580, N2107);
nor NOR4 (N7977, N7930, N7249, N7952, N7318);
nand NAND2 (N7978, N7974, N4193);
nand NAND2 (N7979, N7948, N2645);
and AND2 (N7980, N7975, N5224);
buf BUF1 (N7981, N7970);
nor NOR2 (N7982, N7979, N6666);
or OR4 (N7983, N7978, N5170, N4807, N7375);
xor XOR2 (N7984, N7971, N2790);
not NOT1 (N7985, N7980);
nand NAND4 (N7986, N7976, N7730, N5408, N7138);
nand NAND2 (N7987, N7981, N7903);
nand NAND4 (N7988, N7977, N3806, N3464, N5101);
not NOT1 (N7989, N7982);
not NOT1 (N7990, N7988);
xor XOR2 (N7991, N7986, N34);
nand NAND4 (N7992, N7972, N3447, N1482, N1583);
nor NOR3 (N7993, N7965, N3567, N953);
not NOT1 (N7994, N7987);
not NOT1 (N7995, N7973);
xor XOR2 (N7996, N7984, N6197);
nor NOR3 (N7997, N7993, N6951, N2371);
nand NAND2 (N7998, N7995, N6315);
and AND2 (N7999, N7997, N950);
and AND2 (N8000, N7994, N6028);
not NOT1 (N8001, N8000);
or OR2 (N8002, N7985, N6088);
not NOT1 (N8003, N7983);
nand NAND3 (N8004, N7989, N2236, N7142);
xor XOR2 (N8005, N8002, N863);
buf BUF1 (N8006, N8004);
and AND4 (N8007, N8005, N4584, N5157, N5550);
or OR4 (N8008, N7990, N3978, N1661, N2685);
xor XOR2 (N8009, N7996, N2634);
and AND4 (N8010, N8007, N1062, N3702, N7303);
endmodule