// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N512,N510,N484,N491,N511,N485,N513,N507,N514,N515;

nor NOR4 (N16, N6, N6, N1, N8);
xor XOR2 (N17, N12, N14);
and AND2 (N18, N14, N14);
nand NAND3 (N19, N6, N13, N12);
buf BUF1 (N20, N9);
or OR2 (N21, N7, N2);
and AND3 (N22, N5, N21, N3);
nand NAND2 (N23, N13, N2);
xor XOR2 (N24, N16, N23);
and AND4 (N25, N13, N1, N17, N4);
xor XOR2 (N26, N4, N20);
nand NAND4 (N27, N5, N8, N26, N14);
nor NOR4 (N28, N9, N25, N26, N26);
or OR2 (N29, N17, N15);
nand NAND4 (N30, N21, N5, N28, N14);
nor NOR4 (N31, N15, N30, N13, N11);
not NOT1 (N32, N3);
not NOT1 (N33, N15);
or OR4 (N34, N13, N26, N4, N16);
xor XOR2 (N35, N27, N5);
not NOT1 (N36, N24);
and AND2 (N37, N32, N13);
buf BUF1 (N38, N36);
not NOT1 (N39, N22);
not NOT1 (N40, N37);
xor XOR2 (N41, N18, N16);
buf BUF1 (N42, N41);
or OR3 (N43, N35, N15, N12);
or OR4 (N44, N31, N3, N34, N2);
nand NAND4 (N45, N38, N31, N44, N43);
nand NAND4 (N46, N9, N31, N27, N16);
buf BUF1 (N47, N44);
nand NAND3 (N48, N47, N22, N3);
nor NOR4 (N49, N1, N11, N2, N25);
buf BUF1 (N50, N49);
nor NOR4 (N51, N19, N14, N5, N25);
buf BUF1 (N52, N33);
not NOT1 (N53, N29);
xor XOR2 (N54, N42, N3);
nand NAND4 (N55, N39, N42, N35, N32);
xor XOR2 (N56, N50, N55);
and AND2 (N57, N50, N11);
not NOT1 (N58, N57);
buf BUF1 (N59, N54);
buf BUF1 (N60, N58);
buf BUF1 (N61, N56);
nand NAND2 (N62, N45, N46);
buf BUF1 (N63, N61);
or OR4 (N64, N49, N62, N39, N32);
not NOT1 (N65, N48);
buf BUF1 (N66, N45);
nand NAND3 (N67, N63, N5, N9);
or OR4 (N68, N59, N23, N54, N54);
nand NAND3 (N69, N66, N4, N56);
buf BUF1 (N70, N69);
nor NOR4 (N71, N52, N5, N8, N53);
buf BUF1 (N72, N64);
not NOT1 (N73, N39);
nand NAND4 (N74, N65, N24, N28, N72);
buf BUF1 (N75, N22);
buf BUF1 (N76, N60);
nand NAND4 (N77, N71, N29, N32, N66);
and AND3 (N78, N73, N55, N14);
buf BUF1 (N79, N68);
and AND2 (N80, N78, N43);
nand NAND2 (N81, N77, N3);
buf BUF1 (N82, N67);
or OR4 (N83, N51, N16, N5, N17);
and AND4 (N84, N76, N32, N11, N59);
buf BUF1 (N85, N83);
and AND3 (N86, N79, N51, N59);
nand NAND3 (N87, N75, N83, N54);
nor NOR4 (N88, N85, N68, N75, N62);
xor XOR2 (N89, N88, N35);
nor NOR2 (N90, N86, N58);
or OR2 (N91, N87, N83);
nor NOR3 (N92, N89, N59, N14);
buf BUF1 (N93, N84);
nand NAND4 (N94, N40, N6, N52, N68);
nor NOR2 (N95, N74, N79);
not NOT1 (N96, N90);
and AND3 (N97, N96, N52, N16);
buf BUF1 (N98, N70);
not NOT1 (N99, N93);
xor XOR2 (N100, N94, N96);
buf BUF1 (N101, N100);
and AND4 (N102, N97, N20, N85, N26);
or OR4 (N103, N98, N47, N88, N50);
and AND3 (N104, N81, N16, N41);
not NOT1 (N105, N104);
xor XOR2 (N106, N103, N71);
buf BUF1 (N107, N92);
and AND3 (N108, N102, N41, N72);
buf BUF1 (N109, N108);
and AND4 (N110, N95, N54, N64, N101);
xor XOR2 (N111, N89, N89);
and AND3 (N112, N110, N41, N72);
or OR4 (N113, N82, N36, N4, N79);
and AND3 (N114, N107, N108, N86);
or OR3 (N115, N114, N111, N34);
nor NOR2 (N116, N85, N54);
not NOT1 (N117, N106);
nand NAND4 (N118, N116, N33, N90, N30);
nand NAND3 (N119, N115, N87, N104);
nand NAND3 (N120, N91, N110, N30);
not NOT1 (N121, N113);
nor NOR2 (N122, N99, N2);
or OR3 (N123, N118, N3, N67);
buf BUF1 (N124, N120);
and AND3 (N125, N105, N52, N84);
buf BUF1 (N126, N124);
nor NOR3 (N127, N80, N72, N115);
not NOT1 (N128, N127);
or OR4 (N129, N121, N62, N101, N52);
xor XOR2 (N130, N117, N108);
or OR2 (N131, N126, N65);
or OR3 (N132, N119, N43, N28);
and AND3 (N133, N130, N75, N24);
nand NAND4 (N134, N112, N71, N69, N34);
and AND4 (N135, N134, N64, N115, N104);
or OR3 (N136, N132, N23, N101);
nand NAND4 (N137, N136, N11, N31, N87);
buf BUF1 (N138, N128);
and AND2 (N139, N138, N51);
or OR4 (N140, N139, N97, N117, N64);
or OR4 (N141, N135, N102, N54, N65);
xor XOR2 (N142, N123, N10);
not NOT1 (N143, N109);
not NOT1 (N144, N141);
or OR3 (N145, N125, N50, N64);
not NOT1 (N146, N145);
or OR2 (N147, N142, N58);
and AND3 (N148, N137, N138, N34);
not NOT1 (N149, N140);
xor XOR2 (N150, N149, N114);
nand NAND4 (N151, N122, N10, N83, N58);
nand NAND4 (N152, N146, N136, N123, N18);
nor NOR2 (N153, N147, N27);
not NOT1 (N154, N148);
or OR3 (N155, N152, N37, N154);
buf BUF1 (N156, N143);
xor XOR2 (N157, N47, N26);
buf BUF1 (N158, N156);
buf BUF1 (N159, N158);
and AND2 (N160, N150, N3);
not NOT1 (N161, N133);
and AND4 (N162, N159, N11, N140, N18);
nand NAND4 (N163, N161, N106, N56, N150);
nand NAND2 (N164, N160, N145);
or OR3 (N165, N153, N84, N71);
nor NOR2 (N166, N129, N66);
buf BUF1 (N167, N144);
nor NOR3 (N168, N164, N48, N161);
nand NAND3 (N169, N151, N145, N58);
xor XOR2 (N170, N131, N155);
not NOT1 (N171, N151);
buf BUF1 (N172, N163);
nor NOR3 (N173, N168, N61, N33);
nor NOR4 (N174, N157, N43, N107, N158);
nand NAND3 (N175, N174, N76, N57);
buf BUF1 (N176, N173);
nor NOR2 (N177, N167, N81);
and AND3 (N178, N172, N162, N36);
buf BUF1 (N179, N128);
xor XOR2 (N180, N170, N132);
xor XOR2 (N181, N180, N15);
nand NAND2 (N182, N177, N65);
or OR4 (N183, N165, N145, N20, N76);
buf BUF1 (N184, N175);
nand NAND2 (N185, N166, N136);
not NOT1 (N186, N179);
buf BUF1 (N187, N181);
nor NOR3 (N188, N178, N178, N120);
not NOT1 (N189, N184);
or OR3 (N190, N176, N177, N133);
nand NAND3 (N191, N187, N190, N189);
xor XOR2 (N192, N117, N23);
buf BUF1 (N193, N6);
not NOT1 (N194, N183);
buf BUF1 (N195, N193);
nand NAND2 (N196, N185, N116);
or OR4 (N197, N169, N125, N39, N162);
not NOT1 (N198, N197);
not NOT1 (N199, N188);
nor NOR2 (N200, N192, N41);
nand NAND4 (N201, N186, N13, N118, N180);
or OR4 (N202, N199, N130, N45, N197);
and AND3 (N203, N182, N172, N145);
and AND4 (N204, N198, N157, N181, N66);
xor XOR2 (N205, N196, N183);
nor NOR2 (N206, N191, N49);
or OR2 (N207, N200, N72);
buf BUF1 (N208, N204);
or OR2 (N209, N194, N199);
buf BUF1 (N210, N207);
or OR2 (N211, N209, N64);
or OR2 (N212, N210, N63);
or OR2 (N213, N205, N4);
buf BUF1 (N214, N201);
not NOT1 (N215, N202);
not NOT1 (N216, N215);
buf BUF1 (N217, N206);
and AND4 (N218, N216, N152, N88, N79);
and AND3 (N219, N195, N25, N117);
or OR3 (N220, N218, N178, N45);
xor XOR2 (N221, N171, N103);
and AND2 (N222, N221, N155);
not NOT1 (N223, N203);
xor XOR2 (N224, N211, N206);
buf BUF1 (N225, N212);
nor NOR2 (N226, N214, N116);
or OR4 (N227, N213, N148, N219, N53);
not NOT1 (N228, N184);
buf BUF1 (N229, N208);
nand NAND3 (N230, N225, N20, N15);
buf BUF1 (N231, N226);
buf BUF1 (N232, N229);
buf BUF1 (N233, N232);
nand NAND3 (N234, N233, N88, N73);
buf BUF1 (N235, N223);
not NOT1 (N236, N234);
nand NAND2 (N237, N222, N112);
xor XOR2 (N238, N228, N85);
buf BUF1 (N239, N230);
nand NAND4 (N240, N217, N217, N5, N220);
xor XOR2 (N241, N147, N40);
nor NOR4 (N242, N231, N227, N219, N83);
nand NAND3 (N243, N47, N158, N22);
nor NOR3 (N244, N236, N198, N74);
nor NOR4 (N245, N239, N211, N85, N3);
xor XOR2 (N246, N237, N131);
and AND3 (N247, N246, N74, N67);
nand NAND4 (N248, N240, N146, N34, N129);
nand NAND4 (N249, N244, N222, N113, N121);
buf BUF1 (N250, N242);
buf BUF1 (N251, N224);
buf BUF1 (N252, N238);
or OR2 (N253, N241, N178);
xor XOR2 (N254, N247, N45);
xor XOR2 (N255, N254, N109);
nand NAND3 (N256, N255, N35, N13);
or OR2 (N257, N256, N234);
nor NOR3 (N258, N257, N218, N83);
not NOT1 (N259, N243);
xor XOR2 (N260, N252, N89);
and AND3 (N261, N260, N110, N171);
nand NAND3 (N262, N250, N9, N149);
buf BUF1 (N263, N261);
and AND3 (N264, N251, N81, N115);
nand NAND4 (N265, N262, N164, N131, N28);
not NOT1 (N266, N263);
and AND3 (N267, N245, N133, N144);
nand NAND4 (N268, N248, N31, N221, N95);
xor XOR2 (N269, N264, N92);
and AND3 (N270, N265, N215, N71);
and AND2 (N271, N267, N56);
not NOT1 (N272, N258);
or OR2 (N273, N270, N123);
or OR2 (N274, N272, N51);
nand NAND4 (N275, N273, N80, N52, N141);
nor NOR2 (N276, N253, N255);
xor XOR2 (N277, N269, N36);
buf BUF1 (N278, N275);
nand NAND3 (N279, N259, N176, N212);
and AND3 (N280, N278, N212, N146);
and AND3 (N281, N249, N261, N16);
nor NOR2 (N282, N271, N270);
or OR4 (N283, N277, N44, N211, N247);
or OR3 (N284, N266, N182, N66);
not NOT1 (N285, N274);
xor XOR2 (N286, N235, N198);
xor XOR2 (N287, N281, N253);
or OR2 (N288, N276, N152);
buf BUF1 (N289, N280);
xor XOR2 (N290, N284, N130);
not NOT1 (N291, N288);
not NOT1 (N292, N287);
nor NOR3 (N293, N282, N193, N272);
and AND4 (N294, N292, N11, N221, N116);
and AND3 (N295, N294, N234, N44);
or OR4 (N296, N279, N250, N283, N142);
xor XOR2 (N297, N203, N196);
not NOT1 (N298, N293);
and AND2 (N299, N286, N71);
nand NAND4 (N300, N289, N15, N149, N161);
not NOT1 (N301, N295);
nor NOR4 (N302, N300, N226, N245, N113);
buf BUF1 (N303, N301);
or OR4 (N304, N299, N106, N124, N23);
nor NOR3 (N305, N291, N301, N109);
buf BUF1 (N306, N285);
nor NOR3 (N307, N303, N30, N238);
nor NOR2 (N308, N268, N21);
and AND4 (N309, N296, N187, N186, N172);
or OR4 (N310, N305, N109, N182, N186);
or OR4 (N311, N308, N21, N28, N52);
nand NAND2 (N312, N307, N41);
not NOT1 (N313, N306);
nor NOR4 (N314, N311, N241, N167, N50);
nand NAND4 (N315, N298, N110, N112, N103);
not NOT1 (N316, N309);
buf BUF1 (N317, N290);
xor XOR2 (N318, N310, N200);
nor NOR3 (N319, N312, N17, N64);
or OR3 (N320, N313, N159, N160);
and AND3 (N321, N317, N145, N236);
not NOT1 (N322, N320);
and AND3 (N323, N322, N1, N162);
nand NAND2 (N324, N323, N237);
not NOT1 (N325, N319);
nand NAND2 (N326, N304, N180);
not NOT1 (N327, N314);
or OR3 (N328, N321, N296, N249);
or OR2 (N329, N302, N3);
buf BUF1 (N330, N315);
buf BUF1 (N331, N318);
and AND3 (N332, N329, N137, N299);
not NOT1 (N333, N324);
nor NOR4 (N334, N330, N183, N70, N220);
not NOT1 (N335, N325);
and AND4 (N336, N328, N250, N243, N189);
and AND3 (N337, N297, N166, N209);
xor XOR2 (N338, N332, N220);
xor XOR2 (N339, N334, N232);
nand NAND4 (N340, N326, N311, N193, N117);
xor XOR2 (N341, N333, N36);
and AND3 (N342, N327, N253, N164);
nor NOR3 (N343, N335, N49, N267);
not NOT1 (N344, N341);
nand NAND2 (N345, N331, N272);
and AND2 (N346, N345, N117);
or OR3 (N347, N343, N66, N224);
nor NOR4 (N348, N344, N109, N141, N246);
or OR3 (N349, N316, N319, N266);
buf BUF1 (N350, N349);
or OR3 (N351, N342, N70, N193);
xor XOR2 (N352, N339, N212);
xor XOR2 (N353, N338, N298);
buf BUF1 (N354, N337);
nand NAND4 (N355, N347, N267, N123, N93);
and AND2 (N356, N336, N13);
and AND4 (N357, N356, N224, N180, N93);
and AND3 (N358, N351, N113, N307);
not NOT1 (N359, N354);
buf BUF1 (N360, N346);
buf BUF1 (N361, N350);
nor NOR2 (N362, N348, N13);
not NOT1 (N363, N361);
nor NOR4 (N364, N358, N62, N235, N133);
and AND3 (N365, N364, N133, N330);
nor NOR3 (N366, N357, N362, N146);
not NOT1 (N367, N21);
nor NOR2 (N368, N352, N53);
or OR3 (N369, N368, N292, N159);
or OR2 (N370, N365, N169);
and AND2 (N371, N353, N59);
buf BUF1 (N372, N369);
xor XOR2 (N373, N359, N92);
not NOT1 (N374, N372);
nand NAND3 (N375, N366, N39, N286);
nor NOR4 (N376, N360, N240, N174, N36);
nor NOR4 (N377, N355, N304, N95, N229);
buf BUF1 (N378, N375);
buf BUF1 (N379, N340);
nand NAND2 (N380, N379, N81);
xor XOR2 (N381, N376, N297);
nand NAND4 (N382, N373, N112, N301, N137);
nand NAND2 (N383, N380, N235);
buf BUF1 (N384, N374);
xor XOR2 (N385, N370, N12);
xor XOR2 (N386, N371, N343);
not NOT1 (N387, N386);
or OR3 (N388, N367, N257, N203);
xor XOR2 (N389, N363, N105);
or OR3 (N390, N388, N294, N189);
and AND4 (N391, N390, N265, N66, N266);
nor NOR3 (N392, N383, N33, N292);
or OR4 (N393, N378, N390, N390, N92);
and AND4 (N394, N377, N230, N294, N385);
or OR2 (N395, N52, N320);
or OR4 (N396, N387, N306, N10, N204);
nor NOR3 (N397, N392, N51, N136);
nand NAND3 (N398, N395, N373, N256);
nor NOR2 (N399, N389, N172);
not NOT1 (N400, N381);
xor XOR2 (N401, N399, N82);
nand NAND4 (N402, N384, N111, N393, N226);
nor NOR4 (N403, N397, N252, N236, N151);
not NOT1 (N404, N236);
nor NOR4 (N405, N394, N248, N254, N397);
nand NAND3 (N406, N396, N365, N184);
or OR2 (N407, N405, N183);
buf BUF1 (N408, N402);
nor NOR3 (N409, N406, N169, N22);
nand NAND2 (N410, N408, N357);
and AND3 (N411, N401, N236, N212);
nor NOR3 (N412, N382, N65, N100);
or OR2 (N413, N404, N350);
nor NOR3 (N414, N400, N15, N156);
nor NOR3 (N415, N411, N90, N228);
or OR4 (N416, N410, N411, N182, N211);
not NOT1 (N417, N415);
buf BUF1 (N418, N391);
or OR4 (N419, N418, N355, N418, N262);
nand NAND4 (N420, N409, N59, N177, N137);
nand NAND3 (N421, N416, N378, N115);
not NOT1 (N422, N414);
and AND4 (N423, N398, N299, N291, N275);
nand NAND3 (N424, N403, N246, N6);
and AND2 (N425, N423, N279);
and AND3 (N426, N425, N24, N172);
not NOT1 (N427, N412);
nand NAND3 (N428, N427, N50, N33);
nor NOR4 (N429, N419, N335, N426, N388);
not NOT1 (N430, N190);
not NOT1 (N431, N421);
nor NOR4 (N432, N424, N164, N79, N25);
not NOT1 (N433, N413);
and AND3 (N434, N422, N72, N198);
nand NAND3 (N435, N407, N300, N434);
nor NOR4 (N436, N185, N48, N265, N316);
nor NOR2 (N437, N428, N428);
buf BUF1 (N438, N431);
or OR2 (N439, N435, N228);
buf BUF1 (N440, N430);
nand NAND3 (N441, N432, N17, N329);
not NOT1 (N442, N437);
xor XOR2 (N443, N438, N412);
and AND2 (N444, N433, N305);
nand NAND4 (N445, N436, N386, N392, N192);
not NOT1 (N446, N439);
not NOT1 (N447, N417);
nor NOR2 (N448, N444, N301);
xor XOR2 (N449, N441, N436);
or OR3 (N450, N448, N306, N70);
nand NAND2 (N451, N449, N146);
buf BUF1 (N452, N445);
xor XOR2 (N453, N446, N250);
and AND4 (N454, N429, N403, N94, N92);
or OR3 (N455, N450, N192, N287);
nand NAND4 (N456, N440, N310, N359, N123);
buf BUF1 (N457, N455);
xor XOR2 (N458, N442, N380);
not NOT1 (N459, N443);
nand NAND3 (N460, N447, N357, N116);
not NOT1 (N461, N456);
not NOT1 (N462, N454);
nand NAND3 (N463, N459, N316, N433);
buf BUF1 (N464, N462);
xor XOR2 (N465, N460, N115);
and AND4 (N466, N458, N463, N139, N121);
nor NOR2 (N467, N101, N462);
not NOT1 (N468, N461);
or OR2 (N469, N452, N272);
xor XOR2 (N470, N469, N457);
and AND2 (N471, N61, N60);
or OR3 (N472, N465, N458, N186);
and AND4 (N473, N471, N62, N262, N101);
or OR4 (N474, N453, N172, N302, N83);
nand NAND4 (N475, N451, N215, N375, N346);
or OR3 (N476, N474, N374, N183);
nor NOR3 (N477, N470, N133, N294);
or OR3 (N478, N475, N159, N365);
buf BUF1 (N479, N466);
and AND3 (N480, N473, N464, N8);
or OR4 (N481, N460, N26, N359, N22);
buf BUF1 (N482, N468);
not NOT1 (N483, N480);
buf BUF1 (N484, N467);
or OR3 (N485, N479, N275, N20);
not NOT1 (N486, N476);
nand NAND2 (N487, N420, N119);
or OR4 (N488, N482, N182, N149, N282);
nand NAND3 (N489, N478, N209, N153);
nand NAND3 (N490, N489, N117, N122);
buf BUF1 (N491, N490);
xor XOR2 (N492, N477, N434);
xor XOR2 (N493, N487, N423);
xor XOR2 (N494, N481, N372);
or OR4 (N495, N483, N117, N293, N353);
buf BUF1 (N496, N472);
not NOT1 (N497, N486);
nor NOR4 (N498, N493, N354, N407, N339);
buf BUF1 (N499, N497);
not NOT1 (N500, N488);
nor NOR2 (N501, N494, N495);
nor NOR2 (N502, N298, N346);
or OR3 (N503, N492, N99, N282);
xor XOR2 (N504, N502, N241);
or OR3 (N505, N501, N343, N220);
nor NOR2 (N506, N498, N97);
nor NOR4 (N507, N505, N458, N229, N417);
not NOT1 (N508, N504);
nand NAND4 (N509, N496, N409, N104, N418);
buf BUF1 (N510, N499);
not NOT1 (N511, N506);
xor XOR2 (N512, N500, N325);
or OR2 (N513, N509, N44);
nand NAND4 (N514, N503, N508, N395, N124);
buf BUF1 (N515, N470);
endmodule