// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N1601,N1617,N1613,N1607,N1612,N1615,N1610,N1608,N1616,N1618;

or OR4 (N19, N1, N16, N18, N16);
buf BUF1 (N20, N16);
and AND3 (N21, N3, N11, N17);
or OR3 (N22, N6, N7, N13);
nand NAND3 (N23, N8, N20, N20);
or OR3 (N24, N17, N8, N16);
and AND4 (N25, N21, N2, N20, N14);
nand NAND3 (N26, N17, N12, N5);
or OR4 (N27, N6, N17, N4, N7);
buf BUF1 (N28, N13);
buf BUF1 (N29, N9);
nor NOR4 (N30, N1, N2, N28, N2);
buf BUF1 (N31, N18);
and AND4 (N32, N29, N8, N21, N6);
nand NAND2 (N33, N24, N1);
buf BUF1 (N34, N25);
buf BUF1 (N35, N23);
nand NAND3 (N36, N27, N34, N8);
and AND4 (N37, N10, N13, N4, N10);
xor XOR2 (N38, N36, N32);
nand NAND4 (N39, N25, N32, N32, N10);
nand NAND4 (N40, N39, N33, N1, N26);
not NOT1 (N41, N6);
nand NAND2 (N42, N34, N29);
buf BUF1 (N43, N38);
nand NAND3 (N44, N41, N14, N6);
xor XOR2 (N45, N19, N23);
and AND4 (N46, N35, N28, N32, N1);
or OR4 (N47, N45, N35, N23, N8);
buf BUF1 (N48, N46);
nor NOR3 (N49, N48, N27, N46);
and AND3 (N50, N22, N6, N11);
or OR4 (N51, N43, N4, N33, N14);
and AND3 (N52, N47, N41, N10);
nand NAND2 (N53, N37, N28);
not NOT1 (N54, N40);
buf BUF1 (N55, N50);
buf BUF1 (N56, N53);
not NOT1 (N57, N55);
and AND3 (N58, N56, N12, N19);
buf BUF1 (N59, N31);
not NOT1 (N60, N51);
nand NAND2 (N61, N44, N38);
and AND3 (N62, N58, N25, N3);
nand NAND4 (N63, N49, N1, N49, N7);
and AND2 (N64, N57, N55);
and AND2 (N65, N63, N55);
and AND4 (N66, N52, N15, N40, N3);
nor NOR2 (N67, N42, N8);
not NOT1 (N68, N54);
xor XOR2 (N69, N61, N2);
nand NAND3 (N70, N59, N39, N66);
or OR3 (N71, N70, N38, N51);
or OR2 (N72, N51, N70);
not NOT1 (N73, N62);
buf BUF1 (N74, N67);
or OR3 (N75, N64, N25, N33);
or OR4 (N76, N71, N53, N41, N31);
xor XOR2 (N77, N30, N45);
xor XOR2 (N78, N76, N7);
not NOT1 (N79, N72);
nor NOR4 (N80, N68, N14, N58, N26);
buf BUF1 (N81, N78);
not NOT1 (N82, N73);
and AND3 (N83, N80, N11, N70);
nor NOR4 (N84, N77, N44, N42, N79);
xor XOR2 (N85, N39, N73);
nand NAND4 (N86, N69, N76, N59, N81);
or OR4 (N87, N9, N50, N56, N37);
and AND3 (N88, N85, N50, N50);
xor XOR2 (N89, N74, N1);
buf BUF1 (N90, N75);
nand NAND4 (N91, N65, N67, N7, N65);
not NOT1 (N92, N87);
or OR4 (N93, N60, N34, N84, N53);
nand NAND4 (N94, N41, N66, N5, N93);
nor NOR4 (N95, N39, N12, N48, N74);
nand NAND4 (N96, N94, N85, N57, N14);
buf BUF1 (N97, N86);
nand NAND3 (N98, N95, N22, N28);
or OR2 (N99, N97, N91);
or OR3 (N100, N48, N84, N78);
or OR4 (N101, N83, N80, N93, N90);
nand NAND3 (N102, N77, N1, N65);
buf BUF1 (N103, N98);
nand NAND3 (N104, N99, N80, N48);
nor NOR2 (N105, N103, N85);
nand NAND4 (N106, N102, N101, N31, N95);
xor XOR2 (N107, N31, N73);
buf BUF1 (N108, N88);
or OR3 (N109, N108, N83, N75);
and AND2 (N110, N92, N100);
or OR2 (N111, N101, N28);
and AND2 (N112, N107, N108);
or OR3 (N113, N109, N111, N106);
buf BUF1 (N114, N24);
or OR2 (N115, N47, N8);
buf BUF1 (N116, N112);
not NOT1 (N117, N110);
or OR2 (N118, N82, N33);
and AND3 (N119, N96, N13, N15);
xor XOR2 (N120, N89, N73);
or OR2 (N121, N119, N61);
xor XOR2 (N122, N104, N111);
or OR3 (N123, N122, N77, N53);
nor NOR2 (N124, N113, N4);
buf BUF1 (N125, N115);
xor XOR2 (N126, N118, N119);
and AND2 (N127, N116, N34);
nand NAND3 (N128, N120, N90, N120);
or OR4 (N129, N114, N124, N25, N75);
buf BUF1 (N130, N56);
nand NAND4 (N131, N129, N23, N52, N82);
nand NAND3 (N132, N121, N83, N21);
or OR3 (N133, N105, N18, N93);
buf BUF1 (N134, N125);
buf BUF1 (N135, N123);
nor NOR4 (N136, N133, N6, N54, N11);
buf BUF1 (N137, N135);
nor NOR4 (N138, N134, N115, N108, N7);
xor XOR2 (N139, N137, N86);
and AND3 (N140, N139, N130, N5);
buf BUF1 (N141, N15);
not NOT1 (N142, N140);
nor NOR2 (N143, N132, N62);
or OR3 (N144, N138, N133, N138);
and AND3 (N145, N131, N63, N3);
not NOT1 (N146, N128);
not NOT1 (N147, N142);
buf BUF1 (N148, N144);
buf BUF1 (N149, N143);
nor NOR3 (N150, N147, N73, N28);
nand NAND3 (N151, N146, N5, N85);
nor NOR4 (N152, N126, N126, N83, N1);
or OR4 (N153, N152, N64, N44, N74);
or OR3 (N154, N151, N36, N124);
nor NOR3 (N155, N150, N87, N117);
not NOT1 (N156, N65);
nand NAND2 (N157, N154, N20);
xor XOR2 (N158, N148, N78);
or OR3 (N159, N153, N150, N98);
buf BUF1 (N160, N157);
and AND2 (N161, N156, N15);
buf BUF1 (N162, N136);
and AND3 (N163, N127, N95, N52);
not NOT1 (N164, N145);
nand NAND4 (N165, N149, N44, N140, N4);
not NOT1 (N166, N155);
xor XOR2 (N167, N165, N113);
not NOT1 (N168, N163);
buf BUF1 (N169, N160);
buf BUF1 (N170, N169);
xor XOR2 (N171, N158, N94);
xor XOR2 (N172, N162, N138);
xor XOR2 (N173, N159, N95);
xor XOR2 (N174, N166, N5);
buf BUF1 (N175, N167);
nor NOR4 (N176, N141, N113, N138, N129);
buf BUF1 (N177, N168);
not NOT1 (N178, N164);
xor XOR2 (N179, N176, N103);
buf BUF1 (N180, N179);
nor NOR2 (N181, N174, N70);
nand NAND4 (N182, N175, N14, N51, N19);
xor XOR2 (N183, N178, N177);
not NOT1 (N184, N49);
nor NOR2 (N185, N170, N92);
nand NAND3 (N186, N183, N38, N183);
nand NAND3 (N187, N172, N72, N161);
not NOT1 (N188, N10);
or OR2 (N189, N185, N89);
nor NOR2 (N190, N181, N144);
not NOT1 (N191, N190);
not NOT1 (N192, N187);
buf BUF1 (N193, N186);
not NOT1 (N194, N193);
or OR4 (N195, N184, N22, N160, N175);
xor XOR2 (N196, N171, N94);
nand NAND4 (N197, N191, N162, N19, N176);
xor XOR2 (N198, N189, N24);
nand NAND4 (N199, N195, N34, N46, N10);
not NOT1 (N200, N182);
not NOT1 (N201, N194);
or OR3 (N202, N196, N159, N64);
xor XOR2 (N203, N199, N74);
buf BUF1 (N204, N192);
not NOT1 (N205, N180);
nand NAND2 (N206, N197, N10);
and AND2 (N207, N188, N52);
and AND4 (N208, N203, N196, N194, N46);
nand NAND2 (N209, N208, N4);
xor XOR2 (N210, N201, N59);
xor XOR2 (N211, N207, N6);
nand NAND4 (N212, N206, N49, N48, N2);
nor NOR3 (N213, N202, N88, N144);
nor NOR3 (N214, N212, N64, N202);
buf BUF1 (N215, N173);
not NOT1 (N216, N210);
xor XOR2 (N217, N204, N169);
xor XOR2 (N218, N198, N8);
buf BUF1 (N219, N218);
nor NOR4 (N220, N209, N187, N9, N214);
buf BUF1 (N221, N150);
xor XOR2 (N222, N216, N118);
xor XOR2 (N223, N211, N107);
or OR4 (N224, N205, N32, N219, N185);
nand NAND2 (N225, N39, N55);
and AND3 (N226, N213, N137, N217);
or OR4 (N227, N107, N102, N163, N140);
nor NOR2 (N228, N215, N180);
and AND3 (N229, N225, N163, N215);
buf BUF1 (N230, N200);
nand NAND2 (N231, N227, N24);
nor NOR3 (N232, N231, N177, N65);
xor XOR2 (N233, N221, N224);
buf BUF1 (N234, N84);
nor NOR3 (N235, N230, N143, N213);
buf BUF1 (N236, N228);
and AND2 (N237, N229, N23);
nor NOR4 (N238, N232, N151, N179, N210);
nor NOR2 (N239, N233, N41);
nand NAND3 (N240, N222, N172, N183);
nor NOR4 (N241, N235, N187, N83, N197);
and AND4 (N242, N234, N137, N183, N178);
and AND3 (N243, N237, N5, N102);
nor NOR4 (N244, N238, N63, N223, N23);
or OR2 (N245, N74, N219);
xor XOR2 (N246, N220, N81);
buf BUF1 (N247, N239);
and AND2 (N248, N243, N70);
and AND2 (N249, N240, N7);
or OR2 (N250, N242, N143);
buf BUF1 (N251, N249);
buf BUF1 (N252, N247);
xor XOR2 (N253, N244, N68);
buf BUF1 (N254, N226);
buf BUF1 (N255, N246);
or OR2 (N256, N250, N124);
and AND3 (N257, N248, N106, N184);
nand NAND4 (N258, N257, N249, N234, N18);
not NOT1 (N259, N254);
nand NAND4 (N260, N241, N243, N14, N247);
buf BUF1 (N261, N236);
nand NAND2 (N262, N251, N217);
buf BUF1 (N263, N262);
or OR4 (N264, N259, N245, N210, N255);
nand NAND3 (N265, N194, N163, N254);
xor XOR2 (N266, N145, N18);
nand NAND2 (N267, N266, N210);
and AND3 (N268, N264, N247, N136);
buf BUF1 (N269, N260);
nor NOR3 (N270, N253, N131, N102);
or OR4 (N271, N265, N65, N151, N30);
not NOT1 (N272, N267);
nor NOR4 (N273, N269, N58, N268, N156);
not NOT1 (N274, N154);
or OR2 (N275, N271, N24);
xor XOR2 (N276, N272, N147);
or OR3 (N277, N276, N121, N249);
nand NAND4 (N278, N263, N205, N135, N84);
xor XOR2 (N279, N273, N38);
nor NOR3 (N280, N275, N74, N60);
xor XOR2 (N281, N280, N59);
not NOT1 (N282, N261);
buf BUF1 (N283, N281);
xor XOR2 (N284, N278, N128);
buf BUF1 (N285, N274);
not NOT1 (N286, N270);
nor NOR2 (N287, N279, N52);
and AND2 (N288, N283, N82);
nor NOR3 (N289, N287, N47, N266);
not NOT1 (N290, N258);
nor NOR2 (N291, N252, N153);
not NOT1 (N292, N277);
nand NAND4 (N293, N285, N45, N217, N130);
and AND2 (N294, N291, N224);
or OR2 (N295, N292, N263);
or OR2 (N296, N284, N279);
xor XOR2 (N297, N293, N188);
xor XOR2 (N298, N282, N73);
and AND4 (N299, N298, N273, N28, N202);
nor NOR3 (N300, N297, N23, N235);
nand NAND3 (N301, N294, N216, N223);
not NOT1 (N302, N295);
nand NAND2 (N303, N299, N200);
and AND2 (N304, N290, N134);
nand NAND4 (N305, N286, N242, N84, N58);
and AND3 (N306, N296, N272, N27);
buf BUF1 (N307, N288);
nand NAND3 (N308, N302, N192, N265);
nor NOR3 (N309, N303, N293, N164);
not NOT1 (N310, N309);
not NOT1 (N311, N300);
and AND4 (N312, N301, N270, N63, N23);
buf BUF1 (N313, N307);
and AND3 (N314, N256, N253, N189);
not NOT1 (N315, N306);
buf BUF1 (N316, N310);
and AND4 (N317, N305, N217, N141, N141);
and AND4 (N318, N312, N73, N81, N289);
not NOT1 (N319, N203);
not NOT1 (N320, N315);
buf BUF1 (N321, N317);
or OR3 (N322, N316, N200, N178);
nand NAND4 (N323, N318, N223, N305, N319);
buf BUF1 (N324, N96);
xor XOR2 (N325, N322, N213);
xor XOR2 (N326, N324, N179);
or OR4 (N327, N326, N59, N163, N207);
xor XOR2 (N328, N314, N327);
not NOT1 (N329, N301);
buf BUF1 (N330, N323);
nor NOR3 (N331, N320, N130, N96);
nor NOR4 (N332, N325, N298, N127, N83);
xor XOR2 (N333, N329, N206);
xor XOR2 (N334, N304, N319);
nand NAND2 (N335, N333, N200);
not NOT1 (N336, N330);
not NOT1 (N337, N311);
and AND4 (N338, N308, N102, N71, N170);
or OR4 (N339, N321, N139, N118, N330);
nand NAND2 (N340, N331, N195);
or OR3 (N341, N339, N6, N266);
or OR3 (N342, N341, N151, N297);
or OR4 (N343, N334, N33, N217, N234);
nor NOR3 (N344, N336, N99, N92);
nor NOR2 (N345, N335, N168);
buf BUF1 (N346, N337);
nor NOR3 (N347, N346, N141, N285);
xor XOR2 (N348, N332, N134);
not NOT1 (N349, N328);
not NOT1 (N350, N349);
nor NOR3 (N351, N313, N235, N68);
not NOT1 (N352, N345);
or OR2 (N353, N342, N225);
xor XOR2 (N354, N340, N268);
nor NOR2 (N355, N351, N26);
nand NAND2 (N356, N338, N144);
buf BUF1 (N357, N354);
and AND3 (N358, N343, N315, N108);
xor XOR2 (N359, N357, N278);
nand NAND2 (N360, N352, N245);
or OR4 (N361, N348, N107, N237, N319);
nand NAND3 (N362, N353, N310, N52);
nand NAND2 (N363, N350, N31);
nor NOR4 (N364, N363, N129, N115, N296);
and AND3 (N365, N356, N226, N276);
nand NAND4 (N366, N362, N48, N341, N358);
or OR2 (N367, N204, N22);
xor XOR2 (N368, N360, N355);
buf BUF1 (N369, N260);
not NOT1 (N370, N365);
and AND3 (N371, N368, N257, N273);
and AND3 (N372, N371, N6, N20);
xor XOR2 (N373, N347, N5);
xor XOR2 (N374, N359, N17);
not NOT1 (N375, N344);
not NOT1 (N376, N373);
or OR3 (N377, N367, N217, N146);
and AND2 (N378, N366, N113);
or OR4 (N379, N376, N305, N317, N276);
nand NAND2 (N380, N361, N162);
not NOT1 (N381, N377);
or OR3 (N382, N372, N279, N7);
not NOT1 (N383, N380);
nand NAND4 (N384, N379, N138, N289, N94);
buf BUF1 (N385, N378);
and AND3 (N386, N381, N205, N170);
buf BUF1 (N387, N384);
not NOT1 (N388, N385);
nand NAND4 (N389, N370, N7, N113, N141);
or OR4 (N390, N387, N156, N22, N220);
nor NOR2 (N391, N390, N230);
or OR4 (N392, N388, N226, N334, N361);
nor NOR4 (N393, N392, N367, N82, N228);
buf BUF1 (N394, N374);
not NOT1 (N395, N382);
not NOT1 (N396, N364);
xor XOR2 (N397, N386, N16);
nand NAND4 (N398, N395, N330, N34, N238);
xor XOR2 (N399, N383, N12);
nand NAND2 (N400, N375, N94);
not NOT1 (N401, N398);
nor NOR4 (N402, N389, N224, N317, N120);
not NOT1 (N403, N396);
not NOT1 (N404, N397);
and AND2 (N405, N369, N285);
or OR3 (N406, N401, N345, N341);
nor NOR2 (N407, N394, N149);
nor NOR2 (N408, N406, N127);
and AND3 (N409, N402, N18, N322);
and AND2 (N410, N404, N398);
nand NAND4 (N411, N393, N69, N59, N315);
buf BUF1 (N412, N408);
or OR3 (N413, N410, N246, N213);
nand NAND2 (N414, N411, N135);
or OR2 (N415, N414, N189);
buf BUF1 (N416, N391);
xor XOR2 (N417, N416, N38);
or OR2 (N418, N407, N332);
buf BUF1 (N419, N413);
or OR2 (N420, N400, N272);
nor NOR2 (N421, N420, N312);
or OR4 (N422, N409, N368, N413, N51);
not NOT1 (N423, N417);
buf BUF1 (N424, N423);
or OR4 (N425, N419, N106, N278, N294);
buf BUF1 (N426, N421);
nor NOR4 (N427, N399, N206, N310, N186);
nand NAND4 (N428, N426, N215, N104, N42);
and AND2 (N429, N428, N146);
or OR3 (N430, N412, N413, N202);
not NOT1 (N431, N430);
or OR2 (N432, N424, N169);
buf BUF1 (N433, N432);
or OR3 (N434, N429, N39, N155);
or OR2 (N435, N422, N227);
and AND3 (N436, N433, N346, N58);
not NOT1 (N437, N434);
and AND3 (N438, N418, N81, N312);
and AND2 (N439, N403, N218);
not NOT1 (N440, N431);
or OR2 (N441, N439, N410);
not NOT1 (N442, N435);
buf BUF1 (N443, N437);
buf BUF1 (N444, N436);
buf BUF1 (N445, N442);
xor XOR2 (N446, N438, N9);
and AND4 (N447, N443, N355, N230, N316);
or OR3 (N448, N444, N44, N203);
nor NOR3 (N449, N446, N311, N293);
xor XOR2 (N450, N440, N239);
and AND3 (N451, N445, N293, N186);
xor XOR2 (N452, N449, N195);
or OR2 (N453, N451, N297);
nand NAND4 (N454, N427, N371, N382, N189);
and AND3 (N455, N448, N366, N426);
xor XOR2 (N456, N450, N296);
or OR2 (N457, N456, N151);
nor NOR2 (N458, N447, N220);
xor XOR2 (N459, N425, N14);
nor NOR4 (N460, N459, N108, N43, N221);
not NOT1 (N461, N458);
not NOT1 (N462, N457);
not NOT1 (N463, N461);
buf BUF1 (N464, N415);
not NOT1 (N465, N455);
buf BUF1 (N466, N452);
xor XOR2 (N467, N405, N48);
nand NAND3 (N468, N465, N112, N248);
and AND3 (N469, N468, N394, N250);
xor XOR2 (N470, N464, N76);
not NOT1 (N471, N470);
buf BUF1 (N472, N471);
not NOT1 (N473, N441);
buf BUF1 (N474, N454);
buf BUF1 (N475, N473);
buf BUF1 (N476, N467);
nand NAND4 (N477, N475, N310, N144, N227);
or OR4 (N478, N460, N409, N160, N266);
nor NOR3 (N479, N476, N252, N219);
not NOT1 (N480, N474);
and AND2 (N481, N472, N235);
xor XOR2 (N482, N466, N351);
not NOT1 (N483, N453);
nand NAND2 (N484, N469, N467);
not NOT1 (N485, N481);
and AND4 (N486, N478, N113, N99, N278);
nand NAND4 (N487, N484, N418, N69, N112);
nor NOR4 (N488, N483, N121, N241, N157);
not NOT1 (N489, N477);
and AND2 (N490, N462, N233);
and AND4 (N491, N485, N6, N34, N404);
and AND2 (N492, N479, N458);
not NOT1 (N493, N491);
or OR3 (N494, N488, N284, N297);
nor NOR2 (N495, N490, N424);
buf BUF1 (N496, N480);
not NOT1 (N497, N487);
buf BUF1 (N498, N489);
and AND2 (N499, N486, N74);
buf BUF1 (N500, N492);
and AND3 (N501, N496, N210, N446);
and AND3 (N502, N501, N192, N46);
buf BUF1 (N503, N497);
xor XOR2 (N504, N495, N185);
nand NAND2 (N505, N503, N10);
nand NAND4 (N506, N463, N495, N298, N122);
or OR4 (N507, N505, N198, N131, N29);
nor NOR4 (N508, N482, N26, N201, N284);
and AND2 (N509, N499, N329);
and AND2 (N510, N502, N43);
not NOT1 (N511, N504);
or OR3 (N512, N494, N508, N125);
or OR3 (N513, N51, N424, N360);
xor XOR2 (N514, N498, N431);
or OR2 (N515, N511, N402);
and AND2 (N516, N515, N478);
not NOT1 (N517, N507);
nor NOR4 (N518, N506, N171, N234, N267);
nand NAND4 (N519, N509, N347, N275, N216);
or OR3 (N520, N519, N482, N83);
xor XOR2 (N521, N520, N134);
nand NAND3 (N522, N512, N257, N429);
and AND4 (N523, N493, N363, N183, N88);
xor XOR2 (N524, N514, N284);
and AND4 (N525, N510, N359, N257, N204);
or OR4 (N526, N516, N292, N159, N143);
buf BUF1 (N527, N500);
not NOT1 (N528, N527);
xor XOR2 (N529, N522, N506);
and AND3 (N530, N529, N371, N73);
nand NAND4 (N531, N526, N58, N251, N464);
or OR3 (N532, N530, N80, N327);
nand NAND2 (N533, N528, N329);
nor NOR4 (N534, N517, N522, N191, N135);
not NOT1 (N535, N533);
xor XOR2 (N536, N524, N235);
nand NAND4 (N537, N521, N329, N479, N317);
buf BUF1 (N538, N535);
nor NOR2 (N539, N532, N306);
nand NAND2 (N540, N525, N36);
xor XOR2 (N541, N534, N22);
xor XOR2 (N542, N523, N420);
nand NAND2 (N543, N542, N288);
and AND3 (N544, N543, N1, N534);
xor XOR2 (N545, N518, N18);
buf BUF1 (N546, N537);
and AND2 (N547, N536, N102);
buf BUF1 (N548, N541);
nand NAND4 (N549, N548, N325, N105, N99);
xor XOR2 (N550, N545, N351);
nand NAND2 (N551, N539, N429);
nor NOR3 (N552, N538, N520, N104);
xor XOR2 (N553, N547, N278);
nand NAND2 (N554, N550, N293);
nand NAND2 (N555, N551, N513);
and AND4 (N556, N212, N38, N257, N404);
nand NAND3 (N557, N531, N90, N271);
and AND4 (N558, N540, N434, N445, N94);
not NOT1 (N559, N552);
nor NOR3 (N560, N559, N541, N478);
not NOT1 (N561, N558);
xor XOR2 (N562, N549, N502);
not NOT1 (N563, N555);
and AND4 (N564, N553, N109, N181, N361);
and AND2 (N565, N556, N240);
or OR2 (N566, N565, N98);
nand NAND3 (N567, N564, N308, N80);
and AND4 (N568, N560, N52, N192, N558);
xor XOR2 (N569, N567, N494);
xor XOR2 (N570, N566, N176);
buf BUF1 (N571, N544);
or OR3 (N572, N568, N387, N84);
or OR2 (N573, N570, N41);
and AND3 (N574, N573, N38, N324);
nor NOR2 (N575, N571, N276);
or OR4 (N576, N575, N324, N300, N144);
not NOT1 (N577, N569);
or OR3 (N578, N574, N27, N227);
and AND2 (N579, N557, N319);
buf BUF1 (N580, N563);
xor XOR2 (N581, N579, N293);
nand NAND2 (N582, N578, N350);
nand NAND4 (N583, N576, N404, N195, N267);
nor NOR3 (N584, N546, N337, N308);
and AND4 (N585, N572, N345, N273, N265);
buf BUF1 (N586, N581);
and AND2 (N587, N586, N526);
or OR2 (N588, N561, N16);
xor XOR2 (N589, N580, N288);
xor XOR2 (N590, N588, N374);
or OR3 (N591, N585, N404, N236);
buf BUF1 (N592, N582);
not NOT1 (N593, N590);
buf BUF1 (N594, N587);
or OR2 (N595, N594, N3);
nor NOR4 (N596, N584, N76, N591, N588);
or OR2 (N597, N281, N234);
not NOT1 (N598, N583);
buf BUF1 (N599, N554);
nand NAND2 (N600, N596, N39);
nor NOR3 (N601, N592, N460, N349);
and AND3 (N602, N593, N128, N367);
nor NOR2 (N603, N598, N77);
and AND3 (N604, N602, N57, N108);
xor XOR2 (N605, N589, N168);
not NOT1 (N606, N600);
not NOT1 (N607, N597);
and AND2 (N608, N606, N441);
not NOT1 (N609, N604);
not NOT1 (N610, N577);
not NOT1 (N611, N562);
nand NAND3 (N612, N610, N364, N512);
buf BUF1 (N613, N605);
nand NAND4 (N614, N612, N114, N46, N608);
buf BUF1 (N615, N519);
xor XOR2 (N616, N613, N374);
nor NOR2 (N617, N603, N140);
xor XOR2 (N618, N609, N158);
nand NAND3 (N619, N595, N517, N31);
not NOT1 (N620, N611);
xor XOR2 (N621, N618, N217);
and AND3 (N622, N601, N2, N485);
nor NOR2 (N623, N616, N300);
or OR2 (N624, N617, N335);
nor NOR2 (N625, N599, N27);
xor XOR2 (N626, N621, N498);
xor XOR2 (N627, N622, N193);
not NOT1 (N628, N627);
buf BUF1 (N629, N615);
and AND4 (N630, N614, N99, N155, N86);
xor XOR2 (N631, N623, N142);
nor NOR2 (N632, N630, N2);
nor NOR2 (N633, N624, N505);
and AND4 (N634, N628, N498, N463, N120);
nor NOR2 (N635, N619, N91);
and AND2 (N636, N634, N490);
not NOT1 (N637, N636);
not NOT1 (N638, N631);
and AND4 (N639, N629, N520, N517, N491);
nand NAND4 (N640, N637, N638, N139, N106);
and AND2 (N641, N504, N533);
nor NOR4 (N642, N626, N240, N190, N453);
nor NOR2 (N643, N635, N455);
buf BUF1 (N644, N607);
not NOT1 (N645, N633);
xor XOR2 (N646, N640, N473);
xor XOR2 (N647, N620, N640);
buf BUF1 (N648, N642);
not NOT1 (N649, N625);
not NOT1 (N650, N646);
or OR2 (N651, N650, N543);
and AND2 (N652, N651, N108);
or OR3 (N653, N641, N333, N308);
and AND2 (N654, N644, N246);
or OR2 (N655, N653, N152);
nand NAND4 (N656, N648, N438, N17, N510);
xor XOR2 (N657, N647, N54);
or OR2 (N658, N655, N132);
nor NOR3 (N659, N649, N289, N128);
nand NAND2 (N660, N643, N86);
and AND3 (N661, N652, N520, N250);
nor NOR2 (N662, N659, N9);
nand NAND2 (N663, N658, N80);
and AND2 (N664, N663, N642);
not NOT1 (N665, N645);
or OR4 (N666, N662, N388, N397, N273);
xor XOR2 (N667, N639, N648);
or OR4 (N668, N665, N562, N475, N311);
xor XOR2 (N669, N664, N498);
or OR4 (N670, N667, N163, N290, N603);
buf BUF1 (N671, N660);
nand NAND4 (N672, N671, N585, N454, N319);
and AND2 (N673, N672, N669);
not NOT1 (N674, N2);
nand NAND4 (N675, N632, N66, N664, N13);
and AND2 (N676, N666, N503);
xor XOR2 (N677, N654, N392);
nor NOR3 (N678, N656, N446, N435);
and AND4 (N679, N674, N646, N646, N463);
nand NAND4 (N680, N679, N633, N325, N561);
nand NAND3 (N681, N668, N416, N52);
and AND3 (N682, N681, N568, N315);
and AND4 (N683, N676, N454, N361, N598);
not NOT1 (N684, N677);
or OR3 (N685, N657, N669, N229);
buf BUF1 (N686, N678);
nor NOR4 (N687, N685, N600, N326, N173);
buf BUF1 (N688, N684);
or OR2 (N689, N673, N63);
not NOT1 (N690, N689);
or OR4 (N691, N661, N538, N103, N365);
buf BUF1 (N692, N680);
not NOT1 (N693, N692);
not NOT1 (N694, N690);
nand NAND4 (N695, N691, N298, N28, N629);
and AND2 (N696, N683, N408);
and AND3 (N697, N670, N271, N125);
nand NAND4 (N698, N688, N609, N25, N511);
nor NOR2 (N699, N694, N693);
and AND3 (N700, N573, N369, N632);
nor NOR4 (N701, N686, N53, N667, N265);
xor XOR2 (N702, N697, N603);
not NOT1 (N703, N699);
nor NOR2 (N704, N703, N68);
nor NOR3 (N705, N700, N266, N75);
buf BUF1 (N706, N687);
buf BUF1 (N707, N701);
nand NAND2 (N708, N706, N587);
xor XOR2 (N709, N675, N589);
not NOT1 (N710, N704);
buf BUF1 (N711, N702);
and AND2 (N712, N708, N87);
xor XOR2 (N713, N696, N116);
nand NAND4 (N714, N698, N486, N162, N635);
nor NOR4 (N715, N682, N400, N211, N39);
xor XOR2 (N716, N705, N359);
nand NAND4 (N717, N712, N681, N601, N712);
and AND3 (N718, N709, N455, N156);
xor XOR2 (N719, N714, N275);
xor XOR2 (N720, N715, N154);
xor XOR2 (N721, N717, N680);
buf BUF1 (N722, N720);
nor NOR4 (N723, N707, N245, N585, N630);
or OR4 (N724, N716, N710, N30, N404);
xor XOR2 (N725, N366, N661);
nor NOR3 (N726, N721, N613, N723);
xor XOR2 (N727, N152, N171);
and AND3 (N728, N725, N410, N377);
xor XOR2 (N729, N728, N443);
and AND4 (N730, N718, N241, N376, N656);
and AND4 (N731, N726, N579, N585, N223);
xor XOR2 (N732, N730, N67);
nand NAND2 (N733, N724, N247);
not NOT1 (N734, N729);
or OR4 (N735, N719, N168, N124, N731);
nand NAND3 (N736, N559, N286, N637);
and AND2 (N737, N727, N385);
buf BUF1 (N738, N736);
and AND3 (N739, N722, N350, N495);
not NOT1 (N740, N735);
not NOT1 (N741, N737);
and AND3 (N742, N713, N720, N687);
xor XOR2 (N743, N711, N81);
or OR2 (N744, N742, N32);
and AND2 (N745, N744, N736);
not NOT1 (N746, N745);
buf BUF1 (N747, N738);
or OR2 (N748, N732, N57);
not NOT1 (N749, N695);
buf BUF1 (N750, N748);
not NOT1 (N751, N743);
nand NAND4 (N752, N751, N289, N435, N625);
xor XOR2 (N753, N747, N614);
buf BUF1 (N754, N734);
xor XOR2 (N755, N749, N309);
not NOT1 (N756, N755);
and AND3 (N757, N733, N518, N639);
nand NAND2 (N758, N750, N480);
or OR2 (N759, N753, N645);
and AND3 (N760, N752, N549, N146);
or OR2 (N761, N756, N250);
nor NOR2 (N762, N760, N542);
buf BUF1 (N763, N739);
or OR3 (N764, N759, N456, N594);
nor NOR3 (N765, N762, N74, N124);
buf BUF1 (N766, N741);
xor XOR2 (N767, N758, N412);
buf BUF1 (N768, N764);
not NOT1 (N769, N754);
xor XOR2 (N770, N740, N316);
nand NAND4 (N771, N765, N549, N726, N317);
nand NAND3 (N772, N769, N732, N613);
nor NOR4 (N773, N763, N575, N766, N459);
buf BUF1 (N774, N275);
nor NOR4 (N775, N746, N765, N406, N491);
buf BUF1 (N776, N770);
buf BUF1 (N777, N773);
nand NAND2 (N778, N757, N155);
and AND3 (N779, N771, N375, N206);
buf BUF1 (N780, N779);
and AND3 (N781, N761, N288, N330);
and AND2 (N782, N774, N738);
nand NAND2 (N783, N775, N87);
nor NOR3 (N784, N783, N124, N245);
xor XOR2 (N785, N784, N39);
buf BUF1 (N786, N768);
buf BUF1 (N787, N785);
not NOT1 (N788, N782);
nor NOR4 (N789, N777, N183, N625, N336);
xor XOR2 (N790, N780, N175);
not NOT1 (N791, N788);
buf BUF1 (N792, N791);
or OR3 (N793, N792, N687, N68);
xor XOR2 (N794, N787, N169);
nand NAND4 (N795, N781, N537, N55, N317);
nor NOR3 (N796, N790, N75, N658);
buf BUF1 (N797, N776);
xor XOR2 (N798, N797, N27);
or OR4 (N799, N772, N715, N651, N633);
buf BUF1 (N800, N786);
xor XOR2 (N801, N793, N13);
nand NAND4 (N802, N799, N601, N59, N73);
buf BUF1 (N803, N778);
nor NOR3 (N804, N794, N16, N375);
and AND2 (N805, N796, N349);
not NOT1 (N806, N800);
nand NAND2 (N807, N798, N225);
buf BUF1 (N808, N801);
buf BUF1 (N809, N802);
not NOT1 (N810, N805);
or OR4 (N811, N795, N773, N744, N687);
xor XOR2 (N812, N804, N574);
nor NOR3 (N813, N809, N131, N726);
nor NOR3 (N814, N767, N744, N574);
nor NOR4 (N815, N806, N595, N753, N8);
xor XOR2 (N816, N808, N575);
and AND3 (N817, N810, N414, N645);
not NOT1 (N818, N817);
nand NAND2 (N819, N816, N103);
buf BUF1 (N820, N807);
and AND3 (N821, N811, N623, N501);
xor XOR2 (N822, N789, N419);
nor NOR2 (N823, N821, N557);
xor XOR2 (N824, N820, N241);
buf BUF1 (N825, N812);
xor XOR2 (N826, N825, N76);
xor XOR2 (N827, N826, N372);
not NOT1 (N828, N822);
or OR2 (N829, N803, N338);
nor NOR4 (N830, N829, N333, N255, N353);
nor NOR4 (N831, N828, N125, N101, N11);
xor XOR2 (N832, N814, N304);
or OR3 (N833, N818, N182, N576);
not NOT1 (N834, N823);
nand NAND4 (N835, N830, N415, N386, N606);
and AND4 (N836, N819, N467, N693, N189);
or OR2 (N837, N831, N8);
nor NOR2 (N838, N813, N733);
or OR2 (N839, N824, N116);
nor NOR4 (N840, N833, N809, N73, N784);
nand NAND3 (N841, N827, N157, N207);
or OR4 (N842, N834, N266, N740, N388);
or OR2 (N843, N838, N718);
and AND2 (N844, N839, N410);
and AND2 (N845, N815, N706);
nor NOR2 (N846, N841, N678);
and AND2 (N847, N845, N296);
nor NOR2 (N848, N842, N436);
and AND4 (N849, N844, N347, N197, N298);
and AND4 (N850, N849, N274, N113, N361);
or OR2 (N851, N848, N329);
or OR3 (N852, N843, N505, N527);
xor XOR2 (N853, N851, N238);
or OR3 (N854, N837, N331, N139);
and AND4 (N855, N846, N848, N292, N480);
or OR2 (N856, N847, N5);
buf BUF1 (N857, N853);
not NOT1 (N858, N835);
and AND4 (N859, N840, N837, N600, N853);
xor XOR2 (N860, N854, N397);
buf BUF1 (N861, N855);
not NOT1 (N862, N836);
not NOT1 (N863, N860);
nand NAND4 (N864, N856, N527, N243, N412);
or OR2 (N865, N862, N13);
and AND2 (N866, N864, N580);
not NOT1 (N867, N852);
buf BUF1 (N868, N863);
buf BUF1 (N869, N850);
or OR4 (N870, N861, N301, N539, N315);
xor XOR2 (N871, N865, N106);
buf BUF1 (N872, N866);
xor XOR2 (N873, N832, N226);
and AND3 (N874, N872, N569, N460);
not NOT1 (N875, N869);
or OR3 (N876, N857, N711, N177);
nor NOR3 (N877, N867, N96, N22);
or OR2 (N878, N870, N680);
and AND3 (N879, N871, N658, N75);
buf BUF1 (N880, N876);
nor NOR2 (N881, N868, N241);
xor XOR2 (N882, N874, N567);
nor NOR4 (N883, N877, N95, N206, N138);
buf BUF1 (N884, N879);
nand NAND4 (N885, N878, N284, N399, N658);
or OR4 (N886, N875, N443, N24, N387);
nand NAND4 (N887, N859, N511, N76, N177);
and AND2 (N888, N884, N637);
xor XOR2 (N889, N886, N672);
nor NOR3 (N890, N889, N5, N67);
and AND4 (N891, N858, N503, N149, N491);
xor XOR2 (N892, N887, N544);
nor NOR4 (N893, N891, N457, N760, N833);
buf BUF1 (N894, N883);
buf BUF1 (N895, N894);
buf BUF1 (N896, N885);
nor NOR2 (N897, N896, N118);
and AND3 (N898, N895, N631, N34);
and AND2 (N899, N880, N313);
nand NAND4 (N900, N893, N59, N157, N129);
nor NOR2 (N901, N890, N313);
xor XOR2 (N902, N892, N136);
xor XOR2 (N903, N881, N613);
nand NAND3 (N904, N902, N758, N510);
and AND4 (N905, N900, N245, N321, N816);
or OR3 (N906, N901, N652, N626);
nor NOR2 (N907, N903, N260);
nand NAND3 (N908, N904, N132, N769);
nor NOR4 (N909, N898, N614, N82, N614);
and AND2 (N910, N899, N377);
or OR4 (N911, N882, N379, N156, N190);
and AND4 (N912, N911, N216, N766, N288);
buf BUF1 (N913, N873);
or OR4 (N914, N906, N105, N194, N537);
buf BUF1 (N915, N914);
xor XOR2 (N916, N908, N894);
nor NOR3 (N917, N913, N372, N820);
nand NAND2 (N918, N909, N242);
not NOT1 (N919, N888);
nand NAND3 (N920, N919, N887, N737);
xor XOR2 (N921, N905, N827);
buf BUF1 (N922, N915);
not NOT1 (N923, N897);
nor NOR2 (N924, N912, N654);
or OR2 (N925, N917, N751);
buf BUF1 (N926, N924);
not NOT1 (N927, N916);
nor NOR4 (N928, N920, N621, N699, N385);
nand NAND2 (N929, N928, N672);
not NOT1 (N930, N927);
buf BUF1 (N931, N926);
or OR4 (N932, N910, N159, N713, N893);
and AND4 (N933, N918, N613, N399, N226);
not NOT1 (N934, N922);
buf BUF1 (N935, N930);
nand NAND2 (N936, N933, N248);
or OR2 (N937, N935, N348);
not NOT1 (N938, N907);
buf BUF1 (N939, N929);
or OR2 (N940, N932, N24);
nor NOR4 (N941, N923, N599, N656, N700);
not NOT1 (N942, N934);
buf BUF1 (N943, N937);
or OR4 (N944, N938, N521, N482, N603);
and AND3 (N945, N941, N763, N370);
xor XOR2 (N946, N925, N231);
buf BUF1 (N947, N945);
not NOT1 (N948, N942);
not NOT1 (N949, N946);
not NOT1 (N950, N921);
nor NOR3 (N951, N947, N255, N548);
nor NOR2 (N952, N940, N637);
or OR2 (N953, N950, N254);
nand NAND4 (N954, N939, N256, N371, N372);
buf BUF1 (N955, N953);
and AND3 (N956, N954, N652, N20);
nand NAND2 (N957, N948, N553);
not NOT1 (N958, N955);
or OR3 (N959, N936, N506, N41);
and AND2 (N960, N959, N793);
nor NOR2 (N961, N952, N910);
nand NAND3 (N962, N931, N765, N400);
xor XOR2 (N963, N951, N266);
nor NOR2 (N964, N949, N665);
or OR4 (N965, N943, N387, N781, N807);
xor XOR2 (N966, N965, N493);
or OR3 (N967, N958, N192, N737);
not NOT1 (N968, N962);
not NOT1 (N969, N957);
nand NAND2 (N970, N969, N188);
nand NAND2 (N971, N944, N61);
not NOT1 (N972, N971);
nand NAND4 (N973, N960, N760, N81, N951);
nand NAND2 (N974, N963, N492);
and AND3 (N975, N967, N712, N241);
xor XOR2 (N976, N956, N108);
not NOT1 (N977, N966);
buf BUF1 (N978, N968);
nor NOR3 (N979, N976, N166, N601);
xor XOR2 (N980, N973, N558);
nand NAND4 (N981, N977, N421, N745, N450);
not NOT1 (N982, N979);
buf BUF1 (N983, N981);
buf BUF1 (N984, N974);
or OR2 (N985, N964, N118);
nand NAND4 (N986, N984, N454, N95, N973);
and AND2 (N987, N986, N885);
and AND3 (N988, N982, N386, N321);
nor NOR3 (N989, N978, N739, N667);
and AND3 (N990, N961, N436, N907);
not NOT1 (N991, N988);
or OR3 (N992, N987, N619, N863);
xor XOR2 (N993, N989, N928);
nand NAND2 (N994, N972, N189);
not NOT1 (N995, N994);
nor NOR3 (N996, N975, N878, N356);
xor XOR2 (N997, N991, N755);
xor XOR2 (N998, N993, N190);
nand NAND2 (N999, N998, N657);
nand NAND2 (N1000, N995, N399);
and AND4 (N1001, N1000, N407, N682, N937);
nor NOR3 (N1002, N990, N245, N819);
nor NOR4 (N1003, N1001, N759, N785, N751);
or OR2 (N1004, N996, N571);
buf BUF1 (N1005, N985);
or OR3 (N1006, N1004, N984, N636);
nor NOR3 (N1007, N1002, N354, N951);
nand NAND4 (N1008, N980, N521, N201, N652);
xor XOR2 (N1009, N997, N378);
or OR4 (N1010, N1003, N330, N906, N222);
nor NOR3 (N1011, N970, N348, N537);
nor NOR3 (N1012, N1005, N908, N856);
nand NAND4 (N1013, N1012, N987, N699, N82);
buf BUF1 (N1014, N1010);
buf BUF1 (N1015, N1006);
xor XOR2 (N1016, N1007, N217);
buf BUF1 (N1017, N983);
xor XOR2 (N1018, N999, N311);
buf BUF1 (N1019, N1014);
not NOT1 (N1020, N1018);
and AND2 (N1021, N1019, N867);
nor NOR4 (N1022, N1009, N920, N635, N40);
buf BUF1 (N1023, N1008);
buf BUF1 (N1024, N1016);
nand NAND3 (N1025, N1013, N121, N656);
nand NAND2 (N1026, N1011, N468);
xor XOR2 (N1027, N1023, N912);
buf BUF1 (N1028, N1021);
nor NOR3 (N1029, N1024, N488, N73);
or OR3 (N1030, N1025, N936, N443);
nor NOR4 (N1031, N1020, N3, N930, N835);
and AND4 (N1032, N1017, N203, N639, N572);
nor NOR3 (N1033, N1026, N866, N426);
nor NOR2 (N1034, N1030, N15);
nor NOR4 (N1035, N1028, N75, N693, N1006);
xor XOR2 (N1036, N1035, N786);
or OR2 (N1037, N1027, N74);
nor NOR3 (N1038, N992, N755, N955);
xor XOR2 (N1039, N1037, N108);
xor XOR2 (N1040, N1032, N684);
xor XOR2 (N1041, N1036, N140);
xor XOR2 (N1042, N1031, N358);
and AND4 (N1043, N1015, N38, N87, N146);
buf BUF1 (N1044, N1029);
not NOT1 (N1045, N1034);
not NOT1 (N1046, N1039);
nand NAND4 (N1047, N1042, N261, N981, N636);
nand NAND4 (N1048, N1033, N34, N384, N1002);
and AND4 (N1049, N1045, N683, N992, N901);
not NOT1 (N1050, N1047);
or OR2 (N1051, N1043, N958);
and AND3 (N1052, N1038, N1050, N103);
nand NAND3 (N1053, N600, N595, N381);
and AND2 (N1054, N1049, N622);
and AND4 (N1055, N1041, N704, N583, N868);
or OR2 (N1056, N1055, N292);
or OR3 (N1057, N1022, N513, N73);
xor XOR2 (N1058, N1053, N687);
and AND3 (N1059, N1057, N698, N118);
xor XOR2 (N1060, N1044, N274);
and AND4 (N1061, N1058, N831, N106, N259);
buf BUF1 (N1062, N1046);
xor XOR2 (N1063, N1056, N408);
not NOT1 (N1064, N1048);
xor XOR2 (N1065, N1061, N100);
or OR2 (N1066, N1060, N508);
or OR2 (N1067, N1065, N217);
nor NOR3 (N1068, N1040, N794, N373);
and AND4 (N1069, N1052, N906, N896, N635);
nor NOR3 (N1070, N1064, N814, N315);
buf BUF1 (N1071, N1070);
or OR4 (N1072, N1062, N24, N754, N1001);
xor XOR2 (N1073, N1069, N178);
and AND4 (N1074, N1063, N1058, N865, N128);
nor NOR4 (N1075, N1068, N334, N743, N827);
xor XOR2 (N1076, N1054, N158);
nor NOR2 (N1077, N1075, N1030);
buf BUF1 (N1078, N1076);
not NOT1 (N1079, N1077);
or OR3 (N1080, N1071, N562, N13);
nand NAND3 (N1081, N1080, N963, N892);
xor XOR2 (N1082, N1079, N996);
nand NAND2 (N1083, N1081, N969);
nand NAND2 (N1084, N1078, N436);
not NOT1 (N1085, N1073);
buf BUF1 (N1086, N1082);
nor NOR4 (N1087, N1059, N268, N759, N129);
nor NOR2 (N1088, N1051, N129);
nor NOR2 (N1089, N1074, N74);
buf BUF1 (N1090, N1067);
and AND3 (N1091, N1086, N450, N365);
buf BUF1 (N1092, N1085);
buf BUF1 (N1093, N1091);
nand NAND3 (N1094, N1088, N437, N187);
not NOT1 (N1095, N1083);
not NOT1 (N1096, N1084);
not NOT1 (N1097, N1094);
xor XOR2 (N1098, N1092, N272);
buf BUF1 (N1099, N1093);
xor XOR2 (N1100, N1089, N917);
or OR4 (N1101, N1097, N668, N1076, N1056);
and AND2 (N1102, N1099, N148);
nand NAND3 (N1103, N1090, N474, N143);
and AND2 (N1104, N1102, N565);
nor NOR4 (N1105, N1104, N818, N976, N811);
nand NAND2 (N1106, N1087, N1029);
nor NOR4 (N1107, N1066, N681, N996, N905);
or OR2 (N1108, N1095, N1094);
or OR3 (N1109, N1072, N477, N977);
and AND2 (N1110, N1096, N1093);
not NOT1 (N1111, N1105);
nor NOR4 (N1112, N1098, N280, N954, N1075);
xor XOR2 (N1113, N1107, N361);
not NOT1 (N1114, N1111);
nand NAND4 (N1115, N1108, N331, N32, N1096);
nor NOR4 (N1116, N1114, N458, N703, N786);
and AND2 (N1117, N1106, N504);
and AND2 (N1118, N1100, N309);
buf BUF1 (N1119, N1110);
not NOT1 (N1120, N1116);
nor NOR3 (N1121, N1120, N207, N873);
or OR2 (N1122, N1118, N490);
nand NAND2 (N1123, N1112, N989);
or OR2 (N1124, N1122, N7);
buf BUF1 (N1125, N1124);
buf BUF1 (N1126, N1103);
xor XOR2 (N1127, N1121, N637);
buf BUF1 (N1128, N1127);
nand NAND3 (N1129, N1109, N1081, N139);
nand NAND3 (N1130, N1115, N103, N622);
and AND2 (N1131, N1125, N28);
xor XOR2 (N1132, N1129, N213);
or OR3 (N1133, N1126, N856, N692);
not NOT1 (N1134, N1113);
nor NOR4 (N1135, N1131, N696, N496, N584);
buf BUF1 (N1136, N1132);
buf BUF1 (N1137, N1134);
not NOT1 (N1138, N1137);
and AND4 (N1139, N1138, N1061, N167, N626);
not NOT1 (N1140, N1117);
nor NOR2 (N1141, N1119, N100);
and AND4 (N1142, N1123, N55, N476, N505);
nand NAND3 (N1143, N1133, N95, N581);
nor NOR4 (N1144, N1136, N133, N209, N1051);
not NOT1 (N1145, N1140);
and AND3 (N1146, N1130, N989, N898);
buf BUF1 (N1147, N1128);
nor NOR2 (N1148, N1135, N830);
buf BUF1 (N1149, N1142);
or OR3 (N1150, N1145, N2, N189);
xor XOR2 (N1151, N1148, N294);
nand NAND3 (N1152, N1141, N462, N846);
xor XOR2 (N1153, N1143, N1080);
not NOT1 (N1154, N1144);
nand NAND4 (N1155, N1139, N166, N297, N444);
buf BUF1 (N1156, N1152);
or OR2 (N1157, N1153, N760);
xor XOR2 (N1158, N1146, N218);
xor XOR2 (N1159, N1156, N620);
or OR2 (N1160, N1155, N431);
not NOT1 (N1161, N1150);
nor NOR2 (N1162, N1147, N168);
and AND2 (N1163, N1158, N392);
not NOT1 (N1164, N1161);
buf BUF1 (N1165, N1101);
nand NAND4 (N1166, N1162, N209, N16, N321);
or OR2 (N1167, N1160, N1097);
xor XOR2 (N1168, N1164, N514);
or OR4 (N1169, N1163, N203, N1050, N507);
nor NOR2 (N1170, N1165, N301);
buf BUF1 (N1171, N1151);
or OR3 (N1172, N1166, N748, N1070);
nor NOR2 (N1173, N1149, N700);
not NOT1 (N1174, N1159);
and AND2 (N1175, N1167, N369);
xor XOR2 (N1176, N1170, N160);
or OR2 (N1177, N1168, N105);
nand NAND4 (N1178, N1174, N1141, N992, N554);
and AND3 (N1179, N1169, N167, N925);
and AND2 (N1180, N1154, N867);
nand NAND3 (N1181, N1180, N1150, N344);
not NOT1 (N1182, N1175);
not NOT1 (N1183, N1176);
xor XOR2 (N1184, N1178, N134);
buf BUF1 (N1185, N1179);
nand NAND3 (N1186, N1183, N953, N986);
nor NOR3 (N1187, N1182, N178, N303);
and AND3 (N1188, N1186, N1066, N205);
nor NOR3 (N1189, N1173, N1055, N746);
nand NAND4 (N1190, N1187, N473, N434, N85);
not NOT1 (N1191, N1189);
not NOT1 (N1192, N1185);
not NOT1 (N1193, N1184);
buf BUF1 (N1194, N1177);
buf BUF1 (N1195, N1194);
buf BUF1 (N1196, N1190);
or OR2 (N1197, N1157, N69);
and AND4 (N1198, N1192, N561, N600, N1023);
nor NOR3 (N1199, N1198, N373, N136);
or OR4 (N1200, N1196, N570, N1146, N18);
buf BUF1 (N1201, N1172);
nor NOR3 (N1202, N1191, N813, N1151);
nand NAND2 (N1203, N1188, N421);
buf BUF1 (N1204, N1193);
or OR2 (N1205, N1201, N674);
nand NAND2 (N1206, N1200, N431);
not NOT1 (N1207, N1181);
or OR3 (N1208, N1207, N1014, N944);
not NOT1 (N1209, N1195);
and AND3 (N1210, N1203, N871, N210);
xor XOR2 (N1211, N1209, N997);
xor XOR2 (N1212, N1171, N892);
buf BUF1 (N1213, N1204);
and AND3 (N1214, N1212, N811, N652);
xor XOR2 (N1215, N1202, N931);
nand NAND3 (N1216, N1199, N462, N1077);
not NOT1 (N1217, N1208);
xor XOR2 (N1218, N1215, N1048);
or OR3 (N1219, N1205, N1041, N1096);
nand NAND4 (N1220, N1217, N375, N420, N899);
nand NAND4 (N1221, N1210, N519, N160, N106);
buf BUF1 (N1222, N1218);
xor XOR2 (N1223, N1220, N152);
buf BUF1 (N1224, N1219);
or OR2 (N1225, N1214, N1170);
and AND2 (N1226, N1222, N183);
nand NAND3 (N1227, N1221, N724, N59);
or OR2 (N1228, N1223, N558);
or OR3 (N1229, N1213, N1016, N265);
nor NOR2 (N1230, N1227, N106);
nor NOR4 (N1231, N1225, N809, N126, N197);
buf BUF1 (N1232, N1216);
nor NOR3 (N1233, N1224, N554, N551);
and AND3 (N1234, N1211, N1118, N593);
nand NAND4 (N1235, N1226, N935, N384, N704);
not NOT1 (N1236, N1197);
nor NOR4 (N1237, N1236, N1167, N1065, N514);
and AND2 (N1238, N1235, N405);
and AND4 (N1239, N1238, N889, N966, N57);
not NOT1 (N1240, N1232);
nand NAND4 (N1241, N1239, N1176, N657, N572);
and AND3 (N1242, N1229, N1086, N806);
buf BUF1 (N1243, N1241);
not NOT1 (N1244, N1230);
nor NOR3 (N1245, N1233, N37, N968);
nand NAND2 (N1246, N1237, N178);
buf BUF1 (N1247, N1243);
and AND3 (N1248, N1231, N1032, N290);
buf BUF1 (N1249, N1245);
buf BUF1 (N1250, N1234);
or OR2 (N1251, N1206, N644);
xor XOR2 (N1252, N1250, N1069);
or OR3 (N1253, N1249, N992, N976);
nand NAND4 (N1254, N1252, N78, N615, N209);
or OR3 (N1255, N1251, N176, N79);
buf BUF1 (N1256, N1253);
nand NAND3 (N1257, N1255, N694, N1058);
nand NAND3 (N1258, N1246, N253, N238);
or OR4 (N1259, N1258, N790, N1021, N636);
not NOT1 (N1260, N1254);
nand NAND2 (N1261, N1242, N902);
nand NAND2 (N1262, N1228, N887);
xor XOR2 (N1263, N1244, N333);
and AND2 (N1264, N1263, N608);
buf BUF1 (N1265, N1259);
nor NOR4 (N1266, N1256, N562, N62, N1036);
buf BUF1 (N1267, N1247);
buf BUF1 (N1268, N1240);
not NOT1 (N1269, N1267);
or OR3 (N1270, N1248, N146, N558);
or OR3 (N1271, N1265, N264, N1105);
and AND3 (N1272, N1262, N111, N1099);
or OR2 (N1273, N1272, N483);
buf BUF1 (N1274, N1266);
nor NOR4 (N1275, N1269, N231, N157, N446);
and AND4 (N1276, N1257, N909, N223, N177);
xor XOR2 (N1277, N1268, N918);
or OR3 (N1278, N1264, N911, N1052);
nor NOR2 (N1279, N1271, N1110);
buf BUF1 (N1280, N1278);
xor XOR2 (N1281, N1280, N149);
or OR4 (N1282, N1260, N392, N1256, N356);
xor XOR2 (N1283, N1281, N1039);
nor NOR3 (N1284, N1261, N1188, N185);
xor XOR2 (N1285, N1277, N1095);
not NOT1 (N1286, N1284);
not NOT1 (N1287, N1274);
buf BUF1 (N1288, N1270);
nand NAND3 (N1289, N1273, N521, N1203);
and AND2 (N1290, N1286, N603);
and AND4 (N1291, N1276, N1180, N1027, N314);
not NOT1 (N1292, N1282);
nor NOR3 (N1293, N1287, N1002, N1211);
buf BUF1 (N1294, N1288);
buf BUF1 (N1295, N1293);
or OR4 (N1296, N1275, N850, N901, N815);
nor NOR2 (N1297, N1292, N355);
nor NOR3 (N1298, N1289, N979, N793);
nor NOR4 (N1299, N1295, N1038, N609, N228);
not NOT1 (N1300, N1290);
nor NOR4 (N1301, N1283, N737, N542, N1263);
not NOT1 (N1302, N1285);
xor XOR2 (N1303, N1279, N767);
nor NOR4 (N1304, N1303, N1245, N563, N290);
nand NAND4 (N1305, N1296, N1217, N125, N1093);
buf BUF1 (N1306, N1301);
and AND4 (N1307, N1291, N95, N1081, N890);
nand NAND3 (N1308, N1294, N606, N898);
xor XOR2 (N1309, N1306, N828);
or OR3 (N1310, N1297, N1164, N1294);
xor XOR2 (N1311, N1299, N726);
and AND2 (N1312, N1309, N1208);
and AND4 (N1313, N1302, N21, N458, N17);
and AND3 (N1314, N1310, N652, N741);
nor NOR3 (N1315, N1304, N165, N290);
not NOT1 (N1316, N1314);
buf BUF1 (N1317, N1300);
or OR2 (N1318, N1308, N331);
xor XOR2 (N1319, N1311, N938);
buf BUF1 (N1320, N1316);
and AND2 (N1321, N1320, N368);
nor NOR2 (N1322, N1298, N1103);
not NOT1 (N1323, N1307);
nor NOR3 (N1324, N1321, N1053, N1250);
xor XOR2 (N1325, N1324, N120);
and AND2 (N1326, N1322, N424);
or OR3 (N1327, N1315, N812, N72);
not NOT1 (N1328, N1326);
nor NOR3 (N1329, N1319, N542, N480);
or OR4 (N1330, N1317, N185, N935, N1314);
or OR4 (N1331, N1328, N599, N634, N282);
nor NOR3 (N1332, N1305, N811, N670);
nor NOR3 (N1333, N1332, N829, N921);
buf BUF1 (N1334, N1330);
nand NAND4 (N1335, N1318, N1041, N898, N777);
not NOT1 (N1336, N1325);
or OR4 (N1337, N1313, N73, N872, N342);
xor XOR2 (N1338, N1336, N336);
not NOT1 (N1339, N1329);
nand NAND2 (N1340, N1339, N553);
xor XOR2 (N1341, N1334, N972);
not NOT1 (N1342, N1327);
buf BUF1 (N1343, N1331);
and AND3 (N1344, N1333, N618, N108);
or OR2 (N1345, N1340, N442);
nand NAND4 (N1346, N1323, N527, N805, N130);
or OR2 (N1347, N1337, N898);
nand NAND3 (N1348, N1347, N1189, N644);
or OR3 (N1349, N1348, N104, N1071);
or OR2 (N1350, N1344, N1250);
or OR3 (N1351, N1335, N471, N1002);
nor NOR3 (N1352, N1345, N861, N882);
nand NAND2 (N1353, N1341, N804);
nand NAND2 (N1354, N1343, N1295);
xor XOR2 (N1355, N1351, N270);
buf BUF1 (N1356, N1342);
not NOT1 (N1357, N1346);
not NOT1 (N1358, N1354);
and AND3 (N1359, N1338, N941, N503);
nor NOR4 (N1360, N1359, N684, N402, N1197);
nor NOR2 (N1361, N1356, N683);
xor XOR2 (N1362, N1358, N466);
buf BUF1 (N1363, N1362);
not NOT1 (N1364, N1355);
buf BUF1 (N1365, N1312);
xor XOR2 (N1366, N1363, N1235);
nor NOR3 (N1367, N1352, N44, N921);
nand NAND3 (N1368, N1365, N1208, N715);
xor XOR2 (N1369, N1350, N1018);
not NOT1 (N1370, N1357);
nor NOR2 (N1371, N1364, N925);
xor XOR2 (N1372, N1369, N1172);
nor NOR4 (N1373, N1368, N75, N430, N574);
not NOT1 (N1374, N1372);
not NOT1 (N1375, N1374);
nor NOR4 (N1376, N1360, N46, N494, N1148);
buf BUF1 (N1377, N1371);
and AND4 (N1378, N1377, N620, N93, N981);
and AND2 (N1379, N1378, N580);
nand NAND4 (N1380, N1379, N800, N406, N79);
and AND4 (N1381, N1353, N725, N116, N243);
xor XOR2 (N1382, N1370, N508);
not NOT1 (N1383, N1380);
or OR4 (N1384, N1381, N936, N1031, N1045);
and AND4 (N1385, N1366, N499, N49, N951);
xor XOR2 (N1386, N1376, N975);
nand NAND2 (N1387, N1367, N44);
nor NOR3 (N1388, N1382, N567, N1074);
or OR3 (N1389, N1375, N1076, N642);
or OR3 (N1390, N1383, N396, N68);
or OR2 (N1391, N1385, N648);
not NOT1 (N1392, N1384);
and AND3 (N1393, N1361, N41, N1014);
buf BUF1 (N1394, N1389);
nand NAND2 (N1395, N1394, N414);
xor XOR2 (N1396, N1349, N898);
xor XOR2 (N1397, N1373, N291);
and AND2 (N1398, N1396, N1379);
nor NOR4 (N1399, N1391, N945, N873, N576);
and AND3 (N1400, N1386, N523, N361);
buf BUF1 (N1401, N1398);
buf BUF1 (N1402, N1399);
not NOT1 (N1403, N1397);
nand NAND3 (N1404, N1400, N262, N1100);
nor NOR3 (N1405, N1388, N492, N198);
nor NOR3 (N1406, N1403, N579, N1051);
buf BUF1 (N1407, N1406);
or OR4 (N1408, N1387, N981, N723, N607);
not NOT1 (N1409, N1405);
buf BUF1 (N1410, N1409);
not NOT1 (N1411, N1390);
nand NAND3 (N1412, N1393, N1260, N91);
nand NAND4 (N1413, N1407, N113, N107, N1406);
or OR2 (N1414, N1411, N700);
or OR3 (N1415, N1408, N374, N963);
not NOT1 (N1416, N1401);
and AND2 (N1417, N1414, N1235);
xor XOR2 (N1418, N1417, N1233);
and AND4 (N1419, N1416, N259, N1321, N370);
and AND2 (N1420, N1402, N1240);
buf BUF1 (N1421, N1404);
or OR4 (N1422, N1413, N121, N1217, N1185);
not NOT1 (N1423, N1418);
xor XOR2 (N1424, N1410, N1069);
or OR4 (N1425, N1423, N348, N1219, N187);
nor NOR4 (N1426, N1420, N592, N186, N286);
nor NOR2 (N1427, N1412, N1321);
or OR4 (N1428, N1426, N933, N516, N847);
buf BUF1 (N1429, N1422);
xor XOR2 (N1430, N1424, N1274);
and AND4 (N1431, N1395, N191, N981, N385);
nor NOR2 (N1432, N1425, N1082);
xor XOR2 (N1433, N1392, N106);
and AND3 (N1434, N1429, N891, N608);
and AND4 (N1435, N1430, N894, N501, N991);
and AND4 (N1436, N1433, N77, N1007, N474);
not NOT1 (N1437, N1435);
buf BUF1 (N1438, N1427);
nor NOR4 (N1439, N1432, N566, N1223, N769);
or OR3 (N1440, N1437, N395, N463);
nand NAND2 (N1441, N1431, N118);
xor XOR2 (N1442, N1419, N292);
not NOT1 (N1443, N1428);
xor XOR2 (N1444, N1421, N842);
buf BUF1 (N1445, N1439);
xor XOR2 (N1446, N1441, N89);
buf BUF1 (N1447, N1444);
xor XOR2 (N1448, N1442, N408);
buf BUF1 (N1449, N1415);
not NOT1 (N1450, N1436);
buf BUF1 (N1451, N1438);
or OR2 (N1452, N1446, N219);
or OR3 (N1453, N1434, N385, N574);
xor XOR2 (N1454, N1445, N1367);
and AND2 (N1455, N1453, N1101);
nor NOR3 (N1456, N1449, N754, N1101);
not NOT1 (N1457, N1454);
xor XOR2 (N1458, N1440, N898);
nor NOR4 (N1459, N1443, N196, N125, N1374);
and AND4 (N1460, N1456, N919, N970, N578);
nand NAND2 (N1461, N1452, N72);
xor XOR2 (N1462, N1457, N1317);
not NOT1 (N1463, N1455);
or OR4 (N1464, N1447, N939, N393, N621);
nand NAND2 (N1465, N1459, N308);
xor XOR2 (N1466, N1460, N469);
or OR4 (N1467, N1464, N1248, N5, N716);
xor XOR2 (N1468, N1450, N737);
or OR2 (N1469, N1451, N1332);
nor NOR2 (N1470, N1448, N536);
and AND2 (N1471, N1469, N431);
xor XOR2 (N1472, N1463, N264);
buf BUF1 (N1473, N1468);
buf BUF1 (N1474, N1458);
xor XOR2 (N1475, N1466, N584);
xor XOR2 (N1476, N1462, N67);
nor NOR4 (N1477, N1474, N1418, N722, N537);
nand NAND3 (N1478, N1461, N774, N1453);
nor NOR2 (N1479, N1467, N959);
or OR2 (N1480, N1476, N284);
nand NAND3 (N1481, N1480, N1461, N1031);
nor NOR4 (N1482, N1478, N19, N947, N1474);
or OR3 (N1483, N1481, N689, N1051);
and AND2 (N1484, N1470, N1451);
buf BUF1 (N1485, N1479);
nand NAND3 (N1486, N1485, N433, N465);
or OR4 (N1487, N1486, N955, N163, N436);
not NOT1 (N1488, N1472);
buf BUF1 (N1489, N1488);
nor NOR2 (N1490, N1482, N829);
buf BUF1 (N1491, N1490);
xor XOR2 (N1492, N1471, N640);
or OR3 (N1493, N1484, N904, N1396);
xor XOR2 (N1494, N1465, N258);
or OR3 (N1495, N1477, N1280, N66);
and AND2 (N1496, N1483, N239);
buf BUF1 (N1497, N1489);
or OR4 (N1498, N1496, N761, N633, N327);
or OR4 (N1499, N1493, N550, N1395, N210);
xor XOR2 (N1500, N1497, N1457);
xor XOR2 (N1501, N1473, N1000);
or OR3 (N1502, N1487, N256, N1013);
xor XOR2 (N1503, N1492, N842);
or OR3 (N1504, N1499, N600, N1468);
or OR3 (N1505, N1498, N1430, N443);
not NOT1 (N1506, N1475);
buf BUF1 (N1507, N1503);
or OR2 (N1508, N1501, N256);
or OR2 (N1509, N1507, N14);
nand NAND2 (N1510, N1505, N802);
not NOT1 (N1511, N1510);
nor NOR3 (N1512, N1506, N1082, N427);
nand NAND3 (N1513, N1511, N1370, N1374);
nand NAND2 (N1514, N1500, N863);
nor NOR3 (N1515, N1508, N1021, N688);
xor XOR2 (N1516, N1512, N1290);
and AND4 (N1517, N1516, N129, N836, N752);
not NOT1 (N1518, N1517);
or OR2 (N1519, N1491, N424);
not NOT1 (N1520, N1518);
and AND3 (N1521, N1515, N205, N1398);
not NOT1 (N1522, N1504);
and AND3 (N1523, N1520, N1392, N335);
xor XOR2 (N1524, N1494, N1512);
xor XOR2 (N1525, N1495, N841);
nand NAND4 (N1526, N1509, N686, N1507, N1446);
nand NAND3 (N1527, N1522, N1284, N628);
not NOT1 (N1528, N1527);
nor NOR2 (N1529, N1524, N1517);
nand NAND4 (N1530, N1513, N71, N581, N1305);
nor NOR3 (N1531, N1519, N1344, N1331);
xor XOR2 (N1532, N1514, N763);
buf BUF1 (N1533, N1502);
nand NAND3 (N1534, N1525, N132, N265);
buf BUF1 (N1535, N1528);
nor NOR3 (N1536, N1523, N1267, N93);
nand NAND4 (N1537, N1532, N1496, N1490, N457);
xor XOR2 (N1538, N1537, N1489);
not NOT1 (N1539, N1521);
nor NOR2 (N1540, N1526, N305);
or OR2 (N1541, N1539, N139);
xor XOR2 (N1542, N1540, N182);
and AND4 (N1543, N1542, N202, N800, N1198);
nor NOR3 (N1544, N1531, N445, N1227);
nor NOR4 (N1545, N1541, N1090, N654, N158);
or OR4 (N1546, N1536, N919, N657, N971);
and AND3 (N1547, N1544, N955, N1068);
nor NOR3 (N1548, N1543, N1398, N351);
or OR2 (N1549, N1538, N842);
not NOT1 (N1550, N1545);
and AND2 (N1551, N1546, N82);
buf BUF1 (N1552, N1548);
buf BUF1 (N1553, N1550);
or OR3 (N1554, N1547, N145, N537);
nand NAND4 (N1555, N1530, N729, N1422, N370);
nand NAND3 (N1556, N1552, N789, N1062);
buf BUF1 (N1557, N1533);
nor NOR4 (N1558, N1534, N352, N1525, N886);
nor NOR4 (N1559, N1556, N701, N553, N1410);
not NOT1 (N1560, N1558);
or OR3 (N1561, N1560, N310, N797);
xor XOR2 (N1562, N1529, N892);
xor XOR2 (N1563, N1549, N1127);
or OR2 (N1564, N1555, N429);
and AND2 (N1565, N1562, N238);
xor XOR2 (N1566, N1557, N1021);
nand NAND4 (N1567, N1554, N725, N975, N769);
xor XOR2 (N1568, N1535, N911);
xor XOR2 (N1569, N1559, N1175);
or OR3 (N1570, N1551, N1262, N816);
not NOT1 (N1571, N1565);
or OR4 (N1572, N1570, N433, N323, N1085);
nand NAND4 (N1573, N1561, N556, N130, N295);
or OR2 (N1574, N1564, N1185);
or OR2 (N1575, N1569, N461);
xor XOR2 (N1576, N1567, N536);
nand NAND3 (N1577, N1553, N134, N481);
xor XOR2 (N1578, N1576, N1387);
nor NOR4 (N1579, N1578, N900, N1294, N82);
nand NAND2 (N1580, N1571, N1019);
xor XOR2 (N1581, N1575, N940);
or OR3 (N1582, N1566, N68, N1533);
and AND3 (N1583, N1580, N588, N435);
nor NOR4 (N1584, N1583, N1181, N33, N366);
and AND2 (N1585, N1573, N206);
xor XOR2 (N1586, N1585, N866);
nand NAND4 (N1587, N1563, N779, N412, N1145);
buf BUF1 (N1588, N1577);
nand NAND2 (N1589, N1581, N1418);
or OR2 (N1590, N1588, N1290);
not NOT1 (N1591, N1587);
xor XOR2 (N1592, N1568, N1500);
buf BUF1 (N1593, N1591);
not NOT1 (N1594, N1572);
nor NOR2 (N1595, N1584, N1016);
or OR3 (N1596, N1589, N314, N1543);
and AND3 (N1597, N1579, N477, N232);
or OR3 (N1598, N1593, N686, N704);
and AND2 (N1599, N1598, N479);
buf BUF1 (N1600, N1595);
not NOT1 (N1601, N1599);
not NOT1 (N1602, N1597);
not NOT1 (N1603, N1592);
xor XOR2 (N1604, N1586, N1007);
xor XOR2 (N1605, N1603, N800);
and AND3 (N1606, N1596, N1211, N227);
nand NAND3 (N1607, N1606, N1155, N1457);
nand NAND4 (N1608, N1582, N474, N586, N1005);
buf BUF1 (N1609, N1600);
and AND4 (N1610, N1594, N1461, N389, N1581);
not NOT1 (N1611, N1605);
xor XOR2 (N1612, N1590, N345);
and AND2 (N1613, N1609, N1542);
and AND3 (N1614, N1602, N60, N1229);
not NOT1 (N1615, N1574);
buf BUF1 (N1616, N1614);
and AND2 (N1617, N1604, N1286);
and AND2 (N1618, N1611, N265);
endmodule