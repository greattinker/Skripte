// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N6398,N6410,N6416,N6413,N6409,N6407,N6395,N6404,N6414,N6417;

nand NAND3 (N18, N12, N3, N12);
xor XOR2 (N19, N8, N2);
nand NAND3 (N20, N15, N4, N4);
xor XOR2 (N21, N17, N2);
or OR3 (N22, N12, N15, N12);
nor NOR4 (N23, N6, N13, N5, N11);
nor NOR4 (N24, N19, N11, N12, N18);
or OR2 (N25, N23, N4);
buf BUF1 (N26, N25);
or OR4 (N27, N25, N26, N5, N4);
buf BUF1 (N28, N10);
buf BUF1 (N29, N17);
nand NAND3 (N30, N7, N3, N8);
nor NOR4 (N31, N28, N2, N25, N4);
nor NOR2 (N32, N29, N24);
not NOT1 (N33, N15);
nand NAND3 (N34, N25, N3, N22);
xor XOR2 (N35, N5, N28);
buf BUF1 (N36, N34);
xor XOR2 (N37, N4, N36);
nor NOR3 (N38, N16, N22, N31);
nand NAND2 (N39, N30, N6);
or OR2 (N40, N9, N20);
or OR3 (N41, N19, N36, N40);
buf BUF1 (N42, N39);
nand NAND3 (N43, N29, N37, N4);
not NOT1 (N44, N19);
nand NAND3 (N45, N33, N41, N16);
or OR2 (N46, N42, N28);
buf BUF1 (N47, N24);
buf BUF1 (N48, N21);
not NOT1 (N49, N43);
and AND3 (N50, N38, N30, N23);
not NOT1 (N51, N46);
not NOT1 (N52, N32);
nand NAND3 (N53, N47, N11, N36);
nand NAND4 (N54, N48, N50, N49, N13);
xor XOR2 (N55, N38, N39);
xor XOR2 (N56, N46, N11);
nor NOR4 (N57, N53, N22, N38, N16);
and AND4 (N58, N35, N44, N4, N55);
or OR3 (N59, N23, N53, N41);
or OR3 (N60, N49, N36, N25);
xor XOR2 (N61, N57, N5);
nor NOR2 (N62, N56, N19);
or OR3 (N63, N54, N22, N33);
nand NAND4 (N64, N52, N51, N35, N36);
or OR4 (N65, N25, N40, N34, N58);
nor NOR4 (N66, N53, N3, N28, N62);
not NOT1 (N67, N37);
and AND3 (N68, N65, N9, N8);
not NOT1 (N69, N68);
nand NAND4 (N70, N64, N46, N5, N47);
xor XOR2 (N71, N60, N65);
nand NAND2 (N72, N67, N20);
or OR2 (N73, N72, N12);
not NOT1 (N74, N66);
xor XOR2 (N75, N70, N32);
xor XOR2 (N76, N71, N26);
nand NAND4 (N77, N76, N27, N41, N53);
or OR4 (N78, N58, N57, N69, N52);
or OR2 (N79, N40, N19);
and AND2 (N80, N63, N48);
and AND3 (N81, N74, N14, N42);
and AND4 (N82, N75, N15, N78, N54);
buf BUF1 (N83, N24);
nand NAND3 (N84, N61, N62, N2);
nor NOR4 (N85, N77, N9, N32, N5);
and AND3 (N86, N79, N78, N11);
or OR3 (N87, N82, N80, N32);
nor NOR4 (N88, N44, N18, N64, N1);
and AND4 (N89, N86, N26, N85, N41);
xor XOR2 (N90, N89, N51);
and AND2 (N91, N77, N75);
and AND4 (N92, N88, N53, N41, N3);
xor XOR2 (N93, N59, N90);
not NOT1 (N94, N13);
nand NAND2 (N95, N73, N42);
not NOT1 (N96, N84);
buf BUF1 (N97, N45);
or OR2 (N98, N87, N15);
buf BUF1 (N99, N81);
xor XOR2 (N100, N93, N74);
and AND2 (N101, N91, N94);
and AND3 (N102, N101, N74, N39);
nand NAND3 (N103, N56, N58, N13);
xor XOR2 (N104, N103, N31);
and AND3 (N105, N102, N11, N25);
and AND4 (N106, N105, N37, N100, N99);
buf BUF1 (N107, N50);
not NOT1 (N108, N39);
nor NOR4 (N109, N92, N48, N101, N13);
nand NAND2 (N110, N95, N41);
xor XOR2 (N111, N107, N95);
nor NOR2 (N112, N109, N68);
buf BUF1 (N113, N83);
not NOT1 (N114, N97);
or OR2 (N115, N111, N89);
and AND4 (N116, N108, N41, N107, N56);
xor XOR2 (N117, N110, N4);
and AND2 (N118, N98, N60);
nor NOR2 (N119, N106, N20);
nor NOR2 (N120, N118, N30);
or OR4 (N121, N114, N115, N113, N112);
buf BUF1 (N122, N84);
and AND2 (N123, N22, N32);
xor XOR2 (N124, N25, N78);
buf BUF1 (N125, N117);
buf BUF1 (N126, N123);
not NOT1 (N127, N116);
xor XOR2 (N128, N125, N25);
xor XOR2 (N129, N104, N65);
nor NOR4 (N130, N129, N35, N57, N105);
or OR3 (N131, N130, N36, N72);
nand NAND4 (N132, N120, N39, N77, N92);
buf BUF1 (N133, N119);
or OR3 (N134, N127, N97, N105);
buf BUF1 (N135, N124);
and AND2 (N136, N128, N90);
nand NAND3 (N137, N134, N128, N124);
nor NOR3 (N138, N133, N41, N52);
and AND4 (N139, N135, N23, N112, N6);
and AND2 (N140, N131, N101);
xor XOR2 (N141, N132, N97);
and AND2 (N142, N141, N62);
nor NOR2 (N143, N140, N141);
not NOT1 (N144, N143);
not NOT1 (N145, N126);
and AND2 (N146, N145, N126);
xor XOR2 (N147, N137, N69);
nor NOR3 (N148, N146, N52, N76);
or OR4 (N149, N96, N87, N40, N88);
or OR3 (N150, N122, N116, N70);
buf BUF1 (N151, N142);
xor XOR2 (N152, N121, N3);
nor NOR2 (N153, N152, N30);
xor XOR2 (N154, N138, N10);
or OR3 (N155, N149, N60, N5);
xor XOR2 (N156, N148, N103);
nand NAND2 (N157, N151, N132);
buf BUF1 (N158, N156);
or OR3 (N159, N155, N151, N16);
and AND4 (N160, N159, N138, N26, N69);
nand NAND4 (N161, N158, N140, N24, N147);
and AND3 (N162, N106, N57, N154);
not NOT1 (N163, N146);
not NOT1 (N164, N139);
or OR3 (N165, N136, N117, N66);
and AND4 (N166, N144, N58, N76, N82);
xor XOR2 (N167, N161, N47);
and AND3 (N168, N153, N152, N128);
xor XOR2 (N169, N157, N84);
and AND2 (N170, N165, N97);
nor NOR2 (N171, N170, N75);
or OR3 (N172, N169, N53, N107);
nand NAND4 (N173, N172, N56, N85, N30);
nor NOR3 (N174, N160, N103, N116);
nand NAND4 (N175, N174, N69, N78, N172);
or OR4 (N176, N167, N78, N83, N165);
nor NOR2 (N177, N171, N101);
xor XOR2 (N178, N164, N62);
or OR2 (N179, N173, N81);
nor NOR2 (N180, N150, N74);
nand NAND3 (N181, N166, N82, N36);
and AND4 (N182, N176, N175, N66, N138);
or OR3 (N183, N177, N182, N141);
or OR3 (N184, N43, N143, N166);
and AND2 (N185, N24, N17);
nor NOR2 (N186, N168, N54);
nand NAND3 (N187, N183, N57, N50);
buf BUF1 (N188, N184);
or OR2 (N189, N163, N98);
nand NAND2 (N190, N180, N37);
or OR2 (N191, N188, N60);
or OR2 (N192, N189, N71);
or OR2 (N193, N181, N132);
or OR3 (N194, N187, N16, N42);
buf BUF1 (N195, N186);
xor XOR2 (N196, N195, N46);
not NOT1 (N197, N178);
not NOT1 (N198, N185);
nor NOR2 (N199, N193, N75);
buf BUF1 (N200, N191);
buf BUF1 (N201, N198);
nor NOR3 (N202, N162, N157, N116);
or OR2 (N203, N199, N110);
and AND3 (N204, N197, N38, N104);
nand NAND3 (N205, N179, N85, N53);
buf BUF1 (N206, N192);
not NOT1 (N207, N203);
nand NAND4 (N208, N190, N164, N54, N12);
nor NOR4 (N209, N206, N32, N171, N189);
buf BUF1 (N210, N202);
xor XOR2 (N211, N208, N4);
not NOT1 (N212, N205);
or OR2 (N213, N201, N71);
not NOT1 (N214, N204);
not NOT1 (N215, N213);
buf BUF1 (N216, N212);
xor XOR2 (N217, N196, N172);
nand NAND2 (N218, N214, N143);
or OR4 (N219, N215, N149, N16, N198);
nor NOR4 (N220, N200, N141, N21, N113);
not NOT1 (N221, N209);
not NOT1 (N222, N211);
buf BUF1 (N223, N221);
nand NAND3 (N224, N218, N151, N126);
and AND3 (N225, N210, N107, N7);
nand NAND2 (N226, N224, N223);
or OR4 (N227, N225, N181, N58, N178);
not NOT1 (N228, N29);
nand NAND3 (N229, N228, N8, N92);
buf BUF1 (N230, N217);
or OR2 (N231, N220, N112);
nor NOR4 (N232, N219, N112, N52, N77);
not NOT1 (N233, N222);
and AND3 (N234, N207, N210, N147);
or OR3 (N235, N194, N101, N166);
xor XOR2 (N236, N227, N118);
xor XOR2 (N237, N236, N89);
buf BUF1 (N238, N232);
xor XOR2 (N239, N230, N155);
and AND4 (N240, N234, N96, N33, N190);
and AND2 (N241, N239, N215);
or OR4 (N242, N240, N54, N67, N98);
buf BUF1 (N243, N231);
not NOT1 (N244, N237);
nand NAND3 (N245, N241, N84, N215);
nand NAND4 (N246, N216, N113, N58, N46);
or OR3 (N247, N246, N59, N99);
nand NAND4 (N248, N247, N18, N148, N30);
nand NAND3 (N249, N245, N192, N241);
and AND3 (N250, N226, N168, N41);
not NOT1 (N251, N249);
and AND3 (N252, N248, N110, N242);
nor NOR3 (N253, N71, N187, N241);
nor NOR2 (N254, N251, N13);
not NOT1 (N255, N229);
and AND2 (N256, N253, N207);
and AND3 (N257, N235, N246, N172);
and AND3 (N258, N257, N117, N211);
buf BUF1 (N259, N243);
or OR4 (N260, N259, N220, N46, N167);
buf BUF1 (N261, N244);
or OR2 (N262, N261, N251);
or OR4 (N263, N262, N203, N31, N106);
or OR2 (N264, N256, N161);
buf BUF1 (N265, N238);
nor NOR4 (N266, N255, N89, N69, N231);
and AND4 (N267, N233, N49, N174, N25);
nor NOR2 (N268, N264, N190);
or OR4 (N269, N268, N97, N174, N193);
nor NOR4 (N270, N269, N11, N165, N247);
buf BUF1 (N271, N266);
not NOT1 (N272, N265);
xor XOR2 (N273, N263, N236);
buf BUF1 (N274, N270);
xor XOR2 (N275, N274, N140);
not NOT1 (N276, N260);
buf BUF1 (N277, N252);
xor XOR2 (N278, N277, N59);
or OR4 (N279, N272, N7, N228, N188);
or OR4 (N280, N250, N174, N266, N145);
buf BUF1 (N281, N276);
xor XOR2 (N282, N278, N163);
not NOT1 (N283, N280);
buf BUF1 (N284, N273);
or OR4 (N285, N279, N235, N180, N12);
nor NOR2 (N286, N254, N1);
or OR3 (N287, N284, N258, N39);
nand NAND3 (N288, N153, N242, N50);
or OR4 (N289, N271, N250, N7, N214);
nor NOR3 (N290, N283, N264, N234);
and AND3 (N291, N285, N185, N237);
xor XOR2 (N292, N289, N238);
not NOT1 (N293, N275);
xor XOR2 (N294, N282, N45);
not NOT1 (N295, N281);
not NOT1 (N296, N294);
nor NOR2 (N297, N288, N4);
not NOT1 (N298, N295);
or OR3 (N299, N291, N72, N294);
not NOT1 (N300, N292);
xor XOR2 (N301, N290, N227);
buf BUF1 (N302, N293);
nand NAND2 (N303, N296, N73);
nor NOR3 (N304, N286, N246, N283);
or OR4 (N305, N297, N253, N91, N182);
not NOT1 (N306, N299);
buf BUF1 (N307, N287);
and AND3 (N308, N306, N101, N201);
xor XOR2 (N309, N307, N228);
nand NAND2 (N310, N267, N206);
nand NAND3 (N311, N303, N280, N270);
nand NAND4 (N312, N301, N197, N109, N2);
and AND3 (N313, N309, N33, N61);
xor XOR2 (N314, N313, N204);
xor XOR2 (N315, N302, N118);
nor NOR3 (N316, N305, N271, N61);
nor NOR4 (N317, N304, N52, N110, N129);
nand NAND2 (N318, N317, N276);
nor NOR2 (N319, N315, N317);
and AND3 (N320, N316, N58, N237);
nor NOR4 (N321, N319, N187, N253, N186);
xor XOR2 (N322, N321, N119);
nor NOR3 (N323, N308, N222, N35);
buf BUF1 (N324, N298);
and AND4 (N325, N300, N153, N154, N319);
buf BUF1 (N326, N311);
and AND3 (N327, N312, N154, N62);
nor NOR3 (N328, N326, N72, N234);
nor NOR2 (N329, N327, N72);
nand NAND3 (N330, N324, N77, N231);
or OR3 (N331, N322, N312, N221);
nand NAND3 (N332, N328, N168, N187);
and AND2 (N333, N318, N56);
nor NOR3 (N334, N310, N1, N290);
not NOT1 (N335, N333);
or OR2 (N336, N331, N236);
not NOT1 (N337, N330);
not NOT1 (N338, N325);
nand NAND3 (N339, N329, N329, N201);
buf BUF1 (N340, N314);
not NOT1 (N341, N340);
and AND3 (N342, N320, N310, N114);
nand NAND4 (N343, N341, N175, N28, N174);
nand NAND3 (N344, N323, N312, N206);
or OR4 (N345, N334, N129, N267, N33);
nand NAND4 (N346, N345, N225, N276, N15);
xor XOR2 (N347, N338, N202);
xor XOR2 (N348, N347, N100);
nand NAND4 (N349, N348, N307, N340, N33);
buf BUF1 (N350, N335);
nor NOR3 (N351, N350, N283, N67);
nor NOR2 (N352, N349, N39);
and AND4 (N353, N344, N261, N350, N35);
nand NAND3 (N354, N342, N319, N253);
nand NAND2 (N355, N337, N28);
nand NAND4 (N356, N332, N284, N273, N302);
not NOT1 (N357, N354);
nand NAND3 (N358, N355, N271, N328);
and AND3 (N359, N356, N332, N18);
and AND2 (N360, N336, N183);
and AND3 (N361, N359, N34, N291);
or OR4 (N362, N353, N210, N221, N248);
or OR4 (N363, N360, N279, N167, N159);
xor XOR2 (N364, N357, N257);
xor XOR2 (N365, N364, N145);
buf BUF1 (N366, N346);
nor NOR4 (N367, N358, N219, N55, N38);
and AND3 (N368, N362, N321, N364);
xor XOR2 (N369, N366, N193);
and AND3 (N370, N365, N245, N36);
or OR3 (N371, N369, N84, N244);
or OR2 (N372, N351, N102);
or OR2 (N373, N361, N353);
xor XOR2 (N374, N371, N118);
xor XOR2 (N375, N363, N366);
and AND3 (N376, N375, N247, N110);
nand NAND3 (N377, N370, N8, N180);
xor XOR2 (N378, N377, N162);
not NOT1 (N379, N367);
or OR2 (N380, N374, N212);
not NOT1 (N381, N372);
xor XOR2 (N382, N380, N337);
nor NOR3 (N383, N373, N244, N310);
nand NAND2 (N384, N381, N370);
nand NAND4 (N385, N383, N122, N372, N76);
or OR3 (N386, N368, N253, N126);
buf BUF1 (N387, N379);
not NOT1 (N388, N376);
or OR2 (N389, N382, N379);
buf BUF1 (N390, N384);
nor NOR3 (N391, N388, N126, N219);
buf BUF1 (N392, N378);
nand NAND2 (N393, N387, N87);
not NOT1 (N394, N389);
nor NOR4 (N395, N392, N161, N98, N191);
nor NOR3 (N396, N391, N12, N300);
and AND3 (N397, N385, N164, N81);
buf BUF1 (N398, N386);
nand NAND2 (N399, N394, N151);
xor XOR2 (N400, N343, N360);
buf BUF1 (N401, N398);
xor XOR2 (N402, N390, N86);
xor XOR2 (N403, N400, N157);
buf BUF1 (N404, N403);
nor NOR2 (N405, N399, N344);
and AND2 (N406, N396, N153);
nor NOR3 (N407, N393, N175, N219);
nand NAND2 (N408, N395, N227);
and AND2 (N409, N352, N34);
nor NOR2 (N410, N401, N248);
xor XOR2 (N411, N397, N88);
xor XOR2 (N412, N339, N390);
and AND4 (N413, N404, N186, N384, N114);
and AND2 (N414, N406, N174);
or OR4 (N415, N412, N414, N47, N358);
xor XOR2 (N416, N357, N172);
nor NOR3 (N417, N402, N208, N228);
and AND3 (N418, N405, N173, N177);
xor XOR2 (N419, N409, N101);
xor XOR2 (N420, N416, N74);
buf BUF1 (N421, N407);
nor NOR4 (N422, N411, N320, N147, N403);
xor XOR2 (N423, N410, N174);
nand NAND3 (N424, N417, N330, N365);
nor NOR3 (N425, N424, N86, N112);
not NOT1 (N426, N408);
nor NOR2 (N427, N422, N194);
nand NAND3 (N428, N423, N347, N73);
nand NAND3 (N429, N419, N130, N71);
and AND2 (N430, N429, N243);
and AND2 (N431, N418, N174);
buf BUF1 (N432, N415);
buf BUF1 (N433, N427);
buf BUF1 (N434, N425);
or OR3 (N435, N433, N311, N355);
buf BUF1 (N436, N420);
buf BUF1 (N437, N434);
nand NAND3 (N438, N413, N231, N34);
xor XOR2 (N439, N438, N88);
or OR4 (N440, N421, N115, N98, N21);
not NOT1 (N441, N426);
buf BUF1 (N442, N432);
nand NAND2 (N443, N442, N140);
or OR4 (N444, N435, N31, N332, N134);
nor NOR3 (N445, N441, N369, N255);
xor XOR2 (N446, N437, N276);
or OR4 (N447, N428, N392, N172, N98);
xor XOR2 (N448, N446, N212);
nand NAND4 (N449, N443, N379, N136, N56);
xor XOR2 (N450, N445, N398);
nor NOR4 (N451, N440, N252, N342, N345);
and AND4 (N452, N436, N115, N294, N260);
nand NAND3 (N453, N449, N337, N165);
or OR3 (N454, N431, N105, N74);
not NOT1 (N455, N447);
xor XOR2 (N456, N453, N58);
xor XOR2 (N457, N452, N341);
and AND4 (N458, N454, N80, N176, N31);
or OR3 (N459, N457, N331, N360);
buf BUF1 (N460, N430);
nand NAND2 (N461, N458, N241);
not NOT1 (N462, N439);
and AND3 (N463, N459, N87, N10);
and AND2 (N464, N461, N313);
and AND2 (N465, N462, N86);
buf BUF1 (N466, N456);
not NOT1 (N467, N444);
or OR4 (N468, N466, N51, N36, N405);
and AND4 (N469, N463, N355, N410, N453);
nor NOR2 (N470, N448, N365);
and AND4 (N471, N469, N186, N105, N20);
or OR2 (N472, N450, N59);
buf BUF1 (N473, N460);
nand NAND2 (N474, N455, N439);
nand NAND2 (N475, N467, N118);
nand NAND2 (N476, N472, N396);
or OR4 (N477, N475, N98, N130, N253);
not NOT1 (N478, N474);
buf BUF1 (N479, N470);
buf BUF1 (N480, N476);
not NOT1 (N481, N465);
or OR2 (N482, N451, N323);
not NOT1 (N483, N464);
xor XOR2 (N484, N478, N18);
and AND3 (N485, N471, N436, N152);
not NOT1 (N486, N473);
or OR4 (N487, N482, N394, N129, N224);
xor XOR2 (N488, N483, N431);
not NOT1 (N489, N481);
xor XOR2 (N490, N477, N158);
not NOT1 (N491, N488);
or OR4 (N492, N491, N326, N116, N304);
or OR4 (N493, N492, N258, N432, N369);
nand NAND2 (N494, N487, N378);
and AND2 (N495, N468, N77);
xor XOR2 (N496, N480, N146);
buf BUF1 (N497, N486);
nor NOR2 (N498, N497, N379);
nand NAND3 (N499, N494, N282, N95);
xor XOR2 (N500, N490, N457);
xor XOR2 (N501, N479, N431);
nor NOR2 (N502, N500, N324);
nand NAND4 (N503, N493, N324, N90, N324);
or OR2 (N504, N484, N212);
and AND2 (N505, N498, N430);
not NOT1 (N506, N501);
xor XOR2 (N507, N496, N400);
xor XOR2 (N508, N502, N38);
not NOT1 (N509, N507);
buf BUF1 (N510, N504);
and AND2 (N511, N503, N192);
and AND3 (N512, N499, N371, N299);
or OR3 (N513, N485, N386, N7);
buf BUF1 (N514, N495);
nand NAND4 (N515, N506, N115, N354, N374);
and AND3 (N516, N510, N7, N484);
nor NOR4 (N517, N511, N111, N37, N237);
xor XOR2 (N518, N515, N117);
nor NOR4 (N519, N517, N247, N135, N210);
nand NAND3 (N520, N489, N482, N467);
or OR3 (N521, N519, N511, N491);
nand NAND2 (N522, N521, N190);
buf BUF1 (N523, N522);
or OR3 (N524, N516, N412, N99);
xor XOR2 (N525, N523, N485);
or OR2 (N526, N508, N123);
and AND2 (N527, N526, N499);
not NOT1 (N528, N513);
nor NOR2 (N529, N505, N511);
or OR2 (N530, N514, N125);
buf BUF1 (N531, N528);
nand NAND4 (N532, N527, N438, N524, N529);
nand NAND3 (N533, N218, N371, N398);
nand NAND3 (N534, N150, N181, N451);
buf BUF1 (N535, N530);
not NOT1 (N536, N520);
and AND4 (N537, N525, N303, N142, N335);
and AND3 (N538, N531, N321, N326);
nor NOR4 (N539, N509, N187, N505, N538);
not NOT1 (N540, N318);
xor XOR2 (N541, N539, N337);
and AND4 (N542, N518, N282, N170, N277);
nor NOR3 (N543, N541, N29, N463);
nand NAND2 (N544, N536, N284);
nand NAND4 (N545, N534, N17, N400, N445);
or OR4 (N546, N512, N94, N253, N204);
and AND2 (N547, N543, N167);
nand NAND2 (N548, N540, N390);
or OR2 (N549, N532, N471);
and AND4 (N550, N533, N322, N89, N439);
nor NOR3 (N551, N548, N243, N330);
buf BUF1 (N552, N542);
not NOT1 (N553, N551);
xor XOR2 (N554, N553, N405);
not NOT1 (N555, N535);
xor XOR2 (N556, N537, N194);
nor NOR3 (N557, N550, N498, N41);
buf BUF1 (N558, N549);
and AND4 (N559, N545, N449, N503, N391);
nor NOR3 (N560, N556, N454, N481);
or OR4 (N561, N560, N304, N335, N494);
and AND3 (N562, N547, N142, N3);
buf BUF1 (N563, N558);
nor NOR3 (N564, N554, N387, N206);
not NOT1 (N565, N555);
buf BUF1 (N566, N563);
buf BUF1 (N567, N561);
nor NOR3 (N568, N567, N216, N210);
buf BUF1 (N569, N564);
or OR2 (N570, N557, N526);
buf BUF1 (N571, N544);
and AND4 (N572, N559, N66, N231, N251);
nand NAND3 (N573, N571, N261, N238);
nand NAND2 (N574, N565, N141);
and AND4 (N575, N570, N476, N402, N451);
buf BUF1 (N576, N575);
buf BUF1 (N577, N562);
xor XOR2 (N578, N568, N141);
xor XOR2 (N579, N569, N174);
and AND2 (N580, N576, N74);
nor NOR2 (N581, N566, N403);
buf BUF1 (N582, N546);
nand NAND2 (N583, N580, N168);
and AND2 (N584, N582, N474);
or OR3 (N585, N573, N541, N113);
and AND3 (N586, N572, N39, N269);
and AND2 (N587, N583, N169);
nand NAND4 (N588, N586, N435, N451, N230);
or OR4 (N589, N584, N482, N94, N400);
buf BUF1 (N590, N589);
nor NOR3 (N591, N574, N555, N485);
and AND4 (N592, N588, N38, N227, N124);
not NOT1 (N593, N578);
not NOT1 (N594, N591);
nor NOR4 (N595, N577, N111, N221, N282);
nand NAND3 (N596, N579, N209, N129);
xor XOR2 (N597, N592, N403);
xor XOR2 (N598, N587, N408);
xor XOR2 (N599, N590, N30);
not NOT1 (N600, N594);
buf BUF1 (N601, N597);
not NOT1 (N602, N599);
nor NOR2 (N603, N602, N27);
or OR3 (N604, N581, N36, N42);
nand NAND4 (N605, N593, N560, N395, N520);
and AND3 (N606, N552, N470, N418);
or OR3 (N607, N596, N495, N461);
xor XOR2 (N608, N600, N90);
nand NAND4 (N609, N604, N179, N193, N478);
or OR2 (N610, N598, N502);
or OR3 (N611, N610, N429, N297);
and AND3 (N612, N606, N439, N498);
nor NOR4 (N613, N605, N272, N247, N285);
buf BUF1 (N614, N609);
or OR4 (N615, N603, N552, N213, N102);
nor NOR3 (N616, N614, N551, N63);
buf BUF1 (N617, N595);
nor NOR4 (N618, N611, N586, N387, N56);
not NOT1 (N619, N615);
not NOT1 (N620, N607);
or OR3 (N621, N618, N74, N113);
not NOT1 (N622, N608);
and AND2 (N623, N620, N22);
buf BUF1 (N624, N612);
xor XOR2 (N625, N619, N37);
nor NOR2 (N626, N616, N384);
xor XOR2 (N627, N621, N79);
nand NAND3 (N628, N622, N183, N588);
not NOT1 (N629, N601);
nand NAND2 (N630, N627, N559);
or OR3 (N631, N624, N610, N87);
not NOT1 (N632, N628);
not NOT1 (N633, N631);
nor NOR4 (N634, N633, N386, N363, N302);
or OR3 (N635, N629, N165, N297);
buf BUF1 (N636, N626);
not NOT1 (N637, N623);
xor XOR2 (N638, N637, N492);
buf BUF1 (N639, N585);
and AND3 (N640, N632, N627, N236);
buf BUF1 (N641, N625);
or OR2 (N642, N640, N378);
buf BUF1 (N643, N617);
and AND3 (N644, N634, N89, N70);
xor XOR2 (N645, N613, N571);
nand NAND4 (N646, N635, N208, N166, N225);
nor NOR3 (N647, N646, N619, N645);
nand NAND2 (N648, N5, N332);
and AND4 (N649, N642, N171, N447, N607);
nand NAND2 (N650, N641, N482);
xor XOR2 (N651, N636, N594);
buf BUF1 (N652, N650);
buf BUF1 (N653, N644);
nand NAND4 (N654, N643, N177, N488, N229);
or OR3 (N655, N648, N267, N410);
xor XOR2 (N656, N630, N213);
and AND2 (N657, N655, N509);
buf BUF1 (N658, N638);
not NOT1 (N659, N656);
not NOT1 (N660, N647);
nor NOR4 (N661, N651, N250, N200, N656);
nand NAND3 (N662, N658, N210, N91);
nor NOR3 (N663, N649, N596, N287);
nor NOR2 (N664, N653, N566);
not NOT1 (N665, N663);
not NOT1 (N666, N659);
not NOT1 (N667, N664);
not NOT1 (N668, N639);
xor XOR2 (N669, N668, N534);
nand NAND2 (N670, N662, N374);
buf BUF1 (N671, N666);
xor XOR2 (N672, N657, N214);
and AND3 (N673, N661, N640, N87);
or OR4 (N674, N670, N466, N36, N114);
nor NOR2 (N675, N673, N597);
and AND2 (N676, N654, N579);
nand NAND3 (N677, N667, N365, N488);
not NOT1 (N678, N677);
not NOT1 (N679, N674);
nand NAND2 (N680, N669, N588);
not NOT1 (N681, N678);
and AND2 (N682, N665, N66);
not NOT1 (N683, N652);
and AND4 (N684, N682, N499, N225, N654);
or OR2 (N685, N675, N296);
nor NOR4 (N686, N676, N542, N79, N73);
and AND3 (N687, N672, N441, N40);
nand NAND2 (N688, N660, N239);
xor XOR2 (N689, N681, N575);
nor NOR2 (N690, N686, N299);
or OR2 (N691, N687, N408);
nand NAND3 (N692, N688, N198, N136);
not NOT1 (N693, N679);
nand NAND3 (N694, N692, N667, N74);
nand NAND2 (N695, N691, N446);
xor XOR2 (N696, N684, N260);
nand NAND2 (N697, N671, N534);
nand NAND2 (N698, N689, N395);
nor NOR2 (N699, N693, N143);
not NOT1 (N700, N685);
and AND2 (N701, N696, N134);
buf BUF1 (N702, N701);
nand NAND3 (N703, N698, N52, N473);
not NOT1 (N704, N690);
nor NOR2 (N705, N680, N295);
nor NOR3 (N706, N702, N104, N145);
not NOT1 (N707, N703);
or OR2 (N708, N699, N133);
or OR2 (N709, N700, N623);
or OR4 (N710, N704, N173, N649, N366);
or OR4 (N711, N707, N576, N124, N598);
or OR3 (N712, N695, N172, N143);
nor NOR3 (N713, N709, N649, N383);
not NOT1 (N714, N710);
or OR3 (N715, N683, N358, N477);
nor NOR3 (N716, N706, N154, N652);
not NOT1 (N717, N714);
buf BUF1 (N718, N717);
or OR4 (N719, N712, N61, N524, N25);
and AND2 (N720, N694, N328);
or OR3 (N721, N697, N33, N293);
nand NAND2 (N722, N718, N238);
nand NAND2 (N723, N713, N127);
not NOT1 (N724, N723);
or OR4 (N725, N708, N234, N184, N525);
and AND4 (N726, N720, N520, N144, N498);
not NOT1 (N727, N711);
xor XOR2 (N728, N715, N598);
and AND2 (N729, N727, N47);
not NOT1 (N730, N719);
buf BUF1 (N731, N726);
nor NOR4 (N732, N728, N142, N380, N173);
nand NAND3 (N733, N724, N169, N702);
or OR3 (N734, N721, N415, N731);
xor XOR2 (N735, N629, N356);
xor XOR2 (N736, N735, N719);
nor NOR2 (N737, N734, N639);
xor XOR2 (N738, N736, N575);
nand NAND4 (N739, N738, N394, N220, N670);
or OR4 (N740, N733, N188, N734, N664);
xor XOR2 (N741, N739, N105);
or OR2 (N742, N741, N665);
not NOT1 (N743, N722);
nand NAND3 (N744, N705, N197, N578);
or OR4 (N745, N740, N58, N651, N73);
and AND3 (N746, N743, N421, N552);
nor NOR4 (N747, N737, N391, N575, N39);
or OR4 (N748, N745, N320, N144, N675);
not NOT1 (N749, N748);
not NOT1 (N750, N747);
buf BUF1 (N751, N742);
and AND4 (N752, N729, N547, N441, N470);
nand NAND2 (N753, N716, N42);
or OR4 (N754, N732, N120, N705, N492);
buf BUF1 (N755, N730);
nand NAND4 (N756, N746, N55, N748, N253);
or OR3 (N757, N725, N582, N678);
nor NOR2 (N758, N753, N83);
or OR4 (N759, N758, N475, N639, N492);
nor NOR2 (N760, N759, N578);
and AND2 (N761, N757, N341);
xor XOR2 (N762, N760, N210);
xor XOR2 (N763, N762, N507);
nor NOR4 (N764, N763, N759, N388, N90);
nor NOR4 (N765, N752, N163, N64, N420);
not NOT1 (N766, N749);
buf BUF1 (N767, N756);
and AND4 (N768, N751, N168, N684, N764);
and AND2 (N769, N444, N479);
xor XOR2 (N770, N755, N586);
not NOT1 (N771, N770);
or OR2 (N772, N771, N307);
or OR3 (N773, N766, N121, N469);
buf BUF1 (N774, N772);
or OR2 (N775, N744, N231);
nor NOR2 (N776, N769, N240);
or OR3 (N777, N750, N302, N79);
xor XOR2 (N778, N776, N400);
and AND3 (N779, N774, N722, N443);
xor XOR2 (N780, N761, N34);
and AND3 (N781, N768, N375, N161);
nand NAND3 (N782, N779, N606, N636);
nand NAND4 (N783, N754, N579, N509, N737);
nand NAND4 (N784, N782, N670, N19, N472);
and AND3 (N785, N784, N220, N199);
or OR4 (N786, N777, N391, N234, N361);
or OR4 (N787, N773, N722, N518, N233);
and AND4 (N788, N781, N190, N310, N336);
nand NAND2 (N789, N775, N740);
and AND2 (N790, N780, N363);
or OR4 (N791, N783, N654, N480, N221);
xor XOR2 (N792, N788, N26);
and AND3 (N793, N791, N22, N635);
nand NAND4 (N794, N786, N526, N274, N571);
and AND3 (N795, N767, N74, N703);
nor NOR3 (N796, N789, N123, N711);
not NOT1 (N797, N787);
and AND4 (N798, N795, N590, N525, N505);
or OR4 (N799, N797, N447, N580, N58);
nor NOR2 (N800, N798, N380);
xor XOR2 (N801, N794, N575);
nor NOR2 (N802, N796, N494);
not NOT1 (N803, N785);
nand NAND2 (N804, N803, N784);
not NOT1 (N805, N765);
nor NOR4 (N806, N799, N746, N229, N459);
nand NAND4 (N807, N801, N514, N387, N183);
nand NAND3 (N808, N793, N185, N176);
and AND3 (N809, N802, N734, N562);
and AND4 (N810, N800, N329, N43, N70);
not NOT1 (N811, N805);
nand NAND2 (N812, N804, N786);
not NOT1 (N813, N811);
buf BUF1 (N814, N813);
nor NOR2 (N815, N807, N100);
xor XOR2 (N816, N814, N154);
and AND3 (N817, N815, N489, N124);
or OR2 (N818, N816, N454);
buf BUF1 (N819, N818);
and AND4 (N820, N809, N265, N639, N383);
or OR2 (N821, N806, N492);
and AND2 (N822, N790, N265);
or OR4 (N823, N812, N264, N129, N305);
or OR2 (N824, N820, N750);
buf BUF1 (N825, N822);
or OR3 (N826, N823, N685, N783);
nor NOR3 (N827, N819, N383, N227);
buf BUF1 (N828, N827);
nor NOR2 (N829, N826, N8);
xor XOR2 (N830, N828, N334);
or OR3 (N831, N810, N674, N718);
nand NAND4 (N832, N792, N75, N371, N623);
buf BUF1 (N833, N831);
nor NOR3 (N834, N817, N550, N101);
xor XOR2 (N835, N832, N710);
and AND2 (N836, N833, N732);
or OR3 (N837, N835, N204, N611);
and AND3 (N838, N830, N28, N612);
nand NAND4 (N839, N824, N528, N664, N239);
nand NAND4 (N840, N825, N706, N475, N15);
and AND2 (N841, N821, N147);
not NOT1 (N842, N836);
nor NOR3 (N843, N839, N165, N711);
nor NOR2 (N844, N778, N377);
nor NOR4 (N845, N841, N60, N40, N350);
xor XOR2 (N846, N829, N808);
buf BUF1 (N847, N401);
xor XOR2 (N848, N845, N627);
or OR3 (N849, N843, N152, N507);
xor XOR2 (N850, N849, N132);
or OR3 (N851, N837, N391, N122);
not NOT1 (N852, N846);
buf BUF1 (N853, N851);
nand NAND3 (N854, N848, N416, N786);
buf BUF1 (N855, N834);
nor NOR2 (N856, N838, N357);
buf BUF1 (N857, N854);
xor XOR2 (N858, N840, N210);
nand NAND4 (N859, N852, N737, N89, N788);
buf BUF1 (N860, N850);
or OR3 (N861, N844, N187, N778);
not NOT1 (N862, N856);
xor XOR2 (N863, N860, N804);
nor NOR3 (N864, N842, N36, N321);
xor XOR2 (N865, N864, N716);
not NOT1 (N866, N857);
and AND2 (N867, N861, N315);
nor NOR3 (N868, N865, N828, N127);
xor XOR2 (N869, N855, N610);
nor NOR3 (N870, N847, N748, N196);
nor NOR3 (N871, N863, N774, N156);
nand NAND2 (N872, N853, N787);
not NOT1 (N873, N866);
buf BUF1 (N874, N869);
and AND2 (N875, N867, N295);
or OR3 (N876, N872, N62, N780);
xor XOR2 (N877, N862, N681);
nand NAND4 (N878, N875, N464, N863, N397);
or OR4 (N879, N876, N639, N361, N519);
or OR3 (N880, N870, N582, N798);
nor NOR3 (N881, N871, N555, N229);
xor XOR2 (N882, N877, N98);
nand NAND3 (N883, N880, N493, N544);
nor NOR4 (N884, N882, N828, N819, N878);
nor NOR4 (N885, N599, N235, N434, N390);
xor XOR2 (N886, N873, N827);
buf BUF1 (N887, N886);
xor XOR2 (N888, N858, N522);
buf BUF1 (N889, N887);
and AND3 (N890, N879, N457, N2);
nor NOR3 (N891, N890, N26, N97);
nand NAND3 (N892, N883, N556, N232);
and AND3 (N893, N888, N398, N577);
buf BUF1 (N894, N891);
buf BUF1 (N895, N884);
nor NOR2 (N896, N874, N816);
and AND2 (N897, N885, N206);
not NOT1 (N898, N896);
and AND2 (N899, N894, N441);
and AND3 (N900, N868, N468, N412);
xor XOR2 (N901, N897, N730);
buf BUF1 (N902, N889);
xor XOR2 (N903, N902, N232);
nand NAND2 (N904, N898, N739);
buf BUF1 (N905, N859);
nor NOR3 (N906, N901, N531, N815);
buf BUF1 (N907, N899);
nand NAND4 (N908, N893, N309, N498, N273);
xor XOR2 (N909, N892, N709);
buf BUF1 (N910, N900);
nand NAND3 (N911, N903, N674, N886);
nor NOR4 (N912, N905, N390, N710, N345);
and AND4 (N913, N881, N280, N373, N332);
nand NAND4 (N914, N912, N369, N727, N692);
nor NOR3 (N915, N909, N501, N884);
not NOT1 (N916, N904);
or OR4 (N917, N895, N699, N285, N603);
or OR2 (N918, N917, N416);
nor NOR2 (N919, N906, N291);
nor NOR2 (N920, N914, N170);
nor NOR4 (N921, N919, N371, N831, N639);
or OR2 (N922, N911, N800);
or OR3 (N923, N908, N177, N59);
nand NAND2 (N924, N916, N509);
buf BUF1 (N925, N923);
not NOT1 (N926, N924);
nor NOR2 (N927, N915, N754);
not NOT1 (N928, N926);
xor XOR2 (N929, N922, N810);
nor NOR2 (N930, N929, N394);
buf BUF1 (N931, N907);
nor NOR3 (N932, N918, N327, N370);
nor NOR2 (N933, N927, N11);
xor XOR2 (N934, N933, N815);
nand NAND3 (N935, N930, N621, N925);
not NOT1 (N936, N610);
and AND3 (N937, N934, N470, N737);
nand NAND4 (N938, N937, N443, N162, N110);
buf BUF1 (N939, N938);
or OR3 (N940, N932, N830, N392);
nor NOR2 (N941, N931, N685);
or OR2 (N942, N940, N395);
not NOT1 (N943, N928);
and AND2 (N944, N910, N204);
nor NOR3 (N945, N920, N689, N32);
nand NAND3 (N946, N936, N643, N534);
xor XOR2 (N947, N942, N686);
buf BUF1 (N948, N913);
or OR2 (N949, N935, N23);
or OR4 (N950, N939, N132, N409, N216);
or OR2 (N951, N945, N396);
and AND3 (N952, N943, N238, N217);
xor XOR2 (N953, N921, N54);
not NOT1 (N954, N953);
or OR2 (N955, N949, N493);
nor NOR4 (N956, N950, N620, N553, N452);
nand NAND4 (N957, N956, N2, N153, N140);
and AND2 (N958, N946, N429);
or OR4 (N959, N951, N352, N577, N30);
nand NAND3 (N960, N952, N67, N945);
buf BUF1 (N961, N944);
nor NOR3 (N962, N958, N552, N269);
or OR4 (N963, N948, N691, N576, N709);
nand NAND2 (N964, N963, N945);
buf BUF1 (N965, N954);
buf BUF1 (N966, N961);
nand NAND3 (N967, N957, N522, N386);
not NOT1 (N968, N965);
xor XOR2 (N969, N947, N899);
nand NAND4 (N970, N962, N226, N897, N832);
and AND4 (N971, N964, N497, N301, N17);
buf BUF1 (N972, N970);
and AND3 (N973, N959, N240, N550);
or OR2 (N974, N968, N136);
xor XOR2 (N975, N955, N203);
xor XOR2 (N976, N960, N697);
xor XOR2 (N977, N966, N452);
or OR3 (N978, N976, N712, N231);
buf BUF1 (N979, N941);
buf BUF1 (N980, N979);
nor NOR2 (N981, N980, N47);
buf BUF1 (N982, N972);
or OR2 (N983, N969, N649);
xor XOR2 (N984, N982, N111);
buf BUF1 (N985, N967);
and AND3 (N986, N971, N390, N144);
not NOT1 (N987, N986);
nor NOR4 (N988, N975, N309, N580, N780);
xor XOR2 (N989, N988, N547);
nor NOR4 (N990, N987, N717, N818, N140);
buf BUF1 (N991, N989);
xor XOR2 (N992, N974, N476);
nor NOR3 (N993, N983, N104, N398);
nor NOR3 (N994, N978, N369, N901);
buf BUF1 (N995, N994);
and AND4 (N996, N990, N670, N733, N518);
or OR2 (N997, N995, N723);
and AND3 (N998, N985, N350, N119);
xor XOR2 (N999, N996, N385);
or OR3 (N1000, N984, N595, N196);
nand NAND4 (N1001, N999, N949, N132, N994);
not NOT1 (N1002, N998);
not NOT1 (N1003, N981);
nor NOR2 (N1004, N1001, N703);
nand NAND4 (N1005, N993, N414, N723, N385);
buf BUF1 (N1006, N997);
nand NAND4 (N1007, N1005, N644, N86, N741);
nand NAND4 (N1008, N1003, N487, N811, N649);
buf BUF1 (N1009, N1006);
or OR3 (N1010, N1004, N684, N837);
and AND4 (N1011, N977, N450, N680, N839);
xor XOR2 (N1012, N1000, N209);
xor XOR2 (N1013, N1012, N836);
nor NOR2 (N1014, N973, N299);
or OR4 (N1015, N1010, N914, N292, N92);
xor XOR2 (N1016, N992, N363);
or OR2 (N1017, N1007, N963);
xor XOR2 (N1018, N1014, N353);
and AND3 (N1019, N1008, N92, N248);
and AND4 (N1020, N1015, N182, N85, N996);
not NOT1 (N1021, N1002);
nand NAND4 (N1022, N1017, N472, N242, N702);
and AND2 (N1023, N991, N170);
and AND3 (N1024, N1020, N757, N442);
nand NAND2 (N1025, N1016, N347);
nor NOR3 (N1026, N1024, N817, N702);
and AND3 (N1027, N1022, N266, N564);
nand NAND4 (N1028, N1018, N318, N523, N73);
not NOT1 (N1029, N1013);
nor NOR3 (N1030, N1025, N456, N75);
buf BUF1 (N1031, N1028);
buf BUF1 (N1032, N1019);
or OR2 (N1033, N1027, N900);
nand NAND2 (N1034, N1033, N836);
nand NAND3 (N1035, N1011, N412, N442);
nand NAND4 (N1036, N1009, N582, N869, N864);
nand NAND2 (N1037, N1026, N294);
or OR2 (N1038, N1032, N34);
buf BUF1 (N1039, N1023);
nor NOR4 (N1040, N1034, N462, N926, N647);
not NOT1 (N1041, N1030);
not NOT1 (N1042, N1040);
nand NAND4 (N1043, N1035, N498, N127, N938);
or OR2 (N1044, N1031, N684);
and AND3 (N1045, N1041, N172, N124);
xor XOR2 (N1046, N1029, N103);
and AND2 (N1047, N1042, N632);
nor NOR4 (N1048, N1043, N991, N348, N122);
xor XOR2 (N1049, N1046, N611);
not NOT1 (N1050, N1044);
nand NAND3 (N1051, N1038, N376, N7);
nand NAND4 (N1052, N1051, N87, N490, N77);
nand NAND4 (N1053, N1047, N105, N153, N479);
nand NAND4 (N1054, N1053, N425, N475, N470);
nor NOR4 (N1055, N1049, N436, N729, N739);
or OR3 (N1056, N1021, N1020, N960);
or OR2 (N1057, N1045, N317);
buf BUF1 (N1058, N1037);
nor NOR2 (N1059, N1050, N408);
and AND4 (N1060, N1048, N88, N137, N990);
not NOT1 (N1061, N1058);
or OR4 (N1062, N1061, N987, N278, N810);
and AND4 (N1063, N1056, N6, N179, N636);
nand NAND4 (N1064, N1059, N396, N1045, N396);
xor XOR2 (N1065, N1057, N321);
nand NAND3 (N1066, N1060, N913, N122);
buf BUF1 (N1067, N1039);
and AND4 (N1068, N1052, N98, N674, N868);
nor NOR3 (N1069, N1064, N463, N22);
nand NAND3 (N1070, N1055, N372, N806);
nand NAND4 (N1071, N1068, N11, N930, N433);
nor NOR2 (N1072, N1069, N426);
buf BUF1 (N1073, N1072);
buf BUF1 (N1074, N1036);
buf BUF1 (N1075, N1073);
not NOT1 (N1076, N1063);
nor NOR2 (N1077, N1071, N883);
nand NAND2 (N1078, N1077, N320);
or OR2 (N1079, N1065, N395);
nor NOR4 (N1080, N1067, N299, N876, N834);
nand NAND3 (N1081, N1062, N152, N791);
not NOT1 (N1082, N1081);
and AND3 (N1083, N1070, N45, N1075);
nand NAND3 (N1084, N925, N339, N550);
nor NOR3 (N1085, N1079, N658, N215);
nor NOR3 (N1086, N1083, N4, N1023);
nand NAND3 (N1087, N1066, N694, N272);
nand NAND2 (N1088, N1080, N1047);
nor NOR2 (N1089, N1054, N25);
not NOT1 (N1090, N1076);
nor NOR2 (N1091, N1090, N61);
or OR3 (N1092, N1088, N991, N117);
nor NOR4 (N1093, N1082, N920, N644, N967);
nand NAND4 (N1094, N1085, N948, N816, N661);
not NOT1 (N1095, N1094);
xor XOR2 (N1096, N1084, N349);
nor NOR3 (N1097, N1087, N591, N477);
and AND2 (N1098, N1089, N233);
and AND2 (N1099, N1097, N529);
not NOT1 (N1100, N1095);
buf BUF1 (N1101, N1092);
xor XOR2 (N1102, N1074, N569);
xor XOR2 (N1103, N1102, N84);
and AND4 (N1104, N1096, N457, N369, N741);
xor XOR2 (N1105, N1103, N280);
buf BUF1 (N1106, N1105);
and AND4 (N1107, N1101, N309, N711, N1049);
buf BUF1 (N1108, N1099);
buf BUF1 (N1109, N1091);
and AND2 (N1110, N1104, N122);
and AND2 (N1111, N1110, N651);
or OR4 (N1112, N1086, N403, N93, N900);
nor NOR3 (N1113, N1109, N779, N41);
xor XOR2 (N1114, N1078, N137);
or OR4 (N1115, N1107, N894, N1017, N1055);
not NOT1 (N1116, N1112);
xor XOR2 (N1117, N1115, N459);
nand NAND2 (N1118, N1100, N254);
and AND4 (N1119, N1114, N88, N591, N784);
or OR3 (N1120, N1116, N78, N497);
nand NAND4 (N1121, N1117, N770, N675, N362);
nand NAND2 (N1122, N1120, N118);
nor NOR3 (N1123, N1121, N931, N64);
and AND4 (N1124, N1108, N1123, N457, N645);
nand NAND2 (N1125, N138, N628);
xor XOR2 (N1126, N1098, N743);
nand NAND4 (N1127, N1106, N60, N471, N293);
and AND2 (N1128, N1113, N809);
or OR3 (N1129, N1118, N323, N1047);
xor XOR2 (N1130, N1126, N657);
nand NAND2 (N1131, N1129, N275);
nand NAND2 (N1132, N1128, N1048);
nand NAND4 (N1133, N1130, N164, N7, N902);
not NOT1 (N1134, N1133);
nand NAND2 (N1135, N1134, N1078);
and AND2 (N1136, N1124, N600);
or OR4 (N1137, N1135, N381, N970, N389);
not NOT1 (N1138, N1122);
nor NOR3 (N1139, N1132, N7, N488);
nand NAND2 (N1140, N1127, N732);
buf BUF1 (N1141, N1137);
or OR2 (N1142, N1138, N568);
or OR3 (N1143, N1111, N311, N1094);
xor XOR2 (N1144, N1125, N958);
nor NOR2 (N1145, N1119, N1036);
nor NOR4 (N1146, N1143, N683, N464, N1015);
or OR4 (N1147, N1093, N697, N773, N138);
xor XOR2 (N1148, N1140, N311);
buf BUF1 (N1149, N1145);
nand NAND2 (N1150, N1131, N1030);
xor XOR2 (N1151, N1150, N1042);
not NOT1 (N1152, N1139);
and AND3 (N1153, N1142, N250, N415);
nand NAND3 (N1154, N1148, N832, N977);
buf BUF1 (N1155, N1151);
xor XOR2 (N1156, N1154, N602);
xor XOR2 (N1157, N1136, N747);
xor XOR2 (N1158, N1141, N922);
buf BUF1 (N1159, N1152);
and AND3 (N1160, N1144, N524, N993);
not NOT1 (N1161, N1160);
nor NOR4 (N1162, N1149, N56, N1042, N426);
not NOT1 (N1163, N1162);
nor NOR3 (N1164, N1155, N1143, N567);
buf BUF1 (N1165, N1153);
nor NOR3 (N1166, N1159, N1152, N231);
not NOT1 (N1167, N1163);
or OR2 (N1168, N1161, N907);
nor NOR3 (N1169, N1157, N926, N1076);
nor NOR2 (N1170, N1156, N792);
or OR3 (N1171, N1164, N487, N236);
nor NOR2 (N1172, N1171, N1146);
nor NOR4 (N1173, N840, N867, N59, N635);
or OR2 (N1174, N1166, N379);
not NOT1 (N1175, N1165);
and AND2 (N1176, N1168, N122);
and AND3 (N1177, N1158, N641, N400);
or OR2 (N1178, N1147, N20);
and AND4 (N1179, N1176, N882, N25, N1096);
and AND4 (N1180, N1174, N574, N441, N217);
xor XOR2 (N1181, N1172, N1064);
and AND3 (N1182, N1177, N357, N888);
xor XOR2 (N1183, N1173, N555);
nand NAND2 (N1184, N1183, N214);
nor NOR2 (N1185, N1170, N530);
or OR2 (N1186, N1182, N841);
or OR3 (N1187, N1186, N498, N558);
and AND2 (N1188, N1184, N524);
xor XOR2 (N1189, N1188, N994);
nor NOR2 (N1190, N1169, N741);
and AND3 (N1191, N1178, N492, N989);
nand NAND4 (N1192, N1167, N258, N592, N33);
and AND2 (N1193, N1192, N357);
nand NAND3 (N1194, N1189, N330, N615);
nor NOR2 (N1195, N1175, N1074);
nand NAND2 (N1196, N1193, N615);
nand NAND3 (N1197, N1181, N781, N519);
nor NOR4 (N1198, N1187, N458, N342, N1009);
buf BUF1 (N1199, N1190);
or OR4 (N1200, N1180, N556, N614, N234);
nor NOR3 (N1201, N1185, N715, N451);
nor NOR3 (N1202, N1199, N633, N60);
not NOT1 (N1203, N1198);
or OR2 (N1204, N1195, N179);
nor NOR2 (N1205, N1201, N1055);
and AND4 (N1206, N1200, N547, N1001, N124);
nand NAND3 (N1207, N1206, N873, N547);
not NOT1 (N1208, N1203);
not NOT1 (N1209, N1205);
or OR3 (N1210, N1197, N328, N68);
and AND4 (N1211, N1196, N864, N754, N15);
xor XOR2 (N1212, N1211, N1176);
not NOT1 (N1213, N1212);
nor NOR3 (N1214, N1208, N840, N1179);
xor XOR2 (N1215, N710, N352);
or OR3 (N1216, N1210, N603, N303);
xor XOR2 (N1217, N1207, N342);
nand NAND2 (N1218, N1209, N568);
xor XOR2 (N1219, N1202, N1105);
xor XOR2 (N1220, N1204, N908);
nand NAND3 (N1221, N1191, N413, N195);
and AND4 (N1222, N1194, N172, N677, N1104);
or OR2 (N1223, N1214, N1124);
xor XOR2 (N1224, N1222, N851);
xor XOR2 (N1225, N1218, N525);
nand NAND4 (N1226, N1217, N1034, N1054, N534);
xor XOR2 (N1227, N1224, N672);
nand NAND3 (N1228, N1223, N507, N707);
nor NOR2 (N1229, N1226, N290);
and AND4 (N1230, N1228, N799, N245, N28);
nand NAND2 (N1231, N1230, N851);
xor XOR2 (N1232, N1215, N1060);
not NOT1 (N1233, N1227);
xor XOR2 (N1234, N1229, N42);
not NOT1 (N1235, N1234);
buf BUF1 (N1236, N1220);
nand NAND4 (N1237, N1231, N1089, N845, N597);
nor NOR4 (N1238, N1225, N1125, N822, N1076);
not NOT1 (N1239, N1235);
buf BUF1 (N1240, N1236);
xor XOR2 (N1241, N1219, N355);
buf BUF1 (N1242, N1216);
buf BUF1 (N1243, N1213);
and AND4 (N1244, N1232, N511, N771, N991);
or OR2 (N1245, N1241, N992);
or OR2 (N1246, N1239, N1038);
or OR4 (N1247, N1246, N559, N730, N639);
or OR3 (N1248, N1243, N521, N442);
not NOT1 (N1249, N1245);
and AND3 (N1250, N1237, N132, N1022);
buf BUF1 (N1251, N1248);
nor NOR2 (N1252, N1250, N873);
nand NAND3 (N1253, N1242, N1119, N669);
or OR2 (N1254, N1244, N1166);
and AND3 (N1255, N1254, N772, N193);
nand NAND2 (N1256, N1253, N73);
and AND4 (N1257, N1256, N613, N152, N809);
and AND3 (N1258, N1247, N578, N299);
nand NAND4 (N1259, N1221, N1241, N912, N824);
nand NAND3 (N1260, N1240, N1125, N26);
or OR4 (N1261, N1257, N1206, N1223, N467);
xor XOR2 (N1262, N1238, N815);
nand NAND3 (N1263, N1262, N414, N591);
nor NOR3 (N1264, N1260, N918, N807);
xor XOR2 (N1265, N1258, N162);
or OR3 (N1266, N1261, N629, N559);
xor XOR2 (N1267, N1251, N558);
or OR2 (N1268, N1264, N403);
buf BUF1 (N1269, N1263);
xor XOR2 (N1270, N1233, N605);
buf BUF1 (N1271, N1265);
nor NOR2 (N1272, N1252, N658);
not NOT1 (N1273, N1249);
or OR4 (N1274, N1273, N51, N1250, N151);
not NOT1 (N1275, N1266);
nand NAND2 (N1276, N1272, N596);
or OR3 (N1277, N1270, N128, N140);
nor NOR2 (N1278, N1255, N805);
nand NAND4 (N1279, N1267, N1100, N1008, N837);
and AND3 (N1280, N1274, N407, N942);
nand NAND2 (N1281, N1279, N383);
xor XOR2 (N1282, N1259, N718);
buf BUF1 (N1283, N1268);
nor NOR2 (N1284, N1283, N1247);
and AND4 (N1285, N1281, N719, N321, N567);
buf BUF1 (N1286, N1271);
not NOT1 (N1287, N1286);
xor XOR2 (N1288, N1284, N881);
nand NAND4 (N1289, N1280, N136, N620, N83);
and AND2 (N1290, N1278, N1133);
not NOT1 (N1291, N1277);
nand NAND2 (N1292, N1269, N73);
buf BUF1 (N1293, N1291);
buf BUF1 (N1294, N1287);
or OR3 (N1295, N1293, N334, N611);
and AND2 (N1296, N1275, N813);
nand NAND4 (N1297, N1289, N990, N1175, N472);
not NOT1 (N1298, N1292);
xor XOR2 (N1299, N1290, N228);
or OR3 (N1300, N1298, N343, N771);
nand NAND2 (N1301, N1288, N1195);
not NOT1 (N1302, N1282);
not NOT1 (N1303, N1301);
not NOT1 (N1304, N1299);
not NOT1 (N1305, N1303);
not NOT1 (N1306, N1304);
not NOT1 (N1307, N1276);
buf BUF1 (N1308, N1306);
or OR3 (N1309, N1302, N360, N342);
nand NAND4 (N1310, N1309, N293, N772, N852);
not NOT1 (N1311, N1307);
or OR2 (N1312, N1294, N1288);
nand NAND3 (N1313, N1295, N1076, N436);
buf BUF1 (N1314, N1300);
and AND2 (N1315, N1310, N724);
or OR2 (N1316, N1314, N1220);
or OR3 (N1317, N1311, N869, N487);
nor NOR2 (N1318, N1285, N712);
and AND2 (N1319, N1296, N373);
or OR3 (N1320, N1313, N11, N531);
or OR2 (N1321, N1305, N933);
or OR3 (N1322, N1317, N194, N377);
not NOT1 (N1323, N1308);
buf BUF1 (N1324, N1312);
or OR3 (N1325, N1315, N947, N384);
nand NAND3 (N1326, N1320, N1229, N1001);
xor XOR2 (N1327, N1323, N375);
nor NOR2 (N1328, N1322, N513);
xor XOR2 (N1329, N1316, N56);
buf BUF1 (N1330, N1319);
nor NOR2 (N1331, N1329, N955);
nand NAND4 (N1332, N1321, N570, N1068, N784);
nand NAND3 (N1333, N1324, N276, N1220);
nor NOR4 (N1334, N1333, N11, N558, N1221);
buf BUF1 (N1335, N1332);
not NOT1 (N1336, N1335);
nand NAND2 (N1337, N1297, N739);
buf BUF1 (N1338, N1331);
nor NOR3 (N1339, N1318, N554, N824);
not NOT1 (N1340, N1338);
or OR3 (N1341, N1340, N159, N213);
buf BUF1 (N1342, N1326);
xor XOR2 (N1343, N1334, N1109);
nor NOR3 (N1344, N1328, N635, N1246);
not NOT1 (N1345, N1342);
nand NAND3 (N1346, N1325, N698, N612);
nor NOR4 (N1347, N1339, N1226, N432, N751);
nor NOR2 (N1348, N1337, N1171);
xor XOR2 (N1349, N1344, N1328);
and AND2 (N1350, N1347, N1291);
buf BUF1 (N1351, N1341);
xor XOR2 (N1352, N1351, N979);
nand NAND2 (N1353, N1345, N868);
not NOT1 (N1354, N1336);
and AND4 (N1355, N1350, N1279, N126, N1032);
buf BUF1 (N1356, N1353);
or OR4 (N1357, N1330, N929, N1098, N826);
nor NOR4 (N1358, N1354, N771, N632, N380);
or OR3 (N1359, N1352, N1208, N391);
buf BUF1 (N1360, N1327);
nor NOR2 (N1361, N1356, N539);
buf BUF1 (N1362, N1343);
nand NAND4 (N1363, N1359, N448, N251, N724);
or OR4 (N1364, N1360, N419, N208, N608);
or OR2 (N1365, N1348, N486);
not NOT1 (N1366, N1349);
nand NAND3 (N1367, N1362, N105, N1315);
or OR3 (N1368, N1346, N585, N824);
not NOT1 (N1369, N1357);
buf BUF1 (N1370, N1363);
xor XOR2 (N1371, N1367, N1090);
nor NOR2 (N1372, N1355, N349);
and AND3 (N1373, N1361, N547, N297);
buf BUF1 (N1374, N1358);
nand NAND3 (N1375, N1373, N959, N896);
buf BUF1 (N1376, N1369);
xor XOR2 (N1377, N1366, N972);
and AND2 (N1378, N1365, N783);
nor NOR3 (N1379, N1371, N917, N397);
xor XOR2 (N1380, N1364, N780);
buf BUF1 (N1381, N1379);
nor NOR2 (N1382, N1380, N1037);
not NOT1 (N1383, N1382);
nand NAND3 (N1384, N1375, N162, N427);
xor XOR2 (N1385, N1376, N780);
not NOT1 (N1386, N1377);
nand NAND4 (N1387, N1384, N576, N574, N11);
xor XOR2 (N1388, N1370, N188);
or OR2 (N1389, N1372, N389);
nor NOR3 (N1390, N1385, N829, N895);
nor NOR4 (N1391, N1389, N921, N404, N1046);
or OR4 (N1392, N1378, N1065, N1148, N648);
nand NAND3 (N1393, N1383, N1198, N675);
or OR4 (N1394, N1381, N516, N831, N420);
buf BUF1 (N1395, N1390);
buf BUF1 (N1396, N1374);
nand NAND2 (N1397, N1395, N991);
xor XOR2 (N1398, N1391, N1145);
nor NOR4 (N1399, N1397, N820, N529, N1279);
nand NAND4 (N1400, N1387, N433, N1236, N802);
xor XOR2 (N1401, N1393, N490);
not NOT1 (N1402, N1368);
and AND2 (N1403, N1401, N861);
xor XOR2 (N1404, N1396, N206);
and AND4 (N1405, N1400, N275, N724, N1247);
buf BUF1 (N1406, N1404);
buf BUF1 (N1407, N1392);
nor NOR2 (N1408, N1402, N208);
nor NOR3 (N1409, N1407, N552, N519);
buf BUF1 (N1410, N1386);
xor XOR2 (N1411, N1398, N452);
or OR2 (N1412, N1406, N1090);
or OR4 (N1413, N1408, N922, N29, N1342);
not NOT1 (N1414, N1394);
and AND3 (N1415, N1411, N1342, N1127);
buf BUF1 (N1416, N1388);
not NOT1 (N1417, N1403);
xor XOR2 (N1418, N1399, N101);
buf BUF1 (N1419, N1405);
xor XOR2 (N1420, N1413, N351);
not NOT1 (N1421, N1416);
not NOT1 (N1422, N1417);
not NOT1 (N1423, N1419);
and AND2 (N1424, N1410, N443);
xor XOR2 (N1425, N1421, N784);
nor NOR2 (N1426, N1423, N918);
nor NOR4 (N1427, N1422, N116, N823, N1379);
not NOT1 (N1428, N1409);
and AND2 (N1429, N1424, N631);
or OR2 (N1430, N1418, N1207);
nor NOR3 (N1431, N1429, N768, N1143);
xor XOR2 (N1432, N1431, N1018);
not NOT1 (N1433, N1426);
not NOT1 (N1434, N1428);
nand NAND3 (N1435, N1427, N71, N515);
nor NOR4 (N1436, N1435, N993, N262, N1284);
and AND2 (N1437, N1425, N70);
or OR2 (N1438, N1414, N368);
not NOT1 (N1439, N1436);
nor NOR3 (N1440, N1420, N464, N890);
nand NAND3 (N1441, N1430, N690, N417);
buf BUF1 (N1442, N1441);
or OR2 (N1443, N1432, N754);
nor NOR3 (N1444, N1443, N665, N828);
and AND4 (N1445, N1439, N985, N707, N1214);
not NOT1 (N1446, N1434);
buf BUF1 (N1447, N1445);
and AND4 (N1448, N1440, N866, N106, N1288);
xor XOR2 (N1449, N1438, N180);
or OR3 (N1450, N1448, N934, N1195);
or OR3 (N1451, N1447, N842, N1443);
not NOT1 (N1452, N1444);
buf BUF1 (N1453, N1446);
and AND4 (N1454, N1433, N469, N1146, N262);
buf BUF1 (N1455, N1452);
nand NAND2 (N1456, N1454, N355);
nor NOR2 (N1457, N1450, N1306);
not NOT1 (N1458, N1437);
and AND2 (N1459, N1457, N590);
buf BUF1 (N1460, N1453);
buf BUF1 (N1461, N1451);
and AND3 (N1462, N1460, N1350, N1387);
buf BUF1 (N1463, N1462);
not NOT1 (N1464, N1458);
buf BUF1 (N1465, N1415);
buf BUF1 (N1466, N1464);
or OR3 (N1467, N1442, N504, N1183);
and AND2 (N1468, N1465, N1457);
xor XOR2 (N1469, N1467, N538);
nor NOR2 (N1470, N1466, N711);
or OR4 (N1471, N1455, N1197, N474, N1195);
and AND2 (N1472, N1461, N760);
nor NOR3 (N1473, N1459, N260, N1469);
nand NAND3 (N1474, N848, N983, N118);
nand NAND3 (N1475, N1463, N364, N659);
buf BUF1 (N1476, N1456);
nor NOR4 (N1477, N1412, N1088, N994, N1166);
and AND2 (N1478, N1477, N53);
xor XOR2 (N1479, N1468, N361);
and AND4 (N1480, N1472, N282, N1134, N498);
or OR3 (N1481, N1449, N30, N1176);
xor XOR2 (N1482, N1470, N1055);
not NOT1 (N1483, N1478);
buf BUF1 (N1484, N1473);
nand NAND3 (N1485, N1483, N1418, N1188);
or OR3 (N1486, N1485, N1052, N61);
nand NAND3 (N1487, N1484, N103, N747);
nor NOR3 (N1488, N1482, N595, N422);
nand NAND4 (N1489, N1481, N320, N1023, N349);
nor NOR3 (N1490, N1475, N1361, N513);
not NOT1 (N1491, N1488);
nand NAND4 (N1492, N1476, N1465, N1308, N433);
xor XOR2 (N1493, N1489, N1073);
and AND4 (N1494, N1491, N233, N572, N262);
not NOT1 (N1495, N1490);
buf BUF1 (N1496, N1487);
nand NAND4 (N1497, N1486, N538, N442, N1206);
buf BUF1 (N1498, N1471);
or OR2 (N1499, N1479, N1495);
nand NAND4 (N1500, N750, N854, N1013, N550);
not NOT1 (N1501, N1498);
or OR2 (N1502, N1501, N617);
or OR3 (N1503, N1493, N578, N212);
not NOT1 (N1504, N1500);
nand NAND4 (N1505, N1499, N1263, N1055, N1289);
buf BUF1 (N1506, N1505);
and AND2 (N1507, N1503, N462);
xor XOR2 (N1508, N1506, N1108);
buf BUF1 (N1509, N1497);
xor XOR2 (N1510, N1508, N347);
xor XOR2 (N1511, N1507, N82);
xor XOR2 (N1512, N1510, N632);
and AND2 (N1513, N1480, N630);
or OR2 (N1514, N1513, N554);
and AND2 (N1515, N1502, N623);
not NOT1 (N1516, N1494);
buf BUF1 (N1517, N1516);
nand NAND4 (N1518, N1496, N1503, N1077, N43);
not NOT1 (N1519, N1492);
not NOT1 (N1520, N1474);
and AND4 (N1521, N1518, N402, N1453, N516);
nand NAND2 (N1522, N1517, N388);
nand NAND3 (N1523, N1521, N441, N49);
and AND3 (N1524, N1519, N1424, N174);
not NOT1 (N1525, N1523);
xor XOR2 (N1526, N1512, N337);
not NOT1 (N1527, N1524);
or OR2 (N1528, N1526, N1074);
and AND4 (N1529, N1515, N374, N598, N518);
not NOT1 (N1530, N1528);
and AND4 (N1531, N1509, N1048, N424, N680);
and AND2 (N1532, N1525, N527);
nor NOR4 (N1533, N1531, N620, N1397, N824);
xor XOR2 (N1534, N1522, N129);
nor NOR4 (N1535, N1527, N391, N1184, N1188);
or OR4 (N1536, N1535, N1524, N276, N1328);
not NOT1 (N1537, N1520);
nor NOR2 (N1538, N1533, N669);
buf BUF1 (N1539, N1530);
xor XOR2 (N1540, N1534, N1309);
and AND2 (N1541, N1514, N517);
and AND3 (N1542, N1511, N201, N1341);
xor XOR2 (N1543, N1532, N1114);
nand NAND2 (N1544, N1541, N1068);
nand NAND4 (N1545, N1529, N198, N1484, N263);
or OR3 (N1546, N1539, N581, N319);
or OR3 (N1547, N1537, N1052, N633);
nand NAND2 (N1548, N1545, N297);
not NOT1 (N1549, N1536);
and AND4 (N1550, N1538, N314, N273, N128);
buf BUF1 (N1551, N1546);
and AND2 (N1552, N1551, N343);
not NOT1 (N1553, N1544);
and AND3 (N1554, N1547, N283, N487);
or OR4 (N1555, N1550, N529, N995, N286);
xor XOR2 (N1556, N1504, N1259);
or OR4 (N1557, N1556, N917, N1504, N1532);
or OR2 (N1558, N1542, N691);
nand NAND2 (N1559, N1553, N142);
nor NOR2 (N1560, N1548, N1166);
or OR4 (N1561, N1559, N710, N429, N1342);
nor NOR4 (N1562, N1555, N1088, N481, N860);
nor NOR2 (N1563, N1554, N517);
xor XOR2 (N1564, N1557, N602);
and AND4 (N1565, N1558, N1289, N307, N544);
xor XOR2 (N1566, N1563, N459);
nor NOR3 (N1567, N1562, N1499, N352);
and AND2 (N1568, N1540, N119);
and AND2 (N1569, N1564, N854);
buf BUF1 (N1570, N1543);
not NOT1 (N1571, N1561);
nor NOR3 (N1572, N1560, N546, N681);
nor NOR3 (N1573, N1570, N748, N1027);
not NOT1 (N1574, N1572);
and AND4 (N1575, N1573, N1397, N1346, N36);
buf BUF1 (N1576, N1574);
not NOT1 (N1577, N1549);
not NOT1 (N1578, N1577);
nor NOR2 (N1579, N1575, N179);
nor NOR2 (N1580, N1552, N1048);
nor NOR3 (N1581, N1576, N962, N1003);
not NOT1 (N1582, N1578);
and AND3 (N1583, N1567, N26, N1501);
buf BUF1 (N1584, N1571);
not NOT1 (N1585, N1568);
xor XOR2 (N1586, N1582, N791);
nand NAND2 (N1587, N1586, N1449);
buf BUF1 (N1588, N1581);
and AND4 (N1589, N1566, N781, N584, N885);
buf BUF1 (N1590, N1587);
or OR4 (N1591, N1583, N163, N317, N1206);
nand NAND3 (N1592, N1584, N657, N452);
xor XOR2 (N1593, N1591, N175);
and AND2 (N1594, N1565, N175);
not NOT1 (N1595, N1593);
not NOT1 (N1596, N1569);
xor XOR2 (N1597, N1596, N1549);
nand NAND2 (N1598, N1585, N502);
xor XOR2 (N1599, N1589, N361);
nor NOR4 (N1600, N1595, N530, N413, N1096);
and AND2 (N1601, N1580, N282);
nor NOR2 (N1602, N1599, N538);
xor XOR2 (N1603, N1590, N35);
nand NAND3 (N1604, N1588, N131, N377);
buf BUF1 (N1605, N1579);
and AND2 (N1606, N1592, N1134);
buf BUF1 (N1607, N1604);
xor XOR2 (N1608, N1602, N707);
nand NAND2 (N1609, N1601, N802);
buf BUF1 (N1610, N1603);
nand NAND2 (N1611, N1607, N66);
nand NAND3 (N1612, N1606, N1370, N1472);
nand NAND4 (N1613, N1594, N500, N916, N322);
or OR2 (N1614, N1608, N1352);
or OR3 (N1615, N1609, N1110, N833);
nor NOR3 (N1616, N1614, N334, N1234);
xor XOR2 (N1617, N1611, N680);
and AND4 (N1618, N1617, N1540, N415, N370);
not NOT1 (N1619, N1598);
or OR4 (N1620, N1610, N311, N1560, N1559);
nor NOR3 (N1621, N1618, N1403, N1251);
or OR2 (N1622, N1619, N1210);
xor XOR2 (N1623, N1620, N1349);
and AND4 (N1624, N1615, N408, N610, N744);
buf BUF1 (N1625, N1624);
nor NOR2 (N1626, N1597, N1038);
and AND2 (N1627, N1605, N206);
not NOT1 (N1628, N1622);
nor NOR4 (N1629, N1626, N195, N179, N501);
or OR4 (N1630, N1629, N963, N1502, N152);
and AND3 (N1631, N1621, N330, N1214);
nand NAND3 (N1632, N1616, N750, N1586);
or OR2 (N1633, N1628, N357);
nor NOR4 (N1634, N1613, N446, N1268, N1502);
or OR3 (N1635, N1632, N259, N1125);
nand NAND4 (N1636, N1600, N422, N741, N926);
nand NAND2 (N1637, N1635, N868);
not NOT1 (N1638, N1636);
buf BUF1 (N1639, N1612);
not NOT1 (N1640, N1634);
or OR3 (N1641, N1637, N188, N1071);
or OR4 (N1642, N1630, N1187, N704, N174);
nand NAND2 (N1643, N1627, N1172);
buf BUF1 (N1644, N1643);
xor XOR2 (N1645, N1642, N1284);
nand NAND2 (N1646, N1641, N1094);
nor NOR3 (N1647, N1646, N880, N671);
or OR2 (N1648, N1638, N1058);
or OR2 (N1649, N1631, N272);
not NOT1 (N1650, N1647);
or OR3 (N1651, N1649, N592, N828);
not NOT1 (N1652, N1651);
and AND4 (N1653, N1625, N1350, N1522, N749);
buf BUF1 (N1654, N1648);
not NOT1 (N1655, N1650);
nand NAND4 (N1656, N1655, N1609, N1024, N1096);
buf BUF1 (N1657, N1639);
or OR2 (N1658, N1653, N767);
or OR2 (N1659, N1656, N1107);
and AND2 (N1660, N1654, N578);
and AND2 (N1661, N1633, N729);
xor XOR2 (N1662, N1652, N1445);
and AND3 (N1663, N1657, N1550, N624);
and AND3 (N1664, N1663, N1124, N1097);
xor XOR2 (N1665, N1660, N145);
nor NOR3 (N1666, N1645, N1086, N546);
xor XOR2 (N1667, N1665, N450);
nor NOR2 (N1668, N1667, N1602);
and AND2 (N1669, N1662, N104);
nand NAND4 (N1670, N1644, N200, N858, N1592);
nor NOR3 (N1671, N1659, N807, N1348);
not NOT1 (N1672, N1670);
not NOT1 (N1673, N1668);
xor XOR2 (N1674, N1666, N1230);
buf BUF1 (N1675, N1669);
and AND4 (N1676, N1672, N1672, N957, N356);
not NOT1 (N1677, N1664);
buf BUF1 (N1678, N1671);
xor XOR2 (N1679, N1673, N404);
nand NAND4 (N1680, N1674, N1466, N1307, N1323);
and AND4 (N1681, N1640, N1245, N1466, N1110);
buf BUF1 (N1682, N1658);
or OR4 (N1683, N1623, N1317, N1339, N724);
nand NAND2 (N1684, N1679, N1603);
not NOT1 (N1685, N1675);
or OR4 (N1686, N1683, N561, N772, N983);
and AND4 (N1687, N1685, N266, N1632, N1152);
nand NAND3 (N1688, N1684, N944, N1658);
xor XOR2 (N1689, N1678, N468);
nor NOR4 (N1690, N1680, N382, N1416, N663);
and AND4 (N1691, N1681, N376, N265, N1066);
or OR2 (N1692, N1691, N1353);
nor NOR3 (N1693, N1689, N447, N719);
and AND4 (N1694, N1693, N1502, N898, N1208);
not NOT1 (N1695, N1687);
buf BUF1 (N1696, N1661);
and AND3 (N1697, N1677, N623, N1492);
not NOT1 (N1698, N1695);
xor XOR2 (N1699, N1697, N1081);
nand NAND4 (N1700, N1698, N509, N1654, N1190);
and AND3 (N1701, N1700, N62, N1623);
nor NOR4 (N1702, N1699, N348, N1068, N980);
or OR3 (N1703, N1686, N1269, N1244);
xor XOR2 (N1704, N1701, N436);
or OR2 (N1705, N1694, N477);
nor NOR3 (N1706, N1705, N1037, N324);
and AND4 (N1707, N1688, N138, N1263, N1575);
nor NOR3 (N1708, N1702, N371, N57);
nand NAND4 (N1709, N1696, N107, N785, N652);
nand NAND3 (N1710, N1708, N1480, N1031);
or OR4 (N1711, N1710, N1445, N1575, N1696);
xor XOR2 (N1712, N1676, N1707);
xor XOR2 (N1713, N371, N1204);
xor XOR2 (N1714, N1706, N444);
nand NAND2 (N1715, N1704, N766);
or OR4 (N1716, N1715, N1340, N365, N1092);
or OR2 (N1717, N1703, N1565);
buf BUF1 (N1718, N1713);
and AND4 (N1719, N1692, N469, N1290, N341);
not NOT1 (N1720, N1690);
nand NAND3 (N1721, N1719, N1494, N863);
nand NAND2 (N1722, N1716, N44);
and AND3 (N1723, N1721, N146, N736);
buf BUF1 (N1724, N1723);
buf BUF1 (N1725, N1722);
nor NOR3 (N1726, N1682, N792, N375);
buf BUF1 (N1727, N1717);
and AND2 (N1728, N1712, N1512);
xor XOR2 (N1729, N1728, N1165);
nor NOR2 (N1730, N1724, N211);
not NOT1 (N1731, N1725);
xor XOR2 (N1732, N1718, N763);
nor NOR4 (N1733, N1731, N1017, N1174, N722);
nand NAND4 (N1734, N1727, N510, N1584, N823);
nor NOR2 (N1735, N1714, N1446);
and AND2 (N1736, N1735, N531);
or OR2 (N1737, N1736, N483);
nand NAND3 (N1738, N1726, N1477, N711);
or OR4 (N1739, N1730, N961, N925, N1710);
buf BUF1 (N1740, N1733);
and AND3 (N1741, N1738, N1275, N98);
nor NOR2 (N1742, N1737, N694);
xor XOR2 (N1743, N1720, N810);
xor XOR2 (N1744, N1741, N542);
nand NAND4 (N1745, N1740, N960, N983, N1695);
not NOT1 (N1746, N1709);
xor XOR2 (N1747, N1729, N755);
nor NOR2 (N1748, N1732, N408);
not NOT1 (N1749, N1748);
or OR4 (N1750, N1739, N1317, N941, N987);
nand NAND3 (N1751, N1750, N1571, N1094);
nor NOR2 (N1752, N1742, N1695);
buf BUF1 (N1753, N1745);
or OR3 (N1754, N1752, N1185, N701);
and AND3 (N1755, N1753, N1286, N1739);
nand NAND2 (N1756, N1711, N1564);
and AND3 (N1757, N1756, N460, N834);
nor NOR3 (N1758, N1749, N646, N616);
nand NAND3 (N1759, N1743, N189, N1066);
nand NAND3 (N1760, N1751, N650, N506);
nand NAND4 (N1761, N1744, N881, N150, N60);
xor XOR2 (N1762, N1760, N135);
and AND4 (N1763, N1755, N1156, N1408, N1746);
buf BUF1 (N1764, N731);
xor XOR2 (N1765, N1762, N222);
nor NOR3 (N1766, N1764, N1326, N369);
or OR4 (N1767, N1763, N83, N1304, N1609);
xor XOR2 (N1768, N1757, N181);
xor XOR2 (N1769, N1765, N214);
or OR2 (N1770, N1761, N167);
and AND2 (N1771, N1758, N107);
and AND2 (N1772, N1770, N421);
buf BUF1 (N1773, N1766);
and AND4 (N1774, N1734, N57, N371, N1279);
buf BUF1 (N1775, N1747);
or OR3 (N1776, N1769, N1000, N1596);
xor XOR2 (N1777, N1776, N630);
not NOT1 (N1778, N1767);
or OR4 (N1779, N1768, N825, N828, N542);
buf BUF1 (N1780, N1771);
nand NAND3 (N1781, N1779, N299, N1718);
nand NAND2 (N1782, N1780, N984);
nor NOR3 (N1783, N1774, N777, N1434);
nor NOR4 (N1784, N1759, N608, N731, N1202);
xor XOR2 (N1785, N1772, N553);
buf BUF1 (N1786, N1754);
nand NAND2 (N1787, N1782, N211);
xor XOR2 (N1788, N1786, N447);
not NOT1 (N1789, N1784);
nor NOR2 (N1790, N1787, N313);
buf BUF1 (N1791, N1785);
not NOT1 (N1792, N1773);
not NOT1 (N1793, N1778);
buf BUF1 (N1794, N1783);
and AND4 (N1795, N1793, N1115, N1293, N1705);
or OR3 (N1796, N1791, N11, N556);
buf BUF1 (N1797, N1795);
nand NAND4 (N1798, N1796, N204, N1641, N799);
and AND3 (N1799, N1789, N597, N1543);
not NOT1 (N1800, N1790);
nor NOR4 (N1801, N1797, N1127, N127, N573);
buf BUF1 (N1802, N1798);
buf BUF1 (N1803, N1788);
not NOT1 (N1804, N1801);
and AND4 (N1805, N1781, N1368, N148, N1755);
or OR2 (N1806, N1777, N1404);
buf BUF1 (N1807, N1806);
buf BUF1 (N1808, N1804);
not NOT1 (N1809, N1794);
buf BUF1 (N1810, N1809);
buf BUF1 (N1811, N1808);
nand NAND2 (N1812, N1775, N1381);
buf BUF1 (N1813, N1792);
nor NOR3 (N1814, N1805, N1301, N185);
nand NAND2 (N1815, N1812, N529);
xor XOR2 (N1816, N1814, N47);
and AND2 (N1817, N1803, N1477);
xor XOR2 (N1818, N1811, N1341);
xor XOR2 (N1819, N1813, N1517);
buf BUF1 (N1820, N1810);
xor XOR2 (N1821, N1815, N21);
buf BUF1 (N1822, N1821);
nand NAND4 (N1823, N1822, N606, N1733, N642);
or OR3 (N1824, N1816, N48, N426);
nor NOR3 (N1825, N1800, N554, N517);
nand NAND3 (N1826, N1807, N773, N741);
or OR3 (N1827, N1820, N1349, N1525);
buf BUF1 (N1828, N1827);
and AND4 (N1829, N1802, N1061, N33, N158);
not NOT1 (N1830, N1829);
xor XOR2 (N1831, N1828, N1073);
nand NAND2 (N1832, N1817, N1286);
not NOT1 (N1833, N1819);
buf BUF1 (N1834, N1830);
and AND3 (N1835, N1799, N1438, N716);
not NOT1 (N1836, N1835);
or OR2 (N1837, N1818, N478);
xor XOR2 (N1838, N1831, N1325);
xor XOR2 (N1839, N1832, N1492);
xor XOR2 (N1840, N1833, N1201);
and AND4 (N1841, N1825, N1798, N1470, N966);
xor XOR2 (N1842, N1838, N1695);
not NOT1 (N1843, N1840);
nand NAND2 (N1844, N1836, N914);
xor XOR2 (N1845, N1839, N1476);
and AND4 (N1846, N1842, N1011, N745, N84);
or OR2 (N1847, N1823, N823);
buf BUF1 (N1848, N1824);
xor XOR2 (N1849, N1844, N764);
xor XOR2 (N1850, N1841, N1221);
not NOT1 (N1851, N1834);
nor NOR3 (N1852, N1845, N1005, N1465);
nand NAND4 (N1853, N1851, N834, N454, N1332);
nor NOR4 (N1854, N1853, N717, N94, N122);
not NOT1 (N1855, N1854);
or OR3 (N1856, N1850, N159, N762);
or OR4 (N1857, N1847, N202, N248, N190);
and AND3 (N1858, N1826, N1087, N239);
nor NOR2 (N1859, N1852, N616);
buf BUF1 (N1860, N1846);
xor XOR2 (N1861, N1837, N1409);
xor XOR2 (N1862, N1843, N850);
buf BUF1 (N1863, N1860);
or OR4 (N1864, N1861, N576, N795, N40);
not NOT1 (N1865, N1864);
buf BUF1 (N1866, N1855);
xor XOR2 (N1867, N1865, N1335);
and AND4 (N1868, N1859, N593, N1017, N843);
or OR4 (N1869, N1862, N422, N1379, N258);
buf BUF1 (N1870, N1856);
buf BUF1 (N1871, N1849);
buf BUF1 (N1872, N1867);
buf BUF1 (N1873, N1866);
xor XOR2 (N1874, N1848, N619);
and AND3 (N1875, N1870, N1842, N827);
buf BUF1 (N1876, N1863);
and AND2 (N1877, N1869, N725);
nand NAND4 (N1878, N1876, N934, N226, N319);
or OR3 (N1879, N1874, N348, N1033);
not NOT1 (N1880, N1879);
or OR2 (N1881, N1875, N320);
not NOT1 (N1882, N1857);
buf BUF1 (N1883, N1858);
and AND2 (N1884, N1873, N1831);
or OR3 (N1885, N1882, N1410, N1171);
or OR2 (N1886, N1883, N959);
nand NAND4 (N1887, N1877, N1347, N1367, N446);
xor XOR2 (N1888, N1872, N560);
buf BUF1 (N1889, N1885);
buf BUF1 (N1890, N1886);
not NOT1 (N1891, N1888);
or OR2 (N1892, N1871, N552);
or OR4 (N1893, N1889, N756, N862, N564);
not NOT1 (N1894, N1893);
nor NOR2 (N1895, N1881, N641);
and AND4 (N1896, N1887, N1276, N1034, N94);
not NOT1 (N1897, N1894);
or OR2 (N1898, N1880, N916);
or OR2 (N1899, N1895, N406);
and AND4 (N1900, N1897, N1008, N178, N1342);
nand NAND4 (N1901, N1868, N958, N806, N788);
or OR3 (N1902, N1900, N1004, N895);
buf BUF1 (N1903, N1896);
and AND2 (N1904, N1902, N234);
xor XOR2 (N1905, N1899, N1533);
nor NOR4 (N1906, N1884, N745, N1872, N1568);
xor XOR2 (N1907, N1904, N1127);
or OR4 (N1908, N1892, N324, N992, N1040);
and AND2 (N1909, N1906, N1139);
xor XOR2 (N1910, N1908, N1267);
buf BUF1 (N1911, N1898);
not NOT1 (N1912, N1901);
xor XOR2 (N1913, N1907, N1467);
xor XOR2 (N1914, N1911, N206);
not NOT1 (N1915, N1912);
xor XOR2 (N1916, N1913, N175);
xor XOR2 (N1917, N1890, N293);
nor NOR4 (N1918, N1891, N245, N379, N516);
buf BUF1 (N1919, N1916);
buf BUF1 (N1920, N1878);
buf BUF1 (N1921, N1910);
xor XOR2 (N1922, N1903, N1640);
or OR4 (N1923, N1917, N1335, N863, N1265);
nand NAND3 (N1924, N1920, N546, N1667);
xor XOR2 (N1925, N1909, N1152);
xor XOR2 (N1926, N1918, N689);
or OR3 (N1927, N1922, N926, N468);
not NOT1 (N1928, N1921);
xor XOR2 (N1929, N1915, N1189);
not NOT1 (N1930, N1924);
nor NOR3 (N1931, N1923, N1540, N596);
not NOT1 (N1932, N1914);
xor XOR2 (N1933, N1931, N1252);
buf BUF1 (N1934, N1929);
and AND3 (N1935, N1927, N137, N21);
nor NOR4 (N1936, N1930, N861, N1003, N628);
nor NOR3 (N1937, N1934, N1221, N1445);
nand NAND3 (N1938, N1905, N1358, N1688);
nand NAND2 (N1939, N1933, N668);
xor XOR2 (N1940, N1919, N664);
nand NAND4 (N1941, N1937, N1511, N164, N686);
nor NOR4 (N1942, N1925, N922, N421, N1166);
or OR4 (N1943, N1932, N771, N1884, N626);
nor NOR4 (N1944, N1940, N1152, N1303, N1039);
buf BUF1 (N1945, N1936);
nor NOR3 (N1946, N1945, N547, N1760);
nand NAND4 (N1947, N1944, N1811, N601, N1211);
or OR4 (N1948, N1938, N473, N1616, N561);
not NOT1 (N1949, N1926);
nand NAND3 (N1950, N1942, N1398, N236);
and AND4 (N1951, N1946, N1563, N1546, N295);
nor NOR3 (N1952, N1951, N1070, N1634);
or OR2 (N1953, N1952, N828);
or OR3 (N1954, N1943, N632, N1805);
buf BUF1 (N1955, N1948);
or OR2 (N1956, N1954, N417);
nand NAND3 (N1957, N1935, N133, N680);
xor XOR2 (N1958, N1928, N1776);
nand NAND3 (N1959, N1958, N1105, N1502);
and AND4 (N1960, N1941, N1490, N1039, N923);
xor XOR2 (N1961, N1959, N1835);
xor XOR2 (N1962, N1939, N203);
not NOT1 (N1963, N1947);
xor XOR2 (N1964, N1960, N531);
buf BUF1 (N1965, N1955);
xor XOR2 (N1966, N1949, N1723);
or OR2 (N1967, N1966, N997);
not NOT1 (N1968, N1957);
buf BUF1 (N1969, N1953);
buf BUF1 (N1970, N1962);
and AND2 (N1971, N1967, N1620);
nor NOR3 (N1972, N1956, N469, N1174);
or OR3 (N1973, N1950, N1310, N1585);
and AND3 (N1974, N1965, N687, N1790);
buf BUF1 (N1975, N1968);
nand NAND4 (N1976, N1974, N1913, N236, N1818);
and AND2 (N1977, N1963, N394);
buf BUF1 (N1978, N1972);
xor XOR2 (N1979, N1973, N286);
not NOT1 (N1980, N1961);
and AND3 (N1981, N1980, N502, N1554);
nand NAND3 (N1982, N1976, N770, N1570);
or OR4 (N1983, N1975, N552, N1189, N1904);
not NOT1 (N1984, N1982);
nor NOR2 (N1985, N1981, N1457);
not NOT1 (N1986, N1970);
nor NOR2 (N1987, N1984, N1050);
not NOT1 (N1988, N1969);
or OR4 (N1989, N1987, N783, N463, N457);
nand NAND2 (N1990, N1989, N932);
buf BUF1 (N1991, N1977);
not NOT1 (N1992, N1991);
nor NOR2 (N1993, N1971, N1424);
and AND2 (N1994, N1983, N1170);
and AND2 (N1995, N1985, N1840);
nor NOR2 (N1996, N1986, N223);
nand NAND4 (N1997, N1995, N213, N388, N1792);
and AND3 (N1998, N1988, N1890, N795);
buf BUF1 (N1999, N1998);
and AND3 (N2000, N1992, N971, N1357);
buf BUF1 (N2001, N1990);
xor XOR2 (N2002, N1993, N1080);
or OR3 (N2003, N1978, N903, N1183);
xor XOR2 (N2004, N2000, N639);
or OR4 (N2005, N2004, N1983, N143, N466);
nand NAND4 (N2006, N1979, N642, N1493, N954);
or OR2 (N2007, N1999, N426);
or OR2 (N2008, N1997, N695);
buf BUF1 (N2009, N2006);
xor XOR2 (N2010, N2001, N513);
nor NOR2 (N2011, N2007, N185);
not NOT1 (N2012, N2011);
xor XOR2 (N2013, N2009, N853);
buf BUF1 (N2014, N2008);
xor XOR2 (N2015, N2005, N1764);
and AND2 (N2016, N1994, N849);
xor XOR2 (N2017, N2014, N741);
buf BUF1 (N2018, N2012);
nor NOR2 (N2019, N2017, N1198);
buf BUF1 (N2020, N2002);
and AND4 (N2021, N1996, N449, N252, N1289);
not NOT1 (N2022, N2013);
or OR3 (N2023, N2019, N1691, N197);
or OR2 (N2024, N2016, N1596);
xor XOR2 (N2025, N2023, N1605);
buf BUF1 (N2026, N2025);
nand NAND4 (N2027, N2026, N257, N160, N267);
xor XOR2 (N2028, N2020, N756);
not NOT1 (N2029, N2015);
or OR3 (N2030, N2028, N751, N1322);
nand NAND3 (N2031, N2022, N1788, N1612);
xor XOR2 (N2032, N2029, N894);
or OR2 (N2033, N2021, N895);
and AND4 (N2034, N2033, N400, N1679, N1982);
nand NAND3 (N2035, N2027, N188, N1255);
and AND3 (N2036, N2010, N806, N306);
xor XOR2 (N2037, N2024, N2000);
nor NOR3 (N2038, N2037, N970, N1246);
xor XOR2 (N2039, N2018, N1301);
not NOT1 (N2040, N2003);
buf BUF1 (N2041, N2040);
or OR4 (N2042, N2031, N719, N70, N1919);
or OR2 (N2043, N2039, N1363);
not NOT1 (N2044, N2043);
nor NOR2 (N2045, N2030, N2015);
nand NAND3 (N2046, N1964, N1282, N398);
nand NAND2 (N2047, N2041, N475);
not NOT1 (N2048, N2047);
and AND4 (N2049, N2042, N595, N343, N2036);
xor XOR2 (N2050, N456, N220);
not NOT1 (N2051, N2034);
or OR2 (N2052, N2051, N744);
not NOT1 (N2053, N2044);
not NOT1 (N2054, N2050);
xor XOR2 (N2055, N2053, N844);
and AND3 (N2056, N2032, N38, N981);
nor NOR4 (N2057, N2045, N988, N1343, N542);
not NOT1 (N2058, N2054);
nor NOR3 (N2059, N2049, N1961, N941);
nand NAND4 (N2060, N2048, N1334, N1026, N1126);
buf BUF1 (N2061, N2046);
nor NOR3 (N2062, N2055, N1893, N1496);
and AND2 (N2063, N2062, N961);
not NOT1 (N2064, N2057);
nor NOR4 (N2065, N2035, N1340, N719, N576);
buf BUF1 (N2066, N2063);
and AND4 (N2067, N2059, N1455, N329, N805);
or OR2 (N2068, N2061, N240);
buf BUF1 (N2069, N2064);
nand NAND3 (N2070, N2056, N1658, N305);
nor NOR3 (N2071, N2052, N1736, N615);
nor NOR3 (N2072, N2068, N1851, N322);
or OR2 (N2073, N2066, N626);
or OR4 (N2074, N2060, N1728, N1686, N304);
buf BUF1 (N2075, N2038);
xor XOR2 (N2076, N2058, N35);
or OR4 (N2077, N2072, N1462, N1364, N1801);
or OR2 (N2078, N2069, N1560);
nor NOR3 (N2079, N2074, N1078, N1885);
and AND4 (N2080, N2070, N679, N590, N20);
buf BUF1 (N2081, N2078);
and AND4 (N2082, N2073, N202, N1428, N1936);
nand NAND4 (N2083, N2081, N1527, N53, N1409);
or OR3 (N2084, N2079, N1881, N110);
or OR2 (N2085, N2084, N234);
nand NAND4 (N2086, N2082, N1928, N1902, N974);
and AND4 (N2087, N2076, N270, N230, N898);
buf BUF1 (N2088, N2065);
nor NOR2 (N2089, N2087, N747);
not NOT1 (N2090, N2067);
not NOT1 (N2091, N2089);
not NOT1 (N2092, N2071);
xor XOR2 (N2093, N2085, N1350);
or OR3 (N2094, N2075, N1546, N1857);
nand NAND2 (N2095, N2092, N2069);
nor NOR3 (N2096, N2094, N1347, N1963);
and AND4 (N2097, N2088, N462, N392, N1476);
and AND4 (N2098, N2090, N1933, N2016, N1763);
not NOT1 (N2099, N2091);
xor XOR2 (N2100, N2096, N1465);
xor XOR2 (N2101, N2099, N450);
and AND2 (N2102, N2086, N1335);
or OR3 (N2103, N2102, N648, N162);
buf BUF1 (N2104, N2093);
and AND2 (N2105, N2104, N1643);
xor XOR2 (N2106, N2100, N371);
not NOT1 (N2107, N2105);
and AND4 (N2108, N2107, N1541, N649, N1677);
and AND3 (N2109, N2106, N1600, N83);
and AND3 (N2110, N2077, N994, N1180);
or OR4 (N2111, N2098, N973, N749, N563);
nor NOR4 (N2112, N2083, N339, N702, N378);
xor XOR2 (N2113, N2101, N636);
xor XOR2 (N2114, N2110, N798);
and AND3 (N2115, N2108, N678, N127);
xor XOR2 (N2116, N2103, N559);
buf BUF1 (N2117, N2097);
or OR3 (N2118, N2114, N1226, N2049);
and AND4 (N2119, N2115, N1619, N1469, N1654);
and AND3 (N2120, N2119, N717, N963);
xor XOR2 (N2121, N2109, N223);
nand NAND4 (N2122, N2080, N1542, N920, N1856);
not NOT1 (N2123, N2112);
nand NAND3 (N2124, N2117, N1536, N1726);
not NOT1 (N2125, N2118);
nand NAND4 (N2126, N2121, N175, N197, N2086);
or OR3 (N2127, N2116, N1194, N435);
nand NAND4 (N2128, N2111, N1048, N925, N192);
or OR3 (N2129, N2120, N2050, N489);
buf BUF1 (N2130, N2124);
buf BUF1 (N2131, N2113);
xor XOR2 (N2132, N2095, N513);
nor NOR4 (N2133, N2122, N572, N352, N441);
nor NOR4 (N2134, N2128, N284, N707, N1525);
buf BUF1 (N2135, N2134);
xor XOR2 (N2136, N2131, N161);
not NOT1 (N2137, N2123);
and AND4 (N2138, N2129, N1666, N1439, N1698);
or OR2 (N2139, N2132, N1217);
xor XOR2 (N2140, N2126, N718);
or OR4 (N2141, N2130, N249, N410, N271);
not NOT1 (N2142, N2133);
or OR2 (N2143, N2136, N687);
or OR4 (N2144, N2142, N685, N516, N282);
not NOT1 (N2145, N2127);
nor NOR2 (N2146, N2143, N15);
buf BUF1 (N2147, N2138);
nand NAND2 (N2148, N2140, N664);
and AND3 (N2149, N2137, N1386, N432);
nor NOR2 (N2150, N2141, N712);
or OR2 (N2151, N2125, N1885);
nor NOR2 (N2152, N2145, N1728);
nand NAND2 (N2153, N2144, N2034);
not NOT1 (N2154, N2148);
nand NAND3 (N2155, N2153, N736, N1235);
not NOT1 (N2156, N2146);
not NOT1 (N2157, N2150);
nor NOR4 (N2158, N2135, N1397, N1817, N645);
not NOT1 (N2159, N2149);
not NOT1 (N2160, N2139);
nor NOR4 (N2161, N2160, N1301, N344, N1517);
and AND3 (N2162, N2157, N1208, N486);
nor NOR3 (N2163, N2159, N1462, N166);
buf BUF1 (N2164, N2161);
or OR2 (N2165, N2155, N1187);
not NOT1 (N2166, N2158);
nand NAND3 (N2167, N2156, N1303, N1702);
nand NAND3 (N2168, N2167, N577, N523);
xor XOR2 (N2169, N2168, N365);
nor NOR3 (N2170, N2154, N684, N1860);
xor XOR2 (N2171, N2166, N1664);
or OR2 (N2172, N2152, N744);
and AND3 (N2173, N2164, N11, N709);
nor NOR3 (N2174, N2170, N880, N858);
and AND2 (N2175, N2147, N1463);
buf BUF1 (N2176, N2169);
not NOT1 (N2177, N2165);
nor NOR4 (N2178, N2173, N1685, N1367, N141);
or OR2 (N2179, N2174, N1756);
xor XOR2 (N2180, N2162, N1709);
buf BUF1 (N2181, N2172);
buf BUF1 (N2182, N2181);
xor XOR2 (N2183, N2178, N2075);
and AND3 (N2184, N2177, N1568, N1428);
nand NAND4 (N2185, N2171, N338, N1691, N1452);
nand NAND4 (N2186, N2180, N169, N45, N874);
xor XOR2 (N2187, N2186, N1186);
xor XOR2 (N2188, N2163, N574);
and AND2 (N2189, N2184, N1670);
or OR2 (N2190, N2179, N848);
buf BUF1 (N2191, N2188);
nor NOR3 (N2192, N2185, N1931, N1551);
nor NOR3 (N2193, N2192, N1889, N801);
nor NOR3 (N2194, N2193, N1637, N880);
not NOT1 (N2195, N2176);
not NOT1 (N2196, N2151);
xor XOR2 (N2197, N2191, N1969);
xor XOR2 (N2198, N2197, N1442);
or OR2 (N2199, N2189, N1301);
xor XOR2 (N2200, N2195, N962);
and AND3 (N2201, N2182, N1067, N520);
not NOT1 (N2202, N2196);
and AND3 (N2203, N2190, N1628, N1367);
buf BUF1 (N2204, N2198);
buf BUF1 (N2205, N2201);
nor NOR3 (N2206, N2194, N499, N1037);
nor NOR3 (N2207, N2199, N408, N292);
buf BUF1 (N2208, N2206);
nor NOR2 (N2209, N2175, N1083);
or OR3 (N2210, N2200, N524, N1952);
not NOT1 (N2211, N2207);
buf BUF1 (N2212, N2187);
nor NOR4 (N2213, N2209, N2035, N2190, N1724);
nor NOR2 (N2214, N2208, N246);
or OR3 (N2215, N2203, N986, N26);
nand NAND2 (N2216, N2213, N1003);
xor XOR2 (N2217, N2210, N165);
and AND2 (N2218, N2214, N271);
nor NOR2 (N2219, N2204, N1107);
nand NAND4 (N2220, N2215, N1130, N843, N589);
nor NOR3 (N2221, N2212, N711, N471);
or OR4 (N2222, N2183, N1327, N530, N933);
buf BUF1 (N2223, N2202);
xor XOR2 (N2224, N2220, N1937);
nor NOR4 (N2225, N2223, N1527, N252, N199);
xor XOR2 (N2226, N2221, N418);
nand NAND2 (N2227, N2205, N1325);
xor XOR2 (N2228, N2227, N1974);
and AND2 (N2229, N2216, N816);
xor XOR2 (N2230, N2218, N510);
nand NAND3 (N2231, N2226, N120, N799);
nand NAND2 (N2232, N2225, N613);
nand NAND3 (N2233, N2224, N338, N1695);
xor XOR2 (N2234, N2229, N1136);
xor XOR2 (N2235, N2234, N775);
or OR3 (N2236, N2228, N357, N738);
nand NAND2 (N2237, N2231, N1062);
buf BUF1 (N2238, N2235);
xor XOR2 (N2239, N2238, N328);
nand NAND4 (N2240, N2219, N314, N565, N1650);
nand NAND4 (N2241, N2240, N1752, N2141, N1755);
buf BUF1 (N2242, N2233);
and AND3 (N2243, N2211, N384, N1835);
not NOT1 (N2244, N2222);
nand NAND3 (N2245, N2232, N408, N1977);
xor XOR2 (N2246, N2243, N297);
or OR2 (N2247, N2245, N273);
xor XOR2 (N2248, N2236, N382);
buf BUF1 (N2249, N2241);
nand NAND4 (N2250, N2217, N1249, N1634, N2213);
and AND2 (N2251, N2244, N1919);
buf BUF1 (N2252, N2250);
buf BUF1 (N2253, N2251);
nand NAND3 (N2254, N2247, N617, N1896);
nor NOR3 (N2255, N2254, N949, N1646);
xor XOR2 (N2256, N2239, N109);
buf BUF1 (N2257, N2242);
xor XOR2 (N2258, N2237, N2060);
and AND4 (N2259, N2258, N2223, N2138, N2227);
nor NOR4 (N2260, N2249, N560, N2073, N609);
buf BUF1 (N2261, N2230);
buf BUF1 (N2262, N2257);
nor NOR3 (N2263, N2246, N1540, N244);
buf BUF1 (N2264, N2262);
nand NAND3 (N2265, N2259, N361, N860);
nor NOR3 (N2266, N2253, N1533, N890);
not NOT1 (N2267, N2261);
and AND2 (N2268, N2256, N416);
not NOT1 (N2269, N2264);
nand NAND3 (N2270, N2266, N956, N1173);
not NOT1 (N2271, N2269);
and AND3 (N2272, N2270, N783, N538);
nor NOR4 (N2273, N2271, N276, N1954, N341);
buf BUF1 (N2274, N2272);
xor XOR2 (N2275, N2255, N568);
and AND4 (N2276, N2273, N1127, N375, N1432);
not NOT1 (N2277, N2274);
buf BUF1 (N2278, N2248);
nor NOR4 (N2279, N2265, N979, N1930, N197);
or OR3 (N2280, N2267, N1637, N2259);
or OR3 (N2281, N2276, N1320, N902);
buf BUF1 (N2282, N2281);
and AND2 (N2283, N2278, N1662);
buf BUF1 (N2284, N2260);
not NOT1 (N2285, N2277);
nor NOR3 (N2286, N2279, N829, N310);
buf BUF1 (N2287, N2284);
not NOT1 (N2288, N2287);
xor XOR2 (N2289, N2263, N641);
xor XOR2 (N2290, N2282, N711);
and AND2 (N2291, N2275, N1940);
xor XOR2 (N2292, N2280, N135);
xor XOR2 (N2293, N2288, N1375);
buf BUF1 (N2294, N2293);
not NOT1 (N2295, N2268);
nand NAND4 (N2296, N2285, N1675, N532, N2089);
not NOT1 (N2297, N2290);
xor XOR2 (N2298, N2295, N945);
xor XOR2 (N2299, N2252, N1552);
buf BUF1 (N2300, N2296);
buf BUF1 (N2301, N2298);
not NOT1 (N2302, N2294);
and AND2 (N2303, N2301, N524);
nand NAND4 (N2304, N2300, N763, N927, N530);
buf BUF1 (N2305, N2291);
nor NOR3 (N2306, N2289, N1229, N1124);
buf BUF1 (N2307, N2303);
not NOT1 (N2308, N2302);
and AND4 (N2309, N2286, N547, N2121, N1850);
xor XOR2 (N2310, N2283, N1887);
nand NAND4 (N2311, N2297, N1465, N1625, N748);
nor NOR2 (N2312, N2306, N554);
and AND3 (N2313, N2309, N2265, N2079);
and AND3 (N2314, N2313, N156, N1373);
not NOT1 (N2315, N2307);
not NOT1 (N2316, N2299);
xor XOR2 (N2317, N2310, N1874);
and AND4 (N2318, N2314, N40, N450, N198);
xor XOR2 (N2319, N2308, N1544);
or OR2 (N2320, N2317, N2004);
xor XOR2 (N2321, N2304, N412);
or OR4 (N2322, N2320, N836, N998, N891);
nor NOR4 (N2323, N2321, N1194, N324, N1833);
xor XOR2 (N2324, N2311, N1276);
nand NAND2 (N2325, N2318, N691);
nand NAND2 (N2326, N2323, N1235);
nor NOR2 (N2327, N2324, N1686);
or OR3 (N2328, N2292, N616, N992);
nor NOR2 (N2329, N2328, N1219);
not NOT1 (N2330, N2326);
not NOT1 (N2331, N2319);
not NOT1 (N2332, N2327);
not NOT1 (N2333, N2331);
nand NAND4 (N2334, N2312, N1445, N1239, N1729);
and AND2 (N2335, N2332, N1278);
and AND2 (N2336, N2334, N95);
xor XOR2 (N2337, N2336, N1712);
nor NOR2 (N2338, N2337, N1705);
or OR3 (N2339, N2315, N1741, N90);
buf BUF1 (N2340, N2339);
buf BUF1 (N2341, N2330);
not NOT1 (N2342, N2316);
nand NAND4 (N2343, N2325, N1430, N1171, N2269);
not NOT1 (N2344, N2341);
not NOT1 (N2345, N2344);
or OR3 (N2346, N2345, N1108, N485);
nand NAND2 (N2347, N2322, N687);
and AND3 (N2348, N2342, N616, N2263);
nor NOR3 (N2349, N2343, N1204, N2007);
not NOT1 (N2350, N2335);
or OR4 (N2351, N2329, N505, N699, N2060);
or OR2 (N2352, N2348, N2018);
buf BUF1 (N2353, N2347);
nor NOR4 (N2354, N2353, N1947, N1317, N1050);
nor NOR2 (N2355, N2346, N739);
not NOT1 (N2356, N2352);
xor XOR2 (N2357, N2305, N1553);
and AND2 (N2358, N2333, N240);
not NOT1 (N2359, N2357);
or OR3 (N2360, N2349, N1606, N76);
nor NOR2 (N2361, N2350, N1934);
nor NOR4 (N2362, N2361, N1259, N466, N1720);
nor NOR2 (N2363, N2356, N1178);
and AND4 (N2364, N2351, N1607, N227, N1685);
not NOT1 (N2365, N2355);
not NOT1 (N2366, N2360);
nand NAND4 (N2367, N2359, N2174, N1480, N249);
not NOT1 (N2368, N2358);
nand NAND3 (N2369, N2365, N29, N1521);
nand NAND2 (N2370, N2340, N1977);
xor XOR2 (N2371, N2338, N2349);
nand NAND2 (N2372, N2366, N179);
or OR2 (N2373, N2371, N1772);
not NOT1 (N2374, N2370);
nor NOR3 (N2375, N2368, N1691, N245);
or OR2 (N2376, N2369, N335);
buf BUF1 (N2377, N2374);
and AND3 (N2378, N2377, N2323, N978);
nor NOR3 (N2379, N2375, N1788, N1194);
nand NAND2 (N2380, N2362, N2021);
nand NAND4 (N2381, N2380, N2046, N2103, N1427);
buf BUF1 (N2382, N2376);
nor NOR3 (N2383, N2367, N1299, N1918);
and AND2 (N2384, N2382, N334);
and AND4 (N2385, N2373, N1981, N1599, N351);
or OR3 (N2386, N2381, N1660, N1249);
not NOT1 (N2387, N2385);
not NOT1 (N2388, N2354);
and AND3 (N2389, N2386, N1911, N2154);
nand NAND4 (N2390, N2379, N1367, N2221, N1224);
nor NOR2 (N2391, N2387, N490);
xor XOR2 (N2392, N2363, N549);
nor NOR2 (N2393, N2372, N1405);
or OR4 (N2394, N2393, N565, N495, N409);
and AND4 (N2395, N2389, N1529, N1169, N373);
xor XOR2 (N2396, N2392, N1143);
or OR4 (N2397, N2391, N1883, N1080, N404);
or OR3 (N2398, N2395, N2287, N976);
nand NAND2 (N2399, N2398, N2123);
xor XOR2 (N2400, N2378, N231);
nor NOR3 (N2401, N2396, N253, N1692);
buf BUF1 (N2402, N2388);
xor XOR2 (N2403, N2364, N1561);
buf BUF1 (N2404, N2401);
and AND3 (N2405, N2403, N505, N1331);
nor NOR3 (N2406, N2384, N1908, N641);
buf BUF1 (N2407, N2406);
xor XOR2 (N2408, N2407, N1927);
buf BUF1 (N2409, N2397);
not NOT1 (N2410, N2399);
buf BUF1 (N2411, N2402);
nor NOR4 (N2412, N2410, N166, N2228, N223);
or OR2 (N2413, N2409, N1779);
not NOT1 (N2414, N2400);
not NOT1 (N2415, N2413);
nor NOR2 (N2416, N2390, N1635);
nor NOR3 (N2417, N2383, N1682, N1668);
xor XOR2 (N2418, N2411, N614);
buf BUF1 (N2419, N2416);
nand NAND2 (N2420, N2418, N1794);
nor NOR4 (N2421, N2420, N1765, N168, N1219);
not NOT1 (N2422, N2414);
and AND3 (N2423, N2408, N219, N281);
and AND3 (N2424, N2405, N130, N660);
xor XOR2 (N2425, N2424, N1175);
nor NOR2 (N2426, N2394, N488);
not NOT1 (N2427, N2426);
xor XOR2 (N2428, N2417, N833);
or OR4 (N2429, N2412, N558, N1239, N1317);
not NOT1 (N2430, N2415);
buf BUF1 (N2431, N2421);
xor XOR2 (N2432, N2430, N488);
buf BUF1 (N2433, N2404);
nor NOR4 (N2434, N2428, N773, N385, N387);
nor NOR2 (N2435, N2433, N709);
xor XOR2 (N2436, N2429, N1947);
nor NOR3 (N2437, N2434, N1669, N1743);
nor NOR4 (N2438, N2437, N1084, N544, N432);
and AND3 (N2439, N2427, N1426, N1376);
nand NAND3 (N2440, N2435, N2018, N1383);
buf BUF1 (N2441, N2440);
nor NOR3 (N2442, N2438, N1444, N190);
and AND4 (N2443, N2425, N1806, N1848, N1333);
buf BUF1 (N2444, N2442);
and AND3 (N2445, N2441, N257, N313);
nor NOR2 (N2446, N2439, N1167);
and AND3 (N2447, N2445, N292, N1744);
and AND3 (N2448, N2423, N2425, N1813);
xor XOR2 (N2449, N2436, N202);
xor XOR2 (N2450, N2446, N970);
buf BUF1 (N2451, N2450);
nor NOR3 (N2452, N2449, N47, N2154);
nor NOR2 (N2453, N2432, N337);
buf BUF1 (N2454, N2431);
nand NAND3 (N2455, N2447, N354, N1850);
or OR4 (N2456, N2454, N1793, N1143, N1158);
and AND3 (N2457, N2422, N1747, N2332);
and AND4 (N2458, N2419, N1613, N1331, N1975);
nor NOR4 (N2459, N2444, N1200, N1207, N2024);
nor NOR3 (N2460, N2451, N658, N2449);
not NOT1 (N2461, N2448);
nand NAND2 (N2462, N2460, N1670);
xor XOR2 (N2463, N2458, N1858);
xor XOR2 (N2464, N2456, N1532);
not NOT1 (N2465, N2463);
buf BUF1 (N2466, N2455);
not NOT1 (N2467, N2466);
not NOT1 (N2468, N2453);
xor XOR2 (N2469, N2465, N1768);
nor NOR3 (N2470, N2468, N95, N1505);
xor XOR2 (N2471, N2461, N61);
and AND3 (N2472, N2464, N2406, N1854);
and AND4 (N2473, N2452, N1772, N367, N721);
buf BUF1 (N2474, N2467);
nor NOR3 (N2475, N2473, N730, N295);
not NOT1 (N2476, N2474);
and AND2 (N2477, N2443, N2444);
and AND2 (N2478, N2476, N774);
not NOT1 (N2479, N2469);
buf BUF1 (N2480, N2462);
xor XOR2 (N2481, N2480, N1877);
and AND4 (N2482, N2475, N1332, N1894, N1586);
not NOT1 (N2483, N2471);
and AND2 (N2484, N2481, N2007);
not NOT1 (N2485, N2459);
nor NOR4 (N2486, N2482, N1556, N1412, N1811);
nand NAND2 (N2487, N2470, N1897);
nand NAND2 (N2488, N2485, N1319);
nand NAND4 (N2489, N2477, N1721, N65, N2448);
and AND2 (N2490, N2484, N2242);
or OR2 (N2491, N2479, N1254);
buf BUF1 (N2492, N2488);
or OR3 (N2493, N2490, N708, N1180);
xor XOR2 (N2494, N2487, N549);
and AND4 (N2495, N2494, N92, N1889, N730);
nand NAND2 (N2496, N2457, N1956);
xor XOR2 (N2497, N2495, N624);
xor XOR2 (N2498, N2491, N492);
or OR3 (N2499, N2483, N1901, N1509);
or OR2 (N2500, N2499, N2111);
or OR4 (N2501, N2492, N1967, N246, N1243);
xor XOR2 (N2502, N2496, N1260);
xor XOR2 (N2503, N2472, N2259);
buf BUF1 (N2504, N2498);
not NOT1 (N2505, N2486);
xor XOR2 (N2506, N2501, N966);
and AND2 (N2507, N2504, N1691);
nor NOR3 (N2508, N2500, N1222, N1595);
xor XOR2 (N2509, N2497, N1656);
and AND2 (N2510, N2489, N940);
not NOT1 (N2511, N2509);
and AND4 (N2512, N2493, N547, N1276, N396);
buf BUF1 (N2513, N2507);
or OR3 (N2514, N2506, N725, N1045);
nor NOR3 (N2515, N2503, N719, N583);
or OR2 (N2516, N2505, N1714);
not NOT1 (N2517, N2516);
xor XOR2 (N2518, N2502, N2269);
nor NOR2 (N2519, N2518, N2277);
and AND2 (N2520, N2519, N2203);
and AND3 (N2521, N2514, N1509, N74);
not NOT1 (N2522, N2511);
nand NAND4 (N2523, N2515, N2342, N1733, N216);
or OR3 (N2524, N2521, N40, N1363);
and AND4 (N2525, N2524, N1674, N1882, N872);
not NOT1 (N2526, N2510);
xor XOR2 (N2527, N2525, N558);
and AND4 (N2528, N2508, N98, N1919, N2454);
and AND2 (N2529, N2520, N2126);
not NOT1 (N2530, N2528);
not NOT1 (N2531, N2529);
and AND3 (N2532, N2523, N2377, N2383);
not NOT1 (N2533, N2527);
and AND3 (N2534, N2533, N820, N1459);
and AND4 (N2535, N2513, N555, N479, N2157);
not NOT1 (N2536, N2526);
buf BUF1 (N2537, N2536);
or OR3 (N2538, N2537, N1069, N1145);
xor XOR2 (N2539, N2534, N443);
or OR2 (N2540, N2512, N2340);
or OR4 (N2541, N2522, N1194, N1780, N1962);
and AND3 (N2542, N2517, N119, N1160);
xor XOR2 (N2543, N2532, N1250);
not NOT1 (N2544, N2541);
nor NOR4 (N2545, N2544, N2411, N2115, N728);
or OR4 (N2546, N2538, N2450, N634, N605);
buf BUF1 (N2547, N2545);
and AND3 (N2548, N2546, N1406, N1017);
and AND2 (N2549, N2547, N849);
xor XOR2 (N2550, N2530, N1700);
nand NAND4 (N2551, N2535, N57, N821, N1138);
or OR2 (N2552, N2550, N42);
buf BUF1 (N2553, N2542);
buf BUF1 (N2554, N2531);
not NOT1 (N2555, N2552);
xor XOR2 (N2556, N2549, N597);
and AND2 (N2557, N2556, N214);
nand NAND2 (N2558, N2540, N1870);
and AND4 (N2559, N2553, N484, N1991, N2359);
and AND2 (N2560, N2548, N1512);
nor NOR3 (N2561, N2543, N1125, N1528);
and AND3 (N2562, N2560, N2095, N1904);
xor XOR2 (N2563, N2559, N683);
nand NAND4 (N2564, N2478, N1225, N234, N302);
buf BUF1 (N2565, N2539);
buf BUF1 (N2566, N2555);
or OR2 (N2567, N2558, N731);
nor NOR2 (N2568, N2563, N1022);
and AND4 (N2569, N2566, N692, N1483, N507);
nor NOR4 (N2570, N2554, N248, N2203, N337);
and AND3 (N2571, N2569, N2096, N2215);
and AND4 (N2572, N2561, N2433, N1653, N90);
nand NAND4 (N2573, N2571, N1887, N1292, N1935);
xor XOR2 (N2574, N2572, N2193);
xor XOR2 (N2575, N2562, N1677);
nand NAND2 (N2576, N2567, N2362);
xor XOR2 (N2577, N2557, N2068);
and AND2 (N2578, N2564, N198);
xor XOR2 (N2579, N2575, N1953);
not NOT1 (N2580, N2579);
nor NOR3 (N2581, N2570, N434, N1979);
or OR3 (N2582, N2581, N2344, N2166);
or OR3 (N2583, N2576, N1547, N659);
not NOT1 (N2584, N2582);
buf BUF1 (N2585, N2565);
nand NAND4 (N2586, N2583, N2084, N122, N302);
xor XOR2 (N2587, N2584, N405);
not NOT1 (N2588, N2568);
buf BUF1 (N2589, N2578);
or OR3 (N2590, N2574, N126, N53);
not NOT1 (N2591, N2577);
xor XOR2 (N2592, N2586, N2358);
nand NAND4 (N2593, N2585, N1358, N1991, N797);
nand NAND3 (N2594, N2573, N618, N2475);
or OR2 (N2595, N2589, N226);
nand NAND4 (N2596, N2592, N1746, N2232, N871);
and AND3 (N2597, N2580, N2236, N1650);
or OR3 (N2598, N2596, N2354, N221);
buf BUF1 (N2599, N2590);
and AND4 (N2600, N2588, N1194, N429, N767);
nand NAND2 (N2601, N2600, N356);
xor XOR2 (N2602, N2598, N1657);
not NOT1 (N2603, N2594);
and AND2 (N2604, N2595, N2245);
nand NAND2 (N2605, N2593, N707);
nor NOR4 (N2606, N2602, N757, N2076, N1631);
xor XOR2 (N2607, N2606, N483);
or OR3 (N2608, N2591, N2300, N575);
not NOT1 (N2609, N2601);
or OR4 (N2610, N2607, N1934, N1857, N1316);
not NOT1 (N2611, N2608);
not NOT1 (N2612, N2551);
and AND4 (N2613, N2604, N2367, N430, N2083);
or OR3 (N2614, N2609, N26, N1581);
and AND2 (N2615, N2597, N335);
not NOT1 (N2616, N2605);
not NOT1 (N2617, N2616);
nand NAND3 (N2618, N2614, N1101, N1829);
buf BUF1 (N2619, N2615);
nor NOR4 (N2620, N2610, N2200, N961, N927);
and AND2 (N2621, N2619, N358);
and AND4 (N2622, N2603, N1062, N2003, N1687);
nor NOR4 (N2623, N2618, N2253, N18, N1771);
nand NAND2 (N2624, N2587, N1576);
or OR4 (N2625, N2613, N823, N1443, N2506);
buf BUF1 (N2626, N2622);
buf BUF1 (N2627, N2599);
nand NAND3 (N2628, N2623, N57, N1993);
nand NAND2 (N2629, N2628, N583);
nor NOR4 (N2630, N2611, N2324, N2102, N1909);
or OR4 (N2631, N2612, N455, N212, N2494);
xor XOR2 (N2632, N2624, N2550);
not NOT1 (N2633, N2630);
or OR3 (N2634, N2626, N960, N1685);
xor XOR2 (N2635, N2617, N2401);
nand NAND2 (N2636, N2629, N2341);
nand NAND3 (N2637, N2634, N2536, N850);
and AND2 (N2638, N2637, N2146);
xor XOR2 (N2639, N2635, N1128);
and AND3 (N2640, N2639, N1748, N2616);
nand NAND2 (N2641, N2638, N1187);
nor NOR3 (N2642, N2636, N1563, N11);
nor NOR3 (N2643, N2620, N2044, N1626);
or OR2 (N2644, N2625, N949);
buf BUF1 (N2645, N2633);
nor NOR4 (N2646, N2621, N2001, N2552, N2291);
xor XOR2 (N2647, N2646, N1505);
xor XOR2 (N2648, N2632, N2033);
xor XOR2 (N2649, N2627, N816);
or OR3 (N2650, N2643, N1277, N921);
nand NAND2 (N2651, N2631, N1623);
or OR4 (N2652, N2651, N1645, N1492, N1795);
nand NAND3 (N2653, N2642, N435, N1805);
and AND3 (N2654, N2645, N431, N2653);
xor XOR2 (N2655, N157, N2156);
xor XOR2 (N2656, N2652, N817);
not NOT1 (N2657, N2648);
xor XOR2 (N2658, N2641, N1760);
not NOT1 (N2659, N2656);
or OR2 (N2660, N2655, N937);
nand NAND2 (N2661, N2657, N60);
nor NOR3 (N2662, N2659, N1740, N275);
nor NOR2 (N2663, N2650, N1242);
or OR2 (N2664, N2640, N272);
xor XOR2 (N2665, N2663, N64);
xor XOR2 (N2666, N2664, N735);
nand NAND4 (N2667, N2665, N857, N2051, N1126);
not NOT1 (N2668, N2654);
xor XOR2 (N2669, N2668, N1690);
or OR2 (N2670, N2658, N492);
nor NOR3 (N2671, N2647, N1270, N1329);
buf BUF1 (N2672, N2644);
nand NAND4 (N2673, N2666, N256, N1080, N136);
not NOT1 (N2674, N2661);
or OR4 (N2675, N2674, N1830, N1145, N2638);
or OR2 (N2676, N2669, N765);
or OR2 (N2677, N2672, N486);
not NOT1 (N2678, N2671);
or OR3 (N2679, N2678, N1298, N1330);
not NOT1 (N2680, N2673);
nor NOR2 (N2681, N2667, N2219);
nor NOR4 (N2682, N2676, N636, N2003, N2583);
nand NAND4 (N2683, N2677, N1402, N2129, N2669);
not NOT1 (N2684, N2662);
buf BUF1 (N2685, N2649);
nand NAND2 (N2686, N2681, N508);
and AND3 (N2687, N2682, N2278, N368);
buf BUF1 (N2688, N2670);
buf BUF1 (N2689, N2686);
and AND4 (N2690, N2689, N1998, N2477, N2413);
not NOT1 (N2691, N2688);
not NOT1 (N2692, N2680);
not NOT1 (N2693, N2685);
buf BUF1 (N2694, N2693);
or OR2 (N2695, N2675, N935);
and AND2 (N2696, N2679, N2583);
or OR2 (N2697, N2684, N267);
xor XOR2 (N2698, N2690, N515);
nor NOR4 (N2699, N2660, N2460, N2285, N1694);
buf BUF1 (N2700, N2697);
or OR3 (N2701, N2698, N2436, N254);
or OR4 (N2702, N2683, N718, N1388, N1055);
buf BUF1 (N2703, N2691);
or OR2 (N2704, N2687, N1998);
xor XOR2 (N2705, N2700, N2660);
nor NOR3 (N2706, N2705, N1369, N850);
buf BUF1 (N2707, N2702);
or OR3 (N2708, N2699, N2455, N252);
not NOT1 (N2709, N2694);
and AND2 (N2710, N2692, N515);
not NOT1 (N2711, N2710);
xor XOR2 (N2712, N2708, N212);
xor XOR2 (N2713, N2707, N2685);
xor XOR2 (N2714, N2711, N178);
buf BUF1 (N2715, N2703);
nand NAND2 (N2716, N2696, N992);
xor XOR2 (N2717, N2714, N1970);
or OR4 (N2718, N2695, N1510, N2182, N2328);
and AND4 (N2719, N2701, N2417, N2413, N534);
and AND4 (N2720, N2715, N203, N1337, N2401);
or OR3 (N2721, N2716, N1133, N58);
nor NOR4 (N2722, N2704, N2426, N370, N514);
or OR4 (N2723, N2718, N2559, N2181, N2079);
xor XOR2 (N2724, N2721, N1089);
xor XOR2 (N2725, N2706, N1448);
nand NAND2 (N2726, N2724, N843);
and AND2 (N2727, N2722, N2646);
xor XOR2 (N2728, N2717, N770);
nor NOR2 (N2729, N2713, N734);
nor NOR3 (N2730, N2729, N2560, N195);
not NOT1 (N2731, N2726);
nand NAND4 (N2732, N2709, N2004, N2290, N643);
buf BUF1 (N2733, N2728);
xor XOR2 (N2734, N2725, N45);
buf BUF1 (N2735, N2733);
xor XOR2 (N2736, N2720, N2452);
and AND2 (N2737, N2736, N1787);
not NOT1 (N2738, N2737);
or OR4 (N2739, N2712, N182, N1284, N2477);
nand NAND3 (N2740, N2735, N1078, N777);
buf BUF1 (N2741, N2740);
xor XOR2 (N2742, N2727, N1405);
not NOT1 (N2743, N2723);
nand NAND2 (N2744, N2742, N8);
and AND3 (N2745, N2744, N671, N2352);
buf BUF1 (N2746, N2732);
buf BUF1 (N2747, N2743);
or OR2 (N2748, N2739, N86);
or OR3 (N2749, N2738, N615, N2156);
nand NAND2 (N2750, N2747, N740);
not NOT1 (N2751, N2750);
and AND3 (N2752, N2741, N2010, N729);
not NOT1 (N2753, N2719);
or OR3 (N2754, N2751, N798, N1080);
xor XOR2 (N2755, N2734, N1158);
xor XOR2 (N2756, N2745, N1849);
and AND3 (N2757, N2752, N1244, N271);
and AND3 (N2758, N2730, N2260, N1078);
and AND4 (N2759, N2748, N194, N2417, N2443);
nand NAND3 (N2760, N2746, N548, N2174);
and AND3 (N2761, N2758, N845, N351);
nand NAND4 (N2762, N2755, N36, N1590, N2723);
nor NOR4 (N2763, N2731, N2507, N2623, N245);
and AND4 (N2764, N2761, N1392, N1092, N1169);
and AND4 (N2765, N2763, N582, N95, N1684);
buf BUF1 (N2766, N2760);
nor NOR4 (N2767, N2765, N1593, N1673, N2283);
nor NOR3 (N2768, N2759, N713, N2123);
xor XOR2 (N2769, N2764, N904);
nor NOR2 (N2770, N2757, N1606);
buf BUF1 (N2771, N2770);
and AND4 (N2772, N2749, N1976, N2042, N1737);
or OR4 (N2773, N2768, N1253, N2362, N450);
and AND2 (N2774, N2773, N1529);
nor NOR2 (N2775, N2762, N1809);
buf BUF1 (N2776, N2756);
or OR4 (N2777, N2776, N1697, N2273, N2259);
nand NAND3 (N2778, N2769, N1455, N2282);
xor XOR2 (N2779, N2753, N1115);
and AND4 (N2780, N2766, N2395, N1441, N1250);
xor XOR2 (N2781, N2780, N344);
not NOT1 (N2782, N2778);
xor XOR2 (N2783, N2775, N2476);
and AND2 (N2784, N2774, N1045);
nor NOR2 (N2785, N2781, N1836);
nor NOR2 (N2786, N2771, N2193);
nor NOR4 (N2787, N2785, N7, N249, N636);
or OR2 (N2788, N2782, N2678);
nor NOR3 (N2789, N2754, N645, N1596);
xor XOR2 (N2790, N2777, N293);
not NOT1 (N2791, N2788);
or OR2 (N2792, N2779, N638);
nand NAND2 (N2793, N2787, N441);
buf BUF1 (N2794, N2791);
buf BUF1 (N2795, N2772);
buf BUF1 (N2796, N2783);
nor NOR3 (N2797, N2784, N621, N89);
buf BUF1 (N2798, N2795);
nand NAND4 (N2799, N2798, N2245, N1019, N2251);
nor NOR4 (N2800, N2793, N604, N2421, N1120);
buf BUF1 (N2801, N2786);
nor NOR3 (N2802, N2796, N543, N2402);
or OR4 (N2803, N2790, N2084, N1492, N2360);
and AND4 (N2804, N2803, N920, N556, N2711);
nor NOR2 (N2805, N2789, N2540);
nor NOR2 (N2806, N2805, N2238);
nor NOR4 (N2807, N2794, N693, N2725, N1705);
buf BUF1 (N2808, N2797);
not NOT1 (N2809, N2802);
or OR2 (N2810, N2800, N2700);
nor NOR4 (N2811, N2767, N1775, N2306, N1987);
nor NOR2 (N2812, N2808, N1859);
and AND3 (N2813, N2809, N178, N1835);
nand NAND4 (N2814, N2810, N799, N1474, N602);
or OR4 (N2815, N2814, N712, N1744, N221);
nor NOR4 (N2816, N2806, N1313, N1133, N523);
nand NAND2 (N2817, N2801, N2813);
buf BUF1 (N2818, N358);
xor XOR2 (N2819, N2799, N797);
buf BUF1 (N2820, N2815);
not NOT1 (N2821, N2817);
or OR3 (N2822, N2792, N2141, N912);
buf BUF1 (N2823, N2804);
buf BUF1 (N2824, N2816);
buf BUF1 (N2825, N2823);
xor XOR2 (N2826, N2818, N807);
buf BUF1 (N2827, N2821);
xor XOR2 (N2828, N2825, N2724);
nand NAND3 (N2829, N2819, N2157, N1324);
xor XOR2 (N2830, N2822, N1712);
buf BUF1 (N2831, N2812);
not NOT1 (N2832, N2820);
and AND3 (N2833, N2826, N1246, N326);
or OR2 (N2834, N2811, N495);
not NOT1 (N2835, N2827);
or OR3 (N2836, N2832, N604, N1438);
nand NAND4 (N2837, N2829, N1465, N882, N1934);
nand NAND4 (N2838, N2835, N1669, N1325, N1112);
nor NOR2 (N2839, N2837, N227);
buf BUF1 (N2840, N2836);
nand NAND4 (N2841, N2839, N2038, N1261, N454);
or OR3 (N2842, N2828, N321, N1239);
nor NOR2 (N2843, N2840, N1454);
xor XOR2 (N2844, N2833, N2066);
or OR4 (N2845, N2838, N963, N598, N1137);
or OR4 (N2846, N2830, N1738, N241, N864);
not NOT1 (N2847, N2831);
and AND4 (N2848, N2824, N2737, N2065, N2679);
nor NOR2 (N2849, N2841, N1886);
xor XOR2 (N2850, N2848, N391);
buf BUF1 (N2851, N2842);
and AND2 (N2852, N2849, N109);
xor XOR2 (N2853, N2846, N286);
not NOT1 (N2854, N2843);
buf BUF1 (N2855, N2845);
not NOT1 (N2856, N2834);
nand NAND3 (N2857, N2854, N2841, N1619);
and AND4 (N2858, N2807, N715, N1169, N930);
not NOT1 (N2859, N2858);
nand NAND4 (N2860, N2850, N687, N727, N1917);
not NOT1 (N2861, N2857);
xor XOR2 (N2862, N2853, N2247);
not NOT1 (N2863, N2844);
not NOT1 (N2864, N2851);
xor XOR2 (N2865, N2852, N1519);
nand NAND3 (N2866, N2856, N619, N1645);
or OR4 (N2867, N2864, N541, N435, N681);
and AND4 (N2868, N2860, N1176, N2418, N1800);
xor XOR2 (N2869, N2863, N1463);
xor XOR2 (N2870, N2855, N2412);
xor XOR2 (N2871, N2870, N658);
and AND2 (N2872, N2868, N1564);
nand NAND4 (N2873, N2862, N1655, N1537, N1189);
not NOT1 (N2874, N2871);
buf BUF1 (N2875, N2869);
or OR4 (N2876, N2867, N2502, N2406, N1790);
xor XOR2 (N2877, N2873, N2283);
nand NAND4 (N2878, N2877, N1304, N2045, N867);
or OR3 (N2879, N2859, N1365, N1549);
nor NOR4 (N2880, N2847, N2503, N1639, N2383);
buf BUF1 (N2881, N2880);
nand NAND4 (N2882, N2878, N850, N2219, N128);
nand NAND3 (N2883, N2876, N537, N2795);
and AND3 (N2884, N2861, N1300, N1204);
nand NAND4 (N2885, N2882, N1938, N2228, N2231);
and AND4 (N2886, N2885, N394, N2476, N123);
nand NAND2 (N2887, N2886, N567);
not NOT1 (N2888, N2865);
and AND3 (N2889, N2875, N2246, N2805);
nor NOR2 (N2890, N2887, N1062);
buf BUF1 (N2891, N2872);
nand NAND3 (N2892, N2881, N1952, N2377);
buf BUF1 (N2893, N2883);
not NOT1 (N2894, N2874);
nor NOR2 (N2895, N2894, N248);
buf BUF1 (N2896, N2889);
nor NOR3 (N2897, N2866, N2753, N358);
nand NAND4 (N2898, N2884, N1548, N2445, N403);
not NOT1 (N2899, N2879);
and AND2 (N2900, N2897, N829);
not NOT1 (N2901, N2891);
buf BUF1 (N2902, N2898);
not NOT1 (N2903, N2896);
buf BUF1 (N2904, N2902);
xor XOR2 (N2905, N2890, N106);
and AND4 (N2906, N2904, N2490, N135, N1057);
not NOT1 (N2907, N2899);
nand NAND4 (N2908, N2901, N2318, N1040, N2600);
not NOT1 (N2909, N2908);
nor NOR2 (N2910, N2893, N1329);
not NOT1 (N2911, N2910);
and AND4 (N2912, N2909, N1043, N249, N471);
nor NOR3 (N2913, N2912, N1085, N2230);
nor NOR2 (N2914, N2888, N627);
buf BUF1 (N2915, N2911);
or OR3 (N2916, N2892, N381, N1308);
nor NOR2 (N2917, N2914, N1098);
buf BUF1 (N2918, N2913);
not NOT1 (N2919, N2900);
and AND2 (N2920, N2919, N14);
or OR3 (N2921, N2920, N1628, N761);
not NOT1 (N2922, N2921);
not NOT1 (N2923, N2895);
and AND4 (N2924, N2906, N2003, N1419, N1772);
buf BUF1 (N2925, N2915);
and AND3 (N2926, N2907, N361, N520);
or OR3 (N2927, N2905, N2527, N216);
and AND2 (N2928, N2916, N1406);
or OR4 (N2929, N2926, N545, N2763, N1797);
or OR4 (N2930, N2918, N2729, N348, N1874);
xor XOR2 (N2931, N2930, N356);
xor XOR2 (N2932, N2903, N986);
xor XOR2 (N2933, N2927, N1898);
xor XOR2 (N2934, N2917, N1171);
or OR4 (N2935, N2923, N2245, N2727, N20);
not NOT1 (N2936, N2931);
buf BUF1 (N2937, N2934);
nor NOR2 (N2938, N2924, N2092);
xor XOR2 (N2939, N2935, N751);
and AND3 (N2940, N2929, N501, N2801);
or OR4 (N2941, N2938, N298, N1782, N949);
not NOT1 (N2942, N2933);
or OR4 (N2943, N2928, N1490, N666, N2513);
nor NOR2 (N2944, N2939, N1700);
buf BUF1 (N2945, N2932);
xor XOR2 (N2946, N2925, N552);
nand NAND4 (N2947, N2946, N1310, N1231, N884);
and AND4 (N2948, N2936, N1245, N695, N2475);
buf BUF1 (N2949, N2944);
or OR2 (N2950, N2942, N2474);
or OR3 (N2951, N2937, N1255, N1418);
nand NAND3 (N2952, N2945, N389, N2833);
buf BUF1 (N2953, N2941);
buf BUF1 (N2954, N2943);
and AND2 (N2955, N2940, N2933);
or OR2 (N2956, N2952, N45);
and AND2 (N2957, N2954, N2948);
buf BUF1 (N2958, N689);
and AND2 (N2959, N2922, N1736);
buf BUF1 (N2960, N2947);
nand NAND3 (N2961, N2953, N361, N1554);
nand NAND2 (N2962, N2949, N2225);
nand NAND4 (N2963, N2951, N2437, N2568, N162);
not NOT1 (N2964, N2963);
not NOT1 (N2965, N2961);
or OR2 (N2966, N2965, N2438);
and AND4 (N2967, N2957, N1076, N366, N1998);
or OR2 (N2968, N2956, N2198);
nand NAND3 (N2969, N2968, N687, N2492);
and AND4 (N2970, N2950, N567, N2145, N2456);
nand NAND4 (N2971, N2960, N986, N2747, N1508);
or OR3 (N2972, N2967, N1922, N1622);
xor XOR2 (N2973, N2970, N2606);
or OR3 (N2974, N2973, N2420, N162);
nor NOR2 (N2975, N2966, N2005);
not NOT1 (N2976, N2975);
not NOT1 (N2977, N2972);
and AND3 (N2978, N2959, N168, N2779);
not NOT1 (N2979, N2958);
xor XOR2 (N2980, N2964, N1795);
and AND3 (N2981, N2977, N1145, N2604);
xor XOR2 (N2982, N2962, N2500);
nor NOR3 (N2983, N2955, N2754, N508);
nand NAND2 (N2984, N2983, N2503);
not NOT1 (N2985, N2981);
nor NOR2 (N2986, N2984, N2810);
or OR4 (N2987, N2979, N735, N2036, N976);
or OR4 (N2988, N2969, N1812, N2804, N81);
xor XOR2 (N2989, N2982, N2644);
xor XOR2 (N2990, N2988, N2775);
xor XOR2 (N2991, N2971, N297);
and AND3 (N2992, N2974, N2890, N460);
buf BUF1 (N2993, N2980);
and AND4 (N2994, N2993, N2658, N2260, N796);
buf BUF1 (N2995, N2976);
and AND2 (N2996, N2978, N166);
xor XOR2 (N2997, N2996, N1597);
xor XOR2 (N2998, N2986, N2208);
nor NOR3 (N2999, N2992, N156, N2368);
and AND3 (N3000, N2999, N1214, N2749);
xor XOR2 (N3001, N2989, N433);
xor XOR2 (N3002, N3000, N2023);
not NOT1 (N3003, N2998);
xor XOR2 (N3004, N2991, N259);
and AND4 (N3005, N3001, N1830, N1502, N2637);
and AND3 (N3006, N2995, N2214, N316);
buf BUF1 (N3007, N3002);
nor NOR3 (N3008, N2987, N995, N2602);
and AND2 (N3009, N3008, N1053);
not NOT1 (N3010, N2997);
nor NOR4 (N3011, N2994, N1249, N2170, N284);
buf BUF1 (N3012, N3004);
not NOT1 (N3013, N3010);
xor XOR2 (N3014, N3003, N1087);
or OR4 (N3015, N3011, N2138, N878, N994);
buf BUF1 (N3016, N3012);
and AND3 (N3017, N3016, N1991, N2508);
xor XOR2 (N3018, N3006, N380);
nor NOR3 (N3019, N3017, N2151, N184);
or OR4 (N3020, N3005, N1497, N1929, N2075);
not NOT1 (N3021, N2985);
xor XOR2 (N3022, N3013, N1076);
and AND4 (N3023, N3014, N2709, N2337, N424);
or OR2 (N3024, N3022, N581);
or OR2 (N3025, N3007, N900);
nand NAND4 (N3026, N3019, N1433, N2780, N2826);
buf BUF1 (N3027, N3020);
or OR3 (N3028, N3027, N2321, N1355);
nor NOR2 (N3029, N3025, N2422);
nand NAND2 (N3030, N3021, N473);
or OR4 (N3031, N3026, N1378, N983, N238);
not NOT1 (N3032, N3009);
not NOT1 (N3033, N3031);
and AND2 (N3034, N3033, N2667);
xor XOR2 (N3035, N3029, N794);
buf BUF1 (N3036, N3028);
nor NOR4 (N3037, N3018, N2673, N2835, N1061);
not NOT1 (N3038, N3034);
buf BUF1 (N3039, N3024);
nor NOR2 (N3040, N3036, N1744);
xor XOR2 (N3041, N3037, N846);
not NOT1 (N3042, N3041);
xor XOR2 (N3043, N3035, N2203);
buf BUF1 (N3044, N3042);
nor NOR3 (N3045, N3032, N2181, N1163);
nor NOR4 (N3046, N3043, N2749, N607, N2922);
nor NOR4 (N3047, N3045, N430, N1226, N1433);
nor NOR3 (N3048, N3023, N1815, N116);
or OR2 (N3049, N3048, N2273);
xor XOR2 (N3050, N3044, N2770);
nand NAND2 (N3051, N3050, N2760);
or OR4 (N3052, N3040, N1704, N2794, N1327);
buf BUF1 (N3053, N3046);
buf BUF1 (N3054, N3015);
xor XOR2 (N3055, N3030, N122);
nor NOR3 (N3056, N3047, N2326, N1573);
and AND4 (N3057, N3039, N1527, N652, N1130);
and AND2 (N3058, N3054, N3033);
or OR3 (N3059, N2990, N354, N2001);
nor NOR4 (N3060, N3038, N2110, N908, N112);
and AND4 (N3061, N3060, N750, N1969, N2929);
xor XOR2 (N3062, N3058, N2544);
xor XOR2 (N3063, N3051, N2211);
and AND2 (N3064, N3055, N554);
nor NOR2 (N3065, N3062, N1589);
nor NOR4 (N3066, N3063, N687, N293, N299);
xor XOR2 (N3067, N3065, N922);
nor NOR4 (N3068, N3053, N1578, N1819, N1259);
nor NOR2 (N3069, N3061, N466);
xor XOR2 (N3070, N3066, N2500);
or OR4 (N3071, N3068, N2526, N1007, N2826);
nand NAND2 (N3072, N3071, N2134);
or OR2 (N3073, N3059, N2540);
or OR4 (N3074, N3069, N1763, N1253, N609);
nand NAND4 (N3075, N3067, N887, N2630, N1283);
xor XOR2 (N3076, N3070, N1946);
buf BUF1 (N3077, N3072);
and AND3 (N3078, N3056, N2429, N486);
and AND3 (N3079, N3078, N435, N1582);
not NOT1 (N3080, N3076);
and AND4 (N3081, N3064, N1524, N1948, N1673);
xor XOR2 (N3082, N3075, N1839);
not NOT1 (N3083, N3081);
and AND4 (N3084, N3082, N1918, N1846, N781);
or OR2 (N3085, N3080, N1997);
nor NOR4 (N3086, N3052, N403, N1662, N1592);
not NOT1 (N3087, N3057);
buf BUF1 (N3088, N3085);
or OR3 (N3089, N3073, N921, N2942);
xor XOR2 (N3090, N3088, N1645);
or OR3 (N3091, N3083, N2677, N1702);
or OR4 (N3092, N3086, N1212, N842, N1139);
or OR3 (N3093, N3049, N364, N2339);
and AND3 (N3094, N3074, N1080, N2878);
nand NAND3 (N3095, N3090, N1857, N771);
or OR2 (N3096, N3079, N1056);
nand NAND3 (N3097, N3095, N1790, N877);
not NOT1 (N3098, N3093);
and AND2 (N3099, N3092, N2317);
buf BUF1 (N3100, N3099);
not NOT1 (N3101, N3094);
and AND3 (N3102, N3087, N530, N1712);
or OR2 (N3103, N3089, N2768);
and AND4 (N3104, N3103, N261, N3087, N2652);
nor NOR4 (N3105, N3104, N1798, N2215, N1007);
buf BUF1 (N3106, N3100);
nor NOR3 (N3107, N3102, N330, N338);
or OR4 (N3108, N3107, N843, N2001, N87);
nor NOR3 (N3109, N3077, N1823, N481);
or OR2 (N3110, N3105, N164);
and AND2 (N3111, N3101, N2793);
or OR3 (N3112, N3109, N1020, N3047);
not NOT1 (N3113, N3098);
nand NAND2 (N3114, N3113, N2147);
not NOT1 (N3115, N3108);
nor NOR3 (N3116, N3112, N808, N1684);
not NOT1 (N3117, N3096);
and AND2 (N3118, N3114, N2106);
nand NAND3 (N3119, N3091, N789, N2293);
nand NAND4 (N3120, N3118, N795, N244, N1082);
nand NAND4 (N3121, N3110, N2791, N1231, N1070);
not NOT1 (N3122, N3111);
and AND4 (N3123, N3122, N524, N1800, N2196);
and AND3 (N3124, N3106, N2712, N956);
and AND2 (N3125, N3115, N2728);
nor NOR3 (N3126, N3124, N366, N1528);
nand NAND4 (N3127, N3123, N214, N2096, N2123);
buf BUF1 (N3128, N3097);
or OR3 (N3129, N3119, N3028, N3058);
buf BUF1 (N3130, N3116);
nand NAND2 (N3131, N3117, N791);
buf BUF1 (N3132, N3084);
or OR4 (N3133, N3126, N2952, N1329, N3042);
buf BUF1 (N3134, N3131);
nor NOR2 (N3135, N3133, N1950);
nor NOR3 (N3136, N3129, N2317, N724);
buf BUF1 (N3137, N3121);
xor XOR2 (N3138, N3136, N788);
or OR2 (N3139, N3128, N2126);
not NOT1 (N3140, N3134);
not NOT1 (N3141, N3140);
or OR4 (N3142, N3130, N1759, N1206, N1878);
nand NAND3 (N3143, N3125, N2866, N2150);
and AND4 (N3144, N3139, N2990, N2364, N1085);
and AND3 (N3145, N3141, N1875, N309);
xor XOR2 (N3146, N3137, N1564);
nand NAND3 (N3147, N3127, N2286, N2812);
or OR2 (N3148, N3142, N2285);
not NOT1 (N3149, N3120);
not NOT1 (N3150, N3132);
xor XOR2 (N3151, N3145, N1226);
xor XOR2 (N3152, N3150, N1083);
buf BUF1 (N3153, N3147);
buf BUF1 (N3154, N3152);
nor NOR4 (N3155, N3143, N1569, N3031, N411);
nand NAND3 (N3156, N3155, N738, N841);
xor XOR2 (N3157, N3154, N1791);
not NOT1 (N3158, N3151);
or OR4 (N3159, N3148, N286, N2551, N313);
and AND3 (N3160, N3156, N1005, N1855);
buf BUF1 (N3161, N3146);
not NOT1 (N3162, N3159);
and AND4 (N3163, N3158, N1453, N2628, N603);
or OR3 (N3164, N3135, N2815, N1374);
xor XOR2 (N3165, N3149, N1312);
xor XOR2 (N3166, N3162, N2869);
xor XOR2 (N3167, N3138, N1752);
nor NOR4 (N3168, N3164, N1416, N2269, N2919);
not NOT1 (N3169, N3167);
nor NOR4 (N3170, N3144, N1947, N2819, N310);
or OR2 (N3171, N3169, N1741);
buf BUF1 (N3172, N3166);
xor XOR2 (N3173, N3168, N2646);
not NOT1 (N3174, N3153);
buf BUF1 (N3175, N3170);
and AND2 (N3176, N3163, N2298);
or OR2 (N3177, N3173, N2042);
nand NAND3 (N3178, N3177, N882, N923);
xor XOR2 (N3179, N3161, N1909);
buf BUF1 (N3180, N3165);
and AND4 (N3181, N3175, N1566, N33, N1509);
buf BUF1 (N3182, N3174);
and AND3 (N3183, N3171, N2732, N2738);
not NOT1 (N3184, N3179);
and AND2 (N3185, N3182, N1055);
nor NOR4 (N3186, N3184, N2356, N1008, N1319);
buf BUF1 (N3187, N3172);
nand NAND4 (N3188, N3176, N2275, N1414, N763);
and AND3 (N3189, N3188, N3053, N143);
buf BUF1 (N3190, N3157);
not NOT1 (N3191, N3187);
or OR2 (N3192, N3160, N1906);
nand NAND3 (N3193, N3189, N198, N2594);
buf BUF1 (N3194, N3180);
xor XOR2 (N3195, N3181, N2039);
nor NOR2 (N3196, N3195, N2325);
or OR2 (N3197, N3191, N1604);
xor XOR2 (N3198, N3178, N1258);
nor NOR3 (N3199, N3192, N631, N907);
buf BUF1 (N3200, N3186);
xor XOR2 (N3201, N3198, N2277);
and AND4 (N3202, N3193, N913, N2670, N1860);
xor XOR2 (N3203, N3202, N1322);
and AND3 (N3204, N3203, N1789, N339);
not NOT1 (N3205, N3199);
nand NAND4 (N3206, N3194, N280, N801, N648);
buf BUF1 (N3207, N3185);
nand NAND2 (N3208, N3190, N1413);
and AND2 (N3209, N3205, N839);
nor NOR2 (N3210, N3209, N142);
buf BUF1 (N3211, N3206);
nor NOR3 (N3212, N3208, N2681, N2473);
not NOT1 (N3213, N3196);
not NOT1 (N3214, N3210);
xor XOR2 (N3215, N3183, N1131);
and AND2 (N3216, N3213, N2072);
or OR4 (N3217, N3216, N784, N946, N1455);
and AND2 (N3218, N3204, N1672);
xor XOR2 (N3219, N3207, N1362);
and AND2 (N3220, N3212, N1958);
not NOT1 (N3221, N3200);
and AND4 (N3222, N3201, N1752, N588, N828);
or OR2 (N3223, N3219, N2532);
or OR4 (N3224, N3218, N1585, N1274, N2740);
buf BUF1 (N3225, N3211);
not NOT1 (N3226, N3215);
not NOT1 (N3227, N3226);
or OR4 (N3228, N3197, N1321, N1645, N1968);
nor NOR3 (N3229, N3223, N2879, N1924);
or OR2 (N3230, N3227, N2457);
not NOT1 (N3231, N3230);
nor NOR2 (N3232, N3224, N378);
nor NOR3 (N3233, N3222, N1283, N364);
nand NAND2 (N3234, N3225, N2044);
xor XOR2 (N3235, N3220, N2904);
or OR3 (N3236, N3232, N733, N1992);
xor XOR2 (N3237, N3236, N1333);
and AND3 (N3238, N3214, N3041, N3156);
not NOT1 (N3239, N3229);
nand NAND4 (N3240, N3237, N2285, N1766, N735);
xor XOR2 (N3241, N3231, N1960);
and AND4 (N3242, N3217, N2024, N1918, N3213);
not NOT1 (N3243, N3239);
not NOT1 (N3244, N3221);
nor NOR3 (N3245, N3233, N1441, N2924);
nor NOR3 (N3246, N3234, N1529, N201);
buf BUF1 (N3247, N3244);
nand NAND2 (N3248, N3240, N1191);
nand NAND3 (N3249, N3228, N643, N350);
not NOT1 (N3250, N3238);
nand NAND4 (N3251, N3243, N2310, N2420, N2449);
nand NAND4 (N3252, N3242, N1497, N2107, N3232);
not NOT1 (N3253, N3245);
nor NOR2 (N3254, N3241, N40);
buf BUF1 (N3255, N3251);
buf BUF1 (N3256, N3250);
nand NAND3 (N3257, N3255, N2560, N2918);
nand NAND4 (N3258, N3246, N275, N1452, N2447);
or OR3 (N3259, N3254, N1778, N2723);
not NOT1 (N3260, N3256);
not NOT1 (N3261, N3253);
xor XOR2 (N3262, N3235, N956);
or OR3 (N3263, N3260, N1621, N1147);
nor NOR4 (N3264, N3249, N2763, N1079, N978);
and AND3 (N3265, N3257, N1497, N2457);
not NOT1 (N3266, N3259);
not NOT1 (N3267, N3248);
not NOT1 (N3268, N3265);
nand NAND2 (N3269, N3247, N3092);
and AND4 (N3270, N3258, N1747, N1894, N2350);
xor XOR2 (N3271, N3268, N1920);
nor NOR2 (N3272, N3264, N704);
xor XOR2 (N3273, N3271, N272);
nand NAND4 (N3274, N3270, N1475, N1880, N997);
or OR2 (N3275, N3262, N2292);
nand NAND4 (N3276, N3275, N1062, N1613, N572);
not NOT1 (N3277, N3273);
or OR2 (N3278, N3274, N2374);
xor XOR2 (N3279, N3278, N3046);
nor NOR2 (N3280, N3272, N3207);
buf BUF1 (N3281, N3279);
or OR4 (N3282, N3269, N466, N2391, N1216);
nor NOR4 (N3283, N3252, N1806, N795, N2081);
not NOT1 (N3284, N3281);
or OR4 (N3285, N3263, N1980, N58, N1642);
or OR4 (N3286, N3267, N1335, N1805, N2061);
not NOT1 (N3287, N3285);
buf BUF1 (N3288, N3286);
not NOT1 (N3289, N3283);
nand NAND4 (N3290, N3261, N922, N2887, N3199);
xor XOR2 (N3291, N3288, N1601);
buf BUF1 (N3292, N3289);
nor NOR2 (N3293, N3280, N74);
xor XOR2 (N3294, N3276, N2949);
nor NOR3 (N3295, N3290, N1315, N768);
not NOT1 (N3296, N3284);
buf BUF1 (N3297, N3296);
nand NAND3 (N3298, N3287, N1025, N810);
nand NAND2 (N3299, N3297, N3052);
nand NAND3 (N3300, N3277, N2928, N648);
nand NAND2 (N3301, N3294, N2432);
nand NAND4 (N3302, N3301, N2720, N1368, N2569);
nand NAND3 (N3303, N3292, N2459, N947);
buf BUF1 (N3304, N3293);
nor NOR3 (N3305, N3302, N2969, N567);
or OR4 (N3306, N3300, N667, N1518, N1598);
buf BUF1 (N3307, N3266);
buf BUF1 (N3308, N3295);
or OR2 (N3309, N3291, N2769);
nand NAND2 (N3310, N3299, N1439);
nand NAND2 (N3311, N3307, N2214);
or OR2 (N3312, N3308, N1298);
or OR4 (N3313, N3282, N3032, N2705, N1446);
nand NAND3 (N3314, N3312, N387, N2492);
and AND4 (N3315, N3313, N238, N700, N2798);
nand NAND4 (N3316, N3306, N1255, N1497, N1841);
nand NAND3 (N3317, N3305, N1372, N2946);
nand NAND2 (N3318, N3311, N1528);
and AND2 (N3319, N3303, N831);
nor NOR2 (N3320, N3304, N2883);
or OR3 (N3321, N3314, N670, N1825);
buf BUF1 (N3322, N3318);
xor XOR2 (N3323, N3321, N2208);
buf BUF1 (N3324, N3319);
and AND2 (N3325, N3298, N1233);
not NOT1 (N3326, N3322);
and AND2 (N3327, N3326, N2559);
nand NAND3 (N3328, N3320, N2632, N2300);
xor XOR2 (N3329, N3328, N856);
or OR3 (N3330, N3329, N1520, N789);
or OR2 (N3331, N3315, N2716);
xor XOR2 (N3332, N3330, N2354);
nand NAND2 (N3333, N3331, N1234);
nand NAND3 (N3334, N3317, N2227, N2803);
nand NAND3 (N3335, N3324, N2196, N1007);
or OR4 (N3336, N3327, N775, N1537, N1626);
buf BUF1 (N3337, N3333);
xor XOR2 (N3338, N3335, N1788);
not NOT1 (N3339, N3332);
not NOT1 (N3340, N3339);
or OR4 (N3341, N3337, N820, N7, N1668);
nand NAND3 (N3342, N3316, N2306, N602);
buf BUF1 (N3343, N3323);
not NOT1 (N3344, N3338);
not NOT1 (N3345, N3325);
or OR4 (N3346, N3344, N2378, N1693, N1668);
buf BUF1 (N3347, N3336);
nor NOR2 (N3348, N3309, N1065);
nor NOR2 (N3349, N3343, N2254);
nand NAND4 (N3350, N3342, N1812, N202, N1964);
or OR4 (N3351, N3346, N2215, N1511, N2279);
or OR4 (N3352, N3349, N1458, N995, N1717);
or OR2 (N3353, N3310, N671);
not NOT1 (N3354, N3345);
nand NAND2 (N3355, N3352, N566);
buf BUF1 (N3356, N3355);
buf BUF1 (N3357, N3354);
nor NOR3 (N3358, N3357, N1608, N2454);
not NOT1 (N3359, N3347);
buf BUF1 (N3360, N3341);
nor NOR4 (N3361, N3360, N398, N1513, N2853);
or OR3 (N3362, N3359, N2970, N1473);
buf BUF1 (N3363, N3362);
not NOT1 (N3364, N3353);
not NOT1 (N3365, N3364);
nand NAND3 (N3366, N3340, N3293, N622);
and AND3 (N3367, N3366, N2946, N1786);
xor XOR2 (N3368, N3361, N2447);
and AND2 (N3369, N3358, N1902);
nand NAND2 (N3370, N3369, N765);
and AND2 (N3371, N3334, N964);
xor XOR2 (N3372, N3370, N963);
nor NOR2 (N3373, N3365, N1557);
and AND3 (N3374, N3373, N836, N1517);
not NOT1 (N3375, N3372);
nand NAND3 (N3376, N3368, N2685, N2222);
not NOT1 (N3377, N3367);
not NOT1 (N3378, N3363);
or OR3 (N3379, N3350, N311, N798);
nand NAND3 (N3380, N3376, N1726, N2658);
and AND2 (N3381, N3378, N1932);
or OR4 (N3382, N3377, N783, N729, N603);
nand NAND4 (N3383, N3374, N1693, N1862, N1428);
nand NAND3 (N3384, N3383, N697, N3361);
nor NOR4 (N3385, N3384, N3009, N954, N1692);
nor NOR4 (N3386, N3351, N1148, N1185, N3199);
xor XOR2 (N3387, N3382, N1594);
not NOT1 (N3388, N3386);
xor XOR2 (N3389, N3356, N1031);
xor XOR2 (N3390, N3385, N2294);
and AND4 (N3391, N3381, N446, N170, N2800);
or OR3 (N3392, N3380, N934, N3279);
or OR4 (N3393, N3371, N2084, N49, N1905);
xor XOR2 (N3394, N3390, N350);
xor XOR2 (N3395, N3392, N3313);
or OR4 (N3396, N3375, N437, N238, N1993);
nor NOR2 (N3397, N3394, N2697);
buf BUF1 (N3398, N3389);
nand NAND4 (N3399, N3398, N1845, N2152, N835);
not NOT1 (N3400, N3393);
not NOT1 (N3401, N3348);
nand NAND4 (N3402, N3401, N1414, N1596, N1303);
not NOT1 (N3403, N3400);
and AND2 (N3404, N3399, N2304);
not NOT1 (N3405, N3404);
buf BUF1 (N3406, N3379);
xor XOR2 (N3407, N3403, N743);
buf BUF1 (N3408, N3407);
or OR3 (N3409, N3387, N1766, N1832);
or OR4 (N3410, N3391, N601, N1273, N646);
or OR3 (N3411, N3402, N3186, N813);
buf BUF1 (N3412, N3396);
or OR4 (N3413, N3406, N1725, N3407, N2993);
not NOT1 (N3414, N3395);
nor NOR3 (N3415, N3414, N1402, N2681);
or OR4 (N3416, N3408, N1097, N1754, N3150);
and AND3 (N3417, N3415, N1590, N168);
xor XOR2 (N3418, N3411, N869);
xor XOR2 (N3419, N3409, N887);
or OR2 (N3420, N3410, N1058);
and AND4 (N3421, N3418, N1183, N2958, N816);
and AND2 (N3422, N3405, N1757);
nand NAND4 (N3423, N3388, N1603, N1499, N870);
nor NOR2 (N3424, N3413, N1439);
xor XOR2 (N3425, N3412, N1384);
buf BUF1 (N3426, N3419);
buf BUF1 (N3427, N3397);
or OR4 (N3428, N3425, N1561, N1676, N1958);
xor XOR2 (N3429, N3421, N1909);
nand NAND4 (N3430, N3423, N1419, N2217, N509);
and AND2 (N3431, N3427, N453);
nor NOR3 (N3432, N3416, N727, N312);
nand NAND4 (N3433, N3422, N1037, N63, N1665);
not NOT1 (N3434, N3432);
xor XOR2 (N3435, N3417, N1899);
xor XOR2 (N3436, N3426, N733);
buf BUF1 (N3437, N3434);
buf BUF1 (N3438, N3428);
not NOT1 (N3439, N3420);
buf BUF1 (N3440, N3424);
and AND3 (N3441, N3430, N2428, N1166);
not NOT1 (N3442, N3440);
or OR3 (N3443, N3442, N160, N2958);
nor NOR3 (N3444, N3433, N588, N1750);
nand NAND4 (N3445, N3437, N208, N1311, N1310);
nor NOR2 (N3446, N3445, N2594);
nor NOR4 (N3447, N3444, N1037, N2623, N1364);
nand NAND3 (N3448, N3441, N994, N2141);
not NOT1 (N3449, N3439);
nand NAND2 (N3450, N3446, N311);
buf BUF1 (N3451, N3447);
not NOT1 (N3452, N3443);
nor NOR4 (N3453, N3452, N1034, N9, N558);
nor NOR2 (N3454, N3431, N259);
and AND2 (N3455, N3435, N3039);
nor NOR3 (N3456, N3454, N1543, N1367);
or OR2 (N3457, N3429, N2559);
or OR4 (N3458, N3455, N1382, N2058, N3341);
buf BUF1 (N3459, N3448);
or OR2 (N3460, N3450, N386);
xor XOR2 (N3461, N3438, N2192);
not NOT1 (N3462, N3456);
xor XOR2 (N3463, N3453, N3314);
nor NOR2 (N3464, N3463, N1590);
nor NOR2 (N3465, N3457, N1706);
and AND4 (N3466, N3458, N3177, N2014, N1160);
nor NOR2 (N3467, N3460, N3319);
xor XOR2 (N3468, N3466, N2176);
xor XOR2 (N3469, N3461, N2774);
not NOT1 (N3470, N3449);
or OR2 (N3471, N3451, N1366);
and AND4 (N3472, N3436, N2531, N460, N2036);
and AND2 (N3473, N3469, N3081);
not NOT1 (N3474, N3464);
buf BUF1 (N3475, N3473);
xor XOR2 (N3476, N3475, N621);
not NOT1 (N3477, N3471);
and AND3 (N3478, N3468, N3461, N879);
nand NAND4 (N3479, N3476, N606, N575, N417);
xor XOR2 (N3480, N3477, N755);
buf BUF1 (N3481, N3459);
buf BUF1 (N3482, N3465);
nand NAND4 (N3483, N3474, N2709, N2808, N573);
buf BUF1 (N3484, N3478);
xor XOR2 (N3485, N3482, N989);
and AND4 (N3486, N3480, N345, N770, N1209);
or OR3 (N3487, N3486, N2179, N281);
nand NAND4 (N3488, N3484, N2601, N2400, N631);
nor NOR4 (N3489, N3462, N258, N2925, N2126);
not NOT1 (N3490, N3479);
buf BUF1 (N3491, N3472);
nor NOR4 (N3492, N3483, N3151, N3277, N935);
or OR3 (N3493, N3467, N3005, N556);
and AND3 (N3494, N3491, N1799, N1672);
nor NOR3 (N3495, N3492, N944, N3362);
or OR3 (N3496, N3485, N2049, N2194);
nand NAND4 (N3497, N3496, N1269, N23, N3125);
and AND3 (N3498, N3488, N3255, N2113);
xor XOR2 (N3499, N3470, N1408);
buf BUF1 (N3500, N3497);
xor XOR2 (N3501, N3487, N2975);
buf BUF1 (N3502, N3481);
not NOT1 (N3503, N3499);
nor NOR4 (N3504, N3502, N1438, N2618, N3389);
buf BUF1 (N3505, N3501);
nand NAND3 (N3506, N3494, N2697, N3338);
xor XOR2 (N3507, N3500, N2806);
nor NOR4 (N3508, N3493, N895, N2029, N688);
not NOT1 (N3509, N3504);
xor XOR2 (N3510, N3508, N1568);
or OR4 (N3511, N3505, N3094, N1507, N1984);
buf BUF1 (N3512, N3506);
and AND2 (N3513, N3498, N1237);
nand NAND2 (N3514, N3513, N3471);
or OR4 (N3515, N3511, N3160, N2578, N823);
nor NOR3 (N3516, N3495, N3163, N2839);
buf BUF1 (N3517, N3490);
buf BUF1 (N3518, N3489);
nand NAND3 (N3519, N3517, N51, N3129);
and AND2 (N3520, N3503, N94);
or OR3 (N3521, N3507, N1771, N2002);
or OR4 (N3522, N3510, N1781, N245, N3071);
nor NOR2 (N3523, N3516, N2025);
nand NAND3 (N3524, N3519, N420, N1149);
buf BUF1 (N3525, N3512);
buf BUF1 (N3526, N3520);
nor NOR2 (N3527, N3521, N1030);
or OR4 (N3528, N3509, N1482, N2028, N2639);
nand NAND2 (N3529, N3514, N2469);
and AND2 (N3530, N3524, N703);
or OR3 (N3531, N3530, N109, N2929);
buf BUF1 (N3532, N3518);
xor XOR2 (N3533, N3525, N1437);
nor NOR3 (N3534, N3529, N2874, N2668);
or OR3 (N3535, N3532, N3302, N110);
and AND4 (N3536, N3534, N518, N2986, N1676);
and AND4 (N3537, N3526, N2772, N1351, N2954);
nand NAND3 (N3538, N3536, N3322, N2965);
not NOT1 (N3539, N3528);
nor NOR3 (N3540, N3515, N483, N3190);
xor XOR2 (N3541, N3538, N968);
buf BUF1 (N3542, N3539);
and AND2 (N3543, N3522, N1342);
nand NAND3 (N3544, N3523, N2154, N771);
nor NOR3 (N3545, N3533, N921, N3087);
and AND3 (N3546, N3540, N1984, N507);
buf BUF1 (N3547, N3527);
not NOT1 (N3548, N3541);
nor NOR2 (N3549, N3531, N3537);
and AND2 (N3550, N3281, N459);
buf BUF1 (N3551, N3545);
buf BUF1 (N3552, N3549);
xor XOR2 (N3553, N3551, N2593);
xor XOR2 (N3554, N3543, N124);
xor XOR2 (N3555, N3542, N2820);
not NOT1 (N3556, N3548);
nor NOR2 (N3557, N3556, N1614);
and AND4 (N3558, N3547, N1302, N3214, N2540);
nor NOR2 (N3559, N3546, N1774);
nand NAND2 (N3560, N3559, N1182);
or OR2 (N3561, N3557, N2589);
or OR4 (N3562, N3558, N1967, N3474, N2910);
or OR2 (N3563, N3554, N1655);
or OR2 (N3564, N3552, N3273);
not NOT1 (N3565, N3562);
not NOT1 (N3566, N3561);
or OR4 (N3567, N3535, N524, N3543, N672);
not NOT1 (N3568, N3565);
xor XOR2 (N3569, N3563, N3366);
xor XOR2 (N3570, N3568, N3354);
nor NOR4 (N3571, N3553, N2078, N2230, N827);
nor NOR3 (N3572, N3566, N53, N3153);
and AND3 (N3573, N3560, N1006, N730);
or OR4 (N3574, N3544, N433, N2472, N1005);
buf BUF1 (N3575, N3574);
and AND4 (N3576, N3567, N3362, N2933, N2356);
buf BUF1 (N3577, N3573);
and AND3 (N3578, N3577, N1474, N166);
or OR4 (N3579, N3576, N1330, N110, N3292);
not NOT1 (N3580, N3571);
buf BUF1 (N3581, N3580);
nor NOR4 (N3582, N3569, N1354, N2822, N1097);
nor NOR2 (N3583, N3575, N461);
buf BUF1 (N3584, N3581);
xor XOR2 (N3585, N3584, N2420);
or OR2 (N3586, N3550, N1548);
xor XOR2 (N3587, N3570, N2280);
nand NAND3 (N3588, N3585, N3529, N2515);
not NOT1 (N3589, N3587);
nand NAND3 (N3590, N3578, N1522, N3409);
not NOT1 (N3591, N3590);
buf BUF1 (N3592, N3564);
buf BUF1 (N3593, N3555);
buf BUF1 (N3594, N3572);
xor XOR2 (N3595, N3593, N1310);
buf BUF1 (N3596, N3595);
and AND3 (N3597, N3579, N1146, N3512);
not NOT1 (N3598, N3582);
or OR4 (N3599, N3586, N267, N2818, N830);
or OR2 (N3600, N3592, N680);
or OR3 (N3601, N3594, N3239, N2653);
xor XOR2 (N3602, N3597, N3577);
xor XOR2 (N3603, N3588, N3256);
nand NAND4 (N3604, N3602, N1203, N2376, N380);
not NOT1 (N3605, N3583);
not NOT1 (N3606, N3601);
or OR3 (N3607, N3604, N1664, N160);
xor XOR2 (N3608, N3605, N3597);
buf BUF1 (N3609, N3608);
not NOT1 (N3610, N3589);
not NOT1 (N3611, N3610);
not NOT1 (N3612, N3611);
nand NAND3 (N3613, N3612, N1214, N1179);
buf BUF1 (N3614, N3609);
or OR2 (N3615, N3591, N2398);
nor NOR3 (N3616, N3596, N831, N1036);
or OR3 (N3617, N3613, N2282, N2564);
not NOT1 (N3618, N3603);
and AND3 (N3619, N3616, N2473, N2619);
not NOT1 (N3620, N3615);
and AND3 (N3621, N3618, N1667, N1318);
buf BUF1 (N3622, N3607);
not NOT1 (N3623, N3598);
or OR3 (N3624, N3606, N3078, N2957);
or OR4 (N3625, N3600, N2410, N639, N934);
and AND4 (N3626, N3614, N1225, N987, N1452);
not NOT1 (N3627, N3624);
buf BUF1 (N3628, N3599);
nor NOR4 (N3629, N3625, N1288, N1057, N3528);
xor XOR2 (N3630, N3623, N875);
not NOT1 (N3631, N3622);
not NOT1 (N3632, N3619);
xor XOR2 (N3633, N3626, N978);
not NOT1 (N3634, N3627);
not NOT1 (N3635, N3617);
not NOT1 (N3636, N3621);
buf BUF1 (N3637, N3633);
or OR4 (N3638, N3630, N3028, N2773, N155);
not NOT1 (N3639, N3629);
nand NAND2 (N3640, N3628, N2057);
xor XOR2 (N3641, N3638, N2837);
nor NOR4 (N3642, N3637, N1254, N3191, N3326);
or OR3 (N3643, N3640, N3593, N578);
not NOT1 (N3644, N3643);
and AND3 (N3645, N3620, N1297, N784);
and AND4 (N3646, N3631, N806, N1634, N2081);
nor NOR3 (N3647, N3632, N2420, N1263);
nor NOR2 (N3648, N3634, N264);
nor NOR3 (N3649, N3645, N1771, N691);
nand NAND3 (N3650, N3646, N1917, N3207);
and AND3 (N3651, N3635, N2317, N1699);
xor XOR2 (N3652, N3649, N2436);
xor XOR2 (N3653, N3647, N360);
or OR4 (N3654, N3642, N3470, N3106, N228);
not NOT1 (N3655, N3652);
nand NAND3 (N3656, N3639, N2861, N3605);
not NOT1 (N3657, N3653);
xor XOR2 (N3658, N3655, N1080);
nor NOR2 (N3659, N3648, N2378);
nor NOR2 (N3660, N3651, N1700);
not NOT1 (N3661, N3650);
xor XOR2 (N3662, N3659, N1255);
not NOT1 (N3663, N3660);
or OR2 (N3664, N3658, N3046);
not NOT1 (N3665, N3641);
nor NOR2 (N3666, N3636, N2631);
xor XOR2 (N3667, N3657, N3004);
not NOT1 (N3668, N3656);
buf BUF1 (N3669, N3665);
nor NOR2 (N3670, N3663, N1738);
nand NAND3 (N3671, N3661, N2805, N210);
and AND4 (N3672, N3662, N541, N2776, N2192);
not NOT1 (N3673, N3644);
nand NAND2 (N3674, N3666, N3459);
not NOT1 (N3675, N3671);
buf BUF1 (N3676, N3670);
xor XOR2 (N3677, N3654, N3526);
nand NAND4 (N3678, N3669, N1836, N2587, N1318);
not NOT1 (N3679, N3674);
xor XOR2 (N3680, N3677, N875);
not NOT1 (N3681, N3667);
nand NAND4 (N3682, N3680, N1045, N2244, N872);
nor NOR2 (N3683, N3668, N1089);
nand NAND2 (N3684, N3676, N2446);
and AND4 (N3685, N3664, N3303, N3513, N3187);
or OR3 (N3686, N3684, N3482, N1029);
and AND4 (N3687, N3672, N802, N3021, N1121);
and AND2 (N3688, N3686, N2809);
xor XOR2 (N3689, N3675, N2427);
and AND3 (N3690, N3689, N2968, N183);
or OR2 (N3691, N3683, N1274);
nor NOR4 (N3692, N3681, N1068, N1686, N1714);
not NOT1 (N3693, N3678);
not NOT1 (N3694, N3692);
or OR3 (N3695, N3693, N2037, N838);
or OR2 (N3696, N3688, N3002);
and AND2 (N3697, N3694, N2974);
xor XOR2 (N3698, N3690, N851);
buf BUF1 (N3699, N3682);
buf BUF1 (N3700, N3697);
nand NAND2 (N3701, N3700, N538);
nand NAND2 (N3702, N3698, N2149);
and AND3 (N3703, N3696, N2096, N514);
buf BUF1 (N3704, N3687);
xor XOR2 (N3705, N3695, N630);
nand NAND4 (N3706, N3685, N3003, N238, N1342);
and AND3 (N3707, N3702, N310, N3451);
not NOT1 (N3708, N3707);
not NOT1 (N3709, N3706);
nor NOR3 (N3710, N3705, N1402, N66);
nand NAND3 (N3711, N3691, N874, N1568);
nor NOR3 (N3712, N3673, N587, N2007);
and AND4 (N3713, N3709, N2173, N866, N2764);
or OR4 (N3714, N3703, N870, N2078, N2459);
nand NAND2 (N3715, N3701, N2551);
and AND2 (N3716, N3715, N3505);
xor XOR2 (N3717, N3714, N2943);
nand NAND2 (N3718, N3699, N2409);
nor NOR2 (N3719, N3704, N2030);
buf BUF1 (N3720, N3710);
nand NAND2 (N3721, N3718, N171);
or OR3 (N3722, N3708, N2257, N1006);
nand NAND4 (N3723, N3717, N1688, N2873, N2879);
and AND2 (N3724, N3679, N314);
xor XOR2 (N3725, N3712, N2533);
or OR3 (N3726, N3713, N819, N1196);
buf BUF1 (N3727, N3711);
nand NAND4 (N3728, N3721, N3671, N3295, N1760);
buf BUF1 (N3729, N3724);
or OR3 (N3730, N3720, N189, N1564);
and AND2 (N3731, N3723, N282);
nand NAND2 (N3732, N3719, N2890);
not NOT1 (N3733, N3726);
or OR4 (N3734, N3729, N1276, N2404, N609);
not NOT1 (N3735, N3716);
or OR4 (N3736, N3732, N2974, N473, N2903);
buf BUF1 (N3737, N3727);
nor NOR3 (N3738, N3737, N102, N2275);
nand NAND4 (N3739, N3722, N2573, N1809, N1225);
xor XOR2 (N3740, N3734, N351);
nand NAND4 (N3741, N3728, N1879, N3138, N1111);
buf BUF1 (N3742, N3725);
or OR3 (N3743, N3735, N1532, N3293);
or OR4 (N3744, N3741, N396, N436, N2255);
or OR4 (N3745, N3730, N1997, N1958, N2898);
or OR4 (N3746, N3743, N1715, N1450, N2212);
not NOT1 (N3747, N3731);
buf BUF1 (N3748, N3744);
and AND3 (N3749, N3736, N447, N1944);
and AND4 (N3750, N3749, N517, N2177, N3685);
nand NAND4 (N3751, N3742, N3705, N1105, N348);
buf BUF1 (N3752, N3746);
nand NAND4 (N3753, N3733, N2781, N2231, N3692);
xor XOR2 (N3754, N3752, N16);
or OR3 (N3755, N3753, N610, N1690);
not NOT1 (N3756, N3750);
nor NOR2 (N3757, N3740, N1599);
buf BUF1 (N3758, N3739);
not NOT1 (N3759, N3738);
not NOT1 (N3760, N3758);
and AND3 (N3761, N3759, N337, N936);
nor NOR4 (N3762, N3755, N2295, N2197, N667);
nor NOR4 (N3763, N3748, N1259, N253, N1495);
nand NAND4 (N3764, N3757, N2952, N2350, N844);
nor NOR3 (N3765, N3762, N3183, N2380);
buf BUF1 (N3766, N3756);
nand NAND4 (N3767, N3766, N3151, N2226, N520);
not NOT1 (N3768, N3760);
nand NAND3 (N3769, N3745, N41, N3592);
or OR4 (N3770, N3769, N2053, N1177, N2788);
nand NAND3 (N3771, N3747, N3308, N3112);
nor NOR3 (N3772, N3770, N2277, N2778);
and AND2 (N3773, N3763, N1959);
nor NOR4 (N3774, N3767, N3, N1858, N327);
xor XOR2 (N3775, N3774, N1628);
not NOT1 (N3776, N3751);
and AND3 (N3777, N3776, N3355, N1986);
nand NAND3 (N3778, N3777, N3763, N1121);
buf BUF1 (N3779, N3765);
not NOT1 (N3780, N3778);
nor NOR2 (N3781, N3764, N2919);
xor XOR2 (N3782, N3775, N1493);
nor NOR3 (N3783, N3768, N900, N243);
xor XOR2 (N3784, N3780, N448);
nor NOR2 (N3785, N3784, N316);
xor XOR2 (N3786, N3761, N323);
nor NOR3 (N3787, N3754, N2734, N2889);
not NOT1 (N3788, N3787);
nor NOR4 (N3789, N3781, N3032, N1837, N2984);
xor XOR2 (N3790, N3789, N3533);
xor XOR2 (N3791, N3771, N2553);
and AND3 (N3792, N3790, N3209, N1123);
buf BUF1 (N3793, N3779);
xor XOR2 (N3794, N3786, N1545);
not NOT1 (N3795, N3791);
and AND3 (N3796, N3782, N1646, N2048);
and AND4 (N3797, N3796, N573, N59, N3371);
xor XOR2 (N3798, N3785, N2202);
or OR3 (N3799, N3798, N2838, N745);
or OR4 (N3800, N3795, N1009, N3155, N440);
xor XOR2 (N3801, N3800, N1107);
and AND2 (N3802, N3794, N720);
buf BUF1 (N3803, N3799);
nor NOR4 (N3804, N3803, N2869, N2582, N3465);
xor XOR2 (N3805, N3792, N2168);
or OR2 (N3806, N3772, N2094);
nand NAND3 (N3807, N3788, N877, N1253);
xor XOR2 (N3808, N3783, N768);
buf BUF1 (N3809, N3773);
not NOT1 (N3810, N3806);
nor NOR3 (N3811, N3810, N1195, N2196);
not NOT1 (N3812, N3793);
or OR2 (N3813, N3797, N527);
not NOT1 (N3814, N3813);
xor XOR2 (N3815, N3809, N2282);
or OR4 (N3816, N3807, N481, N3560, N1731);
not NOT1 (N3817, N3808);
nand NAND3 (N3818, N3805, N3686, N3127);
not NOT1 (N3819, N3804);
not NOT1 (N3820, N3814);
and AND4 (N3821, N3820, N69, N3447, N1917);
buf BUF1 (N3822, N3818);
nand NAND3 (N3823, N3802, N3694, N3415);
not NOT1 (N3824, N3816);
not NOT1 (N3825, N3821);
nand NAND3 (N3826, N3824, N1199, N3183);
nand NAND3 (N3827, N3811, N507, N2151);
nor NOR2 (N3828, N3815, N2656);
not NOT1 (N3829, N3812);
nor NOR4 (N3830, N3822, N1392, N1414, N1842);
xor XOR2 (N3831, N3825, N2879);
nor NOR3 (N3832, N3828, N508, N1065);
xor XOR2 (N3833, N3823, N1911);
buf BUF1 (N3834, N3832);
buf BUF1 (N3835, N3826);
and AND4 (N3836, N3833, N2705, N2908, N2253);
nor NOR2 (N3837, N3827, N1407);
not NOT1 (N3838, N3836);
buf BUF1 (N3839, N3819);
or OR4 (N3840, N3831, N3725, N759, N3681);
nor NOR2 (N3841, N3835, N2168);
or OR4 (N3842, N3801, N1846, N2910, N3296);
not NOT1 (N3843, N3837);
not NOT1 (N3844, N3843);
nor NOR3 (N3845, N3817, N3502, N2447);
and AND3 (N3846, N3845, N2279, N223);
nand NAND3 (N3847, N3838, N685, N121);
buf BUF1 (N3848, N3834);
buf BUF1 (N3849, N3844);
xor XOR2 (N3850, N3830, N3337);
nor NOR4 (N3851, N3842, N1592, N3022, N2191);
xor XOR2 (N3852, N3846, N1743);
buf BUF1 (N3853, N3849);
or OR2 (N3854, N3839, N2715);
buf BUF1 (N3855, N3840);
or OR3 (N3856, N3852, N2663, N2428);
xor XOR2 (N3857, N3829, N2156);
not NOT1 (N3858, N3857);
nor NOR4 (N3859, N3856, N1649, N2396, N1922);
xor XOR2 (N3860, N3848, N2904);
nand NAND3 (N3861, N3851, N884, N1396);
xor XOR2 (N3862, N3858, N3743);
nor NOR4 (N3863, N3847, N1320, N429, N2857);
nand NAND4 (N3864, N3853, N2593, N1714, N3615);
nor NOR4 (N3865, N3860, N1420, N2473, N3295);
and AND2 (N3866, N3841, N694);
and AND3 (N3867, N3866, N1775, N615);
xor XOR2 (N3868, N3863, N2279);
and AND2 (N3869, N3862, N3132);
xor XOR2 (N3870, N3867, N858);
not NOT1 (N3871, N3868);
nor NOR2 (N3872, N3864, N1791);
not NOT1 (N3873, N3871);
nor NOR4 (N3874, N3870, N3689, N862, N3286);
nor NOR4 (N3875, N3854, N3667, N1243, N182);
and AND4 (N3876, N3872, N1713, N1366, N1857);
or OR3 (N3877, N3869, N1350, N3653);
buf BUF1 (N3878, N3861);
nor NOR3 (N3879, N3876, N1290, N2985);
nor NOR4 (N3880, N3855, N1769, N822, N736);
buf BUF1 (N3881, N3875);
xor XOR2 (N3882, N3879, N1988);
xor XOR2 (N3883, N3880, N1702);
nand NAND4 (N3884, N3877, N2031, N632, N1688);
nor NOR3 (N3885, N3884, N2008, N469);
or OR4 (N3886, N3859, N2289, N2527, N3082);
nand NAND2 (N3887, N3874, N2053);
and AND2 (N3888, N3886, N236);
buf BUF1 (N3889, N3865);
nor NOR3 (N3890, N3883, N2275, N1044);
not NOT1 (N3891, N3882);
and AND3 (N3892, N3887, N2740, N1895);
not NOT1 (N3893, N3889);
or OR4 (N3894, N3873, N1759, N258, N2023);
xor XOR2 (N3895, N3891, N1632);
not NOT1 (N3896, N3893);
nand NAND4 (N3897, N3892, N1690, N2185, N2814);
or OR3 (N3898, N3897, N1508, N2988);
buf BUF1 (N3899, N3895);
nand NAND4 (N3900, N3894, N1205, N2690, N1033);
or OR2 (N3901, N3878, N2563);
buf BUF1 (N3902, N3890);
nand NAND4 (N3903, N3896, N467, N2534, N1892);
not NOT1 (N3904, N3902);
not NOT1 (N3905, N3881);
and AND3 (N3906, N3901, N1231, N3431);
and AND2 (N3907, N3888, N2445);
nand NAND2 (N3908, N3903, N3678);
xor XOR2 (N3909, N3905, N117);
nor NOR3 (N3910, N3908, N1234, N3793);
nand NAND4 (N3911, N3898, N172, N1049, N1597);
or OR3 (N3912, N3899, N3198, N1198);
buf BUF1 (N3913, N3906);
or OR2 (N3914, N3913, N2099);
nand NAND3 (N3915, N3909, N1270, N3553);
xor XOR2 (N3916, N3885, N3136);
and AND3 (N3917, N3916, N3334, N1383);
and AND4 (N3918, N3904, N3381, N3376, N1251);
not NOT1 (N3919, N3910);
xor XOR2 (N3920, N3911, N2126);
not NOT1 (N3921, N3918);
buf BUF1 (N3922, N3907);
nand NAND3 (N3923, N3912, N3508, N1250);
buf BUF1 (N3924, N3923);
nand NAND2 (N3925, N3924, N3545);
nor NOR4 (N3926, N3922, N2880, N2231, N1838);
nand NAND3 (N3927, N3915, N911, N2433);
or OR4 (N3928, N3926, N677, N3615, N903);
nor NOR2 (N3929, N3914, N1525);
not NOT1 (N3930, N3850);
buf BUF1 (N3931, N3900);
or OR4 (N3932, N3930, N3490, N3009, N1868);
xor XOR2 (N3933, N3932, N213);
nor NOR2 (N3934, N3921, N1520);
nor NOR4 (N3935, N3934, N3640, N1916, N3174);
buf BUF1 (N3936, N3920);
buf BUF1 (N3937, N3929);
nand NAND4 (N3938, N3919, N1624, N1663, N282);
or OR3 (N3939, N3935, N1791, N1760);
buf BUF1 (N3940, N3925);
not NOT1 (N3941, N3940);
nor NOR4 (N3942, N3937, N3402, N1804, N3301);
nand NAND4 (N3943, N3938, N2855, N345, N2223);
not NOT1 (N3944, N3939);
and AND4 (N3945, N3943, N631, N868, N2301);
or OR4 (N3946, N3933, N997, N517, N3237);
and AND3 (N3947, N3936, N306, N3934);
xor XOR2 (N3948, N3944, N2136);
nand NAND3 (N3949, N3945, N91, N3037);
nand NAND2 (N3950, N3931, N410);
buf BUF1 (N3951, N3947);
xor XOR2 (N3952, N3946, N267);
or OR3 (N3953, N3928, N3268, N1325);
xor XOR2 (N3954, N3950, N808);
not NOT1 (N3955, N3948);
buf BUF1 (N3956, N3949);
or OR3 (N3957, N3956, N3787, N3667);
and AND2 (N3958, N3955, N3267);
not NOT1 (N3959, N3957);
buf BUF1 (N3960, N3952);
not NOT1 (N3961, N3954);
nor NOR2 (N3962, N3951, N2419);
and AND3 (N3963, N3941, N2511, N279);
nor NOR4 (N3964, N3961, N3748, N1890, N2606);
nor NOR4 (N3965, N3960, N2025, N742, N3441);
nor NOR2 (N3966, N3942, N2542);
xor XOR2 (N3967, N3966, N1887);
nand NAND3 (N3968, N3962, N1403, N3229);
nor NOR3 (N3969, N3953, N466, N382);
nand NAND4 (N3970, N3964, N368, N187, N583);
and AND2 (N3971, N3969, N2525);
or OR4 (N3972, N3959, N3062, N3114, N823);
buf BUF1 (N3973, N3972);
or OR3 (N3974, N3973, N85, N3473);
nor NOR2 (N3975, N3927, N1818);
buf BUF1 (N3976, N3968);
xor XOR2 (N3977, N3971, N3599);
or OR2 (N3978, N3975, N1843);
and AND2 (N3979, N3965, N1510);
nor NOR4 (N3980, N3979, N1838, N2538, N2695);
buf BUF1 (N3981, N3963);
and AND2 (N3982, N3977, N2560);
xor XOR2 (N3983, N3982, N3417);
buf BUF1 (N3984, N3974);
or OR4 (N3985, N3917, N731, N369, N299);
and AND4 (N3986, N3958, N3644, N865, N2387);
not NOT1 (N3987, N3983);
nor NOR4 (N3988, N3976, N2202, N161, N1140);
and AND4 (N3989, N3970, N3838, N2487, N3422);
or OR3 (N3990, N3986, N1450, N780);
buf BUF1 (N3991, N3985);
nand NAND4 (N3992, N3987, N2500, N1245, N2591);
nand NAND3 (N3993, N3981, N399, N2804);
not NOT1 (N3994, N3984);
or OR2 (N3995, N3990, N2541);
nand NAND4 (N3996, N3967, N2745, N3262, N1651);
nand NAND2 (N3997, N3995, N2830);
buf BUF1 (N3998, N3989);
nor NOR2 (N3999, N3993, N1671);
and AND2 (N4000, N3999, N2841);
buf BUF1 (N4001, N3998);
nor NOR3 (N4002, N3988, N3201, N284);
nor NOR3 (N4003, N3978, N2100, N487);
buf BUF1 (N4004, N4002);
or OR4 (N4005, N4004, N3176, N212, N2024);
or OR3 (N4006, N4000, N2975, N2355);
xor XOR2 (N4007, N3994, N3063);
buf BUF1 (N4008, N4007);
or OR2 (N4009, N4006, N222);
xor XOR2 (N4010, N3992, N573);
nand NAND2 (N4011, N4009, N2204);
xor XOR2 (N4012, N4003, N928);
xor XOR2 (N4013, N3997, N2165);
buf BUF1 (N4014, N4013);
or OR2 (N4015, N3980, N2502);
or OR2 (N4016, N3991, N3603);
not NOT1 (N4017, N4001);
or OR4 (N4018, N4005, N572, N189, N1613);
nor NOR4 (N4019, N4011, N2125, N1380, N70);
buf BUF1 (N4020, N4008);
buf BUF1 (N4021, N4010);
nor NOR2 (N4022, N4021, N562);
or OR3 (N4023, N4018, N2844, N2352);
buf BUF1 (N4024, N4012);
or OR3 (N4025, N4020, N1219, N1141);
nand NAND3 (N4026, N4017, N3374, N538);
xor XOR2 (N4027, N4024, N33);
nor NOR3 (N4028, N4026, N1320, N98);
not NOT1 (N4029, N4014);
nand NAND4 (N4030, N4022, N2963, N530, N3177);
and AND4 (N4031, N4025, N2293, N3190, N256);
and AND3 (N4032, N4031, N1298, N2021);
not NOT1 (N4033, N4028);
xor XOR2 (N4034, N4029, N3664);
and AND2 (N4035, N3996, N836);
not NOT1 (N4036, N4015);
and AND3 (N4037, N4032, N800, N1500);
not NOT1 (N4038, N4037);
nand NAND2 (N4039, N4023, N497);
and AND2 (N4040, N4035, N1097);
nor NOR3 (N4041, N4027, N2294, N3859);
or OR3 (N4042, N4019, N2503, N372);
xor XOR2 (N4043, N4042, N2669);
or OR3 (N4044, N4036, N1814, N2492);
and AND4 (N4045, N4039, N1039, N3417, N1524);
and AND3 (N4046, N4041, N1986, N1780);
nor NOR4 (N4047, N4040, N3953, N1482, N1479);
xor XOR2 (N4048, N4046, N584);
and AND3 (N4049, N4033, N2784, N1243);
nor NOR2 (N4050, N4045, N3797);
nand NAND4 (N4051, N4016, N2918, N659, N2543);
or OR3 (N4052, N4049, N1617, N3281);
nor NOR3 (N4053, N4047, N2254, N2194);
buf BUF1 (N4054, N4052);
buf BUF1 (N4055, N4044);
nor NOR2 (N4056, N4050, N954);
buf BUF1 (N4057, N4051);
nand NAND3 (N4058, N4056, N3054, N3957);
nand NAND4 (N4059, N4058, N893, N949, N3030);
nor NOR3 (N4060, N4030, N253, N855);
buf BUF1 (N4061, N4054);
not NOT1 (N4062, N4038);
nand NAND3 (N4063, N4059, N2786, N2164);
xor XOR2 (N4064, N4063, N879);
or OR4 (N4065, N4057, N1965, N2615, N1148);
or OR4 (N4066, N4060, N1140, N2297, N149);
or OR4 (N4067, N4034, N618, N1898, N4020);
and AND3 (N4068, N4062, N3297, N1719);
and AND4 (N4069, N4055, N959, N237, N165);
or OR4 (N4070, N4066, N1740, N4015, N1372);
nor NOR2 (N4071, N4064, N2580);
nor NOR2 (N4072, N4070, N279);
nor NOR2 (N4073, N4069, N105);
nor NOR3 (N4074, N4061, N3061, N3178);
nand NAND4 (N4075, N4072, N3386, N886, N1841);
xor XOR2 (N4076, N4053, N2956);
nor NOR3 (N4077, N4067, N3731, N3098);
or OR3 (N4078, N4073, N1794, N2366);
nand NAND4 (N4079, N4071, N802, N2824, N4015);
nand NAND2 (N4080, N4048, N3771);
xor XOR2 (N4081, N4068, N2217);
buf BUF1 (N4082, N4078);
nand NAND2 (N4083, N4082, N1509);
nand NAND2 (N4084, N4074, N414);
buf BUF1 (N4085, N4079);
buf BUF1 (N4086, N4084);
xor XOR2 (N4087, N4076, N2487);
not NOT1 (N4088, N4085);
and AND3 (N4089, N4081, N1288, N3960);
nor NOR2 (N4090, N4043, N2627);
xor XOR2 (N4091, N4083, N3481);
nor NOR4 (N4092, N4065, N3686, N1574, N3671);
xor XOR2 (N4093, N4088, N2243);
nand NAND3 (N4094, N4089, N2965, N1873);
buf BUF1 (N4095, N4077);
and AND2 (N4096, N4093, N552);
and AND4 (N4097, N4087, N3423, N1702, N2038);
and AND2 (N4098, N4090, N1544);
and AND3 (N4099, N4098, N3225, N1191);
buf BUF1 (N4100, N4095);
not NOT1 (N4101, N4094);
buf BUF1 (N4102, N4100);
nor NOR4 (N4103, N4075, N2728, N1801, N487);
buf BUF1 (N4104, N4086);
nor NOR4 (N4105, N4097, N1735, N2687, N3839);
and AND2 (N4106, N4104, N2179);
not NOT1 (N4107, N4101);
or OR4 (N4108, N4080, N4013, N3828, N2944);
not NOT1 (N4109, N4107);
not NOT1 (N4110, N4105);
xor XOR2 (N4111, N4103, N285);
and AND3 (N4112, N4108, N3265, N422);
not NOT1 (N4113, N4092);
nand NAND4 (N4114, N4096, N932, N3229, N1773);
not NOT1 (N4115, N4091);
and AND3 (N4116, N4109, N2995, N3411);
nor NOR4 (N4117, N4106, N2664, N550, N1158);
not NOT1 (N4118, N4116);
nand NAND4 (N4119, N4110, N1128, N3350, N1412);
or OR2 (N4120, N4114, N1529);
not NOT1 (N4121, N4120);
and AND4 (N4122, N4119, N3396, N1341, N1667);
xor XOR2 (N4123, N4102, N3835);
and AND2 (N4124, N4115, N3793);
xor XOR2 (N4125, N4123, N3775);
nor NOR4 (N4126, N4113, N1113, N1385, N1560);
nor NOR2 (N4127, N4126, N62);
nand NAND2 (N4128, N4122, N678);
and AND2 (N4129, N4121, N547);
nand NAND4 (N4130, N4124, N107, N2177, N3212);
nand NAND2 (N4131, N4111, N3497);
or OR2 (N4132, N4131, N3971);
xor XOR2 (N4133, N4130, N1023);
buf BUF1 (N4134, N4133);
not NOT1 (N4135, N4127);
xor XOR2 (N4136, N4135, N1831);
xor XOR2 (N4137, N4112, N2154);
not NOT1 (N4138, N4099);
nand NAND4 (N4139, N4129, N321, N2543, N711);
buf BUF1 (N4140, N4136);
nand NAND2 (N4141, N4139, N442);
or OR3 (N4142, N4118, N266, N1385);
or OR2 (N4143, N4117, N2016);
xor XOR2 (N4144, N4141, N1769);
buf BUF1 (N4145, N4144);
nor NOR3 (N4146, N4143, N2094, N1963);
nor NOR3 (N4147, N4138, N1403, N504);
buf BUF1 (N4148, N4145);
xor XOR2 (N4149, N4128, N4131);
not NOT1 (N4150, N4149);
buf BUF1 (N4151, N4148);
not NOT1 (N4152, N4147);
xor XOR2 (N4153, N4132, N3195);
xor XOR2 (N4154, N4153, N1195);
buf BUF1 (N4155, N4125);
or OR3 (N4156, N4140, N1225, N3877);
buf BUF1 (N4157, N4155);
buf BUF1 (N4158, N4156);
nor NOR3 (N4159, N4137, N1259, N575);
or OR4 (N4160, N4142, N4155, N1639, N1141);
and AND2 (N4161, N4146, N4136);
nand NAND4 (N4162, N4157, N1701, N2651, N3560);
nand NAND3 (N4163, N4160, N610, N821);
and AND3 (N4164, N4159, N2741, N457);
or OR4 (N4165, N4158, N2286, N365, N2683);
not NOT1 (N4166, N4152);
nor NOR2 (N4167, N4151, N1691);
and AND2 (N4168, N4154, N2186);
or OR3 (N4169, N4165, N2652, N606);
not NOT1 (N4170, N4167);
not NOT1 (N4171, N4161);
xor XOR2 (N4172, N4168, N256);
xor XOR2 (N4173, N4163, N1391);
not NOT1 (N4174, N4169);
xor XOR2 (N4175, N4162, N856);
xor XOR2 (N4176, N4166, N2983);
nor NOR4 (N4177, N4176, N2963, N132, N3106);
buf BUF1 (N4178, N4134);
or OR3 (N4179, N4171, N3608, N758);
nor NOR2 (N4180, N4178, N3256);
buf BUF1 (N4181, N4170);
and AND3 (N4182, N4174, N3174, N2052);
and AND4 (N4183, N4164, N116, N447, N741);
xor XOR2 (N4184, N4181, N208);
or OR4 (N4185, N4183, N3542, N1126, N3162);
and AND2 (N4186, N4179, N1374);
and AND2 (N4187, N4177, N3142);
nand NAND4 (N4188, N4175, N3072, N1229, N358);
nor NOR4 (N4189, N4150, N3257, N191, N2729);
not NOT1 (N4190, N4184);
xor XOR2 (N4191, N4182, N2554);
or OR2 (N4192, N4172, N448);
buf BUF1 (N4193, N4186);
buf BUF1 (N4194, N4193);
or OR4 (N4195, N4173, N4184, N3285, N188);
nor NOR4 (N4196, N4188, N397, N3168, N3606);
not NOT1 (N4197, N4189);
not NOT1 (N4198, N4185);
buf BUF1 (N4199, N4198);
nand NAND3 (N4200, N4196, N2604, N2126);
nand NAND2 (N4201, N4180, N465);
nor NOR2 (N4202, N4187, N2649);
and AND2 (N4203, N4195, N3115);
nand NAND2 (N4204, N4190, N2720);
and AND4 (N4205, N4201, N2554, N866, N1061);
nand NAND4 (N4206, N4204, N922, N1015, N3802);
buf BUF1 (N4207, N4205);
not NOT1 (N4208, N4207);
nor NOR2 (N4209, N4199, N2498);
buf BUF1 (N4210, N4197);
buf BUF1 (N4211, N4203);
xor XOR2 (N4212, N4208, N3197);
xor XOR2 (N4213, N4206, N3340);
xor XOR2 (N4214, N4211, N327);
nand NAND4 (N4215, N4194, N3054, N804, N440);
xor XOR2 (N4216, N4192, N1206);
nand NAND2 (N4217, N4213, N654);
and AND3 (N4218, N4209, N1017, N3443);
and AND3 (N4219, N4200, N2821, N726);
or OR3 (N4220, N4215, N868, N1586);
xor XOR2 (N4221, N4214, N4009);
and AND4 (N4222, N4210, N1800, N2677, N3753);
nor NOR4 (N4223, N4212, N3879, N3772, N2549);
buf BUF1 (N4224, N4222);
not NOT1 (N4225, N4191);
nand NAND4 (N4226, N4225, N238, N3549, N2928);
xor XOR2 (N4227, N4221, N351);
xor XOR2 (N4228, N4226, N228);
and AND2 (N4229, N4202, N3189);
buf BUF1 (N4230, N4217);
buf BUF1 (N4231, N4220);
buf BUF1 (N4232, N4219);
xor XOR2 (N4233, N4216, N3425);
or OR2 (N4234, N4230, N503);
buf BUF1 (N4235, N4223);
xor XOR2 (N4236, N4228, N1629);
nand NAND2 (N4237, N4229, N344);
buf BUF1 (N4238, N4227);
not NOT1 (N4239, N4235);
and AND3 (N4240, N4236, N104, N2478);
or OR4 (N4241, N4232, N1367, N2350, N805);
nor NOR2 (N4242, N4231, N2320);
nor NOR4 (N4243, N4238, N2926, N1372, N2637);
nand NAND3 (N4244, N4233, N3037, N1681);
xor XOR2 (N4245, N4241, N1195);
not NOT1 (N4246, N4218);
buf BUF1 (N4247, N4242);
nand NAND2 (N4248, N4245, N2935);
or OR2 (N4249, N4224, N1246);
not NOT1 (N4250, N4244);
or OR4 (N4251, N4240, N2213, N1068, N2328);
buf BUF1 (N4252, N4248);
nor NOR2 (N4253, N4249, N2150);
buf BUF1 (N4254, N4237);
nor NOR3 (N4255, N4254, N1117, N1376);
not NOT1 (N4256, N4251);
nand NAND2 (N4257, N4256, N3692);
nand NAND3 (N4258, N4247, N750, N3334);
or OR4 (N4259, N4239, N3284, N81, N2873);
xor XOR2 (N4260, N4258, N695);
xor XOR2 (N4261, N4234, N807);
and AND3 (N4262, N4253, N2474, N340);
nor NOR3 (N4263, N4252, N2173, N3422);
nand NAND3 (N4264, N4262, N3508, N436);
nor NOR2 (N4265, N4255, N1032);
or OR4 (N4266, N4260, N1652, N2162, N1931);
nor NOR2 (N4267, N4257, N73);
and AND4 (N4268, N4246, N2659, N1783, N379);
nand NAND3 (N4269, N4268, N4012, N386);
not NOT1 (N4270, N4266);
nand NAND2 (N4271, N4243, N278);
or OR3 (N4272, N4271, N2248, N843);
not NOT1 (N4273, N4250);
not NOT1 (N4274, N4272);
nor NOR4 (N4275, N4274, N1415, N1290, N2191);
nor NOR3 (N4276, N4275, N3988, N2752);
or OR3 (N4277, N4264, N3268, N840);
or OR4 (N4278, N4259, N2194, N1274, N2556);
nor NOR3 (N4279, N4269, N2551, N1103);
not NOT1 (N4280, N4261);
nand NAND2 (N4281, N4270, N2840);
buf BUF1 (N4282, N4276);
not NOT1 (N4283, N4281);
and AND4 (N4284, N4273, N299, N1236, N2359);
nand NAND2 (N4285, N4263, N3925);
and AND4 (N4286, N4267, N36, N3396, N1026);
xor XOR2 (N4287, N4278, N1863);
xor XOR2 (N4288, N4286, N519);
nand NAND2 (N4289, N4277, N512);
buf BUF1 (N4290, N4289);
or OR3 (N4291, N4288, N3163, N2579);
xor XOR2 (N4292, N4279, N909);
and AND3 (N4293, N4290, N447, N1174);
or OR2 (N4294, N4265, N69);
nand NAND2 (N4295, N4292, N952);
or OR4 (N4296, N4294, N4234, N3625, N3245);
not NOT1 (N4297, N4280);
not NOT1 (N4298, N4296);
xor XOR2 (N4299, N4282, N2453);
buf BUF1 (N4300, N4297);
not NOT1 (N4301, N4298);
or OR3 (N4302, N4299, N1190, N1516);
buf BUF1 (N4303, N4291);
buf BUF1 (N4304, N4293);
xor XOR2 (N4305, N4285, N895);
nand NAND2 (N4306, N4303, N217);
and AND4 (N4307, N4301, N3331, N3042, N4044);
buf BUF1 (N4308, N4304);
nand NAND4 (N4309, N4283, N4019, N3516, N1004);
and AND2 (N4310, N4302, N1027);
not NOT1 (N4311, N4308);
buf BUF1 (N4312, N4287);
nor NOR2 (N4313, N4300, N4108);
not NOT1 (N4314, N4307);
nand NAND2 (N4315, N4312, N2088);
nand NAND2 (N4316, N4311, N3040);
not NOT1 (N4317, N4315);
nor NOR3 (N4318, N4310, N3783, N737);
not NOT1 (N4319, N4316);
nand NAND3 (N4320, N4295, N3868, N735);
nand NAND3 (N4321, N4318, N3207, N2574);
not NOT1 (N4322, N4306);
nor NOR2 (N4323, N4317, N2459);
and AND4 (N4324, N4314, N2256, N1694, N2352);
not NOT1 (N4325, N4324);
xor XOR2 (N4326, N4284, N3386);
buf BUF1 (N4327, N4313);
nand NAND4 (N4328, N4320, N398, N3729, N3293);
and AND2 (N4329, N4325, N3537);
and AND4 (N4330, N4329, N2149, N3306, N2371);
buf BUF1 (N4331, N4319);
and AND2 (N4332, N4309, N3871);
buf BUF1 (N4333, N4326);
nand NAND4 (N4334, N4321, N966, N396, N4300);
nand NAND2 (N4335, N4323, N4057);
or OR4 (N4336, N4305, N324, N3617, N3187);
buf BUF1 (N4337, N4336);
and AND4 (N4338, N4330, N886, N2625, N2205);
buf BUF1 (N4339, N4327);
and AND2 (N4340, N4338, N2874);
not NOT1 (N4341, N4335);
or OR4 (N4342, N4341, N1827, N969, N1948);
not NOT1 (N4343, N4322);
xor XOR2 (N4344, N4328, N345);
xor XOR2 (N4345, N4337, N1917);
buf BUF1 (N4346, N4339);
buf BUF1 (N4347, N4332);
or OR4 (N4348, N4344, N3017, N1172, N3288);
nand NAND3 (N4349, N4342, N3812, N4061);
not NOT1 (N4350, N4349);
nor NOR4 (N4351, N4343, N1655, N2447, N1656);
and AND4 (N4352, N4345, N1441, N2926, N309);
not NOT1 (N4353, N4351);
nand NAND3 (N4354, N4333, N1601, N2084);
buf BUF1 (N4355, N4354);
and AND2 (N4356, N4331, N4238);
xor XOR2 (N4357, N4346, N3050);
not NOT1 (N4358, N4340);
not NOT1 (N4359, N4358);
not NOT1 (N4360, N4357);
or OR2 (N4361, N4356, N932);
xor XOR2 (N4362, N4355, N2869);
nand NAND3 (N4363, N4360, N4067, N378);
and AND3 (N4364, N4334, N1576, N2559);
and AND4 (N4365, N4364, N239, N863, N3601);
xor XOR2 (N4366, N4353, N2064);
not NOT1 (N4367, N4362);
buf BUF1 (N4368, N4366);
nor NOR3 (N4369, N4361, N1117, N2508);
buf BUF1 (N4370, N4368);
nand NAND2 (N4371, N4363, N75);
or OR3 (N4372, N4367, N3808, N1096);
nor NOR2 (N4373, N4348, N1006);
not NOT1 (N4374, N4365);
or OR2 (N4375, N4352, N1403);
buf BUF1 (N4376, N4370);
nand NAND3 (N4377, N4347, N4091, N20);
and AND4 (N4378, N4376, N129, N2832, N2003);
nand NAND4 (N4379, N4374, N3244, N3264, N1541);
nor NOR4 (N4380, N4377, N3216, N2746, N2011);
nor NOR2 (N4381, N4359, N3168);
and AND3 (N4382, N4378, N2358, N1780);
or OR3 (N4383, N4372, N4290, N2707);
nor NOR3 (N4384, N4375, N87, N524);
buf BUF1 (N4385, N4371);
or OR2 (N4386, N4383, N28);
and AND2 (N4387, N4386, N2709);
nor NOR2 (N4388, N4369, N3569);
xor XOR2 (N4389, N4381, N761);
or OR3 (N4390, N4350, N1916, N3432);
buf BUF1 (N4391, N4390);
or OR3 (N4392, N4391, N70, N4374);
xor XOR2 (N4393, N4379, N2346);
and AND3 (N4394, N4388, N1141, N4202);
and AND4 (N4395, N4387, N2324, N3635, N2547);
and AND2 (N4396, N4384, N3267);
nor NOR4 (N4397, N4394, N1117, N2938, N865);
buf BUF1 (N4398, N4380);
buf BUF1 (N4399, N4385);
or OR4 (N4400, N4399, N1603, N425, N738);
not NOT1 (N4401, N4382);
not NOT1 (N4402, N4397);
xor XOR2 (N4403, N4389, N2229);
and AND2 (N4404, N4398, N825);
not NOT1 (N4405, N4373);
and AND4 (N4406, N4393, N1459, N3270, N3992);
or OR4 (N4407, N4405, N4284, N3920, N284);
and AND2 (N4408, N4395, N2187);
or OR2 (N4409, N4396, N418);
or OR2 (N4410, N4409, N2694);
not NOT1 (N4411, N4403);
xor XOR2 (N4412, N4408, N2553);
not NOT1 (N4413, N4412);
or OR4 (N4414, N4400, N625, N1895, N4200);
or OR4 (N4415, N4410, N4384, N1592, N2773);
buf BUF1 (N4416, N4402);
or OR3 (N4417, N4406, N3919, N2070);
xor XOR2 (N4418, N4415, N614);
and AND4 (N4419, N4404, N8, N3115, N4210);
nand NAND2 (N4420, N4413, N1672);
not NOT1 (N4421, N4411);
xor XOR2 (N4422, N4401, N1015);
nor NOR2 (N4423, N4420, N3744);
nand NAND3 (N4424, N4419, N3140, N3465);
or OR3 (N4425, N4392, N1904, N350);
not NOT1 (N4426, N4424);
and AND3 (N4427, N4426, N2295, N2953);
nand NAND4 (N4428, N4423, N3119, N1800, N3213);
buf BUF1 (N4429, N4425);
nand NAND4 (N4430, N4428, N3285, N1094, N1802);
or OR3 (N4431, N4422, N4180, N1200);
and AND3 (N4432, N4427, N1565, N1209);
and AND3 (N4433, N4418, N3877, N253);
not NOT1 (N4434, N4407);
and AND4 (N4435, N4429, N3850, N944, N2202);
buf BUF1 (N4436, N4432);
nor NOR4 (N4437, N4433, N4029, N800, N3471);
not NOT1 (N4438, N4431);
xor XOR2 (N4439, N4416, N3757);
buf BUF1 (N4440, N4436);
xor XOR2 (N4441, N4430, N2903);
not NOT1 (N4442, N4440);
nor NOR2 (N4443, N4437, N3295);
and AND2 (N4444, N4438, N3667);
nand NAND4 (N4445, N4421, N300, N4400, N4191);
and AND4 (N4446, N4445, N3878, N2257, N2829);
or OR2 (N4447, N4435, N1871);
and AND4 (N4448, N4443, N1870, N3682, N1689);
nor NOR3 (N4449, N4447, N2287, N2151);
not NOT1 (N4450, N4449);
buf BUF1 (N4451, N4442);
and AND4 (N4452, N4451, N3807, N1759, N115);
xor XOR2 (N4453, N4441, N263);
nor NOR4 (N4454, N4452, N788, N323, N4226);
buf BUF1 (N4455, N4448);
xor XOR2 (N4456, N4414, N2903);
and AND3 (N4457, N4446, N3686, N919);
buf BUF1 (N4458, N4444);
and AND2 (N4459, N4439, N3074);
nand NAND3 (N4460, N4434, N3332, N3652);
nor NOR2 (N4461, N4455, N514);
and AND3 (N4462, N4453, N1593, N1801);
or OR2 (N4463, N4458, N2456);
buf BUF1 (N4464, N4463);
buf BUF1 (N4465, N4460);
and AND3 (N4466, N4457, N2281, N2080);
and AND2 (N4467, N4450, N775);
buf BUF1 (N4468, N4456);
buf BUF1 (N4469, N4461);
not NOT1 (N4470, N4459);
xor XOR2 (N4471, N4462, N3164);
not NOT1 (N4472, N4468);
or OR3 (N4473, N4466, N1564, N3657);
not NOT1 (N4474, N4465);
and AND3 (N4475, N4467, N3408, N3562);
nand NAND4 (N4476, N4417, N4354, N3155, N3200);
or OR4 (N4477, N4475, N3330, N1973, N228);
not NOT1 (N4478, N4471);
xor XOR2 (N4479, N4476, N3124);
not NOT1 (N4480, N4469);
nand NAND3 (N4481, N4478, N56, N1160);
xor XOR2 (N4482, N4477, N3845);
nor NOR4 (N4483, N4479, N4124, N464, N2654);
not NOT1 (N4484, N4480);
nor NOR4 (N4485, N4484, N2913, N4383, N3132);
or OR3 (N4486, N4485, N823, N1000);
nand NAND2 (N4487, N4481, N2850);
nand NAND3 (N4488, N4487, N3694, N3318);
not NOT1 (N4489, N4486);
nor NOR2 (N4490, N4483, N2836);
nand NAND3 (N4491, N4474, N3428, N2170);
nor NOR3 (N4492, N4491, N3444, N3925);
or OR3 (N4493, N4473, N2384, N1563);
buf BUF1 (N4494, N4472);
buf BUF1 (N4495, N4490);
or OR4 (N4496, N4494, N3984, N3735, N1979);
nor NOR2 (N4497, N4495, N1716);
not NOT1 (N4498, N4497);
xor XOR2 (N4499, N4470, N1241);
xor XOR2 (N4500, N4482, N1264);
xor XOR2 (N4501, N4464, N2185);
nor NOR3 (N4502, N4454, N2215, N4150);
and AND3 (N4503, N4502, N2170, N4226);
not NOT1 (N4504, N4498);
or OR3 (N4505, N4496, N583, N1521);
and AND2 (N4506, N4493, N1085);
nand NAND4 (N4507, N4499, N3420, N542, N3773);
not NOT1 (N4508, N4507);
nor NOR4 (N4509, N4488, N418, N2175, N1907);
buf BUF1 (N4510, N4504);
xor XOR2 (N4511, N4501, N3605);
buf BUF1 (N4512, N4510);
buf BUF1 (N4513, N4506);
nor NOR3 (N4514, N4500, N2625, N2212);
or OR2 (N4515, N4492, N642);
and AND2 (N4516, N4503, N308);
nor NOR2 (N4517, N4513, N202);
nand NAND3 (N4518, N4511, N3921, N2497);
nor NOR3 (N4519, N4517, N3457, N3625);
not NOT1 (N4520, N4514);
nand NAND4 (N4521, N4505, N3952, N2916, N1200);
nor NOR4 (N4522, N4521, N443, N588, N352);
nor NOR4 (N4523, N4518, N3370, N1145, N865);
nand NAND4 (N4524, N4522, N3100, N1898, N4290);
nand NAND4 (N4525, N4515, N282, N819, N774);
and AND3 (N4526, N4516, N3170, N445);
and AND4 (N4527, N4489, N3641, N3736, N2418);
nand NAND4 (N4528, N4523, N774, N1714, N195);
nand NAND2 (N4529, N4512, N350);
or OR4 (N4530, N4520, N109, N2266, N3953);
not NOT1 (N4531, N4528);
nor NOR4 (N4532, N4519, N2537, N3256, N3912);
or OR4 (N4533, N4509, N4313, N4297, N4435);
nand NAND2 (N4534, N4532, N772);
not NOT1 (N4535, N4530);
nor NOR3 (N4536, N4535, N3485, N442);
nand NAND3 (N4537, N4525, N2318, N2364);
xor XOR2 (N4538, N4524, N954);
not NOT1 (N4539, N4538);
nand NAND2 (N4540, N4526, N1216);
not NOT1 (N4541, N4527);
or OR3 (N4542, N4531, N3066, N1610);
and AND3 (N4543, N4539, N1965, N719);
and AND4 (N4544, N4536, N4103, N2848, N1540);
buf BUF1 (N4545, N4544);
buf BUF1 (N4546, N4537);
and AND2 (N4547, N4529, N3389);
not NOT1 (N4548, N4541);
or OR2 (N4549, N4533, N1156);
and AND2 (N4550, N4548, N4057);
nand NAND2 (N4551, N4545, N1550);
or OR3 (N4552, N4542, N4323, N1);
nand NAND4 (N4553, N4551, N1659, N126, N1536);
or OR3 (N4554, N4552, N1265, N1749);
not NOT1 (N4555, N4546);
buf BUF1 (N4556, N4547);
buf BUF1 (N4557, N4550);
nor NOR2 (N4558, N4556, N4547);
or OR2 (N4559, N4555, N335);
xor XOR2 (N4560, N4554, N1429);
nor NOR4 (N4561, N4549, N1515, N1083, N2375);
or OR4 (N4562, N4558, N3887, N2343, N3995);
or OR4 (N4563, N4560, N1309, N3863, N1782);
or OR3 (N4564, N4561, N2706, N2264);
not NOT1 (N4565, N4553);
and AND4 (N4566, N4540, N4525, N4300, N4225);
nand NAND2 (N4567, N4543, N3354);
and AND3 (N4568, N4567, N1088, N3067);
nand NAND3 (N4569, N4562, N2548, N2335);
nand NAND3 (N4570, N4566, N311, N1907);
and AND4 (N4571, N4564, N4162, N2665, N1826);
nor NOR4 (N4572, N4534, N125, N2325, N498);
not NOT1 (N4573, N4568);
not NOT1 (N4574, N4573);
xor XOR2 (N4575, N4569, N3747);
nand NAND3 (N4576, N4575, N3031, N3565);
or OR2 (N4577, N4576, N3219);
xor XOR2 (N4578, N4570, N446);
xor XOR2 (N4579, N4572, N4049);
or OR2 (N4580, N4563, N3059);
nand NAND3 (N4581, N4557, N2208, N2156);
nor NOR2 (N4582, N4580, N340);
nand NAND4 (N4583, N4578, N230, N3061, N304);
buf BUF1 (N4584, N4582);
xor XOR2 (N4585, N4577, N2848);
and AND4 (N4586, N4571, N3156, N1258, N3551);
nand NAND4 (N4587, N4574, N1281, N1962, N2237);
and AND3 (N4588, N4584, N4452, N2253);
not NOT1 (N4589, N4559);
xor XOR2 (N4590, N4579, N3784);
or OR2 (N4591, N4585, N338);
xor XOR2 (N4592, N4591, N225);
or OR3 (N4593, N4565, N1997, N2115);
nand NAND4 (N4594, N4586, N3994, N3563, N3547);
or OR2 (N4595, N4592, N2758);
not NOT1 (N4596, N4508);
xor XOR2 (N4597, N4583, N1601);
nand NAND3 (N4598, N4593, N4076, N2695);
buf BUF1 (N4599, N4590);
or OR4 (N4600, N4589, N1694, N4142, N1405);
nand NAND4 (N4601, N4588, N2410, N2244, N206);
not NOT1 (N4602, N4596);
and AND4 (N4603, N4587, N348, N2923, N580);
nor NOR3 (N4604, N4594, N2406, N737);
and AND2 (N4605, N4602, N3228);
or OR4 (N4606, N4599, N584, N1544, N3280);
buf BUF1 (N4607, N4595);
xor XOR2 (N4608, N4606, N3853);
nor NOR4 (N4609, N4603, N2215, N1924, N2728);
and AND3 (N4610, N4607, N1139, N4379);
and AND3 (N4611, N4598, N2132, N826);
buf BUF1 (N4612, N4609);
nor NOR2 (N4613, N4612, N3454);
nand NAND2 (N4614, N4608, N527);
or OR3 (N4615, N4597, N2102, N3870);
nor NOR4 (N4616, N4615, N4436, N1223, N243);
or OR2 (N4617, N4613, N3866);
not NOT1 (N4618, N4604);
buf BUF1 (N4619, N4581);
buf BUF1 (N4620, N4611);
nor NOR4 (N4621, N4614, N2921, N3971, N2313);
not NOT1 (N4622, N4619);
and AND3 (N4623, N4621, N1366, N229);
buf BUF1 (N4624, N4620);
buf BUF1 (N4625, N4610);
nor NOR3 (N4626, N4625, N454, N3119);
nor NOR4 (N4627, N4626, N1100, N860, N4574);
not NOT1 (N4628, N4617);
nor NOR2 (N4629, N4616, N4588);
and AND3 (N4630, N4622, N2208, N3583);
and AND4 (N4631, N4601, N4301, N1481, N2986);
buf BUF1 (N4632, N4630);
and AND4 (N4633, N4605, N4023, N1153, N2592);
nor NOR4 (N4634, N4624, N3760, N3309, N1200);
and AND4 (N4635, N4623, N2337, N3390, N2377);
buf BUF1 (N4636, N4627);
xor XOR2 (N4637, N4636, N4389);
and AND2 (N4638, N4629, N2527);
not NOT1 (N4639, N4600);
nand NAND2 (N4640, N4631, N4558);
not NOT1 (N4641, N4634);
not NOT1 (N4642, N4633);
nor NOR3 (N4643, N4628, N1985, N4570);
not NOT1 (N4644, N4641);
nand NAND4 (N4645, N4640, N2344, N1379, N4307);
and AND4 (N4646, N4642, N3363, N4386, N2109);
not NOT1 (N4647, N4646);
xor XOR2 (N4648, N4644, N1427);
not NOT1 (N4649, N4647);
nand NAND2 (N4650, N4635, N2754);
buf BUF1 (N4651, N4632);
buf BUF1 (N4652, N4618);
and AND4 (N4653, N4650, N2235, N2755, N1200);
nor NOR4 (N4654, N4639, N266, N4368, N1063);
buf BUF1 (N4655, N4651);
or OR4 (N4656, N4655, N2686, N3898, N1607);
nor NOR4 (N4657, N4645, N652, N4115, N962);
and AND3 (N4658, N4657, N4083, N920);
nor NOR2 (N4659, N4638, N4374);
buf BUF1 (N4660, N4654);
nor NOR3 (N4661, N4652, N993, N813);
or OR3 (N4662, N4660, N2480, N3586);
buf BUF1 (N4663, N4659);
and AND4 (N4664, N4653, N699, N3684, N2101);
not NOT1 (N4665, N4661);
and AND2 (N4666, N4656, N1421);
buf BUF1 (N4667, N4665);
xor XOR2 (N4668, N4666, N1831);
nand NAND3 (N4669, N4637, N473, N2959);
nand NAND3 (N4670, N4648, N916, N3418);
nand NAND2 (N4671, N4663, N1188);
xor XOR2 (N4672, N4668, N813);
nor NOR4 (N4673, N4664, N1359, N3431, N4638);
buf BUF1 (N4674, N4649);
buf BUF1 (N4675, N4643);
and AND3 (N4676, N4673, N4221, N581);
and AND4 (N4677, N4674, N3824, N2355, N973);
xor XOR2 (N4678, N4672, N1249);
not NOT1 (N4679, N4678);
not NOT1 (N4680, N4671);
buf BUF1 (N4681, N4675);
nor NOR2 (N4682, N4681, N2268);
nand NAND4 (N4683, N4669, N470, N2437, N2348);
nor NOR2 (N4684, N4676, N3449);
or OR4 (N4685, N4679, N1249, N3197, N4554);
nor NOR4 (N4686, N4658, N2628, N4651, N2115);
xor XOR2 (N4687, N4685, N94);
nand NAND2 (N4688, N4682, N1608);
xor XOR2 (N4689, N4670, N73);
xor XOR2 (N4690, N4662, N3181);
nand NAND4 (N4691, N4689, N4058, N3619, N2091);
and AND4 (N4692, N4667, N3463, N2557, N4120);
and AND3 (N4693, N4677, N2973, N209);
xor XOR2 (N4694, N4690, N888);
not NOT1 (N4695, N4686);
nor NOR3 (N4696, N4694, N3416, N1840);
xor XOR2 (N4697, N4687, N1715);
xor XOR2 (N4698, N4695, N948);
nand NAND2 (N4699, N4696, N1807);
nand NAND4 (N4700, N4688, N3502, N2469, N1200);
not NOT1 (N4701, N4684);
and AND2 (N4702, N4697, N3651);
xor XOR2 (N4703, N4692, N4436);
not NOT1 (N4704, N4698);
not NOT1 (N4705, N4683);
not NOT1 (N4706, N4700);
xor XOR2 (N4707, N4701, N3439);
or OR4 (N4708, N4702, N3657, N1561, N1993);
not NOT1 (N4709, N4706);
not NOT1 (N4710, N4708);
and AND4 (N4711, N4705, N2662, N2098, N2671);
nand NAND3 (N4712, N4704, N4153, N2412);
nand NAND2 (N4713, N4710, N4576);
xor XOR2 (N4714, N4713, N2148);
and AND3 (N4715, N4703, N3569, N3237);
xor XOR2 (N4716, N4712, N2297);
not NOT1 (N4717, N4714);
nand NAND2 (N4718, N4699, N353);
xor XOR2 (N4719, N4716, N834);
xor XOR2 (N4720, N4691, N4095);
nand NAND3 (N4721, N4720, N2703, N2367);
nand NAND3 (N4722, N4707, N232, N596);
xor XOR2 (N4723, N4722, N530);
and AND4 (N4724, N4718, N3167, N223, N3588);
nor NOR2 (N4725, N4721, N901);
nor NOR4 (N4726, N4680, N3744, N345, N1347);
not NOT1 (N4727, N4717);
nor NOR4 (N4728, N4711, N2323, N1692, N2058);
nor NOR4 (N4729, N4728, N3808, N2677, N4123);
and AND3 (N4730, N4729, N742, N1243);
nor NOR4 (N4731, N4723, N3309, N452, N2506);
nor NOR2 (N4732, N4730, N2348);
not NOT1 (N4733, N4693);
or OR2 (N4734, N4727, N61);
nand NAND4 (N4735, N4731, N992, N453, N3327);
and AND2 (N4736, N4735, N1664);
or OR2 (N4737, N4733, N4404);
or OR2 (N4738, N4725, N3780);
buf BUF1 (N4739, N4738);
buf BUF1 (N4740, N4726);
nand NAND4 (N4741, N4737, N4296, N1416, N2112);
xor XOR2 (N4742, N4709, N4433);
or OR2 (N4743, N4724, N517);
nand NAND4 (N4744, N4715, N2281, N1810, N2529);
not NOT1 (N4745, N4739);
or OR3 (N4746, N4719, N3920, N4428);
not NOT1 (N4747, N4746);
xor XOR2 (N4748, N4743, N675);
not NOT1 (N4749, N4745);
buf BUF1 (N4750, N4748);
or OR4 (N4751, N4750, N121, N1058, N4265);
or OR2 (N4752, N4736, N640);
buf BUF1 (N4753, N4747);
nor NOR2 (N4754, N4744, N840);
nor NOR4 (N4755, N4734, N3450, N96, N3544);
nand NAND4 (N4756, N4740, N2024, N68, N1251);
not NOT1 (N4757, N4751);
and AND2 (N4758, N4749, N1016);
xor XOR2 (N4759, N4732, N3959);
buf BUF1 (N4760, N4759);
or OR3 (N4761, N4754, N117, N4464);
buf BUF1 (N4762, N4756);
and AND3 (N4763, N4742, N3256, N2986);
and AND4 (N4764, N4758, N972, N4348, N2624);
and AND3 (N4765, N4757, N3035, N1602);
nand NAND2 (N4766, N4764, N4272);
buf BUF1 (N4767, N4761);
nor NOR2 (N4768, N4753, N1030);
nor NOR3 (N4769, N4755, N4061, N3112);
nor NOR3 (N4770, N4752, N1363, N4575);
xor XOR2 (N4771, N4766, N878);
nand NAND3 (N4772, N4741, N1744, N3174);
xor XOR2 (N4773, N4760, N3835);
and AND4 (N4774, N4767, N1620, N2072, N641);
buf BUF1 (N4775, N4762);
and AND2 (N4776, N4773, N1389);
nor NOR2 (N4777, N4763, N2483);
xor XOR2 (N4778, N4776, N1211);
or OR2 (N4779, N4771, N2908);
nor NOR3 (N4780, N4774, N2153, N2244);
nand NAND2 (N4781, N4778, N159);
not NOT1 (N4782, N4770);
xor XOR2 (N4783, N4775, N2236);
not NOT1 (N4784, N4765);
buf BUF1 (N4785, N4783);
and AND4 (N4786, N4768, N1037, N1838, N4557);
and AND4 (N4787, N4780, N1408, N2028, N1767);
nand NAND3 (N4788, N4769, N831, N122);
nor NOR2 (N4789, N4784, N3760);
nor NOR4 (N4790, N4782, N2723, N609, N1851);
not NOT1 (N4791, N4779);
or OR2 (N4792, N4777, N1483);
and AND4 (N4793, N4781, N3601, N4094, N1719);
buf BUF1 (N4794, N4772);
xor XOR2 (N4795, N4788, N1128);
not NOT1 (N4796, N4791);
and AND4 (N4797, N4792, N2220, N2086, N2685);
or OR2 (N4798, N4786, N1512);
nor NOR3 (N4799, N4795, N2688, N731);
nand NAND3 (N4800, N4790, N2696, N916);
or OR2 (N4801, N4785, N1909);
not NOT1 (N4802, N4801);
or OR2 (N4803, N4793, N1629);
or OR2 (N4804, N4787, N3800);
or OR2 (N4805, N4797, N842);
xor XOR2 (N4806, N4794, N44);
nor NOR4 (N4807, N4806, N4131, N1140, N2336);
xor XOR2 (N4808, N4807, N1856);
or OR2 (N4809, N4789, N1440);
or OR2 (N4810, N4805, N3680);
buf BUF1 (N4811, N4796);
not NOT1 (N4812, N4808);
xor XOR2 (N4813, N4803, N3841);
xor XOR2 (N4814, N4812, N2720);
not NOT1 (N4815, N4814);
xor XOR2 (N4816, N4802, N4251);
and AND2 (N4817, N4800, N1578);
and AND2 (N4818, N4815, N4607);
xor XOR2 (N4819, N4799, N2850);
xor XOR2 (N4820, N4813, N4341);
not NOT1 (N4821, N4798);
nor NOR4 (N4822, N4811, N4014, N3212, N1143);
or OR4 (N4823, N4809, N1714, N2826, N1079);
nor NOR2 (N4824, N4818, N1375);
or OR4 (N4825, N4817, N3488, N1774, N3586);
xor XOR2 (N4826, N4819, N2184);
buf BUF1 (N4827, N4816);
or OR2 (N4828, N4827, N4247);
nor NOR4 (N4829, N4810, N4706, N2240, N1624);
or OR4 (N4830, N4822, N4624, N3662, N1342);
not NOT1 (N4831, N4825);
and AND3 (N4832, N4823, N509, N4211);
nand NAND2 (N4833, N4824, N348);
xor XOR2 (N4834, N4829, N2670);
buf BUF1 (N4835, N4831);
not NOT1 (N4836, N4804);
buf BUF1 (N4837, N4820);
nor NOR4 (N4838, N4830, N3825, N87, N1923);
xor XOR2 (N4839, N4821, N2864);
xor XOR2 (N4840, N4833, N2686);
nor NOR2 (N4841, N4834, N13);
buf BUF1 (N4842, N4840);
buf BUF1 (N4843, N4832);
buf BUF1 (N4844, N4837);
and AND4 (N4845, N4843, N1627, N3523, N3393);
not NOT1 (N4846, N4841);
not NOT1 (N4847, N4846);
not NOT1 (N4848, N4844);
not NOT1 (N4849, N4838);
and AND3 (N4850, N4828, N4429, N1413);
xor XOR2 (N4851, N4847, N2340);
buf BUF1 (N4852, N4826);
buf BUF1 (N4853, N4839);
nor NOR2 (N4854, N4848, N2941);
nand NAND2 (N4855, N4853, N1574);
or OR3 (N4856, N4836, N3302, N684);
or OR3 (N4857, N4850, N4147, N631);
buf BUF1 (N4858, N4845);
nor NOR3 (N4859, N4842, N3086, N3708);
nand NAND4 (N4860, N4849, N1522, N229, N3525);
nor NOR3 (N4861, N4855, N3176, N4542);
not NOT1 (N4862, N4851);
nand NAND2 (N4863, N4862, N1061);
xor XOR2 (N4864, N4863, N4532);
not NOT1 (N4865, N4859);
buf BUF1 (N4866, N4852);
xor XOR2 (N4867, N4860, N3858);
not NOT1 (N4868, N4854);
nand NAND3 (N4869, N4835, N2623, N2954);
nor NOR2 (N4870, N4861, N333);
xor XOR2 (N4871, N4865, N3376);
nand NAND4 (N4872, N4866, N2676, N1511, N3723);
or OR2 (N4873, N4871, N2942);
buf BUF1 (N4874, N4870);
nor NOR4 (N4875, N4872, N1884, N4731, N3991);
nand NAND2 (N4876, N4867, N4608);
and AND3 (N4877, N4858, N3487, N2247);
nor NOR4 (N4878, N4875, N156, N2514, N2859);
buf BUF1 (N4879, N4878);
and AND2 (N4880, N4868, N229);
buf BUF1 (N4881, N4876);
or OR4 (N4882, N4880, N1875, N597, N2224);
not NOT1 (N4883, N4882);
nand NAND4 (N4884, N4877, N2696, N1285, N1501);
nand NAND2 (N4885, N4857, N3666);
buf BUF1 (N4886, N4884);
nor NOR2 (N4887, N4886, N1222);
xor XOR2 (N4888, N4869, N410);
and AND4 (N4889, N4874, N4838, N1363, N2931);
nand NAND2 (N4890, N4888, N871);
and AND2 (N4891, N4856, N442);
or OR4 (N4892, N4873, N1902, N180, N519);
not NOT1 (N4893, N4883);
nor NOR3 (N4894, N4889, N742, N1218);
nor NOR3 (N4895, N4891, N4024, N3888);
buf BUF1 (N4896, N4895);
and AND2 (N4897, N4885, N1540);
or OR4 (N4898, N4881, N4613, N3446, N2452);
nor NOR4 (N4899, N4864, N1667, N3567, N1068);
not NOT1 (N4900, N4879);
xor XOR2 (N4901, N4890, N595);
nor NOR4 (N4902, N4887, N3809, N2171, N3836);
buf BUF1 (N4903, N4893);
and AND2 (N4904, N4897, N3910);
or OR2 (N4905, N4899, N3688);
buf BUF1 (N4906, N4905);
xor XOR2 (N4907, N4894, N1358);
not NOT1 (N4908, N4892);
and AND3 (N4909, N4898, N2564, N364);
buf BUF1 (N4910, N4909);
or OR2 (N4911, N4910, N1546);
nand NAND2 (N4912, N4906, N3311);
nand NAND3 (N4913, N4912, N1031, N866);
or OR4 (N4914, N4896, N4388, N3102, N1454);
nand NAND4 (N4915, N4901, N1141, N4239, N1844);
nand NAND3 (N4916, N4908, N1044, N4083);
not NOT1 (N4917, N4916);
nand NAND2 (N4918, N4914, N3757);
nor NOR3 (N4919, N4918, N1371, N3627);
nor NOR3 (N4920, N4919, N980, N178);
or OR4 (N4921, N4907, N3266, N1058, N1194);
nor NOR2 (N4922, N4913, N1926);
not NOT1 (N4923, N4920);
and AND4 (N4924, N4917, N4137, N4538, N3385);
buf BUF1 (N4925, N4911);
nand NAND2 (N4926, N4902, N2727);
xor XOR2 (N4927, N4900, N974);
or OR2 (N4928, N4903, N1270);
or OR2 (N4929, N4924, N4521);
buf BUF1 (N4930, N4926);
nor NOR3 (N4931, N4929, N949, N2126);
buf BUF1 (N4932, N4925);
nand NAND4 (N4933, N4921, N329, N1253, N241);
xor XOR2 (N4934, N4931, N1390);
not NOT1 (N4935, N4904);
and AND3 (N4936, N4930, N3619, N933);
not NOT1 (N4937, N4922);
nand NAND3 (N4938, N4928, N4620, N1754);
or OR2 (N4939, N4936, N3226);
or OR4 (N4940, N4923, N938, N3312, N2147);
and AND2 (N4941, N4915, N3230);
not NOT1 (N4942, N4940);
and AND3 (N4943, N4933, N4906, N4377);
and AND2 (N4944, N4943, N4496);
buf BUF1 (N4945, N4944);
buf BUF1 (N4946, N4932);
buf BUF1 (N4947, N4937);
nor NOR4 (N4948, N4938, N2832, N3087, N2848);
not NOT1 (N4949, N4945);
nand NAND3 (N4950, N4941, N1647, N3258);
not NOT1 (N4951, N4942);
nor NOR3 (N4952, N4946, N2045, N2053);
buf BUF1 (N4953, N4952);
buf BUF1 (N4954, N4927);
xor XOR2 (N4955, N4949, N1764);
and AND4 (N4956, N4947, N2241, N1929, N2969);
and AND2 (N4957, N4953, N4252);
xor XOR2 (N4958, N4939, N1827);
and AND3 (N4959, N4955, N3985, N1136);
xor XOR2 (N4960, N4956, N2812);
buf BUF1 (N4961, N4959);
xor XOR2 (N4962, N4948, N735);
nand NAND4 (N4963, N4958, N58, N1102, N897);
and AND2 (N4964, N4962, N1480);
buf BUF1 (N4965, N4934);
or OR4 (N4966, N4954, N1665, N1071, N255);
not NOT1 (N4967, N4950);
buf BUF1 (N4968, N4957);
nand NAND2 (N4969, N4965, N2192);
buf BUF1 (N4970, N4935);
not NOT1 (N4971, N4970);
nand NAND2 (N4972, N4968, N4151);
not NOT1 (N4973, N4964);
buf BUF1 (N4974, N4961);
not NOT1 (N4975, N4951);
nand NAND3 (N4976, N4974, N4051, N2158);
nand NAND2 (N4977, N4973, N1048);
nand NAND4 (N4978, N4972, N4504, N2033, N4219);
buf BUF1 (N4979, N4967);
xor XOR2 (N4980, N4979, N3536);
xor XOR2 (N4981, N4969, N3795);
not NOT1 (N4982, N4975);
nor NOR4 (N4983, N4980, N3692, N2395, N4665);
not NOT1 (N4984, N4981);
xor XOR2 (N4985, N4982, N1540);
buf BUF1 (N4986, N4960);
buf BUF1 (N4987, N4978);
xor XOR2 (N4988, N4966, N4211);
not NOT1 (N4989, N4976);
nor NOR2 (N4990, N4987, N706);
buf BUF1 (N4991, N4985);
not NOT1 (N4992, N4984);
or OR3 (N4993, N4971, N3354, N2372);
nor NOR3 (N4994, N4990, N3993, N1188);
or OR4 (N4995, N4992, N3169, N4059, N147);
nor NOR3 (N4996, N4989, N2174, N4476);
or OR3 (N4997, N4963, N1376, N4554);
nor NOR3 (N4998, N4986, N2965, N2340);
and AND2 (N4999, N4988, N3912);
nor NOR3 (N5000, N4998, N2722, N4437);
and AND3 (N5001, N4993, N4460, N4889);
xor XOR2 (N5002, N4999, N2832);
and AND4 (N5003, N4995, N2715, N1218, N4617);
buf BUF1 (N5004, N4996);
nor NOR4 (N5005, N4991, N858, N4372, N4411);
nor NOR3 (N5006, N5005, N884, N3924);
and AND2 (N5007, N5006, N2410);
nor NOR4 (N5008, N5004, N2957, N2045, N4306);
xor XOR2 (N5009, N5008, N3178);
buf BUF1 (N5010, N4997);
not NOT1 (N5011, N5003);
not NOT1 (N5012, N4977);
xor XOR2 (N5013, N5010, N1761);
and AND2 (N5014, N4994, N255);
and AND4 (N5015, N5012, N4233, N1737, N938);
or OR3 (N5016, N4983, N2418, N4803);
nor NOR4 (N5017, N5011, N4448, N165, N282);
not NOT1 (N5018, N5017);
not NOT1 (N5019, N5016);
buf BUF1 (N5020, N5015);
xor XOR2 (N5021, N5009, N3190);
nand NAND2 (N5022, N5019, N3912);
not NOT1 (N5023, N5002);
not NOT1 (N5024, N5013);
and AND2 (N5025, N5021, N2284);
not NOT1 (N5026, N5001);
nor NOR4 (N5027, N5018, N3514, N1523, N3731);
and AND2 (N5028, N5025, N3278);
nor NOR3 (N5029, N5020, N3783, N3366);
buf BUF1 (N5030, N5027);
not NOT1 (N5031, N5022);
nand NAND4 (N5032, N5026, N2222, N1653, N2440);
not NOT1 (N5033, N5030);
nand NAND3 (N5034, N5023, N1516, N2060);
xor XOR2 (N5035, N5014, N2544);
nand NAND3 (N5036, N5000, N4168, N3371);
or OR2 (N5037, N5033, N3585);
buf BUF1 (N5038, N5036);
nor NOR2 (N5039, N5031, N4536);
or OR3 (N5040, N5037, N3623, N4823);
xor XOR2 (N5041, N5035, N3353);
and AND4 (N5042, N5039, N563, N333, N2532);
nand NAND3 (N5043, N5040, N912, N2237);
and AND2 (N5044, N5043, N1815);
buf BUF1 (N5045, N5042);
not NOT1 (N5046, N5041);
xor XOR2 (N5047, N5024, N599);
or OR4 (N5048, N5047, N2658, N1952, N739);
not NOT1 (N5049, N5046);
nand NAND2 (N5050, N5048, N698);
nand NAND2 (N5051, N5050, N2617);
nor NOR3 (N5052, N5028, N718, N807);
nand NAND3 (N5053, N5032, N581, N1977);
and AND2 (N5054, N5053, N1672);
nand NAND3 (N5055, N5054, N2127, N2544);
nor NOR3 (N5056, N5045, N4122, N4618);
xor XOR2 (N5057, N5044, N1596);
xor XOR2 (N5058, N5052, N4967);
nand NAND3 (N5059, N5034, N4788, N3847);
buf BUF1 (N5060, N5038);
xor XOR2 (N5061, N5056, N2964);
nor NOR3 (N5062, N5057, N688, N3351);
nor NOR3 (N5063, N5062, N1584, N12);
not NOT1 (N5064, N5051);
not NOT1 (N5065, N5059);
buf BUF1 (N5066, N5060);
buf BUF1 (N5067, N5063);
nand NAND2 (N5068, N5065, N1602);
buf BUF1 (N5069, N5068);
and AND4 (N5070, N5055, N2241, N2835, N2945);
not NOT1 (N5071, N5049);
not NOT1 (N5072, N5064);
xor XOR2 (N5073, N5066, N2339);
or OR2 (N5074, N5071, N1078);
not NOT1 (N5075, N5074);
buf BUF1 (N5076, N5070);
xor XOR2 (N5077, N5061, N2354);
nor NOR4 (N5078, N5029, N2372, N3173, N2248);
and AND3 (N5079, N5076, N595, N4918);
nor NOR4 (N5080, N5069, N3840, N772, N1703);
buf BUF1 (N5081, N5058);
nand NAND2 (N5082, N5073, N4263);
and AND4 (N5083, N5079, N2249, N68, N872);
not NOT1 (N5084, N5081);
nand NAND4 (N5085, N5082, N154, N2341, N3402);
xor XOR2 (N5086, N5007, N3127);
buf BUF1 (N5087, N5084);
nor NOR2 (N5088, N5083, N3886);
and AND4 (N5089, N5087, N1258, N1056, N3009);
and AND3 (N5090, N5075, N3227, N4870);
nand NAND4 (N5091, N5089, N2763, N2092, N1270);
buf BUF1 (N5092, N5086);
not NOT1 (N5093, N5092);
not NOT1 (N5094, N5091);
nor NOR2 (N5095, N5093, N4724);
nor NOR3 (N5096, N5085, N1922, N3464);
buf BUF1 (N5097, N5072);
and AND3 (N5098, N5078, N3206, N693);
not NOT1 (N5099, N5077);
not NOT1 (N5100, N5090);
xor XOR2 (N5101, N5096, N2364);
or OR2 (N5102, N5100, N2448);
or OR4 (N5103, N5088, N2997, N3218, N2493);
or OR3 (N5104, N5103, N1347, N288);
not NOT1 (N5105, N5099);
not NOT1 (N5106, N5094);
nor NOR2 (N5107, N5105, N1515);
and AND2 (N5108, N5102, N553);
nand NAND2 (N5109, N5098, N2366);
or OR4 (N5110, N5104, N888, N3182, N4292);
and AND4 (N5111, N5095, N4974, N4210, N4505);
not NOT1 (N5112, N5109);
xor XOR2 (N5113, N5106, N506);
and AND2 (N5114, N5110, N2102);
not NOT1 (N5115, N5107);
nor NOR4 (N5116, N5111, N3389, N64, N4608);
and AND4 (N5117, N5067, N1073, N4299, N967);
xor XOR2 (N5118, N5115, N1625);
buf BUF1 (N5119, N5114);
xor XOR2 (N5120, N5112, N320);
not NOT1 (N5121, N5113);
and AND2 (N5122, N5120, N2387);
not NOT1 (N5123, N5122);
nor NOR3 (N5124, N5108, N537, N3116);
and AND4 (N5125, N5080, N3107, N1405, N1673);
not NOT1 (N5126, N5117);
xor XOR2 (N5127, N5121, N3589);
buf BUF1 (N5128, N5126);
nor NOR3 (N5129, N5123, N548, N1394);
or OR3 (N5130, N5118, N1004, N608);
nor NOR2 (N5131, N5125, N3072);
xor XOR2 (N5132, N5127, N3503);
not NOT1 (N5133, N5129);
xor XOR2 (N5134, N5101, N280);
xor XOR2 (N5135, N5131, N2447);
and AND3 (N5136, N5119, N3703, N3138);
or OR3 (N5137, N5124, N3006, N3387);
not NOT1 (N5138, N5137);
or OR3 (N5139, N5136, N3489, N3376);
nand NAND2 (N5140, N5116, N2636);
nor NOR3 (N5141, N5130, N2444, N4525);
or OR4 (N5142, N5128, N2970, N3724, N1293);
nor NOR4 (N5143, N5097, N4902, N1726, N424);
xor XOR2 (N5144, N5138, N5120);
or OR4 (N5145, N5135, N3380, N2910, N1685);
and AND3 (N5146, N5134, N4227, N2764);
nand NAND4 (N5147, N5141, N1140, N1182, N1753);
nor NOR4 (N5148, N5144, N4360, N2580, N2419);
not NOT1 (N5149, N5140);
buf BUF1 (N5150, N5132);
buf BUF1 (N5151, N5139);
nand NAND2 (N5152, N5133, N1158);
xor XOR2 (N5153, N5151, N54);
nand NAND3 (N5154, N5152, N1280, N1695);
and AND4 (N5155, N5145, N2261, N2933, N4822);
nand NAND4 (N5156, N5154, N10, N3848, N400);
buf BUF1 (N5157, N5142);
xor XOR2 (N5158, N5147, N4989);
nand NAND2 (N5159, N5143, N3292);
nor NOR4 (N5160, N5148, N3341, N3758, N3889);
nand NAND2 (N5161, N5146, N1378);
xor XOR2 (N5162, N5149, N4712);
buf BUF1 (N5163, N5157);
nand NAND3 (N5164, N5159, N4121, N3294);
nor NOR2 (N5165, N5155, N921);
xor XOR2 (N5166, N5160, N4524);
buf BUF1 (N5167, N5165);
nor NOR4 (N5168, N5158, N4945, N3972, N2109);
not NOT1 (N5169, N5167);
xor XOR2 (N5170, N5150, N2497);
nand NAND3 (N5171, N5156, N2987, N4585);
nand NAND4 (N5172, N5162, N4659, N2678, N4705);
nor NOR2 (N5173, N5166, N2070);
buf BUF1 (N5174, N5170);
or OR3 (N5175, N5153, N5005, N191);
or OR3 (N5176, N5161, N1806, N1437);
buf BUF1 (N5177, N5164);
or OR2 (N5178, N5177, N3241);
nand NAND4 (N5179, N5175, N4283, N2156, N4768);
or OR4 (N5180, N5173, N2466, N4907, N2184);
not NOT1 (N5181, N5169);
xor XOR2 (N5182, N5179, N4950);
nor NOR3 (N5183, N5176, N1691, N1684);
nor NOR4 (N5184, N5168, N1908, N351, N4001);
nor NOR3 (N5185, N5178, N2996, N4148);
or OR4 (N5186, N5182, N5169, N5005, N3107);
and AND4 (N5187, N5185, N5154, N552, N4322);
buf BUF1 (N5188, N5184);
xor XOR2 (N5189, N5188, N4044);
not NOT1 (N5190, N5172);
nor NOR4 (N5191, N5171, N5059, N4111, N3475);
xor XOR2 (N5192, N5190, N3298);
or OR2 (N5193, N5191, N2364);
or OR4 (N5194, N5187, N5124, N2956, N2517);
and AND3 (N5195, N5193, N3955, N2147);
xor XOR2 (N5196, N5163, N1498);
buf BUF1 (N5197, N5194);
and AND2 (N5198, N5183, N1940);
nand NAND2 (N5199, N5180, N4125);
not NOT1 (N5200, N5195);
and AND4 (N5201, N5196, N2251, N4687, N3327);
nor NOR3 (N5202, N5198, N2587, N3186);
or OR3 (N5203, N5174, N818, N3697);
not NOT1 (N5204, N5200);
not NOT1 (N5205, N5201);
not NOT1 (N5206, N5192);
nor NOR2 (N5207, N5202, N485);
nand NAND2 (N5208, N5203, N5109);
or OR3 (N5209, N5204, N301, N2019);
or OR4 (N5210, N5208, N611, N2245, N718);
buf BUF1 (N5211, N5205);
not NOT1 (N5212, N5199);
xor XOR2 (N5213, N5211, N3322);
or OR3 (N5214, N5209, N771, N1619);
nor NOR4 (N5215, N5197, N4642, N3562, N2551);
or OR2 (N5216, N5215, N655);
or OR3 (N5217, N5214, N1205, N4463);
buf BUF1 (N5218, N5210);
nor NOR2 (N5219, N5213, N689);
buf BUF1 (N5220, N5219);
xor XOR2 (N5221, N5189, N1155);
buf BUF1 (N5222, N5216);
xor XOR2 (N5223, N5212, N55);
not NOT1 (N5224, N5220);
xor XOR2 (N5225, N5207, N720);
buf BUF1 (N5226, N5223);
buf BUF1 (N5227, N5217);
or OR2 (N5228, N5226, N2030);
not NOT1 (N5229, N5221);
nor NOR3 (N5230, N5225, N23, N4934);
xor XOR2 (N5231, N5206, N288);
nand NAND3 (N5232, N5229, N3204, N2511);
nor NOR3 (N5233, N5227, N1403, N1526);
and AND4 (N5234, N5181, N50, N4324, N1843);
not NOT1 (N5235, N5231);
nand NAND3 (N5236, N5233, N2506, N2732);
xor XOR2 (N5237, N5232, N254);
and AND4 (N5238, N5186, N2927, N566, N3954);
or OR4 (N5239, N5218, N895, N4654, N2185);
and AND2 (N5240, N5238, N1814);
xor XOR2 (N5241, N5224, N4878);
or OR2 (N5242, N5241, N4522);
buf BUF1 (N5243, N5236);
and AND4 (N5244, N5239, N1370, N3037, N320);
and AND4 (N5245, N5240, N4892, N5111, N810);
xor XOR2 (N5246, N5234, N3325);
or OR3 (N5247, N5245, N804, N632);
and AND4 (N5248, N5246, N945, N1893, N4846);
or OR3 (N5249, N5230, N1205, N4826);
or OR3 (N5250, N5249, N4194, N4116);
xor XOR2 (N5251, N5237, N3832);
and AND3 (N5252, N5243, N2082, N1624);
or OR2 (N5253, N5244, N3474);
nand NAND4 (N5254, N5251, N1488, N4111, N4380);
nand NAND2 (N5255, N5222, N975);
not NOT1 (N5256, N5242);
xor XOR2 (N5257, N5252, N3506);
not NOT1 (N5258, N5255);
buf BUF1 (N5259, N5248);
xor XOR2 (N5260, N5235, N1720);
and AND4 (N5261, N5257, N3953, N2529, N874);
nor NOR2 (N5262, N5250, N4671);
xor XOR2 (N5263, N5253, N3006);
not NOT1 (N5264, N5260);
or OR3 (N5265, N5256, N711, N2744);
buf BUF1 (N5266, N5263);
nand NAND4 (N5267, N5261, N4929, N2648, N2724);
or OR2 (N5268, N5259, N676);
or OR3 (N5269, N5267, N5136, N4963);
and AND4 (N5270, N5247, N867, N1974, N1077);
nor NOR4 (N5271, N5265, N3879, N4309, N5167);
buf BUF1 (N5272, N5254);
or OR3 (N5273, N5228, N3593, N3168);
nand NAND3 (N5274, N5268, N1480, N2233);
nor NOR4 (N5275, N5270, N1415, N1594, N4040);
and AND4 (N5276, N5271, N1594, N3962, N4782);
xor XOR2 (N5277, N5258, N2406);
or OR4 (N5278, N5273, N2166, N2167, N612);
xor XOR2 (N5279, N5266, N2607);
or OR4 (N5280, N5277, N3722, N1851, N2239);
or OR2 (N5281, N5278, N3703);
buf BUF1 (N5282, N5281);
xor XOR2 (N5283, N5269, N1198);
or OR4 (N5284, N5274, N2630, N1890, N4739);
or OR3 (N5285, N5284, N962, N4559);
nor NOR2 (N5286, N5283, N3962);
nand NAND3 (N5287, N5272, N1530, N2446);
or OR2 (N5288, N5287, N4594);
xor XOR2 (N5289, N5285, N5125);
and AND3 (N5290, N5280, N339, N4718);
buf BUF1 (N5291, N5282);
buf BUF1 (N5292, N5286);
and AND3 (N5293, N5291, N4509, N4752);
not NOT1 (N5294, N5289);
and AND2 (N5295, N5279, N275);
xor XOR2 (N5296, N5276, N3797);
buf BUF1 (N5297, N5262);
nor NOR3 (N5298, N5290, N3593, N4449);
buf BUF1 (N5299, N5298);
xor XOR2 (N5300, N5293, N3682);
and AND2 (N5301, N5292, N2377);
nor NOR2 (N5302, N5264, N1956);
or OR3 (N5303, N5299, N4590, N4141);
buf BUF1 (N5304, N5301);
buf BUF1 (N5305, N5303);
nand NAND2 (N5306, N5304, N1649);
nor NOR2 (N5307, N5294, N1881);
buf BUF1 (N5308, N5295);
nor NOR4 (N5309, N5288, N3777, N4702, N5240);
or OR4 (N5310, N5296, N3863, N2625, N1700);
nand NAND2 (N5311, N5306, N199);
buf BUF1 (N5312, N5305);
xor XOR2 (N5313, N5297, N1348);
and AND4 (N5314, N5307, N3324, N3280, N83);
and AND3 (N5315, N5300, N5271, N255);
or OR2 (N5316, N5313, N418);
or OR3 (N5317, N5310, N3269, N3776);
not NOT1 (N5318, N5302);
nand NAND4 (N5319, N5318, N4409, N1414, N3475);
nand NAND4 (N5320, N5308, N322, N541, N542);
not NOT1 (N5321, N5314);
not NOT1 (N5322, N5315);
nand NAND2 (N5323, N5322, N3284);
xor XOR2 (N5324, N5311, N345);
or OR2 (N5325, N5275, N3593);
and AND2 (N5326, N5320, N3698);
buf BUF1 (N5327, N5319);
and AND3 (N5328, N5324, N4685, N1086);
buf BUF1 (N5329, N5321);
or OR2 (N5330, N5317, N3337);
or OR3 (N5331, N5325, N726, N3179);
nor NOR3 (N5332, N5328, N4000, N428);
and AND2 (N5333, N5332, N4628);
and AND4 (N5334, N5333, N4041, N1502, N3771);
and AND2 (N5335, N5309, N3330);
xor XOR2 (N5336, N5329, N1808);
buf BUF1 (N5337, N5331);
buf BUF1 (N5338, N5326);
or OR2 (N5339, N5336, N3594);
xor XOR2 (N5340, N5327, N160);
nor NOR2 (N5341, N5338, N688);
nand NAND2 (N5342, N5340, N1358);
or OR2 (N5343, N5339, N5233);
and AND3 (N5344, N5337, N991, N2638);
not NOT1 (N5345, N5312);
and AND3 (N5346, N5345, N4145, N2483);
xor XOR2 (N5347, N5323, N682);
nor NOR3 (N5348, N5330, N569, N1189);
not NOT1 (N5349, N5334);
nand NAND2 (N5350, N5348, N4933);
not NOT1 (N5351, N5347);
nand NAND4 (N5352, N5335, N1326, N1912, N435);
xor XOR2 (N5353, N5343, N2636);
or OR4 (N5354, N5351, N1648, N4664, N666);
and AND2 (N5355, N5341, N4663);
or OR4 (N5356, N5355, N644, N3202, N131);
nor NOR2 (N5357, N5346, N4760);
xor XOR2 (N5358, N5353, N2313);
not NOT1 (N5359, N5350);
nand NAND4 (N5360, N5359, N2250, N3426, N3444);
or OR4 (N5361, N5342, N2072, N1763, N1891);
and AND2 (N5362, N5361, N1270);
xor XOR2 (N5363, N5354, N4540);
nor NOR4 (N5364, N5356, N2459, N1336, N246);
nand NAND4 (N5365, N5349, N787, N3328, N2707);
nand NAND2 (N5366, N5363, N5108);
and AND4 (N5367, N5360, N2492, N567, N1019);
buf BUF1 (N5368, N5352);
not NOT1 (N5369, N5365);
nor NOR3 (N5370, N5364, N312, N3618);
nor NOR4 (N5371, N5316, N810, N4427, N444);
nor NOR3 (N5372, N5367, N2803, N1068);
or OR3 (N5373, N5372, N2864, N324);
not NOT1 (N5374, N5371);
buf BUF1 (N5375, N5344);
not NOT1 (N5376, N5374);
not NOT1 (N5377, N5369);
nor NOR3 (N5378, N5370, N4104, N4948);
nand NAND3 (N5379, N5357, N1114, N2710);
buf BUF1 (N5380, N5362);
or OR4 (N5381, N5375, N4719, N2077, N2554);
xor XOR2 (N5382, N5366, N5041);
and AND3 (N5383, N5358, N2949, N1309);
buf BUF1 (N5384, N5376);
nor NOR4 (N5385, N5377, N2001, N4213, N3260);
buf BUF1 (N5386, N5384);
buf BUF1 (N5387, N5386);
and AND2 (N5388, N5383, N1503);
xor XOR2 (N5389, N5385, N2024);
not NOT1 (N5390, N5380);
xor XOR2 (N5391, N5373, N4672);
or OR4 (N5392, N5381, N3753, N4782, N2971);
not NOT1 (N5393, N5382);
buf BUF1 (N5394, N5379);
or OR2 (N5395, N5390, N2230);
or OR4 (N5396, N5389, N5279, N4981, N2190);
not NOT1 (N5397, N5391);
not NOT1 (N5398, N5395);
not NOT1 (N5399, N5394);
not NOT1 (N5400, N5387);
nand NAND4 (N5401, N5392, N4936, N825, N1708);
not NOT1 (N5402, N5400);
not NOT1 (N5403, N5396);
xor XOR2 (N5404, N5378, N1430);
buf BUF1 (N5405, N5403);
or OR2 (N5406, N5368, N1360);
or OR2 (N5407, N5397, N1108);
nor NOR3 (N5408, N5406, N3337, N832);
nor NOR3 (N5409, N5405, N5221, N5093);
nand NAND2 (N5410, N5398, N2940);
nand NAND3 (N5411, N5402, N586, N428);
or OR4 (N5412, N5411, N949, N1493, N1757);
nand NAND2 (N5413, N5401, N2858);
buf BUF1 (N5414, N5413);
nor NOR3 (N5415, N5393, N4228, N4621);
or OR3 (N5416, N5412, N4417, N722);
nor NOR2 (N5417, N5414, N1984);
xor XOR2 (N5418, N5399, N1736);
and AND3 (N5419, N5410, N1776, N387);
nand NAND3 (N5420, N5418, N3042, N1071);
and AND3 (N5421, N5409, N2880, N2146);
nand NAND4 (N5422, N5415, N2450, N2216, N3117);
nand NAND4 (N5423, N5421, N5236, N2194, N3727);
buf BUF1 (N5424, N5422);
and AND2 (N5425, N5423, N645);
or OR4 (N5426, N5424, N2235, N5112, N5341);
xor XOR2 (N5427, N5426, N2368);
or OR2 (N5428, N5425, N4143);
not NOT1 (N5429, N5420);
buf BUF1 (N5430, N5407);
nor NOR4 (N5431, N5429, N2543, N696, N2992);
buf BUF1 (N5432, N5428);
xor XOR2 (N5433, N5427, N995);
not NOT1 (N5434, N5431);
nor NOR4 (N5435, N5434, N3042, N3018, N908);
buf BUF1 (N5436, N5417);
or OR4 (N5437, N5435, N2870, N1260, N2197);
or OR3 (N5438, N5436, N2621, N4678);
or OR3 (N5439, N5433, N1887, N2193);
or OR4 (N5440, N5432, N1643, N3529, N3227);
buf BUF1 (N5441, N5404);
and AND2 (N5442, N5408, N5290);
and AND2 (N5443, N5438, N2439);
not NOT1 (N5444, N5443);
nand NAND2 (N5445, N5430, N2063);
or OR2 (N5446, N5419, N2167);
buf BUF1 (N5447, N5441);
or OR2 (N5448, N5444, N548);
nor NOR4 (N5449, N5448, N1539, N2945, N1343);
and AND2 (N5450, N5446, N1674);
nor NOR4 (N5451, N5440, N3804, N658, N1825);
nand NAND2 (N5452, N5437, N3390);
or OR2 (N5453, N5445, N2263);
or OR4 (N5454, N5388, N4128, N1230, N4338);
buf BUF1 (N5455, N5453);
not NOT1 (N5456, N5439);
xor XOR2 (N5457, N5447, N338);
buf BUF1 (N5458, N5456);
not NOT1 (N5459, N5451);
xor XOR2 (N5460, N5416, N3461);
or OR3 (N5461, N5457, N3035, N4002);
buf BUF1 (N5462, N5455);
or OR2 (N5463, N5462, N929);
or OR2 (N5464, N5463, N878);
or OR4 (N5465, N5454, N2494, N3791, N1036);
nor NOR4 (N5466, N5460, N1439, N129, N4586);
nand NAND4 (N5467, N5449, N4425, N48, N2808);
buf BUF1 (N5468, N5458);
buf BUF1 (N5469, N5467);
buf BUF1 (N5470, N5469);
not NOT1 (N5471, N5468);
not NOT1 (N5472, N5461);
or OR3 (N5473, N5464, N941, N4393);
and AND3 (N5474, N5472, N3775, N2000);
not NOT1 (N5475, N5459);
and AND4 (N5476, N5473, N3854, N3637, N4860);
nand NAND4 (N5477, N5471, N769, N5353, N5176);
xor XOR2 (N5478, N5470, N1934);
nand NAND3 (N5479, N5475, N200, N5136);
not NOT1 (N5480, N5479);
nor NOR3 (N5481, N5442, N474, N340);
nor NOR3 (N5482, N5476, N4069, N3979);
xor XOR2 (N5483, N5480, N2934);
or OR4 (N5484, N5478, N1698, N629, N2243);
nand NAND4 (N5485, N5483, N1533, N482, N5004);
not NOT1 (N5486, N5482);
not NOT1 (N5487, N5450);
buf BUF1 (N5488, N5477);
or OR2 (N5489, N5452, N3655);
nand NAND2 (N5490, N5481, N824);
or OR4 (N5491, N5465, N4783, N2847, N4909);
and AND2 (N5492, N5486, N3746);
nor NOR3 (N5493, N5466, N4022, N4886);
and AND3 (N5494, N5490, N100, N3642);
nand NAND4 (N5495, N5488, N103, N2861, N1527);
or OR2 (N5496, N5485, N974);
nor NOR2 (N5497, N5492, N1859);
nor NOR3 (N5498, N5497, N1080, N4844);
xor XOR2 (N5499, N5496, N271);
buf BUF1 (N5500, N5499);
xor XOR2 (N5501, N5474, N2653);
xor XOR2 (N5502, N5495, N4079);
and AND3 (N5503, N5501, N3869, N1508);
xor XOR2 (N5504, N5502, N4409);
nand NAND4 (N5505, N5493, N5417, N4917, N5031);
and AND2 (N5506, N5503, N785);
nand NAND2 (N5507, N5504, N5057);
xor XOR2 (N5508, N5487, N5473);
xor XOR2 (N5509, N5489, N4053);
not NOT1 (N5510, N5508);
and AND2 (N5511, N5510, N4723);
buf BUF1 (N5512, N5500);
or OR2 (N5513, N5512, N1357);
buf BUF1 (N5514, N5491);
nand NAND2 (N5515, N5509, N1533);
or OR3 (N5516, N5505, N3416, N640);
not NOT1 (N5517, N5484);
and AND2 (N5518, N5507, N3730);
not NOT1 (N5519, N5513);
not NOT1 (N5520, N5514);
or OR3 (N5521, N5516, N5163, N599);
not NOT1 (N5522, N5517);
and AND3 (N5523, N5498, N536, N5183);
and AND4 (N5524, N5520, N3240, N1988, N4307);
not NOT1 (N5525, N5515);
nor NOR2 (N5526, N5511, N3898);
not NOT1 (N5527, N5522);
nor NOR2 (N5528, N5524, N3219);
and AND3 (N5529, N5506, N2821, N3839);
and AND3 (N5530, N5521, N2985, N3845);
or OR2 (N5531, N5519, N1942);
xor XOR2 (N5532, N5494, N2539);
nand NAND2 (N5533, N5528, N133);
not NOT1 (N5534, N5526);
buf BUF1 (N5535, N5529);
or OR3 (N5536, N5530, N2626, N2122);
not NOT1 (N5537, N5533);
xor XOR2 (N5538, N5532, N663);
buf BUF1 (N5539, N5535);
buf BUF1 (N5540, N5531);
and AND2 (N5541, N5537, N3239);
xor XOR2 (N5542, N5518, N2637);
not NOT1 (N5543, N5536);
nand NAND2 (N5544, N5543, N3136);
nor NOR2 (N5545, N5544, N122);
nand NAND2 (N5546, N5527, N5397);
and AND4 (N5547, N5538, N1622, N3676, N434);
buf BUF1 (N5548, N5534);
nand NAND3 (N5549, N5547, N1984, N886);
and AND2 (N5550, N5542, N1880);
not NOT1 (N5551, N5540);
buf BUF1 (N5552, N5546);
xor XOR2 (N5553, N5545, N4666);
buf BUF1 (N5554, N5541);
or OR3 (N5555, N5539, N3845, N3809);
not NOT1 (N5556, N5552);
and AND4 (N5557, N5556, N1962, N3274, N973);
and AND3 (N5558, N5550, N3418, N4943);
xor XOR2 (N5559, N5548, N2962);
or OR2 (N5560, N5555, N2772);
buf BUF1 (N5561, N5560);
buf BUF1 (N5562, N5561);
and AND2 (N5563, N5551, N1853);
or OR2 (N5564, N5562, N4824);
not NOT1 (N5565, N5563);
and AND3 (N5566, N5553, N4874, N2248);
or OR3 (N5567, N5523, N2720, N364);
nor NOR3 (N5568, N5559, N2854, N4659);
buf BUF1 (N5569, N5564);
xor XOR2 (N5570, N5567, N4933);
xor XOR2 (N5571, N5549, N4882);
and AND2 (N5572, N5568, N1828);
nor NOR4 (N5573, N5572, N1079, N4079, N5188);
nand NAND4 (N5574, N5554, N3582, N1464, N445);
nor NOR2 (N5575, N5573, N5263);
or OR4 (N5576, N5574, N3105, N4894, N871);
xor XOR2 (N5577, N5525, N1358);
not NOT1 (N5578, N5577);
nor NOR3 (N5579, N5575, N2359, N3993);
xor XOR2 (N5580, N5578, N4594);
or OR4 (N5581, N5571, N4799, N5158, N646);
buf BUF1 (N5582, N5557);
nand NAND2 (N5583, N5580, N3068);
or OR4 (N5584, N5581, N5016, N241, N3863);
buf BUF1 (N5585, N5569);
nor NOR3 (N5586, N5576, N3973, N5447);
xor XOR2 (N5587, N5565, N3677);
nor NOR2 (N5588, N5566, N2212);
buf BUF1 (N5589, N5583);
not NOT1 (N5590, N5588);
and AND4 (N5591, N5584, N1472, N465, N3969);
not NOT1 (N5592, N5582);
or OR4 (N5593, N5589, N1150, N1779, N4525);
not NOT1 (N5594, N5593);
not NOT1 (N5595, N5585);
nand NAND4 (N5596, N5586, N5594, N5082, N1907);
xor XOR2 (N5597, N3197, N618);
nand NAND4 (N5598, N5579, N2825, N2435, N5169);
nor NOR4 (N5599, N5592, N3002, N1702, N1119);
nor NOR4 (N5600, N5587, N5049, N905, N1797);
not NOT1 (N5601, N5591);
nand NAND4 (N5602, N5596, N4462, N4492, N4866);
or OR2 (N5603, N5599, N2683);
not NOT1 (N5604, N5590);
not NOT1 (N5605, N5570);
and AND4 (N5606, N5600, N3269, N551, N2016);
nand NAND2 (N5607, N5605, N5485);
not NOT1 (N5608, N5606);
xor XOR2 (N5609, N5558, N2508);
buf BUF1 (N5610, N5598);
nand NAND4 (N5611, N5608, N4758, N4149, N472);
xor XOR2 (N5612, N5611, N157);
xor XOR2 (N5613, N5612, N314);
or OR4 (N5614, N5613, N5609, N3390, N1664);
nand NAND3 (N5615, N524, N2316, N3803);
and AND2 (N5616, N5602, N2284);
buf BUF1 (N5617, N5601);
nand NAND4 (N5618, N5615, N3472, N168, N2528);
buf BUF1 (N5619, N5603);
nand NAND3 (N5620, N5604, N2080, N2815);
buf BUF1 (N5621, N5614);
xor XOR2 (N5622, N5619, N2239);
not NOT1 (N5623, N5622);
buf BUF1 (N5624, N5597);
buf BUF1 (N5625, N5610);
and AND4 (N5626, N5620, N4223, N1351, N407);
buf BUF1 (N5627, N5625);
nand NAND4 (N5628, N5624, N2595, N5427, N2073);
nand NAND2 (N5629, N5617, N736);
and AND3 (N5630, N5623, N4445, N416);
or OR2 (N5631, N5629, N2392);
nand NAND4 (N5632, N5621, N2242, N4297, N1075);
or OR4 (N5633, N5616, N2970, N3049, N907);
buf BUF1 (N5634, N5633);
not NOT1 (N5635, N5607);
nand NAND4 (N5636, N5634, N47, N5040, N3954);
or OR4 (N5637, N5626, N1845, N834, N4810);
and AND4 (N5638, N5595, N3604, N2179, N3698);
and AND4 (N5639, N5635, N4686, N2284, N3891);
xor XOR2 (N5640, N5631, N713);
and AND3 (N5641, N5628, N1203, N4226);
xor XOR2 (N5642, N5636, N5267);
nor NOR2 (N5643, N5642, N1261);
xor XOR2 (N5644, N5618, N2359);
not NOT1 (N5645, N5643);
buf BUF1 (N5646, N5638);
not NOT1 (N5647, N5645);
buf BUF1 (N5648, N5646);
nor NOR2 (N5649, N5639, N3656);
nor NOR4 (N5650, N5632, N1368, N4391, N2185);
nor NOR2 (N5651, N5644, N3941);
not NOT1 (N5652, N5648);
and AND2 (N5653, N5627, N1534);
buf BUF1 (N5654, N5650);
xor XOR2 (N5655, N5651, N1447);
and AND4 (N5656, N5654, N5119, N461, N145);
nor NOR4 (N5657, N5630, N2555, N3650, N3425);
nor NOR3 (N5658, N5655, N4874, N4266);
nor NOR3 (N5659, N5653, N1562, N4750);
nand NAND4 (N5660, N5658, N1540, N3472, N4679);
or OR3 (N5661, N5640, N724, N599);
and AND4 (N5662, N5659, N4241, N5437, N1650);
nand NAND3 (N5663, N5652, N3649, N310);
nor NOR4 (N5664, N5649, N5152, N4365, N1409);
nor NOR4 (N5665, N5664, N4536, N894, N246);
nand NAND2 (N5666, N5662, N3006);
or OR3 (N5667, N5641, N4048, N5231);
not NOT1 (N5668, N5656);
nand NAND2 (N5669, N5637, N5198);
nand NAND2 (N5670, N5657, N3954);
nand NAND4 (N5671, N5667, N3916, N161, N686);
nand NAND2 (N5672, N5669, N1902);
xor XOR2 (N5673, N5663, N1559);
xor XOR2 (N5674, N5673, N921);
or OR3 (N5675, N5660, N4301, N1957);
nor NOR2 (N5676, N5668, N4833);
xor XOR2 (N5677, N5670, N2359);
nor NOR3 (N5678, N5672, N4189, N1976);
xor XOR2 (N5679, N5678, N4371);
buf BUF1 (N5680, N5647);
nand NAND3 (N5681, N5679, N297, N4582);
not NOT1 (N5682, N5665);
xor XOR2 (N5683, N5675, N349);
or OR2 (N5684, N5661, N3516);
or OR4 (N5685, N5683, N4008, N1550, N788);
nor NOR3 (N5686, N5676, N1379, N2937);
and AND4 (N5687, N5671, N2347, N1449, N1450);
not NOT1 (N5688, N5681);
nor NOR4 (N5689, N5684, N5360, N3711, N5369);
xor XOR2 (N5690, N5687, N1787);
or OR3 (N5691, N5686, N1851, N3626);
and AND4 (N5692, N5685, N3935, N658, N1436);
and AND3 (N5693, N5682, N2987, N2249);
and AND4 (N5694, N5692, N5638, N4083, N724);
nand NAND3 (N5695, N5689, N3395, N2661);
or OR2 (N5696, N5680, N1040);
xor XOR2 (N5697, N5691, N460);
or OR3 (N5698, N5697, N3257, N3452);
not NOT1 (N5699, N5694);
and AND2 (N5700, N5677, N1578);
and AND4 (N5701, N5688, N2104, N3647, N1579);
xor XOR2 (N5702, N5690, N1552);
nand NAND3 (N5703, N5700, N2761, N1791);
nor NOR3 (N5704, N5698, N1184, N3774);
nand NAND4 (N5705, N5702, N4934, N5306, N3885);
xor XOR2 (N5706, N5704, N2646);
buf BUF1 (N5707, N5701);
not NOT1 (N5708, N5674);
xor XOR2 (N5709, N5703, N1754);
nor NOR3 (N5710, N5705, N2271, N3707);
xor XOR2 (N5711, N5709, N2104);
not NOT1 (N5712, N5699);
and AND2 (N5713, N5712, N1296);
xor XOR2 (N5714, N5711, N5367);
nand NAND2 (N5715, N5693, N5230);
or OR3 (N5716, N5710, N3756, N579);
and AND3 (N5717, N5695, N3054, N305);
xor XOR2 (N5718, N5666, N5600);
buf BUF1 (N5719, N5714);
buf BUF1 (N5720, N5713);
buf BUF1 (N5721, N5696);
buf BUF1 (N5722, N5720);
not NOT1 (N5723, N5722);
buf BUF1 (N5724, N5708);
or OR2 (N5725, N5718, N3719);
not NOT1 (N5726, N5716);
not NOT1 (N5727, N5715);
and AND2 (N5728, N5717, N257);
buf BUF1 (N5729, N5724);
nand NAND4 (N5730, N5721, N1928, N4218, N4650);
nor NOR3 (N5731, N5719, N905, N938);
not NOT1 (N5732, N5728);
not NOT1 (N5733, N5730);
nand NAND3 (N5734, N5729, N4436, N474);
nor NOR4 (N5735, N5727, N4181, N2125, N1313);
nor NOR2 (N5736, N5732, N1064);
and AND4 (N5737, N5733, N3932, N2884, N282);
and AND4 (N5738, N5723, N852, N3726, N2659);
nor NOR2 (N5739, N5706, N1954);
xor XOR2 (N5740, N5726, N2899);
xor XOR2 (N5741, N5731, N3434);
xor XOR2 (N5742, N5738, N3683);
not NOT1 (N5743, N5736);
not NOT1 (N5744, N5743);
or OR3 (N5745, N5737, N2785, N2895);
and AND3 (N5746, N5734, N3553, N2972);
buf BUF1 (N5747, N5725);
buf BUF1 (N5748, N5746);
nand NAND4 (N5749, N5744, N4354, N4946, N5567);
not NOT1 (N5750, N5742);
and AND2 (N5751, N5748, N4591);
and AND2 (N5752, N5747, N2077);
buf BUF1 (N5753, N5750);
not NOT1 (N5754, N5751);
buf BUF1 (N5755, N5735);
xor XOR2 (N5756, N5707, N3054);
xor XOR2 (N5757, N5745, N1341);
or OR3 (N5758, N5755, N4207, N4811);
or OR3 (N5759, N5741, N4088, N843);
buf BUF1 (N5760, N5754);
xor XOR2 (N5761, N5753, N3018);
nand NAND4 (N5762, N5759, N1319, N496, N1155);
or OR4 (N5763, N5756, N4256, N3095, N4325);
not NOT1 (N5764, N5763);
or OR3 (N5765, N5752, N805, N2952);
nand NAND4 (N5766, N5758, N3884, N4537, N3521);
nor NOR3 (N5767, N5757, N3457, N3338);
or OR4 (N5768, N5765, N5156, N5137, N1761);
and AND4 (N5769, N5762, N999, N4526, N4680);
buf BUF1 (N5770, N5739);
buf BUF1 (N5771, N5766);
xor XOR2 (N5772, N5767, N3787);
not NOT1 (N5773, N5769);
xor XOR2 (N5774, N5761, N2615);
not NOT1 (N5775, N5740);
xor XOR2 (N5776, N5760, N3117);
or OR2 (N5777, N5764, N1624);
nor NOR2 (N5778, N5777, N2874);
or OR3 (N5779, N5770, N4715, N3105);
not NOT1 (N5780, N5768);
nand NAND3 (N5781, N5775, N4794, N4492);
xor XOR2 (N5782, N5771, N4837);
not NOT1 (N5783, N5779);
nand NAND4 (N5784, N5776, N836, N2906, N1674);
buf BUF1 (N5785, N5781);
nor NOR4 (N5786, N5749, N2063, N850, N4626);
not NOT1 (N5787, N5782);
xor XOR2 (N5788, N5772, N1525);
nor NOR4 (N5789, N5780, N656, N5172, N3400);
xor XOR2 (N5790, N5786, N4883);
and AND2 (N5791, N5788, N4360);
or OR3 (N5792, N5783, N69, N2252);
nor NOR2 (N5793, N5790, N2902);
buf BUF1 (N5794, N5774);
not NOT1 (N5795, N5794);
not NOT1 (N5796, N5795);
nand NAND2 (N5797, N5787, N5326);
and AND3 (N5798, N5785, N2517, N1745);
nor NOR2 (N5799, N5796, N5598);
buf BUF1 (N5800, N5791);
or OR4 (N5801, N5784, N706, N3004, N3299);
nand NAND4 (N5802, N5773, N564, N3162, N2723);
nor NOR3 (N5803, N5789, N3594, N5606);
xor XOR2 (N5804, N5802, N3858);
xor XOR2 (N5805, N5778, N5163);
nand NAND2 (N5806, N5793, N1704);
and AND2 (N5807, N5803, N5706);
xor XOR2 (N5808, N5797, N646);
nand NAND2 (N5809, N5792, N3279);
nand NAND3 (N5810, N5807, N1147, N1704);
nor NOR4 (N5811, N5808, N5499, N1278, N279);
or OR2 (N5812, N5804, N887);
not NOT1 (N5813, N5812);
not NOT1 (N5814, N5813);
nor NOR2 (N5815, N5814, N906);
and AND3 (N5816, N5809, N4592, N2890);
nand NAND2 (N5817, N5811, N1099);
not NOT1 (N5818, N5801);
buf BUF1 (N5819, N5800);
or OR3 (N5820, N5810, N5819, N1877);
nor NOR2 (N5821, N2221, N2947);
xor XOR2 (N5822, N5817, N2155);
or OR4 (N5823, N5818, N1622, N2897, N2725);
xor XOR2 (N5824, N5816, N1027);
nand NAND3 (N5825, N5824, N4627, N4476);
or OR3 (N5826, N5823, N3521, N2606);
or OR4 (N5827, N5815, N4282, N3049, N4934);
nor NOR2 (N5828, N5826, N2563);
xor XOR2 (N5829, N5821, N1353);
nor NOR2 (N5830, N5820, N686);
or OR3 (N5831, N5825, N5743, N5133);
and AND3 (N5832, N5798, N3722, N4541);
not NOT1 (N5833, N5822);
buf BUF1 (N5834, N5828);
and AND4 (N5835, N5834, N4539, N4944, N945);
and AND2 (N5836, N5827, N2279);
nand NAND2 (N5837, N5799, N2932);
nor NOR3 (N5838, N5832, N492, N2339);
nor NOR3 (N5839, N5833, N123, N5065);
not NOT1 (N5840, N5838);
and AND4 (N5841, N5835, N213, N4904, N2749);
and AND2 (N5842, N5806, N2264);
not NOT1 (N5843, N5841);
nor NOR2 (N5844, N5836, N4954);
not NOT1 (N5845, N5831);
not NOT1 (N5846, N5843);
and AND4 (N5847, N5839, N4131, N5346, N4402);
or OR3 (N5848, N5837, N3490, N3770);
not NOT1 (N5849, N5844);
or OR2 (N5850, N5842, N5082);
and AND4 (N5851, N5829, N3734, N4916, N5073);
xor XOR2 (N5852, N5830, N2124);
not NOT1 (N5853, N5805);
not NOT1 (N5854, N5846);
buf BUF1 (N5855, N5850);
xor XOR2 (N5856, N5853, N1421);
not NOT1 (N5857, N5849);
or OR3 (N5858, N5857, N1885, N5011);
xor XOR2 (N5859, N5851, N1605);
and AND3 (N5860, N5856, N2399, N2021);
xor XOR2 (N5861, N5852, N1531);
nor NOR3 (N5862, N5855, N2453, N4236);
nand NAND2 (N5863, N5848, N2218);
nand NAND2 (N5864, N5859, N4859);
not NOT1 (N5865, N5861);
nor NOR2 (N5866, N5863, N4648);
xor XOR2 (N5867, N5860, N3260);
xor XOR2 (N5868, N5845, N4192);
and AND2 (N5869, N5858, N4916);
or OR4 (N5870, N5862, N3232, N3149, N2783);
nor NOR4 (N5871, N5869, N999, N955, N4956);
buf BUF1 (N5872, N5870);
buf BUF1 (N5873, N5865);
xor XOR2 (N5874, N5866, N3386);
xor XOR2 (N5875, N5868, N5439);
nor NOR4 (N5876, N5847, N5565, N2836, N4078);
buf BUF1 (N5877, N5872);
xor XOR2 (N5878, N5840, N4525);
buf BUF1 (N5879, N5873);
or OR4 (N5880, N5879, N870, N1242, N3676);
nor NOR4 (N5881, N5878, N5302, N1587, N4426);
buf BUF1 (N5882, N5876);
nor NOR4 (N5883, N5874, N1822, N4613, N5105);
nor NOR2 (N5884, N5871, N4102);
and AND4 (N5885, N5867, N139, N2326, N104);
not NOT1 (N5886, N5877);
buf BUF1 (N5887, N5886);
or OR2 (N5888, N5883, N5075);
or OR2 (N5889, N5887, N3416);
and AND4 (N5890, N5884, N4187, N5223, N2189);
buf BUF1 (N5891, N5880);
or OR2 (N5892, N5891, N626);
buf BUF1 (N5893, N5885);
and AND3 (N5894, N5882, N434, N2660);
nor NOR3 (N5895, N5881, N422, N4473);
xor XOR2 (N5896, N5895, N4123);
not NOT1 (N5897, N5888);
buf BUF1 (N5898, N5892);
nand NAND2 (N5899, N5893, N3875);
or OR2 (N5900, N5896, N5205);
xor XOR2 (N5901, N5889, N4526);
not NOT1 (N5902, N5854);
xor XOR2 (N5903, N5897, N241);
xor XOR2 (N5904, N5901, N2490);
nor NOR4 (N5905, N5890, N885, N3224, N811);
buf BUF1 (N5906, N5864);
nand NAND3 (N5907, N5898, N4333, N3995);
not NOT1 (N5908, N5894);
xor XOR2 (N5909, N5907, N1735);
and AND4 (N5910, N5903, N516, N3946, N1610);
and AND2 (N5911, N5900, N5346);
buf BUF1 (N5912, N5909);
not NOT1 (N5913, N5906);
or OR4 (N5914, N5899, N5752, N5676, N2609);
or OR4 (N5915, N5914, N1783, N2691, N103);
xor XOR2 (N5916, N5905, N3285);
and AND2 (N5917, N5913, N1472);
nand NAND3 (N5918, N5916, N4763, N3491);
nor NOR4 (N5919, N5912, N1880, N1179, N2547);
and AND3 (N5920, N5904, N2965, N1913);
and AND4 (N5921, N5917, N2887, N4776, N3614);
and AND2 (N5922, N5910, N4400);
nor NOR2 (N5923, N5915, N361);
nand NAND3 (N5924, N5921, N3098, N485);
or OR4 (N5925, N5922, N1715, N2356, N4568);
buf BUF1 (N5926, N5923);
buf BUF1 (N5927, N5918);
buf BUF1 (N5928, N5920);
xor XOR2 (N5929, N5927, N3615);
not NOT1 (N5930, N5925);
or OR2 (N5931, N5924, N2596);
xor XOR2 (N5932, N5931, N215);
or OR2 (N5933, N5932, N2618);
xor XOR2 (N5934, N5902, N1979);
xor XOR2 (N5935, N5875, N519);
xor XOR2 (N5936, N5933, N5469);
nand NAND3 (N5937, N5928, N5501, N4489);
or OR4 (N5938, N5911, N2196, N1571, N46);
xor XOR2 (N5939, N5937, N5477);
not NOT1 (N5940, N5926);
nand NAND3 (N5941, N5929, N4, N4863);
nor NOR3 (N5942, N5936, N1162, N273);
nor NOR4 (N5943, N5935, N5560, N687, N3568);
buf BUF1 (N5944, N5908);
and AND4 (N5945, N5944, N2223, N1903, N4001);
nand NAND3 (N5946, N5919, N1845, N2386);
not NOT1 (N5947, N5930);
nor NOR3 (N5948, N5934, N919, N2729);
nand NAND4 (N5949, N5941, N3857, N73, N2826);
xor XOR2 (N5950, N5938, N34);
nand NAND2 (N5951, N5948, N4542);
buf BUF1 (N5952, N5949);
not NOT1 (N5953, N5940);
nand NAND3 (N5954, N5946, N897, N1245);
and AND4 (N5955, N5953, N818, N5794, N3768);
xor XOR2 (N5956, N5943, N2474);
xor XOR2 (N5957, N5952, N4281);
buf BUF1 (N5958, N5950);
or OR4 (N5959, N5958, N3822, N2696, N2176);
not NOT1 (N5960, N5956);
nand NAND4 (N5961, N5957, N1712, N1398, N891);
xor XOR2 (N5962, N5951, N3055);
xor XOR2 (N5963, N5961, N3276);
xor XOR2 (N5964, N5939, N441);
or OR3 (N5965, N5964, N836, N2022);
xor XOR2 (N5966, N5945, N4420);
not NOT1 (N5967, N5962);
and AND2 (N5968, N5960, N906);
nand NAND2 (N5969, N5965, N2952);
xor XOR2 (N5970, N5968, N344);
nand NAND4 (N5971, N5959, N5751, N955, N2378);
not NOT1 (N5972, N5955);
and AND4 (N5973, N5972, N3014, N5871, N4677);
nor NOR3 (N5974, N5963, N557, N994);
nor NOR3 (N5975, N5970, N4733, N1898);
or OR2 (N5976, N5967, N608);
nand NAND2 (N5977, N5973, N21);
nor NOR2 (N5978, N5974, N5332);
xor XOR2 (N5979, N5942, N1632);
or OR4 (N5980, N5979, N5420, N2537, N3977);
nor NOR2 (N5981, N5971, N2115);
or OR2 (N5982, N5954, N3462);
nor NOR4 (N5983, N5947, N5764, N3050, N4930);
nor NOR3 (N5984, N5982, N2929, N3397);
buf BUF1 (N5985, N5984);
and AND4 (N5986, N5978, N1219, N4591, N3836);
or OR2 (N5987, N5985, N3855);
nor NOR2 (N5988, N5966, N4404);
and AND3 (N5989, N5977, N4518, N236);
and AND3 (N5990, N5983, N4749, N2010);
or OR2 (N5991, N5987, N977);
nor NOR2 (N5992, N5988, N2008);
buf BUF1 (N5993, N5992);
and AND2 (N5994, N5981, N215);
or OR2 (N5995, N5975, N168);
and AND2 (N5996, N5993, N1674);
nor NOR4 (N5997, N5969, N3003, N5410, N3084);
nor NOR3 (N5998, N5986, N3971, N2748);
or OR4 (N5999, N5995, N1839, N1060, N5648);
and AND3 (N6000, N5976, N4295, N5014);
or OR3 (N6001, N6000, N1758, N1360);
and AND4 (N6002, N5999, N5437, N3962, N2909);
or OR3 (N6003, N5980, N143, N5065);
nor NOR4 (N6004, N6002, N788, N2268, N3110);
nand NAND4 (N6005, N5997, N736, N5275, N582);
not NOT1 (N6006, N5998);
xor XOR2 (N6007, N6003, N606);
buf BUF1 (N6008, N5990);
and AND2 (N6009, N5994, N4383);
xor XOR2 (N6010, N6007, N1824);
xor XOR2 (N6011, N5989, N2451);
or OR2 (N6012, N6008, N4321);
or OR2 (N6013, N6001, N5045);
nor NOR4 (N6014, N6006, N5392, N1161, N4612);
xor XOR2 (N6015, N6014, N371);
or OR2 (N6016, N5991, N5400);
nand NAND4 (N6017, N6009, N742, N3225, N3370);
xor XOR2 (N6018, N6016, N4620);
nand NAND2 (N6019, N6012, N1967);
or OR2 (N6020, N5996, N4277);
buf BUF1 (N6021, N6005);
buf BUF1 (N6022, N6011);
nand NAND2 (N6023, N6015, N1671);
or OR4 (N6024, N6019, N2278, N4881, N3562);
not NOT1 (N6025, N6013);
xor XOR2 (N6026, N6020, N4606);
and AND2 (N6027, N6025, N177);
buf BUF1 (N6028, N6018);
and AND4 (N6029, N6026, N1669, N4906, N3562);
and AND2 (N6030, N6004, N1897);
and AND3 (N6031, N6029, N462, N4773);
xor XOR2 (N6032, N6031, N1796);
nor NOR4 (N6033, N6017, N5119, N4250, N5932);
xor XOR2 (N6034, N6027, N5707);
nor NOR3 (N6035, N6022, N5321, N4042);
nand NAND2 (N6036, N6028, N5971);
xor XOR2 (N6037, N6021, N1110);
buf BUF1 (N6038, N6035);
or OR2 (N6039, N6036, N1585);
xor XOR2 (N6040, N6037, N990);
not NOT1 (N6041, N6040);
nor NOR2 (N6042, N6041, N3969);
buf BUF1 (N6043, N6034);
xor XOR2 (N6044, N6042, N5156);
buf BUF1 (N6045, N6033);
buf BUF1 (N6046, N6032);
nand NAND2 (N6047, N6045, N548);
or OR3 (N6048, N6044, N5974, N4305);
and AND4 (N6049, N6010, N322, N4570, N2379);
xor XOR2 (N6050, N6038, N621);
or OR4 (N6051, N6023, N2252, N5055, N5507);
buf BUF1 (N6052, N6048);
buf BUF1 (N6053, N6050);
not NOT1 (N6054, N6046);
or OR2 (N6055, N6053, N1930);
nand NAND3 (N6056, N6047, N4821, N5941);
buf BUF1 (N6057, N6030);
nor NOR4 (N6058, N6055, N2382, N3026, N4849);
nor NOR2 (N6059, N6058, N1943);
xor XOR2 (N6060, N6057, N212);
buf BUF1 (N6061, N6060);
not NOT1 (N6062, N6024);
xor XOR2 (N6063, N6039, N5657);
nand NAND4 (N6064, N6062, N1821, N3464, N1013);
and AND2 (N6065, N6043, N1840);
buf BUF1 (N6066, N6059);
not NOT1 (N6067, N6065);
nor NOR4 (N6068, N6064, N1146, N3211, N1800);
xor XOR2 (N6069, N6068, N4318);
buf BUF1 (N6070, N6054);
nor NOR4 (N6071, N6063, N3337, N4245, N5930);
not NOT1 (N6072, N6061);
buf BUF1 (N6073, N6071);
or OR3 (N6074, N6073, N3665, N543);
nand NAND2 (N6075, N6051, N4654);
nor NOR3 (N6076, N6066, N3367, N4194);
nand NAND2 (N6077, N6075, N5272);
or OR2 (N6078, N6072, N136);
xor XOR2 (N6079, N6049, N4771);
and AND2 (N6080, N6070, N4388);
nor NOR3 (N6081, N6078, N4069, N1906);
or OR3 (N6082, N6052, N3713, N3939);
nor NOR2 (N6083, N6079, N2315);
or OR3 (N6084, N6074, N2038, N431);
nor NOR2 (N6085, N6083, N443);
xor XOR2 (N6086, N6056, N4724);
buf BUF1 (N6087, N6086);
or OR4 (N6088, N6085, N3284, N1776, N5516);
nor NOR2 (N6089, N6081, N170);
or OR4 (N6090, N6087, N2829, N1773, N4339);
not NOT1 (N6091, N6088);
buf BUF1 (N6092, N6090);
buf BUF1 (N6093, N6091);
or OR3 (N6094, N6093, N161, N150);
or OR4 (N6095, N6094, N4993, N3191, N230);
or OR3 (N6096, N6082, N647, N1265);
or OR2 (N6097, N6069, N4544);
and AND4 (N6098, N6080, N4104, N4369, N5309);
nand NAND2 (N6099, N6089, N1608);
nand NAND4 (N6100, N6084, N47, N4081, N5307);
and AND3 (N6101, N6100, N1692, N5155);
nand NAND2 (N6102, N6095, N3410);
nand NAND2 (N6103, N6097, N5884);
not NOT1 (N6104, N6076);
nand NAND2 (N6105, N6067, N1112);
nor NOR3 (N6106, N6077, N2432, N3548);
and AND3 (N6107, N6092, N3366, N5699);
xor XOR2 (N6108, N6106, N1868);
or OR4 (N6109, N6101, N4419, N1378, N3088);
buf BUF1 (N6110, N6102);
and AND2 (N6111, N6098, N1179);
or OR2 (N6112, N6111, N5898);
nand NAND3 (N6113, N6096, N2138, N5354);
nor NOR3 (N6114, N6103, N4657, N2019);
buf BUF1 (N6115, N6105);
not NOT1 (N6116, N6109);
nor NOR3 (N6117, N6112, N5940, N2537);
and AND3 (N6118, N6110, N2018, N5325);
or OR2 (N6119, N6107, N5033);
xor XOR2 (N6120, N6108, N5444);
or OR3 (N6121, N6104, N1587, N4747);
buf BUF1 (N6122, N6116);
and AND3 (N6123, N6099, N3458, N3226);
nand NAND3 (N6124, N6114, N4637, N5151);
buf BUF1 (N6125, N6113);
xor XOR2 (N6126, N6123, N560);
buf BUF1 (N6127, N6117);
buf BUF1 (N6128, N6124);
xor XOR2 (N6129, N6126, N21);
and AND3 (N6130, N6119, N4552, N4346);
buf BUF1 (N6131, N6127);
and AND3 (N6132, N6129, N3110, N2164);
or OR4 (N6133, N6131, N1150, N3235, N1922);
xor XOR2 (N6134, N6128, N2066);
xor XOR2 (N6135, N6125, N2906);
buf BUF1 (N6136, N6132);
not NOT1 (N6137, N6134);
or OR4 (N6138, N6120, N1718, N2189, N2919);
and AND3 (N6139, N6121, N5879, N3873);
buf BUF1 (N6140, N6138);
or OR3 (N6141, N6130, N21, N3703);
xor XOR2 (N6142, N6135, N3956);
nor NOR2 (N6143, N6142, N4103);
nor NOR3 (N6144, N6140, N1031, N3338);
nand NAND3 (N6145, N6143, N4614, N4605);
and AND2 (N6146, N6133, N5833);
and AND3 (N6147, N6145, N4631, N3263);
and AND3 (N6148, N6115, N2321, N3813);
and AND2 (N6149, N6122, N5096);
buf BUF1 (N6150, N6147);
xor XOR2 (N6151, N6137, N5873);
buf BUF1 (N6152, N6146);
or OR4 (N6153, N6152, N2259, N2114, N2215);
buf BUF1 (N6154, N6144);
or OR4 (N6155, N6154, N4440, N1881, N5373);
and AND4 (N6156, N6155, N5859, N2093, N4181);
and AND3 (N6157, N6136, N4984, N3059);
nor NOR2 (N6158, N6149, N1895);
and AND4 (N6159, N6150, N5526, N4081, N2681);
nor NOR4 (N6160, N6118, N5252, N4671, N2469);
nor NOR4 (N6161, N6141, N5265, N5251, N3038);
and AND2 (N6162, N6156, N910);
nor NOR3 (N6163, N6160, N2393, N3985);
not NOT1 (N6164, N6153);
xor XOR2 (N6165, N6148, N4189);
buf BUF1 (N6166, N6164);
xor XOR2 (N6167, N6157, N3167);
buf BUF1 (N6168, N6158);
and AND2 (N6169, N6162, N3650);
nor NOR2 (N6170, N6169, N3275);
not NOT1 (N6171, N6170);
and AND3 (N6172, N6167, N3556, N679);
buf BUF1 (N6173, N6161);
buf BUF1 (N6174, N6172);
buf BUF1 (N6175, N6174);
buf BUF1 (N6176, N6171);
not NOT1 (N6177, N6168);
not NOT1 (N6178, N6139);
or OR2 (N6179, N6159, N3349);
or OR4 (N6180, N6173, N1265, N202, N2154);
nand NAND4 (N6181, N6151, N569, N109, N2559);
not NOT1 (N6182, N6177);
not NOT1 (N6183, N6166);
nor NOR2 (N6184, N6181, N2984);
nor NOR2 (N6185, N6175, N2596);
nor NOR2 (N6186, N6180, N4024);
nand NAND3 (N6187, N6179, N1382, N3964);
buf BUF1 (N6188, N6186);
buf BUF1 (N6189, N6188);
not NOT1 (N6190, N6187);
nor NOR3 (N6191, N6189, N5113, N2495);
or OR2 (N6192, N6183, N2473);
nor NOR2 (N6193, N6192, N944);
xor XOR2 (N6194, N6191, N4090);
xor XOR2 (N6195, N6182, N2794);
or OR3 (N6196, N6165, N6100, N1287);
and AND2 (N6197, N6178, N887);
nand NAND2 (N6198, N6190, N2951);
and AND3 (N6199, N6176, N4349, N227);
or OR2 (N6200, N6185, N615);
and AND2 (N6201, N6193, N4446);
not NOT1 (N6202, N6163);
not NOT1 (N6203, N6197);
nand NAND2 (N6204, N6200, N4011);
nor NOR2 (N6205, N6203, N4479);
not NOT1 (N6206, N6199);
nand NAND3 (N6207, N6184, N5910, N3075);
nand NAND2 (N6208, N6205, N5646);
xor XOR2 (N6209, N6201, N830);
nand NAND3 (N6210, N6202, N2356, N2213);
nor NOR2 (N6211, N6210, N5515);
nand NAND3 (N6212, N6211, N5480, N4642);
nor NOR2 (N6213, N6196, N4050);
buf BUF1 (N6214, N6206);
xor XOR2 (N6215, N6194, N5098);
not NOT1 (N6216, N6204);
nor NOR4 (N6217, N6214, N3095, N6121, N2947);
xor XOR2 (N6218, N6208, N1446);
nor NOR4 (N6219, N6195, N1052, N5098, N5093);
buf BUF1 (N6220, N6217);
buf BUF1 (N6221, N6212);
not NOT1 (N6222, N6215);
nor NOR4 (N6223, N6198, N480, N3103, N5102);
xor XOR2 (N6224, N6207, N1848);
not NOT1 (N6225, N6209);
buf BUF1 (N6226, N6224);
or OR2 (N6227, N6221, N3971);
xor XOR2 (N6228, N6219, N1766);
nand NAND2 (N6229, N6222, N676);
not NOT1 (N6230, N6223);
or OR3 (N6231, N6229, N1284, N4525);
and AND2 (N6232, N6230, N1752);
xor XOR2 (N6233, N6225, N1291);
or OR2 (N6234, N6216, N335);
buf BUF1 (N6235, N6226);
buf BUF1 (N6236, N6227);
or OR2 (N6237, N6218, N5250);
nand NAND2 (N6238, N6236, N2684);
nor NOR3 (N6239, N6231, N541, N4909);
not NOT1 (N6240, N6220);
or OR2 (N6241, N6235, N973);
xor XOR2 (N6242, N6213, N4559);
xor XOR2 (N6243, N6237, N3097);
not NOT1 (N6244, N6228);
not NOT1 (N6245, N6243);
buf BUF1 (N6246, N6242);
not NOT1 (N6247, N6232);
nand NAND4 (N6248, N6246, N5284, N836, N4465);
nor NOR4 (N6249, N6233, N737, N1448, N4458);
or OR4 (N6250, N6241, N1578, N6241, N5774);
or OR3 (N6251, N6249, N3258, N330);
nand NAND4 (N6252, N6239, N5885, N324, N6110);
nor NOR2 (N6253, N6252, N4218);
or OR3 (N6254, N6251, N4416, N3480);
nor NOR3 (N6255, N6245, N4266, N1065);
nand NAND2 (N6256, N6254, N5341);
and AND2 (N6257, N6255, N3575);
not NOT1 (N6258, N6247);
nand NAND4 (N6259, N6258, N3169, N515, N4483);
xor XOR2 (N6260, N6253, N4427);
not NOT1 (N6261, N6259);
and AND3 (N6262, N6240, N5258, N928);
and AND3 (N6263, N6238, N3505, N3010);
and AND4 (N6264, N6248, N2038, N5564, N6202);
nand NAND3 (N6265, N6257, N1175, N4046);
and AND3 (N6266, N6250, N4451, N4586);
nor NOR4 (N6267, N6265, N745, N3890, N2766);
not NOT1 (N6268, N6244);
not NOT1 (N6269, N6262);
xor XOR2 (N6270, N6264, N3335);
buf BUF1 (N6271, N6234);
or OR2 (N6272, N6260, N4635);
buf BUF1 (N6273, N6268);
xor XOR2 (N6274, N6272, N3477);
or OR4 (N6275, N6266, N4109, N3288, N4152);
or OR4 (N6276, N6267, N5786, N1742, N1924);
xor XOR2 (N6277, N6271, N1081);
nor NOR2 (N6278, N6277, N6221);
nor NOR3 (N6279, N6275, N4908, N4874);
nor NOR2 (N6280, N6261, N1775);
nand NAND4 (N6281, N6279, N4194, N917, N3778);
and AND2 (N6282, N6269, N2394);
and AND2 (N6283, N6281, N1262);
nand NAND3 (N6284, N6273, N3076, N6158);
xor XOR2 (N6285, N6280, N3352);
or OR2 (N6286, N6285, N5362);
and AND2 (N6287, N6276, N5669);
nand NAND3 (N6288, N6287, N3770, N4005);
nand NAND3 (N6289, N6274, N3383, N6228);
and AND3 (N6290, N6263, N2655, N880);
nor NOR2 (N6291, N6286, N3869);
xor XOR2 (N6292, N6289, N6086);
and AND3 (N6293, N6282, N4433, N3627);
or OR2 (N6294, N6290, N5411);
nor NOR4 (N6295, N6291, N3011, N6111, N480);
xor XOR2 (N6296, N6256, N2061);
or OR2 (N6297, N6296, N880);
xor XOR2 (N6298, N6288, N2166);
nor NOR4 (N6299, N6292, N1750, N1760, N5809);
not NOT1 (N6300, N6294);
or OR2 (N6301, N6298, N2876);
and AND2 (N6302, N6300, N3776);
nor NOR3 (N6303, N6284, N5827, N4426);
or OR4 (N6304, N6278, N3957, N4409, N50);
not NOT1 (N6305, N6297);
nor NOR4 (N6306, N6270, N3849, N3469, N4496);
xor XOR2 (N6307, N6295, N2967);
and AND2 (N6308, N6283, N379);
buf BUF1 (N6309, N6301);
buf BUF1 (N6310, N6304);
or OR4 (N6311, N6305, N2791, N6264, N365);
buf BUF1 (N6312, N6310);
xor XOR2 (N6313, N6312, N1079);
nor NOR4 (N6314, N6311, N3219, N3642, N674);
nand NAND3 (N6315, N6302, N5545, N4112);
buf BUF1 (N6316, N6303);
buf BUF1 (N6317, N6314);
nand NAND2 (N6318, N6306, N815);
xor XOR2 (N6319, N6315, N3219);
or OR3 (N6320, N6308, N3416, N2882);
and AND3 (N6321, N6317, N3247, N1943);
or OR2 (N6322, N6313, N682);
xor XOR2 (N6323, N6293, N3527);
nor NOR3 (N6324, N6318, N3325, N5983);
or OR2 (N6325, N6319, N5593);
or OR3 (N6326, N6316, N1268, N380);
not NOT1 (N6327, N6307);
nand NAND2 (N6328, N6309, N5278);
xor XOR2 (N6329, N6322, N5874);
buf BUF1 (N6330, N6329);
not NOT1 (N6331, N6330);
nand NAND2 (N6332, N6331, N473);
nor NOR3 (N6333, N6324, N372, N235);
nand NAND2 (N6334, N6299, N4522);
not NOT1 (N6335, N6321);
nand NAND2 (N6336, N6326, N635);
xor XOR2 (N6337, N6323, N894);
buf BUF1 (N6338, N6333);
and AND4 (N6339, N6320, N5655, N4735, N3077);
not NOT1 (N6340, N6338);
or OR3 (N6341, N6336, N3356, N4403);
buf BUF1 (N6342, N6340);
or OR2 (N6343, N6335, N4909);
not NOT1 (N6344, N6328);
not NOT1 (N6345, N6344);
buf BUF1 (N6346, N6332);
or OR2 (N6347, N6345, N4039);
and AND3 (N6348, N6347, N1524, N3876);
nand NAND3 (N6349, N6327, N2760, N3794);
not NOT1 (N6350, N6334);
not NOT1 (N6351, N6339);
nor NOR4 (N6352, N6351, N6251, N1945, N2227);
not NOT1 (N6353, N6337);
not NOT1 (N6354, N6343);
xor XOR2 (N6355, N6348, N5215);
and AND4 (N6356, N6352, N4439, N2320, N1365);
xor XOR2 (N6357, N6325, N1271);
xor XOR2 (N6358, N6349, N2980);
and AND4 (N6359, N6357, N2824, N4144, N2285);
and AND3 (N6360, N6342, N1858, N6337);
and AND4 (N6361, N6354, N159, N2564, N297);
buf BUF1 (N6362, N6353);
xor XOR2 (N6363, N6355, N4930);
and AND2 (N6364, N6363, N1196);
or OR4 (N6365, N6364, N4737, N231, N6354);
not NOT1 (N6366, N6358);
and AND2 (N6367, N6361, N5854);
xor XOR2 (N6368, N6362, N4843);
xor XOR2 (N6369, N6368, N3339);
nor NOR4 (N6370, N6366, N2830, N6168, N4955);
or OR3 (N6371, N6346, N6054, N5576);
or OR3 (N6372, N6370, N276, N4982);
not NOT1 (N6373, N6356);
and AND4 (N6374, N6350, N6338, N3608, N909);
xor XOR2 (N6375, N6372, N2140);
buf BUF1 (N6376, N6359);
buf BUF1 (N6377, N6373);
nor NOR4 (N6378, N6374, N4370, N2066, N4810);
nor NOR3 (N6379, N6360, N6096, N5095);
xor XOR2 (N6380, N6379, N1262);
or OR2 (N6381, N6371, N2074);
nand NAND2 (N6382, N6365, N3548);
nor NOR2 (N6383, N6380, N6115);
nor NOR2 (N6384, N6369, N5750);
nor NOR4 (N6385, N6375, N947, N1783, N122);
nand NAND3 (N6386, N6341, N530, N3652);
buf BUF1 (N6387, N6377);
and AND2 (N6388, N6382, N3891);
not NOT1 (N6389, N6381);
nor NOR3 (N6390, N6367, N6241, N2539);
or OR3 (N6391, N6376, N1126, N6346);
xor XOR2 (N6392, N6385, N2166);
buf BUF1 (N6393, N6386);
nand NAND4 (N6394, N6383, N5680, N62, N208);
not NOT1 (N6395, N6393);
xor XOR2 (N6396, N6391, N1330);
buf BUF1 (N6397, N6390);
not NOT1 (N6398, N6384);
nor NOR4 (N6399, N6389, N4561, N5190, N417);
nand NAND3 (N6400, N6388, N5210, N4661);
nand NAND2 (N6401, N6397, N5561);
buf BUF1 (N6402, N6392);
nand NAND2 (N6403, N6402, N3622);
nand NAND4 (N6404, N6400, N1797, N2066, N562);
xor XOR2 (N6405, N6387, N4236);
nand NAND2 (N6406, N6399, N2305);
nor NOR3 (N6407, N6396, N140, N1949);
xor XOR2 (N6408, N6403, N500);
and AND3 (N6409, N6394, N3487, N3424);
nand NAND2 (N6410, N6408, N3016);
nor NOR4 (N6411, N6378, N3136, N6332, N4414);
not NOT1 (N6412, N6401);
xor XOR2 (N6413, N6405, N3996);
buf BUF1 (N6414, N6406);
or OR3 (N6415, N6411, N428, N5948);
not NOT1 (N6416, N6415);
and AND3 (N6417, N6412, N6019, N6268);
endmodule