// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N418,N416,N409,N378,N420,N419,N414,N415,N413,N421;

buf BUF1 (N22, N14);
nand NAND4 (N23, N4, N11, N12, N18);
nor NOR2 (N24, N6, N18);
or OR4 (N25, N12, N2, N16, N5);
not NOT1 (N26, N8);
nand NAND2 (N27, N14, N3);
not NOT1 (N28, N24);
and AND4 (N29, N3, N3, N26, N10);
xor XOR2 (N30, N6, N28);
or OR3 (N31, N5, N7, N10);
not NOT1 (N32, N28);
nor NOR4 (N33, N19, N11, N20, N26);
or OR2 (N34, N24, N4);
buf BUF1 (N35, N22);
nand NAND2 (N36, N31, N32);
or OR2 (N37, N30, N29);
buf BUF1 (N38, N22);
xor XOR2 (N39, N34, N9);
nor NOR4 (N40, N24, N38, N31, N16);
and AND2 (N41, N34, N17);
nand NAND3 (N42, N36, N29, N10);
nand NAND4 (N43, N33, N3, N3, N33);
nor NOR2 (N44, N23, N8);
nor NOR2 (N45, N43, N38);
nor NOR4 (N46, N37, N6, N1, N33);
and AND3 (N47, N35, N34, N13);
or OR2 (N48, N42, N32);
nand NAND4 (N49, N40, N36, N30, N32);
not NOT1 (N50, N39);
nor NOR4 (N51, N44, N13, N11, N3);
buf BUF1 (N52, N45);
and AND2 (N53, N27, N3);
buf BUF1 (N54, N48);
not NOT1 (N55, N52);
not NOT1 (N56, N55);
or OR3 (N57, N25, N2, N53);
not NOT1 (N58, N20);
xor XOR2 (N59, N46, N48);
or OR4 (N60, N57, N21, N43, N18);
nor NOR2 (N61, N49, N55);
not NOT1 (N62, N54);
nand NAND3 (N63, N58, N13, N10);
nor NOR4 (N64, N41, N53, N62, N38);
not NOT1 (N65, N42);
nor NOR2 (N66, N65, N43);
or OR4 (N67, N66, N62, N27, N64);
xor XOR2 (N68, N9, N33);
not NOT1 (N69, N47);
nand NAND2 (N70, N63, N31);
nand NAND4 (N71, N68, N10, N35, N61);
xor XOR2 (N72, N61, N38);
nor NOR4 (N73, N56, N36, N47, N57);
buf BUF1 (N74, N69);
buf BUF1 (N75, N74);
xor XOR2 (N76, N71, N46);
nor NOR2 (N77, N75, N47);
xor XOR2 (N78, N51, N59);
buf BUF1 (N79, N73);
nand NAND4 (N80, N47, N67, N30, N11);
buf BUF1 (N81, N62);
nand NAND2 (N82, N76, N79);
not NOT1 (N83, N60);
and AND4 (N84, N16, N26, N65, N23);
or OR4 (N85, N50, N64, N32, N29);
or OR2 (N86, N77, N50);
nand NAND3 (N87, N81, N75, N47);
nor NOR2 (N88, N83, N18);
and AND4 (N89, N78, N72, N57, N70);
or OR4 (N90, N1, N88, N54, N57);
nand NAND4 (N91, N8, N37, N58, N26);
not NOT1 (N92, N61);
not NOT1 (N93, N80);
and AND3 (N94, N86, N84, N89);
not NOT1 (N95, N1);
and AND4 (N96, N49, N39, N43, N68);
or OR4 (N97, N82, N69, N21, N24);
not NOT1 (N98, N97);
not NOT1 (N99, N96);
and AND3 (N100, N95, N66, N83);
and AND2 (N101, N85, N5);
nand NAND3 (N102, N99, N39, N84);
and AND2 (N103, N101, N62);
nor NOR4 (N104, N93, N91, N92, N22);
buf BUF1 (N105, N21);
nor NOR3 (N106, N66, N80, N85);
buf BUF1 (N107, N103);
nor NOR3 (N108, N107, N84, N33);
nor NOR4 (N109, N106, N29, N2, N33);
buf BUF1 (N110, N87);
xor XOR2 (N111, N94, N61);
nor NOR2 (N112, N102, N3);
and AND2 (N113, N112, N73);
xor XOR2 (N114, N105, N28);
nor NOR3 (N115, N109, N36, N52);
or OR2 (N116, N115, N70);
and AND4 (N117, N100, N113, N16, N48);
not NOT1 (N118, N103);
nand NAND3 (N119, N117, N61, N12);
nor NOR3 (N120, N116, N119, N24);
xor XOR2 (N121, N86, N21);
nor NOR3 (N122, N114, N14, N81);
not NOT1 (N123, N110);
nor NOR3 (N124, N108, N24, N54);
or OR3 (N125, N90, N58, N91);
not NOT1 (N126, N122);
or OR4 (N127, N111, N105, N95, N117);
nor NOR2 (N128, N121, N93);
or OR4 (N129, N104, N75, N26, N55);
not NOT1 (N130, N128);
nand NAND3 (N131, N98, N39, N109);
buf BUF1 (N132, N131);
nor NOR3 (N133, N124, N31, N27);
buf BUF1 (N134, N126);
buf BUF1 (N135, N133);
xor XOR2 (N136, N134, N100);
xor XOR2 (N137, N123, N126);
buf BUF1 (N138, N135);
or OR3 (N139, N125, N128, N29);
nor NOR3 (N140, N120, N43, N138);
nor NOR2 (N141, N23, N73);
nor NOR2 (N142, N132, N49);
xor XOR2 (N143, N118, N28);
nor NOR3 (N144, N137, N41, N110);
or OR3 (N145, N144, N31, N139);
nand NAND2 (N146, N56, N121);
and AND3 (N147, N145, N38, N19);
nor NOR3 (N148, N146, N131, N62);
nor NOR4 (N149, N142, N89, N133, N37);
nand NAND2 (N150, N148, N95);
buf BUF1 (N151, N143);
or OR3 (N152, N130, N31, N45);
nor NOR4 (N153, N149, N94, N113, N114);
nand NAND3 (N154, N153, N96, N59);
and AND4 (N155, N151, N50, N40, N6);
buf BUF1 (N156, N152);
not NOT1 (N157, N150);
buf BUF1 (N158, N155);
nor NOR2 (N159, N157, N24);
or OR4 (N160, N127, N26, N11, N101);
or OR4 (N161, N136, N66, N143, N94);
buf BUF1 (N162, N160);
xor XOR2 (N163, N162, N156);
nand NAND2 (N164, N37, N108);
not NOT1 (N165, N147);
nand NAND3 (N166, N129, N164, N165);
not NOT1 (N167, N59);
nand NAND3 (N168, N76, N125, N57);
or OR4 (N169, N166, N10, N142, N28);
xor XOR2 (N170, N168, N10);
nor NOR3 (N171, N154, N140, N127);
and AND3 (N172, N134, N133, N56);
and AND4 (N173, N158, N83, N12, N163);
and AND4 (N174, N126, N63, N69, N62);
buf BUF1 (N175, N173);
or OR2 (N176, N169, N56);
nor NOR4 (N177, N141, N109, N99, N70);
not NOT1 (N178, N159);
not NOT1 (N179, N174);
nor NOR4 (N180, N161, N75, N63, N105);
nor NOR3 (N181, N167, N62, N110);
nor NOR3 (N182, N170, N137, N153);
nand NAND3 (N183, N181, N83, N60);
not NOT1 (N184, N183);
nand NAND4 (N185, N180, N64, N170, N37);
and AND4 (N186, N178, N139, N160, N81);
xor XOR2 (N187, N186, N79);
nand NAND2 (N188, N187, N124);
nand NAND3 (N189, N175, N80, N33);
xor XOR2 (N190, N185, N175);
or OR2 (N191, N176, N143);
nand NAND2 (N192, N171, N20);
nand NAND3 (N193, N189, N29, N144);
or OR4 (N194, N188, N97, N31, N113);
xor XOR2 (N195, N192, N23);
not NOT1 (N196, N193);
nor NOR3 (N197, N195, N155, N75);
or OR3 (N198, N196, N75, N105);
nand NAND4 (N199, N184, N97, N181, N133);
nor NOR4 (N200, N199, N164, N139, N181);
xor XOR2 (N201, N200, N56);
and AND3 (N202, N201, N27, N117);
not NOT1 (N203, N191);
or OR3 (N204, N203, N117, N52);
and AND2 (N205, N204, N41);
buf BUF1 (N206, N202);
xor XOR2 (N207, N179, N37);
nor NOR2 (N208, N206, N173);
and AND4 (N209, N208, N123, N29, N119);
nor NOR2 (N210, N209, N129);
or OR3 (N211, N210, N56, N67);
nand NAND4 (N212, N211, N83, N105, N69);
and AND2 (N213, N172, N112);
not NOT1 (N214, N212);
xor XOR2 (N215, N213, N123);
xor XOR2 (N216, N215, N169);
nor NOR3 (N217, N197, N92, N190);
nand NAND2 (N218, N18, N142);
nor NOR4 (N219, N194, N67, N79, N179);
or OR2 (N220, N216, N105);
and AND3 (N221, N218, N10, N52);
not NOT1 (N222, N182);
not NOT1 (N223, N217);
and AND3 (N224, N205, N93, N15);
nor NOR3 (N225, N224, N120, N204);
or OR3 (N226, N221, N73, N215);
or OR2 (N227, N207, N49);
and AND3 (N228, N198, N183, N76);
nor NOR3 (N229, N177, N180, N161);
nand NAND2 (N230, N219, N6);
and AND4 (N231, N223, N73, N145, N100);
buf BUF1 (N232, N227);
nand NAND3 (N233, N232, N81, N72);
and AND3 (N234, N231, N9, N25);
xor XOR2 (N235, N228, N61);
and AND2 (N236, N230, N197);
nand NAND2 (N237, N214, N142);
nand NAND2 (N238, N229, N35);
not NOT1 (N239, N226);
xor XOR2 (N240, N225, N156);
and AND2 (N241, N220, N232);
and AND3 (N242, N235, N134, N135);
buf BUF1 (N243, N240);
and AND2 (N244, N239, N163);
xor XOR2 (N245, N244, N224);
or OR3 (N246, N234, N187, N52);
nand NAND2 (N247, N233, N125);
buf BUF1 (N248, N236);
buf BUF1 (N249, N242);
nor NOR3 (N250, N249, N115, N223);
nand NAND2 (N251, N246, N2);
or OR4 (N252, N222, N102, N154, N223);
nand NAND3 (N253, N243, N34, N146);
not NOT1 (N254, N252);
xor XOR2 (N255, N247, N1);
not NOT1 (N256, N238);
not NOT1 (N257, N254);
nor NOR2 (N258, N253, N4);
xor XOR2 (N259, N248, N12);
or OR4 (N260, N251, N13, N78, N13);
or OR3 (N261, N250, N193, N56);
xor XOR2 (N262, N245, N141);
nor NOR3 (N263, N237, N132, N149);
and AND2 (N264, N257, N225);
nor NOR4 (N265, N263, N109, N263, N236);
buf BUF1 (N266, N259);
nor NOR2 (N267, N241, N213);
nand NAND3 (N268, N255, N172, N114);
nand NAND4 (N269, N261, N230, N61, N61);
nand NAND2 (N270, N258, N25);
not NOT1 (N271, N262);
nand NAND2 (N272, N268, N185);
and AND4 (N273, N266, N116, N202, N167);
buf BUF1 (N274, N265);
xor XOR2 (N275, N273, N53);
buf BUF1 (N276, N269);
nand NAND4 (N277, N264, N270, N160, N123);
buf BUF1 (N278, N8);
nor NOR2 (N279, N256, N248);
not NOT1 (N280, N260);
nor NOR3 (N281, N279, N156, N109);
nor NOR2 (N282, N277, N141);
xor XOR2 (N283, N281, N197);
and AND4 (N284, N282, N142, N92, N242);
not NOT1 (N285, N283);
and AND4 (N286, N280, N122, N44, N44);
or OR4 (N287, N285, N226, N62, N201);
nor NOR4 (N288, N276, N238, N17, N200);
and AND4 (N289, N278, N105, N147, N263);
not NOT1 (N290, N267);
xor XOR2 (N291, N272, N31);
not NOT1 (N292, N286);
buf BUF1 (N293, N274);
not NOT1 (N294, N288);
not NOT1 (N295, N275);
or OR2 (N296, N293, N252);
or OR4 (N297, N289, N200, N88, N2);
nand NAND4 (N298, N271, N158, N234, N136);
and AND3 (N299, N294, N100, N18);
xor XOR2 (N300, N284, N71);
xor XOR2 (N301, N300, N172);
or OR2 (N302, N287, N60);
not NOT1 (N303, N296);
buf BUF1 (N304, N299);
and AND3 (N305, N297, N74, N245);
xor XOR2 (N306, N290, N213);
nand NAND3 (N307, N305, N138, N263);
xor XOR2 (N308, N303, N50);
xor XOR2 (N309, N298, N26);
nand NAND3 (N310, N302, N300, N130);
buf BUF1 (N311, N308);
xor XOR2 (N312, N292, N7);
nor NOR3 (N313, N311, N300, N275);
not NOT1 (N314, N306);
and AND2 (N315, N304, N82);
not NOT1 (N316, N309);
or OR2 (N317, N307, N161);
nor NOR3 (N318, N312, N156, N52);
and AND2 (N319, N291, N316);
nand NAND3 (N320, N140, N225, N16);
not NOT1 (N321, N313);
nor NOR3 (N322, N295, N4, N11);
and AND4 (N323, N318, N213, N25, N207);
or OR2 (N324, N315, N168);
or OR2 (N325, N317, N250);
nand NAND2 (N326, N319, N266);
nor NOR2 (N327, N326, N244);
nand NAND4 (N328, N321, N191, N40, N106);
xor XOR2 (N329, N328, N108);
not NOT1 (N330, N323);
buf BUF1 (N331, N329);
or OR2 (N332, N322, N304);
nor NOR3 (N333, N314, N54, N268);
not NOT1 (N334, N333);
or OR4 (N335, N330, N94, N136, N49);
buf BUF1 (N336, N324);
nor NOR2 (N337, N320, N261);
xor XOR2 (N338, N337, N173);
xor XOR2 (N339, N334, N245);
and AND3 (N340, N325, N231, N137);
or OR2 (N341, N335, N30);
nand NAND4 (N342, N338, N148, N124, N290);
not NOT1 (N343, N340);
xor XOR2 (N344, N327, N201);
buf BUF1 (N345, N331);
nand NAND2 (N346, N332, N98);
nand NAND2 (N347, N346, N335);
xor XOR2 (N348, N345, N176);
nand NAND3 (N349, N343, N133, N313);
nand NAND3 (N350, N310, N216, N103);
or OR2 (N351, N341, N96);
nor NOR4 (N352, N348, N35, N146, N301);
nor NOR3 (N353, N30, N86, N327);
nor NOR2 (N354, N350, N139);
nand NAND4 (N355, N347, N309, N59, N271);
or OR4 (N356, N352, N41, N293, N78);
xor XOR2 (N357, N336, N302);
xor XOR2 (N358, N351, N171);
nor NOR2 (N359, N354, N354);
buf BUF1 (N360, N339);
or OR3 (N361, N349, N44, N173);
buf BUF1 (N362, N344);
not NOT1 (N363, N355);
buf BUF1 (N364, N361);
buf BUF1 (N365, N358);
or OR4 (N366, N364, N331, N204, N232);
buf BUF1 (N367, N362);
or OR4 (N368, N342, N236, N93, N184);
nand NAND2 (N369, N356, N338);
not NOT1 (N370, N369);
not NOT1 (N371, N363);
nor NOR3 (N372, N370, N302, N232);
and AND4 (N373, N371, N194, N341, N122);
xor XOR2 (N374, N365, N173);
buf BUF1 (N375, N368);
nor NOR2 (N376, N353, N160);
nor NOR3 (N377, N357, N78, N100);
buf BUF1 (N378, N366);
xor XOR2 (N379, N374, N322);
not NOT1 (N380, N379);
buf BUF1 (N381, N367);
nor NOR2 (N382, N381, N343);
not NOT1 (N383, N380);
and AND3 (N384, N372, N348, N258);
nor NOR4 (N385, N376, N306, N212, N261);
xor XOR2 (N386, N375, N128);
buf BUF1 (N387, N383);
xor XOR2 (N388, N359, N382);
not NOT1 (N389, N272);
or OR3 (N390, N360, N7, N371);
not NOT1 (N391, N377);
nor NOR4 (N392, N384, N233, N152, N136);
and AND3 (N393, N389, N304, N339);
nor NOR4 (N394, N390, N309, N379, N145);
xor XOR2 (N395, N386, N150);
nor NOR4 (N396, N393, N233, N19, N205);
nor NOR3 (N397, N391, N162, N199);
buf BUF1 (N398, N392);
nor NOR4 (N399, N385, N333, N251, N185);
buf BUF1 (N400, N388);
nand NAND4 (N401, N387, N212, N14, N375);
or OR2 (N402, N400, N372);
nand NAND2 (N403, N399, N373);
and AND3 (N404, N396, N355, N269);
or OR4 (N405, N11, N65, N280, N221);
not NOT1 (N406, N402);
buf BUF1 (N407, N395);
and AND4 (N408, N406, N256, N184, N405);
nand NAND3 (N409, N242, N333, N118);
buf BUF1 (N410, N408);
buf BUF1 (N411, N407);
or OR4 (N412, N394, N354, N381, N172);
buf BUF1 (N413, N397);
xor XOR2 (N414, N404, N339);
not NOT1 (N415, N403);
not NOT1 (N416, N412);
nand NAND3 (N417, N411, N402, N373);
and AND2 (N418, N410, N359);
or OR2 (N419, N417, N158);
or OR2 (N420, N401, N174);
xor XOR2 (N421, N398, N81);
endmodule