// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N1505,N1506,N1498,N1510,N1508,N1499,N1511,N1513,N1503,N1514;

nand NAND3 (N15, N2, N9, N11);
and AND2 (N16, N7, N10);
and AND3 (N17, N12, N12, N2);
and AND2 (N18, N4, N8);
buf BUF1 (N19, N10);
or OR3 (N20, N2, N9, N3);
and AND2 (N21, N9, N13);
buf BUF1 (N22, N4);
nor NOR2 (N23, N15, N14);
nand NAND2 (N24, N16, N5);
nor NOR2 (N25, N19, N4);
or OR3 (N26, N1, N17, N17);
not NOT1 (N27, N25);
nand NAND3 (N28, N10, N15, N5);
or OR3 (N29, N27, N28, N9);
or OR3 (N30, N27, N20, N17);
not NOT1 (N31, N4);
nand NAND4 (N32, N7, N26, N26, N14);
nand NAND2 (N33, N10, N1);
buf BUF1 (N34, N32);
nand NAND3 (N35, N23, N30, N6);
nor NOR4 (N36, N29, N21, N31, N24);
buf BUF1 (N37, N1);
nand NAND3 (N38, N13, N32, N29);
buf BUF1 (N39, N19);
not NOT1 (N40, N36);
nor NOR2 (N41, N19, N18);
buf BUF1 (N42, N14);
nand NAND2 (N43, N34, N40);
or OR4 (N44, N25, N18, N43, N40);
xor XOR2 (N45, N44, N9);
or OR4 (N46, N21, N27, N36, N45);
or OR4 (N47, N19, N46, N32, N1);
and AND2 (N48, N6, N26);
or OR2 (N49, N47, N43);
not NOT1 (N50, N33);
or OR2 (N51, N38, N16);
xor XOR2 (N52, N41, N25);
nor NOR2 (N53, N51, N28);
nor NOR2 (N54, N50, N21);
xor XOR2 (N55, N35, N24);
nor NOR2 (N56, N55, N30);
and AND3 (N57, N52, N32, N35);
nand NAND3 (N58, N42, N3, N44);
nand NAND2 (N59, N56, N28);
nand NAND2 (N60, N58, N49);
nand NAND3 (N61, N58, N26, N21);
not NOT1 (N62, N57);
nand NAND3 (N63, N39, N51, N16);
xor XOR2 (N64, N60, N8);
xor XOR2 (N65, N61, N6);
nor NOR2 (N66, N59, N11);
buf BUF1 (N67, N65);
or OR2 (N68, N64, N13);
and AND4 (N69, N37, N2, N25, N30);
nor NOR3 (N70, N48, N24, N34);
xor XOR2 (N71, N53, N8);
not NOT1 (N72, N63);
or OR2 (N73, N68, N72);
or OR4 (N74, N11, N16, N63, N23);
nor NOR2 (N75, N62, N38);
nand NAND2 (N76, N73, N45);
not NOT1 (N77, N69);
nand NAND4 (N78, N77, N54, N26, N20);
nand NAND2 (N79, N64, N18);
or OR2 (N80, N70, N51);
and AND2 (N81, N76, N3);
buf BUF1 (N82, N67);
nor NOR2 (N83, N66, N75);
nor NOR3 (N84, N11, N41, N80);
xor XOR2 (N85, N1, N29);
nor NOR3 (N86, N83, N61, N68);
nor NOR2 (N87, N85, N81);
or OR3 (N88, N11, N2, N79);
not NOT1 (N89, N46);
nor NOR4 (N90, N89, N48, N66, N46);
buf BUF1 (N91, N22);
or OR4 (N92, N88, N33, N78, N85);
not NOT1 (N93, N85);
nand NAND2 (N94, N87, N13);
and AND4 (N95, N93, N49, N5, N15);
or OR4 (N96, N71, N4, N89, N92);
or OR4 (N97, N24, N89, N38, N41);
or OR3 (N98, N96, N42, N14);
or OR3 (N99, N86, N74, N25);
nand NAND3 (N100, N61, N12, N73);
nand NAND2 (N101, N95, N99);
or OR2 (N102, N89, N101);
nand NAND3 (N103, N55, N60, N80);
not NOT1 (N104, N90);
not NOT1 (N105, N82);
or OR3 (N106, N105, N43, N40);
nand NAND3 (N107, N91, N65, N81);
nand NAND4 (N108, N103, N67, N105, N42);
nand NAND2 (N109, N104, N49);
nor NOR4 (N110, N109, N86, N77, N11);
buf BUF1 (N111, N84);
and AND4 (N112, N97, N23, N92, N18);
nor NOR3 (N113, N94, N19, N11);
not NOT1 (N114, N112);
nand NAND2 (N115, N107, N50);
not NOT1 (N116, N114);
not NOT1 (N117, N111);
xor XOR2 (N118, N116, N98);
nor NOR4 (N119, N74, N94, N38, N15);
nor NOR3 (N120, N106, N61, N85);
buf BUF1 (N121, N102);
nor NOR2 (N122, N117, N81);
and AND3 (N123, N115, N100, N117);
buf BUF1 (N124, N47);
buf BUF1 (N125, N121);
nand NAND3 (N126, N120, N81, N118);
and AND4 (N127, N73, N35, N55, N5);
buf BUF1 (N128, N125);
nand NAND2 (N129, N126, N90);
and AND3 (N130, N119, N79, N123);
buf BUF1 (N131, N22);
xor XOR2 (N132, N131, N36);
not NOT1 (N133, N128);
buf BUF1 (N134, N133);
xor XOR2 (N135, N129, N37);
xor XOR2 (N136, N134, N50);
nand NAND2 (N137, N113, N120);
not NOT1 (N138, N130);
nor NOR4 (N139, N135, N11, N10, N81);
buf BUF1 (N140, N137);
xor XOR2 (N141, N140, N37);
xor XOR2 (N142, N122, N45);
buf BUF1 (N143, N142);
and AND3 (N144, N141, N124, N37);
or OR3 (N145, N48, N95, N30);
not NOT1 (N146, N144);
xor XOR2 (N147, N110, N54);
xor XOR2 (N148, N139, N56);
buf BUF1 (N149, N132);
nand NAND3 (N150, N108, N75, N53);
buf BUF1 (N151, N127);
nor NOR2 (N152, N146, N135);
or OR2 (N153, N145, N51);
buf BUF1 (N154, N143);
xor XOR2 (N155, N150, N82);
xor XOR2 (N156, N151, N127);
or OR4 (N157, N149, N114, N122, N36);
buf BUF1 (N158, N157);
buf BUF1 (N159, N155);
buf BUF1 (N160, N156);
buf BUF1 (N161, N147);
or OR2 (N162, N152, N64);
xor XOR2 (N163, N158, N84);
and AND4 (N164, N138, N31, N120, N149);
not NOT1 (N165, N136);
nor NOR2 (N166, N153, N128);
xor XOR2 (N167, N161, N90);
or OR4 (N168, N159, N16, N71, N89);
nor NOR4 (N169, N163, N65, N48, N163);
and AND2 (N170, N166, N72);
nor NOR3 (N171, N169, N158, N121);
and AND3 (N172, N167, N33, N82);
xor XOR2 (N173, N171, N105);
nor NOR4 (N174, N173, N52, N166, N31);
buf BUF1 (N175, N148);
nand NAND3 (N176, N164, N48, N38);
buf BUF1 (N177, N154);
nor NOR3 (N178, N174, N54, N78);
and AND2 (N179, N160, N18);
xor XOR2 (N180, N170, N44);
nor NOR3 (N181, N165, N38, N7);
or OR4 (N182, N175, N52, N101, N116);
nor NOR3 (N183, N180, N33, N45);
xor XOR2 (N184, N172, N64);
buf BUF1 (N185, N181);
buf BUF1 (N186, N162);
nand NAND3 (N187, N183, N105, N81);
buf BUF1 (N188, N179);
nor NOR4 (N189, N182, N160, N182, N13);
and AND2 (N190, N186, N183);
buf BUF1 (N191, N189);
nor NOR2 (N192, N184, N41);
not NOT1 (N193, N176);
not NOT1 (N194, N185);
xor XOR2 (N195, N192, N154);
not NOT1 (N196, N177);
not NOT1 (N197, N191);
xor XOR2 (N198, N197, N57);
nand NAND3 (N199, N178, N125, N42);
xor XOR2 (N200, N188, N119);
and AND3 (N201, N193, N163, N196);
nor NOR2 (N202, N144, N91);
xor XOR2 (N203, N199, N166);
buf BUF1 (N204, N201);
nor NOR3 (N205, N198, N31, N181);
not NOT1 (N206, N205);
or OR2 (N207, N206, N92);
and AND3 (N208, N200, N110, N46);
buf BUF1 (N209, N203);
or OR2 (N210, N209, N95);
or OR2 (N211, N204, N70);
and AND4 (N212, N202, N109, N159, N55);
or OR3 (N213, N190, N73, N39);
nor NOR3 (N214, N187, N76, N195);
buf BUF1 (N215, N42);
nor NOR2 (N216, N211, N114);
xor XOR2 (N217, N213, N89);
not NOT1 (N218, N212);
or OR2 (N219, N214, N178);
and AND4 (N220, N218, N50, N29, N106);
or OR2 (N221, N219, N164);
not NOT1 (N222, N194);
buf BUF1 (N223, N208);
nand NAND4 (N224, N215, N50, N212, N145);
and AND3 (N225, N224, N97, N114);
nor NOR3 (N226, N216, N91, N67);
not NOT1 (N227, N222);
not NOT1 (N228, N221);
nand NAND4 (N229, N227, N126, N34, N51);
nand NAND3 (N230, N207, N49, N14);
and AND2 (N231, N230, N5);
nand NAND3 (N232, N223, N157, N72);
xor XOR2 (N233, N231, N148);
xor XOR2 (N234, N220, N41);
nand NAND4 (N235, N210, N174, N178, N115);
or OR2 (N236, N229, N16);
buf BUF1 (N237, N225);
not NOT1 (N238, N233);
nor NOR3 (N239, N226, N8, N16);
buf BUF1 (N240, N232);
xor XOR2 (N241, N228, N228);
nor NOR4 (N242, N237, N81, N240, N70);
and AND3 (N243, N146, N119, N16);
nor NOR2 (N244, N239, N177);
not NOT1 (N245, N235);
not NOT1 (N246, N244);
buf BUF1 (N247, N217);
and AND3 (N248, N246, N29, N226);
or OR2 (N249, N234, N39);
buf BUF1 (N250, N249);
and AND4 (N251, N242, N63, N97, N109);
nor NOR3 (N252, N243, N164, N187);
buf BUF1 (N253, N238);
or OR4 (N254, N252, N34, N142, N239);
nor NOR4 (N255, N253, N101, N146, N234);
nor NOR2 (N256, N248, N31);
nor NOR4 (N257, N236, N133, N138, N102);
xor XOR2 (N258, N168, N131);
not NOT1 (N259, N250);
or OR4 (N260, N259, N3, N183, N169);
nand NAND2 (N261, N257, N150);
or OR4 (N262, N256, N30, N228, N261);
not NOT1 (N263, N17);
buf BUF1 (N264, N254);
nor NOR4 (N265, N251, N228, N95, N219);
not NOT1 (N266, N245);
buf BUF1 (N267, N266);
xor XOR2 (N268, N267, N60);
not NOT1 (N269, N264);
not NOT1 (N270, N262);
and AND4 (N271, N265, N211, N184, N240);
buf BUF1 (N272, N263);
buf BUF1 (N273, N260);
or OR4 (N274, N241, N83, N262, N243);
buf BUF1 (N275, N268);
or OR4 (N276, N275, N217, N263, N200);
and AND3 (N277, N274, N53, N212);
not NOT1 (N278, N277);
nand NAND3 (N279, N278, N77, N270);
buf BUF1 (N280, N106);
buf BUF1 (N281, N255);
xor XOR2 (N282, N271, N54);
nor NOR3 (N283, N247, N257, N218);
or OR2 (N284, N279, N231);
buf BUF1 (N285, N272);
and AND4 (N286, N284, N7, N34, N270);
buf BUF1 (N287, N273);
buf BUF1 (N288, N281);
not NOT1 (N289, N288);
nor NOR4 (N290, N289, N113, N83, N66);
nand NAND2 (N291, N258, N67);
and AND4 (N292, N285, N147, N180, N162);
and AND4 (N293, N291, N62, N126, N104);
nor NOR3 (N294, N276, N270, N88);
not NOT1 (N295, N286);
nor NOR3 (N296, N293, N228, N245);
xor XOR2 (N297, N294, N103);
buf BUF1 (N298, N283);
nor NOR4 (N299, N295, N195, N50, N186);
not NOT1 (N300, N287);
nor NOR3 (N301, N299, N58, N156);
nor NOR3 (N302, N301, N163, N169);
nor NOR4 (N303, N290, N145, N75, N260);
nand NAND4 (N304, N303, N38, N137, N86);
not NOT1 (N305, N302);
and AND4 (N306, N305, N297, N51, N129);
buf BUF1 (N307, N34);
buf BUF1 (N308, N298);
or OR2 (N309, N292, N103);
or OR2 (N310, N269, N225);
buf BUF1 (N311, N282);
nor NOR4 (N312, N311, N239, N2, N266);
or OR3 (N313, N312, N202, N40);
buf BUF1 (N314, N280);
buf BUF1 (N315, N314);
buf BUF1 (N316, N313);
buf BUF1 (N317, N315);
and AND4 (N318, N306, N316, N81, N173);
not NOT1 (N319, N65);
nor NOR4 (N320, N308, N10, N75, N27);
not NOT1 (N321, N300);
nor NOR2 (N322, N320, N240);
buf BUF1 (N323, N321);
and AND4 (N324, N307, N240, N115, N240);
nor NOR4 (N325, N319, N236, N104, N223);
nor NOR4 (N326, N318, N242, N318, N157);
or OR3 (N327, N310, N74, N317);
xor XOR2 (N328, N167, N220);
nor NOR3 (N329, N324, N235, N127);
nor NOR4 (N330, N328, N165, N206, N68);
and AND4 (N331, N296, N56, N204, N116);
xor XOR2 (N332, N327, N240);
nand NAND4 (N333, N331, N155, N234, N58);
nand NAND2 (N334, N304, N233);
nand NAND2 (N335, N334, N10);
or OR4 (N336, N326, N265, N324, N47);
xor XOR2 (N337, N335, N251);
nor NOR3 (N338, N323, N54, N174);
xor XOR2 (N339, N325, N231);
and AND3 (N340, N336, N322, N198);
not NOT1 (N341, N293);
or OR3 (N342, N309, N69, N244);
and AND3 (N343, N339, N58, N135);
buf BUF1 (N344, N337);
not NOT1 (N345, N333);
not NOT1 (N346, N345);
nor NOR3 (N347, N329, N159, N131);
nor NOR2 (N348, N347, N226);
not NOT1 (N349, N330);
nand NAND3 (N350, N343, N334, N203);
nor NOR4 (N351, N349, N170, N233, N67);
not NOT1 (N352, N351);
xor XOR2 (N353, N341, N96);
buf BUF1 (N354, N340);
nor NOR2 (N355, N354, N321);
nor NOR2 (N356, N332, N130);
or OR2 (N357, N350, N206);
not NOT1 (N358, N346);
not NOT1 (N359, N358);
not NOT1 (N360, N353);
and AND2 (N361, N360, N56);
nor NOR4 (N362, N352, N251, N256, N271);
nor NOR4 (N363, N359, N213, N252, N334);
and AND3 (N364, N344, N270, N350);
and AND4 (N365, N357, N185, N30, N254);
nor NOR2 (N366, N361, N124);
not NOT1 (N367, N366);
nand NAND2 (N368, N356, N158);
nor NOR3 (N369, N368, N122, N256);
nand NAND2 (N370, N348, N91);
xor XOR2 (N371, N342, N168);
buf BUF1 (N372, N367);
and AND4 (N373, N370, N186, N357, N194);
nor NOR3 (N374, N362, N2, N138);
or OR2 (N375, N364, N123);
nor NOR3 (N376, N338, N183, N329);
nand NAND4 (N377, N376, N370, N305, N166);
and AND3 (N378, N371, N250, N174);
or OR2 (N379, N373, N192);
or OR4 (N380, N379, N170, N267, N124);
or OR2 (N381, N363, N14);
xor XOR2 (N382, N369, N175);
nor NOR4 (N383, N378, N197, N307, N160);
or OR4 (N384, N382, N319, N23, N144);
or OR3 (N385, N374, N322, N224);
or OR3 (N386, N372, N330, N47);
nor NOR3 (N387, N386, N374, N223);
or OR3 (N388, N355, N310, N323);
nor NOR2 (N389, N388, N236);
or OR2 (N390, N365, N23);
nand NAND2 (N391, N390, N37);
and AND3 (N392, N385, N45, N1);
nand NAND4 (N393, N381, N51, N345, N248);
xor XOR2 (N394, N392, N342);
buf BUF1 (N395, N375);
not NOT1 (N396, N395);
xor XOR2 (N397, N389, N46);
nand NAND2 (N398, N384, N162);
nor NOR2 (N399, N391, N360);
nand NAND3 (N400, N383, N120, N192);
xor XOR2 (N401, N377, N12);
buf BUF1 (N402, N393);
buf BUF1 (N403, N402);
nand NAND2 (N404, N401, N107);
and AND2 (N405, N403, N324);
nor NOR2 (N406, N394, N46);
nand NAND4 (N407, N406, N146, N270, N13);
buf BUF1 (N408, N398);
and AND2 (N409, N404, N29);
xor XOR2 (N410, N387, N175);
nor NOR2 (N411, N405, N105);
buf BUF1 (N412, N411);
or OR4 (N413, N407, N81, N205, N405);
xor XOR2 (N414, N397, N168);
nor NOR2 (N415, N396, N329);
xor XOR2 (N416, N409, N294);
xor XOR2 (N417, N400, N186);
buf BUF1 (N418, N380);
nand NAND2 (N419, N415, N266);
nor NOR4 (N420, N399, N309, N411, N57);
and AND3 (N421, N408, N161, N51);
and AND2 (N422, N412, N291);
and AND3 (N423, N410, N381, N54);
or OR2 (N424, N419, N214);
xor XOR2 (N425, N421, N337);
nand NAND4 (N426, N413, N1, N61, N218);
not NOT1 (N427, N414);
or OR2 (N428, N422, N85);
nand NAND2 (N429, N420, N242);
nor NOR2 (N430, N428, N114);
nand NAND2 (N431, N423, N281);
xor XOR2 (N432, N427, N381);
nand NAND4 (N433, N416, N347, N193, N77);
xor XOR2 (N434, N425, N142);
buf BUF1 (N435, N433);
xor XOR2 (N436, N424, N28);
or OR2 (N437, N436, N263);
nand NAND3 (N438, N426, N306, N220);
or OR3 (N439, N435, N371, N134);
and AND4 (N440, N437, N262, N177, N307);
buf BUF1 (N441, N417);
not NOT1 (N442, N430);
buf BUF1 (N443, N431);
buf BUF1 (N444, N434);
xor XOR2 (N445, N444, N58);
xor XOR2 (N446, N445, N154);
and AND4 (N447, N438, N182, N414, N240);
or OR3 (N448, N429, N53, N197);
not NOT1 (N449, N439);
or OR4 (N450, N440, N430, N230, N116);
and AND3 (N451, N442, N149, N392);
buf BUF1 (N452, N450);
not NOT1 (N453, N447);
or OR3 (N454, N443, N294, N345);
xor XOR2 (N455, N449, N206);
and AND4 (N456, N441, N446, N9, N349);
or OR4 (N457, N347, N234, N363, N193);
not NOT1 (N458, N452);
buf BUF1 (N459, N432);
and AND4 (N460, N418, N336, N128, N179);
and AND3 (N461, N455, N141, N329);
not NOT1 (N462, N456);
buf BUF1 (N463, N461);
not NOT1 (N464, N463);
or OR4 (N465, N451, N132, N443, N423);
nor NOR4 (N466, N459, N50, N44, N250);
or OR4 (N467, N460, N222, N404, N22);
and AND2 (N468, N448, N315);
and AND4 (N469, N457, N246, N158, N72);
and AND3 (N470, N468, N202, N414);
nor NOR2 (N471, N453, N411);
nand NAND3 (N472, N471, N246, N412);
xor XOR2 (N473, N454, N386);
nor NOR2 (N474, N469, N366);
nand NAND3 (N475, N473, N178, N382);
or OR2 (N476, N464, N139);
and AND3 (N477, N476, N461, N330);
nand NAND4 (N478, N474, N143, N121, N216);
buf BUF1 (N479, N465);
buf BUF1 (N480, N466);
buf BUF1 (N481, N458);
or OR4 (N482, N479, N453, N209, N116);
not NOT1 (N483, N472);
buf BUF1 (N484, N470);
not NOT1 (N485, N478);
nor NOR3 (N486, N477, N435, N437);
and AND3 (N487, N483, N170, N394);
nor NOR2 (N488, N462, N377);
buf BUF1 (N489, N485);
and AND2 (N490, N475, N485);
buf BUF1 (N491, N484);
buf BUF1 (N492, N486);
buf BUF1 (N493, N467);
nor NOR4 (N494, N493, N158, N196, N429);
xor XOR2 (N495, N488, N224);
and AND4 (N496, N481, N452, N92, N78);
xor XOR2 (N497, N495, N330);
and AND3 (N498, N490, N384, N73);
nand NAND2 (N499, N496, N14);
and AND4 (N500, N494, N6, N332, N414);
and AND4 (N501, N499, N17, N73, N500);
and AND3 (N502, N161, N292, N75);
nor NOR4 (N503, N487, N424, N173, N270);
xor XOR2 (N504, N492, N175);
and AND3 (N505, N482, N376, N193);
or OR3 (N506, N504, N476, N459);
nor NOR3 (N507, N505, N74, N41);
and AND3 (N508, N498, N389, N298);
nand NAND3 (N509, N501, N300, N444);
nand NAND2 (N510, N508, N443);
nand NAND3 (N511, N510, N347, N448);
nor NOR2 (N512, N489, N164);
nand NAND2 (N513, N511, N316);
and AND3 (N514, N502, N416, N341);
not NOT1 (N515, N503);
and AND3 (N516, N507, N188, N105);
xor XOR2 (N517, N516, N418);
xor XOR2 (N518, N514, N156);
buf BUF1 (N519, N517);
nand NAND3 (N520, N480, N234, N328);
nand NAND2 (N521, N518, N383);
nor NOR2 (N522, N520, N242);
xor XOR2 (N523, N506, N75);
and AND4 (N524, N497, N235, N508, N126);
or OR4 (N525, N509, N127, N162, N244);
or OR2 (N526, N522, N245);
not NOT1 (N527, N513);
nand NAND3 (N528, N526, N176, N357);
nor NOR3 (N529, N491, N361, N26);
or OR3 (N530, N515, N308, N314);
buf BUF1 (N531, N521);
or OR3 (N532, N512, N72, N64);
nor NOR2 (N533, N523, N145);
not NOT1 (N534, N533);
nand NAND2 (N535, N532, N248);
or OR2 (N536, N529, N100);
nor NOR3 (N537, N519, N411, N18);
buf BUF1 (N538, N525);
buf BUF1 (N539, N531);
buf BUF1 (N540, N539);
and AND4 (N541, N528, N91, N352, N26);
nor NOR2 (N542, N538, N419);
nor NOR3 (N543, N530, N166, N93);
not NOT1 (N544, N527);
or OR2 (N545, N543, N157);
xor XOR2 (N546, N545, N485);
nand NAND3 (N547, N536, N125, N351);
nor NOR3 (N548, N547, N311, N209);
and AND4 (N549, N541, N466, N421, N303);
buf BUF1 (N550, N534);
or OR4 (N551, N546, N168, N212, N126);
nand NAND3 (N552, N550, N258, N339);
or OR2 (N553, N540, N105);
or OR2 (N554, N542, N298);
nand NAND3 (N555, N544, N392, N161);
nand NAND2 (N556, N553, N389);
and AND4 (N557, N555, N350, N225, N467);
and AND3 (N558, N548, N520, N47);
buf BUF1 (N559, N535);
and AND3 (N560, N551, N74, N174);
or OR2 (N561, N549, N280);
xor XOR2 (N562, N558, N413);
nor NOR4 (N563, N559, N60, N517, N356);
and AND2 (N564, N537, N78);
nor NOR2 (N565, N562, N278);
nor NOR2 (N566, N564, N123);
not NOT1 (N567, N566);
not NOT1 (N568, N567);
or OR4 (N569, N556, N428, N347, N4);
nand NAND4 (N570, N563, N3, N26, N241);
buf BUF1 (N571, N554);
nor NOR3 (N572, N569, N266, N399);
nand NAND3 (N573, N557, N541, N485);
nand NAND3 (N574, N568, N323, N30);
nor NOR2 (N575, N561, N398);
or OR3 (N576, N552, N48, N119);
xor XOR2 (N577, N572, N154);
xor XOR2 (N578, N577, N250);
buf BUF1 (N579, N578);
or OR4 (N580, N576, N451, N8, N242);
nor NOR2 (N581, N580, N552);
or OR3 (N582, N573, N335, N297);
xor XOR2 (N583, N570, N70);
or OR3 (N584, N571, N276, N407);
nor NOR3 (N585, N575, N276, N219);
and AND3 (N586, N583, N303, N166);
xor XOR2 (N587, N581, N146);
nor NOR3 (N588, N585, N386, N568);
xor XOR2 (N589, N574, N104);
not NOT1 (N590, N579);
nor NOR4 (N591, N589, N138, N111, N12);
or OR3 (N592, N588, N246, N120);
or OR2 (N593, N586, N96);
or OR2 (N594, N593, N372);
and AND3 (N595, N582, N550, N20);
nand NAND4 (N596, N560, N355, N264, N228);
and AND2 (N597, N595, N222);
xor XOR2 (N598, N565, N233);
and AND4 (N599, N597, N588, N273, N338);
xor XOR2 (N600, N592, N90);
nand NAND4 (N601, N598, N303, N335, N236);
nand NAND3 (N602, N587, N552, N472);
buf BUF1 (N603, N584);
or OR4 (N604, N596, N523, N271, N328);
and AND3 (N605, N601, N45, N220);
or OR4 (N606, N524, N263, N595, N564);
and AND2 (N607, N591, N572);
and AND4 (N608, N606, N115, N58, N362);
and AND3 (N609, N603, N308, N465);
nor NOR3 (N610, N608, N550, N374);
and AND4 (N611, N604, N588, N541, N357);
nand NAND4 (N612, N599, N553, N528, N92);
or OR2 (N613, N590, N224);
or OR2 (N614, N610, N181);
not NOT1 (N615, N602);
not NOT1 (N616, N605);
buf BUF1 (N617, N600);
not NOT1 (N618, N594);
and AND4 (N619, N614, N308, N5, N334);
nand NAND3 (N620, N616, N554, N467);
or OR3 (N621, N611, N416, N393);
or OR3 (N622, N619, N57, N418);
and AND3 (N623, N609, N495, N19);
or OR2 (N624, N623, N127);
or OR3 (N625, N624, N524, N616);
not NOT1 (N626, N622);
nand NAND3 (N627, N613, N177, N374);
nor NOR2 (N628, N626, N259);
buf BUF1 (N629, N628);
xor XOR2 (N630, N615, N298);
not NOT1 (N631, N617);
xor XOR2 (N632, N625, N339);
and AND4 (N633, N612, N480, N235, N446);
or OR3 (N634, N621, N222, N201);
not NOT1 (N635, N632);
xor XOR2 (N636, N635, N463);
buf BUF1 (N637, N620);
nor NOR2 (N638, N637, N456);
not NOT1 (N639, N607);
or OR2 (N640, N618, N4);
nor NOR2 (N641, N634, N635);
buf BUF1 (N642, N636);
nor NOR2 (N643, N638, N385);
and AND3 (N644, N639, N430, N462);
xor XOR2 (N645, N643, N273);
xor XOR2 (N646, N633, N363);
buf BUF1 (N647, N629);
xor XOR2 (N648, N647, N319);
nand NAND3 (N649, N642, N402, N198);
or OR2 (N650, N644, N460);
not NOT1 (N651, N630);
nor NOR2 (N652, N651, N38);
xor XOR2 (N653, N640, N96);
nand NAND2 (N654, N645, N612);
nand NAND4 (N655, N649, N50, N570, N359);
nor NOR3 (N656, N648, N326, N644);
nor NOR3 (N657, N641, N38, N611);
not NOT1 (N658, N654);
not NOT1 (N659, N656);
buf BUF1 (N660, N659);
or OR2 (N661, N652, N373);
nand NAND4 (N662, N660, N127, N173, N501);
xor XOR2 (N663, N657, N536);
not NOT1 (N664, N658);
nor NOR4 (N665, N631, N248, N314, N236);
and AND3 (N666, N653, N425, N286);
nor NOR4 (N667, N664, N173, N135, N422);
not NOT1 (N668, N655);
xor XOR2 (N669, N663, N561);
and AND4 (N670, N646, N561, N511, N248);
or OR3 (N671, N667, N599, N211);
not NOT1 (N672, N669);
nand NAND2 (N673, N672, N1);
and AND3 (N674, N650, N112, N313);
not NOT1 (N675, N673);
not NOT1 (N676, N674);
nor NOR3 (N677, N668, N392, N435);
not NOT1 (N678, N666);
nor NOR4 (N679, N675, N92, N61, N143);
and AND2 (N680, N677, N639);
xor XOR2 (N681, N678, N337);
xor XOR2 (N682, N679, N548);
and AND4 (N683, N662, N213, N672, N273);
nor NOR2 (N684, N676, N103);
not NOT1 (N685, N680);
nor NOR4 (N686, N670, N556, N475, N519);
xor XOR2 (N687, N686, N435);
not NOT1 (N688, N661);
xor XOR2 (N689, N688, N169);
buf BUF1 (N690, N684);
and AND4 (N691, N671, N525, N150, N23);
nor NOR4 (N692, N665, N514, N180, N194);
nand NAND4 (N693, N682, N240, N117, N402);
and AND3 (N694, N691, N281, N13);
or OR4 (N695, N685, N235, N421, N664);
not NOT1 (N696, N694);
or OR4 (N697, N690, N355, N586, N355);
and AND4 (N698, N683, N341, N502, N645);
xor XOR2 (N699, N697, N413);
not NOT1 (N700, N687);
and AND2 (N701, N692, N215);
not NOT1 (N702, N699);
not NOT1 (N703, N700);
nand NAND3 (N704, N702, N621, N351);
or OR4 (N705, N698, N20, N335, N553);
not NOT1 (N706, N704);
xor XOR2 (N707, N703, N225);
not NOT1 (N708, N689);
not NOT1 (N709, N695);
or OR2 (N710, N705, N195);
buf BUF1 (N711, N706);
and AND4 (N712, N711, N321, N653, N276);
and AND2 (N713, N701, N548);
xor XOR2 (N714, N707, N326);
or OR3 (N715, N627, N312, N326);
not NOT1 (N716, N708);
nand NAND3 (N717, N710, N475, N83);
buf BUF1 (N718, N715);
and AND3 (N719, N681, N339, N62);
buf BUF1 (N720, N713);
buf BUF1 (N721, N712);
nand NAND3 (N722, N693, N676, N83);
nor NOR4 (N723, N714, N51, N411, N286);
buf BUF1 (N724, N716);
xor XOR2 (N725, N718, N583);
nand NAND2 (N726, N720, N17);
not NOT1 (N727, N719);
and AND3 (N728, N721, N357, N363);
nand NAND3 (N729, N723, N40, N44);
and AND4 (N730, N696, N255, N438, N538);
nand NAND4 (N731, N722, N442, N686, N264);
not NOT1 (N732, N717);
buf BUF1 (N733, N727);
not NOT1 (N734, N729);
and AND4 (N735, N734, N172, N268, N170);
xor XOR2 (N736, N725, N700);
nor NOR4 (N737, N728, N409, N243, N546);
xor XOR2 (N738, N732, N110);
not NOT1 (N739, N709);
or OR4 (N740, N738, N234, N625, N466);
buf BUF1 (N741, N739);
buf BUF1 (N742, N730);
and AND3 (N743, N733, N392, N19);
nor NOR3 (N744, N726, N268, N84);
xor XOR2 (N745, N744, N187);
and AND3 (N746, N741, N615, N311);
or OR3 (N747, N731, N128, N544);
and AND3 (N748, N746, N63, N625);
buf BUF1 (N749, N743);
nor NOR3 (N750, N740, N98, N379);
buf BUF1 (N751, N748);
nor NOR4 (N752, N750, N343, N272, N154);
not NOT1 (N753, N745);
buf BUF1 (N754, N752);
nand NAND3 (N755, N742, N475, N107);
and AND4 (N756, N755, N529, N515, N510);
nand NAND2 (N757, N724, N693);
not NOT1 (N758, N736);
xor XOR2 (N759, N756, N616);
nor NOR4 (N760, N753, N688, N653, N10);
xor XOR2 (N761, N754, N456);
or OR4 (N762, N735, N272, N600, N476);
nand NAND4 (N763, N758, N180, N478, N196);
buf BUF1 (N764, N751);
nor NOR2 (N765, N762, N674);
and AND4 (N766, N763, N592, N666, N157);
not NOT1 (N767, N766);
or OR3 (N768, N760, N195, N735);
xor XOR2 (N769, N765, N413);
nand NAND4 (N770, N767, N397, N30, N338);
nand NAND3 (N771, N761, N295, N573);
nor NOR3 (N772, N749, N153, N411);
not NOT1 (N773, N737);
not NOT1 (N774, N747);
xor XOR2 (N775, N774, N772);
and AND3 (N776, N176, N535, N80);
xor XOR2 (N777, N768, N608);
or OR3 (N778, N759, N441, N527);
not NOT1 (N779, N769);
not NOT1 (N780, N775);
buf BUF1 (N781, N780);
or OR2 (N782, N764, N366);
xor XOR2 (N783, N781, N151);
nor NOR3 (N784, N778, N574, N405);
not NOT1 (N785, N771);
buf BUF1 (N786, N779);
buf BUF1 (N787, N786);
or OR2 (N788, N757, N189);
and AND3 (N789, N788, N360, N666);
and AND2 (N790, N776, N146);
buf BUF1 (N791, N787);
or OR2 (N792, N791, N170);
nor NOR2 (N793, N783, N576);
nand NAND3 (N794, N773, N642, N526);
nor NOR4 (N795, N793, N616, N197, N665);
nor NOR2 (N796, N777, N471);
nand NAND3 (N797, N792, N504, N180);
nor NOR2 (N798, N785, N80);
not NOT1 (N799, N796);
buf BUF1 (N800, N798);
not NOT1 (N801, N782);
xor XOR2 (N802, N770, N178);
not NOT1 (N803, N799);
xor XOR2 (N804, N802, N701);
nand NAND4 (N805, N790, N328, N762, N611);
not NOT1 (N806, N795);
buf BUF1 (N807, N804);
nand NAND4 (N808, N806, N362, N669, N182);
xor XOR2 (N809, N794, N766);
xor XOR2 (N810, N807, N525);
or OR4 (N811, N784, N109, N30, N309);
nand NAND2 (N812, N810, N164);
and AND2 (N813, N805, N497);
buf BUF1 (N814, N813);
not NOT1 (N815, N797);
not NOT1 (N816, N800);
xor XOR2 (N817, N815, N15);
or OR2 (N818, N789, N564);
buf BUF1 (N819, N811);
nor NOR4 (N820, N803, N311, N22, N557);
xor XOR2 (N821, N819, N145);
buf BUF1 (N822, N816);
not NOT1 (N823, N808);
not NOT1 (N824, N817);
xor XOR2 (N825, N801, N243);
or OR2 (N826, N809, N596);
not NOT1 (N827, N823);
not NOT1 (N828, N820);
buf BUF1 (N829, N814);
and AND4 (N830, N828, N701, N30, N429);
or OR2 (N831, N830, N105);
xor XOR2 (N832, N827, N365);
or OR3 (N833, N829, N61, N616);
buf BUF1 (N834, N831);
xor XOR2 (N835, N825, N375);
and AND3 (N836, N812, N21, N598);
xor XOR2 (N837, N832, N215);
not NOT1 (N838, N834);
nand NAND3 (N839, N833, N245, N813);
or OR2 (N840, N824, N110);
and AND3 (N841, N837, N780, N85);
xor XOR2 (N842, N826, N760);
nand NAND4 (N843, N818, N60, N218, N438);
xor XOR2 (N844, N843, N618);
buf BUF1 (N845, N844);
or OR2 (N846, N838, N466);
buf BUF1 (N847, N822);
buf BUF1 (N848, N840);
buf BUF1 (N849, N847);
nor NOR3 (N850, N848, N85, N117);
nand NAND2 (N851, N841, N495);
and AND2 (N852, N851, N232);
nand NAND4 (N853, N821, N747, N336, N91);
or OR2 (N854, N850, N567);
nand NAND2 (N855, N839, N17);
nand NAND3 (N856, N849, N445, N841);
nand NAND4 (N857, N855, N557, N340, N474);
or OR4 (N858, N835, N531, N518, N674);
buf BUF1 (N859, N852);
nor NOR3 (N860, N858, N229, N702);
buf BUF1 (N861, N853);
nor NOR2 (N862, N857, N777);
and AND3 (N863, N845, N96, N394);
buf BUF1 (N864, N854);
not NOT1 (N865, N861);
nand NAND4 (N866, N856, N846, N361, N582);
xor XOR2 (N867, N95, N381);
and AND3 (N868, N862, N255, N179);
nor NOR3 (N869, N860, N736, N585);
nand NAND3 (N870, N867, N848, N868);
not NOT1 (N871, N654);
nand NAND4 (N872, N864, N133, N160, N767);
or OR2 (N873, N859, N512);
and AND4 (N874, N863, N107, N371, N288);
buf BUF1 (N875, N865);
nor NOR2 (N876, N869, N868);
or OR4 (N877, N870, N127, N649, N683);
or OR2 (N878, N875, N52);
not NOT1 (N879, N878);
not NOT1 (N880, N872);
xor XOR2 (N881, N880, N713);
nor NOR4 (N882, N873, N410, N726, N5);
or OR3 (N883, N882, N16, N390);
nor NOR4 (N884, N881, N779, N49, N399);
nand NAND4 (N885, N842, N169, N625, N512);
buf BUF1 (N886, N871);
or OR3 (N887, N885, N14, N611);
nor NOR3 (N888, N887, N739, N795);
and AND2 (N889, N884, N389);
xor XOR2 (N890, N888, N372);
nand NAND4 (N891, N876, N18, N456, N409);
nor NOR2 (N892, N891, N255);
buf BUF1 (N893, N877);
and AND3 (N894, N893, N832, N680);
buf BUF1 (N895, N883);
and AND3 (N896, N836, N494, N815);
and AND4 (N897, N874, N734, N687, N672);
not NOT1 (N898, N896);
nor NOR2 (N899, N866, N310);
or OR2 (N900, N889, N200);
or OR4 (N901, N886, N119, N861, N780);
buf BUF1 (N902, N890);
buf BUF1 (N903, N895);
xor XOR2 (N904, N879, N844);
not NOT1 (N905, N892);
and AND2 (N906, N905, N656);
not NOT1 (N907, N899);
and AND4 (N908, N900, N619, N318, N445);
and AND2 (N909, N902, N339);
xor XOR2 (N910, N894, N358);
buf BUF1 (N911, N910);
or OR4 (N912, N898, N854, N291, N775);
nor NOR4 (N913, N911, N864, N288, N748);
not NOT1 (N914, N903);
buf BUF1 (N915, N906);
nand NAND4 (N916, N901, N895, N361, N793);
xor XOR2 (N917, N897, N731);
not NOT1 (N918, N913);
buf BUF1 (N919, N914);
xor XOR2 (N920, N915, N714);
nor NOR4 (N921, N907, N219, N252, N115);
or OR2 (N922, N918, N134);
and AND4 (N923, N921, N218, N168, N77);
buf BUF1 (N924, N908);
and AND2 (N925, N922, N593);
xor XOR2 (N926, N919, N527);
xor XOR2 (N927, N904, N225);
not NOT1 (N928, N917);
xor XOR2 (N929, N916, N661);
nor NOR2 (N930, N929, N124);
nor NOR3 (N931, N909, N420, N659);
and AND2 (N932, N927, N294);
and AND3 (N933, N912, N710, N880);
buf BUF1 (N934, N926);
not NOT1 (N935, N934);
nor NOR2 (N936, N923, N854);
buf BUF1 (N937, N925);
or OR4 (N938, N924, N397, N218, N300);
not NOT1 (N939, N935);
and AND2 (N940, N936, N499);
not NOT1 (N941, N930);
xor XOR2 (N942, N941, N430);
nand NAND3 (N943, N940, N209, N510);
xor XOR2 (N944, N928, N151);
not NOT1 (N945, N937);
nand NAND3 (N946, N932, N500, N424);
xor XOR2 (N947, N943, N447);
xor XOR2 (N948, N946, N267);
nand NAND3 (N949, N938, N137, N859);
nor NOR4 (N950, N939, N838, N534, N294);
buf BUF1 (N951, N920);
not NOT1 (N952, N944);
xor XOR2 (N953, N947, N479);
and AND4 (N954, N952, N656, N260, N630);
not NOT1 (N955, N933);
buf BUF1 (N956, N950);
xor XOR2 (N957, N953, N58);
xor XOR2 (N958, N951, N58);
or OR2 (N959, N954, N409);
xor XOR2 (N960, N956, N274);
not NOT1 (N961, N931);
xor XOR2 (N962, N957, N236);
nand NAND3 (N963, N948, N240, N16);
not NOT1 (N964, N963);
buf BUF1 (N965, N961);
buf BUF1 (N966, N965);
not NOT1 (N967, N958);
nand NAND2 (N968, N959, N731);
or OR3 (N969, N945, N730, N833);
nand NAND2 (N970, N967, N967);
nor NOR4 (N971, N968, N874, N729, N738);
and AND3 (N972, N955, N924, N84);
buf BUF1 (N973, N949);
and AND3 (N974, N973, N290, N317);
or OR2 (N975, N960, N715);
not NOT1 (N976, N975);
buf BUF1 (N977, N972);
and AND4 (N978, N976, N71, N359, N606);
nor NOR2 (N979, N942, N150);
not NOT1 (N980, N971);
not NOT1 (N981, N978);
xor XOR2 (N982, N981, N415);
xor XOR2 (N983, N980, N79);
nand NAND2 (N984, N962, N60);
xor XOR2 (N985, N984, N829);
xor XOR2 (N986, N969, N948);
or OR3 (N987, N983, N808, N543);
not NOT1 (N988, N974);
and AND2 (N989, N964, N29);
nand NAND3 (N990, N970, N815, N40);
nor NOR3 (N991, N987, N874, N638);
nand NAND2 (N992, N977, N625);
xor XOR2 (N993, N985, N360);
and AND2 (N994, N986, N590);
and AND4 (N995, N989, N419, N817, N86);
nor NOR2 (N996, N993, N460);
not NOT1 (N997, N991);
not NOT1 (N998, N997);
or OR3 (N999, N992, N55, N891);
not NOT1 (N1000, N995);
not NOT1 (N1001, N966);
xor XOR2 (N1002, N999, N982);
not NOT1 (N1003, N666);
nand NAND3 (N1004, N979, N945, N763);
xor XOR2 (N1005, N1004, N908);
and AND3 (N1006, N1002, N589, N53);
xor XOR2 (N1007, N998, N678);
nand NAND2 (N1008, N1006, N650);
buf BUF1 (N1009, N1005);
nor NOR2 (N1010, N1001, N253);
not NOT1 (N1011, N1009);
buf BUF1 (N1012, N1003);
nor NOR4 (N1013, N1010, N712, N754, N844);
nand NAND2 (N1014, N1013, N959);
not NOT1 (N1015, N988);
and AND2 (N1016, N1000, N122);
buf BUF1 (N1017, N1008);
or OR3 (N1018, N1017, N80, N389);
and AND4 (N1019, N1015, N271, N225, N510);
nor NOR3 (N1020, N1014, N403, N784);
xor XOR2 (N1021, N1007, N365);
nor NOR3 (N1022, N1011, N384, N976);
or OR3 (N1023, N1016, N474, N235);
nand NAND2 (N1024, N990, N646);
nand NAND3 (N1025, N994, N941, N755);
nor NOR4 (N1026, N1023, N427, N796, N8);
and AND4 (N1027, N1012, N389, N465, N570);
nand NAND4 (N1028, N1024, N1010, N996, N515);
not NOT1 (N1029, N573);
and AND3 (N1030, N1028, N343, N815);
buf BUF1 (N1031, N1027);
nand NAND2 (N1032, N1019, N336);
nand NAND4 (N1033, N1022, N545, N961, N365);
nand NAND3 (N1034, N1018, N1001, N404);
not NOT1 (N1035, N1030);
nor NOR3 (N1036, N1025, N378, N118);
not NOT1 (N1037, N1036);
nand NAND2 (N1038, N1026, N464);
xor XOR2 (N1039, N1034, N219);
xor XOR2 (N1040, N1032, N615);
not NOT1 (N1041, N1031);
nand NAND4 (N1042, N1041, N401, N387, N777);
or OR4 (N1043, N1037, N371, N444, N812);
xor XOR2 (N1044, N1021, N849);
xor XOR2 (N1045, N1035, N378);
buf BUF1 (N1046, N1045);
and AND3 (N1047, N1020, N515, N722);
and AND2 (N1048, N1044, N734);
or OR4 (N1049, N1048, N975, N919, N1005);
xor XOR2 (N1050, N1039, N862);
not NOT1 (N1051, N1040);
and AND4 (N1052, N1042, N1015, N949, N853);
xor XOR2 (N1053, N1050, N1014);
and AND2 (N1054, N1051, N953);
not NOT1 (N1055, N1043);
or OR2 (N1056, N1055, N24);
nand NAND3 (N1057, N1033, N573, N166);
buf BUF1 (N1058, N1029);
xor XOR2 (N1059, N1057, N18);
buf BUF1 (N1060, N1058);
nor NOR4 (N1061, N1038, N570, N445, N806);
not NOT1 (N1062, N1047);
or OR3 (N1063, N1059, N525, N722);
or OR4 (N1064, N1049, N1001, N640, N194);
or OR3 (N1065, N1061, N204, N440);
nand NAND4 (N1066, N1052, N602, N33, N407);
xor XOR2 (N1067, N1060, N984);
xor XOR2 (N1068, N1065, N706);
or OR2 (N1069, N1062, N239);
not NOT1 (N1070, N1067);
xor XOR2 (N1071, N1066, N565);
buf BUF1 (N1072, N1053);
xor XOR2 (N1073, N1071, N190);
or OR2 (N1074, N1064, N155);
not NOT1 (N1075, N1069);
xor XOR2 (N1076, N1074, N552);
xor XOR2 (N1077, N1073, N924);
or OR3 (N1078, N1070, N955, N999);
and AND4 (N1079, N1078, N543, N835, N124);
not NOT1 (N1080, N1077);
xor XOR2 (N1081, N1068, N938);
xor XOR2 (N1082, N1080, N33);
nor NOR2 (N1083, N1056, N301);
buf BUF1 (N1084, N1054);
and AND2 (N1085, N1079, N865);
or OR4 (N1086, N1063, N481, N543, N906);
buf BUF1 (N1087, N1084);
or OR3 (N1088, N1081, N186, N141);
nand NAND2 (N1089, N1086, N366);
xor XOR2 (N1090, N1085, N18);
buf BUF1 (N1091, N1083);
or OR3 (N1092, N1076, N817, N274);
nand NAND4 (N1093, N1075, N524, N899, N551);
and AND3 (N1094, N1092, N220, N988);
not NOT1 (N1095, N1093);
buf BUF1 (N1096, N1091);
nor NOR4 (N1097, N1087, N906, N467, N378);
buf BUF1 (N1098, N1089);
nor NOR3 (N1099, N1097, N954, N911);
or OR3 (N1100, N1096, N680, N428);
xor XOR2 (N1101, N1072, N338);
nand NAND2 (N1102, N1082, N1054);
nand NAND3 (N1103, N1098, N563, N219);
not NOT1 (N1104, N1099);
not NOT1 (N1105, N1104);
xor XOR2 (N1106, N1094, N66);
buf BUF1 (N1107, N1101);
and AND3 (N1108, N1095, N561, N144);
buf BUF1 (N1109, N1046);
not NOT1 (N1110, N1107);
not NOT1 (N1111, N1088);
nor NOR3 (N1112, N1106, N54, N814);
nor NOR3 (N1113, N1102, N743, N237);
and AND4 (N1114, N1103, N591, N628, N126);
nor NOR2 (N1115, N1112, N606);
xor XOR2 (N1116, N1105, N667);
or OR3 (N1117, N1109, N648, N983);
nor NOR4 (N1118, N1113, N1095, N550, N1096);
buf BUF1 (N1119, N1108);
nor NOR3 (N1120, N1114, N286, N185);
buf BUF1 (N1121, N1120);
not NOT1 (N1122, N1121);
or OR4 (N1123, N1122, N264, N688, N639);
xor XOR2 (N1124, N1116, N1090);
and AND3 (N1125, N880, N432, N680);
and AND3 (N1126, N1124, N890, N399);
nor NOR3 (N1127, N1115, N812, N599);
or OR4 (N1128, N1111, N470, N176, N897);
or OR4 (N1129, N1127, N243, N1025, N129);
and AND3 (N1130, N1117, N546, N844);
xor XOR2 (N1131, N1130, N368);
or OR4 (N1132, N1129, N885, N176, N656);
or OR4 (N1133, N1125, N971, N846, N894);
buf BUF1 (N1134, N1119);
and AND3 (N1135, N1131, N375, N1075);
nand NAND2 (N1136, N1132, N342);
and AND4 (N1137, N1135, N903, N1119, N171);
and AND2 (N1138, N1100, N90);
not NOT1 (N1139, N1137);
buf BUF1 (N1140, N1136);
not NOT1 (N1141, N1110);
or OR2 (N1142, N1123, N700);
or OR2 (N1143, N1128, N721);
and AND2 (N1144, N1141, N1080);
or OR3 (N1145, N1133, N897, N66);
buf BUF1 (N1146, N1145);
not NOT1 (N1147, N1146);
or OR2 (N1148, N1143, N890);
nor NOR3 (N1149, N1140, N594, N1060);
and AND4 (N1150, N1126, N216, N1118, N123);
or OR4 (N1151, N125, N1080, N93, N292);
xor XOR2 (N1152, N1147, N901);
not NOT1 (N1153, N1150);
xor XOR2 (N1154, N1142, N547);
buf BUF1 (N1155, N1154);
not NOT1 (N1156, N1155);
nor NOR3 (N1157, N1148, N389, N273);
nor NOR3 (N1158, N1153, N575, N475);
xor XOR2 (N1159, N1138, N1107);
xor XOR2 (N1160, N1152, N500);
xor XOR2 (N1161, N1149, N1004);
or OR3 (N1162, N1157, N569, N476);
xor XOR2 (N1163, N1134, N527);
and AND2 (N1164, N1151, N41);
nor NOR2 (N1165, N1160, N1130);
xor XOR2 (N1166, N1156, N450);
nor NOR4 (N1167, N1163, N572, N820, N352);
nor NOR2 (N1168, N1166, N1050);
or OR2 (N1169, N1164, N364);
not NOT1 (N1170, N1144);
not NOT1 (N1171, N1169);
not NOT1 (N1172, N1139);
buf BUF1 (N1173, N1158);
and AND2 (N1174, N1162, N1069);
buf BUF1 (N1175, N1165);
nor NOR4 (N1176, N1173, N868, N470, N177);
or OR4 (N1177, N1176, N507, N187, N559);
or OR2 (N1178, N1171, N610);
not NOT1 (N1179, N1159);
xor XOR2 (N1180, N1170, N419);
nand NAND4 (N1181, N1178, N278, N400, N485);
not NOT1 (N1182, N1180);
buf BUF1 (N1183, N1179);
or OR4 (N1184, N1174, N1123, N479, N927);
or OR4 (N1185, N1161, N574, N187, N493);
nand NAND2 (N1186, N1183, N1170);
nor NOR4 (N1187, N1184, N784, N1162, N896);
xor XOR2 (N1188, N1182, N976);
and AND3 (N1189, N1168, N259, N485);
and AND3 (N1190, N1172, N378, N940);
nand NAND2 (N1191, N1175, N366);
nand NAND3 (N1192, N1177, N396, N981);
nand NAND4 (N1193, N1188, N70, N280, N701);
nand NAND2 (N1194, N1167, N112);
and AND3 (N1195, N1186, N385, N289);
and AND4 (N1196, N1194, N307, N25, N1190);
nand NAND2 (N1197, N612, N481);
and AND4 (N1198, N1187, N279, N162, N887);
buf BUF1 (N1199, N1193);
xor XOR2 (N1200, N1195, N1016);
nand NAND3 (N1201, N1192, N329, N113);
or OR3 (N1202, N1197, N1147, N370);
and AND2 (N1203, N1201, N854);
xor XOR2 (N1204, N1198, N500);
buf BUF1 (N1205, N1203);
and AND4 (N1206, N1185, N590, N476, N881);
xor XOR2 (N1207, N1191, N514);
buf BUF1 (N1208, N1204);
nand NAND2 (N1209, N1202, N619);
xor XOR2 (N1210, N1207, N201);
and AND4 (N1211, N1210, N864, N1096, N957);
buf BUF1 (N1212, N1181);
buf BUF1 (N1213, N1205);
and AND4 (N1214, N1189, N967, N266, N367);
or OR3 (N1215, N1213, N162, N1195);
buf BUF1 (N1216, N1211);
nor NOR3 (N1217, N1206, N1108, N49);
and AND4 (N1218, N1208, N406, N293, N728);
nand NAND3 (N1219, N1212, N23, N287);
xor XOR2 (N1220, N1214, N798);
or OR3 (N1221, N1215, N451, N891);
or OR4 (N1222, N1199, N886, N1177, N671);
not NOT1 (N1223, N1209);
or OR3 (N1224, N1200, N56, N869);
or OR2 (N1225, N1220, N954);
buf BUF1 (N1226, N1222);
or OR3 (N1227, N1225, N449, N275);
buf BUF1 (N1228, N1223);
buf BUF1 (N1229, N1216);
xor XOR2 (N1230, N1218, N840);
or OR4 (N1231, N1227, N220, N400, N407);
not NOT1 (N1232, N1224);
and AND4 (N1233, N1231, N284, N24, N438);
xor XOR2 (N1234, N1217, N1097);
nor NOR4 (N1235, N1233, N1124, N19, N256);
nand NAND2 (N1236, N1235, N374);
and AND3 (N1237, N1234, N805, N1025);
or OR4 (N1238, N1230, N1211, N580, N1128);
buf BUF1 (N1239, N1236);
not NOT1 (N1240, N1239);
not NOT1 (N1241, N1229);
and AND2 (N1242, N1219, N223);
xor XOR2 (N1243, N1226, N554);
xor XOR2 (N1244, N1232, N688);
buf BUF1 (N1245, N1238);
not NOT1 (N1246, N1228);
nor NOR4 (N1247, N1244, N143, N995, N582);
buf BUF1 (N1248, N1245);
xor XOR2 (N1249, N1221, N476);
xor XOR2 (N1250, N1237, N205);
xor XOR2 (N1251, N1249, N200);
xor XOR2 (N1252, N1246, N578);
nand NAND4 (N1253, N1252, N267, N849, N784);
buf BUF1 (N1254, N1250);
xor XOR2 (N1255, N1196, N421);
or OR3 (N1256, N1241, N641, N76);
and AND3 (N1257, N1243, N549, N1028);
buf BUF1 (N1258, N1242);
nand NAND3 (N1259, N1248, N834, N921);
nand NAND2 (N1260, N1255, N555);
buf BUF1 (N1261, N1258);
xor XOR2 (N1262, N1251, N1227);
nand NAND2 (N1263, N1261, N1046);
not NOT1 (N1264, N1247);
or OR4 (N1265, N1240, N1239, N394, N596);
nand NAND4 (N1266, N1259, N51, N318, N596);
or OR4 (N1267, N1263, N252, N1251, N1099);
and AND3 (N1268, N1260, N339, N922);
nor NOR4 (N1269, N1267, N45, N169, N759);
not NOT1 (N1270, N1254);
and AND3 (N1271, N1253, N961, N1130);
buf BUF1 (N1272, N1268);
or OR3 (N1273, N1264, N136, N11);
xor XOR2 (N1274, N1256, N535);
nand NAND4 (N1275, N1271, N986, N958, N95);
xor XOR2 (N1276, N1272, N85);
or OR4 (N1277, N1265, N865, N677, N471);
not NOT1 (N1278, N1277);
nand NAND4 (N1279, N1275, N830, N755, N497);
and AND2 (N1280, N1266, N313);
nor NOR4 (N1281, N1280, N329, N664, N646);
nand NAND2 (N1282, N1262, N1026);
buf BUF1 (N1283, N1257);
nor NOR2 (N1284, N1270, N296);
not NOT1 (N1285, N1284);
xor XOR2 (N1286, N1278, N166);
buf BUF1 (N1287, N1286);
buf BUF1 (N1288, N1273);
nor NOR3 (N1289, N1287, N1155, N835);
xor XOR2 (N1290, N1282, N545);
nand NAND3 (N1291, N1274, N465, N834);
not NOT1 (N1292, N1291);
and AND2 (N1293, N1283, N225);
nand NAND2 (N1294, N1289, N618);
and AND4 (N1295, N1292, N334, N313, N537);
xor XOR2 (N1296, N1293, N782);
nand NAND2 (N1297, N1276, N1146);
and AND2 (N1298, N1297, N909);
not NOT1 (N1299, N1296);
not NOT1 (N1300, N1279);
and AND3 (N1301, N1294, N898, N1259);
buf BUF1 (N1302, N1295);
nand NAND2 (N1303, N1299, N83);
not NOT1 (N1304, N1298);
buf BUF1 (N1305, N1290);
nor NOR3 (N1306, N1269, N1157, N246);
xor XOR2 (N1307, N1285, N724);
nor NOR3 (N1308, N1303, N821, N723);
xor XOR2 (N1309, N1307, N210);
xor XOR2 (N1310, N1288, N1161);
nor NOR2 (N1311, N1310, N573);
buf BUF1 (N1312, N1311);
xor XOR2 (N1313, N1306, N714);
nand NAND2 (N1314, N1309, N374);
or OR4 (N1315, N1313, N89, N41, N632);
and AND3 (N1316, N1302, N384, N895);
xor XOR2 (N1317, N1300, N1032);
and AND2 (N1318, N1317, N190);
and AND2 (N1319, N1305, N373);
buf BUF1 (N1320, N1304);
nand NAND4 (N1321, N1318, N73, N619, N443);
and AND2 (N1322, N1301, N382);
xor XOR2 (N1323, N1314, N793);
xor XOR2 (N1324, N1322, N1023);
and AND2 (N1325, N1321, N120);
and AND2 (N1326, N1315, N356);
not NOT1 (N1327, N1308);
nor NOR2 (N1328, N1326, N760);
nand NAND4 (N1329, N1316, N580, N223, N909);
and AND3 (N1330, N1325, N584, N1175);
nor NOR2 (N1331, N1327, N1040);
xor XOR2 (N1332, N1320, N1112);
xor XOR2 (N1333, N1281, N1260);
buf BUF1 (N1334, N1331);
not NOT1 (N1335, N1323);
or OR4 (N1336, N1335, N129, N504, N680);
and AND4 (N1337, N1334, N468, N288, N1159);
and AND3 (N1338, N1336, N736, N408);
nand NAND4 (N1339, N1332, N275, N485, N737);
buf BUF1 (N1340, N1319);
or OR3 (N1341, N1340, N989, N622);
buf BUF1 (N1342, N1324);
buf BUF1 (N1343, N1333);
buf BUF1 (N1344, N1342);
or OR3 (N1345, N1329, N950, N1074);
and AND4 (N1346, N1341, N1079, N983, N771);
and AND4 (N1347, N1339, N1335, N455, N1344);
xor XOR2 (N1348, N1320, N713);
nand NAND2 (N1349, N1346, N1067);
nand NAND4 (N1350, N1347, N890, N572, N104);
and AND2 (N1351, N1330, N568);
or OR3 (N1352, N1348, N298, N950);
not NOT1 (N1353, N1345);
nand NAND3 (N1354, N1337, N803, N1208);
buf BUF1 (N1355, N1349);
nand NAND2 (N1356, N1352, N1198);
or OR4 (N1357, N1343, N172, N833, N1131);
buf BUF1 (N1358, N1351);
buf BUF1 (N1359, N1312);
nand NAND4 (N1360, N1338, N532, N656, N984);
buf BUF1 (N1361, N1360);
and AND3 (N1362, N1353, N140, N1153);
xor XOR2 (N1363, N1357, N1136);
buf BUF1 (N1364, N1361);
nor NOR3 (N1365, N1328, N1069, N94);
not NOT1 (N1366, N1362);
buf BUF1 (N1367, N1354);
xor XOR2 (N1368, N1355, N986);
not NOT1 (N1369, N1363);
nor NOR3 (N1370, N1356, N180, N128);
nor NOR3 (N1371, N1370, N221, N76);
nor NOR4 (N1372, N1367, N825, N1256, N40);
nor NOR4 (N1373, N1369, N1100, N1112, N714);
nor NOR3 (N1374, N1359, N902, N828);
xor XOR2 (N1375, N1372, N1143);
and AND2 (N1376, N1364, N185);
nor NOR3 (N1377, N1376, N2, N817);
nor NOR4 (N1378, N1368, N140, N1158, N894);
nor NOR4 (N1379, N1371, N1296, N444, N246);
nand NAND3 (N1380, N1375, N1160, N1166);
nor NOR3 (N1381, N1377, N506, N430);
nor NOR2 (N1382, N1366, N1258);
nand NAND2 (N1383, N1350, N1031);
nand NAND3 (N1384, N1358, N466, N972);
not NOT1 (N1385, N1382);
or OR2 (N1386, N1373, N374);
buf BUF1 (N1387, N1385);
xor XOR2 (N1388, N1384, N742);
or OR2 (N1389, N1383, N1232);
or OR4 (N1390, N1378, N1105, N841, N711);
or OR4 (N1391, N1381, N908, N507, N1085);
nor NOR2 (N1392, N1380, N576);
not NOT1 (N1393, N1374);
not NOT1 (N1394, N1393);
not NOT1 (N1395, N1394);
buf BUF1 (N1396, N1391);
buf BUF1 (N1397, N1392);
nor NOR3 (N1398, N1390, N1372, N717);
nand NAND2 (N1399, N1379, N938);
nor NOR4 (N1400, N1396, N183, N251, N1204);
buf BUF1 (N1401, N1399);
nand NAND4 (N1402, N1398, N1351, N508, N422);
xor XOR2 (N1403, N1395, N1360);
nand NAND3 (N1404, N1401, N116, N582);
or OR3 (N1405, N1389, N1256, N698);
and AND4 (N1406, N1402, N540, N878, N1161);
xor XOR2 (N1407, N1397, N656);
xor XOR2 (N1408, N1365, N1064);
or OR4 (N1409, N1405, N412, N1192, N269);
buf BUF1 (N1410, N1388);
and AND3 (N1411, N1386, N858, N796);
buf BUF1 (N1412, N1408);
buf BUF1 (N1413, N1400);
not NOT1 (N1414, N1404);
or OR4 (N1415, N1387, N1149, N1363, N1352);
and AND2 (N1416, N1415, N697);
buf BUF1 (N1417, N1412);
nor NOR2 (N1418, N1403, N185);
and AND2 (N1419, N1417, N464);
or OR3 (N1420, N1414, N1209, N177);
or OR4 (N1421, N1419, N1323, N79, N333);
nor NOR2 (N1422, N1421, N1135);
xor XOR2 (N1423, N1422, N855);
not NOT1 (N1424, N1418);
xor XOR2 (N1425, N1416, N196);
buf BUF1 (N1426, N1423);
buf BUF1 (N1427, N1426);
xor XOR2 (N1428, N1424, N320);
buf BUF1 (N1429, N1428);
buf BUF1 (N1430, N1410);
xor XOR2 (N1431, N1427, N422);
and AND3 (N1432, N1409, N701, N226);
xor XOR2 (N1433, N1431, N1168);
xor XOR2 (N1434, N1406, N721);
nand NAND2 (N1435, N1425, N96);
not NOT1 (N1436, N1413);
xor XOR2 (N1437, N1407, N1362);
and AND3 (N1438, N1437, N1140, N908);
xor XOR2 (N1439, N1432, N348);
nand NAND4 (N1440, N1438, N809, N167, N137);
nand NAND4 (N1441, N1433, N172, N1263, N1356);
not NOT1 (N1442, N1411);
nor NOR3 (N1443, N1439, N1111, N442);
buf BUF1 (N1444, N1434);
not NOT1 (N1445, N1442);
or OR2 (N1446, N1444, N455);
xor XOR2 (N1447, N1443, N1298);
nand NAND3 (N1448, N1447, N1253, N1139);
or OR3 (N1449, N1445, N719, N1002);
or OR4 (N1450, N1435, N1347, N1188, N390);
not NOT1 (N1451, N1436);
nor NOR4 (N1452, N1448, N770, N1122, N878);
not NOT1 (N1453, N1452);
xor XOR2 (N1454, N1429, N721);
nor NOR3 (N1455, N1430, N935, N811);
nor NOR3 (N1456, N1453, N386, N1361);
not NOT1 (N1457, N1449);
not NOT1 (N1458, N1420);
nor NOR2 (N1459, N1446, N152);
not NOT1 (N1460, N1456);
not NOT1 (N1461, N1440);
nor NOR2 (N1462, N1461, N209);
not NOT1 (N1463, N1458);
and AND3 (N1464, N1454, N1099, N267);
or OR3 (N1465, N1450, N591, N1153);
buf BUF1 (N1466, N1464);
nor NOR4 (N1467, N1460, N21, N922, N868);
buf BUF1 (N1468, N1457);
nand NAND2 (N1469, N1463, N665);
nand NAND3 (N1470, N1441, N1151, N1308);
nand NAND3 (N1471, N1466, N1015, N239);
nor NOR4 (N1472, N1462, N1456, N935, N599);
buf BUF1 (N1473, N1468);
not NOT1 (N1474, N1471);
or OR2 (N1475, N1459, N1270);
nand NAND4 (N1476, N1467, N1317, N355, N336);
xor XOR2 (N1477, N1455, N1421);
nor NOR4 (N1478, N1470, N218, N761, N248);
nor NOR4 (N1479, N1476, N1425, N320, N1199);
nor NOR3 (N1480, N1469, N1297, N165);
not NOT1 (N1481, N1451);
nor NOR2 (N1482, N1481, N914);
not NOT1 (N1483, N1473);
nand NAND3 (N1484, N1475, N1457, N1315);
nand NAND4 (N1485, N1465, N990, N773, N554);
buf BUF1 (N1486, N1480);
and AND4 (N1487, N1478, N615, N193, N858);
nor NOR2 (N1488, N1487, N1220);
not NOT1 (N1489, N1479);
nor NOR2 (N1490, N1484, N621);
nor NOR2 (N1491, N1472, N576);
nand NAND3 (N1492, N1490, N788, N1323);
buf BUF1 (N1493, N1486);
and AND2 (N1494, N1488, N590);
buf BUF1 (N1495, N1489);
nand NAND3 (N1496, N1483, N690, N926);
nor NOR3 (N1497, N1493, N808, N621);
and AND3 (N1498, N1474, N1464, N803);
and AND3 (N1499, N1477, N1477, N445);
nand NAND4 (N1500, N1485, N123, N560, N1335);
not NOT1 (N1501, N1494);
nor NOR2 (N1502, N1482, N336);
not NOT1 (N1503, N1491);
not NOT1 (N1504, N1502);
not NOT1 (N1505, N1504);
xor XOR2 (N1506, N1501, N952);
not NOT1 (N1507, N1495);
xor XOR2 (N1508, N1497, N1320);
not NOT1 (N1509, N1496);
nor NOR2 (N1510, N1500, N332);
nand NAND2 (N1511, N1507, N948);
xor XOR2 (N1512, N1492, N218);
not NOT1 (N1513, N1512);
not NOT1 (N1514, N1509);
endmodule