// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N721,N719,N712,N709,N720,N710,N716,N711,N702,N722;

not NOT1 (N23, N12);
nand NAND3 (N24, N17, N10, N9);
not NOT1 (N25, N8);
buf BUF1 (N26, N4);
or OR4 (N27, N9, N18, N18, N18);
xor XOR2 (N28, N19, N7);
xor XOR2 (N29, N15, N1);
xor XOR2 (N30, N16, N28);
nand NAND4 (N31, N22, N29, N12, N3);
nand NAND4 (N32, N2, N17, N15, N16);
not NOT1 (N33, N29);
or OR3 (N34, N22, N31, N16);
nor NOR3 (N35, N8, N10, N25);
not NOT1 (N36, N6);
or OR4 (N37, N30, N11, N14, N26);
not NOT1 (N38, N13);
buf BUF1 (N39, N37);
not NOT1 (N40, N23);
nor NOR2 (N41, N38, N37);
nand NAND2 (N42, N32, N21);
or OR2 (N43, N24, N22);
nor NOR2 (N44, N27, N6);
or OR3 (N45, N33, N3, N36);
nor NOR2 (N46, N17, N25);
nor NOR3 (N47, N45, N28, N19);
not NOT1 (N48, N35);
and AND3 (N49, N41, N42, N24);
or OR4 (N50, N45, N22, N6, N24);
nor NOR4 (N51, N48, N50, N9, N34);
nand NAND2 (N52, N42, N10);
or OR3 (N53, N23, N34, N19);
or OR3 (N54, N52, N33, N32);
nor NOR3 (N55, N51, N38, N47);
and AND2 (N56, N24, N29);
or OR4 (N57, N53, N1, N12, N17);
and AND4 (N58, N55, N46, N24, N40);
or OR4 (N59, N3, N34, N48, N37);
not NOT1 (N60, N40);
not NOT1 (N61, N56);
buf BUF1 (N62, N61);
or OR3 (N63, N57, N45, N33);
nand NAND4 (N64, N44, N27, N39, N5);
nor NOR3 (N65, N61, N34, N54);
nand NAND4 (N66, N30, N50, N14, N4);
nor NOR4 (N67, N49, N51, N9, N17);
nand NAND2 (N68, N66, N58);
nand NAND3 (N69, N48, N5, N34);
nor NOR2 (N70, N60, N16);
or OR2 (N71, N67, N39);
and AND3 (N72, N69, N67, N17);
and AND2 (N73, N63, N69);
xor XOR2 (N74, N70, N41);
xor XOR2 (N75, N64, N71);
nor NOR4 (N76, N26, N10, N34, N12);
or OR3 (N77, N43, N2, N56);
xor XOR2 (N78, N72, N62);
buf BUF1 (N79, N32);
nor NOR3 (N80, N74, N43, N28);
nor NOR3 (N81, N80, N61, N31);
buf BUF1 (N82, N75);
nand NAND4 (N83, N78, N72, N70, N22);
nand NAND2 (N84, N79, N2);
not NOT1 (N85, N59);
not NOT1 (N86, N85);
not NOT1 (N87, N86);
nor NOR4 (N88, N82, N45, N85, N5);
or OR3 (N89, N81, N61, N72);
xor XOR2 (N90, N68, N68);
buf BUF1 (N91, N89);
and AND3 (N92, N91, N68, N31);
nor NOR3 (N93, N84, N55, N49);
xor XOR2 (N94, N73, N44);
and AND2 (N95, N88, N15);
xor XOR2 (N96, N65, N84);
buf BUF1 (N97, N76);
not NOT1 (N98, N83);
nor NOR2 (N99, N92, N13);
xor XOR2 (N100, N94, N86);
nor NOR4 (N101, N100, N47, N56, N36);
not NOT1 (N102, N93);
not NOT1 (N103, N95);
and AND2 (N104, N98, N21);
and AND3 (N105, N96, N64, N37);
and AND3 (N106, N104, N68, N21);
not NOT1 (N107, N102);
not NOT1 (N108, N77);
nand NAND4 (N109, N97, N77, N90, N104);
nor NOR2 (N110, N35, N81);
nor NOR3 (N111, N105, N4, N7);
xor XOR2 (N112, N111, N107);
nor NOR2 (N113, N102, N86);
or OR3 (N114, N110, N73, N81);
buf BUF1 (N115, N112);
and AND4 (N116, N115, N100, N38, N104);
and AND2 (N117, N103, N34);
nand NAND3 (N118, N106, N106, N22);
xor XOR2 (N119, N118, N107);
nand NAND4 (N120, N116, N104, N7, N73);
buf BUF1 (N121, N114);
nor NOR4 (N122, N121, N121, N59, N52);
xor XOR2 (N123, N101, N95);
and AND3 (N124, N113, N93, N81);
or OR3 (N125, N108, N77, N48);
or OR2 (N126, N117, N27);
and AND2 (N127, N119, N28);
nand NAND2 (N128, N126, N64);
nand NAND4 (N129, N128, N120, N95, N23);
buf BUF1 (N130, N91);
and AND3 (N131, N99, N130, N51);
or OR2 (N132, N3, N128);
and AND2 (N133, N87, N117);
xor XOR2 (N134, N125, N32);
buf BUF1 (N135, N132);
and AND4 (N136, N135, N67, N115, N48);
and AND4 (N137, N122, N90, N87, N96);
nor NOR3 (N138, N129, N102, N32);
nand NAND4 (N139, N133, N97, N135, N68);
not NOT1 (N140, N131);
and AND2 (N141, N134, N33);
nand NAND4 (N142, N141, N76, N29, N104);
buf BUF1 (N143, N127);
or OR4 (N144, N138, N107, N110, N116);
buf BUF1 (N145, N139);
nand NAND4 (N146, N144, N119, N45, N32);
or OR3 (N147, N142, N119, N23);
xor XOR2 (N148, N124, N85);
buf BUF1 (N149, N146);
nor NOR2 (N150, N136, N79);
or OR3 (N151, N145, N147, N123);
not NOT1 (N152, N76);
nand NAND3 (N153, N19, N100, N118);
or OR2 (N154, N140, N86);
or OR2 (N155, N154, N6);
nand NAND3 (N156, N151, N75, N111);
nor NOR2 (N157, N149, N97);
xor XOR2 (N158, N157, N4);
nor NOR3 (N159, N152, N141, N87);
or OR3 (N160, N153, N146, N10);
not NOT1 (N161, N137);
buf BUF1 (N162, N148);
nand NAND2 (N163, N156, N51);
or OR2 (N164, N158, N3);
and AND2 (N165, N155, N66);
xor XOR2 (N166, N159, N7);
or OR3 (N167, N160, N66, N149);
nand NAND2 (N168, N164, N125);
nor NOR2 (N169, N166, N51);
and AND4 (N170, N165, N38, N121, N25);
nor NOR4 (N171, N161, N163, N4, N80);
or OR3 (N172, N74, N94, N142);
nand NAND3 (N173, N150, N172, N121);
nand NAND2 (N174, N91, N167);
or OR4 (N175, N73, N48, N114, N9);
nand NAND2 (N176, N169, N130);
buf BUF1 (N177, N175);
or OR3 (N178, N174, N136, N172);
and AND3 (N179, N109, N97, N151);
nand NAND2 (N180, N168, N33);
or OR4 (N181, N162, N49, N43, N144);
nand NAND3 (N182, N179, N14, N5);
not NOT1 (N183, N176);
nand NAND2 (N184, N171, N138);
xor XOR2 (N185, N177, N163);
nor NOR4 (N186, N173, N64, N20, N54);
xor XOR2 (N187, N170, N4);
nand NAND4 (N188, N184, N170, N163, N47);
buf BUF1 (N189, N185);
and AND4 (N190, N181, N158, N100, N72);
buf BUF1 (N191, N188);
and AND3 (N192, N182, N158, N134);
nor NOR2 (N193, N143, N108);
nand NAND4 (N194, N187, N184, N171, N185);
buf BUF1 (N195, N178);
xor XOR2 (N196, N191, N63);
buf BUF1 (N197, N186);
nand NAND4 (N198, N197, N187, N146, N57);
nand NAND2 (N199, N190, N64);
and AND2 (N200, N193, N130);
or OR2 (N201, N196, N125);
or OR2 (N202, N195, N186);
and AND2 (N203, N199, N1);
or OR3 (N204, N183, N82, N21);
or OR2 (N205, N189, N167);
or OR2 (N206, N205, N176);
not NOT1 (N207, N206);
or OR3 (N208, N201, N117, N129);
buf BUF1 (N209, N208);
nor NOR4 (N210, N194, N168, N7, N123);
or OR3 (N211, N203, N47, N57);
buf BUF1 (N212, N180);
and AND4 (N213, N204, N184, N198, N186);
xor XOR2 (N214, N66, N18);
and AND4 (N215, N200, N190, N71, N35);
and AND4 (N216, N211, N30, N159, N61);
nand NAND2 (N217, N207, N174);
nor NOR2 (N218, N212, N87);
nor NOR4 (N219, N202, N120, N121, N136);
buf BUF1 (N220, N192);
and AND2 (N221, N217, N117);
nand NAND4 (N222, N221, N25, N160, N203);
xor XOR2 (N223, N219, N99);
not NOT1 (N224, N220);
or OR2 (N225, N210, N2);
not NOT1 (N226, N214);
nor NOR3 (N227, N215, N56, N80);
xor XOR2 (N228, N222, N163);
and AND3 (N229, N228, N201, N81);
not NOT1 (N230, N218);
nand NAND4 (N231, N229, N103, N211, N54);
not NOT1 (N232, N223);
xor XOR2 (N233, N230, N134);
buf BUF1 (N234, N227);
not NOT1 (N235, N216);
nor NOR3 (N236, N233, N56, N62);
buf BUF1 (N237, N224);
nand NAND3 (N238, N237, N195, N71);
xor XOR2 (N239, N235, N132);
nor NOR2 (N240, N209, N107);
nand NAND4 (N241, N236, N175, N167, N158);
not NOT1 (N242, N231);
not NOT1 (N243, N234);
nor NOR4 (N244, N213, N202, N171, N211);
and AND4 (N245, N240, N93, N149, N170);
nand NAND2 (N246, N226, N183);
and AND2 (N247, N245, N159);
nor NOR4 (N248, N246, N114, N238, N209);
and AND2 (N249, N57, N70);
not NOT1 (N250, N244);
nor NOR2 (N251, N248, N84);
not NOT1 (N252, N247);
or OR3 (N253, N225, N113, N153);
nor NOR2 (N254, N242, N100);
or OR3 (N255, N250, N153, N44);
buf BUF1 (N256, N252);
and AND3 (N257, N243, N31, N159);
buf BUF1 (N258, N256);
nor NOR2 (N259, N239, N70);
xor XOR2 (N260, N254, N219);
or OR4 (N261, N251, N186, N8, N184);
nor NOR2 (N262, N260, N240);
xor XOR2 (N263, N261, N199);
not NOT1 (N264, N249);
buf BUF1 (N265, N262);
and AND2 (N266, N257, N205);
buf BUF1 (N267, N255);
not NOT1 (N268, N266);
or OR4 (N269, N232, N43, N228, N194);
nor NOR4 (N270, N269, N166, N199, N177);
nand NAND2 (N271, N258, N212);
or OR3 (N272, N268, N195, N1);
or OR4 (N273, N265, N110, N209, N57);
and AND4 (N274, N259, N191, N240, N55);
xor XOR2 (N275, N253, N4);
nand NAND2 (N276, N274, N61);
nand NAND3 (N277, N275, N157, N88);
nand NAND3 (N278, N264, N186, N4);
or OR4 (N279, N276, N112, N265, N182);
nand NAND2 (N280, N241, N259);
and AND4 (N281, N280, N162, N277, N259);
xor XOR2 (N282, N42, N196);
or OR4 (N283, N273, N129, N175, N159);
not NOT1 (N284, N272);
nor NOR2 (N285, N283, N33);
buf BUF1 (N286, N278);
nor NOR2 (N287, N281, N55);
not NOT1 (N288, N271);
buf BUF1 (N289, N288);
nand NAND4 (N290, N285, N13, N71, N18);
buf BUF1 (N291, N270);
not NOT1 (N292, N284);
not NOT1 (N293, N289);
xor XOR2 (N294, N291, N273);
or OR2 (N295, N293, N139);
nor NOR4 (N296, N282, N79, N167, N272);
nor NOR2 (N297, N294, N114);
or OR3 (N298, N297, N63, N241);
buf BUF1 (N299, N292);
nor NOR2 (N300, N287, N228);
nand NAND3 (N301, N267, N184, N79);
or OR3 (N302, N295, N172, N295);
nor NOR3 (N303, N302, N7, N258);
or OR2 (N304, N296, N166);
buf BUF1 (N305, N301);
nor NOR2 (N306, N304, N170);
nand NAND2 (N307, N298, N10);
nor NOR3 (N308, N306, N64, N265);
buf BUF1 (N309, N290);
buf BUF1 (N310, N286);
buf BUF1 (N311, N309);
buf BUF1 (N312, N311);
xor XOR2 (N313, N263, N45);
nand NAND4 (N314, N307, N206, N205, N267);
not NOT1 (N315, N312);
nor NOR4 (N316, N315, N263, N52, N174);
and AND3 (N317, N316, N177, N36);
buf BUF1 (N318, N299);
or OR2 (N319, N314, N56);
buf BUF1 (N320, N305);
nor NOR2 (N321, N317, N54);
nor NOR3 (N322, N279, N268, N186);
and AND4 (N323, N321, N122, N99, N61);
nand NAND3 (N324, N320, N226, N97);
or OR2 (N325, N300, N39);
or OR3 (N326, N313, N46, N208);
nor NOR3 (N327, N322, N205, N162);
xor XOR2 (N328, N303, N76);
nor NOR3 (N329, N325, N224, N60);
nand NAND2 (N330, N326, N157);
nor NOR4 (N331, N310, N183, N67, N105);
nand NAND4 (N332, N330, N146, N135, N56);
xor XOR2 (N333, N318, N160);
xor XOR2 (N334, N308, N46);
buf BUF1 (N335, N328);
xor XOR2 (N336, N333, N265);
nand NAND3 (N337, N323, N191, N277);
and AND3 (N338, N324, N108, N56);
xor XOR2 (N339, N327, N116);
buf BUF1 (N340, N319);
nor NOR4 (N341, N336, N64, N95, N150);
nor NOR3 (N342, N337, N308, N41);
xor XOR2 (N343, N331, N62);
and AND3 (N344, N341, N229, N135);
xor XOR2 (N345, N329, N37);
nor NOR3 (N346, N334, N262, N111);
buf BUF1 (N347, N345);
or OR2 (N348, N347, N132);
and AND4 (N349, N348, N329, N120, N287);
and AND3 (N350, N335, N239, N119);
buf BUF1 (N351, N340);
nand NAND3 (N352, N339, N250, N80);
buf BUF1 (N353, N351);
or OR2 (N354, N342, N301);
nand NAND2 (N355, N353, N12);
nand NAND3 (N356, N332, N211, N344);
nor NOR3 (N357, N264, N30, N248);
xor XOR2 (N358, N352, N80);
nand NAND2 (N359, N356, N236);
xor XOR2 (N360, N359, N59);
buf BUF1 (N361, N358);
not NOT1 (N362, N360);
not NOT1 (N363, N349);
and AND3 (N364, N355, N54, N183);
buf BUF1 (N365, N338);
nor NOR2 (N366, N365, N108);
nand NAND2 (N367, N346, N238);
xor XOR2 (N368, N367, N301);
or OR3 (N369, N368, N237, N200);
nand NAND3 (N370, N357, N227, N36);
xor XOR2 (N371, N362, N272);
nor NOR4 (N372, N371, N203, N167, N59);
xor XOR2 (N373, N364, N289);
xor XOR2 (N374, N354, N278);
or OR2 (N375, N343, N45);
not NOT1 (N376, N366);
xor XOR2 (N377, N370, N374);
and AND2 (N378, N334, N246);
nor NOR4 (N379, N376, N220, N30, N191);
xor XOR2 (N380, N363, N101);
not NOT1 (N381, N369);
xor XOR2 (N382, N377, N308);
buf BUF1 (N383, N381);
xor XOR2 (N384, N379, N134);
or OR3 (N385, N373, N163, N14);
and AND3 (N386, N350, N17, N57);
buf BUF1 (N387, N361);
nand NAND3 (N388, N385, N296, N172);
nand NAND3 (N389, N375, N4, N303);
or OR3 (N390, N388, N269, N210);
nand NAND3 (N391, N390, N100, N105);
xor XOR2 (N392, N387, N181);
and AND4 (N393, N383, N262, N243, N250);
nand NAND4 (N394, N378, N239, N312, N177);
nor NOR2 (N395, N394, N9);
not NOT1 (N396, N389);
buf BUF1 (N397, N384);
xor XOR2 (N398, N395, N286);
nand NAND2 (N399, N380, N84);
nor NOR4 (N400, N391, N357, N10, N292);
buf BUF1 (N401, N396);
not NOT1 (N402, N392);
xor XOR2 (N403, N372, N176);
not NOT1 (N404, N393);
and AND3 (N405, N401, N216, N108);
nand NAND4 (N406, N403, N287, N26, N130);
and AND4 (N407, N402, N218, N380, N212);
and AND2 (N408, N397, N130);
nand NAND3 (N409, N406, N192, N34);
or OR2 (N410, N400, N108);
not NOT1 (N411, N407);
buf BUF1 (N412, N399);
and AND2 (N413, N398, N45);
and AND2 (N414, N413, N388);
nand NAND2 (N415, N405, N265);
or OR3 (N416, N412, N147, N58);
buf BUF1 (N417, N415);
not NOT1 (N418, N386);
or OR2 (N419, N382, N222);
or OR3 (N420, N416, N318, N382);
xor XOR2 (N421, N404, N370);
nor NOR3 (N422, N410, N64, N200);
nand NAND3 (N423, N422, N390, N131);
nand NAND2 (N424, N417, N308);
buf BUF1 (N425, N409);
buf BUF1 (N426, N414);
buf BUF1 (N427, N411);
buf BUF1 (N428, N408);
not NOT1 (N429, N427);
nand NAND2 (N430, N421, N381);
not NOT1 (N431, N424);
and AND2 (N432, N419, N53);
nand NAND3 (N433, N428, N416, N61);
buf BUF1 (N434, N429);
xor XOR2 (N435, N433, N350);
buf BUF1 (N436, N425);
buf BUF1 (N437, N434);
and AND4 (N438, N436, N30, N415, N353);
buf BUF1 (N439, N435);
nor NOR4 (N440, N430, N393, N313, N200);
not NOT1 (N441, N432);
and AND3 (N442, N431, N70, N103);
xor XOR2 (N443, N439, N28);
nor NOR3 (N444, N442, N165, N71);
not NOT1 (N445, N437);
or OR2 (N446, N443, N290);
xor XOR2 (N447, N423, N192);
or OR2 (N448, N418, N340);
not NOT1 (N449, N426);
buf BUF1 (N450, N449);
or OR4 (N451, N441, N79, N226, N117);
not NOT1 (N452, N445);
and AND4 (N453, N420, N292, N278, N290);
and AND2 (N454, N440, N407);
not NOT1 (N455, N438);
nor NOR2 (N456, N452, N287);
or OR2 (N457, N444, N430);
xor XOR2 (N458, N456, N442);
nor NOR4 (N459, N458, N241, N127, N353);
and AND3 (N460, N457, N222, N239);
or OR2 (N461, N451, N283);
not NOT1 (N462, N446);
not NOT1 (N463, N460);
not NOT1 (N464, N447);
xor XOR2 (N465, N448, N459);
not NOT1 (N466, N150);
not NOT1 (N467, N462);
or OR4 (N468, N467, N106, N208, N57);
or OR3 (N469, N464, N456, N341);
nand NAND3 (N470, N450, N114, N4);
and AND2 (N471, N469, N78);
nand NAND3 (N472, N461, N245, N16);
and AND2 (N473, N455, N454);
not NOT1 (N474, N155);
or OR2 (N475, N474, N257);
buf BUF1 (N476, N475);
buf BUF1 (N477, N471);
nand NAND2 (N478, N465, N174);
or OR2 (N479, N473, N27);
and AND2 (N480, N478, N328);
or OR3 (N481, N468, N68, N174);
and AND4 (N482, N479, N380, N358, N475);
xor XOR2 (N483, N453, N97);
buf BUF1 (N484, N463);
nand NAND2 (N485, N470, N17);
nand NAND4 (N486, N483, N382, N348, N465);
xor XOR2 (N487, N480, N87);
and AND3 (N488, N484, N150, N206);
xor XOR2 (N489, N488, N337);
and AND4 (N490, N472, N277, N198, N278);
nand NAND2 (N491, N485, N279);
and AND4 (N492, N482, N416, N52, N443);
xor XOR2 (N493, N476, N448);
not NOT1 (N494, N491);
nor NOR3 (N495, N489, N5, N222);
nand NAND2 (N496, N487, N366);
buf BUF1 (N497, N496);
nand NAND4 (N498, N492, N168, N1, N326);
or OR3 (N499, N493, N211, N327);
and AND3 (N500, N499, N44, N386);
buf BUF1 (N501, N481);
xor XOR2 (N502, N486, N189);
xor XOR2 (N503, N490, N214);
or OR3 (N504, N497, N317, N89);
nor NOR2 (N505, N466, N459);
or OR4 (N506, N477, N362, N160, N59);
or OR3 (N507, N501, N480, N306);
nor NOR3 (N508, N506, N468, N11);
or OR2 (N509, N505, N326);
and AND2 (N510, N504, N426);
not NOT1 (N511, N509);
buf BUF1 (N512, N503);
or OR3 (N513, N508, N261, N274);
nor NOR2 (N514, N500, N252);
and AND4 (N515, N512, N435, N304, N103);
not NOT1 (N516, N513);
or OR2 (N517, N510, N329);
and AND2 (N518, N511, N254);
xor XOR2 (N519, N502, N252);
not NOT1 (N520, N494);
buf BUF1 (N521, N518);
or OR2 (N522, N521, N56);
and AND3 (N523, N520, N261, N243);
not NOT1 (N524, N517);
and AND4 (N525, N523, N353, N51, N331);
or OR4 (N526, N524, N234, N363, N81);
buf BUF1 (N527, N495);
nor NOR4 (N528, N522, N402, N206, N464);
nand NAND2 (N529, N528, N412);
xor XOR2 (N530, N519, N471);
buf BUF1 (N531, N514);
nor NOR2 (N532, N525, N457);
nor NOR3 (N533, N530, N102, N62);
nand NAND4 (N534, N533, N447, N233, N77);
not NOT1 (N535, N515);
not NOT1 (N536, N527);
xor XOR2 (N537, N532, N498);
or OR2 (N538, N76, N522);
not NOT1 (N539, N537);
buf BUF1 (N540, N538);
buf BUF1 (N541, N534);
nand NAND3 (N542, N531, N26, N143);
or OR3 (N543, N540, N465, N333);
nor NOR2 (N544, N507, N179);
nand NAND2 (N545, N526, N298);
xor XOR2 (N546, N544, N222);
buf BUF1 (N547, N546);
xor XOR2 (N548, N535, N101);
xor XOR2 (N549, N547, N228);
not NOT1 (N550, N548);
and AND3 (N551, N545, N158, N79);
xor XOR2 (N552, N551, N393);
buf BUF1 (N553, N542);
not NOT1 (N554, N516);
xor XOR2 (N555, N543, N136);
and AND3 (N556, N541, N273, N524);
buf BUF1 (N557, N556);
xor XOR2 (N558, N536, N358);
and AND2 (N559, N550, N501);
and AND4 (N560, N552, N535, N331, N483);
xor XOR2 (N561, N560, N139);
not NOT1 (N562, N558);
and AND4 (N563, N554, N23, N441, N12);
or OR3 (N564, N561, N371, N118);
not NOT1 (N565, N529);
and AND4 (N566, N559, N149, N283, N463);
or OR2 (N567, N539, N563);
xor XOR2 (N568, N18, N145);
not NOT1 (N569, N565);
xor XOR2 (N570, N568, N118);
nor NOR2 (N571, N553, N63);
or OR4 (N572, N566, N122, N328, N203);
or OR3 (N573, N567, N424, N207);
xor XOR2 (N574, N571, N389);
xor XOR2 (N575, N549, N549);
not NOT1 (N576, N573);
xor XOR2 (N577, N562, N413);
and AND3 (N578, N570, N358, N477);
buf BUF1 (N579, N572);
nand NAND3 (N580, N576, N479, N293);
not NOT1 (N581, N579);
buf BUF1 (N582, N557);
xor XOR2 (N583, N577, N117);
not NOT1 (N584, N583);
xor XOR2 (N585, N582, N16);
and AND3 (N586, N581, N78, N153);
nor NOR4 (N587, N564, N263, N74, N25);
and AND4 (N588, N580, N338, N370, N524);
xor XOR2 (N589, N584, N221);
nand NAND3 (N590, N586, N88, N90);
nand NAND2 (N591, N590, N315);
nor NOR3 (N592, N574, N345, N175);
not NOT1 (N593, N578);
nor NOR3 (N594, N555, N592, N209);
and AND2 (N595, N256, N458);
not NOT1 (N596, N593);
or OR2 (N597, N596, N515);
nor NOR4 (N598, N569, N406, N579, N568);
not NOT1 (N599, N575);
not NOT1 (N600, N585);
or OR2 (N601, N600, N218);
not NOT1 (N602, N595);
xor XOR2 (N603, N594, N561);
nand NAND4 (N604, N601, N90, N140, N414);
not NOT1 (N605, N588);
buf BUF1 (N606, N604);
buf BUF1 (N607, N603);
nand NAND3 (N608, N607, N304, N516);
or OR2 (N609, N608, N374);
not NOT1 (N610, N606);
not NOT1 (N611, N609);
not NOT1 (N612, N591);
nor NOR4 (N613, N605, N103, N449, N108);
nor NOR2 (N614, N613, N507);
buf BUF1 (N615, N598);
not NOT1 (N616, N615);
or OR2 (N617, N611, N149);
and AND4 (N618, N610, N138, N152, N153);
or OR4 (N619, N597, N42, N503, N517);
not NOT1 (N620, N619);
or OR3 (N621, N589, N278, N170);
not NOT1 (N622, N599);
buf BUF1 (N623, N621);
and AND4 (N624, N602, N136, N597, N235);
not NOT1 (N625, N612);
buf BUF1 (N626, N587);
xor XOR2 (N627, N620, N502);
not NOT1 (N628, N618);
buf BUF1 (N629, N626);
and AND4 (N630, N628, N204, N205, N453);
not NOT1 (N631, N623);
buf BUF1 (N632, N624);
nor NOR4 (N633, N630, N355, N61, N533);
or OR4 (N634, N614, N172, N497, N242);
or OR4 (N635, N634, N387, N432, N64);
and AND4 (N636, N629, N52, N371, N31);
and AND2 (N637, N616, N515);
nor NOR2 (N638, N622, N385);
or OR3 (N639, N627, N234, N613);
not NOT1 (N640, N637);
not NOT1 (N641, N631);
nor NOR4 (N642, N632, N219, N138, N304);
or OR4 (N643, N636, N149, N509, N249);
buf BUF1 (N644, N638);
nand NAND4 (N645, N641, N415, N526, N554);
buf BUF1 (N646, N644);
and AND4 (N647, N642, N69, N138, N217);
nor NOR4 (N648, N643, N515, N174, N276);
not NOT1 (N649, N625);
and AND3 (N650, N646, N464, N531);
or OR4 (N651, N649, N550, N380, N430);
xor XOR2 (N652, N635, N242);
and AND2 (N653, N639, N564);
buf BUF1 (N654, N648);
buf BUF1 (N655, N652);
or OR4 (N656, N645, N361, N442, N475);
nor NOR2 (N657, N640, N310);
xor XOR2 (N658, N656, N336);
not NOT1 (N659, N633);
xor XOR2 (N660, N658, N261);
or OR2 (N661, N653, N564);
nand NAND3 (N662, N617, N255, N582);
and AND2 (N663, N651, N124);
not NOT1 (N664, N647);
not NOT1 (N665, N662);
xor XOR2 (N666, N657, N481);
or OR2 (N667, N660, N483);
and AND3 (N668, N655, N519, N585);
xor XOR2 (N669, N650, N490);
buf BUF1 (N670, N665);
buf BUF1 (N671, N659);
buf BUF1 (N672, N669);
not NOT1 (N673, N668);
not NOT1 (N674, N661);
xor XOR2 (N675, N654, N162);
or OR2 (N676, N674, N207);
not NOT1 (N677, N673);
not NOT1 (N678, N664);
xor XOR2 (N679, N667, N97);
xor XOR2 (N680, N666, N86);
buf BUF1 (N681, N680);
nor NOR4 (N682, N678, N341, N256, N330);
xor XOR2 (N683, N675, N618);
and AND3 (N684, N681, N407, N30);
buf BUF1 (N685, N672);
not NOT1 (N686, N671);
not NOT1 (N687, N679);
nor NOR4 (N688, N686, N402, N594, N627);
not NOT1 (N689, N685);
not NOT1 (N690, N688);
buf BUF1 (N691, N687);
buf BUF1 (N692, N663);
nor NOR2 (N693, N676, N159);
or OR2 (N694, N692, N382);
buf BUF1 (N695, N684);
nor NOR4 (N696, N689, N122, N230, N641);
nand NAND3 (N697, N696, N414, N591);
and AND3 (N698, N694, N239, N549);
or OR2 (N699, N670, N263);
or OR3 (N700, N691, N412, N42);
nor NOR2 (N701, N683, N433);
nand NAND4 (N702, N677, N33, N487, N201);
nand NAND3 (N703, N698, N374, N66);
or OR2 (N704, N695, N267);
buf BUF1 (N705, N701);
and AND2 (N706, N682, N640);
or OR4 (N707, N703, N400, N636, N29);
or OR3 (N708, N707, N319, N707);
or OR4 (N709, N693, N70, N468, N101);
nand NAND2 (N710, N700, N228);
and AND2 (N711, N705, N268);
and AND4 (N712, N708, N85, N292, N240);
nor NOR2 (N713, N690, N549);
and AND4 (N714, N699, N346, N12, N238);
nand NAND2 (N715, N704, N58);
nand NAND3 (N716, N706, N299, N29);
and AND4 (N717, N713, N200, N340, N488);
not NOT1 (N718, N715);
and AND4 (N719, N714, N220, N364, N465);
buf BUF1 (N720, N697);
and AND4 (N721, N718, N649, N56, N290);
nand NAND4 (N722, N717, N660, N674, N201);
endmodule