// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N3219,N3220,N3214,N3197,N3188,N3211,N3213,N3222,N3210,N3223;

xor XOR2 (N24, N23, N15);
nand NAND3 (N25, N8, N24, N4);
xor XOR2 (N26, N11, N2);
nand NAND2 (N27, N22, N4);
or OR2 (N28, N12, N21);
and AND4 (N29, N23, N16, N26, N25);
and AND2 (N30, N1, N23);
xor XOR2 (N31, N2, N6);
nand NAND4 (N32, N16, N16, N10, N4);
nor NOR4 (N33, N3, N27, N5, N11);
nor NOR2 (N34, N10, N8);
and AND2 (N35, N24, N21);
not NOT1 (N36, N18);
not NOT1 (N37, N6);
and AND3 (N38, N32, N7, N26);
xor XOR2 (N39, N28, N24);
or OR2 (N40, N38, N3);
nor NOR4 (N41, N29, N13, N10, N25);
xor XOR2 (N42, N30, N32);
buf BUF1 (N43, N34);
nor NOR4 (N44, N36, N7, N7, N31);
or OR3 (N45, N11, N34, N17);
nor NOR4 (N46, N33, N23, N5, N29);
nor NOR2 (N47, N45, N32);
xor XOR2 (N48, N47, N26);
xor XOR2 (N49, N48, N25);
or OR3 (N50, N46, N33, N5);
nand NAND2 (N51, N41, N36);
or OR3 (N52, N44, N47, N35);
and AND2 (N53, N9, N4);
xor XOR2 (N54, N49, N50);
or OR3 (N55, N6, N17, N11);
not NOT1 (N56, N52);
nor NOR3 (N57, N42, N18, N4);
nor NOR3 (N58, N55, N6, N20);
not NOT1 (N59, N37);
nor NOR3 (N60, N59, N36, N1);
not NOT1 (N61, N53);
buf BUF1 (N62, N43);
nor NOR3 (N63, N51, N23, N38);
not NOT1 (N64, N60);
nand NAND4 (N65, N40, N24, N17, N32);
and AND2 (N66, N64, N5);
xor XOR2 (N67, N61, N65);
nand NAND4 (N68, N13, N51, N44, N59);
nand NAND3 (N69, N57, N26, N16);
and AND2 (N70, N39, N13);
nand NAND4 (N71, N62, N13, N67, N20);
not NOT1 (N72, N17);
xor XOR2 (N73, N70, N60);
xor XOR2 (N74, N56, N71);
xor XOR2 (N75, N41, N45);
buf BUF1 (N76, N73);
buf BUF1 (N77, N66);
not NOT1 (N78, N58);
and AND3 (N79, N77, N23, N72);
or OR4 (N80, N44, N2, N37, N12);
nand NAND3 (N81, N76, N2, N10);
not NOT1 (N82, N63);
buf BUF1 (N83, N54);
xor XOR2 (N84, N80, N68);
nand NAND4 (N85, N15, N24, N1, N11);
or OR2 (N86, N81, N70);
and AND3 (N87, N75, N47, N23);
and AND2 (N88, N82, N70);
or OR4 (N89, N79, N21, N46, N54);
xor XOR2 (N90, N84, N55);
and AND3 (N91, N90, N30, N9);
xor XOR2 (N92, N74, N90);
not NOT1 (N93, N86);
nand NAND3 (N94, N92, N9, N66);
or OR4 (N95, N89, N67, N89, N80);
or OR3 (N96, N93, N12, N43);
nand NAND4 (N97, N88, N11, N81, N54);
and AND4 (N98, N69, N97, N9, N40);
buf BUF1 (N99, N48);
xor XOR2 (N100, N94, N95);
and AND3 (N101, N54, N26, N49);
buf BUF1 (N102, N99);
buf BUF1 (N103, N91);
and AND4 (N104, N102, N74, N22, N32);
xor XOR2 (N105, N100, N23);
buf BUF1 (N106, N105);
or OR2 (N107, N101, N9);
buf BUF1 (N108, N107);
and AND3 (N109, N78, N72, N62);
nor NOR2 (N110, N104, N87);
not NOT1 (N111, N96);
and AND2 (N112, N89, N103);
or OR4 (N113, N49, N33, N17, N13);
nor NOR4 (N114, N112, N46, N80, N105);
nor NOR2 (N115, N83, N68);
xor XOR2 (N116, N113, N49);
xor XOR2 (N117, N85, N22);
xor XOR2 (N118, N116, N96);
buf BUF1 (N119, N106);
buf BUF1 (N120, N109);
nor NOR3 (N121, N111, N36, N72);
buf BUF1 (N122, N115);
nand NAND4 (N123, N117, N115, N14, N59);
nor NOR2 (N124, N108, N1);
nand NAND3 (N125, N118, N100, N108);
or OR3 (N126, N124, N7, N104);
buf BUF1 (N127, N120);
buf BUF1 (N128, N125);
not NOT1 (N129, N127);
nand NAND4 (N130, N110, N105, N94, N11);
nor NOR3 (N131, N121, N77, N64);
buf BUF1 (N132, N131);
nand NAND4 (N133, N123, N3, N23, N104);
buf BUF1 (N134, N133);
or OR4 (N135, N126, N109, N42, N17);
buf BUF1 (N136, N98);
nor NOR2 (N137, N128, N4);
or OR3 (N138, N114, N54, N100);
nand NAND2 (N139, N134, N10);
xor XOR2 (N140, N139, N105);
xor XOR2 (N141, N138, N5);
buf BUF1 (N142, N135);
buf BUF1 (N143, N129);
and AND4 (N144, N130, N72, N85, N86);
xor XOR2 (N145, N141, N105);
buf BUF1 (N146, N136);
nand NAND3 (N147, N145, N143, N66);
or OR4 (N148, N122, N94, N104, N109);
nand NAND4 (N149, N8, N42, N128, N82);
xor XOR2 (N150, N147, N128);
and AND4 (N151, N140, N36, N111, N134);
buf BUF1 (N152, N137);
or OR3 (N153, N148, N19, N7);
xor XOR2 (N154, N152, N71);
nor NOR2 (N155, N146, N68);
nand NAND3 (N156, N132, N99, N123);
nand NAND3 (N157, N149, N124, N129);
not NOT1 (N158, N155);
and AND4 (N159, N153, N96, N75, N43);
buf BUF1 (N160, N150);
xor XOR2 (N161, N154, N98);
or OR3 (N162, N157, N143, N87);
nor NOR2 (N163, N119, N157);
buf BUF1 (N164, N142);
nor NOR3 (N165, N151, N47, N133);
or OR4 (N166, N159, N32, N143, N98);
or OR2 (N167, N164, N165);
buf BUF1 (N168, N56);
buf BUF1 (N169, N163);
not NOT1 (N170, N169);
not NOT1 (N171, N144);
nand NAND3 (N172, N162, N24, N61);
not NOT1 (N173, N172);
or OR4 (N174, N166, N9, N152, N32);
not NOT1 (N175, N167);
nand NAND4 (N176, N171, N110, N161, N52);
buf BUF1 (N177, N44);
nor NOR4 (N178, N176, N62, N77, N96);
and AND3 (N179, N173, N158, N165);
nand NAND3 (N180, N140, N61, N14);
and AND4 (N181, N180, N18, N30, N127);
nor NOR3 (N182, N156, N121, N138);
and AND3 (N183, N168, N173, N180);
nand NAND2 (N184, N160, N144);
or OR2 (N185, N179, N117);
xor XOR2 (N186, N183, N113);
and AND4 (N187, N174, N12, N78, N31);
not NOT1 (N188, N175);
buf BUF1 (N189, N188);
xor XOR2 (N190, N184, N69);
nand NAND4 (N191, N189, N16, N137, N159);
nand NAND2 (N192, N181, N160);
buf BUF1 (N193, N187);
nand NAND4 (N194, N191, N117, N57, N138);
or OR2 (N195, N194, N77);
nand NAND4 (N196, N193, N17, N19, N95);
and AND4 (N197, N192, N87, N91, N51);
nand NAND2 (N198, N190, N195);
and AND4 (N199, N45, N167, N164, N47);
and AND3 (N200, N198, N120, N63);
xor XOR2 (N201, N170, N91);
nand NAND4 (N202, N186, N170, N29, N66);
not NOT1 (N203, N196);
buf BUF1 (N204, N202);
nand NAND3 (N205, N204, N58, N41);
xor XOR2 (N206, N178, N143);
nor NOR4 (N207, N200, N123, N121, N170);
or OR4 (N208, N205, N23, N137, N201);
or OR4 (N209, N196, N183, N113, N29);
buf BUF1 (N210, N208);
not NOT1 (N211, N206);
or OR2 (N212, N197, N178);
buf BUF1 (N213, N182);
not NOT1 (N214, N211);
nor NOR3 (N215, N207, N7, N174);
and AND3 (N216, N199, N150, N107);
buf BUF1 (N217, N203);
xor XOR2 (N218, N216, N191);
or OR3 (N219, N212, N152, N195);
xor XOR2 (N220, N213, N94);
or OR2 (N221, N210, N81);
nor NOR3 (N222, N217, N77, N11);
nand NAND4 (N223, N215, N158, N183, N50);
nand NAND4 (N224, N214, N48, N214, N47);
buf BUF1 (N225, N224);
not NOT1 (N226, N225);
nand NAND4 (N227, N226, N164, N184, N16);
buf BUF1 (N228, N177);
xor XOR2 (N229, N220, N128);
or OR3 (N230, N219, N203, N22);
buf BUF1 (N231, N221);
nand NAND3 (N232, N231, N18, N31);
not NOT1 (N233, N232);
not NOT1 (N234, N218);
xor XOR2 (N235, N228, N115);
not NOT1 (N236, N227);
not NOT1 (N237, N185);
buf BUF1 (N238, N223);
nand NAND3 (N239, N222, N226, N132);
xor XOR2 (N240, N236, N232);
nand NAND3 (N241, N229, N52, N233);
xor XOR2 (N242, N138, N46);
or OR3 (N243, N242, N219, N153);
and AND2 (N244, N209, N184);
nor NOR3 (N245, N234, N172, N180);
or OR3 (N246, N243, N124, N92);
not NOT1 (N247, N237);
not NOT1 (N248, N244);
not NOT1 (N249, N245);
nand NAND2 (N250, N248, N103);
xor XOR2 (N251, N247, N184);
nor NOR2 (N252, N249, N231);
xor XOR2 (N253, N250, N188);
nand NAND3 (N254, N238, N139, N12);
xor XOR2 (N255, N230, N221);
xor XOR2 (N256, N254, N227);
nand NAND3 (N257, N240, N35, N32);
xor XOR2 (N258, N246, N206);
buf BUF1 (N259, N251);
nor NOR4 (N260, N257, N124, N227, N258);
nor NOR4 (N261, N120, N198, N23, N121);
not NOT1 (N262, N259);
or OR4 (N263, N260, N63, N126, N42);
or OR3 (N264, N235, N62, N27);
not NOT1 (N265, N256);
xor XOR2 (N266, N241, N257);
nor NOR2 (N267, N255, N114);
and AND3 (N268, N263, N55, N90);
xor XOR2 (N269, N267, N187);
nand NAND4 (N270, N252, N247, N68, N217);
nor NOR3 (N271, N266, N30, N189);
xor XOR2 (N272, N239, N53);
buf BUF1 (N273, N270);
or OR4 (N274, N261, N54, N8, N206);
nor NOR2 (N275, N272, N246);
or OR4 (N276, N273, N256, N239, N38);
buf BUF1 (N277, N269);
buf BUF1 (N278, N276);
buf BUF1 (N279, N271);
nor NOR4 (N280, N262, N167, N47, N199);
buf BUF1 (N281, N264);
nand NAND4 (N282, N268, N34, N255, N4);
not NOT1 (N283, N253);
not NOT1 (N284, N265);
and AND4 (N285, N283, N146, N103, N179);
buf BUF1 (N286, N277);
and AND4 (N287, N278, N130, N279, N235);
nand NAND3 (N288, N43, N127, N111);
and AND2 (N289, N280, N121);
nand NAND4 (N290, N289, N163, N38, N277);
or OR3 (N291, N275, N227, N287);
nor NOR3 (N292, N67, N128, N87);
buf BUF1 (N293, N291);
not NOT1 (N294, N281);
xor XOR2 (N295, N293, N218);
and AND4 (N296, N290, N209, N87, N247);
and AND4 (N297, N288, N121, N57, N198);
buf BUF1 (N298, N296);
nor NOR4 (N299, N282, N265, N217, N106);
or OR3 (N300, N286, N107, N262);
not NOT1 (N301, N300);
or OR4 (N302, N299, N81, N11, N287);
nand NAND4 (N303, N295, N31, N4, N120);
buf BUF1 (N304, N297);
or OR3 (N305, N274, N100, N10);
nand NAND4 (N306, N294, N293, N214, N205);
or OR2 (N307, N306, N11);
or OR3 (N308, N298, N307, N227);
xor XOR2 (N309, N278, N10);
and AND2 (N310, N285, N82);
nand NAND4 (N311, N304, N309, N253, N147);
nor NOR2 (N312, N269, N74);
not NOT1 (N313, N311);
nand NAND3 (N314, N301, N245, N251);
buf BUF1 (N315, N305);
and AND2 (N316, N310, N102);
nor NOR3 (N317, N303, N280, N239);
not NOT1 (N318, N313);
xor XOR2 (N319, N316, N20);
nand NAND2 (N320, N308, N187);
or OR2 (N321, N318, N252);
xor XOR2 (N322, N317, N216);
not NOT1 (N323, N315);
or OR3 (N324, N292, N183, N204);
nand NAND4 (N325, N312, N175, N88, N234);
or OR3 (N326, N314, N131, N256);
or OR4 (N327, N284, N105, N299, N187);
xor XOR2 (N328, N324, N314);
buf BUF1 (N329, N327);
and AND4 (N330, N329, N228, N93, N76);
and AND4 (N331, N302, N5, N262, N103);
nand NAND4 (N332, N330, N158, N229, N57);
or OR2 (N333, N328, N29);
or OR2 (N334, N326, N205);
xor XOR2 (N335, N322, N97);
buf BUF1 (N336, N335);
or OR4 (N337, N336, N64, N72, N77);
buf BUF1 (N338, N319);
nand NAND2 (N339, N325, N66);
nand NAND2 (N340, N337, N248);
buf BUF1 (N341, N323);
and AND4 (N342, N321, N306, N91, N295);
and AND3 (N343, N334, N171, N12);
or OR2 (N344, N342, N280);
nand NAND2 (N345, N332, N267);
not NOT1 (N346, N338);
buf BUF1 (N347, N331);
nand NAND2 (N348, N339, N32);
and AND2 (N349, N320, N39);
nor NOR4 (N350, N341, N215, N261, N103);
or OR2 (N351, N346, N142);
not NOT1 (N352, N347);
buf BUF1 (N353, N333);
or OR4 (N354, N349, N64, N267, N193);
or OR3 (N355, N352, N149, N147);
buf BUF1 (N356, N355);
nor NOR3 (N357, N344, N168, N297);
and AND4 (N358, N350, N145, N218, N286);
buf BUF1 (N359, N356);
not NOT1 (N360, N359);
not NOT1 (N361, N340);
not NOT1 (N362, N358);
not NOT1 (N363, N357);
not NOT1 (N364, N363);
and AND4 (N365, N354, N77, N331, N331);
or OR2 (N366, N361, N75);
buf BUF1 (N367, N348);
nor NOR2 (N368, N351, N293);
and AND4 (N369, N366, N363, N351, N201);
nor NOR3 (N370, N353, N204, N222);
or OR2 (N371, N362, N82);
or OR3 (N372, N367, N93, N201);
or OR3 (N373, N368, N55, N130);
nor NOR4 (N374, N343, N371, N319, N265);
xor XOR2 (N375, N178, N157);
nand NAND4 (N376, N360, N287, N306, N190);
or OR3 (N377, N370, N173, N107);
xor XOR2 (N378, N375, N366);
nor NOR4 (N379, N364, N318, N255, N20);
or OR2 (N380, N378, N194);
nand NAND4 (N381, N369, N376, N266, N125);
nand NAND3 (N382, N40, N98, N86);
or OR2 (N383, N379, N232);
and AND4 (N384, N380, N67, N274, N292);
or OR4 (N385, N373, N158, N384, N241);
and AND2 (N386, N48, N371);
nand NAND2 (N387, N374, N5);
nor NOR2 (N388, N383, N151);
buf BUF1 (N389, N345);
xor XOR2 (N390, N372, N190);
buf BUF1 (N391, N389);
not NOT1 (N392, N390);
buf BUF1 (N393, N365);
nor NOR2 (N394, N381, N363);
nor NOR2 (N395, N382, N124);
or OR4 (N396, N394, N258, N54, N21);
and AND3 (N397, N386, N291, N45);
nand NAND2 (N398, N393, N203);
buf BUF1 (N399, N398);
and AND2 (N400, N395, N165);
or OR3 (N401, N397, N276, N202);
not NOT1 (N402, N399);
or OR4 (N403, N401, N333, N166, N233);
nand NAND3 (N404, N391, N308, N374);
not NOT1 (N405, N404);
and AND2 (N406, N377, N81);
not NOT1 (N407, N400);
nand NAND3 (N408, N396, N289, N19);
buf BUF1 (N409, N407);
nor NOR2 (N410, N387, N166);
not NOT1 (N411, N409);
xor XOR2 (N412, N385, N314);
and AND2 (N413, N412, N268);
xor XOR2 (N414, N402, N38);
buf BUF1 (N415, N403);
and AND2 (N416, N413, N74);
xor XOR2 (N417, N414, N271);
xor XOR2 (N418, N416, N255);
buf BUF1 (N419, N417);
nand NAND2 (N420, N392, N270);
nand NAND4 (N421, N405, N58, N195, N399);
or OR4 (N422, N411, N72, N313, N297);
not NOT1 (N423, N406);
xor XOR2 (N424, N419, N382);
buf BUF1 (N425, N421);
not NOT1 (N426, N415);
xor XOR2 (N427, N426, N189);
or OR4 (N428, N422, N333, N3, N57);
and AND4 (N429, N418, N45, N376, N314);
nor NOR4 (N430, N410, N128, N258, N281);
not NOT1 (N431, N424);
nand NAND3 (N432, N408, N354, N273);
nor NOR2 (N433, N420, N213);
xor XOR2 (N434, N427, N378);
buf BUF1 (N435, N432);
xor XOR2 (N436, N435, N289);
buf BUF1 (N437, N388);
nor NOR4 (N438, N428, N236, N433, N217);
nor NOR2 (N439, N346, N205);
or OR3 (N440, N438, N260, N67);
nor NOR3 (N441, N440, N39, N234);
and AND3 (N442, N434, N86, N50);
xor XOR2 (N443, N436, N222);
buf BUF1 (N444, N441);
or OR3 (N445, N439, N391, N72);
nor NOR4 (N446, N437, N284, N38, N229);
buf BUF1 (N447, N425);
buf BUF1 (N448, N442);
xor XOR2 (N449, N430, N121);
buf BUF1 (N450, N446);
nand NAND4 (N451, N450, N44, N257, N393);
nor NOR2 (N452, N447, N396);
or OR3 (N453, N452, N174, N427);
nor NOR3 (N454, N423, N333, N282);
or OR4 (N455, N448, N247, N337, N264);
xor XOR2 (N456, N431, N249);
buf BUF1 (N457, N429);
nand NAND3 (N458, N456, N18, N115);
buf BUF1 (N459, N451);
not NOT1 (N460, N444);
or OR2 (N461, N459, N1);
or OR3 (N462, N449, N187, N226);
buf BUF1 (N463, N461);
nand NAND2 (N464, N454, N276);
nand NAND3 (N465, N457, N175, N278);
buf BUF1 (N466, N453);
nand NAND3 (N467, N460, N16, N376);
xor XOR2 (N468, N467, N163);
nor NOR2 (N469, N462, N345);
not NOT1 (N470, N463);
or OR2 (N471, N468, N190);
and AND2 (N472, N470, N131);
or OR2 (N473, N443, N293);
buf BUF1 (N474, N469);
or OR4 (N475, N474, N61, N74, N349);
xor XOR2 (N476, N458, N297);
xor XOR2 (N477, N466, N259);
xor XOR2 (N478, N472, N126);
xor XOR2 (N479, N471, N181);
nand NAND4 (N480, N465, N381, N315, N122);
nor NOR4 (N481, N477, N96, N4, N429);
xor XOR2 (N482, N473, N391);
buf BUF1 (N483, N480);
buf BUF1 (N484, N476);
buf BUF1 (N485, N479);
xor XOR2 (N486, N478, N96);
xor XOR2 (N487, N482, N142);
nor NOR2 (N488, N485, N339);
xor XOR2 (N489, N487, N152);
and AND2 (N490, N475, N91);
and AND3 (N491, N455, N186, N229);
nor NOR2 (N492, N481, N489);
buf BUF1 (N493, N21);
nand NAND4 (N494, N490, N430, N438, N24);
not NOT1 (N495, N493);
nor NOR4 (N496, N488, N192, N471, N301);
nand NAND2 (N497, N486, N348);
and AND3 (N498, N494, N403, N207);
or OR2 (N499, N483, N257);
not NOT1 (N500, N445);
xor XOR2 (N501, N495, N1);
or OR3 (N502, N500, N26, N421);
nor NOR2 (N503, N499, N52);
or OR4 (N504, N491, N78, N405, N97);
xor XOR2 (N505, N501, N47);
buf BUF1 (N506, N502);
and AND4 (N507, N498, N26, N5, N400);
nor NOR2 (N508, N492, N83);
buf BUF1 (N509, N484);
xor XOR2 (N510, N506, N457);
not NOT1 (N511, N464);
or OR3 (N512, N507, N508, N162);
buf BUF1 (N513, N258);
not NOT1 (N514, N504);
not NOT1 (N515, N512);
and AND2 (N516, N497, N314);
xor XOR2 (N517, N513, N132);
nor NOR4 (N518, N517, N300, N9, N141);
xor XOR2 (N519, N515, N204);
and AND4 (N520, N519, N223, N381, N39);
not NOT1 (N521, N503);
and AND2 (N522, N521, N242);
xor XOR2 (N523, N510, N23);
buf BUF1 (N524, N505);
and AND3 (N525, N511, N62, N421);
and AND4 (N526, N523, N193, N440, N116);
nand NAND2 (N527, N516, N266);
nor NOR4 (N528, N509, N430, N115, N161);
or OR4 (N529, N528, N363, N208, N292);
nand NAND3 (N530, N522, N477, N125);
buf BUF1 (N531, N520);
nor NOR4 (N532, N527, N25, N153, N290);
buf BUF1 (N533, N525);
or OR2 (N534, N533, N174);
not NOT1 (N535, N532);
xor XOR2 (N536, N514, N379);
buf BUF1 (N537, N535);
or OR4 (N538, N530, N298, N65, N272);
or OR3 (N539, N537, N193, N9);
xor XOR2 (N540, N538, N89);
xor XOR2 (N541, N539, N462);
nor NOR4 (N542, N540, N189, N231, N483);
or OR2 (N543, N542, N382);
nor NOR4 (N544, N529, N251, N28, N342);
buf BUF1 (N545, N518);
nor NOR3 (N546, N536, N116, N543);
buf BUF1 (N547, N100);
nand NAND4 (N548, N524, N187, N523, N526);
xor XOR2 (N549, N444, N272);
or OR2 (N550, N546, N438);
not NOT1 (N551, N544);
nor NOR3 (N552, N548, N331, N3);
buf BUF1 (N553, N534);
or OR3 (N554, N552, N101, N54);
nor NOR3 (N555, N547, N391, N16);
buf BUF1 (N556, N545);
nand NAND2 (N557, N531, N57);
buf BUF1 (N558, N557);
not NOT1 (N559, N496);
not NOT1 (N560, N550);
nor NOR3 (N561, N558, N449, N458);
xor XOR2 (N562, N559, N307);
not NOT1 (N563, N553);
not NOT1 (N564, N549);
not NOT1 (N565, N555);
nor NOR2 (N566, N554, N268);
nand NAND4 (N567, N566, N186, N273, N511);
nand NAND4 (N568, N541, N243, N55, N252);
nor NOR4 (N569, N551, N159, N140, N511);
or OR2 (N570, N562, N204);
xor XOR2 (N571, N560, N407);
or OR3 (N572, N567, N144, N198);
or OR4 (N573, N563, N435, N495, N94);
and AND2 (N574, N571, N187);
or OR3 (N575, N572, N372, N253);
nor NOR3 (N576, N570, N144, N39);
nand NAND4 (N577, N568, N1, N276, N348);
or OR4 (N578, N577, N125, N216, N394);
nor NOR3 (N579, N564, N126, N60);
and AND4 (N580, N578, N319, N514, N69);
and AND2 (N581, N569, N527);
not NOT1 (N582, N581);
xor XOR2 (N583, N575, N392);
or OR2 (N584, N573, N174);
nor NOR4 (N585, N584, N412, N408, N369);
buf BUF1 (N586, N585);
not NOT1 (N587, N574);
xor XOR2 (N588, N580, N579);
and AND4 (N589, N389, N10, N212, N357);
and AND4 (N590, N556, N300, N220, N78);
and AND3 (N591, N590, N456, N214);
xor XOR2 (N592, N583, N236);
or OR2 (N593, N565, N214);
xor XOR2 (N594, N561, N361);
buf BUF1 (N595, N592);
buf BUF1 (N596, N591);
or OR4 (N597, N594, N556, N396, N130);
and AND4 (N598, N576, N337, N424, N544);
or OR4 (N599, N596, N398, N311, N570);
not NOT1 (N600, N597);
not NOT1 (N601, N599);
not NOT1 (N602, N595);
buf BUF1 (N603, N598);
or OR4 (N604, N593, N489, N567, N559);
not NOT1 (N605, N587);
xor XOR2 (N606, N600, N1);
nor NOR2 (N607, N586, N563);
nor NOR2 (N608, N603, N339);
nand NAND4 (N609, N607, N269, N574, N241);
nor NOR4 (N610, N582, N567, N283, N351);
or OR4 (N611, N589, N570, N391, N579);
not NOT1 (N612, N604);
or OR3 (N613, N602, N336, N60);
and AND3 (N614, N605, N294, N551);
not NOT1 (N615, N610);
and AND3 (N616, N588, N129, N354);
nor NOR3 (N617, N608, N129, N232);
xor XOR2 (N618, N606, N58);
xor XOR2 (N619, N612, N391);
or OR2 (N620, N609, N126);
not NOT1 (N621, N611);
not NOT1 (N622, N618);
xor XOR2 (N623, N621, N325);
or OR2 (N624, N616, N619);
not NOT1 (N625, N357);
xor XOR2 (N626, N620, N413);
and AND4 (N627, N617, N222, N521, N416);
and AND3 (N628, N615, N528, N399);
and AND3 (N629, N626, N466, N628);
and AND3 (N630, N537, N399, N454);
buf BUF1 (N631, N613);
nand NAND4 (N632, N631, N365, N477, N614);
nand NAND4 (N633, N376, N150, N396, N273);
and AND3 (N634, N633, N50, N253);
buf BUF1 (N635, N629);
buf BUF1 (N636, N601);
nor NOR3 (N637, N625, N570, N170);
nand NAND3 (N638, N627, N295, N54);
nor NOR4 (N639, N632, N133, N150, N123);
xor XOR2 (N640, N624, N121);
or OR3 (N641, N640, N103, N422);
not NOT1 (N642, N637);
xor XOR2 (N643, N642, N376);
nand NAND4 (N644, N638, N228, N502, N13);
or OR3 (N645, N644, N556, N395);
or OR4 (N646, N641, N602, N96, N290);
nor NOR4 (N647, N623, N113, N9, N352);
nor NOR4 (N648, N639, N514, N104, N118);
and AND2 (N649, N622, N552);
xor XOR2 (N650, N646, N192);
and AND4 (N651, N634, N350, N479, N341);
xor XOR2 (N652, N648, N50);
and AND3 (N653, N650, N277, N206);
nor NOR2 (N654, N630, N486);
or OR2 (N655, N645, N337);
not NOT1 (N656, N643);
buf BUF1 (N657, N651);
not NOT1 (N658, N649);
nand NAND2 (N659, N654, N140);
and AND2 (N660, N635, N351);
or OR4 (N661, N636, N16, N567, N84);
xor XOR2 (N662, N659, N415);
xor XOR2 (N663, N657, N132);
not NOT1 (N664, N653);
xor XOR2 (N665, N662, N483);
xor XOR2 (N666, N656, N200);
not NOT1 (N667, N652);
or OR2 (N668, N667, N416);
or OR3 (N669, N660, N268, N468);
not NOT1 (N670, N664);
buf BUF1 (N671, N663);
and AND3 (N672, N665, N533, N367);
nor NOR4 (N673, N672, N453, N132, N32);
buf BUF1 (N674, N655);
or OR2 (N675, N668, N402);
and AND2 (N676, N666, N467);
xor XOR2 (N677, N676, N25);
buf BUF1 (N678, N671);
buf BUF1 (N679, N647);
xor XOR2 (N680, N670, N549);
not NOT1 (N681, N658);
and AND2 (N682, N678, N471);
buf BUF1 (N683, N680);
buf BUF1 (N684, N679);
or OR2 (N685, N681, N38);
buf BUF1 (N686, N683);
nor NOR2 (N687, N661, N90);
nand NAND4 (N688, N685, N523, N352, N569);
not NOT1 (N689, N686);
xor XOR2 (N690, N669, N651);
or OR4 (N691, N682, N154, N192, N568);
nand NAND2 (N692, N677, N544);
or OR4 (N693, N689, N256, N626, N590);
or OR2 (N694, N674, N686);
nand NAND2 (N695, N673, N437);
buf BUF1 (N696, N690);
and AND3 (N697, N691, N603, N76);
and AND3 (N698, N693, N677, N590);
nor NOR4 (N699, N687, N99, N222, N101);
not NOT1 (N700, N694);
or OR3 (N701, N675, N334, N12);
nor NOR3 (N702, N684, N203, N148);
nand NAND3 (N703, N700, N337, N694);
nand NAND3 (N704, N698, N384, N564);
or OR4 (N705, N695, N390, N88, N524);
buf BUF1 (N706, N688);
buf BUF1 (N707, N703);
nand NAND2 (N708, N696, N604);
not NOT1 (N709, N692);
nand NAND2 (N710, N708, N587);
nand NAND4 (N711, N704, N355, N111, N165);
and AND2 (N712, N705, N451);
and AND4 (N713, N712, N64, N377, N275);
and AND3 (N714, N711, N156, N586);
or OR4 (N715, N702, N494, N135, N179);
nand NAND4 (N716, N697, N147, N214, N378);
not NOT1 (N717, N706);
xor XOR2 (N718, N716, N653);
not NOT1 (N719, N699);
and AND2 (N720, N710, N710);
nand NAND4 (N721, N719, N694, N611, N129);
not NOT1 (N722, N701);
nor NOR4 (N723, N718, N142, N131, N491);
or OR3 (N724, N707, N470, N326);
nor NOR3 (N725, N717, N640, N88);
or OR3 (N726, N714, N498, N579);
xor XOR2 (N727, N721, N549);
xor XOR2 (N728, N715, N378);
nand NAND4 (N729, N723, N483, N537, N533);
nor NOR3 (N730, N725, N157, N465);
not NOT1 (N731, N726);
or OR3 (N732, N730, N646, N222);
nand NAND2 (N733, N722, N582);
xor XOR2 (N734, N732, N415);
nor NOR3 (N735, N724, N391, N469);
nor NOR4 (N736, N735, N160, N243, N166);
and AND2 (N737, N736, N698);
or OR4 (N738, N737, N41, N368, N382);
xor XOR2 (N739, N731, N613);
xor XOR2 (N740, N739, N446);
and AND4 (N741, N740, N312, N134, N453);
not NOT1 (N742, N741);
or OR4 (N743, N742, N474, N558, N683);
nor NOR2 (N744, N734, N161);
nand NAND2 (N745, N713, N110);
not NOT1 (N746, N727);
or OR4 (N747, N738, N300, N734, N72);
nor NOR3 (N748, N728, N122, N734);
buf BUF1 (N749, N709);
and AND2 (N750, N733, N343);
nor NOR2 (N751, N720, N480);
not NOT1 (N752, N729);
and AND2 (N753, N745, N564);
xor XOR2 (N754, N751, N409);
not NOT1 (N755, N744);
xor XOR2 (N756, N748, N491);
not NOT1 (N757, N743);
buf BUF1 (N758, N747);
or OR3 (N759, N749, N521, N219);
xor XOR2 (N760, N750, N249);
nand NAND2 (N761, N754, N469);
xor XOR2 (N762, N753, N277);
not NOT1 (N763, N761);
nor NOR2 (N764, N755, N71);
nand NAND3 (N765, N756, N19, N230);
and AND2 (N766, N763, N478);
not NOT1 (N767, N766);
buf BUF1 (N768, N767);
nand NAND4 (N769, N760, N42, N65, N662);
and AND4 (N770, N765, N527, N659, N300);
or OR3 (N771, N759, N177, N676);
buf BUF1 (N772, N769);
buf BUF1 (N773, N758);
not NOT1 (N774, N768);
or OR3 (N775, N752, N615, N568);
not NOT1 (N776, N775);
not NOT1 (N777, N770);
buf BUF1 (N778, N764);
or OR2 (N779, N762, N262);
not NOT1 (N780, N778);
nor NOR2 (N781, N773, N591);
or OR4 (N782, N779, N570, N134, N55);
not NOT1 (N783, N777);
xor XOR2 (N784, N772, N2);
and AND2 (N785, N783, N643);
nand NAND2 (N786, N784, N101);
nor NOR4 (N787, N782, N183, N357, N714);
not NOT1 (N788, N757);
and AND2 (N789, N776, N769);
not NOT1 (N790, N780);
or OR3 (N791, N785, N113, N591);
not NOT1 (N792, N781);
buf BUF1 (N793, N791);
or OR4 (N794, N789, N419, N365, N620);
and AND4 (N795, N792, N781, N253, N717);
xor XOR2 (N796, N771, N375);
nand NAND2 (N797, N790, N2);
xor XOR2 (N798, N794, N72);
xor XOR2 (N799, N788, N181);
nor NOR3 (N800, N799, N679, N160);
or OR4 (N801, N800, N361, N66, N353);
nand NAND4 (N802, N786, N254, N154, N445);
nor NOR2 (N803, N801, N590);
or OR3 (N804, N787, N340, N88);
and AND4 (N805, N802, N131, N387, N173);
and AND3 (N806, N774, N337, N792);
nor NOR2 (N807, N793, N691);
nor NOR3 (N808, N803, N705, N286);
or OR4 (N809, N796, N351, N160, N604);
not NOT1 (N810, N808);
and AND3 (N811, N746, N318, N575);
and AND2 (N812, N797, N369);
buf BUF1 (N813, N810);
nor NOR3 (N814, N812, N16, N329);
xor XOR2 (N815, N804, N87);
not NOT1 (N816, N813);
xor XOR2 (N817, N798, N221);
or OR2 (N818, N817, N383);
xor XOR2 (N819, N818, N609);
buf BUF1 (N820, N819);
buf BUF1 (N821, N805);
xor XOR2 (N822, N807, N543);
buf BUF1 (N823, N821);
nand NAND4 (N824, N795, N51, N130, N614);
not NOT1 (N825, N809);
xor XOR2 (N826, N806, N314);
nor NOR4 (N827, N822, N413, N48, N534);
buf BUF1 (N828, N820);
nand NAND4 (N829, N814, N160, N157, N486);
xor XOR2 (N830, N825, N158);
nor NOR4 (N831, N811, N651, N775, N377);
nand NAND2 (N832, N828, N758);
nand NAND3 (N833, N830, N713, N338);
nand NAND2 (N834, N832, N214);
nor NOR3 (N835, N816, N16, N272);
nor NOR4 (N836, N831, N483, N751, N143);
or OR4 (N837, N824, N734, N628, N81);
nor NOR3 (N838, N815, N202, N807);
or OR4 (N839, N834, N134, N467, N306);
or OR2 (N840, N827, N248);
or OR4 (N841, N826, N260, N408, N5);
buf BUF1 (N842, N838);
nand NAND2 (N843, N835, N783);
nor NOR3 (N844, N829, N776, N738);
not NOT1 (N845, N837);
or OR3 (N846, N833, N785, N598);
not NOT1 (N847, N839);
nor NOR2 (N848, N823, N52);
xor XOR2 (N849, N845, N685);
or OR4 (N850, N843, N50, N66, N837);
and AND3 (N851, N842, N547, N844);
or OR2 (N852, N76, N196);
nand NAND2 (N853, N847, N619);
nor NOR4 (N854, N853, N808, N757, N851);
and AND4 (N855, N258, N502, N721, N573);
and AND2 (N856, N855, N664);
or OR4 (N857, N849, N632, N499, N228);
and AND3 (N858, N852, N516, N733);
xor XOR2 (N859, N854, N88);
xor XOR2 (N860, N857, N620);
nor NOR4 (N861, N859, N218, N101, N387);
nand NAND2 (N862, N856, N462);
and AND3 (N863, N862, N688, N496);
or OR3 (N864, N840, N202, N779);
xor XOR2 (N865, N850, N842);
buf BUF1 (N866, N863);
buf BUF1 (N867, N841);
nand NAND4 (N868, N860, N675, N485, N77);
or OR4 (N869, N861, N234, N477, N36);
buf BUF1 (N870, N868);
xor XOR2 (N871, N869, N41);
buf BUF1 (N872, N870);
nor NOR4 (N873, N848, N662, N656, N600);
and AND3 (N874, N846, N601, N38);
nor NOR4 (N875, N858, N351, N195, N142);
not NOT1 (N876, N874);
and AND4 (N877, N865, N32, N330, N485);
and AND4 (N878, N873, N365, N170, N640);
not NOT1 (N879, N872);
nand NAND3 (N880, N864, N536, N755);
xor XOR2 (N881, N867, N541);
xor XOR2 (N882, N880, N341);
or OR2 (N883, N866, N215);
xor XOR2 (N884, N876, N702);
and AND2 (N885, N882, N468);
nor NOR3 (N886, N883, N220, N704);
not NOT1 (N887, N884);
not NOT1 (N888, N875);
buf BUF1 (N889, N886);
not NOT1 (N890, N888);
nand NAND3 (N891, N836, N395, N687);
xor XOR2 (N892, N879, N504);
xor XOR2 (N893, N889, N841);
and AND3 (N894, N881, N446, N684);
not NOT1 (N895, N894);
or OR4 (N896, N871, N71, N428, N794);
and AND3 (N897, N885, N830, N96);
nor NOR4 (N898, N896, N839, N45, N280);
not NOT1 (N899, N891);
or OR2 (N900, N899, N190);
not NOT1 (N901, N900);
not NOT1 (N902, N878);
buf BUF1 (N903, N890);
and AND2 (N904, N898, N563);
not NOT1 (N905, N897);
buf BUF1 (N906, N893);
xor XOR2 (N907, N903, N100);
nor NOR2 (N908, N887, N866);
xor XOR2 (N909, N905, N224);
and AND2 (N910, N892, N20);
buf BUF1 (N911, N904);
and AND2 (N912, N906, N723);
nor NOR4 (N913, N895, N264, N86, N797);
buf BUF1 (N914, N908);
buf BUF1 (N915, N877);
not NOT1 (N916, N901);
buf BUF1 (N917, N910);
xor XOR2 (N918, N913, N426);
nor NOR2 (N919, N902, N380);
nor NOR2 (N920, N918, N517);
and AND2 (N921, N915, N651);
not NOT1 (N922, N912);
or OR3 (N923, N917, N854, N494);
not NOT1 (N924, N921);
xor XOR2 (N925, N920, N162);
and AND3 (N926, N925, N781, N440);
or OR2 (N927, N922, N86);
xor XOR2 (N928, N914, N379);
buf BUF1 (N929, N928);
and AND3 (N930, N919, N812, N439);
nor NOR4 (N931, N924, N896, N924, N816);
xor XOR2 (N932, N907, N837);
or OR2 (N933, N923, N481);
nand NAND3 (N934, N909, N849, N262);
xor XOR2 (N935, N934, N814);
nand NAND2 (N936, N932, N53);
xor XOR2 (N937, N926, N565);
not NOT1 (N938, N933);
and AND2 (N939, N916, N277);
not NOT1 (N940, N929);
and AND4 (N941, N936, N479, N25, N129);
not NOT1 (N942, N939);
nor NOR4 (N943, N942, N446, N367, N552);
xor XOR2 (N944, N911, N838);
xor XOR2 (N945, N935, N847);
nand NAND3 (N946, N941, N387, N866);
and AND3 (N947, N940, N753, N929);
not NOT1 (N948, N927);
nor NOR3 (N949, N938, N741, N242);
and AND3 (N950, N937, N759, N878);
not NOT1 (N951, N948);
buf BUF1 (N952, N946);
not NOT1 (N953, N949);
nor NOR3 (N954, N930, N114, N347);
or OR4 (N955, N952, N693, N679, N433);
buf BUF1 (N956, N953);
xor XOR2 (N957, N955, N808);
nor NOR2 (N958, N956, N622);
xor XOR2 (N959, N954, N656);
nor NOR2 (N960, N943, N22);
and AND2 (N961, N945, N282);
buf BUF1 (N962, N961);
xor XOR2 (N963, N947, N2);
nand NAND4 (N964, N931, N299, N64, N146);
not NOT1 (N965, N959);
nand NAND3 (N966, N962, N43, N860);
buf BUF1 (N967, N958);
and AND2 (N968, N960, N176);
not NOT1 (N969, N967);
not NOT1 (N970, N964);
xor XOR2 (N971, N969, N655);
or OR4 (N972, N970, N8, N688, N336);
nor NOR2 (N973, N968, N841);
nor NOR4 (N974, N944, N71, N305, N356);
or OR4 (N975, N972, N565, N231, N707);
or OR4 (N976, N975, N552, N156, N149);
xor XOR2 (N977, N974, N507);
and AND2 (N978, N977, N642);
xor XOR2 (N979, N957, N850);
not NOT1 (N980, N966);
and AND4 (N981, N980, N347, N177, N367);
and AND4 (N982, N973, N149, N883, N405);
xor XOR2 (N983, N965, N136);
or OR3 (N984, N963, N803, N790);
xor XOR2 (N985, N983, N600);
nor NOR2 (N986, N971, N643);
xor XOR2 (N987, N951, N101);
nand NAND2 (N988, N987, N975);
not NOT1 (N989, N984);
buf BUF1 (N990, N988);
or OR2 (N991, N990, N396);
buf BUF1 (N992, N991);
or OR2 (N993, N976, N86);
buf BUF1 (N994, N982);
not NOT1 (N995, N989);
and AND4 (N996, N986, N842, N770, N309);
xor XOR2 (N997, N950, N844);
nand NAND2 (N998, N995, N627);
nand NAND3 (N999, N994, N657, N305);
not NOT1 (N1000, N998);
or OR4 (N1001, N997, N208, N29, N551);
xor XOR2 (N1002, N1000, N538);
nand NAND3 (N1003, N992, N304, N3);
nand NAND4 (N1004, N999, N351, N2, N763);
xor XOR2 (N1005, N985, N868);
nand NAND4 (N1006, N1001, N525, N408, N688);
xor XOR2 (N1007, N1004, N589);
buf BUF1 (N1008, N993);
nand NAND4 (N1009, N1003, N375, N333, N577);
nand NAND2 (N1010, N1008, N50);
buf BUF1 (N1011, N1010);
xor XOR2 (N1012, N1005, N313);
and AND4 (N1013, N1011, N947, N182, N593);
nand NAND4 (N1014, N1006, N743, N684, N667);
xor XOR2 (N1015, N1007, N303);
and AND2 (N1016, N1013, N722);
nor NOR2 (N1017, N979, N773);
or OR4 (N1018, N1014, N557, N403, N864);
and AND4 (N1019, N1016, N684, N134, N147);
xor XOR2 (N1020, N1009, N953);
buf BUF1 (N1021, N1020);
not NOT1 (N1022, N996);
buf BUF1 (N1023, N1019);
nand NAND3 (N1024, N1023, N157, N676);
xor XOR2 (N1025, N1015, N1011);
or OR4 (N1026, N978, N783, N1013, N998);
nand NAND2 (N1027, N1024, N928);
xor XOR2 (N1028, N1002, N865);
nand NAND2 (N1029, N1012, N188);
xor XOR2 (N1030, N1026, N214);
nand NAND2 (N1031, N1029, N741);
xor XOR2 (N1032, N1030, N863);
nand NAND4 (N1033, N1031, N247, N89, N871);
nor NOR3 (N1034, N1033, N449, N733);
and AND2 (N1035, N1021, N97);
nand NAND3 (N1036, N1035, N131, N571);
or OR2 (N1037, N1025, N949);
nand NAND2 (N1038, N1028, N548);
nor NOR3 (N1039, N1036, N597, N59);
not NOT1 (N1040, N981);
nor NOR2 (N1041, N1037, N174);
or OR3 (N1042, N1027, N360, N48);
and AND3 (N1043, N1041, N261, N461);
xor XOR2 (N1044, N1043, N232);
nand NAND4 (N1045, N1042, N575, N284, N542);
xor XOR2 (N1046, N1022, N328);
buf BUF1 (N1047, N1045);
buf BUF1 (N1048, N1039);
or OR4 (N1049, N1032, N100, N227, N853);
nor NOR4 (N1050, N1044, N958, N966, N387);
xor XOR2 (N1051, N1049, N696);
nor NOR2 (N1052, N1047, N129);
buf BUF1 (N1053, N1051);
and AND3 (N1054, N1046, N736, N202);
xor XOR2 (N1055, N1018, N918);
buf BUF1 (N1056, N1017);
and AND4 (N1057, N1052, N26, N941, N519);
buf BUF1 (N1058, N1040);
or OR3 (N1059, N1053, N1035, N754);
buf BUF1 (N1060, N1048);
not NOT1 (N1061, N1055);
or OR4 (N1062, N1050, N1031, N64, N1004);
and AND2 (N1063, N1062, N277);
not NOT1 (N1064, N1059);
nor NOR3 (N1065, N1054, N333, N860);
or OR4 (N1066, N1060, N334, N381, N579);
xor XOR2 (N1067, N1034, N720);
not NOT1 (N1068, N1058);
not NOT1 (N1069, N1067);
or OR2 (N1070, N1066, N432);
buf BUF1 (N1071, N1057);
xor XOR2 (N1072, N1069, N747);
xor XOR2 (N1073, N1038, N948);
nand NAND3 (N1074, N1056, N764, N249);
not NOT1 (N1075, N1074);
nor NOR4 (N1076, N1071, N283, N241, N706);
nand NAND4 (N1077, N1063, N680, N749, N779);
xor XOR2 (N1078, N1064, N684);
xor XOR2 (N1079, N1077, N211);
xor XOR2 (N1080, N1065, N985);
and AND3 (N1081, N1068, N681, N668);
buf BUF1 (N1082, N1081);
and AND3 (N1083, N1076, N684, N528);
or OR4 (N1084, N1079, N1024, N998, N967);
and AND2 (N1085, N1082, N736);
buf BUF1 (N1086, N1073);
or OR3 (N1087, N1080, N770, N398);
not NOT1 (N1088, N1070);
nor NOR2 (N1089, N1075, N627);
xor XOR2 (N1090, N1061, N140);
nand NAND4 (N1091, N1072, N846, N370, N1078);
xor XOR2 (N1092, N15, N807);
or OR3 (N1093, N1089, N982, N673);
and AND4 (N1094, N1093, N309, N580, N498);
and AND2 (N1095, N1086, N1033);
nor NOR2 (N1096, N1094, N30);
xor XOR2 (N1097, N1090, N1037);
not NOT1 (N1098, N1087);
nor NOR2 (N1099, N1092, N79);
buf BUF1 (N1100, N1083);
not NOT1 (N1101, N1088);
or OR4 (N1102, N1091, N221, N787, N1097);
buf BUF1 (N1103, N674);
nor NOR3 (N1104, N1099, N164, N760);
not NOT1 (N1105, N1096);
not NOT1 (N1106, N1095);
xor XOR2 (N1107, N1098, N1006);
buf BUF1 (N1108, N1084);
nand NAND4 (N1109, N1100, N471, N800, N764);
or OR3 (N1110, N1085, N676, N323);
nor NOR4 (N1111, N1106, N664, N537, N354);
and AND2 (N1112, N1101, N150);
buf BUF1 (N1113, N1105);
xor XOR2 (N1114, N1109, N849);
nor NOR3 (N1115, N1114, N80, N727);
buf BUF1 (N1116, N1115);
xor XOR2 (N1117, N1104, N477);
nand NAND3 (N1118, N1103, N123, N1009);
xor XOR2 (N1119, N1117, N94);
or OR3 (N1120, N1111, N637, N851);
and AND2 (N1121, N1108, N651);
buf BUF1 (N1122, N1112);
xor XOR2 (N1123, N1102, N93);
xor XOR2 (N1124, N1107, N181);
or OR4 (N1125, N1124, N766, N309, N1117);
nor NOR4 (N1126, N1125, N357, N1017, N147);
xor XOR2 (N1127, N1123, N1082);
nor NOR2 (N1128, N1110, N182);
and AND4 (N1129, N1127, N831, N519, N430);
or OR3 (N1130, N1118, N472, N70);
nand NAND4 (N1131, N1113, N556, N477, N90);
xor XOR2 (N1132, N1128, N776);
nor NOR4 (N1133, N1132, N832, N639, N394);
not NOT1 (N1134, N1119);
buf BUF1 (N1135, N1131);
not NOT1 (N1136, N1130);
or OR4 (N1137, N1121, N525, N1022, N970);
nor NOR4 (N1138, N1126, N452, N197, N40);
buf BUF1 (N1139, N1120);
xor XOR2 (N1140, N1129, N702);
nor NOR2 (N1141, N1137, N571);
not NOT1 (N1142, N1141);
or OR3 (N1143, N1122, N1122, N34);
nand NAND2 (N1144, N1133, N918);
buf BUF1 (N1145, N1116);
buf BUF1 (N1146, N1145);
and AND4 (N1147, N1146, N1012, N209, N678);
nand NAND4 (N1148, N1135, N1071, N290, N916);
xor XOR2 (N1149, N1148, N920);
nand NAND3 (N1150, N1139, N251, N708);
xor XOR2 (N1151, N1144, N236);
not NOT1 (N1152, N1142);
xor XOR2 (N1153, N1150, N343);
and AND2 (N1154, N1138, N703);
buf BUF1 (N1155, N1140);
and AND3 (N1156, N1149, N652, N700);
xor XOR2 (N1157, N1156, N910);
or OR3 (N1158, N1143, N98, N812);
not NOT1 (N1159, N1158);
buf BUF1 (N1160, N1157);
buf BUF1 (N1161, N1153);
nand NAND2 (N1162, N1151, N693);
nor NOR3 (N1163, N1161, N397, N1034);
and AND3 (N1164, N1159, N332, N406);
buf BUF1 (N1165, N1147);
nand NAND3 (N1166, N1163, N1006, N926);
buf BUF1 (N1167, N1134);
buf BUF1 (N1168, N1164);
xor XOR2 (N1169, N1155, N407);
xor XOR2 (N1170, N1136, N951);
nand NAND3 (N1171, N1169, N567, N122);
or OR4 (N1172, N1152, N897, N1070, N986);
nand NAND4 (N1173, N1162, N937, N1151, N760);
or OR4 (N1174, N1166, N612, N254, N1160);
buf BUF1 (N1175, N1073);
or OR2 (N1176, N1171, N930);
buf BUF1 (N1177, N1170);
nand NAND4 (N1178, N1173, N412, N774, N314);
nand NAND4 (N1179, N1174, N523, N35, N146);
nand NAND4 (N1180, N1154, N352, N897, N91);
buf BUF1 (N1181, N1172);
and AND2 (N1182, N1175, N475);
or OR3 (N1183, N1167, N98, N155);
xor XOR2 (N1184, N1181, N970);
buf BUF1 (N1185, N1178);
xor XOR2 (N1186, N1183, N350);
nand NAND4 (N1187, N1185, N1026, N39, N556);
not NOT1 (N1188, N1180);
xor XOR2 (N1189, N1188, N695);
or OR4 (N1190, N1176, N113, N569, N309);
and AND3 (N1191, N1182, N77, N628);
nand NAND4 (N1192, N1189, N940, N1135, N69);
nand NAND4 (N1193, N1191, N1001, N202, N351);
nand NAND4 (N1194, N1179, N1187, N28, N236);
nand NAND3 (N1195, N1160, N1043, N770);
nand NAND4 (N1196, N1165, N1048, N521, N52);
xor XOR2 (N1197, N1196, N383);
nor NOR2 (N1198, N1168, N192);
nor NOR2 (N1199, N1198, N854);
not NOT1 (N1200, N1194);
xor XOR2 (N1201, N1186, N913);
or OR3 (N1202, N1195, N1184, N188);
nor NOR2 (N1203, N274, N315);
and AND4 (N1204, N1201, N699, N212, N1118);
buf BUF1 (N1205, N1203);
or OR3 (N1206, N1202, N1127, N1076);
or OR4 (N1207, N1205, N1014, N830, N1131);
not NOT1 (N1208, N1193);
nand NAND3 (N1209, N1200, N1095, N394);
nand NAND2 (N1210, N1208, N53);
or OR4 (N1211, N1209, N597, N1042, N1116);
nor NOR2 (N1212, N1197, N5);
nand NAND3 (N1213, N1192, N1009, N674);
or OR4 (N1214, N1190, N522, N454, N309);
buf BUF1 (N1215, N1207);
buf BUF1 (N1216, N1206);
buf BUF1 (N1217, N1204);
buf BUF1 (N1218, N1217);
not NOT1 (N1219, N1218);
or OR4 (N1220, N1210, N1022, N1036, N1004);
buf BUF1 (N1221, N1220);
not NOT1 (N1222, N1199);
buf BUF1 (N1223, N1214);
or OR2 (N1224, N1222, N1172);
not NOT1 (N1225, N1212);
and AND2 (N1226, N1223, N1013);
and AND4 (N1227, N1224, N958, N245, N877);
nor NOR3 (N1228, N1225, N543, N550);
xor XOR2 (N1229, N1227, N1013);
nor NOR3 (N1230, N1216, N379, N1154);
and AND3 (N1231, N1211, N113, N411);
and AND4 (N1232, N1226, N1058, N439, N81);
and AND3 (N1233, N1219, N610, N182);
nor NOR3 (N1234, N1232, N10, N396);
nor NOR3 (N1235, N1228, N1148, N1188);
xor XOR2 (N1236, N1221, N22);
not NOT1 (N1237, N1213);
xor XOR2 (N1238, N1237, N984);
xor XOR2 (N1239, N1235, N583);
nand NAND2 (N1240, N1236, N408);
nor NOR2 (N1241, N1240, N688);
or OR3 (N1242, N1238, N403, N98);
and AND2 (N1243, N1230, N258);
xor XOR2 (N1244, N1241, N466);
nand NAND2 (N1245, N1233, N1185);
nand NAND3 (N1246, N1244, N927, N580);
nor NOR4 (N1247, N1242, N495, N369, N367);
and AND4 (N1248, N1239, N288, N717, N1064);
or OR4 (N1249, N1248, N915, N1195, N290);
nor NOR4 (N1250, N1177, N655, N369, N491);
and AND2 (N1251, N1231, N998);
nor NOR3 (N1252, N1249, N952, N1029);
nand NAND2 (N1253, N1229, N821);
nor NOR4 (N1254, N1250, N814, N77, N385);
nor NOR4 (N1255, N1254, N1218, N43, N891);
nor NOR3 (N1256, N1252, N997, N545);
and AND3 (N1257, N1251, N34, N569);
buf BUF1 (N1258, N1246);
not NOT1 (N1259, N1258);
nand NAND3 (N1260, N1247, N649, N24);
or OR3 (N1261, N1256, N769, N348);
buf BUF1 (N1262, N1253);
buf BUF1 (N1263, N1255);
or OR4 (N1264, N1215, N259, N60, N546);
xor XOR2 (N1265, N1262, N38);
or OR3 (N1266, N1245, N343, N121);
and AND3 (N1267, N1264, N1112, N444);
or OR2 (N1268, N1234, N727);
and AND3 (N1269, N1243, N417, N1122);
xor XOR2 (N1270, N1268, N1059);
not NOT1 (N1271, N1259);
buf BUF1 (N1272, N1261);
or OR4 (N1273, N1257, N127, N225, N224);
nand NAND2 (N1274, N1273, N827);
and AND2 (N1275, N1263, N402);
or OR4 (N1276, N1260, N823, N1238, N90);
nor NOR3 (N1277, N1267, N662, N415);
nand NAND2 (N1278, N1271, N221);
nor NOR4 (N1279, N1277, N315, N97, N879);
and AND4 (N1280, N1270, N689, N599, N119);
nand NAND4 (N1281, N1278, N430, N855, N66);
not NOT1 (N1282, N1275);
or OR3 (N1283, N1272, N1195, N699);
nor NOR2 (N1284, N1280, N1080);
nor NOR4 (N1285, N1265, N629, N742, N416);
not NOT1 (N1286, N1266);
and AND2 (N1287, N1279, N1111);
and AND3 (N1288, N1286, N1168, N1227);
xor XOR2 (N1289, N1269, N418);
not NOT1 (N1290, N1282);
buf BUF1 (N1291, N1281);
nand NAND3 (N1292, N1284, N1223, N939);
buf BUF1 (N1293, N1274);
not NOT1 (N1294, N1285);
nand NAND2 (N1295, N1283, N1224);
buf BUF1 (N1296, N1294);
nor NOR2 (N1297, N1296, N602);
or OR3 (N1298, N1289, N481, N384);
or OR3 (N1299, N1297, N151, N80);
and AND4 (N1300, N1291, N1141, N1133, N988);
xor XOR2 (N1301, N1276, N704);
not NOT1 (N1302, N1290);
nand NAND3 (N1303, N1302, N341, N797);
buf BUF1 (N1304, N1293);
nor NOR2 (N1305, N1303, N1254);
not NOT1 (N1306, N1295);
xor XOR2 (N1307, N1292, N338);
nor NOR4 (N1308, N1307, N434, N739, N161);
and AND3 (N1309, N1308, N1013, N381);
and AND4 (N1310, N1306, N681, N774, N1289);
not NOT1 (N1311, N1304);
and AND2 (N1312, N1309, N673);
not NOT1 (N1313, N1300);
not NOT1 (N1314, N1298);
not NOT1 (N1315, N1305);
nor NOR2 (N1316, N1310, N927);
nand NAND2 (N1317, N1315, N750);
nor NOR4 (N1318, N1288, N1197, N588, N906);
nand NAND3 (N1319, N1312, N234, N748);
nor NOR2 (N1320, N1318, N518);
xor XOR2 (N1321, N1301, N487);
nor NOR2 (N1322, N1317, N86);
xor XOR2 (N1323, N1313, N484);
nand NAND3 (N1324, N1319, N659, N735);
and AND3 (N1325, N1320, N1059, N221);
or OR3 (N1326, N1287, N1125, N53);
nor NOR4 (N1327, N1299, N342, N1060, N554);
xor XOR2 (N1328, N1316, N311);
or OR3 (N1329, N1311, N962, N85);
nor NOR3 (N1330, N1323, N1187, N1293);
xor XOR2 (N1331, N1330, N858);
nor NOR2 (N1332, N1329, N1105);
buf BUF1 (N1333, N1327);
or OR3 (N1334, N1332, N612, N1261);
not NOT1 (N1335, N1325);
or OR4 (N1336, N1335, N360, N1234, N430);
nor NOR3 (N1337, N1321, N1005, N1289);
not NOT1 (N1338, N1336);
buf BUF1 (N1339, N1333);
nand NAND4 (N1340, N1334, N715, N38, N524);
or OR2 (N1341, N1314, N456);
xor XOR2 (N1342, N1324, N637);
or OR2 (N1343, N1328, N454);
nand NAND2 (N1344, N1338, N1062);
nand NAND4 (N1345, N1322, N552, N1255, N1082);
buf BUF1 (N1346, N1337);
buf BUF1 (N1347, N1326);
not NOT1 (N1348, N1343);
not NOT1 (N1349, N1345);
and AND2 (N1350, N1344, N687);
and AND3 (N1351, N1346, N612, N1091);
or OR2 (N1352, N1339, N504);
not NOT1 (N1353, N1342);
or OR4 (N1354, N1347, N611, N1174, N398);
or OR2 (N1355, N1354, N1246);
and AND2 (N1356, N1331, N60);
nand NAND4 (N1357, N1348, N1349, N1034, N962);
nor NOR4 (N1358, N1008, N386, N1171, N68);
nand NAND4 (N1359, N1358, N848, N1061, N1228);
xor XOR2 (N1360, N1355, N21);
buf BUF1 (N1361, N1350);
not NOT1 (N1362, N1353);
nand NAND4 (N1363, N1360, N903, N432, N830);
xor XOR2 (N1364, N1341, N842);
nand NAND4 (N1365, N1356, N391, N522, N901);
xor XOR2 (N1366, N1352, N888);
nand NAND4 (N1367, N1366, N313, N1122, N1220);
nor NOR2 (N1368, N1357, N425);
and AND3 (N1369, N1351, N637, N164);
or OR2 (N1370, N1367, N553);
nand NAND2 (N1371, N1370, N697);
nor NOR3 (N1372, N1361, N887, N1333);
buf BUF1 (N1373, N1359);
and AND2 (N1374, N1340, N454);
buf BUF1 (N1375, N1369);
nand NAND3 (N1376, N1365, N1252, N1300);
nand NAND4 (N1377, N1375, N540, N36, N1336);
buf BUF1 (N1378, N1374);
and AND2 (N1379, N1373, N891);
buf BUF1 (N1380, N1376);
or OR3 (N1381, N1379, N393, N691);
nor NOR3 (N1382, N1381, N108, N104);
not NOT1 (N1383, N1368);
or OR2 (N1384, N1372, N241);
not NOT1 (N1385, N1383);
not NOT1 (N1386, N1384);
or OR3 (N1387, N1378, N929, N1204);
and AND3 (N1388, N1362, N1154, N972);
nand NAND2 (N1389, N1371, N1336);
not NOT1 (N1390, N1389);
nand NAND4 (N1391, N1377, N726, N582, N127);
buf BUF1 (N1392, N1380);
nand NAND4 (N1393, N1363, N392, N81, N545);
and AND2 (N1394, N1386, N541);
and AND4 (N1395, N1392, N1051, N889, N972);
xor XOR2 (N1396, N1391, N387);
nand NAND3 (N1397, N1390, N541, N681);
xor XOR2 (N1398, N1394, N950);
not NOT1 (N1399, N1364);
or OR3 (N1400, N1398, N1304, N1138);
nor NOR3 (N1401, N1396, N761, N319);
nand NAND4 (N1402, N1400, N1069, N388, N640);
nor NOR3 (N1403, N1382, N1139, N1079);
xor XOR2 (N1404, N1388, N122);
xor XOR2 (N1405, N1402, N485);
and AND3 (N1406, N1405, N1401, N1359);
nor NOR3 (N1407, N308, N1100, N826);
xor XOR2 (N1408, N1387, N491);
xor XOR2 (N1409, N1403, N595);
xor XOR2 (N1410, N1407, N584);
nor NOR2 (N1411, N1406, N139);
xor XOR2 (N1412, N1395, N1313);
and AND4 (N1413, N1393, N12, N531, N275);
nand NAND3 (N1414, N1412, N120, N105);
nor NOR3 (N1415, N1413, N1409, N903);
and AND3 (N1416, N326, N71, N624);
and AND4 (N1417, N1414, N259, N530, N995);
nor NOR3 (N1418, N1385, N118, N954);
or OR3 (N1419, N1410, N759, N436);
buf BUF1 (N1420, N1411);
xor XOR2 (N1421, N1417, N667);
xor XOR2 (N1422, N1420, N1395);
nor NOR2 (N1423, N1418, N1250);
and AND3 (N1424, N1404, N737, N597);
or OR2 (N1425, N1397, N363);
not NOT1 (N1426, N1422);
not NOT1 (N1427, N1419);
not NOT1 (N1428, N1421);
nor NOR2 (N1429, N1425, N35);
buf BUF1 (N1430, N1423);
and AND3 (N1431, N1430, N415, N649);
xor XOR2 (N1432, N1428, N1285);
nand NAND3 (N1433, N1432, N1227, N625);
buf BUF1 (N1434, N1399);
and AND2 (N1435, N1415, N1356);
nor NOR4 (N1436, N1408, N411, N1082, N297);
nand NAND2 (N1437, N1426, N1017);
or OR2 (N1438, N1435, N970);
not NOT1 (N1439, N1416);
nand NAND4 (N1440, N1439, N853, N456, N566);
xor XOR2 (N1441, N1436, N280);
or OR2 (N1442, N1433, N1136);
nand NAND4 (N1443, N1431, N1092, N776, N323);
xor XOR2 (N1444, N1440, N215);
or OR2 (N1445, N1434, N554);
and AND3 (N1446, N1438, N430, N1143);
or OR3 (N1447, N1445, N216, N1340);
or OR2 (N1448, N1441, N1077);
or OR4 (N1449, N1427, N685, N687, N156);
and AND2 (N1450, N1446, N494);
buf BUF1 (N1451, N1447);
xor XOR2 (N1452, N1451, N1380);
nor NOR3 (N1453, N1443, N934, N19);
buf BUF1 (N1454, N1448);
and AND4 (N1455, N1453, N317, N24, N575);
not NOT1 (N1456, N1454);
nand NAND3 (N1457, N1449, N47, N45);
not NOT1 (N1458, N1450);
not NOT1 (N1459, N1424);
and AND4 (N1460, N1455, N214, N426, N72);
nor NOR4 (N1461, N1460, N388, N977, N708);
nor NOR4 (N1462, N1452, N1361, N858, N724);
and AND4 (N1463, N1437, N572, N923, N866);
not NOT1 (N1464, N1458);
nand NAND2 (N1465, N1462, N473);
or OR4 (N1466, N1463, N1387, N88, N1088);
nor NOR2 (N1467, N1429, N824);
nor NOR4 (N1468, N1457, N1009, N611, N643);
or OR2 (N1469, N1442, N567);
nand NAND3 (N1470, N1459, N159, N104);
or OR3 (N1471, N1468, N635, N1222);
not NOT1 (N1472, N1461);
buf BUF1 (N1473, N1470);
or OR4 (N1474, N1467, N50, N1078, N264);
not NOT1 (N1475, N1464);
not NOT1 (N1476, N1469);
and AND4 (N1477, N1476, N372, N752, N252);
not NOT1 (N1478, N1477);
nand NAND2 (N1479, N1474, N608);
not NOT1 (N1480, N1466);
not NOT1 (N1481, N1475);
xor XOR2 (N1482, N1479, N1220);
nand NAND4 (N1483, N1465, N133, N1305, N85);
and AND4 (N1484, N1456, N317, N474, N475);
nand NAND3 (N1485, N1444, N481, N240);
xor XOR2 (N1486, N1472, N541);
xor XOR2 (N1487, N1484, N1374);
buf BUF1 (N1488, N1485);
nand NAND3 (N1489, N1471, N39, N1014);
or OR2 (N1490, N1478, N142);
and AND3 (N1491, N1490, N901, N628);
or OR3 (N1492, N1482, N1327, N1438);
not NOT1 (N1493, N1491);
nand NAND3 (N1494, N1480, N690, N1464);
and AND3 (N1495, N1473, N991, N1113);
nor NOR3 (N1496, N1486, N665, N902);
buf BUF1 (N1497, N1487);
or OR2 (N1498, N1493, N1246);
not NOT1 (N1499, N1498);
nand NAND3 (N1500, N1497, N674, N339);
not NOT1 (N1501, N1496);
nor NOR2 (N1502, N1481, N178);
not NOT1 (N1503, N1494);
and AND2 (N1504, N1500, N1110);
nor NOR2 (N1505, N1499, N802);
nor NOR2 (N1506, N1483, N1062);
buf BUF1 (N1507, N1506);
nor NOR2 (N1508, N1507, N18);
nor NOR4 (N1509, N1502, N108, N374, N804);
nor NOR4 (N1510, N1495, N846, N628, N1000);
nor NOR4 (N1511, N1505, N1243, N203, N1499);
and AND4 (N1512, N1509, N524, N602, N1326);
nand NAND3 (N1513, N1492, N1479, N532);
not NOT1 (N1514, N1512);
not NOT1 (N1515, N1501);
or OR4 (N1516, N1488, N320, N937, N476);
xor XOR2 (N1517, N1510, N621);
and AND3 (N1518, N1489, N821, N310);
or OR3 (N1519, N1518, N980, N498);
and AND2 (N1520, N1519, N375);
buf BUF1 (N1521, N1513);
xor XOR2 (N1522, N1517, N914);
or OR4 (N1523, N1515, N561, N699, N320);
not NOT1 (N1524, N1520);
and AND4 (N1525, N1508, N773, N1147, N215);
not NOT1 (N1526, N1525);
not NOT1 (N1527, N1503);
not NOT1 (N1528, N1514);
xor XOR2 (N1529, N1527, N40);
nand NAND3 (N1530, N1511, N501, N827);
xor XOR2 (N1531, N1528, N854);
and AND3 (N1532, N1529, N1373, N1072);
buf BUF1 (N1533, N1504);
xor XOR2 (N1534, N1522, N503);
and AND4 (N1535, N1516, N1382, N175, N961);
nand NAND4 (N1536, N1532, N572, N323, N1137);
nand NAND2 (N1537, N1523, N1039);
nor NOR2 (N1538, N1524, N599);
buf BUF1 (N1539, N1526);
nor NOR2 (N1540, N1539, N1296);
xor XOR2 (N1541, N1538, N1065);
buf BUF1 (N1542, N1533);
nor NOR4 (N1543, N1535, N603, N870, N1020);
nand NAND2 (N1544, N1543, N1161);
and AND3 (N1545, N1534, N202, N673);
xor XOR2 (N1546, N1542, N1108);
and AND2 (N1547, N1546, N1186);
or OR4 (N1548, N1545, N74, N1358, N1041);
and AND2 (N1549, N1548, N1112);
xor XOR2 (N1550, N1537, N445);
xor XOR2 (N1551, N1547, N1384);
not NOT1 (N1552, N1551);
and AND3 (N1553, N1552, N904, N169);
or OR3 (N1554, N1521, N202, N70);
xor XOR2 (N1555, N1541, N1168);
not NOT1 (N1556, N1536);
xor XOR2 (N1557, N1554, N1397);
buf BUF1 (N1558, N1555);
nand NAND3 (N1559, N1550, N1550, N311);
and AND3 (N1560, N1531, N1096, N499);
or OR4 (N1561, N1556, N299, N286, N1122);
or OR4 (N1562, N1561, N256, N366, N655);
buf BUF1 (N1563, N1557);
and AND3 (N1564, N1530, N364, N862);
not NOT1 (N1565, N1560);
or OR3 (N1566, N1562, N1476, N753);
or OR3 (N1567, N1566, N367, N1143);
or OR3 (N1568, N1567, N396, N1158);
nand NAND3 (N1569, N1558, N299, N507);
nand NAND4 (N1570, N1553, N641, N1317, N1123);
nor NOR3 (N1571, N1559, N516, N1308);
nor NOR3 (N1572, N1570, N481, N241);
not NOT1 (N1573, N1572);
and AND3 (N1574, N1540, N406, N1357);
nand NAND3 (N1575, N1544, N1285, N36);
buf BUF1 (N1576, N1564);
and AND2 (N1577, N1565, N16);
not NOT1 (N1578, N1575);
not NOT1 (N1579, N1571);
and AND4 (N1580, N1569, N154, N367, N230);
nand NAND3 (N1581, N1577, N184, N303);
not NOT1 (N1582, N1580);
xor XOR2 (N1583, N1574, N662);
nand NAND2 (N1584, N1573, N368);
not NOT1 (N1585, N1578);
not NOT1 (N1586, N1581);
not NOT1 (N1587, N1549);
and AND4 (N1588, N1586, N1494, N980, N1353);
nor NOR2 (N1589, N1563, N886);
and AND2 (N1590, N1588, N73);
nand NAND2 (N1591, N1584, N1151);
xor XOR2 (N1592, N1590, N213);
or OR2 (N1593, N1582, N423);
nand NAND3 (N1594, N1592, N338, N612);
or OR3 (N1595, N1591, N687, N73);
or OR3 (N1596, N1568, N991, N50);
and AND2 (N1597, N1596, N1338);
not NOT1 (N1598, N1587);
xor XOR2 (N1599, N1585, N921);
not NOT1 (N1600, N1595);
xor XOR2 (N1601, N1576, N1260);
xor XOR2 (N1602, N1599, N720);
or OR3 (N1603, N1601, N10, N448);
or OR3 (N1604, N1583, N1501, N854);
or OR2 (N1605, N1589, N12);
xor XOR2 (N1606, N1593, N920);
and AND3 (N1607, N1605, N1012, N1497);
nand NAND4 (N1608, N1598, N21, N950, N346);
nor NOR4 (N1609, N1594, N1419, N379, N361);
not NOT1 (N1610, N1597);
xor XOR2 (N1611, N1600, N635);
or OR4 (N1612, N1610, N831, N379, N1377);
xor XOR2 (N1613, N1612, N714);
and AND4 (N1614, N1606, N280, N1380, N1404);
and AND4 (N1615, N1602, N1373, N1000, N379);
buf BUF1 (N1616, N1614);
not NOT1 (N1617, N1607);
buf BUF1 (N1618, N1608);
or OR4 (N1619, N1618, N1432, N1595, N862);
not NOT1 (N1620, N1617);
not NOT1 (N1621, N1615);
and AND2 (N1622, N1604, N393);
nor NOR3 (N1623, N1616, N53, N903);
buf BUF1 (N1624, N1623);
xor XOR2 (N1625, N1624, N1366);
and AND4 (N1626, N1603, N500, N624, N898);
and AND2 (N1627, N1619, N526);
or OR3 (N1628, N1622, N232, N140);
buf BUF1 (N1629, N1611);
nand NAND4 (N1630, N1579, N1594, N682, N1629);
not NOT1 (N1631, N1378);
not NOT1 (N1632, N1613);
and AND2 (N1633, N1626, N1600);
and AND4 (N1634, N1632, N280, N383, N860);
nand NAND4 (N1635, N1625, N235, N675, N1076);
and AND2 (N1636, N1634, N24);
xor XOR2 (N1637, N1633, N321);
and AND2 (N1638, N1609, N134);
nand NAND4 (N1639, N1620, N614, N1208, N880);
not NOT1 (N1640, N1639);
xor XOR2 (N1641, N1640, N278);
not NOT1 (N1642, N1630);
buf BUF1 (N1643, N1637);
or OR3 (N1644, N1642, N1360, N768);
buf BUF1 (N1645, N1621);
not NOT1 (N1646, N1645);
nand NAND2 (N1647, N1627, N386);
nand NAND2 (N1648, N1638, N1300);
nor NOR2 (N1649, N1636, N544);
buf BUF1 (N1650, N1628);
and AND4 (N1651, N1646, N231, N252, N1344);
nand NAND4 (N1652, N1647, N1272, N911, N365);
not NOT1 (N1653, N1649);
nand NAND2 (N1654, N1652, N1395);
buf BUF1 (N1655, N1635);
nor NOR2 (N1656, N1650, N1259);
xor XOR2 (N1657, N1654, N1124);
nand NAND4 (N1658, N1657, N1296, N970, N1205);
nor NOR4 (N1659, N1658, N1225, N224, N876);
buf BUF1 (N1660, N1656);
xor XOR2 (N1661, N1651, N20);
xor XOR2 (N1662, N1660, N1433);
xor XOR2 (N1663, N1655, N275);
buf BUF1 (N1664, N1643);
or OR4 (N1665, N1641, N995, N34, N879);
and AND2 (N1666, N1663, N245);
and AND2 (N1667, N1662, N1391);
buf BUF1 (N1668, N1644);
not NOT1 (N1669, N1664);
buf BUF1 (N1670, N1648);
nor NOR2 (N1671, N1659, N844);
nand NAND2 (N1672, N1671, N1121);
xor XOR2 (N1673, N1669, N1082);
nand NAND4 (N1674, N1631, N401, N734, N1383);
or OR4 (N1675, N1674, N1193, N1279, N1316);
xor XOR2 (N1676, N1675, N800);
or OR4 (N1677, N1667, N145, N800, N1511);
nand NAND3 (N1678, N1661, N1228, N518);
buf BUF1 (N1679, N1677);
nor NOR3 (N1680, N1673, N203, N1139);
nor NOR2 (N1681, N1670, N183);
buf BUF1 (N1682, N1666);
nor NOR4 (N1683, N1653, N496, N1041, N946);
not NOT1 (N1684, N1678);
xor XOR2 (N1685, N1681, N1600);
and AND3 (N1686, N1676, N143, N1499);
and AND2 (N1687, N1686, N1587);
nor NOR4 (N1688, N1672, N186, N1487, N865);
nand NAND3 (N1689, N1682, N1678, N1287);
not NOT1 (N1690, N1668);
nand NAND4 (N1691, N1679, N342, N707, N1602);
nand NAND4 (N1692, N1665, N1364, N1379, N855);
nand NAND3 (N1693, N1689, N874, N1479);
or OR3 (N1694, N1690, N956, N1293);
or OR2 (N1695, N1688, N427);
or OR2 (N1696, N1693, N402);
not NOT1 (N1697, N1685);
or OR3 (N1698, N1696, N986, N912);
xor XOR2 (N1699, N1694, N126);
xor XOR2 (N1700, N1680, N1054);
xor XOR2 (N1701, N1698, N103);
or OR2 (N1702, N1684, N279);
or OR3 (N1703, N1699, N860, N326);
not NOT1 (N1704, N1703);
and AND3 (N1705, N1702, N1161, N247);
nor NOR2 (N1706, N1691, N488);
buf BUF1 (N1707, N1701);
xor XOR2 (N1708, N1704, N394);
xor XOR2 (N1709, N1708, N12);
buf BUF1 (N1710, N1700);
nand NAND3 (N1711, N1683, N1663, N1668);
xor XOR2 (N1712, N1705, N709);
and AND2 (N1713, N1712, N295);
nor NOR4 (N1714, N1695, N1217, N1394, N1225);
nor NOR4 (N1715, N1697, N1076, N296, N1173);
not NOT1 (N1716, N1709);
buf BUF1 (N1717, N1711);
nor NOR4 (N1718, N1713, N33, N1075, N1106);
xor XOR2 (N1719, N1714, N1355);
not NOT1 (N1720, N1710);
xor XOR2 (N1721, N1717, N1059);
not NOT1 (N1722, N1719);
nand NAND3 (N1723, N1721, N1060, N1661);
xor XOR2 (N1724, N1715, N119);
xor XOR2 (N1725, N1718, N1108);
nand NAND4 (N1726, N1687, N1470, N964, N456);
buf BUF1 (N1727, N1722);
and AND2 (N1728, N1725, N1341);
and AND3 (N1729, N1723, N1098, N325);
xor XOR2 (N1730, N1716, N1508);
nand NAND2 (N1731, N1730, N309);
nor NOR4 (N1732, N1729, N1609, N1083, N281);
nor NOR2 (N1733, N1724, N957);
and AND2 (N1734, N1728, N176);
or OR4 (N1735, N1707, N522, N778, N384);
and AND3 (N1736, N1692, N511, N1017);
and AND2 (N1737, N1733, N234);
nor NOR4 (N1738, N1736, N188, N901, N661);
and AND4 (N1739, N1737, N1116, N1251, N1017);
and AND4 (N1740, N1727, N1094, N1603, N1554);
buf BUF1 (N1741, N1731);
xor XOR2 (N1742, N1732, N555);
or OR2 (N1743, N1720, N803);
nand NAND2 (N1744, N1740, N1128);
nor NOR4 (N1745, N1706, N1293, N1121, N201);
xor XOR2 (N1746, N1741, N768);
not NOT1 (N1747, N1744);
nor NOR4 (N1748, N1747, N1499, N691, N479);
nand NAND2 (N1749, N1739, N892);
nor NOR3 (N1750, N1742, N1340, N1108);
nand NAND2 (N1751, N1748, N1038);
xor XOR2 (N1752, N1735, N799);
not NOT1 (N1753, N1751);
and AND4 (N1754, N1746, N1212, N401, N200);
buf BUF1 (N1755, N1750);
and AND4 (N1756, N1745, N1471, N1212, N1345);
nor NOR2 (N1757, N1726, N816);
nor NOR2 (N1758, N1738, N919);
not NOT1 (N1759, N1752);
buf BUF1 (N1760, N1734);
buf BUF1 (N1761, N1758);
and AND3 (N1762, N1756, N435, N233);
xor XOR2 (N1763, N1762, N648);
not NOT1 (N1764, N1763);
or OR2 (N1765, N1754, N1609);
nor NOR3 (N1766, N1755, N1502, N1119);
nand NAND3 (N1767, N1764, N1332, N1540);
or OR4 (N1768, N1765, N359, N1124, N72);
nor NOR3 (N1769, N1766, N1257, N654);
xor XOR2 (N1770, N1759, N86);
xor XOR2 (N1771, N1768, N1435);
xor XOR2 (N1772, N1761, N1106);
nor NOR4 (N1773, N1743, N1156, N293, N381);
nand NAND2 (N1774, N1749, N822);
xor XOR2 (N1775, N1769, N1113);
xor XOR2 (N1776, N1774, N1008);
buf BUF1 (N1777, N1757);
or OR3 (N1778, N1775, N122, N1346);
nand NAND3 (N1779, N1773, N606, N1041);
nand NAND4 (N1780, N1778, N1753, N394, N1577);
buf BUF1 (N1781, N1032);
and AND2 (N1782, N1760, N1448);
or OR2 (N1783, N1771, N1743);
buf BUF1 (N1784, N1779);
nor NOR2 (N1785, N1784, N761);
or OR4 (N1786, N1767, N1745, N1294, N1340);
and AND4 (N1787, N1780, N1327, N568, N463);
or OR3 (N1788, N1781, N1387, N531);
or OR3 (N1789, N1777, N1502, N117);
not NOT1 (N1790, N1782);
buf BUF1 (N1791, N1790);
or OR4 (N1792, N1783, N1101, N383, N456);
nor NOR3 (N1793, N1786, N1462, N1534);
nand NAND4 (N1794, N1776, N820, N75, N1327);
and AND2 (N1795, N1770, N1567);
xor XOR2 (N1796, N1794, N810);
xor XOR2 (N1797, N1788, N103);
and AND2 (N1798, N1789, N416);
and AND3 (N1799, N1793, N375, N776);
xor XOR2 (N1800, N1792, N102);
buf BUF1 (N1801, N1797);
and AND4 (N1802, N1800, N145, N649, N801);
and AND3 (N1803, N1772, N942, N18);
and AND4 (N1804, N1795, N1306, N768, N406);
xor XOR2 (N1805, N1803, N800);
or OR4 (N1806, N1801, N732, N708, N1391);
buf BUF1 (N1807, N1796);
xor XOR2 (N1808, N1787, N478);
nand NAND2 (N1809, N1785, N1167);
xor XOR2 (N1810, N1799, N395);
not NOT1 (N1811, N1809);
not NOT1 (N1812, N1804);
xor XOR2 (N1813, N1808, N1311);
not NOT1 (N1814, N1813);
or OR2 (N1815, N1814, N1647);
nand NAND2 (N1816, N1815, N788);
or OR3 (N1817, N1807, N1423, N1796);
buf BUF1 (N1818, N1806);
xor XOR2 (N1819, N1791, N447);
nor NOR4 (N1820, N1816, N270, N53, N491);
buf BUF1 (N1821, N1798);
and AND4 (N1822, N1818, N729, N1151, N648);
buf BUF1 (N1823, N1811);
not NOT1 (N1824, N1817);
not NOT1 (N1825, N1820);
nor NOR3 (N1826, N1823, N1770, N1086);
nand NAND2 (N1827, N1812, N1248);
and AND3 (N1828, N1826, N1066, N1025);
xor XOR2 (N1829, N1819, N1196);
or OR3 (N1830, N1829, N1521, N1693);
nor NOR4 (N1831, N1830, N1140, N56, N1068);
and AND4 (N1832, N1805, N303, N798, N1213);
not NOT1 (N1833, N1828);
and AND3 (N1834, N1833, N1190, N1644);
xor XOR2 (N1835, N1822, N546);
nand NAND4 (N1836, N1821, N282, N1025, N93);
nand NAND3 (N1837, N1836, N285, N438);
nor NOR3 (N1838, N1832, N484, N1277);
buf BUF1 (N1839, N1837);
not NOT1 (N1840, N1824);
nor NOR3 (N1841, N1840, N1592, N531);
nor NOR3 (N1842, N1831, N1735, N203);
or OR4 (N1843, N1839, N1782, N137, N628);
or OR3 (N1844, N1838, N942, N1286);
nor NOR4 (N1845, N1802, N15, N1829, N564);
xor XOR2 (N1846, N1834, N1777);
not NOT1 (N1847, N1844);
or OR4 (N1848, N1841, N1234, N244, N1728);
nand NAND3 (N1849, N1835, N1142, N230);
not NOT1 (N1850, N1849);
not NOT1 (N1851, N1810);
not NOT1 (N1852, N1846);
not NOT1 (N1853, N1852);
nand NAND2 (N1854, N1825, N878);
or OR2 (N1855, N1842, N138);
xor XOR2 (N1856, N1851, N42);
xor XOR2 (N1857, N1843, N1297);
buf BUF1 (N1858, N1848);
nand NAND2 (N1859, N1858, N130);
nor NOR3 (N1860, N1850, N1323, N1013);
and AND2 (N1861, N1860, N309);
xor XOR2 (N1862, N1853, N417);
or OR2 (N1863, N1854, N1463);
or OR2 (N1864, N1855, N1551);
nand NAND2 (N1865, N1827, N1124);
nor NOR3 (N1866, N1864, N1242, N509);
or OR3 (N1867, N1857, N681, N848);
nor NOR3 (N1868, N1865, N299, N849);
buf BUF1 (N1869, N1866);
xor XOR2 (N1870, N1867, N594);
and AND2 (N1871, N1859, N1206);
nor NOR2 (N1872, N1862, N1280);
nor NOR2 (N1873, N1847, N181);
nor NOR4 (N1874, N1868, N776, N994, N1019);
xor XOR2 (N1875, N1871, N1155);
nor NOR3 (N1876, N1872, N1207, N939);
or OR2 (N1877, N1845, N1672);
buf BUF1 (N1878, N1869);
and AND3 (N1879, N1878, N73, N901);
xor XOR2 (N1880, N1879, N82);
or OR4 (N1881, N1870, N328, N1005, N1175);
xor XOR2 (N1882, N1874, N16);
xor XOR2 (N1883, N1877, N1849);
nand NAND4 (N1884, N1861, N865, N1054, N454);
buf BUF1 (N1885, N1882);
or OR2 (N1886, N1885, N373);
nand NAND4 (N1887, N1886, N775, N1105, N788);
and AND3 (N1888, N1863, N428, N719);
not NOT1 (N1889, N1883);
nand NAND4 (N1890, N1856, N383, N1218, N833);
nor NOR2 (N1891, N1880, N1583);
xor XOR2 (N1892, N1884, N932);
or OR4 (N1893, N1875, N340, N1696, N226);
buf BUF1 (N1894, N1873);
nand NAND4 (N1895, N1881, N1033, N39, N102);
nor NOR2 (N1896, N1893, N264);
nand NAND2 (N1897, N1889, N188);
xor XOR2 (N1898, N1895, N43);
and AND4 (N1899, N1887, N1084, N185, N680);
xor XOR2 (N1900, N1896, N25);
not NOT1 (N1901, N1899);
not NOT1 (N1902, N1898);
buf BUF1 (N1903, N1876);
or OR3 (N1904, N1897, N229, N1262);
xor XOR2 (N1905, N1903, N196);
nor NOR2 (N1906, N1900, N142);
not NOT1 (N1907, N1888);
not NOT1 (N1908, N1891);
xor XOR2 (N1909, N1894, N1857);
nand NAND2 (N1910, N1902, N269);
buf BUF1 (N1911, N1906);
and AND2 (N1912, N1905, N762);
not NOT1 (N1913, N1890);
buf BUF1 (N1914, N1911);
nand NAND3 (N1915, N1914, N1716, N1016);
xor XOR2 (N1916, N1912, N300);
nor NOR4 (N1917, N1909, N1905, N1783, N1895);
xor XOR2 (N1918, N1907, N1244);
buf BUF1 (N1919, N1918);
nand NAND2 (N1920, N1916, N1121);
nor NOR2 (N1921, N1910, N489);
xor XOR2 (N1922, N1919, N824);
nand NAND4 (N1923, N1922, N975, N217, N570);
not NOT1 (N1924, N1901);
nand NAND3 (N1925, N1913, N1750, N1579);
nand NAND3 (N1926, N1920, N961, N956);
and AND4 (N1927, N1921, N1534, N520, N1623);
and AND2 (N1928, N1926, N1340);
buf BUF1 (N1929, N1923);
xor XOR2 (N1930, N1927, N1554);
or OR3 (N1931, N1892, N1085, N1808);
and AND2 (N1932, N1929, N1781);
xor XOR2 (N1933, N1932, N967);
or OR3 (N1934, N1930, N346, N1110);
and AND2 (N1935, N1931, N699);
not NOT1 (N1936, N1908);
buf BUF1 (N1937, N1936);
or OR4 (N1938, N1935, N1292, N1709, N115);
xor XOR2 (N1939, N1938, N1848);
nor NOR4 (N1940, N1928, N1590, N553, N1278);
xor XOR2 (N1941, N1940, N1083);
buf BUF1 (N1942, N1924);
nor NOR3 (N1943, N1939, N1174, N985);
nor NOR2 (N1944, N1934, N886);
or OR3 (N1945, N1944, N1852, N157);
xor XOR2 (N1946, N1904, N1349);
or OR3 (N1947, N1942, N779, N1201);
and AND3 (N1948, N1945, N456, N576);
xor XOR2 (N1949, N1917, N1395);
nand NAND3 (N1950, N1925, N44, N917);
not NOT1 (N1951, N1941);
or OR3 (N1952, N1950, N1595, N1303);
nand NAND4 (N1953, N1946, N1494, N488, N353);
nand NAND2 (N1954, N1915, N271);
or OR3 (N1955, N1933, N1160, N357);
buf BUF1 (N1956, N1952);
buf BUF1 (N1957, N1948);
or OR3 (N1958, N1951, N682, N882);
not NOT1 (N1959, N1956);
not NOT1 (N1960, N1937);
buf BUF1 (N1961, N1947);
nor NOR2 (N1962, N1953, N502);
and AND4 (N1963, N1955, N1407, N1554, N1547);
or OR4 (N1964, N1963, N976, N606, N1485);
or OR2 (N1965, N1949, N360);
or OR2 (N1966, N1958, N1388);
not NOT1 (N1967, N1954);
buf BUF1 (N1968, N1957);
or OR2 (N1969, N1959, N276);
not NOT1 (N1970, N1965);
nand NAND3 (N1971, N1966, N1925, N316);
buf BUF1 (N1972, N1961);
xor XOR2 (N1973, N1972, N68);
nand NAND2 (N1974, N1970, N525);
not NOT1 (N1975, N1968);
nand NAND4 (N1976, N1969, N1077, N1297, N513);
not NOT1 (N1977, N1976);
not NOT1 (N1978, N1977);
nor NOR3 (N1979, N1962, N1479, N1644);
not NOT1 (N1980, N1971);
buf BUF1 (N1981, N1974);
or OR4 (N1982, N1973, N123, N1789, N1323);
nand NAND4 (N1983, N1980, N975, N200, N1542);
and AND4 (N1984, N1960, N245, N654, N296);
xor XOR2 (N1985, N1975, N1290);
nor NOR2 (N1986, N1978, N595);
xor XOR2 (N1987, N1979, N152);
xor XOR2 (N1988, N1943, N1606);
xor XOR2 (N1989, N1988, N1610);
buf BUF1 (N1990, N1987);
or OR3 (N1991, N1984, N1887, N382);
nor NOR4 (N1992, N1989, N953, N1560, N45);
nand NAND2 (N1993, N1967, N851);
xor XOR2 (N1994, N1964, N1266);
buf BUF1 (N1995, N1983);
or OR3 (N1996, N1992, N1994, N1507);
or OR4 (N1997, N1564, N1583, N1297, N1159);
xor XOR2 (N1998, N1997, N1833);
nand NAND2 (N1999, N1982, N1288);
not NOT1 (N2000, N1985);
buf BUF1 (N2001, N1986);
buf BUF1 (N2002, N1996);
or OR2 (N2003, N2001, N1560);
not NOT1 (N2004, N1993);
or OR3 (N2005, N1995, N1879, N339);
or OR3 (N2006, N2004, N1296, N181);
buf BUF1 (N2007, N2003);
nor NOR3 (N2008, N1998, N1034, N396);
or OR2 (N2009, N2007, N1343);
xor XOR2 (N2010, N1999, N1826);
or OR2 (N2011, N2000, N1889);
buf BUF1 (N2012, N2002);
and AND2 (N2013, N2010, N886);
or OR4 (N2014, N2012, N1466, N1048, N903);
nor NOR3 (N2015, N1991, N377, N1051);
and AND2 (N2016, N2009, N100);
or OR3 (N2017, N2006, N1445, N171);
and AND2 (N2018, N2005, N1311);
nor NOR4 (N2019, N2017, N1194, N482, N1695);
buf BUF1 (N2020, N2014);
nand NAND2 (N2021, N2016, N677);
xor XOR2 (N2022, N2019, N1117);
xor XOR2 (N2023, N2020, N1671);
nand NAND2 (N2024, N1981, N228);
nor NOR3 (N2025, N2024, N324, N1832);
xor XOR2 (N2026, N2018, N67);
xor XOR2 (N2027, N2011, N670);
nor NOR4 (N2028, N2013, N1449, N139, N420);
or OR2 (N2029, N2026, N764);
buf BUF1 (N2030, N1990);
xor XOR2 (N2031, N2015, N1900);
or OR4 (N2032, N2030, N1146, N1493, N402);
nand NAND3 (N2033, N2028, N336, N627);
not NOT1 (N2034, N2033);
xor XOR2 (N2035, N2029, N1933);
and AND2 (N2036, N2022, N1087);
xor XOR2 (N2037, N2023, N1443);
and AND2 (N2038, N2032, N1052);
or OR4 (N2039, N2038, N66, N1805, N76);
or OR4 (N2040, N2035, N1754, N1111, N541);
and AND2 (N2041, N2008, N1613);
buf BUF1 (N2042, N2041);
nor NOR3 (N2043, N2037, N1394, N837);
buf BUF1 (N2044, N2040);
not NOT1 (N2045, N2025);
not NOT1 (N2046, N2031);
and AND4 (N2047, N2045, N1884, N1346, N1867);
nand NAND2 (N2048, N2044, N1113);
nor NOR3 (N2049, N2034, N1288, N1892);
nor NOR3 (N2050, N2039, N1470, N366);
or OR4 (N2051, N2036, N1779, N1415, N1030);
not NOT1 (N2052, N2047);
and AND2 (N2053, N2042, N836);
nor NOR4 (N2054, N2046, N953, N1586, N1633);
and AND2 (N2055, N2051, N1926);
or OR3 (N2056, N2043, N394, N443);
not NOT1 (N2057, N2049);
and AND4 (N2058, N2055, N1677, N738, N1198);
or OR4 (N2059, N2054, N76, N260, N1323);
not NOT1 (N2060, N2048);
and AND2 (N2061, N2053, N938);
nor NOR3 (N2062, N2061, N1397, N835);
buf BUF1 (N2063, N2052);
nand NAND2 (N2064, N2056, N1347);
xor XOR2 (N2065, N2059, N147);
or OR4 (N2066, N2058, N1677, N848, N1614);
buf BUF1 (N2067, N2027);
and AND4 (N2068, N2021, N677, N1619, N75);
not NOT1 (N2069, N2063);
nor NOR2 (N2070, N2050, N337);
nor NOR3 (N2071, N2060, N1653, N1487);
and AND2 (N2072, N2070, N1106);
buf BUF1 (N2073, N2068);
buf BUF1 (N2074, N2062);
nand NAND2 (N2075, N2066, N1979);
and AND3 (N2076, N2071, N1506, N1509);
xor XOR2 (N2077, N2067, N926);
not NOT1 (N2078, N2075);
buf BUF1 (N2079, N2064);
and AND2 (N2080, N2079, N1813);
not NOT1 (N2081, N2072);
nand NAND4 (N2082, N2074, N1824, N737, N1800);
nor NOR4 (N2083, N2076, N1153, N1545, N1397);
or OR4 (N2084, N2083, N1978, N1629, N356);
or OR4 (N2085, N2081, N1531, N1978, N188);
nor NOR4 (N2086, N2069, N6, N1664, N1667);
nor NOR2 (N2087, N2065, N155);
xor XOR2 (N2088, N2085, N1735);
buf BUF1 (N2089, N2086);
nor NOR3 (N2090, N2082, N443, N1035);
xor XOR2 (N2091, N2073, N399);
buf BUF1 (N2092, N2084);
xor XOR2 (N2093, N2077, N1993);
nor NOR2 (N2094, N2091, N1044);
buf BUF1 (N2095, N2094);
xor XOR2 (N2096, N2078, N2064);
and AND4 (N2097, N2092, N2060, N975, N744);
buf BUF1 (N2098, N2088);
and AND2 (N2099, N2098, N1308);
not NOT1 (N2100, N2089);
buf BUF1 (N2101, N2057);
nor NOR4 (N2102, N2097, N1187, N1462, N1071);
nand NAND2 (N2103, N2096, N1380);
nor NOR3 (N2104, N2095, N1735, N667);
or OR4 (N2105, N2103, N1675, N1322, N1139);
nand NAND2 (N2106, N2093, N963);
nor NOR3 (N2107, N2106, N1210, N638);
xor XOR2 (N2108, N2090, N1703);
nor NOR4 (N2109, N2102, N1197, N1892, N1861);
xor XOR2 (N2110, N2105, N892);
and AND3 (N2111, N2108, N168, N1138);
buf BUF1 (N2112, N2104);
xor XOR2 (N2113, N2107, N363);
xor XOR2 (N2114, N2113, N388);
nor NOR4 (N2115, N2111, N454, N1832, N1273);
nand NAND4 (N2116, N2100, N874, N1552, N822);
nand NAND2 (N2117, N2116, N344);
nand NAND3 (N2118, N2109, N1268, N1705);
not NOT1 (N2119, N2099);
nor NOR4 (N2120, N2080, N891, N583, N244);
buf BUF1 (N2121, N2118);
and AND2 (N2122, N2110, N310);
xor XOR2 (N2123, N2101, N705);
or OR3 (N2124, N2119, N1093, N1483);
xor XOR2 (N2125, N2114, N651);
nand NAND4 (N2126, N2124, N1111, N344, N229);
not NOT1 (N2127, N2123);
not NOT1 (N2128, N2122);
and AND4 (N2129, N2127, N459, N181, N1227);
buf BUF1 (N2130, N2117);
xor XOR2 (N2131, N2130, N273);
xor XOR2 (N2132, N2115, N1452);
not NOT1 (N2133, N2131);
not NOT1 (N2134, N2128);
not NOT1 (N2135, N2121);
not NOT1 (N2136, N2135);
buf BUF1 (N2137, N2125);
and AND3 (N2138, N2136, N1763, N1318);
nand NAND2 (N2139, N2137, N421);
nand NAND4 (N2140, N2134, N542, N1440, N514);
or OR4 (N2141, N2129, N1776, N732, N1466);
or OR4 (N2142, N2132, N704, N1097, N1259);
nor NOR3 (N2143, N2126, N980, N1526);
and AND4 (N2144, N2112, N893, N1668, N1573);
not NOT1 (N2145, N2138);
nand NAND4 (N2146, N2140, N1287, N1416, N1770);
buf BUF1 (N2147, N2145);
nand NAND4 (N2148, N2144, N1553, N797, N1351);
not NOT1 (N2149, N2087);
not NOT1 (N2150, N2120);
nor NOR4 (N2151, N2141, N741, N506, N2051);
nor NOR4 (N2152, N2146, N2032, N1693, N990);
nand NAND4 (N2153, N2133, N161, N1292, N1308);
nor NOR2 (N2154, N2148, N1147);
nand NAND2 (N2155, N2142, N11);
and AND3 (N2156, N2150, N1441, N1953);
and AND2 (N2157, N2152, N1616);
nor NOR4 (N2158, N2143, N2110, N119, N2098);
nor NOR3 (N2159, N2153, N373, N1813);
xor XOR2 (N2160, N2151, N1007);
xor XOR2 (N2161, N2155, N715);
nor NOR2 (N2162, N2147, N292);
and AND2 (N2163, N2139, N474);
nand NAND3 (N2164, N2159, N1344, N1203);
nor NOR3 (N2165, N2160, N393, N1728);
or OR4 (N2166, N2165, N1521, N843, N1058);
xor XOR2 (N2167, N2158, N1855);
nor NOR4 (N2168, N2154, N408, N2046, N942);
nor NOR4 (N2169, N2157, N236, N1547, N1902);
buf BUF1 (N2170, N2168);
nor NOR4 (N2171, N2166, N2138, N378, N812);
buf BUF1 (N2172, N2169);
nor NOR4 (N2173, N2167, N125, N431, N1975);
buf BUF1 (N2174, N2172);
xor XOR2 (N2175, N2171, N1542);
nand NAND4 (N2176, N2174, N933, N326, N1562);
and AND2 (N2177, N2176, N772);
not NOT1 (N2178, N2175);
not NOT1 (N2179, N2156);
and AND2 (N2180, N2178, N401);
or OR2 (N2181, N2149, N1266);
and AND4 (N2182, N2162, N544, N799, N91);
and AND3 (N2183, N2177, N1087, N1971);
nand NAND4 (N2184, N2182, N300, N20, N1367);
xor XOR2 (N2185, N2163, N659);
or OR4 (N2186, N2183, N2086, N701, N147);
nor NOR3 (N2187, N2173, N2000, N2062);
buf BUF1 (N2188, N2180);
and AND3 (N2189, N2185, N1437, N157);
buf BUF1 (N2190, N2164);
xor XOR2 (N2191, N2181, N1986);
nor NOR4 (N2192, N2189, N1331, N1520, N2129);
not NOT1 (N2193, N2170);
not NOT1 (N2194, N2187);
and AND4 (N2195, N2191, N53, N2066, N102);
not NOT1 (N2196, N2179);
not NOT1 (N2197, N2194);
nor NOR4 (N2198, N2161, N1246, N928, N1908);
or OR3 (N2199, N2193, N335, N2136);
nor NOR3 (N2200, N2198, N675, N50);
nor NOR3 (N2201, N2190, N202, N410);
buf BUF1 (N2202, N2184);
nand NAND2 (N2203, N2195, N1085);
buf BUF1 (N2204, N2192);
xor XOR2 (N2205, N2202, N652);
nand NAND2 (N2206, N2201, N1726);
and AND4 (N2207, N2205, N1605, N448, N828);
buf BUF1 (N2208, N2207);
buf BUF1 (N2209, N2186);
and AND2 (N2210, N2208, N871);
or OR3 (N2211, N2188, N35, N1985);
or OR4 (N2212, N2210, N988, N1492, N1788);
or OR3 (N2213, N2212, N663, N956);
xor XOR2 (N2214, N2204, N798);
or OR3 (N2215, N2209, N167, N1259);
and AND4 (N2216, N2200, N1950, N1911, N646);
buf BUF1 (N2217, N2215);
or OR4 (N2218, N2211, N452, N963, N1270);
nor NOR3 (N2219, N2214, N1164, N654);
and AND4 (N2220, N2206, N1201, N691, N1993);
nor NOR2 (N2221, N2218, N1602);
or OR2 (N2222, N2219, N1023);
nor NOR2 (N2223, N2196, N455);
nand NAND2 (N2224, N2197, N1307);
not NOT1 (N2225, N2224);
buf BUF1 (N2226, N2216);
nand NAND2 (N2227, N2222, N1017);
or OR3 (N2228, N2225, N1697, N824);
buf BUF1 (N2229, N2228);
and AND3 (N2230, N2203, N1100, N2118);
or OR4 (N2231, N2217, N353, N1309, N896);
not NOT1 (N2232, N2227);
buf BUF1 (N2233, N2232);
xor XOR2 (N2234, N2226, N1707);
or OR2 (N2235, N2234, N950);
nand NAND3 (N2236, N2213, N519, N2069);
xor XOR2 (N2237, N2235, N720);
buf BUF1 (N2238, N2231);
buf BUF1 (N2239, N2237);
and AND4 (N2240, N2221, N649, N1167, N42);
xor XOR2 (N2241, N2238, N1880);
xor XOR2 (N2242, N2223, N1746);
nand NAND2 (N2243, N2240, N1445);
and AND4 (N2244, N2233, N1092, N1544, N1337);
nand NAND3 (N2245, N2236, N1179, N883);
not NOT1 (N2246, N2243);
and AND3 (N2247, N2246, N1599, N1098);
xor XOR2 (N2248, N2245, N1532);
buf BUF1 (N2249, N2239);
and AND2 (N2250, N2249, N1473);
nor NOR4 (N2251, N2244, N2081, N1646, N1956);
buf BUF1 (N2252, N2229);
and AND2 (N2253, N2250, N1278);
not NOT1 (N2254, N2253);
or OR4 (N2255, N2199, N1196, N1673, N766);
buf BUF1 (N2256, N2241);
xor XOR2 (N2257, N2254, N941);
xor XOR2 (N2258, N2255, N463);
or OR3 (N2259, N2257, N368, N914);
xor XOR2 (N2260, N2248, N933);
nand NAND3 (N2261, N2230, N1434, N1029);
nand NAND3 (N2262, N2258, N337, N1288);
not NOT1 (N2263, N2242);
not NOT1 (N2264, N2220);
nor NOR2 (N2265, N2264, N1523);
buf BUF1 (N2266, N2247);
nor NOR2 (N2267, N2265, N2066);
not NOT1 (N2268, N2256);
not NOT1 (N2269, N2260);
and AND4 (N2270, N2252, N1846, N193, N906);
not NOT1 (N2271, N2251);
nand NAND2 (N2272, N2270, N2126);
and AND3 (N2273, N2263, N746, N373);
buf BUF1 (N2274, N2266);
nand NAND4 (N2275, N2268, N748, N1913, N1086);
xor XOR2 (N2276, N2271, N1737);
buf BUF1 (N2277, N2274);
buf BUF1 (N2278, N2272);
buf BUF1 (N2279, N2275);
not NOT1 (N2280, N2269);
nor NOR4 (N2281, N2279, N281, N488, N1692);
or OR2 (N2282, N2267, N577);
buf BUF1 (N2283, N2277);
buf BUF1 (N2284, N2259);
xor XOR2 (N2285, N2262, N688);
not NOT1 (N2286, N2285);
buf BUF1 (N2287, N2282);
nand NAND3 (N2288, N2281, N1969, N1345);
nand NAND2 (N2289, N2284, N238);
nor NOR3 (N2290, N2283, N1189, N655);
or OR4 (N2291, N2273, N1355, N1188, N2013);
not NOT1 (N2292, N2290);
or OR2 (N2293, N2288, N1181);
nand NAND4 (N2294, N2292, N911, N2248, N1368);
nor NOR3 (N2295, N2280, N1127, N550);
buf BUF1 (N2296, N2261);
not NOT1 (N2297, N2289);
not NOT1 (N2298, N2278);
not NOT1 (N2299, N2298);
and AND3 (N2300, N2287, N1256, N50);
xor XOR2 (N2301, N2286, N2224);
xor XOR2 (N2302, N2301, N1286);
and AND2 (N2303, N2291, N566);
nor NOR2 (N2304, N2293, N506);
or OR3 (N2305, N2297, N1937, N228);
nor NOR4 (N2306, N2300, N1781, N1688, N113);
nand NAND2 (N2307, N2304, N345);
nor NOR3 (N2308, N2296, N1255, N936);
buf BUF1 (N2309, N2299);
nor NOR2 (N2310, N2309, N215);
nor NOR4 (N2311, N2303, N1071, N712, N36);
buf BUF1 (N2312, N2310);
xor XOR2 (N2313, N2307, N1333);
xor XOR2 (N2314, N2294, N1588);
buf BUF1 (N2315, N2312);
nor NOR4 (N2316, N2306, N1764, N564, N1501);
or OR2 (N2317, N2302, N937);
xor XOR2 (N2318, N2316, N995);
nand NAND2 (N2319, N2305, N1839);
nand NAND3 (N2320, N2319, N1983, N1646);
and AND3 (N2321, N2315, N1048, N281);
and AND3 (N2322, N2318, N1592, N1598);
buf BUF1 (N2323, N2308);
and AND4 (N2324, N2313, N160, N1112, N771);
xor XOR2 (N2325, N2295, N255);
nand NAND4 (N2326, N2322, N1870, N2028, N1613);
nor NOR4 (N2327, N2276, N781, N1514, N871);
not NOT1 (N2328, N2317);
nor NOR3 (N2329, N2326, N1721, N1562);
buf BUF1 (N2330, N2321);
nor NOR3 (N2331, N2323, N140, N1849);
and AND4 (N2332, N2331, N334, N1410, N2104);
xor XOR2 (N2333, N2314, N266);
nand NAND2 (N2334, N2328, N154);
xor XOR2 (N2335, N2329, N224);
nor NOR3 (N2336, N2320, N43, N668);
buf BUF1 (N2337, N2325);
not NOT1 (N2338, N2332);
buf BUF1 (N2339, N2335);
or OR3 (N2340, N2334, N1419, N1625);
xor XOR2 (N2341, N2311, N1393);
or OR4 (N2342, N2336, N1646, N525, N877);
buf BUF1 (N2343, N2338);
nor NOR3 (N2344, N2339, N2329, N462);
not NOT1 (N2345, N2330);
nor NOR2 (N2346, N2345, N130);
not NOT1 (N2347, N2340);
xor XOR2 (N2348, N2344, N1151);
xor XOR2 (N2349, N2327, N724);
nand NAND4 (N2350, N2347, N2102, N80, N1600);
xor XOR2 (N2351, N2333, N1698);
not NOT1 (N2352, N2349);
and AND3 (N2353, N2352, N160, N1516);
or OR2 (N2354, N2343, N831);
buf BUF1 (N2355, N2353);
and AND3 (N2356, N2348, N358, N78);
not NOT1 (N2357, N2356);
and AND4 (N2358, N2351, N1644, N1325, N226);
buf BUF1 (N2359, N2341);
xor XOR2 (N2360, N2346, N2104);
not NOT1 (N2361, N2357);
nor NOR2 (N2362, N2354, N866);
not NOT1 (N2363, N2342);
nand NAND2 (N2364, N2337, N1895);
xor XOR2 (N2365, N2361, N857);
not NOT1 (N2366, N2363);
buf BUF1 (N2367, N2324);
nand NAND2 (N2368, N2366, N1987);
and AND4 (N2369, N2365, N1628, N77, N759);
xor XOR2 (N2370, N2350, N1948);
nand NAND3 (N2371, N2364, N858, N1431);
and AND3 (N2372, N2369, N233, N2052);
nand NAND4 (N2373, N2362, N152, N1194, N958);
or OR2 (N2374, N2360, N1615);
nor NOR3 (N2375, N2370, N49, N1250);
and AND3 (N2376, N2368, N1574, N333);
or OR4 (N2377, N2375, N1076, N2041, N1637);
xor XOR2 (N2378, N2371, N1266);
and AND2 (N2379, N2355, N341);
and AND4 (N2380, N2373, N1604, N984, N662);
nor NOR2 (N2381, N2372, N1870);
xor XOR2 (N2382, N2374, N403);
nand NAND2 (N2383, N2382, N351);
buf BUF1 (N2384, N2376);
not NOT1 (N2385, N2379);
or OR4 (N2386, N2385, N491, N715, N761);
buf BUF1 (N2387, N2358);
xor XOR2 (N2388, N2387, N2099);
and AND3 (N2389, N2359, N1237, N1179);
not NOT1 (N2390, N2381);
xor XOR2 (N2391, N2386, N1057);
nor NOR3 (N2392, N2378, N1338, N1733);
and AND2 (N2393, N2377, N2246);
and AND3 (N2394, N2390, N1633, N1653);
nand NAND2 (N2395, N2393, N949);
not NOT1 (N2396, N2388);
not NOT1 (N2397, N2367);
buf BUF1 (N2398, N2389);
and AND4 (N2399, N2398, N1923, N697, N1707);
nand NAND2 (N2400, N2384, N567);
xor XOR2 (N2401, N2396, N1358);
xor XOR2 (N2402, N2401, N1968);
buf BUF1 (N2403, N2394);
nor NOR3 (N2404, N2380, N1037, N1563);
xor XOR2 (N2405, N2404, N97);
xor XOR2 (N2406, N2383, N79);
nand NAND2 (N2407, N2392, N889);
nor NOR2 (N2408, N2397, N1362);
nor NOR4 (N2409, N2395, N2353, N2330, N1947);
nor NOR3 (N2410, N2405, N1636, N1027);
buf BUF1 (N2411, N2391);
or OR3 (N2412, N2409, N2394, N947);
not NOT1 (N2413, N2402);
buf BUF1 (N2414, N2400);
buf BUF1 (N2415, N2410);
or OR4 (N2416, N2403, N1877, N1434, N964);
nor NOR4 (N2417, N2414, N1919, N2183, N147);
and AND4 (N2418, N2416, N1879, N1953, N917);
not NOT1 (N2419, N2417);
nand NAND3 (N2420, N2418, N276, N938);
nand NAND2 (N2421, N2411, N1745);
nor NOR2 (N2422, N2420, N140);
nor NOR3 (N2423, N2413, N1228, N1187);
not NOT1 (N2424, N2419);
not NOT1 (N2425, N2423);
or OR3 (N2426, N2399, N1925, N873);
nand NAND2 (N2427, N2407, N1163);
or OR2 (N2428, N2408, N177);
or OR3 (N2429, N2424, N2268, N2400);
and AND2 (N2430, N2428, N645);
buf BUF1 (N2431, N2412);
or OR4 (N2432, N2425, N2164, N2016, N1558);
buf BUF1 (N2433, N2426);
xor XOR2 (N2434, N2431, N503);
and AND3 (N2435, N2406, N416, N1630);
buf BUF1 (N2436, N2429);
xor XOR2 (N2437, N2434, N406);
xor XOR2 (N2438, N2435, N828);
and AND3 (N2439, N2438, N1495, N1521);
buf BUF1 (N2440, N2439);
nand NAND2 (N2441, N2437, N361);
nand NAND3 (N2442, N2430, N2026, N2061);
buf BUF1 (N2443, N2422);
and AND4 (N2444, N2427, N1573, N2415, N1122);
xor XOR2 (N2445, N487, N169);
nor NOR4 (N2446, N2443, N578, N1796, N1121);
nand NAND2 (N2447, N2445, N877);
and AND4 (N2448, N2447, N1905, N2080, N1584);
or OR2 (N2449, N2432, N172);
buf BUF1 (N2450, N2449);
nand NAND2 (N2451, N2433, N866);
buf BUF1 (N2452, N2436);
not NOT1 (N2453, N2451);
xor XOR2 (N2454, N2450, N1686);
and AND2 (N2455, N2448, N731);
not NOT1 (N2456, N2452);
not NOT1 (N2457, N2454);
nand NAND3 (N2458, N2457, N756, N1516);
nor NOR4 (N2459, N2440, N2028, N681, N1301);
or OR3 (N2460, N2455, N723, N279);
or OR2 (N2461, N2421, N1969);
nand NAND2 (N2462, N2461, N1949);
buf BUF1 (N2463, N2446);
or OR3 (N2464, N2444, N2037, N1107);
xor XOR2 (N2465, N2458, N2143);
buf BUF1 (N2466, N2463);
or OR4 (N2467, N2453, N733, N1977, N1292);
and AND4 (N2468, N2441, N717, N420, N731);
buf BUF1 (N2469, N2467);
or OR2 (N2470, N2466, N99);
buf BUF1 (N2471, N2459);
nor NOR3 (N2472, N2470, N2142, N953);
or OR4 (N2473, N2465, N340, N2076, N939);
and AND2 (N2474, N2471, N2090);
xor XOR2 (N2475, N2460, N2124);
and AND3 (N2476, N2469, N145, N950);
not NOT1 (N2477, N2476);
nand NAND2 (N2478, N2472, N100);
and AND4 (N2479, N2473, N865, N517, N1217);
buf BUF1 (N2480, N2478);
and AND4 (N2481, N2462, N2334, N203, N1641);
xor XOR2 (N2482, N2456, N1183);
nor NOR2 (N2483, N2477, N25);
not NOT1 (N2484, N2464);
xor XOR2 (N2485, N2483, N496);
xor XOR2 (N2486, N2442, N2191);
buf BUF1 (N2487, N2468);
nand NAND3 (N2488, N2481, N2377, N666);
or OR4 (N2489, N2488, N1415, N536, N1309);
nor NOR4 (N2490, N2480, N2306, N1798, N281);
or OR2 (N2491, N2475, N1455);
nand NAND3 (N2492, N2484, N1888, N1630);
nand NAND4 (N2493, N2492, N1277, N251, N1672);
nand NAND4 (N2494, N2479, N43, N1740, N2256);
xor XOR2 (N2495, N2487, N995);
xor XOR2 (N2496, N2495, N1540);
xor XOR2 (N2497, N2491, N1917);
or OR4 (N2498, N2486, N1025, N164, N2181);
buf BUF1 (N2499, N2485);
or OR3 (N2500, N2499, N1165, N566);
and AND2 (N2501, N2474, N48);
nand NAND3 (N2502, N2497, N2172, N1288);
nand NAND2 (N2503, N2494, N2239);
buf BUF1 (N2504, N2490);
nor NOR4 (N2505, N2503, N1900, N1289, N1346);
nand NAND2 (N2506, N2505, N88);
buf BUF1 (N2507, N2502);
or OR3 (N2508, N2506, N2301, N2220);
or OR2 (N2509, N2501, N1729);
not NOT1 (N2510, N2500);
and AND4 (N2511, N2504, N220, N444, N2005);
xor XOR2 (N2512, N2509, N1975);
buf BUF1 (N2513, N2507);
and AND3 (N2514, N2511, N1767, N1657);
not NOT1 (N2515, N2510);
not NOT1 (N2516, N2489);
buf BUF1 (N2517, N2514);
nand NAND3 (N2518, N2496, N430, N718);
xor XOR2 (N2519, N2517, N241);
and AND3 (N2520, N2508, N2183, N1618);
not NOT1 (N2521, N2498);
xor XOR2 (N2522, N2518, N2466);
or OR4 (N2523, N2515, N2390, N2076, N278);
nand NAND3 (N2524, N2520, N1541, N2357);
not NOT1 (N2525, N2516);
not NOT1 (N2526, N2519);
buf BUF1 (N2527, N2525);
not NOT1 (N2528, N2523);
and AND4 (N2529, N2524, N2054, N267, N542);
not NOT1 (N2530, N2482);
and AND4 (N2531, N2528, N410, N271, N126);
xor XOR2 (N2532, N2521, N54);
and AND3 (N2533, N2529, N1852, N2246);
not NOT1 (N2534, N2522);
xor XOR2 (N2535, N2533, N1795);
xor XOR2 (N2536, N2530, N533);
xor XOR2 (N2537, N2527, N609);
and AND3 (N2538, N2535, N1598, N830);
nand NAND3 (N2539, N2493, N1753, N608);
and AND2 (N2540, N2531, N587);
xor XOR2 (N2541, N2512, N1405);
or OR4 (N2542, N2538, N1932, N2205, N2498);
and AND4 (N2543, N2526, N1048, N2301, N219);
and AND4 (N2544, N2513, N1554, N1435, N699);
or OR3 (N2545, N2539, N1623, N2524);
nor NOR3 (N2546, N2532, N754, N2416);
and AND4 (N2547, N2545, N1802, N642, N1783);
or OR4 (N2548, N2541, N24, N2474, N298);
xor XOR2 (N2549, N2534, N2073);
nand NAND4 (N2550, N2547, N1270, N1567, N2536);
nor NOR2 (N2551, N704, N1116);
and AND4 (N2552, N2540, N2402, N2465, N635);
nand NAND2 (N2553, N2546, N418);
not NOT1 (N2554, N2537);
and AND4 (N2555, N2553, N894, N639, N183);
nor NOR2 (N2556, N2551, N2444);
and AND4 (N2557, N2543, N2503, N548, N463);
nand NAND3 (N2558, N2557, N2324, N2498);
nor NOR3 (N2559, N2544, N2527, N2155);
not NOT1 (N2560, N2550);
or OR4 (N2561, N2559, N2453, N690, N1841);
not NOT1 (N2562, N2560);
nand NAND2 (N2563, N2555, N1566);
or OR4 (N2564, N2563, N1794, N621, N1911);
or OR4 (N2565, N2558, N1397, N1061, N436);
not NOT1 (N2566, N2552);
nor NOR4 (N2567, N2564, N778, N1453, N2196);
xor XOR2 (N2568, N2554, N2011);
or OR3 (N2569, N2565, N2324, N453);
not NOT1 (N2570, N2549);
nand NAND4 (N2571, N2568, N2426, N2530, N1786);
buf BUF1 (N2572, N2571);
xor XOR2 (N2573, N2572, N903);
or OR4 (N2574, N2548, N2170, N1037, N449);
or OR4 (N2575, N2556, N833, N762, N2007);
and AND2 (N2576, N2569, N1226);
or OR4 (N2577, N2575, N1827, N892, N709);
or OR3 (N2578, N2577, N844, N1731);
and AND3 (N2579, N2573, N423, N2390);
or OR3 (N2580, N2567, N1571, N1003);
and AND3 (N2581, N2570, N2423, N2372);
xor XOR2 (N2582, N2581, N1654);
nand NAND2 (N2583, N2574, N768);
nor NOR3 (N2584, N2542, N586, N1201);
or OR4 (N2585, N2561, N508, N1369, N1255);
xor XOR2 (N2586, N2580, N819);
nand NAND2 (N2587, N2583, N1857);
not NOT1 (N2588, N2566);
not NOT1 (N2589, N2585);
or OR2 (N2590, N2578, N2009);
not NOT1 (N2591, N2584);
or OR3 (N2592, N2562, N1474, N1735);
nand NAND2 (N2593, N2591, N320);
nand NAND4 (N2594, N2587, N957, N2531, N155);
and AND3 (N2595, N2586, N2397, N126);
nor NOR4 (N2596, N2576, N2038, N182, N939);
buf BUF1 (N2597, N2589);
nand NAND3 (N2598, N2597, N2081, N1416);
nand NAND2 (N2599, N2595, N1500);
xor XOR2 (N2600, N2596, N432);
not NOT1 (N2601, N2592);
nor NOR2 (N2602, N2590, N2505);
not NOT1 (N2603, N2582);
buf BUF1 (N2604, N2602);
or OR3 (N2605, N2598, N1618, N895);
not NOT1 (N2606, N2603);
or OR2 (N2607, N2593, N1064);
and AND2 (N2608, N2604, N1170);
nor NOR4 (N2609, N2594, N178, N1910, N1793);
buf BUF1 (N2610, N2606);
nand NAND4 (N2611, N2601, N638, N531, N1439);
or OR2 (N2612, N2610, N2466);
nor NOR3 (N2613, N2579, N1385, N1719);
not NOT1 (N2614, N2605);
nor NOR3 (N2615, N2614, N1709, N1608);
nand NAND4 (N2616, N2612, N2276, N1614, N2557);
buf BUF1 (N2617, N2613);
nand NAND2 (N2618, N2611, N461);
and AND3 (N2619, N2607, N1645, N401);
buf BUF1 (N2620, N2609);
or OR4 (N2621, N2588, N648, N2053, N445);
and AND3 (N2622, N2615, N1513, N1140);
xor XOR2 (N2623, N2617, N185);
and AND4 (N2624, N2618, N874, N1994, N1987);
or OR3 (N2625, N2624, N429, N2413);
xor XOR2 (N2626, N2616, N643);
nor NOR2 (N2627, N2625, N1984);
nand NAND4 (N2628, N2623, N1330, N1662, N1201);
not NOT1 (N2629, N2621);
and AND4 (N2630, N2622, N1534, N429, N1693);
xor XOR2 (N2631, N2620, N435);
nand NAND4 (N2632, N2626, N184, N148, N1657);
or OR3 (N2633, N2628, N264, N322);
nand NAND4 (N2634, N2631, N759, N2158, N1173);
nand NAND2 (N2635, N2599, N2479);
nor NOR4 (N2636, N2630, N988, N186, N780);
xor XOR2 (N2637, N2632, N2603);
not NOT1 (N2638, N2635);
or OR2 (N2639, N2627, N2041);
nand NAND3 (N2640, N2638, N1161, N881);
nor NOR3 (N2641, N2640, N1250, N1741);
not NOT1 (N2642, N2629);
nand NAND3 (N2643, N2637, N616, N2101);
nand NAND2 (N2644, N2642, N684);
not NOT1 (N2645, N2643);
nand NAND3 (N2646, N2645, N2014, N1964);
or OR3 (N2647, N2608, N1068, N2444);
or OR4 (N2648, N2644, N1732, N362, N480);
nor NOR4 (N2649, N2639, N1218, N2066, N1915);
or OR3 (N2650, N2646, N56, N1899);
xor XOR2 (N2651, N2641, N501);
nor NOR4 (N2652, N2649, N2569, N2463, N329);
nand NAND3 (N2653, N2634, N980, N459);
not NOT1 (N2654, N2652);
nor NOR3 (N2655, N2653, N1999, N364);
buf BUF1 (N2656, N2647);
buf BUF1 (N2657, N2633);
not NOT1 (N2658, N2650);
xor XOR2 (N2659, N2619, N1056);
xor XOR2 (N2660, N2656, N2475);
nor NOR4 (N2661, N2654, N411, N358, N314);
xor XOR2 (N2662, N2658, N189);
nor NOR2 (N2663, N2651, N914);
buf BUF1 (N2664, N2660);
not NOT1 (N2665, N2659);
xor XOR2 (N2666, N2600, N759);
nor NOR3 (N2667, N2666, N1963, N1368);
or OR3 (N2668, N2667, N223, N1601);
buf BUF1 (N2669, N2662);
nand NAND2 (N2670, N2655, N2511);
and AND2 (N2671, N2636, N2394);
and AND4 (N2672, N2665, N575, N357, N2370);
not NOT1 (N2673, N2672);
buf BUF1 (N2674, N2670);
xor XOR2 (N2675, N2669, N396);
not NOT1 (N2676, N2673);
or OR3 (N2677, N2676, N438, N666);
nand NAND3 (N2678, N2677, N734, N1933);
and AND2 (N2679, N2657, N446);
nor NOR4 (N2680, N2664, N47, N1169, N2247);
and AND3 (N2681, N2648, N1065, N2056);
or OR2 (N2682, N2674, N2045);
not NOT1 (N2683, N2682);
not NOT1 (N2684, N2680);
or OR4 (N2685, N2679, N1423, N109, N860);
and AND2 (N2686, N2684, N2262);
nand NAND3 (N2687, N2675, N2158, N1564);
and AND4 (N2688, N2678, N426, N2385, N786);
nand NAND4 (N2689, N2663, N1466, N591, N220);
xor XOR2 (N2690, N2661, N584);
buf BUF1 (N2691, N2688);
nand NAND3 (N2692, N2685, N2528, N584);
nor NOR4 (N2693, N2683, N2285, N593, N777);
xor XOR2 (N2694, N2687, N1537);
or OR4 (N2695, N2692, N1620, N345, N118);
or OR3 (N2696, N2693, N1927, N588);
and AND2 (N2697, N2689, N1000);
xor XOR2 (N2698, N2696, N1469);
nand NAND3 (N2699, N2690, N560, N1223);
xor XOR2 (N2700, N2695, N77);
and AND3 (N2701, N2694, N1852, N507);
xor XOR2 (N2702, N2699, N2566);
not NOT1 (N2703, N2671);
nand NAND2 (N2704, N2686, N1841);
not NOT1 (N2705, N2681);
nand NAND4 (N2706, N2698, N2417, N2051, N1780);
xor XOR2 (N2707, N2697, N2421);
xor XOR2 (N2708, N2702, N218);
nor NOR2 (N2709, N2703, N620);
or OR3 (N2710, N2701, N1306, N799);
and AND3 (N2711, N2691, N1481, N1457);
buf BUF1 (N2712, N2708);
nor NOR3 (N2713, N2705, N1098, N1400);
nor NOR4 (N2714, N2710, N953, N2679, N1245);
buf BUF1 (N2715, N2714);
nor NOR3 (N2716, N2706, N1394, N1389);
buf BUF1 (N2717, N2715);
nor NOR3 (N2718, N2713, N1625, N1880);
buf BUF1 (N2719, N2709);
nand NAND2 (N2720, N2700, N454);
nand NAND4 (N2721, N2704, N1021, N891, N615);
or OR4 (N2722, N2718, N1007, N2463, N2440);
and AND3 (N2723, N2711, N2308, N1255);
buf BUF1 (N2724, N2719);
not NOT1 (N2725, N2668);
nand NAND3 (N2726, N2721, N63, N291);
buf BUF1 (N2727, N2724);
not NOT1 (N2728, N2707);
buf BUF1 (N2729, N2723);
nor NOR3 (N2730, N2729, N1563, N2535);
nor NOR2 (N2731, N2716, N523);
xor XOR2 (N2732, N2722, N909);
or OR3 (N2733, N2731, N354, N2036);
xor XOR2 (N2734, N2728, N438);
nand NAND2 (N2735, N2725, N2332);
or OR2 (N2736, N2717, N1983);
not NOT1 (N2737, N2712);
buf BUF1 (N2738, N2737);
nand NAND2 (N2739, N2736, N1362);
not NOT1 (N2740, N2739);
and AND3 (N2741, N2733, N994, N2264);
not NOT1 (N2742, N2732);
or OR3 (N2743, N2730, N482, N2082);
buf BUF1 (N2744, N2727);
not NOT1 (N2745, N2734);
and AND3 (N2746, N2726, N2421, N2233);
nand NAND3 (N2747, N2740, N2585, N1399);
nor NOR4 (N2748, N2746, N857, N1244, N2254);
not NOT1 (N2749, N2748);
nor NOR4 (N2750, N2735, N1389, N938, N931);
or OR4 (N2751, N2744, N1209, N841, N1766);
nor NOR3 (N2752, N2749, N1869, N1515);
nand NAND3 (N2753, N2741, N1839, N12);
not NOT1 (N2754, N2743);
and AND4 (N2755, N2751, N329, N1281, N2527);
or OR4 (N2756, N2720, N1727, N817, N2405);
not NOT1 (N2757, N2756);
xor XOR2 (N2758, N2738, N1280);
buf BUF1 (N2759, N2752);
nor NOR3 (N2760, N2754, N837, N1189);
and AND4 (N2761, N2750, N1895, N413, N594);
xor XOR2 (N2762, N2745, N1580);
xor XOR2 (N2763, N2762, N17);
and AND3 (N2764, N2753, N557, N1931);
or OR4 (N2765, N2760, N1165, N710, N1294);
buf BUF1 (N2766, N2747);
nand NAND2 (N2767, N2765, N808);
nor NOR2 (N2768, N2742, N2368);
nand NAND3 (N2769, N2768, N285, N1604);
nor NOR3 (N2770, N2763, N1741, N2005);
nand NAND3 (N2771, N2770, N447, N1432);
nor NOR4 (N2772, N2771, N1550, N228, N1550);
or OR3 (N2773, N2758, N2381, N244);
buf BUF1 (N2774, N2772);
not NOT1 (N2775, N2759);
buf BUF1 (N2776, N2774);
xor XOR2 (N2777, N2766, N2474);
buf BUF1 (N2778, N2755);
nor NOR3 (N2779, N2776, N996, N2101);
and AND2 (N2780, N2764, N276);
nand NAND2 (N2781, N2779, N905);
nor NOR3 (N2782, N2769, N1575, N300);
xor XOR2 (N2783, N2781, N2025);
xor XOR2 (N2784, N2773, N1397);
xor XOR2 (N2785, N2777, N1211);
buf BUF1 (N2786, N2785);
nand NAND3 (N2787, N2761, N1846, N1657);
not NOT1 (N2788, N2786);
and AND3 (N2789, N2788, N1792, N2321);
and AND2 (N2790, N2780, N1556);
not NOT1 (N2791, N2790);
or OR2 (N2792, N2757, N2077);
nor NOR2 (N2793, N2787, N1179);
and AND3 (N2794, N2782, N1482, N1642);
xor XOR2 (N2795, N2783, N1834);
nand NAND2 (N2796, N2767, N701);
nand NAND4 (N2797, N2793, N1639, N260, N649);
nor NOR3 (N2798, N2795, N2242, N96);
or OR3 (N2799, N2792, N2585, N527);
nand NAND3 (N2800, N2797, N1337, N1850);
nand NAND3 (N2801, N2784, N1367, N808);
and AND2 (N2802, N2775, N2287);
nand NAND2 (N2803, N2794, N2060);
nor NOR4 (N2804, N2789, N2314, N21, N418);
not NOT1 (N2805, N2800);
nor NOR4 (N2806, N2802, N2484, N828, N1751);
nor NOR2 (N2807, N2803, N964);
buf BUF1 (N2808, N2791);
buf BUF1 (N2809, N2799);
nand NAND4 (N2810, N2798, N633, N120, N787);
or OR2 (N2811, N2804, N2568);
or OR3 (N2812, N2805, N2201, N2605);
and AND3 (N2813, N2801, N503, N2128);
nor NOR3 (N2814, N2806, N1332, N2735);
xor XOR2 (N2815, N2778, N2021);
or OR3 (N2816, N2815, N2094, N1929);
and AND2 (N2817, N2816, N1913);
nand NAND3 (N2818, N2811, N866, N2272);
not NOT1 (N2819, N2796);
and AND2 (N2820, N2817, N242);
xor XOR2 (N2821, N2810, N1184);
nand NAND2 (N2822, N2813, N1439);
nand NAND4 (N2823, N2812, N34, N1527, N1048);
nor NOR3 (N2824, N2818, N1623, N2610);
nand NAND2 (N2825, N2823, N347);
nand NAND2 (N2826, N2814, N800);
not NOT1 (N2827, N2820);
buf BUF1 (N2828, N2809);
xor XOR2 (N2829, N2827, N1231);
nor NOR4 (N2830, N2829, N1725, N428, N1223);
nand NAND2 (N2831, N2808, N2405);
not NOT1 (N2832, N2828);
buf BUF1 (N2833, N2819);
not NOT1 (N2834, N2825);
buf BUF1 (N2835, N2832);
and AND4 (N2836, N2831, N1443, N1804, N524);
or OR4 (N2837, N2830, N2342, N1803, N2564);
or OR2 (N2838, N2833, N722);
and AND4 (N2839, N2821, N1369, N659, N599);
or OR2 (N2840, N2837, N1223);
buf BUF1 (N2841, N2839);
not NOT1 (N2842, N2840);
nand NAND3 (N2843, N2834, N203, N493);
nor NOR3 (N2844, N2843, N713, N2105);
not NOT1 (N2845, N2841);
and AND2 (N2846, N2844, N329);
or OR3 (N2847, N2846, N849, N1483);
not NOT1 (N2848, N2845);
nor NOR4 (N2849, N2835, N1527, N1407, N1696);
xor XOR2 (N2850, N2847, N2469);
buf BUF1 (N2851, N2836);
xor XOR2 (N2852, N2851, N152);
and AND2 (N2853, N2822, N1128);
and AND3 (N2854, N2826, N753, N2732);
and AND2 (N2855, N2854, N1047);
buf BUF1 (N2856, N2824);
xor XOR2 (N2857, N2842, N496);
nand NAND2 (N2858, N2857, N1008);
and AND3 (N2859, N2853, N993, N2154);
nor NOR4 (N2860, N2850, N712, N1705, N2588);
and AND4 (N2861, N2848, N1692, N2816, N1280);
not NOT1 (N2862, N2855);
nand NAND2 (N2863, N2838, N1750);
nor NOR2 (N2864, N2861, N112);
and AND4 (N2865, N2849, N555, N921, N2165);
or OR4 (N2866, N2865, N194, N1831, N1201);
buf BUF1 (N2867, N2866);
not NOT1 (N2868, N2859);
and AND4 (N2869, N2852, N127, N2090, N401);
or OR2 (N2870, N2862, N2317);
buf BUF1 (N2871, N2860);
nand NAND3 (N2872, N2858, N2642, N2718);
nand NAND4 (N2873, N2863, N2232, N388, N100);
not NOT1 (N2874, N2871);
nand NAND4 (N2875, N2864, N1596, N1582, N1577);
or OR3 (N2876, N2867, N1077, N582);
nand NAND2 (N2877, N2868, N583);
nand NAND4 (N2878, N2875, N74, N359, N721);
nor NOR3 (N2879, N2874, N2853, N157);
not NOT1 (N2880, N2872);
buf BUF1 (N2881, N2879);
nor NOR3 (N2882, N2869, N695, N2560);
buf BUF1 (N2883, N2876);
or OR3 (N2884, N2856, N869, N2517);
nand NAND3 (N2885, N2881, N776, N609);
nand NAND2 (N2886, N2880, N2493);
not NOT1 (N2887, N2885);
and AND4 (N2888, N2884, N1962, N38, N2790);
not NOT1 (N2889, N2877);
or OR3 (N2890, N2807, N194, N2690);
xor XOR2 (N2891, N2882, N339);
xor XOR2 (N2892, N2873, N954);
nor NOR2 (N2893, N2883, N762);
xor XOR2 (N2894, N2870, N1891);
nand NAND2 (N2895, N2893, N1123);
xor XOR2 (N2896, N2887, N2338);
buf BUF1 (N2897, N2892);
nand NAND3 (N2898, N2886, N526, N225);
not NOT1 (N2899, N2897);
buf BUF1 (N2900, N2896);
nor NOR3 (N2901, N2891, N876, N1);
buf BUF1 (N2902, N2878);
and AND2 (N2903, N2898, N547);
nand NAND3 (N2904, N2901, N1602, N2299);
nor NOR2 (N2905, N2904, N691);
nor NOR4 (N2906, N2903, N1131, N1361, N1312);
buf BUF1 (N2907, N2894);
or OR2 (N2908, N2906, N673);
nand NAND2 (N2909, N2899, N2838);
and AND4 (N2910, N2889, N2225, N2807, N806);
nor NOR4 (N2911, N2890, N120, N2227, N2566);
nor NOR3 (N2912, N2902, N891, N960);
nand NAND3 (N2913, N2910, N2701, N2815);
buf BUF1 (N2914, N2908);
buf BUF1 (N2915, N2907);
and AND4 (N2916, N2915, N1766, N850, N1383);
xor XOR2 (N2917, N2911, N822);
or OR4 (N2918, N2888, N242, N777, N1856);
or OR3 (N2919, N2895, N2106, N1365);
or OR4 (N2920, N2913, N2332, N624, N1159);
nor NOR3 (N2921, N2914, N1523, N2126);
buf BUF1 (N2922, N2917);
and AND3 (N2923, N2909, N2607, N704);
or OR3 (N2924, N2919, N804, N438);
nor NOR2 (N2925, N2916, N2711);
not NOT1 (N2926, N2925);
and AND3 (N2927, N2918, N1345, N414);
and AND2 (N2928, N2924, N981);
nand NAND3 (N2929, N2920, N1426, N2051);
xor XOR2 (N2930, N2926, N2260);
buf BUF1 (N2931, N2928);
nand NAND3 (N2932, N2912, N2040, N505);
or OR2 (N2933, N2922, N1061);
nor NOR4 (N2934, N2933, N544, N269, N2637);
and AND2 (N2935, N2921, N1243);
nand NAND3 (N2936, N2935, N2340, N2296);
and AND2 (N2937, N2936, N2898);
not NOT1 (N2938, N2937);
not NOT1 (N2939, N2900);
and AND4 (N2940, N2938, N341, N1916, N1506);
nor NOR4 (N2941, N2927, N224, N1326, N2236);
nand NAND4 (N2942, N2932, N277, N507, N145);
nor NOR3 (N2943, N2929, N935, N2604);
and AND4 (N2944, N2941, N718, N1179, N2530);
xor XOR2 (N2945, N2940, N1824);
not NOT1 (N2946, N2944);
and AND4 (N2947, N2923, N2284, N918, N11);
or OR3 (N2948, N2931, N88, N523);
and AND3 (N2949, N2930, N1237, N2899);
nand NAND3 (N2950, N2947, N268, N2310);
or OR3 (N2951, N2934, N1994, N1065);
or OR4 (N2952, N2943, N2572, N396, N602);
or OR2 (N2953, N2946, N1219);
not NOT1 (N2954, N2950);
nand NAND4 (N2955, N2953, N1278, N2158, N434);
or OR4 (N2956, N2951, N358, N912, N1360);
buf BUF1 (N2957, N2948);
and AND4 (N2958, N2942, N1310, N95, N2032);
or OR3 (N2959, N2954, N762, N2766);
and AND4 (N2960, N2952, N882, N709, N2880);
nor NOR4 (N2961, N2945, N799, N2689, N2960);
nor NOR4 (N2962, N1411, N199, N1220, N1503);
not NOT1 (N2963, N2958);
or OR3 (N2964, N2905, N2426, N1276);
nor NOR3 (N2965, N2963, N638, N2708);
not NOT1 (N2966, N2957);
or OR3 (N2967, N2956, N945, N383);
and AND2 (N2968, N2961, N2856);
buf BUF1 (N2969, N2966);
not NOT1 (N2970, N2964);
and AND4 (N2971, N2970, N660, N2789, N2883);
nor NOR2 (N2972, N2969, N787);
xor XOR2 (N2973, N2968, N399);
xor XOR2 (N2974, N2972, N1579);
nand NAND4 (N2975, N2955, N1493, N505, N2449);
buf BUF1 (N2976, N2965);
or OR3 (N2977, N2949, N2611, N91);
and AND2 (N2978, N2976, N1760);
xor XOR2 (N2979, N2959, N2440);
and AND3 (N2980, N2967, N216, N888);
nand NAND4 (N2981, N2973, N2212, N1284, N133);
buf BUF1 (N2982, N2981);
or OR2 (N2983, N2978, N101);
xor XOR2 (N2984, N2975, N2852);
nand NAND4 (N2985, N2939, N2235, N1063, N2477);
or OR4 (N2986, N2979, N2736, N399, N1158);
xor XOR2 (N2987, N2985, N2429);
nand NAND2 (N2988, N2982, N1784);
not NOT1 (N2989, N2962);
xor XOR2 (N2990, N2989, N1994);
nand NAND2 (N2991, N2977, N1179);
buf BUF1 (N2992, N2983);
not NOT1 (N2993, N2988);
and AND3 (N2994, N2980, N1696, N152);
nor NOR2 (N2995, N2974, N876);
not NOT1 (N2996, N2971);
xor XOR2 (N2997, N2992, N2399);
or OR3 (N2998, N2995, N1842, N2932);
nor NOR4 (N2999, N2994, N2532, N922, N1221);
and AND3 (N3000, N2997, N2579, N2064);
nor NOR4 (N3001, N2993, N1508, N1713, N1822);
buf BUF1 (N3002, N3001);
and AND4 (N3003, N2984, N2802, N1268, N1426);
nor NOR2 (N3004, N3002, N1967);
and AND4 (N3005, N2991, N622, N912, N1231);
xor XOR2 (N3006, N2987, N1795);
or OR3 (N3007, N2986, N2370, N2466);
not NOT1 (N3008, N3005);
xor XOR2 (N3009, N3007, N1211);
buf BUF1 (N3010, N3008);
and AND3 (N3011, N3004, N1920, N1601);
not NOT1 (N3012, N2996);
and AND3 (N3013, N3000, N2291, N908);
and AND2 (N3014, N3009, N2627);
not NOT1 (N3015, N3011);
buf BUF1 (N3016, N2998);
not NOT1 (N3017, N3015);
or OR4 (N3018, N3016, N3014, N2595, N2285);
nor NOR4 (N3019, N2224, N2682, N2877, N1835);
or OR3 (N3020, N2999, N2501, N1810);
or OR2 (N3021, N2990, N1342);
and AND4 (N3022, N3006, N782, N2100, N1176);
buf BUF1 (N3023, N3018);
and AND2 (N3024, N3021, N1982);
or OR2 (N3025, N3010, N1650);
not NOT1 (N3026, N3003);
nand NAND4 (N3027, N3026, N993, N1835, N2264);
nor NOR4 (N3028, N3023, N2314, N410, N547);
or OR2 (N3029, N3013, N2289);
buf BUF1 (N3030, N3025);
xor XOR2 (N3031, N3028, N360);
nand NAND2 (N3032, N3030, N2983);
nor NOR4 (N3033, N3012, N2887, N778, N2117);
not NOT1 (N3034, N3024);
xor XOR2 (N3035, N3027, N2900);
nand NAND3 (N3036, N3017, N2323, N1430);
or OR2 (N3037, N3022, N2378);
or OR4 (N3038, N3029, N2277, N815, N2681);
not NOT1 (N3039, N3038);
and AND4 (N3040, N3036, N1889, N2397, N263);
not NOT1 (N3041, N3032);
not NOT1 (N3042, N3040);
or OR3 (N3043, N3037, N1748, N318);
nor NOR2 (N3044, N3043, N1077);
buf BUF1 (N3045, N3034);
xor XOR2 (N3046, N3033, N491);
nand NAND3 (N3047, N3019, N2055, N376);
nand NAND4 (N3048, N3045, N1140, N1239, N2571);
and AND3 (N3049, N3035, N530, N1317);
nor NOR2 (N3050, N3044, N494);
not NOT1 (N3051, N3042);
nand NAND3 (N3052, N3049, N2917, N3);
and AND4 (N3053, N3051, N706, N1901, N2933);
xor XOR2 (N3054, N3020, N1319);
and AND3 (N3055, N3039, N2473, N1498);
nor NOR2 (N3056, N3047, N1728);
nand NAND2 (N3057, N3050, N2858);
xor XOR2 (N3058, N3041, N528);
xor XOR2 (N3059, N3055, N2176);
nor NOR3 (N3060, N3057, N1842, N923);
and AND4 (N3061, N3054, N2352, N2351, N1256);
or OR3 (N3062, N3060, N1681, N276);
buf BUF1 (N3063, N3052);
nor NOR2 (N3064, N3058, N629);
xor XOR2 (N3065, N3064, N2935);
buf BUF1 (N3066, N3065);
not NOT1 (N3067, N3061);
nor NOR4 (N3068, N3046, N1264, N2514, N1966);
buf BUF1 (N3069, N3059);
nor NOR3 (N3070, N3031, N2694, N1087);
xor XOR2 (N3071, N3069, N2723);
nand NAND4 (N3072, N3048, N886, N2995, N2299);
buf BUF1 (N3073, N3066);
xor XOR2 (N3074, N3070, N91);
xor XOR2 (N3075, N3073, N793);
nor NOR2 (N3076, N3068, N2029);
or OR3 (N3077, N3075, N361, N601);
nand NAND2 (N3078, N3072, N2290);
not NOT1 (N3079, N3067);
and AND2 (N3080, N3076, N196);
or OR4 (N3081, N3062, N667, N497, N824);
or OR3 (N3082, N3074, N2477, N1102);
or OR2 (N3083, N3081, N728);
nand NAND2 (N3084, N3080, N2725);
not NOT1 (N3085, N3078);
and AND3 (N3086, N3083, N437, N1483);
not NOT1 (N3087, N3086);
xor XOR2 (N3088, N3077, N282);
nand NAND2 (N3089, N3079, N2138);
nor NOR4 (N3090, N3087, N694, N942, N2494);
nor NOR4 (N3091, N3082, N2900, N1632, N2284);
nand NAND2 (N3092, N3090, N1360);
xor XOR2 (N3093, N3071, N975);
nand NAND4 (N3094, N3092, N497, N1045, N1621);
and AND4 (N3095, N3093, N218, N941, N2540);
or OR4 (N3096, N3094, N1350, N1088, N2659);
xor XOR2 (N3097, N3088, N2037);
and AND4 (N3098, N3091, N713, N182, N1197);
xor XOR2 (N3099, N3056, N1962);
or OR4 (N3100, N3053, N2363, N2153, N1005);
and AND3 (N3101, N3098, N2098, N645);
or OR4 (N3102, N3101, N1679, N2677, N27);
not NOT1 (N3103, N3097);
xor XOR2 (N3104, N3102, N732);
nor NOR4 (N3105, N3095, N2761, N1945, N2953);
buf BUF1 (N3106, N3105);
or OR4 (N3107, N3099, N426, N1835, N2913);
nor NOR4 (N3108, N3085, N2239, N2550, N2258);
xor XOR2 (N3109, N3100, N1291);
xor XOR2 (N3110, N3103, N2058);
nor NOR3 (N3111, N3110, N1515, N2190);
nand NAND2 (N3112, N3096, N852);
xor XOR2 (N3113, N3106, N2000);
xor XOR2 (N3114, N3089, N300);
and AND4 (N3115, N3113, N437, N2420, N2363);
xor XOR2 (N3116, N3104, N2165);
or OR3 (N3117, N3107, N3062, N1369);
xor XOR2 (N3118, N3115, N1677);
not NOT1 (N3119, N3116);
and AND4 (N3120, N3114, N1715, N996, N1963);
nand NAND3 (N3121, N3108, N968, N2937);
nand NAND2 (N3122, N3112, N1554);
nor NOR4 (N3123, N3109, N1721, N1377, N830);
xor XOR2 (N3124, N3120, N1035);
not NOT1 (N3125, N3118);
nor NOR3 (N3126, N3125, N1686, N1771);
nand NAND3 (N3127, N3122, N746, N1518);
not NOT1 (N3128, N3063);
nor NOR2 (N3129, N3127, N301);
not NOT1 (N3130, N3128);
nand NAND3 (N3131, N3084, N2933, N3122);
buf BUF1 (N3132, N3121);
not NOT1 (N3133, N3131);
not NOT1 (N3134, N3123);
nor NOR2 (N3135, N3129, N264);
and AND3 (N3136, N3124, N1336, N2406);
not NOT1 (N3137, N3117);
nor NOR4 (N3138, N3126, N1218, N1624, N1452);
and AND4 (N3139, N3130, N1154, N3023, N1058);
or OR4 (N3140, N3136, N2338, N2510, N1983);
and AND3 (N3141, N3140, N2589, N2303);
not NOT1 (N3142, N3132);
buf BUF1 (N3143, N3138);
xor XOR2 (N3144, N3111, N1092);
nand NAND2 (N3145, N3135, N2252);
and AND4 (N3146, N3134, N1494, N2556, N2268);
nand NAND3 (N3147, N3141, N1881, N83);
or OR3 (N3148, N3133, N2479, N1400);
nand NAND3 (N3149, N3139, N2740, N2498);
nand NAND4 (N3150, N3146, N1745, N625, N861);
buf BUF1 (N3151, N3145);
or OR2 (N3152, N3137, N608);
nor NOR4 (N3153, N3119, N2530, N3147, N691);
buf BUF1 (N3154, N523);
not NOT1 (N3155, N3152);
or OR2 (N3156, N3149, N1829);
xor XOR2 (N3157, N3156, N837);
buf BUF1 (N3158, N3154);
not NOT1 (N3159, N3153);
and AND4 (N3160, N3144, N2117, N2502, N1998);
and AND4 (N3161, N3157, N1965, N2220, N271);
xor XOR2 (N3162, N3159, N484);
not NOT1 (N3163, N3142);
and AND4 (N3164, N3161, N1326, N1963, N3094);
not NOT1 (N3165, N3160);
nand NAND2 (N3166, N3158, N723);
buf BUF1 (N3167, N3148);
and AND3 (N3168, N3162, N181, N633);
and AND4 (N3169, N3155, N1766, N2690, N276);
nand NAND4 (N3170, N3168, N2445, N2728, N2722);
or OR3 (N3171, N3169, N2193, N829);
buf BUF1 (N3172, N3171);
and AND3 (N3173, N3165, N1699, N535);
or OR2 (N3174, N3164, N1616);
buf BUF1 (N3175, N3150);
not NOT1 (N3176, N3151);
not NOT1 (N3177, N3174);
xor XOR2 (N3178, N3172, N3111);
or OR4 (N3179, N3176, N607, N3039, N126);
and AND4 (N3180, N3167, N1003, N2856, N583);
and AND2 (N3181, N3163, N3115);
buf BUF1 (N3182, N3181);
nand NAND4 (N3183, N3179, N3024, N2126, N2510);
xor XOR2 (N3184, N3178, N337);
xor XOR2 (N3185, N3183, N258);
nor NOR3 (N3186, N3173, N2711, N2822);
buf BUF1 (N3187, N3184);
buf BUF1 (N3188, N3180);
or OR3 (N3189, N3186, N135, N1239);
nand NAND3 (N3190, N3187, N2429, N3003);
buf BUF1 (N3191, N3143);
xor XOR2 (N3192, N3189, N2554);
nor NOR4 (N3193, N3170, N1711, N1981, N1087);
nand NAND4 (N3194, N3166, N488, N2940, N354);
xor XOR2 (N3195, N3182, N2217);
not NOT1 (N3196, N3194);
and AND4 (N3197, N3175, N1769, N2851, N137);
buf BUF1 (N3198, N3190);
or OR2 (N3199, N3195, N1619);
buf BUF1 (N3200, N3199);
buf BUF1 (N3201, N3192);
and AND4 (N3202, N3177, N2194, N1822, N549);
buf BUF1 (N3203, N3191);
buf BUF1 (N3204, N3201);
or OR3 (N3205, N3185, N2931, N2880);
not NOT1 (N3206, N3193);
buf BUF1 (N3207, N3196);
or OR3 (N3208, N3207, N3149, N256);
or OR3 (N3209, N3205, N1716, N273);
nor NOR4 (N3210, N3200, N676, N238, N2470);
and AND3 (N3211, N3208, N785, N1187);
nor NOR3 (N3212, N3209, N2750, N2849);
nand NAND4 (N3213, N3206, N1265, N2460, N2514);
buf BUF1 (N3214, N3203);
and AND4 (N3215, N3202, N2350, N2130, N867);
buf BUF1 (N3216, N3212);
and AND3 (N3217, N3215, N2637, N816);
not NOT1 (N3218, N3217);
xor XOR2 (N3219, N3218, N2321);
nand NAND4 (N3220, N3198, N738, N2174, N1359);
xor XOR2 (N3221, N3216, N1869);
nand NAND4 (N3222, N3204, N8, N348, N2176);
not NOT1 (N3223, N3221);
endmodule