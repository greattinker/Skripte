// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N518,N500,N517,N506,N521,N514,N520,N519,N492,N522;

or OR3 (N23, N21, N11, N14);
xor XOR2 (N24, N22, N16);
buf BUF1 (N25, N6);
nor NOR2 (N26, N13, N4);
buf BUF1 (N27, N20);
not NOT1 (N28, N23);
buf BUF1 (N29, N17);
buf BUF1 (N30, N15);
nor NOR4 (N31, N5, N24, N4, N21);
nor NOR3 (N32, N1, N10, N5);
nand NAND3 (N33, N31, N9, N18);
or OR4 (N34, N6, N16, N31, N30);
buf BUF1 (N35, N16);
and AND3 (N36, N23, N13, N8);
or OR3 (N37, N26, N16, N14);
nor NOR2 (N38, N37, N35);
and AND3 (N39, N9, N4, N13);
nor NOR4 (N40, N25, N25, N30, N10);
or OR2 (N41, N36, N27);
not NOT1 (N42, N27);
nor NOR4 (N43, N41, N37, N8, N22);
xor XOR2 (N44, N42, N27);
nand NAND4 (N45, N40, N33, N7, N36);
or OR2 (N46, N11, N15);
nor NOR3 (N47, N46, N33, N42);
or OR2 (N48, N45, N31);
nand NAND3 (N49, N28, N40, N13);
buf BUF1 (N50, N38);
or OR2 (N51, N32, N50);
xor XOR2 (N52, N2, N30);
or OR3 (N53, N49, N5, N43);
not NOT1 (N54, N27);
buf BUF1 (N55, N48);
not NOT1 (N56, N54);
or OR4 (N57, N53, N32, N4, N32);
nand NAND2 (N58, N47, N40);
buf BUF1 (N59, N58);
not NOT1 (N60, N59);
xor XOR2 (N61, N57, N50);
buf BUF1 (N62, N51);
buf BUF1 (N63, N44);
or OR3 (N64, N52, N32, N8);
xor XOR2 (N65, N29, N29);
and AND2 (N66, N62, N47);
nor NOR4 (N67, N60, N52, N11, N10);
buf BUF1 (N68, N65);
nor NOR4 (N69, N68, N5, N36, N67);
or OR2 (N70, N19, N43);
nor NOR3 (N71, N66, N48, N47);
nand NAND3 (N72, N61, N54, N69);
nand NAND4 (N73, N50, N59, N60, N2);
nand NAND4 (N74, N63, N25, N62, N29);
xor XOR2 (N75, N56, N44);
nor NOR2 (N76, N34, N40);
nand NAND4 (N77, N64, N30, N72, N75);
buf BUF1 (N78, N67);
xor XOR2 (N79, N10, N70);
and AND3 (N80, N30, N27, N2);
nand NAND2 (N81, N74, N26);
or OR4 (N82, N78, N2, N8, N33);
not NOT1 (N83, N73);
nand NAND2 (N84, N83, N65);
not NOT1 (N85, N84);
and AND2 (N86, N76, N64);
buf BUF1 (N87, N71);
or OR4 (N88, N55, N49, N68, N27);
nor NOR2 (N89, N77, N80);
buf BUF1 (N90, N15);
nand NAND2 (N91, N86, N35);
buf BUF1 (N92, N85);
buf BUF1 (N93, N90);
or OR4 (N94, N39, N66, N8, N69);
or OR3 (N95, N79, N41, N47);
nor NOR4 (N96, N93, N9, N56, N34);
nand NAND2 (N97, N82, N89);
buf BUF1 (N98, N5);
nor NOR4 (N99, N96, N6, N26, N48);
nand NAND3 (N100, N94, N54, N16);
or OR3 (N101, N88, N44, N50);
or OR3 (N102, N97, N36, N1);
and AND3 (N103, N99, N41, N16);
and AND4 (N104, N95, N33, N84, N79);
nand NAND2 (N105, N100, N19);
not NOT1 (N106, N98);
nand NAND2 (N107, N91, N62);
buf BUF1 (N108, N92);
nand NAND4 (N109, N103, N3, N33, N106);
or OR3 (N110, N2, N74, N10);
not NOT1 (N111, N102);
not NOT1 (N112, N110);
not NOT1 (N113, N87);
xor XOR2 (N114, N108, N70);
nand NAND4 (N115, N109, N3, N112, N45);
and AND4 (N116, N86, N31, N19, N11);
nor NOR4 (N117, N105, N76, N52, N85);
or OR2 (N118, N113, N26);
xor XOR2 (N119, N101, N102);
nor NOR4 (N120, N119, N110, N35, N28);
buf BUF1 (N121, N104);
buf BUF1 (N122, N111);
not NOT1 (N123, N121);
and AND3 (N124, N81, N73, N113);
or OR2 (N125, N120, N63);
buf BUF1 (N126, N124);
not NOT1 (N127, N116);
not NOT1 (N128, N126);
buf BUF1 (N129, N107);
not NOT1 (N130, N123);
nand NAND4 (N131, N114, N40, N68, N96);
xor XOR2 (N132, N127, N109);
and AND2 (N133, N128, N33);
nor NOR2 (N134, N130, N71);
nand NAND3 (N135, N125, N20, N106);
buf BUF1 (N136, N135);
or OR2 (N137, N129, N121);
and AND2 (N138, N117, N123);
nand NAND4 (N139, N137, N126, N56, N113);
nor NOR2 (N140, N122, N64);
and AND2 (N141, N132, N73);
or OR2 (N142, N141, N13);
not NOT1 (N143, N134);
xor XOR2 (N144, N139, N16);
nor NOR2 (N145, N118, N48);
nor NOR3 (N146, N142, N9, N13);
and AND2 (N147, N144, N138);
and AND2 (N148, N72, N91);
nand NAND2 (N149, N147, N6);
nand NAND2 (N150, N115, N68);
nor NOR3 (N151, N140, N52, N134);
nor NOR3 (N152, N131, N82, N46);
xor XOR2 (N153, N149, N55);
or OR3 (N154, N146, N151, N36);
nand NAND4 (N155, N45, N49, N7, N15);
or OR3 (N156, N143, N143, N45);
nor NOR4 (N157, N153, N28, N61, N126);
or OR3 (N158, N150, N73, N101);
nor NOR3 (N159, N155, N87, N91);
and AND2 (N160, N154, N72);
not NOT1 (N161, N148);
nand NAND4 (N162, N133, N28, N17, N86);
xor XOR2 (N163, N162, N148);
and AND3 (N164, N136, N92, N128);
xor XOR2 (N165, N152, N49);
not NOT1 (N166, N158);
xor XOR2 (N167, N145, N121);
nor NOR4 (N168, N160, N110, N59, N73);
nor NOR2 (N169, N159, N152);
xor XOR2 (N170, N166, N166);
nand NAND4 (N171, N163, N42, N66, N23);
and AND4 (N172, N171, N169, N35, N34);
nand NAND4 (N173, N52, N48, N150, N153);
and AND4 (N174, N156, N98, N51, N23);
buf BUF1 (N175, N167);
or OR4 (N176, N164, N138, N109, N150);
or OR2 (N177, N168, N163);
not NOT1 (N178, N174);
or OR3 (N179, N172, N172, N132);
nor NOR4 (N180, N170, N70, N10, N46);
nor NOR4 (N181, N180, N56, N164, N78);
nor NOR2 (N182, N157, N37);
xor XOR2 (N183, N165, N125);
nand NAND4 (N184, N176, N3, N160, N130);
or OR2 (N185, N182, N139);
buf BUF1 (N186, N184);
xor XOR2 (N187, N161, N169);
not NOT1 (N188, N178);
not NOT1 (N189, N177);
not NOT1 (N190, N185);
xor XOR2 (N191, N188, N58);
not NOT1 (N192, N186);
nand NAND4 (N193, N192, N73, N98, N158);
or OR2 (N194, N193, N54);
buf BUF1 (N195, N187);
xor XOR2 (N196, N194, N53);
not NOT1 (N197, N183);
nand NAND3 (N198, N181, N112, N87);
nand NAND2 (N199, N196, N48);
or OR2 (N200, N189, N176);
nor NOR4 (N201, N195, N189, N84, N12);
buf BUF1 (N202, N179);
nand NAND3 (N203, N190, N185, N67);
not NOT1 (N204, N200);
buf BUF1 (N205, N199);
not NOT1 (N206, N203);
nor NOR2 (N207, N204, N205);
or OR3 (N208, N83, N22, N43);
or OR2 (N209, N208, N83);
not NOT1 (N210, N197);
nor NOR2 (N211, N206, N102);
buf BUF1 (N212, N202);
or OR3 (N213, N173, N144, N201);
nor NOR2 (N214, N47, N150);
or OR2 (N215, N214, N44);
buf BUF1 (N216, N213);
buf BUF1 (N217, N207);
buf BUF1 (N218, N175);
nor NOR4 (N219, N198, N119, N134, N67);
xor XOR2 (N220, N209, N118);
buf BUF1 (N221, N210);
buf BUF1 (N222, N212);
nor NOR2 (N223, N215, N67);
and AND2 (N224, N219, N159);
or OR3 (N225, N211, N217, N156);
buf BUF1 (N226, N109);
not NOT1 (N227, N218);
buf BUF1 (N228, N221);
nor NOR2 (N229, N191, N191);
buf BUF1 (N230, N224);
not NOT1 (N231, N222);
nor NOR2 (N232, N231, N147);
not NOT1 (N233, N223);
or OR3 (N234, N225, N35, N98);
not NOT1 (N235, N216);
buf BUF1 (N236, N230);
not NOT1 (N237, N234);
not NOT1 (N238, N228);
and AND4 (N239, N229, N21, N58, N222);
not NOT1 (N240, N226);
not NOT1 (N241, N233);
buf BUF1 (N242, N241);
xor XOR2 (N243, N220, N150);
nor NOR4 (N244, N243, N120, N102, N195);
or OR2 (N245, N242, N59);
nand NAND2 (N246, N227, N239);
and AND3 (N247, N236, N117, N233);
or OR4 (N248, N142, N203, N82, N40);
xor XOR2 (N249, N240, N26);
nor NOR3 (N250, N247, N18, N125);
or OR4 (N251, N250, N235, N170, N82);
buf BUF1 (N252, N95);
buf BUF1 (N253, N249);
and AND4 (N254, N245, N129, N66, N169);
buf BUF1 (N255, N237);
not NOT1 (N256, N255);
xor XOR2 (N257, N238, N202);
and AND4 (N258, N254, N167, N29, N154);
xor XOR2 (N259, N258, N77);
buf BUF1 (N260, N256);
nand NAND4 (N261, N248, N88, N49, N42);
nand NAND3 (N262, N246, N69, N178);
or OR3 (N263, N232, N254, N108);
buf BUF1 (N264, N263);
xor XOR2 (N265, N252, N68);
and AND4 (N266, N265, N244, N45, N83);
not NOT1 (N267, N107);
nand NAND2 (N268, N266, N34);
xor XOR2 (N269, N264, N79);
xor XOR2 (N270, N257, N120);
or OR4 (N271, N269, N217, N193, N92);
xor XOR2 (N272, N260, N38);
and AND3 (N273, N267, N149, N67);
nand NAND3 (N274, N273, N151, N206);
or OR4 (N275, N271, N249, N226, N131);
buf BUF1 (N276, N270);
nor NOR3 (N277, N259, N8, N175);
buf BUF1 (N278, N272);
nor NOR3 (N279, N274, N225, N7);
nor NOR4 (N280, N268, N136, N108, N16);
nor NOR2 (N281, N262, N85);
nor NOR3 (N282, N278, N23, N265);
not NOT1 (N283, N261);
not NOT1 (N284, N281);
nand NAND3 (N285, N279, N64, N65);
and AND4 (N286, N253, N149, N115, N155);
nor NOR4 (N287, N282, N261, N72, N264);
and AND3 (N288, N286, N176, N116);
not NOT1 (N289, N251);
not NOT1 (N290, N285);
or OR3 (N291, N275, N174, N97);
not NOT1 (N292, N277);
or OR2 (N293, N290, N262);
nor NOR4 (N294, N283, N198, N245, N1);
nor NOR2 (N295, N280, N108);
xor XOR2 (N296, N276, N21);
nand NAND4 (N297, N294, N234, N117, N115);
nand NAND3 (N298, N293, N254, N217);
not NOT1 (N299, N296);
buf BUF1 (N300, N297);
or OR2 (N301, N299, N297);
xor XOR2 (N302, N291, N140);
xor XOR2 (N303, N288, N65);
or OR3 (N304, N287, N229, N227);
buf BUF1 (N305, N292);
nor NOR4 (N306, N300, N254, N136, N106);
and AND3 (N307, N301, N226, N143);
or OR3 (N308, N306, N202, N291);
nor NOR4 (N309, N302, N122, N261, N273);
nor NOR3 (N310, N303, N149, N8);
or OR3 (N311, N307, N163, N54);
buf BUF1 (N312, N309);
nor NOR3 (N313, N298, N263, N259);
not NOT1 (N314, N308);
and AND4 (N315, N304, N159, N143, N261);
xor XOR2 (N316, N311, N104);
buf BUF1 (N317, N284);
not NOT1 (N318, N314);
and AND4 (N319, N315, N278, N17, N33);
not NOT1 (N320, N317);
xor XOR2 (N321, N318, N143);
xor XOR2 (N322, N320, N277);
not NOT1 (N323, N319);
nand NAND3 (N324, N305, N130, N72);
nand NAND3 (N325, N323, N167, N55);
not NOT1 (N326, N321);
not NOT1 (N327, N325);
not NOT1 (N328, N322);
nand NAND3 (N329, N328, N314, N301);
nor NOR2 (N330, N324, N137);
and AND3 (N331, N316, N322, N4);
not NOT1 (N332, N330);
nand NAND2 (N333, N310, N237);
not NOT1 (N334, N295);
and AND3 (N335, N329, N182, N281);
nor NOR3 (N336, N327, N195, N9);
and AND3 (N337, N326, N72, N57);
nand NAND4 (N338, N337, N325, N146, N170);
nor NOR4 (N339, N338, N58, N128, N279);
buf BUF1 (N340, N333);
not NOT1 (N341, N334);
or OR2 (N342, N335, N326);
not NOT1 (N343, N331);
nor NOR3 (N344, N341, N80, N5);
not NOT1 (N345, N332);
nand NAND3 (N346, N342, N14, N44);
nand NAND3 (N347, N313, N122, N94);
not NOT1 (N348, N339);
not NOT1 (N349, N347);
or OR2 (N350, N348, N68);
and AND4 (N351, N345, N349, N331, N286);
buf BUF1 (N352, N231);
buf BUF1 (N353, N343);
and AND2 (N354, N340, N32);
nor NOR2 (N355, N312, N140);
not NOT1 (N356, N336);
and AND3 (N357, N352, N134, N14);
xor XOR2 (N358, N350, N330);
buf BUF1 (N359, N289);
xor XOR2 (N360, N354, N342);
xor XOR2 (N361, N356, N187);
xor XOR2 (N362, N344, N85);
xor XOR2 (N363, N358, N262);
not NOT1 (N364, N359);
buf BUF1 (N365, N357);
and AND4 (N366, N353, N329, N68, N167);
nor NOR3 (N367, N360, N321, N49);
not NOT1 (N368, N346);
nand NAND2 (N369, N361, N223);
buf BUF1 (N370, N363);
or OR3 (N371, N366, N15, N85);
or OR3 (N372, N355, N296, N344);
not NOT1 (N373, N365);
nor NOR3 (N374, N367, N278, N125);
or OR3 (N375, N374, N310, N293);
or OR4 (N376, N364, N350, N19, N284);
and AND3 (N377, N370, N150, N47);
xor XOR2 (N378, N373, N105);
and AND3 (N379, N377, N78, N150);
and AND2 (N380, N362, N366);
nor NOR2 (N381, N375, N36);
buf BUF1 (N382, N376);
nor NOR3 (N383, N351, N216, N152);
and AND2 (N384, N372, N61);
not NOT1 (N385, N380);
nand NAND3 (N386, N371, N68, N217);
nor NOR4 (N387, N386, N288, N208, N219);
not NOT1 (N388, N369);
or OR3 (N389, N383, N257, N309);
nand NAND4 (N390, N387, N347, N89, N301);
xor XOR2 (N391, N368, N235);
or OR2 (N392, N379, N194);
not NOT1 (N393, N388);
xor XOR2 (N394, N391, N22);
nor NOR4 (N395, N382, N223, N84, N327);
not NOT1 (N396, N392);
nand NAND2 (N397, N390, N254);
buf BUF1 (N398, N396);
nor NOR3 (N399, N381, N385, N351);
nor NOR2 (N400, N395, N293);
or OR4 (N401, N98, N119, N344, N335);
nand NAND2 (N402, N397, N138);
and AND3 (N403, N389, N177, N378);
not NOT1 (N404, N257);
buf BUF1 (N405, N403);
and AND4 (N406, N401, N401, N113, N358);
or OR4 (N407, N398, N361, N348, N272);
buf BUF1 (N408, N402);
and AND2 (N409, N400, N10);
xor XOR2 (N410, N409, N92);
not NOT1 (N411, N406);
not NOT1 (N412, N399);
not NOT1 (N413, N393);
nand NAND3 (N414, N384, N394, N192);
and AND2 (N415, N264, N365);
not NOT1 (N416, N414);
nand NAND2 (N417, N413, N23);
not NOT1 (N418, N411);
xor XOR2 (N419, N412, N132);
xor XOR2 (N420, N419, N117);
or OR3 (N421, N415, N81, N358);
or OR4 (N422, N410, N207, N296, N111);
or OR2 (N423, N407, N402);
xor XOR2 (N424, N422, N96);
not NOT1 (N425, N418);
and AND3 (N426, N420, N70, N418);
buf BUF1 (N427, N423);
buf BUF1 (N428, N426);
and AND3 (N429, N404, N165, N317);
or OR3 (N430, N425, N195, N270);
buf BUF1 (N431, N430);
xor XOR2 (N432, N416, N143);
not NOT1 (N433, N428);
and AND4 (N434, N431, N377, N346, N271);
not NOT1 (N435, N421);
not NOT1 (N436, N424);
not NOT1 (N437, N405);
buf BUF1 (N438, N436);
not NOT1 (N439, N427);
nor NOR4 (N440, N438, N86, N30, N337);
not NOT1 (N441, N440);
nand NAND4 (N442, N437, N397, N400, N64);
xor XOR2 (N443, N435, N243);
or OR4 (N444, N429, N109, N156, N159);
xor XOR2 (N445, N444, N238);
nor NOR2 (N446, N445, N143);
or OR3 (N447, N443, N10, N114);
and AND2 (N448, N433, N195);
nand NAND4 (N449, N442, N299, N306, N366);
buf BUF1 (N450, N441);
not NOT1 (N451, N432);
nand NAND4 (N452, N417, N357, N183, N312);
nor NOR4 (N453, N450, N435, N196, N348);
nor NOR3 (N454, N447, N332, N152);
nor NOR4 (N455, N446, N442, N323, N307);
and AND4 (N456, N449, N157, N441, N173);
or OR2 (N457, N434, N168);
and AND2 (N458, N456, N78);
not NOT1 (N459, N439);
nor NOR2 (N460, N451, N190);
or OR4 (N461, N454, N24, N207, N164);
nand NAND4 (N462, N458, N380, N9, N423);
xor XOR2 (N463, N461, N206);
nor NOR3 (N464, N448, N113, N453);
not NOT1 (N465, N370);
not NOT1 (N466, N455);
nand NAND2 (N467, N462, N217);
and AND2 (N468, N465, N356);
or OR3 (N469, N460, N99, N370);
or OR3 (N470, N457, N418, N469);
xor XOR2 (N471, N245, N93);
and AND2 (N472, N463, N107);
or OR4 (N473, N452, N20, N326, N249);
or OR4 (N474, N408, N53, N230, N450);
and AND3 (N475, N471, N319, N78);
buf BUF1 (N476, N468);
nor NOR3 (N477, N464, N1, N2);
or OR3 (N478, N470, N177, N54);
and AND4 (N479, N459, N139, N86, N114);
nand NAND3 (N480, N478, N149, N155);
nand NAND4 (N481, N474, N130, N338, N32);
nand NAND3 (N482, N472, N415, N431);
and AND4 (N483, N476, N199, N196, N192);
nand NAND3 (N484, N466, N141, N160);
or OR2 (N485, N483, N415);
buf BUF1 (N486, N477);
not NOT1 (N487, N484);
nand NAND3 (N488, N487, N220, N210);
and AND2 (N489, N481, N348);
not NOT1 (N490, N486);
or OR2 (N491, N485, N388);
buf BUF1 (N492, N467);
nor NOR3 (N493, N473, N86, N110);
not NOT1 (N494, N480);
xor XOR2 (N495, N489, N120);
and AND3 (N496, N482, N171, N429);
nor NOR4 (N497, N479, N325, N367, N48);
nand NAND3 (N498, N497, N107, N113);
buf BUF1 (N499, N493);
and AND4 (N500, N494, N371, N53, N448);
buf BUF1 (N501, N495);
xor XOR2 (N502, N490, N263);
nand NAND3 (N503, N498, N86, N266);
and AND3 (N504, N499, N480, N106);
nor NOR4 (N505, N502, N112, N144, N3);
not NOT1 (N506, N501);
buf BUF1 (N507, N503);
xor XOR2 (N508, N507, N190);
or OR3 (N509, N475, N485, N178);
buf BUF1 (N510, N509);
not NOT1 (N511, N504);
buf BUF1 (N512, N488);
nor NOR2 (N513, N510, N234);
not NOT1 (N514, N496);
nand NAND3 (N515, N491, N18, N283);
nand NAND2 (N516, N513, N347);
xor XOR2 (N517, N512, N211);
and AND3 (N518, N508, N489, N290);
nand NAND3 (N519, N516, N17, N330);
not NOT1 (N520, N515);
not NOT1 (N521, N505);
and AND4 (N522, N511, N85, N289, N134);
endmodule