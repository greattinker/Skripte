// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N3507,N3515,N3503,N3512,N3502,N3509,N3510,N3506,N3514,N3516;

nand NAND2 (N17, N2, N14);
nor NOR3 (N18, N5, N13, N3);
xor XOR2 (N19, N16, N18);
and AND2 (N20, N2, N7);
or OR4 (N21, N5, N7, N13, N13);
or OR4 (N22, N20, N14, N4, N18);
xor XOR2 (N23, N16, N21);
or OR3 (N24, N17, N17, N16);
buf BUF1 (N25, N11);
buf BUF1 (N26, N4);
and AND4 (N27, N24, N2, N2, N13);
nand NAND4 (N28, N25, N16, N11, N8);
nor NOR3 (N29, N2, N7, N8);
or OR2 (N30, N23, N3);
or OR3 (N31, N19, N18, N16);
xor XOR2 (N32, N9, N18);
nand NAND2 (N33, N6, N15);
nand NAND3 (N34, N14, N15, N22);
buf BUF1 (N35, N15);
not NOT1 (N36, N28);
and AND4 (N37, N27, N20, N11, N1);
not NOT1 (N38, N36);
xor XOR2 (N39, N33, N19);
and AND3 (N40, N35, N33, N30);
buf BUF1 (N41, N22);
not NOT1 (N42, N34);
nor NOR3 (N43, N31, N38, N11);
not NOT1 (N44, N6);
or OR2 (N45, N42, N28);
not NOT1 (N46, N41);
or OR4 (N47, N45, N1, N23, N31);
buf BUF1 (N48, N40);
buf BUF1 (N49, N44);
and AND4 (N50, N43, N43, N47, N28);
buf BUF1 (N51, N12);
nand NAND2 (N52, N37, N30);
nand NAND4 (N53, N51, N17, N22, N19);
xor XOR2 (N54, N26, N38);
and AND4 (N55, N52, N27, N12, N51);
xor XOR2 (N56, N49, N4);
not NOT1 (N57, N46);
not NOT1 (N58, N56);
or OR4 (N59, N54, N11, N28, N13);
nor NOR4 (N60, N59, N47, N10, N36);
or OR3 (N61, N50, N21, N19);
or OR3 (N62, N32, N3, N60);
nor NOR4 (N63, N16, N16, N61, N52);
nand NAND2 (N64, N63, N1);
nor NOR4 (N65, N56, N32, N7, N17);
or OR3 (N66, N65, N5, N51);
nor NOR2 (N67, N66, N27);
and AND4 (N68, N53, N16, N29, N1);
not NOT1 (N69, N63);
or OR4 (N70, N39, N59, N1, N39);
not NOT1 (N71, N58);
xor XOR2 (N72, N69, N56);
xor XOR2 (N73, N67, N33);
and AND4 (N74, N55, N16, N10, N16);
nor NOR3 (N75, N62, N13, N22);
not NOT1 (N76, N74);
nor NOR4 (N77, N64, N56, N11, N74);
nand NAND4 (N78, N48, N28, N13, N69);
buf BUF1 (N79, N73);
and AND3 (N80, N75, N75, N54);
or OR3 (N81, N77, N64, N42);
buf BUF1 (N82, N76);
or OR3 (N83, N79, N41, N27);
or OR3 (N84, N68, N18, N70);
nand NAND4 (N85, N46, N45, N79, N16);
or OR2 (N86, N81, N27);
nor NOR2 (N87, N78, N53);
buf BUF1 (N88, N80);
xor XOR2 (N89, N87, N88);
nand NAND2 (N90, N34, N48);
xor XOR2 (N91, N84, N58);
nand NAND3 (N92, N72, N79, N87);
not NOT1 (N93, N92);
not NOT1 (N94, N82);
or OR4 (N95, N86, N7, N57, N19);
nor NOR2 (N96, N31, N74);
nor NOR2 (N97, N91, N53);
buf BUF1 (N98, N83);
xor XOR2 (N99, N93, N22);
not NOT1 (N100, N94);
nor NOR3 (N101, N89, N73, N83);
buf BUF1 (N102, N90);
nand NAND3 (N103, N102, N76, N88);
nor NOR2 (N104, N85, N63);
buf BUF1 (N105, N95);
nand NAND3 (N106, N98, N96, N77);
xor XOR2 (N107, N85, N44);
or OR3 (N108, N103, N72, N56);
or OR4 (N109, N97, N6, N74, N85);
buf BUF1 (N110, N109);
nand NAND3 (N111, N99, N18, N22);
not NOT1 (N112, N106);
nor NOR2 (N113, N108, N41);
buf BUF1 (N114, N110);
buf BUF1 (N115, N114);
nor NOR4 (N116, N71, N78, N92, N22);
xor XOR2 (N117, N107, N25);
and AND4 (N118, N116, N43, N92, N56);
not NOT1 (N119, N118);
nand NAND2 (N120, N112, N73);
nor NOR4 (N121, N115, N51, N105, N65);
and AND2 (N122, N39, N92);
not NOT1 (N123, N117);
nand NAND4 (N124, N120, N57, N3, N111);
and AND4 (N125, N81, N123, N73, N43);
nor NOR4 (N126, N8, N107, N7, N106);
nor NOR2 (N127, N100, N51);
nand NAND3 (N128, N121, N97, N115);
nor NOR2 (N129, N113, N23);
nor NOR4 (N130, N127, N76, N115, N39);
nor NOR4 (N131, N101, N37, N45, N98);
xor XOR2 (N132, N124, N70);
buf BUF1 (N133, N129);
nand NAND4 (N134, N122, N26, N13, N102);
and AND2 (N135, N126, N75);
not NOT1 (N136, N130);
not NOT1 (N137, N132);
nor NOR2 (N138, N133, N117);
buf BUF1 (N139, N125);
nand NAND2 (N140, N139, N63);
buf BUF1 (N141, N119);
or OR3 (N142, N140, N78, N120);
not NOT1 (N143, N104);
xor XOR2 (N144, N143, N50);
and AND2 (N145, N136, N17);
nand NAND2 (N146, N141, N37);
nor NOR3 (N147, N131, N32, N84);
nand NAND4 (N148, N147, N81, N77, N135);
buf BUF1 (N149, N61);
not NOT1 (N150, N144);
or OR2 (N151, N148, N150);
or OR3 (N152, N134, N16, N92);
not NOT1 (N153, N47);
nand NAND4 (N154, N128, N136, N100, N28);
or OR4 (N155, N151, N114, N78, N62);
and AND4 (N156, N155, N106, N43, N125);
xor XOR2 (N157, N149, N26);
xor XOR2 (N158, N146, N19);
nor NOR2 (N159, N137, N110);
and AND2 (N160, N154, N85);
or OR2 (N161, N152, N127);
xor XOR2 (N162, N158, N160);
buf BUF1 (N163, N37);
nand NAND4 (N164, N138, N35, N115, N116);
nor NOR3 (N165, N162, N84, N143);
or OR4 (N166, N161, N71, N117, N98);
nor NOR2 (N167, N159, N114);
or OR3 (N168, N167, N164, N149);
buf BUF1 (N169, N109);
or OR3 (N170, N145, N91, N68);
buf BUF1 (N171, N170);
nor NOR3 (N172, N166, N15, N80);
not NOT1 (N173, N169);
xor XOR2 (N174, N165, N169);
buf BUF1 (N175, N172);
and AND3 (N176, N171, N95, N28);
not NOT1 (N177, N163);
or OR2 (N178, N142, N161);
xor XOR2 (N179, N177, N57);
xor XOR2 (N180, N153, N112);
nand NAND2 (N181, N156, N62);
nor NOR4 (N182, N174, N47, N1, N52);
or OR4 (N183, N168, N9, N171, N107);
nor NOR2 (N184, N176, N132);
and AND2 (N185, N181, N66);
or OR4 (N186, N184, N150, N98, N119);
buf BUF1 (N187, N157);
and AND2 (N188, N173, N35);
nor NOR2 (N189, N187, N114);
xor XOR2 (N190, N186, N9);
buf BUF1 (N191, N180);
not NOT1 (N192, N182);
buf BUF1 (N193, N190);
buf BUF1 (N194, N175);
buf BUF1 (N195, N192);
xor XOR2 (N196, N179, N49);
xor XOR2 (N197, N191, N195);
nor NOR3 (N198, N176, N122, N172);
nand NAND4 (N199, N196, N168, N28, N46);
nand NAND4 (N200, N185, N101, N77, N114);
xor XOR2 (N201, N193, N87);
xor XOR2 (N202, N197, N60);
or OR2 (N203, N198, N89);
not NOT1 (N204, N199);
buf BUF1 (N205, N178);
buf BUF1 (N206, N189);
or OR3 (N207, N202, N109, N39);
xor XOR2 (N208, N201, N10);
nand NAND2 (N209, N205, N142);
xor XOR2 (N210, N188, N59);
nor NOR3 (N211, N210, N209, N1);
and AND3 (N212, N74, N137, N4);
nand NAND2 (N213, N194, N149);
xor XOR2 (N214, N206, N156);
buf BUF1 (N215, N204);
xor XOR2 (N216, N214, N41);
and AND3 (N217, N207, N198, N165);
xor XOR2 (N218, N208, N178);
and AND4 (N219, N213, N62, N37, N100);
xor XOR2 (N220, N218, N134);
buf BUF1 (N221, N211);
buf BUF1 (N222, N216);
xor XOR2 (N223, N203, N130);
xor XOR2 (N224, N223, N100);
not NOT1 (N225, N215);
or OR4 (N226, N183, N51, N91, N155);
or OR4 (N227, N221, N162, N96, N48);
xor XOR2 (N228, N227, N153);
buf BUF1 (N229, N200);
nand NAND3 (N230, N226, N25, N27);
buf BUF1 (N231, N219);
nor NOR4 (N232, N220, N219, N170, N65);
buf BUF1 (N233, N225);
nor NOR2 (N234, N217, N224);
nor NOR3 (N235, N49, N8, N48);
xor XOR2 (N236, N231, N88);
or OR2 (N237, N212, N49);
buf BUF1 (N238, N235);
not NOT1 (N239, N236);
buf BUF1 (N240, N229);
nand NAND4 (N241, N232, N128, N152, N125);
nand NAND2 (N242, N230, N152);
buf BUF1 (N243, N237);
nand NAND3 (N244, N242, N36, N212);
nand NAND4 (N245, N233, N242, N104, N191);
nor NOR2 (N246, N243, N53);
nand NAND4 (N247, N240, N226, N233, N201);
nand NAND4 (N248, N246, N11, N199, N52);
or OR4 (N249, N247, N207, N72, N185);
buf BUF1 (N250, N239);
not NOT1 (N251, N249);
and AND4 (N252, N250, N24, N249, N137);
nor NOR4 (N253, N244, N54, N132, N82);
nor NOR4 (N254, N252, N194, N145, N84);
not NOT1 (N255, N245);
xor XOR2 (N256, N241, N42);
nand NAND2 (N257, N255, N154);
not NOT1 (N258, N248);
and AND3 (N259, N234, N119, N214);
and AND3 (N260, N222, N110, N19);
or OR4 (N261, N238, N40, N49, N40);
xor XOR2 (N262, N258, N256);
xor XOR2 (N263, N145, N135);
or OR3 (N264, N257, N158, N187);
nor NOR3 (N265, N253, N232, N118);
nor NOR3 (N266, N259, N83, N151);
or OR4 (N267, N265, N76, N144, N67);
not NOT1 (N268, N267);
nor NOR4 (N269, N268, N257, N11, N256);
nor NOR3 (N270, N263, N180, N170);
not NOT1 (N271, N260);
xor XOR2 (N272, N264, N205);
not NOT1 (N273, N270);
and AND2 (N274, N271, N14);
or OR4 (N275, N262, N150, N11, N80);
and AND3 (N276, N274, N63, N135);
nand NAND2 (N277, N276, N121);
and AND2 (N278, N277, N220);
buf BUF1 (N279, N273);
or OR4 (N280, N278, N276, N86, N251);
xor XOR2 (N281, N247, N131);
nor NOR3 (N282, N228, N69, N127);
buf BUF1 (N283, N272);
and AND2 (N284, N266, N136);
buf BUF1 (N285, N284);
buf BUF1 (N286, N280);
and AND3 (N287, N283, N167, N284);
xor XOR2 (N288, N281, N38);
nor NOR2 (N289, N269, N51);
nand NAND3 (N290, N289, N59, N197);
buf BUF1 (N291, N288);
not NOT1 (N292, N286);
or OR2 (N293, N282, N286);
nand NAND2 (N294, N290, N206);
buf BUF1 (N295, N279);
nand NAND2 (N296, N293, N140);
nor NOR4 (N297, N285, N97, N219, N176);
buf BUF1 (N298, N295);
nor NOR2 (N299, N294, N160);
not NOT1 (N300, N297);
nand NAND4 (N301, N296, N293, N28, N185);
nor NOR4 (N302, N292, N295, N140, N177);
nand NAND4 (N303, N302, N169, N65, N205);
xor XOR2 (N304, N298, N159);
xor XOR2 (N305, N291, N128);
and AND2 (N306, N299, N80);
nand NAND4 (N307, N305, N278, N104, N36);
xor XOR2 (N308, N275, N184);
not NOT1 (N309, N303);
xor XOR2 (N310, N300, N128);
buf BUF1 (N311, N254);
nand NAND2 (N312, N308, N274);
buf BUF1 (N313, N301);
buf BUF1 (N314, N311);
and AND4 (N315, N313, N104, N108, N21);
xor XOR2 (N316, N309, N315);
nor NOR4 (N317, N268, N316, N184, N145);
xor XOR2 (N318, N155, N209);
xor XOR2 (N319, N304, N86);
nor NOR3 (N320, N306, N248, N190);
nor NOR4 (N321, N310, N269, N148, N206);
or OR3 (N322, N319, N8, N231);
buf BUF1 (N323, N318);
not NOT1 (N324, N312);
xor XOR2 (N325, N261, N155);
and AND3 (N326, N314, N235, N209);
not NOT1 (N327, N326);
buf BUF1 (N328, N327);
xor XOR2 (N329, N321, N199);
nand NAND4 (N330, N317, N122, N90, N229);
nor NOR2 (N331, N325, N296);
or OR3 (N332, N331, N21, N268);
and AND3 (N333, N322, N279, N148);
not NOT1 (N334, N307);
buf BUF1 (N335, N320);
nand NAND3 (N336, N330, N192, N160);
and AND2 (N337, N334, N315);
not NOT1 (N338, N323);
nand NAND2 (N339, N338, N115);
or OR3 (N340, N332, N2, N299);
xor XOR2 (N341, N324, N307);
xor XOR2 (N342, N335, N322);
not NOT1 (N343, N341);
buf BUF1 (N344, N340);
nand NAND3 (N345, N344, N62, N74);
buf BUF1 (N346, N328);
or OR4 (N347, N337, N95, N279, N245);
and AND3 (N348, N336, N310, N38);
nor NOR2 (N349, N329, N282);
nand NAND3 (N350, N339, N10, N140);
not NOT1 (N351, N343);
nor NOR2 (N352, N346, N102);
xor XOR2 (N353, N333, N310);
xor XOR2 (N354, N349, N221);
xor XOR2 (N355, N348, N20);
xor XOR2 (N356, N345, N119);
and AND3 (N357, N354, N22, N140);
xor XOR2 (N358, N287, N223);
buf BUF1 (N359, N357);
buf BUF1 (N360, N356);
nand NAND3 (N361, N351, N88, N202);
nand NAND2 (N362, N350, N119);
nand NAND3 (N363, N359, N353, N188);
nand NAND3 (N364, N283, N286, N253);
nor NOR2 (N365, N360, N133);
not NOT1 (N366, N342);
nor NOR4 (N367, N352, N301, N80, N246);
nand NAND3 (N368, N365, N235, N28);
buf BUF1 (N369, N366);
xor XOR2 (N370, N355, N165);
and AND2 (N371, N367, N366);
or OR2 (N372, N361, N145);
and AND3 (N373, N347, N5, N206);
not NOT1 (N374, N370);
nand NAND2 (N375, N373, N61);
nor NOR3 (N376, N358, N7, N322);
nand NAND4 (N377, N376, N276, N114, N324);
nand NAND3 (N378, N362, N313, N106);
nor NOR3 (N379, N378, N211, N20);
not NOT1 (N380, N379);
and AND3 (N381, N371, N252, N314);
and AND4 (N382, N369, N160, N95, N163);
buf BUF1 (N383, N380);
or OR2 (N384, N381, N234);
buf BUF1 (N385, N363);
not NOT1 (N386, N372);
and AND3 (N387, N384, N296, N144);
and AND4 (N388, N383, N131, N319, N263);
nor NOR3 (N389, N385, N383, N289);
not NOT1 (N390, N364);
xor XOR2 (N391, N386, N265);
buf BUF1 (N392, N374);
not NOT1 (N393, N387);
or OR2 (N394, N377, N180);
nor NOR3 (N395, N382, N150, N146);
nor NOR3 (N396, N390, N383, N178);
or OR4 (N397, N396, N76, N128, N140);
xor XOR2 (N398, N375, N256);
buf BUF1 (N399, N389);
xor XOR2 (N400, N391, N259);
xor XOR2 (N401, N397, N28);
nor NOR4 (N402, N368, N401, N6, N95);
and AND4 (N403, N108, N346, N218, N310);
and AND3 (N404, N388, N315, N14);
buf BUF1 (N405, N394);
nor NOR2 (N406, N403, N116);
not NOT1 (N407, N393);
not NOT1 (N408, N405);
nand NAND2 (N409, N404, N102);
nand NAND4 (N410, N399, N335, N53, N347);
buf BUF1 (N411, N398);
or OR2 (N412, N407, N323);
buf BUF1 (N413, N406);
not NOT1 (N414, N410);
nand NAND2 (N415, N414, N33);
or OR2 (N416, N392, N263);
xor XOR2 (N417, N408, N286);
nand NAND3 (N418, N402, N162, N273);
nand NAND2 (N419, N409, N195);
and AND2 (N420, N400, N3);
xor XOR2 (N421, N419, N344);
nand NAND2 (N422, N416, N244);
nor NOR2 (N423, N421, N192);
not NOT1 (N424, N412);
or OR2 (N425, N411, N61);
not NOT1 (N426, N415);
nor NOR2 (N427, N420, N300);
buf BUF1 (N428, N424);
nand NAND2 (N429, N423, N309);
nor NOR2 (N430, N425, N255);
buf BUF1 (N431, N413);
nor NOR2 (N432, N427, N7);
or OR3 (N433, N422, N365, N342);
and AND3 (N434, N395, N136, N101);
and AND3 (N435, N418, N409, N310);
not NOT1 (N436, N426);
xor XOR2 (N437, N430, N362);
xor XOR2 (N438, N433, N5);
nor NOR4 (N439, N436, N397, N17, N102);
and AND2 (N440, N435, N165);
and AND3 (N441, N431, N346, N415);
buf BUF1 (N442, N429);
xor XOR2 (N443, N434, N361);
nand NAND4 (N444, N437, N222, N204, N373);
nand NAND4 (N445, N439, N341, N60, N119);
not NOT1 (N446, N445);
or OR2 (N447, N446, N179);
not NOT1 (N448, N444);
not NOT1 (N449, N440);
buf BUF1 (N450, N449);
or OR4 (N451, N442, N351, N300, N296);
and AND3 (N452, N428, N187, N303);
nand NAND2 (N453, N443, N246);
and AND2 (N454, N453, N438);
nor NOR4 (N455, N5, N425, N98, N299);
buf BUF1 (N456, N441);
nand NAND2 (N457, N447, N34);
xor XOR2 (N458, N457, N216);
or OR4 (N459, N454, N270, N428, N362);
and AND2 (N460, N432, N295);
and AND4 (N461, N459, N250, N213, N301);
xor XOR2 (N462, N456, N80);
nor NOR4 (N463, N461, N399, N81, N299);
nor NOR2 (N464, N452, N10);
nor NOR2 (N465, N417, N257);
and AND4 (N466, N451, N228, N51, N375);
or OR3 (N467, N460, N40, N205);
nor NOR3 (N468, N448, N342, N395);
xor XOR2 (N469, N458, N237);
nand NAND2 (N470, N467, N31);
xor XOR2 (N471, N466, N113);
nand NAND2 (N472, N469, N42);
xor XOR2 (N473, N463, N264);
nor NOR3 (N474, N464, N17, N109);
and AND4 (N475, N468, N182, N356, N7);
xor XOR2 (N476, N450, N155);
not NOT1 (N477, N470);
nor NOR3 (N478, N475, N403, N288);
xor XOR2 (N479, N474, N57);
and AND4 (N480, N465, N211, N346, N113);
xor XOR2 (N481, N472, N437);
or OR4 (N482, N476, N46, N185, N8);
not NOT1 (N483, N478);
or OR3 (N484, N473, N88, N372);
and AND2 (N485, N471, N355);
and AND4 (N486, N462, N58, N226, N258);
nand NAND3 (N487, N455, N357, N102);
nor NOR2 (N488, N479, N150);
and AND4 (N489, N484, N404, N17, N348);
xor XOR2 (N490, N489, N216);
and AND4 (N491, N485, N17, N223, N448);
nor NOR3 (N492, N481, N336, N416);
and AND3 (N493, N477, N94, N260);
nand NAND2 (N494, N490, N140);
nor NOR3 (N495, N482, N491, N418);
xor XOR2 (N496, N335, N287);
nand NAND4 (N497, N488, N299, N314, N362);
or OR4 (N498, N496, N192, N330, N28);
not NOT1 (N499, N492);
or OR2 (N500, N483, N50);
or OR2 (N501, N486, N450);
not NOT1 (N502, N480);
nand NAND3 (N503, N500, N313, N176);
or OR4 (N504, N501, N412, N104, N459);
not NOT1 (N505, N494);
not NOT1 (N506, N504);
nand NAND4 (N507, N503, N375, N16, N303);
xor XOR2 (N508, N502, N280);
or OR2 (N509, N499, N124);
and AND2 (N510, N495, N190);
not NOT1 (N511, N493);
not NOT1 (N512, N508);
xor XOR2 (N513, N510, N247);
and AND3 (N514, N511, N163, N267);
or OR2 (N515, N505, N22);
or OR2 (N516, N514, N428);
or OR4 (N517, N506, N390, N468, N437);
nand NAND4 (N518, N517, N472, N517, N479);
nor NOR4 (N519, N512, N232, N114, N201);
nor NOR3 (N520, N507, N393, N302);
buf BUF1 (N521, N487);
xor XOR2 (N522, N515, N442);
and AND4 (N523, N521, N174, N429, N515);
xor XOR2 (N524, N522, N402);
nand NAND2 (N525, N524, N485);
xor XOR2 (N526, N497, N506);
nand NAND2 (N527, N498, N183);
nand NAND3 (N528, N526, N365, N471);
nand NAND3 (N529, N523, N223, N514);
not NOT1 (N530, N529);
buf BUF1 (N531, N519);
nor NOR2 (N532, N525, N184);
nor NOR3 (N533, N530, N307, N155);
nand NAND3 (N534, N520, N495, N357);
buf BUF1 (N535, N533);
xor XOR2 (N536, N527, N464);
buf BUF1 (N537, N516);
nand NAND4 (N538, N537, N191, N362, N454);
xor XOR2 (N539, N531, N469);
nand NAND2 (N540, N534, N376);
xor XOR2 (N541, N532, N45);
buf BUF1 (N542, N518);
or OR3 (N543, N536, N174, N183);
or OR3 (N544, N543, N3, N238);
buf BUF1 (N545, N538);
nor NOR2 (N546, N539, N325);
xor XOR2 (N547, N528, N153);
and AND2 (N548, N541, N81);
or OR2 (N549, N544, N239);
nand NAND2 (N550, N535, N491);
not NOT1 (N551, N509);
xor XOR2 (N552, N545, N543);
xor XOR2 (N553, N540, N1);
not NOT1 (N554, N550);
not NOT1 (N555, N548);
or OR3 (N556, N552, N337, N289);
nand NAND3 (N557, N546, N429, N379);
not NOT1 (N558, N556);
nand NAND4 (N559, N547, N34, N438, N352);
nor NOR3 (N560, N542, N551, N12);
buf BUF1 (N561, N53);
nand NAND3 (N562, N560, N552, N393);
or OR4 (N563, N549, N283, N231, N558);
nand NAND2 (N564, N464, N159);
nor NOR3 (N565, N564, N558, N563);
not NOT1 (N566, N403);
and AND4 (N567, N566, N387, N512, N371);
nor NOR2 (N568, N555, N159);
or OR4 (N569, N562, N213, N338, N353);
buf BUF1 (N570, N553);
or OR2 (N571, N557, N537);
or OR2 (N572, N570, N507);
xor XOR2 (N573, N568, N306);
and AND3 (N574, N573, N535, N517);
or OR3 (N575, N554, N159, N225);
buf BUF1 (N576, N561);
nand NAND4 (N577, N559, N277, N221, N102);
not NOT1 (N578, N571);
or OR4 (N579, N574, N285, N250, N254);
nand NAND2 (N580, N572, N554);
or OR4 (N581, N567, N227, N208, N34);
or OR4 (N582, N579, N494, N176, N312);
nor NOR2 (N583, N577, N552);
xor XOR2 (N584, N513, N3);
buf BUF1 (N585, N580);
not NOT1 (N586, N583);
nand NAND3 (N587, N582, N439, N490);
not NOT1 (N588, N565);
xor XOR2 (N589, N588, N149);
not NOT1 (N590, N576);
nor NOR2 (N591, N578, N507);
buf BUF1 (N592, N575);
not NOT1 (N593, N569);
nand NAND4 (N594, N587, N53, N257, N473);
or OR3 (N595, N581, N285, N471);
nor NOR4 (N596, N584, N38, N570, N398);
nand NAND4 (N597, N595, N145, N524, N283);
not NOT1 (N598, N591);
xor XOR2 (N599, N592, N204);
not NOT1 (N600, N599);
or OR2 (N601, N596, N40);
not NOT1 (N602, N593);
and AND4 (N603, N602, N291, N539, N308);
nand NAND4 (N604, N597, N594, N536, N11);
nand NAND2 (N605, N351, N352);
buf BUF1 (N606, N603);
and AND3 (N607, N604, N262, N383);
nor NOR3 (N608, N598, N532, N594);
nand NAND4 (N609, N605, N210, N193, N218);
nand NAND2 (N610, N585, N606);
xor XOR2 (N611, N475, N192);
or OR4 (N612, N600, N386, N407, N370);
nor NOR3 (N613, N586, N230, N531);
buf BUF1 (N614, N610);
xor XOR2 (N615, N614, N571);
or OR3 (N616, N612, N391, N242);
xor XOR2 (N617, N607, N250);
xor XOR2 (N618, N617, N313);
buf BUF1 (N619, N616);
and AND4 (N620, N609, N484, N57, N506);
and AND4 (N621, N611, N452, N364, N403);
nand NAND4 (N622, N590, N73, N478, N326);
xor XOR2 (N623, N613, N375);
and AND4 (N624, N615, N65, N76, N202);
nor NOR3 (N625, N608, N97, N501);
not NOT1 (N626, N601);
not NOT1 (N627, N624);
nand NAND3 (N628, N621, N230, N504);
xor XOR2 (N629, N627, N292);
xor XOR2 (N630, N589, N603);
or OR4 (N631, N630, N593, N504, N599);
nand NAND3 (N632, N622, N336, N560);
or OR3 (N633, N618, N281, N597);
buf BUF1 (N634, N628);
buf BUF1 (N635, N629);
nand NAND3 (N636, N635, N602, N393);
xor XOR2 (N637, N631, N261);
nand NAND2 (N638, N637, N556);
buf BUF1 (N639, N620);
nand NAND2 (N640, N639, N609);
or OR3 (N641, N619, N441, N586);
nand NAND2 (N642, N625, N470);
buf BUF1 (N643, N623);
nand NAND2 (N644, N636, N529);
xor XOR2 (N645, N640, N445);
nand NAND3 (N646, N638, N328, N266);
not NOT1 (N647, N644);
buf BUF1 (N648, N634);
or OR3 (N649, N626, N526, N430);
nand NAND2 (N650, N646, N466);
nand NAND3 (N651, N632, N560, N194);
nand NAND2 (N652, N633, N172);
and AND3 (N653, N651, N160, N170);
xor XOR2 (N654, N647, N652);
nand NAND4 (N655, N113, N10, N270, N619);
xor XOR2 (N656, N643, N344);
and AND4 (N657, N655, N121, N143, N340);
and AND4 (N658, N650, N251, N467, N74);
xor XOR2 (N659, N657, N59);
nor NOR3 (N660, N654, N12, N495);
nor NOR2 (N661, N660, N348);
and AND2 (N662, N649, N55);
buf BUF1 (N663, N642);
buf BUF1 (N664, N648);
buf BUF1 (N665, N645);
buf BUF1 (N666, N663);
buf BUF1 (N667, N662);
nor NOR2 (N668, N665, N41);
buf BUF1 (N669, N664);
xor XOR2 (N670, N658, N624);
xor XOR2 (N671, N641, N562);
and AND2 (N672, N669, N376);
nand NAND4 (N673, N661, N166, N576, N404);
nor NOR3 (N674, N672, N668, N53);
and AND2 (N675, N304, N81);
and AND4 (N676, N667, N609, N370, N476);
or OR2 (N677, N675, N271);
buf BUF1 (N678, N677);
and AND4 (N679, N666, N92, N575, N259);
not NOT1 (N680, N678);
nor NOR2 (N681, N679, N493);
and AND3 (N682, N673, N192, N6);
xor XOR2 (N683, N656, N556);
or OR2 (N684, N671, N615);
nand NAND3 (N685, N681, N93, N643);
or OR4 (N686, N676, N455, N208, N243);
nor NOR4 (N687, N659, N175, N441, N577);
buf BUF1 (N688, N685);
nand NAND3 (N689, N682, N626, N511);
buf BUF1 (N690, N653);
or OR3 (N691, N670, N54, N102);
not NOT1 (N692, N684);
buf BUF1 (N693, N683);
and AND2 (N694, N687, N564);
and AND4 (N695, N694, N611, N171, N563);
xor XOR2 (N696, N690, N680);
buf BUF1 (N697, N580);
xor XOR2 (N698, N696, N634);
nand NAND4 (N699, N698, N354, N590, N89);
or OR4 (N700, N689, N608, N661, N36);
nor NOR2 (N701, N674, N268);
xor XOR2 (N702, N688, N486);
buf BUF1 (N703, N692);
not NOT1 (N704, N700);
buf BUF1 (N705, N701);
not NOT1 (N706, N695);
xor XOR2 (N707, N704, N674);
and AND2 (N708, N693, N155);
nand NAND4 (N709, N691, N583, N707, N461);
nor NOR3 (N710, N377, N673, N179);
not NOT1 (N711, N706);
not NOT1 (N712, N699);
or OR4 (N713, N697, N671, N426, N238);
and AND2 (N714, N711, N15);
buf BUF1 (N715, N702);
nand NAND2 (N716, N708, N134);
not NOT1 (N717, N703);
not NOT1 (N718, N709);
or OR4 (N719, N716, N512, N710, N65);
or OR3 (N720, N642, N458, N256);
nor NOR3 (N721, N705, N495, N696);
nand NAND4 (N722, N715, N340, N58, N397);
buf BUF1 (N723, N718);
nor NOR2 (N724, N714, N161);
and AND4 (N725, N717, N416, N51, N118);
or OR3 (N726, N724, N647, N413);
buf BUF1 (N727, N723);
xor XOR2 (N728, N722, N487);
not NOT1 (N729, N726);
not NOT1 (N730, N729);
nand NAND4 (N731, N686, N679, N28, N641);
nor NOR2 (N732, N713, N322);
xor XOR2 (N733, N727, N480);
not NOT1 (N734, N730);
buf BUF1 (N735, N731);
nor NOR3 (N736, N719, N493, N329);
or OR4 (N737, N712, N657, N628, N385);
or OR3 (N738, N734, N247, N323);
xor XOR2 (N739, N720, N108);
xor XOR2 (N740, N739, N525);
and AND4 (N741, N735, N345, N395, N739);
and AND2 (N742, N741, N125);
nand NAND3 (N743, N736, N94, N185);
not NOT1 (N744, N742);
and AND4 (N745, N744, N409, N490, N484);
or OR4 (N746, N728, N443, N563, N713);
not NOT1 (N747, N743);
xor XOR2 (N748, N745, N510);
nand NAND2 (N749, N737, N225);
nand NAND4 (N750, N749, N165, N477, N300);
buf BUF1 (N751, N733);
and AND2 (N752, N750, N75);
buf BUF1 (N753, N748);
and AND2 (N754, N738, N626);
not NOT1 (N755, N751);
buf BUF1 (N756, N732);
nand NAND4 (N757, N755, N281, N329, N90);
xor XOR2 (N758, N721, N556);
buf BUF1 (N759, N746);
or OR4 (N760, N757, N207, N510, N383);
buf BUF1 (N761, N725);
nor NOR3 (N762, N754, N175, N629);
nand NAND2 (N763, N761, N709);
not NOT1 (N764, N760);
xor XOR2 (N765, N740, N328);
nor NOR2 (N766, N762, N207);
not NOT1 (N767, N763);
and AND2 (N768, N759, N78);
xor XOR2 (N769, N756, N213);
nand NAND2 (N770, N768, N6);
or OR4 (N771, N747, N526, N40, N568);
nor NOR4 (N772, N758, N658, N316, N53);
or OR3 (N773, N770, N506, N665);
nand NAND4 (N774, N766, N161, N42, N164);
xor XOR2 (N775, N752, N574);
buf BUF1 (N776, N765);
buf BUF1 (N777, N776);
xor XOR2 (N778, N773, N347);
buf BUF1 (N779, N767);
buf BUF1 (N780, N772);
or OR2 (N781, N769, N698);
nand NAND2 (N782, N779, N286);
xor XOR2 (N783, N780, N781);
nor NOR2 (N784, N501, N631);
and AND4 (N785, N764, N468, N165, N342);
nand NAND4 (N786, N782, N47, N560, N413);
or OR4 (N787, N775, N137, N496, N530);
not NOT1 (N788, N771);
nor NOR2 (N789, N788, N761);
and AND3 (N790, N753, N724, N139);
and AND4 (N791, N790, N554, N570, N680);
buf BUF1 (N792, N784);
buf BUF1 (N793, N777);
buf BUF1 (N794, N778);
xor XOR2 (N795, N794, N788);
nand NAND3 (N796, N793, N291, N740);
not NOT1 (N797, N783);
or OR3 (N798, N797, N724, N682);
and AND3 (N799, N791, N202, N32);
nor NOR3 (N800, N789, N73, N423);
buf BUF1 (N801, N774);
or OR2 (N802, N796, N190);
or OR3 (N803, N802, N345, N167);
not NOT1 (N804, N803);
nand NAND4 (N805, N800, N337, N114, N159);
and AND2 (N806, N798, N325);
xor XOR2 (N807, N806, N73);
xor XOR2 (N808, N799, N200);
xor XOR2 (N809, N795, N622);
and AND4 (N810, N801, N112, N184, N148);
nand NAND4 (N811, N809, N690, N383, N402);
and AND3 (N812, N785, N614, N117);
and AND4 (N813, N804, N404, N509, N807);
not NOT1 (N814, N786);
nand NAND2 (N815, N307, N258);
buf BUF1 (N816, N814);
not NOT1 (N817, N816);
and AND4 (N818, N812, N381, N269, N779);
and AND2 (N819, N787, N411);
not NOT1 (N820, N813);
buf BUF1 (N821, N811);
not NOT1 (N822, N819);
xor XOR2 (N823, N808, N679);
not NOT1 (N824, N805);
or OR4 (N825, N792, N624, N338, N741);
xor XOR2 (N826, N823, N251);
xor XOR2 (N827, N820, N465);
nand NAND3 (N828, N817, N671, N687);
or OR4 (N829, N824, N554, N637, N406);
nor NOR4 (N830, N827, N130, N444, N95);
xor XOR2 (N831, N830, N800);
not NOT1 (N832, N829);
nor NOR4 (N833, N828, N285, N443, N177);
not NOT1 (N834, N818);
not NOT1 (N835, N821);
not NOT1 (N836, N810);
xor XOR2 (N837, N822, N834);
and AND2 (N838, N287, N356);
buf BUF1 (N839, N833);
not NOT1 (N840, N838);
and AND3 (N841, N839, N749, N687);
buf BUF1 (N842, N840);
xor XOR2 (N843, N825, N705);
not NOT1 (N844, N815);
nand NAND4 (N845, N826, N805, N183, N620);
buf BUF1 (N846, N835);
nand NAND2 (N847, N841, N615);
nor NOR4 (N848, N843, N255, N153, N10);
not NOT1 (N849, N846);
buf BUF1 (N850, N832);
and AND3 (N851, N848, N481, N622);
not NOT1 (N852, N845);
and AND4 (N853, N849, N229, N250, N88);
not NOT1 (N854, N837);
or OR2 (N855, N844, N391);
not NOT1 (N856, N853);
xor XOR2 (N857, N836, N426);
buf BUF1 (N858, N854);
xor XOR2 (N859, N831, N549);
nand NAND2 (N860, N850, N480);
buf BUF1 (N861, N847);
and AND3 (N862, N852, N721, N362);
buf BUF1 (N863, N856);
not NOT1 (N864, N862);
buf BUF1 (N865, N851);
not NOT1 (N866, N858);
xor XOR2 (N867, N857, N161);
nor NOR3 (N868, N859, N824, N588);
or OR4 (N869, N868, N58, N717, N688);
or OR4 (N870, N867, N276, N652, N28);
not NOT1 (N871, N870);
nor NOR3 (N872, N864, N762, N677);
or OR4 (N873, N863, N813, N251, N640);
buf BUF1 (N874, N865);
or OR3 (N875, N860, N534, N268);
and AND4 (N876, N875, N142, N372, N35);
not NOT1 (N877, N874);
nor NOR3 (N878, N866, N331, N534);
nor NOR4 (N879, N878, N412, N101, N711);
nand NAND4 (N880, N879, N571, N288, N566);
buf BUF1 (N881, N842);
and AND4 (N882, N871, N7, N303, N567);
buf BUF1 (N883, N861);
or OR4 (N884, N869, N191, N187, N250);
and AND3 (N885, N877, N178, N553);
or OR3 (N886, N880, N500, N847);
nor NOR4 (N887, N883, N53, N645, N819);
nor NOR2 (N888, N873, N687);
and AND3 (N889, N881, N287, N397);
and AND4 (N890, N855, N486, N179, N311);
or OR3 (N891, N890, N410, N880);
not NOT1 (N892, N886);
not NOT1 (N893, N892);
or OR3 (N894, N888, N247, N161);
nand NAND4 (N895, N891, N104, N555, N564);
not NOT1 (N896, N882);
not NOT1 (N897, N872);
nand NAND4 (N898, N889, N709, N560, N267);
nand NAND4 (N899, N887, N891, N673, N513);
not NOT1 (N900, N894);
buf BUF1 (N901, N898);
buf BUF1 (N902, N876);
not NOT1 (N903, N902);
buf BUF1 (N904, N901);
buf BUF1 (N905, N893);
or OR4 (N906, N896, N467, N71, N114);
nor NOR3 (N907, N899, N805, N520);
and AND3 (N908, N905, N516, N288);
not NOT1 (N909, N907);
buf BUF1 (N910, N885);
buf BUF1 (N911, N906);
not NOT1 (N912, N897);
buf BUF1 (N913, N911);
nand NAND4 (N914, N903, N602, N258, N328);
buf BUF1 (N915, N909);
not NOT1 (N916, N913);
or OR3 (N917, N904, N275, N131);
not NOT1 (N918, N917);
xor XOR2 (N919, N916, N9);
and AND4 (N920, N914, N146, N258, N409);
nand NAND3 (N921, N910, N135, N792);
nand NAND4 (N922, N912, N447, N714, N544);
nand NAND3 (N923, N920, N752, N742);
nor NOR2 (N924, N884, N465);
and AND3 (N925, N919, N631, N511);
nand NAND2 (N926, N925, N468);
and AND2 (N927, N924, N728);
nand NAND2 (N928, N915, N234);
buf BUF1 (N929, N900);
not NOT1 (N930, N928);
xor XOR2 (N931, N930, N593);
and AND4 (N932, N929, N920, N819, N879);
buf BUF1 (N933, N908);
nand NAND3 (N934, N922, N607, N795);
not NOT1 (N935, N895);
nand NAND2 (N936, N933, N467);
nor NOR3 (N937, N936, N330, N820);
nor NOR3 (N938, N923, N818, N453);
or OR2 (N939, N918, N506);
nand NAND4 (N940, N938, N236, N306, N866);
nor NOR2 (N941, N935, N580);
nor NOR2 (N942, N940, N570);
nand NAND2 (N943, N921, N416);
xor XOR2 (N944, N934, N414);
xor XOR2 (N945, N931, N284);
and AND2 (N946, N937, N823);
buf BUF1 (N947, N941);
buf BUF1 (N948, N946);
buf BUF1 (N949, N939);
xor XOR2 (N950, N943, N652);
buf BUF1 (N951, N948);
and AND2 (N952, N926, N496);
xor XOR2 (N953, N927, N762);
or OR3 (N954, N945, N913, N698);
nor NOR3 (N955, N952, N101, N635);
nand NAND2 (N956, N950, N768);
xor XOR2 (N957, N944, N418);
or OR3 (N958, N947, N940, N876);
nand NAND4 (N959, N949, N338, N388, N560);
xor XOR2 (N960, N958, N166);
and AND3 (N961, N953, N400, N449);
buf BUF1 (N962, N957);
buf BUF1 (N963, N959);
or OR4 (N964, N942, N888, N607, N807);
and AND3 (N965, N951, N176, N452);
buf BUF1 (N966, N964);
or OR3 (N967, N961, N172, N656);
not NOT1 (N968, N955);
nand NAND4 (N969, N968, N293, N888, N628);
or OR3 (N970, N969, N739, N368);
nor NOR4 (N971, N954, N515, N512, N305);
nand NAND2 (N972, N932, N88);
or OR2 (N973, N971, N9);
nand NAND4 (N974, N965, N121, N938, N543);
or OR2 (N975, N956, N685);
or OR3 (N976, N960, N247, N334);
nand NAND2 (N977, N967, N730);
or OR2 (N978, N976, N522);
nand NAND2 (N979, N978, N248);
or OR2 (N980, N975, N399);
or OR4 (N981, N972, N296, N319, N162);
nand NAND4 (N982, N977, N944, N355, N90);
or OR2 (N983, N982, N430);
not NOT1 (N984, N966);
or OR2 (N985, N979, N222);
or OR4 (N986, N963, N311, N126, N973);
nand NAND2 (N987, N141, N948);
nor NOR2 (N988, N984, N486);
nor NOR2 (N989, N980, N495);
and AND4 (N990, N962, N361, N188, N274);
or OR4 (N991, N985, N819, N740, N842);
nand NAND4 (N992, N989, N588, N366, N788);
not NOT1 (N993, N986);
not NOT1 (N994, N981);
nor NOR2 (N995, N990, N200);
not NOT1 (N996, N974);
nor NOR4 (N997, N994, N392, N172, N706);
nand NAND3 (N998, N983, N356, N111);
xor XOR2 (N999, N996, N444);
xor XOR2 (N1000, N987, N944);
nor NOR3 (N1001, N997, N374, N254);
buf BUF1 (N1002, N1001);
and AND2 (N1003, N998, N873);
nor NOR3 (N1004, N1002, N956, N503);
xor XOR2 (N1005, N1003, N990);
and AND2 (N1006, N1000, N511);
or OR4 (N1007, N993, N289, N306, N560);
and AND3 (N1008, N995, N449, N777);
nand NAND2 (N1009, N1004, N621);
xor XOR2 (N1010, N999, N288);
nand NAND2 (N1011, N1009, N762);
not NOT1 (N1012, N970);
xor XOR2 (N1013, N992, N171);
nor NOR4 (N1014, N1005, N27, N204, N733);
nand NAND4 (N1015, N1013, N659, N259, N214);
nand NAND2 (N1016, N1014, N757);
nor NOR4 (N1017, N1006, N801, N424, N125);
not NOT1 (N1018, N1010);
or OR2 (N1019, N1012, N1006);
not NOT1 (N1020, N1019);
xor XOR2 (N1021, N1011, N420);
nor NOR2 (N1022, N1021, N211);
xor XOR2 (N1023, N1007, N478);
or OR3 (N1024, N1023, N436, N527);
not NOT1 (N1025, N991);
nand NAND3 (N1026, N1008, N637, N570);
nand NAND4 (N1027, N1026, N735, N902, N483);
and AND2 (N1028, N1027, N1002);
nand NAND3 (N1029, N1016, N198, N1009);
nor NOR4 (N1030, N1015, N538, N592, N848);
xor XOR2 (N1031, N1020, N94);
nand NAND4 (N1032, N1024, N587, N1006, N8);
and AND2 (N1033, N988, N168);
buf BUF1 (N1034, N1030);
or OR4 (N1035, N1017, N447, N779, N285);
and AND3 (N1036, N1031, N15, N56);
not NOT1 (N1037, N1025);
or OR2 (N1038, N1036, N674);
and AND2 (N1039, N1033, N504);
nand NAND4 (N1040, N1028, N139, N996, N918);
nor NOR3 (N1041, N1039, N321, N271);
nor NOR4 (N1042, N1041, N905, N938, N1);
and AND3 (N1043, N1042, N963, N614);
nor NOR4 (N1044, N1040, N496, N235, N331);
buf BUF1 (N1045, N1035);
nor NOR2 (N1046, N1032, N327);
or OR3 (N1047, N1046, N617, N46);
nand NAND3 (N1048, N1022, N510, N739);
or OR4 (N1049, N1029, N288, N979, N854);
not NOT1 (N1050, N1044);
and AND3 (N1051, N1034, N556, N415);
and AND2 (N1052, N1038, N173);
xor XOR2 (N1053, N1043, N521);
nor NOR3 (N1054, N1045, N952, N285);
not NOT1 (N1055, N1018);
nand NAND4 (N1056, N1049, N791, N852, N911);
nand NAND4 (N1057, N1047, N641, N770, N709);
not NOT1 (N1058, N1057);
nand NAND4 (N1059, N1048, N127, N179, N1022);
buf BUF1 (N1060, N1052);
not NOT1 (N1061, N1055);
nand NAND3 (N1062, N1050, N490, N46);
nand NAND4 (N1063, N1056, N560, N601, N916);
or OR3 (N1064, N1062, N876, N760);
and AND3 (N1065, N1060, N992, N1012);
buf BUF1 (N1066, N1064);
or OR3 (N1067, N1037, N77, N1);
nand NAND3 (N1068, N1058, N570, N562);
not NOT1 (N1069, N1065);
xor XOR2 (N1070, N1063, N876);
nand NAND3 (N1071, N1051, N987, N264);
not NOT1 (N1072, N1061);
nor NOR3 (N1073, N1067, N95, N105);
and AND2 (N1074, N1053, N859);
not NOT1 (N1075, N1071);
or OR3 (N1076, N1066, N864, N29);
nor NOR3 (N1077, N1076, N91, N787);
not NOT1 (N1078, N1077);
or OR4 (N1079, N1068, N1004, N34, N997);
buf BUF1 (N1080, N1069);
nand NAND3 (N1081, N1070, N341, N334);
not NOT1 (N1082, N1080);
nor NOR2 (N1083, N1079, N813);
nand NAND3 (N1084, N1078, N980, N662);
buf BUF1 (N1085, N1054);
or OR3 (N1086, N1083, N524, N696);
nand NAND2 (N1087, N1085, N20);
nand NAND2 (N1088, N1059, N938);
nor NOR3 (N1089, N1073, N488, N417);
nor NOR3 (N1090, N1082, N444, N186);
xor XOR2 (N1091, N1089, N647);
and AND4 (N1092, N1088, N851, N456, N566);
and AND2 (N1093, N1091, N603);
not NOT1 (N1094, N1090);
not NOT1 (N1095, N1075);
not NOT1 (N1096, N1084);
buf BUF1 (N1097, N1074);
nand NAND4 (N1098, N1072, N199, N49, N579);
nor NOR3 (N1099, N1087, N236, N661);
and AND4 (N1100, N1097, N248, N467, N758);
buf BUF1 (N1101, N1096);
buf BUF1 (N1102, N1100);
nor NOR4 (N1103, N1094, N631, N815, N796);
nand NAND4 (N1104, N1092, N329, N853, N551);
nand NAND2 (N1105, N1099, N869);
buf BUF1 (N1106, N1086);
and AND4 (N1107, N1101, N670, N267, N377);
buf BUF1 (N1108, N1098);
or OR3 (N1109, N1107, N101, N821);
not NOT1 (N1110, N1104);
xor XOR2 (N1111, N1105, N469);
not NOT1 (N1112, N1081);
buf BUF1 (N1113, N1095);
nor NOR4 (N1114, N1103, N408, N171, N459);
xor XOR2 (N1115, N1106, N582);
xor XOR2 (N1116, N1112, N586);
xor XOR2 (N1117, N1111, N54);
xor XOR2 (N1118, N1109, N733);
nand NAND4 (N1119, N1118, N82, N935, N1001);
or OR4 (N1120, N1119, N425, N19, N272);
buf BUF1 (N1121, N1102);
or OR4 (N1122, N1113, N1092, N160, N335);
and AND3 (N1123, N1114, N436, N1096);
nand NAND3 (N1124, N1110, N934, N779);
or OR3 (N1125, N1123, N141, N915);
or OR3 (N1126, N1124, N11, N479);
not NOT1 (N1127, N1126);
buf BUF1 (N1128, N1120);
not NOT1 (N1129, N1117);
not NOT1 (N1130, N1121);
xor XOR2 (N1131, N1127, N548);
buf BUF1 (N1132, N1116);
xor XOR2 (N1133, N1131, N1102);
nor NOR2 (N1134, N1130, N958);
nand NAND4 (N1135, N1122, N1015, N401, N750);
or OR2 (N1136, N1132, N635);
nand NAND4 (N1137, N1115, N789, N977, N911);
and AND3 (N1138, N1108, N769, N263);
not NOT1 (N1139, N1128);
or OR4 (N1140, N1137, N869, N523, N596);
or OR2 (N1141, N1093, N90);
nor NOR3 (N1142, N1140, N780, N588);
not NOT1 (N1143, N1125);
nand NAND2 (N1144, N1139, N342);
not NOT1 (N1145, N1129);
and AND4 (N1146, N1133, N166, N621, N1024);
not NOT1 (N1147, N1142);
nand NAND3 (N1148, N1144, N734, N159);
buf BUF1 (N1149, N1146);
or OR3 (N1150, N1136, N107, N91);
and AND4 (N1151, N1134, N376, N390, N877);
nor NOR4 (N1152, N1150, N512, N929, N43);
not NOT1 (N1153, N1151);
or OR4 (N1154, N1145, N745, N143, N625);
nor NOR3 (N1155, N1153, N20, N87);
nor NOR4 (N1156, N1135, N478, N1001, N669);
nor NOR4 (N1157, N1154, N869, N199, N323);
or OR4 (N1158, N1147, N529, N481, N187);
xor XOR2 (N1159, N1141, N605);
nor NOR2 (N1160, N1157, N65);
nand NAND3 (N1161, N1160, N1023, N988);
nor NOR2 (N1162, N1152, N170);
or OR2 (N1163, N1158, N290);
xor XOR2 (N1164, N1155, N6);
xor XOR2 (N1165, N1161, N392);
not NOT1 (N1166, N1143);
nand NAND4 (N1167, N1162, N31, N278, N750);
or OR2 (N1168, N1164, N279);
or OR4 (N1169, N1138, N63, N866, N729);
or OR3 (N1170, N1156, N406, N690);
xor XOR2 (N1171, N1166, N466);
nor NOR2 (N1172, N1171, N87);
nor NOR3 (N1173, N1165, N166, N142);
buf BUF1 (N1174, N1168);
nor NOR3 (N1175, N1149, N570, N545);
nor NOR4 (N1176, N1175, N213, N96, N154);
buf BUF1 (N1177, N1170);
and AND4 (N1178, N1167, N469, N126, N222);
nor NOR2 (N1179, N1169, N751);
not NOT1 (N1180, N1176);
xor XOR2 (N1181, N1148, N869);
nor NOR3 (N1182, N1159, N314, N105);
not NOT1 (N1183, N1174);
xor XOR2 (N1184, N1172, N242);
or OR2 (N1185, N1183, N254);
nand NAND2 (N1186, N1163, N343);
nor NOR3 (N1187, N1185, N769, N126);
nand NAND4 (N1188, N1181, N192, N267, N369);
nor NOR4 (N1189, N1173, N69, N597, N497);
nor NOR3 (N1190, N1180, N424, N195);
buf BUF1 (N1191, N1179);
nor NOR3 (N1192, N1190, N1051, N110);
nand NAND4 (N1193, N1192, N1083, N568, N993);
or OR2 (N1194, N1189, N349);
or OR4 (N1195, N1177, N882, N896, N702);
nor NOR2 (N1196, N1187, N150);
nand NAND3 (N1197, N1193, N283, N964);
nor NOR2 (N1198, N1186, N863);
and AND4 (N1199, N1195, N554, N89, N965);
and AND3 (N1200, N1198, N16, N75);
nand NAND2 (N1201, N1178, N429);
not NOT1 (N1202, N1194);
xor XOR2 (N1203, N1188, N473);
buf BUF1 (N1204, N1182);
nand NAND4 (N1205, N1184, N385, N679, N438);
not NOT1 (N1206, N1201);
xor XOR2 (N1207, N1200, N7);
not NOT1 (N1208, N1205);
nor NOR3 (N1209, N1197, N920, N127);
or OR4 (N1210, N1203, N739, N815, N102);
or OR2 (N1211, N1206, N739);
buf BUF1 (N1212, N1191);
not NOT1 (N1213, N1204);
nand NAND3 (N1214, N1210, N738, N606);
not NOT1 (N1215, N1208);
and AND2 (N1216, N1212, N86);
xor XOR2 (N1217, N1207, N811);
or OR2 (N1218, N1209, N671);
nand NAND3 (N1219, N1199, N343, N497);
nor NOR3 (N1220, N1196, N653, N1019);
nand NAND2 (N1221, N1218, N694);
xor XOR2 (N1222, N1220, N109);
and AND4 (N1223, N1215, N721, N1098, N167);
or OR2 (N1224, N1211, N598);
and AND4 (N1225, N1202, N1004, N38, N360);
not NOT1 (N1226, N1221);
xor XOR2 (N1227, N1214, N124);
nor NOR3 (N1228, N1225, N637, N973);
buf BUF1 (N1229, N1224);
and AND2 (N1230, N1228, N532);
not NOT1 (N1231, N1222);
xor XOR2 (N1232, N1230, N1151);
buf BUF1 (N1233, N1217);
buf BUF1 (N1234, N1226);
not NOT1 (N1235, N1231);
or OR2 (N1236, N1234, N472);
and AND4 (N1237, N1235, N291, N992, N453);
buf BUF1 (N1238, N1236);
xor XOR2 (N1239, N1219, N781);
or OR3 (N1240, N1213, N195, N1017);
or OR4 (N1241, N1232, N165, N650, N726);
nand NAND2 (N1242, N1241, N1025);
and AND3 (N1243, N1237, N1100, N611);
or OR3 (N1244, N1229, N1133, N536);
nor NOR3 (N1245, N1238, N637, N1040);
buf BUF1 (N1246, N1227);
and AND4 (N1247, N1239, N496, N516, N1117);
buf BUF1 (N1248, N1242);
xor XOR2 (N1249, N1243, N192);
nor NOR2 (N1250, N1246, N403);
buf BUF1 (N1251, N1233);
not NOT1 (N1252, N1251);
nor NOR4 (N1253, N1247, N780, N754, N933);
or OR2 (N1254, N1250, N744);
not NOT1 (N1255, N1253);
xor XOR2 (N1256, N1254, N748);
and AND4 (N1257, N1240, N205, N987, N479);
not NOT1 (N1258, N1248);
and AND3 (N1259, N1223, N337, N950);
and AND4 (N1260, N1249, N1219, N139, N630);
buf BUF1 (N1261, N1245);
nand NAND4 (N1262, N1259, N495, N541, N707);
not NOT1 (N1263, N1257);
and AND2 (N1264, N1260, N708);
nor NOR3 (N1265, N1216, N1036, N693);
nor NOR2 (N1266, N1263, N741);
nor NOR2 (N1267, N1244, N978);
buf BUF1 (N1268, N1258);
nor NOR2 (N1269, N1252, N674);
nand NAND3 (N1270, N1265, N29, N57);
and AND4 (N1271, N1255, N165, N262, N45);
nand NAND2 (N1272, N1271, N1062);
not NOT1 (N1273, N1272);
not NOT1 (N1274, N1266);
and AND3 (N1275, N1264, N181, N507);
buf BUF1 (N1276, N1275);
buf BUF1 (N1277, N1269);
buf BUF1 (N1278, N1276);
nor NOR2 (N1279, N1268, N742);
nor NOR4 (N1280, N1256, N1160, N1184, N293);
nor NOR2 (N1281, N1267, N1016);
not NOT1 (N1282, N1277);
or OR3 (N1283, N1279, N748, N331);
not NOT1 (N1284, N1281);
buf BUF1 (N1285, N1274);
buf BUF1 (N1286, N1283);
not NOT1 (N1287, N1262);
nor NOR4 (N1288, N1286, N168, N674, N996);
not NOT1 (N1289, N1261);
or OR2 (N1290, N1285, N314);
not NOT1 (N1291, N1289);
nand NAND3 (N1292, N1288, N959, N1233);
not NOT1 (N1293, N1290);
nor NOR3 (N1294, N1287, N124, N168);
nand NAND4 (N1295, N1293, N1268, N438, N126);
xor XOR2 (N1296, N1284, N10);
nand NAND2 (N1297, N1270, N946);
or OR2 (N1298, N1296, N180);
or OR3 (N1299, N1278, N1035, N523);
nand NAND2 (N1300, N1280, N970);
and AND2 (N1301, N1300, N508);
and AND4 (N1302, N1291, N877, N1071, N313);
or OR3 (N1303, N1302, N261, N220);
nor NOR4 (N1304, N1301, N1044, N1031, N269);
nor NOR3 (N1305, N1303, N794, N369);
xor XOR2 (N1306, N1292, N418);
nand NAND2 (N1307, N1282, N682);
and AND3 (N1308, N1307, N1206, N1186);
or OR3 (N1309, N1308, N1237, N159);
buf BUF1 (N1310, N1299);
or OR4 (N1311, N1309, N1002, N936, N421);
xor XOR2 (N1312, N1306, N1002);
nand NAND3 (N1313, N1312, N576, N677);
not NOT1 (N1314, N1313);
xor XOR2 (N1315, N1294, N149);
or OR4 (N1316, N1273, N319, N735, N566);
nand NAND2 (N1317, N1316, N81);
nand NAND3 (N1318, N1305, N297, N303);
xor XOR2 (N1319, N1304, N978);
and AND2 (N1320, N1298, N587);
nor NOR2 (N1321, N1317, N5);
nand NAND4 (N1322, N1319, N645, N126, N879);
or OR3 (N1323, N1297, N219, N1162);
nand NAND4 (N1324, N1320, N590, N346, N234);
nor NOR2 (N1325, N1322, N1030);
or OR4 (N1326, N1310, N851, N676, N736);
or OR3 (N1327, N1324, N471, N193);
buf BUF1 (N1328, N1295);
nor NOR3 (N1329, N1311, N274, N439);
or OR3 (N1330, N1328, N137, N1315);
nor NOR2 (N1331, N762, N421);
buf BUF1 (N1332, N1331);
and AND3 (N1333, N1327, N1117, N748);
xor XOR2 (N1334, N1314, N363);
buf BUF1 (N1335, N1325);
or OR2 (N1336, N1335, N983);
nor NOR4 (N1337, N1323, N1163, N1164, N203);
or OR4 (N1338, N1329, N511, N384, N1295);
buf BUF1 (N1339, N1333);
nor NOR2 (N1340, N1336, N391);
or OR3 (N1341, N1326, N339, N1261);
or OR2 (N1342, N1340, N205);
nor NOR2 (N1343, N1318, N93);
and AND4 (N1344, N1321, N341, N618, N248);
nor NOR2 (N1345, N1338, N449);
nor NOR4 (N1346, N1341, N983, N698, N333);
xor XOR2 (N1347, N1334, N526);
not NOT1 (N1348, N1345);
or OR3 (N1349, N1347, N325, N421);
and AND4 (N1350, N1342, N8, N913, N1188);
buf BUF1 (N1351, N1349);
and AND3 (N1352, N1346, N790, N658);
xor XOR2 (N1353, N1343, N40);
not NOT1 (N1354, N1352);
nor NOR4 (N1355, N1350, N416, N426, N877);
buf BUF1 (N1356, N1339);
buf BUF1 (N1357, N1332);
nor NOR3 (N1358, N1356, N744, N90);
nand NAND3 (N1359, N1353, N824, N195);
nand NAND4 (N1360, N1359, N495, N1011, N171);
or OR3 (N1361, N1355, N882, N507);
and AND3 (N1362, N1351, N1041, N144);
not NOT1 (N1363, N1358);
xor XOR2 (N1364, N1348, N278);
not NOT1 (N1365, N1344);
not NOT1 (N1366, N1361);
not NOT1 (N1367, N1362);
not NOT1 (N1368, N1357);
nand NAND2 (N1369, N1364, N1032);
nand NAND3 (N1370, N1365, N290, N906);
or OR2 (N1371, N1368, N1134);
not NOT1 (N1372, N1370);
or OR3 (N1373, N1372, N398, N1184);
and AND3 (N1374, N1354, N655, N172);
not NOT1 (N1375, N1373);
xor XOR2 (N1376, N1369, N287);
or OR3 (N1377, N1330, N538, N1368);
nor NOR2 (N1378, N1366, N1102);
xor XOR2 (N1379, N1374, N271);
not NOT1 (N1380, N1367);
not NOT1 (N1381, N1377);
buf BUF1 (N1382, N1376);
not NOT1 (N1383, N1360);
nor NOR4 (N1384, N1382, N546, N864, N1189);
xor XOR2 (N1385, N1379, N748);
xor XOR2 (N1386, N1378, N806);
nor NOR2 (N1387, N1380, N405);
or OR2 (N1388, N1387, N1076);
not NOT1 (N1389, N1388);
and AND3 (N1390, N1381, N1316, N354);
nor NOR3 (N1391, N1337, N501, N904);
and AND4 (N1392, N1383, N1151, N1257, N1194);
not NOT1 (N1393, N1386);
or OR4 (N1394, N1393, N489, N230, N1361);
or OR4 (N1395, N1392, N82, N643, N461);
or OR2 (N1396, N1391, N1127);
not NOT1 (N1397, N1385);
not NOT1 (N1398, N1375);
xor XOR2 (N1399, N1371, N1099);
not NOT1 (N1400, N1363);
or OR4 (N1401, N1394, N872, N1064, N28);
buf BUF1 (N1402, N1397);
not NOT1 (N1403, N1390);
buf BUF1 (N1404, N1400);
buf BUF1 (N1405, N1398);
or OR4 (N1406, N1402, N700, N828, N978);
and AND2 (N1407, N1405, N599);
xor XOR2 (N1408, N1395, N196);
or OR4 (N1409, N1404, N847, N1341, N1116);
nand NAND4 (N1410, N1401, N499, N474, N1209);
buf BUF1 (N1411, N1389);
nand NAND3 (N1412, N1408, N697, N1365);
nor NOR3 (N1413, N1406, N954, N63);
buf BUF1 (N1414, N1384);
nor NOR2 (N1415, N1399, N75);
and AND4 (N1416, N1411, N1268, N1380, N345);
or OR4 (N1417, N1410, N851, N648, N212);
or OR2 (N1418, N1412, N424);
not NOT1 (N1419, N1416);
buf BUF1 (N1420, N1415);
not NOT1 (N1421, N1407);
nand NAND4 (N1422, N1421, N1134, N658, N1257);
nor NOR4 (N1423, N1422, N428, N146, N988);
not NOT1 (N1424, N1409);
buf BUF1 (N1425, N1419);
not NOT1 (N1426, N1418);
or OR2 (N1427, N1423, N952);
nand NAND3 (N1428, N1413, N81, N1266);
nand NAND4 (N1429, N1417, N1189, N595, N96);
xor XOR2 (N1430, N1414, N824);
buf BUF1 (N1431, N1427);
buf BUF1 (N1432, N1426);
or OR2 (N1433, N1425, N303);
buf BUF1 (N1434, N1433);
not NOT1 (N1435, N1420);
buf BUF1 (N1436, N1428);
and AND2 (N1437, N1430, N1135);
and AND4 (N1438, N1424, N567, N47, N679);
and AND4 (N1439, N1431, N1359, N748, N1116);
nor NOR4 (N1440, N1436, N861, N170, N867);
nand NAND3 (N1441, N1403, N40, N213);
and AND3 (N1442, N1437, N1285, N775);
nor NOR4 (N1443, N1438, N1422, N1212, N110);
or OR4 (N1444, N1429, N1427, N1222, N197);
nand NAND3 (N1445, N1443, N691, N776);
nand NAND2 (N1446, N1434, N67);
xor XOR2 (N1447, N1446, N241);
buf BUF1 (N1448, N1396);
buf BUF1 (N1449, N1432);
or OR3 (N1450, N1442, N820, N1395);
xor XOR2 (N1451, N1439, N241);
xor XOR2 (N1452, N1447, N145);
or OR4 (N1453, N1449, N461, N1305, N248);
nand NAND3 (N1454, N1451, N1221, N216);
or OR4 (N1455, N1453, N19, N43, N915);
nor NOR3 (N1456, N1441, N621, N475);
and AND2 (N1457, N1452, N391);
or OR4 (N1458, N1454, N1006, N412, N875);
nand NAND3 (N1459, N1444, N455, N891);
nor NOR2 (N1460, N1456, N574);
buf BUF1 (N1461, N1450);
xor XOR2 (N1462, N1461, N841);
and AND3 (N1463, N1448, N442, N86);
xor XOR2 (N1464, N1458, N1050);
buf BUF1 (N1465, N1455);
nor NOR4 (N1466, N1440, N1339, N657, N868);
xor XOR2 (N1467, N1463, N1132);
nor NOR3 (N1468, N1462, N961, N200);
and AND3 (N1469, N1435, N1297, N349);
nand NAND2 (N1470, N1457, N201);
xor XOR2 (N1471, N1469, N810);
and AND3 (N1472, N1470, N599, N911);
not NOT1 (N1473, N1459);
nor NOR2 (N1474, N1467, N707);
or OR2 (N1475, N1471, N1414);
xor XOR2 (N1476, N1472, N1048);
and AND4 (N1477, N1464, N1229, N1196, N446);
nand NAND3 (N1478, N1476, N78, N817);
buf BUF1 (N1479, N1466);
buf BUF1 (N1480, N1468);
nor NOR4 (N1481, N1465, N1426, N637, N940);
and AND3 (N1482, N1474, N165, N1319);
xor XOR2 (N1483, N1481, N1233);
not NOT1 (N1484, N1479);
and AND2 (N1485, N1473, N505);
or OR4 (N1486, N1475, N1235, N237, N1473);
nor NOR2 (N1487, N1460, N1060);
and AND3 (N1488, N1486, N718, N20);
and AND4 (N1489, N1484, N595, N390, N1217);
xor XOR2 (N1490, N1445, N530);
nand NAND4 (N1491, N1485, N1078, N966, N379);
xor XOR2 (N1492, N1490, N213);
or OR4 (N1493, N1480, N1310, N101, N497);
or OR2 (N1494, N1493, N358);
or OR3 (N1495, N1487, N1206, N236);
or OR4 (N1496, N1492, N949, N796, N703);
xor XOR2 (N1497, N1496, N1299);
and AND3 (N1498, N1495, N17, N1390);
nor NOR3 (N1499, N1497, N847, N225);
nand NAND4 (N1500, N1483, N42, N194, N371);
xor XOR2 (N1501, N1498, N515);
buf BUF1 (N1502, N1478);
xor XOR2 (N1503, N1502, N452);
nor NOR4 (N1504, N1501, N1218, N776, N260);
buf BUF1 (N1505, N1489);
not NOT1 (N1506, N1488);
and AND3 (N1507, N1500, N1343, N706);
xor XOR2 (N1508, N1503, N1106);
xor XOR2 (N1509, N1499, N755);
and AND2 (N1510, N1506, N757);
buf BUF1 (N1511, N1504);
or OR4 (N1512, N1509, N636, N465, N638);
nand NAND4 (N1513, N1491, N707, N1059, N530);
xor XOR2 (N1514, N1477, N718);
xor XOR2 (N1515, N1513, N1344);
not NOT1 (N1516, N1512);
nand NAND4 (N1517, N1505, N479, N1204, N932);
or OR3 (N1518, N1494, N380, N1141);
xor XOR2 (N1519, N1507, N636);
not NOT1 (N1520, N1510);
not NOT1 (N1521, N1516);
nand NAND3 (N1522, N1519, N782, N29);
or OR2 (N1523, N1520, N739);
and AND2 (N1524, N1517, N434);
xor XOR2 (N1525, N1508, N1152);
buf BUF1 (N1526, N1524);
nand NAND4 (N1527, N1522, N776, N1343, N342);
nand NAND2 (N1528, N1514, N675);
buf BUF1 (N1529, N1528);
xor XOR2 (N1530, N1527, N122);
and AND4 (N1531, N1515, N1087, N1180, N485);
or OR3 (N1532, N1518, N793, N650);
and AND3 (N1533, N1529, N1228, N289);
or OR3 (N1534, N1530, N703, N816);
and AND3 (N1535, N1523, N443, N689);
or OR3 (N1536, N1521, N1010, N334);
nand NAND2 (N1537, N1526, N404);
or OR4 (N1538, N1531, N1404, N1245, N1449);
nor NOR2 (N1539, N1537, N1455);
buf BUF1 (N1540, N1538);
xor XOR2 (N1541, N1535, N553);
or OR2 (N1542, N1511, N1081);
not NOT1 (N1543, N1525);
not NOT1 (N1544, N1542);
xor XOR2 (N1545, N1482, N1132);
xor XOR2 (N1546, N1543, N1262);
xor XOR2 (N1547, N1533, N1170);
nor NOR4 (N1548, N1534, N63, N1406, N164);
and AND3 (N1549, N1540, N1364, N280);
buf BUF1 (N1550, N1547);
buf BUF1 (N1551, N1545);
buf BUF1 (N1552, N1546);
not NOT1 (N1553, N1548);
or OR2 (N1554, N1536, N593);
nand NAND3 (N1555, N1539, N1311, N99);
or OR2 (N1556, N1553, N328);
and AND4 (N1557, N1556, N13, N443, N101);
xor XOR2 (N1558, N1532, N900);
nand NAND4 (N1559, N1551, N1391, N1428, N513);
nor NOR3 (N1560, N1550, N45, N545);
nor NOR2 (N1561, N1554, N43);
not NOT1 (N1562, N1549);
nor NOR3 (N1563, N1541, N1091, N1108);
buf BUF1 (N1564, N1544);
buf BUF1 (N1565, N1559);
nor NOR4 (N1566, N1552, N1362, N231, N1167);
or OR2 (N1567, N1558, N1183);
buf BUF1 (N1568, N1555);
or OR3 (N1569, N1567, N1213, N667);
xor XOR2 (N1570, N1568, N643);
nand NAND4 (N1571, N1566, N375, N435, N968);
xor XOR2 (N1572, N1564, N1021);
and AND2 (N1573, N1570, N1404);
buf BUF1 (N1574, N1563);
nand NAND4 (N1575, N1560, N608, N336, N1125);
and AND4 (N1576, N1561, N1263, N680, N178);
not NOT1 (N1577, N1575);
xor XOR2 (N1578, N1574, N396);
xor XOR2 (N1579, N1577, N340);
buf BUF1 (N1580, N1557);
nand NAND4 (N1581, N1572, N808, N1007, N212);
xor XOR2 (N1582, N1578, N1085);
and AND4 (N1583, N1573, N1093, N1069, N453);
and AND4 (N1584, N1582, N616, N1381, N1485);
not NOT1 (N1585, N1584);
nor NOR3 (N1586, N1576, N780, N1266);
not NOT1 (N1587, N1562);
xor XOR2 (N1588, N1581, N1205);
not NOT1 (N1589, N1588);
or OR2 (N1590, N1569, N732);
xor XOR2 (N1591, N1590, N1424);
or OR3 (N1592, N1580, N1207, N858);
not NOT1 (N1593, N1591);
and AND3 (N1594, N1583, N59, N782);
nor NOR2 (N1595, N1592, N843);
nor NOR2 (N1596, N1593, N939);
buf BUF1 (N1597, N1579);
nor NOR2 (N1598, N1594, N1232);
nand NAND3 (N1599, N1586, N259, N417);
or OR2 (N1600, N1598, N1391);
nand NAND2 (N1601, N1571, N119);
nand NAND3 (N1602, N1600, N1032, N454);
or OR2 (N1603, N1596, N1111);
not NOT1 (N1604, N1587);
buf BUF1 (N1605, N1601);
nand NAND2 (N1606, N1604, N1067);
nor NOR4 (N1607, N1585, N271, N182, N938);
not NOT1 (N1608, N1599);
not NOT1 (N1609, N1606);
buf BUF1 (N1610, N1609);
and AND4 (N1611, N1602, N1585, N954, N989);
not NOT1 (N1612, N1603);
xor XOR2 (N1613, N1608, N879);
xor XOR2 (N1614, N1607, N1544);
nand NAND3 (N1615, N1614, N371, N1392);
xor XOR2 (N1616, N1612, N255);
or OR4 (N1617, N1611, N830, N1216, N1427);
buf BUF1 (N1618, N1617);
buf BUF1 (N1619, N1618);
buf BUF1 (N1620, N1595);
xor XOR2 (N1621, N1619, N1553);
or OR3 (N1622, N1589, N1317, N556);
and AND2 (N1623, N1622, N665);
xor XOR2 (N1624, N1615, N1335);
not NOT1 (N1625, N1610);
or OR2 (N1626, N1625, N1078);
buf BUF1 (N1627, N1623);
buf BUF1 (N1628, N1620);
not NOT1 (N1629, N1621);
not NOT1 (N1630, N1629);
or OR2 (N1631, N1624, N186);
buf BUF1 (N1632, N1565);
or OR2 (N1633, N1613, N154);
buf BUF1 (N1634, N1597);
xor XOR2 (N1635, N1632, N249);
not NOT1 (N1636, N1630);
or OR3 (N1637, N1635, N867, N1568);
nand NAND2 (N1638, N1633, N40);
not NOT1 (N1639, N1638);
not NOT1 (N1640, N1631);
buf BUF1 (N1641, N1640);
nor NOR3 (N1642, N1637, N1584, N758);
not NOT1 (N1643, N1626);
xor XOR2 (N1644, N1628, N897);
or OR2 (N1645, N1634, N132);
xor XOR2 (N1646, N1641, N340);
or OR4 (N1647, N1646, N1628, N1389, N1558);
and AND4 (N1648, N1605, N816, N1, N283);
nand NAND2 (N1649, N1636, N1116);
or OR2 (N1650, N1642, N1556);
nand NAND3 (N1651, N1645, N984, N338);
buf BUF1 (N1652, N1616);
xor XOR2 (N1653, N1650, N568);
xor XOR2 (N1654, N1643, N1113);
nand NAND2 (N1655, N1639, N1482);
and AND4 (N1656, N1649, N688, N1120, N444);
and AND2 (N1657, N1654, N1431);
xor XOR2 (N1658, N1657, N210);
not NOT1 (N1659, N1648);
buf BUF1 (N1660, N1644);
buf BUF1 (N1661, N1647);
xor XOR2 (N1662, N1661, N1329);
and AND2 (N1663, N1627, N723);
nor NOR4 (N1664, N1653, N1345, N840, N717);
nand NAND2 (N1665, N1652, N720);
and AND3 (N1666, N1655, N190, N613);
or OR4 (N1667, N1651, N1640, N593, N1021);
nand NAND2 (N1668, N1659, N210);
and AND2 (N1669, N1662, N1572);
nor NOR4 (N1670, N1667, N1506, N268, N1301);
not NOT1 (N1671, N1668);
or OR2 (N1672, N1660, N1473);
not NOT1 (N1673, N1666);
buf BUF1 (N1674, N1669);
or OR3 (N1675, N1658, N1184, N884);
buf BUF1 (N1676, N1671);
not NOT1 (N1677, N1665);
and AND2 (N1678, N1656, N1421);
xor XOR2 (N1679, N1675, N743);
xor XOR2 (N1680, N1672, N326);
or OR3 (N1681, N1676, N960, N1464);
nand NAND2 (N1682, N1673, N854);
buf BUF1 (N1683, N1678);
nor NOR4 (N1684, N1682, N437, N682, N45);
xor XOR2 (N1685, N1679, N288);
buf BUF1 (N1686, N1685);
not NOT1 (N1687, N1681);
buf BUF1 (N1688, N1674);
xor XOR2 (N1689, N1688, N567);
and AND3 (N1690, N1677, N407, N1004);
xor XOR2 (N1691, N1670, N709);
buf BUF1 (N1692, N1690);
or OR3 (N1693, N1663, N1114, N994);
xor XOR2 (N1694, N1687, N258);
or OR4 (N1695, N1693, N106, N1297, N1213);
or OR3 (N1696, N1691, N52, N1597);
or OR2 (N1697, N1683, N983);
nor NOR2 (N1698, N1692, N568);
nor NOR3 (N1699, N1696, N1054, N1142);
xor XOR2 (N1700, N1664, N1645);
not NOT1 (N1701, N1686);
buf BUF1 (N1702, N1701);
xor XOR2 (N1703, N1695, N110);
and AND3 (N1704, N1700, N367, N619);
buf BUF1 (N1705, N1697);
or OR2 (N1706, N1694, N1339);
nor NOR3 (N1707, N1705, N186, N636);
nand NAND3 (N1708, N1699, N811, N705);
or OR4 (N1709, N1708, N694, N864, N691);
and AND3 (N1710, N1706, N752, N1650);
or OR2 (N1711, N1710, N639);
buf BUF1 (N1712, N1698);
xor XOR2 (N1713, N1712, N1105);
xor XOR2 (N1714, N1684, N1175);
not NOT1 (N1715, N1680);
nor NOR2 (N1716, N1702, N1173);
nor NOR3 (N1717, N1716, N1535, N1545);
not NOT1 (N1718, N1715);
nor NOR3 (N1719, N1704, N241, N1206);
and AND4 (N1720, N1709, N431, N1699, N1066);
and AND4 (N1721, N1713, N88, N356, N544);
nor NOR3 (N1722, N1689, N1592, N1701);
xor XOR2 (N1723, N1703, N997);
nor NOR3 (N1724, N1723, N667, N1074);
xor XOR2 (N1725, N1720, N1451);
nor NOR4 (N1726, N1724, N758, N913, N1000);
and AND4 (N1727, N1714, N738, N50, N917);
xor XOR2 (N1728, N1707, N1138);
or OR2 (N1729, N1728, N1154);
nor NOR2 (N1730, N1719, N543);
nand NAND4 (N1731, N1722, N1624, N901, N733);
nand NAND2 (N1732, N1718, N374);
xor XOR2 (N1733, N1732, N688);
nor NOR2 (N1734, N1731, N1140);
nor NOR2 (N1735, N1734, N176);
buf BUF1 (N1736, N1711);
buf BUF1 (N1737, N1725);
nor NOR4 (N1738, N1733, N1004, N170, N629);
not NOT1 (N1739, N1730);
nand NAND4 (N1740, N1726, N1195, N898, N1307);
or OR4 (N1741, N1740, N249, N1671, N26);
and AND4 (N1742, N1739, N601, N1589, N254);
and AND3 (N1743, N1738, N755, N424);
not NOT1 (N1744, N1735);
or OR4 (N1745, N1727, N1445, N1292, N740);
and AND4 (N1746, N1717, N771, N308, N796);
not NOT1 (N1747, N1744);
not NOT1 (N1748, N1743);
and AND4 (N1749, N1746, N328, N1692, N925);
not NOT1 (N1750, N1741);
or OR4 (N1751, N1745, N1038, N1550, N964);
and AND3 (N1752, N1750, N1454, N228);
or OR2 (N1753, N1752, N240);
not NOT1 (N1754, N1736);
not NOT1 (N1755, N1747);
and AND2 (N1756, N1729, N1044);
or OR2 (N1757, N1754, N1663);
or OR3 (N1758, N1756, N991, N134);
or OR4 (N1759, N1753, N796, N607, N445);
not NOT1 (N1760, N1759);
nand NAND4 (N1761, N1748, N53, N1248, N11);
and AND4 (N1762, N1721, N1604, N973, N1013);
and AND3 (N1763, N1761, N842, N15);
nor NOR2 (N1764, N1755, N905);
not NOT1 (N1765, N1760);
not NOT1 (N1766, N1762);
or OR3 (N1767, N1757, N1290, N1161);
nand NAND4 (N1768, N1767, N239, N1391, N499);
nor NOR2 (N1769, N1749, N1181);
xor XOR2 (N1770, N1765, N134);
not NOT1 (N1771, N1768);
xor XOR2 (N1772, N1770, N167);
buf BUF1 (N1773, N1758);
xor XOR2 (N1774, N1763, N1057);
buf BUF1 (N1775, N1764);
and AND3 (N1776, N1774, N1289, N535);
nor NOR3 (N1777, N1742, N816, N980);
nor NOR4 (N1778, N1766, N1179, N606, N662);
not NOT1 (N1779, N1775);
nand NAND2 (N1780, N1777, N1525);
or OR3 (N1781, N1771, N540, N839);
or OR2 (N1782, N1779, N927);
nand NAND3 (N1783, N1737, N901, N372);
buf BUF1 (N1784, N1780);
buf BUF1 (N1785, N1778);
not NOT1 (N1786, N1769);
nor NOR3 (N1787, N1783, N107, N1528);
nor NOR3 (N1788, N1784, N1163, N69);
buf BUF1 (N1789, N1776);
nand NAND3 (N1790, N1781, N1667, N1653);
or OR4 (N1791, N1786, N923, N1667, N1377);
buf BUF1 (N1792, N1788);
xor XOR2 (N1793, N1792, N257);
xor XOR2 (N1794, N1793, N608);
xor XOR2 (N1795, N1791, N296);
not NOT1 (N1796, N1785);
xor XOR2 (N1797, N1790, N380);
buf BUF1 (N1798, N1797);
or OR4 (N1799, N1789, N1750, N943, N1728);
or OR4 (N1800, N1799, N1578, N1225, N1535);
or OR4 (N1801, N1782, N631, N1162, N1133);
buf BUF1 (N1802, N1751);
nor NOR2 (N1803, N1795, N1072);
nand NAND4 (N1804, N1794, N394, N75, N865);
nor NOR4 (N1805, N1803, N92, N971, N1576);
not NOT1 (N1806, N1800);
xor XOR2 (N1807, N1773, N1678);
or OR3 (N1808, N1807, N109, N1391);
or OR3 (N1809, N1798, N262, N1066);
and AND3 (N1810, N1808, N1718, N1199);
nor NOR4 (N1811, N1809, N284, N91, N1650);
nand NAND2 (N1812, N1810, N854);
nor NOR2 (N1813, N1806, N976);
not NOT1 (N1814, N1801);
and AND2 (N1815, N1804, N820);
nor NOR3 (N1816, N1772, N300, N1291);
not NOT1 (N1817, N1787);
and AND2 (N1818, N1811, N156);
nand NAND2 (N1819, N1815, N123);
nand NAND2 (N1820, N1817, N450);
nor NOR2 (N1821, N1814, N1550);
xor XOR2 (N1822, N1805, N720);
not NOT1 (N1823, N1819);
and AND2 (N1824, N1813, N164);
buf BUF1 (N1825, N1818);
buf BUF1 (N1826, N1822);
nand NAND4 (N1827, N1826, N1331, N308, N997);
or OR4 (N1828, N1820, N1304, N474, N1627);
buf BUF1 (N1829, N1802);
not NOT1 (N1830, N1824);
and AND3 (N1831, N1796, N605, N559);
xor XOR2 (N1832, N1825, N325);
buf BUF1 (N1833, N1812);
nand NAND3 (N1834, N1827, N1449, N1415);
nor NOR3 (N1835, N1834, N687, N51);
nand NAND2 (N1836, N1821, N355);
xor XOR2 (N1837, N1829, N779);
and AND2 (N1838, N1836, N303);
xor XOR2 (N1839, N1816, N749);
nand NAND4 (N1840, N1839, N1727, N1478, N640);
not NOT1 (N1841, N1837);
buf BUF1 (N1842, N1835);
or OR3 (N1843, N1842, N1396, N1680);
or OR2 (N1844, N1833, N662);
and AND4 (N1845, N1843, N1645, N1598, N733);
or OR4 (N1846, N1823, N417, N414, N698);
xor XOR2 (N1847, N1846, N96);
not NOT1 (N1848, N1840);
buf BUF1 (N1849, N1832);
buf BUF1 (N1850, N1848);
or OR4 (N1851, N1847, N1569, N1672, N5);
nand NAND2 (N1852, N1831, N1479);
and AND2 (N1853, N1828, N39);
or OR4 (N1854, N1845, N1178, N1364, N1711);
xor XOR2 (N1855, N1853, N1571);
nand NAND4 (N1856, N1830, N1766, N24, N924);
xor XOR2 (N1857, N1854, N1314);
or OR2 (N1858, N1852, N1836);
nor NOR2 (N1859, N1838, N817);
nor NOR3 (N1860, N1859, N100, N583);
nor NOR4 (N1861, N1844, N262, N883, N474);
and AND4 (N1862, N1855, N1458, N1094, N744);
xor XOR2 (N1863, N1849, N1593);
xor XOR2 (N1864, N1858, N480);
and AND3 (N1865, N1860, N846, N1575);
and AND3 (N1866, N1865, N1746, N1661);
and AND2 (N1867, N1866, N1773);
nand NAND3 (N1868, N1856, N927, N16);
nor NOR2 (N1869, N1868, N1808);
not NOT1 (N1870, N1851);
xor XOR2 (N1871, N1870, N1645);
nand NAND2 (N1872, N1864, N1259);
or OR3 (N1873, N1862, N1482, N729);
nand NAND3 (N1874, N1841, N1685, N1361);
xor XOR2 (N1875, N1874, N528);
nand NAND4 (N1876, N1875, N715, N1779, N1772);
or OR2 (N1877, N1871, N502);
not NOT1 (N1878, N1850);
and AND4 (N1879, N1872, N637, N494, N973);
not NOT1 (N1880, N1869);
nand NAND3 (N1881, N1863, N54, N771);
or OR3 (N1882, N1876, N696, N138);
buf BUF1 (N1883, N1877);
xor XOR2 (N1884, N1867, N1175);
or OR4 (N1885, N1873, N1039, N904, N79);
not NOT1 (N1886, N1879);
buf BUF1 (N1887, N1881);
and AND2 (N1888, N1878, N470);
xor XOR2 (N1889, N1882, N1216);
nand NAND3 (N1890, N1884, N972, N331);
xor XOR2 (N1891, N1883, N174);
nand NAND3 (N1892, N1857, N1437, N1080);
and AND4 (N1893, N1890, N559, N1885, N1663);
xor XOR2 (N1894, N472, N473);
nand NAND2 (N1895, N1891, N725);
nor NOR3 (N1896, N1894, N1852, N1055);
and AND3 (N1897, N1893, N1334, N102);
buf BUF1 (N1898, N1861);
buf BUF1 (N1899, N1892);
xor XOR2 (N1900, N1897, N523);
buf BUF1 (N1901, N1896);
not NOT1 (N1902, N1880);
and AND4 (N1903, N1898, N1466, N924, N4);
and AND4 (N1904, N1886, N966, N984, N1759);
xor XOR2 (N1905, N1901, N1567);
buf BUF1 (N1906, N1900);
buf BUF1 (N1907, N1906);
nand NAND2 (N1908, N1887, N1069);
xor XOR2 (N1909, N1895, N431);
buf BUF1 (N1910, N1889);
nor NOR2 (N1911, N1907, N82);
nor NOR2 (N1912, N1911, N1653);
xor XOR2 (N1913, N1904, N1579);
and AND4 (N1914, N1888, N126, N32, N1773);
nand NAND2 (N1915, N1913, N1486);
xor XOR2 (N1916, N1899, N830);
xor XOR2 (N1917, N1909, N1897);
nor NOR4 (N1918, N1910, N1282, N1279, N687);
buf BUF1 (N1919, N1916);
buf BUF1 (N1920, N1905);
nand NAND4 (N1921, N1902, N1058, N422, N1908);
buf BUF1 (N1922, N1017);
and AND4 (N1923, N1918, N961, N811, N1357);
not NOT1 (N1924, N1921);
buf BUF1 (N1925, N1912);
or OR4 (N1926, N1914, N370, N538, N659);
and AND3 (N1927, N1920, N136, N824);
nand NAND2 (N1928, N1922, N37);
nand NAND3 (N1929, N1925, N1538, N244);
or OR2 (N1930, N1903, N383);
and AND2 (N1931, N1924, N554);
xor XOR2 (N1932, N1926, N1765);
xor XOR2 (N1933, N1932, N886);
buf BUF1 (N1934, N1933);
nand NAND4 (N1935, N1923, N505, N640, N1225);
nor NOR4 (N1936, N1935, N423, N1907, N30);
and AND2 (N1937, N1915, N1380);
xor XOR2 (N1938, N1929, N293);
nand NAND3 (N1939, N1938, N1372, N1210);
not NOT1 (N1940, N1934);
not NOT1 (N1941, N1917);
or OR3 (N1942, N1936, N1070, N319);
xor XOR2 (N1943, N1942, N889);
not NOT1 (N1944, N1919);
nor NOR3 (N1945, N1931, N420, N1299);
nor NOR3 (N1946, N1944, N1739, N1496);
nor NOR2 (N1947, N1930, N1595);
or OR3 (N1948, N1945, N1343, N1885);
not NOT1 (N1949, N1927);
not NOT1 (N1950, N1940);
not NOT1 (N1951, N1948);
and AND4 (N1952, N1939, N1627, N1393, N1618);
nor NOR4 (N1953, N1928, N734, N232, N1145);
xor XOR2 (N1954, N1937, N1335);
not NOT1 (N1955, N1950);
nand NAND2 (N1956, N1946, N1410);
not NOT1 (N1957, N1949);
buf BUF1 (N1958, N1947);
nand NAND4 (N1959, N1953, N1618, N857, N1249);
buf BUF1 (N1960, N1958);
xor XOR2 (N1961, N1952, N641);
xor XOR2 (N1962, N1943, N46);
xor XOR2 (N1963, N1959, N1003);
or OR3 (N1964, N1957, N1311, N1110);
nor NOR3 (N1965, N1941, N1900, N1677);
nand NAND3 (N1966, N1961, N504, N1758);
nor NOR4 (N1967, N1960, N1672, N821, N1939);
not NOT1 (N1968, N1964);
or OR3 (N1969, N1951, N468, N481);
not NOT1 (N1970, N1955);
nor NOR3 (N1971, N1968, N1165, N1441);
xor XOR2 (N1972, N1967, N1172);
buf BUF1 (N1973, N1956);
or OR4 (N1974, N1963, N1100, N1755, N1531);
not NOT1 (N1975, N1973);
xor XOR2 (N1976, N1974, N1417);
xor XOR2 (N1977, N1965, N1922);
xor XOR2 (N1978, N1972, N1129);
buf BUF1 (N1979, N1969);
nand NAND3 (N1980, N1970, N1317, N1075);
nor NOR2 (N1981, N1976, N320);
and AND4 (N1982, N1954, N1625, N952, N745);
or OR3 (N1983, N1982, N1390, N84);
and AND4 (N1984, N1981, N873, N394, N58);
xor XOR2 (N1985, N1984, N1581);
buf BUF1 (N1986, N1985);
nand NAND4 (N1987, N1975, N524, N1980, N641);
or OR4 (N1988, N1939, N1366, N597, N1692);
or OR3 (N1989, N1987, N1919, N1179);
nand NAND3 (N1990, N1962, N539, N1119);
xor XOR2 (N1991, N1983, N29);
and AND3 (N1992, N1966, N1331, N652);
and AND4 (N1993, N1986, N837, N611, N403);
nor NOR2 (N1994, N1993, N1074);
nand NAND4 (N1995, N1977, N1540, N725, N707);
and AND2 (N1996, N1971, N645);
nand NAND2 (N1997, N1990, N944);
and AND3 (N1998, N1978, N931, N232);
not NOT1 (N1999, N1997);
and AND3 (N2000, N1994, N42, N762);
or OR3 (N2001, N1988, N1723, N499);
not NOT1 (N2002, N1998);
xor XOR2 (N2003, N2002, N1553);
xor XOR2 (N2004, N2000, N1393);
and AND3 (N2005, N2003, N1907, N1530);
xor XOR2 (N2006, N1979, N503);
xor XOR2 (N2007, N2005, N284);
or OR2 (N2008, N2004, N343);
nand NAND4 (N2009, N2006, N339, N246, N12);
buf BUF1 (N2010, N1999);
nand NAND3 (N2011, N1992, N1662, N891);
xor XOR2 (N2012, N2001, N1434);
nor NOR3 (N2013, N1991, N1902, N1901);
and AND2 (N2014, N1996, N1601);
nand NAND4 (N2015, N2011, N10, N1508, N1211);
not NOT1 (N2016, N1995);
nand NAND3 (N2017, N2008, N1657, N202);
xor XOR2 (N2018, N2012, N532);
or OR2 (N2019, N2009, N1739);
nor NOR3 (N2020, N2015, N285, N221);
xor XOR2 (N2021, N2013, N1339);
not NOT1 (N2022, N2007);
buf BUF1 (N2023, N2019);
buf BUF1 (N2024, N2014);
and AND2 (N2025, N2024, N454);
not NOT1 (N2026, N2020);
or OR2 (N2027, N2026, N166);
not NOT1 (N2028, N2027);
not NOT1 (N2029, N2022);
nor NOR3 (N2030, N1989, N1996, N762);
nor NOR3 (N2031, N2016, N938, N1836);
buf BUF1 (N2032, N2023);
nand NAND2 (N2033, N2032, N170);
buf BUF1 (N2034, N2010);
and AND2 (N2035, N2017, N1435);
nor NOR4 (N2036, N2031, N110, N1768, N1996);
or OR4 (N2037, N2036, N784, N911, N755);
not NOT1 (N2038, N2018);
not NOT1 (N2039, N2025);
not NOT1 (N2040, N2034);
xor XOR2 (N2041, N2030, N1768);
nand NAND4 (N2042, N2029, N1137, N1056, N1835);
nand NAND2 (N2043, N2041, N1809);
nor NOR4 (N2044, N2039, N2011, N1222, N1525);
and AND3 (N2045, N2033, N363, N1897);
xor XOR2 (N2046, N2028, N1350);
nor NOR4 (N2047, N2043, N330, N747, N941);
xor XOR2 (N2048, N2035, N274);
or OR2 (N2049, N2046, N113);
and AND4 (N2050, N2047, N1244, N1254, N371);
not NOT1 (N2051, N2049);
buf BUF1 (N2052, N2048);
and AND2 (N2053, N2052, N189);
not NOT1 (N2054, N2050);
or OR4 (N2055, N2038, N84, N1815, N147);
xor XOR2 (N2056, N2053, N1648);
xor XOR2 (N2057, N2051, N177);
xor XOR2 (N2058, N2021, N1387);
buf BUF1 (N2059, N2057);
xor XOR2 (N2060, N2055, N331);
not NOT1 (N2061, N2060);
not NOT1 (N2062, N2059);
nor NOR2 (N2063, N2054, N144);
and AND2 (N2064, N2037, N1614);
and AND3 (N2065, N2042, N422, N367);
nor NOR3 (N2066, N2062, N284, N1044);
not NOT1 (N2067, N2064);
nor NOR4 (N2068, N2045, N89, N904, N1341);
buf BUF1 (N2069, N2063);
nand NAND4 (N2070, N2056, N22, N1060, N415);
and AND4 (N2071, N2069, N687, N1700, N56);
nor NOR3 (N2072, N2044, N1354, N293);
buf BUF1 (N2073, N2067);
not NOT1 (N2074, N2061);
not NOT1 (N2075, N2071);
buf BUF1 (N2076, N2040);
nor NOR2 (N2077, N2074, N1651);
and AND2 (N2078, N2068, N1437);
xor XOR2 (N2079, N2058, N475);
not NOT1 (N2080, N2070);
and AND4 (N2081, N2073, N1739, N372, N1889);
not NOT1 (N2082, N2078);
nor NOR3 (N2083, N2075, N1322, N1266);
nor NOR4 (N2084, N2065, N1412, N1148, N864);
xor XOR2 (N2085, N2072, N1520);
or OR2 (N2086, N2081, N1815);
or OR3 (N2087, N2077, N842, N530);
not NOT1 (N2088, N2087);
or OR4 (N2089, N2085, N1648, N959, N809);
or OR2 (N2090, N2082, N106);
nand NAND3 (N2091, N2079, N1387, N538);
and AND3 (N2092, N2090, N10, N702);
nor NOR2 (N2093, N2089, N1194);
and AND4 (N2094, N2076, N1175, N1803, N1688);
or OR4 (N2095, N2094, N751, N1027, N399);
xor XOR2 (N2096, N2083, N1196);
and AND3 (N2097, N2080, N115, N1974);
buf BUF1 (N2098, N2086);
not NOT1 (N2099, N2066);
or OR3 (N2100, N2091, N1282, N589);
nand NAND3 (N2101, N2093, N1432, N216);
and AND4 (N2102, N2097, N542, N142, N1790);
or OR3 (N2103, N2084, N551, N1242);
not NOT1 (N2104, N2098);
xor XOR2 (N2105, N2096, N1550);
buf BUF1 (N2106, N2101);
buf BUF1 (N2107, N2100);
xor XOR2 (N2108, N2103, N1971);
and AND2 (N2109, N2099, N1287);
buf BUF1 (N2110, N2104);
nand NAND4 (N2111, N2092, N1447, N1113, N1670);
not NOT1 (N2112, N2102);
nand NAND4 (N2113, N2109, N1500, N2096, N1128);
xor XOR2 (N2114, N2107, N1947);
or OR3 (N2115, N2112, N1621, N2098);
not NOT1 (N2116, N2111);
buf BUF1 (N2117, N2114);
buf BUF1 (N2118, N2110);
buf BUF1 (N2119, N2108);
or OR4 (N2120, N2095, N1967, N1876, N63);
buf BUF1 (N2121, N2118);
nand NAND2 (N2122, N2105, N746);
or OR2 (N2123, N2088, N1099);
nand NAND4 (N2124, N2121, N1591, N907, N823);
and AND2 (N2125, N2106, N1319);
nor NOR4 (N2126, N2117, N2054, N326, N1640);
nand NAND2 (N2127, N2116, N175);
buf BUF1 (N2128, N2119);
and AND3 (N2129, N2128, N536, N1805);
xor XOR2 (N2130, N2125, N914);
nor NOR2 (N2131, N2123, N274);
nand NAND3 (N2132, N2120, N715, N966);
or OR4 (N2133, N2129, N705, N1750, N842);
nand NAND4 (N2134, N2115, N234, N1522, N54);
or OR3 (N2135, N2130, N1025, N987);
not NOT1 (N2136, N2126);
and AND2 (N2137, N2132, N895);
nor NOR4 (N2138, N2137, N475, N1632, N1385);
nand NAND3 (N2139, N2134, N1034, N350);
nand NAND2 (N2140, N2113, N124);
or OR2 (N2141, N2127, N1693);
or OR2 (N2142, N2133, N1487);
nand NAND2 (N2143, N2139, N910);
buf BUF1 (N2144, N2138);
or OR4 (N2145, N2142, N1250, N1194, N1413);
or OR3 (N2146, N2140, N844, N1510);
or OR3 (N2147, N2144, N1203, N1620);
buf BUF1 (N2148, N2131);
nand NAND4 (N2149, N2122, N1304, N929, N543);
or OR3 (N2150, N2148, N434, N519);
not NOT1 (N2151, N2145);
and AND4 (N2152, N2151, N981, N830, N54);
buf BUF1 (N2153, N2136);
not NOT1 (N2154, N2147);
nor NOR3 (N2155, N2149, N2094, N2047);
and AND2 (N2156, N2155, N1663);
not NOT1 (N2157, N2141);
or OR4 (N2158, N2146, N1337, N1701, N1533);
xor XOR2 (N2159, N2152, N1380);
nor NOR3 (N2160, N2154, N2130, N1517);
buf BUF1 (N2161, N2160);
nand NAND3 (N2162, N2158, N710, N628);
buf BUF1 (N2163, N2161);
or OR3 (N2164, N2153, N545, N1812);
xor XOR2 (N2165, N2159, N1748);
nand NAND2 (N2166, N2162, N1478);
or OR4 (N2167, N2135, N1666, N714, N2062);
xor XOR2 (N2168, N2165, N578);
xor XOR2 (N2169, N2156, N527);
buf BUF1 (N2170, N2150);
nor NOR3 (N2171, N2143, N311, N525);
nor NOR4 (N2172, N2163, N1184, N1794, N413);
xor XOR2 (N2173, N2157, N1965);
nor NOR3 (N2174, N2172, N971, N1019);
or OR4 (N2175, N2166, N1487, N1790, N1728);
and AND4 (N2176, N2168, N805, N1368, N1938);
buf BUF1 (N2177, N2170);
buf BUF1 (N2178, N2176);
and AND4 (N2179, N2169, N1192, N28, N941);
or OR2 (N2180, N2171, N485);
nor NOR2 (N2181, N2174, N208);
nand NAND2 (N2182, N2179, N328);
and AND4 (N2183, N2181, N1861, N798, N590);
and AND4 (N2184, N2175, N706, N102, N1561);
not NOT1 (N2185, N2173);
buf BUF1 (N2186, N2167);
nor NOR3 (N2187, N2178, N1440, N20);
buf BUF1 (N2188, N2164);
and AND3 (N2189, N2180, N539, N2037);
xor XOR2 (N2190, N2177, N1180);
and AND4 (N2191, N2190, N1824, N1685, N1336);
buf BUF1 (N2192, N2188);
xor XOR2 (N2193, N2192, N170);
and AND2 (N2194, N2189, N680);
and AND2 (N2195, N2194, N2001);
and AND4 (N2196, N2186, N1780, N384, N1511);
nand NAND3 (N2197, N2191, N1327, N652);
nand NAND4 (N2198, N2185, N1005, N1124, N486);
xor XOR2 (N2199, N2183, N1207);
buf BUF1 (N2200, N2196);
or OR3 (N2201, N2184, N199, N444);
xor XOR2 (N2202, N2200, N508);
and AND3 (N2203, N2198, N464, N1295);
nor NOR3 (N2204, N2202, N1514, N574);
nor NOR3 (N2205, N2197, N1763, N348);
or OR4 (N2206, N2201, N1540, N1336, N1374);
xor XOR2 (N2207, N2187, N1779);
buf BUF1 (N2208, N2203);
xor XOR2 (N2209, N2182, N2148);
or OR3 (N2210, N2199, N685, N354);
not NOT1 (N2211, N2210);
not NOT1 (N2212, N2209);
nand NAND4 (N2213, N2193, N1824, N1186, N1478);
buf BUF1 (N2214, N2213);
or OR2 (N2215, N2204, N124);
not NOT1 (N2216, N2205);
and AND4 (N2217, N2124, N1590, N1309, N1665);
or OR4 (N2218, N2208, N802, N2132, N1112);
nor NOR4 (N2219, N2214, N20, N1959, N523);
buf BUF1 (N2220, N2216);
nor NOR3 (N2221, N2215, N1620, N884);
nand NAND2 (N2222, N2217, N834);
not NOT1 (N2223, N2207);
and AND2 (N2224, N2221, N1705);
xor XOR2 (N2225, N2223, N439);
and AND4 (N2226, N2224, N1126, N798, N1685);
not NOT1 (N2227, N2220);
not NOT1 (N2228, N2212);
or OR4 (N2229, N2228, N240, N269, N486);
or OR2 (N2230, N2225, N507);
buf BUF1 (N2231, N2206);
and AND2 (N2232, N2219, N80);
or OR3 (N2233, N2227, N1865, N1620);
not NOT1 (N2234, N2218);
not NOT1 (N2235, N2233);
nor NOR4 (N2236, N2232, N1482, N2043, N513);
not NOT1 (N2237, N2234);
nand NAND3 (N2238, N2231, N619, N595);
nor NOR3 (N2239, N2195, N523, N377);
not NOT1 (N2240, N2237);
nand NAND3 (N2241, N2230, N1010, N1427);
and AND2 (N2242, N2235, N1825);
nand NAND4 (N2243, N2222, N2035, N1615, N955);
nand NAND4 (N2244, N2226, N1559, N1737, N1956);
buf BUF1 (N2245, N2244);
not NOT1 (N2246, N2241);
nor NOR2 (N2247, N2238, N763);
and AND2 (N2248, N2243, N380);
nor NOR4 (N2249, N2245, N790, N2054, N366);
buf BUF1 (N2250, N2236);
not NOT1 (N2251, N2246);
nand NAND4 (N2252, N2239, N1178, N437, N1918);
nor NOR4 (N2253, N2240, N2064, N1559, N1369);
xor XOR2 (N2254, N2250, N191);
and AND4 (N2255, N2247, N186, N1062, N1906);
buf BUF1 (N2256, N2249);
xor XOR2 (N2257, N2256, N2202);
not NOT1 (N2258, N2257);
nand NAND3 (N2259, N2258, N1712, N1653);
nand NAND3 (N2260, N2251, N6, N2048);
xor XOR2 (N2261, N2248, N1588);
nor NOR4 (N2262, N2253, N292, N683, N278);
nand NAND4 (N2263, N2211, N1109, N92, N501);
xor XOR2 (N2264, N2229, N1381);
not NOT1 (N2265, N2262);
xor XOR2 (N2266, N2242, N497);
buf BUF1 (N2267, N2254);
or OR3 (N2268, N2259, N2058, N1913);
nor NOR4 (N2269, N2264, N1523, N698, N1592);
nor NOR3 (N2270, N2267, N947, N388);
or OR3 (N2271, N2266, N2079, N918);
nor NOR4 (N2272, N2265, N765, N978, N1863);
not NOT1 (N2273, N2271);
nor NOR2 (N2274, N2270, N242);
and AND3 (N2275, N2269, N1026, N1829);
xor XOR2 (N2276, N2263, N2062);
and AND3 (N2277, N2275, N1444, N1510);
or OR3 (N2278, N2255, N2203, N1354);
buf BUF1 (N2279, N2252);
nand NAND3 (N2280, N2278, N1045, N1091);
xor XOR2 (N2281, N2274, N1868);
and AND4 (N2282, N2273, N123, N1703, N1549);
buf BUF1 (N2283, N2268);
not NOT1 (N2284, N2261);
not NOT1 (N2285, N2283);
and AND2 (N2286, N2279, N2267);
and AND2 (N2287, N2281, N1312);
or OR3 (N2288, N2287, N1905, N1799);
nor NOR2 (N2289, N2280, N1050);
nor NOR2 (N2290, N2277, N2029);
xor XOR2 (N2291, N2276, N1861);
and AND3 (N2292, N2285, N2183, N2042);
nor NOR4 (N2293, N2289, N874, N1134, N1502);
xor XOR2 (N2294, N2293, N246);
nand NAND4 (N2295, N2282, N724, N496, N1715);
nand NAND2 (N2296, N2286, N1418);
not NOT1 (N2297, N2272);
and AND4 (N2298, N2295, N1447, N460, N2229);
xor XOR2 (N2299, N2260, N976);
nor NOR4 (N2300, N2294, N869, N1853, N60);
nor NOR4 (N2301, N2299, N231, N1012, N1873);
xor XOR2 (N2302, N2288, N2046);
buf BUF1 (N2303, N2284);
or OR2 (N2304, N2297, N1241);
or OR3 (N2305, N2302, N722, N1291);
not NOT1 (N2306, N2292);
nand NAND4 (N2307, N2303, N1811, N1711, N805);
buf BUF1 (N2308, N2301);
or OR4 (N2309, N2307, N1026, N275, N1391);
xor XOR2 (N2310, N2309, N1039);
nor NOR2 (N2311, N2290, N1883);
nand NAND3 (N2312, N2304, N2138, N1309);
nor NOR3 (N2313, N2311, N171, N1928);
or OR3 (N2314, N2291, N1600, N1338);
xor XOR2 (N2315, N2298, N571);
nand NAND4 (N2316, N2305, N496, N1783, N2299);
buf BUF1 (N2317, N2315);
and AND3 (N2318, N2314, N368, N1812);
nor NOR4 (N2319, N2316, N875, N555, N2207);
nand NAND4 (N2320, N2312, N1343, N61, N436);
xor XOR2 (N2321, N2313, N1356);
nand NAND2 (N2322, N2306, N1023);
and AND3 (N2323, N2318, N260, N1201);
and AND3 (N2324, N2317, N1219, N486);
nand NAND4 (N2325, N2308, N1121, N1094, N1179);
not NOT1 (N2326, N2324);
nand NAND2 (N2327, N2310, N910);
nor NOR2 (N2328, N2323, N373);
nand NAND3 (N2329, N2322, N2255, N848);
xor XOR2 (N2330, N2296, N2201);
buf BUF1 (N2331, N2327);
xor XOR2 (N2332, N2326, N440);
or OR3 (N2333, N2320, N2024, N1480);
not NOT1 (N2334, N2328);
nand NAND4 (N2335, N2325, N994, N490, N244);
or OR2 (N2336, N2319, N643);
xor XOR2 (N2337, N2333, N1641);
nand NAND2 (N2338, N2334, N1402);
or OR2 (N2339, N2330, N937);
nor NOR4 (N2340, N2329, N263, N1946, N951);
buf BUF1 (N2341, N2335);
nand NAND3 (N2342, N2321, N439, N616);
xor XOR2 (N2343, N2342, N1116);
xor XOR2 (N2344, N2341, N862);
xor XOR2 (N2345, N2340, N1395);
nand NAND2 (N2346, N2300, N796);
or OR4 (N2347, N2338, N898, N1649, N613);
or OR4 (N2348, N2343, N1284, N1979, N2152);
and AND3 (N2349, N2337, N118, N2008);
buf BUF1 (N2350, N2332);
nand NAND3 (N2351, N2350, N1625, N973);
or OR4 (N2352, N2344, N1371, N1164, N1970);
xor XOR2 (N2353, N2336, N995);
nand NAND2 (N2354, N2331, N1338);
nor NOR4 (N2355, N2351, N2065, N645, N1599);
buf BUF1 (N2356, N2349);
buf BUF1 (N2357, N2356);
buf BUF1 (N2358, N2347);
nand NAND4 (N2359, N2352, N228, N1887, N2309);
not NOT1 (N2360, N2353);
nand NAND3 (N2361, N2357, N1537, N1574);
xor XOR2 (N2362, N2345, N1582);
buf BUF1 (N2363, N2358);
nand NAND3 (N2364, N2354, N856, N1434);
buf BUF1 (N2365, N2355);
nand NAND3 (N2366, N2362, N1550, N1326);
xor XOR2 (N2367, N2361, N1969);
not NOT1 (N2368, N2346);
xor XOR2 (N2369, N2366, N1623);
or OR3 (N2370, N2368, N586, N1885);
nand NAND3 (N2371, N2369, N1701, N471);
nand NAND4 (N2372, N2348, N1776, N1269, N1758);
xor XOR2 (N2373, N2339, N2291);
or OR3 (N2374, N2360, N158, N671);
buf BUF1 (N2375, N2359);
and AND2 (N2376, N2367, N1762);
nand NAND3 (N2377, N2371, N2063, N675);
buf BUF1 (N2378, N2372);
not NOT1 (N2379, N2377);
nor NOR3 (N2380, N2378, N1680, N81);
not NOT1 (N2381, N2370);
xor XOR2 (N2382, N2376, N1354);
or OR2 (N2383, N2380, N1964);
not NOT1 (N2384, N2374);
and AND2 (N2385, N2382, N1137);
nor NOR4 (N2386, N2385, N1343, N1743, N806);
not NOT1 (N2387, N2383);
nand NAND3 (N2388, N2375, N1481, N2193);
buf BUF1 (N2389, N2365);
or OR4 (N2390, N2388, N626, N1201, N1064);
not NOT1 (N2391, N2387);
nor NOR3 (N2392, N2379, N49, N21);
not NOT1 (N2393, N2381);
xor XOR2 (N2394, N2363, N1312);
not NOT1 (N2395, N2392);
or OR4 (N2396, N2386, N571, N1084, N1999);
or OR2 (N2397, N2390, N657);
nor NOR4 (N2398, N2393, N855, N954, N60);
and AND3 (N2399, N2397, N2063, N2161);
nand NAND4 (N2400, N2395, N436, N2219, N1605);
or OR4 (N2401, N2394, N1827, N1519, N2050);
xor XOR2 (N2402, N2389, N2153);
or OR2 (N2403, N2398, N1469);
or OR4 (N2404, N2403, N528, N1659, N1761);
nand NAND3 (N2405, N2384, N2128, N735);
and AND3 (N2406, N2402, N202, N1301);
nand NAND2 (N2407, N2396, N124);
buf BUF1 (N2408, N2404);
or OR2 (N2409, N2364, N1121);
nand NAND2 (N2410, N2400, N1403);
or OR4 (N2411, N2408, N959, N1254, N482);
nor NOR3 (N2412, N2373, N1650, N593);
buf BUF1 (N2413, N2409);
not NOT1 (N2414, N2406);
buf BUF1 (N2415, N2407);
xor XOR2 (N2416, N2405, N2359);
not NOT1 (N2417, N2413);
buf BUF1 (N2418, N2416);
buf BUF1 (N2419, N2414);
not NOT1 (N2420, N2391);
buf BUF1 (N2421, N2399);
not NOT1 (N2422, N2411);
nand NAND3 (N2423, N2412, N1496, N1233);
or OR3 (N2424, N2423, N1729, N111);
and AND4 (N2425, N2415, N1133, N977, N125);
not NOT1 (N2426, N2424);
and AND3 (N2427, N2410, N67, N92);
not NOT1 (N2428, N2417);
nand NAND4 (N2429, N2419, N823, N474, N1833);
and AND4 (N2430, N2422, N2417, N2329, N2391);
xor XOR2 (N2431, N2420, N82);
or OR3 (N2432, N2425, N1437, N1282);
xor XOR2 (N2433, N2431, N1414);
xor XOR2 (N2434, N2429, N1072);
and AND2 (N2435, N2401, N2013);
nand NAND3 (N2436, N2427, N421, N949);
not NOT1 (N2437, N2421);
nor NOR4 (N2438, N2432, N1754, N1819, N2097);
or OR2 (N2439, N2430, N1040);
buf BUF1 (N2440, N2437);
or OR2 (N2441, N2436, N2012);
xor XOR2 (N2442, N2439, N2164);
nor NOR3 (N2443, N2434, N944, N1357);
nand NAND2 (N2444, N2441, N2414);
xor XOR2 (N2445, N2418, N1352);
or OR4 (N2446, N2433, N1112, N1336, N706);
buf BUF1 (N2447, N2438);
nor NOR4 (N2448, N2435, N1705, N1671, N1612);
and AND3 (N2449, N2445, N495, N2172);
xor XOR2 (N2450, N2442, N268);
xor XOR2 (N2451, N2450, N2229);
not NOT1 (N2452, N2444);
xor XOR2 (N2453, N2449, N1302);
and AND3 (N2454, N2452, N1555, N1192);
xor XOR2 (N2455, N2440, N558);
and AND3 (N2456, N2451, N2024, N1882);
not NOT1 (N2457, N2443);
not NOT1 (N2458, N2428);
nand NAND3 (N2459, N2453, N1711, N293);
nor NOR4 (N2460, N2447, N1381, N1805, N16);
or OR2 (N2461, N2459, N343);
buf BUF1 (N2462, N2457);
nand NAND2 (N2463, N2454, N1048);
xor XOR2 (N2464, N2460, N1293);
or OR4 (N2465, N2455, N394, N2035, N982);
and AND4 (N2466, N2461, N1383, N2185, N134);
and AND2 (N2467, N2426, N960);
and AND2 (N2468, N2463, N1472);
buf BUF1 (N2469, N2465);
buf BUF1 (N2470, N2466);
buf BUF1 (N2471, N2448);
buf BUF1 (N2472, N2464);
or OR3 (N2473, N2468, N1921, N2323);
buf BUF1 (N2474, N2467);
buf BUF1 (N2475, N2462);
not NOT1 (N2476, N2475);
nor NOR4 (N2477, N2470, N554, N1082, N514);
not NOT1 (N2478, N2458);
nor NOR3 (N2479, N2474, N2338, N700);
buf BUF1 (N2480, N2478);
xor XOR2 (N2481, N2446, N1193);
nor NOR4 (N2482, N2473, N807, N880, N1618);
nor NOR3 (N2483, N2472, N2327, N838);
xor XOR2 (N2484, N2480, N1925);
xor XOR2 (N2485, N2477, N1165);
xor XOR2 (N2486, N2482, N1137);
xor XOR2 (N2487, N2476, N1539);
and AND4 (N2488, N2479, N849, N389, N959);
nor NOR3 (N2489, N2487, N1606, N2090);
nand NAND3 (N2490, N2485, N497, N2327);
nor NOR2 (N2491, N2481, N780);
xor XOR2 (N2492, N2484, N1809);
not NOT1 (N2493, N2492);
nor NOR4 (N2494, N2493, N2217, N277, N467);
nor NOR3 (N2495, N2490, N2346, N116);
buf BUF1 (N2496, N2456);
not NOT1 (N2497, N2491);
nand NAND4 (N2498, N2486, N1722, N638, N2496);
or OR4 (N2499, N750, N1536, N837, N283);
buf BUF1 (N2500, N2471);
and AND4 (N2501, N2495, N2147, N1147, N2242);
xor XOR2 (N2502, N2469, N1133);
nand NAND2 (N2503, N2489, N2088);
and AND2 (N2504, N2500, N1980);
xor XOR2 (N2505, N2497, N1297);
buf BUF1 (N2506, N2488);
nor NOR4 (N2507, N2501, N1532, N987, N1765);
or OR2 (N2508, N2504, N1450);
buf BUF1 (N2509, N2494);
and AND2 (N2510, N2498, N2206);
xor XOR2 (N2511, N2508, N2282);
and AND3 (N2512, N2509, N1060, N2366);
and AND4 (N2513, N2483, N264, N597, N1262);
or OR2 (N2514, N2511, N385);
nand NAND4 (N2515, N2503, N370, N1127, N591);
not NOT1 (N2516, N2510);
not NOT1 (N2517, N2514);
xor XOR2 (N2518, N2505, N1567);
xor XOR2 (N2519, N2513, N1576);
not NOT1 (N2520, N2506);
nor NOR4 (N2521, N2512, N1270, N2063, N1168);
nor NOR4 (N2522, N2516, N1666, N1871, N552);
and AND4 (N2523, N2522, N871, N833, N1195);
xor XOR2 (N2524, N2517, N247);
buf BUF1 (N2525, N2519);
and AND4 (N2526, N2507, N1505, N1089, N2294);
nand NAND3 (N2527, N2499, N779, N2264);
nand NAND3 (N2528, N2527, N545, N2507);
or OR4 (N2529, N2523, N484, N1457, N183);
nor NOR2 (N2530, N2515, N744);
buf BUF1 (N2531, N2520);
not NOT1 (N2532, N2530);
or OR4 (N2533, N2528, N2101, N1973, N575);
and AND2 (N2534, N2529, N577);
buf BUF1 (N2535, N2526);
buf BUF1 (N2536, N2535);
nor NOR2 (N2537, N2525, N1022);
nand NAND2 (N2538, N2524, N1492);
nor NOR3 (N2539, N2533, N1574, N1766);
and AND2 (N2540, N2502, N141);
not NOT1 (N2541, N2536);
and AND2 (N2542, N2534, N2305);
and AND4 (N2543, N2521, N303, N817, N1258);
buf BUF1 (N2544, N2540);
buf BUF1 (N2545, N2541);
or OR4 (N2546, N2539, N52, N588, N405);
xor XOR2 (N2547, N2532, N2146);
nand NAND2 (N2548, N2543, N1460);
nor NOR4 (N2549, N2546, N1936, N585, N115);
xor XOR2 (N2550, N2544, N88);
or OR2 (N2551, N2537, N529);
xor XOR2 (N2552, N2551, N1400);
nand NAND4 (N2553, N2542, N758, N2414, N246);
and AND4 (N2554, N2538, N1474, N961, N2442);
xor XOR2 (N2555, N2552, N1012);
and AND2 (N2556, N2554, N1298);
or OR4 (N2557, N2545, N451, N2544, N1578);
and AND3 (N2558, N2553, N1715, N784);
nor NOR4 (N2559, N2548, N2170, N1484, N1697);
buf BUF1 (N2560, N2549);
nor NOR3 (N2561, N2555, N794, N453);
nand NAND4 (N2562, N2550, N948, N1724, N1038);
buf BUF1 (N2563, N2556);
not NOT1 (N2564, N2560);
buf BUF1 (N2565, N2558);
xor XOR2 (N2566, N2562, N885);
xor XOR2 (N2567, N2547, N981);
and AND2 (N2568, N2563, N1551);
not NOT1 (N2569, N2518);
buf BUF1 (N2570, N2566);
nor NOR2 (N2571, N2570, N1028);
nor NOR3 (N2572, N2567, N1325, N320);
not NOT1 (N2573, N2559);
nor NOR4 (N2574, N2557, N245, N111, N697);
nand NAND2 (N2575, N2573, N2093);
nand NAND4 (N2576, N2568, N1279, N512, N2255);
not NOT1 (N2577, N2561);
nor NOR3 (N2578, N2572, N2561, N388);
buf BUF1 (N2579, N2575);
or OR3 (N2580, N2579, N621, N1004);
or OR4 (N2581, N2574, N668, N1034, N301);
buf BUF1 (N2582, N2578);
xor XOR2 (N2583, N2581, N636);
nand NAND4 (N2584, N2565, N872, N2088, N1227);
nor NOR2 (N2585, N2531, N2350);
or OR2 (N2586, N2564, N1702);
and AND4 (N2587, N2576, N2186, N98, N2165);
not NOT1 (N2588, N2586);
or OR4 (N2589, N2582, N427, N1124, N2427);
buf BUF1 (N2590, N2577);
not NOT1 (N2591, N2587);
nor NOR4 (N2592, N2571, N410, N1945, N795);
nor NOR2 (N2593, N2583, N861);
nor NOR3 (N2594, N2585, N334, N1008);
or OR3 (N2595, N2588, N2329, N270);
nand NAND3 (N2596, N2569, N214, N267);
not NOT1 (N2597, N2584);
or OR4 (N2598, N2580, N2502, N2088, N760);
xor XOR2 (N2599, N2589, N630);
xor XOR2 (N2600, N2595, N2121);
not NOT1 (N2601, N2596);
not NOT1 (N2602, N2599);
nand NAND4 (N2603, N2594, N1005, N40, N1531);
buf BUF1 (N2604, N2590);
nor NOR2 (N2605, N2603, N1528);
xor XOR2 (N2606, N2602, N2337);
not NOT1 (N2607, N2606);
xor XOR2 (N2608, N2598, N512);
or OR2 (N2609, N2601, N1041);
nor NOR3 (N2610, N2592, N1574, N1530);
nand NAND4 (N2611, N2600, N526, N1509, N725);
nand NAND2 (N2612, N2591, N470);
or OR3 (N2613, N2608, N65, N829);
buf BUF1 (N2614, N2610);
not NOT1 (N2615, N2605);
not NOT1 (N2616, N2611);
and AND2 (N2617, N2607, N31);
xor XOR2 (N2618, N2617, N1597);
xor XOR2 (N2619, N2613, N1849);
nand NAND4 (N2620, N2615, N1099, N1717, N2250);
xor XOR2 (N2621, N2614, N304);
buf BUF1 (N2622, N2593);
nand NAND4 (N2623, N2616, N2124, N977, N240);
and AND2 (N2624, N2622, N1020);
xor XOR2 (N2625, N2621, N274);
not NOT1 (N2626, N2609);
or OR2 (N2627, N2624, N461);
buf BUF1 (N2628, N2597);
not NOT1 (N2629, N2604);
and AND2 (N2630, N2627, N601);
not NOT1 (N2631, N2628);
buf BUF1 (N2632, N2625);
nor NOR2 (N2633, N2631, N1034);
not NOT1 (N2634, N2620);
xor XOR2 (N2635, N2629, N2368);
buf BUF1 (N2636, N2630);
nand NAND4 (N2637, N2626, N118, N1970, N2236);
nor NOR2 (N2638, N2634, N1094);
nor NOR3 (N2639, N2623, N1533, N120);
nand NAND4 (N2640, N2618, N437, N1787, N641);
and AND4 (N2641, N2612, N677, N309, N779);
nand NAND2 (N2642, N2636, N819);
or OR2 (N2643, N2638, N1364);
not NOT1 (N2644, N2633);
and AND3 (N2645, N2635, N225, N591);
and AND2 (N2646, N2639, N1235);
buf BUF1 (N2647, N2641);
not NOT1 (N2648, N2645);
nor NOR2 (N2649, N2646, N1000);
xor XOR2 (N2650, N2640, N2332);
nor NOR2 (N2651, N2619, N468);
not NOT1 (N2652, N2637);
buf BUF1 (N2653, N2649);
or OR4 (N2654, N2651, N1959, N2175, N576);
and AND3 (N2655, N2652, N809, N2480);
not NOT1 (N2656, N2648);
xor XOR2 (N2657, N2650, N214);
buf BUF1 (N2658, N2654);
and AND2 (N2659, N2643, N1034);
and AND3 (N2660, N2655, N236, N1339);
not NOT1 (N2661, N2642);
or OR2 (N2662, N2658, N1717);
nand NAND2 (N2663, N2661, N804);
and AND3 (N2664, N2656, N537, N2590);
not NOT1 (N2665, N2657);
and AND4 (N2666, N2660, N1566, N868, N199);
and AND2 (N2667, N2647, N847);
xor XOR2 (N2668, N2665, N2032);
buf BUF1 (N2669, N2666);
nor NOR2 (N2670, N2632, N1067);
nor NOR4 (N2671, N2669, N2191, N2126, N2309);
nor NOR2 (N2672, N2644, N1902);
or OR4 (N2673, N2671, N1675, N1850, N1666);
nor NOR3 (N2674, N2668, N1848, N420);
buf BUF1 (N2675, N2659);
or OR3 (N2676, N2662, N1306, N181);
not NOT1 (N2677, N2676);
and AND2 (N2678, N2673, N281);
buf BUF1 (N2679, N2678);
and AND2 (N2680, N2677, N165);
nor NOR4 (N2681, N2664, N1476, N1531, N765);
or OR2 (N2682, N2667, N1341);
xor XOR2 (N2683, N2680, N1380);
buf BUF1 (N2684, N2674);
not NOT1 (N2685, N2663);
and AND4 (N2686, N2685, N599, N1804, N398);
buf BUF1 (N2687, N2684);
and AND3 (N2688, N2683, N260, N2219);
not NOT1 (N2689, N2679);
nor NOR4 (N2690, N2682, N2397, N2223, N384);
xor XOR2 (N2691, N2675, N282);
buf BUF1 (N2692, N2653);
not NOT1 (N2693, N2670);
nand NAND4 (N2694, N2692, N597, N1367, N652);
buf BUF1 (N2695, N2672);
nand NAND4 (N2696, N2688, N559, N959, N2235);
nand NAND4 (N2697, N2687, N1603, N484, N90);
or OR4 (N2698, N2686, N813, N1081, N502);
xor XOR2 (N2699, N2694, N487);
nor NOR4 (N2700, N2681, N1312, N2458, N1997);
nor NOR3 (N2701, N2700, N277, N283);
xor XOR2 (N2702, N2693, N2284);
or OR4 (N2703, N2691, N1817, N2591, N34);
and AND3 (N2704, N2701, N522, N1051);
nor NOR2 (N2705, N2695, N485);
nor NOR3 (N2706, N2696, N1774, N1463);
nor NOR3 (N2707, N2697, N1274, N1074);
buf BUF1 (N2708, N2704);
xor XOR2 (N2709, N2708, N1637);
xor XOR2 (N2710, N2689, N1156);
buf BUF1 (N2711, N2709);
nor NOR3 (N2712, N2699, N1513, N237);
or OR2 (N2713, N2702, N790);
and AND2 (N2714, N2705, N1664);
or OR3 (N2715, N2690, N2337, N2668);
and AND3 (N2716, N2715, N650, N2431);
nand NAND4 (N2717, N2711, N1675, N1294, N168);
nand NAND4 (N2718, N2707, N285, N2387, N1166);
xor XOR2 (N2719, N2703, N551);
xor XOR2 (N2720, N2706, N650);
and AND3 (N2721, N2714, N2615, N1487);
xor XOR2 (N2722, N2698, N862);
nand NAND2 (N2723, N2713, N239);
buf BUF1 (N2724, N2719);
and AND3 (N2725, N2720, N2300, N1410);
buf BUF1 (N2726, N2721);
buf BUF1 (N2727, N2717);
nor NOR3 (N2728, N2710, N1328, N552);
xor XOR2 (N2729, N2728, N392);
not NOT1 (N2730, N2718);
nor NOR2 (N2731, N2729, N967);
nor NOR3 (N2732, N2731, N1929, N794);
xor XOR2 (N2733, N2724, N63);
or OR2 (N2734, N2722, N1814);
nand NAND3 (N2735, N2723, N269, N1371);
nand NAND4 (N2736, N2727, N1303, N2301, N1887);
or OR4 (N2737, N2730, N1745, N1162, N2059);
buf BUF1 (N2738, N2712);
not NOT1 (N2739, N2738);
xor XOR2 (N2740, N2725, N754);
not NOT1 (N2741, N2737);
nor NOR3 (N2742, N2736, N1926, N1316);
nor NOR2 (N2743, N2732, N1845);
nor NOR2 (N2744, N2742, N757);
or OR4 (N2745, N2740, N60, N1042, N1149);
and AND4 (N2746, N2716, N107, N1036, N1392);
or OR4 (N2747, N2741, N2131, N72, N1215);
nand NAND2 (N2748, N2746, N135);
and AND4 (N2749, N2748, N2036, N601, N1461);
not NOT1 (N2750, N2743);
buf BUF1 (N2751, N2726);
buf BUF1 (N2752, N2744);
or OR4 (N2753, N2747, N76, N1565, N1317);
and AND4 (N2754, N2739, N2296, N877, N826);
or OR2 (N2755, N2750, N389);
buf BUF1 (N2756, N2735);
and AND3 (N2757, N2734, N2149, N79);
nand NAND4 (N2758, N2745, N4, N1733, N599);
nand NAND2 (N2759, N2755, N1500);
or OR2 (N2760, N2758, N1270);
nand NAND4 (N2761, N2760, N1723, N2490, N125);
nor NOR3 (N2762, N2753, N259, N119);
buf BUF1 (N2763, N2761);
or OR2 (N2764, N2757, N1672);
nor NOR3 (N2765, N2762, N489, N1436);
nand NAND2 (N2766, N2759, N1788);
and AND3 (N2767, N2751, N71, N2548);
not NOT1 (N2768, N2749);
or OR4 (N2769, N2764, N2686, N448, N1768);
buf BUF1 (N2770, N2763);
nor NOR2 (N2771, N2752, N1290);
and AND4 (N2772, N2770, N804, N2307, N1122);
and AND2 (N2773, N2769, N634);
not NOT1 (N2774, N2733);
or OR4 (N2775, N2768, N2570, N2255, N1403);
and AND2 (N2776, N2774, N1308);
or OR3 (N2777, N2766, N2605, N32);
nor NOR2 (N2778, N2765, N1967);
buf BUF1 (N2779, N2767);
nor NOR4 (N2780, N2775, N1909, N2725, N1040);
and AND3 (N2781, N2777, N197, N186);
xor XOR2 (N2782, N2756, N802);
nand NAND3 (N2783, N2778, N253, N910);
xor XOR2 (N2784, N2754, N1931);
and AND2 (N2785, N2780, N1128);
or OR4 (N2786, N2776, N2195, N1724, N1297);
and AND4 (N2787, N2772, N1016, N53, N264);
not NOT1 (N2788, N2783);
and AND2 (N2789, N2779, N1206);
nor NOR2 (N2790, N2785, N1213);
xor XOR2 (N2791, N2790, N440);
nor NOR4 (N2792, N2788, N1904, N1353, N1327);
and AND2 (N2793, N2782, N1692);
nand NAND3 (N2794, N2789, N16, N2247);
buf BUF1 (N2795, N2787);
and AND4 (N2796, N2781, N771, N1576, N2445);
buf BUF1 (N2797, N2786);
buf BUF1 (N2798, N2771);
and AND3 (N2799, N2795, N936, N1821);
nand NAND3 (N2800, N2791, N2284, N1775);
nand NAND3 (N2801, N2797, N1314, N921);
buf BUF1 (N2802, N2793);
xor XOR2 (N2803, N2794, N1296);
buf BUF1 (N2804, N2792);
buf BUF1 (N2805, N2796);
or OR4 (N2806, N2773, N1915, N576, N689);
nor NOR2 (N2807, N2804, N583);
nor NOR3 (N2808, N2801, N2685, N2669);
or OR2 (N2809, N2803, N2085);
nor NOR4 (N2810, N2784, N1213, N648, N1545);
nand NAND2 (N2811, N2810, N2600);
or OR3 (N2812, N2805, N2662, N1448);
buf BUF1 (N2813, N2807);
or OR2 (N2814, N2802, N929);
not NOT1 (N2815, N2800);
xor XOR2 (N2816, N2814, N257);
xor XOR2 (N2817, N2806, N1390);
nor NOR2 (N2818, N2811, N1395);
nand NAND3 (N2819, N2809, N2278, N520);
xor XOR2 (N2820, N2808, N1666);
and AND2 (N2821, N2813, N2779);
xor XOR2 (N2822, N2817, N1655);
buf BUF1 (N2823, N2816);
or OR3 (N2824, N2815, N212, N631);
or OR3 (N2825, N2798, N1191, N534);
xor XOR2 (N2826, N2812, N984);
buf BUF1 (N2827, N2825);
buf BUF1 (N2828, N2824);
nand NAND3 (N2829, N2822, N1531, N2368);
xor XOR2 (N2830, N2828, N2253);
and AND4 (N2831, N2823, N2343, N1181, N1376);
not NOT1 (N2832, N2830);
xor XOR2 (N2833, N2819, N1769);
nand NAND3 (N2834, N2820, N2558, N1967);
not NOT1 (N2835, N2832);
xor XOR2 (N2836, N2821, N80);
xor XOR2 (N2837, N2834, N1492);
or OR4 (N2838, N2831, N1606, N1560, N246);
xor XOR2 (N2839, N2826, N2211);
not NOT1 (N2840, N2837);
xor XOR2 (N2841, N2833, N298);
or OR4 (N2842, N2835, N1922, N1090, N173);
nand NAND4 (N2843, N2841, N2480, N188, N2371);
or OR3 (N2844, N2840, N2762, N328);
and AND2 (N2845, N2838, N1650);
or OR3 (N2846, N2818, N418, N2780);
xor XOR2 (N2847, N2839, N1819);
not NOT1 (N2848, N2847);
nand NAND2 (N2849, N2799, N1005);
and AND3 (N2850, N2842, N2346, N682);
and AND3 (N2851, N2845, N1879, N1914);
nor NOR3 (N2852, N2846, N311, N1305);
buf BUF1 (N2853, N2836);
nor NOR2 (N2854, N2829, N2255);
not NOT1 (N2855, N2848);
buf BUF1 (N2856, N2855);
xor XOR2 (N2857, N2843, N2140);
buf BUF1 (N2858, N2849);
buf BUF1 (N2859, N2827);
or OR4 (N2860, N2851, N634, N1743, N1109);
nand NAND2 (N2861, N2857, N1078);
and AND2 (N2862, N2856, N1410);
buf BUF1 (N2863, N2861);
not NOT1 (N2864, N2862);
nor NOR3 (N2865, N2852, N1350, N2711);
xor XOR2 (N2866, N2860, N620);
not NOT1 (N2867, N2865);
not NOT1 (N2868, N2844);
and AND2 (N2869, N2850, N1898);
xor XOR2 (N2870, N2866, N2745);
buf BUF1 (N2871, N2863);
nor NOR2 (N2872, N2853, N2099);
nor NOR3 (N2873, N2868, N279, N151);
buf BUF1 (N2874, N2859);
buf BUF1 (N2875, N2854);
and AND2 (N2876, N2873, N1118);
nand NAND3 (N2877, N2876, N719, N1511);
not NOT1 (N2878, N2864);
and AND4 (N2879, N2878, N268, N1977, N85);
nor NOR4 (N2880, N2875, N703, N826, N925);
or OR4 (N2881, N2871, N595, N1766, N449);
not NOT1 (N2882, N2874);
or OR3 (N2883, N2877, N204, N1654);
or OR2 (N2884, N2870, N2650);
nor NOR2 (N2885, N2858, N594);
buf BUF1 (N2886, N2869);
nand NAND3 (N2887, N2884, N2757, N1141);
or OR4 (N2888, N2880, N2434, N969, N500);
nor NOR3 (N2889, N2867, N1018, N1178);
xor XOR2 (N2890, N2872, N2830);
buf BUF1 (N2891, N2879);
nor NOR4 (N2892, N2886, N722, N759, N710);
xor XOR2 (N2893, N2888, N2442);
nor NOR3 (N2894, N2890, N264, N661);
not NOT1 (N2895, N2887);
buf BUF1 (N2896, N2882);
nor NOR3 (N2897, N2885, N1496, N80);
buf BUF1 (N2898, N2894);
or OR4 (N2899, N2892, N519, N901, N2261);
or OR3 (N2900, N2896, N995, N1330);
xor XOR2 (N2901, N2883, N847);
nor NOR2 (N2902, N2898, N2680);
or OR2 (N2903, N2895, N1168);
nand NAND3 (N2904, N2893, N1181, N2051);
or OR2 (N2905, N2881, N4);
and AND2 (N2906, N2891, N2035);
nor NOR3 (N2907, N2901, N2406, N2141);
or OR4 (N2908, N2902, N830, N1628, N262);
buf BUF1 (N2909, N2897);
xor XOR2 (N2910, N2907, N1090);
or OR4 (N2911, N2910, N1769, N2340, N2564);
nor NOR3 (N2912, N2903, N1685, N2569);
or OR4 (N2913, N2889, N1694, N429, N824);
or OR3 (N2914, N2899, N1225, N2425);
xor XOR2 (N2915, N2908, N424);
xor XOR2 (N2916, N2915, N1176);
nand NAND3 (N2917, N2916, N956, N618);
xor XOR2 (N2918, N2913, N2225);
not NOT1 (N2919, N2911);
nor NOR2 (N2920, N2909, N135);
not NOT1 (N2921, N2900);
nand NAND3 (N2922, N2921, N53, N1902);
not NOT1 (N2923, N2912);
nand NAND3 (N2924, N2918, N2604, N2294);
not NOT1 (N2925, N2920);
buf BUF1 (N2926, N2919);
or OR2 (N2927, N2914, N1706);
nor NOR4 (N2928, N2924, N33, N2238, N2479);
and AND4 (N2929, N2906, N2342, N860, N188);
not NOT1 (N2930, N2925);
xor XOR2 (N2931, N2926, N2295);
not NOT1 (N2932, N2922);
xor XOR2 (N2933, N2929, N2841);
not NOT1 (N2934, N2928);
nand NAND4 (N2935, N2904, N775, N2474, N405);
or OR4 (N2936, N2933, N2867, N1554, N1405);
and AND3 (N2937, N2935, N151, N663);
or OR2 (N2938, N2930, N600);
or OR2 (N2939, N2934, N2899);
buf BUF1 (N2940, N2905);
and AND3 (N2941, N2931, N1997, N1066);
xor XOR2 (N2942, N2927, N2256);
not NOT1 (N2943, N2939);
nand NAND2 (N2944, N2937, N1221);
nand NAND2 (N2945, N2917, N1287);
nor NOR4 (N2946, N2945, N1576, N1018, N470);
not NOT1 (N2947, N2942);
nand NAND4 (N2948, N2943, N1608, N2439, N2853);
nor NOR3 (N2949, N2940, N1095, N1894);
or OR4 (N2950, N2944, N7, N2092, N410);
or OR4 (N2951, N2950, N834, N1726, N1307);
xor XOR2 (N2952, N2923, N995);
xor XOR2 (N2953, N2936, N2121);
or OR4 (N2954, N2938, N2007, N1785, N2512);
nand NAND4 (N2955, N2954, N2010, N818, N84);
nor NOR2 (N2956, N2947, N173);
buf BUF1 (N2957, N2953);
and AND4 (N2958, N2952, N2033, N1465, N1108);
not NOT1 (N2959, N2957);
or OR2 (N2960, N2959, N2106);
not NOT1 (N2961, N2951);
nand NAND4 (N2962, N2956, N2465, N2471, N30);
nand NAND4 (N2963, N2962, N1690, N2467, N1202);
buf BUF1 (N2964, N2960);
nor NOR3 (N2965, N2941, N2882, N2513);
and AND4 (N2966, N2948, N1915, N2415, N890);
buf BUF1 (N2967, N2963);
nand NAND2 (N2968, N2964, N2844);
and AND3 (N2969, N2967, N1011, N2627);
buf BUF1 (N2970, N2965);
not NOT1 (N2971, N2966);
nor NOR4 (N2972, N2969, N1841, N259, N1347);
nor NOR4 (N2973, N2972, N1882, N718, N724);
buf BUF1 (N2974, N2968);
or OR4 (N2975, N2932, N2391, N1482, N2507);
and AND4 (N2976, N2955, N2007, N2491, N1058);
nor NOR2 (N2977, N2975, N302);
buf BUF1 (N2978, N2971);
nand NAND2 (N2979, N2977, N50);
nand NAND2 (N2980, N2974, N1576);
buf BUF1 (N2981, N2979);
not NOT1 (N2982, N2980);
xor XOR2 (N2983, N2982, N1740);
buf BUF1 (N2984, N2958);
not NOT1 (N2985, N2961);
nor NOR3 (N2986, N2984, N1866, N1237);
or OR4 (N2987, N2946, N704, N1910, N2162);
not NOT1 (N2988, N2973);
nor NOR3 (N2989, N2985, N688, N1773);
and AND2 (N2990, N2988, N853);
and AND2 (N2991, N2949, N979);
and AND4 (N2992, N2986, N613, N2866, N1239);
xor XOR2 (N2993, N2989, N919);
not NOT1 (N2994, N2976);
and AND3 (N2995, N2993, N2278, N2174);
and AND2 (N2996, N2994, N2366);
nand NAND3 (N2997, N2983, N2484, N2022);
xor XOR2 (N2998, N2997, N566);
or OR4 (N2999, N2996, N333, N2339, N1457);
not NOT1 (N3000, N2991);
or OR2 (N3001, N2995, N1030);
or OR3 (N3002, N2987, N1348, N2621);
nand NAND4 (N3003, N2998, N2525, N1439, N2300);
nor NOR2 (N3004, N2999, N1155);
nand NAND4 (N3005, N2981, N437, N1189, N373);
nor NOR3 (N3006, N3000, N327, N1032);
or OR4 (N3007, N3003, N2546, N2047, N1720);
nand NAND4 (N3008, N3004, N923, N1426, N2033);
nand NAND3 (N3009, N2970, N494, N1968);
and AND3 (N3010, N2990, N833, N106);
buf BUF1 (N3011, N3009);
nor NOR3 (N3012, N3006, N1035, N2252);
xor XOR2 (N3013, N3007, N3012);
or OR4 (N3014, N2921, N1687, N1550, N2709);
not NOT1 (N3015, N3001);
and AND3 (N3016, N3002, N920, N2663);
and AND4 (N3017, N3014, N945, N2649, N1685);
buf BUF1 (N3018, N3008);
xor XOR2 (N3019, N3013, N2876);
or OR4 (N3020, N3017, N274, N1344, N133);
nand NAND3 (N3021, N3015, N691, N847);
buf BUF1 (N3022, N3010);
and AND4 (N3023, N2992, N651, N1024, N2056);
not NOT1 (N3024, N2978);
and AND3 (N3025, N3024, N1903, N1196);
and AND3 (N3026, N3019, N172, N580);
not NOT1 (N3027, N3023);
or OR4 (N3028, N3025, N1961, N415, N2569);
nor NOR2 (N3029, N3027, N2320);
or OR3 (N3030, N3028, N2617, N1342);
or OR3 (N3031, N3020, N2562, N2011);
nor NOR3 (N3032, N3022, N1559, N2505);
and AND4 (N3033, N3030, N76, N2812, N2344);
and AND2 (N3034, N3026, N886);
or OR4 (N3035, N3011, N2173, N1155, N1334);
buf BUF1 (N3036, N3035);
buf BUF1 (N3037, N3031);
and AND4 (N3038, N3033, N2872, N2871, N1891);
xor XOR2 (N3039, N3037, N942);
or OR3 (N3040, N3029, N2120, N861);
or OR2 (N3041, N3032, N3002);
and AND2 (N3042, N3036, N2100);
buf BUF1 (N3043, N3042);
or OR3 (N3044, N3018, N1139, N1033);
xor XOR2 (N3045, N3039, N2048);
nor NOR3 (N3046, N3005, N2203, N2420);
not NOT1 (N3047, N3034);
nand NAND3 (N3048, N3038, N975, N1690);
buf BUF1 (N3049, N3021);
xor XOR2 (N3050, N3044, N1401);
nand NAND2 (N3051, N3047, N1030);
and AND4 (N3052, N3043, N883, N2295, N2677);
not NOT1 (N3053, N3049);
not NOT1 (N3054, N3041);
xor XOR2 (N3055, N3046, N2132);
and AND4 (N3056, N3053, N299, N1617, N216);
not NOT1 (N3057, N3045);
xor XOR2 (N3058, N3050, N1745);
nand NAND2 (N3059, N3051, N2600);
nand NAND3 (N3060, N3040, N1972, N2344);
nor NOR2 (N3061, N3054, N1466);
buf BUF1 (N3062, N3055);
not NOT1 (N3063, N3062);
buf BUF1 (N3064, N3052);
nor NOR2 (N3065, N3061, N1747);
not NOT1 (N3066, N3048);
nor NOR3 (N3067, N3060, N642, N2774);
nand NAND3 (N3068, N3064, N438, N2352);
or OR2 (N3069, N3057, N1812);
nor NOR4 (N3070, N3069, N1099, N1033, N1982);
nand NAND2 (N3071, N3067, N319);
and AND2 (N3072, N3056, N1394);
buf BUF1 (N3073, N3068);
xor XOR2 (N3074, N3063, N250);
buf BUF1 (N3075, N3065);
or OR2 (N3076, N3059, N21);
not NOT1 (N3077, N3070);
nor NOR2 (N3078, N3016, N995);
or OR3 (N3079, N3073, N64, N1336);
or OR3 (N3080, N3077, N1475, N439);
or OR2 (N3081, N3058, N1107);
and AND4 (N3082, N3074, N2299, N1598, N1040);
buf BUF1 (N3083, N3078);
nor NOR2 (N3084, N3082, N2174);
nor NOR2 (N3085, N3080, N2574);
nand NAND3 (N3086, N3072, N1168, N40);
and AND4 (N3087, N3084, N2173, N1648, N2067);
and AND2 (N3088, N3079, N930);
or OR3 (N3089, N3081, N2939, N740);
and AND2 (N3090, N3088, N1211);
nand NAND3 (N3091, N3090, N767, N1693);
buf BUF1 (N3092, N3087);
or OR3 (N3093, N3083, N2641, N906);
nand NAND2 (N3094, N3066, N2916);
xor XOR2 (N3095, N3075, N674);
xor XOR2 (N3096, N3071, N608);
not NOT1 (N3097, N3096);
not NOT1 (N3098, N3076);
not NOT1 (N3099, N3091);
or OR4 (N3100, N3092, N751, N2913, N1708);
nand NAND4 (N3101, N3097, N453, N995, N2387);
or OR4 (N3102, N3100, N543, N2369, N46);
nand NAND4 (N3103, N3101, N235, N2865, N601);
not NOT1 (N3104, N3085);
and AND3 (N3105, N3103, N84, N1122);
nor NOR4 (N3106, N3102, N1204, N111, N1935);
xor XOR2 (N3107, N3099, N1834);
xor XOR2 (N3108, N3095, N2870);
or OR3 (N3109, N3093, N1488, N1484);
not NOT1 (N3110, N3098);
buf BUF1 (N3111, N3107);
nor NOR4 (N3112, N3105, N3092, N1709, N307);
xor XOR2 (N3113, N3111, N1443);
buf BUF1 (N3114, N3089);
nor NOR2 (N3115, N3094, N1471);
nand NAND3 (N3116, N3109, N1626, N1032);
and AND4 (N3117, N3116, N158, N1407, N46);
buf BUF1 (N3118, N3108);
buf BUF1 (N3119, N3112);
or OR4 (N3120, N3110, N2236, N1026, N676);
nand NAND2 (N3121, N3086, N2008);
nand NAND2 (N3122, N3117, N2485);
buf BUF1 (N3123, N3120);
buf BUF1 (N3124, N3123);
nor NOR3 (N3125, N3114, N310, N500);
nor NOR2 (N3126, N3124, N2788);
and AND2 (N3127, N3125, N748);
or OR2 (N3128, N3115, N1653);
not NOT1 (N3129, N3106);
not NOT1 (N3130, N3104);
nor NOR3 (N3131, N3128, N1542, N247);
and AND2 (N3132, N3129, N203);
nand NAND2 (N3133, N3132, N2672);
xor XOR2 (N3134, N3122, N1587);
and AND2 (N3135, N3134, N1668);
or OR2 (N3136, N3131, N516);
and AND2 (N3137, N3118, N919);
buf BUF1 (N3138, N3113);
nand NAND3 (N3139, N3136, N1785, N911);
nor NOR3 (N3140, N3126, N2434, N1961);
buf BUF1 (N3141, N3135);
buf BUF1 (N3142, N3137);
xor XOR2 (N3143, N3133, N21);
buf BUF1 (N3144, N3141);
nor NOR2 (N3145, N3144, N2982);
buf BUF1 (N3146, N3139);
buf BUF1 (N3147, N3121);
nor NOR2 (N3148, N3138, N2757);
and AND2 (N3149, N3130, N2608);
xor XOR2 (N3150, N3143, N983);
nand NAND2 (N3151, N3119, N1713);
nand NAND3 (N3152, N3148, N1896, N2951);
or OR4 (N3153, N3146, N1463, N1215, N179);
buf BUF1 (N3154, N3149);
nor NOR2 (N3155, N3153, N617);
xor XOR2 (N3156, N3150, N1462);
nor NOR3 (N3157, N3156, N365, N2665);
not NOT1 (N3158, N3127);
not NOT1 (N3159, N3152);
nor NOR3 (N3160, N3147, N888, N821);
buf BUF1 (N3161, N3145);
xor XOR2 (N3162, N3155, N276);
and AND3 (N3163, N3142, N428, N2075);
nand NAND2 (N3164, N3154, N412);
xor XOR2 (N3165, N3151, N3021);
nand NAND3 (N3166, N3157, N409, N323);
nand NAND4 (N3167, N3162, N941, N295, N3080);
buf BUF1 (N3168, N3163);
buf BUF1 (N3169, N3164);
buf BUF1 (N3170, N3158);
and AND2 (N3171, N3167, N1068);
and AND3 (N3172, N3160, N2918, N106);
not NOT1 (N3173, N3140);
xor XOR2 (N3174, N3159, N835);
or OR4 (N3175, N3168, N203, N3123, N2819);
and AND2 (N3176, N3169, N2721);
nor NOR3 (N3177, N3176, N1080, N2931);
and AND3 (N3178, N3177, N793, N3050);
or OR3 (N3179, N3178, N1809, N537);
and AND4 (N3180, N3161, N3147, N223, N677);
or OR4 (N3181, N3171, N1637, N775, N2201);
not NOT1 (N3182, N3180);
xor XOR2 (N3183, N3165, N2217);
nor NOR3 (N3184, N3175, N2362, N2516);
buf BUF1 (N3185, N3179);
or OR4 (N3186, N3183, N384, N1312, N2855);
buf BUF1 (N3187, N3184);
and AND3 (N3188, N3186, N1292, N2293);
xor XOR2 (N3189, N3174, N3175);
xor XOR2 (N3190, N3181, N1105);
or OR2 (N3191, N3166, N569);
nor NOR2 (N3192, N3190, N2252);
not NOT1 (N3193, N3185);
and AND2 (N3194, N3189, N484);
or OR4 (N3195, N3173, N1945, N2106, N2792);
buf BUF1 (N3196, N3182);
xor XOR2 (N3197, N3172, N1092);
xor XOR2 (N3198, N3195, N417);
not NOT1 (N3199, N3170);
not NOT1 (N3200, N3196);
not NOT1 (N3201, N3193);
or OR4 (N3202, N3198, N1213, N224, N2356);
not NOT1 (N3203, N3188);
nor NOR3 (N3204, N3199, N747, N3071);
nand NAND2 (N3205, N3192, N647);
nand NAND4 (N3206, N3191, N1610, N355, N287);
not NOT1 (N3207, N3205);
not NOT1 (N3208, N3207);
xor XOR2 (N3209, N3194, N1259);
nor NOR4 (N3210, N3204, N980, N1487, N66);
or OR3 (N3211, N3203, N1873, N2581);
xor XOR2 (N3212, N3187, N2196);
nor NOR4 (N3213, N3208, N2647, N2829, N1716);
nand NAND3 (N3214, N3209, N2789, N636);
nor NOR4 (N3215, N3202, N2958, N613, N2391);
or OR3 (N3216, N3212, N1976, N797);
nor NOR4 (N3217, N3201, N2618, N2346, N2932);
nor NOR3 (N3218, N3211, N455, N1316);
not NOT1 (N3219, N3200);
not NOT1 (N3220, N3214);
buf BUF1 (N3221, N3215);
buf BUF1 (N3222, N3221);
xor XOR2 (N3223, N3222, N1465);
or OR4 (N3224, N3218, N2841, N2971, N1658);
xor XOR2 (N3225, N3223, N2896);
or OR2 (N3226, N3217, N570);
buf BUF1 (N3227, N3197);
nand NAND3 (N3228, N3206, N66, N1717);
buf BUF1 (N3229, N3216);
xor XOR2 (N3230, N3210, N2630);
xor XOR2 (N3231, N3225, N3164);
nor NOR4 (N3232, N3229, N1601, N1124, N2369);
buf BUF1 (N3233, N3220);
nor NOR3 (N3234, N3219, N514, N1095);
buf BUF1 (N3235, N3213);
not NOT1 (N3236, N3235);
nor NOR3 (N3237, N3231, N1834, N254);
xor XOR2 (N3238, N3224, N3193);
and AND2 (N3239, N3238, N2877);
xor XOR2 (N3240, N3228, N245);
not NOT1 (N3241, N3230);
xor XOR2 (N3242, N3240, N2112);
nand NAND2 (N3243, N3233, N2870);
buf BUF1 (N3244, N3226);
nor NOR3 (N3245, N3234, N2040, N1983);
not NOT1 (N3246, N3243);
buf BUF1 (N3247, N3239);
buf BUF1 (N3248, N3232);
nor NOR2 (N3249, N3245, N749);
nor NOR3 (N3250, N3237, N243, N934);
not NOT1 (N3251, N3250);
xor XOR2 (N3252, N3248, N2011);
not NOT1 (N3253, N3241);
not NOT1 (N3254, N3253);
buf BUF1 (N3255, N3244);
not NOT1 (N3256, N3227);
xor XOR2 (N3257, N3255, N2748);
not NOT1 (N3258, N3254);
and AND2 (N3259, N3242, N1911);
buf BUF1 (N3260, N3247);
not NOT1 (N3261, N3256);
or OR2 (N3262, N3246, N143);
and AND2 (N3263, N3251, N1148);
and AND2 (N3264, N3236, N1418);
nand NAND4 (N3265, N3260, N645, N553, N1909);
xor XOR2 (N3266, N3257, N2096);
not NOT1 (N3267, N3259);
or OR4 (N3268, N3267, N1792, N1607, N1770);
and AND4 (N3269, N3252, N1739, N6, N2390);
not NOT1 (N3270, N3264);
and AND4 (N3271, N3270, N2130, N689, N188);
xor XOR2 (N3272, N3261, N2843);
nand NAND4 (N3273, N3266, N1067, N2090, N1587);
buf BUF1 (N3274, N3262);
nand NAND2 (N3275, N3258, N630);
or OR2 (N3276, N3249, N663);
not NOT1 (N3277, N3275);
xor XOR2 (N3278, N3273, N814);
nor NOR3 (N3279, N3277, N2947, N2617);
nand NAND2 (N3280, N3276, N3081);
xor XOR2 (N3281, N3272, N2334);
and AND4 (N3282, N3278, N3251, N368, N543);
xor XOR2 (N3283, N3280, N3242);
xor XOR2 (N3284, N3263, N2383);
or OR4 (N3285, N3271, N1826, N1796, N1073);
not NOT1 (N3286, N3285);
or OR4 (N3287, N3286, N374, N1250, N2022);
or OR4 (N3288, N3281, N1814, N1454, N2726);
or OR4 (N3289, N3274, N2670, N680, N2077);
nor NOR3 (N3290, N3284, N2718, N2532);
and AND4 (N3291, N3288, N2883, N2644, N3145);
or OR4 (N3292, N3289, N1986, N861, N2680);
nor NOR4 (N3293, N3287, N1199, N1312, N2238);
not NOT1 (N3294, N3269);
nand NAND3 (N3295, N3294, N2003, N2452);
nor NOR2 (N3296, N3265, N2701);
not NOT1 (N3297, N3283);
nor NOR4 (N3298, N3296, N2311, N1213, N1526);
nand NAND2 (N3299, N3298, N772);
not NOT1 (N3300, N3291);
nand NAND3 (N3301, N3299, N262, N1407);
not NOT1 (N3302, N3301);
nor NOR3 (N3303, N3282, N1640, N1492);
buf BUF1 (N3304, N3300);
nor NOR2 (N3305, N3295, N1941);
nand NAND4 (N3306, N3303, N2398, N1181, N647);
not NOT1 (N3307, N3305);
xor XOR2 (N3308, N3302, N385);
buf BUF1 (N3309, N3290);
and AND4 (N3310, N3307, N2522, N2342, N2859);
nand NAND3 (N3311, N3304, N1952, N150);
nor NOR2 (N3312, N3292, N348);
nor NOR4 (N3313, N3293, N1305, N566, N213);
buf BUF1 (N3314, N3310);
buf BUF1 (N3315, N3308);
and AND4 (N3316, N3297, N1783, N2174, N851);
and AND2 (N3317, N3314, N1900);
nor NOR3 (N3318, N3315, N2644, N969);
xor XOR2 (N3319, N3306, N163);
xor XOR2 (N3320, N3316, N498);
nor NOR4 (N3321, N3320, N2111, N2683, N1306);
not NOT1 (N3322, N3312);
buf BUF1 (N3323, N3318);
or OR3 (N3324, N3317, N1619, N3239);
xor XOR2 (N3325, N3323, N487);
nor NOR4 (N3326, N3309, N956, N663, N2420);
xor XOR2 (N3327, N3324, N2736);
nand NAND3 (N3328, N3311, N104, N3110);
or OR2 (N3329, N3268, N335);
buf BUF1 (N3330, N3327);
nand NAND2 (N3331, N3330, N2181);
nand NAND3 (N3332, N3319, N537, N2350);
xor XOR2 (N3333, N3321, N1031);
nor NOR3 (N3334, N3328, N2284, N1160);
buf BUF1 (N3335, N3333);
or OR3 (N3336, N3279, N1838, N315);
and AND2 (N3337, N3335, N867);
not NOT1 (N3338, N3313);
and AND3 (N3339, N3338, N3029, N2591);
or OR4 (N3340, N3337, N2630, N492, N2448);
or OR4 (N3341, N3326, N361, N1300, N1038);
nor NOR4 (N3342, N3336, N779, N65, N1874);
and AND4 (N3343, N3331, N1621, N1222, N1179);
nor NOR3 (N3344, N3334, N3244, N1439);
buf BUF1 (N3345, N3339);
buf BUF1 (N3346, N3343);
not NOT1 (N3347, N3342);
nor NOR4 (N3348, N3325, N714, N2746, N2052);
buf BUF1 (N3349, N3329);
and AND3 (N3350, N3332, N1832, N3349);
nor NOR2 (N3351, N1013, N380);
nand NAND3 (N3352, N3348, N1547, N2995);
buf BUF1 (N3353, N3350);
xor XOR2 (N3354, N3341, N1096);
and AND2 (N3355, N3345, N1697);
xor XOR2 (N3356, N3344, N1079);
nand NAND2 (N3357, N3356, N173);
buf BUF1 (N3358, N3355);
nor NOR2 (N3359, N3322, N476);
and AND4 (N3360, N3347, N1111, N1026, N1863);
not NOT1 (N3361, N3360);
or OR2 (N3362, N3361, N3241);
buf BUF1 (N3363, N3351);
nand NAND2 (N3364, N3358, N554);
not NOT1 (N3365, N3363);
nand NAND3 (N3366, N3352, N2983, N2822);
and AND3 (N3367, N3346, N912, N2588);
buf BUF1 (N3368, N3366);
xor XOR2 (N3369, N3354, N1975);
not NOT1 (N3370, N3359);
not NOT1 (N3371, N3353);
or OR2 (N3372, N3357, N2445);
not NOT1 (N3373, N3371);
or OR2 (N3374, N3368, N1729);
buf BUF1 (N3375, N3369);
xor XOR2 (N3376, N3372, N1024);
nor NOR3 (N3377, N3362, N3313, N1623);
nand NAND2 (N3378, N3340, N2135);
xor XOR2 (N3379, N3365, N2254);
nand NAND4 (N3380, N3376, N39, N1307, N1803);
not NOT1 (N3381, N3379);
nor NOR4 (N3382, N3374, N610, N2636, N2540);
buf BUF1 (N3383, N3370);
nand NAND2 (N3384, N3380, N2697);
xor XOR2 (N3385, N3378, N229);
nor NOR3 (N3386, N3381, N897, N2953);
not NOT1 (N3387, N3375);
not NOT1 (N3388, N3385);
nand NAND4 (N3389, N3388, N3249, N3028, N3094);
not NOT1 (N3390, N3382);
buf BUF1 (N3391, N3389);
buf BUF1 (N3392, N3377);
nor NOR3 (N3393, N3391, N1099, N1949);
not NOT1 (N3394, N3390);
xor XOR2 (N3395, N3387, N1102);
buf BUF1 (N3396, N3386);
nor NOR2 (N3397, N3393, N985);
not NOT1 (N3398, N3392);
buf BUF1 (N3399, N3383);
xor XOR2 (N3400, N3384, N2477);
or OR4 (N3401, N3367, N1063, N1912, N1876);
or OR3 (N3402, N3394, N810, N1417);
or OR3 (N3403, N3400, N3383, N3287);
nand NAND4 (N3404, N3364, N1272, N2283, N2405);
or OR3 (N3405, N3404, N3091, N587);
nor NOR2 (N3406, N3373, N2259);
nor NOR2 (N3407, N3396, N2898);
and AND4 (N3408, N3401, N3168, N3130, N810);
nand NAND4 (N3409, N3408, N2719, N1678, N1888);
xor XOR2 (N3410, N3405, N1021);
or OR3 (N3411, N3410, N2708, N1886);
buf BUF1 (N3412, N3411);
xor XOR2 (N3413, N3406, N2047);
or OR3 (N3414, N3402, N2287, N1969);
buf BUF1 (N3415, N3412);
not NOT1 (N3416, N3409);
not NOT1 (N3417, N3413);
nor NOR4 (N3418, N3395, N2700, N89, N2049);
buf BUF1 (N3419, N3418);
nor NOR2 (N3420, N3417, N2413);
not NOT1 (N3421, N3415);
nor NOR2 (N3422, N3419, N2037);
not NOT1 (N3423, N3399);
or OR4 (N3424, N3422, N2014, N1204, N2964);
or OR4 (N3425, N3421, N1505, N2590, N1658);
buf BUF1 (N3426, N3424);
not NOT1 (N3427, N3423);
not NOT1 (N3428, N3416);
buf BUF1 (N3429, N3427);
buf BUF1 (N3430, N3429);
and AND4 (N3431, N3420, N580, N2334, N869);
nand NAND2 (N3432, N3430, N639);
or OR3 (N3433, N3426, N1046, N2189);
xor XOR2 (N3434, N3403, N3098);
or OR4 (N3435, N3414, N3335, N589, N2400);
and AND4 (N3436, N3428, N356, N1669, N770);
buf BUF1 (N3437, N3435);
nand NAND4 (N3438, N3425, N183, N172, N2789);
nor NOR2 (N3439, N3407, N751);
buf BUF1 (N3440, N3432);
xor XOR2 (N3441, N3437, N796);
and AND2 (N3442, N3439, N2761);
xor XOR2 (N3443, N3434, N327);
not NOT1 (N3444, N3433);
and AND4 (N3445, N3397, N2773, N438, N2676);
not NOT1 (N3446, N3444);
nor NOR2 (N3447, N3441, N2114);
or OR3 (N3448, N3442, N624, N2706);
nor NOR4 (N3449, N3446, N3151, N2934, N2067);
buf BUF1 (N3450, N3445);
and AND3 (N3451, N3447, N644, N1032);
buf BUF1 (N3452, N3449);
nand NAND3 (N3453, N3431, N3171, N1767);
xor XOR2 (N3454, N3440, N2721);
nand NAND2 (N3455, N3438, N505);
and AND2 (N3456, N3450, N864);
xor XOR2 (N3457, N3453, N2428);
buf BUF1 (N3458, N3457);
xor XOR2 (N3459, N3398, N2844);
or OR3 (N3460, N3448, N925, N1778);
nor NOR2 (N3461, N3454, N627);
nand NAND4 (N3462, N3461, N2608, N2898, N1600);
not NOT1 (N3463, N3459);
not NOT1 (N3464, N3462);
not NOT1 (N3465, N3455);
xor XOR2 (N3466, N3443, N380);
and AND2 (N3467, N3463, N2134);
or OR2 (N3468, N3464, N1882);
nand NAND2 (N3469, N3456, N2430);
or OR2 (N3470, N3458, N3122);
and AND4 (N3471, N3460, N1007, N2852, N1922);
or OR2 (N3472, N3467, N1203);
or OR4 (N3473, N3451, N1678, N146, N1290);
not NOT1 (N3474, N3472);
not NOT1 (N3475, N3465);
not NOT1 (N3476, N3469);
nor NOR3 (N3477, N3436, N2004, N2263);
buf BUF1 (N3478, N3452);
not NOT1 (N3479, N3470);
nor NOR2 (N3480, N3468, N1232);
nand NAND2 (N3481, N3479, N510);
nor NOR4 (N3482, N3478, N612, N3465, N1601);
or OR4 (N3483, N3480, N1074, N3168, N874);
xor XOR2 (N3484, N3482, N1379);
not NOT1 (N3485, N3474);
xor XOR2 (N3486, N3483, N1428);
not NOT1 (N3487, N3476);
or OR2 (N3488, N3475, N1346);
not NOT1 (N3489, N3481);
or OR4 (N3490, N3473, N943, N1292, N1749);
xor XOR2 (N3491, N3485, N649);
and AND4 (N3492, N3490, N678, N410, N1615);
nor NOR4 (N3493, N3488, N1451, N3157, N649);
nand NAND3 (N3494, N3466, N1219, N215);
xor XOR2 (N3495, N3493, N81);
not NOT1 (N3496, N3491);
buf BUF1 (N3497, N3492);
or OR2 (N3498, N3496, N1014);
not NOT1 (N3499, N3498);
not NOT1 (N3500, N3499);
not NOT1 (N3501, N3495);
and AND3 (N3502, N3494, N3316, N782);
buf BUF1 (N3503, N3500);
xor XOR2 (N3504, N3486, N2363);
nor NOR2 (N3505, N3497, N2230);
nor NOR4 (N3506, N3489, N142, N1451, N3059);
xor XOR2 (N3507, N3487, N3322);
buf BUF1 (N3508, N3484);
nand NAND4 (N3509, N3501, N898, N379, N2065);
not NOT1 (N3510, N3504);
or OR2 (N3511, N3471, N1066);
or OR3 (N3512, N3508, N3168, N365);
nor NOR3 (N3513, N3511, N2806, N2042);
nor NOR2 (N3514, N3477, N2393);
and AND3 (N3515, N3513, N224, N2018);
or OR3 (N3516, N3505, N768, N936);
endmodule