// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N712,N707,N710,N708,N711,N706,N705,N698,N709,N713;

nor NOR2 (N14, N12, N13);
nor NOR2 (N15, N8, N13);
nor NOR3 (N16, N9, N7, N9);
and AND2 (N17, N14, N4);
and AND4 (N18, N3, N9, N1, N12);
or OR2 (N19, N7, N18);
not NOT1 (N20, N10);
buf BUF1 (N21, N5);
or OR3 (N22, N3, N9, N10);
nor NOR2 (N23, N10, N8);
buf BUF1 (N24, N16);
nand NAND2 (N25, N6, N16);
xor XOR2 (N26, N9, N12);
nor NOR2 (N27, N19, N12);
not NOT1 (N28, N21);
nand NAND3 (N29, N15, N17, N10);
and AND2 (N30, N7, N19);
not NOT1 (N31, N20);
not NOT1 (N32, N30);
and AND4 (N33, N25, N15, N9, N21);
nor NOR3 (N34, N22, N17, N24);
not NOT1 (N35, N4);
nand NAND2 (N36, N34, N2);
buf BUF1 (N37, N35);
buf BUF1 (N38, N33);
nand NAND2 (N39, N37, N20);
and AND3 (N40, N29, N25, N9);
or OR3 (N41, N36, N18, N21);
and AND3 (N42, N41, N28, N14);
not NOT1 (N43, N26);
nor NOR4 (N44, N23, N22, N20, N8);
nand NAND2 (N45, N31, N30);
xor XOR2 (N46, N6, N28);
buf BUF1 (N47, N40);
or OR3 (N48, N45, N46, N29);
or OR3 (N49, N37, N18, N30);
buf BUF1 (N50, N48);
and AND2 (N51, N49, N47);
nand NAND3 (N52, N7, N41, N11);
not NOT1 (N53, N42);
and AND3 (N54, N52, N12, N3);
xor XOR2 (N55, N54, N35);
not NOT1 (N56, N43);
buf BUF1 (N57, N44);
nand NAND2 (N58, N51, N9);
buf BUF1 (N59, N56);
or OR2 (N60, N59, N54);
not NOT1 (N61, N27);
xor XOR2 (N62, N38, N35);
nand NAND3 (N63, N39, N58, N7);
nor NOR3 (N64, N30, N6, N33);
xor XOR2 (N65, N57, N36);
and AND4 (N66, N61, N53, N18, N49);
buf BUF1 (N67, N61);
not NOT1 (N68, N66);
xor XOR2 (N69, N55, N43);
and AND3 (N70, N60, N21, N14);
or OR3 (N71, N62, N53, N21);
and AND4 (N72, N71, N62, N69, N62);
and AND4 (N73, N60, N28, N28, N66);
not NOT1 (N74, N72);
xor XOR2 (N75, N70, N60);
or OR2 (N76, N65, N39);
and AND4 (N77, N63, N40, N75, N71);
and AND2 (N78, N39, N24);
or OR3 (N79, N74, N53, N47);
xor XOR2 (N80, N50, N43);
not NOT1 (N81, N78);
nor NOR4 (N82, N77, N1, N11, N29);
and AND4 (N83, N73, N72, N68, N31);
nor NOR2 (N84, N49, N72);
and AND2 (N85, N64, N5);
xor XOR2 (N86, N67, N14);
nand NAND2 (N87, N83, N56);
and AND2 (N88, N87, N32);
and AND3 (N89, N2, N1, N26);
buf BUF1 (N90, N80);
nand NAND4 (N91, N85, N52, N90, N67);
not NOT1 (N92, N13);
or OR4 (N93, N89, N47, N57, N60);
buf BUF1 (N94, N93);
nor NOR3 (N95, N82, N36, N88);
nor NOR2 (N96, N79, N45);
buf BUF1 (N97, N61);
buf BUF1 (N98, N76);
not NOT1 (N99, N97);
buf BUF1 (N100, N81);
or OR3 (N101, N98, N19, N60);
xor XOR2 (N102, N96, N86);
nor NOR4 (N103, N13, N31, N88, N46);
not NOT1 (N104, N102);
nor NOR3 (N105, N104, N99, N14);
nand NAND3 (N106, N6, N73, N94);
and AND3 (N107, N42, N86, N85);
or OR3 (N108, N84, N20, N58);
buf BUF1 (N109, N92);
and AND2 (N110, N91, N66);
not NOT1 (N111, N101);
nor NOR3 (N112, N111, N20, N96);
or OR3 (N113, N103, N48, N81);
or OR3 (N114, N113, N21, N14);
not NOT1 (N115, N109);
and AND3 (N116, N108, N2, N88);
nand NAND4 (N117, N105, N68, N6, N110);
and AND3 (N118, N87, N77, N86);
not NOT1 (N119, N100);
or OR3 (N120, N112, N100, N102);
not NOT1 (N121, N95);
buf BUF1 (N122, N116);
buf BUF1 (N123, N120);
nand NAND4 (N124, N114, N49, N8, N62);
or OR3 (N125, N107, N56, N22);
buf BUF1 (N126, N121);
not NOT1 (N127, N115);
buf BUF1 (N128, N122);
buf BUF1 (N129, N106);
or OR3 (N130, N119, N114, N1);
buf BUF1 (N131, N129);
not NOT1 (N132, N131);
nor NOR3 (N133, N127, N53, N115);
nand NAND2 (N134, N124, N95);
not NOT1 (N135, N134);
or OR3 (N136, N123, N32, N9);
xor XOR2 (N137, N136, N92);
or OR4 (N138, N118, N59, N115, N4);
or OR3 (N139, N128, N101, N35);
and AND4 (N140, N135, N128, N75, N72);
not NOT1 (N141, N125);
buf BUF1 (N142, N139);
and AND4 (N143, N140, N52, N50, N124);
buf BUF1 (N144, N142);
or OR4 (N145, N130, N82, N71, N96);
or OR4 (N146, N145, N97, N23, N127);
or OR3 (N147, N117, N140, N70);
not NOT1 (N148, N132);
xor XOR2 (N149, N148, N60);
and AND4 (N150, N133, N50, N8, N18);
nand NAND4 (N151, N150, N72, N26, N83);
or OR2 (N152, N138, N94);
nor NOR4 (N153, N151, N55, N6, N35);
and AND3 (N154, N141, N33, N103);
and AND3 (N155, N137, N102, N124);
not NOT1 (N156, N149);
nor NOR3 (N157, N153, N7, N135);
xor XOR2 (N158, N154, N20);
nor NOR3 (N159, N147, N96, N82);
not NOT1 (N160, N126);
not NOT1 (N161, N155);
buf BUF1 (N162, N161);
buf BUF1 (N163, N157);
and AND3 (N164, N160, N22, N158);
xor XOR2 (N165, N124, N2);
nand NAND2 (N166, N162, N88);
nor NOR3 (N167, N156, N157, N113);
and AND4 (N168, N143, N9, N152, N95);
xor XOR2 (N169, N119, N60);
and AND3 (N170, N163, N60, N51);
and AND2 (N171, N170, N142);
not NOT1 (N172, N166);
or OR4 (N173, N172, N29, N16, N26);
not NOT1 (N174, N165);
nor NOR4 (N175, N174, N118, N90, N140);
nand NAND4 (N176, N164, N35, N166, N132);
nor NOR3 (N177, N169, N135, N44);
nor NOR4 (N178, N175, N63, N117, N169);
nand NAND4 (N179, N144, N136, N147, N116);
buf BUF1 (N180, N177);
and AND2 (N181, N179, N92);
xor XOR2 (N182, N180, N179);
xor XOR2 (N183, N167, N20);
xor XOR2 (N184, N181, N104);
or OR4 (N185, N168, N180, N174, N81);
or OR3 (N186, N173, N145, N168);
xor XOR2 (N187, N186, N163);
xor XOR2 (N188, N182, N156);
and AND2 (N189, N176, N112);
nor NOR3 (N190, N159, N30, N83);
or OR2 (N191, N188, N167);
xor XOR2 (N192, N187, N94);
and AND2 (N193, N183, N65);
nor NOR2 (N194, N189, N141);
nor NOR3 (N195, N171, N189, N24);
or OR4 (N196, N194, N138, N31, N6);
nand NAND2 (N197, N195, N145);
buf BUF1 (N198, N146);
xor XOR2 (N199, N178, N18);
nor NOR4 (N200, N199, N10, N112, N137);
nor NOR4 (N201, N192, N122, N64, N114);
nor NOR2 (N202, N201, N80);
buf BUF1 (N203, N193);
nor NOR4 (N204, N191, N55, N106, N112);
nor NOR4 (N205, N200, N24, N44, N132);
nand NAND4 (N206, N203, N199, N130, N126);
xor XOR2 (N207, N202, N40);
nor NOR4 (N208, N197, N185, N91, N47);
xor XOR2 (N209, N206, N6);
buf BUF1 (N210, N149);
buf BUF1 (N211, N198);
xor XOR2 (N212, N210, N12);
nor NOR4 (N213, N204, N17, N137, N24);
not NOT1 (N214, N196);
nand NAND2 (N215, N208, N140);
and AND3 (N216, N184, N58, N131);
xor XOR2 (N217, N213, N117);
nor NOR2 (N218, N211, N52);
xor XOR2 (N219, N218, N78);
xor XOR2 (N220, N215, N93);
or OR2 (N221, N190, N175);
not NOT1 (N222, N216);
xor XOR2 (N223, N221, N3);
nor NOR4 (N224, N214, N145, N11, N49);
or OR4 (N225, N205, N13, N146, N89);
not NOT1 (N226, N223);
nand NAND2 (N227, N220, N72);
or OR3 (N228, N226, N85, N114);
xor XOR2 (N229, N227, N210);
nor NOR2 (N230, N228, N157);
xor XOR2 (N231, N217, N20);
nand NAND3 (N232, N229, N202, N185);
nor NOR4 (N233, N224, N50, N221, N142);
nand NAND4 (N234, N222, N65, N191, N99);
not NOT1 (N235, N212);
nor NOR3 (N236, N219, N16, N41);
nand NAND3 (N237, N230, N93, N126);
or OR4 (N238, N209, N59, N20, N26);
nand NAND3 (N239, N236, N79, N211);
nor NOR3 (N240, N239, N148, N46);
xor XOR2 (N241, N207, N116);
xor XOR2 (N242, N240, N216);
nand NAND3 (N243, N237, N155, N161);
or OR3 (N244, N231, N223, N159);
xor XOR2 (N245, N233, N46);
and AND4 (N246, N232, N165, N18, N198);
nand NAND2 (N247, N225, N149);
buf BUF1 (N248, N244);
nor NOR4 (N249, N242, N122, N152, N221);
and AND4 (N250, N246, N148, N213, N198);
nand NAND4 (N251, N238, N87, N174, N131);
not NOT1 (N252, N250);
or OR4 (N253, N247, N105, N194, N83);
nor NOR2 (N254, N253, N84);
or OR2 (N255, N249, N158);
buf BUF1 (N256, N243);
nor NOR2 (N257, N241, N113);
xor XOR2 (N258, N234, N202);
and AND4 (N259, N252, N221, N158, N148);
nor NOR3 (N260, N257, N80, N117);
nand NAND2 (N261, N256, N214);
and AND4 (N262, N254, N54, N1, N73);
xor XOR2 (N263, N245, N185);
xor XOR2 (N264, N255, N181);
and AND2 (N265, N263, N76);
not NOT1 (N266, N251);
and AND3 (N267, N248, N48, N33);
and AND3 (N268, N264, N81, N182);
not NOT1 (N269, N266);
xor XOR2 (N270, N268, N73);
nand NAND2 (N271, N258, N59);
or OR4 (N272, N262, N193, N203, N131);
nand NAND4 (N273, N269, N199, N114, N7);
and AND4 (N274, N259, N212, N19, N96);
buf BUF1 (N275, N265);
nor NOR3 (N276, N273, N10, N214);
nor NOR2 (N277, N271, N156);
not NOT1 (N278, N267);
and AND2 (N279, N270, N133);
or OR2 (N280, N277, N87);
not NOT1 (N281, N260);
xor XOR2 (N282, N279, N185);
buf BUF1 (N283, N272);
or OR3 (N284, N282, N29, N55);
not NOT1 (N285, N274);
or OR2 (N286, N283, N169);
not NOT1 (N287, N285);
and AND3 (N288, N261, N185, N11);
buf BUF1 (N289, N281);
nand NAND3 (N290, N280, N247, N111);
or OR4 (N291, N290, N44, N142, N254);
xor XOR2 (N292, N278, N143);
nor NOR3 (N293, N235, N68, N127);
or OR3 (N294, N284, N151, N111);
xor XOR2 (N295, N294, N93);
not NOT1 (N296, N295);
or OR2 (N297, N276, N240);
nand NAND3 (N298, N292, N20, N278);
or OR3 (N299, N298, N106, N3);
nand NAND3 (N300, N289, N298, N276);
xor XOR2 (N301, N300, N8);
not NOT1 (N302, N297);
xor XOR2 (N303, N286, N45);
and AND3 (N304, N302, N299, N152);
nor NOR4 (N305, N77, N187, N96, N261);
nand NAND4 (N306, N296, N214, N28, N267);
xor XOR2 (N307, N287, N275);
xor XOR2 (N308, N204, N163);
not NOT1 (N309, N306);
xor XOR2 (N310, N305, N38);
xor XOR2 (N311, N304, N161);
buf BUF1 (N312, N293);
buf BUF1 (N313, N312);
buf BUF1 (N314, N303);
nor NOR4 (N315, N314, N48, N71, N295);
not NOT1 (N316, N301);
and AND2 (N317, N308, N38);
nand NAND4 (N318, N310, N88, N228, N239);
nand NAND3 (N319, N318, N11, N158);
and AND3 (N320, N288, N131, N315);
and AND2 (N321, N162, N42);
not NOT1 (N322, N291);
buf BUF1 (N323, N322);
nand NAND3 (N324, N319, N112, N216);
nor NOR4 (N325, N323, N139, N35, N265);
nand NAND3 (N326, N313, N72, N29);
and AND3 (N327, N316, N265, N265);
xor XOR2 (N328, N327, N268);
nand NAND3 (N329, N307, N89, N63);
and AND4 (N330, N326, N262, N142, N318);
xor XOR2 (N331, N325, N26);
buf BUF1 (N332, N330);
not NOT1 (N333, N321);
nand NAND4 (N334, N333, N37, N225, N325);
nor NOR3 (N335, N320, N121, N54);
nand NAND4 (N336, N332, N305, N332, N314);
or OR4 (N337, N334, N325, N237, N257);
or OR3 (N338, N336, N104, N256);
not NOT1 (N339, N311);
or OR2 (N340, N309, N337);
or OR4 (N341, N203, N3, N172, N46);
and AND4 (N342, N340, N25, N75, N102);
not NOT1 (N343, N342);
nor NOR2 (N344, N331, N248);
buf BUF1 (N345, N343);
nand NAND4 (N346, N341, N166, N224, N65);
not NOT1 (N347, N324);
and AND2 (N348, N339, N162);
buf BUF1 (N349, N329);
nand NAND2 (N350, N347, N328);
buf BUF1 (N351, N24);
buf BUF1 (N352, N317);
nand NAND2 (N353, N338, N308);
and AND3 (N354, N345, N65, N336);
nor NOR2 (N355, N344, N251);
or OR3 (N356, N335, N165, N30);
nand NAND4 (N357, N351, N247, N260, N65);
nor NOR4 (N358, N357, N189, N199, N130);
xor XOR2 (N359, N349, N256);
and AND4 (N360, N356, N141, N197, N185);
or OR4 (N361, N346, N320, N127, N267);
or OR3 (N362, N361, N240, N245);
buf BUF1 (N363, N348);
nand NAND2 (N364, N353, N219);
xor XOR2 (N365, N360, N170);
nand NAND3 (N366, N352, N313, N117);
or OR3 (N367, N355, N252, N222);
or OR2 (N368, N367, N71);
nand NAND4 (N369, N365, N230, N189, N60);
buf BUF1 (N370, N366);
buf BUF1 (N371, N364);
or OR2 (N372, N350, N343);
and AND4 (N373, N363, N127, N181, N102);
nor NOR4 (N374, N370, N193, N50, N4);
nor NOR4 (N375, N354, N269, N49, N242);
buf BUF1 (N376, N375);
buf BUF1 (N377, N371);
and AND3 (N378, N359, N135, N30);
or OR2 (N379, N368, N195);
nor NOR3 (N380, N369, N355, N363);
not NOT1 (N381, N372);
not NOT1 (N382, N362);
and AND4 (N383, N374, N187, N62, N229);
buf BUF1 (N384, N379);
xor XOR2 (N385, N381, N155);
nand NAND2 (N386, N376, N155);
nand NAND4 (N387, N373, N101, N241, N192);
nor NOR4 (N388, N384, N304, N242, N71);
or OR2 (N389, N377, N291);
or OR2 (N390, N388, N377);
not NOT1 (N391, N386);
and AND4 (N392, N380, N56, N381, N147);
or OR2 (N393, N387, N35);
not NOT1 (N394, N385);
and AND4 (N395, N389, N333, N162, N371);
not NOT1 (N396, N358);
and AND2 (N397, N391, N85);
nor NOR3 (N398, N390, N308, N148);
or OR4 (N399, N382, N308, N255, N364);
and AND2 (N400, N397, N170);
or OR3 (N401, N396, N151, N294);
xor XOR2 (N402, N400, N393);
and AND3 (N403, N6, N367, N105);
not NOT1 (N404, N398);
or OR4 (N405, N401, N313, N201, N332);
and AND2 (N406, N392, N116);
nand NAND4 (N407, N394, N311, N335, N110);
and AND4 (N408, N405, N35, N186, N243);
nor NOR3 (N409, N395, N387, N28);
xor XOR2 (N410, N406, N170);
and AND3 (N411, N408, N44, N184);
buf BUF1 (N412, N399);
nand NAND2 (N413, N383, N20);
not NOT1 (N414, N412);
nor NOR3 (N415, N409, N197, N372);
not NOT1 (N416, N415);
not NOT1 (N417, N414);
or OR2 (N418, N378, N33);
nand NAND2 (N419, N404, N322);
or OR3 (N420, N416, N235, N254);
and AND4 (N421, N403, N396, N12, N325);
not NOT1 (N422, N411);
nor NOR4 (N423, N419, N243, N360, N27);
or OR2 (N424, N407, N130);
xor XOR2 (N425, N418, N396);
nor NOR2 (N426, N425, N361);
nor NOR2 (N427, N417, N321);
xor XOR2 (N428, N427, N6);
nand NAND3 (N429, N413, N334, N147);
nand NAND3 (N430, N422, N143, N423);
xor XOR2 (N431, N176, N352);
nor NOR3 (N432, N424, N327, N428);
or OR3 (N433, N260, N70, N132);
buf BUF1 (N434, N410);
buf BUF1 (N435, N420);
nand NAND2 (N436, N426, N149);
not NOT1 (N437, N436);
nand NAND4 (N438, N432, N368, N221, N379);
buf BUF1 (N439, N431);
nor NOR3 (N440, N429, N77, N289);
or OR4 (N441, N439, N212, N78, N229);
or OR3 (N442, N421, N283, N62);
nor NOR2 (N443, N438, N352);
and AND4 (N444, N433, N19, N72, N18);
buf BUF1 (N445, N430);
nand NAND4 (N446, N437, N415, N43, N175);
nor NOR3 (N447, N444, N339, N323);
buf BUF1 (N448, N446);
nor NOR4 (N449, N443, N440, N409, N48);
and AND3 (N450, N272, N278, N404);
or OR3 (N451, N449, N16, N184);
nand NAND4 (N452, N448, N126, N398, N334);
nor NOR3 (N453, N445, N247, N35);
or OR2 (N454, N450, N37);
xor XOR2 (N455, N441, N298);
xor XOR2 (N456, N451, N129);
nand NAND2 (N457, N447, N375);
or OR2 (N458, N456, N358);
nor NOR3 (N459, N453, N351, N373);
nor NOR2 (N460, N435, N95);
xor XOR2 (N461, N452, N394);
or OR3 (N462, N434, N414, N12);
nor NOR2 (N463, N460, N19);
nor NOR4 (N464, N402, N422, N381, N160);
nor NOR3 (N465, N457, N440, N393);
and AND3 (N466, N462, N441, N419);
or OR2 (N467, N458, N299);
nor NOR3 (N468, N461, N152, N209);
buf BUF1 (N469, N465);
or OR2 (N470, N459, N63);
or OR4 (N471, N455, N66, N260, N228);
nor NOR2 (N472, N463, N407);
and AND4 (N473, N467, N453, N16, N446);
not NOT1 (N474, N454);
nand NAND4 (N475, N464, N256, N447, N42);
or OR3 (N476, N469, N463, N44);
or OR3 (N477, N472, N146, N60);
buf BUF1 (N478, N471);
xor XOR2 (N479, N470, N131);
nor NOR3 (N480, N477, N66, N91);
buf BUF1 (N481, N466);
or OR2 (N482, N479, N101);
and AND3 (N483, N473, N87, N481);
nor NOR4 (N484, N132, N117, N428, N336);
not NOT1 (N485, N442);
or OR4 (N486, N468, N73, N171, N351);
buf BUF1 (N487, N480);
or OR3 (N488, N486, N423, N225);
not NOT1 (N489, N483);
and AND3 (N490, N488, N337, N406);
nor NOR3 (N491, N484, N116, N377);
and AND3 (N492, N478, N109, N125);
buf BUF1 (N493, N491);
nor NOR4 (N494, N492, N310, N10, N456);
and AND4 (N495, N494, N303, N192, N255);
xor XOR2 (N496, N493, N219);
xor XOR2 (N497, N485, N366);
or OR4 (N498, N489, N128, N158, N223);
or OR2 (N499, N487, N170);
not NOT1 (N500, N499);
nand NAND4 (N501, N476, N240, N438, N88);
nand NAND4 (N502, N501, N64, N265, N219);
buf BUF1 (N503, N482);
xor XOR2 (N504, N496, N369);
nor NOR3 (N505, N502, N301, N153);
nor NOR4 (N506, N503, N33, N455, N368);
xor XOR2 (N507, N506, N187);
xor XOR2 (N508, N495, N465);
not NOT1 (N509, N490);
nor NOR2 (N510, N504, N390);
buf BUF1 (N511, N509);
not NOT1 (N512, N475);
not NOT1 (N513, N498);
not NOT1 (N514, N512);
not NOT1 (N515, N511);
xor XOR2 (N516, N513, N287);
or OR4 (N517, N505, N462, N377, N470);
buf BUF1 (N518, N474);
xor XOR2 (N519, N518, N468);
or OR4 (N520, N497, N486, N132, N91);
and AND3 (N521, N500, N23, N283);
xor XOR2 (N522, N520, N481);
nor NOR2 (N523, N507, N262);
xor XOR2 (N524, N514, N154);
xor XOR2 (N525, N510, N55);
nor NOR2 (N526, N523, N40);
buf BUF1 (N527, N517);
xor XOR2 (N528, N519, N302);
and AND2 (N529, N515, N461);
buf BUF1 (N530, N527);
or OR2 (N531, N528, N108);
buf BUF1 (N532, N516);
not NOT1 (N533, N525);
nand NAND4 (N534, N532, N260, N57, N363);
nand NAND3 (N535, N531, N523, N112);
buf BUF1 (N536, N533);
and AND3 (N537, N522, N350, N242);
or OR4 (N538, N526, N187, N246, N305);
nor NOR4 (N539, N537, N502, N147, N383);
nor NOR2 (N540, N535, N245);
buf BUF1 (N541, N540);
not NOT1 (N542, N529);
nor NOR4 (N543, N536, N70, N273, N90);
buf BUF1 (N544, N534);
nand NAND2 (N545, N538, N356);
buf BUF1 (N546, N543);
or OR4 (N547, N544, N482, N541, N132);
nand NAND3 (N548, N302, N145, N537);
nand NAND4 (N549, N524, N500, N402, N352);
nor NOR4 (N550, N549, N59, N174, N529);
nor NOR2 (N551, N547, N138);
nor NOR4 (N552, N548, N299, N223, N237);
not NOT1 (N553, N539);
xor XOR2 (N554, N508, N383);
nand NAND3 (N555, N521, N415, N413);
buf BUF1 (N556, N545);
nand NAND4 (N557, N555, N413, N419, N318);
or OR3 (N558, N530, N343, N28);
or OR2 (N559, N552, N365);
xor XOR2 (N560, N554, N173);
not NOT1 (N561, N553);
nand NAND2 (N562, N558, N371);
nor NOR3 (N563, N551, N201, N325);
buf BUF1 (N564, N546);
not NOT1 (N565, N562);
not NOT1 (N566, N542);
or OR2 (N567, N563, N392);
xor XOR2 (N568, N559, N239);
buf BUF1 (N569, N564);
buf BUF1 (N570, N565);
or OR4 (N571, N568, N247, N525, N404);
not NOT1 (N572, N567);
xor XOR2 (N573, N569, N268);
nor NOR4 (N574, N556, N534, N569, N569);
not NOT1 (N575, N573);
xor XOR2 (N576, N560, N566);
nand NAND4 (N577, N90, N301, N544, N351);
or OR4 (N578, N561, N214, N400, N181);
nand NAND2 (N579, N574, N339);
buf BUF1 (N580, N576);
xor XOR2 (N581, N550, N464);
xor XOR2 (N582, N579, N530);
nor NOR3 (N583, N577, N299, N351);
xor XOR2 (N584, N571, N522);
or OR2 (N585, N584, N311);
or OR3 (N586, N582, N313, N343);
buf BUF1 (N587, N570);
or OR4 (N588, N585, N515, N21, N299);
nand NAND2 (N589, N580, N546);
xor XOR2 (N590, N587, N76);
and AND2 (N591, N578, N54);
buf BUF1 (N592, N586);
nor NOR4 (N593, N590, N3, N14, N443);
or OR2 (N594, N591, N395);
nor NOR3 (N595, N589, N273, N466);
and AND4 (N596, N583, N188, N79, N110);
nand NAND4 (N597, N581, N548, N550, N556);
nand NAND3 (N598, N575, N358, N227);
nor NOR2 (N599, N572, N464);
nand NAND4 (N600, N588, N186, N313, N354);
not NOT1 (N601, N599);
and AND3 (N602, N600, N349, N531);
nor NOR2 (N603, N596, N9);
buf BUF1 (N604, N593);
nand NAND4 (N605, N594, N12, N94, N476);
nor NOR4 (N606, N602, N430, N410, N73);
nor NOR4 (N607, N603, N434, N78, N152);
nor NOR4 (N608, N597, N543, N469, N523);
nand NAND3 (N609, N604, N389, N204);
or OR4 (N610, N601, N10, N72, N38);
buf BUF1 (N611, N592);
xor XOR2 (N612, N598, N450);
or OR2 (N613, N557, N216);
and AND3 (N614, N607, N517, N298);
not NOT1 (N615, N610);
not NOT1 (N616, N605);
or OR2 (N617, N616, N411);
nor NOR2 (N618, N615, N253);
not NOT1 (N619, N606);
nor NOR2 (N620, N609, N584);
or OR4 (N621, N595, N556, N31, N488);
buf BUF1 (N622, N614);
nor NOR3 (N623, N613, N408, N484);
xor XOR2 (N624, N618, N590);
not NOT1 (N625, N623);
xor XOR2 (N626, N611, N93);
buf BUF1 (N627, N626);
and AND4 (N628, N624, N305, N35, N349);
not NOT1 (N629, N619);
nand NAND3 (N630, N612, N241, N504);
xor XOR2 (N631, N620, N540);
nand NAND3 (N632, N630, N224, N37);
xor XOR2 (N633, N621, N179);
or OR3 (N634, N633, N145, N385);
nand NAND2 (N635, N622, N157);
nor NOR4 (N636, N608, N292, N477, N615);
buf BUF1 (N637, N629);
or OR2 (N638, N637, N578);
and AND2 (N639, N635, N322);
xor XOR2 (N640, N638, N589);
buf BUF1 (N641, N631);
buf BUF1 (N642, N617);
xor XOR2 (N643, N628, N546);
not NOT1 (N644, N636);
nand NAND2 (N645, N640, N386);
nand NAND4 (N646, N627, N510, N87, N115);
xor XOR2 (N647, N645, N325);
and AND2 (N648, N643, N375);
and AND3 (N649, N641, N27, N23);
nor NOR3 (N650, N632, N582, N138);
and AND4 (N651, N644, N279, N79, N200);
xor XOR2 (N652, N642, N317);
or OR2 (N653, N639, N256);
xor XOR2 (N654, N653, N649);
buf BUF1 (N655, N150);
nor NOR2 (N656, N646, N153);
buf BUF1 (N657, N634);
or OR2 (N658, N647, N506);
xor XOR2 (N659, N655, N464);
nor NOR2 (N660, N657, N442);
not NOT1 (N661, N654);
not NOT1 (N662, N658);
xor XOR2 (N663, N625, N342);
buf BUF1 (N664, N650);
not NOT1 (N665, N651);
nand NAND2 (N666, N663, N166);
nor NOR2 (N667, N652, N627);
not NOT1 (N668, N661);
not NOT1 (N669, N668);
xor XOR2 (N670, N656, N540);
and AND3 (N671, N669, N132, N171);
nor NOR4 (N672, N666, N593, N119, N24);
xor XOR2 (N673, N659, N63);
xor XOR2 (N674, N667, N141);
nor NOR2 (N675, N660, N287);
or OR3 (N676, N672, N148, N188);
nand NAND2 (N677, N671, N615);
nor NOR3 (N678, N648, N214, N479);
nand NAND2 (N679, N664, N137);
buf BUF1 (N680, N677);
nand NAND4 (N681, N680, N318, N82, N655);
buf BUF1 (N682, N670);
and AND2 (N683, N662, N511);
nand NAND2 (N684, N673, N263);
buf BUF1 (N685, N684);
buf BUF1 (N686, N665);
or OR2 (N687, N679, N606);
xor XOR2 (N688, N676, N73);
nor NOR4 (N689, N688, N227, N142, N634);
and AND2 (N690, N689, N620);
xor XOR2 (N691, N687, N222);
buf BUF1 (N692, N690);
and AND4 (N693, N674, N66, N470, N652);
xor XOR2 (N694, N693, N60);
or OR3 (N695, N681, N180, N626);
not NOT1 (N696, N695);
xor XOR2 (N697, N686, N411);
nand NAND4 (N698, N694, N439, N626, N30);
nand NAND4 (N699, N685, N218, N238, N156);
and AND2 (N700, N683, N94);
buf BUF1 (N701, N691);
buf BUF1 (N702, N696);
xor XOR2 (N703, N697, N15);
xor XOR2 (N704, N703, N278);
nand NAND4 (N705, N678, N690, N496, N684);
nand NAND4 (N706, N702, N496, N365, N490);
not NOT1 (N707, N675);
xor XOR2 (N708, N682, N535);
or OR2 (N709, N704, N132);
xor XOR2 (N710, N701, N113);
nor NOR2 (N711, N692, N217);
or OR3 (N712, N699, N305, N643);
buf BUF1 (N713, N700);
endmodule