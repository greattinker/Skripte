// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N12810,N12811,N12807,N12812,N12796,N12813,N12805,N12814,N12806,N12815;

not NOT1 (N16, N12);
and AND3 (N17, N14, N5, N9);
not NOT1 (N18, N15);
and AND3 (N19, N10, N13, N14);
nand NAND2 (N20, N10, N4);
nand NAND3 (N21, N20, N16, N2);
buf BUF1 (N22, N9);
buf BUF1 (N23, N6);
buf BUF1 (N24, N2);
not NOT1 (N25, N9);
nor NOR3 (N26, N3, N12, N19);
xor XOR2 (N27, N14, N9);
or OR3 (N28, N4, N7, N1);
and AND2 (N29, N17, N14);
not NOT1 (N30, N29);
nand NAND4 (N31, N18, N17, N27, N29);
not NOT1 (N32, N16);
not NOT1 (N33, N30);
or OR2 (N34, N26, N33);
or OR3 (N35, N19, N30, N8);
nand NAND3 (N36, N25, N28, N28);
or OR3 (N37, N15, N7, N15);
xor XOR2 (N38, N21, N19);
nand NAND4 (N39, N23, N11, N8, N6);
buf BUF1 (N40, N37);
buf BUF1 (N41, N31);
xor XOR2 (N42, N34, N19);
not NOT1 (N43, N40);
and AND2 (N44, N35, N20);
xor XOR2 (N45, N32, N30);
and AND2 (N46, N22, N17);
nand NAND3 (N47, N44, N14, N30);
or OR3 (N48, N46, N2, N46);
not NOT1 (N49, N36);
and AND2 (N50, N42, N44);
not NOT1 (N51, N24);
buf BUF1 (N52, N48);
and AND2 (N53, N49, N10);
nor NOR2 (N54, N50, N27);
buf BUF1 (N55, N41);
not NOT1 (N56, N39);
xor XOR2 (N57, N43, N41);
xor XOR2 (N58, N53, N32);
nand NAND2 (N59, N55, N7);
xor XOR2 (N60, N59, N12);
buf BUF1 (N61, N51);
xor XOR2 (N62, N38, N8);
and AND4 (N63, N62, N47, N40, N35);
xor XOR2 (N64, N32, N25);
not NOT1 (N65, N64);
and AND3 (N66, N60, N24, N46);
or OR4 (N67, N54, N4, N61, N5);
xor XOR2 (N68, N61, N41);
nand NAND4 (N69, N66, N33, N67, N41);
nor NOR2 (N70, N44, N23);
or OR2 (N71, N56, N64);
xor XOR2 (N72, N45, N12);
or OR2 (N73, N71, N52);
not NOT1 (N74, N62);
buf BUF1 (N75, N69);
not NOT1 (N76, N57);
xor XOR2 (N77, N68, N39);
not NOT1 (N78, N58);
nor NOR3 (N79, N72, N75, N32);
nor NOR3 (N80, N15, N49, N8);
and AND2 (N81, N74, N38);
and AND4 (N82, N73, N77, N43, N62);
xor XOR2 (N83, N30, N79);
and AND2 (N84, N42, N52);
buf BUF1 (N85, N82);
not NOT1 (N86, N85);
nor NOR2 (N87, N78, N61);
or OR3 (N88, N76, N38, N81);
nand NAND2 (N89, N9, N38);
not NOT1 (N90, N70);
buf BUF1 (N91, N84);
buf BUF1 (N92, N80);
or OR3 (N93, N65, N57, N57);
buf BUF1 (N94, N91);
xor XOR2 (N95, N93, N84);
and AND4 (N96, N88, N75, N31, N42);
nor NOR3 (N97, N63, N12, N66);
buf BUF1 (N98, N94);
or OR2 (N99, N92, N17);
buf BUF1 (N100, N98);
buf BUF1 (N101, N90);
buf BUF1 (N102, N96);
and AND4 (N103, N102, N84, N8, N44);
or OR2 (N104, N103, N63);
and AND4 (N105, N97, N11, N43, N40);
nor NOR4 (N106, N101, N61, N90, N34);
xor XOR2 (N107, N83, N1);
buf BUF1 (N108, N104);
xor XOR2 (N109, N86, N80);
nor NOR4 (N110, N87, N102, N23, N109);
buf BUF1 (N111, N74);
or OR2 (N112, N111, N53);
buf BUF1 (N113, N107);
and AND2 (N114, N95, N76);
buf BUF1 (N115, N108);
nand NAND4 (N116, N106, N38, N73, N61);
nand NAND3 (N117, N112, N49, N72);
and AND2 (N118, N113, N88);
xor XOR2 (N119, N89, N45);
and AND3 (N120, N118, N28, N103);
and AND3 (N121, N114, N53, N22);
not NOT1 (N122, N119);
nor NOR4 (N123, N116, N32, N67, N74);
nand NAND4 (N124, N123, N21, N42, N25);
buf BUF1 (N125, N120);
xor XOR2 (N126, N121, N28);
nand NAND4 (N127, N110, N102, N104, N83);
and AND2 (N128, N124, N22);
buf BUF1 (N129, N99);
nor NOR2 (N130, N105, N117);
and AND2 (N131, N86, N84);
and AND3 (N132, N130, N47, N32);
and AND2 (N133, N122, N76);
buf BUF1 (N134, N129);
nand NAND4 (N135, N126, N19, N42, N118);
nand NAND4 (N136, N125, N32, N73, N124);
xor XOR2 (N137, N136, N107);
or OR2 (N138, N131, N2);
xor XOR2 (N139, N128, N35);
nand NAND4 (N140, N138, N122, N108, N7);
nor NOR4 (N141, N133, N99, N72, N53);
or OR2 (N142, N132, N100);
not NOT1 (N143, N20);
not NOT1 (N144, N140);
and AND4 (N145, N143, N100, N30, N99);
xor XOR2 (N146, N139, N24);
buf BUF1 (N147, N144);
nand NAND4 (N148, N134, N90, N76, N9);
or OR3 (N149, N135, N32, N8);
or OR3 (N150, N115, N70, N14);
or OR4 (N151, N148, N47, N92, N137);
nor NOR3 (N152, N33, N92, N97);
nand NAND3 (N153, N150, N136, N44);
xor XOR2 (N154, N141, N106);
and AND4 (N155, N147, N35, N17, N129);
xor XOR2 (N156, N127, N6);
not NOT1 (N157, N154);
nand NAND3 (N158, N157, N124, N116);
xor XOR2 (N159, N156, N128);
nand NAND4 (N160, N149, N94, N44, N68);
and AND2 (N161, N151, N17);
xor XOR2 (N162, N161, N56);
or OR3 (N163, N158, N105, N132);
nand NAND2 (N164, N153, N121);
and AND4 (N165, N162, N110, N134, N50);
buf BUF1 (N166, N142);
not NOT1 (N167, N155);
nand NAND2 (N168, N146, N55);
or OR4 (N169, N152, N63, N9, N152);
or OR3 (N170, N164, N60, N24);
or OR4 (N171, N166, N25, N125, N46);
xor XOR2 (N172, N159, N40);
or OR4 (N173, N163, N134, N105, N135);
buf BUF1 (N174, N165);
nor NOR2 (N175, N169, N170);
or OR2 (N176, N43, N162);
buf BUF1 (N177, N168);
nand NAND4 (N178, N175, N86, N7, N164);
and AND4 (N179, N167, N77, N58, N133);
nand NAND4 (N180, N172, N68, N95, N139);
xor XOR2 (N181, N145, N150);
and AND2 (N182, N160, N166);
nand NAND4 (N183, N174, N48, N85, N166);
nor NOR4 (N184, N173, N53, N179, N17);
xor XOR2 (N185, N159, N29);
nand NAND4 (N186, N177, N22, N25, N151);
and AND4 (N187, N180, N184, N177, N186);
xor XOR2 (N188, N10, N26);
or OR3 (N189, N19, N28, N138);
buf BUF1 (N190, N187);
not NOT1 (N191, N178);
or OR2 (N192, N182, N12);
nand NAND3 (N193, N192, N157, N131);
nor NOR4 (N194, N191, N40, N44, N77);
xor XOR2 (N195, N171, N80);
or OR4 (N196, N183, N115, N58, N62);
nor NOR4 (N197, N193, N2, N9, N115);
xor XOR2 (N198, N185, N157);
and AND2 (N199, N176, N183);
or OR2 (N200, N194, N105);
nor NOR3 (N201, N200, N44, N169);
and AND4 (N202, N181, N44, N53, N23);
buf BUF1 (N203, N189);
buf BUF1 (N204, N201);
not NOT1 (N205, N197);
nor NOR3 (N206, N190, N4, N55);
nor NOR3 (N207, N195, N192, N187);
buf BUF1 (N208, N188);
or OR2 (N209, N207, N6);
nand NAND2 (N210, N206, N45);
or OR2 (N211, N196, N192);
and AND2 (N212, N198, N202);
buf BUF1 (N213, N158);
and AND4 (N214, N208, N206, N210, N89);
or OR2 (N215, N75, N115);
not NOT1 (N216, N214);
and AND4 (N217, N212, N169, N163, N82);
xor XOR2 (N218, N217, N198);
or OR2 (N219, N205, N144);
or OR4 (N220, N218, N10, N102, N24);
not NOT1 (N221, N211);
xor XOR2 (N222, N209, N149);
buf BUF1 (N223, N222);
nor NOR2 (N224, N203, N125);
nor NOR4 (N225, N220, N168, N156, N125);
xor XOR2 (N226, N215, N191);
xor XOR2 (N227, N199, N25);
nor NOR2 (N228, N224, N212);
not NOT1 (N229, N216);
xor XOR2 (N230, N227, N172);
nor NOR3 (N231, N221, N107, N23);
nand NAND2 (N232, N230, N6);
xor XOR2 (N233, N219, N192);
nand NAND4 (N234, N229, N219, N11, N202);
nand NAND3 (N235, N226, N132, N177);
xor XOR2 (N236, N213, N50);
xor XOR2 (N237, N234, N143);
xor XOR2 (N238, N236, N220);
xor XOR2 (N239, N225, N156);
buf BUF1 (N240, N233);
and AND4 (N241, N240, N22, N27, N239);
buf BUF1 (N242, N86);
nor NOR3 (N243, N223, N169, N96);
or OR4 (N244, N235, N146, N66, N105);
and AND4 (N245, N237, N20, N191, N217);
not NOT1 (N246, N241);
and AND3 (N247, N246, N159, N28);
buf BUF1 (N248, N231);
buf BUF1 (N249, N245);
and AND2 (N250, N204, N49);
nand NAND4 (N251, N250, N167, N176, N180);
nand NAND2 (N252, N232, N102);
nand NAND3 (N253, N243, N175, N165);
buf BUF1 (N254, N238);
or OR3 (N255, N251, N154, N90);
not NOT1 (N256, N255);
buf BUF1 (N257, N252);
xor XOR2 (N258, N253, N147);
xor XOR2 (N259, N249, N107);
or OR2 (N260, N259, N10);
nor NOR2 (N261, N256, N19);
buf BUF1 (N262, N258);
or OR2 (N263, N242, N116);
nand NAND2 (N264, N263, N166);
nand NAND2 (N265, N248, N240);
and AND3 (N266, N247, N78, N86);
xor XOR2 (N267, N254, N93);
or OR4 (N268, N257, N238, N92, N236);
and AND4 (N269, N267, N217, N220, N67);
buf BUF1 (N270, N261);
nor NOR4 (N271, N269, N175, N85, N4);
or OR4 (N272, N264, N30, N172, N160);
nor NOR4 (N273, N271, N176, N18, N217);
buf BUF1 (N274, N262);
or OR3 (N275, N265, N29, N203);
buf BUF1 (N276, N270);
or OR2 (N277, N266, N163);
nand NAND2 (N278, N275, N128);
not NOT1 (N279, N260);
or OR4 (N280, N278, N165, N55, N223);
and AND3 (N281, N244, N243, N101);
nand NAND4 (N282, N276, N135, N224, N200);
or OR2 (N283, N280, N244);
xor XOR2 (N284, N279, N237);
and AND3 (N285, N277, N198, N184);
nand NAND3 (N286, N284, N70, N148);
and AND2 (N287, N274, N264);
not NOT1 (N288, N287);
and AND3 (N289, N286, N148, N4);
and AND2 (N290, N273, N118);
or OR3 (N291, N272, N215, N172);
xor XOR2 (N292, N228, N19);
nor NOR3 (N293, N288, N134, N22);
nand NAND3 (N294, N285, N222, N36);
xor XOR2 (N295, N283, N45);
nor NOR3 (N296, N290, N1, N46);
nor NOR3 (N297, N292, N88, N136);
xor XOR2 (N298, N294, N192);
nand NAND4 (N299, N293, N77, N59, N282);
nor NOR4 (N300, N58, N128, N18, N230);
not NOT1 (N301, N268);
or OR4 (N302, N299, N88, N183, N167);
or OR4 (N303, N289, N161, N151, N53);
xor XOR2 (N304, N297, N86);
nand NAND3 (N305, N296, N205, N25);
nand NAND3 (N306, N295, N56, N268);
or OR2 (N307, N306, N64);
and AND4 (N308, N303, N109, N177, N13);
xor XOR2 (N309, N308, N75);
nor NOR3 (N310, N281, N72, N105);
xor XOR2 (N311, N298, N38);
and AND3 (N312, N304, N276, N206);
xor XOR2 (N313, N305, N129);
nand NAND4 (N314, N310, N290, N150, N275);
and AND3 (N315, N302, N83, N67);
not NOT1 (N316, N309);
nor NOR4 (N317, N312, N211, N119, N259);
and AND4 (N318, N291, N216, N89, N269);
not NOT1 (N319, N317);
nor NOR3 (N320, N316, N116, N220);
and AND4 (N321, N313, N237, N61, N3);
and AND2 (N322, N311, N41);
or OR3 (N323, N300, N25, N126);
buf BUF1 (N324, N307);
or OR4 (N325, N321, N226, N43, N309);
nor NOR4 (N326, N323, N75, N294, N195);
xor XOR2 (N327, N325, N10);
or OR3 (N328, N318, N161, N199);
nor NOR3 (N329, N327, N208, N183);
nor NOR2 (N330, N315, N87);
buf BUF1 (N331, N319);
nand NAND2 (N332, N330, N202);
buf BUF1 (N333, N320);
not NOT1 (N334, N331);
xor XOR2 (N335, N334, N320);
or OR3 (N336, N333, N269, N95);
or OR3 (N337, N335, N25, N200);
buf BUF1 (N338, N326);
buf BUF1 (N339, N314);
buf BUF1 (N340, N336);
or OR4 (N341, N340, N144, N110, N175);
nor NOR4 (N342, N329, N216, N203, N191);
nand NAND3 (N343, N301, N293, N243);
xor XOR2 (N344, N337, N275);
not NOT1 (N345, N338);
buf BUF1 (N346, N324);
xor XOR2 (N347, N344, N310);
buf BUF1 (N348, N342);
not NOT1 (N349, N328);
and AND3 (N350, N348, N249, N51);
and AND4 (N351, N350, N69, N38, N62);
nor NOR4 (N352, N322, N15, N140, N255);
xor XOR2 (N353, N346, N79);
and AND2 (N354, N353, N95);
buf BUF1 (N355, N354);
not NOT1 (N356, N343);
not NOT1 (N357, N332);
or OR2 (N358, N347, N233);
or OR3 (N359, N349, N352, N330);
xor XOR2 (N360, N201, N221);
or OR4 (N361, N358, N204, N43, N159);
nor NOR3 (N362, N341, N252, N12);
nor NOR3 (N363, N360, N68, N84);
not NOT1 (N364, N363);
and AND4 (N365, N351, N122, N200, N150);
not NOT1 (N366, N361);
nand NAND3 (N367, N366, N307, N75);
nor NOR4 (N368, N365, N312, N205, N89);
or OR2 (N369, N367, N182);
buf BUF1 (N370, N369);
xor XOR2 (N371, N357, N9);
nand NAND4 (N372, N339, N326, N64, N324);
and AND2 (N373, N371, N112);
and AND2 (N374, N362, N301);
not NOT1 (N375, N368);
xor XOR2 (N376, N345, N273);
xor XOR2 (N377, N374, N278);
nand NAND2 (N378, N376, N222);
nand NAND4 (N379, N375, N40, N361, N354);
not NOT1 (N380, N379);
and AND2 (N381, N378, N26);
nor NOR3 (N382, N359, N372, N219);
buf BUF1 (N383, N45);
nor NOR4 (N384, N382, N137, N16, N248);
and AND3 (N385, N364, N159, N89);
nand NAND3 (N386, N370, N305, N57);
buf BUF1 (N387, N385);
and AND3 (N388, N377, N162, N45);
xor XOR2 (N389, N380, N132);
xor XOR2 (N390, N387, N259);
nor NOR3 (N391, N383, N25, N210);
nand NAND2 (N392, N388, N75);
and AND2 (N393, N391, N67);
nand NAND3 (N394, N355, N61, N159);
nand NAND2 (N395, N356, N161);
or OR2 (N396, N394, N56);
not NOT1 (N397, N373);
xor XOR2 (N398, N393, N151);
buf BUF1 (N399, N386);
or OR2 (N400, N396, N291);
not NOT1 (N401, N389);
nor NOR4 (N402, N400, N393, N83, N241);
not NOT1 (N403, N399);
nand NAND3 (N404, N392, N170, N250);
not NOT1 (N405, N404);
and AND2 (N406, N381, N85);
and AND2 (N407, N395, N285);
and AND2 (N408, N403, N304);
xor XOR2 (N409, N407, N2);
xor XOR2 (N410, N408, N218);
nor NOR4 (N411, N405, N15, N176, N149);
nand NAND3 (N412, N384, N60, N58);
buf BUF1 (N413, N410);
or OR2 (N414, N409, N73);
xor XOR2 (N415, N401, N4);
or OR4 (N416, N412, N9, N63, N14);
buf BUF1 (N417, N397);
nand NAND3 (N418, N414, N285, N383);
not NOT1 (N419, N398);
and AND3 (N420, N390, N21, N73);
nor NOR3 (N421, N411, N279, N253);
buf BUF1 (N422, N420);
xor XOR2 (N423, N421, N13);
xor XOR2 (N424, N419, N206);
xor XOR2 (N425, N422, N173);
and AND2 (N426, N415, N189);
nand NAND2 (N427, N416, N323);
not NOT1 (N428, N425);
or OR3 (N429, N427, N156, N305);
and AND2 (N430, N406, N235);
buf BUF1 (N431, N402);
or OR2 (N432, N424, N152);
nand NAND3 (N433, N431, N402, N219);
xor XOR2 (N434, N430, N366);
not NOT1 (N435, N426);
nor NOR4 (N436, N433, N60, N432, N328);
and AND2 (N437, N378, N29);
nand NAND3 (N438, N437, N45, N118);
nor NOR3 (N439, N435, N197, N426);
not NOT1 (N440, N438);
and AND2 (N441, N423, N289);
or OR2 (N442, N439, N225);
nand NAND3 (N443, N436, N280, N114);
or OR2 (N444, N434, N107);
nand NAND2 (N445, N441, N301);
nand NAND2 (N446, N428, N96);
nand NAND3 (N447, N445, N282, N8);
xor XOR2 (N448, N444, N406);
not NOT1 (N449, N413);
and AND4 (N450, N429, N131, N275, N81);
xor XOR2 (N451, N418, N42);
buf BUF1 (N452, N417);
nor NOR4 (N453, N449, N49, N89, N249);
xor XOR2 (N454, N440, N71);
not NOT1 (N455, N443);
and AND2 (N456, N442, N301);
xor XOR2 (N457, N455, N81);
not NOT1 (N458, N446);
nand NAND2 (N459, N448, N118);
not NOT1 (N460, N459);
buf BUF1 (N461, N460);
not NOT1 (N462, N450);
or OR3 (N463, N461, N171, N275);
or OR3 (N464, N452, N446, N190);
or OR2 (N465, N454, N195);
buf BUF1 (N466, N456);
nor NOR3 (N467, N464, N34, N243);
nor NOR4 (N468, N466, N351, N39, N154);
nand NAND3 (N469, N453, N204, N386);
buf BUF1 (N470, N458);
nand NAND3 (N471, N457, N120, N170);
buf BUF1 (N472, N470);
or OR3 (N473, N472, N422, N287);
nand NAND2 (N474, N468, N155);
nor NOR3 (N475, N471, N305, N338);
not NOT1 (N476, N462);
or OR3 (N477, N473, N415, N53);
and AND2 (N478, N477, N397);
not NOT1 (N479, N447);
xor XOR2 (N480, N451, N305);
or OR2 (N481, N463, N185);
and AND4 (N482, N481, N184, N302, N314);
nand NAND3 (N483, N476, N300, N28);
xor XOR2 (N484, N469, N50);
nor NOR3 (N485, N465, N279, N335);
buf BUF1 (N486, N482);
not NOT1 (N487, N484);
buf BUF1 (N488, N480);
nor NOR4 (N489, N487, N352, N67, N474);
not NOT1 (N490, N103);
xor XOR2 (N491, N490, N92);
nor NOR4 (N492, N479, N286, N402, N482);
nor NOR2 (N493, N486, N162);
nor NOR2 (N494, N483, N417);
nor NOR4 (N495, N478, N114, N104, N77);
or OR2 (N496, N492, N176);
and AND3 (N497, N491, N51, N425);
buf BUF1 (N498, N467);
nand NAND4 (N499, N497, N460, N428, N405);
not NOT1 (N500, N498);
xor XOR2 (N501, N489, N27);
not NOT1 (N502, N475);
nor NOR2 (N503, N485, N145);
not NOT1 (N504, N493);
and AND2 (N505, N500, N401);
xor XOR2 (N506, N505, N167);
buf BUF1 (N507, N503);
buf BUF1 (N508, N494);
or OR4 (N509, N502, N491, N220, N408);
and AND3 (N510, N495, N54, N454);
nand NAND3 (N511, N510, N249, N292);
buf BUF1 (N512, N508);
and AND2 (N513, N507, N409);
nand NAND3 (N514, N509, N476, N113);
nor NOR4 (N515, N511, N347, N489, N233);
xor XOR2 (N516, N496, N32);
nand NAND2 (N517, N516, N461);
and AND2 (N518, N506, N434);
buf BUF1 (N519, N515);
nor NOR2 (N520, N501, N181);
not NOT1 (N521, N499);
xor XOR2 (N522, N518, N367);
nand NAND4 (N523, N512, N202, N63, N342);
or OR2 (N524, N488, N263);
nand NAND2 (N525, N524, N216);
or OR3 (N526, N523, N206, N504);
buf BUF1 (N527, N434);
nor NOR2 (N528, N526, N172);
and AND3 (N529, N525, N456, N68);
and AND4 (N530, N517, N12, N240, N347);
nor NOR2 (N531, N529, N358);
and AND2 (N532, N521, N263);
or OR4 (N533, N513, N23, N425, N275);
and AND3 (N534, N514, N145, N249);
or OR3 (N535, N533, N449, N190);
or OR3 (N536, N528, N141, N143);
buf BUF1 (N537, N531);
not NOT1 (N538, N520);
nor NOR4 (N539, N530, N123, N217, N187);
not NOT1 (N540, N538);
nand NAND4 (N541, N527, N270, N118, N366);
not NOT1 (N542, N537);
nand NAND4 (N543, N540, N423, N212, N421);
and AND3 (N544, N534, N175, N303);
nor NOR4 (N545, N532, N247, N191, N195);
not NOT1 (N546, N544);
nor NOR4 (N547, N535, N66, N498, N542);
nand NAND2 (N548, N451, N267);
or OR2 (N549, N548, N69);
buf BUF1 (N550, N547);
and AND3 (N551, N546, N447, N257);
nor NOR2 (N552, N543, N39);
nor NOR3 (N553, N539, N255, N61);
nand NAND2 (N554, N545, N187);
and AND3 (N555, N536, N147, N83);
not NOT1 (N556, N550);
and AND3 (N557, N554, N149, N50);
xor XOR2 (N558, N556, N224);
xor XOR2 (N559, N551, N7);
or OR2 (N560, N559, N351);
xor XOR2 (N561, N555, N308);
nor NOR4 (N562, N541, N412, N265, N494);
or OR2 (N563, N558, N542);
xor XOR2 (N564, N560, N222);
and AND2 (N565, N561, N308);
and AND2 (N566, N563, N69);
or OR2 (N567, N562, N353);
and AND3 (N568, N564, N152, N195);
nor NOR4 (N569, N567, N112, N214, N383);
or OR2 (N570, N522, N318);
and AND2 (N571, N553, N42);
and AND3 (N572, N519, N416, N366);
or OR2 (N573, N569, N255);
buf BUF1 (N574, N566);
nor NOR4 (N575, N549, N209, N479, N528);
xor XOR2 (N576, N570, N98);
or OR2 (N577, N574, N507);
or OR4 (N578, N577, N496, N180, N304);
and AND3 (N579, N573, N230, N373);
and AND4 (N580, N579, N548, N484, N410);
buf BUF1 (N581, N552);
or OR4 (N582, N576, N520, N30, N76);
xor XOR2 (N583, N572, N276);
nor NOR2 (N584, N568, N345);
and AND3 (N585, N557, N152, N79);
nand NAND3 (N586, N581, N151, N372);
and AND2 (N587, N582, N430);
nand NAND4 (N588, N580, N317, N111, N327);
nor NOR4 (N589, N571, N464, N191, N465);
and AND3 (N590, N589, N419, N188);
not NOT1 (N591, N584);
nor NOR3 (N592, N586, N348, N478);
and AND4 (N593, N575, N451, N367, N183);
nand NAND4 (N594, N585, N342, N28, N239);
and AND2 (N595, N583, N374);
or OR4 (N596, N594, N571, N576, N200);
nand NAND2 (N597, N588, N198);
nand NAND2 (N598, N587, N177);
not NOT1 (N599, N592);
nand NAND2 (N600, N597, N459);
nand NAND4 (N601, N591, N45, N264, N383);
and AND2 (N602, N599, N179);
and AND2 (N603, N595, N240);
nor NOR2 (N604, N578, N115);
and AND3 (N605, N604, N445, N215);
xor XOR2 (N606, N590, N104);
nor NOR4 (N607, N605, N58, N83, N253);
nor NOR3 (N608, N601, N152, N218);
and AND2 (N609, N607, N65);
nand NAND3 (N610, N603, N202, N597);
buf BUF1 (N611, N609);
xor XOR2 (N612, N593, N199);
xor XOR2 (N613, N602, N393);
nand NAND4 (N614, N613, N419, N200, N589);
nand NAND2 (N615, N600, N226);
nand NAND4 (N616, N596, N325, N605, N53);
and AND2 (N617, N606, N350);
and AND2 (N618, N616, N209);
or OR2 (N619, N618, N220);
nor NOR3 (N620, N608, N134, N243);
buf BUF1 (N621, N612);
nand NAND4 (N622, N617, N328, N577, N609);
and AND2 (N623, N614, N234);
nand NAND3 (N624, N610, N165, N198);
nand NAND3 (N625, N624, N83, N141);
buf BUF1 (N626, N620);
xor XOR2 (N627, N626, N278);
nand NAND2 (N628, N611, N57);
nand NAND4 (N629, N622, N389, N480, N468);
xor XOR2 (N630, N623, N527);
xor XOR2 (N631, N628, N10);
xor XOR2 (N632, N627, N265);
or OR3 (N633, N565, N432, N603);
nand NAND4 (N634, N633, N310, N562, N382);
buf BUF1 (N635, N621);
buf BUF1 (N636, N634);
not NOT1 (N637, N630);
buf BUF1 (N638, N625);
nor NOR3 (N639, N637, N495, N361);
xor XOR2 (N640, N598, N122);
not NOT1 (N641, N619);
nor NOR2 (N642, N632, N558);
buf BUF1 (N643, N642);
or OR2 (N644, N615, N546);
nor NOR2 (N645, N639, N481);
nor NOR2 (N646, N638, N151);
not NOT1 (N647, N635);
and AND2 (N648, N644, N91);
not NOT1 (N649, N631);
buf BUF1 (N650, N640);
nor NOR3 (N651, N641, N288, N213);
and AND4 (N652, N650, N560, N321, N174);
and AND4 (N653, N636, N439, N579, N371);
or OR2 (N654, N645, N352);
nor NOR2 (N655, N647, N220);
buf BUF1 (N656, N655);
not NOT1 (N657, N656);
buf BUF1 (N658, N652);
xor XOR2 (N659, N658, N236);
nor NOR2 (N660, N657, N190);
and AND3 (N661, N648, N532, N429);
nand NAND3 (N662, N629, N199, N73);
and AND3 (N663, N643, N374, N371);
and AND4 (N664, N651, N150, N158, N192);
buf BUF1 (N665, N659);
xor XOR2 (N666, N660, N638);
nand NAND2 (N667, N666, N642);
not NOT1 (N668, N667);
nand NAND2 (N669, N663, N514);
or OR3 (N670, N669, N165, N436);
not NOT1 (N671, N661);
buf BUF1 (N672, N649);
or OR4 (N673, N653, N495, N601, N359);
nor NOR2 (N674, N672, N294);
nor NOR3 (N675, N654, N76, N510);
and AND4 (N676, N673, N441, N449, N653);
and AND2 (N677, N664, N638);
not NOT1 (N678, N665);
and AND2 (N679, N674, N500);
nand NAND2 (N680, N646, N522);
nor NOR3 (N681, N662, N577, N555);
not NOT1 (N682, N671);
xor XOR2 (N683, N678, N123);
xor XOR2 (N684, N680, N507);
or OR3 (N685, N668, N302, N631);
nand NAND2 (N686, N682, N348);
not NOT1 (N687, N686);
or OR3 (N688, N675, N363, N402);
or OR3 (N689, N688, N613, N19);
buf BUF1 (N690, N684);
or OR2 (N691, N670, N605);
and AND3 (N692, N685, N689, N119);
nor NOR2 (N693, N648, N142);
nand NAND2 (N694, N692, N192);
xor XOR2 (N695, N693, N41);
buf BUF1 (N696, N691);
buf BUF1 (N697, N696);
nor NOR2 (N698, N694, N246);
or OR4 (N699, N681, N515, N494, N656);
or OR3 (N700, N698, N507, N664);
not NOT1 (N701, N677);
nand NAND4 (N702, N701, N61, N323, N471);
or OR2 (N703, N676, N619);
nand NAND2 (N704, N697, N159);
not NOT1 (N705, N699);
nor NOR4 (N706, N695, N356, N401, N75);
nor NOR4 (N707, N702, N197, N424, N578);
or OR4 (N708, N683, N564, N519, N29);
nand NAND4 (N709, N679, N582, N502, N478);
nand NAND3 (N710, N703, N674, N453);
nand NAND3 (N711, N687, N535, N570);
nand NAND3 (N712, N710, N223, N251);
and AND3 (N713, N705, N288, N286);
nor NOR2 (N714, N708, N345);
not NOT1 (N715, N706);
or OR2 (N716, N690, N354);
and AND4 (N717, N716, N75, N234, N256);
nor NOR4 (N718, N715, N425, N228, N262);
not NOT1 (N719, N700);
and AND2 (N720, N711, N587);
or OR4 (N721, N704, N543, N390, N540);
nand NAND4 (N722, N714, N344, N124, N618);
or OR4 (N723, N712, N540, N74, N270);
xor XOR2 (N724, N721, N64);
nor NOR3 (N725, N724, N570, N564);
nand NAND3 (N726, N723, N450, N513);
and AND2 (N727, N709, N276);
xor XOR2 (N728, N727, N66);
nand NAND2 (N729, N725, N568);
buf BUF1 (N730, N713);
xor XOR2 (N731, N722, N570);
nor NOR4 (N732, N719, N409, N614, N686);
nand NAND4 (N733, N718, N197, N596, N481);
and AND2 (N734, N733, N663);
nor NOR4 (N735, N730, N228, N640, N376);
xor XOR2 (N736, N717, N629);
or OR2 (N737, N734, N397);
nor NOR4 (N738, N736, N157, N42, N686);
xor XOR2 (N739, N726, N662);
and AND2 (N740, N735, N636);
or OR2 (N741, N731, N37);
not NOT1 (N742, N739);
buf BUF1 (N743, N738);
buf BUF1 (N744, N728);
nand NAND4 (N745, N741, N582, N299, N575);
buf BUF1 (N746, N740);
buf BUF1 (N747, N732);
nor NOR2 (N748, N729, N109);
buf BUF1 (N749, N746);
nand NAND4 (N750, N707, N440, N17, N380);
nand NAND3 (N751, N745, N199, N306);
nand NAND4 (N752, N751, N598, N190, N260);
xor XOR2 (N753, N749, N37);
xor XOR2 (N754, N750, N93);
xor XOR2 (N755, N748, N245);
xor XOR2 (N756, N720, N541);
nor NOR3 (N757, N752, N513, N185);
or OR4 (N758, N753, N288, N153, N232);
nand NAND4 (N759, N754, N29, N159, N118);
nor NOR2 (N760, N756, N612);
nand NAND2 (N761, N758, N201);
nor NOR3 (N762, N757, N257, N495);
and AND2 (N763, N744, N251);
and AND3 (N764, N759, N235, N249);
not NOT1 (N765, N747);
and AND2 (N766, N762, N351);
or OR3 (N767, N764, N86, N700);
and AND3 (N768, N763, N59, N437);
buf BUF1 (N769, N743);
nand NAND4 (N770, N769, N331, N692, N49);
buf BUF1 (N771, N767);
buf BUF1 (N772, N765);
buf BUF1 (N773, N742);
and AND2 (N774, N772, N291);
xor XOR2 (N775, N770, N436);
xor XOR2 (N776, N774, N397);
buf BUF1 (N777, N761);
buf BUF1 (N778, N775);
and AND2 (N779, N737, N393);
not NOT1 (N780, N755);
xor XOR2 (N781, N771, N113);
nand NAND2 (N782, N777, N160);
xor XOR2 (N783, N778, N720);
and AND3 (N784, N783, N111, N370);
nor NOR3 (N785, N760, N610, N170);
and AND3 (N786, N785, N633, N601);
xor XOR2 (N787, N779, N774);
xor XOR2 (N788, N784, N385);
buf BUF1 (N789, N780);
nor NOR4 (N790, N773, N382, N132, N425);
nand NAND3 (N791, N768, N54, N587);
and AND4 (N792, N787, N151, N194, N722);
buf BUF1 (N793, N790);
nor NOR4 (N794, N766, N308, N103, N274);
buf BUF1 (N795, N794);
not NOT1 (N796, N793);
and AND2 (N797, N792, N563);
or OR2 (N798, N791, N206);
buf BUF1 (N799, N789);
nor NOR4 (N800, N796, N71, N365, N509);
or OR3 (N801, N800, N645, N72);
or OR4 (N802, N781, N539, N515, N418);
xor XOR2 (N803, N797, N5);
not NOT1 (N804, N795);
or OR2 (N805, N804, N772);
nand NAND4 (N806, N798, N685, N53, N575);
not NOT1 (N807, N782);
or OR2 (N808, N803, N750);
nor NOR2 (N809, N786, N377);
buf BUF1 (N810, N802);
not NOT1 (N811, N805);
and AND4 (N812, N809, N775, N623, N681);
xor XOR2 (N813, N788, N74);
and AND4 (N814, N807, N285, N233, N595);
and AND4 (N815, N811, N319, N344, N367);
nor NOR2 (N816, N808, N28);
and AND4 (N817, N810, N799, N616, N47);
not NOT1 (N818, N744);
and AND2 (N819, N776, N271);
nor NOR3 (N820, N801, N124, N426);
xor XOR2 (N821, N814, N26);
not NOT1 (N822, N813);
buf BUF1 (N823, N821);
nor NOR4 (N824, N816, N288, N52, N27);
not NOT1 (N825, N823);
or OR3 (N826, N806, N774, N762);
nor NOR3 (N827, N812, N640, N649);
buf BUF1 (N828, N819);
and AND4 (N829, N815, N277, N185, N230);
xor XOR2 (N830, N824, N495);
not NOT1 (N831, N830);
or OR3 (N832, N817, N740, N406);
nor NOR2 (N833, N826, N168);
xor XOR2 (N834, N825, N635);
nor NOR4 (N835, N834, N740, N567, N376);
nand NAND2 (N836, N829, N719);
and AND4 (N837, N836, N663, N146, N121);
not NOT1 (N838, N818);
and AND3 (N839, N837, N794, N227);
buf BUF1 (N840, N820);
not NOT1 (N841, N828);
or OR4 (N842, N831, N167, N611, N839);
nand NAND2 (N843, N78, N192);
nand NAND2 (N844, N822, N535);
xor XOR2 (N845, N827, N402);
nand NAND2 (N846, N840, N816);
nand NAND2 (N847, N838, N301);
and AND4 (N848, N841, N728, N87, N830);
buf BUF1 (N849, N848);
not NOT1 (N850, N844);
or OR3 (N851, N833, N244, N230);
and AND3 (N852, N843, N795, N580);
not NOT1 (N853, N845);
or OR4 (N854, N853, N768, N781, N105);
or OR3 (N855, N854, N341, N167);
nand NAND3 (N856, N842, N152, N20);
and AND4 (N857, N856, N680, N735, N362);
nor NOR4 (N858, N857, N792, N665, N830);
buf BUF1 (N859, N850);
buf BUF1 (N860, N847);
and AND2 (N861, N859, N681);
not NOT1 (N862, N851);
or OR3 (N863, N860, N621, N430);
buf BUF1 (N864, N846);
xor XOR2 (N865, N832, N844);
not NOT1 (N866, N855);
nand NAND3 (N867, N835, N831, N476);
buf BUF1 (N868, N866);
buf BUF1 (N869, N849);
buf BUF1 (N870, N864);
nand NAND2 (N871, N865, N793);
nand NAND3 (N872, N869, N842, N211);
or OR3 (N873, N852, N163, N730);
not NOT1 (N874, N861);
and AND2 (N875, N874, N381);
not NOT1 (N876, N873);
not NOT1 (N877, N875);
nand NAND2 (N878, N867, N508);
or OR2 (N879, N872, N736);
not NOT1 (N880, N877);
nor NOR4 (N881, N876, N15, N639, N451);
not NOT1 (N882, N862);
not NOT1 (N883, N880);
not NOT1 (N884, N879);
buf BUF1 (N885, N878);
and AND2 (N886, N868, N319);
and AND3 (N887, N871, N543, N204);
nor NOR4 (N888, N882, N346, N490, N152);
nor NOR4 (N889, N888, N769, N314, N785);
nor NOR2 (N890, N889, N398);
not NOT1 (N891, N884);
buf BUF1 (N892, N870);
buf BUF1 (N893, N890);
and AND2 (N894, N893, N282);
not NOT1 (N895, N886);
or OR4 (N896, N887, N370, N366, N367);
nor NOR2 (N897, N881, N530);
or OR3 (N898, N858, N99, N894);
or OR4 (N899, N272, N197, N499, N587);
buf BUF1 (N900, N885);
nand NAND2 (N901, N900, N454);
buf BUF1 (N902, N895);
and AND4 (N903, N897, N191, N802, N151);
nand NAND4 (N904, N902, N765, N137, N803);
nor NOR3 (N905, N883, N464, N83);
and AND4 (N906, N905, N246, N606, N614);
xor XOR2 (N907, N904, N555);
not NOT1 (N908, N863);
buf BUF1 (N909, N898);
xor XOR2 (N910, N908, N450);
and AND4 (N911, N903, N849, N478, N482);
and AND3 (N912, N901, N56, N830);
not NOT1 (N913, N912);
or OR2 (N914, N909, N724);
or OR3 (N915, N910, N299, N255);
or OR4 (N916, N896, N518, N732, N620);
nand NAND3 (N917, N906, N129, N910);
buf BUF1 (N918, N892);
not NOT1 (N919, N917);
or OR3 (N920, N914, N266, N573);
nand NAND2 (N921, N916, N613);
or OR2 (N922, N913, N134);
buf BUF1 (N923, N899);
buf BUF1 (N924, N918);
buf BUF1 (N925, N921);
or OR3 (N926, N922, N406, N143);
or OR4 (N927, N925, N771, N850, N621);
buf BUF1 (N928, N907);
not NOT1 (N929, N923);
nor NOR4 (N930, N927, N893, N567, N122);
and AND4 (N931, N924, N414, N678, N501);
nand NAND3 (N932, N931, N156, N798);
xor XOR2 (N933, N930, N743);
nand NAND2 (N934, N920, N437);
and AND2 (N935, N926, N664);
xor XOR2 (N936, N915, N824);
xor XOR2 (N937, N928, N504);
nor NOR4 (N938, N911, N220, N456, N625);
and AND3 (N939, N891, N406, N299);
or OR4 (N940, N933, N183, N344, N522);
not NOT1 (N941, N934);
not NOT1 (N942, N929);
buf BUF1 (N943, N941);
and AND4 (N944, N940, N332, N837, N821);
not NOT1 (N945, N943);
and AND3 (N946, N938, N689, N921);
xor XOR2 (N947, N946, N198);
nand NAND3 (N948, N947, N911, N514);
and AND4 (N949, N948, N580, N434, N782);
xor XOR2 (N950, N944, N801);
not NOT1 (N951, N932);
nand NAND3 (N952, N936, N465, N283);
and AND3 (N953, N950, N665, N44);
nor NOR4 (N954, N949, N924, N366, N314);
nor NOR4 (N955, N953, N194, N224, N145);
or OR4 (N956, N954, N531, N354, N731);
nor NOR2 (N957, N955, N97);
xor XOR2 (N958, N956, N661);
or OR3 (N959, N942, N576, N99);
nand NAND3 (N960, N935, N213, N475);
nor NOR2 (N961, N952, N678);
buf BUF1 (N962, N959);
nor NOR3 (N963, N939, N631, N567);
buf BUF1 (N964, N937);
nor NOR3 (N965, N957, N913, N885);
not NOT1 (N966, N965);
xor XOR2 (N967, N966, N660);
nand NAND2 (N968, N945, N212);
nand NAND3 (N969, N958, N559, N781);
or OR2 (N970, N961, N467);
buf BUF1 (N971, N962);
and AND2 (N972, N963, N338);
or OR2 (N973, N919, N756);
not NOT1 (N974, N971);
not NOT1 (N975, N951);
buf BUF1 (N976, N968);
or OR2 (N977, N976, N328);
and AND3 (N978, N970, N251, N823);
and AND3 (N979, N977, N528, N334);
not NOT1 (N980, N975);
buf BUF1 (N981, N974);
buf BUF1 (N982, N973);
and AND3 (N983, N969, N888, N879);
nor NOR4 (N984, N982, N73, N18, N960);
or OR2 (N985, N694, N489);
buf BUF1 (N986, N981);
buf BUF1 (N987, N964);
buf BUF1 (N988, N985);
nand NAND2 (N989, N980, N382);
nor NOR4 (N990, N989, N9, N287, N404);
and AND2 (N991, N967, N920);
nand NAND4 (N992, N978, N851, N979, N156);
or OR3 (N993, N85, N369, N608);
and AND2 (N994, N990, N880);
not NOT1 (N995, N993);
and AND3 (N996, N984, N510, N915);
nor NOR3 (N997, N986, N173, N155);
nor NOR3 (N998, N992, N84, N65);
and AND2 (N999, N994, N9);
nor NOR2 (N1000, N987, N765);
buf BUF1 (N1001, N991);
not NOT1 (N1002, N1000);
nand NAND3 (N1003, N972, N433, N791);
and AND4 (N1004, N1002, N610, N872, N473);
nand NAND2 (N1005, N998, N14);
not NOT1 (N1006, N1004);
not NOT1 (N1007, N995);
not NOT1 (N1008, N983);
not NOT1 (N1009, N1006);
or OR3 (N1010, N999, N132, N226);
or OR2 (N1011, N1001, N376);
and AND3 (N1012, N1009, N165, N56);
nand NAND2 (N1013, N1008, N651);
nor NOR4 (N1014, N988, N249, N518, N531);
not NOT1 (N1015, N1003);
and AND2 (N1016, N997, N88);
xor XOR2 (N1017, N1012, N479);
nand NAND2 (N1018, N1016, N11);
xor XOR2 (N1019, N1010, N323);
nor NOR3 (N1020, N1015, N237, N354);
nor NOR4 (N1021, N1011, N429, N230, N303);
not NOT1 (N1022, N1014);
nand NAND2 (N1023, N1017, N260);
xor XOR2 (N1024, N1013, N184);
nand NAND3 (N1025, N1018, N777, N521);
not NOT1 (N1026, N1021);
xor XOR2 (N1027, N1019, N177);
buf BUF1 (N1028, N1027);
xor XOR2 (N1029, N1022, N588);
nor NOR3 (N1030, N1007, N379, N739);
or OR2 (N1031, N1024, N830);
and AND4 (N1032, N1005, N428, N664, N315);
xor XOR2 (N1033, N1032, N301);
nor NOR4 (N1034, N1033, N814, N454, N784);
or OR3 (N1035, N1025, N842, N550);
nor NOR4 (N1036, N1023, N564, N613, N124);
nor NOR2 (N1037, N1026, N372);
buf BUF1 (N1038, N1031);
or OR3 (N1039, N1037, N489, N984);
nand NAND2 (N1040, N996, N43);
nor NOR4 (N1041, N1034, N382, N51, N814);
or OR3 (N1042, N1029, N590, N977);
buf BUF1 (N1043, N1039);
nor NOR3 (N1044, N1035, N51, N680);
and AND2 (N1045, N1028, N481);
and AND4 (N1046, N1040, N241, N468, N227);
xor XOR2 (N1047, N1041, N231);
buf BUF1 (N1048, N1038);
or OR4 (N1049, N1045, N75, N257, N519);
and AND4 (N1050, N1044, N242, N489, N218);
xor XOR2 (N1051, N1030, N445);
nand NAND4 (N1052, N1036, N1049, N195, N964);
not NOT1 (N1053, N197);
buf BUF1 (N1054, N1052);
xor XOR2 (N1055, N1050, N279);
nand NAND4 (N1056, N1046, N699, N1001, N626);
and AND2 (N1057, N1020, N63);
and AND2 (N1058, N1043, N27);
nand NAND4 (N1059, N1051, N141, N29, N881);
not NOT1 (N1060, N1042);
buf BUF1 (N1061, N1059);
and AND3 (N1062, N1060, N302, N521);
buf BUF1 (N1063, N1053);
xor XOR2 (N1064, N1054, N52);
xor XOR2 (N1065, N1063, N678);
buf BUF1 (N1066, N1056);
buf BUF1 (N1067, N1064);
xor XOR2 (N1068, N1067, N268);
or OR2 (N1069, N1066, N152);
not NOT1 (N1070, N1061);
nor NOR3 (N1071, N1062, N336, N603);
not NOT1 (N1072, N1068);
nand NAND2 (N1073, N1057, N1004);
or OR4 (N1074, N1058, N45, N117, N1053);
or OR4 (N1075, N1055, N649, N928, N116);
not NOT1 (N1076, N1074);
nor NOR2 (N1077, N1048, N748);
buf BUF1 (N1078, N1077);
not NOT1 (N1079, N1065);
not NOT1 (N1080, N1069);
buf BUF1 (N1081, N1047);
xor XOR2 (N1082, N1079, N688);
not NOT1 (N1083, N1080);
nor NOR3 (N1084, N1072, N925, N961);
not NOT1 (N1085, N1076);
nand NAND4 (N1086, N1073, N271, N933, N106);
xor XOR2 (N1087, N1071, N732);
xor XOR2 (N1088, N1081, N1009);
and AND2 (N1089, N1084, N661);
nand NAND4 (N1090, N1086, N492, N62, N378);
nand NAND2 (N1091, N1070, N69);
nand NAND2 (N1092, N1088, N175);
not NOT1 (N1093, N1083);
xor XOR2 (N1094, N1090, N1044);
nand NAND2 (N1095, N1087, N226);
buf BUF1 (N1096, N1082);
buf BUF1 (N1097, N1075);
nor NOR2 (N1098, N1091, N282);
or OR4 (N1099, N1093, N823, N43, N374);
nor NOR2 (N1100, N1085, N137);
not NOT1 (N1101, N1078);
xor XOR2 (N1102, N1094, N76);
xor XOR2 (N1103, N1097, N221);
buf BUF1 (N1104, N1092);
not NOT1 (N1105, N1089);
nand NAND2 (N1106, N1102, N211);
buf BUF1 (N1107, N1103);
nand NAND2 (N1108, N1098, N443);
nand NAND2 (N1109, N1104, N865);
or OR2 (N1110, N1107, N839);
or OR4 (N1111, N1096, N1028, N153, N1075);
nor NOR3 (N1112, N1109, N543, N327);
buf BUF1 (N1113, N1100);
nor NOR2 (N1114, N1101, N75);
buf BUF1 (N1115, N1108);
xor XOR2 (N1116, N1110, N812);
buf BUF1 (N1117, N1116);
nand NAND2 (N1118, N1114, N476);
nand NAND3 (N1119, N1113, N714, N1016);
xor XOR2 (N1120, N1112, N221);
and AND4 (N1121, N1099, N55, N615, N307);
buf BUF1 (N1122, N1111);
or OR3 (N1123, N1121, N397, N353);
nand NAND4 (N1124, N1118, N509, N1035, N1048);
nor NOR2 (N1125, N1117, N574);
buf BUF1 (N1126, N1119);
not NOT1 (N1127, N1106);
buf BUF1 (N1128, N1127);
not NOT1 (N1129, N1105);
not NOT1 (N1130, N1128);
nand NAND2 (N1131, N1126, N212);
or OR3 (N1132, N1122, N365, N686);
buf BUF1 (N1133, N1132);
xor XOR2 (N1134, N1129, N852);
nand NAND3 (N1135, N1131, N1049, N329);
buf BUF1 (N1136, N1133);
or OR3 (N1137, N1130, N376, N859);
not NOT1 (N1138, N1125);
nor NOR4 (N1139, N1123, N446, N26, N262);
nand NAND3 (N1140, N1095, N647, N460);
nand NAND4 (N1141, N1138, N383, N824, N818);
nor NOR2 (N1142, N1141, N345);
or OR2 (N1143, N1139, N272);
and AND4 (N1144, N1115, N676, N136, N207);
nand NAND3 (N1145, N1142, N363, N345);
and AND4 (N1146, N1140, N256, N739, N202);
xor XOR2 (N1147, N1120, N385);
nor NOR4 (N1148, N1136, N573, N518, N586);
buf BUF1 (N1149, N1143);
or OR2 (N1150, N1124, N320);
and AND3 (N1151, N1144, N410, N311);
nor NOR3 (N1152, N1135, N748, N323);
and AND3 (N1153, N1151, N538, N949);
nand NAND2 (N1154, N1146, N542);
nor NOR2 (N1155, N1147, N684);
buf BUF1 (N1156, N1149);
or OR3 (N1157, N1150, N1053, N664);
or OR4 (N1158, N1137, N958, N626, N349);
nor NOR4 (N1159, N1155, N370, N1085, N476);
not NOT1 (N1160, N1145);
or OR4 (N1161, N1156, N1013, N1076, N1069);
nor NOR3 (N1162, N1148, N853, N539);
nand NAND3 (N1163, N1154, N443, N489);
and AND3 (N1164, N1160, N239, N930);
xor XOR2 (N1165, N1164, N68);
nand NAND2 (N1166, N1134, N840);
and AND2 (N1167, N1157, N967);
xor XOR2 (N1168, N1163, N44);
nor NOR3 (N1169, N1167, N504, N204);
buf BUF1 (N1170, N1152);
or OR2 (N1171, N1166, N79);
buf BUF1 (N1172, N1169);
and AND4 (N1173, N1158, N1021, N568, N1037);
nand NAND2 (N1174, N1153, N28);
nand NAND3 (N1175, N1172, N745, N1071);
buf BUF1 (N1176, N1159);
nand NAND4 (N1177, N1162, N394, N445, N112);
and AND4 (N1178, N1173, N760, N456, N541);
buf BUF1 (N1179, N1171);
nor NOR4 (N1180, N1178, N327, N994, N1084);
buf BUF1 (N1181, N1161);
nor NOR4 (N1182, N1175, N992, N78, N93);
nor NOR4 (N1183, N1176, N941, N1058, N268);
or OR4 (N1184, N1181, N103, N1067, N1044);
buf BUF1 (N1185, N1177);
not NOT1 (N1186, N1170);
xor XOR2 (N1187, N1165, N603);
or OR3 (N1188, N1184, N682, N599);
and AND2 (N1189, N1188, N931);
and AND2 (N1190, N1168, N678);
xor XOR2 (N1191, N1185, N79);
and AND4 (N1192, N1179, N890, N893, N76);
not NOT1 (N1193, N1192);
or OR3 (N1194, N1182, N552, N724);
nand NAND3 (N1195, N1193, N190, N722);
xor XOR2 (N1196, N1189, N589);
and AND4 (N1197, N1180, N3, N297, N477);
xor XOR2 (N1198, N1183, N1179);
nor NOR2 (N1199, N1197, N964);
not NOT1 (N1200, N1198);
not NOT1 (N1201, N1191);
buf BUF1 (N1202, N1200);
nand NAND3 (N1203, N1202, N237, N428);
and AND4 (N1204, N1194, N277, N679, N645);
nor NOR2 (N1205, N1187, N156);
not NOT1 (N1206, N1205);
nor NOR3 (N1207, N1195, N140, N630);
nor NOR3 (N1208, N1206, N1030, N852);
nand NAND2 (N1209, N1208, N584);
xor XOR2 (N1210, N1199, N578);
not NOT1 (N1211, N1210);
nand NAND3 (N1212, N1174, N402, N313);
nand NAND3 (N1213, N1196, N233, N329);
or OR4 (N1214, N1211, N373, N874, N283);
and AND3 (N1215, N1201, N369, N814);
nand NAND2 (N1216, N1203, N601);
buf BUF1 (N1217, N1212);
xor XOR2 (N1218, N1209, N543);
not NOT1 (N1219, N1217);
or OR4 (N1220, N1219, N669, N470, N6);
or OR4 (N1221, N1213, N1154, N563, N867);
nand NAND3 (N1222, N1190, N707, N1219);
buf BUF1 (N1223, N1204);
xor XOR2 (N1224, N1186, N582);
nor NOR2 (N1225, N1207, N255);
or OR3 (N1226, N1223, N389, N808);
xor XOR2 (N1227, N1225, N684);
not NOT1 (N1228, N1216);
buf BUF1 (N1229, N1220);
nor NOR2 (N1230, N1227, N217);
buf BUF1 (N1231, N1221);
not NOT1 (N1232, N1224);
nor NOR3 (N1233, N1232, N814, N561);
not NOT1 (N1234, N1228);
buf BUF1 (N1235, N1222);
or OR4 (N1236, N1233, N31, N445, N875);
and AND4 (N1237, N1229, N901, N1033, N911);
nor NOR3 (N1238, N1214, N907, N404);
nand NAND2 (N1239, N1215, N18);
nor NOR2 (N1240, N1238, N1191);
nand NAND2 (N1241, N1231, N51);
buf BUF1 (N1242, N1241);
nand NAND3 (N1243, N1218, N260, N298);
or OR2 (N1244, N1234, N470);
buf BUF1 (N1245, N1240);
not NOT1 (N1246, N1239);
and AND3 (N1247, N1242, N1057, N1004);
nor NOR3 (N1248, N1235, N337, N429);
nor NOR2 (N1249, N1236, N116);
nor NOR2 (N1250, N1244, N926);
not NOT1 (N1251, N1237);
xor XOR2 (N1252, N1245, N709);
buf BUF1 (N1253, N1243);
or OR4 (N1254, N1248, N1015, N379, N389);
xor XOR2 (N1255, N1250, N46);
xor XOR2 (N1256, N1226, N584);
xor XOR2 (N1257, N1255, N556);
buf BUF1 (N1258, N1246);
buf BUF1 (N1259, N1258);
buf BUF1 (N1260, N1252);
not NOT1 (N1261, N1249);
or OR3 (N1262, N1251, N1066, N794);
nor NOR4 (N1263, N1254, N94, N1258, N675);
or OR4 (N1264, N1260, N895, N103, N323);
nor NOR2 (N1265, N1264, N866);
nand NAND4 (N1266, N1256, N514, N135, N212);
nand NAND3 (N1267, N1262, N140, N448);
buf BUF1 (N1268, N1263);
and AND3 (N1269, N1266, N1014, N159);
nor NOR4 (N1270, N1247, N250, N435, N1025);
nand NAND3 (N1271, N1253, N642, N247);
xor XOR2 (N1272, N1261, N134);
nor NOR4 (N1273, N1269, N877, N585, N450);
nor NOR2 (N1274, N1230, N855);
or OR3 (N1275, N1267, N937, N1126);
and AND4 (N1276, N1272, N666, N243, N1157);
and AND3 (N1277, N1270, N325, N718);
buf BUF1 (N1278, N1265);
and AND3 (N1279, N1276, N210, N1097);
or OR2 (N1280, N1257, N510);
or OR2 (N1281, N1268, N76);
and AND2 (N1282, N1281, N753);
and AND3 (N1283, N1280, N711, N339);
nand NAND4 (N1284, N1274, N301, N407, N813);
buf BUF1 (N1285, N1284);
nand NAND4 (N1286, N1279, N54, N1250, N1200);
buf BUF1 (N1287, N1282);
buf BUF1 (N1288, N1277);
or OR4 (N1289, N1259, N634, N1200, N20);
buf BUF1 (N1290, N1278);
buf BUF1 (N1291, N1286);
or OR3 (N1292, N1291, N452, N539);
xor XOR2 (N1293, N1275, N1104);
not NOT1 (N1294, N1290);
not NOT1 (N1295, N1287);
or OR4 (N1296, N1271, N1163, N897, N1240);
nand NAND3 (N1297, N1289, N183, N925);
buf BUF1 (N1298, N1294);
nor NOR3 (N1299, N1295, N301, N881);
not NOT1 (N1300, N1298);
xor XOR2 (N1301, N1273, N14);
or OR3 (N1302, N1296, N754, N373);
not NOT1 (N1303, N1301);
buf BUF1 (N1304, N1288);
nand NAND2 (N1305, N1292, N610);
or OR4 (N1306, N1293, N317, N16, N1237);
not NOT1 (N1307, N1303);
xor XOR2 (N1308, N1304, N204);
and AND4 (N1309, N1306, N320, N867, N1142);
buf BUF1 (N1310, N1305);
and AND2 (N1311, N1300, N486);
nor NOR2 (N1312, N1302, N794);
or OR4 (N1313, N1308, N605, N299, N657);
nor NOR2 (N1314, N1297, N285);
nor NOR2 (N1315, N1285, N231);
xor XOR2 (N1316, N1313, N363);
nand NAND2 (N1317, N1315, N801);
or OR3 (N1318, N1311, N351, N1068);
nor NOR2 (N1319, N1299, N1009);
nand NAND3 (N1320, N1307, N1259, N308);
xor XOR2 (N1321, N1309, N860);
buf BUF1 (N1322, N1312);
or OR3 (N1323, N1317, N761, N212);
not NOT1 (N1324, N1321);
or OR3 (N1325, N1310, N121, N1120);
buf BUF1 (N1326, N1314);
buf BUF1 (N1327, N1319);
nor NOR3 (N1328, N1323, N1198, N1251);
nand NAND2 (N1329, N1327, N65);
or OR3 (N1330, N1326, N1080, N575);
or OR2 (N1331, N1318, N994);
not NOT1 (N1332, N1322);
nor NOR4 (N1333, N1316, N1158, N518, N1142);
xor XOR2 (N1334, N1320, N223);
and AND2 (N1335, N1329, N11);
nor NOR3 (N1336, N1333, N1203, N482);
nor NOR4 (N1337, N1335, N190, N684, N614);
or OR4 (N1338, N1337, N104, N263, N821);
or OR2 (N1339, N1338, N463);
and AND2 (N1340, N1325, N954);
nor NOR4 (N1341, N1328, N142, N1025, N1097);
nand NAND4 (N1342, N1339, N140, N398, N436);
xor XOR2 (N1343, N1332, N944);
xor XOR2 (N1344, N1343, N72);
nor NOR2 (N1345, N1324, N1040);
buf BUF1 (N1346, N1331);
nand NAND4 (N1347, N1346, N824, N335, N109);
or OR4 (N1348, N1342, N1230, N763, N1237);
nor NOR2 (N1349, N1334, N287);
nand NAND3 (N1350, N1347, N572, N216);
not NOT1 (N1351, N1341);
nor NOR3 (N1352, N1351, N490, N1181);
buf BUF1 (N1353, N1336);
not NOT1 (N1354, N1350);
or OR2 (N1355, N1348, N416);
xor XOR2 (N1356, N1283, N1062);
buf BUF1 (N1357, N1344);
buf BUF1 (N1358, N1355);
nor NOR2 (N1359, N1354, N386);
buf BUF1 (N1360, N1357);
and AND2 (N1361, N1352, N1351);
or OR2 (N1362, N1340, N1225);
or OR3 (N1363, N1345, N297, N775);
nor NOR2 (N1364, N1356, N775);
and AND2 (N1365, N1359, N1220);
nor NOR3 (N1366, N1364, N463, N1106);
nor NOR4 (N1367, N1349, N656, N650, N326);
nand NAND4 (N1368, N1330, N670, N88, N1302);
nand NAND4 (N1369, N1358, N1206, N1214, N1019);
buf BUF1 (N1370, N1360);
xor XOR2 (N1371, N1362, N207);
buf BUF1 (N1372, N1367);
and AND4 (N1373, N1368, N658, N863, N703);
buf BUF1 (N1374, N1361);
and AND4 (N1375, N1373, N86, N1290, N525);
not NOT1 (N1376, N1369);
and AND2 (N1377, N1374, N966);
xor XOR2 (N1378, N1353, N146);
or OR3 (N1379, N1372, N542, N187);
or OR3 (N1380, N1379, N354, N1041);
xor XOR2 (N1381, N1370, N1322);
and AND4 (N1382, N1366, N1187, N541, N513);
or OR4 (N1383, N1371, N618, N601, N954);
nand NAND3 (N1384, N1382, N1256, N700);
not NOT1 (N1385, N1384);
not NOT1 (N1386, N1377);
buf BUF1 (N1387, N1365);
nor NOR4 (N1388, N1381, N929, N1303, N970);
not NOT1 (N1389, N1375);
nand NAND4 (N1390, N1378, N422, N439, N951);
nand NAND3 (N1391, N1385, N1365, N590);
nor NOR4 (N1392, N1391, N179, N348, N392);
nand NAND4 (N1393, N1389, N380, N104, N1263);
xor XOR2 (N1394, N1383, N417);
nor NOR4 (N1395, N1387, N688, N874, N1361);
buf BUF1 (N1396, N1392);
nor NOR4 (N1397, N1394, N1373, N1300, N981);
xor XOR2 (N1398, N1363, N157);
and AND2 (N1399, N1386, N820);
nor NOR3 (N1400, N1399, N1109, N49);
xor XOR2 (N1401, N1400, N341);
or OR2 (N1402, N1398, N227);
or OR2 (N1403, N1395, N1137);
xor XOR2 (N1404, N1390, N1012);
nor NOR4 (N1405, N1380, N253, N758, N668);
nand NAND4 (N1406, N1397, N701, N732, N21);
not NOT1 (N1407, N1405);
not NOT1 (N1408, N1401);
buf BUF1 (N1409, N1404);
not NOT1 (N1410, N1407);
xor XOR2 (N1411, N1410, N132);
nor NOR2 (N1412, N1406, N636);
and AND2 (N1413, N1409, N632);
and AND2 (N1414, N1412, N751);
buf BUF1 (N1415, N1402);
nor NOR3 (N1416, N1376, N1321, N30);
xor XOR2 (N1417, N1416, N1139);
xor XOR2 (N1418, N1414, N1307);
nor NOR4 (N1419, N1403, N404, N387, N1238);
nor NOR3 (N1420, N1419, N56, N1353);
nor NOR2 (N1421, N1411, N1406);
buf BUF1 (N1422, N1420);
nand NAND2 (N1423, N1422, N56);
buf BUF1 (N1424, N1418);
not NOT1 (N1425, N1396);
buf BUF1 (N1426, N1388);
buf BUF1 (N1427, N1415);
nand NAND2 (N1428, N1423, N402);
and AND2 (N1429, N1425, N774);
not NOT1 (N1430, N1426);
and AND3 (N1431, N1428, N161, N629);
and AND2 (N1432, N1429, N335);
and AND2 (N1433, N1417, N655);
not NOT1 (N1434, N1433);
buf BUF1 (N1435, N1393);
nand NAND2 (N1436, N1431, N964);
not NOT1 (N1437, N1408);
nand NAND3 (N1438, N1432, N1249, N150);
nor NOR3 (N1439, N1434, N406, N1008);
or OR4 (N1440, N1413, N529, N1427, N96);
or OR4 (N1441, N1247, N200, N1217, N472);
nand NAND4 (N1442, N1441, N169, N1170, N300);
buf BUF1 (N1443, N1438);
and AND2 (N1444, N1442, N1238);
nand NAND3 (N1445, N1421, N474, N881);
xor XOR2 (N1446, N1439, N688);
nand NAND2 (N1447, N1430, N1428);
buf BUF1 (N1448, N1445);
buf BUF1 (N1449, N1440);
nor NOR3 (N1450, N1443, N1009, N1211);
buf BUF1 (N1451, N1437);
or OR4 (N1452, N1436, N429, N1115, N339);
xor XOR2 (N1453, N1444, N1310);
nor NOR4 (N1454, N1451, N632, N665, N585);
nor NOR3 (N1455, N1453, N456, N71);
buf BUF1 (N1456, N1424);
nor NOR4 (N1457, N1449, N993, N1021, N715);
xor XOR2 (N1458, N1450, N1161);
or OR3 (N1459, N1458, N47, N566);
or OR3 (N1460, N1457, N1095, N1371);
nor NOR4 (N1461, N1454, N539, N436, N343);
and AND4 (N1462, N1460, N797, N645, N402);
or OR3 (N1463, N1446, N1400, N1416);
not NOT1 (N1464, N1459);
buf BUF1 (N1465, N1461);
buf BUF1 (N1466, N1448);
nor NOR3 (N1467, N1464, N1463, N926);
nand NAND2 (N1468, N302, N1162);
xor XOR2 (N1469, N1468, N494);
nand NAND3 (N1470, N1435, N14, N400);
nand NAND2 (N1471, N1462, N1072);
not NOT1 (N1472, N1466);
and AND2 (N1473, N1472, N650);
and AND4 (N1474, N1447, N1224, N203, N871);
buf BUF1 (N1475, N1465);
or OR2 (N1476, N1467, N544);
buf BUF1 (N1477, N1471);
not NOT1 (N1478, N1469);
nor NOR2 (N1479, N1473, N1053);
nand NAND2 (N1480, N1475, N1411);
or OR4 (N1481, N1480, N74, N995, N1221);
and AND2 (N1482, N1476, N595);
not NOT1 (N1483, N1479);
or OR4 (N1484, N1452, N1289, N977, N361);
not NOT1 (N1485, N1481);
nor NOR4 (N1486, N1485, N779, N750, N666);
or OR3 (N1487, N1455, N496, N98);
and AND3 (N1488, N1487, N758, N1414);
and AND3 (N1489, N1477, N45, N227);
not NOT1 (N1490, N1474);
or OR4 (N1491, N1484, N809, N1249, N1232);
and AND2 (N1492, N1488, N1337);
or OR4 (N1493, N1456, N535, N1453, N529);
xor XOR2 (N1494, N1482, N629);
nor NOR2 (N1495, N1486, N475);
or OR4 (N1496, N1492, N454, N479, N1293);
nor NOR4 (N1497, N1478, N302, N940, N1486);
nor NOR4 (N1498, N1493, N333, N1284, N33);
nor NOR3 (N1499, N1497, N313, N1037);
buf BUF1 (N1500, N1489);
and AND3 (N1501, N1491, N1105, N1050);
xor XOR2 (N1502, N1483, N55);
nor NOR4 (N1503, N1498, N1189, N1366, N353);
nor NOR2 (N1504, N1502, N311);
nand NAND4 (N1505, N1500, N77, N215, N1502);
not NOT1 (N1506, N1470);
or OR2 (N1507, N1504, N1194);
nand NAND4 (N1508, N1494, N218, N973, N380);
nor NOR3 (N1509, N1507, N694, N1086);
not NOT1 (N1510, N1503);
and AND2 (N1511, N1501, N152);
not NOT1 (N1512, N1499);
not NOT1 (N1513, N1495);
and AND2 (N1514, N1510, N637);
xor XOR2 (N1515, N1511, N1408);
or OR4 (N1516, N1509, N319, N414, N1503);
xor XOR2 (N1517, N1512, N686);
nand NAND3 (N1518, N1514, N199, N381);
nand NAND4 (N1519, N1490, N1093, N1069, N1484);
nor NOR3 (N1520, N1517, N1324, N493);
xor XOR2 (N1521, N1508, N1184);
and AND3 (N1522, N1506, N389, N357);
not NOT1 (N1523, N1520);
nor NOR2 (N1524, N1516, N7);
buf BUF1 (N1525, N1515);
and AND3 (N1526, N1525, N1025, N82);
or OR3 (N1527, N1518, N720, N71);
buf BUF1 (N1528, N1519);
and AND3 (N1529, N1524, N901, N3);
nor NOR4 (N1530, N1528, N319, N176, N1215);
nor NOR2 (N1531, N1521, N342);
or OR3 (N1532, N1513, N53, N473);
or OR4 (N1533, N1527, N267, N235, N402);
nor NOR3 (N1534, N1522, N883, N1011);
and AND2 (N1535, N1532, N19);
or OR3 (N1536, N1529, N994, N1507);
buf BUF1 (N1537, N1534);
xor XOR2 (N1538, N1530, N429);
xor XOR2 (N1539, N1505, N1511);
nand NAND4 (N1540, N1536, N650, N953, N266);
nor NOR3 (N1541, N1535, N493, N933);
and AND3 (N1542, N1540, N273, N1115);
buf BUF1 (N1543, N1523);
and AND3 (N1544, N1533, N1119, N1161);
nand NAND2 (N1545, N1531, N975);
and AND2 (N1546, N1537, N882);
nand NAND2 (N1547, N1546, N55);
or OR2 (N1548, N1538, N1407);
not NOT1 (N1549, N1547);
nand NAND3 (N1550, N1542, N551, N526);
and AND3 (N1551, N1545, N230, N393);
buf BUF1 (N1552, N1544);
buf BUF1 (N1553, N1550);
xor XOR2 (N1554, N1553, N160);
xor XOR2 (N1555, N1496, N1455);
or OR3 (N1556, N1543, N1470, N1521);
not NOT1 (N1557, N1556);
buf BUF1 (N1558, N1557);
xor XOR2 (N1559, N1555, N1521);
nor NOR2 (N1560, N1551, N642);
and AND3 (N1561, N1558, N1154, N843);
nor NOR2 (N1562, N1552, N1332);
nor NOR2 (N1563, N1549, N124);
xor XOR2 (N1564, N1539, N901);
or OR4 (N1565, N1541, N1377, N830, N1273);
nand NAND4 (N1566, N1560, N542, N20, N529);
nand NAND3 (N1567, N1561, N559, N281);
nor NOR2 (N1568, N1548, N1053);
nand NAND2 (N1569, N1564, N774);
buf BUF1 (N1570, N1554);
not NOT1 (N1571, N1526);
xor XOR2 (N1572, N1568, N1020);
and AND3 (N1573, N1567, N1494, N519);
nand NAND4 (N1574, N1562, N404, N192, N969);
nor NOR2 (N1575, N1559, N1344);
buf BUF1 (N1576, N1566);
buf BUF1 (N1577, N1573);
xor XOR2 (N1578, N1570, N79);
nor NOR4 (N1579, N1572, N431, N357, N935);
not NOT1 (N1580, N1576);
not NOT1 (N1581, N1578);
xor XOR2 (N1582, N1571, N396);
or OR4 (N1583, N1563, N294, N1044, N566);
xor XOR2 (N1584, N1565, N1320);
and AND4 (N1585, N1580, N1297, N1356, N1106);
nor NOR3 (N1586, N1579, N278, N292);
xor XOR2 (N1587, N1575, N153);
xor XOR2 (N1588, N1581, N1171);
nor NOR4 (N1589, N1574, N95, N1005, N1500);
nor NOR2 (N1590, N1586, N984);
buf BUF1 (N1591, N1585);
buf BUF1 (N1592, N1569);
nand NAND3 (N1593, N1584, N1435, N693);
nand NAND2 (N1594, N1589, N1083);
not NOT1 (N1595, N1577);
nand NAND3 (N1596, N1588, N1111, N957);
or OR3 (N1597, N1591, N457, N17);
xor XOR2 (N1598, N1594, N200);
or OR4 (N1599, N1596, N709, N574, N850);
xor XOR2 (N1600, N1593, N277);
and AND4 (N1601, N1587, N1374, N390, N1282);
and AND3 (N1602, N1600, N1201, N1312);
and AND2 (N1603, N1590, N84);
buf BUF1 (N1604, N1595);
not NOT1 (N1605, N1601);
not NOT1 (N1606, N1592);
nor NOR4 (N1607, N1597, N790, N1293, N1180);
xor XOR2 (N1608, N1607, N303);
not NOT1 (N1609, N1583);
nor NOR3 (N1610, N1604, N1448, N458);
xor XOR2 (N1611, N1582, N308);
not NOT1 (N1612, N1611);
nor NOR4 (N1613, N1603, N704, N903, N1257);
or OR4 (N1614, N1609, N984, N1359, N1095);
nor NOR2 (N1615, N1608, N693);
nor NOR3 (N1616, N1606, N1016, N1223);
nor NOR3 (N1617, N1616, N611, N222);
and AND3 (N1618, N1614, N1198, N1342);
and AND2 (N1619, N1615, N958);
nand NAND3 (N1620, N1617, N1347, N647);
buf BUF1 (N1621, N1599);
xor XOR2 (N1622, N1618, N1218);
nand NAND4 (N1623, N1619, N1148, N266, N989);
nor NOR4 (N1624, N1621, N1552, N1327, N358);
or OR3 (N1625, N1602, N748, N964);
not NOT1 (N1626, N1622);
nand NAND4 (N1627, N1612, N393, N772, N900);
nor NOR2 (N1628, N1623, N929);
nand NAND2 (N1629, N1598, N729);
or OR2 (N1630, N1627, N1375);
and AND4 (N1631, N1624, N995, N1040, N1322);
nor NOR4 (N1632, N1628, N1444, N1575, N1047);
nand NAND4 (N1633, N1626, N4, N950, N942);
or OR3 (N1634, N1633, N1371, N1432);
xor XOR2 (N1635, N1630, N661);
and AND4 (N1636, N1632, N1622, N248, N728);
or OR3 (N1637, N1613, N167, N1117);
and AND2 (N1638, N1620, N657);
not NOT1 (N1639, N1637);
or OR3 (N1640, N1636, N1534, N1223);
nor NOR4 (N1641, N1605, N178, N826, N265);
buf BUF1 (N1642, N1634);
not NOT1 (N1643, N1631);
not NOT1 (N1644, N1629);
xor XOR2 (N1645, N1644, N904);
nand NAND4 (N1646, N1641, N1386, N853, N606);
nor NOR3 (N1647, N1642, N11, N481);
xor XOR2 (N1648, N1638, N353);
nand NAND2 (N1649, N1647, N37);
not NOT1 (N1650, N1635);
nand NAND2 (N1651, N1640, N1070);
not NOT1 (N1652, N1643);
buf BUF1 (N1653, N1645);
buf BUF1 (N1654, N1649);
nand NAND2 (N1655, N1651, N469);
or OR4 (N1656, N1610, N923, N1436, N183);
nand NAND4 (N1657, N1639, N1334, N1370, N1017);
nand NAND2 (N1658, N1655, N583);
not NOT1 (N1659, N1657);
nand NAND3 (N1660, N1652, N251, N1528);
xor XOR2 (N1661, N1625, N1443);
buf BUF1 (N1662, N1658);
buf BUF1 (N1663, N1662);
nor NOR3 (N1664, N1663, N376, N771);
and AND4 (N1665, N1656, N806, N93, N1362);
nand NAND3 (N1666, N1654, N1269, N1578);
nor NOR4 (N1667, N1664, N1520, N127, N1488);
buf BUF1 (N1668, N1650);
nor NOR4 (N1669, N1665, N671, N147, N1221);
not NOT1 (N1670, N1667);
and AND2 (N1671, N1646, N804);
nand NAND3 (N1672, N1668, N336, N1305);
nand NAND4 (N1673, N1672, N433, N1369, N405);
not NOT1 (N1674, N1648);
nor NOR4 (N1675, N1669, N1201, N631, N758);
nand NAND3 (N1676, N1674, N778, N1264);
nand NAND2 (N1677, N1659, N89);
not NOT1 (N1678, N1666);
nand NAND2 (N1679, N1673, N1546);
xor XOR2 (N1680, N1660, N378);
or OR3 (N1681, N1677, N318, N631);
nor NOR4 (N1682, N1676, N651, N1018, N882);
buf BUF1 (N1683, N1670);
nor NOR4 (N1684, N1680, N549, N816, N538);
xor XOR2 (N1685, N1671, N20);
not NOT1 (N1686, N1661);
xor XOR2 (N1687, N1686, N1183);
nor NOR2 (N1688, N1684, N899);
not NOT1 (N1689, N1688);
buf BUF1 (N1690, N1653);
xor XOR2 (N1691, N1689, N1619);
or OR3 (N1692, N1678, N618, N1592);
or OR2 (N1693, N1692, N1410);
and AND3 (N1694, N1682, N1481, N496);
and AND4 (N1695, N1694, N1553, N1262, N790);
or OR3 (N1696, N1695, N261, N766);
nand NAND2 (N1697, N1691, N117);
not NOT1 (N1698, N1693);
nor NOR3 (N1699, N1690, N1545, N1412);
or OR2 (N1700, N1699, N80);
nor NOR2 (N1701, N1687, N703);
and AND3 (N1702, N1696, N989, N1544);
nand NAND4 (N1703, N1698, N777, N914, N266);
xor XOR2 (N1704, N1700, N300);
xor XOR2 (N1705, N1697, N189);
xor XOR2 (N1706, N1683, N1032);
and AND3 (N1707, N1703, N1488, N102);
nand NAND4 (N1708, N1675, N1685, N1345, N1521);
and AND2 (N1709, N692, N977);
xor XOR2 (N1710, N1708, N1692);
and AND2 (N1711, N1702, N1411);
and AND2 (N1712, N1679, N1105);
xor XOR2 (N1713, N1706, N257);
not NOT1 (N1714, N1709);
buf BUF1 (N1715, N1705);
nor NOR3 (N1716, N1715, N1542, N614);
nor NOR4 (N1717, N1707, N689, N743, N1255);
nor NOR3 (N1718, N1681, N1577, N1026);
not NOT1 (N1719, N1701);
nor NOR3 (N1720, N1711, N438, N811);
and AND2 (N1721, N1710, N330);
nand NAND3 (N1722, N1714, N33, N942);
xor XOR2 (N1723, N1719, N1700);
not NOT1 (N1724, N1721);
and AND2 (N1725, N1723, N1003);
or OR4 (N1726, N1704, N1178, N1076, N1615);
nor NOR3 (N1727, N1725, N424, N1046);
or OR2 (N1728, N1713, N75);
or OR4 (N1729, N1724, N295, N1663, N1726);
or OR2 (N1730, N69, N152);
and AND3 (N1731, N1716, N1054, N804);
or OR2 (N1732, N1729, N1429);
and AND2 (N1733, N1720, N1389);
not NOT1 (N1734, N1712);
or OR3 (N1735, N1718, N1217, N396);
not NOT1 (N1736, N1735);
not NOT1 (N1737, N1728);
buf BUF1 (N1738, N1734);
nor NOR2 (N1739, N1733, N111);
xor XOR2 (N1740, N1717, N333);
buf BUF1 (N1741, N1730);
not NOT1 (N1742, N1722);
and AND2 (N1743, N1739, N513);
nand NAND4 (N1744, N1736, N689, N1220, N42);
buf BUF1 (N1745, N1727);
and AND3 (N1746, N1738, N157, N217);
xor XOR2 (N1747, N1745, N419);
nor NOR3 (N1748, N1743, N1268, N1263);
xor XOR2 (N1749, N1732, N1508);
nand NAND2 (N1750, N1731, N1358);
nor NOR3 (N1751, N1744, N875, N426);
xor XOR2 (N1752, N1749, N311);
buf BUF1 (N1753, N1742);
nand NAND4 (N1754, N1741, N939, N1584, N157);
and AND3 (N1755, N1750, N1540, N410);
nor NOR4 (N1756, N1753, N1652, N1088, N1053);
xor XOR2 (N1757, N1740, N1209);
xor XOR2 (N1758, N1747, N366);
not NOT1 (N1759, N1757);
xor XOR2 (N1760, N1758, N89);
or OR2 (N1761, N1737, N1640);
nand NAND3 (N1762, N1756, N1240, N1512);
xor XOR2 (N1763, N1755, N374);
or OR4 (N1764, N1752, N141, N1363, N13);
nor NOR3 (N1765, N1761, N350, N137);
xor XOR2 (N1766, N1763, N969);
nand NAND4 (N1767, N1759, N460, N508, N396);
buf BUF1 (N1768, N1748);
xor XOR2 (N1769, N1746, N614);
nor NOR2 (N1770, N1768, N884);
xor XOR2 (N1771, N1767, N1403);
nand NAND3 (N1772, N1771, N648, N1513);
nand NAND3 (N1773, N1764, N1148, N1109);
not NOT1 (N1774, N1754);
xor XOR2 (N1775, N1769, N1165);
and AND3 (N1776, N1766, N976, N288);
or OR4 (N1777, N1775, N264, N848, N1549);
not NOT1 (N1778, N1777);
nand NAND4 (N1779, N1774, N499, N1421, N395);
xor XOR2 (N1780, N1773, N1316);
and AND4 (N1781, N1770, N1723, N1758, N1498);
xor XOR2 (N1782, N1779, N672);
or OR2 (N1783, N1776, N654);
nand NAND3 (N1784, N1751, N131, N962);
or OR3 (N1785, N1760, N429, N623);
nor NOR2 (N1786, N1780, N569);
nand NAND3 (N1787, N1785, N1126, N602);
not NOT1 (N1788, N1787);
not NOT1 (N1789, N1786);
not NOT1 (N1790, N1765);
or OR2 (N1791, N1772, N1070);
not NOT1 (N1792, N1788);
or OR4 (N1793, N1784, N1701, N233, N1361);
nor NOR3 (N1794, N1792, N1432, N1139);
nor NOR4 (N1795, N1790, N1148, N1611, N904);
or OR2 (N1796, N1794, N1032);
or OR3 (N1797, N1782, N197, N433);
not NOT1 (N1798, N1797);
or OR2 (N1799, N1793, N1276);
and AND3 (N1800, N1798, N586, N573);
xor XOR2 (N1801, N1791, N1275);
or OR3 (N1802, N1789, N292, N956);
xor XOR2 (N1803, N1762, N1679);
not NOT1 (N1804, N1795);
not NOT1 (N1805, N1796);
nand NAND4 (N1806, N1783, N97, N276, N1554);
buf BUF1 (N1807, N1803);
and AND4 (N1808, N1799, N111, N766, N273);
and AND4 (N1809, N1805, N254, N1759, N375);
not NOT1 (N1810, N1809);
not NOT1 (N1811, N1800);
or OR3 (N1812, N1804, N1406, N1110);
xor XOR2 (N1813, N1806, N1066);
xor XOR2 (N1814, N1802, N781);
xor XOR2 (N1815, N1781, N1635);
or OR3 (N1816, N1811, N361, N158);
xor XOR2 (N1817, N1778, N980);
xor XOR2 (N1818, N1812, N1399);
nand NAND2 (N1819, N1807, N640);
and AND2 (N1820, N1818, N1417);
buf BUF1 (N1821, N1819);
or OR4 (N1822, N1814, N1540, N1077, N1245);
not NOT1 (N1823, N1820);
nor NOR2 (N1824, N1813, N105);
nand NAND3 (N1825, N1816, N536, N1085);
and AND3 (N1826, N1810, N19, N1227);
or OR4 (N1827, N1824, N1606, N6, N1752);
and AND3 (N1828, N1823, N918, N1712);
buf BUF1 (N1829, N1801);
not NOT1 (N1830, N1826);
or OR4 (N1831, N1821, N602, N725, N1767);
and AND4 (N1832, N1825, N1104, N145, N24);
not NOT1 (N1833, N1817);
buf BUF1 (N1834, N1815);
buf BUF1 (N1835, N1822);
nand NAND3 (N1836, N1828, N1300, N704);
or OR3 (N1837, N1833, N609, N1660);
nor NOR2 (N1838, N1827, N1107);
buf BUF1 (N1839, N1838);
buf BUF1 (N1840, N1836);
or OR4 (N1841, N1835, N1118, N204, N1479);
nor NOR4 (N1842, N1808, N620, N911, N131);
nand NAND4 (N1843, N1830, N1393, N1115, N38);
nor NOR2 (N1844, N1831, N1000);
xor XOR2 (N1845, N1837, N136);
xor XOR2 (N1846, N1834, N948);
nand NAND3 (N1847, N1841, N339, N119);
or OR2 (N1848, N1842, N989);
buf BUF1 (N1849, N1839);
and AND3 (N1850, N1849, N9, N1702);
nand NAND4 (N1851, N1848, N799, N1580, N709);
not NOT1 (N1852, N1840);
not NOT1 (N1853, N1832);
xor XOR2 (N1854, N1845, N1052);
buf BUF1 (N1855, N1843);
not NOT1 (N1856, N1853);
buf BUF1 (N1857, N1829);
and AND3 (N1858, N1846, N1299, N584);
and AND4 (N1859, N1850, N1543, N1619, N334);
xor XOR2 (N1860, N1855, N446);
xor XOR2 (N1861, N1844, N1674);
and AND2 (N1862, N1847, N651);
nand NAND3 (N1863, N1851, N185, N1116);
nor NOR3 (N1864, N1856, N1574, N1473);
buf BUF1 (N1865, N1861);
buf BUF1 (N1866, N1862);
and AND4 (N1867, N1857, N213, N418, N1806);
not NOT1 (N1868, N1858);
xor XOR2 (N1869, N1860, N1763);
buf BUF1 (N1870, N1867);
xor XOR2 (N1871, N1869, N404);
buf BUF1 (N1872, N1859);
nor NOR4 (N1873, N1866, N1663, N601, N436);
and AND2 (N1874, N1852, N620);
not NOT1 (N1875, N1872);
buf BUF1 (N1876, N1873);
xor XOR2 (N1877, N1868, N1070);
or OR4 (N1878, N1877, N726, N353, N69);
buf BUF1 (N1879, N1878);
buf BUF1 (N1880, N1875);
not NOT1 (N1881, N1863);
nand NAND4 (N1882, N1870, N1756, N881, N957);
and AND4 (N1883, N1882, N1641, N1550, N536);
not NOT1 (N1884, N1864);
and AND3 (N1885, N1854, N528, N1131);
nor NOR2 (N1886, N1865, N321);
buf BUF1 (N1887, N1876);
or OR4 (N1888, N1874, N224, N379, N1840);
nor NOR2 (N1889, N1871, N1501);
xor XOR2 (N1890, N1887, N733);
and AND2 (N1891, N1886, N653);
or OR4 (N1892, N1885, N1293, N1313, N1887);
not NOT1 (N1893, N1880);
nand NAND2 (N1894, N1892, N1429);
nor NOR3 (N1895, N1884, N1798, N217);
buf BUF1 (N1896, N1883);
or OR3 (N1897, N1890, N285, N869);
xor XOR2 (N1898, N1891, N1609);
not NOT1 (N1899, N1879);
nor NOR3 (N1900, N1894, N526, N11);
nor NOR3 (N1901, N1896, N1073, N237);
and AND2 (N1902, N1889, N1482);
nor NOR4 (N1903, N1897, N914, N172, N1649);
xor XOR2 (N1904, N1893, N280);
or OR4 (N1905, N1899, N105, N1872, N52);
and AND2 (N1906, N1881, N1794);
and AND3 (N1907, N1906, N1018, N1739);
or OR2 (N1908, N1901, N1798);
nand NAND4 (N1909, N1895, N1222, N866, N1004);
and AND3 (N1910, N1902, N963, N1583);
nor NOR3 (N1911, N1908, N39, N1638);
xor XOR2 (N1912, N1888, N1744);
nand NAND2 (N1913, N1903, N1802);
nor NOR3 (N1914, N1913, N207, N1226);
not NOT1 (N1915, N1900);
nand NAND2 (N1916, N1912, N440);
or OR4 (N1917, N1915, N1088, N1584, N1808);
and AND4 (N1918, N1909, N840, N1352, N1615);
not NOT1 (N1919, N1917);
or OR3 (N1920, N1919, N1248, N440);
buf BUF1 (N1921, N1910);
xor XOR2 (N1922, N1920, N683);
not NOT1 (N1923, N1898);
and AND3 (N1924, N1921, N338, N864);
not NOT1 (N1925, N1914);
buf BUF1 (N1926, N1904);
nor NOR4 (N1927, N1926, N334, N232, N333);
not NOT1 (N1928, N1925);
buf BUF1 (N1929, N1923);
not NOT1 (N1930, N1927);
and AND3 (N1931, N1911, N1563, N155);
buf BUF1 (N1932, N1907);
and AND4 (N1933, N1924, N697, N275, N152);
and AND2 (N1934, N1932, N589);
xor XOR2 (N1935, N1934, N671);
or OR4 (N1936, N1933, N1224, N1792, N1632);
and AND3 (N1937, N1928, N29, N1218);
and AND3 (N1938, N1935, N1218, N1485);
and AND3 (N1939, N1929, N705, N742);
buf BUF1 (N1940, N1918);
not NOT1 (N1941, N1940);
or OR4 (N1942, N1905, N978, N522, N1504);
xor XOR2 (N1943, N1936, N539);
nand NAND3 (N1944, N1930, N46, N496);
not NOT1 (N1945, N1916);
and AND4 (N1946, N1939, N513, N1529, N652);
buf BUF1 (N1947, N1937);
nand NAND3 (N1948, N1943, N987, N221);
nand NAND3 (N1949, N1947, N1346, N1592);
or OR3 (N1950, N1941, N1532, N1662);
nand NAND4 (N1951, N1942, N1561, N1371, N724);
buf BUF1 (N1952, N1948);
and AND4 (N1953, N1922, N1938, N529, N1218);
not NOT1 (N1954, N885);
and AND3 (N1955, N1946, N1485, N725);
or OR2 (N1956, N1950, N1575);
nor NOR4 (N1957, N1951, N13, N886, N1851);
and AND3 (N1958, N1949, N1238, N1449);
xor XOR2 (N1959, N1957, N1536);
not NOT1 (N1960, N1931);
and AND2 (N1961, N1955, N54);
not NOT1 (N1962, N1959);
not NOT1 (N1963, N1958);
nor NOR4 (N1964, N1960, N1392, N1458, N1233);
nor NOR3 (N1965, N1963, N609, N1830);
not NOT1 (N1966, N1944);
xor XOR2 (N1967, N1945, N1177);
nand NAND4 (N1968, N1965, N1410, N1370, N1126);
not NOT1 (N1969, N1962);
not NOT1 (N1970, N1966);
not NOT1 (N1971, N1956);
and AND4 (N1972, N1961, N538, N804, N609);
nand NAND4 (N1973, N1971, N1913, N1755, N555);
or OR3 (N1974, N1972, N710, N1687);
nand NAND3 (N1975, N1968, N1774, N1793);
and AND4 (N1976, N1964, N4, N1901, N1803);
buf BUF1 (N1977, N1952);
buf BUF1 (N1978, N1953);
xor XOR2 (N1979, N1976, N1498);
buf BUF1 (N1980, N1969);
xor XOR2 (N1981, N1967, N569);
and AND4 (N1982, N1981, N1404, N1359, N1423);
not NOT1 (N1983, N1982);
not NOT1 (N1984, N1978);
nand NAND2 (N1985, N1973, N1110);
and AND2 (N1986, N1977, N1089);
not NOT1 (N1987, N1954);
not NOT1 (N1988, N1984);
and AND3 (N1989, N1985, N1523, N1790);
nor NOR4 (N1990, N1974, N47, N883, N1404);
xor XOR2 (N1991, N1988, N745);
buf BUF1 (N1992, N1989);
or OR3 (N1993, N1979, N1282, N539);
or OR2 (N1994, N1987, N1977);
nor NOR2 (N1995, N1994, N1855);
or OR3 (N1996, N1990, N1462, N1830);
nor NOR3 (N1997, N1983, N1106, N1095);
xor XOR2 (N1998, N1975, N1713);
and AND2 (N1999, N1997, N651);
and AND4 (N2000, N1992, N181, N683, N246);
buf BUF1 (N2001, N1980);
and AND2 (N2002, N1995, N325);
xor XOR2 (N2003, N1970, N252);
xor XOR2 (N2004, N1993, N1080);
nor NOR2 (N2005, N1986, N1105);
not NOT1 (N2006, N2002);
nor NOR3 (N2007, N1998, N327, N1525);
nor NOR4 (N2008, N2004, N408, N1728, N1705);
xor XOR2 (N2009, N1991, N1302);
buf BUF1 (N2010, N2007);
buf BUF1 (N2011, N1996);
nor NOR2 (N2012, N1999, N915);
not NOT1 (N2013, N2008);
buf BUF1 (N2014, N2006);
and AND2 (N2015, N2000, N494);
nor NOR2 (N2016, N2001, N1013);
nand NAND3 (N2017, N2011, N1529, N1374);
nand NAND3 (N2018, N2013, N371, N1355);
buf BUF1 (N2019, N2014);
buf BUF1 (N2020, N2017);
nor NOR2 (N2021, N2005, N1235);
or OR3 (N2022, N2003, N488, N681);
and AND2 (N2023, N2016, N746);
nor NOR2 (N2024, N2012, N76);
nor NOR2 (N2025, N2019, N1833);
buf BUF1 (N2026, N2010);
xor XOR2 (N2027, N2024, N142);
not NOT1 (N2028, N2023);
buf BUF1 (N2029, N2026);
xor XOR2 (N2030, N2021, N1685);
and AND2 (N2031, N2029, N257);
xor XOR2 (N2032, N2031, N1560);
or OR2 (N2033, N2022, N1254);
not NOT1 (N2034, N2027);
nand NAND3 (N2035, N2028, N1852, N1912);
xor XOR2 (N2036, N2030, N366);
not NOT1 (N2037, N2032);
and AND4 (N2038, N2020, N1566, N452, N231);
and AND4 (N2039, N2038, N1487, N1676, N372);
xor XOR2 (N2040, N2033, N838);
xor XOR2 (N2041, N2039, N97);
nor NOR2 (N2042, N2018, N534);
nand NAND4 (N2043, N2034, N1384, N1400, N1454);
nor NOR4 (N2044, N2040, N1604, N1381, N1105);
xor XOR2 (N2045, N2042, N1963);
buf BUF1 (N2046, N2035);
nor NOR2 (N2047, N2046, N1882);
nor NOR4 (N2048, N2009, N593, N232, N1050);
nand NAND4 (N2049, N2047, N828, N771, N741);
and AND3 (N2050, N2048, N1350, N1334);
or OR3 (N2051, N2015, N428, N1054);
or OR4 (N2052, N2045, N369, N246, N619);
buf BUF1 (N2053, N2044);
nor NOR3 (N2054, N2025, N1617, N996);
or OR4 (N2055, N2051, N2047, N419, N1779);
or OR4 (N2056, N2041, N1104, N934, N74);
xor XOR2 (N2057, N2036, N1903);
not NOT1 (N2058, N2037);
nand NAND3 (N2059, N2053, N905, N1534);
or OR4 (N2060, N2050, N1220, N1206, N290);
and AND4 (N2061, N2052, N2015, N1219, N37);
and AND2 (N2062, N2060, N1005);
buf BUF1 (N2063, N2054);
nor NOR2 (N2064, N2056, N1019);
nand NAND2 (N2065, N2062, N1797);
nor NOR3 (N2066, N2064, N1749, N2054);
nor NOR3 (N2067, N2043, N11, N1951);
nand NAND2 (N2068, N2067, N1813);
and AND2 (N2069, N2049, N992);
xor XOR2 (N2070, N2068, N1453);
not NOT1 (N2071, N2058);
buf BUF1 (N2072, N2070);
buf BUF1 (N2073, N2059);
nor NOR3 (N2074, N2072, N197, N1488);
xor XOR2 (N2075, N2074, N1857);
and AND3 (N2076, N2063, N671, N1209);
nor NOR2 (N2077, N2069, N1511);
not NOT1 (N2078, N2071);
or OR4 (N2079, N2066, N100, N1823, N776);
and AND2 (N2080, N2073, N773);
not NOT1 (N2081, N2055);
nand NAND3 (N2082, N2075, N1492, N475);
xor XOR2 (N2083, N2081, N1014);
xor XOR2 (N2084, N2080, N1222);
buf BUF1 (N2085, N2061);
nand NAND4 (N2086, N2078, N343, N1014, N252);
nand NAND4 (N2087, N2065, N1233, N614, N898);
and AND4 (N2088, N2057, N1853, N96, N2044);
or OR3 (N2089, N2086, N283, N1396);
nor NOR2 (N2090, N2089, N67);
nand NAND3 (N2091, N2087, N1734, N1069);
or OR2 (N2092, N2082, N600);
or OR3 (N2093, N2088, N1942, N87);
and AND4 (N2094, N2093, N68, N1018, N940);
or OR3 (N2095, N2094, N1667, N1159);
not NOT1 (N2096, N2090);
buf BUF1 (N2097, N2091);
nor NOR3 (N2098, N2084, N1872, N1242);
not NOT1 (N2099, N2095);
xor XOR2 (N2100, N2079, N1753);
not NOT1 (N2101, N2076);
and AND4 (N2102, N2100, N858, N1147, N1868);
buf BUF1 (N2103, N2096);
nor NOR4 (N2104, N2099, N1000, N1591, N742);
xor XOR2 (N2105, N2097, N606);
not NOT1 (N2106, N2105);
buf BUF1 (N2107, N2106);
xor XOR2 (N2108, N2102, N1231);
xor XOR2 (N2109, N2077, N1407);
nor NOR4 (N2110, N2107, N1956, N1526, N1224);
and AND2 (N2111, N2103, N836);
nor NOR2 (N2112, N2101, N2057);
and AND3 (N2113, N2112, N595, N599);
xor XOR2 (N2114, N2113, N1183);
and AND4 (N2115, N2098, N830, N693, N35);
or OR3 (N2116, N2111, N539, N1726);
or OR4 (N2117, N2116, N1898, N153, N2018);
or OR2 (N2118, N2117, N1709);
buf BUF1 (N2119, N2115);
or OR2 (N2120, N2104, N1045);
nand NAND2 (N2121, N2109, N1372);
or OR3 (N2122, N2083, N1111, N1658);
or OR4 (N2123, N2114, N257, N1167, N404);
or OR2 (N2124, N2121, N677);
buf BUF1 (N2125, N2092);
or OR4 (N2126, N2123, N1981, N989, N1848);
nand NAND3 (N2127, N2125, N1633, N2100);
nand NAND3 (N2128, N2127, N621, N1139);
buf BUF1 (N2129, N2124);
nor NOR3 (N2130, N2122, N1458, N1082);
or OR3 (N2131, N2128, N1358, N416);
or OR4 (N2132, N2085, N2024, N889, N1938);
or OR4 (N2133, N2131, N204, N556, N1772);
nand NAND3 (N2134, N2126, N1171, N887);
nand NAND3 (N2135, N2132, N656, N1764);
buf BUF1 (N2136, N2108);
not NOT1 (N2137, N2129);
xor XOR2 (N2138, N2137, N1707);
nand NAND4 (N2139, N2138, N577, N20, N1306);
nor NOR2 (N2140, N2135, N350);
nand NAND3 (N2141, N2130, N687, N1593);
buf BUF1 (N2142, N2110);
or OR2 (N2143, N2133, N402);
not NOT1 (N2144, N2139);
and AND4 (N2145, N2141, N2128, N1078, N1158);
xor XOR2 (N2146, N2120, N2023);
nand NAND4 (N2147, N2142, N1022, N418, N428);
not NOT1 (N2148, N2144);
xor XOR2 (N2149, N2136, N287);
nor NOR4 (N2150, N2143, N2083, N855, N1650);
nand NAND4 (N2151, N2140, N544, N1092, N519);
not NOT1 (N2152, N2149);
and AND3 (N2153, N2152, N83, N649);
and AND2 (N2154, N2147, N1513);
buf BUF1 (N2155, N2151);
buf BUF1 (N2156, N2153);
buf BUF1 (N2157, N2146);
nand NAND2 (N2158, N2145, N1980);
xor XOR2 (N2159, N2158, N456);
or OR2 (N2160, N2157, N72);
nand NAND2 (N2161, N2119, N1015);
buf BUF1 (N2162, N2150);
nor NOR4 (N2163, N2154, N585, N392, N2016);
not NOT1 (N2164, N2134);
and AND4 (N2165, N2163, N1381, N558, N1131);
or OR2 (N2166, N2164, N108);
nand NAND3 (N2167, N2166, N1603, N1312);
buf BUF1 (N2168, N2156);
xor XOR2 (N2169, N2165, N1573);
or OR2 (N2170, N2161, N812);
nand NAND2 (N2171, N2155, N2061);
xor XOR2 (N2172, N2170, N1517);
buf BUF1 (N2173, N2118);
nand NAND4 (N2174, N2167, N2162, N1957, N1756);
nand NAND4 (N2175, N983, N1277, N1175, N600);
or OR2 (N2176, N2168, N1288);
nand NAND3 (N2177, N2160, N396, N2068);
and AND3 (N2178, N2148, N893, N1203);
xor XOR2 (N2179, N2169, N722);
and AND3 (N2180, N2178, N183, N902);
nand NAND2 (N2181, N2173, N1130);
or OR4 (N2182, N2179, N256, N261, N1758);
xor XOR2 (N2183, N2181, N1834);
xor XOR2 (N2184, N2171, N92);
buf BUF1 (N2185, N2184);
not NOT1 (N2186, N2176);
or OR4 (N2187, N2185, N1660, N1558, N358);
not NOT1 (N2188, N2187);
not NOT1 (N2189, N2180);
and AND3 (N2190, N2172, N1064, N306);
xor XOR2 (N2191, N2177, N303);
not NOT1 (N2192, N2159);
xor XOR2 (N2193, N2192, N1315);
buf BUF1 (N2194, N2174);
nor NOR3 (N2195, N2186, N2177, N625);
xor XOR2 (N2196, N2191, N2);
not NOT1 (N2197, N2189);
and AND2 (N2198, N2194, N1089);
buf BUF1 (N2199, N2198);
nor NOR4 (N2200, N2190, N744, N1433, N973);
and AND4 (N2201, N2188, N1082, N1710, N1320);
or OR3 (N2202, N2200, N791, N1889);
and AND2 (N2203, N2183, N1241);
not NOT1 (N2204, N2193);
and AND2 (N2205, N2203, N1085);
nor NOR4 (N2206, N2197, N802, N1374, N1374);
nor NOR2 (N2207, N2182, N2124);
or OR4 (N2208, N2207, N1874, N1119, N872);
buf BUF1 (N2209, N2199);
not NOT1 (N2210, N2196);
or OR3 (N2211, N2202, N872, N550);
and AND2 (N2212, N2209, N2156);
nand NAND2 (N2213, N2208, N637);
and AND3 (N2214, N2213, N1157, N1751);
buf BUF1 (N2215, N2211);
nand NAND4 (N2216, N2204, N1348, N2135, N922);
nand NAND3 (N2217, N2215, N1623, N723);
nand NAND4 (N2218, N2201, N1195, N2181, N2108);
or OR4 (N2219, N2214, N1678, N2140, N170);
nor NOR4 (N2220, N2217, N1538, N1728, N199);
not NOT1 (N2221, N2175);
or OR3 (N2222, N2219, N1095, N367);
buf BUF1 (N2223, N2218);
buf BUF1 (N2224, N2210);
buf BUF1 (N2225, N2224);
or OR2 (N2226, N2222, N1479);
not NOT1 (N2227, N2212);
and AND2 (N2228, N2225, N39);
nor NOR3 (N2229, N2228, N1617, N1919);
buf BUF1 (N2230, N2195);
buf BUF1 (N2231, N2221);
nand NAND4 (N2232, N2216, N380, N660, N95);
nand NAND3 (N2233, N2229, N370, N1893);
buf BUF1 (N2234, N2231);
or OR4 (N2235, N2234, N2135, N329, N995);
nand NAND4 (N2236, N2235, N289, N99, N2219);
buf BUF1 (N2237, N2223);
xor XOR2 (N2238, N2206, N73);
nor NOR4 (N2239, N2238, N1902, N1968, N423);
or OR3 (N2240, N2227, N14, N71);
not NOT1 (N2241, N2226);
nor NOR4 (N2242, N2240, N417, N825, N1705);
nor NOR4 (N2243, N2242, N316, N1132, N1045);
nor NOR3 (N2244, N2205, N150, N2178);
not NOT1 (N2245, N2243);
or OR3 (N2246, N2237, N1048, N475);
buf BUF1 (N2247, N2236);
and AND4 (N2248, N2244, N1651, N1979, N206);
xor XOR2 (N2249, N2248, N379);
or OR2 (N2250, N2233, N1596);
buf BUF1 (N2251, N2247);
or OR3 (N2252, N2249, N1844, N393);
xor XOR2 (N2253, N2220, N1287);
and AND2 (N2254, N2251, N1012);
not NOT1 (N2255, N2241);
or OR2 (N2256, N2230, N1856);
nor NOR4 (N2257, N2256, N1913, N64, N1875);
and AND3 (N2258, N2252, N249, N1839);
nand NAND2 (N2259, N2258, N2241);
xor XOR2 (N2260, N2259, N1008);
buf BUF1 (N2261, N2253);
and AND3 (N2262, N2246, N907, N1281);
buf BUF1 (N2263, N2257);
and AND4 (N2264, N2262, N773, N117, N797);
or OR4 (N2265, N2264, N1316, N2232, N600);
nand NAND4 (N2266, N1958, N207, N138, N641);
nor NOR2 (N2267, N2260, N893);
not NOT1 (N2268, N2254);
xor XOR2 (N2269, N2255, N549);
or OR2 (N2270, N2265, N1475);
or OR2 (N2271, N2239, N614);
not NOT1 (N2272, N2261);
nor NOR2 (N2273, N2272, N1020);
nand NAND2 (N2274, N2263, N912);
nand NAND4 (N2275, N2270, N1060, N1666, N826);
or OR3 (N2276, N2245, N1802, N1468);
or OR4 (N2277, N2273, N222, N925, N1028);
buf BUF1 (N2278, N2271);
not NOT1 (N2279, N2277);
buf BUF1 (N2280, N2274);
or OR4 (N2281, N2267, N1568, N1318, N288);
nand NAND3 (N2282, N2276, N950, N1517);
or OR2 (N2283, N2278, N335);
not NOT1 (N2284, N2266);
not NOT1 (N2285, N2279);
xor XOR2 (N2286, N2284, N64);
nand NAND3 (N2287, N2281, N123, N880);
nor NOR2 (N2288, N2268, N1672);
buf BUF1 (N2289, N2269);
not NOT1 (N2290, N2250);
and AND4 (N2291, N2289, N2040, N1404, N496);
not NOT1 (N2292, N2282);
not NOT1 (N2293, N2291);
and AND4 (N2294, N2283, N444, N143, N906);
buf BUF1 (N2295, N2287);
buf BUF1 (N2296, N2285);
buf BUF1 (N2297, N2292);
buf BUF1 (N2298, N2290);
and AND4 (N2299, N2288, N342, N1127, N736);
not NOT1 (N2300, N2280);
and AND3 (N2301, N2275, N2273, N1519);
buf BUF1 (N2302, N2293);
nand NAND3 (N2303, N2301, N349, N1983);
nor NOR4 (N2304, N2300, N447, N577, N1085);
buf BUF1 (N2305, N2302);
not NOT1 (N2306, N2294);
nor NOR2 (N2307, N2298, N1422);
xor XOR2 (N2308, N2295, N1878);
buf BUF1 (N2309, N2299);
or OR4 (N2310, N2304, N81, N2073, N1319);
nand NAND3 (N2311, N2303, N1951, N432);
or OR2 (N2312, N2297, N16);
not NOT1 (N2313, N2311);
and AND2 (N2314, N2312, N772);
or OR4 (N2315, N2310, N1118, N951, N717);
nor NOR4 (N2316, N2305, N1402, N315, N618);
and AND3 (N2317, N2316, N442, N1684);
xor XOR2 (N2318, N2286, N1675);
or OR2 (N2319, N2306, N1105);
nor NOR3 (N2320, N2317, N1425, N1368);
xor XOR2 (N2321, N2320, N1345);
not NOT1 (N2322, N2296);
not NOT1 (N2323, N2308);
xor XOR2 (N2324, N2314, N1967);
nand NAND2 (N2325, N2324, N1833);
xor XOR2 (N2326, N2325, N1338);
and AND3 (N2327, N2326, N114, N261);
and AND4 (N2328, N2318, N2024, N1105, N717);
nand NAND2 (N2329, N2315, N200);
and AND3 (N2330, N2323, N1494, N990);
nor NOR2 (N2331, N2327, N2);
nor NOR4 (N2332, N2307, N2111, N1694, N2105);
nand NAND4 (N2333, N2330, N232, N990, N1412);
nand NAND2 (N2334, N2332, N120);
buf BUF1 (N2335, N2322);
nor NOR3 (N2336, N2321, N1564, N1151);
xor XOR2 (N2337, N2313, N1611);
or OR3 (N2338, N2319, N1690, N2126);
not NOT1 (N2339, N2333);
and AND3 (N2340, N2338, N2122, N30);
and AND3 (N2341, N2339, N772, N196);
nand NAND3 (N2342, N2328, N1579, N18);
and AND4 (N2343, N2309, N566, N427, N675);
or OR3 (N2344, N2334, N1646, N1116);
or OR2 (N2345, N2342, N775);
or OR3 (N2346, N2337, N1998, N661);
or OR3 (N2347, N2344, N153, N386);
nor NOR2 (N2348, N2346, N1293);
nand NAND4 (N2349, N2340, N2029, N1367, N1680);
not NOT1 (N2350, N2347);
xor XOR2 (N2351, N2341, N1652);
not NOT1 (N2352, N2343);
not NOT1 (N2353, N2352);
and AND3 (N2354, N2349, N276, N826);
not NOT1 (N2355, N2331);
or OR3 (N2356, N2329, N1151, N1968);
and AND3 (N2357, N2351, N1559, N38);
buf BUF1 (N2358, N2357);
buf BUF1 (N2359, N2335);
or OR4 (N2360, N2356, N199, N78, N1686);
xor XOR2 (N2361, N2348, N1423);
buf BUF1 (N2362, N2353);
or OR2 (N2363, N2360, N2324);
xor XOR2 (N2364, N2350, N238);
nand NAND3 (N2365, N2362, N555, N59);
nand NAND2 (N2366, N2361, N411);
and AND2 (N2367, N2345, N1647);
buf BUF1 (N2368, N2355);
and AND2 (N2369, N2363, N423);
xor XOR2 (N2370, N2365, N1706);
buf BUF1 (N2371, N2370);
and AND4 (N2372, N2354, N1894, N558, N1125);
nor NOR4 (N2373, N2367, N905, N374, N1441);
or OR2 (N2374, N2369, N2150);
buf BUF1 (N2375, N2368);
not NOT1 (N2376, N2371);
nand NAND3 (N2377, N2373, N1965, N1775);
or OR4 (N2378, N2366, N874, N1967, N457);
buf BUF1 (N2379, N2358);
nand NAND2 (N2380, N2377, N1102);
xor XOR2 (N2381, N2376, N1124);
nor NOR3 (N2382, N2374, N746, N1412);
not NOT1 (N2383, N2372);
nand NAND4 (N2384, N2359, N1457, N1112, N17);
buf BUF1 (N2385, N2375);
not NOT1 (N2386, N2384);
xor XOR2 (N2387, N2386, N1164);
nand NAND2 (N2388, N2387, N502);
or OR3 (N2389, N2382, N466, N941);
nor NOR3 (N2390, N2389, N1854, N2187);
nor NOR4 (N2391, N2381, N1934, N1948, N247);
or OR4 (N2392, N2364, N1637, N813, N1913);
nor NOR3 (N2393, N2379, N1398, N825);
nor NOR2 (N2394, N2385, N78);
nor NOR3 (N2395, N2378, N2392, N1782);
nand NAND3 (N2396, N2085, N1641, N1929);
and AND3 (N2397, N2390, N140, N1060);
xor XOR2 (N2398, N2391, N1112);
and AND3 (N2399, N2393, N1876, N383);
or OR4 (N2400, N2388, N396, N899, N1369);
nor NOR2 (N2401, N2380, N475);
or OR4 (N2402, N2399, N12, N528, N1711);
xor XOR2 (N2403, N2394, N1656);
or OR3 (N2404, N2397, N1459, N1417);
buf BUF1 (N2405, N2398);
nor NOR4 (N2406, N2403, N1864, N10, N1673);
not NOT1 (N2407, N2395);
and AND2 (N2408, N2405, N950);
nand NAND2 (N2409, N2383, N1591);
nor NOR4 (N2410, N2400, N2119, N2218, N26);
nand NAND2 (N2411, N2406, N1530);
xor XOR2 (N2412, N2407, N1275);
xor XOR2 (N2413, N2404, N1232);
not NOT1 (N2414, N2412);
buf BUF1 (N2415, N2410);
not NOT1 (N2416, N2411);
or OR4 (N2417, N2409, N700, N807, N627);
and AND4 (N2418, N2401, N1365, N908, N1077);
not NOT1 (N2419, N2336);
buf BUF1 (N2420, N2419);
buf BUF1 (N2421, N2402);
nand NAND4 (N2422, N2417, N375, N1768, N1044);
xor XOR2 (N2423, N2413, N1232);
nand NAND2 (N2424, N2396, N1043);
nand NAND2 (N2425, N2416, N1599);
and AND4 (N2426, N2418, N806, N1888, N1873);
nand NAND4 (N2427, N2426, N1183, N2215, N2338);
and AND3 (N2428, N2425, N872, N1627);
not NOT1 (N2429, N2420);
buf BUF1 (N2430, N2421);
not NOT1 (N2431, N2424);
buf BUF1 (N2432, N2408);
nand NAND4 (N2433, N2422, N2176, N454, N776);
not NOT1 (N2434, N2429);
nand NAND4 (N2435, N2428, N1162, N976, N1537);
or OR3 (N2436, N2423, N467, N1832);
nand NAND4 (N2437, N2432, N1013, N2434, N1902);
nand NAND2 (N2438, N189, N641);
not NOT1 (N2439, N2433);
not NOT1 (N2440, N2438);
nand NAND4 (N2441, N2439, N161, N330, N2231);
and AND2 (N2442, N2427, N1104);
and AND3 (N2443, N2441, N1214, N761);
nor NOR3 (N2444, N2415, N2168, N1919);
and AND3 (N2445, N2414, N1936, N1629);
and AND3 (N2446, N2437, N1412, N878);
xor XOR2 (N2447, N2436, N286);
nor NOR4 (N2448, N2443, N1152, N2424, N2298);
buf BUF1 (N2449, N2445);
not NOT1 (N2450, N2444);
and AND3 (N2451, N2447, N253, N159);
nand NAND4 (N2452, N2449, N1843, N624, N1669);
nand NAND4 (N2453, N2448, N1353, N1679, N604);
nor NOR2 (N2454, N2451, N497);
xor XOR2 (N2455, N2435, N523);
or OR4 (N2456, N2450, N1279, N2352, N265);
not NOT1 (N2457, N2456);
or OR3 (N2458, N2446, N748, N1854);
buf BUF1 (N2459, N2440);
xor XOR2 (N2460, N2452, N240);
buf BUF1 (N2461, N2460);
nand NAND2 (N2462, N2442, N2217);
xor XOR2 (N2463, N2455, N169);
buf BUF1 (N2464, N2430);
nor NOR2 (N2465, N2458, N2140);
and AND2 (N2466, N2464, N272);
xor XOR2 (N2467, N2459, N519);
buf BUF1 (N2468, N2461);
xor XOR2 (N2469, N2465, N967);
or OR2 (N2470, N2453, N1182);
xor XOR2 (N2471, N2467, N1218);
buf BUF1 (N2472, N2457);
and AND4 (N2473, N2469, N834, N2083, N1626);
not NOT1 (N2474, N2466);
buf BUF1 (N2475, N2454);
xor XOR2 (N2476, N2470, N2225);
xor XOR2 (N2477, N2473, N1700);
xor XOR2 (N2478, N2476, N339);
or OR3 (N2479, N2474, N1093, N1950);
xor XOR2 (N2480, N2471, N1212);
not NOT1 (N2481, N2468);
xor XOR2 (N2482, N2480, N2076);
buf BUF1 (N2483, N2481);
nand NAND2 (N2484, N2472, N1819);
not NOT1 (N2485, N2462);
not NOT1 (N2486, N2479);
nor NOR3 (N2487, N2478, N504, N1176);
nand NAND4 (N2488, N2487, N1873, N1911, N2085);
not NOT1 (N2489, N2482);
or OR2 (N2490, N2483, N1977);
xor XOR2 (N2491, N2486, N181);
xor XOR2 (N2492, N2485, N2399);
not NOT1 (N2493, N2492);
nand NAND3 (N2494, N2490, N1614, N426);
xor XOR2 (N2495, N2463, N1876);
not NOT1 (N2496, N2488);
or OR3 (N2497, N2431, N341, N634);
or OR3 (N2498, N2497, N2319, N394);
or OR2 (N2499, N2491, N1418);
nor NOR3 (N2500, N2477, N792, N1665);
xor XOR2 (N2501, N2475, N1862);
not NOT1 (N2502, N2501);
buf BUF1 (N2503, N2496);
nor NOR2 (N2504, N2503, N1205);
and AND3 (N2505, N2500, N71, N1529);
xor XOR2 (N2506, N2504, N1545);
buf BUF1 (N2507, N2506);
and AND2 (N2508, N2507, N1237);
and AND3 (N2509, N2498, N663, N1669);
nand NAND3 (N2510, N2499, N83, N1356);
not NOT1 (N2511, N2502);
nor NOR2 (N2512, N2489, N1976);
and AND4 (N2513, N2484, N1253, N1306, N2252);
or OR2 (N2514, N2505, N2339);
not NOT1 (N2515, N2511);
nor NOR3 (N2516, N2513, N347, N681);
not NOT1 (N2517, N2509);
or OR3 (N2518, N2515, N249, N1641);
nor NOR2 (N2519, N2514, N2099);
and AND2 (N2520, N2510, N769);
nand NAND2 (N2521, N2518, N69);
not NOT1 (N2522, N2495);
xor XOR2 (N2523, N2494, N819);
buf BUF1 (N2524, N2522);
nor NOR4 (N2525, N2519, N2178, N315, N1927);
nor NOR4 (N2526, N2493, N612, N637, N262);
or OR3 (N2527, N2523, N582, N2199);
nand NAND3 (N2528, N2508, N2363, N1400);
nand NAND4 (N2529, N2520, N141, N2091, N837);
xor XOR2 (N2530, N2517, N1094);
or OR2 (N2531, N2516, N83);
or OR4 (N2532, N2527, N2352, N1836, N965);
not NOT1 (N2533, N2528);
not NOT1 (N2534, N2531);
buf BUF1 (N2535, N2526);
buf BUF1 (N2536, N2533);
nor NOR3 (N2537, N2524, N1136, N88);
or OR2 (N2538, N2512, N501);
or OR2 (N2539, N2521, N602);
nand NAND4 (N2540, N2538, N1105, N400, N293);
buf BUF1 (N2541, N2530);
nand NAND2 (N2542, N2535, N1029);
nor NOR2 (N2543, N2529, N474);
or OR3 (N2544, N2537, N581, N2024);
not NOT1 (N2545, N2534);
xor XOR2 (N2546, N2545, N937);
and AND2 (N2547, N2532, N1234);
or OR2 (N2548, N2540, N2533);
xor XOR2 (N2549, N2539, N361);
or OR3 (N2550, N2541, N2023, N1469);
nand NAND3 (N2551, N2536, N1667, N1638);
and AND3 (N2552, N2548, N827, N1019);
nor NOR2 (N2553, N2551, N1229);
and AND3 (N2554, N2547, N907, N2283);
buf BUF1 (N2555, N2542);
not NOT1 (N2556, N2554);
nand NAND2 (N2557, N2544, N833);
and AND2 (N2558, N2550, N159);
nand NAND3 (N2559, N2525, N2102, N2427);
not NOT1 (N2560, N2555);
buf BUF1 (N2561, N2543);
not NOT1 (N2562, N2552);
xor XOR2 (N2563, N2553, N1037);
xor XOR2 (N2564, N2556, N2409);
nor NOR4 (N2565, N2557, N1319, N754, N1579);
nand NAND4 (N2566, N2564, N272, N905, N801);
nor NOR2 (N2567, N2546, N547);
or OR3 (N2568, N2558, N508, N2092);
nor NOR2 (N2569, N2563, N1434);
and AND2 (N2570, N2566, N991);
not NOT1 (N2571, N2559);
xor XOR2 (N2572, N2567, N847);
nor NOR3 (N2573, N2570, N1802, N395);
buf BUF1 (N2574, N2568);
or OR2 (N2575, N2565, N83);
and AND3 (N2576, N2560, N2097, N214);
nand NAND4 (N2577, N2575, N574, N2246, N2436);
xor XOR2 (N2578, N2572, N1171);
nand NAND3 (N2579, N2561, N2536, N61);
not NOT1 (N2580, N2576);
nand NAND4 (N2581, N2579, N2252, N478, N555);
buf BUF1 (N2582, N2580);
and AND3 (N2583, N2574, N1449, N1888);
or OR3 (N2584, N2582, N1777, N1208);
nand NAND4 (N2585, N2583, N1545, N1682, N1838);
xor XOR2 (N2586, N2581, N1949);
or OR3 (N2587, N2578, N423, N1809);
nand NAND3 (N2588, N2585, N284, N476);
nand NAND2 (N2589, N2571, N2428);
not NOT1 (N2590, N2562);
xor XOR2 (N2591, N2549, N1000);
nand NAND4 (N2592, N2589, N1720, N2380, N712);
buf BUF1 (N2593, N2573);
buf BUF1 (N2594, N2569);
xor XOR2 (N2595, N2584, N1336);
not NOT1 (N2596, N2577);
nand NAND3 (N2597, N2587, N1720, N1384);
or OR2 (N2598, N2594, N1445);
xor XOR2 (N2599, N2593, N2594);
buf BUF1 (N2600, N2591);
nor NOR4 (N2601, N2599, N878, N1039, N1037);
and AND3 (N2602, N2596, N2490, N1000);
buf BUF1 (N2603, N2586);
nor NOR3 (N2604, N2602, N1685, N750);
buf BUF1 (N2605, N2603);
or OR2 (N2606, N2605, N1162);
or OR3 (N2607, N2588, N2172, N2528);
nand NAND4 (N2608, N2595, N1674, N1331, N88);
not NOT1 (N2609, N2604);
xor XOR2 (N2610, N2592, N1213);
or OR4 (N2611, N2597, N19, N2556, N1327);
and AND4 (N2612, N2608, N481, N163, N1184);
nor NOR2 (N2613, N2609, N1982);
buf BUF1 (N2614, N2600);
nor NOR3 (N2615, N2601, N690, N1879);
nand NAND3 (N2616, N2613, N785, N532);
nor NOR3 (N2617, N2614, N2359, N1077);
nand NAND3 (N2618, N2615, N221, N1958);
and AND3 (N2619, N2616, N1786, N1474);
xor XOR2 (N2620, N2617, N653);
or OR2 (N2621, N2619, N2419);
nor NOR4 (N2622, N2598, N1095, N1484, N1542);
buf BUF1 (N2623, N2590);
not NOT1 (N2624, N2612);
nand NAND3 (N2625, N2610, N2209, N1486);
and AND3 (N2626, N2622, N2153, N592);
nor NOR3 (N2627, N2621, N683, N55);
nor NOR3 (N2628, N2611, N535, N378);
xor XOR2 (N2629, N2624, N1736);
and AND4 (N2630, N2620, N2297, N2546, N1896);
not NOT1 (N2631, N2623);
xor XOR2 (N2632, N2631, N528);
not NOT1 (N2633, N2606);
or OR2 (N2634, N2629, N1213);
xor XOR2 (N2635, N2628, N823);
or OR3 (N2636, N2626, N1736, N2628);
or OR3 (N2637, N2636, N362, N675);
not NOT1 (N2638, N2633);
nand NAND4 (N2639, N2627, N234, N71, N2510);
or OR4 (N2640, N2630, N1889, N186, N621);
nand NAND2 (N2641, N2638, N1411);
not NOT1 (N2642, N2618);
not NOT1 (N2643, N2635);
buf BUF1 (N2644, N2643);
and AND3 (N2645, N2637, N163, N557);
or OR4 (N2646, N2641, N463, N611, N655);
nand NAND2 (N2647, N2640, N2618);
xor XOR2 (N2648, N2645, N1268);
buf BUF1 (N2649, N2648);
or OR3 (N2650, N2647, N1803, N1333);
and AND2 (N2651, N2646, N1873);
and AND4 (N2652, N2642, N919, N760, N2154);
and AND3 (N2653, N2651, N1342, N2242);
nand NAND4 (N2654, N2632, N1331, N1307, N305);
buf BUF1 (N2655, N2653);
xor XOR2 (N2656, N2644, N1694);
xor XOR2 (N2657, N2652, N2572);
not NOT1 (N2658, N2656);
buf BUF1 (N2659, N2649);
buf BUF1 (N2660, N2625);
buf BUF1 (N2661, N2658);
xor XOR2 (N2662, N2655, N193);
nor NOR2 (N2663, N2634, N379);
nand NAND2 (N2664, N2661, N1304);
not NOT1 (N2665, N2659);
xor XOR2 (N2666, N2663, N1229);
nand NAND2 (N2667, N2657, N267);
not NOT1 (N2668, N2639);
nor NOR3 (N2669, N2666, N418, N1253);
nor NOR2 (N2670, N2669, N2494);
nor NOR3 (N2671, N2667, N91, N232);
not NOT1 (N2672, N2671);
or OR2 (N2673, N2664, N2089);
buf BUF1 (N2674, N2662);
nor NOR2 (N2675, N2607, N1795);
buf BUF1 (N2676, N2672);
nand NAND3 (N2677, N2674, N2511, N1352);
xor XOR2 (N2678, N2670, N1343);
or OR3 (N2679, N2665, N1095, N1444);
nor NOR3 (N2680, N2677, N1664, N1547);
or OR4 (N2681, N2675, N372, N999, N1760);
buf BUF1 (N2682, N2673);
nand NAND2 (N2683, N2668, N2470);
and AND2 (N2684, N2660, N2490);
xor XOR2 (N2685, N2654, N466);
xor XOR2 (N2686, N2679, N595);
not NOT1 (N2687, N2650);
and AND3 (N2688, N2683, N2292, N1361);
not NOT1 (N2689, N2681);
buf BUF1 (N2690, N2676);
not NOT1 (N2691, N2684);
or OR3 (N2692, N2682, N738, N1291);
xor XOR2 (N2693, N2685, N1082);
xor XOR2 (N2694, N2690, N1154);
or OR2 (N2695, N2689, N53);
nand NAND4 (N2696, N2686, N719, N2025, N1668);
buf BUF1 (N2697, N2691);
nand NAND3 (N2698, N2696, N1024, N781);
buf BUF1 (N2699, N2678);
and AND4 (N2700, N2698, N1542, N1756, N699);
or OR4 (N2701, N2692, N1027, N107, N812);
nand NAND2 (N2702, N2695, N830);
buf BUF1 (N2703, N2694);
and AND2 (N2704, N2703, N2325);
nand NAND4 (N2705, N2697, N578, N1513, N2166);
and AND2 (N2706, N2687, N1998);
xor XOR2 (N2707, N2706, N1233);
or OR3 (N2708, N2707, N2322, N496);
and AND4 (N2709, N2680, N2251, N519, N949);
not NOT1 (N2710, N2700);
or OR3 (N2711, N2710, N1174, N1042);
buf BUF1 (N2712, N2701);
nand NAND4 (N2713, N2708, N1976, N1180, N1988);
nor NOR3 (N2714, N2688, N1219, N1736);
and AND3 (N2715, N2704, N9, N2567);
not NOT1 (N2716, N2714);
not NOT1 (N2717, N2702);
buf BUF1 (N2718, N2693);
nor NOR3 (N2719, N2718, N2120, N1258);
nor NOR4 (N2720, N2717, N2083, N425, N1011);
xor XOR2 (N2721, N2699, N558);
buf BUF1 (N2722, N2721);
or OR4 (N2723, N2719, N2535, N2467, N1700);
nand NAND2 (N2724, N2715, N353);
or OR4 (N2725, N2709, N723, N1903, N1305);
xor XOR2 (N2726, N2711, N1438);
nand NAND3 (N2727, N2716, N878, N613);
not NOT1 (N2728, N2722);
nor NOR4 (N2729, N2725, N1786, N686, N2462);
not NOT1 (N2730, N2728);
not NOT1 (N2731, N2712);
nand NAND2 (N2732, N2731, N937);
not NOT1 (N2733, N2713);
xor XOR2 (N2734, N2733, N2386);
or OR4 (N2735, N2705, N1656, N1715, N1593);
not NOT1 (N2736, N2730);
nand NAND2 (N2737, N2723, N235);
nor NOR2 (N2738, N2735, N623);
nor NOR2 (N2739, N2724, N2698);
or OR4 (N2740, N2737, N2051, N1634, N1011);
nor NOR4 (N2741, N2738, N217, N2009, N1210);
or OR4 (N2742, N2740, N194, N1172, N1713);
xor XOR2 (N2743, N2742, N755);
nor NOR4 (N2744, N2732, N1720, N1836, N1600);
not NOT1 (N2745, N2734);
or OR2 (N2746, N2739, N1452);
or OR2 (N2747, N2741, N1911);
and AND2 (N2748, N2747, N220);
or OR4 (N2749, N2743, N2551, N933, N396);
nor NOR2 (N2750, N2727, N689);
buf BUF1 (N2751, N2746);
buf BUF1 (N2752, N2729);
nand NAND2 (N2753, N2749, N2023);
not NOT1 (N2754, N2726);
or OR2 (N2755, N2751, N170);
buf BUF1 (N2756, N2753);
or OR2 (N2757, N2756, N2432);
or OR4 (N2758, N2748, N683, N1774, N2529);
and AND3 (N2759, N2736, N1575, N170);
nand NAND2 (N2760, N2744, N2259);
xor XOR2 (N2761, N2759, N1109);
nand NAND4 (N2762, N2752, N55, N2125, N1136);
nor NOR3 (N2763, N2750, N93, N1575);
buf BUF1 (N2764, N2762);
nor NOR2 (N2765, N2761, N2222);
or OR3 (N2766, N2765, N429, N973);
buf BUF1 (N2767, N2764);
buf BUF1 (N2768, N2757);
nand NAND3 (N2769, N2763, N1835, N662);
xor XOR2 (N2770, N2758, N552);
and AND4 (N2771, N2767, N574, N820, N2280);
nor NOR3 (N2772, N2755, N2371, N976);
or OR4 (N2773, N2754, N1234, N2564, N1816);
xor XOR2 (N2774, N2770, N591);
nor NOR4 (N2775, N2768, N765, N1777, N1398);
and AND4 (N2776, N2774, N2704, N1429, N1296);
nor NOR3 (N2777, N2771, N1545, N874);
and AND3 (N2778, N2769, N955, N1667);
xor XOR2 (N2779, N2777, N1489);
xor XOR2 (N2780, N2760, N2212);
nor NOR4 (N2781, N2720, N1801, N1562, N1283);
not NOT1 (N2782, N2773);
xor XOR2 (N2783, N2766, N546);
buf BUF1 (N2784, N2783);
not NOT1 (N2785, N2780);
and AND3 (N2786, N2779, N1715, N1094);
buf BUF1 (N2787, N2745);
nor NOR4 (N2788, N2782, N1511, N1427, N2776);
buf BUF1 (N2789, N221);
xor XOR2 (N2790, N2778, N2170);
or OR3 (N2791, N2781, N99, N2329);
and AND3 (N2792, N2791, N727, N723);
buf BUF1 (N2793, N2775);
xor XOR2 (N2794, N2789, N1295);
xor XOR2 (N2795, N2785, N2188);
not NOT1 (N2796, N2790);
buf BUF1 (N2797, N2794);
and AND4 (N2798, N2796, N1300, N167, N2405);
nand NAND4 (N2799, N2798, N1780, N2393, N362);
and AND4 (N2800, N2793, N2316, N1160, N1315);
or OR3 (N2801, N2788, N685, N1039);
not NOT1 (N2802, N2792);
buf BUF1 (N2803, N2787);
or OR2 (N2804, N2795, N1953);
and AND3 (N2805, N2804, N2445, N427);
and AND2 (N2806, N2802, N1542);
and AND4 (N2807, N2801, N2509, N1226, N1130);
nand NAND3 (N2808, N2799, N1300, N1685);
buf BUF1 (N2809, N2808);
and AND3 (N2810, N2806, N380, N2417);
and AND2 (N2811, N2797, N2140);
nand NAND4 (N2812, N2786, N2709, N1660, N1272);
and AND4 (N2813, N2809, N2613, N211, N1976);
nor NOR3 (N2814, N2811, N540, N1537);
nor NOR3 (N2815, N2784, N2578, N715);
or OR2 (N2816, N2810, N1406);
nor NOR3 (N2817, N2800, N2589, N827);
or OR3 (N2818, N2807, N750, N1866);
xor XOR2 (N2819, N2815, N1092);
nor NOR4 (N2820, N2812, N2413, N1609, N2458);
nand NAND4 (N2821, N2818, N64, N2260, N2408);
not NOT1 (N2822, N2821);
and AND4 (N2823, N2803, N9, N1361, N632);
nor NOR4 (N2824, N2817, N1102, N1949, N992);
xor XOR2 (N2825, N2814, N2814);
buf BUF1 (N2826, N2823);
xor XOR2 (N2827, N2805, N1767);
not NOT1 (N2828, N2816);
and AND2 (N2829, N2772, N296);
or OR3 (N2830, N2826, N945, N1484);
nor NOR4 (N2831, N2825, N1068, N2170, N2233);
buf BUF1 (N2832, N2830);
buf BUF1 (N2833, N2828);
xor XOR2 (N2834, N2820, N929);
not NOT1 (N2835, N2819);
not NOT1 (N2836, N2824);
nand NAND2 (N2837, N2822, N827);
not NOT1 (N2838, N2833);
and AND4 (N2839, N2831, N2048, N591, N2674);
nor NOR4 (N2840, N2834, N1918, N1254, N2329);
or OR3 (N2841, N2832, N1401, N2524);
xor XOR2 (N2842, N2839, N470);
buf BUF1 (N2843, N2827);
nor NOR3 (N2844, N2842, N1974, N126);
or OR2 (N2845, N2840, N1401);
or OR2 (N2846, N2843, N2559);
and AND3 (N2847, N2836, N2758, N1455);
xor XOR2 (N2848, N2829, N311);
buf BUF1 (N2849, N2837);
not NOT1 (N2850, N2846);
xor XOR2 (N2851, N2845, N2396);
or OR4 (N2852, N2841, N2797, N1104, N1927);
not NOT1 (N2853, N2844);
or OR3 (N2854, N2813, N27, N2310);
nor NOR4 (N2855, N2850, N2347, N470, N365);
not NOT1 (N2856, N2853);
nand NAND2 (N2857, N2849, N1179);
buf BUF1 (N2858, N2847);
and AND4 (N2859, N2854, N2156, N2264, N2633);
buf BUF1 (N2860, N2855);
or OR3 (N2861, N2852, N2212, N2342);
nand NAND4 (N2862, N2859, N1117, N1032, N304);
xor XOR2 (N2863, N2862, N1592);
buf BUF1 (N2864, N2856);
not NOT1 (N2865, N2838);
or OR4 (N2866, N2860, N1218, N1976, N2577);
and AND2 (N2867, N2866, N575);
xor XOR2 (N2868, N2863, N767);
or OR4 (N2869, N2865, N2405, N40, N1947);
xor XOR2 (N2870, N2835, N1298);
not NOT1 (N2871, N2858);
nand NAND4 (N2872, N2868, N679, N2111, N665);
xor XOR2 (N2873, N2869, N1357);
or OR3 (N2874, N2851, N1926, N57);
buf BUF1 (N2875, N2872);
nand NAND4 (N2876, N2867, N2437, N458, N2788);
and AND2 (N2877, N2848, N1543);
buf BUF1 (N2878, N2857);
xor XOR2 (N2879, N2870, N1297);
not NOT1 (N2880, N2861);
not NOT1 (N2881, N2878);
not NOT1 (N2882, N2864);
nor NOR3 (N2883, N2871, N436, N2638);
nand NAND3 (N2884, N2879, N884, N1725);
xor XOR2 (N2885, N2875, N2714);
buf BUF1 (N2886, N2877);
nor NOR4 (N2887, N2876, N700, N488, N2753);
xor XOR2 (N2888, N2882, N2382);
not NOT1 (N2889, N2873);
and AND4 (N2890, N2887, N430, N2671, N2091);
buf BUF1 (N2891, N2889);
xor XOR2 (N2892, N2874, N2269);
nand NAND2 (N2893, N2880, N1378);
nor NOR4 (N2894, N2890, N1616, N2241, N2634);
not NOT1 (N2895, N2883);
and AND4 (N2896, N2893, N641, N647, N1652);
not NOT1 (N2897, N2888);
not NOT1 (N2898, N2892);
not NOT1 (N2899, N2895);
not NOT1 (N2900, N2891);
and AND3 (N2901, N2900, N567, N176);
and AND2 (N2902, N2885, N2609);
not NOT1 (N2903, N2884);
nand NAND4 (N2904, N2886, N1810, N1347, N1427);
xor XOR2 (N2905, N2894, N2546);
and AND2 (N2906, N2904, N8);
or OR3 (N2907, N2897, N1124, N2711);
nor NOR2 (N2908, N2901, N298);
xor XOR2 (N2909, N2906, N2773);
nor NOR4 (N2910, N2881, N1772, N2559, N2516);
and AND2 (N2911, N2905, N599);
or OR3 (N2912, N2899, N2910, N2911);
or OR3 (N2913, N1693, N2704, N410);
and AND2 (N2914, N2896, N2421);
or OR2 (N2915, N1109, N1263);
and AND2 (N2916, N2907, N2447);
not NOT1 (N2917, N2914);
and AND4 (N2918, N2909, N616, N301, N897);
nor NOR2 (N2919, N2917, N1487);
not NOT1 (N2920, N2918);
and AND3 (N2921, N2915, N2625, N183);
not NOT1 (N2922, N2908);
or OR2 (N2923, N2913, N224);
or OR2 (N2924, N2898, N342);
and AND3 (N2925, N2922, N2025, N2278);
nand NAND3 (N2926, N2921, N23, N472);
and AND2 (N2927, N2902, N2902);
xor XOR2 (N2928, N2903, N2009);
xor XOR2 (N2929, N2912, N1447);
and AND2 (N2930, N2927, N1708);
or OR4 (N2931, N2929, N1467, N2564, N1293);
nor NOR3 (N2932, N2924, N818, N786);
nand NAND2 (N2933, N2928, N266);
xor XOR2 (N2934, N2926, N563);
nor NOR4 (N2935, N2933, N1814, N803, N2785);
or OR2 (N2936, N2931, N1641);
or OR3 (N2937, N2919, N22, N172);
nand NAND2 (N2938, N2930, N2769);
buf BUF1 (N2939, N2935);
and AND3 (N2940, N2934, N2569, N2213);
buf BUF1 (N2941, N2916);
nand NAND2 (N2942, N2940, N2813);
nor NOR2 (N2943, N2939, N500);
nand NAND2 (N2944, N2942, N2776);
xor XOR2 (N2945, N2938, N1589);
buf BUF1 (N2946, N2923);
nand NAND2 (N2947, N2932, N2018);
nand NAND2 (N2948, N2936, N794);
buf BUF1 (N2949, N2937);
not NOT1 (N2950, N2947);
xor XOR2 (N2951, N2950, N1804);
and AND2 (N2952, N2920, N2488);
and AND3 (N2953, N2943, N1638, N820);
xor XOR2 (N2954, N2953, N2046);
not NOT1 (N2955, N2941);
or OR4 (N2956, N2949, N1869, N1883, N2225);
not NOT1 (N2957, N2948);
and AND2 (N2958, N2955, N1144);
nor NOR2 (N2959, N2946, N1017);
nand NAND3 (N2960, N2957, N1697, N2359);
and AND2 (N2961, N2954, N2711);
or OR2 (N2962, N2960, N742);
nand NAND3 (N2963, N2925, N992, N2257);
nor NOR2 (N2964, N2958, N1694);
xor XOR2 (N2965, N2959, N664);
nor NOR4 (N2966, N2951, N1406, N2447, N670);
xor XOR2 (N2967, N2945, N1235);
nor NOR4 (N2968, N2967, N2565, N1894, N2884);
nor NOR4 (N2969, N2964, N1321, N2904, N3);
nand NAND2 (N2970, N2956, N1156);
not NOT1 (N2971, N2966);
buf BUF1 (N2972, N2963);
or OR2 (N2973, N2944, N107);
buf BUF1 (N2974, N2969);
nor NOR2 (N2975, N2952, N2291);
xor XOR2 (N2976, N2971, N1905);
nand NAND3 (N2977, N2968, N1686, N1745);
or OR3 (N2978, N2976, N603, N59);
xor XOR2 (N2979, N2973, N2876);
nor NOR4 (N2980, N2961, N977, N571, N376);
nand NAND2 (N2981, N2979, N2163);
nor NOR2 (N2982, N2970, N874);
xor XOR2 (N2983, N2982, N2032);
or OR4 (N2984, N2962, N1988, N2271, N2198);
nor NOR3 (N2985, N2965, N2025, N1244);
nand NAND4 (N2986, N2981, N1557, N2313, N1647);
nor NOR4 (N2987, N2977, N2149, N2116, N2655);
and AND4 (N2988, N2987, N2319, N2892, N1143);
or OR2 (N2989, N2978, N951);
xor XOR2 (N2990, N2985, N1015);
or OR4 (N2991, N2972, N48, N89, N2952);
buf BUF1 (N2992, N2991);
buf BUF1 (N2993, N2992);
not NOT1 (N2994, N2975);
nor NOR4 (N2995, N2988, N2375, N1585, N1592);
xor XOR2 (N2996, N2986, N967);
nor NOR3 (N2997, N2994, N2054, N2224);
not NOT1 (N2998, N2995);
nand NAND3 (N2999, N2997, N2252, N1168);
or OR3 (N3000, N2999, N1044, N2834);
or OR2 (N3001, N2974, N2450);
and AND4 (N3002, N2996, N587, N2002, N1502);
nor NOR2 (N3003, N2998, N2074);
nand NAND4 (N3004, N2993, N1627, N2847, N760);
and AND2 (N3005, N2983, N2307);
not NOT1 (N3006, N3001);
and AND2 (N3007, N2989, N2944);
buf BUF1 (N3008, N3006);
xor XOR2 (N3009, N2980, N168);
and AND3 (N3010, N3005, N2339, N2805);
nor NOR4 (N3011, N2990, N1310, N1642, N1308);
buf BUF1 (N3012, N2984);
nor NOR2 (N3013, N3007, N2317);
buf BUF1 (N3014, N3011);
xor XOR2 (N3015, N3008, N1578);
or OR4 (N3016, N3004, N2239, N2182, N629);
xor XOR2 (N3017, N3013, N370);
nand NAND4 (N3018, N3000, N1291, N2723, N75);
not NOT1 (N3019, N3015);
and AND3 (N3020, N3014, N306, N188);
xor XOR2 (N3021, N3016, N2826);
nor NOR3 (N3022, N3003, N2265, N1037);
buf BUF1 (N3023, N3017);
or OR3 (N3024, N3002, N954, N39);
nor NOR3 (N3025, N3010, N1220, N53);
xor XOR2 (N3026, N3020, N67);
and AND3 (N3027, N3023, N251, N520);
or OR4 (N3028, N3012, N2450, N2021, N2841);
xor XOR2 (N3029, N3009, N207);
nand NAND4 (N3030, N3026, N2203, N941, N1287);
nand NAND4 (N3031, N3027, N2416, N2919, N2784);
buf BUF1 (N3032, N3021);
buf BUF1 (N3033, N3025);
buf BUF1 (N3034, N3019);
xor XOR2 (N3035, N3030, N707);
buf BUF1 (N3036, N3032);
xor XOR2 (N3037, N3034, N418);
nor NOR2 (N3038, N3035, N2413);
or OR2 (N3039, N3031, N51);
nor NOR2 (N3040, N3022, N411);
buf BUF1 (N3041, N3039);
not NOT1 (N3042, N3036);
nand NAND3 (N3043, N3033, N1215, N1838);
nor NOR2 (N3044, N3037, N2907);
xor XOR2 (N3045, N3041, N1748);
or OR2 (N3046, N3024, N467);
and AND3 (N3047, N3040, N2197, N2440);
or OR4 (N3048, N3047, N40, N1124, N1499);
buf BUF1 (N3049, N3029);
or OR4 (N3050, N3046, N492, N2760, N2098);
nor NOR4 (N3051, N3049, N919, N1545, N2707);
nand NAND4 (N3052, N3044, N2774, N1041, N2872);
or OR2 (N3053, N3038, N2631);
xor XOR2 (N3054, N3051, N956);
buf BUF1 (N3055, N3028);
nand NAND3 (N3056, N3045, N1982, N992);
not NOT1 (N3057, N3055);
buf BUF1 (N3058, N3054);
or OR3 (N3059, N3056, N518, N1411);
nand NAND3 (N3060, N3057, N274, N1880);
nor NOR2 (N3061, N3042, N487);
xor XOR2 (N3062, N3018, N2503);
xor XOR2 (N3063, N3053, N1052);
not NOT1 (N3064, N3058);
buf BUF1 (N3065, N3063);
nor NOR4 (N3066, N3043, N135, N100, N446);
and AND3 (N3067, N3059, N1474, N1613);
xor XOR2 (N3068, N3060, N1542);
nor NOR3 (N3069, N3068, N1546, N2341);
and AND4 (N3070, N3061, N700, N2906, N723);
xor XOR2 (N3071, N3067, N4);
and AND3 (N3072, N3066, N2381, N2026);
and AND3 (N3073, N3069, N2638, N1504);
and AND4 (N3074, N3064, N1091, N1572, N2870);
buf BUF1 (N3075, N3070);
and AND2 (N3076, N3074, N1494);
nand NAND2 (N3077, N3052, N634);
buf BUF1 (N3078, N3073);
or OR4 (N3079, N3065, N1812, N1411, N1044);
not NOT1 (N3080, N3072);
nor NOR4 (N3081, N3076, N364, N1579, N1679);
nor NOR2 (N3082, N3079, N504);
buf BUF1 (N3083, N3082);
not NOT1 (N3084, N3078);
buf BUF1 (N3085, N3062);
buf BUF1 (N3086, N3080);
nand NAND4 (N3087, N3084, N48, N1492, N2849);
and AND2 (N3088, N3085, N2413);
not NOT1 (N3089, N3081);
or OR4 (N3090, N3077, N2168, N707, N2396);
not NOT1 (N3091, N3087);
or OR4 (N3092, N3050, N853, N2486, N767);
and AND2 (N3093, N3086, N2999);
and AND2 (N3094, N3071, N417);
buf BUF1 (N3095, N3092);
xor XOR2 (N3096, N3095, N1146);
not NOT1 (N3097, N3094);
xor XOR2 (N3098, N3097, N1428);
and AND3 (N3099, N3090, N1408, N1133);
nor NOR3 (N3100, N3091, N1828, N2110);
nor NOR4 (N3101, N3098, N2239, N2715, N942);
nand NAND4 (N3102, N3093, N9, N686, N1542);
not NOT1 (N3103, N3075);
not NOT1 (N3104, N3096);
or OR4 (N3105, N3101, N270, N2457, N314);
xor XOR2 (N3106, N3099, N2650);
xor XOR2 (N3107, N3106, N2295);
nor NOR4 (N3108, N3103, N2917, N1138, N1799);
not NOT1 (N3109, N3102);
nor NOR4 (N3110, N3104, N233, N1181, N677);
nand NAND2 (N3111, N3110, N1717);
nor NOR2 (N3112, N3111, N410);
nand NAND4 (N3113, N3089, N187, N2156, N1957);
or OR3 (N3114, N3083, N1271, N289);
not NOT1 (N3115, N3100);
xor XOR2 (N3116, N3109, N2231);
or OR4 (N3117, N3088, N2092, N966, N2835);
buf BUF1 (N3118, N3115);
not NOT1 (N3119, N3105);
nor NOR2 (N3120, N3118, N379);
and AND3 (N3121, N3116, N223, N1800);
xor XOR2 (N3122, N3107, N203);
or OR2 (N3123, N3120, N959);
or OR3 (N3124, N3108, N19, N2379);
nand NAND3 (N3125, N3048, N1238, N2209);
or OR2 (N3126, N3113, N2480);
nand NAND2 (N3127, N3119, N1668);
or OR4 (N3128, N3124, N401, N861, N734);
xor XOR2 (N3129, N3122, N736);
nor NOR2 (N3130, N3117, N90);
nand NAND4 (N3131, N3121, N2622, N1345, N89);
xor XOR2 (N3132, N3112, N1168);
or OR2 (N3133, N3129, N26);
not NOT1 (N3134, N3127);
nand NAND2 (N3135, N3130, N837);
not NOT1 (N3136, N3132);
not NOT1 (N3137, N3136);
not NOT1 (N3138, N3134);
buf BUF1 (N3139, N3128);
not NOT1 (N3140, N3135);
and AND2 (N3141, N3131, N900);
nor NOR4 (N3142, N3126, N1597, N1192, N426);
nor NOR4 (N3143, N3133, N1842, N2347, N2833);
and AND3 (N3144, N3142, N733, N305);
and AND2 (N3145, N3140, N1381);
or OR2 (N3146, N3125, N2937);
buf BUF1 (N3147, N3143);
nor NOR3 (N3148, N3146, N2561, N2637);
and AND2 (N3149, N3147, N2671);
not NOT1 (N3150, N3145);
nor NOR4 (N3151, N3144, N755, N957, N518);
or OR4 (N3152, N3148, N1051, N2120, N283);
or OR3 (N3153, N3138, N706, N3007);
buf BUF1 (N3154, N3137);
nor NOR4 (N3155, N3149, N436, N2154, N623);
and AND4 (N3156, N3114, N2523, N970, N613);
not NOT1 (N3157, N3151);
nor NOR4 (N3158, N3154, N3066, N1215, N439);
or OR2 (N3159, N3152, N2566);
xor XOR2 (N3160, N3123, N2079);
buf BUF1 (N3161, N3150);
buf BUF1 (N3162, N3139);
xor XOR2 (N3163, N3162, N548);
or OR3 (N3164, N3161, N637, N1352);
or OR3 (N3165, N3153, N1780, N1754);
buf BUF1 (N3166, N3163);
buf BUF1 (N3167, N3156);
or OR4 (N3168, N3160, N1846, N317, N153);
or OR3 (N3169, N3167, N2050, N217);
or OR2 (N3170, N3141, N404);
not NOT1 (N3171, N3157);
not NOT1 (N3172, N3155);
and AND2 (N3173, N3166, N1963);
and AND2 (N3174, N3165, N316);
not NOT1 (N3175, N3168);
xor XOR2 (N3176, N3172, N1880);
buf BUF1 (N3177, N3170);
nand NAND4 (N3178, N3173, N1351, N998, N1992);
not NOT1 (N3179, N3178);
nor NOR3 (N3180, N3158, N1860, N2260);
nor NOR2 (N3181, N3169, N728);
or OR2 (N3182, N3181, N2307);
not NOT1 (N3183, N3164);
nand NAND4 (N3184, N3171, N2336, N507, N2467);
xor XOR2 (N3185, N3179, N3018);
nand NAND3 (N3186, N3176, N2691, N2957);
nor NOR2 (N3187, N3185, N1128);
nor NOR2 (N3188, N3183, N2147);
and AND2 (N3189, N3188, N935);
nor NOR2 (N3190, N3159, N2845);
nor NOR4 (N3191, N3180, N3102, N713, N318);
nand NAND4 (N3192, N3184, N874, N966, N1079);
and AND2 (N3193, N3174, N691);
nand NAND4 (N3194, N3191, N2174, N757, N1786);
buf BUF1 (N3195, N3194);
nand NAND3 (N3196, N3187, N208, N1743);
nand NAND4 (N3197, N3177, N1340, N3053, N30);
nand NAND2 (N3198, N3190, N3038);
nand NAND2 (N3199, N3186, N2709);
nor NOR3 (N3200, N3192, N1132, N1529);
xor XOR2 (N3201, N3196, N2207);
buf BUF1 (N3202, N3199);
and AND2 (N3203, N3197, N1166);
nand NAND3 (N3204, N3195, N47, N1006);
or OR2 (N3205, N3193, N97);
xor XOR2 (N3206, N3182, N2016);
buf BUF1 (N3207, N3202);
not NOT1 (N3208, N3203);
nand NAND3 (N3209, N3207, N1195, N151);
or OR4 (N3210, N3201, N898, N2845, N1803);
xor XOR2 (N3211, N3200, N783);
not NOT1 (N3212, N3211);
buf BUF1 (N3213, N3210);
buf BUF1 (N3214, N3209);
and AND3 (N3215, N3212, N1653, N2282);
xor XOR2 (N3216, N3175, N1189);
or OR4 (N3217, N3215, N2322, N59, N1119);
or OR2 (N3218, N3208, N305);
and AND4 (N3219, N3204, N2914, N1427, N651);
xor XOR2 (N3220, N3219, N1392);
buf BUF1 (N3221, N3213);
nor NOR2 (N3222, N3206, N421);
nor NOR3 (N3223, N3214, N2025, N254);
buf BUF1 (N3224, N3223);
or OR2 (N3225, N3189, N2132);
not NOT1 (N3226, N3221);
buf BUF1 (N3227, N3224);
nand NAND3 (N3228, N3217, N1597, N1328);
or OR2 (N3229, N3216, N3192);
buf BUF1 (N3230, N3225);
nand NAND2 (N3231, N3220, N1097);
not NOT1 (N3232, N3227);
buf BUF1 (N3233, N3228);
and AND2 (N3234, N3222, N2787);
not NOT1 (N3235, N3232);
xor XOR2 (N3236, N3205, N63);
or OR2 (N3237, N3218, N2989);
and AND3 (N3238, N3231, N1287, N2321);
nor NOR3 (N3239, N3234, N2333, N2552);
nor NOR2 (N3240, N3233, N792);
buf BUF1 (N3241, N3235);
buf BUF1 (N3242, N3198);
buf BUF1 (N3243, N3239);
buf BUF1 (N3244, N3243);
xor XOR2 (N3245, N3229, N61);
nand NAND4 (N3246, N3236, N571, N630, N3093);
and AND2 (N3247, N3245, N179);
xor XOR2 (N3248, N3244, N2861);
buf BUF1 (N3249, N3230);
buf BUF1 (N3250, N3246);
not NOT1 (N3251, N3237);
buf BUF1 (N3252, N3250);
xor XOR2 (N3253, N3251, N1453);
not NOT1 (N3254, N3226);
nor NOR2 (N3255, N3252, N3185);
or OR3 (N3256, N3238, N394, N1879);
nor NOR4 (N3257, N3255, N3146, N1964, N3138);
xor XOR2 (N3258, N3256, N631);
or OR2 (N3259, N3254, N2127);
nand NAND3 (N3260, N3253, N2763, N1328);
nor NOR3 (N3261, N3258, N2142, N2578);
nand NAND2 (N3262, N3242, N1318);
and AND3 (N3263, N3247, N2923, N1554);
buf BUF1 (N3264, N3259);
nand NAND2 (N3265, N3257, N400);
nor NOR3 (N3266, N3262, N2575, N1697);
or OR4 (N3267, N3266, N2896, N224, N2685);
buf BUF1 (N3268, N3240);
not NOT1 (N3269, N3268);
nand NAND3 (N3270, N3261, N640, N2877);
not NOT1 (N3271, N3270);
and AND2 (N3272, N3241, N2912);
nor NOR3 (N3273, N3260, N2289, N1856);
nand NAND4 (N3274, N3273, N715, N2940, N2043);
buf BUF1 (N3275, N3269);
xor XOR2 (N3276, N3267, N2947);
nand NAND2 (N3277, N3274, N100);
nor NOR2 (N3278, N3276, N1595);
nand NAND4 (N3279, N3272, N50, N1283, N492);
xor XOR2 (N3280, N3263, N3196);
nand NAND3 (N3281, N3248, N1956, N3098);
buf BUF1 (N3282, N3277);
nor NOR4 (N3283, N3271, N1668, N1154, N2537);
or OR3 (N3284, N3280, N3279, N1921);
or OR2 (N3285, N981, N2602);
or OR3 (N3286, N3265, N2075, N249);
nor NOR3 (N3287, N3285, N340, N2740);
not NOT1 (N3288, N3283);
nor NOR3 (N3289, N3249, N557, N2298);
or OR3 (N3290, N3281, N913, N2370);
nor NOR4 (N3291, N3289, N532, N2382, N892);
or OR2 (N3292, N3275, N2039);
nand NAND3 (N3293, N3287, N1018, N270);
xor XOR2 (N3294, N3291, N832);
nand NAND4 (N3295, N3290, N2073, N1324, N1634);
and AND4 (N3296, N3292, N810, N1683, N1494);
not NOT1 (N3297, N3296);
buf BUF1 (N3298, N3286);
not NOT1 (N3299, N3282);
and AND2 (N3300, N3264, N2300);
buf BUF1 (N3301, N3299);
not NOT1 (N3302, N3288);
xor XOR2 (N3303, N3301, N2984);
buf BUF1 (N3304, N3293);
nor NOR4 (N3305, N3278, N1625, N2134, N539);
and AND3 (N3306, N3294, N3166, N1426);
nor NOR2 (N3307, N3295, N3260);
or OR4 (N3308, N3300, N1791, N640, N172);
or OR4 (N3309, N3302, N383, N797, N2231);
not NOT1 (N3310, N3298);
nor NOR3 (N3311, N3306, N3182, N2387);
nor NOR4 (N3312, N3303, N672, N1387, N273);
buf BUF1 (N3313, N3305);
and AND3 (N3314, N3297, N2545, N2590);
nor NOR2 (N3315, N3308, N848);
buf BUF1 (N3316, N3315);
nor NOR4 (N3317, N3311, N2370, N1426, N2174);
not NOT1 (N3318, N3317);
buf BUF1 (N3319, N3313);
or OR2 (N3320, N3307, N1467);
not NOT1 (N3321, N3319);
nor NOR2 (N3322, N3314, N204);
and AND3 (N3323, N3321, N1642, N1015);
xor XOR2 (N3324, N3323, N2814);
buf BUF1 (N3325, N3316);
nor NOR4 (N3326, N3320, N2656, N779, N3129);
nand NAND3 (N3327, N3325, N2104, N443);
buf BUF1 (N3328, N3312);
xor XOR2 (N3329, N3318, N813);
not NOT1 (N3330, N3324);
nand NAND4 (N3331, N3310, N2424, N194, N866);
buf BUF1 (N3332, N3309);
not NOT1 (N3333, N3326);
and AND4 (N3334, N3329, N2626, N2489, N1526);
or OR2 (N3335, N3284, N1599);
or OR4 (N3336, N3328, N3032, N772, N836);
xor XOR2 (N3337, N3336, N2482);
buf BUF1 (N3338, N3331);
or OR3 (N3339, N3330, N2485, N61);
nor NOR3 (N3340, N3322, N1206, N916);
not NOT1 (N3341, N3327);
not NOT1 (N3342, N3333);
or OR4 (N3343, N3339, N942, N1811, N1271);
nor NOR3 (N3344, N3332, N1333, N314);
nor NOR3 (N3345, N3342, N1649, N1823);
and AND3 (N3346, N3338, N2569, N528);
or OR3 (N3347, N3344, N2382, N617);
xor XOR2 (N3348, N3340, N1900);
xor XOR2 (N3349, N3341, N2171);
buf BUF1 (N3350, N3337);
or OR3 (N3351, N3345, N1671, N1217);
nand NAND3 (N3352, N3343, N1892, N1857);
nor NOR2 (N3353, N3350, N2814);
xor XOR2 (N3354, N3335, N1130);
buf BUF1 (N3355, N3353);
not NOT1 (N3356, N3355);
nor NOR4 (N3357, N3351, N1953, N1669, N2610);
nand NAND4 (N3358, N3352, N3235, N704, N747);
buf BUF1 (N3359, N3346);
nor NOR3 (N3360, N3354, N708, N2099);
nor NOR3 (N3361, N3348, N846, N2222);
nand NAND2 (N3362, N3356, N1899);
and AND2 (N3363, N3304, N183);
or OR3 (N3364, N3358, N2786, N1995);
xor XOR2 (N3365, N3349, N210);
buf BUF1 (N3366, N3360);
nor NOR4 (N3367, N3365, N1480, N3122, N3232);
nor NOR4 (N3368, N3366, N2947, N474, N3244);
buf BUF1 (N3369, N3347);
xor XOR2 (N3370, N3362, N594);
not NOT1 (N3371, N3368);
buf BUF1 (N3372, N3363);
xor XOR2 (N3373, N3367, N95);
buf BUF1 (N3374, N3334);
nand NAND4 (N3375, N3371, N1934, N1620, N3101);
and AND4 (N3376, N3374, N1715, N2169, N983);
and AND4 (N3377, N3361, N2539, N2143, N2145);
buf BUF1 (N3378, N3370);
nand NAND2 (N3379, N3378, N3045);
xor XOR2 (N3380, N3359, N2167);
nand NAND3 (N3381, N3377, N1499, N3127);
or OR4 (N3382, N3381, N1958, N1413, N533);
nor NOR2 (N3383, N3369, N1279);
not NOT1 (N3384, N3376);
or OR3 (N3385, N3383, N950, N660);
nor NOR2 (N3386, N3380, N1976);
nor NOR3 (N3387, N3385, N2314, N1243);
buf BUF1 (N3388, N3375);
and AND4 (N3389, N3388, N859, N2770, N3359);
nand NAND4 (N3390, N3384, N3379, N539, N889);
not NOT1 (N3391, N498);
xor XOR2 (N3392, N3372, N1103);
nand NAND2 (N3393, N3389, N1789);
nor NOR2 (N3394, N3382, N3011);
buf BUF1 (N3395, N3386);
not NOT1 (N3396, N3392);
buf BUF1 (N3397, N3396);
xor XOR2 (N3398, N3357, N2462);
not NOT1 (N3399, N3387);
buf BUF1 (N3400, N3373);
buf BUF1 (N3401, N3400);
nand NAND4 (N3402, N3391, N186, N3111, N501);
nor NOR3 (N3403, N3395, N2029, N1790);
and AND4 (N3404, N3399, N2171, N3278, N18);
not NOT1 (N3405, N3402);
nor NOR2 (N3406, N3394, N2417);
xor XOR2 (N3407, N3397, N2483);
or OR3 (N3408, N3403, N2537, N706);
and AND2 (N3409, N3406, N2791);
or OR2 (N3410, N3364, N2558);
buf BUF1 (N3411, N3408);
nor NOR3 (N3412, N3404, N479, N1911);
and AND3 (N3413, N3405, N1421, N1873);
or OR2 (N3414, N3398, N1624);
or OR4 (N3415, N3393, N1044, N1255, N2662);
xor XOR2 (N3416, N3412, N564);
or OR2 (N3417, N3416, N3065);
or OR3 (N3418, N3401, N40, N2339);
nor NOR4 (N3419, N3410, N2014, N2076, N1072);
or OR2 (N3420, N3415, N525);
buf BUF1 (N3421, N3418);
and AND3 (N3422, N3409, N724, N514);
nand NAND2 (N3423, N3417, N1508);
buf BUF1 (N3424, N3413);
xor XOR2 (N3425, N3422, N1419);
not NOT1 (N3426, N3421);
and AND3 (N3427, N3420, N129, N2262);
nor NOR3 (N3428, N3424, N3156, N1882);
nor NOR4 (N3429, N3411, N343, N1403, N1295);
nor NOR4 (N3430, N3426, N102, N1872, N2679);
xor XOR2 (N3431, N3414, N2160);
xor XOR2 (N3432, N3419, N3387);
and AND3 (N3433, N3427, N1540, N2965);
nor NOR3 (N3434, N3425, N1818, N298);
not NOT1 (N3435, N3429);
nor NOR4 (N3436, N3423, N3093, N3163, N148);
buf BUF1 (N3437, N3435);
buf BUF1 (N3438, N3431);
or OR2 (N3439, N3436, N1220);
not NOT1 (N3440, N3439);
or OR4 (N3441, N3438, N1981, N1304, N1355);
nand NAND3 (N3442, N3407, N2321, N1147);
and AND2 (N3443, N3432, N3221);
nor NOR4 (N3444, N3442, N328, N1368, N121);
nor NOR4 (N3445, N3428, N2846, N220, N159);
or OR3 (N3446, N3430, N2512, N316);
and AND2 (N3447, N3434, N3274);
nor NOR2 (N3448, N3447, N260);
buf BUF1 (N3449, N3390);
nand NAND3 (N3450, N3445, N203, N1146);
or OR2 (N3451, N3443, N348);
and AND3 (N3452, N3448, N2930, N3122);
or OR3 (N3453, N3433, N3343, N966);
nor NOR3 (N3454, N3446, N199, N2331);
buf BUF1 (N3455, N3453);
not NOT1 (N3456, N3444);
or OR3 (N3457, N3437, N97, N3433);
xor XOR2 (N3458, N3449, N836);
nand NAND3 (N3459, N3450, N953, N2847);
nand NAND2 (N3460, N3457, N2982);
nand NAND4 (N3461, N3456, N2981, N664, N2187);
nand NAND4 (N3462, N3441, N1337, N815, N1137);
nor NOR2 (N3463, N3452, N420);
not NOT1 (N3464, N3454);
or OR2 (N3465, N3461, N3203);
nand NAND4 (N3466, N3440, N197, N3144, N2648);
nand NAND3 (N3467, N3460, N1242, N3284);
not NOT1 (N3468, N3465);
or OR2 (N3469, N3464, N2865);
nor NOR3 (N3470, N3468, N3447, N315);
or OR3 (N3471, N3459, N417, N3294);
and AND3 (N3472, N3458, N130, N256);
nand NAND4 (N3473, N3463, N432, N849, N3109);
not NOT1 (N3474, N3467);
and AND2 (N3475, N3471, N982);
and AND3 (N3476, N3466, N338, N2985);
xor XOR2 (N3477, N3473, N1519);
or OR4 (N3478, N3455, N1067, N280, N883);
not NOT1 (N3479, N3462);
not NOT1 (N3480, N3475);
buf BUF1 (N3481, N3474);
and AND2 (N3482, N3477, N1382);
or OR2 (N3483, N3479, N1957);
xor XOR2 (N3484, N3483, N1161);
buf BUF1 (N3485, N3478);
xor XOR2 (N3486, N3476, N138);
nor NOR2 (N3487, N3481, N907);
buf BUF1 (N3488, N3470);
and AND4 (N3489, N3480, N2846, N3147, N558);
nand NAND2 (N3490, N3482, N862);
not NOT1 (N3491, N3489);
and AND3 (N3492, N3469, N1146, N2072);
and AND2 (N3493, N3490, N1774);
nor NOR2 (N3494, N3493, N465);
or OR3 (N3495, N3488, N183, N1535);
xor XOR2 (N3496, N3491, N625);
and AND4 (N3497, N3451, N708, N1018, N222);
not NOT1 (N3498, N3494);
nor NOR4 (N3499, N3496, N958, N518, N1933);
not NOT1 (N3500, N3497);
or OR4 (N3501, N3499, N2915, N1375, N1683);
xor XOR2 (N3502, N3472, N3209);
xor XOR2 (N3503, N3486, N2291);
nand NAND4 (N3504, N3485, N3432, N2147, N2368);
nand NAND4 (N3505, N3503, N445, N1578, N3310);
xor XOR2 (N3506, N3504, N3302);
and AND4 (N3507, N3498, N2255, N2230, N556);
xor XOR2 (N3508, N3492, N136);
not NOT1 (N3509, N3487);
or OR2 (N3510, N3500, N2940);
and AND2 (N3511, N3505, N1216);
or OR3 (N3512, N3495, N3123, N1222);
and AND3 (N3513, N3507, N3226, N797);
and AND2 (N3514, N3508, N2752);
nor NOR3 (N3515, N3506, N3382, N2770);
or OR2 (N3516, N3515, N1642);
nor NOR2 (N3517, N3502, N1003);
buf BUF1 (N3518, N3510);
or OR4 (N3519, N3518, N2364, N2760, N2824);
not NOT1 (N3520, N3509);
xor XOR2 (N3521, N3514, N3003);
nor NOR3 (N3522, N3519, N1825, N2836);
and AND4 (N3523, N3516, N3162, N538, N910);
xor XOR2 (N3524, N3522, N1319);
or OR2 (N3525, N3501, N2241);
buf BUF1 (N3526, N3511);
and AND3 (N3527, N3513, N585, N2830);
or OR2 (N3528, N3517, N2571);
nor NOR2 (N3529, N3520, N2118);
buf BUF1 (N3530, N3512);
or OR4 (N3531, N3529, N1369, N3132, N2854);
nor NOR4 (N3532, N3484, N955, N1077, N140);
or OR2 (N3533, N3523, N2300);
and AND4 (N3534, N3525, N2918, N2901, N754);
or OR3 (N3535, N3526, N3411, N2937);
or OR4 (N3536, N3524, N3468, N1335, N910);
nor NOR4 (N3537, N3533, N2850, N3386, N1545);
nand NAND2 (N3538, N3527, N3493);
nor NOR4 (N3539, N3537, N1309, N2235, N3202);
nand NAND2 (N3540, N3539, N2610);
and AND3 (N3541, N3536, N1518, N921);
nor NOR2 (N3542, N3531, N3480);
or OR3 (N3543, N3538, N2637, N3111);
buf BUF1 (N3544, N3534);
nand NAND2 (N3545, N3541, N530);
not NOT1 (N3546, N3544);
nor NOR4 (N3547, N3540, N481, N3034, N1208);
not NOT1 (N3548, N3547);
nor NOR3 (N3549, N3542, N848, N948);
not NOT1 (N3550, N3549);
and AND4 (N3551, N3532, N986, N2704, N126);
nor NOR4 (N3552, N3551, N673, N226, N1311);
or OR2 (N3553, N3545, N2716);
nor NOR3 (N3554, N3546, N1509, N2984);
and AND4 (N3555, N3550, N2978, N3314, N2912);
xor XOR2 (N3556, N3535, N3249);
xor XOR2 (N3557, N3554, N1428);
or OR4 (N3558, N3528, N1527, N1267, N2108);
nor NOR2 (N3559, N3548, N1694);
not NOT1 (N3560, N3553);
nand NAND3 (N3561, N3556, N315, N2474);
nand NAND3 (N3562, N3558, N1466, N428);
xor XOR2 (N3563, N3562, N1168);
buf BUF1 (N3564, N3555);
buf BUF1 (N3565, N3560);
not NOT1 (N3566, N3521);
or OR2 (N3567, N3561, N3501);
not NOT1 (N3568, N3567);
nor NOR4 (N3569, N3559, N552, N3511, N2951);
nand NAND2 (N3570, N3530, N1790);
and AND4 (N3571, N3569, N786, N3363, N2724);
or OR2 (N3572, N3543, N2258);
nand NAND3 (N3573, N3552, N2225, N2310);
nand NAND2 (N3574, N3564, N1629);
not NOT1 (N3575, N3571);
not NOT1 (N3576, N3574);
xor XOR2 (N3577, N3576, N889);
nand NAND4 (N3578, N3568, N795, N1403, N3036);
or OR3 (N3579, N3577, N3515, N1164);
not NOT1 (N3580, N3557);
buf BUF1 (N3581, N3570);
nand NAND2 (N3582, N3563, N1317);
nand NAND2 (N3583, N3582, N271);
not NOT1 (N3584, N3578);
and AND4 (N3585, N3575, N2937, N2864, N2477);
nand NAND4 (N3586, N3584, N1845, N3413, N1444);
and AND3 (N3587, N3586, N614, N498);
xor XOR2 (N3588, N3579, N447);
xor XOR2 (N3589, N3588, N2908);
xor XOR2 (N3590, N3587, N3372);
buf BUF1 (N3591, N3566);
not NOT1 (N3592, N3591);
xor XOR2 (N3593, N3583, N202);
not NOT1 (N3594, N3589);
and AND3 (N3595, N3581, N3563, N3476);
nor NOR4 (N3596, N3592, N2264, N1619, N2374);
buf BUF1 (N3597, N3572);
or OR4 (N3598, N3597, N3187, N2604, N3429);
not NOT1 (N3599, N3565);
and AND2 (N3600, N3590, N221);
xor XOR2 (N3601, N3595, N3206);
buf BUF1 (N3602, N3601);
and AND3 (N3603, N3593, N386, N1619);
xor XOR2 (N3604, N3573, N1043);
or OR3 (N3605, N3585, N3411, N2906);
not NOT1 (N3606, N3603);
nand NAND3 (N3607, N3599, N1609, N1574);
buf BUF1 (N3608, N3604);
xor XOR2 (N3609, N3606, N3551);
or OR2 (N3610, N3607, N2418);
xor XOR2 (N3611, N3610, N371);
buf BUF1 (N3612, N3598);
nand NAND4 (N3613, N3594, N287, N2006, N641);
or OR3 (N3614, N3613, N1800, N2186);
not NOT1 (N3615, N3580);
not NOT1 (N3616, N3609);
xor XOR2 (N3617, N3602, N3146);
nand NAND3 (N3618, N3608, N27, N3579);
and AND4 (N3619, N3615, N2598, N1509, N2380);
xor XOR2 (N3620, N3618, N3604);
xor XOR2 (N3621, N3611, N470);
xor XOR2 (N3622, N3617, N630);
nand NAND4 (N3623, N3616, N358, N84, N2716);
nand NAND3 (N3624, N3605, N2561, N2467);
or OR3 (N3625, N3620, N3291, N2981);
nand NAND3 (N3626, N3619, N321, N890);
xor XOR2 (N3627, N3612, N331);
xor XOR2 (N3628, N3614, N42);
nor NOR4 (N3629, N3600, N1583, N2025, N2460);
nand NAND2 (N3630, N3622, N549);
buf BUF1 (N3631, N3630);
xor XOR2 (N3632, N3629, N203);
or OR3 (N3633, N3596, N2102, N3596);
nand NAND4 (N3634, N3626, N2421, N489, N1992);
buf BUF1 (N3635, N3633);
not NOT1 (N3636, N3627);
nand NAND3 (N3637, N3635, N111, N230);
nor NOR4 (N3638, N3624, N1585, N445, N3524);
nor NOR4 (N3639, N3631, N1482, N565, N3607);
and AND3 (N3640, N3639, N2583, N2402);
nor NOR4 (N3641, N3636, N1922, N3275, N2828);
or OR3 (N3642, N3638, N1490, N3017);
or OR4 (N3643, N3628, N1427, N583, N3511);
nor NOR3 (N3644, N3637, N2331, N929);
buf BUF1 (N3645, N3643);
nor NOR4 (N3646, N3623, N1513, N2503, N1166);
buf BUF1 (N3647, N3632);
buf BUF1 (N3648, N3647);
nand NAND3 (N3649, N3648, N2439, N3027);
xor XOR2 (N3650, N3644, N1856);
or OR4 (N3651, N3650, N1605, N2329, N982);
xor XOR2 (N3652, N3642, N536);
nor NOR3 (N3653, N3645, N3560, N2500);
nor NOR2 (N3654, N3646, N2781);
or OR3 (N3655, N3634, N1501, N663);
nor NOR3 (N3656, N3641, N1010, N1801);
nor NOR3 (N3657, N3655, N970, N2364);
nor NOR2 (N3658, N3649, N3570);
nor NOR2 (N3659, N3658, N987);
or OR4 (N3660, N3621, N1904, N2823, N168);
nand NAND4 (N3661, N3653, N410, N808, N1462);
not NOT1 (N3662, N3659);
buf BUF1 (N3663, N3656);
nor NOR4 (N3664, N3661, N592, N3253, N3119);
xor XOR2 (N3665, N3652, N1483);
and AND3 (N3666, N3640, N701, N1825);
xor XOR2 (N3667, N3654, N1712);
nor NOR2 (N3668, N3667, N1517);
or OR3 (N3669, N3664, N539, N1546);
nor NOR3 (N3670, N3625, N1393, N791);
and AND4 (N3671, N3665, N1636, N3128, N284);
not NOT1 (N3672, N3662);
nor NOR4 (N3673, N3651, N3394, N1069, N3115);
xor XOR2 (N3674, N3663, N2680);
nor NOR2 (N3675, N3672, N279);
or OR2 (N3676, N3674, N3175);
nand NAND3 (N3677, N3668, N2613, N3573);
or OR2 (N3678, N3673, N1961);
buf BUF1 (N3679, N3671);
not NOT1 (N3680, N3679);
buf BUF1 (N3681, N3669);
buf BUF1 (N3682, N3678);
and AND4 (N3683, N3676, N2922, N2557, N2247);
not NOT1 (N3684, N3682);
nor NOR2 (N3685, N3666, N3449);
not NOT1 (N3686, N3684);
buf BUF1 (N3687, N3670);
nand NAND4 (N3688, N3687, N2798, N3346, N1850);
nor NOR2 (N3689, N3675, N3435);
nor NOR4 (N3690, N3677, N1603, N61, N2589);
not NOT1 (N3691, N3683);
buf BUF1 (N3692, N3660);
nand NAND4 (N3693, N3689, N920, N776, N2722);
buf BUF1 (N3694, N3691);
nand NAND3 (N3695, N3690, N3516, N2719);
or OR3 (N3696, N3688, N3451, N2929);
nor NOR2 (N3697, N3696, N2948);
buf BUF1 (N3698, N3692);
nor NOR3 (N3699, N3680, N2449, N3673);
or OR4 (N3700, N3697, N2436, N2695, N2003);
nor NOR4 (N3701, N3695, N409, N1074, N1831);
and AND2 (N3702, N3693, N282);
nor NOR4 (N3703, N3657, N1912, N1296, N843);
nand NAND2 (N3704, N3685, N1525);
and AND2 (N3705, N3701, N3125);
xor XOR2 (N3706, N3703, N187);
nor NOR3 (N3707, N3699, N849, N2217);
and AND4 (N3708, N3706, N1195, N2241, N679);
nand NAND3 (N3709, N3700, N333, N2374);
xor XOR2 (N3710, N3681, N3631);
or OR4 (N3711, N3709, N332, N3242, N1736);
xor XOR2 (N3712, N3694, N1840);
nor NOR4 (N3713, N3705, N755, N2008, N1868);
not NOT1 (N3714, N3712);
nor NOR3 (N3715, N3702, N1607, N1964);
nor NOR4 (N3716, N3711, N2786, N1852, N1240);
and AND2 (N3717, N3698, N739);
nor NOR3 (N3718, N3714, N1997, N1697);
nand NAND4 (N3719, N3717, N3060, N3034, N600);
or OR4 (N3720, N3704, N2149, N3518, N2430);
nor NOR3 (N3721, N3713, N2510, N29);
xor XOR2 (N3722, N3686, N481);
buf BUF1 (N3723, N3716);
xor XOR2 (N3724, N3719, N3006);
and AND4 (N3725, N3715, N3616, N3003, N2622);
not NOT1 (N3726, N3721);
nor NOR2 (N3727, N3724, N983);
buf BUF1 (N3728, N3718);
nor NOR3 (N3729, N3728, N3267, N2129);
nor NOR2 (N3730, N3710, N1937);
buf BUF1 (N3731, N3726);
nor NOR4 (N3732, N3729, N2492, N2545, N3495);
nand NAND3 (N3733, N3722, N219, N2265);
or OR3 (N3734, N3733, N2124, N63);
and AND2 (N3735, N3731, N1372);
xor XOR2 (N3736, N3720, N518);
or OR3 (N3737, N3734, N3260, N228);
nand NAND3 (N3738, N3723, N1389, N456);
or OR3 (N3739, N3730, N50, N1209);
buf BUF1 (N3740, N3737);
nor NOR2 (N3741, N3736, N2918);
xor XOR2 (N3742, N3740, N2904);
xor XOR2 (N3743, N3742, N1058);
nand NAND4 (N3744, N3708, N2223, N640, N3740);
or OR4 (N3745, N3725, N3085, N135, N2131);
buf BUF1 (N3746, N3739);
xor XOR2 (N3747, N3743, N1414);
xor XOR2 (N3748, N3727, N2570);
xor XOR2 (N3749, N3735, N1506);
or OR4 (N3750, N3707, N3638, N880, N341);
buf BUF1 (N3751, N3749);
or OR4 (N3752, N3732, N1733, N3561, N3103);
or OR4 (N3753, N3750, N2501, N571, N3444);
nor NOR3 (N3754, N3745, N696, N3673);
nor NOR4 (N3755, N3754, N1029, N2868, N2625);
xor XOR2 (N3756, N3755, N1270);
nor NOR3 (N3757, N3752, N738, N1135);
or OR4 (N3758, N3746, N3353, N3626, N2031);
nor NOR4 (N3759, N3756, N3592, N1778, N164);
or OR3 (N3760, N3751, N1802, N3344);
nor NOR3 (N3761, N3738, N1063, N3402);
nor NOR3 (N3762, N3747, N1683, N3632);
xor XOR2 (N3763, N3757, N3410);
and AND4 (N3764, N3744, N1461, N1030, N2836);
xor XOR2 (N3765, N3764, N2393);
nand NAND3 (N3766, N3763, N512, N432);
buf BUF1 (N3767, N3762);
nand NAND3 (N3768, N3760, N1745, N1690);
or OR3 (N3769, N3765, N413, N844);
xor XOR2 (N3770, N3766, N2347);
or OR3 (N3771, N3767, N106, N908);
not NOT1 (N3772, N3758);
nor NOR2 (N3773, N3771, N282);
and AND2 (N3774, N3753, N427);
or OR3 (N3775, N3774, N2585, N2030);
buf BUF1 (N3776, N3759);
not NOT1 (N3777, N3768);
nor NOR4 (N3778, N3772, N3454, N1397, N3164);
nand NAND2 (N3779, N3777, N1302);
or OR3 (N3780, N3769, N3394, N2786);
not NOT1 (N3781, N3779);
buf BUF1 (N3782, N3741);
nand NAND3 (N3783, N3780, N1448, N1881);
not NOT1 (N3784, N3761);
nor NOR4 (N3785, N3748, N3743, N836, N418);
and AND3 (N3786, N3773, N188, N3099);
nand NAND3 (N3787, N3786, N1880, N1579);
not NOT1 (N3788, N3783);
nor NOR4 (N3789, N3785, N620, N3555, N755);
nand NAND2 (N3790, N3789, N504);
not NOT1 (N3791, N3782);
xor XOR2 (N3792, N3787, N137);
xor XOR2 (N3793, N3791, N493);
and AND4 (N3794, N3775, N2136, N3668, N2588);
nor NOR3 (N3795, N3776, N3284, N1430);
buf BUF1 (N3796, N3770);
buf BUF1 (N3797, N3795);
and AND4 (N3798, N3797, N3740, N2146, N3669);
nor NOR3 (N3799, N3793, N1848, N159);
xor XOR2 (N3800, N3798, N3690);
nor NOR3 (N3801, N3799, N3260, N488);
not NOT1 (N3802, N3794);
or OR4 (N3803, N3802, N1690, N2926, N2047);
not NOT1 (N3804, N3792);
and AND3 (N3805, N3801, N3587, N3060);
not NOT1 (N3806, N3788);
not NOT1 (N3807, N3806);
nor NOR4 (N3808, N3790, N1471, N386, N2070);
or OR3 (N3809, N3807, N2640, N771);
buf BUF1 (N3810, N3805);
nand NAND3 (N3811, N3781, N767, N3271);
and AND3 (N3812, N3784, N980, N998);
nor NOR2 (N3813, N3778, N854);
nand NAND3 (N3814, N3809, N1718, N1955);
or OR3 (N3815, N3800, N3228, N1963);
or OR4 (N3816, N3813, N643, N1418, N3437);
and AND4 (N3817, N3803, N2559, N3222, N1662);
and AND3 (N3818, N3814, N8, N923);
buf BUF1 (N3819, N3812);
not NOT1 (N3820, N3808);
buf BUF1 (N3821, N3817);
nand NAND4 (N3822, N3821, N2987, N3303, N847);
nor NOR3 (N3823, N3804, N220, N1527);
nand NAND3 (N3824, N3820, N910, N894);
nand NAND2 (N3825, N3818, N3514);
nor NOR3 (N3826, N3796, N3301, N1736);
and AND3 (N3827, N3810, N2384, N1220);
nor NOR2 (N3828, N3816, N13);
nand NAND3 (N3829, N3815, N3211, N820);
xor XOR2 (N3830, N3811, N383);
and AND2 (N3831, N3822, N934);
buf BUF1 (N3832, N3828);
or OR2 (N3833, N3829, N2346);
xor XOR2 (N3834, N3819, N705);
nand NAND2 (N3835, N3833, N1268);
and AND2 (N3836, N3830, N2725);
nor NOR3 (N3837, N3823, N530, N2508);
nor NOR3 (N3838, N3832, N277, N502);
nand NAND3 (N3839, N3836, N3304, N1291);
xor XOR2 (N3840, N3834, N238);
not NOT1 (N3841, N3826);
or OR4 (N3842, N3841, N3359, N209, N3344);
or OR2 (N3843, N3835, N1552);
nor NOR3 (N3844, N3840, N3202, N2042);
and AND4 (N3845, N3844, N734, N192, N2162);
and AND3 (N3846, N3839, N2502, N2163);
nand NAND4 (N3847, N3831, N1599, N2330, N2753);
or OR3 (N3848, N3838, N2007, N2815);
or OR2 (N3849, N3843, N3115);
nand NAND4 (N3850, N3837, N430, N2229, N839);
buf BUF1 (N3851, N3845);
buf BUF1 (N3852, N3848);
nand NAND3 (N3853, N3846, N497, N887);
and AND2 (N3854, N3847, N3259);
nand NAND2 (N3855, N3853, N3761);
nor NOR4 (N3856, N3855, N115, N3737, N3346);
and AND2 (N3857, N3825, N2579);
buf BUF1 (N3858, N3849);
not NOT1 (N3859, N3858);
or OR2 (N3860, N3842, N2648);
not NOT1 (N3861, N3857);
xor XOR2 (N3862, N3860, N410);
or OR4 (N3863, N3862, N628, N3070, N1814);
and AND2 (N3864, N3856, N702);
buf BUF1 (N3865, N3827);
and AND2 (N3866, N3859, N2373);
buf BUF1 (N3867, N3824);
and AND4 (N3868, N3867, N3104, N180, N2625);
nor NOR4 (N3869, N3854, N1383, N2394, N3748);
nor NOR4 (N3870, N3865, N2002, N12, N1547);
xor XOR2 (N3871, N3861, N133);
xor XOR2 (N3872, N3869, N530);
xor XOR2 (N3873, N3851, N546);
and AND2 (N3874, N3850, N454);
buf BUF1 (N3875, N3852);
nor NOR2 (N3876, N3875, N3260);
nor NOR2 (N3877, N3868, N2724);
not NOT1 (N3878, N3872);
nand NAND4 (N3879, N3870, N852, N1933, N972);
and AND4 (N3880, N3871, N3166, N3570, N1277);
or OR4 (N3881, N3877, N2508, N2511, N3225);
nand NAND4 (N3882, N3864, N1424, N2251, N2155);
nor NOR4 (N3883, N3866, N2731, N79, N780);
nand NAND2 (N3884, N3873, N1204);
or OR2 (N3885, N3879, N559);
not NOT1 (N3886, N3885);
and AND2 (N3887, N3883, N246);
xor XOR2 (N3888, N3882, N2479);
nor NOR4 (N3889, N3876, N3152, N1037, N2892);
nand NAND4 (N3890, N3884, N3659, N1738, N2964);
xor XOR2 (N3891, N3880, N401);
nand NAND2 (N3892, N3890, N513);
not NOT1 (N3893, N3889);
nor NOR2 (N3894, N3887, N1403);
not NOT1 (N3895, N3874);
nor NOR3 (N3896, N3881, N1427, N1663);
xor XOR2 (N3897, N3894, N1373);
buf BUF1 (N3898, N3878);
buf BUF1 (N3899, N3888);
not NOT1 (N3900, N3863);
nor NOR3 (N3901, N3886, N2532, N3643);
and AND3 (N3902, N3891, N915, N3117);
nand NAND3 (N3903, N3893, N1601, N1755);
xor XOR2 (N3904, N3898, N1910);
buf BUF1 (N3905, N3892);
xor XOR2 (N3906, N3901, N2368);
not NOT1 (N3907, N3902);
xor XOR2 (N3908, N3895, N2354);
or OR3 (N3909, N3903, N506, N2624);
nand NAND4 (N3910, N3906, N1051, N929, N2386);
nor NOR2 (N3911, N3910, N2848);
nor NOR4 (N3912, N3900, N450, N2993, N3792);
buf BUF1 (N3913, N3908);
buf BUF1 (N3914, N3913);
and AND2 (N3915, N3914, N97);
nand NAND2 (N3916, N3907, N2494);
and AND4 (N3917, N3904, N2025, N2591, N2379);
nand NAND2 (N3918, N3911, N3797);
or OR2 (N3919, N3912, N2262);
or OR3 (N3920, N3909, N2859, N2476);
or OR3 (N3921, N3899, N763, N1949);
nor NOR4 (N3922, N3918, N3067, N2031, N1159);
or OR2 (N3923, N3916, N1765);
nand NAND3 (N3924, N3915, N545, N1229);
buf BUF1 (N3925, N3897);
buf BUF1 (N3926, N3924);
nor NOR3 (N3927, N3919, N3555, N1466);
nand NAND4 (N3928, N3896, N3895, N3184, N721);
buf BUF1 (N3929, N3922);
or OR3 (N3930, N3921, N3069, N2819);
and AND2 (N3931, N3917, N2999);
not NOT1 (N3932, N3926);
xor XOR2 (N3933, N3931, N1196);
not NOT1 (N3934, N3932);
buf BUF1 (N3935, N3923);
xor XOR2 (N3936, N3930, N3480);
not NOT1 (N3937, N3933);
or OR3 (N3938, N3936, N1692, N2461);
buf BUF1 (N3939, N3920);
nor NOR3 (N3940, N3937, N1629, N1883);
not NOT1 (N3941, N3929);
not NOT1 (N3942, N3925);
or OR2 (N3943, N3905, N538);
nor NOR3 (N3944, N3938, N3853, N2686);
nand NAND4 (N3945, N3941, N1730, N1370, N3622);
not NOT1 (N3946, N3939);
not NOT1 (N3947, N3927);
or OR2 (N3948, N3935, N964);
nand NAND2 (N3949, N3947, N3928);
nor NOR3 (N3950, N615, N1413, N362);
nor NOR3 (N3951, N3945, N3507, N2767);
buf BUF1 (N3952, N3942);
xor XOR2 (N3953, N3952, N3271);
xor XOR2 (N3954, N3948, N1617);
and AND3 (N3955, N3954, N1059, N2599);
or OR4 (N3956, N3944, N1408, N2254, N1603);
or OR4 (N3957, N3940, N962, N2754, N1263);
buf BUF1 (N3958, N3950);
nor NOR2 (N3959, N3949, N350);
nand NAND2 (N3960, N3953, N2336);
or OR4 (N3961, N3957, N2903, N938, N1745);
and AND3 (N3962, N3946, N1335, N3637);
nor NOR4 (N3963, N3958, N185, N2337, N332);
xor XOR2 (N3964, N3955, N2187);
or OR4 (N3965, N3964, N3214, N952, N713);
or OR4 (N3966, N3960, N1602, N792, N1501);
xor XOR2 (N3967, N3961, N2425);
xor XOR2 (N3968, N3966, N3916);
nand NAND4 (N3969, N3963, N2105, N2467, N2612);
nor NOR3 (N3970, N3968, N2941, N3064);
nand NAND4 (N3971, N3951, N164, N1080, N582);
or OR3 (N3972, N3970, N2145, N2032);
xor XOR2 (N3973, N3956, N1856);
nor NOR2 (N3974, N3973, N2771);
buf BUF1 (N3975, N3967);
buf BUF1 (N3976, N3969);
xor XOR2 (N3977, N3975, N3365);
not NOT1 (N3978, N3972);
nand NAND4 (N3979, N3959, N1037, N1933, N3033);
nor NOR4 (N3980, N3965, N3624, N2776, N1436);
xor XOR2 (N3981, N3977, N3978);
nand NAND2 (N3982, N186, N3004);
xor XOR2 (N3983, N3982, N1651);
buf BUF1 (N3984, N3979);
or OR2 (N3985, N3984, N2602);
buf BUF1 (N3986, N3971);
xor XOR2 (N3987, N3983, N1820);
and AND2 (N3988, N3981, N3381);
nand NAND2 (N3989, N3974, N1626);
nor NOR2 (N3990, N3976, N1358);
xor XOR2 (N3991, N3985, N2887);
not NOT1 (N3992, N3962);
nand NAND3 (N3993, N3990, N1206, N3958);
or OR4 (N3994, N3989, N419, N3751, N3732);
buf BUF1 (N3995, N3993);
buf BUF1 (N3996, N3991);
buf BUF1 (N3997, N3987);
nor NOR4 (N3998, N3986, N2648, N1375, N3615);
buf BUF1 (N3999, N3994);
nand NAND3 (N4000, N3998, N3519, N199);
nand NAND4 (N4001, N3999, N2502, N865, N464);
and AND3 (N4002, N3996, N1149, N2484);
nor NOR2 (N4003, N4002, N3830);
nand NAND2 (N4004, N3995, N2137);
buf BUF1 (N4005, N3980);
xor XOR2 (N4006, N4003, N2433);
xor XOR2 (N4007, N4006, N3524);
not NOT1 (N4008, N4001);
nand NAND2 (N4009, N3943, N261);
and AND3 (N4010, N3988, N198, N1757);
xor XOR2 (N4011, N4005, N931);
nor NOR2 (N4012, N3934, N2924);
nor NOR3 (N4013, N3997, N1586, N3864);
or OR2 (N4014, N4009, N2708);
not NOT1 (N4015, N4011);
xor XOR2 (N4016, N4004, N3790);
buf BUF1 (N4017, N4016);
or OR2 (N4018, N4014, N688);
nand NAND4 (N4019, N4017, N3846, N3370, N1030);
buf BUF1 (N4020, N4007);
nor NOR2 (N4021, N4008, N3766);
nor NOR2 (N4022, N4013, N3075);
buf BUF1 (N4023, N4000);
and AND2 (N4024, N4021, N2922);
or OR2 (N4025, N4024, N2020);
xor XOR2 (N4026, N4023, N3646);
buf BUF1 (N4027, N4025);
nor NOR4 (N4028, N4015, N3046, N197, N1924);
buf BUF1 (N4029, N4022);
nor NOR3 (N4030, N4018, N477, N2031);
and AND4 (N4031, N4030, N2708, N2397, N3726);
buf BUF1 (N4032, N4031);
not NOT1 (N4033, N4029);
or OR4 (N4034, N4027, N577, N268, N2587);
xor XOR2 (N4035, N4020, N2306);
nand NAND4 (N4036, N4010, N3271, N1196, N487);
nand NAND2 (N4037, N4036, N916);
nor NOR4 (N4038, N4033, N3458, N1532, N1888);
nand NAND3 (N4039, N4032, N3261, N357);
nor NOR4 (N4040, N4012, N3266, N2638, N3461);
and AND3 (N4041, N4026, N2182, N1460);
nor NOR4 (N4042, N4037, N968, N1602, N2655);
or OR2 (N4043, N4041, N1006);
not NOT1 (N4044, N4039);
or OR2 (N4045, N4043, N1729);
or OR3 (N4046, N4028, N3419, N1537);
nand NAND2 (N4047, N4044, N1747);
not NOT1 (N4048, N4047);
nand NAND2 (N4049, N4019, N994);
not NOT1 (N4050, N3992);
buf BUF1 (N4051, N4049);
and AND2 (N4052, N4045, N2732);
and AND3 (N4053, N4051, N3897, N840);
not NOT1 (N4054, N4034);
xor XOR2 (N4055, N4046, N1809);
not NOT1 (N4056, N4040);
xor XOR2 (N4057, N4056, N288);
xor XOR2 (N4058, N4035, N3342);
nand NAND2 (N4059, N4055, N1683);
and AND2 (N4060, N4059, N3158);
and AND3 (N4061, N4053, N1160, N3099);
or OR3 (N4062, N4061, N3212, N1887);
buf BUF1 (N4063, N4060);
or OR4 (N4064, N4048, N924, N3407, N1767);
or OR2 (N4065, N4063, N3054);
buf BUF1 (N4066, N4058);
not NOT1 (N4067, N4066);
nor NOR3 (N4068, N4067, N172, N1944);
not NOT1 (N4069, N4050);
xor XOR2 (N4070, N4038, N1127);
not NOT1 (N4071, N4065);
nor NOR2 (N4072, N4071, N1662);
or OR2 (N4073, N4054, N2917);
nand NAND4 (N4074, N4068, N1227, N842, N3717);
buf BUF1 (N4075, N4072);
nand NAND2 (N4076, N4057, N3717);
or OR3 (N4077, N4073, N696, N910);
nor NOR3 (N4078, N4064, N2052, N483);
and AND4 (N4079, N4052, N1303, N3144, N1297);
nand NAND4 (N4080, N4078, N3340, N3750, N199);
buf BUF1 (N4081, N4076);
xor XOR2 (N4082, N4081, N689);
nor NOR4 (N4083, N4080, N3718, N3725, N75);
and AND2 (N4084, N4070, N3288);
and AND2 (N4085, N4079, N1036);
buf BUF1 (N4086, N4085);
and AND2 (N4087, N4062, N1328);
xor XOR2 (N4088, N4086, N597);
and AND4 (N4089, N4087, N2610, N533, N3293);
xor XOR2 (N4090, N4075, N919);
and AND4 (N4091, N4042, N1760, N3001, N3740);
xor XOR2 (N4092, N4089, N3681);
and AND4 (N4093, N4088, N4026, N3165, N572);
nor NOR2 (N4094, N4091, N2947);
not NOT1 (N4095, N4094);
nor NOR2 (N4096, N4074, N312);
nor NOR2 (N4097, N4069, N2793);
or OR3 (N4098, N4095, N43, N2971);
and AND4 (N4099, N4092, N3196, N2988, N3976);
and AND3 (N4100, N4099, N371, N2512);
nor NOR3 (N4101, N4090, N1241, N3038);
not NOT1 (N4102, N4077);
not NOT1 (N4103, N4100);
or OR2 (N4104, N4102, N3688);
or OR3 (N4105, N4098, N2353, N301);
nand NAND4 (N4106, N4096, N2438, N1682, N1304);
buf BUF1 (N4107, N4093);
or OR3 (N4108, N4103, N2730, N830);
or OR2 (N4109, N4106, N3737);
nor NOR4 (N4110, N4083, N2307, N3156, N3536);
xor XOR2 (N4111, N4108, N3234);
or OR4 (N4112, N4104, N3728, N2413, N2021);
nand NAND3 (N4113, N4105, N2218, N3129);
buf BUF1 (N4114, N4082);
nand NAND4 (N4115, N4110, N822, N816, N3622);
or OR4 (N4116, N4109, N3208, N1057, N1168);
nor NOR2 (N4117, N4084, N1452);
buf BUF1 (N4118, N4116);
and AND4 (N4119, N4097, N253, N3148, N422);
nand NAND4 (N4120, N4112, N2209, N4106, N1391);
not NOT1 (N4121, N4107);
or OR2 (N4122, N4101, N3370);
not NOT1 (N4123, N4122);
nand NAND4 (N4124, N4111, N2250, N537, N1231);
buf BUF1 (N4125, N4115);
buf BUF1 (N4126, N4117);
xor XOR2 (N4127, N4113, N3725);
nand NAND3 (N4128, N4120, N1975, N35);
and AND2 (N4129, N4121, N3434);
xor XOR2 (N4130, N4114, N1224);
xor XOR2 (N4131, N4119, N1419);
or OR3 (N4132, N4123, N3723, N3105);
or OR4 (N4133, N4118, N2502, N722, N3904);
and AND2 (N4134, N4129, N857);
xor XOR2 (N4135, N4134, N615);
buf BUF1 (N4136, N4127);
xor XOR2 (N4137, N4132, N1463);
nand NAND3 (N4138, N4133, N3682, N2471);
nand NAND2 (N4139, N4130, N4074);
and AND3 (N4140, N4128, N310, N1502);
not NOT1 (N4141, N4137);
nand NAND3 (N4142, N4136, N2740, N3734);
nand NAND3 (N4143, N4125, N1250, N3447);
not NOT1 (N4144, N4135);
or OR3 (N4145, N4139, N3665, N2535);
buf BUF1 (N4146, N4142);
buf BUF1 (N4147, N4141);
or OR3 (N4148, N4145, N1644, N2526);
not NOT1 (N4149, N4131);
buf BUF1 (N4150, N4148);
xor XOR2 (N4151, N4138, N1819);
xor XOR2 (N4152, N4149, N2327);
not NOT1 (N4153, N4150);
or OR3 (N4154, N4124, N588, N2924);
buf BUF1 (N4155, N4152);
not NOT1 (N4156, N4153);
nor NOR3 (N4157, N4144, N1905, N715);
and AND4 (N4158, N4140, N3265, N95, N2906);
buf BUF1 (N4159, N4156);
not NOT1 (N4160, N4159);
not NOT1 (N4161, N4151);
xor XOR2 (N4162, N4157, N2098);
xor XOR2 (N4163, N4160, N472);
or OR3 (N4164, N4155, N3214, N816);
not NOT1 (N4165, N4161);
buf BUF1 (N4166, N4147);
nand NAND3 (N4167, N4158, N836, N3433);
not NOT1 (N4168, N4143);
nor NOR3 (N4169, N4166, N1134, N40);
not NOT1 (N4170, N4163);
not NOT1 (N4171, N4167);
xor XOR2 (N4172, N4170, N2026);
nor NOR4 (N4173, N4168, N3454, N1876, N2458);
nor NOR4 (N4174, N4173, N705, N2672, N2852);
buf BUF1 (N4175, N4171);
or OR4 (N4176, N4169, N2481, N4054, N2235);
buf BUF1 (N4177, N4175);
buf BUF1 (N4178, N4172);
buf BUF1 (N4179, N4164);
or OR3 (N4180, N4174, N1529, N2901);
and AND2 (N4181, N4154, N2443);
nand NAND3 (N4182, N4178, N1802, N3728);
nand NAND4 (N4183, N4165, N1123, N1710, N21);
and AND3 (N4184, N4176, N1922, N2414);
nand NAND4 (N4185, N4183, N3885, N1968, N3154);
nand NAND4 (N4186, N4146, N98, N1707, N86);
or OR4 (N4187, N4185, N1484, N516, N3461);
nand NAND2 (N4188, N4162, N2504);
and AND2 (N4189, N4180, N3014);
and AND4 (N4190, N4126, N210, N1860, N3238);
xor XOR2 (N4191, N4188, N1649);
xor XOR2 (N4192, N4182, N1022);
and AND4 (N4193, N4186, N3617, N1631, N201);
buf BUF1 (N4194, N4192);
not NOT1 (N4195, N4193);
buf BUF1 (N4196, N4191);
not NOT1 (N4197, N4187);
or OR2 (N4198, N4194, N3760);
xor XOR2 (N4199, N4195, N3329);
nor NOR2 (N4200, N4181, N2555);
not NOT1 (N4201, N4177);
buf BUF1 (N4202, N4200);
not NOT1 (N4203, N4201);
xor XOR2 (N4204, N4198, N903);
nand NAND4 (N4205, N4196, N2190, N716, N2333);
and AND4 (N4206, N4205, N3207, N1764, N1681);
and AND3 (N4207, N4189, N2475, N3978);
xor XOR2 (N4208, N4204, N1979);
not NOT1 (N4209, N4190);
and AND3 (N4210, N4207, N180, N3485);
and AND3 (N4211, N4209, N318, N1990);
not NOT1 (N4212, N4184);
nand NAND4 (N4213, N4206, N2974, N724, N1970);
buf BUF1 (N4214, N4208);
nor NOR2 (N4215, N4202, N632);
xor XOR2 (N4216, N4179, N134);
nor NOR3 (N4217, N4216, N866, N964);
not NOT1 (N4218, N4214);
nor NOR3 (N4219, N4218, N1858, N3396);
buf BUF1 (N4220, N4217);
nor NOR2 (N4221, N4215, N379);
or OR2 (N4222, N4221, N2706);
buf BUF1 (N4223, N4219);
buf BUF1 (N4224, N4199);
xor XOR2 (N4225, N4212, N2722);
nor NOR2 (N4226, N4224, N1350);
nand NAND3 (N4227, N4222, N3449, N2467);
xor XOR2 (N4228, N4225, N1554);
nor NOR2 (N4229, N4211, N2577);
and AND3 (N4230, N4213, N1343, N2923);
and AND4 (N4231, N4197, N1597, N2385, N3090);
nor NOR4 (N4232, N4210, N1624, N313, N3220);
buf BUF1 (N4233, N4227);
or OR3 (N4234, N4223, N2809, N3032);
buf BUF1 (N4235, N4203);
nor NOR3 (N4236, N4232, N2904, N3062);
or OR3 (N4237, N4235, N2485, N618);
xor XOR2 (N4238, N4231, N864);
xor XOR2 (N4239, N4229, N4221);
buf BUF1 (N4240, N4234);
nor NOR2 (N4241, N4220, N1557);
and AND4 (N4242, N4238, N628, N3514, N70);
xor XOR2 (N4243, N4240, N1049);
nand NAND3 (N4244, N4236, N36, N2112);
not NOT1 (N4245, N4230);
not NOT1 (N4246, N4228);
not NOT1 (N4247, N4226);
buf BUF1 (N4248, N4233);
not NOT1 (N4249, N4246);
xor XOR2 (N4250, N4247, N3669);
buf BUF1 (N4251, N4241);
xor XOR2 (N4252, N4248, N467);
and AND2 (N4253, N4244, N1742);
buf BUF1 (N4254, N4253);
and AND2 (N4255, N4250, N2092);
buf BUF1 (N4256, N4243);
and AND3 (N4257, N4255, N2874, N1806);
xor XOR2 (N4258, N4242, N777);
not NOT1 (N4259, N4258);
and AND4 (N4260, N4237, N2094, N1964, N4117);
nand NAND4 (N4261, N4239, N2845, N3933, N2431);
nand NAND2 (N4262, N4261, N3306);
buf BUF1 (N4263, N4257);
xor XOR2 (N4264, N4259, N2444);
nand NAND2 (N4265, N4245, N823);
or OR4 (N4266, N4251, N2761, N3705, N2921);
nand NAND2 (N4267, N4264, N681);
buf BUF1 (N4268, N4266);
buf BUF1 (N4269, N4256);
nand NAND2 (N4270, N4254, N2412);
not NOT1 (N4271, N4252);
xor XOR2 (N4272, N4268, N2718);
buf BUF1 (N4273, N4270);
xor XOR2 (N4274, N4262, N1886);
xor XOR2 (N4275, N4260, N649);
nand NAND3 (N4276, N4274, N629, N1590);
xor XOR2 (N4277, N4265, N2151);
not NOT1 (N4278, N4277);
and AND4 (N4279, N4249, N203, N2535, N2803);
nand NAND4 (N4280, N4275, N1743, N1991, N1330);
not NOT1 (N4281, N4263);
not NOT1 (N4282, N4267);
nand NAND3 (N4283, N4280, N2536, N3381);
buf BUF1 (N4284, N4281);
xor XOR2 (N4285, N4269, N3763);
not NOT1 (N4286, N4276);
or OR3 (N4287, N4285, N3275, N1371);
and AND2 (N4288, N4284, N2977);
or OR4 (N4289, N4279, N3108, N452, N1331);
xor XOR2 (N4290, N4287, N768);
and AND2 (N4291, N4282, N130);
and AND4 (N4292, N4273, N1046, N145, N859);
buf BUF1 (N4293, N4278);
and AND2 (N4294, N4283, N3873);
buf BUF1 (N4295, N4294);
or OR2 (N4296, N4271, N152);
nand NAND3 (N4297, N4286, N2314, N4197);
or OR3 (N4298, N4297, N1625, N683);
nor NOR2 (N4299, N4288, N1512);
and AND2 (N4300, N4291, N529);
and AND3 (N4301, N4290, N985, N1682);
nor NOR2 (N4302, N4300, N2959);
not NOT1 (N4303, N4289);
not NOT1 (N4304, N4293);
buf BUF1 (N4305, N4304);
xor XOR2 (N4306, N4296, N1898);
and AND4 (N4307, N4298, N683, N2556, N3970);
xor XOR2 (N4308, N4272, N1804);
not NOT1 (N4309, N4303);
or OR2 (N4310, N4306, N3581);
nor NOR2 (N4311, N4305, N3633);
not NOT1 (N4312, N4309);
nor NOR3 (N4313, N4301, N3836, N26);
xor XOR2 (N4314, N4292, N3191);
xor XOR2 (N4315, N4313, N3946);
and AND3 (N4316, N4311, N1045, N2454);
not NOT1 (N4317, N4314);
or OR2 (N4318, N4312, N1425);
buf BUF1 (N4319, N4302);
nor NOR4 (N4320, N4299, N1377, N1584, N1428);
nand NAND2 (N4321, N4295, N268);
and AND2 (N4322, N4307, N4032);
buf BUF1 (N4323, N4319);
and AND4 (N4324, N4322, N770, N2176, N1827);
buf BUF1 (N4325, N4320);
or OR3 (N4326, N4308, N222, N2050);
and AND3 (N4327, N4326, N2291, N3195);
buf BUF1 (N4328, N4317);
not NOT1 (N4329, N4310);
or OR3 (N4330, N4328, N2195, N4063);
not NOT1 (N4331, N4330);
or OR3 (N4332, N4325, N22, N4218);
nand NAND4 (N4333, N4318, N3636, N3778, N887);
buf BUF1 (N4334, N4323);
buf BUF1 (N4335, N4331);
nor NOR3 (N4336, N4332, N2201, N3249);
nor NOR2 (N4337, N4336, N2774);
buf BUF1 (N4338, N4316);
and AND3 (N4339, N4329, N3443, N2755);
and AND2 (N4340, N4315, N1084);
and AND4 (N4341, N4337, N3135, N2671, N2735);
buf BUF1 (N4342, N4321);
xor XOR2 (N4343, N4339, N187);
and AND4 (N4344, N4338, N3202, N3032, N2850);
buf BUF1 (N4345, N4344);
nand NAND4 (N4346, N4333, N2557, N1619, N2167);
or OR3 (N4347, N4346, N1017, N1716);
not NOT1 (N4348, N4327);
or OR4 (N4349, N4341, N1741, N2678, N500);
buf BUF1 (N4350, N4334);
nand NAND3 (N4351, N4348, N2422, N1002);
not NOT1 (N4352, N4340);
not NOT1 (N4353, N4351);
xor XOR2 (N4354, N4324, N1940);
nand NAND2 (N4355, N4354, N1108);
and AND3 (N4356, N4345, N1565, N650);
or OR4 (N4357, N4352, N3664, N771, N2637);
not NOT1 (N4358, N4350);
nand NAND3 (N4359, N4349, N2863, N4109);
nand NAND4 (N4360, N4347, N2930, N419, N1823);
nand NAND3 (N4361, N4356, N2426, N2618);
nand NAND2 (N4362, N4342, N2556);
xor XOR2 (N4363, N4355, N1252);
nor NOR2 (N4364, N4359, N2172);
not NOT1 (N4365, N4343);
nand NAND4 (N4366, N4364, N478, N3692, N1086);
and AND3 (N4367, N4366, N2950, N2620);
buf BUF1 (N4368, N4335);
or OR2 (N4369, N4367, N1778);
nand NAND3 (N4370, N4369, N744, N1829);
xor XOR2 (N4371, N4357, N4069);
or OR2 (N4372, N4358, N2015);
xor XOR2 (N4373, N4365, N1166);
xor XOR2 (N4374, N4368, N2722);
buf BUF1 (N4375, N4373);
and AND3 (N4376, N4371, N3289, N296);
or OR4 (N4377, N4360, N1287, N3634, N149);
buf BUF1 (N4378, N4376);
xor XOR2 (N4379, N4362, N2042);
buf BUF1 (N4380, N4374);
nand NAND3 (N4381, N4380, N281, N604);
buf BUF1 (N4382, N4361);
buf BUF1 (N4383, N4382);
nor NOR4 (N4384, N4363, N1046, N117, N3902);
xor XOR2 (N4385, N4370, N4004);
nor NOR4 (N4386, N4377, N4015, N2282, N400);
and AND4 (N4387, N4385, N796, N1786, N3756);
nor NOR2 (N4388, N4378, N3538);
xor XOR2 (N4389, N4388, N665);
and AND4 (N4390, N4353, N3912, N2958, N1777);
not NOT1 (N4391, N4390);
not NOT1 (N4392, N4384);
nand NAND2 (N4393, N4386, N2345);
and AND2 (N4394, N4381, N1825);
buf BUF1 (N4395, N4393);
xor XOR2 (N4396, N4394, N1400);
buf BUF1 (N4397, N4392);
and AND3 (N4398, N4372, N2429, N3905);
buf BUF1 (N4399, N4397);
buf BUF1 (N4400, N4399);
nand NAND4 (N4401, N4396, N1692, N799, N4031);
not NOT1 (N4402, N4395);
xor XOR2 (N4403, N4402, N664);
or OR3 (N4404, N4379, N2465, N4199);
buf BUF1 (N4405, N4404);
or OR4 (N4406, N4398, N2123, N1875, N1014);
and AND2 (N4407, N4403, N2544);
not NOT1 (N4408, N4387);
or OR3 (N4409, N4389, N3671, N1328);
not NOT1 (N4410, N4408);
xor XOR2 (N4411, N4383, N468);
and AND4 (N4412, N4410, N3884, N2835, N2047);
nand NAND4 (N4413, N4401, N1749, N1086, N2480);
buf BUF1 (N4414, N4400);
xor XOR2 (N4415, N4391, N692);
buf BUF1 (N4416, N4413);
nand NAND2 (N4417, N4416, N1982);
or OR3 (N4418, N4412, N3962, N1193);
and AND2 (N4419, N4407, N647);
nor NOR2 (N4420, N4375, N3291);
not NOT1 (N4421, N4418);
and AND4 (N4422, N4405, N1451, N2877, N3195);
xor XOR2 (N4423, N4406, N80);
buf BUF1 (N4424, N4420);
buf BUF1 (N4425, N4424);
or OR4 (N4426, N4422, N1571, N2339, N639);
or OR4 (N4427, N4419, N2601, N3019, N4021);
nor NOR3 (N4428, N4417, N341, N3253);
buf BUF1 (N4429, N4414);
and AND4 (N4430, N4429, N2659, N1548, N10);
xor XOR2 (N4431, N4423, N284);
not NOT1 (N4432, N4427);
or OR2 (N4433, N4432, N220);
xor XOR2 (N4434, N4430, N4068);
nand NAND3 (N4435, N4421, N3744, N3378);
not NOT1 (N4436, N4435);
xor XOR2 (N4437, N4431, N3874);
nor NOR4 (N4438, N4436, N2630, N2269, N3371);
nand NAND3 (N4439, N4434, N347, N3941);
not NOT1 (N4440, N4425);
and AND3 (N4441, N4411, N4409, N600);
buf BUF1 (N4442, N1360);
not NOT1 (N4443, N4442);
nor NOR4 (N4444, N4433, N4434, N1745, N2234);
not NOT1 (N4445, N4440);
xor XOR2 (N4446, N4443, N2527);
nand NAND2 (N4447, N4439, N2103);
and AND2 (N4448, N4441, N2452);
nand NAND3 (N4449, N4415, N1671, N4398);
and AND3 (N4450, N4446, N4045, N2525);
nor NOR2 (N4451, N4448, N3046);
nor NOR3 (N4452, N4451, N1135, N1987);
or OR2 (N4453, N4452, N1082);
and AND4 (N4454, N4426, N495, N1848, N51);
or OR3 (N4455, N4428, N4453, N3584);
nor NOR4 (N4456, N3478, N2550, N919, N1412);
buf BUF1 (N4457, N4456);
buf BUF1 (N4458, N4445);
xor XOR2 (N4459, N4447, N4210);
or OR3 (N4460, N4458, N4128, N155);
buf BUF1 (N4461, N4459);
not NOT1 (N4462, N4460);
not NOT1 (N4463, N4438);
and AND2 (N4464, N4437, N1368);
not NOT1 (N4465, N4444);
buf BUF1 (N4466, N4461);
nand NAND3 (N4467, N4465, N961, N1172);
not NOT1 (N4468, N4466);
or OR2 (N4469, N4455, N3453);
or OR4 (N4470, N4462, N497, N1277, N4180);
not NOT1 (N4471, N4454);
or OR3 (N4472, N4463, N2437, N212);
or OR2 (N4473, N4464, N3902);
or OR3 (N4474, N4449, N3174, N3285);
xor XOR2 (N4475, N4470, N998);
buf BUF1 (N4476, N4467);
not NOT1 (N4477, N4476);
buf BUF1 (N4478, N4469);
or OR4 (N4479, N4457, N774, N4165, N122);
or OR4 (N4480, N4450, N4208, N1735, N2033);
nor NOR3 (N4481, N4479, N1803, N3051);
not NOT1 (N4482, N4471);
or OR2 (N4483, N4481, N353);
xor XOR2 (N4484, N4483, N4042);
and AND3 (N4485, N4478, N1208, N729);
xor XOR2 (N4486, N4480, N1588);
nand NAND4 (N4487, N4468, N144, N4477, N4385);
xor XOR2 (N4488, N4009, N1914);
nand NAND4 (N4489, N4484, N1119, N3723, N1887);
or OR3 (N4490, N4487, N3433, N2553);
not NOT1 (N4491, N4486);
xor XOR2 (N4492, N4488, N1331);
xor XOR2 (N4493, N4472, N3551);
or OR4 (N4494, N4473, N1801, N1578, N873);
buf BUF1 (N4495, N4489);
not NOT1 (N4496, N4490);
or OR3 (N4497, N4491, N227, N3125);
or OR2 (N4498, N4494, N103);
not NOT1 (N4499, N4496);
nand NAND2 (N4500, N4475, N3856);
not NOT1 (N4501, N4497);
and AND4 (N4502, N4492, N1183, N1595, N2689);
not NOT1 (N4503, N4498);
nand NAND2 (N4504, N4474, N3875);
nor NOR4 (N4505, N4485, N3362, N1415, N4318);
not NOT1 (N4506, N4504);
and AND2 (N4507, N4495, N896);
or OR3 (N4508, N4507, N3043, N3048);
or OR4 (N4509, N4503, N2724, N4233, N1098);
xor XOR2 (N4510, N4482, N1315);
not NOT1 (N4511, N4502);
xor XOR2 (N4512, N4511, N465);
or OR2 (N4513, N4510, N3911);
buf BUF1 (N4514, N4509);
or OR2 (N4515, N4514, N1917);
not NOT1 (N4516, N4513);
and AND2 (N4517, N4508, N477);
buf BUF1 (N4518, N4512);
buf BUF1 (N4519, N4517);
buf BUF1 (N4520, N4493);
and AND2 (N4521, N4506, N3639);
or OR2 (N4522, N4516, N1537);
or OR2 (N4523, N4500, N3911);
nor NOR2 (N4524, N4523, N3787);
buf BUF1 (N4525, N4521);
or OR3 (N4526, N4518, N377, N4238);
not NOT1 (N4527, N4522);
buf BUF1 (N4528, N4501);
nor NOR4 (N4529, N4519, N3752, N345, N1296);
or OR2 (N4530, N4526, N4374);
xor XOR2 (N4531, N4515, N3393);
or OR2 (N4532, N4529, N3609);
xor XOR2 (N4533, N4520, N73);
buf BUF1 (N4534, N4533);
buf BUF1 (N4535, N4499);
buf BUF1 (N4536, N4534);
and AND2 (N4537, N4536, N2582);
or OR4 (N4538, N4505, N487, N891, N1591);
or OR2 (N4539, N4527, N3651);
not NOT1 (N4540, N4525);
not NOT1 (N4541, N4524);
buf BUF1 (N4542, N4535);
or OR2 (N4543, N4530, N3438);
nor NOR4 (N4544, N4542, N803, N2542, N2390);
or OR4 (N4545, N4531, N709, N2255, N707);
nand NAND2 (N4546, N4528, N4120);
and AND2 (N4547, N4546, N3920);
nand NAND4 (N4548, N4540, N2996, N487, N1757);
not NOT1 (N4549, N4548);
or OR4 (N4550, N4549, N2828, N614, N3465);
nor NOR4 (N4551, N4547, N2361, N3427, N1529);
xor XOR2 (N4552, N4545, N3255);
nor NOR4 (N4553, N4551, N2382, N2040, N2145);
xor XOR2 (N4554, N4541, N46);
nand NAND2 (N4555, N4554, N565);
buf BUF1 (N4556, N4543);
nand NAND3 (N4557, N4532, N49, N1736);
not NOT1 (N4558, N4539);
not NOT1 (N4559, N4556);
nor NOR2 (N4560, N4553, N1331);
nand NAND4 (N4561, N4557, N4228, N3871, N4243);
and AND3 (N4562, N4538, N992, N3757);
or OR4 (N4563, N4560, N1759, N282, N1139);
not NOT1 (N4564, N4561);
nor NOR3 (N4565, N4552, N1901, N1592);
buf BUF1 (N4566, N4565);
nor NOR4 (N4567, N4537, N4300, N2767, N787);
not NOT1 (N4568, N4563);
nand NAND4 (N4569, N4568, N1940, N2196, N3209);
buf BUF1 (N4570, N4564);
not NOT1 (N4571, N4544);
not NOT1 (N4572, N4550);
nor NOR2 (N4573, N4572, N2007);
buf BUF1 (N4574, N4559);
nor NOR3 (N4575, N4562, N3191, N3498);
not NOT1 (N4576, N4575);
or OR4 (N4577, N4558, N3803, N864, N920);
nand NAND3 (N4578, N4569, N3466, N865);
or OR2 (N4579, N4574, N276);
nand NAND3 (N4580, N4578, N1612, N1265);
and AND2 (N4581, N4573, N1656);
and AND2 (N4582, N4555, N2403);
not NOT1 (N4583, N4582);
or OR3 (N4584, N4579, N3131, N1107);
buf BUF1 (N4585, N4584);
or OR2 (N4586, N4566, N2246);
or OR4 (N4587, N4585, N4236, N2963, N1424);
not NOT1 (N4588, N4586);
buf BUF1 (N4589, N4571);
nor NOR2 (N4590, N4570, N4077);
or OR4 (N4591, N4581, N3490, N2900, N1632);
and AND4 (N4592, N4576, N3915, N1355, N3080);
buf BUF1 (N4593, N4590);
nor NOR2 (N4594, N4580, N1812);
not NOT1 (N4595, N4583);
nor NOR2 (N4596, N4587, N3432);
buf BUF1 (N4597, N4591);
xor XOR2 (N4598, N4592, N2377);
nand NAND3 (N4599, N4593, N3369, N3321);
xor XOR2 (N4600, N4596, N591);
and AND2 (N4601, N4600, N2742);
or OR4 (N4602, N4598, N4158, N2625, N1881);
and AND4 (N4603, N4588, N2436, N3576, N2844);
xor XOR2 (N4604, N4594, N170);
not NOT1 (N4605, N4601);
or OR2 (N4606, N4605, N540);
nor NOR2 (N4607, N4606, N3287);
not NOT1 (N4608, N4599);
nor NOR3 (N4609, N4597, N1457, N2593);
buf BUF1 (N4610, N4577);
nand NAND2 (N4611, N4610, N185);
and AND4 (N4612, N4567, N2904, N2902, N1476);
not NOT1 (N4613, N4595);
not NOT1 (N4614, N4611);
not NOT1 (N4615, N4604);
nand NAND3 (N4616, N4609, N4255, N1095);
not NOT1 (N4617, N4612);
nand NAND3 (N4618, N4617, N1336, N349);
and AND3 (N4619, N4607, N1329, N4113);
buf BUF1 (N4620, N4616);
or OR2 (N4621, N4608, N443);
buf BUF1 (N4622, N4614);
or OR2 (N4623, N4622, N1318);
and AND2 (N4624, N4619, N2166);
and AND3 (N4625, N4615, N2170, N2203);
and AND4 (N4626, N4624, N3348, N63, N3286);
not NOT1 (N4627, N4613);
buf BUF1 (N4628, N4618);
xor XOR2 (N4629, N4589, N854);
and AND3 (N4630, N4621, N1879, N2275);
not NOT1 (N4631, N4629);
not NOT1 (N4632, N4628);
and AND3 (N4633, N4623, N1408, N3780);
and AND2 (N4634, N4627, N3076);
xor XOR2 (N4635, N4633, N3692);
nor NOR2 (N4636, N4632, N4496);
not NOT1 (N4637, N4631);
or OR2 (N4638, N4637, N2683);
or OR4 (N4639, N4602, N1240, N2477, N4327);
nand NAND4 (N4640, N4635, N116, N1838, N766);
nand NAND4 (N4641, N4639, N827, N901, N4075);
xor XOR2 (N4642, N4640, N2264);
nand NAND2 (N4643, N4641, N1100);
nand NAND2 (N4644, N4630, N3563);
or OR3 (N4645, N4626, N1452, N3793);
not NOT1 (N4646, N4625);
nand NAND2 (N4647, N4645, N1385);
nand NAND4 (N4648, N4647, N2160, N2629, N2193);
not NOT1 (N4649, N4620);
or OR3 (N4650, N4636, N676, N3341);
nor NOR2 (N4651, N4642, N39);
buf BUF1 (N4652, N4644);
or OR2 (N4653, N4634, N3748);
nor NOR4 (N4654, N4650, N3658, N1634, N4267);
nor NOR3 (N4655, N4638, N862, N4372);
not NOT1 (N4656, N4651);
buf BUF1 (N4657, N4649);
buf BUF1 (N4658, N4654);
or OR3 (N4659, N4652, N4463, N2015);
xor XOR2 (N4660, N4655, N631);
and AND4 (N4661, N4658, N3750, N3198, N2014);
or OR2 (N4662, N4648, N2339);
xor XOR2 (N4663, N4653, N2351);
nor NOR3 (N4664, N4643, N2071, N3291);
nand NAND3 (N4665, N4661, N3805, N3961);
nor NOR3 (N4666, N4663, N2078, N2308);
nand NAND3 (N4667, N4657, N3412, N3146);
xor XOR2 (N4668, N4646, N1424);
nor NOR4 (N4669, N4660, N259, N2524, N375);
buf BUF1 (N4670, N4659);
buf BUF1 (N4671, N4670);
or OR4 (N4672, N4656, N3269, N454, N4405);
or OR2 (N4673, N4603, N2606);
and AND4 (N4674, N4664, N3536, N3960, N3053);
or OR3 (N4675, N4665, N2731, N2150);
xor XOR2 (N4676, N4675, N4113);
not NOT1 (N4677, N4671);
xor XOR2 (N4678, N4666, N1936);
and AND3 (N4679, N4676, N2210, N2878);
or OR3 (N4680, N4669, N3396, N1705);
nand NAND3 (N4681, N4680, N4216, N2770);
not NOT1 (N4682, N4679);
or OR2 (N4683, N4673, N4369);
and AND4 (N4684, N4662, N3155, N743, N4310);
buf BUF1 (N4685, N4674);
and AND4 (N4686, N4682, N1038, N2575, N3280);
and AND3 (N4687, N4672, N4364, N2209);
or OR2 (N4688, N4685, N442);
or OR2 (N4689, N4668, N4051);
and AND3 (N4690, N4687, N1722, N2995);
buf BUF1 (N4691, N4678);
and AND4 (N4692, N4667, N3950, N40, N2941);
buf BUF1 (N4693, N4683);
and AND4 (N4694, N4688, N4284, N2498, N1302);
nor NOR3 (N4695, N4693, N3079, N935);
xor XOR2 (N4696, N4681, N3487);
xor XOR2 (N4697, N4692, N2676);
buf BUF1 (N4698, N4690);
nand NAND4 (N4699, N4686, N2956, N4014, N624);
buf BUF1 (N4700, N4697);
xor XOR2 (N4701, N4700, N1819);
xor XOR2 (N4702, N4698, N2355);
not NOT1 (N4703, N4684);
nor NOR2 (N4704, N4702, N867);
xor XOR2 (N4705, N4696, N1073);
or OR3 (N4706, N4694, N4489, N3834);
nor NOR4 (N4707, N4701, N2163, N2786, N3482);
nand NAND2 (N4708, N4677, N3638);
or OR2 (N4709, N4699, N880);
buf BUF1 (N4710, N4705);
nand NAND4 (N4711, N4695, N1630, N972, N55);
or OR4 (N4712, N4711, N2789, N1769, N4393);
buf BUF1 (N4713, N4706);
or OR2 (N4714, N4691, N2863);
buf BUF1 (N4715, N4703);
not NOT1 (N4716, N4712);
xor XOR2 (N4717, N4716, N2645);
buf BUF1 (N4718, N4717);
nand NAND2 (N4719, N4707, N3093);
nand NAND3 (N4720, N4713, N3654, N2416);
nor NOR2 (N4721, N4714, N3033);
and AND4 (N4722, N4721, N3068, N2735, N424);
nand NAND2 (N4723, N4710, N269);
not NOT1 (N4724, N4709);
nand NAND3 (N4725, N4723, N796, N1960);
not NOT1 (N4726, N4689);
nor NOR2 (N4727, N4704, N2557);
nand NAND3 (N4728, N4725, N451, N2405);
and AND3 (N4729, N4728, N510, N1100);
xor XOR2 (N4730, N4722, N4717);
nand NAND4 (N4731, N4718, N1760, N3583, N1413);
nor NOR2 (N4732, N4730, N1662);
nand NAND2 (N4733, N4708, N1219);
buf BUF1 (N4734, N4715);
xor XOR2 (N4735, N4727, N394);
nor NOR2 (N4736, N4734, N3971);
nor NOR4 (N4737, N4735, N4666, N1526, N3944);
or OR2 (N4738, N4736, N4204);
or OR4 (N4739, N4726, N4182, N2638, N1258);
nor NOR4 (N4740, N4724, N1243, N1288, N2058);
nand NAND3 (N4741, N4733, N955, N1526);
buf BUF1 (N4742, N4719);
xor XOR2 (N4743, N4720, N1851);
xor XOR2 (N4744, N4740, N2505);
xor XOR2 (N4745, N4737, N2600);
and AND2 (N4746, N4744, N3670);
nor NOR2 (N4747, N4745, N3343);
not NOT1 (N4748, N4741);
not NOT1 (N4749, N4748);
nand NAND3 (N4750, N4732, N141, N1009);
xor XOR2 (N4751, N4729, N1711);
and AND4 (N4752, N4731, N2315, N4190, N3591);
xor XOR2 (N4753, N4750, N338);
xor XOR2 (N4754, N4746, N413);
nand NAND3 (N4755, N4738, N4132, N4575);
nor NOR3 (N4756, N4752, N3098, N705);
or OR2 (N4757, N4756, N195);
and AND3 (N4758, N4757, N1619, N952);
nand NAND4 (N4759, N4742, N1835, N542, N47);
xor XOR2 (N4760, N4755, N2999);
nor NOR2 (N4761, N4751, N1892);
nor NOR4 (N4762, N4754, N3191, N2121, N4095);
xor XOR2 (N4763, N4739, N3007);
nor NOR2 (N4764, N4762, N657);
and AND3 (N4765, N4743, N55, N4525);
or OR3 (N4766, N4763, N3457, N4349);
nor NOR4 (N4767, N4766, N2383, N1441, N2479);
xor XOR2 (N4768, N4749, N1832);
nand NAND2 (N4769, N4759, N3683);
buf BUF1 (N4770, N4753);
nor NOR2 (N4771, N4769, N4283);
and AND2 (N4772, N4770, N4476);
buf BUF1 (N4773, N4761);
buf BUF1 (N4774, N4765);
or OR4 (N4775, N4772, N1057, N2396, N1026);
not NOT1 (N4776, N4764);
nand NAND4 (N4777, N4773, N2743, N1723, N1576);
nand NAND3 (N4778, N4776, N1949, N3635);
not NOT1 (N4779, N4747);
xor XOR2 (N4780, N4767, N4736);
xor XOR2 (N4781, N4778, N1458);
nand NAND4 (N4782, N4760, N1377, N4564, N2672);
nand NAND2 (N4783, N4781, N1992);
xor XOR2 (N4784, N4777, N655);
buf BUF1 (N4785, N4782);
and AND2 (N4786, N4774, N4337);
not NOT1 (N4787, N4779);
not NOT1 (N4788, N4787);
not NOT1 (N4789, N4786);
xor XOR2 (N4790, N4789, N1126);
buf BUF1 (N4791, N4783);
nor NOR2 (N4792, N4790, N2070);
and AND3 (N4793, N4784, N394, N3527);
xor XOR2 (N4794, N4771, N1621);
nand NAND4 (N4795, N4780, N3784, N1086, N1635);
xor XOR2 (N4796, N4788, N4052);
xor XOR2 (N4797, N4794, N239);
not NOT1 (N4798, N4785);
nand NAND3 (N4799, N4798, N2783, N3975);
not NOT1 (N4800, N4792);
nand NAND4 (N4801, N4758, N3427, N1163, N3633);
nand NAND2 (N4802, N4793, N1237);
and AND2 (N4803, N4800, N3284);
buf BUF1 (N4804, N4796);
xor XOR2 (N4805, N4791, N2237);
not NOT1 (N4806, N4802);
buf BUF1 (N4807, N4775);
or OR3 (N4808, N4799, N2547, N1400);
xor XOR2 (N4809, N4808, N310);
buf BUF1 (N4810, N4804);
nor NOR4 (N4811, N4803, N565, N551, N2206);
xor XOR2 (N4812, N4806, N4376);
buf BUF1 (N4813, N4812);
buf BUF1 (N4814, N4768);
nor NOR4 (N4815, N4810, N119, N2024, N3617);
or OR3 (N4816, N4801, N1385, N2734);
nand NAND2 (N4817, N4815, N2929);
buf BUF1 (N4818, N4814);
buf BUF1 (N4819, N4807);
and AND2 (N4820, N4819, N1914);
buf BUF1 (N4821, N4817);
nor NOR2 (N4822, N4821, N2012);
not NOT1 (N4823, N4816);
xor XOR2 (N4824, N4797, N3443);
nand NAND4 (N4825, N4822, N455, N3297, N4259);
nand NAND4 (N4826, N4824, N131, N246, N518);
not NOT1 (N4827, N4823);
or OR4 (N4828, N4811, N2374, N3368, N338);
not NOT1 (N4829, N4826);
nor NOR4 (N4830, N4795, N3344, N1451, N2190);
xor XOR2 (N4831, N4829, N2544);
not NOT1 (N4832, N4818);
not NOT1 (N4833, N4825);
xor XOR2 (N4834, N4813, N1068);
not NOT1 (N4835, N4809);
buf BUF1 (N4836, N4835);
not NOT1 (N4837, N4827);
xor XOR2 (N4838, N4836, N2231);
or OR4 (N4839, N4831, N4833, N486, N2191);
not NOT1 (N4840, N2172);
xor XOR2 (N4841, N4830, N1597);
and AND2 (N4842, N4832, N3639);
nand NAND4 (N4843, N4840, N54, N545, N1512);
and AND2 (N4844, N4839, N4101);
or OR2 (N4845, N4805, N449);
nand NAND2 (N4846, N4842, N3912);
nand NAND2 (N4847, N4837, N2020);
and AND4 (N4848, N4834, N3503, N42, N1269);
xor XOR2 (N4849, N4846, N1945);
nand NAND4 (N4850, N4820, N3008, N1957, N3882);
nor NOR2 (N4851, N4845, N1013);
buf BUF1 (N4852, N4848);
not NOT1 (N4853, N4851);
or OR3 (N4854, N4841, N3950, N2561);
or OR3 (N4855, N4850, N1641, N1731);
or OR3 (N4856, N4847, N3296, N3356);
nand NAND3 (N4857, N4828, N2446, N34);
or OR3 (N4858, N4855, N3245, N4795);
or OR2 (N4859, N4852, N1211);
or OR3 (N4860, N4856, N836, N343);
nand NAND2 (N4861, N4860, N4102);
buf BUF1 (N4862, N4853);
nand NAND4 (N4863, N4844, N1120, N512, N2098);
nor NOR4 (N4864, N4863, N14, N1979, N1551);
not NOT1 (N4865, N4843);
nor NOR3 (N4866, N4865, N2042, N4211);
nand NAND3 (N4867, N4857, N4747, N170);
nor NOR4 (N4868, N4861, N4866, N443, N1352);
or OR3 (N4869, N4679, N1888, N139);
buf BUF1 (N4870, N4858);
not NOT1 (N4871, N4868);
buf BUF1 (N4872, N4864);
buf BUF1 (N4873, N4872);
buf BUF1 (N4874, N4854);
nand NAND3 (N4875, N4838, N547, N3920);
not NOT1 (N4876, N4873);
nand NAND4 (N4877, N4862, N806, N969, N4441);
nor NOR2 (N4878, N4877, N92);
and AND3 (N4879, N4849, N3133, N2577);
nor NOR3 (N4880, N4859, N4041, N2112);
nand NAND2 (N4881, N4867, N2634);
or OR2 (N4882, N4871, N3915);
nor NOR4 (N4883, N4880, N4508, N1619, N4496);
not NOT1 (N4884, N4874);
nor NOR4 (N4885, N4884, N3687, N164, N171);
nor NOR4 (N4886, N4881, N1643, N78, N289);
or OR4 (N4887, N4879, N2349, N301, N4842);
or OR3 (N4888, N4876, N2091, N120);
xor XOR2 (N4889, N4878, N2992);
nand NAND3 (N4890, N4888, N4353, N1957);
buf BUF1 (N4891, N4889);
and AND3 (N4892, N4890, N2590, N4508);
xor XOR2 (N4893, N4891, N3800);
or OR4 (N4894, N4883, N2656, N1292, N4298);
xor XOR2 (N4895, N4870, N1139);
nor NOR3 (N4896, N4886, N2917, N4691);
xor XOR2 (N4897, N4885, N2704);
xor XOR2 (N4898, N4896, N4647);
buf BUF1 (N4899, N4869);
xor XOR2 (N4900, N4895, N536);
xor XOR2 (N4901, N4893, N2188);
not NOT1 (N4902, N4900);
buf BUF1 (N4903, N4894);
xor XOR2 (N4904, N4887, N1138);
nor NOR3 (N4905, N4899, N4435, N1180);
nand NAND4 (N4906, N4903, N1040, N3808, N3940);
nand NAND3 (N4907, N4902, N2753, N3402);
not NOT1 (N4908, N4901);
not NOT1 (N4909, N4905);
not NOT1 (N4910, N4875);
xor XOR2 (N4911, N4904, N1825);
xor XOR2 (N4912, N4906, N2428);
nand NAND2 (N4913, N4911, N2227);
nor NOR3 (N4914, N4909, N2030, N2140);
xor XOR2 (N4915, N4910, N1408);
nand NAND2 (N4916, N4913, N4256);
xor XOR2 (N4917, N4882, N367);
or OR2 (N4918, N4897, N3782);
not NOT1 (N4919, N4912);
not NOT1 (N4920, N4908);
or OR3 (N4921, N4898, N4485, N3554);
buf BUF1 (N4922, N4918);
xor XOR2 (N4923, N4917, N470);
and AND2 (N4924, N4920, N63);
nor NOR4 (N4925, N4919, N814, N1898, N874);
or OR4 (N4926, N4924, N4219, N4755, N3334);
and AND4 (N4927, N4925, N92, N165, N4662);
xor XOR2 (N4928, N4914, N2490);
nand NAND3 (N4929, N4921, N3756, N2092);
nor NOR4 (N4930, N4929, N2728, N689, N3629);
xor XOR2 (N4931, N4892, N3658);
not NOT1 (N4932, N4923);
xor XOR2 (N4933, N4931, N1852);
buf BUF1 (N4934, N4932);
nor NOR2 (N4935, N4926, N2335);
not NOT1 (N4936, N4927);
and AND3 (N4937, N4915, N1046, N440);
not NOT1 (N4938, N4916);
buf BUF1 (N4939, N4907);
not NOT1 (N4940, N4934);
nand NAND4 (N4941, N4930, N3747, N881, N2662);
buf BUF1 (N4942, N4939);
or OR2 (N4943, N4937, N2374);
and AND2 (N4944, N4943, N470);
not NOT1 (N4945, N4940);
nor NOR4 (N4946, N4935, N254, N4458, N1026);
nand NAND2 (N4947, N4936, N429);
not NOT1 (N4948, N4942);
nand NAND3 (N4949, N4944, N2973, N3775);
nor NOR4 (N4950, N4945, N4308, N4222, N2616);
or OR3 (N4951, N4949, N3295, N852);
xor XOR2 (N4952, N4946, N4700);
nor NOR3 (N4953, N4933, N2144, N1119);
buf BUF1 (N4954, N4952);
xor XOR2 (N4955, N4950, N1022);
xor XOR2 (N4956, N4954, N2408);
not NOT1 (N4957, N4951);
or OR3 (N4958, N4947, N1366, N3261);
and AND4 (N4959, N4955, N2155, N3270, N4215);
buf BUF1 (N4960, N4922);
not NOT1 (N4961, N4948);
nor NOR3 (N4962, N4953, N343, N2344);
not NOT1 (N4963, N4928);
xor XOR2 (N4964, N4961, N4962);
or OR3 (N4965, N970, N3338, N3302);
or OR4 (N4966, N4957, N3243, N4339, N3377);
not NOT1 (N4967, N4960);
nor NOR3 (N4968, N4959, N1492, N2479);
buf BUF1 (N4969, N4958);
xor XOR2 (N4970, N4968, N1870);
and AND2 (N4971, N4956, N219);
not NOT1 (N4972, N4941);
not NOT1 (N4973, N4938);
not NOT1 (N4974, N4970);
or OR3 (N4975, N4974, N1703, N1155);
not NOT1 (N4976, N4967);
nand NAND4 (N4977, N4965, N3227, N83, N2135);
nor NOR4 (N4978, N4972, N819, N1261, N4831);
not NOT1 (N4979, N4971);
buf BUF1 (N4980, N4978);
xor XOR2 (N4981, N4980, N763);
buf BUF1 (N4982, N4973);
not NOT1 (N4983, N4976);
not NOT1 (N4984, N4963);
xor XOR2 (N4985, N4977, N2169);
nor NOR2 (N4986, N4964, N2852);
and AND3 (N4987, N4969, N4438, N3586);
or OR2 (N4988, N4986, N4680);
not NOT1 (N4989, N4975);
nand NAND4 (N4990, N4989, N1615, N98, N614);
or OR4 (N4991, N4979, N3554, N1484, N2381);
nor NOR2 (N4992, N4984, N2295);
and AND2 (N4993, N4982, N212);
or OR4 (N4994, N4987, N4472, N4486, N1049);
and AND2 (N4995, N4994, N1821);
or OR4 (N4996, N4985, N3588, N3948, N4717);
and AND2 (N4997, N4988, N959);
nor NOR4 (N4998, N4993, N3394, N1745, N683);
not NOT1 (N4999, N4996);
or OR2 (N5000, N4997, N1290);
buf BUF1 (N5001, N4992);
buf BUF1 (N5002, N4991);
buf BUF1 (N5003, N4998);
buf BUF1 (N5004, N4983);
buf BUF1 (N5005, N5002);
nor NOR2 (N5006, N4966, N1708);
buf BUF1 (N5007, N5003);
or OR3 (N5008, N4990, N1237, N2187);
xor XOR2 (N5009, N5006, N3034);
or OR3 (N5010, N4981, N4651, N2882);
buf BUF1 (N5011, N5000);
buf BUF1 (N5012, N5011);
buf BUF1 (N5013, N5004);
nand NAND3 (N5014, N5013, N2315, N3976);
xor XOR2 (N5015, N5005, N941);
xor XOR2 (N5016, N5007, N4859);
or OR4 (N5017, N5010, N1562, N1432, N4722);
nor NOR4 (N5018, N5016, N878, N1538, N2383);
buf BUF1 (N5019, N5018);
buf BUF1 (N5020, N4999);
xor XOR2 (N5021, N5017, N2191);
not NOT1 (N5022, N5021);
and AND4 (N5023, N5015, N1329, N2234, N2519);
not NOT1 (N5024, N5009);
and AND3 (N5025, N5024, N3281, N2091);
nor NOR2 (N5026, N5019, N5025);
or OR3 (N5027, N182, N72, N802);
buf BUF1 (N5028, N4995);
nor NOR2 (N5029, N5026, N3031);
and AND2 (N5030, N5027, N1553);
or OR4 (N5031, N5028, N2047, N3272, N719);
and AND2 (N5032, N5012, N3420);
and AND2 (N5033, N5030, N3405);
xor XOR2 (N5034, N5020, N1588);
nor NOR4 (N5035, N5029, N3089, N2326, N1686);
xor XOR2 (N5036, N5031, N4194);
nor NOR4 (N5037, N5008, N60, N2891, N3490);
buf BUF1 (N5038, N5032);
xor XOR2 (N5039, N5033, N2501);
or OR2 (N5040, N5038, N226);
and AND2 (N5041, N5040, N4930);
nor NOR4 (N5042, N5041, N5034, N3817, N2850);
or OR4 (N5043, N333, N3665, N4404, N2711);
buf BUF1 (N5044, N5042);
xor XOR2 (N5045, N5001, N2710);
buf BUF1 (N5046, N5045);
nand NAND4 (N5047, N5014, N4334, N2004, N4028);
buf BUF1 (N5048, N5035);
or OR3 (N5049, N5022, N182, N4120);
xor XOR2 (N5050, N5023, N666);
and AND4 (N5051, N5036, N3452, N1971, N3441);
not NOT1 (N5052, N5047);
nor NOR4 (N5053, N5049, N3402, N2697, N3523);
not NOT1 (N5054, N5051);
xor XOR2 (N5055, N5050, N1999);
nand NAND2 (N5056, N5043, N4620);
nand NAND3 (N5057, N5039, N1625, N49);
and AND4 (N5058, N5056, N4416, N457, N3021);
and AND3 (N5059, N5053, N198, N6);
nand NAND2 (N5060, N5055, N46);
nand NAND3 (N5061, N5052, N2682, N2819);
nand NAND2 (N5062, N5060, N2318);
and AND2 (N5063, N5046, N4375);
buf BUF1 (N5064, N5063);
or OR3 (N5065, N5057, N464, N3796);
or OR3 (N5066, N5062, N3095, N4205);
buf BUF1 (N5067, N5054);
buf BUF1 (N5068, N5067);
and AND3 (N5069, N5058, N3442, N3769);
and AND4 (N5070, N5066, N2934, N1018, N3962);
not NOT1 (N5071, N5061);
nand NAND3 (N5072, N5071, N1249, N1804);
nor NOR3 (N5073, N5072, N5037, N115);
buf BUF1 (N5074, N1355);
xor XOR2 (N5075, N5059, N1120);
and AND2 (N5076, N5068, N4066);
nand NAND2 (N5077, N5065, N771);
not NOT1 (N5078, N5076);
and AND3 (N5079, N5048, N2267, N1122);
not NOT1 (N5080, N5073);
not NOT1 (N5081, N5064);
buf BUF1 (N5082, N5080);
buf BUF1 (N5083, N5070);
not NOT1 (N5084, N5044);
not NOT1 (N5085, N5069);
and AND3 (N5086, N5081, N1261, N3978);
nand NAND3 (N5087, N5083, N169, N2958);
nor NOR3 (N5088, N5079, N1360, N2342);
nand NAND3 (N5089, N5074, N3949, N4241);
nor NOR2 (N5090, N5089, N4507);
and AND2 (N5091, N5084, N1651);
nand NAND2 (N5092, N5090, N1455);
buf BUF1 (N5093, N5092);
xor XOR2 (N5094, N5091, N2752);
nand NAND3 (N5095, N5082, N1079, N2347);
not NOT1 (N5096, N5075);
nand NAND4 (N5097, N5078, N2896, N3959, N773);
nand NAND3 (N5098, N5094, N831, N1375);
xor XOR2 (N5099, N5097, N4747);
nor NOR3 (N5100, N5095, N2345, N2878);
or OR2 (N5101, N5093, N31);
buf BUF1 (N5102, N5077);
xor XOR2 (N5103, N5096, N1862);
and AND3 (N5104, N5099, N1935, N2462);
nor NOR2 (N5105, N5088, N2519);
or OR4 (N5106, N5102, N1738, N4067, N4200);
xor XOR2 (N5107, N5087, N1246);
buf BUF1 (N5108, N5106);
not NOT1 (N5109, N5103);
nor NOR4 (N5110, N5086, N3729, N4429, N1573);
or OR2 (N5111, N5110, N3816);
and AND2 (N5112, N5085, N3777);
nor NOR4 (N5113, N5111, N3145, N4305, N4133);
xor XOR2 (N5114, N5098, N3028);
and AND3 (N5115, N5112, N1536, N4549);
xor XOR2 (N5116, N5101, N4503);
nor NOR3 (N5117, N5108, N4712, N2221);
buf BUF1 (N5118, N5114);
and AND3 (N5119, N5116, N91, N397);
nor NOR4 (N5120, N5117, N2218, N2448, N3910);
buf BUF1 (N5121, N5109);
nand NAND2 (N5122, N5120, N3654);
xor XOR2 (N5123, N5118, N118);
buf BUF1 (N5124, N5121);
xor XOR2 (N5125, N5104, N3283);
or OR2 (N5126, N5125, N3800);
xor XOR2 (N5127, N5126, N2929);
not NOT1 (N5128, N5107);
not NOT1 (N5129, N5122);
not NOT1 (N5130, N5119);
nor NOR2 (N5131, N5130, N531);
and AND3 (N5132, N5105, N4794, N4741);
or OR3 (N5133, N5131, N2472, N3785);
and AND4 (N5134, N5129, N2645, N1290, N2358);
buf BUF1 (N5135, N5100);
nand NAND2 (N5136, N5115, N4096);
buf BUF1 (N5137, N5136);
nor NOR4 (N5138, N5132, N4110, N2098, N3729);
nand NAND4 (N5139, N5127, N1114, N3894, N4906);
nor NOR2 (N5140, N5135, N2160);
and AND3 (N5141, N5133, N4016, N1140);
or OR4 (N5142, N5139, N2196, N220, N4623);
buf BUF1 (N5143, N5141);
nor NOR4 (N5144, N5140, N2633, N1748, N3615);
xor XOR2 (N5145, N5143, N3587);
xor XOR2 (N5146, N5145, N3753);
or OR3 (N5147, N5124, N862, N1999);
not NOT1 (N5148, N5142);
buf BUF1 (N5149, N5137);
nand NAND4 (N5150, N5147, N1968, N3425, N1068);
nand NAND2 (N5151, N5144, N3254);
or OR2 (N5152, N5150, N3891);
nand NAND3 (N5153, N5134, N2091, N1410);
nand NAND4 (N5154, N5128, N646, N3069, N689);
nand NAND3 (N5155, N5146, N1935, N4954);
or OR4 (N5156, N5123, N4421, N4990, N2728);
buf BUF1 (N5157, N5154);
and AND3 (N5158, N5148, N3032, N5021);
and AND3 (N5159, N5157, N531, N629);
xor XOR2 (N5160, N5159, N4730);
xor XOR2 (N5161, N5149, N2338);
not NOT1 (N5162, N5155);
not NOT1 (N5163, N5162);
xor XOR2 (N5164, N5153, N4147);
buf BUF1 (N5165, N5164);
buf BUF1 (N5166, N5163);
not NOT1 (N5167, N5165);
nor NOR4 (N5168, N5160, N495, N3674, N5058);
nor NOR4 (N5169, N5138, N4035, N1606, N3598);
or OR2 (N5170, N5161, N1958);
or OR2 (N5171, N5158, N2324);
not NOT1 (N5172, N5113);
not NOT1 (N5173, N5151);
not NOT1 (N5174, N5173);
nand NAND3 (N5175, N5170, N3733, N4907);
nand NAND2 (N5176, N5167, N875);
buf BUF1 (N5177, N5152);
xor XOR2 (N5178, N5156, N1731);
nand NAND4 (N5179, N5176, N1711, N4964, N1444);
xor XOR2 (N5180, N5174, N3227);
or OR4 (N5181, N5166, N2450, N1487, N4912);
nor NOR3 (N5182, N5180, N5168, N695);
nor NOR3 (N5183, N658, N849, N3110);
buf BUF1 (N5184, N5181);
nor NOR4 (N5185, N5178, N2754, N2459, N4713);
and AND3 (N5186, N5179, N3239, N4201);
and AND3 (N5187, N5169, N2955, N2667);
not NOT1 (N5188, N5175);
xor XOR2 (N5189, N5186, N2313);
nand NAND3 (N5190, N5184, N2383, N1967);
not NOT1 (N5191, N5185);
buf BUF1 (N5192, N5171);
not NOT1 (N5193, N5190);
xor XOR2 (N5194, N5182, N2696);
not NOT1 (N5195, N5191);
nor NOR2 (N5196, N5192, N454);
nand NAND3 (N5197, N5196, N3512, N2382);
xor XOR2 (N5198, N5177, N4367);
and AND3 (N5199, N5198, N639, N4627);
nor NOR2 (N5200, N5187, N2893);
not NOT1 (N5201, N5189);
buf BUF1 (N5202, N5183);
or OR4 (N5203, N5188, N3444, N1621, N4420);
nor NOR3 (N5204, N5172, N3083, N1448);
and AND4 (N5205, N5201, N4098, N2145, N2351);
xor XOR2 (N5206, N5204, N2291);
or OR3 (N5207, N5199, N3810, N228);
buf BUF1 (N5208, N5194);
and AND3 (N5209, N5193, N4192, N3109);
xor XOR2 (N5210, N5205, N1870);
not NOT1 (N5211, N5200);
nor NOR2 (N5212, N5207, N1167);
not NOT1 (N5213, N5197);
or OR4 (N5214, N5210, N2558, N387, N2913);
buf BUF1 (N5215, N5212);
not NOT1 (N5216, N5206);
and AND2 (N5217, N5208, N884);
or OR2 (N5218, N5195, N870);
not NOT1 (N5219, N5216);
or OR4 (N5220, N5219, N3763, N1070, N1932);
nand NAND3 (N5221, N5213, N4031, N4257);
nor NOR3 (N5222, N5209, N626, N1547);
buf BUF1 (N5223, N5214);
and AND3 (N5224, N5220, N257, N2176);
buf BUF1 (N5225, N5217);
nand NAND3 (N5226, N5223, N3653, N3015);
and AND2 (N5227, N5203, N3569);
and AND3 (N5228, N5218, N1096, N3550);
nand NAND4 (N5229, N5226, N2351, N4447, N930);
nand NAND3 (N5230, N5224, N3662, N4009);
nand NAND2 (N5231, N5215, N1575);
xor XOR2 (N5232, N5229, N771);
buf BUF1 (N5233, N5228);
not NOT1 (N5234, N5221);
nand NAND3 (N5235, N5234, N3411, N2708);
nand NAND2 (N5236, N5233, N4619);
nand NAND4 (N5237, N5211, N2960, N2595, N3639);
buf BUF1 (N5238, N5237);
nand NAND2 (N5239, N5227, N97);
nor NOR2 (N5240, N5231, N4576);
xor XOR2 (N5241, N5238, N1325);
buf BUF1 (N5242, N5202);
and AND3 (N5243, N5240, N3390, N4441);
nand NAND4 (N5244, N5243, N1692, N2985, N566);
or OR3 (N5245, N5241, N3014, N748);
and AND4 (N5246, N5232, N1631, N2741, N4786);
and AND3 (N5247, N5245, N3106, N4363);
or OR3 (N5248, N5236, N3631, N3793);
nor NOR4 (N5249, N5248, N2406, N259, N4230);
nor NOR2 (N5250, N5225, N3004);
and AND4 (N5251, N5247, N4734, N4985, N1302);
nand NAND3 (N5252, N5235, N4469, N4568);
not NOT1 (N5253, N5250);
and AND4 (N5254, N5230, N4047, N1760, N577);
or OR2 (N5255, N5244, N446);
nand NAND4 (N5256, N5239, N3809, N4282, N4350);
or OR2 (N5257, N5251, N1323);
xor XOR2 (N5258, N5252, N2410);
nand NAND4 (N5259, N5256, N49, N2743, N4116);
and AND4 (N5260, N5258, N2525, N667, N3260);
xor XOR2 (N5261, N5254, N5213);
not NOT1 (N5262, N5253);
not NOT1 (N5263, N5246);
and AND3 (N5264, N5260, N2528, N3846);
or OR3 (N5265, N5222, N1180, N153);
xor XOR2 (N5266, N5259, N2684);
and AND2 (N5267, N5264, N5067);
xor XOR2 (N5268, N5249, N2635);
nand NAND2 (N5269, N5262, N4028);
and AND4 (N5270, N5242, N3126, N4818, N2545);
nor NOR4 (N5271, N5267, N1550, N3500, N2298);
nand NAND4 (N5272, N5263, N690, N2618, N1605);
nand NAND3 (N5273, N5271, N1339, N2338);
and AND2 (N5274, N5266, N3318);
nor NOR2 (N5275, N5268, N4999);
nand NAND2 (N5276, N5261, N3556);
nand NAND4 (N5277, N5257, N2143, N4415, N3618);
not NOT1 (N5278, N5270);
nand NAND4 (N5279, N5277, N3717, N4778, N864);
buf BUF1 (N5280, N5278);
and AND2 (N5281, N5269, N4827);
buf BUF1 (N5282, N5255);
nor NOR2 (N5283, N5265, N4393);
or OR3 (N5284, N5275, N2292, N173);
xor XOR2 (N5285, N5272, N1988);
buf BUF1 (N5286, N5283);
nor NOR2 (N5287, N5281, N5216);
nand NAND4 (N5288, N5284, N2266, N1293, N1692);
xor XOR2 (N5289, N5287, N3081);
nor NOR3 (N5290, N5280, N4851, N453);
nand NAND3 (N5291, N5276, N5277, N4097);
xor XOR2 (N5292, N5290, N4851);
or OR4 (N5293, N5282, N556, N384, N3917);
not NOT1 (N5294, N5273);
buf BUF1 (N5295, N5289);
buf BUF1 (N5296, N5286);
nor NOR2 (N5297, N5288, N5232);
buf BUF1 (N5298, N5274);
or OR2 (N5299, N5297, N5115);
nand NAND4 (N5300, N5285, N4756, N479, N4551);
or OR2 (N5301, N5293, N164);
not NOT1 (N5302, N5295);
nand NAND4 (N5303, N5299, N3971, N1525, N3895);
buf BUF1 (N5304, N5303);
not NOT1 (N5305, N5304);
nand NAND2 (N5306, N5296, N2600);
buf BUF1 (N5307, N5306);
buf BUF1 (N5308, N5301);
and AND4 (N5309, N5307, N2087, N4663, N3501);
buf BUF1 (N5310, N5292);
buf BUF1 (N5311, N5300);
or OR3 (N5312, N5309, N1394, N3318);
not NOT1 (N5313, N5308);
or OR4 (N5314, N5312, N2023, N3918, N321);
buf BUF1 (N5315, N5294);
nor NOR2 (N5316, N5305, N3808);
nand NAND4 (N5317, N5310, N3699, N3096, N603);
not NOT1 (N5318, N5311);
nor NOR4 (N5319, N5313, N1473, N1781, N962);
not NOT1 (N5320, N5314);
xor XOR2 (N5321, N5319, N2083);
and AND2 (N5322, N5298, N4546);
buf BUF1 (N5323, N5322);
or OR2 (N5324, N5321, N3393);
and AND3 (N5325, N5291, N4241, N3323);
buf BUF1 (N5326, N5316);
or OR2 (N5327, N5317, N713);
and AND3 (N5328, N5302, N1476, N3283);
not NOT1 (N5329, N5318);
nor NOR4 (N5330, N5315, N799, N4843, N1217);
buf BUF1 (N5331, N5330);
xor XOR2 (N5332, N5320, N1872);
xor XOR2 (N5333, N5327, N3470);
and AND3 (N5334, N5329, N1812, N3399);
nor NOR2 (N5335, N5326, N3661);
not NOT1 (N5336, N5324);
nand NAND3 (N5337, N5336, N4290, N3841);
not NOT1 (N5338, N5335);
and AND2 (N5339, N5325, N1644);
and AND4 (N5340, N5331, N3997, N3052, N1770);
and AND2 (N5341, N5328, N5209);
or OR4 (N5342, N5334, N1240, N4489, N4619);
buf BUF1 (N5343, N5323);
buf BUF1 (N5344, N5332);
buf BUF1 (N5345, N5343);
and AND3 (N5346, N5333, N4892, N1516);
buf BUF1 (N5347, N5279);
xor XOR2 (N5348, N5345, N4117);
not NOT1 (N5349, N5339);
and AND3 (N5350, N5338, N5035, N2763);
and AND4 (N5351, N5342, N5088, N872, N5031);
nand NAND2 (N5352, N5350, N1702);
and AND4 (N5353, N5346, N2766, N5146, N3484);
and AND3 (N5354, N5353, N3442, N2241);
or OR3 (N5355, N5340, N390, N2421);
nor NOR3 (N5356, N5352, N4696, N5314);
and AND3 (N5357, N5341, N4297, N2626);
buf BUF1 (N5358, N5348);
or OR3 (N5359, N5337, N1666, N5198);
nor NOR3 (N5360, N5354, N1262, N297);
nor NOR2 (N5361, N5360, N2312);
nor NOR2 (N5362, N5358, N4381);
and AND4 (N5363, N5359, N3506, N4959, N2865);
not NOT1 (N5364, N5356);
xor XOR2 (N5365, N5362, N3324);
or OR2 (N5366, N5349, N2783);
nand NAND3 (N5367, N5344, N3465, N1288);
or OR3 (N5368, N5351, N5262, N4638);
and AND3 (N5369, N5363, N892, N4118);
buf BUF1 (N5370, N5355);
xor XOR2 (N5371, N5365, N4866);
nand NAND3 (N5372, N5366, N3747, N4356);
buf BUF1 (N5373, N5357);
and AND4 (N5374, N5347, N155, N231, N2132);
nor NOR4 (N5375, N5371, N3469, N111, N3268);
and AND4 (N5376, N5364, N3227, N2837, N119);
not NOT1 (N5377, N5369);
buf BUF1 (N5378, N5367);
not NOT1 (N5379, N5374);
and AND2 (N5380, N5361, N3682);
nor NOR3 (N5381, N5375, N3133, N2614);
not NOT1 (N5382, N5372);
or OR2 (N5383, N5368, N3493);
or OR4 (N5384, N5382, N2923, N3969, N2143);
nor NOR2 (N5385, N5373, N31);
buf BUF1 (N5386, N5379);
not NOT1 (N5387, N5376);
or OR3 (N5388, N5377, N1372, N4187);
buf BUF1 (N5389, N5380);
nand NAND2 (N5390, N5384, N2837);
xor XOR2 (N5391, N5385, N1755);
buf BUF1 (N5392, N5381);
or OR3 (N5393, N5383, N2651, N3815);
buf BUF1 (N5394, N5393);
nor NOR3 (N5395, N5391, N2884, N2254);
xor XOR2 (N5396, N5388, N4026);
xor XOR2 (N5397, N5394, N446);
not NOT1 (N5398, N5378);
or OR3 (N5399, N5397, N342, N4785);
nor NOR4 (N5400, N5390, N456, N2270, N1025);
nand NAND3 (N5401, N5399, N4532, N1608);
xor XOR2 (N5402, N5398, N5184);
nor NOR3 (N5403, N5401, N546, N4986);
xor XOR2 (N5404, N5389, N2337);
and AND3 (N5405, N5386, N4612, N2539);
nor NOR4 (N5406, N5404, N4441, N1669, N3925);
not NOT1 (N5407, N5387);
buf BUF1 (N5408, N5405);
xor XOR2 (N5409, N5370, N533);
not NOT1 (N5410, N5400);
not NOT1 (N5411, N5408);
buf BUF1 (N5412, N5392);
buf BUF1 (N5413, N5406);
nor NOR4 (N5414, N5413, N2419, N1068, N4434);
or OR4 (N5415, N5407, N2986, N5009, N2737);
and AND2 (N5416, N5411, N995);
buf BUF1 (N5417, N5410);
xor XOR2 (N5418, N5396, N2758);
buf BUF1 (N5419, N5395);
xor XOR2 (N5420, N5403, N5356);
nor NOR3 (N5421, N5409, N3541, N2511);
or OR4 (N5422, N5420, N5188, N2403, N3849);
buf BUF1 (N5423, N5417);
buf BUF1 (N5424, N5423);
not NOT1 (N5425, N5422);
buf BUF1 (N5426, N5421);
and AND2 (N5427, N5419, N204);
and AND3 (N5428, N5414, N1863, N5354);
not NOT1 (N5429, N5425);
not NOT1 (N5430, N5416);
not NOT1 (N5431, N5426);
nand NAND2 (N5432, N5424, N4965);
not NOT1 (N5433, N5415);
nor NOR4 (N5434, N5432, N3969, N2020, N4522);
buf BUF1 (N5435, N5412);
buf BUF1 (N5436, N5434);
or OR2 (N5437, N5427, N505);
not NOT1 (N5438, N5418);
nand NAND4 (N5439, N5437, N368, N3255, N26);
nand NAND3 (N5440, N5436, N1556, N2274);
nor NOR3 (N5441, N5430, N2915, N11);
nand NAND3 (N5442, N5438, N1066, N667);
nand NAND4 (N5443, N5442, N1113, N867, N5337);
not NOT1 (N5444, N5429);
nand NAND4 (N5445, N5402, N4194, N4016, N2734);
buf BUF1 (N5446, N5441);
xor XOR2 (N5447, N5428, N2248);
not NOT1 (N5448, N5446);
not NOT1 (N5449, N5448);
nand NAND4 (N5450, N5433, N887, N3116, N1297);
buf BUF1 (N5451, N5445);
not NOT1 (N5452, N5450);
and AND3 (N5453, N5447, N4191, N4675);
or OR3 (N5454, N5451, N477, N1183);
xor XOR2 (N5455, N5431, N327);
buf BUF1 (N5456, N5435);
nand NAND3 (N5457, N5455, N47, N747);
not NOT1 (N5458, N5449);
and AND4 (N5459, N5444, N1579, N3896, N2986);
nor NOR4 (N5460, N5458, N4879, N4457, N4999);
and AND4 (N5461, N5453, N2377, N1806, N4742);
xor XOR2 (N5462, N5454, N3351);
or OR4 (N5463, N5460, N4187, N4896, N3895);
nand NAND3 (N5464, N5443, N3250, N3853);
nand NAND2 (N5465, N5439, N3563);
not NOT1 (N5466, N5440);
nor NOR4 (N5467, N5456, N3781, N4886, N2317);
or OR4 (N5468, N5459, N1862, N2113, N323);
and AND2 (N5469, N5466, N5225);
nand NAND3 (N5470, N5462, N2743, N392);
nor NOR2 (N5471, N5468, N1977);
xor XOR2 (N5472, N5469, N4383);
nor NOR4 (N5473, N5464, N4814, N2185, N97);
nand NAND2 (N5474, N5471, N1132);
nand NAND4 (N5475, N5474, N3174, N3165, N1693);
buf BUF1 (N5476, N5472);
buf BUF1 (N5477, N5476);
not NOT1 (N5478, N5465);
nor NOR4 (N5479, N5463, N1623, N781, N3772);
xor XOR2 (N5480, N5457, N4717);
xor XOR2 (N5481, N5480, N1852);
buf BUF1 (N5482, N5473);
or OR2 (N5483, N5467, N5253);
nand NAND2 (N5484, N5470, N416);
and AND3 (N5485, N5475, N2196, N3403);
not NOT1 (N5486, N5452);
nand NAND2 (N5487, N5486, N3233);
xor XOR2 (N5488, N5485, N1544);
nand NAND4 (N5489, N5482, N1302, N220, N1454);
and AND4 (N5490, N5461, N3734, N1687, N2372);
and AND3 (N5491, N5483, N3599, N2832);
or OR2 (N5492, N5481, N4300);
or OR3 (N5493, N5487, N5393, N3909);
nand NAND3 (N5494, N5478, N4849, N1969);
nor NOR4 (N5495, N5492, N1633, N5211, N5387);
buf BUF1 (N5496, N5495);
or OR3 (N5497, N5489, N5351, N2548);
buf BUF1 (N5498, N5494);
buf BUF1 (N5499, N5496);
nand NAND4 (N5500, N5497, N2563, N900, N2466);
nand NAND4 (N5501, N5500, N4687, N5212, N3948);
xor XOR2 (N5502, N5490, N3624);
buf BUF1 (N5503, N5477);
buf BUF1 (N5504, N5493);
buf BUF1 (N5505, N5491);
and AND4 (N5506, N5503, N4888, N861, N5211);
or OR2 (N5507, N5501, N473);
and AND3 (N5508, N5498, N576, N4539);
nand NAND4 (N5509, N5506, N2996, N4852, N2004);
nand NAND4 (N5510, N5484, N5003, N657, N4693);
and AND2 (N5511, N5502, N4367);
and AND4 (N5512, N5510, N3013, N5311, N98);
not NOT1 (N5513, N5505);
and AND3 (N5514, N5479, N4289, N3277);
xor XOR2 (N5515, N5512, N5291);
xor XOR2 (N5516, N5504, N1314);
nor NOR3 (N5517, N5508, N5241, N3347);
nand NAND3 (N5518, N5509, N2789, N2198);
or OR3 (N5519, N5514, N377, N4776);
xor XOR2 (N5520, N5519, N2596);
nand NAND4 (N5521, N5513, N2717, N4958, N3239);
buf BUF1 (N5522, N5499);
not NOT1 (N5523, N5521);
not NOT1 (N5524, N5520);
nand NAND2 (N5525, N5524, N116);
and AND2 (N5526, N5525, N1562);
buf BUF1 (N5527, N5507);
nor NOR3 (N5528, N5517, N4971, N4638);
buf BUF1 (N5529, N5527);
nand NAND4 (N5530, N5518, N738, N2348, N4931);
nor NOR2 (N5531, N5511, N4342);
buf BUF1 (N5532, N5526);
buf BUF1 (N5533, N5530);
xor XOR2 (N5534, N5488, N3029);
xor XOR2 (N5535, N5532, N2179);
buf BUF1 (N5536, N5515);
or OR3 (N5537, N5531, N1509, N1805);
or OR4 (N5538, N5523, N1120, N3066, N1366);
or OR2 (N5539, N5538, N1479);
and AND2 (N5540, N5537, N1027);
buf BUF1 (N5541, N5534);
buf BUF1 (N5542, N5529);
not NOT1 (N5543, N5541);
or OR3 (N5544, N5535, N4183, N756);
buf BUF1 (N5545, N5516);
nor NOR2 (N5546, N5522, N1643);
xor XOR2 (N5547, N5543, N3927);
nor NOR3 (N5548, N5528, N4934, N937);
and AND3 (N5549, N5536, N2937, N2679);
buf BUF1 (N5550, N5544);
and AND2 (N5551, N5539, N4631);
xor XOR2 (N5552, N5551, N2668);
or OR4 (N5553, N5546, N845, N4365, N5477);
nor NOR2 (N5554, N5552, N5002);
or OR3 (N5555, N5548, N2451, N368);
nor NOR2 (N5556, N5549, N2846);
not NOT1 (N5557, N5545);
not NOT1 (N5558, N5533);
xor XOR2 (N5559, N5558, N5260);
nand NAND2 (N5560, N5556, N49);
xor XOR2 (N5561, N5542, N2495);
xor XOR2 (N5562, N5560, N469);
or OR2 (N5563, N5562, N4928);
buf BUF1 (N5564, N5540);
xor XOR2 (N5565, N5553, N4335);
buf BUF1 (N5566, N5554);
nor NOR3 (N5567, N5547, N4660, N4638);
nand NAND3 (N5568, N5550, N466, N3775);
nand NAND4 (N5569, N5567, N2638, N531, N1847);
and AND2 (N5570, N5564, N469);
xor XOR2 (N5571, N5561, N303);
nor NOR4 (N5572, N5571, N2121, N2467, N738);
buf BUF1 (N5573, N5559);
and AND4 (N5574, N5570, N1906, N1814, N3158);
buf BUF1 (N5575, N5557);
nor NOR4 (N5576, N5569, N1494, N4388, N2654);
nand NAND4 (N5577, N5566, N491, N3774, N458);
buf BUF1 (N5578, N5577);
nor NOR3 (N5579, N5555, N3014, N2154);
nand NAND4 (N5580, N5565, N5528, N4825, N4946);
nand NAND3 (N5581, N5580, N2306, N4511);
xor XOR2 (N5582, N5575, N4530);
buf BUF1 (N5583, N5568);
and AND4 (N5584, N5581, N4370, N2407, N3257);
or OR2 (N5585, N5583, N79);
or OR4 (N5586, N5584, N4276, N1841, N1244);
nand NAND3 (N5587, N5574, N4891, N4236);
or OR2 (N5588, N5586, N3331);
not NOT1 (N5589, N5578);
or OR4 (N5590, N5587, N2476, N396, N51);
nand NAND2 (N5591, N5590, N1728);
xor XOR2 (N5592, N5591, N307);
and AND3 (N5593, N5573, N5223, N2531);
not NOT1 (N5594, N5576);
xor XOR2 (N5595, N5572, N170);
nor NOR4 (N5596, N5582, N2178, N3080, N1597);
nor NOR4 (N5597, N5579, N2627, N2309, N1711);
xor XOR2 (N5598, N5595, N3715);
or OR2 (N5599, N5598, N3940);
or OR2 (N5600, N5599, N2215);
or OR2 (N5601, N5563, N588);
buf BUF1 (N5602, N5588);
and AND2 (N5603, N5596, N2886);
or OR2 (N5604, N5585, N1166);
and AND3 (N5605, N5597, N2068, N1284);
and AND3 (N5606, N5602, N5234, N1920);
and AND3 (N5607, N5594, N4979, N2153);
nand NAND2 (N5608, N5606, N2149);
buf BUF1 (N5609, N5592);
not NOT1 (N5610, N5600);
or OR2 (N5611, N5605, N4074);
xor XOR2 (N5612, N5610, N4500);
xor XOR2 (N5613, N5609, N1292);
nor NOR3 (N5614, N5604, N1745, N2750);
or OR3 (N5615, N5614, N3308, N856);
xor XOR2 (N5616, N5593, N2534);
nand NAND4 (N5617, N5603, N2354, N1731, N400);
nand NAND2 (N5618, N5612, N4059);
and AND2 (N5619, N5608, N2280);
not NOT1 (N5620, N5601);
xor XOR2 (N5621, N5613, N3115);
and AND4 (N5622, N5616, N3092, N4927, N2146);
xor XOR2 (N5623, N5620, N476);
nor NOR3 (N5624, N5621, N2050, N3019);
and AND4 (N5625, N5622, N2761, N2597, N4321);
nor NOR2 (N5626, N5611, N3837);
or OR2 (N5627, N5619, N4420);
and AND2 (N5628, N5624, N2510);
nand NAND3 (N5629, N5617, N1437, N1972);
not NOT1 (N5630, N5625);
nor NOR2 (N5631, N5589, N1291);
nor NOR2 (N5632, N5618, N2524);
xor XOR2 (N5633, N5628, N2474);
and AND4 (N5634, N5631, N4868, N1030, N1329);
nor NOR2 (N5635, N5627, N5508);
or OR2 (N5636, N5634, N1649);
nand NAND2 (N5637, N5635, N4712);
xor XOR2 (N5638, N5637, N58);
nor NOR3 (N5639, N5623, N1243, N1066);
buf BUF1 (N5640, N5607);
and AND2 (N5641, N5640, N847);
buf BUF1 (N5642, N5630);
and AND2 (N5643, N5642, N238);
and AND3 (N5644, N5632, N1670, N3608);
nor NOR3 (N5645, N5641, N3651, N2423);
xor XOR2 (N5646, N5633, N2905);
not NOT1 (N5647, N5629);
or OR4 (N5648, N5643, N666, N2974, N3610);
buf BUF1 (N5649, N5639);
or OR3 (N5650, N5645, N2336, N857);
nand NAND2 (N5651, N5647, N5516);
nor NOR4 (N5652, N5638, N3263, N2564, N2535);
nor NOR2 (N5653, N5648, N5480);
nand NAND3 (N5654, N5644, N2821, N133);
buf BUF1 (N5655, N5652);
not NOT1 (N5656, N5646);
nor NOR2 (N5657, N5650, N399);
not NOT1 (N5658, N5626);
buf BUF1 (N5659, N5657);
not NOT1 (N5660, N5656);
or OR2 (N5661, N5654, N3636);
xor XOR2 (N5662, N5651, N644);
and AND3 (N5663, N5649, N1651, N3090);
buf BUF1 (N5664, N5659);
xor XOR2 (N5665, N5663, N4384);
buf BUF1 (N5666, N5660);
not NOT1 (N5667, N5658);
and AND4 (N5668, N5653, N1171, N660, N2886);
nor NOR4 (N5669, N5667, N4799, N593, N1935);
or OR4 (N5670, N5666, N1273, N606, N5620);
nand NAND4 (N5671, N5669, N849, N2156, N3255);
nand NAND4 (N5672, N5668, N1834, N3664, N1035);
or OR2 (N5673, N5671, N4682);
xor XOR2 (N5674, N5670, N1512);
buf BUF1 (N5675, N5636);
buf BUF1 (N5676, N5675);
buf BUF1 (N5677, N5672);
and AND3 (N5678, N5665, N2312, N2449);
nand NAND3 (N5679, N5664, N1641, N2263);
or OR4 (N5680, N5662, N3283, N5053, N2743);
or OR2 (N5681, N5661, N4927);
nand NAND2 (N5682, N5674, N5378);
nor NOR4 (N5683, N5679, N4595, N2212, N5260);
xor XOR2 (N5684, N5680, N4418);
not NOT1 (N5685, N5678);
and AND3 (N5686, N5681, N5410, N3114);
not NOT1 (N5687, N5682);
nand NAND3 (N5688, N5673, N3305, N3103);
nand NAND4 (N5689, N5687, N3425, N5323, N3504);
not NOT1 (N5690, N5615);
buf BUF1 (N5691, N5690);
and AND4 (N5692, N5688, N3311, N4198, N1246);
nand NAND3 (N5693, N5676, N3895, N5174);
xor XOR2 (N5694, N5691, N1099);
or OR3 (N5695, N5684, N4516, N3091);
nand NAND3 (N5696, N5694, N514, N839);
xor XOR2 (N5697, N5683, N2836);
buf BUF1 (N5698, N5677);
not NOT1 (N5699, N5697);
xor XOR2 (N5700, N5689, N1901);
xor XOR2 (N5701, N5700, N2689);
not NOT1 (N5702, N5701);
xor XOR2 (N5703, N5693, N108);
nor NOR4 (N5704, N5698, N5342, N3708, N5369);
nand NAND2 (N5705, N5692, N1697);
or OR4 (N5706, N5703, N5268, N279, N598);
not NOT1 (N5707, N5655);
nor NOR4 (N5708, N5699, N2477, N4729, N3642);
or OR3 (N5709, N5696, N823, N4853);
or OR4 (N5710, N5707, N123, N5540, N3607);
nor NOR4 (N5711, N5686, N5652, N1305, N1534);
nor NOR3 (N5712, N5710, N2912, N1318);
not NOT1 (N5713, N5708);
nor NOR3 (N5714, N5711, N77, N883);
or OR3 (N5715, N5714, N2750, N1388);
buf BUF1 (N5716, N5685);
xor XOR2 (N5717, N5715, N4572);
nand NAND2 (N5718, N5704, N1733);
or OR3 (N5719, N5706, N798, N1524);
xor XOR2 (N5720, N5716, N2198);
or OR2 (N5721, N5719, N2169);
or OR3 (N5722, N5695, N817, N1643);
nor NOR4 (N5723, N5720, N1598, N1885, N3816);
not NOT1 (N5724, N5709);
or OR2 (N5725, N5705, N575);
not NOT1 (N5726, N5702);
or OR4 (N5727, N5725, N4003, N4236, N4803);
buf BUF1 (N5728, N5723);
and AND4 (N5729, N5721, N1817, N4658, N2897);
or OR3 (N5730, N5724, N803, N2436);
nand NAND4 (N5731, N5730, N4053, N4352, N5554);
or OR2 (N5732, N5717, N3259);
and AND4 (N5733, N5718, N4598, N1157, N1488);
and AND2 (N5734, N5733, N5209);
xor XOR2 (N5735, N5729, N5061);
and AND2 (N5736, N5728, N3009);
nand NAND4 (N5737, N5722, N5324, N1098, N4896);
buf BUF1 (N5738, N5732);
buf BUF1 (N5739, N5726);
buf BUF1 (N5740, N5734);
xor XOR2 (N5741, N5713, N3729);
nand NAND3 (N5742, N5741, N3206, N2610);
nand NAND2 (N5743, N5727, N5298);
nand NAND4 (N5744, N5736, N727, N1430, N4752);
not NOT1 (N5745, N5737);
xor XOR2 (N5746, N5739, N4793);
xor XOR2 (N5747, N5735, N3942);
not NOT1 (N5748, N5747);
buf BUF1 (N5749, N5746);
or OR2 (N5750, N5749, N3623);
nand NAND3 (N5751, N5745, N3423, N4420);
not NOT1 (N5752, N5731);
or OR2 (N5753, N5744, N2182);
and AND2 (N5754, N5753, N4474);
nor NOR4 (N5755, N5743, N3677, N2548, N2251);
buf BUF1 (N5756, N5755);
or OR3 (N5757, N5712, N1720, N2309);
not NOT1 (N5758, N5756);
or OR3 (N5759, N5751, N3419, N1001);
nor NOR3 (N5760, N5742, N2337, N5205);
nand NAND2 (N5761, N5760, N827);
not NOT1 (N5762, N5740);
xor XOR2 (N5763, N5759, N3477);
nor NOR3 (N5764, N5757, N3983, N2293);
nor NOR3 (N5765, N5750, N644, N5481);
xor XOR2 (N5766, N5748, N3928);
or OR2 (N5767, N5758, N1979);
or OR3 (N5768, N5762, N3649, N5459);
and AND3 (N5769, N5767, N2864, N5346);
and AND4 (N5770, N5738, N4346, N2175, N2015);
nor NOR2 (N5771, N5752, N84);
and AND4 (N5772, N5768, N1910, N2113, N4297);
nor NOR2 (N5773, N5770, N5384);
not NOT1 (N5774, N5765);
xor XOR2 (N5775, N5772, N4544);
and AND3 (N5776, N5769, N3834, N2360);
not NOT1 (N5777, N5771);
nand NAND3 (N5778, N5775, N2769, N2556);
not NOT1 (N5779, N5773);
nand NAND2 (N5780, N5776, N5514);
buf BUF1 (N5781, N5766);
not NOT1 (N5782, N5754);
nand NAND4 (N5783, N5774, N2291, N706, N3258);
not NOT1 (N5784, N5783);
nand NAND4 (N5785, N5777, N206, N1215, N237);
and AND4 (N5786, N5764, N891, N76, N1867);
xor XOR2 (N5787, N5778, N1795);
nor NOR2 (N5788, N5786, N5308);
buf BUF1 (N5789, N5779);
buf BUF1 (N5790, N5787);
not NOT1 (N5791, N5785);
nand NAND4 (N5792, N5761, N5638, N2344, N3004);
nor NOR4 (N5793, N5782, N1712, N274, N3888);
nor NOR3 (N5794, N5792, N5360, N4583);
buf BUF1 (N5795, N5790);
nor NOR2 (N5796, N5794, N3091);
or OR4 (N5797, N5791, N5431, N5281, N5406);
xor XOR2 (N5798, N5789, N3753);
buf BUF1 (N5799, N5781);
and AND4 (N5800, N5788, N2920, N2804, N1490);
or OR4 (N5801, N5797, N2096, N2291, N3158);
buf BUF1 (N5802, N5780);
nand NAND4 (N5803, N5802, N4609, N3319, N5178);
not NOT1 (N5804, N5799);
buf BUF1 (N5805, N5803);
not NOT1 (N5806, N5793);
nor NOR3 (N5807, N5800, N2347, N5417);
buf BUF1 (N5808, N5806);
nor NOR2 (N5809, N5808, N4853);
buf BUF1 (N5810, N5763);
and AND2 (N5811, N5795, N4348);
buf BUF1 (N5812, N5805);
not NOT1 (N5813, N5801);
xor XOR2 (N5814, N5809, N2384);
nand NAND4 (N5815, N5807, N3045, N4619, N2008);
xor XOR2 (N5816, N5815, N5058);
and AND2 (N5817, N5814, N3301);
not NOT1 (N5818, N5804);
not NOT1 (N5819, N5817);
buf BUF1 (N5820, N5811);
not NOT1 (N5821, N5819);
and AND4 (N5822, N5798, N1346, N3993, N3134);
nor NOR2 (N5823, N5784, N1442);
buf BUF1 (N5824, N5812);
buf BUF1 (N5825, N5796);
nor NOR4 (N5826, N5818, N2949, N4781, N3451);
xor XOR2 (N5827, N5826, N4502);
buf BUF1 (N5828, N5827);
nand NAND2 (N5829, N5820, N4177);
or OR2 (N5830, N5823, N2308);
buf BUF1 (N5831, N5813);
and AND4 (N5832, N5810, N4976, N1765, N4607);
and AND3 (N5833, N5816, N1102, N5368);
not NOT1 (N5834, N5828);
nor NOR2 (N5835, N5832, N4978);
not NOT1 (N5836, N5825);
not NOT1 (N5837, N5835);
xor XOR2 (N5838, N5829, N735);
nand NAND3 (N5839, N5834, N4447, N1748);
and AND3 (N5840, N5833, N4334, N5001);
xor XOR2 (N5841, N5836, N347);
buf BUF1 (N5842, N5839);
nor NOR3 (N5843, N5837, N1568, N3514);
or OR2 (N5844, N5831, N251);
and AND2 (N5845, N5844, N4037);
nand NAND2 (N5846, N5830, N2941);
not NOT1 (N5847, N5846);
or OR3 (N5848, N5845, N1609, N4832);
nor NOR3 (N5849, N5847, N377, N531);
or OR4 (N5850, N5821, N1209, N2857, N3823);
not NOT1 (N5851, N5849);
buf BUF1 (N5852, N5841);
nor NOR4 (N5853, N5848, N604, N3159, N3346);
buf BUF1 (N5854, N5851);
and AND4 (N5855, N5852, N2274, N5624, N150);
buf BUF1 (N5856, N5840);
nor NOR4 (N5857, N5850, N2598, N3272, N5056);
nor NOR2 (N5858, N5822, N1449);
not NOT1 (N5859, N5857);
and AND2 (N5860, N5838, N5688);
xor XOR2 (N5861, N5859, N2622);
nand NAND3 (N5862, N5854, N3818, N3429);
or OR2 (N5863, N5842, N4163);
not NOT1 (N5864, N5863);
and AND4 (N5865, N5858, N1882, N4295, N5724);
xor XOR2 (N5866, N5861, N4588);
or OR2 (N5867, N5843, N5533);
nand NAND3 (N5868, N5824, N5644, N3228);
nand NAND4 (N5869, N5864, N2854, N5254, N5707);
or OR3 (N5870, N5866, N2802, N1541);
not NOT1 (N5871, N5868);
and AND4 (N5872, N5855, N4773, N2963, N3555);
or OR3 (N5873, N5870, N4627, N3037);
nand NAND3 (N5874, N5860, N3859, N2898);
and AND3 (N5875, N5865, N5371, N2112);
or OR2 (N5876, N5874, N899);
xor XOR2 (N5877, N5856, N2587);
buf BUF1 (N5878, N5867);
buf BUF1 (N5879, N5871);
xor XOR2 (N5880, N5876, N1458);
not NOT1 (N5881, N5869);
buf BUF1 (N5882, N5877);
nand NAND2 (N5883, N5862, N1925);
nand NAND4 (N5884, N5880, N2277, N180, N5471);
not NOT1 (N5885, N5881);
nor NOR3 (N5886, N5873, N4760, N1298);
and AND4 (N5887, N5883, N1367, N3429, N5791);
buf BUF1 (N5888, N5884);
and AND4 (N5889, N5879, N4644, N49, N4439);
xor XOR2 (N5890, N5885, N4554);
xor XOR2 (N5891, N5888, N4888);
not NOT1 (N5892, N5889);
not NOT1 (N5893, N5882);
and AND3 (N5894, N5890, N166, N3670);
nand NAND4 (N5895, N5894, N546, N72, N5463);
xor XOR2 (N5896, N5878, N3947);
or OR2 (N5897, N5853, N1408);
or OR2 (N5898, N5872, N3207);
xor XOR2 (N5899, N5898, N1354);
nand NAND2 (N5900, N5897, N4086);
not NOT1 (N5901, N5899);
or OR2 (N5902, N5875, N3040);
not NOT1 (N5903, N5893);
and AND3 (N5904, N5896, N2770, N62);
or OR4 (N5905, N5891, N936, N1359, N4396);
and AND2 (N5906, N5895, N169);
or OR3 (N5907, N5903, N2685, N884);
and AND2 (N5908, N5892, N4215);
not NOT1 (N5909, N5907);
buf BUF1 (N5910, N5900);
buf BUF1 (N5911, N5906);
nor NOR3 (N5912, N5887, N5731, N4707);
or OR3 (N5913, N5909, N29, N3040);
not NOT1 (N5914, N5908);
or OR4 (N5915, N5886, N5444, N4879, N2326);
xor XOR2 (N5916, N5915, N3401);
xor XOR2 (N5917, N5901, N1945);
or OR3 (N5918, N5914, N893, N665);
nor NOR4 (N5919, N5917, N3259, N2721, N5500);
or OR3 (N5920, N5916, N4906, N2499);
nand NAND4 (N5921, N5913, N5748, N4589, N2127);
nor NOR4 (N5922, N5918, N465, N3794, N2382);
and AND4 (N5923, N5911, N2909, N5099, N317);
or OR4 (N5924, N5905, N4234, N298, N1172);
not NOT1 (N5925, N5923);
or OR4 (N5926, N5912, N4576, N5754, N4502);
nor NOR4 (N5927, N5924, N519, N4571, N2648);
buf BUF1 (N5928, N5904);
xor XOR2 (N5929, N5920, N4603);
buf BUF1 (N5930, N5921);
buf BUF1 (N5931, N5926);
and AND4 (N5932, N5930, N32, N1364, N1318);
nand NAND2 (N5933, N5928, N3708);
nor NOR2 (N5934, N5931, N5097);
nor NOR2 (N5935, N5933, N3558);
and AND3 (N5936, N5902, N5129, N1394);
and AND4 (N5937, N5936, N2726, N2827, N4407);
not NOT1 (N5938, N5925);
buf BUF1 (N5939, N5937);
not NOT1 (N5940, N5939);
and AND2 (N5941, N5910, N5510);
xor XOR2 (N5942, N5938, N299);
xor XOR2 (N5943, N5940, N158);
or OR2 (N5944, N5919, N3910);
buf BUF1 (N5945, N5944);
or OR3 (N5946, N5922, N2838, N3119);
and AND2 (N5947, N5942, N1814);
not NOT1 (N5948, N5932);
xor XOR2 (N5949, N5935, N4384);
or OR2 (N5950, N5947, N9);
and AND3 (N5951, N5927, N3785, N5836);
and AND3 (N5952, N5950, N1006, N1270);
xor XOR2 (N5953, N5934, N3363);
not NOT1 (N5954, N5945);
and AND2 (N5955, N5948, N241);
or OR3 (N5956, N5929, N755, N173);
nand NAND2 (N5957, N5943, N1871);
and AND2 (N5958, N5957, N2221);
xor XOR2 (N5959, N5952, N1643);
or OR4 (N5960, N5958, N4937, N2476, N1045);
nand NAND2 (N5961, N5953, N3987);
xor XOR2 (N5962, N5955, N5300);
nand NAND2 (N5963, N5960, N3020);
nor NOR4 (N5964, N5961, N1529, N387, N3141);
nor NOR2 (N5965, N5956, N3873);
or OR3 (N5966, N5963, N587, N2372);
nor NOR3 (N5967, N5949, N2693, N5426);
and AND4 (N5968, N5941, N5476, N3105, N711);
xor XOR2 (N5969, N5964, N4638);
xor XOR2 (N5970, N5966, N2354);
not NOT1 (N5971, N5968);
and AND2 (N5972, N5946, N969);
xor XOR2 (N5973, N5951, N3091);
or OR2 (N5974, N5971, N4220);
and AND2 (N5975, N5962, N971);
buf BUF1 (N5976, N5973);
or OR2 (N5977, N5969, N188);
nor NOR3 (N5978, N5970, N5822, N580);
xor XOR2 (N5979, N5978, N437);
nand NAND3 (N5980, N5972, N5518, N2917);
or OR2 (N5981, N5980, N5946);
xor XOR2 (N5982, N5979, N2188);
and AND4 (N5983, N5965, N5119, N2513, N5388);
not NOT1 (N5984, N5975);
buf BUF1 (N5985, N5967);
nor NOR2 (N5986, N5954, N4035);
buf BUF1 (N5987, N5974);
not NOT1 (N5988, N5976);
nand NAND2 (N5989, N5977, N1534);
nor NOR4 (N5990, N5986, N2703, N3176, N3132);
nand NAND3 (N5991, N5959, N544, N4563);
nor NOR4 (N5992, N5991, N1306, N3133, N3638);
nand NAND2 (N5993, N5990, N3484);
buf BUF1 (N5994, N5981);
and AND4 (N5995, N5992, N1232, N2723, N3897);
buf BUF1 (N5996, N5994);
buf BUF1 (N5997, N5989);
xor XOR2 (N5998, N5988, N5500);
or OR2 (N5999, N5998, N2503);
buf BUF1 (N6000, N5982);
nand NAND3 (N6001, N6000, N3830, N2965);
and AND2 (N6002, N6001, N5259);
xor XOR2 (N6003, N5987, N3251);
or OR4 (N6004, N5997, N273, N1040, N740);
or OR2 (N6005, N5995, N1047);
not NOT1 (N6006, N5983);
nand NAND4 (N6007, N6006, N4605, N3042, N431);
not NOT1 (N6008, N6002);
buf BUF1 (N6009, N6004);
xor XOR2 (N6010, N6009, N4662);
or OR3 (N6011, N5993, N1515, N3766);
not NOT1 (N6012, N5999);
buf BUF1 (N6013, N6007);
not NOT1 (N6014, N6003);
and AND3 (N6015, N6005, N1436, N2676);
nor NOR3 (N6016, N6010, N128, N5353);
and AND4 (N6017, N6015, N4276, N3683, N1280);
or OR4 (N6018, N6008, N1543, N445, N448);
nor NOR2 (N6019, N6011, N3590);
nand NAND3 (N6020, N6017, N136, N2922);
or OR2 (N6021, N5985, N5187);
buf BUF1 (N6022, N6013);
nand NAND2 (N6023, N6022, N2403);
buf BUF1 (N6024, N6023);
or OR2 (N6025, N6021, N1418);
nor NOR3 (N6026, N6019, N3948, N3291);
or OR2 (N6027, N6026, N1309);
xor XOR2 (N6028, N6020, N4359);
xor XOR2 (N6029, N6027, N2144);
and AND3 (N6030, N6016, N1513, N5516);
xor XOR2 (N6031, N6030, N1881);
not NOT1 (N6032, N6031);
and AND4 (N6033, N5984, N907, N2224, N2908);
buf BUF1 (N6034, N6025);
nor NOR3 (N6035, N6032, N925, N2803);
xor XOR2 (N6036, N6012, N5863);
or OR4 (N6037, N5996, N3992, N294, N2973);
nand NAND4 (N6038, N6035, N3811, N267, N5872);
xor XOR2 (N6039, N6018, N5903);
xor XOR2 (N6040, N6039, N623);
xor XOR2 (N6041, N6036, N4426);
not NOT1 (N6042, N6028);
xor XOR2 (N6043, N6024, N2137);
or OR3 (N6044, N6041, N1961, N17);
or OR4 (N6045, N6044, N3806, N63, N154);
xor XOR2 (N6046, N6037, N1200);
or OR2 (N6047, N6034, N1048);
or OR4 (N6048, N6047, N5477, N3705, N4848);
or OR2 (N6049, N6042, N2725);
buf BUF1 (N6050, N6038);
not NOT1 (N6051, N6014);
buf BUF1 (N6052, N6043);
nand NAND3 (N6053, N6051, N5079, N3516);
or OR3 (N6054, N6029, N3987, N864);
or OR3 (N6055, N6049, N2276, N279);
nor NOR3 (N6056, N6040, N4763, N931);
nor NOR4 (N6057, N6045, N2665, N5492, N5264);
nor NOR2 (N6058, N6052, N4694);
not NOT1 (N6059, N6048);
not NOT1 (N6060, N6059);
not NOT1 (N6061, N6033);
not NOT1 (N6062, N6054);
nand NAND4 (N6063, N6057, N2409, N3300, N948);
nor NOR4 (N6064, N6058, N5604, N595, N2669);
or OR4 (N6065, N6053, N5930, N1875, N2246);
or OR2 (N6066, N6056, N5913);
nand NAND3 (N6067, N6066, N4380, N1133);
nand NAND3 (N6068, N6060, N4893, N3186);
buf BUF1 (N6069, N6067);
and AND2 (N6070, N6063, N4907);
nor NOR2 (N6071, N6050, N3008);
not NOT1 (N6072, N6068);
and AND2 (N6073, N6071, N1298);
nand NAND4 (N6074, N6069, N521, N1893, N2280);
or OR3 (N6075, N6062, N3689, N2114);
xor XOR2 (N6076, N6055, N2577);
nor NOR4 (N6077, N6073, N3063, N2983, N1448);
xor XOR2 (N6078, N6076, N1731);
nand NAND4 (N6079, N6074, N5899, N324, N3103);
and AND2 (N6080, N6070, N4053);
or OR4 (N6081, N6080, N3453, N1364, N1273);
or OR3 (N6082, N6065, N2196, N4113);
buf BUF1 (N6083, N6046);
and AND3 (N6084, N6061, N5176, N3227);
nor NOR2 (N6085, N6077, N4936);
buf BUF1 (N6086, N6078);
not NOT1 (N6087, N6079);
and AND2 (N6088, N6086, N580);
not NOT1 (N6089, N6064);
or OR2 (N6090, N6088, N3089);
nand NAND4 (N6091, N6075, N2436, N26, N1875);
not NOT1 (N6092, N6090);
and AND3 (N6093, N6087, N4617, N1814);
buf BUF1 (N6094, N6085);
buf BUF1 (N6095, N6091);
nand NAND2 (N6096, N6095, N2317);
nor NOR2 (N6097, N6094, N2144);
or OR3 (N6098, N6081, N1834, N1682);
xor XOR2 (N6099, N6096, N5862);
or OR3 (N6100, N6083, N2172, N3157);
and AND3 (N6101, N6097, N5700, N4708);
or OR4 (N6102, N6089, N2768, N4792, N5348);
and AND4 (N6103, N6072, N1852, N4571, N4547);
not NOT1 (N6104, N6093);
not NOT1 (N6105, N6100);
and AND2 (N6106, N6101, N191);
nand NAND2 (N6107, N6092, N3444);
not NOT1 (N6108, N6104);
nand NAND2 (N6109, N6102, N4534);
and AND2 (N6110, N6107, N1904);
xor XOR2 (N6111, N6084, N2333);
xor XOR2 (N6112, N6105, N4852);
xor XOR2 (N6113, N6106, N4262);
or OR3 (N6114, N6099, N5685, N4091);
not NOT1 (N6115, N6112);
or OR3 (N6116, N6103, N1345, N4485);
nand NAND2 (N6117, N6098, N5937);
xor XOR2 (N6118, N6117, N5534);
nand NAND4 (N6119, N6109, N4532, N5363, N874);
xor XOR2 (N6120, N6113, N1435);
nand NAND2 (N6121, N6108, N3526);
xor XOR2 (N6122, N6118, N5427);
not NOT1 (N6123, N6082);
and AND2 (N6124, N6120, N3133);
not NOT1 (N6125, N6121);
nor NOR3 (N6126, N6122, N4186, N844);
nor NOR4 (N6127, N6114, N4901, N3357, N4583);
nand NAND3 (N6128, N6127, N2683, N438);
or OR3 (N6129, N6123, N2084, N6015);
nand NAND4 (N6130, N6110, N5480, N3625, N727);
and AND2 (N6131, N6116, N2376);
and AND4 (N6132, N6130, N5869, N119, N2263);
nor NOR4 (N6133, N6124, N485, N4879, N934);
xor XOR2 (N6134, N6132, N847);
and AND3 (N6135, N6126, N5525, N1802);
not NOT1 (N6136, N6134);
not NOT1 (N6137, N6115);
nand NAND4 (N6138, N6119, N4688, N2928, N1911);
buf BUF1 (N6139, N6136);
xor XOR2 (N6140, N6131, N4131);
and AND3 (N6141, N6128, N1762, N103);
xor XOR2 (N6142, N6141, N2344);
or OR3 (N6143, N6137, N4055, N4333);
or OR2 (N6144, N6129, N5247);
nor NOR3 (N6145, N6140, N891, N1625);
buf BUF1 (N6146, N6111);
buf BUF1 (N6147, N6143);
or OR3 (N6148, N6144, N5412, N2319);
not NOT1 (N6149, N6135);
or OR2 (N6150, N6145, N1375);
and AND3 (N6151, N6148, N1040, N4222);
nand NAND4 (N6152, N6149, N2362, N3583, N5109);
buf BUF1 (N6153, N6139);
or OR2 (N6154, N6142, N2877);
nand NAND4 (N6155, N6150, N829, N5948, N4218);
xor XOR2 (N6156, N6146, N4017);
and AND4 (N6157, N6153, N995, N5438, N617);
nand NAND4 (N6158, N6138, N3360, N1882, N4207);
nand NAND3 (N6159, N6151, N4640, N364);
nor NOR4 (N6160, N6158, N5546, N2177, N974);
buf BUF1 (N6161, N6156);
and AND2 (N6162, N6154, N1725);
buf BUF1 (N6163, N6162);
xor XOR2 (N6164, N6155, N130);
nor NOR3 (N6165, N6147, N872, N4683);
buf BUF1 (N6166, N6164);
buf BUF1 (N6167, N6125);
xor XOR2 (N6168, N6167, N2087);
and AND2 (N6169, N6160, N4766);
buf BUF1 (N6170, N6165);
nor NOR2 (N6171, N6157, N3171);
buf BUF1 (N6172, N6166);
not NOT1 (N6173, N6163);
nand NAND4 (N6174, N6152, N2711, N5280, N660);
xor XOR2 (N6175, N6161, N3532);
not NOT1 (N6176, N6168);
xor XOR2 (N6177, N6170, N490);
xor XOR2 (N6178, N6174, N2156);
nor NOR2 (N6179, N6133, N5597);
not NOT1 (N6180, N6169);
and AND2 (N6181, N6178, N239);
or OR2 (N6182, N6179, N2506);
nand NAND2 (N6183, N6180, N515);
buf BUF1 (N6184, N6173);
not NOT1 (N6185, N6184);
xor XOR2 (N6186, N6175, N208);
xor XOR2 (N6187, N6186, N1292);
not NOT1 (N6188, N6177);
and AND4 (N6189, N6182, N3690, N1443, N3689);
nor NOR2 (N6190, N6171, N5979);
or OR2 (N6191, N6176, N5395);
nor NOR2 (N6192, N6181, N562);
nand NAND3 (N6193, N6183, N1525, N4647);
not NOT1 (N6194, N6190);
xor XOR2 (N6195, N6191, N5939);
and AND3 (N6196, N6172, N5329, N5248);
or OR4 (N6197, N6196, N3623, N2736, N3547);
and AND3 (N6198, N6195, N1300, N649);
xor XOR2 (N6199, N6198, N5839);
buf BUF1 (N6200, N6189);
xor XOR2 (N6201, N6192, N930);
and AND3 (N6202, N6197, N6062, N3317);
or OR4 (N6203, N6188, N2614, N5207, N1829);
nor NOR3 (N6204, N6159, N5234, N5366);
or OR3 (N6205, N6201, N4772, N1141);
buf BUF1 (N6206, N6204);
buf BUF1 (N6207, N6205);
nand NAND2 (N6208, N6206, N5594);
nand NAND4 (N6209, N6202, N875, N3908, N2281);
xor XOR2 (N6210, N6187, N2246);
xor XOR2 (N6211, N6208, N3342);
xor XOR2 (N6212, N6210, N4311);
nand NAND4 (N6213, N6199, N2540, N5640, N1151);
and AND2 (N6214, N6193, N3188);
and AND4 (N6215, N6200, N3734, N5694, N343);
xor XOR2 (N6216, N6207, N5070);
nor NOR2 (N6217, N6209, N2176);
not NOT1 (N6218, N6213);
buf BUF1 (N6219, N6218);
buf BUF1 (N6220, N6215);
or OR4 (N6221, N6203, N5069, N1258, N4278);
not NOT1 (N6222, N6214);
nand NAND3 (N6223, N6185, N2415, N5652);
nor NOR2 (N6224, N6211, N3172);
buf BUF1 (N6225, N6194);
nor NOR4 (N6226, N6225, N4986, N4687, N5164);
and AND4 (N6227, N6219, N2914, N5691, N92);
not NOT1 (N6228, N6212);
buf BUF1 (N6229, N6221);
not NOT1 (N6230, N6226);
nor NOR4 (N6231, N6229, N3560, N4821, N2882);
not NOT1 (N6232, N6224);
or OR3 (N6233, N6227, N6148, N4147);
not NOT1 (N6234, N6231);
or OR4 (N6235, N6223, N4431, N3894, N4403);
and AND4 (N6236, N6222, N248, N5769, N985);
buf BUF1 (N6237, N6234);
or OR3 (N6238, N6235, N2677, N1740);
xor XOR2 (N6239, N6236, N2841);
not NOT1 (N6240, N6237);
nand NAND2 (N6241, N6239, N2742);
xor XOR2 (N6242, N6230, N3488);
nand NAND4 (N6243, N6233, N4093, N1300, N2535);
xor XOR2 (N6244, N6217, N2720);
xor XOR2 (N6245, N6232, N5954);
nand NAND2 (N6246, N6228, N5316);
nor NOR4 (N6247, N6241, N5181, N5432, N5593);
nand NAND3 (N6248, N6216, N5945, N431);
nand NAND3 (N6249, N6242, N3278, N5864);
and AND3 (N6250, N6243, N3012, N1589);
nand NAND2 (N6251, N6247, N5532);
xor XOR2 (N6252, N6245, N5474);
xor XOR2 (N6253, N6249, N2336);
or OR2 (N6254, N6248, N487);
not NOT1 (N6255, N6244);
or OR2 (N6256, N6251, N266);
and AND2 (N6257, N6254, N5438);
and AND2 (N6258, N6253, N1730);
xor XOR2 (N6259, N6255, N5446);
and AND3 (N6260, N6259, N125, N2671);
nor NOR4 (N6261, N6220, N778, N103, N5378);
and AND4 (N6262, N6256, N126, N134, N4276);
buf BUF1 (N6263, N6258);
nor NOR2 (N6264, N6262, N3802);
nor NOR4 (N6265, N6246, N2477, N3926, N404);
buf BUF1 (N6266, N6240);
xor XOR2 (N6267, N6265, N6160);
nand NAND4 (N6268, N6252, N597, N4953, N2961);
not NOT1 (N6269, N6268);
not NOT1 (N6270, N6261);
and AND3 (N6271, N6269, N2911, N5678);
xor XOR2 (N6272, N6238, N564);
buf BUF1 (N6273, N6257);
xor XOR2 (N6274, N6270, N3828);
nor NOR2 (N6275, N6266, N4568);
or OR3 (N6276, N6273, N4875, N1210);
or OR2 (N6277, N6263, N883);
and AND2 (N6278, N6272, N2570);
and AND2 (N6279, N6278, N3349);
nand NAND2 (N6280, N6267, N1689);
and AND4 (N6281, N6275, N5716, N2951, N3577);
nand NAND2 (N6282, N6250, N5188);
and AND2 (N6283, N6260, N2793);
xor XOR2 (N6284, N6271, N2417);
xor XOR2 (N6285, N6283, N4588);
not NOT1 (N6286, N6281);
not NOT1 (N6287, N6279);
and AND4 (N6288, N6285, N4756, N1475, N3686);
and AND2 (N6289, N6274, N2866);
and AND3 (N6290, N6284, N2291, N1068);
nand NAND2 (N6291, N6277, N2906);
not NOT1 (N6292, N6290);
nand NAND3 (N6293, N6288, N5235, N2941);
buf BUF1 (N6294, N6276);
buf BUF1 (N6295, N6286);
buf BUF1 (N6296, N6292);
and AND4 (N6297, N6289, N4300, N3457, N5891);
not NOT1 (N6298, N6293);
xor XOR2 (N6299, N6264, N16);
and AND3 (N6300, N6296, N5064, N4627);
buf BUF1 (N6301, N6287);
not NOT1 (N6302, N6301);
or OR4 (N6303, N6291, N5452, N1866, N5748);
or OR2 (N6304, N6299, N4116);
or OR2 (N6305, N6304, N185);
not NOT1 (N6306, N6300);
buf BUF1 (N6307, N6282);
not NOT1 (N6308, N6305);
not NOT1 (N6309, N6298);
and AND4 (N6310, N6303, N4748, N2177, N5724);
not NOT1 (N6311, N6306);
nor NOR3 (N6312, N6311, N881, N4095);
nand NAND3 (N6313, N6297, N3969, N1924);
and AND3 (N6314, N6308, N5123, N4996);
not NOT1 (N6315, N6302);
not NOT1 (N6316, N6294);
and AND3 (N6317, N6295, N2677, N836);
or OR4 (N6318, N6309, N805, N2730, N1611);
or OR3 (N6319, N6314, N898, N905);
nand NAND4 (N6320, N6316, N6025, N3369, N4793);
nand NAND2 (N6321, N6318, N4473);
xor XOR2 (N6322, N6317, N6101);
nand NAND3 (N6323, N6307, N2828, N5588);
nor NOR3 (N6324, N6313, N679, N5067);
not NOT1 (N6325, N6322);
nand NAND4 (N6326, N6280, N2070, N5600, N2602);
not NOT1 (N6327, N6320);
and AND2 (N6328, N6323, N2373);
buf BUF1 (N6329, N6319);
xor XOR2 (N6330, N6321, N2990);
nand NAND4 (N6331, N6315, N243, N1674, N3213);
buf BUF1 (N6332, N6324);
and AND3 (N6333, N6328, N4457, N2523);
not NOT1 (N6334, N6312);
or OR2 (N6335, N6333, N2511);
or OR4 (N6336, N6330, N4877, N3689, N2879);
nand NAND4 (N6337, N6327, N6265, N3906, N1524);
not NOT1 (N6338, N6331);
nand NAND3 (N6339, N6326, N4358, N40);
buf BUF1 (N6340, N6329);
not NOT1 (N6341, N6334);
nand NAND4 (N6342, N6341, N2817, N6000, N6146);
not NOT1 (N6343, N6325);
xor XOR2 (N6344, N6339, N600);
xor XOR2 (N6345, N6344, N3680);
nor NOR2 (N6346, N6310, N1020);
and AND4 (N6347, N6335, N366, N3511, N3829);
and AND4 (N6348, N6336, N964, N4152, N3398);
or OR2 (N6349, N6337, N3617);
buf BUF1 (N6350, N6343);
xor XOR2 (N6351, N6350, N2458);
buf BUF1 (N6352, N6345);
or OR3 (N6353, N6346, N1287, N721);
or OR3 (N6354, N6347, N408, N4274);
nand NAND2 (N6355, N6342, N5038);
and AND4 (N6356, N6355, N5205, N194, N5835);
nor NOR4 (N6357, N6352, N1180, N277, N2672);
nand NAND4 (N6358, N6351, N1437, N401, N1364);
buf BUF1 (N6359, N6353);
or OR4 (N6360, N6338, N82, N972, N781);
buf BUF1 (N6361, N6348);
nor NOR2 (N6362, N6356, N2423);
nand NAND3 (N6363, N6358, N1933, N314);
buf BUF1 (N6364, N6362);
and AND4 (N6365, N6354, N3192, N3196, N1392);
nor NOR3 (N6366, N6363, N5731, N2564);
nor NOR3 (N6367, N6332, N5259, N3769);
xor XOR2 (N6368, N6349, N2269);
nand NAND4 (N6369, N6359, N2924, N3528, N2182);
or OR4 (N6370, N6368, N4331, N3176, N5623);
and AND2 (N6371, N6357, N4709);
and AND2 (N6372, N6365, N4693);
buf BUF1 (N6373, N6361);
nand NAND2 (N6374, N6360, N2081);
not NOT1 (N6375, N6367);
not NOT1 (N6376, N6374);
buf BUF1 (N6377, N6366);
nor NOR3 (N6378, N6375, N2557, N3556);
not NOT1 (N6379, N6370);
xor XOR2 (N6380, N6376, N1592);
or OR2 (N6381, N6340, N4039);
or OR3 (N6382, N6377, N6340, N5230);
or OR2 (N6383, N6381, N3789);
xor XOR2 (N6384, N6371, N1609);
and AND4 (N6385, N6372, N3330, N4277, N2049);
not NOT1 (N6386, N6380);
not NOT1 (N6387, N6384);
nand NAND3 (N6388, N6378, N6149, N4519);
nor NOR4 (N6389, N6382, N2380, N2454, N3555);
nor NOR2 (N6390, N6373, N5659);
nor NOR2 (N6391, N6388, N400);
not NOT1 (N6392, N6379);
and AND3 (N6393, N6389, N1712, N5180);
nor NOR4 (N6394, N6369, N3202, N2061, N4623);
or OR3 (N6395, N6385, N5040, N2419);
not NOT1 (N6396, N6395);
xor XOR2 (N6397, N6393, N6132);
buf BUF1 (N6398, N6387);
nor NOR4 (N6399, N6364, N4333, N1841, N5847);
or OR3 (N6400, N6398, N175, N506);
not NOT1 (N6401, N6391);
buf BUF1 (N6402, N6394);
or OR3 (N6403, N6397, N2436, N1376);
not NOT1 (N6404, N6383);
nor NOR2 (N6405, N6399, N841);
nor NOR3 (N6406, N6386, N2648, N6318);
or OR2 (N6407, N6392, N4566);
nand NAND4 (N6408, N6396, N5556, N2277, N4673);
buf BUF1 (N6409, N6390);
and AND2 (N6410, N6400, N1832);
not NOT1 (N6411, N6406);
and AND4 (N6412, N6409, N216, N3470, N2954);
buf BUF1 (N6413, N6401);
not NOT1 (N6414, N6407);
nor NOR4 (N6415, N6408, N3562, N431, N452);
and AND4 (N6416, N6412, N6055, N3914, N489);
and AND4 (N6417, N6402, N2674, N1110, N92);
not NOT1 (N6418, N6403);
xor XOR2 (N6419, N6417, N4861);
xor XOR2 (N6420, N6410, N4907);
and AND4 (N6421, N6413, N3460, N2909, N2191);
or OR2 (N6422, N6411, N2983);
or OR4 (N6423, N6415, N543, N4683, N5215);
nand NAND3 (N6424, N6414, N4331, N4062);
xor XOR2 (N6425, N6416, N734);
and AND2 (N6426, N6418, N796);
buf BUF1 (N6427, N6419);
or OR4 (N6428, N6427, N6255, N4678, N692);
and AND3 (N6429, N6426, N2085, N4470);
not NOT1 (N6430, N6423);
or OR4 (N6431, N6424, N5700, N4185, N5777);
or OR3 (N6432, N6431, N1326, N2079);
and AND3 (N6433, N6425, N2754, N5348);
not NOT1 (N6434, N6429);
xor XOR2 (N6435, N6422, N5720);
xor XOR2 (N6436, N6435, N6238);
and AND4 (N6437, N6436, N214, N1895, N5190);
nor NOR4 (N6438, N6434, N1370, N5181, N478);
xor XOR2 (N6439, N6421, N5920);
and AND2 (N6440, N6430, N575);
buf BUF1 (N6441, N6420);
nor NOR2 (N6442, N6440, N4015);
not NOT1 (N6443, N6439);
xor XOR2 (N6444, N6428, N5387);
or OR3 (N6445, N6441, N41, N3934);
xor XOR2 (N6446, N6438, N245);
nor NOR4 (N6447, N6443, N3451, N5620, N1049);
or OR4 (N6448, N6446, N1695, N1729, N3235);
or OR2 (N6449, N6442, N896);
nor NOR2 (N6450, N6405, N3816);
nand NAND4 (N6451, N6437, N1044, N4890, N1741);
nor NOR2 (N6452, N6432, N5316);
xor XOR2 (N6453, N6445, N734);
nand NAND3 (N6454, N6451, N3778, N1170);
buf BUF1 (N6455, N6444);
xor XOR2 (N6456, N6454, N4844);
buf BUF1 (N6457, N6452);
nor NOR4 (N6458, N6450, N1425, N3476, N2981);
xor XOR2 (N6459, N6456, N31);
buf BUF1 (N6460, N6448);
or OR3 (N6461, N6404, N5658, N3774);
or OR3 (N6462, N6461, N534, N3138);
nor NOR3 (N6463, N6457, N2935, N6421);
nand NAND4 (N6464, N6460, N6397, N5046, N4759);
nand NAND2 (N6465, N6433, N1131);
nand NAND4 (N6466, N6447, N824, N4123, N4007);
nand NAND2 (N6467, N6453, N4808);
not NOT1 (N6468, N6449);
nand NAND4 (N6469, N6463, N5148, N5004, N3335);
not NOT1 (N6470, N6458);
or OR4 (N6471, N6465, N1364, N384, N2046);
nor NOR3 (N6472, N6470, N4465, N4289);
or OR2 (N6473, N6455, N5130);
or OR2 (N6474, N6466, N2365);
nand NAND3 (N6475, N6474, N3830, N1216);
and AND2 (N6476, N6475, N1426);
nor NOR2 (N6477, N6467, N5935);
or OR4 (N6478, N6473, N3512, N3708, N6360);
buf BUF1 (N6479, N6478);
nand NAND3 (N6480, N6468, N972, N4400);
and AND2 (N6481, N6472, N3810);
and AND3 (N6482, N6480, N3695, N2145);
nor NOR2 (N6483, N6477, N2606);
xor XOR2 (N6484, N6471, N4003);
nor NOR4 (N6485, N6469, N4198, N6000, N5132);
buf BUF1 (N6486, N6483);
and AND3 (N6487, N6482, N6279, N5779);
not NOT1 (N6488, N6481);
xor XOR2 (N6489, N6476, N4758);
and AND4 (N6490, N6459, N3936, N4220, N3090);
buf BUF1 (N6491, N6464);
not NOT1 (N6492, N6486);
nor NOR2 (N6493, N6479, N5971);
or OR2 (N6494, N6462, N2472);
xor XOR2 (N6495, N6492, N2292);
buf BUF1 (N6496, N6488);
not NOT1 (N6497, N6487);
or OR3 (N6498, N6485, N3192, N2367);
xor XOR2 (N6499, N6494, N3684);
buf BUF1 (N6500, N6484);
or OR3 (N6501, N6500, N1208, N3618);
not NOT1 (N6502, N6493);
nor NOR3 (N6503, N6499, N1474, N2892);
nand NAND4 (N6504, N6495, N5740, N610, N382);
nor NOR3 (N6505, N6497, N289, N6464);
buf BUF1 (N6506, N6498);
not NOT1 (N6507, N6503);
and AND3 (N6508, N6505, N4313, N4966);
and AND3 (N6509, N6496, N5623, N5132);
not NOT1 (N6510, N6509);
buf BUF1 (N6511, N6502);
nor NOR2 (N6512, N6490, N4512);
nand NAND2 (N6513, N6512, N2052);
or OR4 (N6514, N6506, N1520, N5733, N182);
buf BUF1 (N6515, N6504);
nand NAND4 (N6516, N6513, N1502, N2268, N5810);
buf BUF1 (N6517, N6510);
xor XOR2 (N6518, N6491, N6089);
nor NOR3 (N6519, N6517, N5592, N3744);
nand NAND2 (N6520, N6518, N3716);
or OR2 (N6521, N6515, N4424);
nor NOR2 (N6522, N6511, N6187);
xor XOR2 (N6523, N6521, N2850);
nand NAND3 (N6524, N6520, N2937, N3729);
and AND2 (N6525, N6519, N928);
nor NOR3 (N6526, N6525, N54, N1537);
or OR3 (N6527, N6508, N4382, N4835);
or OR3 (N6528, N6526, N2249, N5669);
buf BUF1 (N6529, N6507);
nand NAND3 (N6530, N6527, N4301, N4185);
and AND3 (N6531, N6524, N2256, N3149);
xor XOR2 (N6532, N6501, N3373);
buf BUF1 (N6533, N6528);
buf BUF1 (N6534, N6514);
xor XOR2 (N6535, N6531, N6217);
xor XOR2 (N6536, N6516, N4114);
nand NAND2 (N6537, N6523, N2834);
or OR2 (N6538, N6533, N5187);
nor NOR4 (N6539, N6538, N2281, N5011, N2153);
or OR2 (N6540, N6532, N5483);
not NOT1 (N6541, N6534);
nand NAND4 (N6542, N6536, N4557, N2033, N5663);
buf BUF1 (N6543, N6535);
and AND3 (N6544, N6540, N5646, N3617);
buf BUF1 (N6545, N6529);
or OR4 (N6546, N6541, N1876, N3973, N1267);
not NOT1 (N6547, N6543);
nand NAND3 (N6548, N6544, N2012, N5692);
nor NOR3 (N6549, N6530, N2375, N3765);
nand NAND2 (N6550, N6545, N4445);
nor NOR3 (N6551, N6546, N3956, N4685);
buf BUF1 (N6552, N6542);
and AND2 (N6553, N6522, N600);
not NOT1 (N6554, N6547);
buf BUF1 (N6555, N6489);
or OR3 (N6556, N6539, N2419, N6474);
or OR2 (N6557, N6556, N3346);
buf BUF1 (N6558, N6555);
nand NAND3 (N6559, N6551, N4500, N829);
not NOT1 (N6560, N6558);
buf BUF1 (N6561, N6549);
nor NOR2 (N6562, N6550, N5492);
xor XOR2 (N6563, N6561, N2885);
and AND2 (N6564, N6563, N5426);
or OR3 (N6565, N6554, N1134, N1730);
not NOT1 (N6566, N6565);
or OR4 (N6567, N6537, N3127, N4403, N5236);
nand NAND3 (N6568, N6560, N413, N654);
buf BUF1 (N6569, N6559);
xor XOR2 (N6570, N6553, N4262);
not NOT1 (N6571, N6567);
xor XOR2 (N6572, N6569, N3997);
buf BUF1 (N6573, N6572);
or OR4 (N6574, N6564, N155, N1127, N5519);
nor NOR3 (N6575, N6573, N426, N5569);
nor NOR2 (N6576, N6566, N5888);
not NOT1 (N6577, N6562);
nand NAND4 (N6578, N6575, N3545, N3109, N4073);
nand NAND4 (N6579, N6557, N2040, N3844, N6553);
buf BUF1 (N6580, N6576);
xor XOR2 (N6581, N6552, N5192);
nand NAND3 (N6582, N6548, N3137, N1401);
and AND3 (N6583, N6582, N744, N4450);
xor XOR2 (N6584, N6579, N6537);
xor XOR2 (N6585, N6568, N2975);
buf BUF1 (N6586, N6581);
and AND2 (N6587, N6586, N796);
nand NAND2 (N6588, N6580, N4786);
not NOT1 (N6589, N6571);
and AND4 (N6590, N6585, N443, N3245, N4631);
or OR2 (N6591, N6587, N2964);
xor XOR2 (N6592, N6570, N5997);
xor XOR2 (N6593, N6589, N6042);
nand NAND3 (N6594, N6591, N3004, N1622);
nor NOR2 (N6595, N6584, N6388);
not NOT1 (N6596, N6577);
nor NOR2 (N6597, N6592, N1101);
not NOT1 (N6598, N6578);
xor XOR2 (N6599, N6593, N3683);
or OR4 (N6600, N6599, N1157, N2098, N4508);
nor NOR4 (N6601, N6588, N5004, N6279, N5659);
nand NAND2 (N6602, N6600, N5350);
xor XOR2 (N6603, N6597, N2192);
not NOT1 (N6604, N6590);
buf BUF1 (N6605, N6594);
not NOT1 (N6606, N6598);
nand NAND3 (N6607, N6604, N4484, N597);
buf BUF1 (N6608, N6602);
or OR2 (N6609, N6596, N3714);
nor NOR2 (N6610, N6601, N3777);
not NOT1 (N6611, N6605);
nor NOR3 (N6612, N6603, N5440, N1251);
nor NOR3 (N6613, N6608, N3262, N2382);
and AND2 (N6614, N6612, N6247);
xor XOR2 (N6615, N6614, N154);
nand NAND3 (N6616, N6611, N4182, N3162);
nor NOR2 (N6617, N6583, N3071);
nand NAND3 (N6618, N6574, N863, N4105);
nand NAND3 (N6619, N6615, N4265, N2679);
not NOT1 (N6620, N6616);
nor NOR3 (N6621, N6610, N4837, N5788);
nand NAND3 (N6622, N6595, N3416, N4010);
and AND4 (N6623, N6613, N4772, N2976, N1378);
not NOT1 (N6624, N6619);
nand NAND2 (N6625, N6606, N2554);
or OR2 (N6626, N6607, N2903);
buf BUF1 (N6627, N6623);
nand NAND2 (N6628, N6627, N3295);
not NOT1 (N6629, N6618);
and AND3 (N6630, N6629, N1647, N4153);
buf BUF1 (N6631, N6625);
and AND4 (N6632, N6621, N3031, N6036, N3597);
buf BUF1 (N6633, N6628);
buf BUF1 (N6634, N6626);
nand NAND2 (N6635, N6632, N4877);
not NOT1 (N6636, N6620);
nor NOR4 (N6637, N6634, N1805, N884, N2941);
buf BUF1 (N6638, N6624);
or OR3 (N6639, N6630, N314, N2146);
nand NAND2 (N6640, N6637, N2908);
and AND3 (N6641, N6631, N4974, N3501);
xor XOR2 (N6642, N6640, N6272);
xor XOR2 (N6643, N6638, N6239);
nand NAND2 (N6644, N6617, N3050);
and AND3 (N6645, N6635, N706, N134);
nand NAND3 (N6646, N6633, N1015, N404);
buf BUF1 (N6647, N6646);
and AND4 (N6648, N6642, N2616, N2064, N3234);
xor XOR2 (N6649, N6644, N3143);
not NOT1 (N6650, N6645);
nor NOR4 (N6651, N6622, N4151, N4674, N4465);
nand NAND4 (N6652, N6609, N2688, N4510, N1673);
buf BUF1 (N6653, N6649);
not NOT1 (N6654, N6647);
or OR3 (N6655, N6648, N4026, N1110);
nor NOR4 (N6656, N6639, N466, N3055, N396);
and AND3 (N6657, N6655, N767, N2157);
xor XOR2 (N6658, N6641, N5938);
buf BUF1 (N6659, N6651);
or OR2 (N6660, N6650, N5536);
xor XOR2 (N6661, N6660, N199);
nand NAND3 (N6662, N6653, N2902, N2403);
xor XOR2 (N6663, N6659, N3524);
nor NOR4 (N6664, N6643, N478, N3814, N1155);
buf BUF1 (N6665, N6662);
or OR2 (N6666, N6654, N1122);
nor NOR3 (N6667, N6663, N5927, N4738);
buf BUF1 (N6668, N6657);
xor XOR2 (N6669, N6667, N6555);
and AND3 (N6670, N6666, N925, N4069);
nor NOR3 (N6671, N6652, N5432, N2160);
or OR3 (N6672, N6665, N4617, N1791);
buf BUF1 (N6673, N6672);
or OR4 (N6674, N6673, N13, N560, N4862);
and AND3 (N6675, N6661, N2320, N139);
nand NAND4 (N6676, N6636, N75, N5376, N5790);
buf BUF1 (N6677, N6668);
nand NAND4 (N6678, N6674, N5622, N1697, N608);
nor NOR4 (N6679, N6669, N3065, N4828, N930);
not NOT1 (N6680, N6671);
xor XOR2 (N6681, N6656, N4913);
buf BUF1 (N6682, N6681);
not NOT1 (N6683, N6678);
nand NAND3 (N6684, N6679, N1333, N78);
buf BUF1 (N6685, N6683);
buf BUF1 (N6686, N6685);
nor NOR3 (N6687, N6684, N4185, N4837);
and AND3 (N6688, N6670, N5433, N1851);
buf BUF1 (N6689, N6682);
nor NOR3 (N6690, N6689, N285, N5377);
buf BUF1 (N6691, N6658);
nand NAND2 (N6692, N6690, N5741);
or OR2 (N6693, N6676, N6405);
or OR2 (N6694, N6693, N412);
and AND4 (N6695, N6686, N6240, N5183, N2280);
nor NOR3 (N6696, N6687, N3026, N4555);
and AND2 (N6697, N6677, N254);
buf BUF1 (N6698, N6691);
nand NAND2 (N6699, N6664, N1432);
not NOT1 (N6700, N6680);
and AND3 (N6701, N6688, N3778, N5421);
and AND2 (N6702, N6696, N6279);
buf BUF1 (N6703, N6702);
or OR2 (N6704, N6699, N1136);
nor NOR3 (N6705, N6694, N2755, N854);
not NOT1 (N6706, N6701);
nand NAND2 (N6707, N6697, N6144);
and AND4 (N6708, N6707, N4067, N5400, N1108);
or OR3 (N6709, N6695, N1861, N4604);
not NOT1 (N6710, N6708);
or OR3 (N6711, N6705, N2810, N4057);
or OR3 (N6712, N6700, N5281, N4257);
or OR4 (N6713, N6710, N3172, N6481, N4616);
buf BUF1 (N6714, N6698);
nand NAND2 (N6715, N6692, N1225);
buf BUF1 (N6716, N6709);
nor NOR2 (N6717, N6703, N5325);
or OR2 (N6718, N6717, N2629);
xor XOR2 (N6719, N6718, N1142);
not NOT1 (N6720, N6675);
nand NAND3 (N6721, N6715, N3816, N6459);
nor NOR4 (N6722, N6713, N3881, N3927, N5546);
not NOT1 (N6723, N6714);
nor NOR4 (N6724, N6719, N3874, N3506, N143);
nand NAND3 (N6725, N6723, N4700, N3735);
nor NOR3 (N6726, N6716, N6328, N5939);
not NOT1 (N6727, N6725);
not NOT1 (N6728, N6724);
and AND4 (N6729, N6711, N3109, N1298, N5859);
xor XOR2 (N6730, N6729, N5221);
or OR4 (N6731, N6722, N2681, N4965, N6253);
and AND2 (N6732, N6704, N3104);
xor XOR2 (N6733, N6721, N468);
xor XOR2 (N6734, N6733, N2654);
and AND2 (N6735, N6731, N6101);
and AND2 (N6736, N6735, N4607);
and AND2 (N6737, N6728, N2518);
buf BUF1 (N6738, N6727);
xor XOR2 (N6739, N6720, N3763);
nor NOR4 (N6740, N6730, N2254, N2359, N2837);
not NOT1 (N6741, N6739);
buf BUF1 (N6742, N6706);
nand NAND3 (N6743, N6738, N369, N1462);
and AND3 (N6744, N6712, N149, N6430);
nand NAND4 (N6745, N6743, N6229, N1650, N4806);
xor XOR2 (N6746, N6734, N5306);
and AND3 (N6747, N6741, N303, N2678);
nor NOR3 (N6748, N6740, N6022, N5907);
xor XOR2 (N6749, N6736, N4290);
xor XOR2 (N6750, N6746, N5226);
buf BUF1 (N6751, N6747);
nor NOR3 (N6752, N6748, N2443, N2305);
xor XOR2 (N6753, N6726, N1748);
xor XOR2 (N6754, N6752, N2079);
not NOT1 (N6755, N6749);
xor XOR2 (N6756, N6750, N3950);
nand NAND3 (N6757, N6751, N2702, N5470);
or OR3 (N6758, N6745, N3307, N1164);
or OR4 (N6759, N6754, N250, N212, N2308);
xor XOR2 (N6760, N6759, N5380);
not NOT1 (N6761, N6742);
buf BUF1 (N6762, N6760);
and AND4 (N6763, N6762, N6461, N1603, N4466);
xor XOR2 (N6764, N6757, N5934);
and AND2 (N6765, N6737, N851);
xor XOR2 (N6766, N6761, N4021);
not NOT1 (N6767, N6756);
nand NAND4 (N6768, N6755, N57, N2723, N6561);
nor NOR2 (N6769, N6765, N2085);
xor XOR2 (N6770, N6753, N1921);
and AND4 (N6771, N6744, N2957, N2096, N6117);
nand NAND4 (N6772, N6764, N4821, N4617, N4911);
nor NOR2 (N6773, N6767, N3367);
nor NOR3 (N6774, N6773, N3837, N746);
and AND3 (N6775, N6771, N5989, N4415);
not NOT1 (N6776, N6763);
not NOT1 (N6777, N6758);
xor XOR2 (N6778, N6768, N4355);
and AND2 (N6779, N6778, N4765);
not NOT1 (N6780, N6766);
or OR2 (N6781, N6776, N4236);
not NOT1 (N6782, N6732);
not NOT1 (N6783, N6777);
buf BUF1 (N6784, N6782);
nand NAND3 (N6785, N6775, N1516, N3197);
xor XOR2 (N6786, N6785, N1950);
not NOT1 (N6787, N6784);
nand NAND4 (N6788, N6774, N1587, N5529, N2278);
and AND3 (N6789, N6770, N2491, N1025);
nand NAND2 (N6790, N6788, N423);
nand NAND2 (N6791, N6783, N3977);
buf BUF1 (N6792, N6787);
buf BUF1 (N6793, N6769);
not NOT1 (N6794, N6789);
buf BUF1 (N6795, N6791);
buf BUF1 (N6796, N6795);
not NOT1 (N6797, N6779);
and AND2 (N6798, N6790, N4682);
and AND2 (N6799, N6798, N3385);
or OR4 (N6800, N6780, N4281, N4997, N3334);
xor XOR2 (N6801, N6796, N2423);
or OR4 (N6802, N6800, N3756, N6649, N4317);
xor XOR2 (N6803, N6793, N2698);
xor XOR2 (N6804, N6803, N2773);
xor XOR2 (N6805, N6781, N847);
buf BUF1 (N6806, N6802);
not NOT1 (N6807, N6805);
and AND3 (N6808, N6786, N5640, N1215);
or OR4 (N6809, N6806, N6209, N955, N4428);
nor NOR4 (N6810, N6794, N2575, N2522, N452);
nor NOR3 (N6811, N6804, N2321, N1883);
and AND4 (N6812, N6810, N6688, N1922, N3911);
xor XOR2 (N6813, N6797, N932);
or OR4 (N6814, N6811, N326, N2890, N701);
and AND3 (N6815, N6807, N5536, N1079);
or OR4 (N6816, N6814, N21, N2350, N5200);
xor XOR2 (N6817, N6816, N5613);
or OR4 (N6818, N6815, N3741, N1388, N294);
and AND2 (N6819, N6817, N6027);
nor NOR2 (N6820, N6818, N3501);
not NOT1 (N6821, N6799);
not NOT1 (N6822, N6820);
and AND4 (N6823, N6808, N5003, N1986, N5444);
nor NOR4 (N6824, N6812, N5379, N696, N1938);
nor NOR2 (N6825, N6819, N4623);
buf BUF1 (N6826, N6821);
nor NOR2 (N6827, N6822, N4459);
or OR2 (N6828, N6772, N4589);
nand NAND3 (N6829, N6801, N1391, N1667);
nor NOR2 (N6830, N6809, N2709);
not NOT1 (N6831, N6813);
nand NAND2 (N6832, N6826, N4554);
xor XOR2 (N6833, N6829, N5494);
nand NAND2 (N6834, N6827, N4627);
not NOT1 (N6835, N6834);
and AND3 (N6836, N6824, N824, N4285);
xor XOR2 (N6837, N6792, N1102);
and AND3 (N6838, N6836, N3242, N2639);
buf BUF1 (N6839, N6833);
and AND4 (N6840, N6823, N149, N6211, N6194);
buf BUF1 (N6841, N6839);
buf BUF1 (N6842, N6825);
or OR4 (N6843, N6831, N4557, N5376, N2272);
nand NAND2 (N6844, N6832, N753);
not NOT1 (N6845, N6843);
nand NAND4 (N6846, N6844, N5114, N6742, N5777);
or OR4 (N6847, N6838, N3873, N6841, N2418);
nor NOR3 (N6848, N783, N2316, N657);
nand NAND3 (N6849, N6840, N6506, N1809);
not NOT1 (N6850, N6828);
xor XOR2 (N6851, N6846, N6042);
not NOT1 (N6852, N6842);
buf BUF1 (N6853, N6852);
and AND2 (N6854, N6851, N4262);
not NOT1 (N6855, N6847);
buf BUF1 (N6856, N6830);
nand NAND2 (N6857, N6854, N388);
xor XOR2 (N6858, N6857, N3064);
nor NOR2 (N6859, N6835, N5983);
buf BUF1 (N6860, N6853);
nor NOR2 (N6861, N6837, N466);
and AND4 (N6862, N6860, N2296, N253, N2438);
and AND2 (N6863, N6862, N2402);
xor XOR2 (N6864, N6849, N4081);
or OR3 (N6865, N6845, N2685, N2504);
and AND4 (N6866, N6848, N2916, N3379, N5614);
xor XOR2 (N6867, N6861, N1797);
not NOT1 (N6868, N6859);
xor XOR2 (N6869, N6850, N4960);
and AND4 (N6870, N6863, N6379, N6390, N2987);
or OR2 (N6871, N6868, N5616);
nand NAND3 (N6872, N6870, N3992, N862);
nand NAND4 (N6873, N6858, N3768, N4210, N5304);
xor XOR2 (N6874, N6871, N2319);
not NOT1 (N6875, N6856);
not NOT1 (N6876, N6872);
xor XOR2 (N6877, N6864, N1018);
nand NAND4 (N6878, N6874, N4078, N1518, N890);
buf BUF1 (N6879, N6875);
nor NOR4 (N6880, N6865, N5729, N3062, N6372);
buf BUF1 (N6881, N6855);
and AND2 (N6882, N6876, N2084);
buf BUF1 (N6883, N6879);
not NOT1 (N6884, N6883);
nand NAND3 (N6885, N6880, N32, N4350);
nor NOR3 (N6886, N6873, N4878, N774);
or OR2 (N6887, N6867, N2499);
not NOT1 (N6888, N6881);
not NOT1 (N6889, N6882);
xor XOR2 (N6890, N6878, N6061);
or OR3 (N6891, N6886, N2970, N5846);
and AND3 (N6892, N6866, N4640, N2861);
buf BUF1 (N6893, N6891);
or OR2 (N6894, N6893, N6462);
nor NOR2 (N6895, N6894, N2463);
buf BUF1 (N6896, N6890);
nor NOR2 (N6897, N6887, N2369);
nand NAND2 (N6898, N6889, N3922);
not NOT1 (N6899, N6898);
and AND2 (N6900, N6888, N5348);
or OR2 (N6901, N6900, N6010);
xor XOR2 (N6902, N6877, N2478);
xor XOR2 (N6903, N6869, N1044);
xor XOR2 (N6904, N6901, N1811);
and AND4 (N6905, N6892, N2320, N5916, N4909);
nand NAND4 (N6906, N6903, N787, N1050, N4067);
xor XOR2 (N6907, N6906, N1620);
not NOT1 (N6908, N6897);
or OR2 (N6909, N6899, N5281);
nor NOR2 (N6910, N6902, N4582);
xor XOR2 (N6911, N6895, N6371);
or OR2 (N6912, N6908, N6348);
nand NAND3 (N6913, N6912, N4064, N5235);
not NOT1 (N6914, N6907);
nor NOR2 (N6915, N6884, N5093);
not NOT1 (N6916, N6905);
or OR2 (N6917, N6909, N277);
and AND2 (N6918, N6917, N1223);
nor NOR4 (N6919, N6904, N6745, N6426, N5215);
not NOT1 (N6920, N6913);
or OR3 (N6921, N6914, N2487, N1350);
xor XOR2 (N6922, N6919, N5848);
xor XOR2 (N6923, N6922, N3217);
not NOT1 (N6924, N6915);
nor NOR2 (N6925, N6923, N2265);
nand NAND4 (N6926, N6918, N2218, N4184, N3001);
and AND3 (N6927, N6920, N6149, N6764);
nand NAND2 (N6928, N6885, N4637);
not NOT1 (N6929, N6896);
nand NAND4 (N6930, N6910, N3800, N5377, N2900);
nand NAND4 (N6931, N6929, N40, N5669, N216);
not NOT1 (N6932, N6930);
and AND3 (N6933, N6927, N6522, N2611);
nor NOR2 (N6934, N6911, N113);
or OR3 (N6935, N6925, N1373, N4799);
or OR3 (N6936, N6935, N6647, N1716);
and AND2 (N6937, N6926, N4064);
nor NOR4 (N6938, N6934, N5732, N6129, N2476);
nand NAND2 (N6939, N6933, N6298);
xor XOR2 (N6940, N6938, N1149);
not NOT1 (N6941, N6939);
nor NOR2 (N6942, N6936, N6302);
or OR2 (N6943, N6928, N934);
or OR2 (N6944, N6943, N94);
xor XOR2 (N6945, N6944, N2614);
not NOT1 (N6946, N6940);
buf BUF1 (N6947, N6924);
not NOT1 (N6948, N6942);
nor NOR4 (N6949, N6937, N2241, N4864, N6655);
not NOT1 (N6950, N6947);
and AND3 (N6951, N6941, N114, N2019);
and AND2 (N6952, N6932, N6233);
buf BUF1 (N6953, N6946);
nand NAND3 (N6954, N6953, N1354, N5836);
nand NAND4 (N6955, N6945, N6816, N2400, N6845);
nor NOR4 (N6956, N6950, N5377, N3951, N2507);
nand NAND2 (N6957, N6916, N4658);
not NOT1 (N6958, N6951);
buf BUF1 (N6959, N6958);
nand NAND3 (N6960, N6956, N4271, N5136);
not NOT1 (N6961, N6921);
xor XOR2 (N6962, N6948, N714);
nor NOR3 (N6963, N6955, N3807, N4394);
or OR3 (N6964, N6957, N1419, N4583);
nor NOR3 (N6965, N6961, N89, N6762);
nor NOR3 (N6966, N6964, N5491, N3726);
or OR3 (N6967, N6962, N2649, N1704);
and AND3 (N6968, N6952, N6548, N6181);
nor NOR4 (N6969, N6965, N4379, N1195, N1291);
buf BUF1 (N6970, N6954);
nor NOR4 (N6971, N6963, N6558, N2605, N5688);
nor NOR3 (N6972, N6959, N5634, N6395);
and AND4 (N6973, N6972, N4180, N3239, N90);
not NOT1 (N6974, N6949);
and AND2 (N6975, N6973, N5611);
nor NOR4 (N6976, N6966, N426, N4144, N6599);
xor XOR2 (N6977, N6974, N2472);
and AND3 (N6978, N6967, N2194, N2061);
xor XOR2 (N6979, N6971, N5610);
or OR2 (N6980, N6977, N436);
nand NAND3 (N6981, N6960, N3528, N3276);
and AND3 (N6982, N6978, N1795, N5893);
xor XOR2 (N6983, N6980, N2944);
xor XOR2 (N6984, N6975, N3818);
not NOT1 (N6985, N6982);
or OR4 (N6986, N6970, N189, N5200, N2675);
or OR2 (N6987, N6986, N2559);
or OR2 (N6988, N6987, N883);
nand NAND3 (N6989, N6985, N2194, N5193);
nand NAND3 (N6990, N6976, N2594, N2414);
and AND4 (N6991, N6981, N6769, N5924, N3395);
buf BUF1 (N6992, N6969);
buf BUF1 (N6993, N6968);
or OR4 (N6994, N6993, N4178, N772, N3321);
nand NAND3 (N6995, N6984, N1829, N6901);
xor XOR2 (N6996, N6988, N3387);
and AND2 (N6997, N6989, N1544);
nor NOR4 (N6998, N6994, N6093, N2725, N2526);
not NOT1 (N6999, N6995);
nor NOR3 (N7000, N6992, N2704, N4274);
xor XOR2 (N7001, N6931, N5474);
not NOT1 (N7002, N6998);
nor NOR4 (N7003, N7001, N1712, N4383, N981);
xor XOR2 (N7004, N7003, N6838);
and AND4 (N7005, N6996, N6103, N5073, N5142);
not NOT1 (N7006, N6990);
not NOT1 (N7007, N6997);
not NOT1 (N7008, N7000);
buf BUF1 (N7009, N6999);
buf BUF1 (N7010, N7005);
not NOT1 (N7011, N7010);
and AND3 (N7012, N7009, N4794, N6905);
nand NAND2 (N7013, N7008, N1357);
and AND4 (N7014, N6979, N4584, N6202, N4732);
buf BUF1 (N7015, N7004);
xor XOR2 (N7016, N7013, N6137);
not NOT1 (N7017, N6991);
buf BUF1 (N7018, N7016);
nor NOR2 (N7019, N7007, N2382);
nand NAND2 (N7020, N7012, N6479);
or OR3 (N7021, N7002, N679, N5340);
and AND2 (N7022, N7021, N254);
buf BUF1 (N7023, N6983);
buf BUF1 (N7024, N7018);
not NOT1 (N7025, N7014);
or OR3 (N7026, N7022, N2058, N3031);
not NOT1 (N7027, N7011);
not NOT1 (N7028, N7026);
not NOT1 (N7029, N7015);
nand NAND4 (N7030, N7017, N5032, N1984, N866);
not NOT1 (N7031, N7023);
buf BUF1 (N7032, N7025);
and AND3 (N7033, N7020, N5243, N1419);
nor NOR3 (N7034, N7030, N3035, N3490);
nand NAND3 (N7035, N7033, N2145, N532);
nor NOR3 (N7036, N7027, N660, N1715);
not NOT1 (N7037, N7031);
nand NAND2 (N7038, N7034, N1937);
nor NOR4 (N7039, N7038, N3128, N5500, N381);
not NOT1 (N7040, N7036);
or OR4 (N7041, N7032, N856, N787, N2135);
nand NAND2 (N7042, N7041, N5620);
not NOT1 (N7043, N7042);
not NOT1 (N7044, N7037);
xor XOR2 (N7045, N7035, N2520);
and AND4 (N7046, N7040, N69, N50, N1364);
xor XOR2 (N7047, N7024, N5144);
not NOT1 (N7048, N7019);
nand NAND2 (N7049, N7045, N5496);
or OR4 (N7050, N7029, N2818, N5752, N224);
or OR2 (N7051, N7050, N5256);
not NOT1 (N7052, N7051);
not NOT1 (N7053, N7006);
not NOT1 (N7054, N7049);
nand NAND4 (N7055, N7044, N4969, N294, N2721);
buf BUF1 (N7056, N7047);
or OR4 (N7057, N7046, N269, N1781, N3039);
xor XOR2 (N7058, N7052, N138);
nor NOR3 (N7059, N7039, N4040, N25);
or OR4 (N7060, N7054, N6696, N1445, N6767);
nor NOR4 (N7061, N7057, N6033, N522, N4023);
nand NAND2 (N7062, N7056, N4539);
nor NOR3 (N7063, N7059, N2783, N6430);
and AND3 (N7064, N7053, N3741, N6584);
nand NAND3 (N7065, N7048, N588, N1857);
nor NOR3 (N7066, N7063, N5727, N6273);
buf BUF1 (N7067, N7060);
nor NOR2 (N7068, N7064, N5112);
not NOT1 (N7069, N7062);
nand NAND4 (N7070, N7028, N2144, N6009, N2710);
not NOT1 (N7071, N7061);
and AND2 (N7072, N7068, N1360);
nor NOR4 (N7073, N7066, N2547, N4064, N4113);
xor XOR2 (N7074, N7065, N4769);
and AND4 (N7075, N7067, N2243, N3015, N694);
nor NOR2 (N7076, N7072, N4468);
not NOT1 (N7077, N7055);
buf BUF1 (N7078, N7075);
or OR4 (N7079, N7076, N4248, N2677, N7070);
xor XOR2 (N7080, N2751, N6241);
buf BUF1 (N7081, N7043);
xor XOR2 (N7082, N7073, N2607);
nand NAND4 (N7083, N7079, N6628, N6642, N4394);
nor NOR3 (N7084, N7083, N2212, N2485);
and AND2 (N7085, N7058, N507);
xor XOR2 (N7086, N7069, N3126);
buf BUF1 (N7087, N7080);
xor XOR2 (N7088, N7081, N6370);
not NOT1 (N7089, N7078);
buf BUF1 (N7090, N7074);
and AND2 (N7091, N7086, N1067);
not NOT1 (N7092, N7085);
nand NAND2 (N7093, N7089, N4715);
nand NAND2 (N7094, N7093, N1797);
and AND2 (N7095, N7088, N5650);
and AND4 (N7096, N7092, N797, N3368, N6547);
or OR2 (N7097, N7096, N4261);
xor XOR2 (N7098, N7095, N3757);
xor XOR2 (N7099, N7097, N6981);
nand NAND4 (N7100, N7077, N2329, N1354, N2968);
nor NOR2 (N7101, N7100, N1633);
nand NAND2 (N7102, N7098, N4636);
not NOT1 (N7103, N7091);
nor NOR4 (N7104, N7087, N2191, N3649, N802);
or OR4 (N7105, N7103, N2002, N1444, N3879);
buf BUF1 (N7106, N7090);
or OR4 (N7107, N7099, N5805, N6331, N2799);
and AND2 (N7108, N7101, N2193);
and AND4 (N7109, N7102, N1970, N717, N7056);
not NOT1 (N7110, N7105);
and AND3 (N7111, N7109, N4742, N979);
xor XOR2 (N7112, N7108, N5234);
or OR3 (N7113, N7106, N5518, N2999);
nand NAND4 (N7114, N7111, N5866, N1098, N5171);
nor NOR2 (N7115, N7114, N6746);
nand NAND2 (N7116, N7071, N2514);
or OR2 (N7117, N7113, N6038);
nor NOR4 (N7118, N7110, N1484, N2948, N6730);
buf BUF1 (N7119, N7084);
not NOT1 (N7120, N7082);
buf BUF1 (N7121, N7112);
nand NAND3 (N7122, N7107, N142, N2671);
not NOT1 (N7123, N7119);
xor XOR2 (N7124, N7123, N4230);
or OR4 (N7125, N7118, N4895, N2464, N5047);
nand NAND3 (N7126, N7122, N6592, N6165);
not NOT1 (N7127, N7124);
buf BUF1 (N7128, N7125);
not NOT1 (N7129, N7128);
xor XOR2 (N7130, N7116, N6232);
xor XOR2 (N7131, N7094, N166);
or OR2 (N7132, N7130, N1469);
buf BUF1 (N7133, N7126);
not NOT1 (N7134, N7115);
xor XOR2 (N7135, N7121, N4535);
not NOT1 (N7136, N7120);
or OR4 (N7137, N7104, N3562, N27, N7074);
xor XOR2 (N7138, N7135, N3540);
xor XOR2 (N7139, N7132, N328);
or OR3 (N7140, N7129, N231, N4503);
or OR3 (N7141, N7138, N3210, N6810);
not NOT1 (N7142, N7139);
nor NOR3 (N7143, N7137, N2742, N1528);
and AND2 (N7144, N7133, N4743);
buf BUF1 (N7145, N7134);
xor XOR2 (N7146, N7140, N6556);
nand NAND3 (N7147, N7117, N1586, N3197);
not NOT1 (N7148, N7127);
and AND4 (N7149, N7145, N4110, N6745, N1347);
not NOT1 (N7150, N7144);
not NOT1 (N7151, N7147);
buf BUF1 (N7152, N7131);
not NOT1 (N7153, N7141);
or OR3 (N7154, N7148, N4778, N6452);
buf BUF1 (N7155, N7136);
xor XOR2 (N7156, N7142, N6548);
nor NOR4 (N7157, N7154, N7089, N1204, N3282);
buf BUF1 (N7158, N7152);
and AND4 (N7159, N7151, N1950, N4462, N6150);
buf BUF1 (N7160, N7155);
nor NOR4 (N7161, N7150, N2948, N463, N6183);
or OR4 (N7162, N7157, N6173, N5842, N2211);
not NOT1 (N7163, N7143);
buf BUF1 (N7164, N7149);
nor NOR3 (N7165, N7164, N592, N3354);
nand NAND2 (N7166, N7161, N5399);
or OR3 (N7167, N7163, N1757, N7098);
or OR3 (N7168, N7162, N1978, N857);
xor XOR2 (N7169, N7156, N177);
not NOT1 (N7170, N7166);
or OR3 (N7171, N7165, N6658, N6029);
xor XOR2 (N7172, N7158, N1508);
xor XOR2 (N7173, N7153, N1463);
nor NOR4 (N7174, N7159, N6915, N1036, N1);
nand NAND4 (N7175, N7173, N1336, N3758, N618);
xor XOR2 (N7176, N7167, N2147);
nor NOR3 (N7177, N7169, N4970, N2549);
and AND4 (N7178, N7176, N6514, N1015, N7011);
nor NOR2 (N7179, N7170, N5465);
or OR3 (N7180, N7168, N1386, N5493);
not NOT1 (N7181, N7174);
or OR4 (N7182, N7178, N2883, N1717, N7144);
xor XOR2 (N7183, N7171, N5541);
buf BUF1 (N7184, N7183);
nor NOR3 (N7185, N7146, N6405, N3135);
and AND4 (N7186, N7179, N1428, N2007, N5088);
or OR2 (N7187, N7180, N402);
nand NAND2 (N7188, N7181, N3866);
or OR3 (N7189, N7187, N379, N1755);
buf BUF1 (N7190, N7185);
nor NOR2 (N7191, N7184, N5894);
nand NAND2 (N7192, N7175, N6578);
xor XOR2 (N7193, N7191, N1439);
buf BUF1 (N7194, N7189);
and AND4 (N7195, N7193, N3364, N7152, N5850);
not NOT1 (N7196, N7192);
xor XOR2 (N7197, N7182, N170);
not NOT1 (N7198, N7186);
and AND2 (N7199, N7196, N4241);
xor XOR2 (N7200, N7177, N32);
nand NAND2 (N7201, N7195, N5782);
buf BUF1 (N7202, N7172);
nor NOR3 (N7203, N7197, N5036, N87);
nand NAND2 (N7204, N7201, N4237);
xor XOR2 (N7205, N7199, N797);
xor XOR2 (N7206, N7194, N6611);
xor XOR2 (N7207, N7190, N2992);
buf BUF1 (N7208, N7198);
and AND2 (N7209, N7208, N3638);
nand NAND4 (N7210, N7206, N1165, N2627, N2714);
not NOT1 (N7211, N7203);
xor XOR2 (N7212, N7202, N179);
nor NOR2 (N7213, N7211, N4441);
buf BUF1 (N7214, N7200);
nor NOR4 (N7215, N7160, N649, N3402, N3066);
or OR3 (N7216, N7204, N6579, N5737);
xor XOR2 (N7217, N7207, N4167);
or OR4 (N7218, N7205, N6667, N5464, N1080);
nand NAND2 (N7219, N7188, N6843);
nor NOR4 (N7220, N7212, N5493, N233, N2249);
buf BUF1 (N7221, N7219);
buf BUF1 (N7222, N7221);
xor XOR2 (N7223, N7216, N858);
xor XOR2 (N7224, N7215, N4923);
not NOT1 (N7225, N7223);
nor NOR2 (N7226, N7214, N2171);
buf BUF1 (N7227, N7224);
buf BUF1 (N7228, N7220);
buf BUF1 (N7229, N7210);
not NOT1 (N7230, N7217);
not NOT1 (N7231, N7222);
nor NOR2 (N7232, N7225, N5150);
or OR4 (N7233, N7213, N1404, N5143, N519);
or OR3 (N7234, N7230, N7136, N4642);
and AND2 (N7235, N7227, N122);
nor NOR3 (N7236, N7218, N5921, N6410);
nand NAND2 (N7237, N7234, N5846);
buf BUF1 (N7238, N7229);
nand NAND3 (N7239, N7209, N6809, N892);
nand NAND3 (N7240, N7232, N5948, N3620);
xor XOR2 (N7241, N7240, N3088);
nand NAND4 (N7242, N7231, N6037, N1316, N1662);
nor NOR2 (N7243, N7242, N4139);
or OR3 (N7244, N7238, N1399, N1206);
nand NAND3 (N7245, N7236, N5153, N910);
xor XOR2 (N7246, N7245, N3136);
or OR4 (N7247, N7243, N3712, N970, N3032);
not NOT1 (N7248, N7247);
not NOT1 (N7249, N7239);
nor NOR3 (N7250, N7237, N2969, N4850);
buf BUF1 (N7251, N7228);
xor XOR2 (N7252, N7244, N4452);
not NOT1 (N7253, N7226);
nand NAND2 (N7254, N7246, N70);
buf BUF1 (N7255, N7235);
nand NAND4 (N7256, N7252, N61, N2970, N2806);
nor NOR2 (N7257, N7255, N4996);
and AND4 (N7258, N7249, N7027, N2115, N1098);
or OR4 (N7259, N7257, N5072, N218, N4832);
not NOT1 (N7260, N7250);
buf BUF1 (N7261, N7233);
xor XOR2 (N7262, N7260, N69);
xor XOR2 (N7263, N7262, N57);
or OR3 (N7264, N7261, N4236, N4117);
or OR4 (N7265, N7254, N1877, N2308, N5675);
nor NOR3 (N7266, N7258, N3846, N4455);
nand NAND3 (N7267, N7251, N6971, N6023);
xor XOR2 (N7268, N7256, N4512);
and AND4 (N7269, N7264, N6992, N6977, N6847);
xor XOR2 (N7270, N7265, N7000);
or OR4 (N7271, N7269, N5371, N1878, N2418);
xor XOR2 (N7272, N7259, N7174);
not NOT1 (N7273, N7271);
nor NOR2 (N7274, N7241, N6154);
buf BUF1 (N7275, N7253);
buf BUF1 (N7276, N7268);
not NOT1 (N7277, N7263);
not NOT1 (N7278, N7274);
not NOT1 (N7279, N7277);
xor XOR2 (N7280, N7278, N5056);
buf BUF1 (N7281, N7270);
not NOT1 (N7282, N7267);
nand NAND2 (N7283, N7266, N2173);
or OR2 (N7284, N7248, N165);
xor XOR2 (N7285, N7282, N6761);
and AND4 (N7286, N7284, N4216, N7247, N6420);
and AND3 (N7287, N7275, N3001, N6329);
nor NOR3 (N7288, N7286, N4164, N4145);
nor NOR2 (N7289, N7285, N1264);
or OR3 (N7290, N7273, N321, N227);
or OR2 (N7291, N7290, N6005);
xor XOR2 (N7292, N7281, N4341);
nor NOR3 (N7293, N7272, N1498, N2793);
and AND3 (N7294, N7291, N16, N1593);
xor XOR2 (N7295, N7292, N6575);
and AND2 (N7296, N7276, N3318);
nor NOR3 (N7297, N7293, N275, N6877);
and AND3 (N7298, N7296, N4319, N4521);
or OR2 (N7299, N7294, N4821);
or OR4 (N7300, N7283, N5272, N3489, N3);
and AND3 (N7301, N7297, N1861, N48);
not NOT1 (N7302, N7279);
not NOT1 (N7303, N7300);
not NOT1 (N7304, N7288);
or OR3 (N7305, N7289, N4570, N6818);
and AND4 (N7306, N7287, N1664, N337, N965);
nor NOR4 (N7307, N7304, N2677, N5526, N7221);
not NOT1 (N7308, N7299);
xor XOR2 (N7309, N7302, N567);
xor XOR2 (N7310, N7308, N3984);
nand NAND2 (N7311, N7307, N434);
xor XOR2 (N7312, N7310, N5473);
buf BUF1 (N7313, N7295);
nor NOR4 (N7314, N7305, N3415, N3175, N1757);
nand NAND4 (N7315, N7313, N3769, N5148, N5498);
nand NAND4 (N7316, N7315, N1112, N2079, N6541);
buf BUF1 (N7317, N7301);
buf BUF1 (N7318, N7314);
nor NOR4 (N7319, N7311, N4400, N4615, N430);
nand NAND4 (N7320, N7298, N6700, N1650, N5718);
nor NOR3 (N7321, N7312, N6857, N5301);
nand NAND3 (N7322, N7318, N2097, N266);
and AND3 (N7323, N7309, N4954, N2519);
nor NOR4 (N7324, N7323, N4826, N6743, N2574);
or OR3 (N7325, N7303, N4530, N5746);
buf BUF1 (N7326, N7321);
xor XOR2 (N7327, N7280, N3577);
and AND3 (N7328, N7322, N1224, N836);
xor XOR2 (N7329, N7317, N2513);
xor XOR2 (N7330, N7327, N174);
buf BUF1 (N7331, N7306);
not NOT1 (N7332, N7331);
nand NAND4 (N7333, N7319, N4346, N1187, N6659);
xor XOR2 (N7334, N7330, N2218);
nor NOR4 (N7335, N7328, N2976, N5578, N3864);
buf BUF1 (N7336, N7325);
and AND3 (N7337, N7329, N7296, N4526);
not NOT1 (N7338, N7334);
or OR4 (N7339, N7338, N6963, N1940, N2899);
xor XOR2 (N7340, N7324, N2581);
nand NAND3 (N7341, N7337, N1643, N7325);
not NOT1 (N7342, N7326);
nand NAND3 (N7343, N7332, N1179, N6454);
and AND2 (N7344, N7335, N3305);
xor XOR2 (N7345, N7333, N1663);
nor NOR4 (N7346, N7320, N6954, N5532, N6188);
xor XOR2 (N7347, N7344, N1862);
nor NOR3 (N7348, N7342, N632, N3361);
xor XOR2 (N7349, N7336, N2632);
or OR4 (N7350, N7346, N4639, N996, N2976);
and AND3 (N7351, N7316, N848, N5968);
and AND3 (N7352, N7345, N2481, N1631);
buf BUF1 (N7353, N7340);
or OR3 (N7354, N7351, N1942, N5950);
nand NAND4 (N7355, N7354, N2855, N5430, N4295);
nand NAND3 (N7356, N7350, N4916, N3635);
not NOT1 (N7357, N7348);
or OR4 (N7358, N7356, N3658, N6115, N2040);
xor XOR2 (N7359, N7357, N1528);
xor XOR2 (N7360, N7347, N227);
not NOT1 (N7361, N7360);
and AND4 (N7362, N7349, N4181, N2408, N270);
nand NAND2 (N7363, N7339, N1878);
not NOT1 (N7364, N7362);
buf BUF1 (N7365, N7363);
and AND2 (N7366, N7358, N6402);
buf BUF1 (N7367, N7352);
xor XOR2 (N7368, N7367, N4744);
nand NAND2 (N7369, N7368, N2007);
not NOT1 (N7370, N7364);
nor NOR2 (N7371, N7370, N6614);
not NOT1 (N7372, N7371);
nor NOR2 (N7373, N7365, N304);
nor NOR3 (N7374, N7353, N4110, N5694);
nor NOR2 (N7375, N7361, N6314);
nand NAND3 (N7376, N7372, N2886, N6006);
buf BUF1 (N7377, N7375);
buf BUF1 (N7378, N7341);
buf BUF1 (N7379, N7355);
or OR2 (N7380, N7378, N6179);
or OR4 (N7381, N7366, N6464, N4373, N6918);
and AND2 (N7382, N7343, N2905);
nand NAND3 (N7383, N7376, N5513, N1750);
not NOT1 (N7384, N7383);
buf BUF1 (N7385, N7369);
or OR3 (N7386, N7382, N4879, N1071);
nand NAND2 (N7387, N7374, N2515);
and AND4 (N7388, N7380, N1702, N292, N1369);
nand NAND3 (N7389, N7388, N803, N1783);
buf BUF1 (N7390, N7386);
and AND4 (N7391, N7359, N6527, N653, N4524);
not NOT1 (N7392, N7377);
or OR2 (N7393, N7373, N6570);
nand NAND2 (N7394, N7389, N4048);
or OR4 (N7395, N7381, N2576, N1640, N3027);
not NOT1 (N7396, N7387);
xor XOR2 (N7397, N7395, N2764);
buf BUF1 (N7398, N7390);
not NOT1 (N7399, N7393);
xor XOR2 (N7400, N7398, N931);
nor NOR4 (N7401, N7392, N4383, N3940, N3190);
nand NAND3 (N7402, N7400, N3350, N5365);
nor NOR3 (N7403, N7402, N1270, N7080);
or OR4 (N7404, N7385, N4727, N620, N2976);
xor XOR2 (N7405, N7397, N7049);
or OR3 (N7406, N7379, N1111, N4601);
nand NAND3 (N7407, N7384, N5321, N3340);
and AND4 (N7408, N7394, N2642, N6581, N3763);
or OR3 (N7409, N7401, N5695, N3439);
or OR4 (N7410, N7403, N4427, N1679, N2456);
not NOT1 (N7411, N7406);
xor XOR2 (N7412, N7409, N4611);
nor NOR3 (N7413, N7410, N6136, N1096);
nand NAND3 (N7414, N7404, N1691, N3001);
and AND2 (N7415, N7396, N1050);
xor XOR2 (N7416, N7414, N5958);
nand NAND2 (N7417, N7407, N1405);
and AND4 (N7418, N7413, N3992, N1105, N3628);
xor XOR2 (N7419, N7411, N910);
nand NAND2 (N7420, N7391, N6991);
buf BUF1 (N7421, N7416);
nand NAND4 (N7422, N7408, N5192, N2004, N1393);
and AND4 (N7423, N7419, N3908, N6049, N4880);
nand NAND3 (N7424, N7415, N3055, N574);
and AND3 (N7425, N7417, N6743, N5284);
not NOT1 (N7426, N7421);
buf BUF1 (N7427, N7405);
or OR2 (N7428, N7425, N3685);
xor XOR2 (N7429, N7412, N2322);
xor XOR2 (N7430, N7428, N4480);
nand NAND4 (N7431, N7427, N7216, N5754, N229);
or OR2 (N7432, N7430, N1405);
buf BUF1 (N7433, N7429);
nor NOR2 (N7434, N7433, N2865);
nor NOR3 (N7435, N7418, N5483, N5786);
not NOT1 (N7436, N7420);
nor NOR4 (N7437, N7436, N2197, N3801, N178);
nand NAND3 (N7438, N7437, N6000, N1238);
not NOT1 (N7439, N7435);
nand NAND4 (N7440, N7422, N4362, N7239, N6137);
not NOT1 (N7441, N7432);
and AND4 (N7442, N7424, N1402, N6302, N3309);
xor XOR2 (N7443, N7442, N4733);
and AND4 (N7444, N7438, N5685, N938, N3219);
buf BUF1 (N7445, N7443);
and AND4 (N7446, N7440, N3591, N5511, N7091);
nor NOR2 (N7447, N7444, N3894);
or OR4 (N7448, N7446, N1491, N1279, N7366);
not NOT1 (N7449, N7441);
not NOT1 (N7450, N7426);
and AND3 (N7451, N7448, N5582, N3132);
nand NAND2 (N7452, N7431, N5886);
not NOT1 (N7453, N7451);
nor NOR4 (N7454, N7423, N2957, N2980, N6418);
buf BUF1 (N7455, N7445);
not NOT1 (N7456, N7453);
nor NOR2 (N7457, N7452, N1513);
and AND4 (N7458, N7434, N5653, N511, N6646);
nor NOR3 (N7459, N7454, N1567, N2944);
nor NOR4 (N7460, N7439, N2403, N5706, N6958);
or OR3 (N7461, N7450, N2174, N746);
nand NAND3 (N7462, N7456, N1379, N7443);
and AND2 (N7463, N7447, N5316);
buf BUF1 (N7464, N7463);
nand NAND3 (N7465, N7458, N838, N5242);
and AND3 (N7466, N7464, N1185, N5454);
not NOT1 (N7467, N7455);
buf BUF1 (N7468, N7461);
nor NOR2 (N7469, N7460, N6007);
nand NAND3 (N7470, N7449, N6417, N1830);
not NOT1 (N7471, N7459);
and AND2 (N7472, N7399, N2905);
xor XOR2 (N7473, N7470, N2406);
nand NAND2 (N7474, N7465, N5121);
nor NOR3 (N7475, N7466, N1150, N25);
and AND4 (N7476, N7473, N3900, N3870, N5141);
and AND4 (N7477, N7467, N5183, N7355, N3940);
buf BUF1 (N7478, N7472);
or OR3 (N7479, N7477, N5080, N6845);
or OR4 (N7480, N7471, N3249, N4380, N6568);
or OR2 (N7481, N7474, N5873);
buf BUF1 (N7482, N7469);
buf BUF1 (N7483, N7479);
and AND2 (N7484, N7483, N1890);
and AND4 (N7485, N7457, N1305, N5462, N2550);
xor XOR2 (N7486, N7468, N2827);
xor XOR2 (N7487, N7486, N5411);
or OR2 (N7488, N7481, N2805);
nor NOR3 (N7489, N7484, N6920, N1965);
buf BUF1 (N7490, N7476);
xor XOR2 (N7491, N7487, N4546);
and AND4 (N7492, N7462, N3314, N1990, N5906);
not NOT1 (N7493, N7491);
or OR4 (N7494, N7480, N7215, N4551, N7245);
nand NAND4 (N7495, N7494, N1896, N6576, N4719);
and AND2 (N7496, N7485, N4215);
nor NOR2 (N7497, N7496, N4917);
nand NAND4 (N7498, N7488, N2446, N7429, N174);
and AND2 (N7499, N7492, N4448);
not NOT1 (N7500, N7497);
xor XOR2 (N7501, N7495, N341);
nor NOR2 (N7502, N7493, N5828);
and AND2 (N7503, N7489, N4268);
and AND4 (N7504, N7503, N3525, N4484, N1532);
and AND2 (N7505, N7482, N2980);
nand NAND4 (N7506, N7475, N211, N4033, N6959);
buf BUF1 (N7507, N7499);
and AND2 (N7508, N7498, N2846);
and AND4 (N7509, N7478, N277, N6217, N4395);
xor XOR2 (N7510, N7509, N6369);
xor XOR2 (N7511, N7508, N3469);
buf BUF1 (N7512, N7490);
nor NOR2 (N7513, N7504, N1704);
and AND4 (N7514, N7511, N2370, N5785, N3452);
xor XOR2 (N7515, N7512, N1266);
nand NAND2 (N7516, N7501, N6815);
buf BUF1 (N7517, N7515);
nand NAND2 (N7518, N7500, N4798);
not NOT1 (N7519, N7502);
xor XOR2 (N7520, N7516, N956);
or OR3 (N7521, N7506, N2513, N5058);
nor NOR4 (N7522, N7513, N6723, N3016, N4213);
and AND4 (N7523, N7519, N5855, N779, N5928);
and AND3 (N7524, N7514, N3864, N77);
and AND2 (N7525, N7522, N5591);
or OR2 (N7526, N7521, N5939);
buf BUF1 (N7527, N7507);
buf BUF1 (N7528, N7505);
nor NOR2 (N7529, N7517, N4961);
and AND2 (N7530, N7525, N5015);
buf BUF1 (N7531, N7524);
not NOT1 (N7532, N7520);
or OR2 (N7533, N7529, N3870);
nand NAND4 (N7534, N7518, N1859, N7166, N2316);
or OR2 (N7535, N7527, N185);
xor XOR2 (N7536, N7531, N1113);
not NOT1 (N7537, N7526);
nand NAND2 (N7538, N7528, N2564);
not NOT1 (N7539, N7537);
and AND3 (N7540, N7510, N6042, N3137);
buf BUF1 (N7541, N7536);
nand NAND4 (N7542, N7532, N7343, N5193, N6965);
nor NOR3 (N7543, N7542, N3237, N1825);
buf BUF1 (N7544, N7540);
nand NAND3 (N7545, N7541, N4485, N6415);
nor NOR4 (N7546, N7535, N687, N6329, N6370);
not NOT1 (N7547, N7534);
or OR2 (N7548, N7543, N6225);
xor XOR2 (N7549, N7548, N1260);
not NOT1 (N7550, N7549);
and AND2 (N7551, N7547, N2970);
or OR2 (N7552, N7550, N1043);
not NOT1 (N7553, N7546);
buf BUF1 (N7554, N7523);
and AND2 (N7555, N7539, N600);
nand NAND3 (N7556, N7538, N5616, N7290);
not NOT1 (N7557, N7545);
nor NOR2 (N7558, N7553, N824);
xor XOR2 (N7559, N7557, N2455);
not NOT1 (N7560, N7559);
and AND3 (N7561, N7551, N1170, N3608);
nand NAND4 (N7562, N7561, N6264, N1916, N289);
nand NAND3 (N7563, N7562, N1291, N4768);
xor XOR2 (N7564, N7558, N2863);
or OR2 (N7565, N7560, N5280);
xor XOR2 (N7566, N7552, N6994);
or OR4 (N7567, N7566, N2520, N1601, N3744);
xor XOR2 (N7568, N7544, N588);
buf BUF1 (N7569, N7563);
nand NAND3 (N7570, N7568, N6197, N2157);
nand NAND4 (N7571, N7533, N7465, N6664, N4877);
xor XOR2 (N7572, N7569, N3558);
or OR2 (N7573, N7565, N3883);
and AND2 (N7574, N7556, N3785);
not NOT1 (N7575, N7564);
nand NAND2 (N7576, N7575, N3544);
and AND4 (N7577, N7571, N6375, N2429, N7189);
xor XOR2 (N7578, N7573, N5539);
xor XOR2 (N7579, N7572, N6430);
or OR2 (N7580, N7570, N4659);
buf BUF1 (N7581, N7577);
not NOT1 (N7582, N7576);
buf BUF1 (N7583, N7579);
xor XOR2 (N7584, N7578, N4569);
nor NOR3 (N7585, N7580, N2895, N1620);
nor NOR4 (N7586, N7574, N3242, N1808, N4624);
nand NAND3 (N7587, N7555, N2154, N4324);
or OR4 (N7588, N7585, N3491, N1502, N1087);
nand NAND2 (N7589, N7586, N3254);
and AND2 (N7590, N7567, N2911);
and AND2 (N7591, N7588, N1425);
buf BUF1 (N7592, N7583);
and AND4 (N7593, N7554, N5136, N6323, N2756);
buf BUF1 (N7594, N7592);
or OR2 (N7595, N7594, N5733);
nor NOR4 (N7596, N7582, N6793, N2861, N3014);
nor NOR4 (N7597, N7587, N5207, N3993, N6832);
and AND4 (N7598, N7530, N307, N1265, N6429);
or OR2 (N7599, N7589, N3185);
or OR3 (N7600, N7599, N2854, N2418);
and AND4 (N7601, N7597, N679, N4848, N5363);
xor XOR2 (N7602, N7596, N1567);
not NOT1 (N7603, N7595);
not NOT1 (N7604, N7603);
xor XOR2 (N7605, N7581, N4465);
nor NOR4 (N7606, N7605, N4021, N624, N1027);
xor XOR2 (N7607, N7591, N795);
buf BUF1 (N7608, N7602);
xor XOR2 (N7609, N7601, N6198);
and AND2 (N7610, N7584, N5489);
buf BUF1 (N7611, N7590);
or OR3 (N7612, N7598, N1793, N4245);
nor NOR2 (N7613, N7610, N99);
xor XOR2 (N7614, N7606, N226);
xor XOR2 (N7615, N7593, N5868);
and AND3 (N7616, N7615, N3265, N1272);
or OR4 (N7617, N7608, N4758, N561, N5550);
or OR4 (N7618, N7604, N6538, N5233, N4811);
or OR4 (N7619, N7611, N6251, N6983, N6084);
or OR3 (N7620, N7612, N6309, N479);
buf BUF1 (N7621, N7617);
or OR4 (N7622, N7616, N1854, N6708, N6300);
xor XOR2 (N7623, N7621, N4213);
not NOT1 (N7624, N7614);
xor XOR2 (N7625, N7618, N3228);
buf BUF1 (N7626, N7607);
nand NAND4 (N7627, N7622, N4793, N2688, N2664);
xor XOR2 (N7628, N7613, N6928);
nor NOR2 (N7629, N7624, N280);
xor XOR2 (N7630, N7620, N424);
not NOT1 (N7631, N7609);
nor NOR2 (N7632, N7628, N5646);
not NOT1 (N7633, N7626);
nor NOR3 (N7634, N7629, N2795, N231);
buf BUF1 (N7635, N7630);
nor NOR4 (N7636, N7600, N1072, N4322, N6925);
xor XOR2 (N7637, N7627, N882);
and AND3 (N7638, N7632, N7105, N7621);
or OR2 (N7639, N7637, N3653);
or OR4 (N7640, N7623, N6985, N5418, N260);
and AND2 (N7641, N7636, N779);
and AND3 (N7642, N7639, N5740, N1472);
and AND2 (N7643, N7640, N340);
and AND4 (N7644, N7642, N5628, N2971, N2094);
and AND2 (N7645, N7638, N1556);
not NOT1 (N7646, N7625);
not NOT1 (N7647, N7641);
not NOT1 (N7648, N7619);
buf BUF1 (N7649, N7644);
nand NAND2 (N7650, N7648, N5965);
or OR3 (N7651, N7645, N733, N2511);
nand NAND3 (N7652, N7634, N3858, N5987);
buf BUF1 (N7653, N7643);
or OR4 (N7654, N7647, N5897, N2350, N4755);
xor XOR2 (N7655, N7649, N5196);
buf BUF1 (N7656, N7633);
not NOT1 (N7657, N7656);
buf BUF1 (N7658, N7646);
xor XOR2 (N7659, N7650, N3363);
not NOT1 (N7660, N7659);
and AND3 (N7661, N7657, N6390, N6522);
buf BUF1 (N7662, N7631);
buf BUF1 (N7663, N7658);
and AND3 (N7664, N7635, N4775, N5042);
and AND2 (N7665, N7655, N9);
nand NAND3 (N7666, N7664, N345, N2913);
nand NAND2 (N7667, N7653, N6466);
or OR2 (N7668, N7666, N3914);
xor XOR2 (N7669, N7662, N360);
nand NAND3 (N7670, N7661, N2935, N863);
xor XOR2 (N7671, N7663, N1291);
and AND4 (N7672, N7671, N7240, N4269, N4670);
buf BUF1 (N7673, N7654);
nand NAND3 (N7674, N7669, N4387, N3835);
buf BUF1 (N7675, N7670);
nand NAND4 (N7676, N7674, N6731, N4783, N4716);
not NOT1 (N7677, N7660);
and AND3 (N7678, N7672, N663, N6643);
xor XOR2 (N7679, N7665, N4488);
buf BUF1 (N7680, N7679);
not NOT1 (N7681, N7680);
xor XOR2 (N7682, N7681, N1406);
and AND3 (N7683, N7673, N4086, N6329);
nor NOR3 (N7684, N7678, N7488, N2537);
not NOT1 (N7685, N7667);
xor XOR2 (N7686, N7684, N7122);
nand NAND4 (N7687, N7668, N7553, N1740, N7334);
not NOT1 (N7688, N7651);
xor XOR2 (N7689, N7686, N7043);
nand NAND3 (N7690, N7676, N2420, N1572);
xor XOR2 (N7691, N7689, N4095);
nand NAND3 (N7692, N7675, N1833, N7103);
nand NAND3 (N7693, N7687, N5779, N7511);
nand NAND4 (N7694, N7683, N6803, N7133, N6556);
buf BUF1 (N7695, N7685);
and AND3 (N7696, N7695, N957, N2713);
not NOT1 (N7697, N7693);
nand NAND4 (N7698, N7688, N7316, N4338, N4545);
and AND4 (N7699, N7692, N134, N6199, N920);
nor NOR2 (N7700, N7690, N7124);
nand NAND4 (N7701, N7698, N4615, N123, N1574);
xor XOR2 (N7702, N7699, N7025);
nand NAND4 (N7703, N7697, N2786, N7210, N4984);
or OR4 (N7704, N7682, N1083, N6060, N1710);
nand NAND3 (N7705, N7704, N4758, N1522);
nor NOR2 (N7706, N7701, N2350);
and AND3 (N7707, N7652, N2195, N3067);
buf BUF1 (N7708, N7700);
buf BUF1 (N7709, N7677);
xor XOR2 (N7710, N7705, N4103);
and AND2 (N7711, N7703, N3701);
xor XOR2 (N7712, N7696, N6721);
nand NAND4 (N7713, N7711, N5391, N1197, N3033);
nand NAND4 (N7714, N7706, N2683, N2860, N1516);
and AND2 (N7715, N7710, N5246);
xor XOR2 (N7716, N7713, N1242);
nor NOR4 (N7717, N7712, N982, N5281, N2828);
not NOT1 (N7718, N7702);
and AND3 (N7719, N7694, N3864, N1528);
nand NAND3 (N7720, N7715, N1436, N6691);
not NOT1 (N7721, N7719);
nand NAND2 (N7722, N7716, N7096);
and AND4 (N7723, N7691, N4804, N2280, N6327);
not NOT1 (N7724, N7717);
and AND2 (N7725, N7709, N5557);
or OR3 (N7726, N7721, N7247, N7671);
not NOT1 (N7727, N7722);
nor NOR4 (N7728, N7708, N3036, N1575, N5133);
not NOT1 (N7729, N7718);
nor NOR2 (N7730, N7728, N4436);
not NOT1 (N7731, N7723);
xor XOR2 (N7732, N7726, N6072);
and AND2 (N7733, N7720, N6970);
and AND2 (N7734, N7707, N2551);
or OR3 (N7735, N7714, N539, N6152);
buf BUF1 (N7736, N7725);
or OR2 (N7737, N7732, N1298);
nand NAND2 (N7738, N7736, N4238);
nand NAND2 (N7739, N7738, N6564);
xor XOR2 (N7740, N7727, N3957);
not NOT1 (N7741, N7729);
nand NAND3 (N7742, N7735, N7205, N2535);
not NOT1 (N7743, N7733);
xor XOR2 (N7744, N7724, N4535);
xor XOR2 (N7745, N7740, N7386);
or OR4 (N7746, N7739, N6458, N5335, N3610);
xor XOR2 (N7747, N7745, N1707);
or OR4 (N7748, N7741, N5606, N6736, N5516);
nand NAND2 (N7749, N7730, N1300);
buf BUF1 (N7750, N7737);
xor XOR2 (N7751, N7747, N2459);
nor NOR4 (N7752, N7731, N5679, N4856, N4745);
or OR2 (N7753, N7749, N4366);
or OR2 (N7754, N7748, N5379);
not NOT1 (N7755, N7734);
not NOT1 (N7756, N7752);
not NOT1 (N7757, N7742);
not NOT1 (N7758, N7746);
and AND4 (N7759, N7743, N4031, N865, N879);
xor XOR2 (N7760, N7759, N2241);
nor NOR3 (N7761, N7750, N1482, N5353);
buf BUF1 (N7762, N7753);
or OR2 (N7763, N7758, N4559);
xor XOR2 (N7764, N7763, N1471);
or OR4 (N7765, N7761, N6936, N3173, N4281);
not NOT1 (N7766, N7755);
xor XOR2 (N7767, N7766, N6460);
nor NOR3 (N7768, N7764, N6605, N5137);
not NOT1 (N7769, N7754);
and AND4 (N7770, N7767, N4895, N1489, N7530);
buf BUF1 (N7771, N7760);
not NOT1 (N7772, N7757);
xor XOR2 (N7773, N7751, N7466);
xor XOR2 (N7774, N7773, N4821);
not NOT1 (N7775, N7772);
xor XOR2 (N7776, N7769, N4416);
nand NAND4 (N7777, N7775, N397, N585, N6853);
or OR3 (N7778, N7744, N601, N2760);
xor XOR2 (N7779, N7770, N218);
xor XOR2 (N7780, N7762, N2444);
xor XOR2 (N7781, N7756, N4076);
nand NAND2 (N7782, N7774, N112);
nor NOR2 (N7783, N7771, N4557);
xor XOR2 (N7784, N7779, N6868);
or OR2 (N7785, N7783, N7720);
nand NAND3 (N7786, N7781, N6488, N5247);
or OR2 (N7787, N7768, N6332);
nand NAND2 (N7788, N7780, N4869);
or OR2 (N7789, N7778, N5593);
nor NOR2 (N7790, N7787, N1082);
xor XOR2 (N7791, N7785, N2475);
and AND3 (N7792, N7790, N4998, N6070);
or OR2 (N7793, N7786, N2934);
xor XOR2 (N7794, N7784, N452);
and AND3 (N7795, N7765, N2516, N126);
buf BUF1 (N7796, N7789);
buf BUF1 (N7797, N7793);
and AND3 (N7798, N7792, N4210, N7309);
xor XOR2 (N7799, N7795, N7596);
and AND2 (N7800, N7799, N4354);
xor XOR2 (N7801, N7776, N961);
buf BUF1 (N7802, N7801);
not NOT1 (N7803, N7794);
buf BUF1 (N7804, N7796);
nor NOR3 (N7805, N7791, N455, N1933);
nor NOR2 (N7806, N7798, N6610);
nor NOR4 (N7807, N7797, N1928, N1139, N5982);
buf BUF1 (N7808, N7806);
and AND2 (N7809, N7802, N3766);
xor XOR2 (N7810, N7809, N7663);
nor NOR4 (N7811, N7808, N2886, N2151, N4852);
and AND3 (N7812, N7782, N1535, N5023);
and AND4 (N7813, N7803, N6060, N296, N3306);
nand NAND4 (N7814, N7811, N1259, N1736, N6943);
not NOT1 (N7815, N7814);
nand NAND4 (N7816, N7777, N2373, N6128, N534);
buf BUF1 (N7817, N7788);
nand NAND2 (N7818, N7810, N71);
xor XOR2 (N7819, N7807, N5464);
buf BUF1 (N7820, N7818);
or OR2 (N7821, N7812, N6156);
not NOT1 (N7822, N7800);
xor XOR2 (N7823, N7816, N4525);
nand NAND4 (N7824, N7823, N4193, N3129, N564);
not NOT1 (N7825, N7804);
not NOT1 (N7826, N7815);
buf BUF1 (N7827, N7822);
buf BUF1 (N7828, N7825);
xor XOR2 (N7829, N7813, N1119);
nand NAND4 (N7830, N7821, N89, N4890, N3050);
and AND4 (N7831, N7820, N6623, N603, N6342);
buf BUF1 (N7832, N7819);
buf BUF1 (N7833, N7829);
nor NOR3 (N7834, N7827, N4667, N7120);
or OR4 (N7835, N7832, N5774, N3773, N3562);
not NOT1 (N7836, N7835);
xor XOR2 (N7837, N7836, N3439);
buf BUF1 (N7838, N7828);
nor NOR2 (N7839, N7837, N5660);
nand NAND3 (N7840, N7833, N2238, N3205);
or OR2 (N7841, N7834, N1196);
nand NAND3 (N7842, N7831, N7111, N3344);
or OR4 (N7843, N7824, N4744, N3628, N6426);
nand NAND2 (N7844, N7843, N5191);
nand NAND3 (N7845, N7840, N205, N3244);
or OR4 (N7846, N7845, N6336, N1194, N4966);
or OR4 (N7847, N7826, N4288, N1784, N6160);
and AND3 (N7848, N7805, N6980, N802);
nand NAND2 (N7849, N7847, N200);
nand NAND2 (N7850, N7817, N6149);
and AND4 (N7851, N7839, N199, N5200, N3176);
nor NOR2 (N7852, N7850, N4491);
xor XOR2 (N7853, N7849, N4920);
or OR2 (N7854, N7844, N1291);
nor NOR2 (N7855, N7848, N7525);
nand NAND4 (N7856, N7854, N1896, N5879, N4674);
and AND4 (N7857, N7846, N5514, N7544, N3021);
buf BUF1 (N7858, N7851);
and AND4 (N7859, N7853, N3765, N6685, N6272);
nor NOR4 (N7860, N7858, N1755, N125, N1389);
buf BUF1 (N7861, N7857);
xor XOR2 (N7862, N7856, N1015);
xor XOR2 (N7863, N7861, N7462);
or OR3 (N7864, N7859, N2493, N2396);
nand NAND2 (N7865, N7841, N5865);
or OR2 (N7866, N7863, N6418);
xor XOR2 (N7867, N7830, N4799);
or OR3 (N7868, N7866, N2393, N3119);
and AND4 (N7869, N7865, N6962, N1623, N5835);
and AND4 (N7870, N7838, N2669, N1277, N4122);
buf BUF1 (N7871, N7855);
xor XOR2 (N7872, N7842, N7415);
buf BUF1 (N7873, N7862);
xor XOR2 (N7874, N7864, N149);
and AND4 (N7875, N7868, N445, N7325, N1376);
not NOT1 (N7876, N7873);
nor NOR3 (N7877, N7876, N1987, N6386);
nor NOR2 (N7878, N7852, N4927);
not NOT1 (N7879, N7860);
not NOT1 (N7880, N7878);
nand NAND4 (N7881, N7872, N127, N6551, N5203);
buf BUF1 (N7882, N7870);
and AND3 (N7883, N7869, N7869, N2040);
and AND4 (N7884, N7879, N6516, N7539, N7169);
nand NAND2 (N7885, N7884, N408);
and AND3 (N7886, N7867, N206, N6604);
and AND4 (N7887, N7874, N1521, N3579, N7386);
buf BUF1 (N7888, N7871);
nor NOR3 (N7889, N7883, N7503, N7257);
nand NAND3 (N7890, N7886, N4086, N5908);
nand NAND2 (N7891, N7888, N3698);
and AND4 (N7892, N7891, N7156, N6207, N6242);
buf BUF1 (N7893, N7877);
nor NOR3 (N7894, N7875, N2210, N3230);
nor NOR3 (N7895, N7890, N7265, N111);
xor XOR2 (N7896, N7880, N1788);
buf BUF1 (N7897, N7896);
xor XOR2 (N7898, N7889, N7344);
buf BUF1 (N7899, N7882);
nand NAND2 (N7900, N7881, N1337);
buf BUF1 (N7901, N7887);
xor XOR2 (N7902, N7895, N7576);
nor NOR2 (N7903, N7897, N7814);
nor NOR4 (N7904, N7893, N3344, N5876, N6455);
buf BUF1 (N7905, N7902);
buf BUF1 (N7906, N7904);
buf BUF1 (N7907, N7903);
xor XOR2 (N7908, N7900, N2433);
xor XOR2 (N7909, N7905, N2237);
nor NOR2 (N7910, N7898, N6685);
not NOT1 (N7911, N7907);
or OR4 (N7912, N7909, N2296, N2032, N4960);
buf BUF1 (N7913, N7911);
not NOT1 (N7914, N7913);
buf BUF1 (N7915, N7901);
nand NAND4 (N7916, N7915, N342, N5562, N1727);
nor NOR4 (N7917, N7885, N2754, N1917, N3047);
or OR3 (N7918, N7906, N1966, N7813);
buf BUF1 (N7919, N7892);
or OR3 (N7920, N7912, N3080, N2277);
and AND4 (N7921, N7899, N558, N6487, N1982);
nand NAND4 (N7922, N7919, N3316, N6768, N933);
xor XOR2 (N7923, N7894, N2603);
nand NAND3 (N7924, N7916, N2303, N3798);
nand NAND3 (N7925, N7910, N7782, N1127);
nand NAND3 (N7926, N7917, N1588, N5640);
buf BUF1 (N7927, N7914);
or OR4 (N7928, N7922, N4226, N7778, N3097);
xor XOR2 (N7929, N7928, N3177);
and AND2 (N7930, N7926, N5871);
buf BUF1 (N7931, N7927);
or OR2 (N7932, N7929, N5486);
xor XOR2 (N7933, N7932, N3334);
xor XOR2 (N7934, N7923, N2176);
nor NOR2 (N7935, N7934, N4441);
xor XOR2 (N7936, N7921, N848);
nand NAND2 (N7937, N7933, N3673);
buf BUF1 (N7938, N7918);
nor NOR4 (N7939, N7935, N5620, N2534, N815);
nand NAND3 (N7940, N7930, N6389, N2068);
nand NAND4 (N7941, N7920, N742, N5258, N2389);
nand NAND4 (N7942, N7908, N7201, N47, N4880);
xor XOR2 (N7943, N7937, N6537);
or OR4 (N7944, N7924, N4430, N2610, N6494);
buf BUF1 (N7945, N7936);
nand NAND2 (N7946, N7945, N5134);
and AND2 (N7947, N7931, N3428);
and AND4 (N7948, N7939, N5988, N6651, N810);
and AND4 (N7949, N7946, N715, N7938, N6288);
not NOT1 (N7950, N6755);
xor XOR2 (N7951, N7947, N183);
nand NAND2 (N7952, N7940, N500);
nand NAND2 (N7953, N7942, N3912);
or OR2 (N7954, N7953, N395);
or OR2 (N7955, N7950, N2921);
xor XOR2 (N7956, N7949, N6779);
nor NOR3 (N7957, N7948, N3868, N3810);
or OR2 (N7958, N7925, N4804);
nand NAND4 (N7959, N7943, N4596, N6218, N4481);
and AND3 (N7960, N7951, N3802, N7448);
nor NOR3 (N7961, N7941, N2888, N2064);
nand NAND2 (N7962, N7955, N3259);
not NOT1 (N7963, N7956);
buf BUF1 (N7964, N7961);
nand NAND3 (N7965, N7954, N5217, N851);
or OR4 (N7966, N7963, N5257, N4360, N6594);
nor NOR2 (N7967, N7965, N5081);
buf BUF1 (N7968, N7957);
or OR2 (N7969, N7959, N2084);
nor NOR2 (N7970, N7966, N5561);
nand NAND4 (N7971, N7964, N3982, N2210, N2422);
nor NOR2 (N7972, N7969, N2935);
nor NOR2 (N7973, N7958, N3602);
nand NAND3 (N7974, N7971, N4082, N5518);
not NOT1 (N7975, N7960);
nand NAND4 (N7976, N7973, N291, N4387, N7557);
xor XOR2 (N7977, N7975, N6234);
buf BUF1 (N7978, N7976);
nor NOR3 (N7979, N7952, N2062, N6065);
nand NAND3 (N7980, N7978, N3307, N6436);
or OR2 (N7981, N7967, N5574);
nand NAND4 (N7982, N7970, N6181, N4343, N2573);
buf BUF1 (N7983, N7974);
buf BUF1 (N7984, N7980);
nor NOR3 (N7985, N7979, N2632, N418);
and AND4 (N7986, N7985, N146, N693, N7725);
buf BUF1 (N7987, N7984);
xor XOR2 (N7988, N7982, N6138);
not NOT1 (N7989, N7944);
xor XOR2 (N7990, N7968, N83);
nand NAND3 (N7991, N7977, N3555, N5360);
nand NAND2 (N7992, N7990, N7284);
nor NOR3 (N7993, N7991, N3303, N5981);
not NOT1 (N7994, N7986);
buf BUF1 (N7995, N7962);
or OR2 (N7996, N7989, N590);
and AND3 (N7997, N7992, N979, N6626);
buf BUF1 (N7998, N7997);
nor NOR2 (N7999, N7987, N3948);
nor NOR4 (N8000, N7981, N5389, N1729, N7109);
nor NOR2 (N8001, N8000, N7932);
not NOT1 (N8002, N7983);
and AND3 (N8003, N7995, N1355, N659);
and AND3 (N8004, N7988, N5049, N3489);
and AND4 (N8005, N7972, N997, N5907, N3641);
and AND2 (N8006, N7996, N7621);
nand NAND4 (N8007, N7993, N4251, N5427, N4276);
buf BUF1 (N8008, N7999);
nand NAND2 (N8009, N8007, N2247);
and AND2 (N8010, N8006, N3490);
nor NOR4 (N8011, N8004, N4541, N397, N7572);
xor XOR2 (N8012, N7998, N6506);
or OR3 (N8013, N8008, N6936, N5261);
nor NOR4 (N8014, N7994, N1932, N6012, N1998);
not NOT1 (N8015, N8013);
nor NOR4 (N8016, N8015, N5705, N597, N436);
nor NOR4 (N8017, N8012, N7689, N5142, N5105);
nand NAND3 (N8018, N8014, N6656, N266);
not NOT1 (N8019, N8001);
not NOT1 (N8020, N8017);
nor NOR2 (N8021, N8011, N7283);
not NOT1 (N8022, N8018);
not NOT1 (N8023, N8010);
xor XOR2 (N8024, N8020, N237);
not NOT1 (N8025, N8002);
and AND4 (N8026, N8005, N2205, N3163, N2739);
nor NOR2 (N8027, N8026, N6684);
nand NAND2 (N8028, N8016, N4162);
nand NAND3 (N8029, N8023, N1998, N7410);
not NOT1 (N8030, N8022);
buf BUF1 (N8031, N8027);
buf BUF1 (N8032, N8031);
buf BUF1 (N8033, N8003);
or OR3 (N8034, N8024, N7470, N3934);
xor XOR2 (N8035, N8033, N2925);
or OR4 (N8036, N8035, N7635, N1975, N4240);
nor NOR2 (N8037, N8032, N6515);
not NOT1 (N8038, N8025);
xor XOR2 (N8039, N8038, N2414);
or OR3 (N8040, N8029, N2505, N6360);
not NOT1 (N8041, N8019);
xor XOR2 (N8042, N8037, N4407);
not NOT1 (N8043, N8009);
xor XOR2 (N8044, N8039, N4845);
and AND4 (N8045, N8021, N4388, N1002, N1938);
xor XOR2 (N8046, N8043, N5080);
or OR2 (N8047, N8041, N1108);
nor NOR2 (N8048, N8046, N4500);
not NOT1 (N8049, N8040);
buf BUF1 (N8050, N8049);
xor XOR2 (N8051, N8047, N1713);
not NOT1 (N8052, N8034);
nand NAND2 (N8053, N8044, N4260);
nand NAND2 (N8054, N8028, N3625);
and AND4 (N8055, N8030, N5860, N2390, N4245);
nand NAND2 (N8056, N8054, N539);
xor XOR2 (N8057, N8036, N7735);
or OR3 (N8058, N8057, N1776, N2040);
and AND4 (N8059, N8052, N7885, N1310, N6767);
or OR2 (N8060, N8059, N6516);
and AND2 (N8061, N8045, N1476);
not NOT1 (N8062, N8058);
xor XOR2 (N8063, N8061, N3789);
buf BUF1 (N8064, N8055);
nor NOR2 (N8065, N8064, N5447);
nor NOR2 (N8066, N8060, N4524);
nor NOR2 (N8067, N8066, N4466);
nor NOR3 (N8068, N8053, N3982, N2202);
buf BUF1 (N8069, N8050);
not NOT1 (N8070, N8042);
or OR2 (N8071, N8063, N4368);
nor NOR4 (N8072, N8062, N1631, N7603, N458);
xor XOR2 (N8073, N8071, N5698);
nand NAND4 (N8074, N8051, N7524, N1731, N5113);
nor NOR2 (N8075, N8065, N7138);
or OR4 (N8076, N8069, N379, N3313, N5860);
nand NAND4 (N8077, N8048, N7481, N2678, N7155);
and AND2 (N8078, N8056, N2221);
and AND3 (N8079, N8077, N4541, N3083);
buf BUF1 (N8080, N8076);
nor NOR4 (N8081, N8073, N3133, N5410, N6858);
nor NOR3 (N8082, N8070, N2376, N2739);
not NOT1 (N8083, N8067);
nor NOR4 (N8084, N8083, N6481, N2272, N184);
buf BUF1 (N8085, N8075);
nand NAND4 (N8086, N8080, N4390, N6737, N808);
nand NAND2 (N8087, N8085, N2306);
xor XOR2 (N8088, N8079, N4973);
xor XOR2 (N8089, N8084, N6999);
and AND2 (N8090, N8086, N5256);
xor XOR2 (N8091, N8089, N2472);
buf BUF1 (N8092, N8078);
or OR3 (N8093, N8072, N7475, N5899);
and AND3 (N8094, N8074, N3710, N4971);
not NOT1 (N8095, N8087);
not NOT1 (N8096, N8088);
buf BUF1 (N8097, N8068);
or OR2 (N8098, N8095, N5456);
nor NOR2 (N8099, N8097, N5092);
and AND3 (N8100, N8091, N5565, N7230);
xor XOR2 (N8101, N8096, N6620);
xor XOR2 (N8102, N8081, N1771);
and AND4 (N8103, N8100, N4325, N1248, N969);
buf BUF1 (N8104, N8099);
xor XOR2 (N8105, N8102, N636);
xor XOR2 (N8106, N8105, N3478);
xor XOR2 (N8107, N8082, N7093);
xor XOR2 (N8108, N8107, N4911);
nand NAND4 (N8109, N8106, N7488, N856, N7869);
nor NOR3 (N8110, N8094, N8067, N3094);
nor NOR4 (N8111, N8104, N6832, N7668, N6053);
xor XOR2 (N8112, N8093, N1854);
nand NAND2 (N8113, N8090, N2666);
xor XOR2 (N8114, N8113, N6616);
xor XOR2 (N8115, N8098, N3929);
and AND2 (N8116, N8103, N503);
and AND3 (N8117, N8116, N2975, N1795);
xor XOR2 (N8118, N8117, N7126);
not NOT1 (N8119, N8112);
nor NOR4 (N8120, N8114, N1094, N3367, N3265);
buf BUF1 (N8121, N8115);
not NOT1 (N8122, N8092);
buf BUF1 (N8123, N8109);
nand NAND4 (N8124, N8120, N2073, N3584, N4414);
or OR4 (N8125, N8110, N1974, N4941, N3479);
xor XOR2 (N8126, N8119, N208);
not NOT1 (N8127, N8111);
and AND4 (N8128, N8127, N2864, N605, N7494);
nand NAND3 (N8129, N8128, N5015, N3780);
and AND4 (N8130, N8129, N1403, N6589, N2089);
not NOT1 (N8131, N8118);
not NOT1 (N8132, N8122);
xor XOR2 (N8133, N8132, N8015);
or OR3 (N8134, N8126, N1397, N5811);
buf BUF1 (N8135, N8134);
nor NOR4 (N8136, N8130, N2063, N5431, N1619);
nand NAND2 (N8137, N8123, N1294);
nor NOR4 (N8138, N8121, N3348, N4578, N4405);
nand NAND3 (N8139, N8133, N7597, N5141);
not NOT1 (N8140, N8124);
not NOT1 (N8141, N8125);
buf BUF1 (N8142, N8138);
not NOT1 (N8143, N8137);
xor XOR2 (N8144, N8136, N2155);
buf BUF1 (N8145, N8101);
nor NOR4 (N8146, N8141, N7151, N3946, N4553);
or OR2 (N8147, N8146, N7898);
or OR2 (N8148, N8143, N485);
not NOT1 (N8149, N8145);
and AND4 (N8150, N8139, N7524, N2645, N5838);
buf BUF1 (N8151, N8131);
not NOT1 (N8152, N8142);
buf BUF1 (N8153, N8149);
xor XOR2 (N8154, N8147, N2707);
nand NAND2 (N8155, N8153, N2157);
or OR2 (N8156, N8108, N1627);
and AND3 (N8157, N8154, N2463, N857);
and AND4 (N8158, N8135, N1473, N2717, N4502);
or OR2 (N8159, N8151, N7718);
xor XOR2 (N8160, N8140, N4400);
nor NOR2 (N8161, N8158, N5740);
not NOT1 (N8162, N8159);
xor XOR2 (N8163, N8157, N457);
xor XOR2 (N8164, N8163, N2862);
buf BUF1 (N8165, N8164);
xor XOR2 (N8166, N8160, N1724);
or OR2 (N8167, N8166, N1297);
not NOT1 (N8168, N8167);
buf BUF1 (N8169, N8161);
not NOT1 (N8170, N8165);
or OR3 (N8171, N8152, N941, N3140);
nor NOR2 (N8172, N8156, N468);
not NOT1 (N8173, N8148);
or OR4 (N8174, N8162, N5560, N2590, N604);
and AND4 (N8175, N8170, N5289, N7263, N1934);
xor XOR2 (N8176, N8172, N5667);
and AND2 (N8177, N8174, N2044);
buf BUF1 (N8178, N8150);
buf BUF1 (N8179, N8169);
or OR2 (N8180, N8173, N5806);
or OR2 (N8181, N8178, N5213);
xor XOR2 (N8182, N8144, N7684);
or OR3 (N8183, N8177, N563, N2844);
buf BUF1 (N8184, N8171);
nor NOR3 (N8185, N8181, N4336, N1493);
or OR3 (N8186, N8182, N3585, N3376);
and AND4 (N8187, N8186, N6707, N3812, N1916);
or OR3 (N8188, N8183, N2512, N7693);
not NOT1 (N8189, N8187);
buf BUF1 (N8190, N8188);
nand NAND2 (N8191, N8185, N516);
and AND3 (N8192, N8191, N6973, N5283);
buf BUF1 (N8193, N8190);
buf BUF1 (N8194, N8175);
nand NAND4 (N8195, N8180, N1421, N6141, N67);
and AND3 (N8196, N8184, N93, N7418);
xor XOR2 (N8197, N8193, N4823);
nand NAND3 (N8198, N8195, N598, N2342);
not NOT1 (N8199, N8194);
nand NAND4 (N8200, N8176, N6662, N4403, N556);
not NOT1 (N8201, N8199);
nor NOR4 (N8202, N8168, N7846, N1906, N7561);
nor NOR3 (N8203, N8189, N952, N4284);
and AND2 (N8204, N8179, N1041);
nor NOR2 (N8205, N8192, N6127);
nand NAND2 (N8206, N8198, N7854);
or OR4 (N8207, N8205, N4696, N3787, N7394);
nor NOR3 (N8208, N8196, N3438, N2028);
xor XOR2 (N8209, N8200, N821);
not NOT1 (N8210, N8204);
buf BUF1 (N8211, N8155);
not NOT1 (N8212, N8207);
buf BUF1 (N8213, N8209);
buf BUF1 (N8214, N8212);
and AND4 (N8215, N8206, N3567, N1728, N4330);
and AND2 (N8216, N8211, N5398);
not NOT1 (N8217, N8214);
nor NOR2 (N8218, N8208, N5139);
buf BUF1 (N8219, N8197);
buf BUF1 (N8220, N8203);
xor XOR2 (N8221, N8219, N3037);
buf BUF1 (N8222, N8201);
nand NAND2 (N8223, N8220, N4921);
or OR4 (N8224, N8216, N2309, N1382, N3798);
and AND2 (N8225, N8215, N5698);
nor NOR2 (N8226, N8218, N2813);
or OR2 (N8227, N8222, N6977);
and AND2 (N8228, N8224, N1468);
nand NAND3 (N8229, N8223, N3475, N1855);
not NOT1 (N8230, N8213);
not NOT1 (N8231, N8226);
not NOT1 (N8232, N8210);
buf BUF1 (N8233, N8230);
xor XOR2 (N8234, N8217, N2386);
nor NOR3 (N8235, N8225, N7322, N3866);
buf BUF1 (N8236, N8234);
or OR2 (N8237, N8231, N2823);
not NOT1 (N8238, N8236);
and AND4 (N8239, N8228, N4381, N4101, N4699);
or OR2 (N8240, N8202, N6943);
and AND3 (N8241, N8240, N2614, N5140);
xor XOR2 (N8242, N8227, N1368);
buf BUF1 (N8243, N8232);
or OR3 (N8244, N8237, N4968, N706);
nor NOR4 (N8245, N8238, N6777, N865, N7296);
xor XOR2 (N8246, N8244, N7527);
or OR2 (N8247, N8239, N1269);
buf BUF1 (N8248, N8233);
nand NAND3 (N8249, N8241, N6528, N1270);
or OR4 (N8250, N8221, N5859, N3807, N4585);
or OR4 (N8251, N8247, N6402, N3594, N6319);
or OR3 (N8252, N8248, N2345, N4758);
xor XOR2 (N8253, N8252, N1537);
xor XOR2 (N8254, N8245, N2818);
xor XOR2 (N8255, N8249, N2530);
xor XOR2 (N8256, N8243, N6898);
xor XOR2 (N8257, N8254, N4937);
nor NOR3 (N8258, N8255, N3484, N4465);
nand NAND4 (N8259, N8235, N6770, N5632, N4142);
or OR3 (N8260, N8257, N7571, N4604);
nor NOR3 (N8261, N8246, N4890, N7890);
buf BUF1 (N8262, N8258);
nor NOR2 (N8263, N8242, N3178);
nor NOR4 (N8264, N8253, N7290, N2452, N3661);
not NOT1 (N8265, N8263);
nand NAND4 (N8266, N8260, N2077, N4439, N5015);
or OR4 (N8267, N8259, N5825, N891, N7436);
buf BUF1 (N8268, N8250);
nand NAND4 (N8269, N8261, N6737, N6374, N5559);
and AND2 (N8270, N8256, N3459);
buf BUF1 (N8271, N8270);
not NOT1 (N8272, N8265);
or OR4 (N8273, N8269, N7826, N2462, N1328);
or OR4 (N8274, N8272, N5132, N3343, N800);
xor XOR2 (N8275, N8229, N2518);
buf BUF1 (N8276, N8273);
nor NOR2 (N8277, N8271, N2295);
or OR2 (N8278, N8276, N3315);
nor NOR3 (N8279, N8266, N7488, N4689);
nand NAND4 (N8280, N8262, N5649, N3991, N526);
nor NOR4 (N8281, N8264, N5094, N1784, N1487);
and AND3 (N8282, N8274, N215, N1614);
or OR3 (N8283, N8278, N2860, N112);
nand NAND4 (N8284, N8279, N4147, N5752, N5737);
xor XOR2 (N8285, N8283, N5619);
buf BUF1 (N8286, N8275);
or OR2 (N8287, N8281, N2403);
and AND2 (N8288, N8287, N2764);
not NOT1 (N8289, N8251);
xor XOR2 (N8290, N8282, N232);
and AND3 (N8291, N8286, N7772, N6273);
or OR2 (N8292, N8284, N904);
not NOT1 (N8293, N8289);
nand NAND4 (N8294, N8288, N698, N3862, N2607);
not NOT1 (N8295, N8280);
nand NAND2 (N8296, N8290, N279);
xor XOR2 (N8297, N8294, N3565);
nor NOR2 (N8298, N8291, N232);
nor NOR2 (N8299, N8277, N4635);
xor XOR2 (N8300, N8295, N8104);
xor XOR2 (N8301, N8298, N8242);
or OR3 (N8302, N8297, N4295, N3455);
or OR2 (N8303, N8292, N1497);
xor XOR2 (N8304, N8299, N7260);
or OR2 (N8305, N8268, N5606);
nand NAND4 (N8306, N8305, N60, N376, N6928);
nand NAND4 (N8307, N8296, N2906, N1900, N1257);
or OR3 (N8308, N8306, N7703, N7649);
and AND4 (N8309, N8308, N7836, N4735, N2922);
or OR4 (N8310, N8303, N1593, N4930, N7068);
and AND3 (N8311, N8301, N4924, N2684);
xor XOR2 (N8312, N8302, N7096);
buf BUF1 (N8313, N8304);
and AND4 (N8314, N8267, N2425, N8308, N3882);
buf BUF1 (N8315, N8300);
buf BUF1 (N8316, N8310);
nor NOR2 (N8317, N8312, N3744);
nand NAND2 (N8318, N8285, N6773);
buf BUF1 (N8319, N8309);
nand NAND3 (N8320, N8307, N6010, N7382);
or OR3 (N8321, N8318, N7974, N7258);
xor XOR2 (N8322, N8293, N5287);
nor NOR3 (N8323, N8315, N811, N2307);
and AND4 (N8324, N8320, N2168, N7862, N1697);
xor XOR2 (N8325, N8316, N4788);
xor XOR2 (N8326, N8313, N6539);
nand NAND2 (N8327, N8317, N606);
not NOT1 (N8328, N8326);
not NOT1 (N8329, N8327);
xor XOR2 (N8330, N8325, N4372);
or OR2 (N8331, N8324, N4396);
not NOT1 (N8332, N8322);
nor NOR2 (N8333, N8319, N7945);
buf BUF1 (N8334, N8328);
nor NOR3 (N8335, N8331, N1071, N6424);
not NOT1 (N8336, N8332);
or OR2 (N8337, N8333, N753);
xor XOR2 (N8338, N8337, N8109);
xor XOR2 (N8339, N8334, N1121);
nand NAND3 (N8340, N8323, N432, N4358);
nor NOR2 (N8341, N8338, N1175);
and AND4 (N8342, N8330, N541, N4159, N8238);
or OR3 (N8343, N8321, N2870, N4595);
not NOT1 (N8344, N8341);
buf BUF1 (N8345, N8342);
and AND4 (N8346, N8314, N1951, N5675, N1709);
nor NOR4 (N8347, N8339, N582, N4324, N3050);
nand NAND3 (N8348, N8311, N1070, N1175);
or OR2 (N8349, N8347, N7166);
nand NAND4 (N8350, N8340, N184, N5657, N709);
or OR2 (N8351, N8329, N6409);
xor XOR2 (N8352, N8343, N3780);
not NOT1 (N8353, N8344);
and AND2 (N8354, N8353, N7834);
nand NAND2 (N8355, N8346, N1904);
or OR2 (N8356, N8348, N3994);
or OR3 (N8357, N8355, N747, N5997);
nor NOR4 (N8358, N8336, N6641, N2561, N216);
nor NOR3 (N8359, N8335, N8048, N7757);
nand NAND2 (N8360, N8351, N5884);
nor NOR4 (N8361, N8345, N388, N6447, N3386);
nor NOR2 (N8362, N8357, N3703);
nor NOR3 (N8363, N8354, N3028, N2604);
xor XOR2 (N8364, N8356, N4965);
nor NOR2 (N8365, N8349, N187);
xor XOR2 (N8366, N8359, N574);
or OR3 (N8367, N8364, N2405, N5126);
and AND4 (N8368, N8365, N8138, N3654, N1810);
and AND2 (N8369, N8350, N873);
nand NAND3 (N8370, N8360, N7217, N2980);
or OR2 (N8371, N8352, N6100);
xor XOR2 (N8372, N8367, N6357);
and AND2 (N8373, N8366, N928);
not NOT1 (N8374, N8371);
or OR3 (N8375, N8361, N1958, N8182);
not NOT1 (N8376, N8370);
or OR4 (N8377, N8375, N1964, N1954, N296);
or OR3 (N8378, N8377, N2567, N771);
nor NOR3 (N8379, N8363, N1103, N3625);
xor XOR2 (N8380, N8373, N1477);
not NOT1 (N8381, N8378);
and AND2 (N8382, N8376, N7815);
or OR3 (N8383, N8358, N3995, N4832);
xor XOR2 (N8384, N8382, N2788);
or OR4 (N8385, N8384, N6163, N6470, N847);
and AND2 (N8386, N8372, N4241);
nor NOR4 (N8387, N8368, N7587, N2561, N3515);
nor NOR2 (N8388, N8381, N5343);
xor XOR2 (N8389, N8362, N2163);
buf BUF1 (N8390, N8386);
not NOT1 (N8391, N8369);
buf BUF1 (N8392, N8390);
buf BUF1 (N8393, N8379);
not NOT1 (N8394, N8393);
nor NOR2 (N8395, N8374, N5187);
nor NOR3 (N8396, N8392, N4018, N1028);
not NOT1 (N8397, N8396);
not NOT1 (N8398, N8391);
or OR3 (N8399, N8395, N3940, N570);
nand NAND2 (N8400, N8387, N3712);
not NOT1 (N8401, N8399);
xor XOR2 (N8402, N8401, N4337);
buf BUF1 (N8403, N8400);
or OR2 (N8404, N8397, N5890);
xor XOR2 (N8405, N8394, N5639);
buf BUF1 (N8406, N8403);
xor XOR2 (N8407, N8398, N3313);
xor XOR2 (N8408, N8405, N457);
or OR3 (N8409, N8380, N6120, N5832);
not NOT1 (N8410, N8389);
or OR3 (N8411, N8383, N6676, N7798);
buf BUF1 (N8412, N8411);
xor XOR2 (N8413, N8409, N4870);
and AND2 (N8414, N8404, N1610);
xor XOR2 (N8415, N8388, N3332);
nand NAND4 (N8416, N8408, N4261, N125, N5744);
buf BUF1 (N8417, N8413);
not NOT1 (N8418, N8406);
not NOT1 (N8419, N8417);
nand NAND3 (N8420, N8416, N8271, N7663);
nand NAND4 (N8421, N8419, N7445, N5092, N4561);
nor NOR3 (N8422, N8421, N6032, N5803);
nand NAND2 (N8423, N8414, N1205);
or OR2 (N8424, N8402, N965);
nor NOR3 (N8425, N8385, N3703, N7198);
buf BUF1 (N8426, N8422);
xor XOR2 (N8427, N8426, N4853);
nor NOR2 (N8428, N8425, N8204);
or OR4 (N8429, N8427, N4820, N1033, N602);
or OR4 (N8430, N8428, N7612, N4537, N941);
nor NOR3 (N8431, N8410, N7640, N7387);
not NOT1 (N8432, N8415);
nor NOR4 (N8433, N8412, N1078, N3619, N1438);
nor NOR2 (N8434, N8423, N6532);
not NOT1 (N8435, N8424);
buf BUF1 (N8436, N8418);
or OR2 (N8437, N8429, N3199);
not NOT1 (N8438, N8430);
not NOT1 (N8439, N8436);
nor NOR4 (N8440, N8431, N1124, N3807, N4932);
nand NAND4 (N8441, N8407, N6235, N1609, N4873);
not NOT1 (N8442, N8438);
or OR2 (N8443, N8442, N626);
nor NOR2 (N8444, N8420, N2857);
and AND4 (N8445, N8433, N8184, N3449, N1391);
xor XOR2 (N8446, N8444, N914);
xor XOR2 (N8447, N8446, N4292);
nor NOR3 (N8448, N8445, N1413, N7994);
nand NAND4 (N8449, N8437, N7131, N2355, N4952);
or OR2 (N8450, N8448, N766);
buf BUF1 (N8451, N8447);
nor NOR2 (N8452, N8451, N228);
xor XOR2 (N8453, N8452, N1696);
nor NOR4 (N8454, N8435, N248, N1747, N4507);
not NOT1 (N8455, N8439);
not NOT1 (N8456, N8450);
nor NOR3 (N8457, N8453, N1273, N4856);
and AND3 (N8458, N8440, N1165, N1471);
and AND2 (N8459, N8455, N5334);
xor XOR2 (N8460, N8459, N3755);
nand NAND3 (N8461, N8449, N4056, N4356);
xor XOR2 (N8462, N8456, N1048);
not NOT1 (N8463, N8458);
and AND2 (N8464, N8461, N2661);
not NOT1 (N8465, N8464);
xor XOR2 (N8466, N8465, N2053);
and AND2 (N8467, N8441, N2638);
xor XOR2 (N8468, N8434, N807);
or OR2 (N8469, N8454, N1550);
not NOT1 (N8470, N8462);
nor NOR2 (N8471, N8460, N8419);
nand NAND2 (N8472, N8470, N3218);
nand NAND3 (N8473, N8463, N3421, N5391);
xor XOR2 (N8474, N8471, N1714);
or OR4 (N8475, N8466, N197, N7561, N4033);
nor NOR4 (N8476, N8469, N38, N7160, N629);
buf BUF1 (N8477, N8474);
not NOT1 (N8478, N8443);
nand NAND4 (N8479, N8468, N7678, N5959, N5663);
or OR4 (N8480, N8457, N108, N5646, N5416);
xor XOR2 (N8481, N8478, N3185);
xor XOR2 (N8482, N8467, N5153);
not NOT1 (N8483, N8473);
nor NOR3 (N8484, N8472, N3924, N3133);
and AND3 (N8485, N8483, N3696, N1770);
and AND2 (N8486, N8480, N5805);
nand NAND3 (N8487, N8479, N8098, N7676);
buf BUF1 (N8488, N8486);
nor NOR4 (N8489, N8488, N7841, N1485, N5497);
or OR4 (N8490, N8485, N2718, N7501, N5471);
or OR4 (N8491, N8477, N80, N5697, N1306);
nor NOR3 (N8492, N8481, N1006, N2939);
nor NOR2 (N8493, N8476, N3702);
not NOT1 (N8494, N8493);
or OR3 (N8495, N8491, N2729, N4214);
nand NAND2 (N8496, N8432, N3929);
nand NAND4 (N8497, N8492, N7926, N6192, N3607);
and AND3 (N8498, N8497, N4091, N8398);
buf BUF1 (N8499, N8490);
or OR3 (N8500, N8489, N7076, N224);
and AND4 (N8501, N8500, N1003, N1436, N4651);
and AND2 (N8502, N8484, N3896);
and AND2 (N8503, N8499, N6633);
xor XOR2 (N8504, N8482, N6691);
nand NAND4 (N8505, N8496, N2529, N7026, N2577);
and AND3 (N8506, N8501, N421, N8150);
nand NAND3 (N8507, N8502, N6642, N5635);
not NOT1 (N8508, N8495);
nand NAND2 (N8509, N8494, N7554);
nor NOR3 (N8510, N8507, N1047, N151);
nor NOR2 (N8511, N8503, N1550);
not NOT1 (N8512, N8506);
and AND3 (N8513, N8504, N4274, N4685);
nor NOR3 (N8514, N8510, N682, N3101);
nor NOR3 (N8515, N8505, N5999, N8010);
buf BUF1 (N8516, N8487);
and AND2 (N8517, N8512, N6234);
nor NOR2 (N8518, N8511, N3145);
or OR4 (N8519, N8516, N402, N1375, N582);
buf BUF1 (N8520, N8514);
nor NOR4 (N8521, N8498, N5137, N5214, N319);
xor XOR2 (N8522, N8509, N2490);
nor NOR3 (N8523, N8518, N5968, N5070);
nor NOR4 (N8524, N8508, N7047, N5062, N7738);
nor NOR3 (N8525, N8523, N4152, N6591);
and AND2 (N8526, N8524, N7624);
buf BUF1 (N8527, N8519);
nor NOR4 (N8528, N8513, N6650, N7060, N4623);
xor XOR2 (N8529, N8522, N4167);
or OR3 (N8530, N8528, N5018, N3611);
and AND3 (N8531, N8527, N2269, N927);
nand NAND3 (N8532, N8530, N1393, N8381);
nand NAND3 (N8533, N8475, N7185, N6049);
xor XOR2 (N8534, N8521, N7163);
and AND2 (N8535, N8515, N942);
or OR3 (N8536, N8529, N3175, N3791);
not NOT1 (N8537, N8535);
nor NOR4 (N8538, N8525, N282, N5973, N5501);
nand NAND3 (N8539, N8532, N2312, N1464);
nand NAND2 (N8540, N8538, N709);
buf BUF1 (N8541, N8517);
not NOT1 (N8542, N8536);
nor NOR3 (N8543, N8537, N5829, N7140);
and AND2 (N8544, N8526, N1212);
and AND4 (N8545, N8539, N227, N4327, N5568);
xor XOR2 (N8546, N8543, N8156);
or OR4 (N8547, N8520, N2735, N7627, N2019);
not NOT1 (N8548, N8546);
and AND3 (N8549, N8540, N4380, N6148);
nand NAND4 (N8550, N8541, N4845, N1269, N2592);
or OR2 (N8551, N8531, N2259);
not NOT1 (N8552, N8547);
xor XOR2 (N8553, N8534, N4121);
not NOT1 (N8554, N8549);
or OR2 (N8555, N8554, N5787);
buf BUF1 (N8556, N8555);
or OR4 (N8557, N8556, N386, N6828, N7732);
xor XOR2 (N8558, N8544, N2265);
not NOT1 (N8559, N8557);
not NOT1 (N8560, N8552);
and AND2 (N8561, N8551, N5344);
nand NAND2 (N8562, N8560, N861);
buf BUF1 (N8563, N8553);
xor XOR2 (N8564, N8561, N7463);
not NOT1 (N8565, N8548);
and AND4 (N8566, N8564, N4821, N131, N5544);
xor XOR2 (N8567, N8566, N6357);
xor XOR2 (N8568, N8559, N1644);
xor XOR2 (N8569, N8558, N2827);
nor NOR3 (N8570, N8533, N2157, N837);
and AND2 (N8571, N8568, N1638);
nor NOR2 (N8572, N8542, N1750);
buf BUF1 (N8573, N8563);
and AND3 (N8574, N8550, N6756, N257);
nor NOR2 (N8575, N8567, N6299);
or OR2 (N8576, N8545, N5017);
not NOT1 (N8577, N8572);
nand NAND2 (N8578, N8574, N6009);
nor NOR2 (N8579, N8575, N7297);
xor XOR2 (N8580, N8565, N2221);
buf BUF1 (N8581, N8580);
nor NOR3 (N8582, N8581, N7030, N4341);
buf BUF1 (N8583, N8570);
nand NAND3 (N8584, N8576, N6033, N5724);
nand NAND2 (N8585, N8584, N7583);
not NOT1 (N8586, N8573);
nand NAND2 (N8587, N8577, N7149);
xor XOR2 (N8588, N8571, N8436);
not NOT1 (N8589, N8569);
buf BUF1 (N8590, N8562);
nand NAND3 (N8591, N8583, N6619, N2666);
xor XOR2 (N8592, N8587, N4064);
xor XOR2 (N8593, N8582, N1428);
not NOT1 (N8594, N8578);
not NOT1 (N8595, N8594);
nor NOR2 (N8596, N8589, N8515);
nand NAND3 (N8597, N8590, N2660, N1932);
and AND3 (N8598, N8579, N3103, N5275);
xor XOR2 (N8599, N8588, N2218);
nand NAND4 (N8600, N8595, N2689, N7156, N6716);
nand NAND4 (N8601, N8600, N7571, N5436, N7241);
buf BUF1 (N8602, N8596);
nand NAND2 (N8603, N8597, N5576);
and AND2 (N8604, N8586, N2829);
not NOT1 (N8605, N8601);
or OR3 (N8606, N8598, N7883, N671);
nor NOR4 (N8607, N8593, N3818, N4092, N3357);
not NOT1 (N8608, N8604);
nor NOR3 (N8609, N8602, N7121, N349);
nand NAND3 (N8610, N8603, N7708, N7261);
and AND3 (N8611, N8599, N5841, N425);
xor XOR2 (N8612, N8610, N5497);
nand NAND4 (N8613, N8608, N5148, N1949, N1500);
or OR3 (N8614, N8606, N7254, N1289);
not NOT1 (N8615, N8585);
or OR2 (N8616, N8613, N4746);
nand NAND4 (N8617, N8592, N5445, N3478, N6568);
xor XOR2 (N8618, N8611, N4581);
or OR3 (N8619, N8618, N8141, N7707);
nand NAND4 (N8620, N8614, N5884, N5675, N6818);
or OR3 (N8621, N8609, N6852, N2887);
xor XOR2 (N8622, N8617, N3802);
buf BUF1 (N8623, N8612);
buf BUF1 (N8624, N8615);
and AND2 (N8625, N8607, N6882);
or OR3 (N8626, N8625, N2865, N5022);
or OR4 (N8627, N8619, N5325, N479, N2700);
buf BUF1 (N8628, N8621);
not NOT1 (N8629, N8591);
or OR3 (N8630, N8626, N596, N5232);
or OR3 (N8631, N8630, N2319, N303);
nor NOR4 (N8632, N8620, N8167, N7705, N4403);
nor NOR3 (N8633, N8624, N2782, N3489);
or OR3 (N8634, N8616, N6711, N293);
or OR2 (N8635, N8627, N756);
and AND3 (N8636, N8605, N2730, N994);
and AND3 (N8637, N8631, N8039, N5844);
nor NOR2 (N8638, N8629, N803);
and AND4 (N8639, N8622, N6174, N5292, N4419);
not NOT1 (N8640, N8633);
xor XOR2 (N8641, N8634, N280);
nor NOR4 (N8642, N8637, N594, N1701, N1552);
nand NAND2 (N8643, N8639, N1469);
nor NOR4 (N8644, N8638, N4609, N731, N5864);
buf BUF1 (N8645, N8643);
or OR3 (N8646, N8636, N2179, N393);
or OR2 (N8647, N8644, N4745);
or OR4 (N8648, N8645, N4268, N3587, N4791);
nand NAND4 (N8649, N8641, N6504, N1497, N1724);
nor NOR3 (N8650, N8642, N6482, N6639);
xor XOR2 (N8651, N8632, N1675);
nand NAND2 (N8652, N8635, N6675);
not NOT1 (N8653, N8651);
or OR2 (N8654, N8653, N1739);
buf BUF1 (N8655, N8646);
not NOT1 (N8656, N8628);
nand NAND2 (N8657, N8647, N383);
xor XOR2 (N8658, N8652, N6771);
not NOT1 (N8659, N8656);
or OR4 (N8660, N8659, N2733, N3828, N8394);
nor NOR2 (N8661, N8660, N8407);
not NOT1 (N8662, N8648);
buf BUF1 (N8663, N8661);
nand NAND4 (N8664, N8650, N4361, N1162, N8436);
or OR2 (N8665, N8654, N3583);
nor NOR4 (N8666, N8665, N4529, N7810, N4245);
xor XOR2 (N8667, N8655, N6);
nor NOR4 (N8668, N8658, N5003, N2684, N5859);
and AND3 (N8669, N8649, N6109, N8353);
nor NOR4 (N8670, N8664, N6275, N5922, N48);
xor XOR2 (N8671, N8669, N3104);
or OR2 (N8672, N8623, N2613);
nand NAND4 (N8673, N8662, N1310, N4238, N8516);
nor NOR4 (N8674, N8668, N4090, N2817, N1978);
and AND2 (N8675, N8667, N5099);
buf BUF1 (N8676, N8640);
or OR3 (N8677, N8671, N5598, N3987);
not NOT1 (N8678, N8670);
nand NAND4 (N8679, N8666, N1077, N4919, N8159);
nor NOR3 (N8680, N8677, N6058, N3084);
not NOT1 (N8681, N8678);
buf BUF1 (N8682, N8663);
xor XOR2 (N8683, N8681, N5476);
and AND3 (N8684, N8672, N6928, N743);
nand NAND3 (N8685, N8676, N8160, N6525);
nor NOR4 (N8686, N8683, N5944, N3893, N73);
not NOT1 (N8687, N8679);
nand NAND4 (N8688, N8674, N4605, N4261, N5979);
xor XOR2 (N8689, N8680, N3798);
buf BUF1 (N8690, N8685);
nand NAND3 (N8691, N8684, N3034, N1362);
nor NOR2 (N8692, N8690, N3253);
nand NAND2 (N8693, N8692, N6400);
or OR2 (N8694, N8675, N2476);
or OR2 (N8695, N8682, N1816);
or OR2 (N8696, N8695, N4463);
and AND4 (N8697, N8694, N1675, N3054, N6586);
xor XOR2 (N8698, N8673, N1998);
buf BUF1 (N8699, N8698);
and AND4 (N8700, N8689, N7896, N1834, N4931);
nand NAND2 (N8701, N8693, N6156);
nand NAND3 (N8702, N8686, N8519, N4016);
not NOT1 (N8703, N8696);
not NOT1 (N8704, N8688);
and AND3 (N8705, N8657, N5389, N3722);
buf BUF1 (N8706, N8697);
or OR4 (N8707, N8700, N741, N1623, N1349);
buf BUF1 (N8708, N8687);
buf BUF1 (N8709, N8703);
nand NAND4 (N8710, N8702, N7996, N2269, N3422);
nor NOR4 (N8711, N8707, N5817, N6191, N7607);
nor NOR4 (N8712, N8710, N6608, N7912, N5581);
and AND2 (N8713, N8711, N6448);
and AND3 (N8714, N8706, N6451, N8209);
or OR3 (N8715, N8699, N7680, N3906);
buf BUF1 (N8716, N8712);
or OR4 (N8717, N8709, N1814, N7767, N6991);
buf BUF1 (N8718, N8714);
buf BUF1 (N8719, N8691);
not NOT1 (N8720, N8719);
xor XOR2 (N8721, N8705, N4027);
or OR4 (N8722, N8717, N3301, N6217, N7717);
not NOT1 (N8723, N8718);
nor NOR4 (N8724, N8720, N5694, N6848, N2875);
or OR4 (N8725, N8721, N7500, N3606, N2154);
nor NOR2 (N8726, N8715, N8441);
and AND3 (N8727, N8701, N7321, N6832);
or OR3 (N8728, N8724, N5329, N853);
not NOT1 (N8729, N8713);
and AND2 (N8730, N8708, N7115);
not NOT1 (N8731, N8723);
and AND2 (N8732, N8722, N7241);
nor NOR2 (N8733, N8729, N5712);
nand NAND2 (N8734, N8732, N2611);
nand NAND3 (N8735, N8731, N7071, N4477);
xor XOR2 (N8736, N8727, N8340);
not NOT1 (N8737, N8704);
nand NAND3 (N8738, N8726, N8451, N1138);
buf BUF1 (N8739, N8730);
nor NOR3 (N8740, N8733, N3638, N7293);
xor XOR2 (N8741, N8740, N4719);
nor NOR2 (N8742, N8741, N4120);
and AND2 (N8743, N8739, N635);
nor NOR4 (N8744, N8728, N387, N2117, N1992);
not NOT1 (N8745, N8743);
or OR3 (N8746, N8735, N5598, N6897);
nor NOR3 (N8747, N8744, N4714, N5962);
not NOT1 (N8748, N8746);
xor XOR2 (N8749, N8738, N4317);
nand NAND4 (N8750, N8748, N3126, N5436, N4143);
nand NAND3 (N8751, N8734, N3261, N1285);
xor XOR2 (N8752, N8745, N4247);
and AND2 (N8753, N8716, N2733);
or OR2 (N8754, N8747, N6320);
xor XOR2 (N8755, N8753, N2264);
or OR3 (N8756, N8752, N3067, N8506);
nand NAND4 (N8757, N8742, N6100, N6527, N7759);
nor NOR2 (N8758, N8754, N8090);
or OR4 (N8759, N8756, N425, N8735, N1933);
not NOT1 (N8760, N8751);
xor XOR2 (N8761, N8749, N4197);
nor NOR4 (N8762, N8736, N6186, N7151, N1258);
and AND2 (N8763, N8755, N104);
or OR3 (N8764, N8762, N4769, N5120);
nand NAND3 (N8765, N8737, N3987, N5792);
and AND4 (N8766, N8758, N1772, N5047, N1197);
and AND4 (N8767, N8766, N4990, N5875, N3133);
nand NAND4 (N8768, N8759, N6910, N2921, N1067);
nand NAND4 (N8769, N8757, N2089, N4869, N5503);
buf BUF1 (N8770, N8769);
nand NAND2 (N8771, N8764, N875);
and AND3 (N8772, N8750, N6886, N5916);
nand NAND2 (N8773, N8763, N1058);
buf BUF1 (N8774, N8773);
or OR2 (N8775, N8725, N1691);
buf BUF1 (N8776, N8775);
nand NAND2 (N8777, N8776, N5160);
nand NAND4 (N8778, N8772, N717, N3664, N2395);
nor NOR3 (N8779, N8774, N5168, N7268);
and AND4 (N8780, N8777, N197, N3475, N6745);
xor XOR2 (N8781, N8770, N6812);
and AND2 (N8782, N8767, N8609);
buf BUF1 (N8783, N8780);
or OR2 (N8784, N8779, N7519);
and AND3 (N8785, N8784, N1872, N2701);
not NOT1 (N8786, N8765);
xor XOR2 (N8787, N8760, N8625);
nor NOR4 (N8788, N8768, N903, N6132, N900);
not NOT1 (N8789, N8781);
nor NOR3 (N8790, N8787, N606, N1317);
nand NAND3 (N8791, N8782, N5908, N1454);
or OR3 (N8792, N8786, N7221, N8702);
nand NAND3 (N8793, N8790, N5945, N3858);
xor XOR2 (N8794, N8771, N5438);
nor NOR3 (N8795, N8778, N6503, N2646);
nor NOR3 (N8796, N8794, N3671, N2781);
or OR3 (N8797, N8788, N5953, N7136);
nand NAND3 (N8798, N8796, N3220, N3119);
xor XOR2 (N8799, N8795, N7796);
xor XOR2 (N8800, N8785, N2345);
xor XOR2 (N8801, N8798, N2456);
nand NAND2 (N8802, N8792, N7876);
nand NAND4 (N8803, N8791, N3484, N1132, N1702);
nand NAND2 (N8804, N8803, N7002);
not NOT1 (N8805, N8804);
nand NAND3 (N8806, N8805, N4664, N337);
buf BUF1 (N8807, N8793);
nand NAND2 (N8808, N8783, N1476);
buf BUF1 (N8809, N8808);
and AND3 (N8810, N8807, N2861, N352);
buf BUF1 (N8811, N8789);
buf BUF1 (N8812, N8802);
xor XOR2 (N8813, N8811, N4153);
buf BUF1 (N8814, N8810);
or OR2 (N8815, N8761, N4006);
not NOT1 (N8816, N8812);
and AND2 (N8817, N8816, N456);
and AND3 (N8818, N8813, N5203, N4777);
and AND4 (N8819, N8799, N4098, N1957, N8090);
and AND3 (N8820, N8819, N3038, N4249);
buf BUF1 (N8821, N8806);
nand NAND2 (N8822, N8821, N3307);
nand NAND3 (N8823, N8801, N8002, N4700);
nand NAND4 (N8824, N8809, N6689, N3320, N6135);
not NOT1 (N8825, N8823);
nand NAND4 (N8826, N8820, N3965, N497, N2743);
nor NOR4 (N8827, N8824, N2226, N4882, N3695);
not NOT1 (N8828, N8817);
nand NAND2 (N8829, N8814, N5809);
or OR2 (N8830, N8822, N3526);
and AND4 (N8831, N8797, N5059, N268, N5827);
or OR3 (N8832, N8826, N8332, N4723);
nand NAND4 (N8833, N8830, N1099, N6981, N6501);
nand NAND4 (N8834, N8818, N25, N5737, N220);
and AND4 (N8835, N8800, N1689, N1158, N8597);
not NOT1 (N8836, N8832);
buf BUF1 (N8837, N8829);
buf BUF1 (N8838, N8831);
or OR2 (N8839, N8827, N1990);
and AND2 (N8840, N8833, N3266);
not NOT1 (N8841, N8839);
nor NOR3 (N8842, N8837, N6071, N569);
not NOT1 (N8843, N8825);
nand NAND4 (N8844, N8815, N5832, N580, N8025);
nand NAND2 (N8845, N8844, N6353);
and AND4 (N8846, N8836, N4903, N636, N5808);
nand NAND3 (N8847, N8841, N8342, N3501);
and AND2 (N8848, N8840, N7592);
not NOT1 (N8849, N8847);
nor NOR2 (N8850, N8845, N6028);
nand NAND3 (N8851, N8850, N6109, N7068);
or OR4 (N8852, N8828, N3307, N1427, N8164);
not NOT1 (N8853, N8834);
or OR3 (N8854, N8852, N3491, N7393);
xor XOR2 (N8855, N8835, N4528);
xor XOR2 (N8856, N8842, N3433);
not NOT1 (N8857, N8843);
nor NOR2 (N8858, N8853, N4698);
nor NOR3 (N8859, N8855, N1882, N4036);
nor NOR4 (N8860, N8854, N1594, N428, N2848);
buf BUF1 (N8861, N8846);
xor XOR2 (N8862, N8858, N2818);
nand NAND3 (N8863, N8851, N7298, N2142);
buf BUF1 (N8864, N8848);
xor XOR2 (N8865, N8859, N8051);
nor NOR3 (N8866, N8857, N2785, N6951);
nand NAND3 (N8867, N8861, N6313, N475);
nand NAND2 (N8868, N8864, N4522);
and AND2 (N8869, N8866, N5082);
buf BUF1 (N8870, N8867);
buf BUF1 (N8871, N8838);
buf BUF1 (N8872, N8862);
and AND4 (N8873, N8860, N6106, N6797, N7534);
buf BUF1 (N8874, N8873);
nand NAND4 (N8875, N8874, N2388, N1439, N3099);
not NOT1 (N8876, N8856);
nor NOR2 (N8877, N8875, N4656);
nor NOR3 (N8878, N8870, N8248, N8249);
nand NAND4 (N8879, N8865, N3416, N2269, N1742);
or OR2 (N8880, N8879, N7232);
nand NAND2 (N8881, N8869, N1173);
not NOT1 (N8882, N8881);
nor NOR3 (N8883, N8880, N5822, N2734);
buf BUF1 (N8884, N8876);
buf BUF1 (N8885, N8871);
not NOT1 (N8886, N8878);
not NOT1 (N8887, N8868);
not NOT1 (N8888, N8849);
and AND3 (N8889, N8884, N3609, N4625);
not NOT1 (N8890, N8883);
nor NOR4 (N8891, N8886, N8075, N325, N1424);
not NOT1 (N8892, N8885);
nor NOR3 (N8893, N8891, N343, N1774);
nand NAND4 (N8894, N8887, N4408, N8685, N1134);
not NOT1 (N8895, N8890);
and AND2 (N8896, N8893, N5265);
or OR3 (N8897, N8888, N5953, N5208);
buf BUF1 (N8898, N8894);
and AND2 (N8899, N8895, N53);
nand NAND3 (N8900, N8872, N7368, N4265);
or OR3 (N8901, N8863, N2089, N2906);
xor XOR2 (N8902, N8889, N5888);
and AND2 (N8903, N8900, N7531);
nand NAND3 (N8904, N8901, N6198, N5368);
nor NOR2 (N8905, N8902, N8201);
xor XOR2 (N8906, N8905, N8216);
nand NAND3 (N8907, N8892, N1742, N4737);
nor NOR4 (N8908, N8906, N3457, N24, N565);
not NOT1 (N8909, N8907);
nor NOR3 (N8910, N8897, N7052, N2530);
xor XOR2 (N8911, N8898, N6798);
and AND3 (N8912, N8899, N4795, N5380);
xor XOR2 (N8913, N8912, N6189);
nand NAND2 (N8914, N8908, N5509);
or OR2 (N8915, N8877, N710);
not NOT1 (N8916, N8911);
xor XOR2 (N8917, N8903, N5572);
xor XOR2 (N8918, N8909, N4383);
nand NAND2 (N8919, N8910, N5559);
buf BUF1 (N8920, N8917);
not NOT1 (N8921, N8904);
buf BUF1 (N8922, N8921);
and AND3 (N8923, N8913, N6593, N5279);
buf BUF1 (N8924, N8916);
not NOT1 (N8925, N8924);
or OR4 (N8926, N8920, N2644, N7852, N2194);
xor XOR2 (N8927, N8914, N4000);
or OR3 (N8928, N8915, N6634, N7087);
buf BUF1 (N8929, N8922);
xor XOR2 (N8930, N8927, N4222);
not NOT1 (N8931, N8925);
and AND3 (N8932, N8882, N116, N447);
xor XOR2 (N8933, N8928, N3445);
and AND4 (N8934, N8918, N4574, N8436, N6370);
or OR4 (N8935, N8934, N2829, N6689, N5475);
and AND2 (N8936, N8931, N1469);
nor NOR2 (N8937, N8936, N53);
not NOT1 (N8938, N8937);
not NOT1 (N8939, N8933);
nand NAND3 (N8940, N8939, N96, N3618);
xor XOR2 (N8941, N8929, N6602);
and AND3 (N8942, N8941, N4538, N4994);
nand NAND4 (N8943, N8940, N7532, N2259, N2335);
and AND2 (N8944, N8930, N7921);
and AND4 (N8945, N8944, N4271, N4536, N7140);
buf BUF1 (N8946, N8932);
xor XOR2 (N8947, N8896, N6803);
nand NAND4 (N8948, N8935, N1945, N2, N3030);
buf BUF1 (N8949, N8948);
nor NOR4 (N8950, N8946, N2684, N4053, N1205);
buf BUF1 (N8951, N8942);
not NOT1 (N8952, N8938);
not NOT1 (N8953, N8919);
nor NOR2 (N8954, N8952, N7239);
or OR3 (N8955, N8923, N5310, N2316);
nor NOR2 (N8956, N8943, N8764);
or OR2 (N8957, N8950, N5299);
or OR2 (N8958, N8951, N4348);
and AND4 (N8959, N8957, N8201, N8697, N514);
nor NOR4 (N8960, N8947, N3474, N1667, N5278);
and AND4 (N8961, N8958, N4183, N441, N377);
not NOT1 (N8962, N8959);
not NOT1 (N8963, N8960);
nand NAND3 (N8964, N8955, N3725, N3705);
nand NAND4 (N8965, N8945, N3855, N636, N832);
xor XOR2 (N8966, N8961, N8692);
nand NAND2 (N8967, N8963, N8686);
nand NAND4 (N8968, N8953, N744, N7698, N2532);
or OR3 (N8969, N8967, N1793, N1780);
and AND3 (N8970, N8956, N4843, N3489);
buf BUF1 (N8971, N8968);
xor XOR2 (N8972, N8962, N5342);
and AND2 (N8973, N8965, N7908);
and AND3 (N8974, N8964, N1712, N8649);
or OR4 (N8975, N8969, N594, N8867, N4953);
nand NAND3 (N8976, N8975, N2872, N7256);
buf BUF1 (N8977, N8949);
nand NAND2 (N8978, N8976, N6305);
not NOT1 (N8979, N8973);
buf BUF1 (N8980, N8979);
nand NAND4 (N8981, N8966, N1985, N8611, N1013);
xor XOR2 (N8982, N8977, N4203);
nor NOR3 (N8983, N8982, N5515, N6204);
not NOT1 (N8984, N8971);
or OR2 (N8985, N8974, N8545);
not NOT1 (N8986, N8954);
nand NAND2 (N8987, N8985, N2452);
and AND4 (N8988, N8980, N7474, N7853, N403);
or OR2 (N8989, N8972, N3144);
buf BUF1 (N8990, N8981);
and AND4 (N8991, N8986, N3524, N2155, N1517);
xor XOR2 (N8992, N8988, N3760);
and AND3 (N8993, N8983, N4948, N5274);
buf BUF1 (N8994, N8926);
buf BUF1 (N8995, N8970);
nor NOR2 (N8996, N8990, N6251);
not NOT1 (N8997, N8995);
buf BUF1 (N8998, N8978);
nand NAND3 (N8999, N8984, N1717, N7226);
buf BUF1 (N9000, N8997);
nor NOR4 (N9001, N8989, N2324, N2919, N1677);
or OR2 (N9002, N9001, N7341);
or OR2 (N9003, N8996, N4998);
buf BUF1 (N9004, N8993);
and AND2 (N9005, N9002, N4318);
xor XOR2 (N9006, N9000, N6652);
nor NOR4 (N9007, N8999, N1402, N3452, N3345);
nor NOR4 (N9008, N8991, N5343, N6845, N2895);
or OR2 (N9009, N9008, N348);
or OR2 (N9010, N9009, N262);
xor XOR2 (N9011, N9007, N2645);
and AND4 (N9012, N8994, N7161, N4547, N8425);
nor NOR3 (N9013, N9003, N1093, N2311);
nor NOR2 (N9014, N9004, N5015);
not NOT1 (N9015, N9010);
xor XOR2 (N9016, N9015, N2176);
xor XOR2 (N9017, N9005, N3693);
not NOT1 (N9018, N9017);
and AND3 (N9019, N9012, N1888, N5705);
not NOT1 (N9020, N9016);
nand NAND4 (N9021, N8998, N2518, N1069, N1888);
not NOT1 (N9022, N9020);
and AND3 (N9023, N9006, N8336, N8438);
buf BUF1 (N9024, N9013);
nand NAND4 (N9025, N9014, N8546, N719, N1145);
nor NOR3 (N9026, N9023, N6488, N1223);
nand NAND3 (N9027, N9011, N5037, N3711);
buf BUF1 (N9028, N9027);
and AND4 (N9029, N9028, N5509, N7252, N8174);
xor XOR2 (N9030, N8992, N1010);
buf BUF1 (N9031, N9018);
and AND4 (N9032, N9030, N1296, N3219, N6829);
nand NAND4 (N9033, N9022, N7576, N2194, N8462);
not NOT1 (N9034, N9025);
nand NAND3 (N9035, N9024, N7152, N5471);
or OR3 (N9036, N9033, N5805, N2795);
xor XOR2 (N9037, N9031, N7174);
not NOT1 (N9038, N8987);
and AND3 (N9039, N9038, N5259, N2850);
not NOT1 (N9040, N9019);
not NOT1 (N9041, N9021);
nor NOR2 (N9042, N9037, N6822);
nor NOR4 (N9043, N9035, N5210, N8185, N556);
buf BUF1 (N9044, N9029);
or OR2 (N9045, N9034, N5943);
or OR3 (N9046, N9045, N478, N6697);
nor NOR4 (N9047, N9044, N1778, N6333, N4812);
nor NOR3 (N9048, N9042, N1146, N1213);
not NOT1 (N9049, N9026);
buf BUF1 (N9050, N9040);
buf BUF1 (N9051, N9050);
buf BUF1 (N9052, N9047);
or OR3 (N9053, N9041, N1860, N1907);
nand NAND2 (N9054, N9046, N296);
not NOT1 (N9055, N9032);
not NOT1 (N9056, N9052);
xor XOR2 (N9057, N9051, N7321);
nand NAND2 (N9058, N9054, N4519);
buf BUF1 (N9059, N9056);
nor NOR4 (N9060, N9048, N5212, N7575, N3957);
not NOT1 (N9061, N9049);
or OR2 (N9062, N9055, N8891);
nor NOR4 (N9063, N9043, N4948, N4557, N4732);
or OR3 (N9064, N9058, N6308, N7825);
and AND4 (N9065, N9036, N2417, N2559, N5289);
and AND4 (N9066, N9064, N1544, N8775, N8920);
or OR4 (N9067, N9063, N4190, N2552, N338);
buf BUF1 (N9068, N9057);
buf BUF1 (N9069, N9060);
nand NAND2 (N9070, N9065, N502);
or OR2 (N9071, N9039, N5882);
or OR4 (N9072, N9053, N7642, N406, N7671);
or OR4 (N9073, N9059, N7380, N5640, N4678);
nand NAND3 (N9074, N9070, N4892, N4346);
xor XOR2 (N9075, N9072, N8091);
nor NOR3 (N9076, N9074, N4381, N8079);
xor XOR2 (N9077, N9062, N5463);
and AND4 (N9078, N9071, N5088, N2748, N8341);
nand NAND3 (N9079, N9077, N264, N5088);
nor NOR2 (N9080, N9068, N6053);
buf BUF1 (N9081, N9073);
xor XOR2 (N9082, N9075, N7549);
or OR4 (N9083, N9076, N2561, N7337, N2831);
nor NOR4 (N9084, N9069, N422, N7615, N6509);
nand NAND4 (N9085, N9081, N5431, N2407, N1330);
xor XOR2 (N9086, N9082, N8652);
nor NOR3 (N9087, N9085, N1641, N2347);
and AND3 (N9088, N9083, N5411, N3987);
not NOT1 (N9089, N9084);
nor NOR3 (N9090, N9078, N217, N6602);
buf BUF1 (N9091, N9061);
nor NOR3 (N9092, N9067, N4559, N3650);
nand NAND4 (N9093, N9087, N6482, N1373, N8306);
nand NAND3 (N9094, N9093, N3876, N338);
nor NOR3 (N9095, N9092, N8151, N7435);
nor NOR3 (N9096, N9094, N2646, N4073);
or OR3 (N9097, N9095, N2376, N5284);
or OR2 (N9098, N9090, N6011);
not NOT1 (N9099, N9079);
nand NAND2 (N9100, N9089, N8434);
nor NOR3 (N9101, N9086, N1540, N2130);
and AND2 (N9102, N9097, N5247);
not NOT1 (N9103, N9091);
or OR4 (N9104, N9102, N7412, N7717, N4111);
nand NAND3 (N9105, N9080, N3016, N8122);
or OR2 (N9106, N9104, N6936);
xor XOR2 (N9107, N9066, N7043);
xor XOR2 (N9108, N9099, N7351);
not NOT1 (N9109, N9101);
nor NOR2 (N9110, N9105, N6420);
buf BUF1 (N9111, N9108);
and AND2 (N9112, N9088, N741);
xor XOR2 (N9113, N9103, N5163);
or OR4 (N9114, N9107, N8635, N7275, N7305);
nor NOR2 (N9115, N9096, N2244);
nor NOR4 (N9116, N9115, N55, N6236, N1437);
xor XOR2 (N9117, N9113, N4885);
not NOT1 (N9118, N9106);
buf BUF1 (N9119, N9116);
nor NOR2 (N9120, N9114, N8218);
nand NAND2 (N9121, N9100, N115);
or OR2 (N9122, N9117, N5567);
or OR3 (N9123, N9119, N7542, N523);
nand NAND4 (N9124, N9122, N4755, N3014, N7300);
buf BUF1 (N9125, N9109);
nor NOR3 (N9126, N9112, N2955, N3451);
nand NAND4 (N9127, N9118, N716, N2519, N8121);
nand NAND3 (N9128, N9123, N974, N7721);
not NOT1 (N9129, N9124);
or OR4 (N9130, N9125, N5686, N2129, N5038);
xor XOR2 (N9131, N9121, N3830);
nand NAND2 (N9132, N9126, N2414);
xor XOR2 (N9133, N9132, N8087);
buf BUF1 (N9134, N9129);
xor XOR2 (N9135, N9131, N3070);
xor XOR2 (N9136, N9133, N95);
nand NAND4 (N9137, N9127, N3948, N6258, N5585);
xor XOR2 (N9138, N9110, N4613);
xor XOR2 (N9139, N9120, N6868);
nand NAND2 (N9140, N9098, N2673);
nand NAND2 (N9141, N9136, N8744);
buf BUF1 (N9142, N9141);
nor NOR4 (N9143, N9134, N5570, N5008, N1108);
not NOT1 (N9144, N9111);
not NOT1 (N9145, N9143);
nor NOR4 (N9146, N9145, N707, N5752, N6929);
nor NOR3 (N9147, N9137, N2528, N4216);
nor NOR2 (N9148, N9142, N3650);
nand NAND4 (N9149, N9130, N4663, N1718, N3002);
nor NOR2 (N9150, N9138, N1008);
buf BUF1 (N9151, N9139);
nand NAND2 (N9152, N9148, N1795);
xor XOR2 (N9153, N9149, N4140);
and AND4 (N9154, N9140, N4347, N3565, N1458);
not NOT1 (N9155, N9146);
not NOT1 (N9156, N9152);
nand NAND2 (N9157, N9147, N8130);
buf BUF1 (N9158, N9144);
and AND3 (N9159, N9153, N4272, N26);
buf BUF1 (N9160, N9155);
buf BUF1 (N9161, N9151);
xor XOR2 (N9162, N9159, N3262);
and AND4 (N9163, N9157, N8839, N8933, N650);
xor XOR2 (N9164, N9158, N3275);
not NOT1 (N9165, N9150);
nand NAND4 (N9166, N9156, N3141, N4261, N4680);
xor XOR2 (N9167, N9160, N6399);
nor NOR2 (N9168, N9165, N2309);
nor NOR3 (N9169, N9168, N712, N902);
xor XOR2 (N9170, N9128, N1359);
and AND3 (N9171, N9154, N8235, N1382);
buf BUF1 (N9172, N9164);
or OR2 (N9173, N9166, N6754);
or OR4 (N9174, N9170, N6889, N3289, N2032);
xor XOR2 (N9175, N9161, N7165);
buf BUF1 (N9176, N9169);
nand NAND2 (N9177, N9172, N1242);
or OR3 (N9178, N9176, N8653, N8736);
not NOT1 (N9179, N9171);
nand NAND3 (N9180, N9177, N1125, N4610);
not NOT1 (N9181, N9167);
and AND4 (N9182, N9162, N485, N2544, N1124);
xor XOR2 (N9183, N9163, N365);
and AND4 (N9184, N9179, N7192, N8071, N8778);
xor XOR2 (N9185, N9173, N3587);
xor XOR2 (N9186, N9175, N5135);
xor XOR2 (N9187, N9182, N878);
or OR3 (N9188, N9135, N8841, N1327);
buf BUF1 (N9189, N9180);
buf BUF1 (N9190, N9188);
not NOT1 (N9191, N9184);
nor NOR3 (N9192, N9189, N2348, N2897);
not NOT1 (N9193, N9185);
buf BUF1 (N9194, N9190);
xor XOR2 (N9195, N9174, N4139);
or OR2 (N9196, N9191, N8538);
or OR4 (N9197, N9181, N5970, N8899, N17);
and AND2 (N9198, N9193, N7573);
buf BUF1 (N9199, N9198);
nand NAND4 (N9200, N9196, N7519, N8576, N7212);
xor XOR2 (N9201, N9194, N747);
or OR2 (N9202, N9186, N636);
not NOT1 (N9203, N9200);
nand NAND3 (N9204, N9199, N5802, N5747);
xor XOR2 (N9205, N9192, N517);
and AND3 (N9206, N9187, N3270, N1245);
not NOT1 (N9207, N9183);
nor NOR2 (N9208, N9205, N3829);
nand NAND4 (N9209, N9207, N3186, N1715, N4280);
nand NAND3 (N9210, N9209, N4931, N3598);
not NOT1 (N9211, N9202);
xor XOR2 (N9212, N9201, N125);
nand NAND2 (N9213, N9204, N7147);
nor NOR3 (N9214, N9208, N7273, N6214);
buf BUF1 (N9215, N9213);
xor XOR2 (N9216, N9212, N668);
not NOT1 (N9217, N9215);
buf BUF1 (N9218, N9197);
xor XOR2 (N9219, N9211, N9185);
or OR3 (N9220, N9217, N8863, N6021);
not NOT1 (N9221, N9206);
nand NAND3 (N9222, N9216, N4212, N7662);
not NOT1 (N9223, N9195);
and AND2 (N9224, N9220, N8195);
buf BUF1 (N9225, N9210);
nor NOR3 (N9226, N9178, N5936, N4955);
nand NAND3 (N9227, N9218, N1986, N2186);
and AND2 (N9228, N9223, N4793);
not NOT1 (N9229, N9219);
xor XOR2 (N9230, N9229, N4903);
nand NAND2 (N9231, N9228, N6718);
and AND2 (N9232, N9226, N6257);
xor XOR2 (N9233, N9222, N4593);
xor XOR2 (N9234, N9203, N3951);
xor XOR2 (N9235, N9234, N1970);
and AND2 (N9236, N9232, N6957);
nor NOR4 (N9237, N9230, N4544, N7865, N5082);
nand NAND3 (N9238, N9214, N7424, N4693);
and AND4 (N9239, N9224, N4782, N8882, N7725);
buf BUF1 (N9240, N9238);
nor NOR4 (N9241, N9225, N4495, N1325, N2702);
not NOT1 (N9242, N9237);
buf BUF1 (N9243, N9231);
and AND3 (N9244, N9235, N6340, N1626);
not NOT1 (N9245, N9242);
nand NAND4 (N9246, N9221, N6025, N135, N5257);
nor NOR3 (N9247, N9243, N4912, N4668);
xor XOR2 (N9248, N9241, N8601);
buf BUF1 (N9249, N9239);
xor XOR2 (N9250, N9245, N6264);
xor XOR2 (N9251, N9250, N2731);
and AND3 (N9252, N9240, N6998, N3963);
not NOT1 (N9253, N9244);
buf BUF1 (N9254, N9248);
nor NOR4 (N9255, N9252, N293, N6917, N6324);
or OR3 (N9256, N9254, N5277, N5169);
not NOT1 (N9257, N9236);
not NOT1 (N9258, N9255);
not NOT1 (N9259, N9256);
buf BUF1 (N9260, N9227);
nand NAND3 (N9261, N9253, N5515, N8254);
and AND2 (N9262, N9261, N3012);
xor XOR2 (N9263, N9262, N4042);
nand NAND4 (N9264, N9246, N4614, N6936, N8779);
nor NOR4 (N9265, N9260, N6182, N8203, N554);
nand NAND3 (N9266, N9264, N1142, N6081);
not NOT1 (N9267, N9251);
not NOT1 (N9268, N9265);
xor XOR2 (N9269, N9247, N6855);
nand NAND4 (N9270, N9267, N5444, N4198, N2335);
xor XOR2 (N9271, N9269, N4807);
xor XOR2 (N9272, N9259, N257);
not NOT1 (N9273, N9258);
nor NOR3 (N9274, N9249, N5575, N3170);
nor NOR2 (N9275, N9274, N8549);
nand NAND2 (N9276, N9272, N2334);
xor XOR2 (N9277, N9266, N2237);
nand NAND2 (N9278, N9233, N915);
and AND2 (N9279, N9257, N7255);
nand NAND3 (N9280, N9279, N7614, N7785);
or OR4 (N9281, N9268, N3018, N499, N4622);
not NOT1 (N9282, N9275);
buf BUF1 (N9283, N9280);
nand NAND4 (N9284, N9263, N8412, N3008, N1811);
xor XOR2 (N9285, N9270, N4575);
or OR3 (N9286, N9276, N2192, N824);
nand NAND3 (N9287, N9273, N4837, N9067);
xor XOR2 (N9288, N9271, N4994);
not NOT1 (N9289, N9281);
xor XOR2 (N9290, N9277, N7199);
nand NAND2 (N9291, N9289, N92);
not NOT1 (N9292, N9288);
or OR3 (N9293, N9283, N2433, N5234);
or OR3 (N9294, N9290, N6825, N2129);
nor NOR4 (N9295, N9287, N1339, N6673, N8476);
or OR2 (N9296, N9285, N7442);
xor XOR2 (N9297, N9278, N3659);
nand NAND3 (N9298, N9296, N1, N3311);
xor XOR2 (N9299, N9291, N8068);
buf BUF1 (N9300, N9295);
xor XOR2 (N9301, N9282, N2987);
buf BUF1 (N9302, N9297);
nor NOR4 (N9303, N9302, N1724, N2336, N3030);
not NOT1 (N9304, N9294);
or OR4 (N9305, N9300, N8990, N5276, N7767);
not NOT1 (N9306, N9286);
nand NAND4 (N9307, N9303, N6607, N2320, N302);
and AND2 (N9308, N9304, N1022);
nand NAND2 (N9309, N9306, N584);
buf BUF1 (N9310, N9284);
or OR4 (N9311, N9299, N6523, N6118, N3106);
nand NAND2 (N9312, N9298, N9082);
not NOT1 (N9313, N9305);
and AND4 (N9314, N9312, N7393, N390, N992);
xor XOR2 (N9315, N9310, N6209);
xor XOR2 (N9316, N9309, N8297);
nor NOR3 (N9317, N9316, N6984, N5229);
nand NAND3 (N9318, N9293, N7259, N6102);
or OR4 (N9319, N9292, N6886, N4735, N1428);
and AND3 (N9320, N9311, N5128, N6772);
xor XOR2 (N9321, N9317, N5357);
and AND3 (N9322, N9315, N6658, N9009);
not NOT1 (N9323, N9321);
or OR4 (N9324, N9314, N4836, N5646, N5734);
not NOT1 (N9325, N9320);
or OR3 (N9326, N9301, N1907, N5186);
or OR3 (N9327, N9326, N8023, N6827);
and AND3 (N9328, N9308, N4746, N7668);
and AND2 (N9329, N9313, N6276);
nor NOR4 (N9330, N9325, N8030, N6666, N7439);
not NOT1 (N9331, N9328);
and AND4 (N9332, N9319, N3941, N7398, N8167);
nor NOR3 (N9333, N9324, N2040, N3165);
buf BUF1 (N9334, N9318);
buf BUF1 (N9335, N9322);
and AND2 (N9336, N9329, N1589);
and AND2 (N9337, N9336, N9187);
or OR2 (N9338, N9331, N6525);
xor XOR2 (N9339, N9335, N186);
nand NAND3 (N9340, N9330, N6772, N95);
nand NAND4 (N9341, N9332, N551, N5517, N1399);
buf BUF1 (N9342, N9340);
nor NOR3 (N9343, N9342, N5621, N638);
nand NAND4 (N9344, N9337, N8467, N1818, N4729);
not NOT1 (N9345, N9344);
and AND3 (N9346, N9333, N8028, N6086);
buf BUF1 (N9347, N9334);
buf BUF1 (N9348, N9345);
xor XOR2 (N9349, N9346, N2054);
nand NAND2 (N9350, N9338, N3999);
and AND2 (N9351, N9348, N6212);
nor NOR2 (N9352, N9351, N1742);
buf BUF1 (N9353, N9341);
and AND3 (N9354, N9347, N8150, N6775);
buf BUF1 (N9355, N9349);
not NOT1 (N9356, N9352);
buf BUF1 (N9357, N9327);
nor NOR3 (N9358, N9355, N5428, N5447);
nand NAND4 (N9359, N9307, N2060, N734, N5064);
not NOT1 (N9360, N9358);
buf BUF1 (N9361, N9343);
and AND3 (N9362, N9354, N4489, N9234);
nand NAND3 (N9363, N9350, N6162, N8893);
or OR4 (N9364, N9353, N5394, N2294, N4435);
xor XOR2 (N9365, N9360, N4481);
buf BUF1 (N9366, N9365);
xor XOR2 (N9367, N9366, N5161);
xor XOR2 (N9368, N9367, N492);
nor NOR3 (N9369, N9356, N8636, N4179);
buf BUF1 (N9370, N9362);
xor XOR2 (N9371, N9323, N5205);
nor NOR2 (N9372, N9359, N1325);
not NOT1 (N9373, N9372);
not NOT1 (N9374, N9373);
xor XOR2 (N9375, N9374, N901);
not NOT1 (N9376, N9357);
nand NAND2 (N9377, N9363, N4804);
buf BUF1 (N9378, N9339);
xor XOR2 (N9379, N9371, N8126);
nand NAND3 (N9380, N9361, N2919, N9123);
nand NAND3 (N9381, N9377, N5576, N7342);
nor NOR4 (N9382, N9376, N916, N5406, N6542);
buf BUF1 (N9383, N9368);
xor XOR2 (N9384, N9381, N4358);
nor NOR3 (N9385, N9375, N8366, N8219);
xor XOR2 (N9386, N9378, N1906);
or OR4 (N9387, N9386, N5186, N7165, N783);
not NOT1 (N9388, N9380);
or OR2 (N9389, N9385, N5037);
and AND2 (N9390, N9388, N9279);
and AND4 (N9391, N9387, N292, N1484, N3059);
nand NAND4 (N9392, N9390, N1360, N544, N6360);
not NOT1 (N9393, N9392);
not NOT1 (N9394, N9369);
buf BUF1 (N9395, N9364);
and AND2 (N9396, N9383, N7928);
and AND2 (N9397, N9394, N1339);
nand NAND2 (N9398, N9397, N5699);
buf BUF1 (N9399, N9396);
xor XOR2 (N9400, N9379, N4077);
nor NOR4 (N9401, N9382, N4954, N2764, N968);
nand NAND2 (N9402, N9395, N841);
nor NOR3 (N9403, N9389, N730, N3666);
not NOT1 (N9404, N9401);
buf BUF1 (N9405, N9404);
nand NAND4 (N9406, N9391, N622, N5532, N602);
xor XOR2 (N9407, N9406, N1552);
or OR4 (N9408, N9403, N3241, N1257, N4288);
buf BUF1 (N9409, N9407);
nand NAND4 (N9410, N9409, N3384, N3341, N6778);
nand NAND3 (N9411, N9370, N3882, N7211);
nor NOR2 (N9412, N9411, N5508);
and AND3 (N9413, N9410, N2429, N7134);
xor XOR2 (N9414, N9393, N3334);
not NOT1 (N9415, N9412);
or OR4 (N9416, N9405, N5839, N8051, N1786);
xor XOR2 (N9417, N9416, N4997);
and AND2 (N9418, N9417, N3554);
buf BUF1 (N9419, N9415);
nor NOR4 (N9420, N9419, N3501, N3747, N3861);
nand NAND2 (N9421, N9420, N1192);
buf BUF1 (N9422, N9418);
and AND4 (N9423, N9421, N8704, N2627, N4430);
or OR4 (N9424, N9398, N1869, N5465, N7346);
or OR3 (N9425, N9400, N8081, N6753);
xor XOR2 (N9426, N9422, N3979);
nor NOR4 (N9427, N9384, N740, N1081, N5470);
and AND3 (N9428, N9426, N9091, N1855);
buf BUF1 (N9429, N9399);
buf BUF1 (N9430, N9427);
not NOT1 (N9431, N9423);
not NOT1 (N9432, N9430);
nor NOR2 (N9433, N9425, N4282);
not NOT1 (N9434, N9433);
xor XOR2 (N9435, N9434, N1241);
nor NOR2 (N9436, N9435, N2315);
not NOT1 (N9437, N9414);
and AND2 (N9438, N9424, N6299);
and AND2 (N9439, N9438, N6112);
not NOT1 (N9440, N9413);
buf BUF1 (N9441, N9408);
buf BUF1 (N9442, N9432);
nor NOR2 (N9443, N9442, N7943);
or OR3 (N9444, N9429, N6015, N4479);
xor XOR2 (N9445, N9402, N8057);
buf BUF1 (N9446, N9445);
buf BUF1 (N9447, N9443);
or OR3 (N9448, N9428, N3311, N8320);
nor NOR2 (N9449, N9440, N8885);
buf BUF1 (N9450, N9436);
nor NOR3 (N9451, N9449, N9012, N6024);
xor XOR2 (N9452, N9451, N2700);
xor XOR2 (N9453, N9448, N3765);
not NOT1 (N9454, N9452);
nor NOR2 (N9455, N9431, N8273);
or OR2 (N9456, N9447, N5537);
nand NAND4 (N9457, N9439, N4951, N4179, N6622);
nand NAND2 (N9458, N9454, N3416);
nor NOR4 (N9459, N9446, N7035, N2751, N4782);
nor NOR3 (N9460, N9453, N1629, N3228);
not NOT1 (N9461, N9459);
nand NAND3 (N9462, N9457, N3194, N8635);
nand NAND4 (N9463, N9458, N6697, N5988, N8916);
nand NAND3 (N9464, N9455, N7698, N5513);
or OR2 (N9465, N9444, N7425);
nor NOR3 (N9466, N9437, N6292, N2240);
and AND3 (N9467, N9462, N3516, N845);
buf BUF1 (N9468, N9467);
xor XOR2 (N9469, N9450, N5408);
not NOT1 (N9470, N9468);
and AND4 (N9471, N9461, N4294, N5951, N6593);
or OR2 (N9472, N9465, N8628);
xor XOR2 (N9473, N9441, N1948);
not NOT1 (N9474, N9473);
and AND2 (N9475, N9466, N630);
nand NAND3 (N9476, N9464, N5352, N7896);
not NOT1 (N9477, N9475);
nand NAND2 (N9478, N9476, N4339);
nor NOR3 (N9479, N9469, N5507, N3702);
or OR3 (N9480, N9463, N3795, N3519);
and AND4 (N9481, N9471, N424, N6411, N2636);
nand NAND2 (N9482, N9460, N7426);
buf BUF1 (N9483, N9474);
xor XOR2 (N9484, N9482, N1891);
nand NAND2 (N9485, N9456, N9293);
nand NAND3 (N9486, N9472, N1545, N7675);
and AND2 (N9487, N9479, N7816);
xor XOR2 (N9488, N9470, N5862);
xor XOR2 (N9489, N9485, N7895);
nand NAND2 (N9490, N9483, N2872);
xor XOR2 (N9491, N9486, N5427);
nor NOR4 (N9492, N9480, N3359, N1070, N2349);
or OR4 (N9493, N9484, N7872, N7496, N7285);
and AND2 (N9494, N9491, N8141);
and AND4 (N9495, N9487, N6140, N8866, N5922);
xor XOR2 (N9496, N9494, N2526);
buf BUF1 (N9497, N9477);
buf BUF1 (N9498, N9497);
nand NAND3 (N9499, N9490, N1404, N1148);
buf BUF1 (N9500, N9495);
not NOT1 (N9501, N9500);
nor NOR2 (N9502, N9489, N4897);
not NOT1 (N9503, N9493);
nand NAND4 (N9504, N9498, N7056, N5155, N6074);
nor NOR4 (N9505, N9501, N3849, N345, N5201);
or OR2 (N9506, N9492, N3088);
and AND2 (N9507, N9478, N6737);
buf BUF1 (N9508, N9488);
buf BUF1 (N9509, N9504);
buf BUF1 (N9510, N9496);
buf BUF1 (N9511, N9502);
buf BUF1 (N9512, N9481);
not NOT1 (N9513, N9511);
or OR3 (N9514, N9508, N4841, N7950);
buf BUF1 (N9515, N9505);
buf BUF1 (N9516, N9509);
xor XOR2 (N9517, N9499, N5608);
xor XOR2 (N9518, N9512, N5835);
nand NAND4 (N9519, N9513, N8806, N3276, N921);
nand NAND3 (N9520, N9519, N1787, N4157);
nor NOR4 (N9521, N9517, N9373, N8145, N3897);
nor NOR3 (N9522, N9506, N6810, N2636);
xor XOR2 (N9523, N9522, N9369);
and AND2 (N9524, N9523, N3894);
or OR3 (N9525, N9503, N8548, N4728);
and AND4 (N9526, N9525, N328, N6102, N9249);
nor NOR3 (N9527, N9516, N3348, N5969);
nand NAND3 (N9528, N9510, N1882, N7398);
nand NAND2 (N9529, N9527, N8513);
buf BUF1 (N9530, N9524);
nor NOR3 (N9531, N9520, N8114, N3710);
and AND3 (N9532, N9507, N3496, N505);
nor NOR3 (N9533, N9530, N7130, N3482);
buf BUF1 (N9534, N9529);
not NOT1 (N9535, N9531);
and AND4 (N9536, N9514, N5952, N6601, N4512);
and AND3 (N9537, N9533, N4159, N2009);
and AND4 (N9538, N9528, N2094, N4171, N3324);
or OR3 (N9539, N9537, N4501, N2449);
not NOT1 (N9540, N9535);
nor NOR2 (N9541, N9532, N4565);
buf BUF1 (N9542, N9521);
buf BUF1 (N9543, N9539);
not NOT1 (N9544, N9540);
or OR3 (N9545, N9526, N6589, N7986);
nand NAND2 (N9546, N9536, N8397);
nor NOR4 (N9547, N9543, N9304, N5530, N1365);
and AND2 (N9548, N9546, N9535);
not NOT1 (N9549, N9541);
and AND2 (N9550, N9534, N6254);
or OR2 (N9551, N9549, N2814);
buf BUF1 (N9552, N9544);
and AND4 (N9553, N9542, N7241, N7887, N7726);
buf BUF1 (N9554, N9547);
or OR3 (N9555, N9554, N2344, N39);
nand NAND3 (N9556, N9550, N619, N5278);
and AND4 (N9557, N9552, N5438, N5917, N7838);
and AND3 (N9558, N9551, N8954, N1180);
and AND2 (N9559, N9538, N7618);
not NOT1 (N9560, N9518);
nor NOR4 (N9561, N9557, N4502, N3257, N1995);
not NOT1 (N9562, N9558);
nor NOR2 (N9563, N9559, N3075);
nand NAND4 (N9564, N9561, N8231, N2413, N1133);
and AND4 (N9565, N9560, N7224, N641, N5320);
not NOT1 (N9566, N9553);
xor XOR2 (N9567, N9556, N2565);
and AND3 (N9568, N9515, N4590, N7146);
nor NOR3 (N9569, N9562, N2466, N8707);
not NOT1 (N9570, N9568);
not NOT1 (N9571, N9548);
or OR2 (N9572, N9571, N3564);
xor XOR2 (N9573, N9563, N1142);
xor XOR2 (N9574, N9570, N5175);
not NOT1 (N9575, N9572);
xor XOR2 (N9576, N9574, N1044);
nor NOR2 (N9577, N9566, N720);
or OR4 (N9578, N9577, N4415, N2818, N30);
or OR4 (N9579, N9564, N6533, N7416, N5730);
and AND3 (N9580, N9565, N8822, N6054);
xor XOR2 (N9581, N9575, N8600);
not NOT1 (N9582, N9569);
nor NOR3 (N9583, N9573, N6997, N1024);
nand NAND4 (N9584, N9579, N3187, N7987, N2279);
xor XOR2 (N9585, N9582, N519);
xor XOR2 (N9586, N9584, N4189);
nand NAND3 (N9587, N9578, N4671, N6031);
or OR4 (N9588, N9545, N3501, N7806, N3124);
or OR4 (N9589, N9583, N604, N8050, N720);
buf BUF1 (N9590, N9586);
not NOT1 (N9591, N9555);
buf BUF1 (N9592, N9567);
nor NOR3 (N9593, N9587, N2176, N8468);
buf BUF1 (N9594, N9592);
nor NOR4 (N9595, N9581, N8077, N4648, N2516);
nor NOR2 (N9596, N9593, N360);
and AND3 (N9597, N9580, N7095, N4469);
buf BUF1 (N9598, N9589);
nand NAND2 (N9599, N9585, N7280);
or OR4 (N9600, N9597, N7074, N6154, N5963);
or OR2 (N9601, N9599, N3863);
nand NAND3 (N9602, N9590, N3424, N138);
nand NAND2 (N9603, N9588, N7131);
nand NAND2 (N9604, N9603, N3775);
or OR4 (N9605, N9602, N5593, N30, N8108);
and AND2 (N9606, N9595, N4799);
and AND2 (N9607, N9604, N2429);
nor NOR2 (N9608, N9601, N6619);
and AND3 (N9609, N9600, N1618, N3772);
nor NOR4 (N9610, N9598, N6342, N5496, N4117);
buf BUF1 (N9611, N9576);
and AND2 (N9612, N9611, N2164);
nor NOR4 (N9613, N9610, N8261, N1368, N7679);
or OR3 (N9614, N9606, N2617, N3799);
buf BUF1 (N9615, N9607);
and AND2 (N9616, N9591, N4569);
not NOT1 (N9617, N9612);
and AND2 (N9618, N9615, N2516);
nand NAND4 (N9619, N9614, N4664, N6277, N6900);
nand NAND2 (N9620, N9594, N9058);
nor NOR2 (N9621, N9613, N2609);
and AND2 (N9622, N9609, N5477);
or OR3 (N9623, N9619, N2516, N3301);
and AND2 (N9624, N9621, N1905);
not NOT1 (N9625, N9618);
and AND3 (N9626, N9616, N5468, N2014);
nor NOR4 (N9627, N9625, N42, N4774, N3163);
nor NOR3 (N9628, N9620, N3060, N6376);
or OR4 (N9629, N9605, N6832, N4282, N6151);
nand NAND4 (N9630, N9629, N5005, N2011, N2839);
and AND3 (N9631, N9623, N8681, N5433);
buf BUF1 (N9632, N9617);
and AND2 (N9633, N9632, N7203);
nand NAND2 (N9634, N9627, N5475);
nand NAND4 (N9635, N9626, N1836, N3582, N2347);
and AND4 (N9636, N9631, N3099, N753, N1929);
xor XOR2 (N9637, N9635, N8271);
not NOT1 (N9638, N9622);
or OR3 (N9639, N9624, N2774, N9039);
nor NOR2 (N9640, N9628, N3703);
xor XOR2 (N9641, N9636, N5573);
nor NOR4 (N9642, N9633, N5091, N8856, N2352);
not NOT1 (N9643, N9630);
buf BUF1 (N9644, N9596);
nand NAND3 (N9645, N9644, N1951, N8852);
not NOT1 (N9646, N9640);
nand NAND3 (N9647, N9638, N8101, N7125);
nand NAND2 (N9648, N9642, N9169);
xor XOR2 (N9649, N9646, N6579);
buf BUF1 (N9650, N9639);
nor NOR4 (N9651, N9648, N9512, N877, N2130);
nand NAND3 (N9652, N9634, N943, N151);
buf BUF1 (N9653, N9608);
or OR4 (N9654, N9651, N7417, N3400, N6983);
xor XOR2 (N9655, N9653, N3071);
xor XOR2 (N9656, N9655, N5866);
buf BUF1 (N9657, N9637);
not NOT1 (N9658, N9657);
xor XOR2 (N9659, N9645, N3853);
not NOT1 (N9660, N9643);
nand NAND2 (N9661, N9649, N464);
nand NAND2 (N9662, N9647, N1349);
buf BUF1 (N9663, N9660);
nand NAND3 (N9664, N9652, N678, N3110);
and AND4 (N9665, N9664, N4670, N3748, N3509);
xor XOR2 (N9666, N9661, N8352);
nor NOR2 (N9667, N9658, N5323);
xor XOR2 (N9668, N9641, N4551);
buf BUF1 (N9669, N9667);
nand NAND2 (N9670, N9650, N6669);
or OR2 (N9671, N9662, N8315);
nor NOR2 (N9672, N9663, N6756);
or OR3 (N9673, N9671, N4724, N2288);
not NOT1 (N9674, N9656);
xor XOR2 (N9675, N9665, N1283);
xor XOR2 (N9676, N9666, N6760);
nor NOR4 (N9677, N9670, N6206, N4692, N7924);
buf BUF1 (N9678, N9668);
and AND2 (N9679, N9676, N7465);
xor XOR2 (N9680, N9654, N2289);
nor NOR4 (N9681, N9674, N5376, N2496, N737);
nand NAND4 (N9682, N9659, N7328, N8906, N8880);
xor XOR2 (N9683, N9680, N3869);
or OR2 (N9684, N9672, N6841);
buf BUF1 (N9685, N9681);
or OR2 (N9686, N9679, N4829);
xor XOR2 (N9687, N9682, N3240);
xor XOR2 (N9688, N9687, N3773);
xor XOR2 (N9689, N9669, N2405);
xor XOR2 (N9690, N9689, N5040);
not NOT1 (N9691, N9684);
nand NAND2 (N9692, N9683, N7646);
and AND4 (N9693, N9685, N1622, N4057, N786);
nand NAND4 (N9694, N9675, N4222, N8861, N7751);
buf BUF1 (N9695, N9677);
or OR2 (N9696, N9678, N5316);
nor NOR2 (N9697, N9693, N4516);
buf BUF1 (N9698, N9696);
and AND3 (N9699, N9694, N8696, N9189);
xor XOR2 (N9700, N9698, N3873);
nand NAND2 (N9701, N9697, N1847);
xor XOR2 (N9702, N9692, N390);
xor XOR2 (N9703, N9673, N8738);
buf BUF1 (N9704, N9699);
or OR3 (N9705, N9690, N8074, N645);
xor XOR2 (N9706, N9702, N8316);
or OR3 (N9707, N9705, N8458, N7642);
buf BUF1 (N9708, N9701);
nand NAND4 (N9709, N9703, N1001, N5993, N4823);
xor XOR2 (N9710, N9700, N9049);
or OR4 (N9711, N9688, N7602, N5777, N4552);
buf BUF1 (N9712, N9709);
nand NAND2 (N9713, N9704, N1245);
buf BUF1 (N9714, N9706);
nand NAND2 (N9715, N9686, N2531);
nand NAND2 (N9716, N9710, N5331);
or OR4 (N9717, N9695, N887, N7230, N8888);
nor NOR4 (N9718, N9714, N552, N485, N6491);
xor XOR2 (N9719, N9711, N3806);
not NOT1 (N9720, N9719);
nand NAND2 (N9721, N9713, N3888);
nand NAND3 (N9722, N9715, N7958, N1840);
or OR2 (N9723, N9721, N2902);
nor NOR2 (N9724, N9708, N336);
or OR2 (N9725, N9712, N7854);
not NOT1 (N9726, N9716);
or OR3 (N9727, N9718, N532, N8601);
not NOT1 (N9728, N9724);
buf BUF1 (N9729, N9727);
nor NOR4 (N9730, N9729, N75, N614, N4955);
nand NAND4 (N9731, N9730, N6683, N7594, N6642);
nor NOR2 (N9732, N9725, N7967);
nand NAND2 (N9733, N9691, N6163);
xor XOR2 (N9734, N9731, N5066);
nor NOR4 (N9735, N9732, N2123, N7922, N3939);
or OR4 (N9736, N9717, N3473, N7611, N3403);
not NOT1 (N9737, N9707);
xor XOR2 (N9738, N9734, N2903);
and AND3 (N9739, N9728, N7249, N5319);
not NOT1 (N9740, N9735);
and AND4 (N9741, N9723, N4728, N725, N6070);
nor NOR3 (N9742, N9740, N2001, N4530);
and AND4 (N9743, N9737, N7332, N5859, N5839);
buf BUF1 (N9744, N9741);
nand NAND2 (N9745, N9744, N4333);
xor XOR2 (N9746, N9726, N9269);
buf BUF1 (N9747, N9736);
nand NAND4 (N9748, N9739, N1489, N5298, N3684);
nand NAND4 (N9749, N9748, N3217, N966, N6205);
xor XOR2 (N9750, N9746, N1566);
and AND4 (N9751, N9722, N2168, N4988, N577);
not NOT1 (N9752, N9747);
not NOT1 (N9753, N9742);
buf BUF1 (N9754, N9720);
or OR2 (N9755, N9750, N4990);
and AND4 (N9756, N9753, N8834, N2253, N1946);
buf BUF1 (N9757, N9738);
and AND2 (N9758, N9756, N1817);
nor NOR2 (N9759, N9754, N627);
or OR3 (N9760, N9759, N2575, N5552);
buf BUF1 (N9761, N9752);
nand NAND2 (N9762, N9751, N8021);
or OR4 (N9763, N9745, N745, N1720, N7398);
and AND4 (N9764, N9749, N4524, N7830, N1578);
nor NOR3 (N9765, N9762, N538, N5199);
nand NAND3 (N9766, N9758, N5279, N6697);
and AND4 (N9767, N9765, N9346, N6004, N3786);
nor NOR4 (N9768, N9755, N3857, N4763, N2680);
not NOT1 (N9769, N9757);
nor NOR4 (N9770, N9733, N6463, N6219, N1401);
not NOT1 (N9771, N9768);
nand NAND2 (N9772, N9771, N6779);
and AND2 (N9773, N9770, N6446);
not NOT1 (N9774, N9760);
not NOT1 (N9775, N9774);
and AND4 (N9776, N9761, N7501, N9761, N4216);
nor NOR4 (N9777, N9773, N6310, N2584, N8535);
and AND2 (N9778, N9764, N8114);
nor NOR4 (N9779, N9766, N5399, N5866, N974);
nor NOR2 (N9780, N9777, N3588);
xor XOR2 (N9781, N9767, N3691);
not NOT1 (N9782, N9769);
buf BUF1 (N9783, N9763);
nor NOR4 (N9784, N9743, N1562, N2398, N9532);
buf BUF1 (N9785, N9782);
and AND2 (N9786, N9785, N870);
xor XOR2 (N9787, N9776, N4489);
not NOT1 (N9788, N9775);
nand NAND3 (N9789, N9781, N1323, N4380);
and AND3 (N9790, N9780, N5327, N380);
nand NAND3 (N9791, N9784, N5024, N5852);
not NOT1 (N9792, N9790);
and AND4 (N9793, N9788, N7281, N3027, N1904);
or OR2 (N9794, N9779, N9334);
not NOT1 (N9795, N9786);
xor XOR2 (N9796, N9783, N1609);
nor NOR2 (N9797, N9789, N1709);
or OR3 (N9798, N9772, N2134, N7960);
nor NOR3 (N9799, N9797, N7329, N9078);
buf BUF1 (N9800, N9778);
and AND4 (N9801, N9795, N1110, N2146, N556);
xor XOR2 (N9802, N9794, N8359);
not NOT1 (N9803, N9792);
buf BUF1 (N9804, N9801);
or OR4 (N9805, N9793, N7159, N7558, N876);
or OR4 (N9806, N9805, N7352, N809, N9736);
nand NAND2 (N9807, N9799, N7838);
not NOT1 (N9808, N9791);
nand NAND2 (N9809, N9804, N9732);
or OR3 (N9810, N9802, N4275, N8981);
nor NOR3 (N9811, N9796, N7249, N5936);
xor XOR2 (N9812, N9811, N576);
buf BUF1 (N9813, N9798);
or OR2 (N9814, N9803, N5176);
nand NAND4 (N9815, N9813, N6501, N3209, N8964);
buf BUF1 (N9816, N9806);
or OR4 (N9817, N9807, N851, N5142, N2485);
nor NOR4 (N9818, N9814, N5935, N3590, N1610);
or OR2 (N9819, N9816, N9400);
buf BUF1 (N9820, N9808);
nand NAND4 (N9821, N9809, N1874, N4273, N1690);
or OR3 (N9822, N9820, N4744, N6810);
nor NOR2 (N9823, N9819, N7119);
or OR4 (N9824, N9822, N2015, N6241, N8314);
and AND3 (N9825, N9823, N6577, N667);
nand NAND4 (N9826, N9815, N3078, N1489, N6610);
and AND2 (N9827, N9812, N5055);
xor XOR2 (N9828, N9827, N3437);
and AND3 (N9829, N9826, N6955, N130);
nand NAND2 (N9830, N9829, N5440);
xor XOR2 (N9831, N9817, N9014);
nand NAND2 (N9832, N9800, N156);
not NOT1 (N9833, N9787);
not NOT1 (N9834, N9825);
xor XOR2 (N9835, N9810, N8138);
or OR3 (N9836, N9818, N3363, N6837);
nand NAND4 (N9837, N9830, N2123, N7207, N2830);
or OR3 (N9838, N9821, N992, N3023);
buf BUF1 (N9839, N9837);
xor XOR2 (N9840, N9824, N1655);
or OR2 (N9841, N9831, N9790);
nand NAND4 (N9842, N9836, N3044, N2213, N8791);
and AND3 (N9843, N9833, N3700, N5416);
or OR4 (N9844, N9842, N9674, N6504, N3277);
buf BUF1 (N9845, N9834);
nor NOR4 (N9846, N9828, N2162, N4548, N9429);
nor NOR3 (N9847, N9844, N2634, N4596);
buf BUF1 (N9848, N9847);
xor XOR2 (N9849, N9843, N7277);
nor NOR4 (N9850, N9832, N6238, N852, N1315);
not NOT1 (N9851, N9845);
not NOT1 (N9852, N9846);
or OR2 (N9853, N9852, N8893);
nand NAND2 (N9854, N9835, N2210);
nor NOR2 (N9855, N9854, N3927);
not NOT1 (N9856, N9838);
buf BUF1 (N9857, N9850);
not NOT1 (N9858, N9840);
nand NAND4 (N9859, N9848, N46, N6822, N3262);
xor XOR2 (N9860, N9857, N5261);
or OR2 (N9861, N9856, N7353);
nor NOR3 (N9862, N9858, N4423, N7730);
buf BUF1 (N9863, N9859);
xor XOR2 (N9864, N9863, N9144);
not NOT1 (N9865, N9839);
nand NAND2 (N9866, N9841, N5116);
or OR2 (N9867, N9853, N8434);
nand NAND3 (N9868, N9849, N1736, N4384);
buf BUF1 (N9869, N9851);
nor NOR3 (N9870, N9866, N8546, N391);
or OR2 (N9871, N9862, N1392);
not NOT1 (N9872, N9865);
not NOT1 (N9873, N9870);
nand NAND4 (N9874, N9871, N5289, N5634, N2554);
buf BUF1 (N9875, N9872);
nor NOR2 (N9876, N9868, N3766);
or OR3 (N9877, N9875, N6440, N9784);
buf BUF1 (N9878, N9874);
nor NOR2 (N9879, N9864, N2785);
or OR3 (N9880, N9867, N420, N8195);
not NOT1 (N9881, N9878);
xor XOR2 (N9882, N9860, N3355);
buf BUF1 (N9883, N9880);
or OR3 (N9884, N9881, N8267, N9836);
or OR4 (N9885, N9884, N2600, N578, N1016);
xor XOR2 (N9886, N9855, N6812);
nor NOR3 (N9887, N9886, N5918, N4346);
or OR2 (N9888, N9877, N7912);
not NOT1 (N9889, N9879);
or OR4 (N9890, N9861, N1035, N3754, N431);
xor XOR2 (N9891, N9888, N394);
nand NAND3 (N9892, N9887, N5179, N1819);
and AND2 (N9893, N9891, N8270);
not NOT1 (N9894, N9869);
and AND2 (N9895, N9893, N9276);
not NOT1 (N9896, N9873);
xor XOR2 (N9897, N9894, N9344);
or OR2 (N9898, N9876, N9877);
nor NOR2 (N9899, N9897, N1454);
xor XOR2 (N9900, N9895, N7441);
and AND4 (N9901, N9900, N7637, N1643, N5344);
xor XOR2 (N9902, N9901, N4945);
not NOT1 (N9903, N9899);
and AND2 (N9904, N9885, N6963);
xor XOR2 (N9905, N9889, N2678);
xor XOR2 (N9906, N9896, N7814);
nor NOR3 (N9907, N9902, N9703, N5121);
or OR3 (N9908, N9904, N7153, N6438);
xor XOR2 (N9909, N9908, N6523);
buf BUF1 (N9910, N9890);
buf BUF1 (N9911, N9883);
not NOT1 (N9912, N9892);
not NOT1 (N9913, N9905);
nand NAND4 (N9914, N9912, N4077, N2359, N5511);
or OR4 (N9915, N9911, N3106, N5693, N4402);
nor NOR3 (N9916, N9914, N8080, N7182);
not NOT1 (N9917, N9906);
nor NOR4 (N9918, N9913, N7267, N1612, N9811);
buf BUF1 (N9919, N9910);
not NOT1 (N9920, N9915);
nor NOR2 (N9921, N9918, N6060);
not NOT1 (N9922, N9882);
and AND3 (N9923, N9903, N4737, N2511);
buf BUF1 (N9924, N9921);
buf BUF1 (N9925, N9920);
buf BUF1 (N9926, N9919);
nor NOR3 (N9927, N9916, N4656, N9698);
nor NOR4 (N9928, N9909, N4766, N2974, N3028);
nand NAND3 (N9929, N9907, N5120, N1049);
and AND2 (N9930, N9926, N1314);
and AND4 (N9931, N9929, N6959, N344, N5087);
nand NAND3 (N9932, N9925, N9793, N5342);
not NOT1 (N9933, N9922);
and AND3 (N9934, N9930, N5989, N179);
not NOT1 (N9935, N9923);
buf BUF1 (N9936, N9917);
buf BUF1 (N9937, N9924);
xor XOR2 (N9938, N9932, N3680);
or OR4 (N9939, N9928, N1711, N6008, N7764);
or OR3 (N9940, N9934, N8365, N8585);
nand NAND2 (N9941, N9936, N304);
nor NOR4 (N9942, N9927, N9940, N9567, N9325);
buf BUF1 (N9943, N7870);
nand NAND3 (N9944, N9943, N4494, N3251);
and AND4 (N9945, N9931, N1862, N1845, N3073);
or OR4 (N9946, N9939, N9269, N5818, N9448);
buf BUF1 (N9947, N9942);
and AND3 (N9948, N9944, N1496, N7687);
and AND4 (N9949, N9946, N9519, N3954, N1932);
xor XOR2 (N9950, N9941, N1872);
not NOT1 (N9951, N9937);
nor NOR2 (N9952, N9951, N5303);
nor NOR4 (N9953, N9938, N9569, N8609, N3845);
xor XOR2 (N9954, N9948, N7719);
nand NAND4 (N9955, N9898, N4588, N1348, N6744);
or OR2 (N9956, N9945, N6081);
not NOT1 (N9957, N9953);
or OR2 (N9958, N9933, N9856);
xor XOR2 (N9959, N9958, N3867);
and AND4 (N9960, N9955, N2198, N4746, N9395);
xor XOR2 (N9961, N9950, N1810);
xor XOR2 (N9962, N9949, N6965);
or OR2 (N9963, N9935, N7);
not NOT1 (N9964, N9957);
not NOT1 (N9965, N9960);
buf BUF1 (N9966, N9963);
buf BUF1 (N9967, N9962);
buf BUF1 (N9968, N9947);
or OR3 (N9969, N9964, N1207, N1139);
buf BUF1 (N9970, N9967);
and AND3 (N9971, N9954, N7702, N4120);
buf BUF1 (N9972, N9966);
xor XOR2 (N9973, N9952, N9786);
buf BUF1 (N9974, N9971);
not NOT1 (N9975, N9972);
not NOT1 (N9976, N9968);
not NOT1 (N9977, N9959);
xor XOR2 (N9978, N9956, N10);
nand NAND3 (N9979, N9974, N8284, N9363);
and AND4 (N9980, N9961, N2128, N564, N9351);
nor NOR4 (N9981, N9978, N5415, N4295, N9356);
nor NOR3 (N9982, N9970, N6441, N7222);
xor XOR2 (N9983, N9973, N9039);
or OR3 (N9984, N9965, N7776, N8018);
and AND3 (N9985, N9975, N6010, N1299);
not NOT1 (N9986, N9969);
nand NAND4 (N9987, N9981, N5221, N988, N7656);
nor NOR4 (N9988, N9982, N9383, N860, N916);
not NOT1 (N9989, N9983);
not NOT1 (N9990, N9976);
and AND3 (N9991, N9985, N1578, N9435);
or OR2 (N9992, N9990, N4888);
xor XOR2 (N9993, N9987, N9990);
nand NAND2 (N9994, N9988, N9845);
or OR2 (N9995, N9980, N5470);
buf BUF1 (N9996, N9989);
nand NAND2 (N9997, N9979, N1006);
xor XOR2 (N9998, N9992, N3717);
and AND2 (N9999, N9995, N7592);
or OR3 (N10000, N9996, N8116, N3622);
not NOT1 (N10001, N9998);
not NOT1 (N10002, N9997);
xor XOR2 (N10003, N9991, N5032);
not NOT1 (N10004, N9977);
and AND4 (N10005, N9993, N5023, N4760, N2962);
nand NAND4 (N10006, N9999, N5428, N1833, N2192);
nor NOR3 (N10007, N10000, N5813, N9529);
nand NAND4 (N10008, N10004, N4540, N6585, N2588);
nand NAND3 (N10009, N9994, N2867, N4369);
and AND4 (N10010, N9986, N1925, N2689, N6837);
xor XOR2 (N10011, N10010, N8774);
buf BUF1 (N10012, N10006);
not NOT1 (N10013, N9984);
and AND2 (N10014, N10007, N6626);
and AND2 (N10015, N10012, N601);
nor NOR4 (N10016, N10001, N6201, N6872, N5649);
not NOT1 (N10017, N10011);
or OR2 (N10018, N10005, N2134);
buf BUF1 (N10019, N10017);
nor NOR2 (N10020, N10002, N4507);
buf BUF1 (N10021, N10018);
xor XOR2 (N10022, N10008, N2252);
buf BUF1 (N10023, N10019);
not NOT1 (N10024, N10003);
or OR2 (N10025, N10023, N5435);
and AND3 (N10026, N10025, N6589, N2638);
buf BUF1 (N10027, N10015);
xor XOR2 (N10028, N10016, N3727);
xor XOR2 (N10029, N10028, N5925);
nor NOR4 (N10030, N10020, N3735, N9079, N5018);
buf BUF1 (N10031, N10013);
nor NOR3 (N10032, N10027, N3260, N2547);
and AND3 (N10033, N10021, N5521, N297);
or OR4 (N10034, N10030, N6209, N7650, N9506);
buf BUF1 (N10035, N10014);
not NOT1 (N10036, N10029);
nor NOR3 (N10037, N10031, N4675, N6095);
nor NOR3 (N10038, N10036, N4673, N5732);
buf BUF1 (N10039, N10024);
nand NAND4 (N10040, N10035, N8340, N4599, N2812);
or OR4 (N10041, N10037, N6428, N1273, N4642);
not NOT1 (N10042, N10022);
or OR3 (N10043, N10039, N8245, N5430);
and AND3 (N10044, N10043, N8572, N9527);
and AND4 (N10045, N10009, N7273, N1457, N2932);
xor XOR2 (N10046, N10044, N8300);
nand NAND2 (N10047, N10034, N8341);
nor NOR2 (N10048, N10042, N999);
and AND4 (N10049, N10041, N5422, N4279, N9405);
or OR3 (N10050, N10040, N8222, N6431);
nor NOR2 (N10051, N10032, N7725);
xor XOR2 (N10052, N10048, N8700);
buf BUF1 (N10053, N10038);
and AND2 (N10054, N10053, N5204);
nand NAND4 (N10055, N10033, N8029, N3336, N6030);
or OR3 (N10056, N10054, N9759, N9921);
or OR2 (N10057, N10047, N5646);
not NOT1 (N10058, N10055);
or OR4 (N10059, N10052, N6880, N10028, N9388);
or OR4 (N10060, N10046, N8329, N4939, N5688);
nor NOR4 (N10061, N10059, N1796, N2984, N6406);
xor XOR2 (N10062, N10049, N2288);
and AND3 (N10063, N10060, N2587, N8766);
not NOT1 (N10064, N10051);
buf BUF1 (N10065, N10050);
nand NAND3 (N10066, N10057, N6798, N4291);
xor XOR2 (N10067, N10065, N2422);
not NOT1 (N10068, N10026);
and AND3 (N10069, N10064, N6503, N8229);
nand NAND4 (N10070, N10062, N5817, N6684, N2519);
nor NOR2 (N10071, N10069, N7779);
xor XOR2 (N10072, N10061, N1875);
nand NAND2 (N10073, N10071, N4756);
nor NOR2 (N10074, N10066, N6037);
xor XOR2 (N10075, N10070, N1320);
nor NOR2 (N10076, N10073, N5356);
not NOT1 (N10077, N10068);
nand NAND4 (N10078, N10063, N3035, N8644, N6461);
nor NOR4 (N10079, N10075, N8024, N5117, N6919);
nor NOR3 (N10080, N10072, N7587, N6946);
and AND2 (N10081, N10045, N61);
xor XOR2 (N10082, N10078, N721);
buf BUF1 (N10083, N10058);
or OR2 (N10084, N10067, N7045);
xor XOR2 (N10085, N10074, N8540);
or OR4 (N10086, N10080, N6962, N10018, N7628);
buf BUF1 (N10087, N10084);
not NOT1 (N10088, N10085);
or OR4 (N10089, N10083, N91, N7514, N1418);
nor NOR4 (N10090, N10089, N8700, N8216, N2192);
and AND2 (N10091, N10082, N9001);
nor NOR3 (N10092, N10086, N9988, N5251);
or OR4 (N10093, N10091, N259, N1891, N8524);
not NOT1 (N10094, N10088);
not NOT1 (N10095, N10081);
nand NAND4 (N10096, N10092, N7554, N9361, N6747);
or OR4 (N10097, N10076, N6259, N916, N6248);
nand NAND2 (N10098, N10093, N243);
xor XOR2 (N10099, N10087, N9126);
or OR4 (N10100, N10056, N4394, N6625, N8454);
or OR3 (N10101, N10079, N9622, N2439);
nor NOR4 (N10102, N10094, N6564, N5457, N6515);
xor XOR2 (N10103, N10097, N3286);
buf BUF1 (N10104, N10099);
xor XOR2 (N10105, N10098, N3047);
or OR2 (N10106, N10104, N5105);
xor XOR2 (N10107, N10106, N8112);
and AND2 (N10108, N10105, N8131);
nor NOR3 (N10109, N10077, N4177, N3055);
xor XOR2 (N10110, N10101, N1387);
nand NAND2 (N10111, N10110, N9053);
not NOT1 (N10112, N10107);
nand NAND2 (N10113, N10095, N5553);
nor NOR2 (N10114, N10100, N2457);
buf BUF1 (N10115, N10108);
not NOT1 (N10116, N10090);
xor XOR2 (N10117, N10115, N6036);
nand NAND4 (N10118, N10103, N2331, N1346, N4515);
buf BUF1 (N10119, N10096);
not NOT1 (N10120, N10111);
not NOT1 (N10121, N10117);
not NOT1 (N10122, N10113);
or OR2 (N10123, N10112, N3907);
xor XOR2 (N10124, N10121, N2761);
or OR2 (N10125, N10120, N1811);
buf BUF1 (N10126, N10118);
nor NOR4 (N10127, N10126, N7223, N3319, N3015);
nand NAND4 (N10128, N10122, N4603, N730, N7187);
not NOT1 (N10129, N10119);
xor XOR2 (N10130, N10123, N7828);
nor NOR4 (N10131, N10125, N5048, N4068, N1449);
nand NAND4 (N10132, N10109, N3723, N3084, N2366);
buf BUF1 (N10133, N10129);
xor XOR2 (N10134, N10133, N7851);
buf BUF1 (N10135, N10128);
nand NAND2 (N10136, N10127, N9719);
and AND3 (N10137, N10124, N8900, N8999);
or OR4 (N10138, N10116, N2367, N5342, N2884);
not NOT1 (N10139, N10114);
nor NOR3 (N10140, N10134, N9005, N9974);
or OR4 (N10141, N10135, N4567, N7016, N2411);
buf BUF1 (N10142, N10137);
xor XOR2 (N10143, N10131, N5857);
nor NOR2 (N10144, N10142, N5426);
nand NAND3 (N10145, N10132, N8118, N4164);
buf BUF1 (N10146, N10136);
nand NAND2 (N10147, N10145, N484);
xor XOR2 (N10148, N10144, N9603);
nand NAND4 (N10149, N10138, N6440, N3233, N9854);
and AND3 (N10150, N10140, N5932, N1980);
buf BUF1 (N10151, N10143);
buf BUF1 (N10152, N10148);
nor NOR3 (N10153, N10130, N6945, N3858);
and AND2 (N10154, N10150, N3608);
nand NAND2 (N10155, N10151, N1005);
or OR3 (N10156, N10154, N4862, N614);
and AND4 (N10157, N10153, N1193, N8545, N1168);
nand NAND2 (N10158, N10141, N828);
xor XOR2 (N10159, N10156, N375);
or OR3 (N10160, N10155, N8001, N1228);
xor XOR2 (N10161, N10139, N4718);
xor XOR2 (N10162, N10161, N5114);
nor NOR3 (N10163, N10152, N4043, N1830);
not NOT1 (N10164, N10149);
buf BUF1 (N10165, N10147);
or OR4 (N10166, N10164, N8518, N775, N8032);
nor NOR4 (N10167, N10158, N7687, N1878, N5786);
nor NOR2 (N10168, N10165, N5855);
xor XOR2 (N10169, N10162, N5764);
nor NOR2 (N10170, N10159, N1057);
xor XOR2 (N10171, N10169, N4261);
nor NOR3 (N10172, N10171, N7028, N5634);
nor NOR2 (N10173, N10172, N986);
xor XOR2 (N10174, N10168, N1293);
or OR2 (N10175, N10102, N5260);
and AND4 (N10176, N10146, N5068, N4367, N5614);
xor XOR2 (N10177, N10174, N2362);
buf BUF1 (N10178, N10170);
buf BUF1 (N10179, N10166);
not NOT1 (N10180, N10173);
xor XOR2 (N10181, N10175, N6956);
xor XOR2 (N10182, N10167, N953);
buf BUF1 (N10183, N10163);
buf BUF1 (N10184, N10182);
buf BUF1 (N10185, N10179);
xor XOR2 (N10186, N10183, N3454);
nor NOR3 (N10187, N10176, N9797, N2208);
and AND4 (N10188, N10186, N8380, N3948, N5024);
buf BUF1 (N10189, N10184);
buf BUF1 (N10190, N10157);
or OR2 (N10191, N10160, N4684);
nand NAND2 (N10192, N10189, N5037);
nor NOR4 (N10193, N10180, N655, N1977, N3727);
or OR4 (N10194, N10178, N7445, N4802, N6149);
nor NOR4 (N10195, N10190, N779, N1906, N5135);
nor NOR4 (N10196, N10187, N8677, N8657, N9248);
nand NAND3 (N10197, N10185, N2087, N8013);
xor XOR2 (N10198, N10188, N2269);
nor NOR2 (N10199, N10181, N9285);
nor NOR4 (N10200, N10191, N4770, N2544, N7932);
nor NOR3 (N10201, N10193, N10119, N1383);
nor NOR2 (N10202, N10177, N6627);
not NOT1 (N10203, N10198);
or OR4 (N10204, N10194, N7975, N9080, N8442);
buf BUF1 (N10205, N10192);
and AND3 (N10206, N10204, N840, N6045);
nand NAND2 (N10207, N10203, N9315);
buf BUF1 (N10208, N10207);
or OR2 (N10209, N10205, N5818);
or OR2 (N10210, N10206, N2512);
and AND2 (N10211, N10197, N10060);
not NOT1 (N10212, N10196);
buf BUF1 (N10213, N10211);
not NOT1 (N10214, N10212);
buf BUF1 (N10215, N10214);
nand NAND4 (N10216, N10201, N5943, N9739, N1111);
not NOT1 (N10217, N10213);
nor NOR4 (N10218, N10209, N6952, N804, N2196);
or OR3 (N10219, N10215, N6276, N6146);
not NOT1 (N10220, N10219);
not NOT1 (N10221, N10218);
not NOT1 (N10222, N10216);
not NOT1 (N10223, N10199);
and AND3 (N10224, N10210, N9173, N1518);
and AND4 (N10225, N10208, N3764, N8922, N7632);
not NOT1 (N10226, N10200);
or OR3 (N10227, N10222, N2201, N4650);
nor NOR3 (N10228, N10225, N3084, N4845);
nor NOR2 (N10229, N10224, N8013);
and AND2 (N10230, N10229, N9458);
nor NOR2 (N10231, N10227, N57);
not NOT1 (N10232, N10202);
xor XOR2 (N10233, N10195, N5944);
xor XOR2 (N10234, N10226, N6241);
and AND4 (N10235, N10220, N10065, N1396, N8837);
xor XOR2 (N10236, N10233, N246);
nor NOR3 (N10237, N10228, N8090, N6588);
not NOT1 (N10238, N10231);
or OR4 (N10239, N10238, N915, N7558, N9807);
not NOT1 (N10240, N10217);
xor XOR2 (N10241, N10237, N1408);
xor XOR2 (N10242, N10240, N5630);
xor XOR2 (N10243, N10234, N2028);
buf BUF1 (N10244, N10230);
xor XOR2 (N10245, N10243, N4646);
nor NOR3 (N10246, N10245, N4624, N625);
nor NOR3 (N10247, N10241, N7947, N2445);
nand NAND4 (N10248, N10223, N606, N1396, N8015);
buf BUF1 (N10249, N10244);
nor NOR4 (N10250, N10242, N2278, N4234, N8673);
nor NOR3 (N10251, N10239, N7996, N6391);
not NOT1 (N10252, N10250);
not NOT1 (N10253, N10221);
xor XOR2 (N10254, N10253, N5547);
nor NOR2 (N10255, N10249, N4268);
buf BUF1 (N10256, N10235);
not NOT1 (N10257, N10236);
xor XOR2 (N10258, N10256, N3632);
xor XOR2 (N10259, N10246, N7349);
xor XOR2 (N10260, N10232, N32);
xor XOR2 (N10261, N10248, N312);
or OR3 (N10262, N10247, N6557, N8297);
or OR2 (N10263, N10252, N4149);
and AND3 (N10264, N10261, N3664, N9885);
and AND4 (N10265, N10255, N2062, N476, N8148);
xor XOR2 (N10266, N10265, N3400);
not NOT1 (N10267, N10254);
buf BUF1 (N10268, N10260);
nand NAND2 (N10269, N10258, N1929);
buf BUF1 (N10270, N10262);
and AND2 (N10271, N10257, N7540);
nor NOR4 (N10272, N10263, N4662, N6791, N6513);
nor NOR4 (N10273, N10272, N7604, N1466, N1069);
xor XOR2 (N10274, N10273, N7194);
xor XOR2 (N10275, N10267, N6846);
xor XOR2 (N10276, N10270, N9856);
not NOT1 (N10277, N10276);
nor NOR4 (N10278, N10259, N1557, N7314, N6146);
and AND4 (N10279, N10264, N7111, N1152, N8044);
nand NAND4 (N10280, N10277, N8701, N8446, N9380);
or OR4 (N10281, N10269, N7237, N147, N5062);
buf BUF1 (N10282, N10268);
and AND2 (N10283, N10251, N5051);
nor NOR4 (N10284, N10281, N4458, N3922, N4070);
nor NOR3 (N10285, N10266, N1330, N6976);
not NOT1 (N10286, N10283);
nor NOR4 (N10287, N10274, N298, N7559, N4372);
buf BUF1 (N10288, N10287);
nor NOR2 (N10289, N10282, N3164);
xor XOR2 (N10290, N10286, N7177);
xor XOR2 (N10291, N10279, N9152);
nand NAND2 (N10292, N10288, N1957);
or OR3 (N10293, N10291, N3696, N2154);
and AND3 (N10294, N10278, N4266, N10155);
xor XOR2 (N10295, N10275, N214);
nand NAND3 (N10296, N10292, N3494, N8167);
and AND3 (N10297, N10271, N4653, N7287);
xor XOR2 (N10298, N10280, N3732);
nand NAND2 (N10299, N10295, N2245);
or OR4 (N10300, N10293, N8774, N108, N7754);
xor XOR2 (N10301, N10285, N9689);
nand NAND4 (N10302, N10296, N6533, N7558, N7759);
and AND3 (N10303, N10297, N2691, N10052);
buf BUF1 (N10304, N10301);
nand NAND2 (N10305, N10304, N5689);
nand NAND2 (N10306, N10294, N6540);
not NOT1 (N10307, N10300);
and AND4 (N10308, N10307, N3717, N3930, N6637);
nand NAND2 (N10309, N10308, N10261);
and AND3 (N10310, N10305, N7289, N1386);
buf BUF1 (N10311, N10303);
not NOT1 (N10312, N10298);
buf BUF1 (N10313, N10290);
nor NOR3 (N10314, N10310, N9328, N10220);
and AND4 (N10315, N10311, N10281, N2611, N4629);
buf BUF1 (N10316, N10299);
nor NOR2 (N10317, N10315, N5254);
nand NAND3 (N10318, N10306, N2411, N4499);
and AND3 (N10319, N10317, N7203, N1774);
and AND3 (N10320, N10319, N4917, N5956);
and AND4 (N10321, N10313, N7436, N6537, N4494);
and AND2 (N10322, N10312, N4422);
nand NAND4 (N10323, N10302, N5128, N3397, N1231);
and AND2 (N10324, N10322, N2675);
and AND2 (N10325, N10309, N6092);
or OR3 (N10326, N10324, N2235, N9029);
not NOT1 (N10327, N10314);
xor XOR2 (N10328, N10318, N10168);
nor NOR4 (N10329, N10328, N7602, N4779, N2566);
not NOT1 (N10330, N10289);
not NOT1 (N10331, N10330);
nor NOR3 (N10332, N10326, N4718, N6582);
nand NAND4 (N10333, N10327, N8282, N1429, N630);
not NOT1 (N10334, N10331);
nor NOR3 (N10335, N10332, N246, N5157);
nand NAND2 (N10336, N10335, N8293);
or OR2 (N10337, N10316, N9581);
nand NAND2 (N10338, N10284, N8130);
buf BUF1 (N10339, N10333);
xor XOR2 (N10340, N10338, N8083);
not NOT1 (N10341, N10325);
not NOT1 (N10342, N10321);
nor NOR4 (N10343, N10342, N8238, N1869, N5225);
nand NAND2 (N10344, N10329, N2098);
xor XOR2 (N10345, N10340, N8794);
buf BUF1 (N10346, N10341);
and AND4 (N10347, N10320, N2460, N2455, N4250);
or OR3 (N10348, N10334, N9285, N2734);
nand NAND2 (N10349, N10344, N3038);
not NOT1 (N10350, N10323);
xor XOR2 (N10351, N10346, N2776);
nor NOR3 (N10352, N10349, N9543, N8403);
xor XOR2 (N10353, N10348, N893);
buf BUF1 (N10354, N10350);
not NOT1 (N10355, N10345);
nor NOR2 (N10356, N10343, N10346);
xor XOR2 (N10357, N10339, N2068);
not NOT1 (N10358, N10354);
and AND3 (N10359, N10356, N9960, N8674);
buf BUF1 (N10360, N10353);
and AND3 (N10361, N10357, N9453, N3249);
or OR4 (N10362, N10358, N7973, N747, N5545);
nand NAND3 (N10363, N10359, N3387, N3000);
not NOT1 (N10364, N10362);
not NOT1 (N10365, N10363);
xor XOR2 (N10366, N10360, N1509);
nand NAND3 (N10367, N10337, N2129, N319);
buf BUF1 (N10368, N10365);
nand NAND2 (N10369, N10355, N2522);
and AND4 (N10370, N10364, N8197, N2315, N4378);
xor XOR2 (N10371, N10336, N9432);
nand NAND3 (N10372, N10369, N3330, N5390);
and AND4 (N10373, N10352, N7125, N4734, N6409);
and AND3 (N10374, N10371, N3790, N5471);
not NOT1 (N10375, N10361);
or OR4 (N10376, N10373, N2400, N8229, N7261);
not NOT1 (N10377, N10376);
not NOT1 (N10378, N10370);
xor XOR2 (N10379, N10351, N2962);
xor XOR2 (N10380, N10374, N10354);
buf BUF1 (N10381, N10377);
and AND2 (N10382, N10372, N54);
and AND2 (N10383, N10375, N209);
not NOT1 (N10384, N10380);
buf BUF1 (N10385, N10379);
and AND2 (N10386, N10366, N5041);
or OR4 (N10387, N10385, N7573, N8302, N5222);
nand NAND4 (N10388, N10382, N6893, N1381, N8254);
buf BUF1 (N10389, N10386);
or OR4 (N10390, N10387, N5878, N4688, N1978);
nand NAND4 (N10391, N10347, N6618, N4015, N2140);
buf BUF1 (N10392, N10384);
nand NAND4 (N10393, N10391, N9160, N10269, N3419);
buf BUF1 (N10394, N10378);
or OR3 (N10395, N10392, N6370, N7046);
and AND2 (N10396, N10393, N1261);
xor XOR2 (N10397, N10381, N6278);
or OR2 (N10398, N10367, N8618);
and AND4 (N10399, N10388, N3685, N8341, N4006);
nor NOR2 (N10400, N10396, N6692);
xor XOR2 (N10401, N10383, N2988);
buf BUF1 (N10402, N10399);
nor NOR3 (N10403, N10400, N9190, N7436);
nor NOR3 (N10404, N10403, N935, N7651);
nor NOR4 (N10405, N10404, N6637, N2902, N3423);
xor XOR2 (N10406, N10405, N9418);
or OR2 (N10407, N10395, N9704);
nand NAND2 (N10408, N10394, N9354);
not NOT1 (N10409, N10397);
not NOT1 (N10410, N10401);
nor NOR2 (N10411, N10406, N5979);
nand NAND2 (N10412, N10390, N10251);
and AND3 (N10413, N10398, N1839, N7182);
and AND2 (N10414, N10407, N4478);
and AND2 (N10415, N10409, N8820);
or OR3 (N10416, N10402, N5299, N6389);
not NOT1 (N10417, N10413);
nand NAND3 (N10418, N10415, N8832, N4860);
nand NAND4 (N10419, N10408, N8157, N2924, N4678);
buf BUF1 (N10420, N10419);
xor XOR2 (N10421, N10411, N3419);
or OR4 (N10422, N10412, N8928, N8127, N5700);
nor NOR2 (N10423, N10389, N4131);
nand NAND2 (N10424, N10416, N7127);
not NOT1 (N10425, N10421);
nor NOR2 (N10426, N10417, N8509);
or OR2 (N10427, N10425, N2194);
xor XOR2 (N10428, N10414, N5428);
not NOT1 (N10429, N10410);
or OR4 (N10430, N10426, N2159, N10229, N9030);
not NOT1 (N10431, N10428);
nand NAND4 (N10432, N10420, N5968, N5857, N3849);
or OR4 (N10433, N10423, N2975, N7471, N5498);
and AND4 (N10434, N10422, N972, N1492, N2474);
xor XOR2 (N10435, N10424, N491);
or OR4 (N10436, N10430, N2670, N899, N1063);
xor XOR2 (N10437, N10433, N4216);
nor NOR3 (N10438, N10436, N6384, N6423);
nor NOR2 (N10439, N10434, N9826);
or OR3 (N10440, N10418, N3769, N300);
or OR2 (N10441, N10431, N2896);
not NOT1 (N10442, N10435);
not NOT1 (N10443, N10440);
buf BUF1 (N10444, N10429);
and AND4 (N10445, N10427, N5358, N2953, N7137);
xor XOR2 (N10446, N10442, N9558);
not NOT1 (N10447, N10443);
nor NOR4 (N10448, N10432, N3522, N546, N6733);
nor NOR2 (N10449, N10445, N9507);
and AND3 (N10450, N10441, N294, N8769);
buf BUF1 (N10451, N10448);
or OR3 (N10452, N10451, N8673, N9703);
or OR4 (N10453, N10368, N4310, N7768, N696);
not NOT1 (N10454, N10447);
not NOT1 (N10455, N10454);
nand NAND2 (N10456, N10450, N6755);
xor XOR2 (N10457, N10456, N434);
nand NAND3 (N10458, N10438, N2216, N9456);
buf BUF1 (N10459, N10453);
not NOT1 (N10460, N10446);
buf BUF1 (N10461, N10457);
or OR4 (N10462, N10444, N6192, N1656, N5797);
buf BUF1 (N10463, N10460);
buf BUF1 (N10464, N10455);
buf BUF1 (N10465, N10437);
or OR3 (N10466, N10461, N111, N6691);
nor NOR3 (N10467, N10466, N4595, N3817);
and AND3 (N10468, N10458, N4463, N8361);
not NOT1 (N10469, N10452);
and AND2 (N10470, N10464, N1872);
xor XOR2 (N10471, N10439, N4681);
nor NOR3 (N10472, N10469, N7518, N8415);
or OR2 (N10473, N10459, N9706);
buf BUF1 (N10474, N10463);
xor XOR2 (N10475, N10473, N302);
buf BUF1 (N10476, N10462);
buf BUF1 (N10477, N10449);
nand NAND2 (N10478, N10470, N674);
nand NAND2 (N10479, N10477, N6515);
not NOT1 (N10480, N10467);
or OR2 (N10481, N10465, N4073);
nor NOR2 (N10482, N10472, N2408);
nor NOR4 (N10483, N10474, N2421, N8528, N5896);
buf BUF1 (N10484, N10471);
nand NAND3 (N10485, N10484, N130, N4973);
and AND4 (N10486, N10482, N8871, N10071, N4039);
or OR4 (N10487, N10483, N9885, N7524, N2976);
nor NOR2 (N10488, N10479, N10422);
not NOT1 (N10489, N10488);
nor NOR2 (N10490, N10478, N6531);
nor NOR2 (N10491, N10489, N9433);
nand NAND4 (N10492, N10490, N3330, N146, N8863);
xor XOR2 (N10493, N10476, N3086);
xor XOR2 (N10494, N10493, N2353);
or OR3 (N10495, N10468, N10139, N2547);
not NOT1 (N10496, N10492);
or OR2 (N10497, N10486, N9981);
nor NOR3 (N10498, N10487, N439, N3556);
not NOT1 (N10499, N10496);
and AND3 (N10500, N10481, N8356, N2475);
and AND3 (N10501, N10499, N8803, N1175);
or OR2 (N10502, N10497, N10137);
xor XOR2 (N10503, N10491, N3832);
nand NAND2 (N10504, N10502, N3963);
or OR3 (N10505, N10485, N4620, N2940);
nand NAND4 (N10506, N10505, N9503, N7068, N3315);
or OR4 (N10507, N10494, N9764, N3719, N3559);
and AND3 (N10508, N10501, N3270, N311);
buf BUF1 (N10509, N10475);
buf BUF1 (N10510, N10498);
or OR2 (N10511, N10510, N8292);
xor XOR2 (N10512, N10507, N1258);
xor XOR2 (N10513, N10506, N5580);
buf BUF1 (N10514, N10508);
or OR2 (N10515, N10495, N7886);
nor NOR2 (N10516, N10515, N5782);
not NOT1 (N10517, N10504);
not NOT1 (N10518, N10480);
not NOT1 (N10519, N10512);
nor NOR2 (N10520, N10513, N5798);
or OR3 (N10521, N10509, N3590, N5889);
or OR3 (N10522, N10514, N8576, N10210);
xor XOR2 (N10523, N10521, N2933);
buf BUF1 (N10524, N10503);
buf BUF1 (N10525, N10518);
and AND3 (N10526, N10523, N5147, N1260);
xor XOR2 (N10527, N10500, N6581);
nand NAND4 (N10528, N10525, N5494, N2299, N9413);
not NOT1 (N10529, N10527);
or OR3 (N10530, N10516, N7770, N6551);
not NOT1 (N10531, N10520);
nand NAND4 (N10532, N10529, N5352, N7862, N2569);
or OR4 (N10533, N10511, N1228, N158, N1921);
xor XOR2 (N10534, N10528, N2140);
or OR2 (N10535, N10533, N10260);
nand NAND2 (N10536, N10535, N278);
nor NOR4 (N10537, N10534, N10032, N2950, N6967);
nand NAND2 (N10538, N10526, N5688);
nor NOR4 (N10539, N10524, N3328, N10360, N3013);
not NOT1 (N10540, N10530);
nor NOR3 (N10541, N10532, N4810, N2574);
or OR2 (N10542, N10541, N5322);
not NOT1 (N10543, N10519);
or OR3 (N10544, N10540, N4251, N3735);
xor XOR2 (N10545, N10544, N9729);
buf BUF1 (N10546, N10536);
not NOT1 (N10547, N10517);
and AND4 (N10548, N10547, N4736, N5993, N1758);
nand NAND4 (N10549, N10539, N5014, N1850, N772);
nand NAND2 (N10550, N10548, N10434);
nand NAND3 (N10551, N10549, N5266, N3428);
and AND2 (N10552, N10538, N3319);
xor XOR2 (N10553, N10522, N10291);
nand NAND2 (N10554, N10551, N5922);
nand NAND2 (N10555, N10543, N86);
xor XOR2 (N10556, N10546, N1218);
not NOT1 (N10557, N10556);
xor XOR2 (N10558, N10557, N9857);
nor NOR4 (N10559, N10550, N6273, N6408, N5208);
nor NOR3 (N10560, N10555, N6063, N2573);
nand NAND2 (N10561, N10552, N7206);
or OR2 (N10562, N10560, N8598);
xor XOR2 (N10563, N10545, N9267);
nand NAND3 (N10564, N10554, N9956, N2810);
and AND2 (N10565, N10542, N8356);
nor NOR2 (N10566, N10561, N9301);
not NOT1 (N10567, N10563);
or OR3 (N10568, N10559, N1194, N7588);
nor NOR3 (N10569, N10553, N2136, N2374);
buf BUF1 (N10570, N10564);
nand NAND3 (N10571, N10537, N5927, N2218);
or OR2 (N10572, N10570, N5372);
not NOT1 (N10573, N10531);
and AND3 (N10574, N10565, N2070, N587);
nor NOR3 (N10575, N10572, N7116, N6938);
not NOT1 (N10576, N10571);
not NOT1 (N10577, N10558);
buf BUF1 (N10578, N10569);
nand NAND4 (N10579, N10576, N8214, N3971, N2825);
buf BUF1 (N10580, N10568);
or OR3 (N10581, N10578, N3237, N6627);
and AND3 (N10582, N10581, N10073, N3646);
nor NOR4 (N10583, N10562, N7990, N4852, N3398);
not NOT1 (N10584, N10575);
xor XOR2 (N10585, N10584, N6603);
or OR3 (N10586, N10577, N7256, N2861);
not NOT1 (N10587, N10580);
not NOT1 (N10588, N10579);
buf BUF1 (N10589, N10566);
and AND3 (N10590, N10585, N959, N6415);
buf BUF1 (N10591, N10590);
and AND2 (N10592, N10586, N3112);
and AND4 (N10593, N10573, N8212, N3587, N4123);
not NOT1 (N10594, N10593);
nand NAND2 (N10595, N10594, N9109);
xor XOR2 (N10596, N10591, N4854);
buf BUF1 (N10597, N10582);
nor NOR3 (N10598, N10597, N10447, N4308);
buf BUF1 (N10599, N10587);
or OR4 (N10600, N10592, N5240, N3382, N1347);
and AND4 (N10601, N10596, N6449, N6948, N5349);
nand NAND2 (N10602, N10588, N1010);
not NOT1 (N10603, N10574);
xor XOR2 (N10604, N10599, N4417);
not NOT1 (N10605, N10567);
nor NOR2 (N10606, N10598, N1075);
not NOT1 (N10607, N10600);
or OR3 (N10608, N10607, N6055, N9692);
nand NAND2 (N10609, N10605, N2619);
nand NAND2 (N10610, N10583, N10474);
nor NOR4 (N10611, N10610, N7515, N7346, N10093);
not NOT1 (N10612, N10602);
and AND4 (N10613, N10609, N2047, N6091, N16);
or OR2 (N10614, N10611, N8025);
nor NOR4 (N10615, N10589, N8387, N137, N984);
and AND3 (N10616, N10608, N2659, N6775);
buf BUF1 (N10617, N10615);
and AND4 (N10618, N10603, N8328, N2532, N8862);
nand NAND4 (N10619, N10618, N2164, N8030, N10260);
nand NAND4 (N10620, N10614, N7737, N9009, N6208);
or OR4 (N10621, N10595, N6605, N4070, N5459);
not NOT1 (N10622, N10616);
buf BUF1 (N10623, N10613);
and AND2 (N10624, N10620, N8288);
and AND3 (N10625, N10604, N4963, N8257);
nand NAND2 (N10626, N10617, N10534);
not NOT1 (N10627, N10622);
buf BUF1 (N10628, N10601);
nand NAND3 (N10629, N10626, N8851, N9914);
buf BUF1 (N10630, N10629);
or OR4 (N10631, N10624, N2810, N1197, N1273);
nor NOR4 (N10632, N10625, N2499, N2268, N6259);
nand NAND2 (N10633, N10621, N62);
nand NAND4 (N10634, N10619, N8460, N8401, N8688);
nand NAND2 (N10635, N10631, N1277);
nand NAND2 (N10636, N10635, N954);
xor XOR2 (N10637, N10636, N2784);
nand NAND3 (N10638, N10632, N10382, N1743);
nor NOR4 (N10639, N10606, N1116, N5418, N907);
or OR3 (N10640, N10634, N1157, N617);
or OR4 (N10641, N10639, N5150, N8773, N8562);
nor NOR4 (N10642, N10633, N1682, N7492, N612);
nand NAND4 (N10643, N10637, N1781, N5429, N6383);
or OR4 (N10644, N10628, N2902, N5826, N8740);
or OR2 (N10645, N10640, N10208);
and AND2 (N10646, N10638, N1217);
nor NOR2 (N10647, N10623, N3706);
not NOT1 (N10648, N10646);
nor NOR4 (N10649, N10612, N1187, N10457, N729);
xor XOR2 (N10650, N10647, N3059);
or OR3 (N10651, N10645, N9575, N7055);
not NOT1 (N10652, N10630);
and AND2 (N10653, N10652, N50);
nand NAND3 (N10654, N10643, N2834, N719);
xor XOR2 (N10655, N10642, N10231);
buf BUF1 (N10656, N10648);
and AND2 (N10657, N10627, N1305);
nor NOR3 (N10658, N10653, N6188, N3688);
nor NOR3 (N10659, N10644, N7669, N6121);
nor NOR4 (N10660, N10651, N7014, N3215, N2651);
nand NAND4 (N10661, N10641, N7743, N9999, N5540);
not NOT1 (N10662, N10659);
not NOT1 (N10663, N10662);
and AND2 (N10664, N10663, N7553);
xor XOR2 (N10665, N10649, N7974);
buf BUF1 (N10666, N10657);
or OR3 (N10667, N10650, N5096, N9297);
or OR3 (N10668, N10666, N9683, N10160);
or OR4 (N10669, N10660, N4736, N7507, N3224);
or OR2 (N10670, N10656, N2372);
nand NAND3 (N10671, N10667, N6896, N2788);
xor XOR2 (N10672, N10661, N1414);
nand NAND3 (N10673, N10672, N10471, N3197);
or OR3 (N10674, N10671, N5704, N4085);
and AND4 (N10675, N10654, N4328, N2695, N4191);
xor XOR2 (N10676, N10669, N7109);
nor NOR2 (N10677, N10673, N354);
or OR4 (N10678, N10655, N5568, N3671, N9202);
nand NAND3 (N10679, N10658, N10431, N8827);
not NOT1 (N10680, N10677);
buf BUF1 (N10681, N10670);
nand NAND2 (N10682, N10679, N6519);
and AND3 (N10683, N10675, N10488, N288);
or OR4 (N10684, N10665, N8695, N3228, N91);
or OR3 (N10685, N10664, N6317, N4968);
and AND4 (N10686, N10683, N5388, N6356, N3587);
buf BUF1 (N10687, N10685);
xor XOR2 (N10688, N10674, N7137);
nand NAND2 (N10689, N10688, N6974);
or OR4 (N10690, N10684, N8904, N3979, N8971);
nand NAND2 (N10691, N10668, N1664);
buf BUF1 (N10692, N10686);
nand NAND3 (N10693, N10678, N8671, N230);
nor NOR4 (N10694, N10682, N4267, N4929, N9028);
nand NAND2 (N10695, N10693, N10614);
or OR3 (N10696, N10689, N8452, N3183);
not NOT1 (N10697, N10690);
xor XOR2 (N10698, N10691, N349);
xor XOR2 (N10699, N10698, N5255);
and AND4 (N10700, N10699, N2713, N1440, N3607);
and AND2 (N10701, N10681, N4582);
nand NAND3 (N10702, N10701, N2334, N8644);
not NOT1 (N10703, N10696);
and AND4 (N10704, N10687, N5079, N2523, N8946);
nand NAND3 (N10705, N10680, N8993, N7205);
not NOT1 (N10706, N10704);
nor NOR3 (N10707, N10694, N5924, N5088);
and AND3 (N10708, N10676, N363, N1122);
or OR4 (N10709, N10705, N9419, N823, N5271);
and AND3 (N10710, N10709, N9757, N5062);
nand NAND4 (N10711, N10703, N6480, N10546, N10673);
or OR4 (N10712, N10708, N6859, N3367, N6278);
and AND2 (N10713, N10702, N1791);
not NOT1 (N10714, N10695);
xor XOR2 (N10715, N10700, N8664);
nor NOR3 (N10716, N10692, N3411, N3728);
and AND4 (N10717, N10710, N4538, N1072, N1223);
not NOT1 (N10718, N10717);
nand NAND3 (N10719, N10697, N7937, N3022);
buf BUF1 (N10720, N10714);
not NOT1 (N10721, N10713);
not NOT1 (N10722, N10716);
and AND3 (N10723, N10718, N10245, N3490);
or OR4 (N10724, N10715, N2671, N9554, N1035);
not NOT1 (N10725, N10707);
and AND3 (N10726, N10720, N10409, N3375);
and AND2 (N10727, N10724, N10114);
and AND3 (N10728, N10712, N1286, N7337);
buf BUF1 (N10729, N10719);
buf BUF1 (N10730, N10729);
and AND4 (N10731, N10725, N820, N5910, N8892);
or OR4 (N10732, N10730, N7926, N464, N3955);
nor NOR4 (N10733, N10731, N6701, N6227, N10353);
nand NAND4 (N10734, N10728, N9225, N2392, N10556);
or OR4 (N10735, N10726, N5278, N8029, N8613);
xor XOR2 (N10736, N10706, N10386);
buf BUF1 (N10737, N10711);
nor NOR3 (N10738, N10734, N1183, N666);
and AND3 (N10739, N10732, N400, N9386);
not NOT1 (N10740, N10721);
nor NOR3 (N10741, N10733, N10267, N2502);
xor XOR2 (N10742, N10739, N3401);
nand NAND3 (N10743, N10740, N6354, N2670);
not NOT1 (N10744, N10742);
and AND2 (N10745, N10744, N262);
xor XOR2 (N10746, N10722, N9760);
not NOT1 (N10747, N10746);
nand NAND2 (N10748, N10727, N4375);
nand NAND2 (N10749, N10747, N3625);
nand NAND3 (N10750, N10735, N9631, N8010);
nand NAND4 (N10751, N10745, N185, N5945, N9200);
buf BUF1 (N10752, N10750);
xor XOR2 (N10753, N10736, N7027);
nand NAND4 (N10754, N10752, N7682, N4208, N4024);
buf BUF1 (N10755, N10753);
and AND4 (N10756, N10754, N4483, N1732, N3821);
nor NOR2 (N10757, N10741, N1534);
and AND4 (N10758, N10738, N4514, N10389, N5427);
or OR4 (N10759, N10751, N10100, N4622, N776);
and AND2 (N10760, N10749, N4208);
or OR4 (N10761, N10723, N380, N850, N1768);
and AND2 (N10762, N10759, N10623);
not NOT1 (N10763, N10758);
not NOT1 (N10764, N10757);
buf BUF1 (N10765, N10756);
nor NOR3 (N10766, N10743, N6479, N573);
nor NOR4 (N10767, N10761, N23, N6362, N8346);
and AND2 (N10768, N10764, N1907);
nor NOR4 (N10769, N10768, N5545, N2750, N10349);
and AND4 (N10770, N10760, N5634, N9992, N9111);
nor NOR4 (N10771, N10737, N4796, N8738, N10493);
nor NOR2 (N10772, N10770, N3826);
buf BUF1 (N10773, N10762);
not NOT1 (N10774, N10771);
nand NAND4 (N10775, N10766, N10188, N4230, N8997);
nand NAND3 (N10776, N10773, N5151, N501);
nor NOR2 (N10777, N10767, N300);
and AND2 (N10778, N10765, N7633);
nand NAND3 (N10779, N10778, N10707, N7051);
not NOT1 (N10780, N10775);
buf BUF1 (N10781, N10755);
xor XOR2 (N10782, N10781, N4102);
buf BUF1 (N10783, N10763);
buf BUF1 (N10784, N10772);
buf BUF1 (N10785, N10780);
nor NOR3 (N10786, N10769, N5633, N9794);
and AND2 (N10787, N10784, N881);
nand NAND3 (N10788, N10782, N9917, N2399);
nor NOR2 (N10789, N10748, N4298);
not NOT1 (N10790, N10785);
and AND3 (N10791, N10789, N132, N398);
buf BUF1 (N10792, N10779);
xor XOR2 (N10793, N10777, N2337);
not NOT1 (N10794, N10776);
nor NOR2 (N10795, N10783, N5589);
and AND4 (N10796, N10774, N8003, N8882, N4308);
and AND4 (N10797, N10790, N6578, N6352, N1267);
not NOT1 (N10798, N10787);
xor XOR2 (N10799, N10796, N3576);
and AND2 (N10800, N10793, N1710);
or OR3 (N10801, N10800, N7825, N6959);
xor XOR2 (N10802, N10794, N2963);
or OR3 (N10803, N10788, N889, N4202);
nor NOR2 (N10804, N10795, N10648);
not NOT1 (N10805, N10804);
and AND2 (N10806, N10798, N3772);
buf BUF1 (N10807, N10805);
buf BUF1 (N10808, N10806);
or OR2 (N10809, N10808, N2901);
xor XOR2 (N10810, N10803, N1515);
buf BUF1 (N10811, N10799);
and AND2 (N10812, N10791, N8563);
and AND2 (N10813, N10792, N6771);
nor NOR2 (N10814, N10810, N3649);
and AND3 (N10815, N10812, N3579, N9881);
buf BUF1 (N10816, N10813);
buf BUF1 (N10817, N10816);
nor NOR3 (N10818, N10809, N745, N3864);
buf BUF1 (N10819, N10815);
nand NAND2 (N10820, N10817, N72);
not NOT1 (N10821, N10820);
nand NAND2 (N10822, N10802, N3654);
nand NAND2 (N10823, N10811, N3203);
nor NOR3 (N10824, N10821, N10033, N9383);
xor XOR2 (N10825, N10823, N5353);
nor NOR2 (N10826, N10818, N568);
not NOT1 (N10827, N10786);
not NOT1 (N10828, N10807);
nand NAND2 (N10829, N10801, N2561);
buf BUF1 (N10830, N10814);
and AND2 (N10831, N10828, N7866);
or OR2 (N10832, N10825, N4944);
not NOT1 (N10833, N10831);
not NOT1 (N10834, N10822);
and AND3 (N10835, N10834, N7820, N7995);
and AND2 (N10836, N10835, N126);
or OR3 (N10837, N10830, N7333, N6296);
nor NOR3 (N10838, N10833, N9925, N8046);
and AND3 (N10839, N10838, N5312, N117);
buf BUF1 (N10840, N10832);
or OR2 (N10841, N10797, N1972);
xor XOR2 (N10842, N10836, N5402);
and AND2 (N10843, N10842, N7518);
buf BUF1 (N10844, N10843);
or OR3 (N10845, N10840, N2411, N2639);
and AND3 (N10846, N10829, N4021, N1010);
buf BUF1 (N10847, N10826);
nor NOR4 (N10848, N10837, N7604, N2768, N29);
and AND2 (N10849, N10848, N9450);
nand NAND2 (N10850, N10839, N2307);
nand NAND4 (N10851, N10846, N9236, N7223, N7974);
not NOT1 (N10852, N10844);
xor XOR2 (N10853, N10852, N4610);
and AND2 (N10854, N10853, N1260);
xor XOR2 (N10855, N10824, N701);
xor XOR2 (N10856, N10841, N2624);
nand NAND3 (N10857, N10819, N6600, N8193);
not NOT1 (N10858, N10856);
nand NAND3 (N10859, N10851, N6504, N1888);
nor NOR3 (N10860, N10857, N3731, N5007);
or OR3 (N10861, N10858, N4464, N10517);
nor NOR2 (N10862, N10845, N9107);
xor XOR2 (N10863, N10849, N2844);
xor XOR2 (N10864, N10847, N5975);
not NOT1 (N10865, N10854);
nand NAND2 (N10866, N10865, N8338);
not NOT1 (N10867, N10859);
or OR3 (N10868, N10860, N6326, N7161);
xor XOR2 (N10869, N10862, N377);
and AND2 (N10870, N10868, N7809);
and AND2 (N10871, N10867, N2032);
not NOT1 (N10872, N10855);
nand NAND2 (N10873, N10869, N9762);
nor NOR3 (N10874, N10873, N3523, N1803);
xor XOR2 (N10875, N10827, N9645);
xor XOR2 (N10876, N10861, N8961);
buf BUF1 (N10877, N10875);
nor NOR3 (N10878, N10866, N6735, N8891);
buf BUF1 (N10879, N10850);
xor XOR2 (N10880, N10876, N7757);
nand NAND2 (N10881, N10864, N9219);
nor NOR3 (N10882, N10877, N9913, N1423);
nor NOR3 (N10883, N10874, N7204, N2008);
xor XOR2 (N10884, N10878, N106);
xor XOR2 (N10885, N10871, N9406);
xor XOR2 (N10886, N10882, N9986);
nor NOR4 (N10887, N10879, N9715, N8619, N341);
xor XOR2 (N10888, N10880, N1890);
buf BUF1 (N10889, N10872);
not NOT1 (N10890, N10885);
nor NOR3 (N10891, N10863, N6394, N593);
or OR2 (N10892, N10883, N2497);
buf BUF1 (N10893, N10870);
xor XOR2 (N10894, N10891, N2972);
or OR2 (N10895, N10888, N10064);
nand NAND4 (N10896, N10881, N797, N398, N2645);
not NOT1 (N10897, N10887);
or OR2 (N10898, N10889, N5716);
nand NAND4 (N10899, N10886, N924, N5997, N4105);
xor XOR2 (N10900, N10890, N6207);
buf BUF1 (N10901, N10898);
buf BUF1 (N10902, N10892);
xor XOR2 (N10903, N10900, N4755);
nor NOR4 (N10904, N10902, N10395, N8032, N2203);
not NOT1 (N10905, N10903);
or OR4 (N10906, N10905, N4183, N956, N7179);
and AND3 (N10907, N10896, N2847, N10544);
nor NOR3 (N10908, N10895, N1570, N4575);
and AND2 (N10909, N10906, N7819);
not NOT1 (N10910, N10897);
not NOT1 (N10911, N10901);
xor XOR2 (N10912, N10893, N4130);
buf BUF1 (N10913, N10894);
not NOT1 (N10914, N10912);
xor XOR2 (N10915, N10913, N10563);
and AND2 (N10916, N10899, N2146);
not NOT1 (N10917, N10914);
or OR4 (N10918, N10915, N1879, N7323, N2711);
nand NAND2 (N10919, N10908, N9767);
xor XOR2 (N10920, N10904, N208);
buf BUF1 (N10921, N10884);
and AND2 (N10922, N10911, N10552);
buf BUF1 (N10923, N10907);
nand NAND4 (N10924, N10916, N1258, N185, N3369);
buf BUF1 (N10925, N10910);
buf BUF1 (N10926, N10920);
nor NOR3 (N10927, N10918, N1174, N4625);
buf BUF1 (N10928, N10923);
nor NOR4 (N10929, N10917, N3872, N8836, N5118);
nand NAND3 (N10930, N10922, N6552, N2445);
nand NAND4 (N10931, N10924, N1293, N7043, N3998);
nand NAND3 (N10932, N10929, N9479, N1561);
nand NAND4 (N10933, N10909, N4670, N8132, N2235);
and AND2 (N10934, N10925, N10053);
nor NOR2 (N10935, N10919, N4771);
or OR2 (N10936, N10927, N2959);
buf BUF1 (N10937, N10936);
and AND4 (N10938, N10937, N5330, N374, N2997);
and AND3 (N10939, N10926, N9304, N4798);
and AND4 (N10940, N10928, N1356, N9994, N8675);
or OR3 (N10941, N10935, N3613, N3084);
or OR4 (N10942, N10921, N7180, N5928, N6904);
and AND3 (N10943, N10938, N5603, N10095);
nor NOR2 (N10944, N10931, N9067);
xor XOR2 (N10945, N10944, N2007);
and AND2 (N10946, N10942, N2744);
or OR4 (N10947, N10940, N2723, N4482, N10535);
buf BUF1 (N10948, N10939);
xor XOR2 (N10949, N10934, N5055);
nor NOR4 (N10950, N10941, N1867, N2504, N9199);
not NOT1 (N10951, N10946);
nor NOR2 (N10952, N10949, N2767);
and AND3 (N10953, N10930, N2141, N1105);
and AND4 (N10954, N10953, N3415, N2033, N1672);
nand NAND4 (N10955, N10933, N1973, N4479, N10914);
nand NAND3 (N10956, N10943, N7788, N3725);
xor XOR2 (N10957, N10932, N246);
not NOT1 (N10958, N10955);
and AND2 (N10959, N10954, N3435);
not NOT1 (N10960, N10957);
and AND4 (N10961, N10956, N14, N30, N6103);
xor XOR2 (N10962, N10959, N3588);
nand NAND2 (N10963, N10960, N3041);
nand NAND3 (N10964, N10958, N6482, N10797);
nor NOR4 (N10965, N10950, N2141, N325, N3905);
or OR3 (N10966, N10947, N10708, N7235);
xor XOR2 (N10967, N10965, N5663);
buf BUF1 (N10968, N10951);
nor NOR3 (N10969, N10961, N1982, N6571);
nand NAND3 (N10970, N10969, N5829, N7558);
not NOT1 (N10971, N10962);
nand NAND3 (N10972, N10966, N3316, N1334);
and AND2 (N10973, N10972, N10820);
nor NOR3 (N10974, N10963, N10010, N6072);
xor XOR2 (N10975, N10971, N6724);
buf BUF1 (N10976, N10974);
xor XOR2 (N10977, N10975, N6229);
nand NAND4 (N10978, N10976, N4277, N9182, N1640);
xor XOR2 (N10979, N10977, N480);
or OR3 (N10980, N10952, N10814, N7798);
not NOT1 (N10981, N10964);
xor XOR2 (N10982, N10978, N5850);
buf BUF1 (N10983, N10980);
and AND3 (N10984, N10981, N8800, N9107);
nand NAND2 (N10985, N10967, N4450);
not NOT1 (N10986, N10970);
nor NOR3 (N10987, N10982, N3704, N5424);
and AND2 (N10988, N10948, N4230);
nand NAND2 (N10989, N10968, N9821);
nor NOR4 (N10990, N10986, N8913, N2460, N9214);
not NOT1 (N10991, N10979);
nor NOR4 (N10992, N10973, N3091, N2790, N6765);
nand NAND4 (N10993, N10983, N3059, N9809, N1236);
or OR2 (N10994, N10985, N7016);
and AND4 (N10995, N10992, N1368, N9948, N8178);
or OR3 (N10996, N10988, N2374, N7658);
xor XOR2 (N10997, N10984, N100);
or OR2 (N10998, N10994, N8001);
or OR3 (N10999, N10997, N5726, N4173);
xor XOR2 (N11000, N10998, N9684);
nor NOR2 (N11001, N11000, N10218);
buf BUF1 (N11002, N10989);
nand NAND2 (N11003, N10999, N10451);
and AND2 (N11004, N10995, N4119);
nor NOR3 (N11005, N10993, N2773, N5784);
not NOT1 (N11006, N11004);
xor XOR2 (N11007, N10945, N4459);
not NOT1 (N11008, N11002);
nor NOR2 (N11009, N10991, N7549);
nor NOR3 (N11010, N10987, N10553, N9934);
xor XOR2 (N11011, N11001, N1204);
buf BUF1 (N11012, N10990);
nand NAND2 (N11013, N11006, N10231);
not NOT1 (N11014, N11011);
buf BUF1 (N11015, N11007);
or OR3 (N11016, N11014, N10712, N9874);
not NOT1 (N11017, N10996);
buf BUF1 (N11018, N11008);
nand NAND3 (N11019, N11015, N1595, N6325);
xor XOR2 (N11020, N11017, N8304);
and AND2 (N11021, N11005, N5141);
and AND3 (N11022, N11018, N5809, N4024);
and AND4 (N11023, N11016, N6383, N7944, N853);
xor XOR2 (N11024, N11003, N1463);
buf BUF1 (N11025, N11010);
xor XOR2 (N11026, N11019, N6989);
and AND4 (N11027, N11020, N4269, N7347, N3574);
xor XOR2 (N11028, N11012, N9385);
nor NOR2 (N11029, N11024, N7150);
not NOT1 (N11030, N11023);
not NOT1 (N11031, N11025);
nor NOR4 (N11032, N11022, N2836, N9726, N6175);
buf BUF1 (N11033, N11013);
and AND4 (N11034, N11021, N664, N2659, N6064);
and AND2 (N11035, N11033, N3834);
xor XOR2 (N11036, N11034, N7859);
and AND3 (N11037, N11030, N83, N2932);
and AND3 (N11038, N11031, N10608, N5781);
not NOT1 (N11039, N11027);
not NOT1 (N11040, N11028);
and AND2 (N11041, N11039, N6068);
nor NOR4 (N11042, N11029, N8249, N3496, N2860);
xor XOR2 (N11043, N11036, N2385);
xor XOR2 (N11044, N11037, N6874);
nand NAND3 (N11045, N11041, N7002, N7909);
and AND3 (N11046, N11035, N478, N2723);
or OR4 (N11047, N11044, N7983, N11027, N3008);
not NOT1 (N11048, N11043);
and AND4 (N11049, N11045, N8648, N6945, N3204);
nand NAND2 (N11050, N11032, N10507);
nor NOR2 (N11051, N11049, N300);
not NOT1 (N11052, N11046);
nand NAND4 (N11053, N11051, N6051, N6147, N5346);
not NOT1 (N11054, N11048);
and AND4 (N11055, N11038, N4622, N2878, N4223);
and AND2 (N11056, N11009, N8948);
and AND4 (N11057, N11047, N2137, N531, N7188);
nor NOR3 (N11058, N11042, N7464, N1286);
nand NAND4 (N11059, N11058, N6875, N10444, N4956);
xor XOR2 (N11060, N11059, N2769);
and AND3 (N11061, N11053, N6033, N7924);
and AND2 (N11062, N11052, N7563);
buf BUF1 (N11063, N11055);
nor NOR2 (N11064, N11060, N3131);
or OR2 (N11065, N11056, N10526);
xor XOR2 (N11066, N11026, N2668);
xor XOR2 (N11067, N11040, N8493);
not NOT1 (N11068, N11065);
xor XOR2 (N11069, N11067, N10980);
buf BUF1 (N11070, N11062);
nand NAND3 (N11071, N11054, N6446, N4835);
buf BUF1 (N11072, N11061);
nor NOR3 (N11073, N11070, N5173, N7681);
nor NOR2 (N11074, N11068, N439);
not NOT1 (N11075, N11073);
not NOT1 (N11076, N11069);
nand NAND4 (N11077, N11050, N4192, N4304, N6070);
nand NAND2 (N11078, N11064, N2728);
or OR2 (N11079, N11071, N10747);
not NOT1 (N11080, N11078);
not NOT1 (N11081, N11063);
nand NAND3 (N11082, N11076, N4908, N9352);
or OR3 (N11083, N11080, N5606, N673);
or OR3 (N11084, N11074, N8359, N7448);
nor NOR3 (N11085, N11072, N2362, N8709);
or OR2 (N11086, N11085, N7606);
nand NAND3 (N11087, N11084, N7912, N8255);
nor NOR2 (N11088, N11081, N8389);
nand NAND3 (N11089, N11082, N9436, N7774);
and AND3 (N11090, N11057, N8055, N954);
not NOT1 (N11091, N11086);
and AND4 (N11092, N11090, N2751, N9327, N10861);
and AND3 (N11093, N11089, N7151, N6744);
or OR3 (N11094, N11077, N768, N2795);
xor XOR2 (N11095, N11079, N6357);
and AND3 (N11096, N11094, N5664, N9963);
not NOT1 (N11097, N11087);
not NOT1 (N11098, N11075);
or OR4 (N11099, N11097, N7601, N7528, N7183);
xor XOR2 (N11100, N11096, N4373);
xor XOR2 (N11101, N11093, N262);
xor XOR2 (N11102, N11095, N2041);
xor XOR2 (N11103, N11088, N6432);
and AND2 (N11104, N11101, N3893);
not NOT1 (N11105, N11103);
nor NOR2 (N11106, N11100, N10833);
xor XOR2 (N11107, N11104, N7815);
nor NOR4 (N11108, N11092, N8568, N1916, N5897);
nor NOR3 (N11109, N11066, N7935, N9139);
not NOT1 (N11110, N11098);
nand NAND2 (N11111, N11099, N4812);
or OR3 (N11112, N11111, N8589, N2257);
nand NAND3 (N11113, N11110, N8868, N6044);
not NOT1 (N11114, N11107);
nor NOR4 (N11115, N11102, N3461, N7444, N8884);
or OR4 (N11116, N11106, N8681, N3605, N5679);
buf BUF1 (N11117, N11114);
nor NOR2 (N11118, N11113, N5437);
not NOT1 (N11119, N11115);
not NOT1 (N11120, N11118);
nor NOR2 (N11121, N11112, N2716);
or OR4 (N11122, N11083, N3548, N2724, N9137);
or OR3 (N11123, N11117, N3099, N11100);
nand NAND3 (N11124, N11116, N9513, N607);
or OR4 (N11125, N11109, N5911, N1955, N9200);
nand NAND4 (N11126, N11091, N609, N5552, N4077);
nand NAND3 (N11127, N11108, N9029, N3242);
and AND3 (N11128, N11119, N4386, N6579);
buf BUF1 (N11129, N11121);
xor XOR2 (N11130, N11124, N8507);
nor NOR2 (N11131, N11123, N4898);
not NOT1 (N11132, N11126);
and AND4 (N11133, N11131, N9399, N3736, N5412);
and AND2 (N11134, N11120, N5583);
nand NAND4 (N11135, N11133, N9420, N562, N4170);
and AND2 (N11136, N11125, N9561);
nor NOR2 (N11137, N11136, N8865);
nand NAND2 (N11138, N11105, N4356);
xor XOR2 (N11139, N11132, N7547);
nand NAND3 (N11140, N11122, N5767, N3121);
not NOT1 (N11141, N11127);
xor XOR2 (N11142, N11134, N7810);
nor NOR4 (N11143, N11139, N9876, N602, N1556);
and AND3 (N11144, N11140, N943, N5968);
not NOT1 (N11145, N11129);
not NOT1 (N11146, N11135);
xor XOR2 (N11147, N11130, N7184);
xor XOR2 (N11148, N11142, N8399);
nor NOR4 (N11149, N11147, N2336, N1523, N4525);
or OR4 (N11150, N11137, N1431, N4710, N5591);
xor XOR2 (N11151, N11145, N6651);
or OR2 (N11152, N11151, N1890);
or OR2 (N11153, N11152, N10353);
and AND2 (N11154, N11150, N8130);
xor XOR2 (N11155, N11149, N8184);
xor XOR2 (N11156, N11144, N8856);
not NOT1 (N11157, N11141);
xor XOR2 (N11158, N11143, N3199);
or OR2 (N11159, N11146, N262);
nand NAND2 (N11160, N11156, N630);
xor XOR2 (N11161, N11159, N2519);
or OR2 (N11162, N11128, N10568);
or OR2 (N11163, N11161, N11094);
buf BUF1 (N11164, N11160);
nand NAND3 (N11165, N11163, N4334, N5869);
buf BUF1 (N11166, N11138);
nor NOR2 (N11167, N11154, N9502);
xor XOR2 (N11168, N11166, N273);
xor XOR2 (N11169, N11164, N10325);
and AND2 (N11170, N11167, N3606);
xor XOR2 (N11171, N11162, N9022);
and AND4 (N11172, N11171, N469, N1415, N100);
nor NOR3 (N11173, N11165, N697, N4194);
nand NAND3 (N11174, N11168, N4260, N4996);
buf BUF1 (N11175, N11158);
xor XOR2 (N11176, N11175, N10826);
nand NAND2 (N11177, N11157, N2277);
nand NAND4 (N11178, N11172, N9016, N2585, N2304);
and AND4 (N11179, N11176, N2504, N4066, N9852);
xor XOR2 (N11180, N11153, N7397);
or OR4 (N11181, N11173, N4268, N5002, N732);
not NOT1 (N11182, N11148);
buf BUF1 (N11183, N11181);
buf BUF1 (N11184, N11183);
or OR4 (N11185, N11155, N9330, N2846, N4901);
or OR4 (N11186, N11180, N4009, N8443, N5508);
or OR2 (N11187, N11186, N8637);
not NOT1 (N11188, N11170);
buf BUF1 (N11189, N11188);
or OR4 (N11190, N11179, N1859, N4806, N1392);
nor NOR4 (N11191, N11182, N10054, N1005, N10219);
and AND2 (N11192, N11178, N6626);
xor XOR2 (N11193, N11174, N5121);
not NOT1 (N11194, N11190);
and AND4 (N11195, N11169, N9755, N4038, N8620);
nor NOR4 (N11196, N11195, N4797, N6282, N299);
buf BUF1 (N11197, N11193);
nand NAND4 (N11198, N11191, N5492, N9700, N7942);
nand NAND2 (N11199, N11185, N3626);
xor XOR2 (N11200, N11189, N3528);
and AND2 (N11201, N11196, N6840);
nor NOR2 (N11202, N11201, N5327);
and AND4 (N11203, N11177, N6803, N6865, N9627);
nand NAND4 (N11204, N11184, N1713, N3090, N10009);
buf BUF1 (N11205, N11194);
and AND2 (N11206, N11198, N9483);
not NOT1 (N11207, N11205);
nand NAND3 (N11208, N11187, N154, N1947);
and AND3 (N11209, N11204, N987, N1996);
or OR4 (N11210, N11206, N7555, N7178, N377);
not NOT1 (N11211, N11200);
or OR2 (N11212, N11210, N6641);
buf BUF1 (N11213, N11208);
not NOT1 (N11214, N11197);
or OR2 (N11215, N11203, N10365);
buf BUF1 (N11216, N11212);
xor XOR2 (N11217, N11214, N907);
and AND3 (N11218, N11216, N911, N1846);
or OR2 (N11219, N11211, N1300);
nor NOR4 (N11220, N11218, N9414, N5931, N9189);
not NOT1 (N11221, N11213);
and AND2 (N11222, N11221, N8460);
or OR3 (N11223, N11207, N9806, N2407);
not NOT1 (N11224, N11209);
nor NOR2 (N11225, N11215, N11085);
and AND3 (N11226, N11202, N1102, N6499);
not NOT1 (N11227, N11217);
and AND2 (N11228, N11224, N9596);
not NOT1 (N11229, N11227);
xor XOR2 (N11230, N11222, N7445);
nand NAND3 (N11231, N11225, N5338, N10214);
not NOT1 (N11232, N11223);
buf BUF1 (N11233, N11230);
and AND4 (N11234, N11220, N2208, N5427, N7882);
and AND3 (N11235, N11199, N5258, N9693);
not NOT1 (N11236, N11219);
and AND4 (N11237, N11233, N2133, N4286, N6259);
buf BUF1 (N11238, N11192);
buf BUF1 (N11239, N11238);
xor XOR2 (N11240, N11235, N5687);
nand NAND4 (N11241, N11232, N1852, N6618, N7846);
and AND4 (N11242, N11236, N3430, N10696, N4163);
or OR4 (N11243, N11241, N7393, N6669, N467);
or OR2 (N11244, N11234, N626);
xor XOR2 (N11245, N11240, N6441);
buf BUF1 (N11246, N11239);
not NOT1 (N11247, N11231);
nand NAND2 (N11248, N11229, N9234);
and AND4 (N11249, N11226, N7467, N44, N2548);
xor XOR2 (N11250, N11242, N6037);
xor XOR2 (N11251, N11250, N6644);
nor NOR3 (N11252, N11237, N1903, N10848);
or OR4 (N11253, N11248, N8640, N7226, N5948);
not NOT1 (N11254, N11228);
and AND3 (N11255, N11251, N9338, N1016);
not NOT1 (N11256, N11245);
nand NAND4 (N11257, N11247, N7291, N5278, N10487);
nand NAND2 (N11258, N11256, N5550);
buf BUF1 (N11259, N11244);
nand NAND2 (N11260, N11243, N3049);
not NOT1 (N11261, N11254);
buf BUF1 (N11262, N11246);
not NOT1 (N11263, N11253);
xor XOR2 (N11264, N11259, N11160);
not NOT1 (N11265, N11264);
and AND3 (N11266, N11257, N6410, N245);
and AND4 (N11267, N11265, N941, N7525, N3806);
buf BUF1 (N11268, N11266);
nand NAND4 (N11269, N11268, N2173, N1992, N5423);
xor XOR2 (N11270, N11261, N207);
and AND2 (N11271, N11270, N7280);
xor XOR2 (N11272, N11267, N424);
not NOT1 (N11273, N11271);
nand NAND3 (N11274, N11249, N9213, N4066);
or OR4 (N11275, N11260, N3989, N7776, N4397);
buf BUF1 (N11276, N11274);
nand NAND4 (N11277, N11272, N4698, N8735, N8783);
or OR2 (N11278, N11273, N479);
or OR2 (N11279, N11277, N2831);
and AND2 (N11280, N11276, N5703);
not NOT1 (N11281, N11263);
not NOT1 (N11282, N11252);
not NOT1 (N11283, N11262);
nor NOR3 (N11284, N11269, N8089, N1392);
or OR2 (N11285, N11284, N1140);
and AND3 (N11286, N11258, N3153, N3593);
and AND4 (N11287, N11279, N2637, N7265, N9316);
buf BUF1 (N11288, N11281);
nand NAND2 (N11289, N11285, N11278);
xor XOR2 (N11290, N1542, N3585);
xor XOR2 (N11291, N11286, N9113);
buf BUF1 (N11292, N11282);
and AND3 (N11293, N11288, N2718, N9923);
or OR3 (N11294, N11289, N5613, N1868);
nand NAND2 (N11295, N11292, N2546);
nor NOR3 (N11296, N11275, N2541, N9136);
xor XOR2 (N11297, N11287, N1103);
nand NAND3 (N11298, N11294, N1616, N4664);
xor XOR2 (N11299, N11297, N1913);
nand NAND3 (N11300, N11296, N8563, N8082);
not NOT1 (N11301, N11255);
nor NOR2 (N11302, N11293, N1589);
not NOT1 (N11303, N11300);
nor NOR4 (N11304, N11291, N1998, N113, N1382);
xor XOR2 (N11305, N11280, N6865);
and AND3 (N11306, N11298, N2313, N1501);
not NOT1 (N11307, N11305);
and AND3 (N11308, N11303, N10323, N10376);
nor NOR2 (N11309, N11290, N1320);
xor XOR2 (N11310, N11307, N419);
nor NOR4 (N11311, N11304, N10873, N4103, N4735);
or OR4 (N11312, N11301, N7984, N9877, N8990);
or OR2 (N11313, N11312, N1873);
or OR4 (N11314, N11309, N5962, N4578, N788);
nand NAND3 (N11315, N11302, N7148, N3869);
or OR4 (N11316, N11314, N426, N7857, N309);
and AND4 (N11317, N11310, N8555, N35, N9383);
or OR2 (N11318, N11299, N9759);
nor NOR4 (N11319, N11306, N3283, N2378, N3126);
or OR2 (N11320, N11317, N1162);
nor NOR4 (N11321, N11319, N3573, N3512, N139);
not NOT1 (N11322, N11283);
nor NOR4 (N11323, N11315, N6063, N1883, N1842);
xor XOR2 (N11324, N11311, N4419);
and AND2 (N11325, N11295, N6262);
and AND4 (N11326, N11318, N9513, N721, N6285);
not NOT1 (N11327, N11313);
buf BUF1 (N11328, N11320);
xor XOR2 (N11329, N11321, N6767);
and AND2 (N11330, N11308, N4261);
nor NOR4 (N11331, N11325, N396, N10525, N7031);
buf BUF1 (N11332, N11327);
xor XOR2 (N11333, N11322, N509);
xor XOR2 (N11334, N11331, N11134);
nand NAND3 (N11335, N11333, N6631, N10199);
nor NOR4 (N11336, N11326, N1069, N210, N3325);
xor XOR2 (N11337, N11328, N891);
not NOT1 (N11338, N11329);
or OR4 (N11339, N11335, N6381, N5145, N5709);
nand NAND2 (N11340, N11323, N3443);
xor XOR2 (N11341, N11338, N6005);
and AND2 (N11342, N11341, N9250);
not NOT1 (N11343, N11337);
and AND3 (N11344, N11332, N7346, N11214);
nor NOR2 (N11345, N11324, N5365);
nor NOR2 (N11346, N11343, N2175);
or OR2 (N11347, N11334, N3764);
or OR3 (N11348, N11340, N8386, N3732);
nor NOR4 (N11349, N11316, N10972, N930, N410);
nor NOR4 (N11350, N11330, N1486, N7551, N6123);
or OR3 (N11351, N11339, N7988, N5945);
buf BUF1 (N11352, N11345);
nor NOR4 (N11353, N11349, N10423, N2600, N11298);
xor XOR2 (N11354, N11347, N8647);
nor NOR2 (N11355, N11348, N546);
and AND2 (N11356, N11355, N1351);
not NOT1 (N11357, N11350);
not NOT1 (N11358, N11352);
and AND3 (N11359, N11356, N9189, N8800);
not NOT1 (N11360, N11357);
not NOT1 (N11361, N11344);
nand NAND3 (N11362, N11342, N9353, N4596);
nor NOR4 (N11363, N11360, N10703, N871, N893);
not NOT1 (N11364, N11353);
nand NAND3 (N11365, N11364, N3600, N8591);
nand NAND4 (N11366, N11354, N7766, N9211, N2611);
not NOT1 (N11367, N11336);
nand NAND4 (N11368, N11361, N11342, N2018, N1508);
or OR3 (N11369, N11346, N5356, N6938);
nand NAND4 (N11370, N11351, N475, N2139, N10086);
nand NAND3 (N11371, N11358, N7239, N11122);
nor NOR3 (N11372, N11370, N5656, N7735);
xor XOR2 (N11373, N11365, N4683);
and AND4 (N11374, N11373, N10508, N3450, N2682);
and AND2 (N11375, N11368, N289);
and AND3 (N11376, N11374, N4784, N8022);
not NOT1 (N11377, N11363);
and AND3 (N11378, N11367, N10148, N647);
xor XOR2 (N11379, N11378, N6031);
xor XOR2 (N11380, N11366, N5039);
buf BUF1 (N11381, N11362);
nor NOR4 (N11382, N11376, N10133, N2058, N9594);
or OR2 (N11383, N11359, N1869);
not NOT1 (N11384, N11375);
nor NOR2 (N11385, N11371, N2594);
xor XOR2 (N11386, N11377, N8160);
not NOT1 (N11387, N11384);
nor NOR2 (N11388, N11380, N6888);
and AND3 (N11389, N11385, N7127, N9509);
not NOT1 (N11390, N11389);
xor XOR2 (N11391, N11386, N6868);
not NOT1 (N11392, N11381);
and AND4 (N11393, N11379, N11251, N1315, N10502);
and AND2 (N11394, N11372, N2636);
nor NOR4 (N11395, N11392, N2856, N8276, N951);
nand NAND4 (N11396, N11394, N3919, N710, N9353);
buf BUF1 (N11397, N11393);
xor XOR2 (N11398, N11388, N2046);
and AND3 (N11399, N11369, N10029, N3316);
or OR3 (N11400, N11396, N3967, N10581);
xor XOR2 (N11401, N11400, N259);
and AND3 (N11402, N11382, N3336, N10355);
xor XOR2 (N11403, N11390, N9699);
nor NOR4 (N11404, N11403, N11295, N9869, N9137);
or OR4 (N11405, N11395, N1176, N7958, N1734);
nand NAND2 (N11406, N11404, N207);
nand NAND4 (N11407, N11398, N1222, N8298, N7730);
nor NOR4 (N11408, N11391, N5145, N1038, N5938);
not NOT1 (N11409, N11387);
or OR4 (N11410, N11409, N5373, N10111, N7471);
nor NOR3 (N11411, N11399, N7401, N1137);
or OR4 (N11412, N11408, N4427, N8874, N7734);
buf BUF1 (N11413, N11412);
or OR2 (N11414, N11383, N7895);
nand NAND2 (N11415, N11405, N755);
nand NAND3 (N11416, N11407, N2913, N9200);
or OR4 (N11417, N11414, N6766, N9969, N33);
and AND2 (N11418, N11417, N7006);
not NOT1 (N11419, N11401);
nand NAND4 (N11420, N11397, N4705, N10678, N2115);
buf BUF1 (N11421, N11416);
or OR4 (N11422, N11413, N9835, N1856, N1388);
not NOT1 (N11423, N11406);
xor XOR2 (N11424, N11418, N8867);
or OR2 (N11425, N11420, N8171);
not NOT1 (N11426, N11421);
or OR4 (N11427, N11425, N3265, N1138, N3094);
nand NAND4 (N11428, N11426, N8872, N235, N4830);
nand NAND3 (N11429, N11424, N9194, N9604);
or OR3 (N11430, N11428, N3568, N7674);
and AND4 (N11431, N11430, N2566, N9122, N7423);
or OR3 (N11432, N11419, N285, N5924);
nand NAND3 (N11433, N11402, N6127, N1495);
xor XOR2 (N11434, N11433, N4884);
not NOT1 (N11435, N11410);
xor XOR2 (N11436, N11415, N11321);
buf BUF1 (N11437, N11411);
buf BUF1 (N11438, N11432);
and AND3 (N11439, N11435, N9154, N10760);
and AND3 (N11440, N11434, N6738, N1608);
buf BUF1 (N11441, N11437);
xor XOR2 (N11442, N11439, N10478);
or OR2 (N11443, N11427, N4605);
nor NOR4 (N11444, N11441, N1061, N8698, N3645);
not NOT1 (N11445, N11438);
and AND4 (N11446, N11429, N2798, N6373, N8407);
buf BUF1 (N11447, N11440);
buf BUF1 (N11448, N11445);
and AND3 (N11449, N11443, N4966, N7035);
buf BUF1 (N11450, N11447);
xor XOR2 (N11451, N11448, N9982);
or OR3 (N11452, N11450, N7226, N2685);
xor XOR2 (N11453, N11444, N6426);
not NOT1 (N11454, N11431);
and AND4 (N11455, N11453, N9107, N2880, N6031);
buf BUF1 (N11456, N11446);
nand NAND2 (N11457, N11451, N1263);
or OR2 (N11458, N11456, N8563);
buf BUF1 (N11459, N11442);
xor XOR2 (N11460, N11449, N10982);
not NOT1 (N11461, N11436);
buf BUF1 (N11462, N11455);
and AND3 (N11463, N11423, N2115, N6826);
and AND4 (N11464, N11452, N5840, N3303, N10772);
nand NAND3 (N11465, N11460, N2890, N1771);
buf BUF1 (N11466, N11458);
and AND3 (N11467, N11457, N978, N1598);
not NOT1 (N11468, N11459);
and AND3 (N11469, N11468, N6427, N11284);
or OR3 (N11470, N11463, N2017, N11407);
xor XOR2 (N11471, N11466, N10106);
nand NAND3 (N11472, N11454, N11261, N2890);
not NOT1 (N11473, N11469);
nand NAND2 (N11474, N11465, N6318);
buf BUF1 (N11475, N11467);
and AND3 (N11476, N11473, N7978, N1291);
buf BUF1 (N11477, N11422);
or OR4 (N11478, N11464, N5526, N312, N4101);
not NOT1 (N11479, N11470);
and AND2 (N11480, N11478, N10648);
or OR4 (N11481, N11462, N656, N4956, N7079);
buf BUF1 (N11482, N11481);
nand NAND2 (N11483, N11475, N7095);
nor NOR2 (N11484, N11477, N9498);
nor NOR2 (N11485, N11479, N4632);
not NOT1 (N11486, N11483);
or OR4 (N11487, N11485, N3919, N7118, N6994);
nand NAND2 (N11488, N11480, N3403);
not NOT1 (N11489, N11482);
not NOT1 (N11490, N11487);
or OR2 (N11491, N11488, N9391);
and AND4 (N11492, N11461, N4454, N8801, N8791);
not NOT1 (N11493, N11490);
or OR3 (N11494, N11492, N7235, N2620);
nor NOR4 (N11495, N11474, N1998, N9542, N4353);
xor XOR2 (N11496, N11491, N1193);
xor XOR2 (N11497, N11489, N8584);
nand NAND2 (N11498, N11476, N3545);
or OR3 (N11499, N11486, N2379, N2314);
or OR2 (N11500, N11484, N11151);
and AND2 (N11501, N11497, N10077);
and AND4 (N11502, N11495, N3613, N9406, N369);
xor XOR2 (N11503, N11472, N5819);
xor XOR2 (N11504, N11498, N404);
xor XOR2 (N11505, N11496, N5560);
buf BUF1 (N11506, N11502);
nand NAND2 (N11507, N11501, N9975);
xor XOR2 (N11508, N11494, N3736);
or OR3 (N11509, N11471, N3002, N661);
nor NOR2 (N11510, N11505, N5149);
or OR2 (N11511, N11510, N691);
not NOT1 (N11512, N11508);
nand NAND4 (N11513, N11493, N4709, N7581, N777);
and AND2 (N11514, N11511, N881);
or OR2 (N11515, N11503, N2597);
xor XOR2 (N11516, N11504, N4621);
not NOT1 (N11517, N11516);
nor NOR3 (N11518, N11506, N9333, N1276);
buf BUF1 (N11519, N11515);
nand NAND3 (N11520, N11507, N10628, N11357);
buf BUF1 (N11521, N11519);
nor NOR3 (N11522, N11513, N3324, N6212);
not NOT1 (N11523, N11521);
and AND3 (N11524, N11522, N310, N144);
nor NOR2 (N11525, N11523, N9166);
buf BUF1 (N11526, N11512);
nand NAND3 (N11527, N11509, N9876, N3500);
or OR2 (N11528, N11524, N9338);
buf BUF1 (N11529, N11525);
not NOT1 (N11530, N11520);
not NOT1 (N11531, N11529);
not NOT1 (N11532, N11528);
and AND3 (N11533, N11526, N8117, N2422);
or OR2 (N11534, N11514, N2339);
buf BUF1 (N11535, N11534);
nor NOR2 (N11536, N11517, N8077);
and AND2 (N11537, N11536, N3959);
not NOT1 (N11538, N11531);
not NOT1 (N11539, N11535);
nor NOR3 (N11540, N11537, N8359, N5937);
not NOT1 (N11541, N11532);
xor XOR2 (N11542, N11533, N1950);
buf BUF1 (N11543, N11530);
not NOT1 (N11544, N11518);
xor XOR2 (N11545, N11544, N3457);
nor NOR4 (N11546, N11527, N8310, N4562, N6716);
nor NOR4 (N11547, N11541, N850, N10519, N8053);
nand NAND3 (N11548, N11538, N4895, N4422);
or OR4 (N11549, N11543, N6591, N3393, N10327);
not NOT1 (N11550, N11540);
not NOT1 (N11551, N11539);
or OR2 (N11552, N11547, N11082);
buf BUF1 (N11553, N11549);
xor XOR2 (N11554, N11553, N1817);
nand NAND3 (N11555, N11554, N3371, N2931);
or OR2 (N11556, N11548, N5915);
nand NAND2 (N11557, N11550, N4347);
or OR2 (N11558, N11557, N8477);
buf BUF1 (N11559, N11558);
xor XOR2 (N11560, N11546, N10845);
nor NOR2 (N11561, N11556, N6769);
not NOT1 (N11562, N11555);
nand NAND4 (N11563, N11560, N8601, N3413, N10883);
buf BUF1 (N11564, N11545);
nor NOR4 (N11565, N11551, N10645, N6182, N9006);
or OR2 (N11566, N11564, N9248);
nor NOR3 (N11567, N11563, N8373, N4140);
and AND4 (N11568, N11561, N3352, N6560, N2343);
and AND4 (N11569, N11559, N782, N6628, N5468);
nor NOR4 (N11570, N11562, N6682, N2598, N9925);
buf BUF1 (N11571, N11500);
or OR4 (N11572, N11567, N7777, N11307, N5428);
or OR4 (N11573, N11570, N3774, N7306, N8224);
or OR3 (N11574, N11571, N11494, N3404);
not NOT1 (N11575, N11499);
buf BUF1 (N11576, N11572);
xor XOR2 (N11577, N11565, N6969);
nor NOR3 (N11578, N11566, N6508, N1157);
xor XOR2 (N11579, N11552, N8466);
buf BUF1 (N11580, N11569);
not NOT1 (N11581, N11568);
xor XOR2 (N11582, N11579, N10740);
xor XOR2 (N11583, N11576, N8661);
nand NAND3 (N11584, N11573, N8380, N9856);
and AND3 (N11585, N11577, N240, N6096);
or OR4 (N11586, N11581, N1920, N11568, N9748);
buf BUF1 (N11587, N11575);
nand NAND3 (N11588, N11587, N3329, N1881);
buf BUF1 (N11589, N11585);
not NOT1 (N11590, N11586);
xor XOR2 (N11591, N11584, N2663);
xor XOR2 (N11592, N11591, N11208);
not NOT1 (N11593, N11582);
buf BUF1 (N11594, N11590);
not NOT1 (N11595, N11588);
xor XOR2 (N11596, N11574, N10643);
xor XOR2 (N11597, N11595, N9366);
or OR2 (N11598, N11589, N7578);
xor XOR2 (N11599, N11596, N1422);
buf BUF1 (N11600, N11597);
buf BUF1 (N11601, N11594);
or OR3 (N11602, N11593, N5924, N389);
nor NOR3 (N11603, N11598, N7923, N8749);
or OR2 (N11604, N11578, N3416);
buf BUF1 (N11605, N11542);
or OR4 (N11606, N11599, N9441, N1261, N1515);
or OR3 (N11607, N11580, N4727, N3101);
xor XOR2 (N11608, N11606, N6746);
xor XOR2 (N11609, N11592, N1122);
not NOT1 (N11610, N11583);
and AND4 (N11611, N11610, N9677, N230, N10757);
xor XOR2 (N11612, N11605, N173);
xor XOR2 (N11613, N11600, N2823);
nand NAND2 (N11614, N11603, N3515);
buf BUF1 (N11615, N11614);
not NOT1 (N11616, N11604);
not NOT1 (N11617, N11608);
not NOT1 (N11618, N11616);
xor XOR2 (N11619, N11618, N4545);
not NOT1 (N11620, N11601);
and AND3 (N11621, N11609, N6246, N4057);
not NOT1 (N11622, N11617);
not NOT1 (N11623, N11613);
not NOT1 (N11624, N11612);
buf BUF1 (N11625, N11619);
xor XOR2 (N11626, N11622, N3116);
or OR3 (N11627, N11626, N10604, N1891);
buf BUF1 (N11628, N11620);
and AND3 (N11629, N11602, N11060, N6493);
buf BUF1 (N11630, N11629);
xor XOR2 (N11631, N11628, N4472);
nor NOR3 (N11632, N11615, N1693, N7407);
nor NOR4 (N11633, N11611, N1594, N6110, N3461);
not NOT1 (N11634, N11631);
nand NAND3 (N11635, N11630, N8460, N6209);
not NOT1 (N11636, N11625);
nand NAND2 (N11637, N11623, N3782);
xor XOR2 (N11638, N11607, N2562);
nor NOR2 (N11639, N11636, N7159);
xor XOR2 (N11640, N11627, N10827);
nand NAND3 (N11641, N11633, N717, N1947);
or OR2 (N11642, N11621, N2151);
nor NOR3 (N11643, N11641, N1056, N6365);
not NOT1 (N11644, N11635);
and AND4 (N11645, N11643, N3443, N6541, N2000);
or OR2 (N11646, N11637, N3557);
nor NOR3 (N11647, N11640, N6873, N10776);
buf BUF1 (N11648, N11624);
not NOT1 (N11649, N11647);
or OR3 (N11650, N11646, N2114, N7548);
xor XOR2 (N11651, N11650, N8635);
and AND3 (N11652, N11651, N3560, N1396);
nand NAND2 (N11653, N11648, N1368);
nand NAND4 (N11654, N11652, N6311, N3819, N7335);
buf BUF1 (N11655, N11645);
not NOT1 (N11656, N11632);
xor XOR2 (N11657, N11642, N101);
nand NAND3 (N11658, N11644, N1346, N8439);
nand NAND3 (N11659, N11654, N2045, N7325);
and AND3 (N11660, N11653, N7502, N7290);
xor XOR2 (N11661, N11655, N6014);
nand NAND2 (N11662, N11656, N9314);
or OR4 (N11663, N11658, N394, N2640, N10687);
buf BUF1 (N11664, N11649);
xor XOR2 (N11665, N11659, N11012);
not NOT1 (N11666, N11660);
nand NAND3 (N11667, N11662, N7152, N9767);
and AND2 (N11668, N11657, N9207);
xor XOR2 (N11669, N11668, N2331);
not NOT1 (N11670, N11669);
xor XOR2 (N11671, N11634, N10430);
nor NOR3 (N11672, N11638, N4107, N677);
nand NAND2 (N11673, N11671, N10550);
xor XOR2 (N11674, N11673, N1588);
nor NOR3 (N11675, N11639, N2658, N3485);
or OR2 (N11676, N11663, N3729);
buf BUF1 (N11677, N11665);
buf BUF1 (N11678, N11670);
nor NOR3 (N11679, N11661, N3416, N3503);
buf BUF1 (N11680, N11677);
nand NAND4 (N11681, N11666, N11203, N1734, N7756);
or OR2 (N11682, N11678, N8102);
not NOT1 (N11683, N11680);
nor NOR3 (N11684, N11672, N2010, N6604);
nand NAND2 (N11685, N11682, N9011);
nand NAND2 (N11686, N11683, N2654);
not NOT1 (N11687, N11667);
or OR3 (N11688, N11676, N175, N9785);
or OR2 (N11689, N11679, N4739);
and AND3 (N11690, N11674, N6548, N1558);
nor NOR4 (N11691, N11684, N7436, N3994, N7309);
or OR2 (N11692, N11686, N8498);
nor NOR4 (N11693, N11681, N5464, N9630, N11617);
nand NAND3 (N11694, N11692, N10544, N3223);
nand NAND2 (N11695, N11675, N6214);
not NOT1 (N11696, N11664);
nor NOR3 (N11697, N11690, N2862, N2407);
nand NAND3 (N11698, N11687, N10875, N2975);
nor NOR2 (N11699, N11685, N1300);
and AND4 (N11700, N11688, N2358, N9059, N1621);
buf BUF1 (N11701, N11689);
not NOT1 (N11702, N11698);
nand NAND2 (N11703, N11700, N1238);
and AND3 (N11704, N11691, N8114, N10580);
not NOT1 (N11705, N11703);
and AND2 (N11706, N11696, N8630);
nand NAND2 (N11707, N11701, N8847);
nand NAND3 (N11708, N11707, N5518, N7424);
not NOT1 (N11709, N11695);
buf BUF1 (N11710, N11694);
nor NOR2 (N11711, N11708, N10414);
and AND2 (N11712, N11709, N5475);
nand NAND3 (N11713, N11706, N3962, N75);
nor NOR2 (N11714, N11711, N4311);
xor XOR2 (N11715, N11693, N2931);
buf BUF1 (N11716, N11714);
not NOT1 (N11717, N11715);
or OR2 (N11718, N11712, N10362);
and AND4 (N11719, N11699, N2141, N7558, N5229);
nor NOR4 (N11720, N11713, N39, N9205, N2837);
nor NOR3 (N11721, N11705, N1724, N7944);
not NOT1 (N11722, N11710);
or OR3 (N11723, N11719, N4406, N10088);
not NOT1 (N11724, N11723);
or OR4 (N11725, N11704, N7985, N7511, N7191);
nor NOR3 (N11726, N11721, N2609, N6728);
and AND2 (N11727, N11722, N486);
nor NOR2 (N11728, N11720, N11035);
nand NAND2 (N11729, N11728, N2065);
and AND4 (N11730, N11697, N5965, N8421, N387);
or OR2 (N11731, N11726, N209);
nand NAND4 (N11732, N11716, N9790, N3001, N2281);
nor NOR3 (N11733, N11731, N8643, N2738);
or OR2 (N11734, N11724, N4867);
buf BUF1 (N11735, N11732);
and AND3 (N11736, N11733, N5013, N8495);
not NOT1 (N11737, N11727);
nor NOR3 (N11738, N11718, N7157, N6032);
nor NOR2 (N11739, N11702, N8704);
not NOT1 (N11740, N11736);
xor XOR2 (N11741, N11739, N2216);
and AND2 (N11742, N11734, N309);
xor XOR2 (N11743, N11740, N679);
nor NOR4 (N11744, N11738, N2970, N7666, N4196);
xor XOR2 (N11745, N11744, N3041);
nand NAND2 (N11746, N11717, N4268);
or OR2 (N11747, N11743, N2599);
nand NAND2 (N11748, N11735, N7232);
buf BUF1 (N11749, N11747);
nor NOR2 (N11750, N11742, N11309);
buf BUF1 (N11751, N11749);
and AND4 (N11752, N11741, N2550, N761, N7771);
xor XOR2 (N11753, N11745, N2222);
nand NAND3 (N11754, N11748, N6689, N10274);
buf BUF1 (N11755, N11751);
nand NAND2 (N11756, N11750, N7288);
not NOT1 (N11757, N11752);
not NOT1 (N11758, N11755);
xor XOR2 (N11759, N11753, N8902);
nand NAND4 (N11760, N11725, N10446, N3458, N9758);
nor NOR3 (N11761, N11759, N10797, N4792);
xor XOR2 (N11762, N11754, N7030);
nand NAND3 (N11763, N11756, N8490, N972);
xor XOR2 (N11764, N11763, N7785);
buf BUF1 (N11765, N11764);
buf BUF1 (N11766, N11758);
buf BUF1 (N11767, N11737);
not NOT1 (N11768, N11761);
or OR3 (N11769, N11768, N2993, N3839);
or OR3 (N11770, N11766, N11522, N9238);
or OR4 (N11771, N11730, N5035, N11120, N4203);
not NOT1 (N11772, N11746);
nor NOR3 (N11773, N11760, N8749, N4108);
nand NAND2 (N11774, N11773, N6850);
nor NOR2 (N11775, N11765, N5231);
nand NAND3 (N11776, N11774, N5188, N7933);
xor XOR2 (N11777, N11762, N9118);
nor NOR3 (N11778, N11771, N5767, N6478);
and AND4 (N11779, N11775, N5763, N3590, N3513);
xor XOR2 (N11780, N11779, N11059);
and AND2 (N11781, N11776, N6305);
or OR3 (N11782, N11757, N5025, N1581);
nand NAND4 (N11783, N11782, N4282, N3609, N6740);
nor NOR4 (N11784, N11767, N7072, N311, N8048);
buf BUF1 (N11785, N11770);
xor XOR2 (N11786, N11781, N994);
and AND3 (N11787, N11772, N1049, N9008);
nor NOR4 (N11788, N11784, N4076, N9925, N9926);
buf BUF1 (N11789, N11786);
and AND2 (N11790, N11789, N5927);
buf BUF1 (N11791, N11787);
and AND4 (N11792, N11783, N4991, N4575, N6055);
or OR3 (N11793, N11780, N9319, N9138);
xor XOR2 (N11794, N11793, N10555);
not NOT1 (N11795, N11769);
buf BUF1 (N11796, N11792);
or OR3 (N11797, N11729, N3638, N7893);
not NOT1 (N11798, N11796);
and AND3 (N11799, N11798, N10606, N7445);
or OR3 (N11800, N11790, N4, N9078);
buf BUF1 (N11801, N11777);
and AND2 (N11802, N11794, N1281);
and AND4 (N11803, N11800, N2429, N7852, N10411);
xor XOR2 (N11804, N11797, N6616);
not NOT1 (N11805, N11801);
buf BUF1 (N11806, N11795);
or OR2 (N11807, N11799, N4856);
xor XOR2 (N11808, N11803, N2972);
nand NAND4 (N11809, N11778, N2938, N6179, N11105);
not NOT1 (N11810, N11805);
and AND3 (N11811, N11804, N11325, N11713);
buf BUF1 (N11812, N11809);
nand NAND4 (N11813, N11810, N7369, N10749, N8637);
nor NOR3 (N11814, N11785, N7877, N3033);
xor XOR2 (N11815, N11806, N3465);
xor XOR2 (N11816, N11814, N3987);
nand NAND2 (N11817, N11791, N8397);
not NOT1 (N11818, N11816);
not NOT1 (N11819, N11813);
not NOT1 (N11820, N11802);
nand NAND3 (N11821, N11817, N4720, N2501);
or OR4 (N11822, N11807, N7610, N1733, N7907);
not NOT1 (N11823, N11812);
or OR2 (N11824, N11820, N10757);
nor NOR4 (N11825, N11819, N1649, N11431, N11422);
and AND2 (N11826, N11824, N4297);
nand NAND3 (N11827, N11788, N5788, N7290);
nand NAND2 (N11828, N11808, N9180);
or OR2 (N11829, N11821, N2592);
and AND3 (N11830, N11825, N9316, N2437);
nand NAND2 (N11831, N11823, N6497);
buf BUF1 (N11832, N11831);
buf BUF1 (N11833, N11829);
and AND2 (N11834, N11815, N3651);
nand NAND4 (N11835, N11827, N9525, N9068, N7500);
xor XOR2 (N11836, N11818, N2582);
nor NOR3 (N11837, N11828, N529, N5753);
nand NAND4 (N11838, N11833, N5897, N10595, N11783);
xor XOR2 (N11839, N11830, N1367);
buf BUF1 (N11840, N11838);
not NOT1 (N11841, N11834);
nand NAND3 (N11842, N11837, N10008, N891);
and AND2 (N11843, N11842, N6903);
or OR3 (N11844, N11822, N7759, N5282);
and AND3 (N11845, N11840, N8912, N3734);
buf BUF1 (N11846, N11832);
and AND3 (N11847, N11844, N4838, N2966);
nand NAND4 (N11848, N11836, N11756, N1689, N3317);
or OR4 (N11849, N11847, N8304, N946, N827);
and AND4 (N11850, N11811, N1838, N10216, N9777);
nand NAND3 (N11851, N11848, N6253, N6686);
nor NOR4 (N11852, N11851, N2220, N9354, N10862);
xor XOR2 (N11853, N11850, N8802);
not NOT1 (N11854, N11843);
nand NAND3 (N11855, N11845, N9651, N2442);
or OR4 (N11856, N11835, N6178, N5797, N8396);
buf BUF1 (N11857, N11853);
nor NOR4 (N11858, N11856, N907, N604, N10684);
and AND4 (N11859, N11841, N5827, N11836, N5872);
xor XOR2 (N11860, N11859, N10733);
not NOT1 (N11861, N11849);
buf BUF1 (N11862, N11854);
buf BUF1 (N11863, N11860);
and AND3 (N11864, N11863, N5346, N1351);
nand NAND3 (N11865, N11826, N9786, N3673);
nor NOR4 (N11866, N11858, N10982, N10810, N2586);
xor XOR2 (N11867, N11839, N4205);
not NOT1 (N11868, N11866);
nand NAND2 (N11869, N11852, N10895);
buf BUF1 (N11870, N11855);
buf BUF1 (N11871, N11846);
nand NAND4 (N11872, N11861, N1455, N2490, N2304);
or OR4 (N11873, N11864, N9586, N7903, N2254);
and AND3 (N11874, N11857, N7347, N5990);
xor XOR2 (N11875, N11868, N7252);
nor NOR2 (N11876, N11872, N6789);
and AND4 (N11877, N11865, N3402, N6649, N9365);
xor XOR2 (N11878, N11870, N1512);
xor XOR2 (N11879, N11869, N9513);
not NOT1 (N11880, N11874);
xor XOR2 (N11881, N11875, N6825);
nor NOR4 (N11882, N11862, N737, N881, N8473);
buf BUF1 (N11883, N11867);
not NOT1 (N11884, N11876);
nand NAND4 (N11885, N11883, N5016, N7358, N10440);
xor XOR2 (N11886, N11884, N2859);
not NOT1 (N11887, N11880);
and AND2 (N11888, N11878, N4636);
nand NAND3 (N11889, N11879, N11836, N2853);
not NOT1 (N11890, N11889);
nor NOR2 (N11891, N11871, N7023);
or OR4 (N11892, N11881, N10900, N6420, N3263);
xor XOR2 (N11893, N11887, N294);
and AND4 (N11894, N11877, N11218, N5746, N8533);
nor NOR4 (N11895, N11894, N1559, N11244, N2480);
nand NAND3 (N11896, N11886, N5795, N4485);
buf BUF1 (N11897, N11893);
not NOT1 (N11898, N11885);
not NOT1 (N11899, N11896);
nor NOR3 (N11900, N11899, N1257, N4582);
xor XOR2 (N11901, N11900, N9850);
buf BUF1 (N11902, N11898);
buf BUF1 (N11903, N11892);
not NOT1 (N11904, N11890);
and AND4 (N11905, N11904, N949, N728, N6648);
and AND2 (N11906, N11901, N1831);
nand NAND2 (N11907, N11905, N9628);
nand NAND3 (N11908, N11903, N11907, N5762);
buf BUF1 (N11909, N4037);
xor XOR2 (N11910, N11882, N7591);
not NOT1 (N11911, N11888);
not NOT1 (N11912, N11910);
xor XOR2 (N11913, N11897, N2803);
not NOT1 (N11914, N11908);
and AND3 (N11915, N11891, N9794, N10896);
nor NOR2 (N11916, N11911, N6610);
xor XOR2 (N11917, N11916, N1953);
nand NAND4 (N11918, N11914, N1216, N2467, N6123);
not NOT1 (N11919, N11918);
nand NAND3 (N11920, N11912, N8117, N3476);
nor NOR4 (N11921, N11895, N10147, N2386, N11472);
and AND4 (N11922, N11902, N924, N11552, N631);
not NOT1 (N11923, N11922);
not NOT1 (N11924, N11921);
not NOT1 (N11925, N11909);
or OR2 (N11926, N11923, N528);
not NOT1 (N11927, N11906);
not NOT1 (N11928, N11917);
or OR2 (N11929, N11919, N831);
or OR4 (N11930, N11915, N11532, N11919, N518);
xor XOR2 (N11931, N11920, N5110);
nand NAND4 (N11932, N11926, N1550, N9801, N2059);
or OR2 (N11933, N11873, N7833);
buf BUF1 (N11934, N11931);
nor NOR2 (N11935, N11934, N9933);
not NOT1 (N11936, N11930);
nor NOR3 (N11937, N11913, N8886, N5640);
or OR4 (N11938, N11936, N8744, N4109, N6396);
or OR2 (N11939, N11924, N8095);
xor XOR2 (N11940, N11929, N4260);
nand NAND2 (N11941, N11937, N4373);
xor XOR2 (N11942, N11935, N8218);
and AND2 (N11943, N11933, N3699);
nand NAND3 (N11944, N11925, N1540, N9215);
not NOT1 (N11945, N11942);
buf BUF1 (N11946, N11944);
xor XOR2 (N11947, N11928, N9688);
nand NAND4 (N11948, N11940, N7632, N7206, N9993);
not NOT1 (N11949, N11939);
not NOT1 (N11950, N11941);
not NOT1 (N11951, N11938);
nor NOR3 (N11952, N11945, N1198, N536);
and AND2 (N11953, N11943, N7532);
xor XOR2 (N11954, N11951, N8923);
buf BUF1 (N11955, N11932);
buf BUF1 (N11956, N11952);
xor XOR2 (N11957, N11947, N8714);
buf BUF1 (N11958, N11953);
nor NOR2 (N11959, N11948, N1374);
xor XOR2 (N11960, N11954, N1548);
nor NOR3 (N11961, N11950, N11852, N9964);
and AND4 (N11962, N11946, N5337, N693, N1309);
nand NAND2 (N11963, N11955, N3602);
nand NAND3 (N11964, N11963, N1963, N3663);
and AND3 (N11965, N11960, N10330, N7995);
not NOT1 (N11966, N11959);
nand NAND3 (N11967, N11958, N8900, N9886);
or OR4 (N11968, N11961, N5677, N8596, N2872);
nand NAND4 (N11969, N11927, N2439, N5407, N159);
xor XOR2 (N11970, N11962, N1760);
buf BUF1 (N11971, N11969);
xor XOR2 (N11972, N11966, N4303);
xor XOR2 (N11973, N11970, N3152);
and AND2 (N11974, N11964, N1869);
and AND3 (N11975, N11971, N8529, N11092);
and AND2 (N11976, N11974, N10405);
nand NAND2 (N11977, N11965, N11752);
and AND4 (N11978, N11957, N4511, N1627, N10342);
xor XOR2 (N11979, N11949, N11186);
nor NOR3 (N11980, N11967, N8619, N5551);
nand NAND2 (N11981, N11978, N5774);
xor XOR2 (N11982, N11977, N5175);
buf BUF1 (N11983, N11968);
and AND2 (N11984, N11981, N7822);
or OR4 (N11985, N11972, N8300, N11574, N9904);
not NOT1 (N11986, N11976);
xor XOR2 (N11987, N11984, N2869);
xor XOR2 (N11988, N11982, N3187);
buf BUF1 (N11989, N11988);
not NOT1 (N11990, N11985);
buf BUF1 (N11991, N11980);
and AND4 (N11992, N11986, N6260, N11023, N10847);
or OR3 (N11993, N11990, N8868, N6033);
not NOT1 (N11994, N11975);
not NOT1 (N11995, N11979);
nand NAND4 (N11996, N11995, N905, N4345, N10507);
or OR4 (N11997, N11987, N10428, N11305, N5152);
buf BUF1 (N11998, N11983);
buf BUF1 (N11999, N11973);
not NOT1 (N12000, N11956);
nand NAND2 (N12001, N11994, N2082);
buf BUF1 (N12002, N11998);
not NOT1 (N12003, N11996);
and AND4 (N12004, N11993, N1590, N8259, N7267);
nor NOR4 (N12005, N11989, N4, N196, N8125);
xor XOR2 (N12006, N12000, N3279);
or OR4 (N12007, N12003, N6117, N10184, N1148);
nor NOR2 (N12008, N11992, N2300);
nand NAND3 (N12009, N11991, N3560, N564);
xor XOR2 (N12010, N12008, N7893);
and AND4 (N12011, N12002, N7723, N8922, N5120);
and AND3 (N12012, N12007, N10443, N6503);
xor XOR2 (N12013, N12009, N6712);
not NOT1 (N12014, N12005);
or OR2 (N12015, N12001, N4559);
nor NOR4 (N12016, N12004, N2436, N2255, N9145);
not NOT1 (N12017, N12013);
nor NOR4 (N12018, N12010, N7422, N2423, N9861);
buf BUF1 (N12019, N12015);
or OR3 (N12020, N12011, N5868, N7744);
or OR2 (N12021, N12019, N1296);
nor NOR4 (N12022, N12018, N201, N3230, N8428);
nor NOR4 (N12023, N12020, N4542, N8722, N10052);
nand NAND2 (N12024, N12017, N7152);
not NOT1 (N12025, N12014);
nand NAND2 (N12026, N11997, N1054);
xor XOR2 (N12027, N12022, N11580);
not NOT1 (N12028, N12024);
buf BUF1 (N12029, N12016);
buf BUF1 (N12030, N12025);
and AND4 (N12031, N11999, N10059, N4106, N6630);
and AND2 (N12032, N12031, N9510);
nor NOR3 (N12033, N12026, N4465, N3967);
buf BUF1 (N12034, N12012);
buf BUF1 (N12035, N12030);
nor NOR4 (N12036, N12027, N8771, N3695, N3743);
not NOT1 (N12037, N12034);
buf BUF1 (N12038, N12032);
buf BUF1 (N12039, N12021);
not NOT1 (N12040, N12029);
nand NAND4 (N12041, N12023, N580, N3131, N6636);
not NOT1 (N12042, N12036);
not NOT1 (N12043, N12038);
and AND2 (N12044, N12042, N10412);
not NOT1 (N12045, N12039);
or OR3 (N12046, N12035, N10321, N1335);
buf BUF1 (N12047, N12041);
nor NOR2 (N12048, N12028, N156);
not NOT1 (N12049, N12037);
and AND4 (N12050, N12046, N5912, N11018, N7149);
xor XOR2 (N12051, N12006, N11875);
xor XOR2 (N12052, N12033, N995);
or OR4 (N12053, N12050, N8620, N11182, N11562);
and AND2 (N12054, N12044, N9689);
and AND4 (N12055, N12053, N2384, N2916, N2453);
or OR3 (N12056, N12048, N2647, N10719);
or OR4 (N12057, N12047, N5010, N4916, N3777);
xor XOR2 (N12058, N12043, N906);
buf BUF1 (N12059, N12057);
not NOT1 (N12060, N12040);
buf BUF1 (N12061, N12056);
or OR2 (N12062, N12052, N379);
nor NOR4 (N12063, N12049, N2832, N4228, N3757);
or OR4 (N12064, N12061, N6368, N3769, N130);
or OR2 (N12065, N12063, N3784);
xor XOR2 (N12066, N12062, N1651);
or OR4 (N12067, N12051, N3057, N10187, N932);
nand NAND4 (N12068, N12054, N7371, N4605, N7040);
nand NAND3 (N12069, N12058, N4996, N6279);
nor NOR4 (N12070, N12060, N8183, N11928, N3283);
and AND4 (N12071, N12045, N9115, N3758, N785);
not NOT1 (N12072, N12069);
nand NAND3 (N12073, N12068, N156, N9255);
xor XOR2 (N12074, N12072, N5899);
and AND2 (N12075, N12067, N4066);
nand NAND2 (N12076, N12070, N11317);
nor NOR4 (N12077, N12074, N6818, N5177, N8155);
nand NAND4 (N12078, N12064, N4718, N2048, N3428);
not NOT1 (N12079, N12065);
xor XOR2 (N12080, N12071, N2503);
nand NAND3 (N12081, N12079, N4400, N8259);
nand NAND4 (N12082, N12081, N7494, N9562, N1578);
nor NOR3 (N12083, N12077, N9367, N8362);
or OR2 (N12084, N12073, N10892);
nor NOR3 (N12085, N12082, N3995, N1237);
buf BUF1 (N12086, N12075);
nand NAND3 (N12087, N12078, N4797, N5699);
and AND4 (N12088, N12085, N1013, N4172, N5329);
nand NAND3 (N12089, N12087, N11073, N8423);
nand NAND3 (N12090, N12084, N4119, N7383);
nor NOR2 (N12091, N12083, N10173);
and AND4 (N12092, N12055, N5780, N8092, N11189);
buf BUF1 (N12093, N12089);
xor XOR2 (N12094, N12076, N9257);
nor NOR2 (N12095, N12092, N11316);
and AND3 (N12096, N12088, N8252, N6988);
not NOT1 (N12097, N12090);
and AND2 (N12098, N12086, N10196);
not NOT1 (N12099, N12093);
and AND2 (N12100, N12099, N10660);
nor NOR4 (N12101, N12091, N606, N11855, N3322);
nor NOR4 (N12102, N12094, N9875, N4641, N10581);
nand NAND2 (N12103, N12096, N10449);
xor XOR2 (N12104, N12097, N9866);
or OR4 (N12105, N12066, N1245, N7382, N7003);
not NOT1 (N12106, N12101);
nor NOR3 (N12107, N12095, N11709, N9725);
nand NAND4 (N12108, N12100, N3965, N2077, N2878);
xor XOR2 (N12109, N12105, N453);
and AND2 (N12110, N12109, N11247);
or OR2 (N12111, N12102, N638);
nand NAND4 (N12112, N12103, N9041, N120, N1628);
and AND2 (N12113, N12104, N10619);
and AND2 (N12114, N12113, N6790);
nor NOR2 (N12115, N12108, N10964);
xor XOR2 (N12116, N12080, N1206);
not NOT1 (N12117, N12110);
and AND2 (N12118, N12107, N5186);
nand NAND4 (N12119, N12118, N6763, N6442, N3066);
and AND2 (N12120, N12116, N2107);
or OR4 (N12121, N12059, N6118, N1346, N4312);
nor NOR2 (N12122, N12121, N10158);
nor NOR2 (N12123, N12098, N2847);
or OR3 (N12124, N12123, N10819, N2860);
not NOT1 (N12125, N12112);
or OR4 (N12126, N12122, N7438, N10495, N6341);
or OR3 (N12127, N12124, N352, N7465);
or OR2 (N12128, N12114, N2614);
and AND2 (N12129, N12111, N734);
nor NOR2 (N12130, N12120, N5609);
nor NOR2 (N12131, N12106, N8680);
and AND2 (N12132, N12128, N1483);
or OR4 (N12133, N12126, N3653, N4375, N10351);
not NOT1 (N12134, N12117);
buf BUF1 (N12135, N12132);
and AND4 (N12136, N12134, N982, N2656, N2262);
and AND2 (N12137, N12125, N5659);
nor NOR4 (N12138, N12137, N5601, N7181, N2054);
not NOT1 (N12139, N12136);
and AND3 (N12140, N12115, N9773, N1238);
nor NOR4 (N12141, N12131, N10370, N10098, N8106);
not NOT1 (N12142, N12130);
xor XOR2 (N12143, N12129, N2315);
xor XOR2 (N12144, N12141, N5759);
nand NAND2 (N12145, N12140, N6986);
not NOT1 (N12146, N12119);
buf BUF1 (N12147, N12127);
buf BUF1 (N12148, N12133);
or OR4 (N12149, N12146, N9807, N6596, N8649);
nand NAND4 (N12150, N12142, N11783, N4235, N4323);
and AND3 (N12151, N12139, N9960, N2098);
nand NAND2 (N12152, N12150, N3513);
and AND3 (N12153, N12138, N7189, N4215);
or OR3 (N12154, N12135, N1455, N2152);
not NOT1 (N12155, N12149);
or OR4 (N12156, N12153, N7516, N6398, N5607);
nor NOR2 (N12157, N12143, N4295);
and AND2 (N12158, N12151, N6254);
or OR3 (N12159, N12158, N2994, N302);
xor XOR2 (N12160, N12144, N5762);
nand NAND2 (N12161, N12152, N1786);
or OR3 (N12162, N12148, N2661, N10846);
nor NOR4 (N12163, N12162, N7055, N5161, N3626);
or OR3 (N12164, N12145, N1925, N1542);
nand NAND2 (N12165, N12156, N2879);
not NOT1 (N12166, N12157);
buf BUF1 (N12167, N12165);
buf BUF1 (N12168, N12167);
xor XOR2 (N12169, N12154, N496);
or OR3 (N12170, N12147, N6992, N10502);
and AND2 (N12171, N12155, N9303);
xor XOR2 (N12172, N12166, N11277);
or OR4 (N12173, N12159, N4818, N10085, N10205);
and AND3 (N12174, N12160, N1871, N1893);
xor XOR2 (N12175, N12173, N8169);
nand NAND3 (N12176, N12172, N3585, N12163);
nand NAND4 (N12177, N7504, N5936, N10582, N10807);
nor NOR2 (N12178, N12161, N6704);
or OR4 (N12179, N12177, N5478, N7797, N4455);
or OR2 (N12180, N12179, N5915);
buf BUF1 (N12181, N12174);
not NOT1 (N12182, N12169);
buf BUF1 (N12183, N12176);
and AND3 (N12184, N12171, N6923, N5008);
or OR3 (N12185, N12183, N6725, N6106);
or OR4 (N12186, N12170, N7685, N4155, N10577);
or OR3 (N12187, N12181, N11956, N8610);
buf BUF1 (N12188, N12168);
nor NOR2 (N12189, N12187, N9942);
buf BUF1 (N12190, N12186);
nand NAND3 (N12191, N12178, N6191, N1072);
nor NOR3 (N12192, N12184, N3989, N1394);
nand NAND4 (N12193, N12180, N7254, N6626, N10486);
and AND2 (N12194, N12188, N5267);
buf BUF1 (N12195, N12185);
and AND3 (N12196, N12189, N5185, N3972);
nor NOR3 (N12197, N12194, N9040, N9198);
nor NOR4 (N12198, N12164, N8502, N10880, N380);
and AND4 (N12199, N12191, N2228, N10898, N7782);
or OR4 (N12200, N12182, N4330, N1408, N7720);
or OR3 (N12201, N12200, N8380, N8617);
buf BUF1 (N12202, N12190);
buf BUF1 (N12203, N12196);
buf BUF1 (N12204, N12203);
or OR4 (N12205, N12197, N4920, N8068, N7751);
nor NOR3 (N12206, N12205, N8542, N1601);
and AND4 (N12207, N12199, N9351, N3102, N404);
or OR4 (N12208, N12201, N4838, N960, N5175);
nand NAND3 (N12209, N12193, N2021, N9419);
not NOT1 (N12210, N12209);
and AND3 (N12211, N12208, N5692, N6571);
and AND4 (N12212, N12206, N3318, N298, N697);
nand NAND4 (N12213, N12198, N11387, N9905, N9958);
xor XOR2 (N12214, N12192, N7500);
nor NOR3 (N12215, N12214, N7805, N10361);
nor NOR2 (N12216, N12202, N6889);
nor NOR4 (N12217, N12215, N5531, N6714, N5982);
nand NAND4 (N12218, N12216, N12093, N8198, N8365);
and AND3 (N12219, N12211, N9335, N10727);
or OR3 (N12220, N12207, N4424, N10062);
or OR2 (N12221, N12212, N3168);
buf BUF1 (N12222, N12213);
nand NAND2 (N12223, N12218, N1181);
and AND2 (N12224, N12195, N2947);
and AND4 (N12225, N12224, N8001, N8605, N10748);
buf BUF1 (N12226, N12222);
or OR2 (N12227, N12217, N9543);
and AND2 (N12228, N12204, N12009);
xor XOR2 (N12229, N12219, N11483);
xor XOR2 (N12230, N12229, N4660);
not NOT1 (N12231, N12225);
and AND4 (N12232, N12220, N9253, N7839, N10807);
nor NOR4 (N12233, N12223, N11389, N2632, N10514);
buf BUF1 (N12234, N12228);
buf BUF1 (N12235, N12227);
nor NOR2 (N12236, N12232, N4730);
nand NAND2 (N12237, N12235, N5615);
xor XOR2 (N12238, N12236, N8810);
and AND4 (N12239, N12221, N9763, N640, N9200);
xor XOR2 (N12240, N12226, N1262);
xor XOR2 (N12241, N12239, N8349);
nor NOR2 (N12242, N12233, N1390);
not NOT1 (N12243, N12175);
and AND3 (N12244, N12241, N1008, N5556);
nor NOR2 (N12245, N12237, N9578);
xor XOR2 (N12246, N12243, N8656);
and AND2 (N12247, N12246, N7969);
xor XOR2 (N12248, N12230, N8963);
not NOT1 (N12249, N12238);
and AND4 (N12250, N12245, N3817, N6631, N11049);
or OR2 (N12251, N12231, N8523);
buf BUF1 (N12252, N12244);
buf BUF1 (N12253, N12234);
nor NOR3 (N12254, N12248, N8744, N3537);
not NOT1 (N12255, N12250);
or OR4 (N12256, N12210, N10492, N10731, N8765);
not NOT1 (N12257, N12253);
not NOT1 (N12258, N12240);
xor XOR2 (N12259, N12255, N446);
buf BUF1 (N12260, N12251);
or OR2 (N12261, N12260, N7532);
and AND2 (N12262, N12252, N7305);
nand NAND3 (N12263, N12257, N3005, N6318);
buf BUF1 (N12264, N12249);
and AND2 (N12265, N12259, N11775);
xor XOR2 (N12266, N12242, N6076);
nand NAND2 (N12267, N12247, N68);
buf BUF1 (N12268, N12267);
xor XOR2 (N12269, N12265, N6368);
nor NOR4 (N12270, N12269, N8334, N5506, N7086);
buf BUF1 (N12271, N12262);
not NOT1 (N12272, N12266);
and AND3 (N12273, N12263, N6635, N10039);
xor XOR2 (N12274, N12270, N8760);
nor NOR3 (N12275, N12261, N4152, N7710);
nand NAND3 (N12276, N12254, N5454, N9535);
nor NOR3 (N12277, N12264, N8720, N11682);
nor NOR3 (N12278, N12268, N7322, N10809);
or OR3 (N12279, N12278, N6630, N9248);
nand NAND3 (N12280, N12271, N1581, N2813);
buf BUF1 (N12281, N12274);
nor NOR2 (N12282, N12281, N10380);
and AND4 (N12283, N12280, N5713, N7747, N8553);
nor NOR3 (N12284, N12272, N4093, N4261);
or OR2 (N12285, N12275, N477);
not NOT1 (N12286, N12277);
or OR2 (N12287, N12256, N2272);
nand NAND4 (N12288, N12273, N3954, N10813, N7396);
and AND2 (N12289, N12279, N3048);
not NOT1 (N12290, N12276);
nand NAND3 (N12291, N12287, N9582, N7637);
and AND3 (N12292, N12285, N9808, N2461);
or OR3 (N12293, N12282, N11513, N2629);
and AND2 (N12294, N12258, N10116);
nor NOR4 (N12295, N12290, N694, N10310, N9614);
nor NOR3 (N12296, N12284, N2763, N1387);
xor XOR2 (N12297, N12286, N6743);
not NOT1 (N12298, N12283);
nand NAND3 (N12299, N12293, N5307, N1007);
nor NOR4 (N12300, N12299, N10763, N11817, N10764);
nor NOR3 (N12301, N12292, N10164, N1910);
buf BUF1 (N12302, N12301);
not NOT1 (N12303, N12300);
or OR2 (N12304, N12296, N10018);
not NOT1 (N12305, N12288);
xor XOR2 (N12306, N12294, N2641);
or OR3 (N12307, N12289, N10963, N6709);
nand NAND4 (N12308, N12297, N6504, N10259, N315);
buf BUF1 (N12309, N12302);
xor XOR2 (N12310, N12309, N7262);
xor XOR2 (N12311, N12310, N1924);
xor XOR2 (N12312, N12306, N6430);
nor NOR2 (N12313, N12305, N5747);
xor XOR2 (N12314, N12313, N4119);
buf BUF1 (N12315, N12303);
nand NAND2 (N12316, N12298, N1806);
or OR3 (N12317, N12307, N9950, N542);
xor XOR2 (N12318, N12311, N8323);
nand NAND3 (N12319, N12295, N2851, N5705);
or OR4 (N12320, N12312, N8411, N4485, N10157);
xor XOR2 (N12321, N12304, N2494);
and AND2 (N12322, N12291, N7534);
nor NOR4 (N12323, N12314, N7434, N8783, N4803);
buf BUF1 (N12324, N12323);
and AND3 (N12325, N12322, N10185, N8456);
or OR4 (N12326, N12317, N4928, N7581, N12042);
nor NOR3 (N12327, N12316, N2272, N792);
xor XOR2 (N12328, N12315, N11602);
and AND3 (N12329, N12327, N5839, N1462);
nand NAND4 (N12330, N12320, N1311, N11796, N9403);
xor XOR2 (N12331, N12326, N5181);
and AND2 (N12332, N12325, N7512);
or OR2 (N12333, N12330, N11368);
and AND4 (N12334, N12329, N11519, N5560, N3419);
nand NAND4 (N12335, N12333, N774, N4293, N5733);
nor NOR3 (N12336, N12332, N8656, N9816);
buf BUF1 (N12337, N12321);
or OR3 (N12338, N12336, N4077, N3173);
or OR2 (N12339, N12335, N5034);
nor NOR4 (N12340, N12334, N1801, N8927, N5564);
xor XOR2 (N12341, N12340, N6809);
buf BUF1 (N12342, N12341);
buf BUF1 (N12343, N12324);
and AND3 (N12344, N12319, N9288, N2403);
nand NAND3 (N12345, N12339, N5332, N2482);
nor NOR2 (N12346, N12345, N11276);
and AND3 (N12347, N12346, N6914, N6183);
nor NOR3 (N12348, N12328, N9705, N3954);
nor NOR4 (N12349, N12347, N6124, N11226, N7758);
and AND3 (N12350, N12349, N6708, N8209);
not NOT1 (N12351, N12337);
and AND3 (N12352, N12351, N11505, N10191);
nor NOR2 (N12353, N12344, N453);
nand NAND2 (N12354, N12350, N5702);
and AND2 (N12355, N12348, N817);
nor NOR3 (N12356, N12353, N9132, N4412);
not NOT1 (N12357, N12352);
buf BUF1 (N12358, N12343);
and AND4 (N12359, N12331, N189, N10442, N11915);
and AND4 (N12360, N12318, N7955, N4551, N2531);
buf BUF1 (N12361, N12357);
and AND3 (N12362, N12359, N10713, N6368);
not NOT1 (N12363, N12308);
nand NAND2 (N12364, N12360, N5186);
and AND2 (N12365, N12363, N10643);
buf BUF1 (N12366, N12361);
and AND3 (N12367, N12342, N5699, N3289);
nand NAND2 (N12368, N12355, N8588);
and AND4 (N12369, N12358, N9757, N7564, N8914);
or OR3 (N12370, N12368, N4589, N4353);
and AND2 (N12371, N12366, N9169);
xor XOR2 (N12372, N12369, N1545);
xor XOR2 (N12373, N12354, N8507);
or OR2 (N12374, N12356, N1300);
xor XOR2 (N12375, N12365, N6885);
xor XOR2 (N12376, N12372, N1089);
or OR3 (N12377, N12364, N5356, N7033);
or OR3 (N12378, N12374, N7945, N6786);
nor NOR4 (N12379, N12377, N7062, N10056, N11004);
or OR4 (N12380, N12376, N4027, N9345, N1170);
and AND2 (N12381, N12362, N666);
xor XOR2 (N12382, N12380, N467);
nand NAND3 (N12383, N12375, N6948, N10909);
buf BUF1 (N12384, N12370);
xor XOR2 (N12385, N12383, N12184);
xor XOR2 (N12386, N12381, N2928);
nor NOR4 (N12387, N12371, N8900, N9, N4090);
nand NAND4 (N12388, N12385, N662, N8062, N41);
not NOT1 (N12389, N12386);
xor XOR2 (N12390, N12388, N6386);
and AND3 (N12391, N12387, N8338, N4075);
and AND2 (N12392, N12384, N10650);
not NOT1 (N12393, N12389);
nor NOR3 (N12394, N12390, N5083, N6719);
buf BUF1 (N12395, N12338);
xor XOR2 (N12396, N12395, N4245);
xor XOR2 (N12397, N12367, N9801);
xor XOR2 (N12398, N12397, N9158);
buf BUF1 (N12399, N12378);
xor XOR2 (N12400, N12391, N4219);
buf BUF1 (N12401, N12392);
not NOT1 (N12402, N12379);
not NOT1 (N12403, N12393);
nor NOR3 (N12404, N12401, N4274, N3082);
buf BUF1 (N12405, N12400);
xor XOR2 (N12406, N12382, N12304);
xor XOR2 (N12407, N12396, N11703);
buf BUF1 (N12408, N12398);
buf BUF1 (N12409, N12399);
not NOT1 (N12410, N12402);
or OR3 (N12411, N12403, N6887, N825);
nor NOR3 (N12412, N12404, N6171, N2431);
not NOT1 (N12413, N12410);
not NOT1 (N12414, N12373);
buf BUF1 (N12415, N12414);
nor NOR4 (N12416, N12415, N7523, N9437, N10866);
xor XOR2 (N12417, N12409, N8452);
nor NOR3 (N12418, N12406, N970, N9612);
and AND2 (N12419, N12408, N9202);
and AND3 (N12420, N12417, N7980, N4419);
nor NOR2 (N12421, N12418, N9720);
and AND2 (N12422, N12394, N765);
nor NOR2 (N12423, N12422, N6633);
and AND2 (N12424, N12421, N9307);
nor NOR4 (N12425, N12411, N9274, N11722, N6751);
and AND3 (N12426, N12420, N11205, N3993);
nand NAND2 (N12427, N12405, N12289);
nand NAND2 (N12428, N12412, N1989);
or OR3 (N12429, N12423, N8172, N7012);
not NOT1 (N12430, N12429);
nand NAND4 (N12431, N12427, N5074, N6557, N4603);
xor XOR2 (N12432, N12407, N10214);
nor NOR3 (N12433, N12424, N2760, N2787);
buf BUF1 (N12434, N12432);
and AND4 (N12435, N12434, N5381, N12409, N11197);
xor XOR2 (N12436, N12430, N6822);
buf BUF1 (N12437, N12416);
and AND3 (N12438, N12431, N882, N10806);
or OR2 (N12439, N12433, N4054);
not NOT1 (N12440, N12438);
not NOT1 (N12441, N12440);
nor NOR3 (N12442, N12437, N939, N9326);
xor XOR2 (N12443, N12425, N11410);
xor XOR2 (N12444, N12419, N10853);
nor NOR3 (N12445, N12428, N10087, N7276);
or OR4 (N12446, N12444, N1926, N718, N605);
or OR2 (N12447, N12436, N599);
buf BUF1 (N12448, N12426);
nand NAND4 (N12449, N12413, N791, N12362, N462);
nand NAND3 (N12450, N12448, N9691, N4133);
nand NAND4 (N12451, N12445, N1903, N6045, N6982);
nor NOR3 (N12452, N12439, N2825, N9628);
nor NOR2 (N12453, N12435, N8488);
xor XOR2 (N12454, N12441, N6011);
or OR3 (N12455, N12449, N2503, N5740);
or OR2 (N12456, N12453, N12189);
buf BUF1 (N12457, N12451);
and AND4 (N12458, N12457, N4560, N9670, N8768);
nor NOR3 (N12459, N12458, N7264, N8476);
nand NAND4 (N12460, N12459, N11315, N7422, N5353);
xor XOR2 (N12461, N12446, N11306);
nor NOR3 (N12462, N12443, N3381, N4722);
and AND2 (N12463, N12461, N11543);
and AND3 (N12464, N12447, N3158, N11034);
nand NAND3 (N12465, N12452, N1468, N150);
nor NOR2 (N12466, N12450, N8239);
buf BUF1 (N12467, N12455);
buf BUF1 (N12468, N12456);
buf BUF1 (N12469, N12467);
nor NOR3 (N12470, N12469, N8368, N7939);
nand NAND4 (N12471, N12454, N6627, N44, N10318);
and AND2 (N12472, N12468, N4049);
or OR2 (N12473, N12471, N5977);
and AND3 (N12474, N12442, N395, N5295);
or OR3 (N12475, N12465, N1376, N519);
xor XOR2 (N12476, N12475, N10082);
buf BUF1 (N12477, N12470);
not NOT1 (N12478, N12473);
nand NAND4 (N12479, N12474, N888, N9462, N3926);
nand NAND4 (N12480, N12463, N9202, N11413, N11726);
buf BUF1 (N12481, N12462);
and AND4 (N12482, N12478, N3364, N1230, N11809);
not NOT1 (N12483, N12479);
not NOT1 (N12484, N12483);
or OR3 (N12485, N12477, N3607, N9896);
nor NOR2 (N12486, N12485, N4940);
or OR2 (N12487, N12481, N3151);
nand NAND4 (N12488, N12472, N5841, N9918, N838);
buf BUF1 (N12489, N12487);
nor NOR2 (N12490, N12480, N2227);
and AND3 (N12491, N12482, N11504, N11001);
nand NAND3 (N12492, N12484, N3597, N11546);
and AND4 (N12493, N12460, N7502, N11204, N1751);
not NOT1 (N12494, N12466);
xor XOR2 (N12495, N12488, N2550);
or OR4 (N12496, N12493, N10084, N4005, N5877);
and AND4 (N12497, N12495, N2938, N11951, N2936);
or OR4 (N12498, N12497, N9010, N7756, N5534);
nor NOR2 (N12499, N12464, N4497);
and AND2 (N12500, N12491, N8191);
not NOT1 (N12501, N12490);
buf BUF1 (N12502, N12500);
or OR3 (N12503, N12502, N8135, N8803);
nor NOR2 (N12504, N12492, N552);
or OR2 (N12505, N12498, N12339);
nor NOR2 (N12506, N12501, N9042);
or OR2 (N12507, N12504, N69);
not NOT1 (N12508, N12505);
nand NAND2 (N12509, N12489, N4776);
xor XOR2 (N12510, N12496, N8715);
buf BUF1 (N12511, N12507);
or OR4 (N12512, N12499, N12151, N11615, N4848);
xor XOR2 (N12513, N12512, N7615);
nor NOR4 (N12514, N12510, N10770, N5773, N373);
not NOT1 (N12515, N12508);
nor NOR2 (N12516, N12486, N6201);
nand NAND3 (N12517, N12503, N1110, N6337);
or OR4 (N12518, N12511, N6954, N2833, N4907);
nor NOR4 (N12519, N12509, N2915, N1453, N11387);
nor NOR3 (N12520, N12476, N5999, N25);
nor NOR3 (N12521, N12519, N12218, N6337);
or OR2 (N12522, N12513, N11173);
nor NOR2 (N12523, N12521, N6775);
nand NAND2 (N12524, N12506, N3122);
or OR3 (N12525, N12522, N2668, N1799);
nor NOR3 (N12526, N12520, N11365, N7279);
or OR4 (N12527, N12518, N3956, N2618, N4473);
buf BUF1 (N12528, N12494);
not NOT1 (N12529, N12516);
nand NAND3 (N12530, N12528, N5598, N3576);
nor NOR3 (N12531, N12523, N7520, N8403);
nor NOR3 (N12532, N12530, N5437, N10227);
or OR4 (N12533, N12525, N9449, N3894, N10718);
or OR2 (N12534, N12533, N7580);
nor NOR2 (N12535, N12532, N12352);
buf BUF1 (N12536, N12517);
nand NAND2 (N12537, N12534, N4235);
xor XOR2 (N12538, N12527, N5598);
or OR2 (N12539, N12514, N5337);
buf BUF1 (N12540, N12536);
and AND3 (N12541, N12539, N7634, N7691);
or OR3 (N12542, N12535, N11306, N9616);
or OR4 (N12543, N12531, N4313, N3850, N10365);
buf BUF1 (N12544, N12543);
buf BUF1 (N12545, N12540);
xor XOR2 (N12546, N12524, N815);
and AND2 (N12547, N12529, N8587);
and AND3 (N12548, N12526, N8879, N11229);
nor NOR2 (N12549, N12515, N4806);
and AND3 (N12550, N12548, N9345, N5683);
nand NAND4 (N12551, N12546, N3616, N1426, N9000);
nor NOR2 (N12552, N12538, N264);
xor XOR2 (N12553, N12549, N9401);
nand NAND2 (N12554, N12544, N856);
nor NOR3 (N12555, N12545, N1440, N6025);
nor NOR2 (N12556, N12554, N10640);
and AND4 (N12557, N12556, N211, N12551, N8326);
and AND2 (N12558, N12279, N4328);
and AND2 (N12559, N12547, N7700);
not NOT1 (N12560, N12550);
buf BUF1 (N12561, N12542);
and AND2 (N12562, N12553, N2380);
nor NOR3 (N12563, N12555, N8355, N2483);
and AND3 (N12564, N12560, N3414, N786);
and AND3 (N12565, N12564, N10699, N2182);
or OR2 (N12566, N12537, N5367);
buf BUF1 (N12567, N12566);
nand NAND3 (N12568, N12552, N538, N8030);
not NOT1 (N12569, N12558);
buf BUF1 (N12570, N12557);
or OR3 (N12571, N12559, N5204, N22);
or OR2 (N12572, N12570, N10878);
or OR4 (N12573, N12562, N11913, N2277, N2935);
nand NAND3 (N12574, N12563, N744, N3354);
nor NOR2 (N12575, N12569, N4076);
nor NOR3 (N12576, N12565, N743, N4413);
not NOT1 (N12577, N12575);
not NOT1 (N12578, N12568);
and AND2 (N12579, N12574, N976);
nor NOR4 (N12580, N12577, N10809, N4843, N12316);
not NOT1 (N12581, N12541);
xor XOR2 (N12582, N12579, N9960);
nor NOR4 (N12583, N12576, N4037, N10330, N11158);
nor NOR4 (N12584, N12567, N4596, N10911, N3547);
buf BUF1 (N12585, N12573);
buf BUF1 (N12586, N12561);
nand NAND3 (N12587, N12580, N6138, N12430);
not NOT1 (N12588, N12578);
or OR2 (N12589, N12585, N229);
nor NOR3 (N12590, N12586, N7389, N3476);
or OR3 (N12591, N12589, N2070, N9752);
xor XOR2 (N12592, N12582, N2914);
or OR3 (N12593, N12584, N11656, N7222);
and AND3 (N12594, N12592, N4705, N4259);
and AND3 (N12595, N12593, N8746, N6859);
or OR3 (N12596, N12571, N8680, N336);
nor NOR3 (N12597, N12588, N9068, N7365);
xor XOR2 (N12598, N12591, N12518);
not NOT1 (N12599, N12597);
xor XOR2 (N12600, N12598, N12153);
buf BUF1 (N12601, N12600);
not NOT1 (N12602, N12583);
nor NOR3 (N12603, N12596, N9389, N3425);
nor NOR2 (N12604, N12602, N12307);
nor NOR2 (N12605, N12601, N9528);
buf BUF1 (N12606, N12605);
nand NAND2 (N12607, N12604, N8984);
nand NAND4 (N12608, N12581, N7405, N3515, N12072);
nor NOR2 (N12609, N12603, N9660);
and AND2 (N12610, N12587, N2647);
nand NAND4 (N12611, N12608, N3800, N9121, N10365);
buf BUF1 (N12612, N12610);
nor NOR4 (N12613, N12612, N7582, N588, N8739);
nand NAND3 (N12614, N12595, N6047, N2229);
and AND3 (N12615, N12599, N5643, N433);
buf BUF1 (N12616, N12613);
not NOT1 (N12617, N12590);
nand NAND3 (N12618, N12572, N1538, N12275);
or OR4 (N12619, N12615, N2596, N1669, N7273);
and AND3 (N12620, N12594, N6990, N1901);
and AND3 (N12621, N12617, N4393, N9365);
nor NOR2 (N12622, N12616, N10332);
or OR2 (N12623, N12620, N11055);
xor XOR2 (N12624, N12622, N9539);
or OR4 (N12625, N12614, N6679, N39, N3041);
nand NAND3 (N12626, N12609, N1895, N2290);
and AND4 (N12627, N12625, N943, N11842, N3991);
or OR2 (N12628, N12626, N4443);
buf BUF1 (N12629, N12606);
xor XOR2 (N12630, N12611, N1081);
or OR4 (N12631, N12623, N5024, N8340, N9400);
and AND3 (N12632, N12628, N6248, N6895);
xor XOR2 (N12633, N12630, N7747);
buf BUF1 (N12634, N12619);
not NOT1 (N12635, N12633);
buf BUF1 (N12636, N12634);
not NOT1 (N12637, N12635);
or OR4 (N12638, N12636, N6874, N3613, N1791);
xor XOR2 (N12639, N12624, N921);
xor XOR2 (N12640, N12618, N9279);
not NOT1 (N12641, N12639);
nor NOR3 (N12642, N12631, N9615, N2756);
nand NAND4 (N12643, N12640, N8906, N4364, N6168);
xor XOR2 (N12644, N12607, N7973);
not NOT1 (N12645, N12642);
xor XOR2 (N12646, N12641, N9202);
and AND3 (N12647, N12646, N2596, N10419);
or OR3 (N12648, N12637, N921, N11697);
xor XOR2 (N12649, N12627, N8408);
nand NAND3 (N12650, N12643, N10454, N10994);
nand NAND4 (N12651, N12638, N2768, N782, N11760);
or OR4 (N12652, N12621, N9212, N770, N10705);
nand NAND3 (N12653, N12645, N9382, N11036);
buf BUF1 (N12654, N12647);
nor NOR4 (N12655, N12649, N8230, N8760, N604);
xor XOR2 (N12656, N12652, N4042);
or OR2 (N12657, N12654, N1332);
nand NAND3 (N12658, N12650, N2660, N5711);
and AND2 (N12659, N12653, N1454);
and AND4 (N12660, N12629, N10477, N2645, N7434);
not NOT1 (N12661, N12632);
or OR3 (N12662, N12648, N1451, N3473);
and AND4 (N12663, N12660, N11428, N4975, N1334);
not NOT1 (N12664, N12663);
buf BUF1 (N12665, N12662);
nand NAND3 (N12666, N12644, N1964, N5956);
not NOT1 (N12667, N12666);
buf BUF1 (N12668, N12664);
and AND3 (N12669, N12658, N3918, N9443);
not NOT1 (N12670, N12655);
or OR4 (N12671, N12665, N11145, N8072, N1327);
xor XOR2 (N12672, N12659, N10617);
and AND2 (N12673, N12661, N11380);
or OR3 (N12674, N12668, N8877, N10767);
or OR2 (N12675, N12669, N11618);
nand NAND2 (N12676, N12672, N6211);
xor XOR2 (N12677, N12651, N6499);
nand NAND4 (N12678, N12670, N5572, N10325, N9200);
nor NOR2 (N12679, N12675, N1155);
nand NAND3 (N12680, N12677, N6302, N580);
xor XOR2 (N12681, N12674, N7852);
nor NOR2 (N12682, N12681, N1742);
not NOT1 (N12683, N12667);
or OR4 (N12684, N12679, N10913, N2132, N9239);
xor XOR2 (N12685, N12656, N2902);
and AND4 (N12686, N12673, N4332, N1451, N2663);
and AND2 (N12687, N12685, N11959);
nand NAND4 (N12688, N12684, N12632, N3160, N11989);
nor NOR2 (N12689, N12682, N12134);
and AND2 (N12690, N12671, N10374);
buf BUF1 (N12691, N12688);
nor NOR4 (N12692, N12678, N6468, N12512, N1274);
xor XOR2 (N12693, N12657, N10519);
nor NOR2 (N12694, N12676, N11252);
nor NOR3 (N12695, N12691, N1498, N6199);
and AND3 (N12696, N12690, N9129, N11956);
nand NAND2 (N12697, N12694, N11642);
and AND4 (N12698, N12680, N7469, N5556, N540);
nand NAND4 (N12699, N12687, N8778, N1212, N2736);
buf BUF1 (N12700, N12689);
not NOT1 (N12701, N12697);
nor NOR4 (N12702, N12698, N2308, N6184, N2846);
not NOT1 (N12703, N12693);
or OR2 (N12704, N12703, N20);
nand NAND4 (N12705, N12701, N3815, N10175, N6888);
nand NAND4 (N12706, N12683, N3703, N3550, N8687);
and AND2 (N12707, N12699, N12315);
xor XOR2 (N12708, N12696, N1528);
buf BUF1 (N12709, N12702);
buf BUF1 (N12710, N12708);
buf BUF1 (N12711, N12706);
buf BUF1 (N12712, N12710);
not NOT1 (N12713, N12704);
buf BUF1 (N12714, N12692);
nor NOR2 (N12715, N12709, N4090);
nor NOR4 (N12716, N12686, N10366, N2725, N5912);
xor XOR2 (N12717, N12695, N2040);
xor XOR2 (N12718, N12716, N3780);
not NOT1 (N12719, N12717);
and AND4 (N12720, N12707, N9749, N9491, N1300);
buf BUF1 (N12721, N12714);
not NOT1 (N12722, N12718);
nor NOR4 (N12723, N12715, N6287, N6902, N7508);
and AND2 (N12724, N12723, N1270);
nand NAND4 (N12725, N12724, N7587, N10002, N4496);
nor NOR3 (N12726, N12700, N4125, N4835);
nor NOR4 (N12727, N12705, N8760, N1145, N1883);
nor NOR4 (N12728, N12721, N2159, N745, N8951);
nand NAND2 (N12729, N12713, N3840);
or OR2 (N12730, N12722, N4110);
not NOT1 (N12731, N12720);
or OR2 (N12732, N12719, N11076);
and AND3 (N12733, N12731, N2720, N9919);
not NOT1 (N12734, N12725);
xor XOR2 (N12735, N12727, N1780);
buf BUF1 (N12736, N12735);
nor NOR2 (N12737, N12729, N956);
xor XOR2 (N12738, N12728, N235);
nor NOR4 (N12739, N12726, N3819, N5015, N2716);
and AND4 (N12740, N12732, N1059, N5309, N4359);
nand NAND4 (N12741, N12737, N136, N7655, N10466);
not NOT1 (N12742, N12739);
buf BUF1 (N12743, N12734);
xor XOR2 (N12744, N12741, N4427);
not NOT1 (N12745, N12742);
buf BUF1 (N12746, N12745);
nor NOR4 (N12747, N12711, N850, N12154, N9500);
nand NAND2 (N12748, N12744, N2091);
nand NAND4 (N12749, N12747, N1513, N10510, N489);
nor NOR2 (N12750, N12738, N8619);
or OR4 (N12751, N12748, N8298, N12061, N12106);
nand NAND3 (N12752, N12750, N5296, N7748);
and AND4 (N12753, N12743, N6719, N7619, N11434);
nand NAND4 (N12754, N12712, N2000, N7619, N5437);
xor XOR2 (N12755, N12754, N4817);
and AND3 (N12756, N12752, N2941, N4818);
and AND3 (N12757, N12733, N4775, N10932);
not NOT1 (N12758, N12756);
xor XOR2 (N12759, N12749, N11828);
or OR3 (N12760, N12753, N3666, N4168);
and AND2 (N12761, N12730, N2175);
xor XOR2 (N12762, N12755, N12113);
xor XOR2 (N12763, N12746, N12380);
nand NAND4 (N12764, N12757, N4380, N340, N5564);
not NOT1 (N12765, N12740);
nor NOR2 (N12766, N12759, N3191);
buf BUF1 (N12767, N12736);
not NOT1 (N12768, N12763);
not NOT1 (N12769, N12766);
xor XOR2 (N12770, N12767, N4530);
nor NOR3 (N12771, N12758, N4849, N12563);
and AND3 (N12772, N12761, N7590, N6096);
or OR2 (N12773, N12764, N7883);
and AND4 (N12774, N12773, N6893, N5370, N10231);
xor XOR2 (N12775, N12770, N8497);
or OR3 (N12776, N12760, N8588, N5729);
xor XOR2 (N12777, N12771, N11743);
buf BUF1 (N12778, N12775);
nor NOR4 (N12779, N12777, N2431, N2111, N11869);
not NOT1 (N12780, N12778);
xor XOR2 (N12781, N12774, N2430);
or OR3 (N12782, N12769, N7483, N8381);
buf BUF1 (N12783, N12768);
xor XOR2 (N12784, N12781, N950);
buf BUF1 (N12785, N12762);
not NOT1 (N12786, N12776);
buf BUF1 (N12787, N12786);
nand NAND4 (N12788, N12779, N3145, N8569, N1627);
not NOT1 (N12789, N12782);
nand NAND2 (N12790, N12780, N9639);
not NOT1 (N12791, N12784);
or OR3 (N12792, N12791, N5608, N1741);
nand NAND4 (N12793, N12785, N4934, N8860, N1999);
buf BUF1 (N12794, N12793);
nor NOR4 (N12795, N12790, N12603, N12679, N2806);
buf BUF1 (N12796, N12772);
xor XOR2 (N12797, N12789, N4477);
and AND3 (N12798, N12792, N5131, N3697);
nor NOR2 (N12799, N12798, N2310);
and AND3 (N12800, N12783, N2883, N9340);
xor XOR2 (N12801, N12794, N6081);
nor NOR2 (N12802, N12799, N5149);
and AND4 (N12803, N12795, N1692, N6181, N3828);
nand NAND4 (N12804, N12788, N2626, N5516, N2046);
nand NAND3 (N12805, N12800, N5127, N5868);
not NOT1 (N12806, N12801);
and AND2 (N12807, N12797, N4825);
buf BUF1 (N12808, N12803);
nand NAND2 (N12809, N12787, N8741);
not NOT1 (N12810, N12751);
nand NAND3 (N12811, N12802, N6098, N6528);
nor NOR3 (N12812, N12808, N11872, N9680);
nor NOR2 (N12813, N12804, N8682);
nor NOR3 (N12814, N12809, N5085, N6091);
nand NAND2 (N12815, N12765, N11454);
endmodule