// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N1602,N1614,N1606,N1604,N1610,N1613,N1609,N1612,N1598,N1615;

buf BUF1 (N16, N3);
nand NAND4 (N17, N8, N2, N15, N9);
buf BUF1 (N18, N3);
not NOT1 (N19, N8);
xor XOR2 (N20, N19, N1);
or OR3 (N21, N6, N7, N19);
nor NOR2 (N22, N1, N16);
nor NOR2 (N23, N21, N19);
or OR4 (N24, N6, N21, N14, N21);
xor XOR2 (N25, N17, N16);
nor NOR4 (N26, N3, N5, N18, N15);
not NOT1 (N27, N18);
buf BUF1 (N28, N12);
or OR2 (N29, N6, N17);
nand NAND3 (N30, N7, N1, N13);
xor XOR2 (N31, N25, N8);
not NOT1 (N32, N20);
xor XOR2 (N33, N23, N6);
nand NAND2 (N34, N31, N30);
nor NOR4 (N35, N32, N16, N19, N31);
nand NAND3 (N36, N15, N16, N35);
nand NAND2 (N37, N21, N14);
xor XOR2 (N38, N29, N18);
nand NAND4 (N39, N37, N23, N8, N27);
not NOT1 (N40, N39);
and AND4 (N41, N39, N40, N16, N28);
nor NOR4 (N42, N25, N16, N23, N40);
or OR4 (N43, N11, N23, N20, N11);
buf BUF1 (N44, N22);
xor XOR2 (N45, N24, N34);
or OR3 (N46, N45, N7, N6);
buf BUF1 (N47, N24);
nand NAND3 (N48, N44, N16, N35);
nand NAND3 (N49, N42, N34, N8);
or OR3 (N50, N26, N30, N33);
or OR4 (N51, N8, N3, N23, N26);
and AND2 (N52, N43, N43);
or OR2 (N53, N51, N15);
xor XOR2 (N54, N46, N39);
not NOT1 (N55, N47);
xor XOR2 (N56, N52, N19);
nand NAND3 (N57, N53, N42, N30);
nand NAND3 (N58, N54, N26, N1);
not NOT1 (N59, N48);
xor XOR2 (N60, N57, N7);
and AND4 (N61, N49, N51, N14, N48);
xor XOR2 (N62, N60, N2);
or OR4 (N63, N38, N40, N46, N43);
buf BUF1 (N64, N55);
and AND2 (N65, N36, N4);
xor XOR2 (N66, N56, N16);
not NOT1 (N67, N61);
and AND2 (N68, N41, N54);
or OR3 (N69, N66, N30, N59);
or OR3 (N70, N25, N60, N56);
or OR4 (N71, N70, N57, N2, N3);
buf BUF1 (N72, N68);
buf BUF1 (N73, N64);
and AND2 (N74, N65, N6);
nor NOR4 (N75, N69, N47, N4, N58);
or OR4 (N76, N42, N17, N18, N20);
xor XOR2 (N77, N76, N70);
nor NOR4 (N78, N67, N9, N8, N6);
buf BUF1 (N79, N77);
nor NOR4 (N80, N79, N31, N36, N51);
not NOT1 (N81, N63);
not NOT1 (N82, N50);
xor XOR2 (N83, N62, N62);
and AND4 (N84, N74, N81, N19, N71);
and AND3 (N85, N45, N65, N39);
nand NAND2 (N86, N75, N32);
nand NAND4 (N87, N40, N44, N29, N49);
and AND4 (N88, N80, N26, N63, N58);
or OR3 (N89, N78, N50, N48);
or OR3 (N90, N87, N8, N74);
buf BUF1 (N91, N88);
xor XOR2 (N92, N90, N47);
nand NAND2 (N93, N82, N58);
nor NOR2 (N94, N86, N84);
nor NOR3 (N95, N9, N59, N5);
and AND3 (N96, N89, N68, N93);
not NOT1 (N97, N96);
xor XOR2 (N98, N62, N16);
nor NOR2 (N99, N91, N35);
or OR2 (N100, N92, N47);
xor XOR2 (N101, N94, N76);
nand NAND3 (N102, N100, N11, N47);
buf BUF1 (N103, N95);
xor XOR2 (N104, N102, N70);
xor XOR2 (N105, N85, N66);
xor XOR2 (N106, N97, N70);
nor NOR4 (N107, N103, N54, N32, N78);
nor NOR3 (N108, N106, N61, N19);
buf BUF1 (N109, N73);
and AND3 (N110, N98, N19, N49);
xor XOR2 (N111, N99, N95);
not NOT1 (N112, N101);
buf BUF1 (N113, N107);
nand NAND2 (N114, N110, N108);
or OR2 (N115, N108, N112);
and AND4 (N116, N89, N100, N73, N1);
nand NAND3 (N117, N109, N28, N40);
xor XOR2 (N118, N117, N102);
and AND3 (N119, N72, N2, N111);
buf BUF1 (N120, N76);
nor NOR3 (N121, N116, N28, N10);
nor NOR2 (N122, N118, N67);
xor XOR2 (N123, N105, N32);
nand NAND2 (N124, N122, N94);
nor NOR3 (N125, N119, N74, N49);
and AND3 (N126, N123, N62, N64);
xor XOR2 (N127, N83, N11);
buf BUF1 (N128, N125);
xor XOR2 (N129, N114, N48);
xor XOR2 (N130, N113, N82);
nand NAND4 (N131, N129, N30, N35, N53);
not NOT1 (N132, N115);
and AND3 (N133, N121, N87, N126);
nor NOR2 (N134, N32, N10);
not NOT1 (N135, N133);
xor XOR2 (N136, N128, N22);
or OR3 (N137, N135, N120, N135);
not NOT1 (N138, N20);
xor XOR2 (N139, N132, N105);
nor NOR3 (N140, N124, N112, N59);
xor XOR2 (N141, N134, N130);
nor NOR2 (N142, N59, N34);
or OR3 (N143, N104, N18, N82);
or OR4 (N144, N136, N54, N95, N14);
nand NAND4 (N145, N142, N45, N25, N16);
or OR4 (N146, N139, N59, N27, N123);
buf BUF1 (N147, N145);
xor XOR2 (N148, N143, N34);
not NOT1 (N149, N140);
nand NAND2 (N150, N149, N139);
xor XOR2 (N151, N150, N111);
buf BUF1 (N152, N148);
xor XOR2 (N153, N146, N105);
xor XOR2 (N154, N153, N24);
xor XOR2 (N155, N137, N45);
nor NOR3 (N156, N154, N123, N13);
and AND3 (N157, N144, N82, N102);
xor XOR2 (N158, N127, N79);
and AND4 (N159, N147, N84, N127, N20);
or OR3 (N160, N159, N9, N21);
not NOT1 (N161, N138);
or OR2 (N162, N131, N53);
or OR2 (N163, N158, N84);
xor XOR2 (N164, N157, N28);
buf BUF1 (N165, N155);
not NOT1 (N166, N141);
buf BUF1 (N167, N160);
and AND3 (N168, N163, N83, N136);
not NOT1 (N169, N151);
or OR4 (N170, N168, N113, N112, N140);
nor NOR3 (N171, N169, N155, N43);
and AND4 (N172, N171, N139, N78, N118);
not NOT1 (N173, N167);
buf BUF1 (N174, N173);
or OR3 (N175, N170, N43, N104);
not NOT1 (N176, N161);
or OR3 (N177, N156, N38, N133);
and AND3 (N178, N164, N48, N146);
not NOT1 (N179, N175);
nand NAND4 (N180, N177, N35, N102, N45);
or OR2 (N181, N165, N11);
buf BUF1 (N182, N176);
nor NOR2 (N183, N178, N17);
and AND2 (N184, N152, N176);
not NOT1 (N185, N184);
nor NOR3 (N186, N179, N13, N147);
or OR2 (N187, N180, N72);
or OR2 (N188, N187, N100);
xor XOR2 (N189, N162, N58);
and AND2 (N190, N185, N2);
not NOT1 (N191, N174);
nand NAND4 (N192, N172, N161, N186, N148);
not NOT1 (N193, N98);
xor XOR2 (N194, N191, N174);
not NOT1 (N195, N182);
nand NAND4 (N196, N183, N95, N129, N23);
nand NAND4 (N197, N190, N191, N114, N99);
and AND3 (N198, N188, N20, N71);
and AND4 (N199, N195, N86, N143, N193);
nand NAND4 (N200, N47, N104, N58, N180);
or OR3 (N201, N166, N170, N169);
nor NOR3 (N202, N197, N106, N26);
not NOT1 (N203, N194);
nand NAND4 (N204, N203, N39, N149, N105);
nand NAND3 (N205, N201, N146, N108);
not NOT1 (N206, N200);
or OR2 (N207, N198, N173);
and AND4 (N208, N206, N198, N152, N175);
nand NAND4 (N209, N192, N11, N144, N180);
buf BUF1 (N210, N207);
or OR4 (N211, N189, N112, N148, N201);
xor XOR2 (N212, N199, N122);
and AND4 (N213, N210, N100, N173, N73);
buf BUF1 (N214, N202);
buf BUF1 (N215, N211);
nor NOR3 (N216, N215, N168, N171);
nor NOR3 (N217, N196, N149, N166);
nand NAND3 (N218, N209, N130, N92);
not NOT1 (N219, N217);
and AND4 (N220, N204, N218, N10, N23);
not NOT1 (N221, N39);
nor NOR2 (N222, N221, N118);
xor XOR2 (N223, N216, N69);
nand NAND3 (N224, N181, N138, N146);
or OR4 (N225, N222, N43, N108, N160);
xor XOR2 (N226, N220, N20);
nor NOR4 (N227, N214, N192, N18, N94);
buf BUF1 (N228, N205);
not NOT1 (N229, N212);
and AND2 (N230, N224, N64);
not NOT1 (N231, N208);
nand NAND3 (N232, N225, N204, N98);
nor NOR2 (N233, N223, N155);
and AND2 (N234, N232, N91);
or OR3 (N235, N229, N21, N122);
xor XOR2 (N236, N219, N96);
not NOT1 (N237, N227);
and AND3 (N238, N234, N179, N165);
xor XOR2 (N239, N236, N135);
nand NAND2 (N240, N228, N123);
xor XOR2 (N241, N230, N1);
or OR3 (N242, N240, N165, N133);
nor NOR2 (N243, N238, N5);
or OR2 (N244, N226, N219);
xor XOR2 (N245, N237, N241);
buf BUF1 (N246, N194);
nor NOR4 (N247, N243, N112, N91, N119);
xor XOR2 (N248, N239, N221);
nor NOR4 (N249, N231, N77, N10, N237);
and AND2 (N250, N246, N167);
and AND2 (N251, N242, N175);
xor XOR2 (N252, N244, N118);
not NOT1 (N253, N252);
nand NAND3 (N254, N235, N250, N133);
nor NOR3 (N255, N54, N45, N8);
buf BUF1 (N256, N255);
or OR3 (N257, N256, N112, N71);
and AND3 (N258, N257, N132, N104);
not NOT1 (N259, N213);
or OR2 (N260, N251, N82);
nor NOR3 (N261, N248, N73, N169);
and AND3 (N262, N247, N163, N105);
xor XOR2 (N263, N260, N77);
xor XOR2 (N264, N254, N83);
or OR2 (N265, N249, N150);
buf BUF1 (N266, N263);
xor XOR2 (N267, N253, N146);
buf BUF1 (N268, N265);
xor XOR2 (N269, N259, N218);
nor NOR2 (N270, N268, N152);
xor XOR2 (N271, N233, N145);
xor XOR2 (N272, N264, N257);
not NOT1 (N273, N262);
nand NAND3 (N274, N261, N201, N179);
and AND3 (N275, N267, N199, N191);
nand NAND3 (N276, N272, N259, N44);
not NOT1 (N277, N266);
buf BUF1 (N278, N258);
or OR4 (N279, N275, N202, N85, N160);
or OR4 (N280, N274, N239, N16, N18);
or OR2 (N281, N270, N119);
buf BUF1 (N282, N273);
nand NAND3 (N283, N276, N147, N20);
and AND4 (N284, N269, N122, N225, N115);
xor XOR2 (N285, N281, N19);
and AND4 (N286, N285, N110, N183, N186);
xor XOR2 (N287, N245, N141);
and AND2 (N288, N283, N213);
or OR2 (N289, N277, N19);
buf BUF1 (N290, N288);
not NOT1 (N291, N290);
nand NAND3 (N292, N282, N99, N110);
or OR2 (N293, N280, N49);
not NOT1 (N294, N279);
and AND4 (N295, N287, N227, N54, N178);
and AND4 (N296, N271, N8, N134, N200);
or OR2 (N297, N292, N296);
nor NOR3 (N298, N59, N39, N28);
not NOT1 (N299, N295);
or OR4 (N300, N291, N271, N273, N85);
or OR4 (N301, N300, N181, N33, N142);
nand NAND3 (N302, N301, N173, N96);
nor NOR2 (N303, N299, N59);
and AND3 (N304, N302, N56, N155);
or OR4 (N305, N298, N36, N100, N232);
or OR3 (N306, N305, N35, N269);
nand NAND2 (N307, N284, N108);
or OR4 (N308, N289, N70, N142, N196);
or OR3 (N309, N297, N271, N84);
nand NAND3 (N310, N293, N116, N303);
not NOT1 (N311, N283);
buf BUF1 (N312, N286);
and AND3 (N313, N278, N2, N43);
and AND2 (N314, N304, N224);
and AND4 (N315, N314, N108, N209, N249);
nand NAND2 (N316, N294, N81);
buf BUF1 (N317, N316);
nor NOR2 (N318, N308, N196);
buf BUF1 (N319, N317);
not NOT1 (N320, N313);
and AND2 (N321, N312, N146);
xor XOR2 (N322, N310, N150);
nor NOR3 (N323, N321, N127, N17);
nor NOR4 (N324, N319, N84, N223, N150);
and AND4 (N325, N306, N163, N127, N235);
xor XOR2 (N326, N320, N124);
nand NAND3 (N327, N322, N21, N152);
nand NAND4 (N328, N311, N2, N149, N167);
nor NOR2 (N329, N327, N155);
not NOT1 (N330, N326);
and AND2 (N331, N330, N56);
buf BUF1 (N332, N309);
not NOT1 (N333, N331);
or OR3 (N334, N324, N32, N255);
and AND2 (N335, N334, N193);
buf BUF1 (N336, N329);
nand NAND3 (N337, N325, N211, N144);
and AND2 (N338, N336, N19);
not NOT1 (N339, N333);
not NOT1 (N340, N315);
or OR2 (N341, N335, N136);
nand NAND3 (N342, N323, N25, N135);
xor XOR2 (N343, N342, N148);
not NOT1 (N344, N338);
nand NAND4 (N345, N343, N170, N292, N336);
nand NAND2 (N346, N345, N269);
buf BUF1 (N347, N339);
xor XOR2 (N348, N337, N314);
nand NAND4 (N349, N346, N84, N126, N222);
or OR4 (N350, N349, N206, N64, N136);
not NOT1 (N351, N307);
xor XOR2 (N352, N350, N71);
not NOT1 (N353, N344);
buf BUF1 (N354, N353);
or OR2 (N355, N351, N272);
and AND3 (N356, N354, N297, N354);
xor XOR2 (N357, N340, N136);
not NOT1 (N358, N348);
not NOT1 (N359, N358);
nor NOR4 (N360, N332, N302, N111, N276);
not NOT1 (N361, N360);
or OR3 (N362, N347, N22, N338);
nor NOR3 (N363, N356, N1, N151);
nand NAND4 (N364, N341, N173, N91, N107);
not NOT1 (N365, N357);
or OR4 (N366, N364, N247, N56, N253);
or OR4 (N367, N361, N34, N57, N167);
not NOT1 (N368, N355);
or OR3 (N369, N367, N172, N306);
or OR3 (N370, N365, N87, N267);
buf BUF1 (N371, N370);
nor NOR4 (N372, N362, N296, N61, N297);
not NOT1 (N373, N352);
buf BUF1 (N374, N363);
not NOT1 (N375, N373);
nand NAND4 (N376, N366, N285, N286, N76);
nand NAND2 (N377, N375, N85);
xor XOR2 (N378, N376, N167);
and AND2 (N379, N318, N110);
not NOT1 (N380, N378);
nand NAND3 (N381, N379, N126, N34);
not NOT1 (N382, N368);
and AND4 (N383, N381, N21, N4, N345);
and AND3 (N384, N371, N370, N317);
not NOT1 (N385, N374);
nor NOR4 (N386, N385, N72, N295, N288);
buf BUF1 (N387, N372);
not NOT1 (N388, N386);
or OR3 (N389, N369, N208, N194);
not NOT1 (N390, N382);
buf BUF1 (N391, N328);
not NOT1 (N392, N389);
nand NAND3 (N393, N359, N245, N65);
not NOT1 (N394, N390);
and AND4 (N395, N391, N155, N182, N237);
nand NAND2 (N396, N388, N254);
nor NOR2 (N397, N384, N103);
not NOT1 (N398, N380);
not NOT1 (N399, N377);
nand NAND4 (N400, N395, N44, N224, N374);
xor XOR2 (N401, N387, N239);
buf BUF1 (N402, N396);
nand NAND3 (N403, N397, N369, N374);
and AND4 (N404, N394, N218, N155, N357);
nand NAND4 (N405, N399, N131, N192, N264);
xor XOR2 (N406, N402, N323);
nor NOR4 (N407, N406, N162, N229, N26);
nand NAND4 (N408, N404, N303, N144, N68);
or OR4 (N409, N403, N14, N372, N395);
and AND2 (N410, N383, N14);
not NOT1 (N411, N407);
xor XOR2 (N412, N393, N20);
xor XOR2 (N413, N412, N72);
nand NAND3 (N414, N413, N338, N354);
not NOT1 (N415, N398);
xor XOR2 (N416, N392, N245);
or OR2 (N417, N410, N217);
not NOT1 (N418, N401);
xor XOR2 (N419, N405, N272);
buf BUF1 (N420, N411);
not NOT1 (N421, N417);
not NOT1 (N422, N419);
and AND4 (N423, N421, N376, N393, N19);
nor NOR3 (N424, N420, N221, N225);
or OR4 (N425, N423, N415, N367, N392);
or OR2 (N426, N420, N304);
not NOT1 (N427, N426);
not NOT1 (N428, N408);
or OR2 (N429, N400, N168);
nand NAND4 (N430, N416, N202, N12, N233);
not NOT1 (N431, N414);
nand NAND4 (N432, N427, N333, N294, N397);
buf BUF1 (N433, N422);
not NOT1 (N434, N424);
xor XOR2 (N435, N409, N189);
not NOT1 (N436, N428);
buf BUF1 (N437, N418);
and AND4 (N438, N429, N351, N18, N192);
or OR4 (N439, N435, N247, N193, N125);
and AND4 (N440, N434, N266, N222, N384);
or OR4 (N441, N436, N105, N268, N60);
and AND3 (N442, N439, N139, N207);
or OR3 (N443, N441, N120, N71);
nor NOR4 (N444, N440, N369, N212, N79);
nor NOR4 (N445, N442, N386, N13, N129);
buf BUF1 (N446, N431);
buf BUF1 (N447, N430);
not NOT1 (N448, N445);
nor NOR4 (N449, N438, N314, N35, N214);
buf BUF1 (N450, N448);
buf BUF1 (N451, N449);
not NOT1 (N452, N451);
nor NOR3 (N453, N443, N104, N70);
and AND3 (N454, N447, N404, N336);
nor NOR3 (N455, N425, N298, N56);
or OR4 (N456, N452, N258, N40, N228);
xor XOR2 (N457, N456, N377);
not NOT1 (N458, N457);
xor XOR2 (N459, N453, N263);
nand NAND3 (N460, N455, N68, N124);
buf BUF1 (N461, N433);
nand NAND4 (N462, N432, N189, N117, N251);
xor XOR2 (N463, N446, N44);
nand NAND2 (N464, N460, N349);
nor NOR4 (N465, N437, N123, N269, N254);
not NOT1 (N466, N459);
xor XOR2 (N467, N463, N331);
not NOT1 (N468, N444);
xor XOR2 (N469, N461, N340);
buf BUF1 (N470, N466);
buf BUF1 (N471, N468);
or OR3 (N472, N467, N154, N432);
buf BUF1 (N473, N458);
buf BUF1 (N474, N454);
nand NAND2 (N475, N462, N380);
xor XOR2 (N476, N465, N180);
nor NOR4 (N477, N471, N45, N391, N467);
and AND4 (N478, N450, N88, N43, N126);
and AND2 (N479, N477, N367);
nand NAND4 (N480, N478, N271, N159, N160);
or OR4 (N481, N474, N53, N18, N72);
buf BUF1 (N482, N476);
xor XOR2 (N483, N480, N370);
nor NOR2 (N484, N479, N303);
buf BUF1 (N485, N482);
buf BUF1 (N486, N481);
nor NOR3 (N487, N484, N154, N13);
or OR3 (N488, N464, N379, N211);
nor NOR2 (N489, N470, N355);
and AND3 (N490, N469, N162, N87);
and AND4 (N491, N488, N19, N151, N10);
and AND2 (N492, N473, N221);
not NOT1 (N493, N486);
not NOT1 (N494, N489);
nand NAND4 (N495, N472, N175, N149, N407);
nand NAND4 (N496, N485, N477, N235, N379);
and AND4 (N497, N487, N415, N7, N8);
and AND2 (N498, N483, N120);
or OR4 (N499, N495, N230, N83, N497);
or OR3 (N500, N48, N312, N15);
not NOT1 (N501, N496);
and AND2 (N502, N494, N377);
and AND2 (N503, N475, N5);
nand NAND3 (N504, N491, N102, N134);
or OR3 (N505, N499, N266, N153);
not NOT1 (N506, N503);
not NOT1 (N507, N498);
buf BUF1 (N508, N504);
not NOT1 (N509, N500);
nor NOR2 (N510, N501, N272);
and AND3 (N511, N505, N295, N498);
not NOT1 (N512, N506);
xor XOR2 (N513, N511, N3);
nor NOR3 (N514, N508, N480, N311);
and AND2 (N515, N502, N356);
not NOT1 (N516, N509);
nand NAND3 (N517, N515, N76, N200);
buf BUF1 (N518, N490);
xor XOR2 (N519, N493, N329);
nor NOR4 (N520, N512, N48, N156, N243);
and AND2 (N521, N510, N193);
or OR2 (N522, N520, N467);
nor NOR3 (N523, N522, N102, N250);
or OR2 (N524, N523, N249);
nor NOR2 (N525, N519, N373);
buf BUF1 (N526, N525);
nand NAND4 (N527, N521, N310, N276, N486);
and AND4 (N528, N513, N309, N256, N415);
or OR2 (N529, N517, N331);
and AND3 (N530, N516, N37, N491);
nand NAND4 (N531, N514, N296, N35, N98);
and AND4 (N532, N492, N411, N396, N102);
and AND4 (N533, N524, N400, N273, N91);
buf BUF1 (N534, N530);
and AND4 (N535, N528, N403, N16, N246);
nand NAND4 (N536, N531, N454, N355, N385);
buf BUF1 (N537, N507);
buf BUF1 (N538, N536);
buf BUF1 (N539, N518);
xor XOR2 (N540, N537, N439);
not NOT1 (N541, N538);
nand NAND2 (N542, N526, N13);
buf BUF1 (N543, N539);
nor NOR3 (N544, N529, N471, N306);
nand NAND2 (N545, N542, N369);
nor NOR4 (N546, N545, N321, N359, N272);
or OR4 (N547, N546, N44, N27, N156);
nand NAND3 (N548, N527, N65, N216);
or OR3 (N549, N543, N240, N235);
or OR2 (N550, N532, N338);
or OR2 (N551, N533, N200);
not NOT1 (N552, N550);
nor NOR3 (N553, N544, N115, N338);
and AND2 (N554, N540, N72);
not NOT1 (N555, N549);
nand NAND3 (N556, N541, N114, N73);
not NOT1 (N557, N548);
and AND3 (N558, N556, N349, N244);
nand NAND2 (N559, N534, N491);
and AND3 (N560, N554, N526, N80);
or OR3 (N561, N552, N322, N535);
not NOT1 (N562, N441);
and AND4 (N563, N551, N400, N541, N423);
nand NAND2 (N564, N557, N121);
nor NOR4 (N565, N564, N299, N388, N336);
nor NOR2 (N566, N560, N121);
xor XOR2 (N567, N547, N350);
or OR2 (N568, N563, N293);
xor XOR2 (N569, N562, N97);
and AND2 (N570, N553, N500);
not NOT1 (N571, N565);
nand NAND2 (N572, N555, N464);
nand NAND3 (N573, N566, N477, N312);
xor XOR2 (N574, N573, N109);
nor NOR4 (N575, N574, N193, N151, N28);
buf BUF1 (N576, N570);
or OR3 (N577, N576, N35, N98);
not NOT1 (N578, N559);
nor NOR3 (N579, N558, N64, N473);
nand NAND4 (N580, N575, N298, N62, N37);
xor XOR2 (N581, N567, N218);
not NOT1 (N582, N580);
xor XOR2 (N583, N577, N55);
and AND3 (N584, N572, N92, N393);
not NOT1 (N585, N579);
not NOT1 (N586, N578);
buf BUF1 (N587, N561);
and AND2 (N588, N582, N158);
buf BUF1 (N589, N568);
buf BUF1 (N590, N571);
nor NOR4 (N591, N583, N572, N546, N400);
or OR2 (N592, N569, N415);
and AND2 (N593, N584, N428);
buf BUF1 (N594, N587);
and AND4 (N595, N594, N177, N441, N264);
and AND3 (N596, N585, N122, N225);
nor NOR4 (N597, N593, N465, N384, N286);
xor XOR2 (N598, N591, N504);
and AND4 (N599, N590, N140, N383, N568);
or OR2 (N600, N599, N357);
xor XOR2 (N601, N592, N83);
buf BUF1 (N602, N586);
buf BUF1 (N603, N589);
not NOT1 (N604, N595);
not NOT1 (N605, N600);
buf BUF1 (N606, N601);
or OR2 (N607, N598, N336);
buf BUF1 (N608, N607);
buf BUF1 (N609, N604);
nand NAND4 (N610, N609, N128, N441, N75);
or OR4 (N611, N603, N530, N238, N218);
nand NAND3 (N612, N597, N504, N395);
xor XOR2 (N613, N605, N502);
and AND3 (N614, N608, N487, N547);
or OR3 (N615, N581, N197, N359);
xor XOR2 (N616, N602, N260);
not NOT1 (N617, N596);
and AND2 (N618, N614, N395);
not NOT1 (N619, N613);
nand NAND3 (N620, N606, N618, N245);
or OR2 (N621, N61, N593);
not NOT1 (N622, N612);
nand NAND2 (N623, N615, N395);
nor NOR2 (N624, N621, N63);
buf BUF1 (N625, N623);
not NOT1 (N626, N616);
nand NAND2 (N627, N622, N468);
xor XOR2 (N628, N619, N569);
nand NAND3 (N629, N588, N41, N153);
nand NAND2 (N630, N617, N470);
and AND3 (N631, N627, N372, N255);
not NOT1 (N632, N610);
or OR4 (N633, N624, N214, N9, N399);
or OR4 (N634, N628, N480, N559, N326);
xor XOR2 (N635, N631, N163);
nand NAND2 (N636, N635, N386);
not NOT1 (N637, N625);
buf BUF1 (N638, N633);
not NOT1 (N639, N629);
nor NOR3 (N640, N626, N246, N555);
not NOT1 (N641, N632);
buf BUF1 (N642, N640);
xor XOR2 (N643, N637, N255);
buf BUF1 (N644, N620);
xor XOR2 (N645, N634, N574);
not NOT1 (N646, N641);
or OR2 (N647, N646, N52);
nor NOR2 (N648, N638, N255);
buf BUF1 (N649, N639);
xor XOR2 (N650, N647, N59);
xor XOR2 (N651, N648, N328);
not NOT1 (N652, N642);
nor NOR2 (N653, N644, N149);
and AND3 (N654, N645, N229, N630);
or OR2 (N655, N461, N555);
not NOT1 (N656, N643);
xor XOR2 (N657, N651, N370);
nand NAND4 (N658, N650, N110, N359, N531);
xor XOR2 (N659, N611, N77);
or OR4 (N660, N659, N333, N61, N509);
nor NOR2 (N661, N660, N582);
xor XOR2 (N662, N654, N429);
nand NAND2 (N663, N656, N588);
xor XOR2 (N664, N636, N33);
not NOT1 (N665, N664);
not NOT1 (N666, N652);
buf BUF1 (N667, N661);
or OR2 (N668, N662, N400);
not NOT1 (N669, N667);
nor NOR4 (N670, N663, N11, N165, N510);
or OR3 (N671, N665, N509, N83);
xor XOR2 (N672, N666, N648);
buf BUF1 (N673, N669);
buf BUF1 (N674, N649);
not NOT1 (N675, N658);
not NOT1 (N676, N670);
nand NAND4 (N677, N675, N228, N19, N30);
buf BUF1 (N678, N657);
buf BUF1 (N679, N671);
xor XOR2 (N680, N676, N613);
not NOT1 (N681, N680);
or OR3 (N682, N678, N612, N27);
nand NAND4 (N683, N677, N190, N194, N272);
or OR2 (N684, N681, N433);
buf BUF1 (N685, N682);
buf BUF1 (N686, N672);
buf BUF1 (N687, N686);
nand NAND2 (N688, N674, N591);
or OR3 (N689, N653, N218, N88);
and AND2 (N690, N685, N163);
nand NAND3 (N691, N689, N545, N547);
xor XOR2 (N692, N673, N338);
buf BUF1 (N693, N687);
xor XOR2 (N694, N688, N259);
and AND2 (N695, N655, N489);
nand NAND3 (N696, N679, N323, N35);
not NOT1 (N697, N695);
or OR2 (N698, N697, N130);
xor XOR2 (N699, N698, N483);
and AND3 (N700, N699, N138, N347);
xor XOR2 (N701, N700, N679);
nor NOR2 (N702, N690, N128);
or OR3 (N703, N693, N119, N690);
not NOT1 (N704, N694);
buf BUF1 (N705, N696);
xor XOR2 (N706, N692, N75);
and AND2 (N707, N668, N504);
xor XOR2 (N708, N684, N259);
buf BUF1 (N709, N702);
buf BUF1 (N710, N703);
nand NAND2 (N711, N705, N482);
nand NAND4 (N712, N707, N270, N156, N98);
nor NOR2 (N713, N709, N405);
not NOT1 (N714, N713);
nand NAND2 (N715, N691, N58);
and AND3 (N716, N715, N492, N584);
not NOT1 (N717, N706);
not NOT1 (N718, N716);
and AND2 (N719, N708, N629);
and AND2 (N720, N719, N459);
or OR4 (N721, N720, N44, N598, N582);
not NOT1 (N722, N704);
nand NAND4 (N723, N683, N332, N463, N123);
nand NAND4 (N724, N710, N236, N355, N228);
nand NAND2 (N725, N717, N397);
nand NAND4 (N726, N722, N573, N462, N510);
and AND3 (N727, N726, N353, N470);
or OR4 (N728, N724, N78, N199, N121);
nand NAND4 (N729, N714, N707, N537, N688);
or OR3 (N730, N728, N381, N294);
not NOT1 (N731, N727);
and AND3 (N732, N729, N568, N383);
xor XOR2 (N733, N701, N72);
or OR2 (N734, N725, N268);
nand NAND4 (N735, N723, N356, N198, N619);
buf BUF1 (N736, N721);
buf BUF1 (N737, N730);
or OR2 (N738, N731, N130);
or OR2 (N739, N733, N40);
xor XOR2 (N740, N735, N297);
xor XOR2 (N741, N732, N165);
not NOT1 (N742, N737);
and AND3 (N743, N741, N366, N130);
nor NOR3 (N744, N742, N668, N434);
or OR2 (N745, N744, N135);
not NOT1 (N746, N734);
nand NAND2 (N747, N718, N637);
or OR3 (N748, N711, N249, N493);
not NOT1 (N749, N745);
nor NOR2 (N750, N740, N616);
xor XOR2 (N751, N748, N204);
nor NOR4 (N752, N712, N159, N219, N449);
xor XOR2 (N753, N743, N52);
not NOT1 (N754, N753);
nand NAND2 (N755, N736, N723);
nor NOR4 (N756, N749, N360, N620, N336);
xor XOR2 (N757, N755, N728);
and AND4 (N758, N746, N614, N19, N313);
nand NAND2 (N759, N738, N701);
xor XOR2 (N760, N759, N38);
not NOT1 (N761, N747);
and AND3 (N762, N761, N556, N132);
and AND3 (N763, N756, N220, N460);
and AND4 (N764, N751, N350, N450, N752);
and AND4 (N765, N683, N66, N468, N229);
buf BUF1 (N766, N765);
or OR4 (N767, N757, N512, N482, N675);
nor NOR3 (N768, N763, N79, N529);
xor XOR2 (N769, N768, N627);
and AND3 (N770, N769, N7, N488);
or OR4 (N771, N766, N161, N225, N424);
nor NOR3 (N772, N762, N270, N684);
buf BUF1 (N773, N750);
not NOT1 (N774, N754);
nor NOR3 (N775, N773, N65, N12);
xor XOR2 (N776, N760, N603);
not NOT1 (N777, N758);
xor XOR2 (N778, N774, N418);
buf BUF1 (N779, N764);
nand NAND2 (N780, N778, N594);
not NOT1 (N781, N779);
xor XOR2 (N782, N781, N292);
or OR3 (N783, N782, N148, N530);
and AND4 (N784, N767, N372, N664, N606);
xor XOR2 (N785, N780, N135);
nand NAND4 (N786, N739, N615, N275, N518);
nand NAND3 (N787, N771, N725, N165);
not NOT1 (N788, N776);
xor XOR2 (N789, N784, N548);
nor NOR2 (N790, N777, N106);
xor XOR2 (N791, N788, N524);
nor NOR2 (N792, N791, N65);
not NOT1 (N793, N775);
and AND3 (N794, N792, N367, N751);
or OR3 (N795, N794, N159, N26);
nand NAND4 (N796, N772, N500, N715, N216);
nor NOR2 (N797, N785, N482);
and AND4 (N798, N790, N419, N586, N390);
nand NAND2 (N799, N798, N160);
or OR2 (N800, N799, N761);
nand NAND2 (N801, N789, N315);
nor NOR3 (N802, N796, N619, N554);
or OR3 (N803, N783, N216, N151);
nor NOR3 (N804, N795, N792, N432);
xor XOR2 (N805, N802, N661);
not NOT1 (N806, N800);
or OR4 (N807, N806, N305, N519, N190);
buf BUF1 (N808, N804);
not NOT1 (N809, N808);
nor NOR4 (N810, N801, N171, N714, N606);
and AND4 (N811, N810, N215, N475, N185);
nand NAND3 (N812, N811, N41, N705);
not NOT1 (N813, N807);
not NOT1 (N814, N812);
nor NOR3 (N815, N809, N199, N151);
not NOT1 (N816, N786);
buf BUF1 (N817, N805);
nand NAND4 (N818, N787, N396, N477, N259);
nand NAND4 (N819, N814, N15, N205, N255);
or OR2 (N820, N817, N476);
and AND4 (N821, N770, N373, N740, N404);
buf BUF1 (N822, N815);
nor NOR3 (N823, N819, N611, N749);
nand NAND3 (N824, N822, N238, N31);
nor NOR2 (N825, N803, N435);
buf BUF1 (N826, N824);
xor XOR2 (N827, N820, N634);
not NOT1 (N828, N821);
and AND3 (N829, N826, N11, N380);
buf BUF1 (N830, N829);
or OR4 (N831, N827, N573, N439, N16);
and AND4 (N832, N797, N383, N615, N48);
and AND4 (N833, N823, N393, N213, N645);
nor NOR4 (N834, N818, N354, N317, N738);
nor NOR4 (N835, N830, N570, N6, N478);
buf BUF1 (N836, N828);
and AND3 (N837, N793, N513, N660);
nand NAND4 (N838, N831, N346, N836, N789);
and AND2 (N839, N357, N86);
xor XOR2 (N840, N834, N357);
or OR2 (N841, N838, N386);
nor NOR4 (N842, N835, N45, N715, N838);
or OR2 (N843, N825, N548);
buf BUF1 (N844, N843);
nor NOR3 (N845, N841, N660, N834);
and AND3 (N846, N816, N498, N756);
xor XOR2 (N847, N839, N578);
nand NAND3 (N848, N842, N281, N115);
buf BUF1 (N849, N813);
and AND4 (N850, N840, N686, N475, N305);
nand NAND3 (N851, N837, N603, N810);
or OR2 (N852, N847, N207);
nor NOR3 (N853, N845, N482, N237);
not NOT1 (N854, N844);
and AND2 (N855, N848, N638);
and AND2 (N856, N846, N152);
not NOT1 (N857, N853);
and AND2 (N858, N855, N36);
buf BUF1 (N859, N851);
nor NOR4 (N860, N832, N70, N3, N585);
or OR3 (N861, N857, N82, N393);
and AND4 (N862, N854, N390, N607, N248);
buf BUF1 (N863, N833);
nor NOR2 (N864, N856, N699);
buf BUF1 (N865, N850);
xor XOR2 (N866, N852, N670);
or OR2 (N867, N866, N501);
buf BUF1 (N868, N858);
nand NAND3 (N869, N862, N722, N381);
nand NAND3 (N870, N863, N737, N75);
nor NOR3 (N871, N861, N41, N441);
nor NOR3 (N872, N864, N137, N320);
and AND3 (N873, N869, N388, N118);
and AND3 (N874, N873, N310, N590);
xor XOR2 (N875, N871, N696);
buf BUF1 (N876, N874);
or OR4 (N877, N865, N668, N290, N63);
nand NAND3 (N878, N870, N140, N273);
or OR2 (N879, N875, N432);
xor XOR2 (N880, N849, N840);
not NOT1 (N881, N867);
nor NOR2 (N882, N868, N284);
and AND4 (N883, N880, N308, N269, N868);
buf BUF1 (N884, N879);
buf BUF1 (N885, N884);
nor NOR4 (N886, N872, N622, N366, N570);
nand NAND2 (N887, N885, N5);
nor NOR3 (N888, N887, N335, N219);
buf BUF1 (N889, N881);
buf BUF1 (N890, N883);
buf BUF1 (N891, N882);
xor XOR2 (N892, N886, N655);
xor XOR2 (N893, N859, N503);
and AND3 (N894, N891, N234, N619);
nor NOR4 (N895, N890, N696, N684, N170);
xor XOR2 (N896, N894, N102);
not NOT1 (N897, N877);
xor XOR2 (N898, N878, N220);
xor XOR2 (N899, N893, N615);
not NOT1 (N900, N896);
nand NAND3 (N901, N898, N134, N681);
buf BUF1 (N902, N901);
or OR4 (N903, N860, N266, N505, N8);
and AND4 (N904, N903, N544, N267, N270);
nand NAND4 (N905, N899, N858, N288, N388);
buf BUF1 (N906, N889);
not NOT1 (N907, N876);
and AND3 (N908, N895, N588, N323);
not NOT1 (N909, N904);
buf BUF1 (N910, N900);
not NOT1 (N911, N908);
xor XOR2 (N912, N907, N841);
not NOT1 (N913, N906);
nor NOR4 (N914, N902, N893, N781, N564);
nand NAND4 (N915, N914, N102, N794, N748);
and AND4 (N916, N892, N782, N219, N615);
buf BUF1 (N917, N912);
nor NOR4 (N918, N916, N452, N828, N400);
xor XOR2 (N919, N909, N531);
and AND3 (N920, N910, N299, N711);
nor NOR4 (N921, N918, N69, N24, N314);
or OR4 (N922, N920, N678, N264, N519);
nand NAND3 (N923, N921, N647, N519);
buf BUF1 (N924, N923);
nor NOR4 (N925, N915, N796, N615, N229);
or OR3 (N926, N917, N781, N781);
buf BUF1 (N927, N888);
nand NAND2 (N928, N926, N364);
xor XOR2 (N929, N925, N890);
or OR3 (N930, N911, N153, N314);
nand NAND4 (N931, N919, N635, N890, N329);
nand NAND4 (N932, N930, N214, N466, N229);
and AND3 (N933, N905, N658, N411);
not NOT1 (N934, N927);
not NOT1 (N935, N897);
or OR4 (N936, N933, N442, N382, N808);
and AND3 (N937, N936, N570, N442);
buf BUF1 (N938, N924);
not NOT1 (N939, N931);
not NOT1 (N940, N939);
nor NOR2 (N941, N934, N477);
and AND4 (N942, N928, N715, N428, N128);
nor NOR3 (N943, N937, N347, N460);
not NOT1 (N944, N932);
or OR2 (N945, N913, N3);
and AND4 (N946, N929, N15, N316, N180);
nand NAND4 (N947, N935, N664, N771, N364);
nor NOR3 (N948, N942, N514, N231);
nor NOR4 (N949, N948, N725, N888, N472);
buf BUF1 (N950, N941);
xor XOR2 (N951, N949, N662);
xor XOR2 (N952, N938, N193);
or OR4 (N953, N950, N102, N951, N449);
nor NOR2 (N954, N75, N134);
buf BUF1 (N955, N940);
buf BUF1 (N956, N947);
and AND2 (N957, N946, N642);
not NOT1 (N958, N957);
or OR3 (N959, N955, N391, N353);
nor NOR3 (N960, N945, N552, N310);
nand NAND2 (N961, N943, N821);
nand NAND4 (N962, N953, N550, N637, N646);
xor XOR2 (N963, N944, N572);
xor XOR2 (N964, N922, N957);
or OR2 (N965, N958, N475);
buf BUF1 (N966, N959);
buf BUF1 (N967, N956);
or OR4 (N968, N952, N102, N450, N502);
not NOT1 (N969, N962);
xor XOR2 (N970, N963, N162);
nand NAND3 (N971, N970, N19, N821);
and AND4 (N972, N965, N399, N960, N909);
nand NAND2 (N973, N40, N341);
not NOT1 (N974, N968);
not NOT1 (N975, N966);
or OR3 (N976, N975, N937, N673);
or OR2 (N977, N967, N544);
buf BUF1 (N978, N973);
nor NOR4 (N979, N969, N426, N70, N463);
nor NOR4 (N980, N977, N769, N742, N77);
nor NOR4 (N981, N961, N548, N777, N612);
or OR3 (N982, N974, N438, N92);
buf BUF1 (N983, N981);
nand NAND3 (N984, N976, N475, N635);
not NOT1 (N985, N980);
and AND4 (N986, N984, N950, N182, N431);
xor XOR2 (N987, N954, N935);
nand NAND3 (N988, N987, N780, N500);
and AND3 (N989, N985, N790, N966);
nand NAND3 (N990, N989, N766, N645);
or OR2 (N991, N972, N96);
and AND3 (N992, N964, N789, N357);
nand NAND2 (N993, N991, N602);
nand NAND4 (N994, N986, N584, N461, N18);
nor NOR4 (N995, N983, N404, N381, N284);
not NOT1 (N996, N995);
nand NAND4 (N997, N971, N742, N632, N809);
nand NAND2 (N998, N996, N543);
or OR2 (N999, N998, N562);
nand NAND3 (N1000, N979, N585, N311);
nor NOR3 (N1001, N999, N723, N938);
xor XOR2 (N1002, N982, N689);
buf BUF1 (N1003, N992);
xor XOR2 (N1004, N990, N260);
xor XOR2 (N1005, N997, N110);
or OR4 (N1006, N1000, N548, N1002, N57);
nand NAND4 (N1007, N567, N282, N161, N162);
xor XOR2 (N1008, N993, N965);
nor NOR2 (N1009, N978, N229);
nor NOR4 (N1010, N1006, N442, N113, N411);
or OR3 (N1011, N1003, N37, N84);
xor XOR2 (N1012, N988, N931);
nor NOR3 (N1013, N1008, N420, N451);
or OR4 (N1014, N1012, N1003, N488, N625);
and AND2 (N1015, N1010, N528);
not NOT1 (N1016, N994);
nand NAND4 (N1017, N1001, N463, N735, N194);
and AND3 (N1018, N1015, N97, N133);
xor XOR2 (N1019, N1005, N844);
nor NOR2 (N1020, N1016, N360);
buf BUF1 (N1021, N1004);
not NOT1 (N1022, N1013);
nor NOR2 (N1023, N1017, N255);
or OR2 (N1024, N1011, N623);
nor NOR3 (N1025, N1022, N544, N882);
and AND3 (N1026, N1007, N534, N910);
buf BUF1 (N1027, N1021);
xor XOR2 (N1028, N1018, N955);
buf BUF1 (N1029, N1026);
not NOT1 (N1030, N1024);
xor XOR2 (N1031, N1023, N124);
nand NAND3 (N1032, N1025, N539, N606);
buf BUF1 (N1033, N1029);
xor XOR2 (N1034, N1027, N372);
buf BUF1 (N1035, N1033);
not NOT1 (N1036, N1032);
xor XOR2 (N1037, N1028, N31);
and AND2 (N1038, N1020, N1034);
not NOT1 (N1039, N896);
buf BUF1 (N1040, N1035);
xor XOR2 (N1041, N1031, N650);
nand NAND2 (N1042, N1038, N286);
buf BUF1 (N1043, N1042);
nand NAND4 (N1044, N1009, N934, N2, N315);
nor NOR2 (N1045, N1036, N883);
xor XOR2 (N1046, N1045, N952);
not NOT1 (N1047, N1014);
and AND3 (N1048, N1041, N512, N646);
and AND2 (N1049, N1043, N600);
not NOT1 (N1050, N1039);
and AND3 (N1051, N1047, N108, N229);
nor NOR3 (N1052, N1030, N297, N116);
not NOT1 (N1053, N1049);
nor NOR2 (N1054, N1048, N573);
and AND3 (N1055, N1019, N957, N1001);
and AND3 (N1056, N1052, N303, N1010);
buf BUF1 (N1057, N1040);
not NOT1 (N1058, N1057);
nor NOR4 (N1059, N1055, N598, N396, N939);
or OR3 (N1060, N1056, N685, N368);
buf BUF1 (N1061, N1051);
and AND3 (N1062, N1037, N256, N573);
xor XOR2 (N1063, N1058, N70);
not NOT1 (N1064, N1059);
buf BUF1 (N1065, N1063);
nand NAND3 (N1066, N1050, N605, N217);
buf BUF1 (N1067, N1062);
buf BUF1 (N1068, N1060);
xor XOR2 (N1069, N1066, N424);
nand NAND3 (N1070, N1053, N789, N185);
or OR2 (N1071, N1065, N645);
not NOT1 (N1072, N1064);
xor XOR2 (N1073, N1072, N161);
or OR2 (N1074, N1069, N740);
not NOT1 (N1075, N1068);
buf BUF1 (N1076, N1067);
or OR2 (N1077, N1074, N307);
buf BUF1 (N1078, N1075);
not NOT1 (N1079, N1046);
nor NOR4 (N1080, N1073, N1019, N480, N803);
xor XOR2 (N1081, N1054, N841);
nand NAND3 (N1082, N1070, N117, N620);
nand NAND3 (N1083, N1044, N574, N54);
or OR3 (N1084, N1071, N650, N954);
nor NOR4 (N1085, N1081, N870, N983, N316);
not NOT1 (N1086, N1061);
and AND4 (N1087, N1080, N548, N814, N316);
or OR3 (N1088, N1086, N180, N816);
not NOT1 (N1089, N1085);
and AND3 (N1090, N1076, N449, N662);
or OR4 (N1091, N1083, N310, N748, N331);
nand NAND4 (N1092, N1088, N569, N827, N672);
buf BUF1 (N1093, N1089);
and AND4 (N1094, N1084, N766, N241, N902);
and AND4 (N1095, N1079, N1062, N1081, N495);
xor XOR2 (N1096, N1091, N381);
or OR4 (N1097, N1094, N113, N289, N207);
nand NAND4 (N1098, N1093, N916, N1074, N556);
nor NOR2 (N1099, N1082, N1057);
nand NAND2 (N1100, N1099, N939);
and AND4 (N1101, N1077, N510, N501, N509);
and AND4 (N1102, N1100, N424, N937, N106);
buf BUF1 (N1103, N1102);
buf BUF1 (N1104, N1078);
xor XOR2 (N1105, N1090, N874);
nor NOR4 (N1106, N1104, N454, N728, N1075);
nand NAND4 (N1107, N1105, N603, N861, N422);
buf BUF1 (N1108, N1087);
or OR2 (N1109, N1092, N213);
nor NOR4 (N1110, N1098, N871, N385, N709);
nor NOR3 (N1111, N1097, N463, N1083);
xor XOR2 (N1112, N1108, N1013);
buf BUF1 (N1113, N1103);
or OR4 (N1114, N1096, N437, N622, N528);
or OR4 (N1115, N1110, N953, N262, N318);
not NOT1 (N1116, N1109);
nor NOR2 (N1117, N1114, N588);
or OR2 (N1118, N1113, N523);
not NOT1 (N1119, N1107);
nor NOR2 (N1120, N1115, N537);
nor NOR2 (N1121, N1117, N232);
or OR4 (N1122, N1118, N668, N233, N560);
or OR2 (N1123, N1122, N766);
not NOT1 (N1124, N1121);
and AND3 (N1125, N1124, N530, N887);
and AND4 (N1126, N1101, N1006, N557, N456);
or OR4 (N1127, N1112, N265, N935, N216);
xor XOR2 (N1128, N1119, N1007);
not NOT1 (N1129, N1123);
not NOT1 (N1130, N1125);
xor XOR2 (N1131, N1128, N1049);
buf BUF1 (N1132, N1126);
buf BUF1 (N1133, N1130);
or OR4 (N1134, N1133, N417, N509, N1006);
or OR2 (N1135, N1129, N402);
not NOT1 (N1136, N1135);
not NOT1 (N1137, N1106);
buf BUF1 (N1138, N1132);
buf BUF1 (N1139, N1127);
and AND3 (N1140, N1116, N578, N378);
nand NAND3 (N1141, N1139, N725, N1076);
nor NOR4 (N1142, N1120, N310, N909, N416);
nor NOR2 (N1143, N1137, N745);
nor NOR3 (N1144, N1095, N742, N1015);
nor NOR2 (N1145, N1141, N981);
nand NAND4 (N1146, N1144, N337, N23, N746);
xor XOR2 (N1147, N1142, N360);
xor XOR2 (N1148, N1143, N516);
buf BUF1 (N1149, N1147);
buf BUF1 (N1150, N1131);
buf BUF1 (N1151, N1150);
not NOT1 (N1152, N1151);
nand NAND4 (N1153, N1148, N587, N970, N1146);
buf BUF1 (N1154, N105);
buf BUF1 (N1155, N1136);
xor XOR2 (N1156, N1155, N679);
nand NAND2 (N1157, N1156, N447);
or OR4 (N1158, N1153, N927, N89, N310);
xor XOR2 (N1159, N1111, N906);
or OR4 (N1160, N1140, N1148, N1085, N1059);
not NOT1 (N1161, N1158);
nor NOR4 (N1162, N1154, N31, N427, N151);
nor NOR4 (N1163, N1134, N969, N655, N176);
xor XOR2 (N1164, N1138, N851);
or OR3 (N1165, N1160, N941, N97);
and AND4 (N1166, N1149, N513, N406, N1142);
nor NOR2 (N1167, N1159, N216);
nor NOR4 (N1168, N1166, N192, N135, N968);
nand NAND4 (N1169, N1152, N196, N37, N926);
buf BUF1 (N1170, N1169);
not NOT1 (N1171, N1163);
or OR4 (N1172, N1167, N867, N1062, N181);
buf BUF1 (N1173, N1172);
or OR2 (N1174, N1173, N293);
nor NOR2 (N1175, N1162, N353);
and AND4 (N1176, N1145, N419, N468, N695);
or OR2 (N1177, N1164, N1000);
nand NAND3 (N1178, N1177, N1160, N904);
nor NOR2 (N1179, N1174, N200);
or OR3 (N1180, N1171, N952, N1100);
or OR2 (N1181, N1180, N203);
or OR4 (N1182, N1178, N1030, N9, N45);
nor NOR2 (N1183, N1157, N298);
or OR4 (N1184, N1165, N121, N1141, N690);
buf BUF1 (N1185, N1182);
buf BUF1 (N1186, N1170);
buf BUF1 (N1187, N1184);
nor NOR2 (N1188, N1179, N232);
xor XOR2 (N1189, N1161, N627);
nor NOR3 (N1190, N1185, N407, N197);
not NOT1 (N1191, N1186);
buf BUF1 (N1192, N1191);
and AND3 (N1193, N1190, N399, N910);
nand NAND3 (N1194, N1189, N805, N708);
nor NOR3 (N1195, N1193, N518, N392);
not NOT1 (N1196, N1175);
xor XOR2 (N1197, N1181, N1187);
nor NOR4 (N1198, N925, N833, N171, N595);
buf BUF1 (N1199, N1183);
xor XOR2 (N1200, N1188, N954);
buf BUF1 (N1201, N1197);
and AND3 (N1202, N1194, N686, N299);
and AND4 (N1203, N1199, N1117, N657, N1176);
or OR2 (N1204, N1166, N1127);
nand NAND3 (N1205, N1198, N937, N207);
buf BUF1 (N1206, N1204);
or OR4 (N1207, N1196, N891, N8, N302);
and AND2 (N1208, N1206, N1062);
buf BUF1 (N1209, N1192);
xor XOR2 (N1210, N1209, N829);
xor XOR2 (N1211, N1205, N171);
and AND2 (N1212, N1201, N863);
nor NOR4 (N1213, N1203, N1001, N606, N238);
and AND4 (N1214, N1213, N963, N532, N403);
not NOT1 (N1215, N1202);
and AND3 (N1216, N1195, N924, N467);
not NOT1 (N1217, N1210);
nand NAND3 (N1218, N1212, N712, N1038);
nand NAND3 (N1219, N1214, N570, N1127);
xor XOR2 (N1220, N1215, N281);
nand NAND2 (N1221, N1220, N1215);
or OR2 (N1222, N1207, N87);
and AND2 (N1223, N1217, N821);
not NOT1 (N1224, N1200);
and AND2 (N1225, N1222, N952);
and AND4 (N1226, N1225, N1149, N888, N61);
nor NOR3 (N1227, N1168, N888, N949);
or OR2 (N1228, N1208, N439);
xor XOR2 (N1229, N1224, N921);
nand NAND4 (N1230, N1219, N1041, N432, N694);
nand NAND4 (N1231, N1223, N507, N726, N830);
xor XOR2 (N1232, N1228, N1228);
and AND2 (N1233, N1231, N905);
buf BUF1 (N1234, N1216);
or OR2 (N1235, N1229, N957);
nand NAND4 (N1236, N1232, N151, N217, N305);
not NOT1 (N1237, N1236);
buf BUF1 (N1238, N1230);
and AND4 (N1239, N1235, N221, N858, N584);
nor NOR4 (N1240, N1211, N728, N374, N1052);
buf BUF1 (N1241, N1234);
nor NOR4 (N1242, N1221, N1156, N1042, N871);
nand NAND2 (N1243, N1226, N1195);
not NOT1 (N1244, N1242);
or OR3 (N1245, N1240, N1242, N418);
and AND2 (N1246, N1243, N624);
xor XOR2 (N1247, N1241, N392);
or OR2 (N1248, N1218, N641);
xor XOR2 (N1249, N1238, N561);
not NOT1 (N1250, N1249);
not NOT1 (N1251, N1227);
or OR3 (N1252, N1246, N736, N804);
and AND3 (N1253, N1244, N846, N785);
not NOT1 (N1254, N1239);
not NOT1 (N1255, N1253);
and AND3 (N1256, N1255, N909, N475);
or OR2 (N1257, N1250, N366);
nor NOR3 (N1258, N1245, N954, N737);
nor NOR2 (N1259, N1256, N45);
or OR4 (N1260, N1248, N774, N1042, N854);
nand NAND3 (N1261, N1259, N520, N251);
nor NOR2 (N1262, N1237, N874);
nand NAND3 (N1263, N1258, N276, N25);
not NOT1 (N1264, N1262);
buf BUF1 (N1265, N1260);
and AND2 (N1266, N1252, N384);
xor XOR2 (N1267, N1266, N829);
xor XOR2 (N1268, N1257, N371);
not NOT1 (N1269, N1265);
buf BUF1 (N1270, N1269);
not NOT1 (N1271, N1267);
not NOT1 (N1272, N1264);
nand NAND3 (N1273, N1270, N398, N646);
not NOT1 (N1274, N1247);
nand NAND3 (N1275, N1268, N708, N1025);
and AND4 (N1276, N1272, N900, N413, N1123);
or OR3 (N1277, N1271, N538, N971);
and AND2 (N1278, N1277, N1177);
and AND4 (N1279, N1274, N837, N313, N248);
not NOT1 (N1280, N1273);
xor XOR2 (N1281, N1251, N402);
not NOT1 (N1282, N1254);
xor XOR2 (N1283, N1233, N972);
nand NAND2 (N1284, N1280, N775);
nor NOR3 (N1285, N1261, N798, N348);
buf BUF1 (N1286, N1284);
or OR4 (N1287, N1282, N1218, N1235, N1145);
not NOT1 (N1288, N1283);
xor XOR2 (N1289, N1278, N792);
nor NOR4 (N1290, N1276, N79, N419, N598);
nand NAND3 (N1291, N1263, N308, N288);
and AND2 (N1292, N1287, N500);
nor NOR4 (N1293, N1286, N1126, N1211, N380);
xor XOR2 (N1294, N1291, N973);
nor NOR3 (N1295, N1288, N680, N799);
nor NOR2 (N1296, N1290, N1131);
xor XOR2 (N1297, N1279, N576);
not NOT1 (N1298, N1289);
xor XOR2 (N1299, N1275, N92);
xor XOR2 (N1300, N1299, N518);
nand NAND4 (N1301, N1292, N993, N640, N416);
buf BUF1 (N1302, N1295);
xor XOR2 (N1303, N1281, N1005);
or OR2 (N1304, N1303, N17);
xor XOR2 (N1305, N1293, N257);
buf BUF1 (N1306, N1296);
xor XOR2 (N1307, N1300, N59);
xor XOR2 (N1308, N1294, N848);
xor XOR2 (N1309, N1307, N8);
nor NOR3 (N1310, N1309, N111, N531);
and AND3 (N1311, N1306, N688, N1228);
nand NAND2 (N1312, N1297, N1054);
not NOT1 (N1313, N1308);
nor NOR4 (N1314, N1304, N642, N365, N1216);
nand NAND4 (N1315, N1310, N718, N120, N1058);
not NOT1 (N1316, N1301);
or OR3 (N1317, N1313, N79, N1175);
nor NOR3 (N1318, N1298, N944, N328);
or OR3 (N1319, N1302, N1152, N504);
nor NOR2 (N1320, N1318, N52);
not NOT1 (N1321, N1311);
or OR4 (N1322, N1317, N375, N1095, N1049);
buf BUF1 (N1323, N1315);
buf BUF1 (N1324, N1285);
not NOT1 (N1325, N1312);
or OR2 (N1326, N1316, N1256);
buf BUF1 (N1327, N1324);
nand NAND4 (N1328, N1326, N589, N779, N738);
buf BUF1 (N1329, N1305);
or OR4 (N1330, N1323, N1155, N960, N124);
or OR2 (N1331, N1322, N42);
or OR4 (N1332, N1329, N433, N15, N589);
buf BUF1 (N1333, N1321);
not NOT1 (N1334, N1330);
nand NAND3 (N1335, N1332, N13, N428);
or OR3 (N1336, N1333, N299, N720);
and AND4 (N1337, N1328, N221, N422, N717);
not NOT1 (N1338, N1337);
buf BUF1 (N1339, N1331);
not NOT1 (N1340, N1339);
and AND2 (N1341, N1335, N747);
not NOT1 (N1342, N1325);
not NOT1 (N1343, N1319);
xor XOR2 (N1344, N1343, N1075);
not NOT1 (N1345, N1341);
nand NAND4 (N1346, N1338, N559, N1088, N965);
buf BUF1 (N1347, N1320);
and AND2 (N1348, N1340, N125);
or OR4 (N1349, N1344, N144, N1169, N446);
or OR4 (N1350, N1327, N480, N490, N1040);
buf BUF1 (N1351, N1342);
buf BUF1 (N1352, N1345);
xor XOR2 (N1353, N1349, N1337);
xor XOR2 (N1354, N1353, N921);
xor XOR2 (N1355, N1351, N868);
not NOT1 (N1356, N1348);
and AND2 (N1357, N1334, N499);
nor NOR4 (N1358, N1336, N58, N818, N710);
or OR2 (N1359, N1357, N392);
and AND3 (N1360, N1358, N1133, N564);
nor NOR3 (N1361, N1354, N898, N21);
buf BUF1 (N1362, N1361);
nor NOR3 (N1363, N1356, N91, N1021);
not NOT1 (N1364, N1359);
or OR3 (N1365, N1355, N824, N17);
nor NOR4 (N1366, N1365, N358, N1096, N102);
and AND2 (N1367, N1362, N271);
not NOT1 (N1368, N1367);
xor XOR2 (N1369, N1346, N242);
not NOT1 (N1370, N1350);
buf BUF1 (N1371, N1366);
nand NAND3 (N1372, N1360, N529, N677);
not NOT1 (N1373, N1363);
xor XOR2 (N1374, N1368, N684);
nor NOR3 (N1375, N1347, N773, N1002);
buf BUF1 (N1376, N1370);
nand NAND2 (N1377, N1371, N471);
nor NOR4 (N1378, N1369, N1082, N1340, N1021);
nand NAND2 (N1379, N1376, N740);
xor XOR2 (N1380, N1364, N718);
not NOT1 (N1381, N1374);
buf BUF1 (N1382, N1372);
buf BUF1 (N1383, N1375);
nor NOR4 (N1384, N1373, N283, N1111, N689);
xor XOR2 (N1385, N1383, N187);
and AND4 (N1386, N1382, N625, N650, N950);
or OR4 (N1387, N1386, N542, N1173, N1178);
nor NOR4 (N1388, N1378, N418, N1351, N292);
buf BUF1 (N1389, N1379);
and AND4 (N1390, N1385, N760, N338, N430);
xor XOR2 (N1391, N1390, N1075);
nor NOR3 (N1392, N1384, N658, N1321);
buf BUF1 (N1393, N1380);
xor XOR2 (N1394, N1388, N105);
buf BUF1 (N1395, N1387);
nor NOR3 (N1396, N1314, N678, N1345);
xor XOR2 (N1397, N1393, N1327);
or OR3 (N1398, N1394, N39, N299);
or OR3 (N1399, N1398, N1344, N1189);
and AND2 (N1400, N1391, N1328);
nor NOR2 (N1401, N1392, N325);
buf BUF1 (N1402, N1399);
nand NAND2 (N1403, N1400, N495);
nand NAND4 (N1404, N1401, N1021, N782, N81);
buf BUF1 (N1405, N1395);
nand NAND4 (N1406, N1404, N392, N1130, N419);
buf BUF1 (N1407, N1406);
buf BUF1 (N1408, N1397);
nor NOR2 (N1409, N1389, N995);
xor XOR2 (N1410, N1381, N614);
and AND3 (N1411, N1402, N772, N250);
buf BUF1 (N1412, N1377);
xor XOR2 (N1413, N1352, N382);
and AND3 (N1414, N1412, N577, N929);
xor XOR2 (N1415, N1405, N887);
not NOT1 (N1416, N1409);
or OR4 (N1417, N1396, N330, N1188, N1268);
and AND3 (N1418, N1407, N331, N1064);
not NOT1 (N1419, N1410);
xor XOR2 (N1420, N1408, N1388);
and AND2 (N1421, N1420, N1344);
or OR2 (N1422, N1403, N563);
nand NAND2 (N1423, N1415, N82);
nor NOR4 (N1424, N1416, N153, N239, N738);
not NOT1 (N1425, N1411);
not NOT1 (N1426, N1417);
and AND4 (N1427, N1422, N323, N1046, N814);
and AND4 (N1428, N1427, N384, N45, N1384);
nand NAND3 (N1429, N1423, N1166, N1322);
and AND2 (N1430, N1421, N246);
xor XOR2 (N1431, N1429, N604);
nor NOR3 (N1432, N1430, N670, N1091);
nor NOR4 (N1433, N1432, N183, N98, N951);
xor XOR2 (N1434, N1418, N433);
nand NAND3 (N1435, N1413, N791, N595);
and AND4 (N1436, N1435, N821, N243, N1229);
and AND2 (N1437, N1426, N504);
not NOT1 (N1438, N1433);
buf BUF1 (N1439, N1419);
nand NAND4 (N1440, N1431, N1179, N1252, N899);
nor NOR3 (N1441, N1424, N350, N949);
and AND3 (N1442, N1437, N952, N333);
or OR4 (N1443, N1425, N882, N679, N301);
xor XOR2 (N1444, N1428, N524);
nor NOR2 (N1445, N1442, N1202);
and AND4 (N1446, N1440, N612, N584, N506);
not NOT1 (N1447, N1434);
nor NOR2 (N1448, N1443, N1080);
and AND4 (N1449, N1414, N1106, N1408, N1131);
nor NOR4 (N1450, N1444, N1162, N1114, N349);
buf BUF1 (N1451, N1436);
buf BUF1 (N1452, N1449);
and AND2 (N1453, N1450, N1177);
nor NOR2 (N1454, N1441, N1401);
xor XOR2 (N1455, N1452, N892);
nand NAND3 (N1456, N1438, N1302, N1426);
buf BUF1 (N1457, N1447);
and AND2 (N1458, N1445, N538);
nand NAND4 (N1459, N1455, N525, N338, N1349);
xor XOR2 (N1460, N1459, N1020);
buf BUF1 (N1461, N1446);
buf BUF1 (N1462, N1461);
or OR3 (N1463, N1456, N332, N1427);
nor NOR3 (N1464, N1457, N978, N904);
and AND3 (N1465, N1463, N475, N654);
or OR3 (N1466, N1460, N1223, N1300);
nand NAND3 (N1467, N1458, N380, N175);
and AND4 (N1468, N1453, N1391, N1379, N504);
nor NOR3 (N1469, N1448, N1220, N1225);
nand NAND3 (N1470, N1451, N1322, N1411);
xor XOR2 (N1471, N1439, N1050);
xor XOR2 (N1472, N1464, N224);
and AND3 (N1473, N1470, N1359, N330);
not NOT1 (N1474, N1468);
nor NOR3 (N1475, N1474, N1099, N1045);
nor NOR3 (N1476, N1475, N140, N1109);
nor NOR2 (N1477, N1471, N843);
nor NOR3 (N1478, N1473, N252, N843);
buf BUF1 (N1479, N1477);
and AND2 (N1480, N1469, N1267);
buf BUF1 (N1481, N1479);
and AND3 (N1482, N1465, N1392, N270);
and AND2 (N1483, N1454, N1155);
not NOT1 (N1484, N1476);
nand NAND3 (N1485, N1484, N766, N604);
nand NAND2 (N1486, N1482, N1339);
not NOT1 (N1487, N1485);
not NOT1 (N1488, N1480);
nand NAND3 (N1489, N1487, N601, N1073);
buf BUF1 (N1490, N1481);
not NOT1 (N1491, N1483);
not NOT1 (N1492, N1472);
nand NAND3 (N1493, N1478, N1292, N1058);
not NOT1 (N1494, N1488);
nand NAND2 (N1495, N1494, N501);
not NOT1 (N1496, N1495);
nor NOR3 (N1497, N1462, N22, N1001);
and AND4 (N1498, N1492, N814, N1006, N704);
xor XOR2 (N1499, N1496, N626);
nor NOR2 (N1500, N1497, N251);
buf BUF1 (N1501, N1499);
and AND3 (N1502, N1489, N333, N1410);
xor XOR2 (N1503, N1467, N962);
buf BUF1 (N1504, N1502);
nand NAND4 (N1505, N1491, N84, N74, N570);
or OR2 (N1506, N1503, N757);
nor NOR4 (N1507, N1500, N1096, N1235, N834);
not NOT1 (N1508, N1504);
and AND4 (N1509, N1505, N235, N1246, N514);
xor XOR2 (N1510, N1509, N864);
buf BUF1 (N1511, N1493);
buf BUF1 (N1512, N1510);
xor XOR2 (N1513, N1506, N697);
or OR2 (N1514, N1490, N900);
nand NAND4 (N1515, N1513, N1028, N825, N585);
and AND2 (N1516, N1486, N256);
xor XOR2 (N1517, N1511, N93);
and AND3 (N1518, N1514, N551, N41);
nand NAND2 (N1519, N1501, N442);
or OR4 (N1520, N1516, N545, N974, N686);
or OR2 (N1521, N1517, N683);
nand NAND4 (N1522, N1498, N787, N410, N1112);
xor XOR2 (N1523, N1520, N606);
and AND4 (N1524, N1522, N238, N1222, N955);
and AND2 (N1525, N1508, N836);
nor NOR2 (N1526, N1507, N763);
or OR2 (N1527, N1521, N977);
not NOT1 (N1528, N1519);
or OR3 (N1529, N1515, N1172, N500);
xor XOR2 (N1530, N1512, N1213);
nor NOR3 (N1531, N1525, N117, N586);
not NOT1 (N1532, N1531);
or OR2 (N1533, N1529, N936);
and AND3 (N1534, N1527, N943, N506);
nand NAND2 (N1535, N1533, N229);
nand NAND3 (N1536, N1523, N1482, N1288);
xor XOR2 (N1537, N1528, N59);
xor XOR2 (N1538, N1537, N768);
nor NOR4 (N1539, N1536, N241, N326, N109);
nor NOR2 (N1540, N1534, N271);
buf BUF1 (N1541, N1535);
xor XOR2 (N1542, N1526, N1025);
or OR4 (N1543, N1532, N851, N275, N1487);
not NOT1 (N1544, N1543);
xor XOR2 (N1545, N1538, N949);
nor NOR2 (N1546, N1539, N1104);
nand NAND2 (N1547, N1544, N893);
nor NOR4 (N1548, N1540, N653, N1199, N703);
and AND3 (N1549, N1548, N466, N872);
and AND2 (N1550, N1547, N585);
and AND3 (N1551, N1466, N766, N760);
nor NOR2 (N1552, N1541, N1130);
nor NOR4 (N1553, N1518, N1122, N1130, N1431);
or OR3 (N1554, N1552, N582, N862);
not NOT1 (N1555, N1551);
not NOT1 (N1556, N1550);
or OR2 (N1557, N1524, N361);
not NOT1 (N1558, N1556);
nand NAND2 (N1559, N1549, N1494);
nand NAND2 (N1560, N1553, N1293);
nor NOR3 (N1561, N1555, N1392, N504);
nand NAND4 (N1562, N1557, N740, N1042, N481);
and AND4 (N1563, N1560, N681, N100, N1348);
buf BUF1 (N1564, N1562);
or OR3 (N1565, N1561, N1341, N508);
xor XOR2 (N1566, N1559, N575);
and AND4 (N1567, N1554, N712, N1357, N1438);
xor XOR2 (N1568, N1546, N1458);
buf BUF1 (N1569, N1564);
not NOT1 (N1570, N1565);
nand NAND4 (N1571, N1567, N261, N34, N652);
or OR4 (N1572, N1563, N203, N587, N740);
nor NOR2 (N1573, N1568, N1308);
xor XOR2 (N1574, N1530, N836);
buf BUF1 (N1575, N1566);
buf BUF1 (N1576, N1574);
xor XOR2 (N1577, N1570, N1203);
and AND2 (N1578, N1545, N1333);
nor NOR3 (N1579, N1576, N246, N98);
xor XOR2 (N1580, N1542, N200);
not NOT1 (N1581, N1580);
not NOT1 (N1582, N1578);
nand NAND3 (N1583, N1575, N867, N258);
nand NAND4 (N1584, N1582, N1000, N533, N1573);
nand NAND2 (N1585, N1546, N966);
not NOT1 (N1586, N1571);
xor XOR2 (N1587, N1584, N1480);
xor XOR2 (N1588, N1585, N339);
or OR4 (N1589, N1569, N822, N789, N1145);
nor NOR2 (N1590, N1587, N528);
nor NOR3 (N1591, N1558, N978, N43);
buf BUF1 (N1592, N1591);
buf BUF1 (N1593, N1592);
buf BUF1 (N1594, N1572);
nand NAND3 (N1595, N1579, N1039, N96);
and AND2 (N1596, N1577, N804);
nor NOR4 (N1597, N1596, N182, N1069, N22);
nand NAND4 (N1598, N1594, N1404, N913, N871);
buf BUF1 (N1599, N1595);
and AND3 (N1600, N1583, N1569, N679);
xor XOR2 (N1601, N1581, N1577);
xor XOR2 (N1602, N1586, N1401);
xor XOR2 (N1603, N1599, N1428);
nor NOR2 (N1604, N1590, N972);
or OR2 (N1605, N1588, N1);
xor XOR2 (N1606, N1589, N330);
nand NAND4 (N1607, N1600, N1050, N714, N293);
xor XOR2 (N1608, N1601, N717);
and AND3 (N1609, N1608, N1096, N181);
nand NAND2 (N1610, N1597, N1210);
buf BUF1 (N1611, N1607);
xor XOR2 (N1612, N1611, N671);
or OR3 (N1613, N1593, N367, N1488);
or OR3 (N1614, N1603, N199, N1031);
or OR4 (N1615, N1605, N209, N300, N327);
endmodule