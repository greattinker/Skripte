// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N12813,N12809,N12787,N12781,N12790,N12812,N12815,N12804,N12800,N12816;

xor XOR2 (N17, N2, N16);
and AND4 (N18, N10, N3, N12, N17);
not NOT1 (N19, N12);
or OR2 (N20, N12, N11);
or OR2 (N21, N15, N8);
buf BUF1 (N22, N21);
not NOT1 (N23, N20);
nor NOR2 (N24, N7, N3);
not NOT1 (N25, N12);
buf BUF1 (N26, N12);
not NOT1 (N27, N13);
or OR4 (N28, N23, N20, N14, N14);
nor NOR4 (N29, N11, N25, N6, N12);
or OR2 (N30, N25, N3);
and AND2 (N31, N12, N24);
not NOT1 (N32, N5);
xor XOR2 (N33, N22, N13);
xor XOR2 (N34, N28, N15);
or OR3 (N35, N34, N13, N26);
or OR3 (N36, N11, N19, N13);
nand NAND3 (N37, N18, N6, N35);
and AND3 (N38, N31, N31, N9);
nor NOR3 (N39, N34, N24, N11);
not NOT1 (N40, N15);
nor NOR2 (N41, N32, N37);
buf BUF1 (N42, N23);
nor NOR2 (N43, N33, N5);
nor NOR2 (N44, N29, N8);
nand NAND3 (N45, N41, N39, N7);
xor XOR2 (N46, N38, N34);
nor NOR4 (N47, N20, N9, N6, N27);
not NOT1 (N48, N25);
nand NAND2 (N49, N40, N15);
or OR4 (N50, N48, N3, N24, N13);
xor XOR2 (N51, N49, N48);
xor XOR2 (N52, N44, N1);
buf BUF1 (N53, N51);
buf BUF1 (N54, N47);
buf BUF1 (N55, N52);
not NOT1 (N56, N53);
not NOT1 (N57, N50);
nand NAND3 (N58, N57, N55, N22);
nand NAND4 (N59, N45, N25, N6, N41);
or OR4 (N60, N21, N8, N45, N18);
nor NOR3 (N61, N30, N22, N37);
nand NAND3 (N62, N58, N41, N30);
xor XOR2 (N63, N61, N23);
and AND3 (N64, N56, N37, N37);
xor XOR2 (N65, N43, N64);
nand NAND2 (N66, N32, N56);
or OR2 (N67, N60, N54);
or OR2 (N68, N44, N15);
nand NAND4 (N69, N67, N34, N21, N54);
and AND4 (N70, N68, N9, N26, N4);
xor XOR2 (N71, N66, N57);
not NOT1 (N72, N63);
or OR4 (N73, N69, N56, N4, N34);
not NOT1 (N74, N65);
xor XOR2 (N75, N42, N55);
buf BUF1 (N76, N62);
buf BUF1 (N77, N70);
nand NAND3 (N78, N72, N22, N60);
not NOT1 (N79, N77);
buf BUF1 (N80, N59);
xor XOR2 (N81, N73, N33);
not NOT1 (N82, N78);
and AND4 (N83, N71, N26, N60, N47);
nor NOR3 (N84, N81, N43, N30);
and AND2 (N85, N83, N42);
not NOT1 (N86, N82);
not NOT1 (N87, N75);
nand NAND2 (N88, N79, N57);
and AND2 (N89, N46, N47);
xor XOR2 (N90, N88, N34);
or OR3 (N91, N36, N23, N55);
and AND4 (N92, N90, N71, N48, N82);
not NOT1 (N93, N85);
not NOT1 (N94, N91);
not NOT1 (N95, N76);
nand NAND2 (N96, N95, N13);
not NOT1 (N97, N94);
and AND3 (N98, N97, N50, N94);
or OR3 (N99, N98, N67, N75);
not NOT1 (N100, N86);
and AND3 (N101, N84, N74, N64);
not NOT1 (N102, N11);
not NOT1 (N103, N100);
not NOT1 (N104, N89);
and AND2 (N105, N102, N64);
not NOT1 (N106, N105);
nand NAND2 (N107, N87, N106);
xor XOR2 (N108, N12, N93);
not NOT1 (N109, N87);
buf BUF1 (N110, N103);
not NOT1 (N111, N99);
nand NAND2 (N112, N96, N49);
and AND2 (N113, N101, N71);
and AND2 (N114, N80, N61);
xor XOR2 (N115, N113, N76);
buf BUF1 (N116, N115);
not NOT1 (N117, N109);
nor NOR4 (N118, N117, N25, N98, N68);
nor NOR2 (N119, N92, N79);
nor NOR3 (N120, N118, N70, N16);
and AND4 (N121, N104, N14, N8, N33);
nand NAND3 (N122, N108, N38, N20);
or OR3 (N123, N116, N16, N111);
xor XOR2 (N124, N73, N81);
buf BUF1 (N125, N122);
and AND4 (N126, N123, N71, N27, N35);
or OR4 (N127, N114, N26, N72, N57);
and AND4 (N128, N112, N6, N2, N77);
buf BUF1 (N129, N121);
or OR2 (N130, N127, N104);
nand NAND2 (N131, N128, N114);
nand NAND4 (N132, N131, N50, N75, N120);
xor XOR2 (N133, N58, N80);
nor NOR2 (N134, N124, N80);
or OR2 (N135, N107, N72);
buf BUF1 (N136, N126);
nor NOR2 (N137, N134, N56);
xor XOR2 (N138, N133, N36);
and AND3 (N139, N119, N75, N10);
not NOT1 (N140, N130);
buf BUF1 (N141, N125);
nor NOR2 (N142, N141, N3);
not NOT1 (N143, N110);
buf BUF1 (N144, N129);
buf BUF1 (N145, N139);
buf BUF1 (N146, N145);
or OR3 (N147, N146, N99, N85);
nand NAND3 (N148, N147, N9, N38);
not NOT1 (N149, N132);
not NOT1 (N150, N136);
or OR3 (N151, N150, N91, N138);
and AND2 (N152, N43, N100);
xor XOR2 (N153, N149, N100);
xor XOR2 (N154, N151, N125);
nand NAND3 (N155, N153, N135, N136);
buf BUF1 (N156, N4);
and AND3 (N157, N148, N71, N108);
nor NOR4 (N158, N152, N97, N21, N52);
or OR2 (N159, N143, N122);
and AND4 (N160, N159, N144, N146, N54);
nand NAND3 (N161, N38, N114, N85);
not NOT1 (N162, N155);
nor NOR2 (N163, N158, N159);
and AND4 (N164, N163, N89, N142, N27);
nor NOR4 (N165, N51, N22, N134, N86);
nor NOR3 (N166, N165, N158, N135);
not NOT1 (N167, N164);
xor XOR2 (N168, N154, N161);
not NOT1 (N169, N20);
or OR2 (N170, N162, N30);
nor NOR4 (N171, N169, N38, N129, N51);
xor XOR2 (N172, N156, N49);
or OR3 (N173, N170, N148, N156);
xor XOR2 (N174, N157, N113);
not NOT1 (N175, N172);
or OR3 (N176, N166, N16, N32);
or OR3 (N177, N140, N115, N29);
buf BUF1 (N178, N174);
nand NAND2 (N179, N173, N115);
xor XOR2 (N180, N167, N129);
nand NAND2 (N181, N179, N1);
buf BUF1 (N182, N171);
and AND4 (N183, N168, N172, N22, N51);
xor XOR2 (N184, N180, N145);
not NOT1 (N185, N137);
nor NOR2 (N186, N160, N171);
or OR2 (N187, N185, N4);
nor NOR4 (N188, N176, N141, N69, N21);
and AND2 (N189, N183, N67);
nand NAND4 (N190, N178, N66, N80, N94);
nand NAND2 (N191, N182, N187);
xor XOR2 (N192, N149, N69);
xor XOR2 (N193, N191, N169);
buf BUF1 (N194, N177);
buf BUF1 (N195, N186);
xor XOR2 (N196, N193, N158);
buf BUF1 (N197, N196);
nand NAND3 (N198, N175, N36, N86);
nor NOR3 (N199, N192, N148, N166);
and AND4 (N200, N195, N181, N130, N33);
buf BUF1 (N201, N54);
nor NOR4 (N202, N190, N192, N109, N52);
or OR2 (N203, N194, N58);
xor XOR2 (N204, N201, N129);
buf BUF1 (N205, N197);
or OR2 (N206, N184, N105);
or OR4 (N207, N205, N8, N172, N60);
xor XOR2 (N208, N188, N177);
nand NAND4 (N209, N198, N203, N136, N116);
or OR2 (N210, N122, N70);
not NOT1 (N211, N204);
xor XOR2 (N212, N211, N50);
nor NOR4 (N213, N189, N40, N137, N48);
or OR4 (N214, N209, N152, N204, N31);
not NOT1 (N215, N212);
and AND2 (N216, N210, N170);
not NOT1 (N217, N208);
not NOT1 (N218, N216);
and AND2 (N219, N214, N51);
xor XOR2 (N220, N219, N78);
buf BUF1 (N221, N213);
nand NAND4 (N222, N220, N89, N47, N186);
nor NOR2 (N223, N202, N8);
or OR2 (N224, N199, N203);
nand NAND3 (N225, N215, N8, N193);
or OR2 (N226, N224, N188);
not NOT1 (N227, N207);
and AND4 (N228, N221, N198, N67, N60);
nor NOR4 (N229, N218, N165, N218, N185);
nor NOR3 (N230, N206, N68, N104);
buf BUF1 (N231, N222);
nor NOR4 (N232, N228, N44, N191, N53);
nor NOR4 (N233, N230, N148, N186, N118);
not NOT1 (N234, N226);
not NOT1 (N235, N223);
nand NAND3 (N236, N229, N225, N48);
not NOT1 (N237, N204);
and AND4 (N238, N232, N202, N234, N16);
and AND2 (N239, N180, N120);
nor NOR4 (N240, N227, N106, N138, N28);
not NOT1 (N241, N233);
nand NAND2 (N242, N237, N76);
buf BUF1 (N243, N241);
buf BUF1 (N244, N200);
nor NOR3 (N245, N242, N38, N91);
buf BUF1 (N246, N238);
buf BUF1 (N247, N235);
nand NAND3 (N248, N240, N148, N211);
nand NAND3 (N249, N239, N66, N138);
nand NAND2 (N250, N249, N51);
nor NOR3 (N251, N236, N18, N12);
not NOT1 (N252, N245);
not NOT1 (N253, N246);
xor XOR2 (N254, N252, N64);
buf BUF1 (N255, N247);
not NOT1 (N256, N253);
xor XOR2 (N257, N255, N30);
not NOT1 (N258, N248);
or OR4 (N259, N254, N246, N29, N130);
or OR3 (N260, N257, N188, N14);
and AND4 (N261, N259, N65, N85, N259);
nand NAND4 (N262, N260, N147, N171, N34);
xor XOR2 (N263, N256, N87);
and AND3 (N264, N263, N199, N112);
nand NAND4 (N265, N250, N167, N31, N132);
or OR2 (N266, N231, N87);
and AND4 (N267, N217, N126, N57, N118);
xor XOR2 (N268, N261, N233);
nand NAND2 (N269, N266, N2);
not NOT1 (N270, N262);
nand NAND3 (N271, N264, N208, N198);
buf BUF1 (N272, N243);
not NOT1 (N273, N268);
and AND3 (N274, N272, N267, N190);
and AND3 (N275, N190, N7, N138);
and AND4 (N276, N273, N247, N5, N7);
buf BUF1 (N277, N275);
nand NAND2 (N278, N258, N157);
or OR3 (N279, N274, N222, N234);
xor XOR2 (N280, N251, N5);
or OR3 (N281, N280, N163, N239);
buf BUF1 (N282, N271);
buf BUF1 (N283, N277);
nand NAND2 (N284, N276, N54);
buf BUF1 (N285, N265);
nand NAND3 (N286, N281, N39, N232);
nand NAND2 (N287, N279, N163);
not NOT1 (N288, N244);
nor NOR4 (N289, N286, N168, N46, N115);
xor XOR2 (N290, N270, N69);
nor NOR3 (N291, N282, N4, N109);
not NOT1 (N292, N285);
and AND4 (N293, N290, N2, N10, N187);
xor XOR2 (N294, N287, N94);
xor XOR2 (N295, N288, N26);
or OR4 (N296, N289, N94, N238, N51);
and AND4 (N297, N278, N97, N106, N285);
not NOT1 (N298, N294);
nand NAND4 (N299, N297, N157, N92, N9);
nand NAND2 (N300, N293, N25);
nor NOR2 (N301, N292, N174);
xor XOR2 (N302, N301, N249);
or OR2 (N303, N296, N79);
buf BUF1 (N304, N300);
or OR2 (N305, N291, N147);
buf BUF1 (N306, N269);
nor NOR4 (N307, N304, N302, N138, N223);
or OR4 (N308, N143, N104, N148, N255);
nor NOR2 (N309, N307, N75);
buf BUF1 (N310, N309);
nand NAND4 (N311, N284, N229, N137, N229);
buf BUF1 (N312, N310);
not NOT1 (N313, N311);
and AND4 (N314, N312, N167, N33, N293);
buf BUF1 (N315, N295);
nor NOR2 (N316, N305, N49);
nand NAND3 (N317, N303, N184, N175);
or OR2 (N318, N299, N231);
xor XOR2 (N319, N317, N60);
nand NAND2 (N320, N315, N214);
nor NOR4 (N321, N313, N138, N221, N191);
or OR3 (N322, N283, N140, N231);
buf BUF1 (N323, N306);
not NOT1 (N324, N308);
and AND3 (N325, N298, N202, N178);
not NOT1 (N326, N325);
or OR2 (N327, N322, N315);
nor NOR2 (N328, N324, N182);
not NOT1 (N329, N327);
nand NAND2 (N330, N329, N80);
nor NOR3 (N331, N319, N189, N128);
nand NAND2 (N332, N318, N309);
not NOT1 (N333, N323);
nand NAND3 (N334, N328, N332, N159);
xor XOR2 (N335, N306, N97);
buf BUF1 (N336, N335);
nor NOR3 (N337, N331, N168, N251);
buf BUF1 (N338, N333);
nand NAND4 (N339, N316, N113, N183, N228);
and AND4 (N340, N326, N221, N50, N152);
buf BUF1 (N341, N338);
or OR3 (N342, N314, N267, N289);
or OR2 (N343, N337, N328);
not NOT1 (N344, N330);
buf BUF1 (N345, N344);
nor NOR3 (N346, N343, N289, N332);
and AND4 (N347, N345, N28, N105, N209);
or OR3 (N348, N339, N111, N6);
not NOT1 (N349, N348);
nand NAND4 (N350, N346, N173, N251, N128);
buf BUF1 (N351, N340);
buf BUF1 (N352, N342);
nand NAND4 (N353, N352, N117, N210, N345);
buf BUF1 (N354, N350);
or OR3 (N355, N354, N329, N200);
or OR3 (N356, N336, N164, N135);
buf BUF1 (N357, N347);
and AND4 (N358, N355, N138, N210, N18);
not NOT1 (N359, N320);
not NOT1 (N360, N358);
and AND3 (N361, N359, N322, N271);
not NOT1 (N362, N361);
and AND3 (N363, N360, N163, N271);
nand NAND3 (N364, N363, N158, N363);
xor XOR2 (N365, N357, N13);
not NOT1 (N366, N349);
xor XOR2 (N367, N365, N14);
nor NOR2 (N368, N341, N290);
xor XOR2 (N369, N321, N263);
nand NAND3 (N370, N367, N70, N308);
nor NOR4 (N371, N366, N351, N339, N69);
xor XOR2 (N372, N100, N204);
xor XOR2 (N373, N370, N91);
or OR2 (N374, N369, N62);
nand NAND4 (N375, N368, N116, N111, N239);
buf BUF1 (N376, N373);
xor XOR2 (N377, N375, N315);
nor NOR2 (N378, N372, N284);
nand NAND3 (N379, N334, N180, N182);
nor NOR3 (N380, N353, N44, N226);
nand NAND3 (N381, N380, N248, N33);
and AND3 (N382, N371, N156, N213);
nor NOR4 (N383, N381, N165, N327, N13);
xor XOR2 (N384, N364, N381);
not NOT1 (N385, N383);
not NOT1 (N386, N385);
or OR2 (N387, N374, N86);
xor XOR2 (N388, N382, N63);
not NOT1 (N389, N378);
nor NOR4 (N390, N377, N312, N236, N229);
xor XOR2 (N391, N376, N83);
nor NOR4 (N392, N386, N139, N129, N31);
buf BUF1 (N393, N391);
buf BUF1 (N394, N387);
xor XOR2 (N395, N362, N82);
or OR4 (N396, N388, N212, N318, N345);
buf BUF1 (N397, N394);
xor XOR2 (N398, N389, N26);
and AND2 (N399, N379, N254);
buf BUF1 (N400, N395);
and AND3 (N401, N397, N263, N11);
and AND3 (N402, N356, N35, N305);
nor NOR4 (N403, N390, N248, N370, N287);
nand NAND3 (N404, N393, N259, N174);
nand NAND2 (N405, N396, N98);
nor NOR3 (N406, N384, N38, N31);
and AND2 (N407, N399, N242);
buf BUF1 (N408, N404);
not NOT1 (N409, N408);
xor XOR2 (N410, N398, N310);
buf BUF1 (N411, N409);
xor XOR2 (N412, N400, N121);
not NOT1 (N413, N402);
or OR4 (N414, N410, N264, N281, N276);
nand NAND2 (N415, N405, N242);
nor NOR4 (N416, N412, N70, N353, N389);
and AND4 (N417, N411, N400, N49, N45);
nor NOR4 (N418, N406, N74, N2, N9);
and AND3 (N419, N414, N383, N247);
nand NAND3 (N420, N407, N113, N377);
or OR4 (N421, N413, N267, N185, N183);
or OR3 (N422, N421, N346, N2);
nand NAND3 (N423, N416, N92, N260);
not NOT1 (N424, N392);
and AND2 (N425, N422, N237);
nand NAND2 (N426, N425, N373);
xor XOR2 (N427, N419, N18);
nand NAND3 (N428, N418, N117, N366);
and AND4 (N429, N417, N50, N389, N277);
xor XOR2 (N430, N403, N26);
and AND2 (N431, N428, N424);
and AND3 (N432, N130, N198, N299);
buf BUF1 (N433, N426);
xor XOR2 (N434, N401, N311);
nor NOR2 (N435, N427, N72);
xor XOR2 (N436, N430, N327);
or OR4 (N437, N434, N417, N298, N231);
and AND2 (N438, N435, N361);
xor XOR2 (N439, N415, N386);
or OR3 (N440, N439, N301, N274);
or OR2 (N441, N429, N268);
buf BUF1 (N442, N437);
buf BUF1 (N443, N433);
nand NAND2 (N444, N436, N238);
and AND2 (N445, N443, N336);
nand NAND3 (N446, N440, N240, N293);
nand NAND3 (N447, N442, N256, N136);
not NOT1 (N448, N423);
xor XOR2 (N449, N438, N340);
not NOT1 (N450, N441);
xor XOR2 (N451, N420, N31);
xor XOR2 (N452, N431, N103);
nor NOR2 (N453, N447, N170);
buf BUF1 (N454, N450);
nor NOR4 (N455, N445, N423, N129, N223);
not NOT1 (N456, N453);
nand NAND2 (N457, N452, N230);
or OR2 (N458, N446, N209);
nor NOR4 (N459, N444, N230, N345, N268);
and AND3 (N460, N457, N172, N325);
nand NAND4 (N461, N451, N150, N228, N83);
and AND2 (N462, N432, N444);
xor XOR2 (N463, N455, N454);
buf BUF1 (N464, N11);
or OR4 (N465, N459, N282, N69, N190);
xor XOR2 (N466, N449, N3);
or OR2 (N467, N456, N371);
and AND2 (N468, N467, N379);
not NOT1 (N469, N461);
or OR4 (N470, N468, N366, N269, N255);
nand NAND3 (N471, N458, N354, N71);
or OR2 (N472, N448, N381);
buf BUF1 (N473, N462);
xor XOR2 (N474, N471, N179);
or OR2 (N475, N473, N222);
nor NOR3 (N476, N464, N39, N264);
or OR3 (N477, N466, N463, N201);
not NOT1 (N478, N208);
xor XOR2 (N479, N476, N318);
not NOT1 (N480, N472);
not NOT1 (N481, N469);
and AND4 (N482, N465, N381, N46, N223);
nand NAND3 (N483, N470, N345, N321);
or OR4 (N484, N460, N49, N38, N20);
or OR4 (N485, N483, N480, N79, N3);
and AND4 (N486, N174, N183, N472, N254);
nand NAND4 (N487, N479, N252, N123, N230);
xor XOR2 (N488, N475, N227);
or OR3 (N489, N487, N309, N255);
nand NAND4 (N490, N474, N18, N93, N430);
nand NAND4 (N491, N482, N10, N387, N329);
nor NOR4 (N492, N488, N153, N218, N455);
not NOT1 (N493, N481);
xor XOR2 (N494, N485, N315);
nand NAND3 (N495, N494, N8, N57);
and AND3 (N496, N492, N54, N212);
xor XOR2 (N497, N496, N275);
nor NOR2 (N498, N493, N112);
buf BUF1 (N499, N478);
buf BUF1 (N500, N489);
xor XOR2 (N501, N500, N265);
and AND4 (N502, N497, N70, N343, N288);
buf BUF1 (N503, N498);
nor NOR3 (N504, N491, N41, N49);
not NOT1 (N505, N495);
nand NAND4 (N506, N490, N464, N209, N136);
or OR4 (N507, N504, N106, N346, N154);
nor NOR2 (N508, N507, N453);
buf BUF1 (N509, N501);
or OR2 (N510, N506, N315);
nand NAND4 (N511, N499, N323, N21, N372);
xor XOR2 (N512, N509, N246);
buf BUF1 (N513, N508);
nor NOR4 (N514, N510, N32, N448, N233);
or OR4 (N515, N477, N506, N465, N228);
buf BUF1 (N516, N513);
nand NAND3 (N517, N514, N507, N93);
xor XOR2 (N518, N502, N13);
or OR2 (N519, N515, N247);
xor XOR2 (N520, N516, N400);
nor NOR3 (N521, N519, N128, N236);
buf BUF1 (N522, N505);
xor XOR2 (N523, N518, N59);
nor NOR4 (N524, N484, N81, N285, N246);
or OR3 (N525, N511, N306, N220);
xor XOR2 (N526, N522, N65);
or OR4 (N527, N524, N436, N486, N280);
or OR2 (N528, N247, N431);
or OR2 (N529, N527, N147);
nand NAND2 (N530, N517, N68);
and AND2 (N531, N530, N121);
or OR4 (N532, N503, N176, N365, N207);
or OR3 (N533, N520, N72, N441);
not NOT1 (N534, N529);
buf BUF1 (N535, N525);
or OR2 (N536, N526, N432);
or OR3 (N537, N531, N11, N328);
nor NOR3 (N538, N536, N92, N61);
nand NAND3 (N539, N532, N450, N269);
nand NAND2 (N540, N512, N62);
not NOT1 (N541, N535);
not NOT1 (N542, N534);
nand NAND4 (N543, N538, N477, N279, N528);
not NOT1 (N544, N163);
not NOT1 (N545, N523);
nand NAND4 (N546, N542, N325, N204, N372);
nor NOR4 (N547, N543, N160, N379, N469);
not NOT1 (N548, N541);
and AND2 (N549, N548, N488);
not NOT1 (N550, N539);
nand NAND2 (N551, N537, N319);
or OR4 (N552, N546, N113, N244, N150);
nand NAND2 (N553, N549, N81);
xor XOR2 (N554, N545, N356);
nor NOR3 (N555, N521, N364, N482);
or OR2 (N556, N553, N544);
xor XOR2 (N557, N465, N165);
or OR2 (N558, N557, N281);
nand NAND2 (N559, N540, N133);
and AND2 (N560, N533, N54);
and AND2 (N561, N547, N307);
buf BUF1 (N562, N552);
or OR2 (N563, N562, N295);
or OR2 (N564, N561, N273);
not NOT1 (N565, N550);
or OR3 (N566, N565, N540, N222);
buf BUF1 (N567, N554);
nor NOR3 (N568, N555, N433, N98);
nand NAND2 (N569, N568, N51);
not NOT1 (N570, N556);
buf BUF1 (N571, N551);
nor NOR3 (N572, N560, N485, N475);
and AND2 (N573, N572, N216);
not NOT1 (N574, N571);
buf BUF1 (N575, N559);
nand NAND3 (N576, N573, N529, N490);
nand NAND2 (N577, N570, N197);
nand NAND3 (N578, N569, N389, N414);
nand NAND4 (N579, N558, N335, N499, N440);
nor NOR3 (N580, N576, N568, N89);
or OR3 (N581, N563, N498, N531);
or OR2 (N582, N578, N204);
buf BUF1 (N583, N574);
nand NAND3 (N584, N581, N215, N138);
nand NAND2 (N585, N582, N455);
and AND4 (N586, N577, N18, N71, N349);
not NOT1 (N587, N586);
not NOT1 (N588, N579);
or OR4 (N589, N584, N322, N337, N397);
not NOT1 (N590, N588);
xor XOR2 (N591, N564, N185);
xor XOR2 (N592, N587, N439);
buf BUF1 (N593, N589);
buf BUF1 (N594, N593);
buf BUF1 (N595, N591);
not NOT1 (N596, N583);
nor NOR2 (N597, N595, N399);
xor XOR2 (N598, N597, N365);
and AND2 (N599, N580, N394);
or OR3 (N600, N566, N73, N398);
xor XOR2 (N601, N592, N65);
nor NOR3 (N602, N598, N455, N228);
not NOT1 (N603, N575);
or OR4 (N604, N594, N182, N130, N136);
and AND2 (N605, N599, N345);
buf BUF1 (N606, N585);
not NOT1 (N607, N605);
nand NAND3 (N608, N606, N606, N177);
nand NAND2 (N609, N608, N537);
and AND2 (N610, N609, N320);
nand NAND2 (N611, N603, N66);
and AND2 (N612, N567, N550);
buf BUF1 (N613, N602);
buf BUF1 (N614, N612);
not NOT1 (N615, N604);
xor XOR2 (N616, N611, N583);
or OR4 (N617, N614, N313, N66, N614);
or OR3 (N618, N616, N531, N540);
not NOT1 (N619, N610);
xor XOR2 (N620, N596, N493);
not NOT1 (N621, N618);
nand NAND4 (N622, N590, N81, N214, N442);
and AND4 (N623, N617, N413, N299, N148);
nor NOR3 (N624, N613, N525, N461);
or OR2 (N625, N600, N285);
nand NAND3 (N626, N620, N305, N501);
buf BUF1 (N627, N619);
not NOT1 (N628, N627);
and AND2 (N629, N622, N46);
nand NAND2 (N630, N629, N552);
or OR4 (N631, N615, N382, N149, N394);
and AND3 (N632, N621, N586, N476);
nand NAND3 (N633, N601, N278, N16);
xor XOR2 (N634, N632, N607);
not NOT1 (N635, N268);
and AND2 (N636, N623, N63);
nor NOR4 (N637, N624, N574, N184, N226);
nand NAND2 (N638, N633, N485);
xor XOR2 (N639, N626, N224);
xor XOR2 (N640, N631, N82);
nor NOR2 (N641, N637, N113);
not NOT1 (N642, N628);
nor NOR4 (N643, N641, N95, N278, N641);
buf BUF1 (N644, N643);
buf BUF1 (N645, N640);
nor NOR3 (N646, N644, N556, N347);
nand NAND4 (N647, N625, N319, N322, N4);
nand NAND3 (N648, N642, N415, N562);
not NOT1 (N649, N645);
not NOT1 (N650, N630);
buf BUF1 (N651, N650);
nand NAND4 (N652, N639, N2, N327, N398);
not NOT1 (N653, N649);
nand NAND2 (N654, N651, N184);
buf BUF1 (N655, N634);
or OR2 (N656, N653, N210);
buf BUF1 (N657, N652);
nor NOR2 (N658, N656, N579);
nor NOR3 (N659, N654, N8, N633);
or OR4 (N660, N635, N352, N424, N220);
nor NOR4 (N661, N657, N80, N57, N464);
and AND2 (N662, N648, N351);
or OR3 (N663, N655, N576, N453);
and AND2 (N664, N646, N414);
or OR4 (N665, N660, N54, N20, N263);
xor XOR2 (N666, N659, N465);
or OR2 (N667, N662, N170);
nand NAND2 (N668, N636, N438);
nor NOR2 (N669, N667, N567);
nand NAND3 (N670, N665, N289, N633);
and AND4 (N671, N663, N553, N604, N495);
nor NOR3 (N672, N638, N628, N317);
xor XOR2 (N673, N647, N361);
buf BUF1 (N674, N658);
nand NAND3 (N675, N669, N349, N523);
xor XOR2 (N676, N673, N626);
nor NOR4 (N677, N672, N496, N648, N187);
nand NAND4 (N678, N676, N248, N529, N239);
or OR4 (N679, N671, N209, N618, N652);
or OR4 (N680, N661, N468, N145, N388);
or OR3 (N681, N668, N595, N431);
xor XOR2 (N682, N677, N572);
nor NOR2 (N683, N680, N415);
nand NAND2 (N684, N678, N343);
or OR4 (N685, N670, N8, N26, N550);
or OR4 (N686, N674, N468, N66, N573);
not NOT1 (N687, N684);
nor NOR2 (N688, N664, N190);
and AND2 (N689, N681, N169);
or OR4 (N690, N688, N99, N439, N146);
or OR4 (N691, N687, N347, N577, N196);
nor NOR2 (N692, N690, N649);
not NOT1 (N693, N685);
and AND2 (N694, N689, N63);
nand NAND4 (N695, N682, N531, N360, N595);
nand NAND4 (N696, N686, N491, N554, N367);
not NOT1 (N697, N691);
xor XOR2 (N698, N679, N245);
xor XOR2 (N699, N697, N509);
or OR4 (N700, N693, N150, N288, N330);
or OR2 (N701, N694, N137);
nor NOR3 (N702, N698, N384, N9);
and AND2 (N703, N699, N366);
xor XOR2 (N704, N696, N590);
nor NOR3 (N705, N704, N642, N491);
not NOT1 (N706, N701);
or OR4 (N707, N666, N438, N534, N530);
and AND4 (N708, N692, N590, N255, N529);
not NOT1 (N709, N708);
or OR2 (N710, N707, N469);
nand NAND4 (N711, N702, N304, N619, N171);
buf BUF1 (N712, N706);
and AND3 (N713, N675, N271, N89);
nor NOR3 (N714, N710, N551, N31);
nand NAND3 (N715, N705, N706, N4);
buf BUF1 (N716, N703);
not NOT1 (N717, N711);
and AND3 (N718, N712, N192, N40);
or OR2 (N719, N717, N653);
xor XOR2 (N720, N719, N173);
nand NAND2 (N721, N700, N412);
not NOT1 (N722, N714);
xor XOR2 (N723, N716, N160);
or OR4 (N724, N713, N442, N648, N101);
or OR2 (N725, N715, N631);
xor XOR2 (N726, N683, N159);
buf BUF1 (N727, N725);
xor XOR2 (N728, N727, N133);
nor NOR4 (N729, N721, N205, N453, N194);
xor XOR2 (N730, N722, N315);
nand NAND4 (N731, N726, N63, N478, N53);
not NOT1 (N732, N718);
or OR2 (N733, N732, N586);
buf BUF1 (N734, N723);
or OR4 (N735, N729, N180, N383, N712);
xor XOR2 (N736, N735, N505);
nand NAND3 (N737, N734, N470, N581);
buf BUF1 (N738, N730);
buf BUF1 (N739, N709);
xor XOR2 (N740, N737, N318);
or OR2 (N741, N733, N426);
nand NAND4 (N742, N728, N464, N317, N296);
or OR2 (N743, N740, N204);
nor NOR3 (N744, N743, N261, N711);
nand NAND2 (N745, N741, N379);
or OR4 (N746, N744, N610, N487, N68);
and AND3 (N747, N739, N573, N492);
buf BUF1 (N748, N695);
or OR2 (N749, N748, N692);
xor XOR2 (N750, N747, N641);
buf BUF1 (N751, N720);
not NOT1 (N752, N750);
nand NAND3 (N753, N745, N30, N47);
buf BUF1 (N754, N736);
nor NOR4 (N755, N751, N89, N111, N280);
and AND2 (N756, N754, N29);
not NOT1 (N757, N746);
buf BUF1 (N758, N753);
xor XOR2 (N759, N752, N697);
not NOT1 (N760, N738);
or OR4 (N761, N731, N426, N100, N659);
xor XOR2 (N762, N742, N493);
nand NAND2 (N763, N755, N342);
xor XOR2 (N764, N756, N487);
nor NOR3 (N765, N763, N680, N600);
nor NOR3 (N766, N760, N539, N291);
buf BUF1 (N767, N757);
xor XOR2 (N768, N759, N579);
or OR2 (N769, N758, N279);
not NOT1 (N770, N766);
nor NOR4 (N771, N749, N424, N292, N744);
not NOT1 (N772, N771);
nor NOR3 (N773, N769, N555, N11);
not NOT1 (N774, N767);
xor XOR2 (N775, N724, N692);
nand NAND4 (N776, N768, N503, N355, N617);
or OR4 (N777, N761, N688, N756, N82);
and AND3 (N778, N775, N280, N110);
buf BUF1 (N779, N770);
nor NOR2 (N780, N773, N650);
xor XOR2 (N781, N776, N32);
buf BUF1 (N782, N762);
buf BUF1 (N783, N765);
xor XOR2 (N784, N782, N85);
xor XOR2 (N785, N764, N377);
nand NAND3 (N786, N780, N531, N651);
nand NAND2 (N787, N785, N64);
nor NOR3 (N788, N774, N658, N396);
buf BUF1 (N789, N778);
nand NAND3 (N790, N788, N472, N704);
not NOT1 (N791, N784);
not NOT1 (N792, N783);
not NOT1 (N793, N789);
and AND4 (N794, N791, N192, N155, N468);
or OR4 (N795, N790, N182, N19, N35);
xor XOR2 (N796, N787, N516);
nor NOR4 (N797, N795, N383, N181, N688);
nand NAND3 (N798, N793, N52, N785);
xor XOR2 (N799, N792, N447);
xor XOR2 (N800, N797, N78);
or OR4 (N801, N777, N646, N761, N520);
nand NAND3 (N802, N772, N23, N281);
and AND4 (N803, N800, N554, N342, N386);
not NOT1 (N804, N779);
or OR2 (N805, N786, N425);
nor NOR2 (N806, N798, N131);
nand NAND3 (N807, N805, N764, N327);
buf BUF1 (N808, N801);
and AND3 (N809, N781, N56, N460);
and AND2 (N810, N808, N377);
and AND2 (N811, N807, N775);
or OR3 (N812, N811, N754, N252);
nor NOR3 (N813, N809, N447, N763);
buf BUF1 (N814, N810);
not NOT1 (N815, N794);
buf BUF1 (N816, N803);
or OR2 (N817, N804, N66);
and AND2 (N818, N806, N236);
xor XOR2 (N819, N815, N616);
not NOT1 (N820, N814);
nand NAND3 (N821, N813, N694, N780);
nand NAND4 (N822, N819, N24, N119, N31);
nand NAND2 (N823, N821, N10);
nor NOR2 (N824, N796, N294);
and AND2 (N825, N818, N84);
nand NAND2 (N826, N817, N162);
or OR3 (N827, N825, N381, N771);
or OR4 (N828, N802, N107, N26, N81);
nor NOR4 (N829, N827, N82, N746, N115);
nand NAND3 (N830, N826, N127, N318);
or OR2 (N831, N799, N476);
buf BUF1 (N832, N812);
xor XOR2 (N833, N820, N102);
not NOT1 (N834, N822);
xor XOR2 (N835, N831, N480);
buf BUF1 (N836, N824);
xor XOR2 (N837, N816, N828);
nor NOR3 (N838, N410, N436, N573);
xor XOR2 (N839, N834, N147);
not NOT1 (N840, N839);
or OR4 (N841, N835, N10, N801, N752);
buf BUF1 (N842, N830);
not NOT1 (N843, N841);
nor NOR2 (N844, N836, N823);
not NOT1 (N845, N636);
nand NAND3 (N846, N838, N347, N563);
nand NAND3 (N847, N842, N358, N307);
not NOT1 (N848, N844);
or OR4 (N849, N832, N125, N140, N696);
buf BUF1 (N850, N843);
nor NOR2 (N851, N840, N87);
buf BUF1 (N852, N849);
buf BUF1 (N853, N846);
and AND2 (N854, N847, N797);
nor NOR3 (N855, N837, N286, N31);
nor NOR2 (N856, N855, N417);
and AND2 (N857, N854, N285);
buf BUF1 (N858, N851);
nand NAND3 (N859, N852, N674, N740);
not NOT1 (N860, N857);
xor XOR2 (N861, N829, N331);
or OR4 (N862, N853, N613, N179, N411);
or OR2 (N863, N862, N150);
buf BUF1 (N864, N858);
buf BUF1 (N865, N856);
buf BUF1 (N866, N859);
nor NOR4 (N867, N845, N670, N188, N281);
and AND4 (N868, N865, N674, N716, N569);
xor XOR2 (N869, N866, N732);
or OR4 (N870, N869, N630, N341, N202);
xor XOR2 (N871, N848, N592);
not NOT1 (N872, N870);
nor NOR2 (N873, N863, N357);
buf BUF1 (N874, N868);
or OR2 (N875, N861, N833);
or OR3 (N876, N90, N639, N611);
or OR2 (N877, N864, N666);
and AND4 (N878, N860, N869, N212, N641);
not NOT1 (N879, N873);
nand NAND2 (N880, N876, N31);
buf BUF1 (N881, N872);
nand NAND2 (N882, N881, N230);
or OR2 (N883, N871, N72);
nor NOR3 (N884, N874, N117, N180);
nand NAND4 (N885, N879, N673, N80, N703);
nor NOR2 (N886, N867, N192);
nand NAND3 (N887, N880, N471, N194);
xor XOR2 (N888, N885, N402);
not NOT1 (N889, N886);
or OR2 (N890, N883, N344);
or OR4 (N891, N875, N544, N793, N87);
buf BUF1 (N892, N884);
xor XOR2 (N893, N888, N827);
nand NAND4 (N894, N878, N121, N185, N217);
xor XOR2 (N895, N892, N878);
not NOT1 (N896, N889);
nand NAND2 (N897, N882, N884);
xor XOR2 (N898, N897, N644);
xor XOR2 (N899, N890, N776);
xor XOR2 (N900, N899, N517);
not NOT1 (N901, N891);
nand NAND3 (N902, N898, N355, N99);
not NOT1 (N903, N850);
xor XOR2 (N904, N893, N833);
nand NAND3 (N905, N896, N241, N880);
or OR3 (N906, N877, N229, N522);
nand NAND4 (N907, N902, N820, N316, N148);
nand NAND4 (N908, N887, N432, N218, N160);
buf BUF1 (N909, N905);
or OR3 (N910, N907, N11, N676);
nor NOR3 (N911, N906, N906, N567);
or OR4 (N912, N904, N315, N160, N702);
not NOT1 (N913, N900);
or OR3 (N914, N913, N523, N284);
not NOT1 (N915, N910);
xor XOR2 (N916, N909, N317);
not NOT1 (N917, N911);
buf BUF1 (N918, N908);
and AND3 (N919, N917, N123, N59);
nor NOR4 (N920, N895, N676, N504, N636);
and AND4 (N921, N916, N719, N149, N152);
nand NAND3 (N922, N920, N491, N888);
or OR4 (N923, N901, N888, N68, N856);
nand NAND4 (N924, N912, N505, N730, N906);
buf BUF1 (N925, N924);
buf BUF1 (N926, N894);
and AND3 (N927, N903, N920, N586);
or OR3 (N928, N923, N793, N446);
nor NOR3 (N929, N918, N478, N135);
nand NAND4 (N930, N928, N152, N109, N645);
xor XOR2 (N931, N922, N680);
nand NAND2 (N932, N927, N600);
or OR4 (N933, N929, N518, N385, N874);
xor XOR2 (N934, N933, N490);
not NOT1 (N935, N930);
nand NAND2 (N936, N935, N369);
or OR3 (N937, N925, N330, N866);
nor NOR2 (N938, N914, N596);
nand NAND3 (N939, N934, N405, N813);
nor NOR4 (N940, N939, N353, N571, N835);
or OR2 (N941, N936, N688);
not NOT1 (N942, N940);
nand NAND3 (N943, N915, N28, N8);
not NOT1 (N944, N937);
buf BUF1 (N945, N938);
nand NAND3 (N946, N931, N318, N72);
xor XOR2 (N947, N943, N20);
or OR2 (N948, N942, N151);
not NOT1 (N949, N921);
nor NOR2 (N950, N949, N469);
nand NAND3 (N951, N932, N511, N841);
nand NAND4 (N952, N946, N60, N59, N7);
xor XOR2 (N953, N950, N759);
buf BUF1 (N954, N952);
buf BUF1 (N955, N951);
xor XOR2 (N956, N953, N528);
not NOT1 (N957, N947);
nand NAND2 (N958, N957, N913);
not NOT1 (N959, N958);
xor XOR2 (N960, N956, N104);
xor XOR2 (N961, N941, N247);
and AND2 (N962, N959, N818);
xor XOR2 (N963, N960, N948);
xor XOR2 (N964, N516, N857);
or OR4 (N965, N954, N584, N419, N182);
xor XOR2 (N966, N944, N270);
nand NAND2 (N967, N919, N657);
xor XOR2 (N968, N961, N957);
or OR3 (N969, N926, N27, N192);
nor NOR3 (N970, N965, N790, N909);
nand NAND3 (N971, N964, N406, N481);
not NOT1 (N972, N971);
nor NOR2 (N973, N945, N898);
or OR3 (N974, N969, N220, N94);
and AND4 (N975, N955, N507, N128, N101);
not NOT1 (N976, N972);
and AND2 (N977, N975, N91);
and AND3 (N978, N977, N970, N412);
not NOT1 (N979, N119);
not NOT1 (N980, N973);
buf BUF1 (N981, N963);
buf BUF1 (N982, N978);
xor XOR2 (N983, N976, N928);
or OR2 (N984, N962, N154);
nand NAND2 (N985, N967, N965);
nor NOR4 (N986, N974, N378, N635, N621);
xor XOR2 (N987, N983, N536);
not NOT1 (N988, N986);
xor XOR2 (N989, N981, N716);
nand NAND4 (N990, N988, N155, N980, N705);
not NOT1 (N991, N89);
nand NAND4 (N992, N979, N145, N810, N646);
or OR4 (N993, N966, N139, N72, N484);
buf BUF1 (N994, N992);
nand NAND3 (N995, N991, N810, N281);
or OR2 (N996, N993, N928);
xor XOR2 (N997, N987, N865);
xor XOR2 (N998, N996, N640);
nor NOR2 (N999, N982, N467);
nand NAND4 (N1000, N985, N512, N765, N902);
and AND3 (N1001, N989, N929, N139);
or OR3 (N1002, N998, N632, N958);
buf BUF1 (N1003, N994);
nand NAND2 (N1004, N1003, N802);
not NOT1 (N1005, N1000);
not NOT1 (N1006, N990);
nand NAND2 (N1007, N1002, N817);
and AND3 (N1008, N995, N522, N726);
or OR3 (N1009, N984, N351, N671);
or OR2 (N1010, N999, N338);
or OR2 (N1011, N1007, N308);
and AND3 (N1012, N1005, N539, N274);
nor NOR4 (N1013, N1011, N554, N393, N51);
buf BUF1 (N1014, N968);
nor NOR3 (N1015, N1010, N892, N923);
or OR2 (N1016, N997, N449);
not NOT1 (N1017, N1008);
and AND3 (N1018, N1017, N812, N192);
or OR3 (N1019, N1016, N336, N154);
buf BUF1 (N1020, N1013);
not NOT1 (N1021, N1014);
nand NAND4 (N1022, N1015, N60, N873, N54);
buf BUF1 (N1023, N1021);
nand NAND4 (N1024, N1018, N1017, N154, N221);
and AND2 (N1025, N1020, N891);
or OR2 (N1026, N1004, N61);
nand NAND3 (N1027, N1009, N902, N1016);
not NOT1 (N1028, N1019);
and AND2 (N1029, N1006, N197);
or OR2 (N1030, N1026, N425);
or OR3 (N1031, N1012, N615, N335);
not NOT1 (N1032, N1027);
and AND3 (N1033, N1022, N456, N238);
or OR3 (N1034, N1031, N419, N899);
or OR2 (N1035, N1023, N761);
xor XOR2 (N1036, N1024, N692);
not NOT1 (N1037, N1025);
or OR3 (N1038, N1029, N865, N817);
nand NAND4 (N1039, N1030, N502, N227, N809);
nor NOR3 (N1040, N1037, N210, N14);
buf BUF1 (N1041, N1035);
or OR2 (N1042, N1039, N805);
nand NAND2 (N1043, N1041, N185);
nor NOR2 (N1044, N1001, N643);
buf BUF1 (N1045, N1033);
xor XOR2 (N1046, N1034, N208);
or OR2 (N1047, N1044, N69);
and AND4 (N1048, N1042, N48, N39, N715);
buf BUF1 (N1049, N1045);
and AND3 (N1050, N1040, N268, N355);
nand NAND3 (N1051, N1047, N520, N28);
not NOT1 (N1052, N1032);
not NOT1 (N1053, N1052);
not NOT1 (N1054, N1038);
and AND4 (N1055, N1036, N1053, N800, N944);
buf BUF1 (N1056, N485);
nand NAND3 (N1057, N1051, N909, N478);
xor XOR2 (N1058, N1050, N231);
nor NOR3 (N1059, N1048, N334, N12);
buf BUF1 (N1060, N1059);
or OR3 (N1061, N1043, N392, N87);
nor NOR3 (N1062, N1056, N350, N1028);
or OR2 (N1063, N677, N1022);
nand NAND2 (N1064, N1063, N1057);
not NOT1 (N1065, N419);
nand NAND4 (N1066, N1060, N900, N46, N466);
buf BUF1 (N1067, N1054);
nor NOR3 (N1068, N1067, N363, N1002);
xor XOR2 (N1069, N1049, N487);
nand NAND3 (N1070, N1061, N360, N813);
nor NOR2 (N1071, N1068, N472);
and AND4 (N1072, N1064, N712, N348, N903);
nand NAND4 (N1073, N1066, N187, N27, N435);
not NOT1 (N1074, N1070);
buf BUF1 (N1075, N1071);
nand NAND4 (N1076, N1058, N555, N645, N594);
nand NAND4 (N1077, N1055, N448, N254, N196);
or OR2 (N1078, N1046, N999);
not NOT1 (N1079, N1065);
and AND2 (N1080, N1072, N983);
nor NOR2 (N1081, N1076, N368);
xor XOR2 (N1082, N1075, N251);
or OR2 (N1083, N1078, N402);
not NOT1 (N1084, N1062);
and AND3 (N1085, N1069, N67, N817);
nor NOR4 (N1086, N1074, N1006, N797, N528);
or OR3 (N1087, N1082, N707, N1);
or OR3 (N1088, N1086, N860, N84);
nand NAND4 (N1089, N1088, N257, N669, N154);
and AND4 (N1090, N1081, N85, N551, N118);
xor XOR2 (N1091, N1085, N231);
xor XOR2 (N1092, N1080, N1077);
or OR3 (N1093, N1035, N150, N723);
xor XOR2 (N1094, N1079, N273);
and AND4 (N1095, N1087, N53, N1053, N658);
or OR3 (N1096, N1090, N409, N744);
nor NOR2 (N1097, N1096, N910);
buf BUF1 (N1098, N1095);
and AND3 (N1099, N1084, N364, N843);
not NOT1 (N1100, N1094);
not NOT1 (N1101, N1098);
not NOT1 (N1102, N1091);
xor XOR2 (N1103, N1097, N18);
and AND2 (N1104, N1100, N337);
xor XOR2 (N1105, N1102, N180);
buf BUF1 (N1106, N1099);
nor NOR2 (N1107, N1101, N939);
nor NOR4 (N1108, N1093, N916, N387, N826);
or OR3 (N1109, N1083, N29, N1105);
not NOT1 (N1110, N549);
buf BUF1 (N1111, N1110);
nor NOR2 (N1112, N1092, N907);
buf BUF1 (N1113, N1104);
buf BUF1 (N1114, N1106);
buf BUF1 (N1115, N1109);
or OR2 (N1116, N1073, N909);
xor XOR2 (N1117, N1107, N1105);
buf BUF1 (N1118, N1108);
and AND3 (N1119, N1111, N688, N508);
not NOT1 (N1120, N1103);
nand NAND4 (N1121, N1119, N1065, N674, N474);
and AND2 (N1122, N1115, N532);
nor NOR2 (N1123, N1089, N830);
or OR4 (N1124, N1117, N867, N1121, N578);
nor NOR4 (N1125, N232, N377, N448, N1088);
nand NAND2 (N1126, N1112, N92);
nor NOR3 (N1127, N1124, N250, N387);
not NOT1 (N1128, N1123);
or OR2 (N1129, N1114, N941);
buf BUF1 (N1130, N1126);
or OR3 (N1131, N1128, N573, N1103);
nand NAND4 (N1132, N1122, N588, N213, N692);
xor XOR2 (N1133, N1118, N417);
not NOT1 (N1134, N1132);
nand NAND2 (N1135, N1116, N537);
and AND2 (N1136, N1134, N40);
xor XOR2 (N1137, N1131, N574);
not NOT1 (N1138, N1130);
or OR3 (N1139, N1136, N531, N1089);
xor XOR2 (N1140, N1127, N827);
nand NAND3 (N1141, N1120, N483, N267);
nor NOR2 (N1142, N1140, N68);
nor NOR4 (N1143, N1135, N378, N181, N320);
buf BUF1 (N1144, N1143);
not NOT1 (N1145, N1125);
or OR3 (N1146, N1138, N841, N25);
not NOT1 (N1147, N1144);
or OR4 (N1148, N1146, N1010, N789, N486);
or OR2 (N1149, N1148, N1085);
nand NAND2 (N1150, N1129, N612);
and AND2 (N1151, N1139, N198);
buf BUF1 (N1152, N1150);
and AND2 (N1153, N1152, N985);
not NOT1 (N1154, N1147);
and AND4 (N1155, N1149, N449, N92, N147);
nor NOR3 (N1156, N1153, N768, N959);
buf BUF1 (N1157, N1154);
buf BUF1 (N1158, N1156);
nor NOR4 (N1159, N1133, N132, N574, N68);
buf BUF1 (N1160, N1158);
xor XOR2 (N1161, N1145, N667);
buf BUF1 (N1162, N1151);
not NOT1 (N1163, N1161);
nor NOR4 (N1164, N1142, N94, N932, N731);
and AND4 (N1165, N1141, N415, N550, N1118);
xor XOR2 (N1166, N1137, N530);
xor XOR2 (N1167, N1162, N405);
xor XOR2 (N1168, N1155, N34);
not NOT1 (N1169, N1159);
or OR4 (N1170, N1163, N880, N126, N172);
and AND2 (N1171, N1168, N759);
nand NAND2 (N1172, N1169, N530);
buf BUF1 (N1173, N1171);
nor NOR4 (N1174, N1173, N420, N79, N632);
xor XOR2 (N1175, N1170, N616);
nand NAND2 (N1176, N1167, N865);
nor NOR4 (N1177, N1160, N939, N65, N1078);
nor NOR4 (N1178, N1176, N306, N439, N111);
nor NOR3 (N1179, N1172, N778, N820);
xor XOR2 (N1180, N1165, N1137);
or OR3 (N1181, N1157, N395, N1090);
and AND3 (N1182, N1164, N1133, N244);
or OR4 (N1183, N1174, N865, N773, N1078);
nor NOR2 (N1184, N1175, N55);
not NOT1 (N1185, N1178);
nor NOR4 (N1186, N1181, N896, N124, N345);
not NOT1 (N1187, N1183);
nor NOR3 (N1188, N1180, N676, N150);
or OR4 (N1189, N1187, N165, N340, N857);
not NOT1 (N1190, N1166);
or OR3 (N1191, N1186, N108, N653);
or OR2 (N1192, N1113, N189);
buf BUF1 (N1193, N1188);
or OR4 (N1194, N1185, N153, N1017, N328);
not NOT1 (N1195, N1192);
or OR4 (N1196, N1189, N1038, N745, N1016);
and AND3 (N1197, N1195, N1017, N1088);
not NOT1 (N1198, N1191);
buf BUF1 (N1199, N1182);
nor NOR4 (N1200, N1196, N1192, N847, N59);
xor XOR2 (N1201, N1200, N892);
not NOT1 (N1202, N1197);
and AND2 (N1203, N1193, N405);
nand NAND3 (N1204, N1198, N1177, N639);
and AND3 (N1205, N99, N877, N988);
xor XOR2 (N1206, N1204, N181);
buf BUF1 (N1207, N1205);
and AND3 (N1208, N1203, N763, N548);
nand NAND3 (N1209, N1179, N1000, N654);
nand NAND4 (N1210, N1209, N137, N172, N840);
and AND4 (N1211, N1207, N1210, N980, N554);
nand NAND4 (N1212, N1081, N6, N1063, N96);
nand NAND2 (N1213, N1208, N670);
and AND3 (N1214, N1184, N822, N79);
xor XOR2 (N1215, N1212, N1057);
nand NAND3 (N1216, N1213, N746, N615);
and AND2 (N1217, N1214, N174);
nand NAND2 (N1218, N1199, N1072);
nor NOR2 (N1219, N1202, N391);
buf BUF1 (N1220, N1194);
nor NOR4 (N1221, N1201, N1064, N1026, N980);
nor NOR2 (N1222, N1217, N60);
buf BUF1 (N1223, N1222);
buf BUF1 (N1224, N1211);
nand NAND2 (N1225, N1223, N231);
nor NOR3 (N1226, N1206, N558, N862);
nor NOR4 (N1227, N1220, N132, N419, N243);
not NOT1 (N1228, N1224);
and AND4 (N1229, N1227, N971, N343, N855);
not NOT1 (N1230, N1228);
and AND2 (N1231, N1225, N1016);
or OR2 (N1232, N1190, N717);
and AND3 (N1233, N1218, N305, N947);
buf BUF1 (N1234, N1229);
xor XOR2 (N1235, N1219, N200);
nor NOR3 (N1236, N1233, N1093, N522);
buf BUF1 (N1237, N1236);
xor XOR2 (N1238, N1234, N646);
and AND3 (N1239, N1237, N226, N129);
nor NOR3 (N1240, N1235, N1137, N605);
xor XOR2 (N1241, N1221, N332);
buf BUF1 (N1242, N1230);
not NOT1 (N1243, N1241);
and AND4 (N1244, N1238, N976, N1144, N449);
buf BUF1 (N1245, N1240);
or OR3 (N1246, N1231, N578, N973);
and AND3 (N1247, N1242, N671, N754);
or OR4 (N1248, N1244, N518, N323, N856);
xor XOR2 (N1249, N1247, N311);
buf BUF1 (N1250, N1246);
or OR2 (N1251, N1249, N681);
not NOT1 (N1252, N1226);
nor NOR4 (N1253, N1243, N688, N9, N1090);
and AND4 (N1254, N1215, N848, N18, N588);
or OR4 (N1255, N1232, N391, N227, N456);
buf BUF1 (N1256, N1255);
nand NAND3 (N1257, N1239, N278, N447);
xor XOR2 (N1258, N1256, N412);
nand NAND4 (N1259, N1216, N581, N1207, N239);
buf BUF1 (N1260, N1257);
xor XOR2 (N1261, N1252, N299);
nand NAND2 (N1262, N1245, N1088);
not NOT1 (N1263, N1251);
buf BUF1 (N1264, N1250);
buf BUF1 (N1265, N1254);
xor XOR2 (N1266, N1261, N83);
xor XOR2 (N1267, N1263, N574);
and AND3 (N1268, N1266, N296, N493);
nand NAND2 (N1269, N1264, N1183);
and AND3 (N1270, N1258, N718, N550);
and AND4 (N1271, N1267, N1085, N168, N105);
xor XOR2 (N1272, N1269, N378);
nor NOR4 (N1273, N1268, N744, N1264, N462);
and AND3 (N1274, N1270, N637, N751);
or OR2 (N1275, N1253, N338);
xor XOR2 (N1276, N1265, N155);
buf BUF1 (N1277, N1259);
nor NOR3 (N1278, N1262, N421, N700);
or OR4 (N1279, N1260, N1071, N616, N798);
nand NAND4 (N1280, N1276, N250, N1246, N281);
nor NOR3 (N1281, N1278, N654, N1235);
or OR2 (N1282, N1275, N899);
and AND2 (N1283, N1277, N235);
or OR3 (N1284, N1281, N995, N1074);
and AND2 (N1285, N1279, N1080);
and AND4 (N1286, N1271, N477, N19, N852);
not NOT1 (N1287, N1272);
nor NOR3 (N1288, N1280, N1204, N149);
nor NOR3 (N1289, N1288, N83, N1183);
nor NOR2 (N1290, N1284, N789);
nand NAND2 (N1291, N1290, N1213);
or OR3 (N1292, N1283, N23, N865);
nand NAND2 (N1293, N1285, N469);
and AND3 (N1294, N1291, N923, N786);
nand NAND4 (N1295, N1289, N841, N176, N720);
or OR4 (N1296, N1293, N151, N958, N670);
nor NOR2 (N1297, N1248, N1250);
nor NOR2 (N1298, N1292, N748);
nor NOR2 (N1299, N1296, N406);
buf BUF1 (N1300, N1295);
nand NAND2 (N1301, N1300, N661);
not NOT1 (N1302, N1294);
not NOT1 (N1303, N1282);
or OR3 (N1304, N1299, N1186, N828);
or OR4 (N1305, N1286, N993, N1033, N970);
or OR4 (N1306, N1274, N850, N987, N350);
buf BUF1 (N1307, N1273);
nor NOR4 (N1308, N1303, N883, N589, N344);
xor XOR2 (N1309, N1304, N242);
buf BUF1 (N1310, N1302);
or OR4 (N1311, N1310, N431, N792, N313);
nand NAND4 (N1312, N1306, N433, N875, N441);
and AND2 (N1313, N1301, N960);
xor XOR2 (N1314, N1312, N1112);
xor XOR2 (N1315, N1297, N57);
not NOT1 (N1316, N1287);
nand NAND3 (N1317, N1309, N119, N685);
or OR2 (N1318, N1308, N1260);
not NOT1 (N1319, N1307);
or OR3 (N1320, N1318, N994, N216);
or OR4 (N1321, N1316, N1141, N286, N100);
or OR4 (N1322, N1311, N789, N550, N345);
and AND3 (N1323, N1317, N498, N272);
nand NAND3 (N1324, N1313, N6, N654);
not NOT1 (N1325, N1319);
nor NOR3 (N1326, N1305, N1275, N892);
buf BUF1 (N1327, N1324);
nand NAND4 (N1328, N1315, N1159, N819, N96);
nor NOR4 (N1329, N1314, N387, N176, N941);
or OR4 (N1330, N1298, N112, N171, N220);
buf BUF1 (N1331, N1322);
or OR2 (N1332, N1325, N173);
xor XOR2 (N1333, N1321, N161);
not NOT1 (N1334, N1332);
nor NOR4 (N1335, N1328, N984, N437, N1231);
or OR2 (N1336, N1320, N640);
nor NOR2 (N1337, N1331, N893);
or OR3 (N1338, N1327, N640, N1307);
or OR4 (N1339, N1326, N468, N353, N625);
nor NOR3 (N1340, N1335, N49, N870);
buf BUF1 (N1341, N1340);
and AND4 (N1342, N1330, N1097, N1274, N718);
xor XOR2 (N1343, N1329, N15);
and AND3 (N1344, N1342, N1026, N1264);
nand NAND3 (N1345, N1344, N968, N1247);
not NOT1 (N1346, N1336);
nand NAND4 (N1347, N1333, N818, N1079, N600);
buf BUF1 (N1348, N1343);
not NOT1 (N1349, N1341);
and AND2 (N1350, N1337, N1104);
nor NOR4 (N1351, N1347, N321, N1247, N244);
buf BUF1 (N1352, N1346);
and AND3 (N1353, N1323, N49, N1285);
or OR2 (N1354, N1349, N1196);
not NOT1 (N1355, N1345);
and AND2 (N1356, N1348, N1267);
nor NOR2 (N1357, N1353, N1143);
not NOT1 (N1358, N1355);
xor XOR2 (N1359, N1334, N471);
buf BUF1 (N1360, N1350);
xor XOR2 (N1361, N1339, N733);
not NOT1 (N1362, N1361);
or OR4 (N1363, N1356, N808, N970, N11);
and AND3 (N1364, N1357, N989, N408);
or OR4 (N1365, N1358, N111, N417, N423);
and AND2 (N1366, N1351, N687);
buf BUF1 (N1367, N1364);
or OR2 (N1368, N1366, N724);
nand NAND2 (N1369, N1352, N743);
xor XOR2 (N1370, N1368, N1355);
nand NAND3 (N1371, N1338, N359, N543);
xor XOR2 (N1372, N1362, N90);
nor NOR2 (N1373, N1359, N35);
buf BUF1 (N1374, N1363);
not NOT1 (N1375, N1374);
nand NAND2 (N1376, N1369, N18);
nor NOR4 (N1377, N1360, N719, N895, N1021);
not NOT1 (N1378, N1354);
buf BUF1 (N1379, N1372);
xor XOR2 (N1380, N1379, N63);
or OR2 (N1381, N1373, N1145);
or OR4 (N1382, N1378, N660, N365, N1054);
buf BUF1 (N1383, N1365);
or OR3 (N1384, N1377, N130, N901);
and AND4 (N1385, N1383, N983, N1166, N470);
xor XOR2 (N1386, N1367, N1087);
buf BUF1 (N1387, N1376);
xor XOR2 (N1388, N1381, N199);
not NOT1 (N1389, N1388);
nor NOR3 (N1390, N1385, N594, N499);
buf BUF1 (N1391, N1370);
buf BUF1 (N1392, N1387);
nor NOR3 (N1393, N1371, N1164, N1230);
buf BUF1 (N1394, N1380);
nor NOR4 (N1395, N1392, N147, N1042, N594);
nor NOR2 (N1396, N1390, N804);
not NOT1 (N1397, N1384);
nor NOR4 (N1398, N1375, N1179, N363, N182);
xor XOR2 (N1399, N1391, N264);
not NOT1 (N1400, N1393);
nor NOR3 (N1401, N1395, N1109, N157);
or OR2 (N1402, N1389, N685);
and AND2 (N1403, N1386, N884);
nand NAND2 (N1404, N1401, N936);
or OR2 (N1405, N1394, N473);
xor XOR2 (N1406, N1397, N212);
xor XOR2 (N1407, N1399, N879);
not NOT1 (N1408, N1382);
and AND3 (N1409, N1403, N918, N419);
xor XOR2 (N1410, N1396, N115);
nand NAND4 (N1411, N1404, N400, N116, N529);
not NOT1 (N1412, N1408);
buf BUF1 (N1413, N1406);
buf BUF1 (N1414, N1410);
buf BUF1 (N1415, N1402);
nand NAND2 (N1416, N1415, N1292);
and AND4 (N1417, N1405, N757, N808, N968);
not NOT1 (N1418, N1409);
nor NOR2 (N1419, N1411, N322);
xor XOR2 (N1420, N1419, N1395);
not NOT1 (N1421, N1412);
nand NAND3 (N1422, N1418, N370, N487);
or OR4 (N1423, N1407, N380, N891, N1012);
xor XOR2 (N1424, N1420, N651);
buf BUF1 (N1425, N1414);
buf BUF1 (N1426, N1417);
nor NOR2 (N1427, N1416, N109);
xor XOR2 (N1428, N1427, N246);
xor XOR2 (N1429, N1428, N547);
and AND4 (N1430, N1423, N99, N414, N827);
or OR2 (N1431, N1413, N793);
xor XOR2 (N1432, N1431, N779);
and AND4 (N1433, N1422, N589, N17, N734);
nand NAND4 (N1434, N1400, N545, N1251, N1311);
and AND3 (N1435, N1424, N487, N259);
or OR3 (N1436, N1430, N313, N13);
and AND3 (N1437, N1421, N1104, N1161);
nand NAND2 (N1438, N1398, N589);
xor XOR2 (N1439, N1425, N875);
not NOT1 (N1440, N1438);
and AND4 (N1441, N1434, N1411, N1181, N1173);
or OR2 (N1442, N1436, N1340);
and AND3 (N1443, N1441, N418, N290);
or OR3 (N1444, N1435, N1010, N649);
nor NOR3 (N1445, N1440, N1094, N1271);
not NOT1 (N1446, N1432);
nand NAND2 (N1447, N1433, N850);
buf BUF1 (N1448, N1442);
nand NAND2 (N1449, N1448, N908);
nor NOR3 (N1450, N1437, N1237, N582);
buf BUF1 (N1451, N1450);
not NOT1 (N1452, N1447);
nor NOR4 (N1453, N1444, N1124, N1406, N670);
and AND3 (N1454, N1443, N554, N1289);
buf BUF1 (N1455, N1426);
nor NOR3 (N1456, N1455, N1104, N207);
xor XOR2 (N1457, N1439, N503);
not NOT1 (N1458, N1449);
xor XOR2 (N1459, N1429, N1028);
and AND3 (N1460, N1454, N1250, N241);
buf BUF1 (N1461, N1446);
xor XOR2 (N1462, N1458, N192);
nor NOR2 (N1463, N1445, N565);
or OR3 (N1464, N1456, N1173, N318);
or OR4 (N1465, N1453, N830, N84, N1250);
xor XOR2 (N1466, N1457, N277);
buf BUF1 (N1467, N1464);
buf BUF1 (N1468, N1461);
nand NAND4 (N1469, N1451, N1305, N1148, N977);
xor XOR2 (N1470, N1460, N803);
nand NAND4 (N1471, N1463, N1193, N1433, N22);
buf BUF1 (N1472, N1468);
or OR2 (N1473, N1471, N675);
xor XOR2 (N1474, N1467, N1361);
and AND3 (N1475, N1473, N137, N1054);
or OR2 (N1476, N1472, N586);
nor NOR2 (N1477, N1475, N215);
buf BUF1 (N1478, N1465);
xor XOR2 (N1479, N1469, N1183);
not NOT1 (N1480, N1477);
nand NAND2 (N1481, N1478, N1300);
nand NAND2 (N1482, N1470, N1351);
nand NAND2 (N1483, N1459, N734);
nor NOR3 (N1484, N1462, N1313, N447);
not NOT1 (N1485, N1480);
xor XOR2 (N1486, N1483, N663);
or OR2 (N1487, N1479, N1211);
and AND4 (N1488, N1474, N1013, N1107, N1387);
or OR2 (N1489, N1481, N1148);
or OR3 (N1490, N1485, N196, N722);
buf BUF1 (N1491, N1484);
or OR2 (N1492, N1466, N174);
and AND2 (N1493, N1492, N427);
nor NOR3 (N1494, N1490, N486, N968);
nor NOR2 (N1495, N1482, N16);
nand NAND2 (N1496, N1489, N1130);
not NOT1 (N1497, N1496);
xor XOR2 (N1498, N1495, N733);
xor XOR2 (N1499, N1491, N814);
and AND2 (N1500, N1493, N830);
nor NOR4 (N1501, N1498, N668, N257, N403);
nor NOR3 (N1502, N1499, N931, N1232);
and AND4 (N1503, N1488, N242, N921, N79);
nor NOR2 (N1504, N1494, N397);
xor XOR2 (N1505, N1502, N693);
or OR3 (N1506, N1504, N815, N1267);
nand NAND2 (N1507, N1503, N216);
xor XOR2 (N1508, N1486, N660);
nand NAND3 (N1509, N1501, N1029, N1202);
nand NAND2 (N1510, N1452, N192);
nand NAND3 (N1511, N1509, N921, N1079);
xor XOR2 (N1512, N1505, N1000);
or OR2 (N1513, N1512, N136);
and AND2 (N1514, N1476, N248);
or OR2 (N1515, N1510, N609);
buf BUF1 (N1516, N1507);
buf BUF1 (N1517, N1515);
nand NAND4 (N1518, N1497, N1028, N1151, N1309);
nor NOR2 (N1519, N1518, N751);
not NOT1 (N1520, N1514);
nor NOR4 (N1521, N1520, N1216, N992, N562);
buf BUF1 (N1522, N1500);
not NOT1 (N1523, N1521);
nand NAND3 (N1524, N1513, N1305, N938);
xor XOR2 (N1525, N1508, N1215);
nand NAND4 (N1526, N1523, N1101, N633, N563);
nor NOR3 (N1527, N1522, N1134, N326);
nand NAND4 (N1528, N1527, N1205, N1083, N1130);
or OR2 (N1529, N1525, N1151);
nor NOR2 (N1530, N1526, N1321);
buf BUF1 (N1531, N1506);
not NOT1 (N1532, N1528);
not NOT1 (N1533, N1524);
nor NOR3 (N1534, N1516, N620, N359);
buf BUF1 (N1535, N1531);
nor NOR4 (N1536, N1535, N724, N732, N1205);
and AND2 (N1537, N1532, N193);
or OR4 (N1538, N1487, N812, N660, N559);
nand NAND2 (N1539, N1519, N617);
buf BUF1 (N1540, N1536);
not NOT1 (N1541, N1511);
not NOT1 (N1542, N1537);
xor XOR2 (N1543, N1529, N221);
not NOT1 (N1544, N1540);
not NOT1 (N1545, N1541);
not NOT1 (N1546, N1517);
buf BUF1 (N1547, N1546);
buf BUF1 (N1548, N1544);
xor XOR2 (N1549, N1542, N1010);
buf BUF1 (N1550, N1533);
nor NOR4 (N1551, N1539, N1208, N318, N1385);
nand NAND3 (N1552, N1530, N201, N1527);
buf BUF1 (N1553, N1551);
nor NOR2 (N1554, N1549, N608);
nor NOR3 (N1555, N1553, N108, N740);
buf BUF1 (N1556, N1545);
nand NAND4 (N1557, N1548, N337, N532, N355);
xor XOR2 (N1558, N1547, N859);
xor XOR2 (N1559, N1556, N1390);
nor NOR4 (N1560, N1555, N443, N325, N493);
nor NOR4 (N1561, N1559, N1527, N180, N1261);
buf BUF1 (N1562, N1538);
nor NOR2 (N1563, N1550, N208);
nor NOR2 (N1564, N1561, N929);
nand NAND2 (N1565, N1560, N212);
or OR4 (N1566, N1552, N1300, N596, N1065);
nor NOR2 (N1567, N1564, N1331);
nor NOR2 (N1568, N1534, N736);
nor NOR3 (N1569, N1563, N13, N893);
nand NAND3 (N1570, N1557, N832, N520);
not NOT1 (N1571, N1562);
xor XOR2 (N1572, N1571, N158);
buf BUF1 (N1573, N1566);
nand NAND3 (N1574, N1565, N179, N311);
nor NOR4 (N1575, N1568, N1107, N1275, N958);
nand NAND4 (N1576, N1567, N145, N621, N1539);
nand NAND2 (N1577, N1569, N291);
buf BUF1 (N1578, N1543);
xor XOR2 (N1579, N1578, N6);
not NOT1 (N1580, N1579);
or OR2 (N1581, N1570, N1453);
and AND2 (N1582, N1577, N212);
nand NAND3 (N1583, N1558, N945, N843);
xor XOR2 (N1584, N1576, N1452);
and AND3 (N1585, N1575, N1120, N519);
not NOT1 (N1586, N1554);
xor XOR2 (N1587, N1574, N755);
not NOT1 (N1588, N1587);
nand NAND4 (N1589, N1585, N1018, N831, N755);
or OR4 (N1590, N1580, N1068, N1529, N1194);
nand NAND2 (N1591, N1572, N668);
and AND3 (N1592, N1573, N170, N795);
buf BUF1 (N1593, N1581);
buf BUF1 (N1594, N1591);
and AND3 (N1595, N1588, N1543, N1431);
nand NAND2 (N1596, N1583, N153);
or OR2 (N1597, N1582, N241);
not NOT1 (N1598, N1586);
nand NAND2 (N1599, N1589, N1275);
or OR4 (N1600, N1597, N1068, N1388, N228);
buf BUF1 (N1601, N1599);
nor NOR4 (N1602, N1598, N219, N994, N1181);
and AND4 (N1603, N1584, N585, N741, N542);
not NOT1 (N1604, N1601);
and AND4 (N1605, N1594, N518, N285, N866);
buf BUF1 (N1606, N1603);
and AND2 (N1607, N1595, N919);
nand NAND2 (N1608, N1600, N1463);
buf BUF1 (N1609, N1604);
nor NOR2 (N1610, N1590, N60);
nor NOR2 (N1611, N1592, N321);
not NOT1 (N1612, N1593);
xor XOR2 (N1613, N1610, N656);
not NOT1 (N1614, N1609);
buf BUF1 (N1615, N1607);
and AND3 (N1616, N1614, N442, N149);
and AND2 (N1617, N1611, N534);
and AND3 (N1618, N1606, N1398, N94);
and AND4 (N1619, N1596, N936, N1537, N383);
nand NAND4 (N1620, N1605, N1453, N63, N790);
xor XOR2 (N1621, N1608, N1008);
not NOT1 (N1622, N1616);
not NOT1 (N1623, N1618);
not NOT1 (N1624, N1621);
not NOT1 (N1625, N1617);
nor NOR4 (N1626, N1625, N1622, N960, N1104);
buf BUF1 (N1627, N632);
not NOT1 (N1628, N1626);
nor NOR3 (N1629, N1615, N718, N1203);
not NOT1 (N1630, N1627);
not NOT1 (N1631, N1612);
xor XOR2 (N1632, N1620, N596);
buf BUF1 (N1633, N1632);
nand NAND4 (N1634, N1623, N549, N93, N949);
buf BUF1 (N1635, N1633);
not NOT1 (N1636, N1628);
and AND2 (N1637, N1630, N866);
xor XOR2 (N1638, N1637, N935);
xor XOR2 (N1639, N1631, N874);
nand NAND2 (N1640, N1619, N1446);
or OR2 (N1641, N1636, N529);
xor XOR2 (N1642, N1634, N1087);
xor XOR2 (N1643, N1613, N1240);
and AND4 (N1644, N1638, N712, N668, N739);
not NOT1 (N1645, N1641);
buf BUF1 (N1646, N1643);
or OR3 (N1647, N1644, N1600, N255);
not NOT1 (N1648, N1642);
buf BUF1 (N1649, N1640);
nor NOR2 (N1650, N1602, N83);
buf BUF1 (N1651, N1629);
nor NOR2 (N1652, N1648, N32);
buf BUF1 (N1653, N1635);
nand NAND4 (N1654, N1646, N585, N276, N409);
nand NAND3 (N1655, N1651, N1568, N23);
and AND2 (N1656, N1645, N206);
and AND2 (N1657, N1649, N1595);
xor XOR2 (N1658, N1657, N358);
and AND2 (N1659, N1624, N1322);
or OR2 (N1660, N1658, N258);
buf BUF1 (N1661, N1660);
not NOT1 (N1662, N1652);
or OR3 (N1663, N1655, N45, N813);
nor NOR3 (N1664, N1659, N955, N1373);
buf BUF1 (N1665, N1639);
nand NAND2 (N1666, N1664, N1440);
not NOT1 (N1667, N1663);
or OR2 (N1668, N1661, N135);
nor NOR4 (N1669, N1647, N1220, N1064, N1403);
and AND4 (N1670, N1668, N565, N568, N359);
nor NOR2 (N1671, N1654, N435);
or OR3 (N1672, N1653, N977, N157);
xor XOR2 (N1673, N1669, N161);
or OR4 (N1674, N1671, N1279, N1539, N190);
not NOT1 (N1675, N1670);
nand NAND2 (N1676, N1656, N1402);
not NOT1 (N1677, N1666);
or OR2 (N1678, N1672, N814);
buf BUF1 (N1679, N1674);
nand NAND4 (N1680, N1676, N1270, N895, N133);
or OR4 (N1681, N1680, N1025, N76, N1029);
and AND3 (N1682, N1650, N714, N1339);
buf BUF1 (N1683, N1682);
buf BUF1 (N1684, N1683);
xor XOR2 (N1685, N1678, N910);
or OR2 (N1686, N1685, N1072);
and AND4 (N1687, N1667, N1014, N287, N1663);
buf BUF1 (N1688, N1665);
xor XOR2 (N1689, N1662, N1168);
and AND2 (N1690, N1686, N1026);
nor NOR3 (N1691, N1673, N612, N509);
xor XOR2 (N1692, N1687, N21);
nor NOR2 (N1693, N1681, N287);
nand NAND2 (N1694, N1684, N93);
nand NAND4 (N1695, N1691, N1186, N566, N1034);
nand NAND4 (N1696, N1688, N341, N137, N1027);
or OR4 (N1697, N1692, N1343, N476, N1609);
or OR3 (N1698, N1679, N1243, N1378);
buf BUF1 (N1699, N1697);
xor XOR2 (N1700, N1677, N463);
or OR3 (N1701, N1690, N488, N809);
nand NAND2 (N1702, N1700, N411);
not NOT1 (N1703, N1699);
buf BUF1 (N1704, N1702);
buf BUF1 (N1705, N1695);
nor NOR4 (N1706, N1694, N1262, N746, N259);
buf BUF1 (N1707, N1675);
nand NAND4 (N1708, N1698, N997, N1649, N1207);
not NOT1 (N1709, N1689);
xor XOR2 (N1710, N1693, N189);
or OR4 (N1711, N1701, N423, N921, N142);
or OR4 (N1712, N1705, N1211, N950, N1589);
nor NOR4 (N1713, N1703, N581, N643, N1519);
nor NOR4 (N1714, N1710, N736, N1131, N1317);
xor XOR2 (N1715, N1712, N1661);
xor XOR2 (N1716, N1696, N1300);
buf BUF1 (N1717, N1714);
nor NOR3 (N1718, N1708, N64, N211);
or OR4 (N1719, N1704, N582, N1537, N1701);
not NOT1 (N1720, N1717);
buf BUF1 (N1721, N1711);
not NOT1 (N1722, N1709);
nor NOR4 (N1723, N1706, N1593, N1301, N746);
xor XOR2 (N1724, N1723, N909);
buf BUF1 (N1725, N1713);
buf BUF1 (N1726, N1722);
or OR2 (N1727, N1707, N1148);
not NOT1 (N1728, N1718);
or OR4 (N1729, N1725, N898, N1177, N396);
or OR3 (N1730, N1719, N412, N1633);
and AND2 (N1731, N1730, N36);
nor NOR3 (N1732, N1726, N889, N1107);
nor NOR3 (N1733, N1732, N799, N1253);
nand NAND4 (N1734, N1716, N838, N1609, N550);
not NOT1 (N1735, N1715);
buf BUF1 (N1736, N1720);
or OR3 (N1737, N1733, N556, N1461);
xor XOR2 (N1738, N1735, N1086);
and AND3 (N1739, N1724, N1371, N1491);
and AND2 (N1740, N1729, N1456);
xor XOR2 (N1741, N1737, N338);
and AND3 (N1742, N1728, N1436, N956);
and AND3 (N1743, N1727, N1692, N1554);
or OR4 (N1744, N1736, N1443, N35, N1034);
or OR2 (N1745, N1741, N903);
nand NAND4 (N1746, N1742, N332, N878, N728);
and AND2 (N1747, N1743, N59);
nor NOR4 (N1748, N1747, N58, N9, N876);
nor NOR3 (N1749, N1734, N735, N61);
buf BUF1 (N1750, N1738);
not NOT1 (N1751, N1750);
xor XOR2 (N1752, N1740, N1006);
nand NAND3 (N1753, N1749, N312, N846);
not NOT1 (N1754, N1721);
xor XOR2 (N1755, N1751, N26);
xor XOR2 (N1756, N1739, N516);
or OR2 (N1757, N1753, N707);
nand NAND4 (N1758, N1754, N1075, N1354, N1392);
not NOT1 (N1759, N1744);
nor NOR2 (N1760, N1731, N1497);
buf BUF1 (N1761, N1752);
buf BUF1 (N1762, N1757);
nand NAND3 (N1763, N1759, N759, N1034);
buf BUF1 (N1764, N1762);
and AND2 (N1765, N1760, N12);
or OR3 (N1766, N1761, N1471, N798);
not NOT1 (N1767, N1745);
not NOT1 (N1768, N1748);
xor XOR2 (N1769, N1767, N1338);
or OR4 (N1770, N1766, N1342, N295, N1059);
nand NAND3 (N1771, N1769, N1522, N532);
not NOT1 (N1772, N1758);
buf BUF1 (N1773, N1772);
nor NOR4 (N1774, N1764, N492, N469, N861);
not NOT1 (N1775, N1756);
nor NOR2 (N1776, N1770, N1228);
nor NOR2 (N1777, N1763, N741);
buf BUF1 (N1778, N1774);
and AND4 (N1779, N1775, N1522, N1265, N96);
nor NOR4 (N1780, N1755, N1573, N117, N778);
xor XOR2 (N1781, N1746, N611);
nand NAND3 (N1782, N1776, N999, N1297);
xor XOR2 (N1783, N1765, N264);
buf BUF1 (N1784, N1782);
or OR3 (N1785, N1773, N1634, N349);
not NOT1 (N1786, N1785);
and AND2 (N1787, N1784, N994);
xor XOR2 (N1788, N1781, N1374);
and AND2 (N1789, N1777, N235);
buf BUF1 (N1790, N1783);
buf BUF1 (N1791, N1789);
and AND4 (N1792, N1787, N333, N684, N1453);
and AND4 (N1793, N1790, N1700, N629, N1753);
or OR4 (N1794, N1768, N770, N1592, N1623);
or OR2 (N1795, N1793, N233);
or OR3 (N1796, N1794, N1049, N133);
nor NOR4 (N1797, N1778, N1567, N1395, N860);
or OR4 (N1798, N1791, N1730, N704, N1735);
and AND3 (N1799, N1795, N1422, N441);
buf BUF1 (N1800, N1771);
and AND4 (N1801, N1779, N815, N1259, N1096);
or OR4 (N1802, N1799, N55, N410, N1127);
buf BUF1 (N1803, N1802);
xor XOR2 (N1804, N1786, N146);
nor NOR2 (N1805, N1804, N813);
or OR2 (N1806, N1798, N1746);
or OR2 (N1807, N1780, N1148);
and AND2 (N1808, N1796, N584);
or OR2 (N1809, N1801, N328);
buf BUF1 (N1810, N1797);
not NOT1 (N1811, N1805);
nor NOR2 (N1812, N1810, N1114);
nor NOR2 (N1813, N1788, N1080);
and AND3 (N1814, N1812, N1664, N1663);
nand NAND4 (N1815, N1809, N42, N1807, N961);
buf BUF1 (N1816, N1321);
buf BUF1 (N1817, N1814);
and AND2 (N1818, N1815, N882);
buf BUF1 (N1819, N1816);
xor XOR2 (N1820, N1808, N1190);
buf BUF1 (N1821, N1818);
nor NOR3 (N1822, N1806, N618, N79);
not NOT1 (N1823, N1811);
nor NOR3 (N1824, N1820, N439, N1766);
nor NOR3 (N1825, N1800, N159, N875);
or OR4 (N1826, N1825, N1014, N914, N1390);
or OR2 (N1827, N1826, N49);
nor NOR4 (N1828, N1792, N1105, N1176, N1180);
or OR2 (N1829, N1817, N1014);
not NOT1 (N1830, N1823);
and AND3 (N1831, N1822, N1726, N1387);
nand NAND3 (N1832, N1831, N69, N563);
or OR3 (N1833, N1819, N631, N1661);
and AND2 (N1834, N1803, N1786);
nor NOR2 (N1835, N1828, N172);
or OR4 (N1836, N1821, N1533, N34, N895);
nand NAND4 (N1837, N1836, N854, N1295, N523);
buf BUF1 (N1838, N1813);
or OR3 (N1839, N1837, N1540, N554);
buf BUF1 (N1840, N1839);
not NOT1 (N1841, N1824);
nand NAND3 (N1842, N1827, N493, N872);
not NOT1 (N1843, N1841);
xor XOR2 (N1844, N1829, N1445);
nor NOR2 (N1845, N1834, N1725);
nand NAND2 (N1846, N1835, N1830);
not NOT1 (N1847, N561);
xor XOR2 (N1848, N1840, N367);
and AND3 (N1849, N1848, N1214, N130);
buf BUF1 (N1850, N1844);
and AND2 (N1851, N1838, N1459);
nor NOR4 (N1852, N1842, N1847, N1112, N921);
nor NOR4 (N1853, N1627, N18, N93, N428);
not NOT1 (N1854, N1850);
or OR3 (N1855, N1843, N1283, N1607);
xor XOR2 (N1856, N1849, N1807);
nor NOR2 (N1857, N1845, N1175);
not NOT1 (N1858, N1853);
buf BUF1 (N1859, N1846);
xor XOR2 (N1860, N1856, N1489);
xor XOR2 (N1861, N1832, N630);
nor NOR2 (N1862, N1859, N1368);
nand NAND4 (N1863, N1854, N1751, N634, N1801);
xor XOR2 (N1864, N1855, N840);
or OR2 (N1865, N1861, N1767);
or OR2 (N1866, N1852, N1477);
buf BUF1 (N1867, N1858);
xor XOR2 (N1868, N1866, N684);
nand NAND2 (N1869, N1860, N1145);
or OR3 (N1870, N1868, N1076, N1650);
and AND4 (N1871, N1867, N62, N166, N1547);
or OR3 (N1872, N1864, N1808, N1616);
nand NAND4 (N1873, N1872, N1641, N401, N721);
nand NAND2 (N1874, N1857, N1176);
xor XOR2 (N1875, N1863, N1189);
not NOT1 (N1876, N1873);
not NOT1 (N1877, N1862);
nand NAND4 (N1878, N1871, N1645, N1170, N677);
buf BUF1 (N1879, N1870);
xor XOR2 (N1880, N1875, N1594);
nand NAND4 (N1881, N1833, N935, N553, N1064);
xor XOR2 (N1882, N1876, N908);
buf BUF1 (N1883, N1881);
not NOT1 (N1884, N1879);
buf BUF1 (N1885, N1869);
nor NOR2 (N1886, N1880, N1863);
buf BUF1 (N1887, N1878);
and AND4 (N1888, N1883, N1146, N293, N465);
buf BUF1 (N1889, N1886);
or OR3 (N1890, N1889, N445, N675);
not NOT1 (N1891, N1888);
buf BUF1 (N1892, N1851);
buf BUF1 (N1893, N1882);
nor NOR4 (N1894, N1893, N1693, N83, N176);
nand NAND4 (N1895, N1887, N108, N558, N1179);
nor NOR4 (N1896, N1894, N320, N1160, N986);
xor XOR2 (N1897, N1865, N524);
not NOT1 (N1898, N1897);
xor XOR2 (N1899, N1884, N209);
not NOT1 (N1900, N1874);
and AND3 (N1901, N1895, N1613, N372);
nand NAND4 (N1902, N1877, N32, N1371, N829);
nand NAND2 (N1903, N1902, N1868);
not NOT1 (N1904, N1901);
not NOT1 (N1905, N1904);
nor NOR2 (N1906, N1892, N889);
and AND2 (N1907, N1890, N372);
not NOT1 (N1908, N1907);
not NOT1 (N1909, N1898);
buf BUF1 (N1910, N1903);
nor NOR4 (N1911, N1896, N1008, N450, N1243);
and AND3 (N1912, N1910, N901, N1096);
or OR3 (N1913, N1906, N1498, N1358);
or OR3 (N1914, N1900, N866, N640);
xor XOR2 (N1915, N1913, N1193);
xor XOR2 (N1916, N1914, N558);
and AND2 (N1917, N1915, N1347);
buf BUF1 (N1918, N1908);
and AND4 (N1919, N1885, N1318, N454, N1552);
or OR3 (N1920, N1919, N1444, N1218);
nor NOR3 (N1921, N1899, N276, N1161);
xor XOR2 (N1922, N1911, N1464);
nor NOR2 (N1923, N1891, N888);
and AND3 (N1924, N1905, N595, N1526);
buf BUF1 (N1925, N1917);
and AND3 (N1926, N1923, N138, N660);
nor NOR2 (N1927, N1921, N830);
nor NOR3 (N1928, N1925, N589, N1875);
or OR3 (N1929, N1927, N747, N286);
or OR2 (N1930, N1926, N1608);
xor XOR2 (N1931, N1909, N1817);
or OR4 (N1932, N1928, N48, N1248, N1536);
nand NAND4 (N1933, N1922, N1022, N1860, N621);
buf BUF1 (N1934, N1929);
buf BUF1 (N1935, N1930);
buf BUF1 (N1936, N1918);
buf BUF1 (N1937, N1916);
xor XOR2 (N1938, N1937, N441);
xor XOR2 (N1939, N1924, N380);
xor XOR2 (N1940, N1936, N650);
xor XOR2 (N1941, N1932, N559);
xor XOR2 (N1942, N1931, N685);
nand NAND2 (N1943, N1938, N1714);
xor XOR2 (N1944, N1943, N37);
nor NOR3 (N1945, N1942, N1467, N314);
buf BUF1 (N1946, N1935);
not NOT1 (N1947, N1946);
not NOT1 (N1948, N1920);
nor NOR3 (N1949, N1940, N379, N1870);
nor NOR3 (N1950, N1934, N423, N1276);
nor NOR4 (N1951, N1912, N1804, N196, N123);
nand NAND3 (N1952, N1950, N989, N1434);
not NOT1 (N1953, N1947);
buf BUF1 (N1954, N1933);
nor NOR3 (N1955, N1951, N469, N225);
xor XOR2 (N1956, N1941, N1072);
buf BUF1 (N1957, N1939);
nand NAND3 (N1958, N1956, N1423, N157);
xor XOR2 (N1959, N1955, N780);
or OR3 (N1960, N1957, N96, N630);
not NOT1 (N1961, N1960);
and AND4 (N1962, N1953, N1132, N49, N504);
not NOT1 (N1963, N1945);
nor NOR4 (N1964, N1952, N194, N1612, N1010);
nand NAND3 (N1965, N1963, N877, N269);
nand NAND2 (N1966, N1944, N1599);
nand NAND3 (N1967, N1958, N473, N552);
or OR4 (N1968, N1965, N1591, N673, N645);
or OR2 (N1969, N1968, N1724);
nand NAND2 (N1970, N1967, N1465);
not NOT1 (N1971, N1948);
xor XOR2 (N1972, N1959, N523);
not NOT1 (N1973, N1961);
nor NOR2 (N1974, N1966, N48);
not NOT1 (N1975, N1949);
buf BUF1 (N1976, N1969);
nand NAND4 (N1977, N1974, N34, N616, N1859);
buf BUF1 (N1978, N1973);
nand NAND4 (N1979, N1972, N880, N34, N825);
xor XOR2 (N1980, N1954, N1308);
nor NOR3 (N1981, N1980, N1077, N1245);
xor XOR2 (N1982, N1977, N215);
xor XOR2 (N1983, N1970, N317);
nor NOR4 (N1984, N1976, N374, N1221, N381);
buf BUF1 (N1985, N1984);
or OR3 (N1986, N1979, N1618, N521);
or OR3 (N1987, N1985, N1455, N1592);
and AND3 (N1988, N1964, N206, N1278);
xor XOR2 (N1989, N1981, N1946);
buf BUF1 (N1990, N1988);
nor NOR3 (N1991, N1982, N802, N1015);
buf BUF1 (N1992, N1978);
nand NAND2 (N1993, N1962, N133);
nand NAND4 (N1994, N1971, N93, N1304, N362);
or OR4 (N1995, N1987, N183, N1008, N730);
nand NAND4 (N1996, N1994, N458, N1389, N1359);
not NOT1 (N1997, N1989);
nor NOR2 (N1998, N1995, N337);
nand NAND2 (N1999, N1975, N1329);
not NOT1 (N2000, N1992);
nor NOR3 (N2001, N1986, N452, N1516);
buf BUF1 (N2002, N2000);
not NOT1 (N2003, N1999);
xor XOR2 (N2004, N1998, N1411);
nor NOR4 (N2005, N2002, N277, N1471, N697);
not NOT1 (N2006, N2005);
and AND2 (N2007, N2001, N1357);
buf BUF1 (N2008, N1993);
buf BUF1 (N2009, N2004);
nor NOR4 (N2010, N2007, N690, N636, N524);
and AND3 (N2011, N1983, N282, N1926);
nor NOR2 (N2012, N1990, N908);
nand NAND2 (N2013, N2009, N736);
xor XOR2 (N2014, N1996, N1444);
not NOT1 (N2015, N2012);
buf BUF1 (N2016, N2015);
buf BUF1 (N2017, N2016);
not NOT1 (N2018, N2008);
nor NOR2 (N2019, N2011, N761);
xor XOR2 (N2020, N2019, N1264);
not NOT1 (N2021, N2003);
buf BUF1 (N2022, N2018);
or OR2 (N2023, N1997, N446);
xor XOR2 (N2024, N2020, N673);
and AND4 (N2025, N2023, N287, N844, N1767);
and AND2 (N2026, N2017, N549);
buf BUF1 (N2027, N2024);
not NOT1 (N2028, N1991);
not NOT1 (N2029, N2010);
xor XOR2 (N2030, N2029, N1813);
buf BUF1 (N2031, N2027);
nand NAND2 (N2032, N2028, N1602);
or OR2 (N2033, N2021, N1592);
not NOT1 (N2034, N2006);
nor NOR3 (N2035, N2034, N1320, N1690);
nand NAND2 (N2036, N2013, N135);
xor XOR2 (N2037, N2033, N873);
and AND3 (N2038, N2035, N292, N1789);
xor XOR2 (N2039, N2038, N780);
or OR3 (N2040, N2031, N1039, N1371);
or OR3 (N2041, N2032, N88, N1729);
nand NAND4 (N2042, N2037, N1857, N1664, N1622);
and AND4 (N2043, N2026, N1767, N267, N808);
not NOT1 (N2044, N2043);
buf BUF1 (N2045, N2044);
and AND3 (N2046, N2041, N1267, N1163);
buf BUF1 (N2047, N2042);
nand NAND3 (N2048, N2022, N198, N1584);
nand NAND3 (N2049, N2048, N1057, N695);
xor XOR2 (N2050, N2045, N514);
nand NAND4 (N2051, N2047, N1997, N58, N4);
nor NOR3 (N2052, N2050, N909, N1120);
nor NOR3 (N2053, N2051, N1402, N594);
nor NOR3 (N2054, N2052, N1574, N1832);
buf BUF1 (N2055, N2014);
or OR3 (N2056, N2039, N1703, N897);
buf BUF1 (N2057, N2055);
not NOT1 (N2058, N2056);
nor NOR2 (N2059, N2030, N772);
nor NOR4 (N2060, N2046, N778, N407, N1297);
xor XOR2 (N2061, N2036, N1994);
buf BUF1 (N2062, N2057);
buf BUF1 (N2063, N2053);
xor XOR2 (N2064, N2062, N59);
xor XOR2 (N2065, N2061, N1028);
buf BUF1 (N2066, N2054);
xor XOR2 (N2067, N2040, N1955);
nor NOR4 (N2068, N2067, N2048, N1714, N544);
nand NAND4 (N2069, N2049, N790, N1971, N65);
and AND4 (N2070, N2059, N1748, N1236, N1124);
or OR4 (N2071, N2058, N441, N463, N451);
or OR3 (N2072, N2065, N895, N587);
nand NAND3 (N2073, N2060, N1877, N375);
nand NAND2 (N2074, N2071, N1628);
nor NOR3 (N2075, N2066, N355, N1930);
and AND2 (N2076, N2068, N2044);
nor NOR3 (N2077, N2075, N63, N991);
nand NAND3 (N2078, N2077, N761, N7);
or OR2 (N2079, N2064, N1166);
nor NOR2 (N2080, N2079, N1266);
or OR3 (N2081, N2070, N1381, N1852);
nor NOR3 (N2082, N2078, N1526, N571);
xor XOR2 (N2083, N2073, N1169);
and AND4 (N2084, N2082, N1896, N1508, N444);
not NOT1 (N2085, N2069);
or OR2 (N2086, N2072, N2037);
xor XOR2 (N2087, N2086, N132);
buf BUF1 (N2088, N2085);
not NOT1 (N2089, N2076);
or OR4 (N2090, N2087, N67, N869, N2069);
nor NOR3 (N2091, N2074, N344, N1017);
not NOT1 (N2092, N2080);
nand NAND2 (N2093, N2092, N1294);
nor NOR3 (N2094, N2084, N1284, N1829);
buf BUF1 (N2095, N2081);
or OR2 (N2096, N2091, N328);
xor XOR2 (N2097, N2090, N1391);
xor XOR2 (N2098, N2093, N1899);
and AND4 (N2099, N2097, N871, N591, N8);
nand NAND4 (N2100, N2095, N391, N1907, N334);
buf BUF1 (N2101, N2063);
or OR4 (N2102, N2096, N1354, N1350, N723);
not NOT1 (N2103, N2102);
and AND4 (N2104, N2100, N1679, N178, N812);
nor NOR2 (N2105, N2101, N856);
xor XOR2 (N2106, N2089, N1630);
buf BUF1 (N2107, N2088);
not NOT1 (N2108, N2104);
nand NAND3 (N2109, N2094, N1678, N1913);
xor XOR2 (N2110, N2025, N2002);
not NOT1 (N2111, N2103);
nand NAND2 (N2112, N2108, N1211);
not NOT1 (N2113, N2110);
xor XOR2 (N2114, N2111, N404);
buf BUF1 (N2115, N2098);
nand NAND3 (N2116, N2109, N275, N1735);
nand NAND2 (N2117, N2113, N817);
xor XOR2 (N2118, N2099, N1175);
xor XOR2 (N2119, N2106, N464);
nand NAND3 (N2120, N2117, N1006, N806);
and AND4 (N2121, N2119, N597, N158, N250);
xor XOR2 (N2122, N2121, N1174);
not NOT1 (N2123, N2118);
and AND2 (N2124, N2083, N92);
or OR2 (N2125, N2124, N291);
and AND3 (N2126, N2114, N1773, N1621);
not NOT1 (N2127, N2122);
or OR3 (N2128, N2112, N723, N1824);
nand NAND4 (N2129, N2125, N1989, N356, N35);
nand NAND3 (N2130, N2105, N2048, N1499);
and AND2 (N2131, N2115, N1536);
buf BUF1 (N2132, N2116);
and AND4 (N2133, N2130, N1019, N1311, N10);
and AND4 (N2134, N2126, N1402, N831, N114);
xor XOR2 (N2135, N2134, N1612);
not NOT1 (N2136, N2131);
not NOT1 (N2137, N2107);
and AND4 (N2138, N2123, N331, N690, N1705);
not NOT1 (N2139, N2133);
nor NOR3 (N2140, N2128, N1843, N1736);
not NOT1 (N2141, N2129);
buf BUF1 (N2142, N2141);
or OR3 (N2143, N2139, N1522, N1337);
buf BUF1 (N2144, N2138);
xor XOR2 (N2145, N2140, N502);
nand NAND3 (N2146, N2120, N412, N342);
xor XOR2 (N2147, N2142, N1715);
buf BUF1 (N2148, N2132);
xor XOR2 (N2149, N2135, N1431);
buf BUF1 (N2150, N2137);
xor XOR2 (N2151, N2143, N1437);
not NOT1 (N2152, N2147);
xor XOR2 (N2153, N2146, N974);
buf BUF1 (N2154, N2145);
or OR3 (N2155, N2136, N470, N2106);
nor NOR2 (N2156, N2151, N1479);
nor NOR2 (N2157, N2148, N1424);
nand NAND2 (N2158, N2152, N1100);
buf BUF1 (N2159, N2153);
and AND3 (N2160, N2154, N2093, N987);
and AND4 (N2161, N2150, N1717, N750, N531);
buf BUF1 (N2162, N2144);
or OR3 (N2163, N2162, N1945, N48);
xor XOR2 (N2164, N2159, N1761);
xor XOR2 (N2165, N2156, N1948);
buf BUF1 (N2166, N2161);
nor NOR4 (N2167, N2158, N1556, N1247, N863);
xor XOR2 (N2168, N2167, N1458);
xor XOR2 (N2169, N2165, N826);
nor NOR2 (N2170, N2149, N2138);
or OR4 (N2171, N2169, N515, N698, N1167);
and AND3 (N2172, N2163, N822, N1056);
and AND2 (N2173, N2160, N1898);
xor XOR2 (N2174, N2127, N1015);
and AND3 (N2175, N2171, N1660, N701);
nand NAND3 (N2176, N2164, N347, N1186);
xor XOR2 (N2177, N2176, N528);
nor NOR4 (N2178, N2166, N691, N1765, N886);
nand NAND3 (N2179, N2177, N1448, N1267);
xor XOR2 (N2180, N2172, N1088);
and AND4 (N2181, N2180, N82, N76, N219);
or OR2 (N2182, N2179, N1226);
or OR2 (N2183, N2181, N926);
not NOT1 (N2184, N2174);
or OR4 (N2185, N2184, N1962, N1214, N321);
nand NAND2 (N2186, N2178, N883);
not NOT1 (N2187, N2183);
or OR3 (N2188, N2168, N1214, N84);
or OR2 (N2189, N2186, N1867);
xor XOR2 (N2190, N2182, N977);
nand NAND2 (N2191, N2175, N636);
or OR3 (N2192, N2173, N2096, N1035);
or OR2 (N2193, N2155, N978);
nor NOR4 (N2194, N2157, N1410, N755, N1753);
and AND3 (N2195, N2189, N1058, N1293);
xor XOR2 (N2196, N2170, N47);
buf BUF1 (N2197, N2187);
nand NAND4 (N2198, N2194, N203, N1107, N1188);
nor NOR2 (N2199, N2196, N83);
nand NAND2 (N2200, N2188, N492);
nand NAND4 (N2201, N2200, N1919, N1339, N849);
buf BUF1 (N2202, N2195);
buf BUF1 (N2203, N2192);
not NOT1 (N2204, N2191);
nand NAND2 (N2205, N2190, N1309);
nor NOR3 (N2206, N2193, N1457, N871);
or OR2 (N2207, N2204, N387);
nand NAND3 (N2208, N2198, N340, N887);
or OR3 (N2209, N2185, N930, N461);
and AND2 (N2210, N2206, N1582);
nor NOR2 (N2211, N2199, N1079);
buf BUF1 (N2212, N2208);
or OR3 (N2213, N2202, N975, N940);
nand NAND3 (N2214, N2213, N1514, N798);
buf BUF1 (N2215, N2209);
not NOT1 (N2216, N2205);
and AND3 (N2217, N2197, N1526, N1457);
and AND2 (N2218, N2216, N1074);
and AND4 (N2219, N2215, N1676, N1836, N1232);
xor XOR2 (N2220, N2207, N1712);
nor NOR4 (N2221, N2211, N1743, N1862, N893);
xor XOR2 (N2222, N2212, N1130);
xor XOR2 (N2223, N2217, N340);
not NOT1 (N2224, N2220);
or OR2 (N2225, N2218, N1138);
or OR4 (N2226, N2203, N778, N501, N1685);
buf BUF1 (N2227, N2210);
nand NAND4 (N2228, N2226, N14, N2164, N1796);
xor XOR2 (N2229, N2228, N472);
not NOT1 (N2230, N2222);
and AND3 (N2231, N2214, N1358, N2158);
nand NAND3 (N2232, N2230, N2094, N592);
nand NAND4 (N2233, N2221, N2150, N1944, N199);
buf BUF1 (N2234, N2201);
nor NOR2 (N2235, N2233, N2112);
and AND3 (N2236, N2231, N613, N1728);
and AND3 (N2237, N2234, N177, N1546);
xor XOR2 (N2238, N2237, N251);
xor XOR2 (N2239, N2229, N1377);
nand NAND4 (N2240, N2219, N971, N1804, N994);
nand NAND2 (N2241, N2232, N1056);
or OR2 (N2242, N2223, N1898);
or OR2 (N2243, N2224, N2144);
nor NOR3 (N2244, N2235, N6, N1455);
buf BUF1 (N2245, N2242);
and AND4 (N2246, N2243, N1455, N231, N183);
nor NOR3 (N2247, N2239, N36, N1802);
or OR3 (N2248, N2238, N1999, N591);
nand NAND2 (N2249, N2225, N801);
nor NOR2 (N2250, N2241, N1783);
xor XOR2 (N2251, N2240, N1307);
and AND2 (N2252, N2248, N290);
or OR3 (N2253, N2244, N2036, N1716);
xor XOR2 (N2254, N2250, N34);
xor XOR2 (N2255, N2247, N947);
not NOT1 (N2256, N2253);
buf BUF1 (N2257, N2236);
or OR3 (N2258, N2256, N930, N2030);
and AND4 (N2259, N2255, N1107, N62, N1405);
and AND4 (N2260, N2249, N696, N1669, N540);
not NOT1 (N2261, N2245);
not NOT1 (N2262, N2261);
nor NOR3 (N2263, N2251, N1184, N507);
nor NOR2 (N2264, N2259, N939);
nand NAND4 (N2265, N2257, N1485, N1669, N2069);
xor XOR2 (N2266, N2258, N1562);
not NOT1 (N2267, N2264);
and AND4 (N2268, N2227, N1859, N1919, N684);
nand NAND3 (N2269, N2265, N1041, N799);
nand NAND3 (N2270, N2260, N1508, N280);
or OR3 (N2271, N2267, N1934, N771);
nand NAND4 (N2272, N2263, N1638, N1408, N1480);
and AND3 (N2273, N2271, N2069, N840);
and AND3 (N2274, N2266, N1531, N1177);
nor NOR2 (N2275, N2273, N1420);
or OR4 (N2276, N2252, N178, N1385, N1188);
xor XOR2 (N2277, N2254, N853);
and AND2 (N2278, N2268, N283);
and AND2 (N2279, N2277, N285);
buf BUF1 (N2280, N2246);
xor XOR2 (N2281, N2270, N465);
and AND3 (N2282, N2274, N193, N2185);
nand NAND4 (N2283, N2272, N1305, N792, N320);
nor NOR4 (N2284, N2282, N814, N316, N944);
nand NAND2 (N2285, N2269, N1346);
nand NAND4 (N2286, N2280, N308, N1545, N891);
and AND3 (N2287, N2279, N353, N1870);
and AND3 (N2288, N2276, N1809, N2129);
buf BUF1 (N2289, N2278);
xor XOR2 (N2290, N2287, N995);
or OR2 (N2291, N2288, N169);
or OR3 (N2292, N2275, N843, N64);
nor NOR2 (N2293, N2262, N717);
buf BUF1 (N2294, N2292);
not NOT1 (N2295, N2286);
nand NAND4 (N2296, N2289, N2092, N1264, N574);
nand NAND2 (N2297, N2284, N639);
nand NAND2 (N2298, N2285, N1467);
xor XOR2 (N2299, N2298, N1261);
nand NAND3 (N2300, N2283, N124, N1429);
not NOT1 (N2301, N2299);
nand NAND2 (N2302, N2296, N2093);
xor XOR2 (N2303, N2301, N2055);
nand NAND3 (N2304, N2295, N957, N1979);
nand NAND4 (N2305, N2303, N337, N14, N2268);
and AND2 (N2306, N2304, N1325);
or OR2 (N2307, N2294, N1272);
and AND2 (N2308, N2302, N138);
not NOT1 (N2309, N2290);
xor XOR2 (N2310, N2308, N1502);
buf BUF1 (N2311, N2291);
not NOT1 (N2312, N2306);
buf BUF1 (N2313, N2305);
nor NOR4 (N2314, N2312, N2154, N148, N487);
and AND4 (N2315, N2313, N464, N1692, N1419);
buf BUF1 (N2316, N2293);
and AND2 (N2317, N2297, N1543);
nand NAND2 (N2318, N2311, N1571);
nor NOR3 (N2319, N2317, N777, N1803);
and AND3 (N2320, N2281, N200, N1084);
nor NOR4 (N2321, N2318, N595, N1025, N838);
nand NAND3 (N2322, N2315, N1774, N513);
nor NOR2 (N2323, N2321, N1001);
buf BUF1 (N2324, N2323);
and AND3 (N2325, N2316, N1895, N2070);
buf BUF1 (N2326, N2300);
not NOT1 (N2327, N2326);
or OR2 (N2328, N2324, N40);
xor XOR2 (N2329, N2314, N1806);
nor NOR3 (N2330, N2319, N2308, N2245);
or OR3 (N2331, N2320, N673, N2155);
nand NAND3 (N2332, N2309, N1555, N725);
nor NOR2 (N2333, N2325, N1355);
or OR3 (N2334, N2307, N786, N2262);
or OR4 (N2335, N2332, N1486, N342, N977);
buf BUF1 (N2336, N2330);
buf BUF1 (N2337, N2329);
nor NOR3 (N2338, N2336, N1157, N24);
or OR4 (N2339, N2331, N2056, N262, N1873);
nand NAND2 (N2340, N2339, N2016);
nor NOR2 (N2341, N2337, N1313);
xor XOR2 (N2342, N2340, N1127);
and AND4 (N2343, N2338, N1909, N1651, N1988);
not NOT1 (N2344, N2341);
nand NAND4 (N2345, N2334, N45, N1683, N392);
not NOT1 (N2346, N2333);
or OR4 (N2347, N2327, N1075, N1146, N2205);
or OR4 (N2348, N2322, N1020, N388, N609);
nand NAND4 (N2349, N2348, N31, N628, N2278);
buf BUF1 (N2350, N2346);
and AND2 (N2351, N2345, N1945);
xor XOR2 (N2352, N2310, N1134);
or OR3 (N2353, N2347, N1773, N1246);
nor NOR4 (N2354, N2343, N502, N1340, N1769);
nand NAND2 (N2355, N2351, N1906);
xor XOR2 (N2356, N2353, N1550);
nor NOR4 (N2357, N2352, N594, N314, N1688);
xor XOR2 (N2358, N2342, N1701);
not NOT1 (N2359, N2357);
nor NOR3 (N2360, N2349, N1948, N786);
not NOT1 (N2361, N2350);
buf BUF1 (N2362, N2328);
buf BUF1 (N2363, N2360);
or OR3 (N2364, N2344, N849, N735);
xor XOR2 (N2365, N2356, N2052);
xor XOR2 (N2366, N2354, N1661);
and AND3 (N2367, N2364, N291, N1324);
or OR3 (N2368, N2363, N1951, N2019);
or OR2 (N2369, N2366, N2296);
or OR4 (N2370, N2335, N463, N924, N1167);
or OR4 (N2371, N2367, N1686, N18, N1485);
xor XOR2 (N2372, N2358, N1094);
nor NOR3 (N2373, N2365, N665, N2127);
or OR2 (N2374, N2369, N1222);
buf BUF1 (N2375, N2374);
or OR3 (N2376, N2359, N497, N59);
nor NOR4 (N2377, N2368, N1105, N296, N1663);
and AND2 (N2378, N2375, N2174);
buf BUF1 (N2379, N2371);
nor NOR3 (N2380, N2377, N938, N1973);
xor XOR2 (N2381, N2361, N776);
nor NOR4 (N2382, N2381, N1354, N1430, N1675);
and AND4 (N2383, N2372, N2235, N1553, N844);
buf BUF1 (N2384, N2370);
xor XOR2 (N2385, N2382, N2256);
buf BUF1 (N2386, N2383);
nand NAND2 (N2387, N2376, N2265);
not NOT1 (N2388, N2378);
not NOT1 (N2389, N2362);
not NOT1 (N2390, N2380);
nand NAND4 (N2391, N2373, N1133, N1411, N1793);
nor NOR3 (N2392, N2390, N1267, N2024);
buf BUF1 (N2393, N2385);
and AND3 (N2394, N2391, N1827, N1303);
and AND4 (N2395, N2392, N42, N2291, N1337);
nor NOR2 (N2396, N2394, N1449);
nor NOR4 (N2397, N2395, N757, N2319, N682);
and AND4 (N2398, N2379, N1183, N1959, N1737);
nand NAND3 (N2399, N2386, N1642, N1180);
and AND4 (N2400, N2389, N1489, N482, N2131);
nor NOR2 (N2401, N2384, N999);
buf BUF1 (N2402, N2398);
nor NOR3 (N2403, N2396, N2208, N307);
nor NOR4 (N2404, N2400, N1290, N1433, N1729);
or OR2 (N2405, N2388, N117);
nor NOR4 (N2406, N2401, N1428, N1847, N1046);
or OR4 (N2407, N2404, N2356, N758, N1580);
nor NOR3 (N2408, N2402, N431, N1088);
nor NOR2 (N2409, N2399, N993);
nand NAND3 (N2410, N2409, N1237, N197);
buf BUF1 (N2411, N2393);
not NOT1 (N2412, N2355);
xor XOR2 (N2413, N2410, N1369);
nand NAND4 (N2414, N2413, N241, N1200, N786);
or OR4 (N2415, N2412, N1409, N2192, N1256);
xor XOR2 (N2416, N2407, N1004);
buf BUF1 (N2417, N2403);
nand NAND3 (N2418, N2406, N260, N986);
or OR3 (N2419, N2416, N1621, N482);
or OR4 (N2420, N2387, N2408, N2388, N455);
or OR4 (N2421, N459, N704, N425, N1019);
not NOT1 (N2422, N2405);
nor NOR2 (N2423, N2421, N1573);
nor NOR3 (N2424, N2418, N791, N974);
not NOT1 (N2425, N2397);
or OR3 (N2426, N2415, N1830, N1089);
not NOT1 (N2427, N2419);
nand NAND4 (N2428, N2414, N406, N26, N384);
nand NAND3 (N2429, N2424, N1878, N1258);
buf BUF1 (N2430, N2411);
buf BUF1 (N2431, N2428);
or OR3 (N2432, N2426, N1774, N1509);
and AND2 (N2433, N2422, N2227);
nor NOR2 (N2434, N2425, N1311);
xor XOR2 (N2435, N2423, N202);
nor NOR2 (N2436, N2435, N1002);
and AND4 (N2437, N2433, N2295, N340, N356);
and AND4 (N2438, N2437, N2166, N2167, N919);
or OR2 (N2439, N2438, N1739);
buf BUF1 (N2440, N2427);
nor NOR3 (N2441, N2436, N604, N296);
nand NAND3 (N2442, N2439, N828, N1767);
and AND2 (N2443, N2431, N707);
buf BUF1 (N2444, N2441);
or OR4 (N2445, N2429, N470, N319, N1665);
or OR4 (N2446, N2444, N1013, N2365, N1505);
or OR4 (N2447, N2417, N158, N1478, N907);
and AND4 (N2448, N2434, N410, N1790, N1189);
not NOT1 (N2449, N2442);
nor NOR2 (N2450, N2446, N1389);
xor XOR2 (N2451, N2432, N125);
not NOT1 (N2452, N2420);
nand NAND3 (N2453, N2430, N574, N939);
xor XOR2 (N2454, N2451, N2381);
buf BUF1 (N2455, N2449);
and AND3 (N2456, N2445, N282, N2024);
xor XOR2 (N2457, N2448, N1093);
nor NOR4 (N2458, N2455, N1237, N607, N167);
not NOT1 (N2459, N2454);
and AND4 (N2460, N2459, N1032, N939, N1202);
or OR2 (N2461, N2456, N948);
not NOT1 (N2462, N2452);
nand NAND3 (N2463, N2457, N1980, N1404);
not NOT1 (N2464, N2453);
or OR4 (N2465, N2440, N2040, N2155, N419);
nand NAND2 (N2466, N2450, N31);
or OR3 (N2467, N2458, N165, N687);
nor NOR4 (N2468, N2461, N1831, N638, N2014);
nand NAND3 (N2469, N2468, N242, N68);
nand NAND3 (N2470, N2462, N214, N964);
not NOT1 (N2471, N2443);
nand NAND2 (N2472, N2460, N1414);
not NOT1 (N2473, N2464);
and AND3 (N2474, N2473, N119, N609);
nor NOR4 (N2475, N2466, N450, N633, N748);
or OR4 (N2476, N2447, N1389, N2344, N775);
or OR2 (N2477, N2465, N1828);
not NOT1 (N2478, N2470);
and AND3 (N2479, N2471, N1883, N124);
not NOT1 (N2480, N2475);
buf BUF1 (N2481, N2467);
buf BUF1 (N2482, N2478);
nand NAND3 (N2483, N2472, N2157, N917);
nand NAND2 (N2484, N2476, N1649);
and AND3 (N2485, N2474, N1017, N1913);
buf BUF1 (N2486, N2484);
nand NAND2 (N2487, N2479, N1241);
nor NOR3 (N2488, N2477, N2246, N1384);
nor NOR3 (N2489, N2487, N1479, N1903);
xor XOR2 (N2490, N2485, N2399);
xor XOR2 (N2491, N2490, N1687);
nor NOR3 (N2492, N2482, N1908, N1458);
nor NOR4 (N2493, N2480, N2197, N627, N1926);
or OR4 (N2494, N2491, N2314, N1588, N426);
buf BUF1 (N2495, N2463);
and AND2 (N2496, N2495, N282);
xor XOR2 (N2497, N2489, N355);
not NOT1 (N2498, N2496);
nor NOR4 (N2499, N2498, N259, N2375, N2481);
or OR4 (N2500, N1668, N1431, N1275, N447);
xor XOR2 (N2501, N2483, N1402);
xor XOR2 (N2502, N2486, N1168);
xor XOR2 (N2503, N2492, N1821);
nor NOR3 (N2504, N2501, N679, N421);
xor XOR2 (N2505, N2497, N1559);
and AND4 (N2506, N2488, N889, N24, N270);
or OR4 (N2507, N2493, N136, N735, N721);
nor NOR4 (N2508, N2504, N325, N1717, N2466);
nor NOR2 (N2509, N2506, N1527);
and AND2 (N2510, N2500, N2491);
nor NOR4 (N2511, N2499, N1309, N6, N933);
and AND4 (N2512, N2494, N966, N1893, N1716);
buf BUF1 (N2513, N2512);
nor NOR3 (N2514, N2510, N292, N88);
buf BUF1 (N2515, N2502);
and AND4 (N2516, N2514, N1801, N2145, N1626);
buf BUF1 (N2517, N2516);
and AND4 (N2518, N2503, N1747, N353, N1933);
or OR3 (N2519, N2518, N289, N390);
xor XOR2 (N2520, N2511, N260);
xor XOR2 (N2521, N2505, N194);
or OR4 (N2522, N2519, N1456, N2438, N1904);
nor NOR2 (N2523, N2520, N2179);
nor NOR2 (N2524, N2521, N2048);
xor XOR2 (N2525, N2517, N1878);
xor XOR2 (N2526, N2513, N2375);
not NOT1 (N2527, N2525);
xor XOR2 (N2528, N2507, N1289);
not NOT1 (N2529, N2509);
or OR3 (N2530, N2469, N894, N2219);
not NOT1 (N2531, N2523);
xor XOR2 (N2532, N2527, N1897);
or OR2 (N2533, N2529, N2036);
not NOT1 (N2534, N2530);
nor NOR2 (N2535, N2515, N131);
xor XOR2 (N2536, N2508, N2447);
and AND4 (N2537, N2534, N2263, N1932, N2317);
not NOT1 (N2538, N2522);
not NOT1 (N2539, N2533);
or OR2 (N2540, N2528, N1233);
buf BUF1 (N2541, N2531);
and AND3 (N2542, N2537, N276, N758);
nor NOR2 (N2543, N2541, N557);
buf BUF1 (N2544, N2543);
not NOT1 (N2545, N2526);
buf BUF1 (N2546, N2544);
nand NAND4 (N2547, N2532, N1359, N380, N1874);
or OR2 (N2548, N2542, N1399);
xor XOR2 (N2549, N2524, N1968);
xor XOR2 (N2550, N2547, N1778);
nand NAND3 (N2551, N2540, N1646, N390);
xor XOR2 (N2552, N2548, N2006);
and AND2 (N2553, N2546, N518);
or OR3 (N2554, N2552, N751, N2171);
nand NAND3 (N2555, N2550, N1187, N2319);
or OR3 (N2556, N2539, N1226, N685);
and AND3 (N2557, N2535, N429, N1694);
and AND4 (N2558, N2549, N203, N2058, N278);
not NOT1 (N2559, N2554);
nand NAND2 (N2560, N2545, N2315);
buf BUF1 (N2561, N2560);
not NOT1 (N2562, N2556);
or OR3 (N2563, N2559, N2496, N454);
nand NAND3 (N2564, N2553, N2505, N622);
or OR2 (N2565, N2536, N310);
nor NOR3 (N2566, N2561, N1290, N298);
nor NOR3 (N2567, N2557, N2463, N2492);
xor XOR2 (N2568, N2558, N1422);
or OR3 (N2569, N2538, N2106, N1716);
nand NAND4 (N2570, N2555, N1915, N674, N2133);
or OR4 (N2571, N2562, N1282, N834, N243);
buf BUF1 (N2572, N2551);
nor NOR3 (N2573, N2563, N1747, N428);
buf BUF1 (N2574, N2573);
nand NAND2 (N2575, N2567, N881);
xor XOR2 (N2576, N2574, N693);
buf BUF1 (N2577, N2572);
and AND3 (N2578, N2570, N1632, N1931);
not NOT1 (N2579, N2565);
nor NOR2 (N2580, N2568, N2415);
xor XOR2 (N2581, N2577, N832);
xor XOR2 (N2582, N2578, N1022);
and AND2 (N2583, N2579, N1098);
nor NOR3 (N2584, N2582, N1578, N1777);
buf BUF1 (N2585, N2584);
or OR3 (N2586, N2583, N998, N1639);
not NOT1 (N2587, N2585);
not NOT1 (N2588, N2580);
nor NOR2 (N2589, N2575, N1671);
nand NAND2 (N2590, N2569, N847);
nor NOR4 (N2591, N2588, N1369, N923, N1517);
buf BUF1 (N2592, N2571);
or OR2 (N2593, N2564, N1622);
nand NAND2 (N2594, N2589, N2302);
not NOT1 (N2595, N2594);
buf BUF1 (N2596, N2581);
buf BUF1 (N2597, N2596);
buf BUF1 (N2598, N2576);
or OR4 (N2599, N2598, N1511, N341, N1781);
nand NAND2 (N2600, N2566, N240);
nand NAND3 (N2601, N2599, N1271, N1587);
buf BUF1 (N2602, N2587);
or OR3 (N2603, N2602, N975, N1879);
xor XOR2 (N2604, N2590, N1932);
nand NAND3 (N2605, N2601, N772, N1108);
nand NAND4 (N2606, N2593, N1895, N2154, N1793);
xor XOR2 (N2607, N2605, N2091);
and AND3 (N2608, N2592, N2185, N831);
nor NOR2 (N2609, N2586, N1610);
nand NAND3 (N2610, N2600, N1698, N730);
not NOT1 (N2611, N2591);
xor XOR2 (N2612, N2610, N983);
not NOT1 (N2613, N2597);
not NOT1 (N2614, N2595);
and AND2 (N2615, N2607, N228);
nand NAND4 (N2616, N2612, N1354, N44, N668);
not NOT1 (N2617, N2616);
xor XOR2 (N2618, N2617, N1563);
nor NOR4 (N2619, N2604, N1748, N2336, N1512);
xor XOR2 (N2620, N2606, N1602);
and AND2 (N2621, N2620, N2370);
not NOT1 (N2622, N2614);
buf BUF1 (N2623, N2619);
buf BUF1 (N2624, N2622);
buf BUF1 (N2625, N2613);
and AND3 (N2626, N2603, N2311, N687);
xor XOR2 (N2627, N2611, N1041);
and AND4 (N2628, N2618, N1870, N189, N2303);
and AND2 (N2629, N2624, N2481);
and AND2 (N2630, N2615, N2484);
nor NOR2 (N2631, N2623, N2003);
nor NOR2 (N2632, N2626, N591);
buf BUF1 (N2633, N2632);
nor NOR3 (N2634, N2628, N250, N2607);
not NOT1 (N2635, N2609);
and AND3 (N2636, N2627, N630, N413);
xor XOR2 (N2637, N2625, N938);
and AND4 (N2638, N2631, N873, N1291, N211);
nand NAND4 (N2639, N2636, N1242, N2069, N2124);
not NOT1 (N2640, N2621);
xor XOR2 (N2641, N2634, N695);
nand NAND2 (N2642, N2641, N839);
xor XOR2 (N2643, N2630, N435);
xor XOR2 (N2644, N2633, N1253);
buf BUF1 (N2645, N2644);
nor NOR2 (N2646, N2642, N2215);
not NOT1 (N2647, N2608);
nand NAND2 (N2648, N2647, N1780);
not NOT1 (N2649, N2645);
nor NOR2 (N2650, N2638, N1637);
buf BUF1 (N2651, N2650);
not NOT1 (N2652, N2651);
nor NOR3 (N2653, N2646, N967, N414);
not NOT1 (N2654, N2640);
and AND4 (N2655, N2637, N1154, N2241, N1205);
not NOT1 (N2656, N2648);
nor NOR3 (N2657, N2654, N1394, N843);
or OR2 (N2658, N2629, N1012);
buf BUF1 (N2659, N2658);
and AND4 (N2660, N2653, N406, N2434, N1634);
xor XOR2 (N2661, N2655, N1983);
xor XOR2 (N2662, N2652, N699);
nor NOR3 (N2663, N2649, N2462, N1961);
or OR2 (N2664, N2657, N2071);
xor XOR2 (N2665, N2664, N421);
xor XOR2 (N2666, N2659, N2440);
or OR3 (N2667, N2663, N1303, N1920);
or OR2 (N2668, N2639, N1600);
xor XOR2 (N2669, N2661, N285);
and AND4 (N2670, N2665, N1613, N1035, N203);
buf BUF1 (N2671, N2643);
nand NAND3 (N2672, N2670, N989, N859);
not NOT1 (N2673, N2671);
buf BUF1 (N2674, N2669);
not NOT1 (N2675, N2666);
nand NAND4 (N2676, N2656, N2397, N1988, N2523);
nand NAND4 (N2677, N2668, N713, N235, N9);
xor XOR2 (N2678, N2660, N415);
buf BUF1 (N2679, N2635);
nor NOR3 (N2680, N2675, N1460, N311);
xor XOR2 (N2681, N2667, N2351);
and AND4 (N2682, N2674, N1808, N1924, N834);
not NOT1 (N2683, N2672);
xor XOR2 (N2684, N2662, N204);
nor NOR3 (N2685, N2681, N2429, N402);
not NOT1 (N2686, N2673);
buf BUF1 (N2687, N2682);
not NOT1 (N2688, N2683);
not NOT1 (N2689, N2680);
nand NAND4 (N2690, N2687, N2519, N1180, N1314);
nand NAND3 (N2691, N2679, N2501, N1647);
nand NAND4 (N2692, N2684, N981, N2517, N715);
not NOT1 (N2693, N2686);
not NOT1 (N2694, N2693);
nand NAND2 (N2695, N2685, N2184);
xor XOR2 (N2696, N2691, N394);
xor XOR2 (N2697, N2676, N306);
or OR4 (N2698, N2690, N2072, N694, N1938);
buf BUF1 (N2699, N2695);
buf BUF1 (N2700, N2689);
not NOT1 (N2701, N2696);
and AND4 (N2702, N2677, N1185, N2404, N1953);
buf BUF1 (N2703, N2692);
or OR2 (N2704, N2699, N795);
or OR2 (N2705, N2694, N1076);
or OR2 (N2706, N2701, N1383);
nand NAND3 (N2707, N2702, N30, N1947);
xor XOR2 (N2708, N2698, N2567);
and AND2 (N2709, N2688, N170);
xor XOR2 (N2710, N2705, N1935);
nor NOR2 (N2711, N2697, N2388);
not NOT1 (N2712, N2704);
or OR2 (N2713, N2678, N201);
and AND4 (N2714, N2706, N1863, N211, N2278);
buf BUF1 (N2715, N2703);
buf BUF1 (N2716, N2713);
nor NOR2 (N2717, N2711, N885);
and AND2 (N2718, N2710, N1151);
not NOT1 (N2719, N2707);
not NOT1 (N2720, N2708);
nand NAND3 (N2721, N2717, N1135, N702);
and AND3 (N2722, N2700, N1566, N1134);
xor XOR2 (N2723, N2719, N508);
buf BUF1 (N2724, N2716);
and AND3 (N2725, N2724, N2088, N865);
nor NOR4 (N2726, N2712, N1738, N562, N1593);
buf BUF1 (N2727, N2720);
or OR2 (N2728, N2721, N834);
not NOT1 (N2729, N2709);
buf BUF1 (N2730, N2714);
not NOT1 (N2731, N2728);
or OR2 (N2732, N2727, N206);
nor NOR2 (N2733, N2723, N585);
buf BUF1 (N2734, N2729);
xor XOR2 (N2735, N2726, N2152);
nor NOR4 (N2736, N2732, N2611, N2133, N2112);
not NOT1 (N2737, N2730);
or OR2 (N2738, N2736, N2615);
nor NOR2 (N2739, N2734, N1681);
buf BUF1 (N2740, N2725);
and AND4 (N2741, N2718, N1382, N1676, N571);
and AND2 (N2742, N2731, N848);
xor XOR2 (N2743, N2722, N1860);
and AND2 (N2744, N2735, N911);
and AND3 (N2745, N2739, N2658, N1607);
buf BUF1 (N2746, N2745);
not NOT1 (N2747, N2746);
nor NOR3 (N2748, N2741, N1181, N2543);
nand NAND4 (N2749, N2740, N96, N2354, N683);
or OR2 (N2750, N2737, N1613);
nor NOR4 (N2751, N2715, N2247, N586, N555);
nand NAND4 (N2752, N2747, N109, N1184, N2144);
nand NAND4 (N2753, N2752, N1983, N1510, N1222);
nand NAND2 (N2754, N2748, N896);
xor XOR2 (N2755, N2742, N2024);
and AND2 (N2756, N2743, N640);
and AND3 (N2757, N2753, N735, N395);
and AND4 (N2758, N2754, N2443, N1074, N146);
buf BUF1 (N2759, N2749);
xor XOR2 (N2760, N2758, N573);
not NOT1 (N2761, N2750);
or OR4 (N2762, N2733, N398, N1219, N2216);
xor XOR2 (N2763, N2759, N1230);
xor XOR2 (N2764, N2744, N2751);
buf BUF1 (N2765, N2653);
xor XOR2 (N2766, N2755, N2392);
buf BUF1 (N2767, N2764);
or OR2 (N2768, N2766, N491);
not NOT1 (N2769, N2763);
and AND2 (N2770, N2756, N2014);
buf BUF1 (N2771, N2757);
not NOT1 (N2772, N2767);
xor XOR2 (N2773, N2769, N2527);
nand NAND3 (N2774, N2770, N1643, N2119);
nor NOR2 (N2775, N2762, N1188);
nand NAND3 (N2776, N2773, N155, N2087);
xor XOR2 (N2777, N2776, N2112);
nand NAND3 (N2778, N2774, N1174, N2033);
xor XOR2 (N2779, N2778, N936);
and AND3 (N2780, N2772, N1763, N1755);
not NOT1 (N2781, N2779);
nand NAND4 (N2782, N2781, N32, N1491, N601);
xor XOR2 (N2783, N2768, N1796);
nor NOR4 (N2784, N2783, N830, N2460, N929);
nor NOR3 (N2785, N2765, N1740, N2044);
buf BUF1 (N2786, N2785);
buf BUF1 (N2787, N2784);
buf BUF1 (N2788, N2780);
xor XOR2 (N2789, N2788, N2204);
xor XOR2 (N2790, N2777, N1904);
nor NOR4 (N2791, N2761, N427, N1117, N269);
or OR2 (N2792, N2738, N689);
or OR4 (N2793, N2760, N526, N1706, N851);
and AND3 (N2794, N2786, N680, N1298);
nor NOR2 (N2795, N2775, N1982);
or OR4 (N2796, N2793, N1525, N776, N695);
nand NAND2 (N2797, N2795, N2626);
and AND4 (N2798, N2789, N1352, N2744, N1392);
not NOT1 (N2799, N2790);
nand NAND4 (N2800, N2792, N2117, N1088, N1261);
nand NAND3 (N2801, N2800, N2776, N1527);
nand NAND2 (N2802, N2796, N1133);
or OR4 (N2803, N2787, N1096, N417, N2050);
and AND2 (N2804, N2799, N2585);
not NOT1 (N2805, N2801);
nand NAND4 (N2806, N2805, N2397, N2021, N1070);
buf BUF1 (N2807, N2804);
and AND2 (N2808, N2797, N9);
nand NAND4 (N2809, N2771, N2138, N1538, N2084);
not NOT1 (N2810, N2782);
not NOT1 (N2811, N2809);
not NOT1 (N2812, N2810);
xor XOR2 (N2813, N2794, N1700);
not NOT1 (N2814, N2791);
nand NAND3 (N2815, N2802, N1153, N2687);
nand NAND3 (N2816, N2814, N645, N1096);
xor XOR2 (N2817, N2812, N427);
nor NOR3 (N2818, N2813, N1738, N2047);
or OR4 (N2819, N2806, N2618, N55, N2705);
nor NOR2 (N2820, N2817, N24);
and AND3 (N2821, N2816, N2688, N1107);
nand NAND2 (N2822, N2803, N1380);
nand NAND3 (N2823, N2811, N1128, N63);
buf BUF1 (N2824, N2822);
and AND2 (N2825, N2808, N2270);
xor XOR2 (N2826, N2819, N1301);
nor NOR4 (N2827, N2815, N1332, N2007, N1806);
buf BUF1 (N2828, N2821);
nor NOR2 (N2829, N2825, N829);
xor XOR2 (N2830, N2798, N900);
buf BUF1 (N2831, N2820);
buf BUF1 (N2832, N2830);
xor XOR2 (N2833, N2832, N69);
xor XOR2 (N2834, N2823, N2296);
or OR3 (N2835, N2831, N1270, N1441);
and AND3 (N2836, N2829, N1232, N2143);
not NOT1 (N2837, N2824);
buf BUF1 (N2838, N2807);
not NOT1 (N2839, N2836);
or OR2 (N2840, N2834, N91);
not NOT1 (N2841, N2826);
nand NAND2 (N2842, N2841, N165);
xor XOR2 (N2843, N2842, N1985);
buf BUF1 (N2844, N2828);
xor XOR2 (N2845, N2843, N959);
not NOT1 (N2846, N2840);
and AND4 (N2847, N2833, N2806, N1572, N882);
buf BUF1 (N2848, N2846);
not NOT1 (N2849, N2837);
and AND3 (N2850, N2839, N2218, N829);
buf BUF1 (N2851, N2847);
xor XOR2 (N2852, N2835, N1238);
and AND2 (N2853, N2838, N2736);
nand NAND3 (N2854, N2849, N582, N1072);
xor XOR2 (N2855, N2827, N1809);
nor NOR4 (N2856, N2854, N903, N1153, N115);
or OR4 (N2857, N2845, N802, N1315, N2622);
buf BUF1 (N2858, N2818);
nor NOR3 (N2859, N2857, N1244, N1165);
nand NAND2 (N2860, N2853, N2194);
or OR4 (N2861, N2859, N2667, N1399, N208);
buf BUF1 (N2862, N2856);
xor XOR2 (N2863, N2852, N2629);
buf BUF1 (N2864, N2850);
buf BUF1 (N2865, N2862);
and AND4 (N2866, N2844, N822, N560, N2761);
buf BUF1 (N2867, N2861);
nor NOR4 (N2868, N2864, N1504, N2612, N1543);
not NOT1 (N2869, N2863);
and AND3 (N2870, N2860, N2485, N352);
not NOT1 (N2871, N2865);
xor XOR2 (N2872, N2855, N1990);
nand NAND4 (N2873, N2848, N1223, N1361, N2643);
buf BUF1 (N2874, N2866);
xor XOR2 (N2875, N2868, N2580);
or OR4 (N2876, N2875, N2560, N49, N2843);
or OR4 (N2877, N2876, N1499, N2764, N1073);
xor XOR2 (N2878, N2851, N95);
buf BUF1 (N2879, N2871);
buf BUF1 (N2880, N2873);
nor NOR3 (N2881, N2869, N2359, N1111);
or OR3 (N2882, N2872, N1561, N199);
xor XOR2 (N2883, N2881, N2781);
buf BUF1 (N2884, N2878);
and AND4 (N2885, N2883, N2200, N101, N2320);
xor XOR2 (N2886, N2880, N2788);
buf BUF1 (N2887, N2885);
xor XOR2 (N2888, N2887, N1776);
and AND3 (N2889, N2884, N1210, N882);
buf BUF1 (N2890, N2870);
not NOT1 (N2891, N2889);
or OR2 (N2892, N2888, N1207);
nor NOR3 (N2893, N2858, N687, N2435);
and AND4 (N2894, N2886, N1801, N2430, N2859);
nand NAND3 (N2895, N2882, N655, N1029);
or OR2 (N2896, N2879, N2494);
not NOT1 (N2897, N2893);
or OR3 (N2898, N2877, N134, N1724);
and AND4 (N2899, N2890, N1415, N1526, N1830);
nor NOR3 (N2900, N2896, N2348, N2050);
nor NOR3 (N2901, N2867, N866, N2007);
or OR3 (N2902, N2892, N670, N201);
xor XOR2 (N2903, N2899, N553);
buf BUF1 (N2904, N2894);
nor NOR4 (N2905, N2904, N1850, N1329, N2723);
or OR2 (N2906, N2905, N1871);
or OR3 (N2907, N2901, N1716, N788);
nand NAND4 (N2908, N2874, N1033, N2215, N1789);
xor XOR2 (N2909, N2891, N2375);
not NOT1 (N2910, N2906);
nand NAND4 (N2911, N2898, N2077, N398, N2192);
xor XOR2 (N2912, N2903, N203);
buf BUF1 (N2913, N2907);
xor XOR2 (N2914, N2911, N2457);
and AND4 (N2915, N2895, N767, N430, N1613);
and AND4 (N2916, N2910, N2329, N1097, N48);
or OR2 (N2917, N2897, N655);
not NOT1 (N2918, N2917);
xor XOR2 (N2919, N2908, N2483);
xor XOR2 (N2920, N2909, N189);
or OR4 (N2921, N2902, N309, N657, N1782);
buf BUF1 (N2922, N2900);
not NOT1 (N2923, N2918);
xor XOR2 (N2924, N2923, N1850);
or OR4 (N2925, N2920, N1758, N2915, N1792);
nor NOR4 (N2926, N1093, N1783, N2354, N745);
nor NOR2 (N2927, N2913, N751);
xor XOR2 (N2928, N2925, N9);
nor NOR2 (N2929, N2912, N2097);
xor XOR2 (N2930, N2916, N830);
and AND2 (N2931, N2919, N722);
or OR3 (N2932, N2928, N1977, N839);
nand NAND2 (N2933, N2914, N1092);
nor NOR2 (N2934, N2932, N2835);
nand NAND3 (N2935, N2933, N2841, N738);
nor NOR3 (N2936, N2922, N829, N1589);
and AND3 (N2937, N2935, N164, N2031);
nand NAND2 (N2938, N2921, N1565);
nor NOR3 (N2939, N2936, N535, N966);
nand NAND4 (N2940, N2930, N967, N2773, N241);
nor NOR4 (N2941, N2938, N216, N1330, N386);
nor NOR2 (N2942, N2941, N927);
buf BUF1 (N2943, N2940);
not NOT1 (N2944, N2924);
or OR2 (N2945, N2944, N2163);
xor XOR2 (N2946, N2926, N2261);
not NOT1 (N2947, N2931);
buf BUF1 (N2948, N2929);
not NOT1 (N2949, N2948);
xor XOR2 (N2950, N2949, N1560);
nand NAND2 (N2951, N2927, N169);
buf BUF1 (N2952, N2934);
and AND2 (N2953, N2939, N2212);
or OR4 (N2954, N2946, N1414, N2054, N933);
buf BUF1 (N2955, N2954);
or OR4 (N2956, N2945, N1361, N1403, N2663);
or OR4 (N2957, N2953, N1226, N2829, N1568);
buf BUF1 (N2958, N2957);
nand NAND3 (N2959, N2937, N2044, N1367);
xor XOR2 (N2960, N2956, N1597);
nor NOR4 (N2961, N2951, N549, N1033, N2468);
nor NOR4 (N2962, N2961, N1897, N1066, N2464);
nand NAND4 (N2963, N2960, N174, N859, N1002);
and AND4 (N2964, N2962, N2627, N2165, N1886);
and AND2 (N2965, N2955, N2014);
buf BUF1 (N2966, N2963);
buf BUF1 (N2967, N2942);
or OR4 (N2968, N2964, N268, N2413, N2234);
xor XOR2 (N2969, N2959, N1136);
nor NOR3 (N2970, N2968, N1470, N109);
xor XOR2 (N2971, N2966, N1228);
buf BUF1 (N2972, N2971);
nor NOR4 (N2973, N2950, N926, N996, N218);
nand NAND2 (N2974, N2969, N175);
or OR3 (N2975, N2952, N564, N2647);
and AND3 (N2976, N2943, N875, N2488);
nor NOR3 (N2977, N2965, N1422, N137);
or OR2 (N2978, N2977, N2066);
nor NOR2 (N2979, N2974, N2878);
and AND3 (N2980, N2958, N1351, N130);
not NOT1 (N2981, N2973);
buf BUF1 (N2982, N2976);
nand NAND4 (N2983, N2972, N1588, N1012, N827);
nor NOR2 (N2984, N2975, N2805);
or OR3 (N2985, N2982, N743, N1978);
or OR4 (N2986, N2978, N564, N1741, N1494);
xor XOR2 (N2987, N2983, N1525);
nand NAND3 (N2988, N2970, N1722, N391);
and AND3 (N2989, N2967, N2389, N871);
or OR3 (N2990, N2989, N2761, N1120);
not NOT1 (N2991, N2979);
xor XOR2 (N2992, N2990, N1230);
or OR2 (N2993, N2980, N1577);
xor XOR2 (N2994, N2984, N456);
or OR3 (N2995, N2994, N1160, N1640);
not NOT1 (N2996, N2981);
or OR2 (N2997, N2985, N1626);
or OR3 (N2998, N2988, N2713, N1640);
and AND2 (N2999, N2998, N683);
nor NOR2 (N3000, N2997, N646);
or OR2 (N3001, N2996, N2368);
and AND3 (N3002, N2995, N2738, N984);
or OR4 (N3003, N2991, N410, N1793, N335);
xor XOR2 (N3004, N2999, N1224);
not NOT1 (N3005, N3004);
and AND3 (N3006, N2947, N801, N544);
not NOT1 (N3007, N2993);
xor XOR2 (N3008, N2992, N1348);
or OR4 (N3009, N2987, N2452, N2702, N1015);
or OR2 (N3010, N3001, N826);
xor XOR2 (N3011, N2986, N2920);
not NOT1 (N3012, N3005);
buf BUF1 (N3013, N3003);
nor NOR2 (N3014, N3002, N1700);
and AND3 (N3015, N3007, N2171, N2561);
and AND4 (N3016, N3011, N1443, N1203, N2093);
not NOT1 (N3017, N3000);
not NOT1 (N3018, N3016);
buf BUF1 (N3019, N3017);
or OR3 (N3020, N3013, N412, N1735);
buf BUF1 (N3021, N3015);
nor NOR2 (N3022, N3014, N24);
buf BUF1 (N3023, N3006);
and AND3 (N3024, N3012, N1699, N2718);
and AND2 (N3025, N3019, N1353);
not NOT1 (N3026, N3018);
not NOT1 (N3027, N3023);
not NOT1 (N3028, N3026);
buf BUF1 (N3029, N3020);
nor NOR3 (N3030, N3022, N2331, N2385);
or OR3 (N3031, N3028, N1836, N1905);
nor NOR2 (N3032, N3021, N977);
buf BUF1 (N3033, N3010);
buf BUF1 (N3034, N3029);
buf BUF1 (N3035, N3031);
xor XOR2 (N3036, N3034, N88);
buf BUF1 (N3037, N3027);
nand NAND3 (N3038, N3024, N1555, N484);
nand NAND4 (N3039, N3025, N2834, N1493, N2600);
or OR2 (N3040, N3030, N1652);
xor XOR2 (N3041, N3037, N1141);
or OR3 (N3042, N3040, N179, N1135);
and AND3 (N3043, N3033, N807, N1919);
and AND3 (N3044, N3009, N1735, N1835);
nand NAND3 (N3045, N3044, N1982, N2147);
and AND4 (N3046, N3032, N664, N2293, N1579);
nand NAND4 (N3047, N3039, N2526, N469, N374);
not NOT1 (N3048, N3042);
nand NAND3 (N3049, N3035, N230, N1567);
xor XOR2 (N3050, N3045, N2867);
and AND3 (N3051, N3041, N2475, N2720);
xor XOR2 (N3052, N3038, N1984);
and AND2 (N3053, N3046, N2729);
xor XOR2 (N3054, N3043, N2973);
not NOT1 (N3055, N3054);
xor XOR2 (N3056, N3050, N2136);
nand NAND2 (N3057, N3056, N2739);
nor NOR2 (N3058, N3048, N1855);
buf BUF1 (N3059, N3051);
nor NOR4 (N3060, N3052, N2943, N1450, N1916);
or OR3 (N3061, N3059, N861, N2950);
xor XOR2 (N3062, N3053, N1219);
or OR2 (N3063, N3049, N2626);
and AND2 (N3064, N3060, N2581);
or OR3 (N3065, N3047, N263, N1435);
not NOT1 (N3066, N3057);
nor NOR4 (N3067, N3065, N1596, N556, N2887);
not NOT1 (N3068, N3062);
and AND3 (N3069, N3008, N2965, N1339);
or OR4 (N3070, N3036, N2230, N364, N434);
xor XOR2 (N3071, N3061, N349);
nand NAND2 (N3072, N3058, N2223);
nand NAND2 (N3073, N3063, N2242);
or OR2 (N3074, N3055, N476);
buf BUF1 (N3075, N3074);
not NOT1 (N3076, N3067);
or OR2 (N3077, N3076, N534);
xor XOR2 (N3078, N3064, N2082);
xor XOR2 (N3079, N3070, N1600);
and AND2 (N3080, N3075, N2163);
buf BUF1 (N3081, N3080);
nand NAND3 (N3082, N3071, N2929, N1110);
not NOT1 (N3083, N3081);
nor NOR2 (N3084, N3073, N643);
nand NAND3 (N3085, N3072, N1403, N925);
or OR4 (N3086, N3082, N260, N380, N892);
and AND2 (N3087, N3083, N390);
not NOT1 (N3088, N3086);
not NOT1 (N3089, N3069);
nand NAND3 (N3090, N3084, N2634, N1513);
or OR3 (N3091, N3079, N590, N1710);
nor NOR2 (N3092, N3087, N2675);
xor XOR2 (N3093, N3077, N2594);
not NOT1 (N3094, N3078);
nand NAND2 (N3095, N3068, N729);
not NOT1 (N3096, N3090);
buf BUF1 (N3097, N3091);
and AND3 (N3098, N3097, N626, N315);
and AND2 (N3099, N3095, N2390);
or OR4 (N3100, N3098, N656, N88, N310);
xor XOR2 (N3101, N3085, N2658);
nor NOR4 (N3102, N3094, N348, N617, N1286);
nand NAND4 (N3103, N3088, N1435, N1195, N548);
nand NAND4 (N3104, N3103, N1545, N1397, N1393);
buf BUF1 (N3105, N3102);
nand NAND3 (N3106, N3096, N2554, N2891);
xor XOR2 (N3107, N3099, N2918);
nor NOR2 (N3108, N3066, N1308);
xor XOR2 (N3109, N3093, N1590);
or OR4 (N3110, N3107, N2681, N276, N1309);
nand NAND3 (N3111, N3100, N813, N1733);
or OR2 (N3112, N3101, N16);
buf BUF1 (N3113, N3108);
nor NOR2 (N3114, N3111, N508);
nand NAND2 (N3115, N3092, N3018);
and AND4 (N3116, N3105, N289, N1750, N2714);
nand NAND3 (N3117, N3106, N2734, N1960);
buf BUF1 (N3118, N3113);
nor NOR3 (N3119, N3110, N2905, N2800);
buf BUF1 (N3120, N3104);
nor NOR3 (N3121, N3114, N864, N855);
buf BUF1 (N3122, N3112);
not NOT1 (N3123, N3117);
nor NOR3 (N3124, N3118, N1029, N2977);
xor XOR2 (N3125, N3120, N687);
not NOT1 (N3126, N3125);
nand NAND4 (N3127, N3089, N2298, N2749, N3078);
nor NOR3 (N3128, N3123, N2068, N1197);
nor NOR3 (N3129, N3115, N2261, N1570);
nor NOR2 (N3130, N3126, N977);
nand NAND2 (N3131, N3119, N2471);
buf BUF1 (N3132, N3109);
not NOT1 (N3133, N3130);
and AND2 (N3134, N3127, N163);
nand NAND2 (N3135, N3121, N2636);
nand NAND3 (N3136, N3128, N1944, N1201);
nor NOR2 (N3137, N3129, N940);
not NOT1 (N3138, N3132);
xor XOR2 (N3139, N3131, N3039);
and AND3 (N3140, N3133, N2645, N947);
buf BUF1 (N3141, N3136);
buf BUF1 (N3142, N3137);
or OR2 (N3143, N3122, N1305);
and AND2 (N3144, N3124, N35);
buf BUF1 (N3145, N3140);
xor XOR2 (N3146, N3141, N1472);
not NOT1 (N3147, N3143);
xor XOR2 (N3148, N3116, N1956);
or OR4 (N3149, N3135, N1549, N2805, N1943);
nor NOR4 (N3150, N3146, N1917, N1081, N2890);
nor NOR2 (N3151, N3142, N1434);
or OR4 (N3152, N3138, N2931, N1834, N2532);
nand NAND4 (N3153, N3139, N222, N1694, N1987);
and AND2 (N3154, N3149, N1627);
or OR3 (N3155, N3144, N1248, N3071);
nand NAND4 (N3156, N3155, N775, N2938, N698);
and AND2 (N3157, N3154, N2042);
nor NOR2 (N3158, N3153, N1642);
buf BUF1 (N3159, N3147);
nand NAND2 (N3160, N3151, N309);
xor XOR2 (N3161, N3156, N338);
nand NAND3 (N3162, N3145, N1248, N3045);
nor NOR3 (N3163, N3158, N2708, N2195);
xor XOR2 (N3164, N3152, N555);
or OR2 (N3165, N3134, N2413);
or OR2 (N3166, N3163, N2873);
nor NOR4 (N3167, N3161, N1893, N2412, N698);
buf BUF1 (N3168, N3165);
nand NAND2 (N3169, N3166, N1807);
not NOT1 (N3170, N3159);
and AND4 (N3171, N3169, N319, N2236, N1160);
or OR3 (N3172, N3150, N1521, N375);
or OR3 (N3173, N3157, N3158, N2215);
and AND3 (N3174, N3162, N1770, N423);
not NOT1 (N3175, N3160);
and AND4 (N3176, N3168, N1562, N1306, N146);
and AND2 (N3177, N3175, N1714);
or OR3 (N3178, N3177, N157, N1025);
nor NOR2 (N3179, N3170, N3137);
or OR3 (N3180, N3167, N1291, N2376);
and AND4 (N3181, N3179, N2593, N96, N1716);
xor XOR2 (N3182, N3164, N1815);
not NOT1 (N3183, N3178);
or OR3 (N3184, N3181, N2238, N1129);
xor XOR2 (N3185, N3184, N2336);
and AND4 (N3186, N3148, N656, N1765, N1569);
buf BUF1 (N3187, N3185);
or OR4 (N3188, N3180, N1640, N2105, N2607);
not NOT1 (N3189, N3182);
nand NAND3 (N3190, N3188, N1964, N673);
nand NAND2 (N3191, N3173, N353);
not NOT1 (N3192, N3191);
buf BUF1 (N3193, N3172);
nor NOR3 (N3194, N3192, N962, N1568);
xor XOR2 (N3195, N3176, N1907);
not NOT1 (N3196, N3195);
nor NOR4 (N3197, N3196, N2166, N628, N1564);
and AND3 (N3198, N3190, N1373, N443);
or OR3 (N3199, N3183, N2764, N2662);
nand NAND3 (N3200, N3186, N37, N2787);
not NOT1 (N3201, N3187);
not NOT1 (N3202, N3198);
not NOT1 (N3203, N3193);
xor XOR2 (N3204, N3171, N352);
xor XOR2 (N3205, N3200, N1327);
buf BUF1 (N3206, N3202);
nor NOR4 (N3207, N3194, N1759, N432, N2988);
or OR2 (N3208, N3204, N923);
or OR4 (N3209, N3206, N2285, N2388, N2781);
nand NAND4 (N3210, N3205, N2009, N2084, N2324);
or OR2 (N3211, N3189, N2948);
xor XOR2 (N3212, N3203, N1912);
or OR2 (N3213, N3199, N333);
and AND3 (N3214, N3197, N1027, N2654);
nor NOR4 (N3215, N3212, N1827, N1910, N1353);
nand NAND3 (N3216, N3209, N639, N2475);
and AND3 (N3217, N3207, N42, N2663);
nor NOR3 (N3218, N3201, N946, N302);
xor XOR2 (N3219, N3213, N228);
or OR4 (N3220, N3214, N508, N1323, N606);
nor NOR3 (N3221, N3211, N3027, N1523);
buf BUF1 (N3222, N3218);
or OR2 (N3223, N3217, N2998);
nor NOR3 (N3224, N3210, N1554, N698);
buf BUF1 (N3225, N3219);
buf BUF1 (N3226, N3174);
not NOT1 (N3227, N3223);
or OR3 (N3228, N3215, N2271, N2320);
or OR3 (N3229, N3222, N2687, N1358);
nand NAND3 (N3230, N3226, N62, N2243);
buf BUF1 (N3231, N3229);
and AND3 (N3232, N3220, N1567, N1133);
buf BUF1 (N3233, N3232);
buf BUF1 (N3234, N3231);
nand NAND4 (N3235, N3234, N490, N2049, N93);
and AND4 (N3236, N3230, N2721, N1774, N2366);
not NOT1 (N3237, N3225);
not NOT1 (N3238, N3227);
nor NOR3 (N3239, N3237, N1456, N25);
nor NOR2 (N3240, N3216, N1991);
nand NAND2 (N3241, N3224, N708);
buf BUF1 (N3242, N3236);
buf BUF1 (N3243, N3228);
xor XOR2 (N3244, N3235, N2929);
and AND3 (N3245, N3241, N336, N1768);
nor NOR3 (N3246, N3208, N141, N2991);
xor XOR2 (N3247, N3245, N2711);
or OR2 (N3248, N3242, N355);
not NOT1 (N3249, N3244);
nor NOR3 (N3250, N3247, N1373, N148);
not NOT1 (N3251, N3239);
nor NOR3 (N3252, N3233, N2891, N606);
or OR2 (N3253, N3248, N1550);
not NOT1 (N3254, N3246);
or OR4 (N3255, N3250, N2781, N1396, N788);
buf BUF1 (N3256, N3255);
nor NOR2 (N3257, N3221, N653);
and AND4 (N3258, N3257, N569, N2814, N2636);
nor NOR3 (N3259, N3253, N2701, N972);
not NOT1 (N3260, N3251);
nand NAND4 (N3261, N3249, N283, N3215, N3153);
xor XOR2 (N3262, N3240, N576);
buf BUF1 (N3263, N3260);
nor NOR2 (N3264, N3238, N900);
buf BUF1 (N3265, N3243);
and AND3 (N3266, N3254, N1192, N1415);
xor XOR2 (N3267, N3261, N590);
and AND4 (N3268, N3262, N2734, N614, N1576);
not NOT1 (N3269, N3265);
not NOT1 (N3270, N3252);
or OR2 (N3271, N3264, N1305);
buf BUF1 (N3272, N3269);
or OR4 (N3273, N3256, N2711, N2530, N531);
xor XOR2 (N3274, N3272, N1546);
not NOT1 (N3275, N3259);
nor NOR3 (N3276, N3263, N2295, N596);
nor NOR2 (N3277, N3271, N993);
buf BUF1 (N3278, N3273);
xor XOR2 (N3279, N3275, N1809);
and AND2 (N3280, N3279, N2447);
and AND4 (N3281, N3270, N2429, N1213, N1892);
and AND3 (N3282, N3268, N894, N1569);
xor XOR2 (N3283, N3277, N2459);
and AND2 (N3284, N3281, N1737);
buf BUF1 (N3285, N3283);
nand NAND3 (N3286, N3284, N1136, N938);
buf BUF1 (N3287, N3286);
nand NAND3 (N3288, N3285, N596, N1597);
buf BUF1 (N3289, N3267);
not NOT1 (N3290, N3278);
and AND4 (N3291, N3290, N2077, N1720, N1964);
nor NOR3 (N3292, N3288, N812, N922);
not NOT1 (N3293, N3266);
buf BUF1 (N3294, N3293);
nor NOR3 (N3295, N3287, N2163, N2899);
xor XOR2 (N3296, N3274, N997);
nand NAND2 (N3297, N3292, N2429);
buf BUF1 (N3298, N3296);
not NOT1 (N3299, N3282);
not NOT1 (N3300, N3291);
nor NOR4 (N3301, N3295, N724, N837, N1978);
buf BUF1 (N3302, N3301);
xor XOR2 (N3303, N3258, N1207);
not NOT1 (N3304, N3299);
and AND3 (N3305, N3298, N1932, N384);
xor XOR2 (N3306, N3304, N360);
or OR4 (N3307, N3306, N2709, N3135, N563);
xor XOR2 (N3308, N3297, N1615);
and AND2 (N3309, N3303, N2945);
xor XOR2 (N3310, N3276, N2514);
buf BUF1 (N3311, N3280);
or OR4 (N3312, N3311, N2873, N1158, N180);
nand NAND4 (N3313, N3312, N2814, N2310, N788);
not NOT1 (N3314, N3310);
and AND3 (N3315, N3305, N1213, N2661);
buf BUF1 (N3316, N3294);
or OR3 (N3317, N3316, N350, N537);
nor NOR4 (N3318, N3300, N504, N288, N2640);
not NOT1 (N3319, N3315);
nor NOR2 (N3320, N3308, N3264);
xor XOR2 (N3321, N3289, N1566);
nor NOR2 (N3322, N3309, N892);
nand NAND3 (N3323, N3317, N2895, N1085);
xor XOR2 (N3324, N3307, N698);
buf BUF1 (N3325, N3314);
or OR2 (N3326, N3323, N1588);
nor NOR3 (N3327, N3321, N1196, N525);
not NOT1 (N3328, N3320);
not NOT1 (N3329, N3324);
buf BUF1 (N3330, N3318);
nand NAND3 (N3331, N3329, N130, N305);
buf BUF1 (N3332, N3319);
nand NAND3 (N3333, N3313, N3237, N997);
and AND2 (N3334, N3332, N3314);
buf BUF1 (N3335, N3325);
or OR2 (N3336, N3322, N2690);
nand NAND2 (N3337, N3335, N1717);
not NOT1 (N3338, N3326);
not NOT1 (N3339, N3336);
xor XOR2 (N3340, N3331, N2661);
and AND3 (N3341, N3340, N3296, N518);
xor XOR2 (N3342, N3334, N1238);
nor NOR4 (N3343, N3333, N896, N2644, N260);
nand NAND3 (N3344, N3337, N2719, N1780);
not NOT1 (N3345, N3338);
and AND2 (N3346, N3302, N2039);
nand NAND3 (N3347, N3339, N918, N3276);
and AND3 (N3348, N3343, N3251, N616);
not NOT1 (N3349, N3327);
or OR2 (N3350, N3328, N1642);
nor NOR2 (N3351, N3350, N757);
and AND3 (N3352, N3351, N894, N1458);
buf BUF1 (N3353, N3346);
nor NOR2 (N3354, N3349, N1190);
not NOT1 (N3355, N3341);
and AND3 (N3356, N3348, N3211, N3271);
and AND4 (N3357, N3355, N2210, N3169, N2659);
nand NAND4 (N3358, N3352, N2776, N605, N959);
nand NAND4 (N3359, N3342, N108, N2960, N2867);
nor NOR3 (N3360, N3357, N2175, N2391);
not NOT1 (N3361, N3345);
nand NAND2 (N3362, N3358, N2665);
xor XOR2 (N3363, N3362, N2885);
buf BUF1 (N3364, N3344);
not NOT1 (N3365, N3360);
nor NOR3 (N3366, N3353, N234, N2725);
not NOT1 (N3367, N3354);
xor XOR2 (N3368, N3361, N336);
or OR2 (N3369, N3367, N947);
and AND3 (N3370, N3347, N2734, N2585);
nor NOR4 (N3371, N3369, N1005, N328, N37);
and AND3 (N3372, N3330, N956, N2777);
not NOT1 (N3373, N3365);
or OR2 (N3374, N3370, N3212);
nand NAND4 (N3375, N3366, N5, N930, N308);
not NOT1 (N3376, N3374);
nand NAND3 (N3377, N3376, N436, N3100);
nor NOR4 (N3378, N3373, N2788, N123, N1371);
nand NAND3 (N3379, N3363, N469, N47);
nor NOR4 (N3380, N3359, N2323, N3017, N1824);
nor NOR3 (N3381, N3377, N2623, N741);
xor XOR2 (N3382, N3356, N1189);
nor NOR2 (N3383, N3381, N1083);
and AND3 (N3384, N3380, N638, N1732);
xor XOR2 (N3385, N3384, N448);
nor NOR3 (N3386, N3383, N1146, N2163);
not NOT1 (N3387, N3379);
not NOT1 (N3388, N3371);
nor NOR4 (N3389, N3386, N1592, N1918, N1063);
xor XOR2 (N3390, N3387, N3201);
nor NOR2 (N3391, N3388, N1456);
nand NAND4 (N3392, N3382, N1301, N1305, N2420);
not NOT1 (N3393, N3364);
not NOT1 (N3394, N3390);
nand NAND3 (N3395, N3378, N703, N879);
not NOT1 (N3396, N3389);
or OR3 (N3397, N3393, N134, N2998);
xor XOR2 (N3398, N3395, N2589);
nand NAND4 (N3399, N3394, N3266, N617, N1741);
nand NAND2 (N3400, N3397, N2125);
not NOT1 (N3401, N3399);
nand NAND4 (N3402, N3391, N2264, N1647, N1229);
not NOT1 (N3403, N3372);
not NOT1 (N3404, N3392);
and AND4 (N3405, N3398, N792, N1462, N2681);
xor XOR2 (N3406, N3400, N68);
nand NAND4 (N3407, N3401, N3207, N465, N1699);
nand NAND3 (N3408, N3406, N2555, N1883);
nor NOR2 (N3409, N3407, N2699);
nand NAND2 (N3410, N3403, N696);
xor XOR2 (N3411, N3385, N779);
xor XOR2 (N3412, N3409, N302);
or OR2 (N3413, N3412, N1743);
and AND3 (N3414, N3375, N2040, N3255);
not NOT1 (N3415, N3396);
xor XOR2 (N3416, N3410, N1700);
and AND4 (N3417, N3413, N2276, N1592, N1503);
buf BUF1 (N3418, N3408);
or OR3 (N3419, N3418, N2914, N858);
and AND2 (N3420, N3417, N2157);
xor XOR2 (N3421, N3402, N1762);
buf BUF1 (N3422, N3405);
xor XOR2 (N3423, N3416, N2671);
or OR4 (N3424, N3422, N3305, N2441, N2874);
nor NOR4 (N3425, N3423, N1635, N903, N3344);
or OR3 (N3426, N3411, N2161, N2480);
xor XOR2 (N3427, N3425, N289);
buf BUF1 (N3428, N3421);
or OR3 (N3429, N3419, N1871, N3241);
and AND2 (N3430, N3404, N3195);
and AND4 (N3431, N3415, N2625, N89, N2951);
not NOT1 (N3432, N3426);
xor XOR2 (N3433, N3368, N3301);
buf BUF1 (N3434, N3433);
not NOT1 (N3435, N3414);
not NOT1 (N3436, N3430);
nor NOR4 (N3437, N3427, N2102, N1374, N3381);
buf BUF1 (N3438, N3436);
buf BUF1 (N3439, N3435);
nand NAND3 (N3440, N3434, N2678, N1032);
nor NOR3 (N3441, N3420, N3043, N1098);
nor NOR3 (N3442, N3429, N493, N1454);
nor NOR2 (N3443, N3439, N2799);
not NOT1 (N3444, N3441);
not NOT1 (N3445, N3424);
not NOT1 (N3446, N3431);
nand NAND4 (N3447, N3438, N1990, N2293, N741);
buf BUF1 (N3448, N3437);
and AND2 (N3449, N3448, N1750);
buf BUF1 (N3450, N3442);
buf BUF1 (N3451, N3428);
or OR3 (N3452, N3447, N505, N1436);
and AND2 (N3453, N3451, N2941);
or OR4 (N3454, N3444, N566, N2755, N1663);
or OR4 (N3455, N3454, N704, N1557, N1485);
xor XOR2 (N3456, N3455, N2253);
nand NAND2 (N3457, N3452, N222);
and AND4 (N3458, N3432, N1971, N486, N1086);
not NOT1 (N3459, N3449);
xor XOR2 (N3460, N3458, N3055);
not NOT1 (N3461, N3443);
and AND3 (N3462, N3440, N333, N467);
not NOT1 (N3463, N3460);
xor XOR2 (N3464, N3456, N2185);
not NOT1 (N3465, N3445);
and AND4 (N3466, N3462, N2072, N1967, N802);
buf BUF1 (N3467, N3457);
nand NAND3 (N3468, N3446, N526, N1881);
buf BUF1 (N3469, N3461);
or OR2 (N3470, N3450, N764);
or OR2 (N3471, N3459, N176);
buf BUF1 (N3472, N3470);
xor XOR2 (N3473, N3467, N2754);
buf BUF1 (N3474, N3472);
buf BUF1 (N3475, N3465);
nand NAND4 (N3476, N3475, N219, N837, N659);
buf BUF1 (N3477, N3466);
nand NAND4 (N3478, N3468, N558, N2797, N549);
nand NAND2 (N3479, N3478, N2438);
buf BUF1 (N3480, N3469);
nand NAND2 (N3481, N3464, N592);
or OR2 (N3482, N3474, N2930);
buf BUF1 (N3483, N3471);
not NOT1 (N3484, N3481);
or OR3 (N3485, N3453, N1372, N1767);
nor NOR2 (N3486, N3477, N640);
buf BUF1 (N3487, N3484);
and AND4 (N3488, N3479, N3414, N1672, N3472);
and AND3 (N3489, N3483, N1144, N1234);
or OR2 (N3490, N3488, N3039);
or OR3 (N3491, N3473, N1725, N523);
buf BUF1 (N3492, N3485);
not NOT1 (N3493, N3490);
or OR3 (N3494, N3476, N567, N3362);
nor NOR2 (N3495, N3487, N1525);
nor NOR2 (N3496, N3463, N1264);
and AND2 (N3497, N3493, N1037);
buf BUF1 (N3498, N3497);
and AND2 (N3499, N3494, N2052);
and AND4 (N3500, N3496, N198, N1524, N2127);
nor NOR4 (N3501, N3500, N1583, N68, N1062);
and AND4 (N3502, N3495, N3331, N258, N536);
and AND2 (N3503, N3480, N3142);
or OR3 (N3504, N3482, N2221, N244);
not NOT1 (N3505, N3503);
nand NAND2 (N3506, N3492, N996);
and AND3 (N3507, N3489, N1086, N395);
buf BUF1 (N3508, N3498);
and AND2 (N3509, N3507, N2495);
nand NAND3 (N3510, N3508, N1082, N2646);
or OR3 (N3511, N3491, N1742, N3174);
xor XOR2 (N3512, N3486, N87);
not NOT1 (N3513, N3506);
nor NOR4 (N3514, N3504, N91, N3280, N2681);
nand NAND2 (N3515, N3505, N571);
buf BUF1 (N3516, N3512);
nor NOR3 (N3517, N3509, N2529, N1662);
nor NOR3 (N3518, N3513, N1206, N137);
nor NOR4 (N3519, N3518, N2763, N1905, N1018);
nor NOR2 (N3520, N3516, N3051);
and AND2 (N3521, N3515, N1858);
or OR3 (N3522, N3520, N3286, N3411);
not NOT1 (N3523, N3517);
buf BUF1 (N3524, N3501);
nor NOR2 (N3525, N3511, N2863);
or OR2 (N3526, N3519, N968);
not NOT1 (N3527, N3524);
buf BUF1 (N3528, N3527);
and AND3 (N3529, N3514, N923, N2947);
nor NOR4 (N3530, N3526, N1604, N984, N918);
buf BUF1 (N3531, N3525);
buf BUF1 (N3532, N3530);
or OR2 (N3533, N3528, N3268);
buf BUF1 (N3534, N3523);
and AND4 (N3535, N3510, N631, N513, N2117);
nor NOR2 (N3536, N3532, N611);
buf BUF1 (N3537, N3531);
xor XOR2 (N3538, N3502, N863);
buf BUF1 (N3539, N3499);
nor NOR2 (N3540, N3537, N1905);
xor XOR2 (N3541, N3533, N952);
or OR4 (N3542, N3539, N2167, N2475, N1713);
not NOT1 (N3543, N3542);
or OR3 (N3544, N3534, N310, N1479);
nand NAND3 (N3545, N3535, N1700, N1068);
xor XOR2 (N3546, N3521, N1756);
nand NAND2 (N3547, N3541, N1354);
or OR3 (N3548, N3522, N1174, N3136);
or OR4 (N3549, N3543, N3038, N461, N3542);
nor NOR2 (N3550, N3536, N1243);
xor XOR2 (N3551, N3538, N2369);
or OR2 (N3552, N3545, N2902);
nand NAND2 (N3553, N3548, N2709);
or OR2 (N3554, N3552, N1677);
nand NAND2 (N3555, N3553, N1297);
nand NAND4 (N3556, N3546, N273, N1351, N1263);
or OR3 (N3557, N3529, N793, N174);
and AND3 (N3558, N3554, N1223, N1016);
nand NAND4 (N3559, N3550, N3414, N1481, N1187);
not NOT1 (N3560, N3549);
nand NAND4 (N3561, N3555, N3511, N1687, N3004);
or OR4 (N3562, N3556, N3393, N473, N2252);
not NOT1 (N3563, N3547);
not NOT1 (N3564, N3560);
and AND2 (N3565, N3540, N1454);
nand NAND4 (N3566, N3561, N395, N658, N772);
or OR3 (N3567, N3557, N3131, N3025);
or OR3 (N3568, N3558, N2825, N1973);
and AND3 (N3569, N3564, N2536, N2423);
nand NAND2 (N3570, N3567, N533);
buf BUF1 (N3571, N3570);
or OR3 (N3572, N3568, N2883, N2276);
nand NAND2 (N3573, N3572, N1882);
and AND4 (N3574, N3562, N3042, N379, N1089);
or OR3 (N3575, N3565, N3335, N1647);
buf BUF1 (N3576, N3551);
and AND3 (N3577, N3573, N2498, N1382);
nor NOR2 (N3578, N3566, N1252);
nand NAND4 (N3579, N3576, N335, N1431, N3362);
xor XOR2 (N3580, N3569, N3132);
not NOT1 (N3581, N3578);
buf BUF1 (N3582, N3559);
buf BUF1 (N3583, N3577);
or OR3 (N3584, N3544, N1675, N3426);
nor NOR4 (N3585, N3581, N150, N2112, N1483);
buf BUF1 (N3586, N3584);
not NOT1 (N3587, N3585);
and AND3 (N3588, N3586, N2716, N2180);
not NOT1 (N3589, N3582);
not NOT1 (N3590, N3579);
buf BUF1 (N3591, N3580);
xor XOR2 (N3592, N3574, N1532);
and AND3 (N3593, N3571, N3182, N1171);
buf BUF1 (N3594, N3592);
nand NAND4 (N3595, N3588, N1080, N380, N3264);
nand NAND2 (N3596, N3589, N3256);
xor XOR2 (N3597, N3596, N1224);
buf BUF1 (N3598, N3591);
nor NOR4 (N3599, N3575, N949, N3041, N1867);
buf BUF1 (N3600, N3594);
buf BUF1 (N3601, N3593);
or OR2 (N3602, N3587, N2707);
nor NOR2 (N3603, N3590, N3549);
buf BUF1 (N3604, N3600);
nor NOR4 (N3605, N3595, N2009, N2334, N2156);
nand NAND3 (N3606, N3599, N2966, N2832);
nand NAND4 (N3607, N3603, N2375, N2880, N1054);
and AND2 (N3608, N3606, N34);
nor NOR3 (N3609, N3563, N496, N2373);
buf BUF1 (N3610, N3607);
or OR3 (N3611, N3597, N1633, N78);
and AND2 (N3612, N3583, N3229);
nor NOR4 (N3613, N3608, N489, N3178, N3104);
or OR3 (N3614, N3612, N648, N1041);
nor NOR2 (N3615, N3613, N1566);
or OR3 (N3616, N3615, N179, N1188);
or OR2 (N3617, N3601, N199);
nor NOR3 (N3618, N3605, N1380, N244);
not NOT1 (N3619, N3618);
or OR4 (N3620, N3616, N205, N3133, N559);
not NOT1 (N3621, N3617);
nor NOR4 (N3622, N3609, N1059, N715, N1514);
buf BUF1 (N3623, N3619);
xor XOR2 (N3624, N3602, N2404);
nor NOR3 (N3625, N3623, N1801, N892);
or OR2 (N3626, N3624, N3561);
nand NAND3 (N3627, N3614, N2985, N3547);
buf BUF1 (N3628, N3610);
or OR3 (N3629, N3626, N1914, N130);
xor XOR2 (N3630, N3611, N115);
nor NOR2 (N3631, N3627, N2675);
or OR3 (N3632, N3630, N615, N1617);
not NOT1 (N3633, N3629);
xor XOR2 (N3634, N3598, N2972);
not NOT1 (N3635, N3628);
and AND4 (N3636, N3620, N22, N2239, N563);
or OR2 (N3637, N3631, N2188);
buf BUF1 (N3638, N3621);
not NOT1 (N3639, N3632);
xor XOR2 (N3640, N3622, N911);
nand NAND4 (N3641, N3604, N539, N2830, N1485);
and AND3 (N3642, N3636, N631, N419);
and AND4 (N3643, N3635, N3470, N3589, N1776);
or OR2 (N3644, N3637, N174);
or OR4 (N3645, N3641, N1127, N2428, N1708);
xor XOR2 (N3646, N3625, N1194);
xor XOR2 (N3647, N3646, N910);
or OR4 (N3648, N3633, N2672, N2486, N2327);
not NOT1 (N3649, N3643);
not NOT1 (N3650, N3642);
not NOT1 (N3651, N3648);
and AND2 (N3652, N3650, N3589);
nand NAND3 (N3653, N3640, N446, N3110);
xor XOR2 (N3654, N3647, N83);
and AND3 (N3655, N3634, N1482, N1589);
buf BUF1 (N3656, N3649);
nor NOR2 (N3657, N3655, N665);
nor NOR2 (N3658, N3644, N3115);
nand NAND2 (N3659, N3657, N825);
buf BUF1 (N3660, N3656);
nand NAND3 (N3661, N3658, N1465, N2376);
nor NOR3 (N3662, N3661, N1553, N363);
and AND3 (N3663, N3653, N1786, N2833);
nand NAND3 (N3664, N3638, N866, N1692);
or OR4 (N3665, N3654, N3455, N2788, N3379);
buf BUF1 (N3666, N3639);
nand NAND3 (N3667, N3659, N1385, N2358);
nor NOR2 (N3668, N3667, N3494);
nor NOR2 (N3669, N3665, N2493);
and AND3 (N3670, N3668, N1272, N616);
nand NAND2 (N3671, N3666, N2428);
and AND4 (N3672, N3660, N1744, N2367, N1382);
xor XOR2 (N3673, N3669, N2885);
and AND2 (N3674, N3662, N1111);
and AND2 (N3675, N3652, N453);
not NOT1 (N3676, N3664);
not NOT1 (N3677, N3672);
or OR3 (N3678, N3676, N2755, N1738);
nor NOR3 (N3679, N3651, N2761, N2610);
nand NAND4 (N3680, N3679, N495, N3625, N148);
not NOT1 (N3681, N3678);
buf BUF1 (N3682, N3671);
or OR4 (N3683, N3645, N1012, N1470, N3186);
xor XOR2 (N3684, N3683, N1311);
or OR2 (N3685, N3680, N3301);
not NOT1 (N3686, N3682);
nand NAND2 (N3687, N3685, N2479);
buf BUF1 (N3688, N3670);
buf BUF1 (N3689, N3675);
xor XOR2 (N3690, N3673, N3309);
buf BUF1 (N3691, N3663);
or OR4 (N3692, N3687, N1839, N130, N1812);
nand NAND4 (N3693, N3686, N2433, N3545, N2972);
nand NAND4 (N3694, N3688, N246, N1246, N1347);
xor XOR2 (N3695, N3689, N2386);
and AND4 (N3696, N3684, N2423, N2134, N1108);
nand NAND3 (N3697, N3696, N1955, N966);
nand NAND4 (N3698, N3691, N1802, N893, N1457);
or OR3 (N3699, N3690, N1076, N2761);
xor XOR2 (N3700, N3695, N3099);
buf BUF1 (N3701, N3700);
xor XOR2 (N3702, N3674, N1765);
buf BUF1 (N3703, N3702);
nor NOR2 (N3704, N3701, N3528);
or OR2 (N3705, N3698, N2426);
xor XOR2 (N3706, N3699, N3489);
not NOT1 (N3707, N3705);
nand NAND2 (N3708, N3692, N203);
or OR4 (N3709, N3707, N2589, N1918, N3224);
not NOT1 (N3710, N3704);
nor NOR3 (N3711, N3708, N1746, N685);
nand NAND4 (N3712, N3706, N1788, N1429, N3662);
buf BUF1 (N3713, N3711);
nand NAND2 (N3714, N3694, N2316);
buf BUF1 (N3715, N3703);
nor NOR4 (N3716, N3712, N1404, N3115, N1919);
nor NOR4 (N3717, N3713, N359, N2401, N1976);
buf BUF1 (N3718, N3677);
and AND2 (N3719, N3718, N713);
buf BUF1 (N3720, N3715);
not NOT1 (N3721, N3681);
and AND2 (N3722, N3717, N402);
nor NOR2 (N3723, N3722, N206);
nor NOR2 (N3724, N3709, N3137);
or OR2 (N3725, N3719, N506);
buf BUF1 (N3726, N3724);
nor NOR3 (N3727, N3697, N3434, N3516);
and AND2 (N3728, N3710, N3601);
not NOT1 (N3729, N3714);
buf BUF1 (N3730, N3725);
nand NAND4 (N3731, N3726, N770, N813, N1811);
nor NOR2 (N3732, N3716, N1894);
not NOT1 (N3733, N3732);
or OR4 (N3734, N3728, N187, N201, N285);
not NOT1 (N3735, N3723);
xor XOR2 (N3736, N3721, N791);
nand NAND2 (N3737, N3730, N3493);
and AND2 (N3738, N3720, N2691);
xor XOR2 (N3739, N3738, N1756);
nor NOR4 (N3740, N3734, N3552, N974, N510);
nor NOR4 (N3741, N3729, N2149, N3382, N751);
nand NAND2 (N3742, N3739, N2232);
nor NOR2 (N3743, N3693, N2555);
buf BUF1 (N3744, N3736);
or OR3 (N3745, N3737, N2385, N1311);
nand NAND2 (N3746, N3742, N969);
or OR4 (N3747, N3733, N3709, N2209, N1893);
and AND2 (N3748, N3746, N3120);
and AND3 (N3749, N3743, N3424, N311);
or OR4 (N3750, N3735, N3176, N301, N1645);
nand NAND4 (N3751, N3750, N1591, N1372, N3211);
not NOT1 (N3752, N3745);
nand NAND2 (N3753, N3747, N2976);
xor XOR2 (N3754, N3751, N1970);
nand NAND4 (N3755, N3740, N669, N1990, N2905);
xor XOR2 (N3756, N3744, N606);
nor NOR3 (N3757, N3754, N1650, N2344);
or OR2 (N3758, N3749, N164);
nand NAND3 (N3759, N3758, N613, N2093);
xor XOR2 (N3760, N3759, N365);
or OR4 (N3761, N3727, N3343, N1634, N1790);
nor NOR2 (N3762, N3752, N406);
and AND3 (N3763, N3753, N2344, N1082);
not NOT1 (N3764, N3755);
or OR2 (N3765, N3760, N195);
nor NOR4 (N3766, N3748, N3144, N789, N2337);
nand NAND2 (N3767, N3757, N2489);
or OR4 (N3768, N3767, N2438, N259, N121);
nor NOR2 (N3769, N3768, N991);
not NOT1 (N3770, N3763);
and AND2 (N3771, N3761, N249);
and AND3 (N3772, N3764, N1027, N1620);
xor XOR2 (N3773, N3741, N373);
or OR4 (N3774, N3756, N1405, N1141, N1771);
nor NOR2 (N3775, N3762, N3603);
not NOT1 (N3776, N3770);
xor XOR2 (N3777, N3765, N171);
and AND3 (N3778, N3772, N1332, N587);
nor NOR3 (N3779, N3778, N1350, N7);
buf BUF1 (N3780, N3769);
not NOT1 (N3781, N3774);
nor NOR2 (N3782, N3766, N2771);
not NOT1 (N3783, N3780);
nand NAND4 (N3784, N3781, N3751, N2164, N2528);
xor XOR2 (N3785, N3784, N843);
or OR3 (N3786, N3773, N2398, N2530);
or OR2 (N3787, N3779, N782);
nor NOR3 (N3788, N3771, N111, N1047);
and AND2 (N3789, N3787, N1901);
nand NAND4 (N3790, N3789, N3406, N3483, N1923);
nor NOR2 (N3791, N3783, N1576);
or OR4 (N3792, N3788, N1388, N662, N2635);
xor XOR2 (N3793, N3790, N3789);
nand NAND2 (N3794, N3782, N2693);
not NOT1 (N3795, N3793);
buf BUF1 (N3796, N3785);
nand NAND3 (N3797, N3777, N2791, N1841);
not NOT1 (N3798, N3796);
nand NAND3 (N3799, N3795, N1312, N755);
buf BUF1 (N3800, N3786);
buf BUF1 (N3801, N3799);
buf BUF1 (N3802, N3776);
or OR3 (N3803, N3801, N1604, N2314);
nand NAND2 (N3804, N3803, N3687);
and AND2 (N3805, N3797, N246);
xor XOR2 (N3806, N3791, N222);
or OR3 (N3807, N3731, N1705, N3583);
and AND3 (N3808, N3798, N2286, N129);
nor NOR3 (N3809, N3800, N2527, N3799);
and AND4 (N3810, N3805, N3365, N390, N3210);
nor NOR3 (N3811, N3808, N1909, N473);
nor NOR2 (N3812, N3804, N557);
and AND4 (N3813, N3807, N959, N2969, N3431);
and AND2 (N3814, N3792, N454);
not NOT1 (N3815, N3806);
not NOT1 (N3816, N3811);
nor NOR3 (N3817, N3812, N2431, N1242);
nand NAND4 (N3818, N3816, N261, N2568, N2015);
or OR2 (N3819, N3794, N532);
nand NAND2 (N3820, N3814, N441);
buf BUF1 (N3821, N3820);
buf BUF1 (N3822, N3810);
xor XOR2 (N3823, N3775, N3112);
nand NAND4 (N3824, N3817, N2087, N2770, N1294);
and AND3 (N3825, N3822, N3062, N3677);
nor NOR2 (N3826, N3825, N2354);
nor NOR3 (N3827, N3821, N3169, N2395);
not NOT1 (N3828, N3819);
and AND3 (N3829, N3813, N1779, N864);
xor XOR2 (N3830, N3815, N3386);
xor XOR2 (N3831, N3823, N3264);
nand NAND4 (N3832, N3827, N2237, N3728, N438);
and AND4 (N3833, N3824, N3279, N751, N3359);
nor NOR2 (N3834, N3826, N2711);
or OR2 (N3835, N3828, N811);
nor NOR3 (N3836, N3830, N2525, N74);
xor XOR2 (N3837, N3833, N465);
not NOT1 (N3838, N3835);
or OR2 (N3839, N3818, N1438);
buf BUF1 (N3840, N3832);
not NOT1 (N3841, N3839);
buf BUF1 (N3842, N3837);
not NOT1 (N3843, N3831);
or OR2 (N3844, N3809, N3207);
nand NAND3 (N3845, N3840, N2314, N2688);
and AND4 (N3846, N3843, N1584, N2725, N3793);
buf BUF1 (N3847, N3802);
and AND2 (N3848, N3841, N3202);
and AND2 (N3849, N3834, N1045);
not NOT1 (N3850, N3844);
or OR2 (N3851, N3845, N947);
not NOT1 (N3852, N3849);
and AND4 (N3853, N3850, N1062, N2121, N3125);
nand NAND4 (N3854, N3829, N2504, N2783, N3176);
or OR3 (N3855, N3848, N2815, N136);
and AND4 (N3856, N3854, N1340, N1882, N1162);
nand NAND2 (N3857, N3855, N2967);
xor XOR2 (N3858, N3851, N1087);
or OR4 (N3859, N3838, N1898, N1403, N449);
xor XOR2 (N3860, N3836, N3313);
and AND3 (N3861, N3842, N1489, N2433);
not NOT1 (N3862, N3857);
xor XOR2 (N3863, N3862, N1649);
nand NAND2 (N3864, N3859, N768);
not NOT1 (N3865, N3861);
nand NAND3 (N3866, N3852, N3681, N2329);
nor NOR4 (N3867, N3863, N2692, N227, N706);
nor NOR4 (N3868, N3866, N2061, N935, N94);
xor XOR2 (N3869, N3860, N2907);
not NOT1 (N3870, N3858);
nand NAND2 (N3871, N3864, N3631);
buf BUF1 (N3872, N3868);
nor NOR3 (N3873, N3853, N2109, N3558);
xor XOR2 (N3874, N3867, N1256);
buf BUF1 (N3875, N3846);
or OR4 (N3876, N3856, N2249, N2843, N3290);
or OR2 (N3877, N3865, N1881);
nor NOR3 (N3878, N3871, N1469, N3470);
buf BUF1 (N3879, N3869);
nor NOR3 (N3880, N3847, N155, N2934);
not NOT1 (N3881, N3873);
nand NAND4 (N3882, N3878, N2829, N403, N2209);
xor XOR2 (N3883, N3877, N2988);
nand NAND3 (N3884, N3876, N1370, N1318);
not NOT1 (N3885, N3882);
and AND4 (N3886, N3881, N1933, N2383, N1837);
nor NOR4 (N3887, N3884, N128, N528, N3710);
and AND4 (N3888, N3870, N3001, N2419, N2161);
nand NAND2 (N3889, N3883, N2177);
buf BUF1 (N3890, N3875);
and AND4 (N3891, N3887, N1074, N579, N1705);
nor NOR2 (N3892, N3872, N3027);
or OR2 (N3893, N3889, N1748);
or OR4 (N3894, N3880, N2950, N3851, N213);
nand NAND2 (N3895, N3891, N2654);
xor XOR2 (N3896, N3886, N1059);
or OR3 (N3897, N3892, N2607, N48);
xor XOR2 (N3898, N3896, N355);
or OR2 (N3899, N3897, N3876);
nor NOR3 (N3900, N3898, N2380, N3285);
or OR3 (N3901, N3888, N3301, N3524);
nand NAND3 (N3902, N3885, N2038, N3270);
or OR2 (N3903, N3893, N3024);
nand NAND3 (N3904, N3902, N2317, N380);
xor XOR2 (N3905, N3903, N2232);
and AND2 (N3906, N3890, N2878);
not NOT1 (N3907, N3901);
and AND3 (N3908, N3900, N277, N1367);
not NOT1 (N3909, N3906);
nand NAND3 (N3910, N3909, N997, N942);
buf BUF1 (N3911, N3910);
xor XOR2 (N3912, N3874, N1331);
xor XOR2 (N3913, N3894, N72);
and AND2 (N3914, N3907, N2135);
not NOT1 (N3915, N3895);
nand NAND3 (N3916, N3905, N912, N472);
nand NAND3 (N3917, N3904, N1601, N1492);
and AND3 (N3918, N3915, N1249, N1839);
nor NOR3 (N3919, N3908, N1551, N2352);
nor NOR2 (N3920, N3916, N8);
not NOT1 (N3921, N3879);
xor XOR2 (N3922, N3917, N1123);
xor XOR2 (N3923, N3913, N588);
and AND3 (N3924, N3919, N3540, N3494);
not NOT1 (N3925, N3911);
and AND2 (N3926, N3923, N3140);
nor NOR2 (N3927, N3914, N1502);
nand NAND2 (N3928, N3899, N373);
nor NOR2 (N3929, N3918, N3309);
xor XOR2 (N3930, N3922, N2376);
and AND2 (N3931, N3929, N920);
nor NOR4 (N3932, N3920, N22, N830, N3702);
buf BUF1 (N3933, N3927);
and AND4 (N3934, N3924, N2548, N3359, N3261);
nor NOR4 (N3935, N3921, N3847, N2633, N396);
or OR2 (N3936, N3925, N3878);
nor NOR4 (N3937, N3932, N607, N1011, N2633);
buf BUF1 (N3938, N3935);
not NOT1 (N3939, N3937);
nor NOR3 (N3940, N3931, N2845, N2733);
or OR3 (N3941, N3930, N158, N3475);
buf BUF1 (N3942, N3941);
buf BUF1 (N3943, N3912);
not NOT1 (N3944, N3940);
and AND4 (N3945, N3943, N2419, N3555, N3446);
or OR4 (N3946, N3942, N466, N290, N2289);
not NOT1 (N3947, N3946);
not NOT1 (N3948, N3928);
buf BUF1 (N3949, N3926);
buf BUF1 (N3950, N3948);
xor XOR2 (N3951, N3945, N2070);
nand NAND2 (N3952, N3947, N200);
xor XOR2 (N3953, N3951, N3337);
nor NOR2 (N3954, N3938, N3173);
buf BUF1 (N3955, N3933);
not NOT1 (N3956, N3939);
buf BUF1 (N3957, N3936);
not NOT1 (N3958, N3950);
buf BUF1 (N3959, N3957);
nand NAND2 (N3960, N3956, N1040);
buf BUF1 (N3961, N3934);
nor NOR2 (N3962, N3953, N1265);
and AND4 (N3963, N3960, N1135, N2899, N2680);
not NOT1 (N3964, N3961);
not NOT1 (N3965, N3952);
xor XOR2 (N3966, N3962, N3463);
nand NAND4 (N3967, N3963, N3271, N214, N2133);
nand NAND2 (N3968, N3959, N2120);
buf BUF1 (N3969, N3968);
and AND4 (N3970, N3965, N451, N3231, N2931);
buf BUF1 (N3971, N3955);
or OR3 (N3972, N3966, N672, N3435);
nand NAND4 (N3973, N3967, N1131, N78, N3897);
nand NAND3 (N3974, N3964, N3153, N1067);
xor XOR2 (N3975, N3973, N2376);
buf BUF1 (N3976, N3949);
nor NOR2 (N3977, N3972, N2760);
or OR2 (N3978, N3944, N1782);
and AND3 (N3979, N3977, N587, N2796);
nor NOR4 (N3980, N3970, N2940, N2732, N2034);
or OR2 (N3981, N3980, N2449);
nor NOR2 (N3982, N3981, N3594);
nor NOR3 (N3983, N3976, N3912, N1231);
xor XOR2 (N3984, N3971, N513);
and AND2 (N3985, N3984, N3866);
and AND4 (N3986, N3969, N3901, N1167, N2424);
nor NOR2 (N3987, N3983, N842);
xor XOR2 (N3988, N3974, N3806);
or OR4 (N3989, N3982, N3655, N2017, N2200);
nand NAND3 (N3990, N3986, N2110, N1711);
or OR3 (N3991, N3988, N1346, N3537);
and AND4 (N3992, N3978, N3207, N287, N2873);
buf BUF1 (N3993, N3979);
and AND4 (N3994, N3989, N365, N1677, N856);
buf BUF1 (N3995, N3991);
or OR2 (N3996, N3994, N3193);
and AND3 (N3997, N3975, N2028, N2890);
nor NOR4 (N3998, N3995, N2270, N3192, N573);
nand NAND3 (N3999, N3990, N2895, N537);
xor XOR2 (N4000, N3958, N1659);
nand NAND3 (N4001, N3992, N30, N2392);
not NOT1 (N4002, N3987);
nand NAND4 (N4003, N3993, N821, N3361, N3529);
nor NOR4 (N4004, N4000, N93, N2210, N676);
nand NAND4 (N4005, N3996, N3310, N558, N1670);
not NOT1 (N4006, N4002);
or OR3 (N4007, N3999, N2070, N3884);
not NOT1 (N4008, N4006);
nand NAND3 (N4009, N4004, N3683, N1706);
or OR4 (N4010, N3997, N896, N2135, N1645);
nor NOR3 (N4011, N4010, N2037, N3676);
nand NAND2 (N4012, N4009, N476);
xor XOR2 (N4013, N4003, N340);
and AND4 (N4014, N4013, N3835, N1260, N3235);
not NOT1 (N4015, N4014);
nand NAND3 (N4016, N3985, N1216, N310);
buf BUF1 (N4017, N4005);
buf BUF1 (N4018, N3954);
xor XOR2 (N4019, N4007, N3827);
not NOT1 (N4020, N4008);
not NOT1 (N4021, N3998);
and AND3 (N4022, N4017, N171, N844);
buf BUF1 (N4023, N4001);
buf BUF1 (N4024, N4015);
nor NOR3 (N4025, N4020, N393, N3183);
buf BUF1 (N4026, N4021);
buf BUF1 (N4027, N4026);
not NOT1 (N4028, N4011);
and AND2 (N4029, N4023, N3562);
not NOT1 (N4030, N4012);
and AND3 (N4031, N4029, N63, N2996);
xor XOR2 (N4032, N4022, N1856);
not NOT1 (N4033, N4018);
and AND2 (N4034, N4033, N2043);
or OR2 (N4035, N4032, N2692);
and AND4 (N4036, N4016, N3903, N802, N1662);
nor NOR3 (N4037, N4034, N943, N1688);
nor NOR2 (N4038, N4030, N2198);
nand NAND4 (N4039, N4038, N2173, N1087, N1678);
and AND4 (N4040, N4031, N828, N2156, N1777);
xor XOR2 (N4041, N4035, N3932);
xor XOR2 (N4042, N4025, N398);
xor XOR2 (N4043, N4024, N3558);
and AND4 (N4044, N4027, N3851, N2265, N2180);
not NOT1 (N4045, N4037);
buf BUF1 (N4046, N4042);
and AND4 (N4047, N4041, N645, N2391, N2189);
and AND2 (N4048, N4019, N943);
or OR4 (N4049, N4044, N2582, N489, N3288);
and AND2 (N4050, N4046, N3826);
buf BUF1 (N4051, N4045);
not NOT1 (N4052, N4040);
not NOT1 (N4053, N4028);
xor XOR2 (N4054, N4052, N1947);
and AND4 (N4055, N4047, N156, N2462, N3660);
xor XOR2 (N4056, N4036, N1458);
or OR4 (N4057, N4050, N2840, N441, N3030);
xor XOR2 (N4058, N4055, N2859);
buf BUF1 (N4059, N4058);
or OR3 (N4060, N4051, N567, N1708);
nor NOR2 (N4061, N4048, N2335);
nand NAND4 (N4062, N4061, N133, N980, N983);
nor NOR3 (N4063, N4060, N3022, N3328);
or OR2 (N4064, N4062, N2521);
xor XOR2 (N4065, N4039, N714);
nand NAND4 (N4066, N4043, N3584, N2809, N2336);
nand NAND2 (N4067, N4049, N104);
nor NOR3 (N4068, N4057, N3257, N2830);
and AND3 (N4069, N4063, N1951, N1049);
and AND3 (N4070, N4056, N3808, N1459);
and AND4 (N4071, N4067, N2938, N636, N3485);
or OR3 (N4072, N4066, N2114, N2528);
xor XOR2 (N4073, N4064, N3955);
nand NAND4 (N4074, N4059, N1970, N1812, N2701);
nand NAND4 (N4075, N4068, N3928, N3955, N3514);
not NOT1 (N4076, N4072);
xor XOR2 (N4077, N4073, N3098);
xor XOR2 (N4078, N4074, N370);
and AND2 (N4079, N4070, N3906);
buf BUF1 (N4080, N4065);
not NOT1 (N4081, N4071);
nor NOR2 (N4082, N4053, N4072);
or OR3 (N4083, N4080, N3920, N1569);
not NOT1 (N4084, N4076);
or OR3 (N4085, N4078, N2226, N1594);
xor XOR2 (N4086, N4081, N2959);
buf BUF1 (N4087, N4086);
and AND4 (N4088, N4083, N275, N820, N2207);
or OR2 (N4089, N4082, N1675);
nor NOR3 (N4090, N4054, N182, N456);
nor NOR2 (N4091, N4075, N3689);
nor NOR2 (N4092, N4084, N3975);
and AND2 (N4093, N4079, N1732);
xor XOR2 (N4094, N4093, N48);
or OR4 (N4095, N4090, N150, N1218, N3477);
nor NOR3 (N4096, N4095, N2133, N984);
buf BUF1 (N4097, N4096);
nand NAND3 (N4098, N4089, N3676, N69);
not NOT1 (N4099, N4087);
buf BUF1 (N4100, N4077);
xor XOR2 (N4101, N4088, N2803);
nor NOR3 (N4102, N4101, N3102, N1223);
nor NOR2 (N4103, N4094, N2853);
buf BUF1 (N4104, N4092);
xor XOR2 (N4105, N4091, N173);
nand NAND2 (N4106, N4097, N361);
xor XOR2 (N4107, N4102, N3174);
and AND4 (N4108, N4103, N4008, N419, N3655);
and AND3 (N4109, N4069, N1384, N55);
or OR2 (N4110, N4106, N375);
not NOT1 (N4111, N4085);
buf BUF1 (N4112, N4107);
nor NOR4 (N4113, N4108, N755, N4024, N35);
buf BUF1 (N4114, N4098);
or OR4 (N4115, N4099, N1078, N3891, N2746);
or OR3 (N4116, N4110, N4103, N116);
xor XOR2 (N4117, N4100, N224);
nand NAND3 (N4118, N4109, N3981, N969);
not NOT1 (N4119, N4116);
not NOT1 (N4120, N4112);
nand NAND3 (N4121, N4114, N3731, N3382);
nand NAND4 (N4122, N4119, N3186, N1440, N552);
or OR2 (N4123, N4117, N123);
xor XOR2 (N4124, N4115, N1205);
buf BUF1 (N4125, N4122);
xor XOR2 (N4126, N4120, N3027);
or OR4 (N4127, N4125, N3533, N2718, N2474);
nor NOR3 (N4128, N4118, N1462, N3999);
buf BUF1 (N4129, N4113);
nor NOR2 (N4130, N4123, N3731);
nand NAND4 (N4131, N4129, N4057, N2422, N4103);
nand NAND3 (N4132, N4126, N1095, N705);
or OR2 (N4133, N4127, N2099);
buf BUF1 (N4134, N4124);
buf BUF1 (N4135, N4133);
nor NOR4 (N4136, N4121, N841, N2617, N355);
or OR3 (N4137, N4135, N2785, N1262);
xor XOR2 (N4138, N4137, N467);
nand NAND4 (N4139, N4136, N2236, N1031, N2333);
and AND3 (N4140, N4128, N1447, N162);
xor XOR2 (N4141, N4139, N2241);
nand NAND2 (N4142, N4104, N1218);
or OR2 (N4143, N4142, N1810);
buf BUF1 (N4144, N4105);
not NOT1 (N4145, N4140);
nor NOR3 (N4146, N4134, N2382, N38);
xor XOR2 (N4147, N4143, N3805);
and AND2 (N4148, N4132, N534);
not NOT1 (N4149, N4138);
nor NOR2 (N4150, N4111, N1615);
or OR3 (N4151, N4148, N2744, N3129);
nand NAND4 (N4152, N4130, N683, N2015, N3966);
and AND3 (N4153, N4147, N3882, N50);
buf BUF1 (N4154, N4152);
nand NAND2 (N4155, N4145, N3060);
nand NAND2 (N4156, N4151, N1494);
xor XOR2 (N4157, N4156, N1566);
or OR4 (N4158, N4144, N1910, N3181, N3626);
and AND3 (N4159, N4146, N2263, N1760);
buf BUF1 (N4160, N4159);
and AND2 (N4161, N4155, N3940);
nor NOR4 (N4162, N4153, N1188, N3297, N3526);
xor XOR2 (N4163, N4158, N3087);
buf BUF1 (N4164, N4149);
not NOT1 (N4165, N4161);
buf BUF1 (N4166, N4141);
nand NAND3 (N4167, N4164, N1498, N3007);
or OR3 (N4168, N4162, N604, N1879);
buf BUF1 (N4169, N4131);
and AND4 (N4170, N4163, N2332, N3174, N1645);
nand NAND2 (N4171, N4165, N3783);
xor XOR2 (N4172, N4168, N4015);
not NOT1 (N4173, N4169);
nor NOR2 (N4174, N4170, N3262);
not NOT1 (N4175, N4171);
nand NAND3 (N4176, N4157, N2197, N1508);
not NOT1 (N4177, N4176);
xor XOR2 (N4178, N4174, N2895);
buf BUF1 (N4179, N4167);
or OR2 (N4180, N4160, N1671);
nor NOR2 (N4181, N4154, N4015);
buf BUF1 (N4182, N4172);
not NOT1 (N4183, N4182);
nand NAND2 (N4184, N4166, N2505);
not NOT1 (N4185, N4150);
or OR2 (N4186, N4181, N2979);
nand NAND4 (N4187, N4186, N935, N2740, N2526);
nand NAND4 (N4188, N4183, N3732, N352, N2771);
buf BUF1 (N4189, N4180);
and AND4 (N4190, N4177, N830, N2751, N2612);
nand NAND2 (N4191, N4173, N3645);
buf BUF1 (N4192, N4184);
buf BUF1 (N4193, N4190);
nor NOR2 (N4194, N4189, N2461);
buf BUF1 (N4195, N4178);
nand NAND3 (N4196, N4193, N2492, N1027);
buf BUF1 (N4197, N4192);
not NOT1 (N4198, N4197);
or OR2 (N4199, N4191, N1690);
nor NOR3 (N4200, N4196, N3207, N687);
nand NAND3 (N4201, N4199, N2384, N1346);
and AND4 (N4202, N4201, N1984, N197, N2063);
buf BUF1 (N4203, N4194);
or OR2 (N4204, N4195, N2682);
not NOT1 (N4205, N4185);
nand NAND4 (N4206, N4198, N2301, N513, N706);
nor NOR2 (N4207, N4202, N425);
buf BUF1 (N4208, N4187);
and AND4 (N4209, N4175, N856, N829, N2901);
xor XOR2 (N4210, N4206, N3254);
xor XOR2 (N4211, N4204, N474);
or OR2 (N4212, N4200, N2743);
buf BUF1 (N4213, N4211);
nor NOR2 (N4214, N4203, N3064);
and AND2 (N4215, N4214, N2223);
xor XOR2 (N4216, N4215, N1237);
xor XOR2 (N4217, N4179, N2585);
nand NAND3 (N4218, N4216, N2061, N2098);
buf BUF1 (N4219, N4217);
and AND3 (N4220, N4188, N1827, N19);
or OR3 (N4221, N4207, N341, N1222);
not NOT1 (N4222, N4209);
nor NOR2 (N4223, N4210, N2830);
and AND4 (N4224, N4205, N3886, N3131, N3715);
xor XOR2 (N4225, N4221, N289);
nor NOR3 (N4226, N4222, N487, N3044);
and AND2 (N4227, N4223, N1875);
or OR4 (N4228, N4227, N900, N2333, N296);
buf BUF1 (N4229, N4213);
and AND2 (N4230, N4228, N3861);
buf BUF1 (N4231, N4208);
buf BUF1 (N4232, N4224);
buf BUF1 (N4233, N4231);
xor XOR2 (N4234, N4218, N1714);
xor XOR2 (N4235, N4219, N2250);
buf BUF1 (N4236, N4230);
nand NAND4 (N4237, N4220, N753, N1441, N574);
and AND4 (N4238, N4212, N1436, N2323, N1362);
not NOT1 (N4239, N4234);
nand NAND4 (N4240, N4233, N1634, N1582, N3901);
nor NOR3 (N4241, N4226, N3413, N1674);
xor XOR2 (N4242, N4240, N2961);
xor XOR2 (N4243, N4242, N3410);
nor NOR2 (N4244, N4238, N1530);
and AND3 (N4245, N4225, N3216, N2270);
xor XOR2 (N4246, N4236, N3317);
xor XOR2 (N4247, N4241, N2256);
or OR4 (N4248, N4246, N1380, N1860, N3567);
or OR4 (N4249, N4237, N3495, N3924, N1892);
nor NOR2 (N4250, N4248, N3951);
or OR2 (N4251, N4245, N983);
xor XOR2 (N4252, N4244, N3875);
nand NAND4 (N4253, N4232, N2737, N961, N1935);
and AND4 (N4254, N4250, N2105, N2863, N3853);
buf BUF1 (N4255, N4239);
nor NOR4 (N4256, N4247, N2333, N713, N4209);
or OR2 (N4257, N4249, N2042);
nor NOR3 (N4258, N4235, N1429, N1086);
xor XOR2 (N4259, N4251, N3140);
not NOT1 (N4260, N4257);
nand NAND4 (N4261, N4229, N2243, N1802, N4073);
not NOT1 (N4262, N4255);
not NOT1 (N4263, N4253);
nand NAND2 (N4264, N4254, N4177);
not NOT1 (N4265, N4258);
not NOT1 (N4266, N4263);
xor XOR2 (N4267, N4260, N1246);
buf BUF1 (N4268, N4259);
not NOT1 (N4269, N4265);
nand NAND3 (N4270, N4256, N1327, N4190);
or OR4 (N4271, N4266, N2821, N2708, N99);
xor XOR2 (N4272, N4267, N1231);
nor NOR3 (N4273, N4271, N1721, N1781);
and AND2 (N4274, N4252, N964);
and AND3 (N4275, N4274, N2801, N3086);
nor NOR2 (N4276, N4261, N4146);
xor XOR2 (N4277, N4268, N2987);
and AND3 (N4278, N4269, N4185, N2209);
and AND4 (N4279, N4270, N3223, N1145, N424);
nor NOR4 (N4280, N4243, N2771, N278, N1994);
buf BUF1 (N4281, N4262);
nor NOR2 (N4282, N4277, N3266);
not NOT1 (N4283, N4276);
not NOT1 (N4284, N4273);
or OR3 (N4285, N4279, N1636, N451);
or OR3 (N4286, N4282, N2770, N1651);
buf BUF1 (N4287, N4281);
and AND4 (N4288, N4280, N3187, N975, N3390);
not NOT1 (N4289, N4275);
or OR3 (N4290, N4278, N578, N2049);
not NOT1 (N4291, N4290);
buf BUF1 (N4292, N4289);
and AND4 (N4293, N4292, N2608, N1702, N3562);
and AND4 (N4294, N4283, N3574, N2667, N1210);
nand NAND3 (N4295, N4287, N1976, N1671);
not NOT1 (N4296, N4286);
nor NOR2 (N4297, N4296, N3963);
nand NAND4 (N4298, N4297, N2172, N824, N468);
nor NOR3 (N4299, N4288, N1191, N3129);
buf BUF1 (N4300, N4295);
not NOT1 (N4301, N4285);
not NOT1 (N4302, N4272);
nor NOR3 (N4303, N4293, N2953, N3106);
buf BUF1 (N4304, N4264);
or OR3 (N4305, N4298, N1390, N1652);
buf BUF1 (N4306, N4302);
nand NAND3 (N4307, N4306, N4069, N2988);
not NOT1 (N4308, N4300);
nor NOR2 (N4309, N4294, N319);
not NOT1 (N4310, N4303);
buf BUF1 (N4311, N4301);
xor XOR2 (N4312, N4311, N3283);
or OR4 (N4313, N4310, N3412, N2754, N1999);
not NOT1 (N4314, N4309);
nand NAND3 (N4315, N4314, N443, N2604);
and AND4 (N4316, N4304, N1407, N100, N2098);
and AND3 (N4317, N4315, N844, N531);
buf BUF1 (N4318, N4305);
buf BUF1 (N4319, N4317);
not NOT1 (N4320, N4307);
and AND3 (N4321, N4316, N3239, N37);
not NOT1 (N4322, N4308);
xor XOR2 (N4323, N4322, N3437);
nor NOR3 (N4324, N4284, N2842, N1863);
nor NOR2 (N4325, N4319, N862);
xor XOR2 (N4326, N4320, N3805);
and AND3 (N4327, N4325, N4248, N3270);
or OR2 (N4328, N4299, N1273);
not NOT1 (N4329, N4326);
buf BUF1 (N4330, N4312);
not NOT1 (N4331, N4323);
nand NAND3 (N4332, N4331, N3089, N1169);
xor XOR2 (N4333, N4324, N2202);
xor XOR2 (N4334, N4313, N2554);
nand NAND3 (N4335, N4328, N765, N3331);
and AND4 (N4336, N4318, N1969, N192, N224);
xor XOR2 (N4337, N4334, N434);
buf BUF1 (N4338, N4336);
and AND4 (N4339, N4338, N2233, N4168, N3623);
xor XOR2 (N4340, N4327, N232);
or OR4 (N4341, N4321, N1392, N2202, N1915);
and AND3 (N4342, N4335, N44, N1126);
nand NAND2 (N4343, N4332, N1855);
and AND4 (N4344, N4339, N1633, N3537, N1056);
or OR2 (N4345, N4342, N219);
nor NOR3 (N4346, N4345, N2368, N3545);
nor NOR4 (N4347, N4333, N3844, N1104, N605);
buf BUF1 (N4348, N4341);
nand NAND2 (N4349, N4340, N3285);
buf BUF1 (N4350, N4291);
nor NOR3 (N4351, N4349, N2387, N1648);
nor NOR3 (N4352, N4348, N2980, N3104);
nand NAND3 (N4353, N4329, N3208, N2556);
not NOT1 (N4354, N4351);
nand NAND4 (N4355, N4343, N2844, N2877, N1455);
not NOT1 (N4356, N4344);
not NOT1 (N4357, N4355);
nor NOR2 (N4358, N4347, N2336);
or OR3 (N4359, N4354, N4290, N3327);
nand NAND3 (N4360, N4346, N910, N2325);
xor XOR2 (N4361, N4350, N41);
and AND3 (N4362, N4360, N2380, N1438);
not NOT1 (N4363, N4352);
buf BUF1 (N4364, N4363);
xor XOR2 (N4365, N4361, N707);
nor NOR3 (N4366, N4330, N1403, N1260);
nor NOR2 (N4367, N4337, N2294);
and AND3 (N4368, N4364, N57, N37);
buf BUF1 (N4369, N4359);
or OR2 (N4370, N4362, N1954);
not NOT1 (N4371, N4356);
buf BUF1 (N4372, N4366);
not NOT1 (N4373, N4370);
or OR4 (N4374, N4367, N3098, N3362, N1773);
buf BUF1 (N4375, N4365);
nand NAND3 (N4376, N4369, N1790, N1188);
buf BUF1 (N4377, N4372);
not NOT1 (N4378, N4357);
nor NOR3 (N4379, N4353, N3925, N3803);
buf BUF1 (N4380, N4377);
buf BUF1 (N4381, N4368);
and AND4 (N4382, N4380, N1527, N1100, N3385);
and AND3 (N4383, N4378, N1093, N2181);
nand NAND4 (N4384, N4381, N3581, N392, N1457);
nor NOR2 (N4385, N4358, N4358);
and AND2 (N4386, N4385, N62);
not NOT1 (N4387, N4379);
buf BUF1 (N4388, N4387);
nand NAND3 (N4389, N4383, N131, N2813);
or OR2 (N4390, N4375, N4195);
or OR2 (N4391, N4388, N3829);
not NOT1 (N4392, N4384);
xor XOR2 (N4393, N4391, N1123);
nor NOR2 (N4394, N4376, N3601);
or OR2 (N4395, N4382, N2679);
xor XOR2 (N4396, N4386, N3407);
or OR2 (N4397, N4394, N2993);
xor XOR2 (N4398, N4390, N2341);
buf BUF1 (N4399, N4397);
or OR3 (N4400, N4399, N1123, N2489);
nor NOR2 (N4401, N4396, N3155);
or OR2 (N4402, N4373, N3908);
buf BUF1 (N4403, N4374);
buf BUF1 (N4404, N4393);
or OR4 (N4405, N4392, N4149, N3251, N2081);
buf BUF1 (N4406, N4400);
nand NAND4 (N4407, N4389, N1142, N3380, N3354);
xor XOR2 (N4408, N4395, N529);
and AND2 (N4409, N4402, N3983);
nor NOR3 (N4410, N4405, N3688, N1160);
xor XOR2 (N4411, N4401, N2096);
not NOT1 (N4412, N4403);
not NOT1 (N4413, N4407);
or OR3 (N4414, N4408, N3725, N992);
nor NOR4 (N4415, N4406, N1918, N2356, N4220);
xor XOR2 (N4416, N4413, N792);
nand NAND3 (N4417, N4404, N1630, N4023);
not NOT1 (N4418, N4412);
nor NOR3 (N4419, N4409, N2294, N3284);
or OR3 (N4420, N4419, N2374, N418);
nor NOR4 (N4421, N4420, N3958, N4222, N3241);
nand NAND3 (N4422, N4410, N1329, N595);
not NOT1 (N4423, N4415);
not NOT1 (N4424, N4414);
xor XOR2 (N4425, N4421, N2628);
or OR2 (N4426, N4411, N3817);
not NOT1 (N4427, N4424);
nor NOR2 (N4428, N4418, N1518);
and AND4 (N4429, N4426, N3029, N4272, N1866);
and AND4 (N4430, N4417, N3972, N2742, N2874);
buf BUF1 (N4431, N4429);
xor XOR2 (N4432, N4428, N1858);
nand NAND2 (N4433, N4416, N3788);
or OR2 (N4434, N4432, N1460);
xor XOR2 (N4435, N4398, N1718);
nor NOR4 (N4436, N4371, N3229, N3110, N2353);
and AND3 (N4437, N4435, N3331, N1320);
buf BUF1 (N4438, N4437);
nor NOR2 (N4439, N4436, N1375);
nand NAND3 (N4440, N4425, N1371, N4276);
and AND4 (N4441, N4434, N4404, N1455, N2902);
and AND3 (N4442, N4422, N65, N983);
nand NAND4 (N4443, N4441, N3694, N2619, N1707);
or OR4 (N4444, N4438, N3093, N2661, N764);
xor XOR2 (N4445, N4423, N1401);
nor NOR4 (N4446, N4427, N1105, N307, N2598);
xor XOR2 (N4447, N4443, N1178);
or OR4 (N4448, N4442, N3898, N2776, N1050);
nor NOR4 (N4449, N4444, N1672, N421, N2018);
not NOT1 (N4450, N4430);
or OR4 (N4451, N4439, N2493, N2595, N1087);
xor XOR2 (N4452, N4445, N3492);
nand NAND4 (N4453, N4452, N964, N126, N834);
and AND4 (N4454, N4446, N3593, N1801, N2278);
xor XOR2 (N4455, N4448, N1876);
xor XOR2 (N4456, N4433, N134);
nor NOR3 (N4457, N4449, N2667, N1903);
and AND4 (N4458, N4451, N2684, N3175, N319);
buf BUF1 (N4459, N4450);
nand NAND2 (N4460, N4457, N3394);
xor XOR2 (N4461, N4454, N1462);
xor XOR2 (N4462, N4460, N3201);
xor XOR2 (N4463, N4456, N1283);
xor XOR2 (N4464, N4447, N2563);
xor XOR2 (N4465, N4458, N1237);
or OR3 (N4466, N4453, N2401, N11);
and AND2 (N4467, N4465, N2095);
buf BUF1 (N4468, N4455);
not NOT1 (N4469, N4467);
nor NOR4 (N4470, N4468, N192, N1956, N2529);
or OR2 (N4471, N4459, N4394);
or OR3 (N4472, N4440, N739, N3734);
and AND3 (N4473, N4463, N3076, N1841);
nor NOR2 (N4474, N4471, N891);
xor XOR2 (N4475, N4431, N3298);
or OR4 (N4476, N4475, N1884, N1718, N2528);
or OR3 (N4477, N4469, N2997, N75);
not NOT1 (N4478, N4464);
and AND3 (N4479, N4472, N1411, N484);
nand NAND2 (N4480, N4470, N2874);
and AND3 (N4481, N4466, N4070, N4009);
nor NOR2 (N4482, N4478, N4361);
nand NAND4 (N4483, N4461, N3013, N202, N3692);
not NOT1 (N4484, N4477);
or OR2 (N4485, N4481, N764);
and AND2 (N4486, N4476, N1175);
xor XOR2 (N4487, N4483, N2848);
not NOT1 (N4488, N4484);
nand NAND4 (N4489, N4479, N875, N4389, N3079);
not NOT1 (N4490, N4462);
nand NAND4 (N4491, N4487, N172, N4031, N1081);
buf BUF1 (N4492, N4488);
not NOT1 (N4493, N4489);
or OR3 (N4494, N4492, N3140, N4255);
nand NAND3 (N4495, N4474, N1329, N4346);
or OR3 (N4496, N4495, N4470, N2774);
xor XOR2 (N4497, N4496, N3528);
not NOT1 (N4498, N4485);
nand NAND3 (N4499, N4491, N1023, N4445);
and AND2 (N4500, N4480, N2707);
buf BUF1 (N4501, N4497);
or OR2 (N4502, N4473, N2203);
buf BUF1 (N4503, N4499);
or OR3 (N4504, N4498, N263, N3497);
xor XOR2 (N4505, N4482, N1890);
or OR4 (N4506, N4490, N1104, N1873, N3666);
nor NOR4 (N4507, N4493, N953, N3192, N1711);
buf BUF1 (N4508, N4505);
and AND4 (N4509, N4504, N3598, N2285, N528);
and AND2 (N4510, N4503, N2328);
nand NAND4 (N4511, N4506, N2069, N1340, N1887);
or OR3 (N4512, N4494, N1557, N3136);
or OR4 (N4513, N4509, N1965, N2687, N3891);
xor XOR2 (N4514, N4507, N4382);
buf BUF1 (N4515, N4511);
buf BUF1 (N4516, N4514);
xor XOR2 (N4517, N4516, N4363);
nand NAND4 (N4518, N4486, N6, N3728, N4076);
nor NOR3 (N4519, N4508, N1562, N4319);
nor NOR2 (N4520, N4519, N3032);
and AND4 (N4521, N4515, N1249, N3237, N1519);
buf BUF1 (N4522, N4512);
or OR2 (N4523, N4520, N857);
or OR4 (N4524, N4510, N3851, N123, N2337);
and AND2 (N4525, N4524, N686);
buf BUF1 (N4526, N4521);
or OR4 (N4527, N4517, N4374, N4339, N2360);
xor XOR2 (N4528, N4523, N1942);
nor NOR3 (N4529, N4500, N1941, N4118);
and AND2 (N4530, N4528, N611);
or OR3 (N4531, N4526, N3834, N871);
nor NOR4 (N4532, N4501, N3378, N1595, N3337);
or OR3 (N4533, N4518, N1475, N389);
and AND4 (N4534, N4532, N1741, N4198, N3582);
or OR3 (N4535, N4502, N406, N4382);
xor XOR2 (N4536, N4529, N3028);
and AND2 (N4537, N4531, N3241);
nand NAND2 (N4538, N4522, N4360);
xor XOR2 (N4539, N4533, N2399);
nand NAND2 (N4540, N4539, N1423);
and AND4 (N4541, N4525, N3659, N2059, N1525);
not NOT1 (N4542, N4527);
xor XOR2 (N4543, N4513, N2064);
nand NAND2 (N4544, N4540, N3663);
not NOT1 (N4545, N4537);
buf BUF1 (N4546, N4538);
and AND3 (N4547, N4542, N2781, N2690);
nand NAND4 (N4548, N4543, N1077, N668, N3320);
xor XOR2 (N4549, N4530, N2647);
not NOT1 (N4550, N4541);
nand NAND3 (N4551, N4546, N401, N696);
or OR2 (N4552, N4548, N1572);
buf BUF1 (N4553, N4551);
and AND2 (N4554, N4545, N2982);
not NOT1 (N4555, N4552);
xor XOR2 (N4556, N4549, N2927);
or OR2 (N4557, N4534, N2184);
xor XOR2 (N4558, N4553, N2956);
nor NOR4 (N4559, N4544, N2526, N569, N103);
not NOT1 (N4560, N4559);
nor NOR3 (N4561, N4550, N1528, N2334);
and AND4 (N4562, N4558, N3910, N1598, N179);
and AND3 (N4563, N4555, N3438, N1286);
buf BUF1 (N4564, N4554);
and AND3 (N4565, N4564, N1231, N258);
nor NOR4 (N4566, N4560, N21, N2124, N3642);
not NOT1 (N4567, N4561);
buf BUF1 (N4568, N4536);
and AND4 (N4569, N4557, N455, N1389, N815);
xor XOR2 (N4570, N4562, N1731);
or OR4 (N4571, N4565, N113, N4175, N14);
nor NOR2 (N4572, N4547, N4272);
buf BUF1 (N4573, N4572);
buf BUF1 (N4574, N4573);
xor XOR2 (N4575, N4569, N119);
nand NAND4 (N4576, N4556, N1096, N1342, N2053);
not NOT1 (N4577, N4576);
buf BUF1 (N4578, N4568);
buf BUF1 (N4579, N4567);
buf BUF1 (N4580, N4575);
nor NOR2 (N4581, N4570, N2037);
and AND4 (N4582, N4535, N2195, N3012, N34);
not NOT1 (N4583, N4566);
buf BUF1 (N4584, N4583);
xor XOR2 (N4585, N4581, N4182);
xor XOR2 (N4586, N4585, N1037);
and AND3 (N4587, N4578, N584, N4564);
not NOT1 (N4588, N4571);
xor XOR2 (N4589, N4563, N2258);
or OR4 (N4590, N4588, N839, N4583, N2994);
nor NOR4 (N4591, N4589, N522, N2570, N1148);
nand NAND2 (N4592, N4580, N2598);
or OR3 (N4593, N4587, N3316, N3533);
nand NAND3 (N4594, N4590, N3726, N4283);
nand NAND3 (N4595, N4574, N4306, N3726);
buf BUF1 (N4596, N4593);
xor XOR2 (N4597, N4586, N1419);
or OR4 (N4598, N4582, N4123, N4253, N11);
not NOT1 (N4599, N4579);
nor NOR3 (N4600, N4594, N3888, N4198);
buf BUF1 (N4601, N4597);
xor XOR2 (N4602, N4600, N1529);
or OR2 (N4603, N4601, N3333);
xor XOR2 (N4604, N4599, N4019);
buf BUF1 (N4605, N4604);
not NOT1 (N4606, N4592);
buf BUF1 (N4607, N4577);
buf BUF1 (N4608, N4584);
nand NAND2 (N4609, N4598, N1141);
nand NAND2 (N4610, N4608, N3113);
and AND4 (N4611, N4602, N1107, N1416, N4127);
buf BUF1 (N4612, N4611);
and AND4 (N4613, N4596, N1409, N1882, N604);
nand NAND2 (N4614, N4595, N1086);
not NOT1 (N4615, N4607);
and AND2 (N4616, N4613, N4266);
buf BUF1 (N4617, N4614);
nand NAND2 (N4618, N4605, N3813);
nand NAND4 (N4619, N4618, N3640, N2114, N168);
or OR3 (N4620, N4610, N1231, N820);
buf BUF1 (N4621, N4591);
not NOT1 (N4622, N4619);
nand NAND2 (N4623, N4612, N2765);
not NOT1 (N4624, N4615);
and AND2 (N4625, N4624, N1974);
xor XOR2 (N4626, N4609, N228);
nand NAND4 (N4627, N4606, N3092, N3704, N123);
or OR4 (N4628, N4617, N3042, N3243, N638);
and AND2 (N4629, N4603, N327);
and AND3 (N4630, N4625, N4273, N2956);
nor NOR3 (N4631, N4621, N660, N3450);
and AND4 (N4632, N4630, N3316, N1564, N1285);
buf BUF1 (N4633, N4631);
and AND4 (N4634, N4626, N1387, N774, N405);
nand NAND2 (N4635, N4632, N410);
xor XOR2 (N4636, N4633, N4559);
or OR2 (N4637, N4628, N1430);
buf BUF1 (N4638, N4634);
buf BUF1 (N4639, N4623);
nor NOR4 (N4640, N4638, N401, N4007, N2347);
and AND4 (N4641, N4627, N4087, N1362, N1335);
nor NOR4 (N4642, N4620, N2938, N578, N3866);
not NOT1 (N4643, N4641);
buf BUF1 (N4644, N4640);
not NOT1 (N4645, N4643);
not NOT1 (N4646, N4616);
and AND4 (N4647, N4637, N421, N1752, N446);
buf BUF1 (N4648, N4622);
and AND3 (N4649, N4644, N4643, N3112);
xor XOR2 (N4650, N4639, N1458);
or OR4 (N4651, N4629, N536, N234, N2584);
buf BUF1 (N4652, N4646);
and AND3 (N4653, N4642, N3586, N3252);
not NOT1 (N4654, N4653);
and AND2 (N4655, N4636, N863);
nand NAND3 (N4656, N4645, N3031, N1836);
and AND2 (N4657, N4656, N1193);
not NOT1 (N4658, N4652);
nand NAND4 (N4659, N4651, N4405, N1065, N294);
and AND4 (N4660, N4635, N2643, N3945, N333);
and AND2 (N4661, N4650, N4101);
and AND3 (N4662, N4659, N2353, N2360);
and AND4 (N4663, N4661, N1087, N3997, N4433);
xor XOR2 (N4664, N4657, N1309);
nand NAND2 (N4665, N4663, N3988);
and AND4 (N4666, N4664, N3994, N66, N860);
or OR2 (N4667, N4655, N3180);
and AND3 (N4668, N4658, N2413, N2413);
not NOT1 (N4669, N4666);
nand NAND2 (N4670, N4662, N3681);
or OR3 (N4671, N4665, N2840, N2990);
or OR4 (N4672, N4648, N512, N3567, N1994);
nor NOR2 (N4673, N4667, N3170);
nand NAND2 (N4674, N4671, N1770);
buf BUF1 (N4675, N4674);
buf BUF1 (N4676, N4654);
nand NAND3 (N4677, N4672, N672, N3691);
nand NAND4 (N4678, N4668, N805, N1934, N425);
buf BUF1 (N4679, N4670);
buf BUF1 (N4680, N4660);
buf BUF1 (N4681, N4678);
not NOT1 (N4682, N4647);
and AND3 (N4683, N4649, N669, N47);
nand NAND2 (N4684, N4682, N2871);
nor NOR2 (N4685, N4677, N669);
not NOT1 (N4686, N4679);
nand NAND4 (N4687, N4685, N893, N1671, N1830);
buf BUF1 (N4688, N4673);
buf BUF1 (N4689, N4684);
not NOT1 (N4690, N4687);
xor XOR2 (N4691, N4689, N1325);
not NOT1 (N4692, N4688);
and AND4 (N4693, N4690, N1616, N3350, N3555);
nor NOR2 (N4694, N4686, N4142);
not NOT1 (N4695, N4675);
nand NAND2 (N4696, N4691, N4417);
nand NAND3 (N4697, N4669, N4425, N150);
nand NAND2 (N4698, N4697, N1119);
or OR4 (N4699, N4696, N4607, N3981, N415);
and AND4 (N4700, N4680, N2539, N668, N4466);
not NOT1 (N4701, N4700);
buf BUF1 (N4702, N4701);
nor NOR2 (N4703, N4693, N3388);
buf BUF1 (N4704, N4703);
buf BUF1 (N4705, N4683);
xor XOR2 (N4706, N4698, N649);
buf BUF1 (N4707, N4681);
and AND2 (N4708, N4694, N4106);
nand NAND3 (N4709, N4699, N2580, N750);
not NOT1 (N4710, N4708);
xor XOR2 (N4711, N4709, N4634);
or OR4 (N4712, N4710, N2108, N3445, N2616);
nor NOR2 (N4713, N4706, N3160);
not NOT1 (N4714, N4702);
not NOT1 (N4715, N4713);
nor NOR3 (N4716, N4707, N647, N4553);
nand NAND3 (N4717, N4705, N4618, N4542);
not NOT1 (N4718, N4692);
nor NOR2 (N4719, N4715, N3201);
nand NAND2 (N4720, N4704, N1020);
and AND3 (N4721, N4720, N4090, N4507);
nand NAND4 (N4722, N4716, N2410, N726, N3365);
nand NAND3 (N4723, N4721, N1316, N703);
not NOT1 (N4724, N4712);
or OR3 (N4725, N4695, N765, N2786);
and AND3 (N4726, N4714, N4676, N3996);
buf BUF1 (N4727, N1613);
xor XOR2 (N4728, N4724, N1053);
and AND4 (N4729, N4723, N1681, N956, N1939);
xor XOR2 (N4730, N4718, N2143);
not NOT1 (N4731, N4717);
not NOT1 (N4732, N4726);
buf BUF1 (N4733, N4727);
nor NOR4 (N4734, N4731, N63, N2019, N3309);
buf BUF1 (N4735, N4722);
xor XOR2 (N4736, N4735, N4488);
or OR4 (N4737, N4733, N3273, N621, N4653);
xor XOR2 (N4738, N4711, N1940);
or OR3 (N4739, N4719, N2, N4312);
and AND2 (N4740, N4738, N2974);
nor NOR2 (N4741, N4732, N2166);
or OR3 (N4742, N4739, N2080, N3480);
or OR3 (N4743, N4729, N4201, N4630);
or OR3 (N4744, N4741, N4028, N566);
nor NOR2 (N4745, N4728, N2930);
xor XOR2 (N4746, N4725, N797);
not NOT1 (N4747, N4746);
not NOT1 (N4748, N4745);
nand NAND4 (N4749, N4736, N260, N907, N1325);
nand NAND3 (N4750, N4740, N4045, N737);
nor NOR4 (N4751, N4747, N9, N447, N1227);
or OR4 (N4752, N4744, N3232, N1939, N1159);
nand NAND3 (N4753, N4749, N3075, N2132);
nand NAND2 (N4754, N4753, N3530);
or OR3 (N4755, N4754, N419, N4292);
nand NAND2 (N4756, N4737, N2403);
xor XOR2 (N4757, N4751, N4491);
not NOT1 (N4758, N4755);
not NOT1 (N4759, N4752);
buf BUF1 (N4760, N4756);
or OR4 (N4761, N4734, N604, N2557, N1644);
xor XOR2 (N4762, N4759, N794);
nor NOR2 (N4763, N4762, N1306);
buf BUF1 (N4764, N4742);
and AND2 (N4765, N4757, N1734);
not NOT1 (N4766, N4758);
not NOT1 (N4767, N4730);
and AND2 (N4768, N4767, N4450);
xor XOR2 (N4769, N4768, N2990);
and AND3 (N4770, N4760, N210, N1001);
or OR2 (N4771, N4764, N1828);
xor XOR2 (N4772, N4765, N4050);
buf BUF1 (N4773, N4771);
nand NAND3 (N4774, N4770, N3213, N25);
buf BUF1 (N4775, N4761);
xor XOR2 (N4776, N4743, N119);
xor XOR2 (N4777, N4775, N544);
xor XOR2 (N4778, N4750, N1732);
nor NOR2 (N4779, N4777, N4170);
and AND2 (N4780, N4763, N600);
xor XOR2 (N4781, N4766, N4045);
nand NAND4 (N4782, N4772, N2335, N2000, N2269);
nand NAND2 (N4783, N4769, N4588);
and AND3 (N4784, N4748, N3879, N315);
nand NAND2 (N4785, N4778, N3941);
and AND3 (N4786, N4782, N4299, N907);
or OR4 (N4787, N4774, N4220, N764, N1297);
nor NOR2 (N4788, N4783, N2763);
nand NAND3 (N4789, N4780, N3798, N2402);
nand NAND2 (N4790, N4784, N4738);
xor XOR2 (N4791, N4773, N3132);
nor NOR2 (N4792, N4790, N367);
not NOT1 (N4793, N4781);
buf BUF1 (N4794, N4776);
not NOT1 (N4795, N4789);
buf BUF1 (N4796, N4787);
nor NOR2 (N4797, N4793, N2296);
nor NOR2 (N4798, N4791, N4668);
or OR2 (N4799, N4794, N1543);
or OR3 (N4800, N4786, N3923, N1099);
buf BUF1 (N4801, N4792);
nor NOR2 (N4802, N4788, N3069);
and AND3 (N4803, N4797, N970, N2357);
nor NOR4 (N4804, N4796, N2750, N2930, N3738);
and AND4 (N4805, N4779, N3064, N1690, N4105);
xor XOR2 (N4806, N4801, N3651);
buf BUF1 (N4807, N4798);
nor NOR2 (N4808, N4802, N3243);
or OR4 (N4809, N4785, N1891, N1189, N424);
buf BUF1 (N4810, N4803);
nand NAND4 (N4811, N4800, N3998, N182, N3484);
buf BUF1 (N4812, N4808);
buf BUF1 (N4813, N4804);
nor NOR4 (N4814, N4806, N1952, N960, N4477);
not NOT1 (N4815, N4805);
or OR3 (N4816, N4812, N3674, N1280);
and AND4 (N4817, N4795, N3002, N206, N2232);
and AND3 (N4818, N4815, N2827, N3238);
and AND4 (N4819, N4809, N3384, N2239, N4015);
xor XOR2 (N4820, N4811, N4436);
nand NAND2 (N4821, N4807, N140);
not NOT1 (N4822, N4821);
xor XOR2 (N4823, N4816, N271);
buf BUF1 (N4824, N4810);
nor NOR3 (N4825, N4824, N4250, N3238);
buf BUF1 (N4826, N4818);
or OR2 (N4827, N4822, N2181);
nor NOR4 (N4828, N4814, N4545, N3480, N1868);
xor XOR2 (N4829, N4827, N4665);
xor XOR2 (N4830, N4826, N1818);
xor XOR2 (N4831, N4820, N4504);
xor XOR2 (N4832, N4817, N1060);
and AND3 (N4833, N4828, N298, N1604);
xor XOR2 (N4834, N4823, N4797);
nand NAND4 (N4835, N4799, N3252, N3008, N2812);
nor NOR4 (N4836, N4831, N1814, N2663, N2648);
not NOT1 (N4837, N4829);
and AND2 (N4838, N4837, N1704);
and AND4 (N4839, N4813, N4577, N676, N4572);
nor NOR2 (N4840, N4819, N2687);
xor XOR2 (N4841, N4833, N4094);
and AND2 (N4842, N4836, N3795);
or OR2 (N4843, N4842, N3563);
buf BUF1 (N4844, N4843);
and AND3 (N4845, N4839, N4408, N4063);
nor NOR2 (N4846, N4838, N4367);
buf BUF1 (N4847, N4844);
or OR2 (N4848, N4830, N4439);
nor NOR2 (N4849, N4847, N2558);
nand NAND3 (N4850, N4832, N1829, N2493);
nand NAND2 (N4851, N4849, N65);
nor NOR3 (N4852, N4840, N1681, N2666);
not NOT1 (N4853, N4834);
xor XOR2 (N4854, N4845, N2133);
or OR4 (N4855, N4825, N2342, N3618, N3103);
buf BUF1 (N4856, N4841);
buf BUF1 (N4857, N4855);
buf BUF1 (N4858, N4851);
not NOT1 (N4859, N4854);
not NOT1 (N4860, N4846);
xor XOR2 (N4861, N4859, N1621);
nor NOR2 (N4862, N4857, N1956);
nor NOR3 (N4863, N4835, N4119, N2624);
not NOT1 (N4864, N4853);
nand NAND2 (N4865, N4864, N209);
nor NOR4 (N4866, N4848, N2460, N2229, N3941);
not NOT1 (N4867, N4863);
nand NAND4 (N4868, N4860, N4007, N2128, N4653);
buf BUF1 (N4869, N4867);
and AND2 (N4870, N4850, N1313);
nor NOR3 (N4871, N4856, N1300, N1872);
not NOT1 (N4872, N4866);
and AND2 (N4873, N4872, N3448);
buf BUF1 (N4874, N4862);
or OR3 (N4875, N4870, N3422, N928);
or OR2 (N4876, N4852, N391);
or OR3 (N4877, N4874, N821, N1681);
or OR4 (N4878, N4871, N4142, N3310, N2805);
nand NAND4 (N4879, N4858, N1277, N759, N4324);
not NOT1 (N4880, N4869);
xor XOR2 (N4881, N4879, N1247);
xor XOR2 (N4882, N4875, N2034);
nand NAND3 (N4883, N4861, N1287, N2477);
nor NOR2 (N4884, N4868, N3247);
or OR2 (N4885, N4877, N2012);
nor NOR4 (N4886, N4882, N3619, N1631, N832);
nor NOR4 (N4887, N4878, N2526, N464, N4878);
xor XOR2 (N4888, N4885, N4005);
buf BUF1 (N4889, N4883);
xor XOR2 (N4890, N4886, N3385);
or OR4 (N4891, N4865, N890, N376, N2536);
nand NAND3 (N4892, N4873, N61, N2743);
xor XOR2 (N4893, N4892, N3329);
buf BUF1 (N4894, N4888);
or OR4 (N4895, N4889, N3968, N3699, N2208);
nand NAND3 (N4896, N4894, N654, N256);
not NOT1 (N4897, N4890);
nor NOR2 (N4898, N4881, N961);
buf BUF1 (N4899, N4880);
or OR2 (N4900, N4896, N4032);
and AND3 (N4901, N4900, N1283, N1926);
nor NOR3 (N4902, N4899, N3170, N2568);
or OR4 (N4903, N4897, N1568, N374, N2041);
buf BUF1 (N4904, N4891);
or OR3 (N4905, N4884, N3320, N2535);
or OR2 (N4906, N4901, N302);
or OR3 (N4907, N4893, N1567, N1382);
nor NOR3 (N4908, N4898, N3478, N1104);
and AND4 (N4909, N4905, N2554, N2295, N2464);
not NOT1 (N4910, N4895);
buf BUF1 (N4911, N4906);
and AND3 (N4912, N4904, N3431, N3165);
nand NAND3 (N4913, N4902, N1404, N2704);
or OR4 (N4914, N4909, N4239, N1900, N1785);
and AND2 (N4915, N4910, N4706);
buf BUF1 (N4916, N4903);
and AND3 (N4917, N4911, N3605, N1181);
nor NOR2 (N4918, N4915, N710);
not NOT1 (N4919, N4916);
nand NAND3 (N4920, N4876, N3038, N2819);
nand NAND2 (N4921, N4913, N2128);
nor NOR3 (N4922, N4918, N2378, N4366);
or OR4 (N4923, N4914, N3275, N2392, N2005);
not NOT1 (N4924, N4908);
and AND2 (N4925, N4907, N4635);
nand NAND4 (N4926, N4921, N2424, N2497, N2549);
buf BUF1 (N4927, N4924);
nor NOR4 (N4928, N4920, N412, N3352, N905);
xor XOR2 (N4929, N4912, N4544);
nand NAND4 (N4930, N4917, N756, N1927, N1058);
or OR2 (N4931, N4925, N1152);
nand NAND4 (N4932, N4927, N1228, N4461, N1378);
and AND2 (N4933, N4930, N2719);
buf BUF1 (N4934, N4919);
not NOT1 (N4935, N4887);
or OR2 (N4936, N4934, N1866);
xor XOR2 (N4937, N4932, N645);
xor XOR2 (N4938, N4935, N2718);
or OR3 (N4939, N4928, N3357, N3597);
xor XOR2 (N4940, N4929, N1627);
buf BUF1 (N4941, N4940);
or OR2 (N4942, N4936, N1110);
not NOT1 (N4943, N4939);
or OR3 (N4944, N4931, N3231, N4798);
and AND4 (N4945, N4933, N3390, N462, N1855);
nor NOR2 (N4946, N4926, N3596);
nor NOR4 (N4947, N4944, N756, N3183, N3572);
buf BUF1 (N4948, N4922);
nor NOR4 (N4949, N4946, N2351, N564, N2764);
buf BUF1 (N4950, N4942);
buf BUF1 (N4951, N4945);
not NOT1 (N4952, N4943);
nor NOR3 (N4953, N4947, N832, N17);
and AND3 (N4954, N4952, N4366, N1455);
and AND3 (N4955, N4941, N187, N1142);
xor XOR2 (N4956, N4948, N4277);
or OR2 (N4957, N4951, N1518);
nand NAND4 (N4958, N4937, N751, N2162, N1766);
nor NOR2 (N4959, N4957, N598);
and AND3 (N4960, N4954, N4660, N1842);
nor NOR4 (N4961, N4950, N2154, N3511, N3595);
and AND4 (N4962, N4956, N3529, N4604, N3113);
xor XOR2 (N4963, N4938, N1555);
not NOT1 (N4964, N4960);
nand NAND3 (N4965, N4949, N3093, N4595);
and AND4 (N4966, N4964, N2680, N3565, N1110);
buf BUF1 (N4967, N4959);
nor NOR2 (N4968, N4958, N1085);
buf BUF1 (N4969, N4966);
xor XOR2 (N4970, N4962, N4004);
xor XOR2 (N4971, N4963, N2201);
not NOT1 (N4972, N4961);
nand NAND3 (N4973, N4965, N219, N3984);
not NOT1 (N4974, N4953);
nand NAND4 (N4975, N4971, N55, N50, N1204);
not NOT1 (N4976, N4969);
nor NOR3 (N4977, N4967, N955, N3032);
not NOT1 (N4978, N4975);
buf BUF1 (N4979, N4978);
and AND4 (N4980, N4923, N4006, N713, N560);
and AND3 (N4981, N4974, N3160, N4229);
nor NOR4 (N4982, N4980, N1220, N1549, N3393);
nor NOR2 (N4983, N4981, N1777);
and AND3 (N4984, N4970, N1637, N2750);
and AND3 (N4985, N4976, N4649, N3120);
xor XOR2 (N4986, N4984, N3251);
nor NOR4 (N4987, N4986, N4324, N4743, N4337);
xor XOR2 (N4988, N4955, N4286);
nor NOR4 (N4989, N4979, N2317, N3162, N2338);
nand NAND2 (N4990, N4977, N2412);
not NOT1 (N4991, N4972);
xor XOR2 (N4992, N4985, N393);
nor NOR3 (N4993, N4988, N1920, N1921);
or OR2 (N4994, N4973, N1477);
buf BUF1 (N4995, N4991);
nor NOR2 (N4996, N4990, N2521);
or OR3 (N4997, N4982, N2566, N3620);
buf BUF1 (N4998, N4983);
not NOT1 (N4999, N4992);
or OR3 (N5000, N4968, N3706, N1868);
not NOT1 (N5001, N4994);
and AND4 (N5002, N4995, N720, N3615, N2991);
xor XOR2 (N5003, N4997, N4844);
nor NOR4 (N5004, N5002, N3728, N4623, N1327);
nor NOR4 (N5005, N4996, N4999, N3304, N571);
nand NAND3 (N5006, N3280, N4160, N4273);
nand NAND2 (N5007, N5005, N1659);
or OR2 (N5008, N5004, N3339);
not NOT1 (N5009, N4989);
or OR2 (N5010, N5006, N399);
buf BUF1 (N5011, N4993);
xor XOR2 (N5012, N5001, N2377);
buf BUF1 (N5013, N4987);
nor NOR4 (N5014, N5007, N3847, N1241, N4295);
buf BUF1 (N5015, N5000);
or OR2 (N5016, N5015, N4150);
xor XOR2 (N5017, N5012, N4553);
xor XOR2 (N5018, N5014, N1716);
nand NAND2 (N5019, N5003, N3718);
not NOT1 (N5020, N5017);
buf BUF1 (N5021, N5020);
buf BUF1 (N5022, N4998);
and AND3 (N5023, N5016, N197, N2751);
nand NAND4 (N5024, N5009, N1879, N484, N1532);
nor NOR4 (N5025, N5023, N270, N764, N979);
and AND2 (N5026, N5025, N734);
xor XOR2 (N5027, N5013, N2035);
or OR2 (N5028, N5024, N4714);
or OR4 (N5029, N5022, N4973, N4713, N4127);
and AND2 (N5030, N5026, N3593);
nand NAND4 (N5031, N5010, N943, N2749, N3063);
or OR4 (N5032, N5011, N1534, N3138, N1);
and AND2 (N5033, N5031, N63);
or OR4 (N5034, N5028, N252, N4884, N1676);
nand NAND2 (N5035, N5021, N2311);
nand NAND3 (N5036, N5032, N2810, N2024);
nor NOR2 (N5037, N5033, N2886);
nor NOR2 (N5038, N5018, N3720);
and AND3 (N5039, N5034, N3213, N2939);
nand NAND3 (N5040, N5036, N1731, N3807);
not NOT1 (N5041, N5029);
not NOT1 (N5042, N5041);
nor NOR3 (N5043, N5040, N2655, N4480);
nand NAND2 (N5044, N5030, N4810);
nor NOR4 (N5045, N5042, N4181, N2848, N3757);
or OR2 (N5046, N5043, N385);
xor XOR2 (N5047, N5038, N2503);
xor XOR2 (N5048, N5019, N76);
xor XOR2 (N5049, N5046, N199);
not NOT1 (N5050, N5008);
buf BUF1 (N5051, N5035);
not NOT1 (N5052, N5048);
and AND3 (N5053, N5037, N76, N401);
buf BUF1 (N5054, N5047);
or OR4 (N5055, N5054, N1646, N1985, N1429);
buf BUF1 (N5056, N5049);
not NOT1 (N5057, N5055);
not NOT1 (N5058, N5044);
not NOT1 (N5059, N5053);
not NOT1 (N5060, N5058);
buf BUF1 (N5061, N5056);
or OR3 (N5062, N5057, N17, N3585);
nand NAND2 (N5063, N5052, N495);
and AND2 (N5064, N5050, N2505);
xor XOR2 (N5065, N5063, N3284);
xor XOR2 (N5066, N5065, N4078);
not NOT1 (N5067, N5064);
buf BUF1 (N5068, N5060);
or OR3 (N5069, N5027, N4417, N4929);
nand NAND2 (N5070, N5069, N2501);
and AND2 (N5071, N5061, N5034);
buf BUF1 (N5072, N5068);
buf BUF1 (N5073, N5045);
or OR2 (N5074, N5062, N942);
nor NOR3 (N5075, N5051, N452, N1489);
or OR2 (N5076, N5070, N3757);
buf BUF1 (N5077, N5072);
buf BUF1 (N5078, N5076);
or OR4 (N5079, N5078, N1680, N1543, N4691);
nor NOR2 (N5080, N5074, N1885);
or OR2 (N5081, N5059, N1759);
and AND3 (N5082, N5039, N1561, N947);
and AND4 (N5083, N5082, N3973, N1979, N1146);
nand NAND3 (N5084, N5081, N934, N1430);
buf BUF1 (N5085, N5067);
and AND4 (N5086, N5080, N4996, N2441, N4027);
not NOT1 (N5087, N5077);
nor NOR4 (N5088, N5086, N1902, N4253, N702);
nor NOR2 (N5089, N5073, N127);
or OR3 (N5090, N5085, N129, N1757);
xor XOR2 (N5091, N5071, N2877);
or OR4 (N5092, N5089, N2397, N574, N306);
xor XOR2 (N5093, N5079, N1644);
and AND2 (N5094, N5066, N563);
buf BUF1 (N5095, N5093);
or OR2 (N5096, N5075, N2126);
not NOT1 (N5097, N5094);
xor XOR2 (N5098, N5090, N4872);
and AND4 (N5099, N5091, N4094, N4907, N1482);
or OR2 (N5100, N5087, N4436);
nand NAND2 (N5101, N5095, N1570);
xor XOR2 (N5102, N5097, N3821);
xor XOR2 (N5103, N5100, N4832);
xor XOR2 (N5104, N5103, N822);
nor NOR2 (N5105, N5083, N2237);
and AND4 (N5106, N5105, N5012, N3225, N1297);
not NOT1 (N5107, N5098);
nand NAND3 (N5108, N5096, N3148, N4117);
xor XOR2 (N5109, N5099, N821);
nor NOR4 (N5110, N5088, N3837, N3665, N1359);
or OR4 (N5111, N5108, N4312, N3557, N3930);
xor XOR2 (N5112, N5084, N4281);
buf BUF1 (N5113, N5104);
and AND2 (N5114, N5113, N123);
buf BUF1 (N5115, N5101);
xor XOR2 (N5116, N5115, N821);
nand NAND2 (N5117, N5109, N2591);
nand NAND2 (N5118, N5106, N3321);
buf BUF1 (N5119, N5102);
xor XOR2 (N5120, N5092, N1148);
nand NAND2 (N5121, N5112, N4537);
xor XOR2 (N5122, N5116, N3693);
buf BUF1 (N5123, N5111);
nand NAND3 (N5124, N5119, N743, N582);
not NOT1 (N5125, N5117);
or OR3 (N5126, N5123, N2932, N918);
or OR4 (N5127, N5114, N4280, N3650, N3179);
nor NOR4 (N5128, N5118, N2072, N127, N734);
or OR4 (N5129, N5107, N1039, N3310, N1601);
xor XOR2 (N5130, N5129, N2459);
not NOT1 (N5131, N5124);
nand NAND2 (N5132, N5110, N4142);
nand NAND4 (N5133, N5128, N970, N2296, N4983);
nor NOR2 (N5134, N5126, N2230);
nor NOR3 (N5135, N5122, N703, N3163);
nand NAND2 (N5136, N5134, N4414);
not NOT1 (N5137, N5131);
buf BUF1 (N5138, N5133);
xor XOR2 (N5139, N5125, N4696);
buf BUF1 (N5140, N5121);
buf BUF1 (N5141, N5139);
not NOT1 (N5142, N5140);
and AND4 (N5143, N5142, N1011, N3869, N461);
xor XOR2 (N5144, N5137, N3093);
nand NAND2 (N5145, N5135, N1672);
not NOT1 (N5146, N5138);
buf BUF1 (N5147, N5146);
xor XOR2 (N5148, N5136, N2878);
xor XOR2 (N5149, N5148, N2448);
and AND2 (N5150, N5130, N3616);
or OR2 (N5151, N5144, N4591);
and AND4 (N5152, N5120, N1565, N4939, N1730);
and AND2 (N5153, N5127, N2707);
not NOT1 (N5154, N5151);
and AND2 (N5155, N5152, N1435);
and AND3 (N5156, N5155, N1887, N4626);
buf BUF1 (N5157, N5147);
xor XOR2 (N5158, N5141, N265);
not NOT1 (N5159, N5153);
nand NAND2 (N5160, N5149, N3486);
and AND2 (N5161, N5157, N612);
and AND3 (N5162, N5156, N1837, N229);
or OR2 (N5163, N5160, N4818);
and AND4 (N5164, N5159, N593, N3671, N4153);
or OR4 (N5165, N5132, N1997, N3431, N3681);
nand NAND2 (N5166, N5161, N4805);
nor NOR3 (N5167, N5158, N3498, N2518);
or OR4 (N5168, N5162, N4075, N174, N101);
and AND4 (N5169, N5167, N3371, N274, N4379);
not NOT1 (N5170, N5169);
not NOT1 (N5171, N5168);
xor XOR2 (N5172, N5164, N2289);
nand NAND2 (N5173, N5166, N1219);
and AND2 (N5174, N5173, N1227);
nor NOR3 (N5175, N5171, N5039, N4003);
or OR3 (N5176, N5175, N1361, N3003);
nand NAND3 (N5177, N5143, N2757, N3338);
not NOT1 (N5178, N5145);
not NOT1 (N5179, N5176);
and AND4 (N5180, N5154, N3291, N5124, N2940);
nor NOR4 (N5181, N5165, N5142, N1756, N1252);
nand NAND3 (N5182, N5150, N4604, N4940);
nand NAND3 (N5183, N5177, N1806, N2667);
buf BUF1 (N5184, N5174);
nand NAND4 (N5185, N5172, N2707, N3683, N269);
xor XOR2 (N5186, N5163, N5170);
xor XOR2 (N5187, N4795, N1627);
nor NOR4 (N5188, N5185, N5155, N2636, N515);
nand NAND2 (N5189, N5181, N4232);
not NOT1 (N5190, N5184);
nand NAND2 (N5191, N5188, N4404);
and AND2 (N5192, N5191, N415);
and AND4 (N5193, N5189, N3937, N4156, N4820);
not NOT1 (N5194, N5186);
and AND2 (N5195, N5179, N650);
xor XOR2 (N5196, N5180, N647);
xor XOR2 (N5197, N5190, N997);
and AND2 (N5198, N5195, N4779);
buf BUF1 (N5199, N5192);
not NOT1 (N5200, N5198);
xor XOR2 (N5201, N5197, N4414);
and AND3 (N5202, N5200, N2960, N3318);
and AND4 (N5203, N5199, N2093, N510, N3404);
nor NOR3 (N5204, N5196, N163, N1827);
buf BUF1 (N5205, N5182);
and AND2 (N5206, N5183, N1304);
not NOT1 (N5207, N5205);
buf BUF1 (N5208, N5206);
and AND4 (N5209, N5194, N2358, N3793, N839);
and AND3 (N5210, N5207, N3993, N3386);
not NOT1 (N5211, N5187);
or OR3 (N5212, N5208, N2064, N5207);
buf BUF1 (N5213, N5210);
nand NAND2 (N5214, N5213, N3336);
buf BUF1 (N5215, N5193);
nor NOR2 (N5216, N5209, N2862);
nor NOR2 (N5217, N5211, N459);
and AND2 (N5218, N5203, N4356);
nor NOR2 (N5219, N5204, N2738);
nor NOR3 (N5220, N5215, N3634, N2533);
nor NOR3 (N5221, N5212, N1759, N4539);
nand NAND3 (N5222, N5201, N4438, N3372);
or OR3 (N5223, N5218, N3949, N653);
xor XOR2 (N5224, N5222, N3988);
nand NAND4 (N5225, N5223, N2276, N894, N2906);
and AND2 (N5226, N5221, N1301);
buf BUF1 (N5227, N5216);
xor XOR2 (N5228, N5220, N4285);
xor XOR2 (N5229, N5227, N1816);
nand NAND3 (N5230, N5226, N4083, N1100);
buf BUF1 (N5231, N5178);
not NOT1 (N5232, N5228);
nand NAND4 (N5233, N5229, N3977, N3468, N3567);
nand NAND4 (N5234, N5230, N5005, N1826, N1549);
nor NOR4 (N5235, N5224, N3730, N3522, N4556);
and AND4 (N5236, N5231, N4443, N4768, N4883);
nand NAND2 (N5237, N5217, N3791);
xor XOR2 (N5238, N5214, N2227);
not NOT1 (N5239, N5225);
not NOT1 (N5240, N5236);
not NOT1 (N5241, N5232);
nor NOR3 (N5242, N5241, N3185, N464);
xor XOR2 (N5243, N5237, N3485);
or OR2 (N5244, N5233, N1487);
and AND3 (N5245, N5239, N2314, N1509);
xor XOR2 (N5246, N5235, N2538);
buf BUF1 (N5247, N5243);
buf BUF1 (N5248, N5247);
not NOT1 (N5249, N5248);
buf BUF1 (N5250, N5219);
and AND2 (N5251, N5240, N4543);
buf BUF1 (N5252, N5202);
buf BUF1 (N5253, N5251);
buf BUF1 (N5254, N5246);
or OR4 (N5255, N5238, N4291, N4937, N2713);
nand NAND3 (N5256, N5244, N2951, N2974);
nor NOR2 (N5257, N5252, N34);
not NOT1 (N5258, N5257);
or OR4 (N5259, N5242, N1973, N470, N2657);
buf BUF1 (N5260, N5250);
and AND4 (N5261, N5253, N5230, N4236, N1960);
and AND3 (N5262, N5249, N1069, N2393);
not NOT1 (N5263, N5261);
nor NOR2 (N5264, N5259, N4003);
xor XOR2 (N5265, N5255, N4138);
buf BUF1 (N5266, N5260);
nand NAND3 (N5267, N5234, N986, N2249);
xor XOR2 (N5268, N5263, N3376);
buf BUF1 (N5269, N5258);
xor XOR2 (N5270, N5262, N4239);
nand NAND4 (N5271, N5265, N2629, N4316, N354);
xor XOR2 (N5272, N5271, N1922);
nand NAND2 (N5273, N5254, N22);
buf BUF1 (N5274, N5272);
or OR3 (N5275, N5266, N5131, N508);
not NOT1 (N5276, N5256);
nor NOR2 (N5277, N5269, N1284);
xor XOR2 (N5278, N5273, N3913);
nand NAND4 (N5279, N5275, N4827, N4076, N931);
nand NAND3 (N5280, N5278, N2231, N1464);
nor NOR3 (N5281, N5279, N3210, N1632);
nand NAND2 (N5282, N5280, N367);
nand NAND4 (N5283, N5245, N1020, N2612, N3624);
nor NOR2 (N5284, N5268, N1313);
nor NOR4 (N5285, N5270, N187, N3841, N5118);
nor NOR2 (N5286, N5277, N3148);
or OR2 (N5287, N5264, N3508);
xor XOR2 (N5288, N5281, N2912);
nor NOR4 (N5289, N5276, N1451, N3103, N1);
nand NAND2 (N5290, N5284, N4291);
xor XOR2 (N5291, N5287, N4883);
not NOT1 (N5292, N5286);
xor XOR2 (N5293, N5288, N3444);
xor XOR2 (N5294, N5293, N1911);
or OR2 (N5295, N5289, N5240);
nor NOR4 (N5296, N5291, N2126, N3885, N4111);
nor NOR2 (N5297, N5290, N4333);
not NOT1 (N5298, N5283);
not NOT1 (N5299, N5282);
xor XOR2 (N5300, N5299, N3443);
nand NAND4 (N5301, N5295, N648, N2409, N4526);
or OR2 (N5302, N5294, N279);
nor NOR2 (N5303, N5301, N897);
and AND3 (N5304, N5267, N3569, N5017);
buf BUF1 (N5305, N5274);
and AND3 (N5306, N5304, N121, N4687);
or OR4 (N5307, N5303, N4204, N4084, N3832);
nor NOR4 (N5308, N5298, N700, N246, N1900);
not NOT1 (N5309, N5307);
nor NOR2 (N5310, N5297, N1387);
and AND4 (N5311, N5310, N4477, N1318, N668);
or OR3 (N5312, N5305, N5226, N1047);
not NOT1 (N5313, N5311);
xor XOR2 (N5314, N5306, N903);
and AND4 (N5315, N5314, N3072, N3414, N896);
nor NOR4 (N5316, N5296, N4119, N5293, N583);
buf BUF1 (N5317, N5308);
nand NAND3 (N5318, N5316, N1521, N762);
nor NOR4 (N5319, N5313, N3035, N506, N5044);
and AND2 (N5320, N5315, N5122);
and AND3 (N5321, N5318, N3480, N4051);
buf BUF1 (N5322, N5292);
nor NOR2 (N5323, N5312, N4936);
nor NOR3 (N5324, N5322, N5198, N5028);
nor NOR2 (N5325, N5319, N3617);
buf BUF1 (N5326, N5302);
and AND4 (N5327, N5326, N5297, N5165, N1015);
nor NOR4 (N5328, N5327, N4261, N3566, N4441);
buf BUF1 (N5329, N5324);
nand NAND2 (N5330, N5285, N3075);
nand NAND4 (N5331, N5309, N1429, N2924, N4457);
or OR3 (N5332, N5300, N1153, N2672);
buf BUF1 (N5333, N5323);
xor XOR2 (N5334, N5331, N4849);
or OR3 (N5335, N5329, N4570, N1291);
buf BUF1 (N5336, N5333);
xor XOR2 (N5337, N5334, N3082);
nand NAND4 (N5338, N5317, N30, N3773, N1234);
or OR3 (N5339, N5330, N1405, N5125);
and AND3 (N5340, N5325, N2986, N262);
not NOT1 (N5341, N5321);
xor XOR2 (N5342, N5337, N3758);
nand NAND2 (N5343, N5335, N4807);
buf BUF1 (N5344, N5332);
or OR2 (N5345, N5320, N3721);
not NOT1 (N5346, N5328);
buf BUF1 (N5347, N5343);
or OR2 (N5348, N5344, N5328);
and AND3 (N5349, N5339, N1291, N2026);
not NOT1 (N5350, N5346);
nor NOR2 (N5351, N5345, N3671);
nor NOR3 (N5352, N5341, N356, N3310);
nor NOR4 (N5353, N5350, N323, N4928, N3686);
and AND4 (N5354, N5349, N4888, N2880, N1293);
nor NOR2 (N5355, N5354, N1598);
xor XOR2 (N5356, N5352, N3475);
not NOT1 (N5357, N5353);
not NOT1 (N5358, N5357);
and AND2 (N5359, N5336, N4307);
and AND4 (N5360, N5351, N3263, N775, N4419);
nor NOR4 (N5361, N5356, N831, N3762, N2344);
and AND3 (N5362, N5347, N1887, N786);
nor NOR3 (N5363, N5338, N1324, N210);
not NOT1 (N5364, N5355);
nand NAND3 (N5365, N5362, N1374, N1143);
or OR4 (N5366, N5342, N2856, N3638, N1559);
or OR2 (N5367, N5366, N2503);
and AND3 (N5368, N5358, N1499, N1724);
and AND2 (N5369, N5364, N817);
nor NOR4 (N5370, N5368, N2521, N1912, N4563);
nand NAND3 (N5371, N5361, N1832, N2506);
xor XOR2 (N5372, N5348, N3445);
nand NAND3 (N5373, N5365, N3115, N1497);
xor XOR2 (N5374, N5373, N4813);
buf BUF1 (N5375, N5360);
xor XOR2 (N5376, N5367, N1381);
and AND3 (N5377, N5369, N3372, N1138);
and AND3 (N5378, N5374, N2976, N46);
nor NOR3 (N5379, N5340, N4427, N5303);
not NOT1 (N5380, N5359);
and AND2 (N5381, N5379, N497);
xor XOR2 (N5382, N5376, N3140);
nand NAND3 (N5383, N5382, N3954, N4190);
not NOT1 (N5384, N5381);
xor XOR2 (N5385, N5372, N5287);
buf BUF1 (N5386, N5378);
buf BUF1 (N5387, N5380);
nand NAND4 (N5388, N5371, N2568, N198, N4668);
nor NOR4 (N5389, N5375, N4926, N1456, N1837);
buf BUF1 (N5390, N5386);
nand NAND2 (N5391, N5383, N4840);
xor XOR2 (N5392, N5390, N4044);
buf BUF1 (N5393, N5370);
not NOT1 (N5394, N5391);
nand NAND3 (N5395, N5387, N315, N596);
xor XOR2 (N5396, N5395, N1327);
nor NOR2 (N5397, N5384, N5141);
xor XOR2 (N5398, N5377, N4752);
not NOT1 (N5399, N5397);
nor NOR4 (N5400, N5363, N812, N891, N3283);
xor XOR2 (N5401, N5393, N3370);
or OR3 (N5402, N5394, N4709, N1232);
xor XOR2 (N5403, N5388, N119);
or OR3 (N5404, N5396, N4609, N4115);
not NOT1 (N5405, N5389);
not NOT1 (N5406, N5403);
nor NOR4 (N5407, N5398, N1065, N457, N4212);
not NOT1 (N5408, N5399);
or OR3 (N5409, N5405, N219, N836);
not NOT1 (N5410, N5407);
or OR4 (N5411, N5401, N2256, N3164, N2240);
and AND4 (N5412, N5406, N3534, N2892, N5410);
nand NAND3 (N5413, N2291, N1340, N4888);
and AND2 (N5414, N5404, N156);
nand NAND4 (N5415, N5411, N70, N514, N2106);
nand NAND3 (N5416, N5415, N3273, N1648);
and AND3 (N5417, N5413, N1922, N5348);
and AND4 (N5418, N5400, N1144, N1829, N742);
and AND2 (N5419, N5402, N3677);
and AND2 (N5420, N5417, N4755);
xor XOR2 (N5421, N5392, N2296);
and AND3 (N5422, N5418, N337, N4117);
or OR2 (N5423, N5419, N4536);
or OR3 (N5424, N5409, N2031, N2311);
buf BUF1 (N5425, N5416);
and AND4 (N5426, N5408, N3228, N1421, N4957);
buf BUF1 (N5427, N5422);
and AND3 (N5428, N5427, N5, N818);
xor XOR2 (N5429, N5421, N4540);
nand NAND4 (N5430, N5385, N5035, N1611, N5063);
buf BUF1 (N5431, N5414);
xor XOR2 (N5432, N5429, N2179);
or OR3 (N5433, N5428, N4504, N4636);
and AND4 (N5434, N5425, N4782, N4410, N4682);
or OR4 (N5435, N5423, N3762, N4837, N4050);
nor NOR4 (N5436, N5433, N2432, N1929, N4157);
or OR2 (N5437, N5431, N5010);
nand NAND3 (N5438, N5424, N2129, N3847);
buf BUF1 (N5439, N5420);
nand NAND2 (N5440, N5437, N2073);
nor NOR3 (N5441, N5430, N4867, N1359);
nand NAND3 (N5442, N5440, N476, N1211);
xor XOR2 (N5443, N5412, N221);
nor NOR3 (N5444, N5426, N884, N1705);
not NOT1 (N5445, N5444);
and AND3 (N5446, N5441, N4396, N2068);
and AND4 (N5447, N5446, N404, N3709, N2058);
xor XOR2 (N5448, N5447, N651);
buf BUF1 (N5449, N5432);
or OR2 (N5450, N5448, N3678);
or OR2 (N5451, N5443, N4661);
nor NOR3 (N5452, N5445, N1081, N1051);
buf BUF1 (N5453, N5438);
or OR2 (N5454, N5435, N3484);
buf BUF1 (N5455, N5434);
nor NOR4 (N5456, N5452, N2577, N2524, N1936);
xor XOR2 (N5457, N5436, N2185);
not NOT1 (N5458, N5450);
xor XOR2 (N5459, N5442, N3244);
xor XOR2 (N5460, N5453, N44);
buf BUF1 (N5461, N5457);
xor XOR2 (N5462, N5460, N5137);
not NOT1 (N5463, N5456);
xor XOR2 (N5464, N5449, N801);
not NOT1 (N5465, N5463);
not NOT1 (N5466, N5439);
or OR4 (N5467, N5465, N3158, N3835, N2078);
buf BUF1 (N5468, N5467);
or OR2 (N5469, N5462, N3637);
buf BUF1 (N5470, N5458);
buf BUF1 (N5471, N5468);
not NOT1 (N5472, N5451);
and AND3 (N5473, N5471, N4457, N814);
xor XOR2 (N5474, N5469, N2631);
not NOT1 (N5475, N5474);
or OR4 (N5476, N5464, N524, N1188, N4280);
nand NAND4 (N5477, N5454, N4975, N711, N252);
nand NAND3 (N5478, N5472, N5130, N4233);
xor XOR2 (N5479, N5478, N3039);
xor XOR2 (N5480, N5459, N1432);
buf BUF1 (N5481, N5475);
xor XOR2 (N5482, N5480, N260);
and AND4 (N5483, N5473, N976, N281, N1003);
and AND3 (N5484, N5476, N5313, N4420);
buf BUF1 (N5485, N5470);
xor XOR2 (N5486, N5461, N1137);
xor XOR2 (N5487, N5455, N1594);
nand NAND4 (N5488, N5479, N333, N1836, N3294);
xor XOR2 (N5489, N5481, N2926);
or OR4 (N5490, N5482, N2337, N1674, N5076);
and AND3 (N5491, N5484, N267, N1170);
not NOT1 (N5492, N5491);
nand NAND2 (N5493, N5486, N3768);
xor XOR2 (N5494, N5490, N1995);
nor NOR2 (N5495, N5488, N4482);
nand NAND4 (N5496, N5494, N1914, N58, N1678);
nand NAND4 (N5497, N5495, N3940, N3251, N2889);
buf BUF1 (N5498, N5485);
xor XOR2 (N5499, N5492, N2209);
buf BUF1 (N5500, N5487);
not NOT1 (N5501, N5498);
and AND2 (N5502, N5496, N1220);
or OR4 (N5503, N5500, N2553, N4423, N2542);
nor NOR2 (N5504, N5502, N2791);
buf BUF1 (N5505, N5466);
or OR2 (N5506, N5505, N3441);
nor NOR3 (N5507, N5503, N4794, N2386);
buf BUF1 (N5508, N5507);
nor NOR3 (N5509, N5504, N1602, N3773);
nand NAND4 (N5510, N5483, N3109, N2657, N1615);
and AND3 (N5511, N5506, N1616, N2973);
or OR3 (N5512, N5489, N3705, N1511);
nand NAND4 (N5513, N5499, N1976, N4872, N4361);
buf BUF1 (N5514, N5513);
or OR2 (N5515, N5511, N393);
buf BUF1 (N5516, N5493);
nor NOR2 (N5517, N5512, N1723);
nor NOR4 (N5518, N5477, N3038, N2138, N1594);
or OR4 (N5519, N5517, N3785, N2192, N1816);
and AND4 (N5520, N5501, N2329, N3952, N4686);
buf BUF1 (N5521, N5497);
not NOT1 (N5522, N5519);
nand NAND3 (N5523, N5521, N2815, N3333);
and AND2 (N5524, N5518, N958);
not NOT1 (N5525, N5516);
buf BUF1 (N5526, N5525);
or OR2 (N5527, N5526, N4690);
not NOT1 (N5528, N5520);
not NOT1 (N5529, N5524);
and AND3 (N5530, N5523, N553, N3533);
nor NOR2 (N5531, N5528, N615);
or OR2 (N5532, N5527, N2784);
and AND4 (N5533, N5515, N4682, N1193, N196);
buf BUF1 (N5534, N5533);
nand NAND2 (N5535, N5531, N2179);
and AND2 (N5536, N5535, N4757);
nor NOR2 (N5537, N5530, N3568);
xor XOR2 (N5538, N5532, N4167);
not NOT1 (N5539, N5534);
nand NAND2 (N5540, N5510, N3303);
xor XOR2 (N5541, N5536, N4657);
not NOT1 (N5542, N5539);
or OR4 (N5543, N5529, N5266, N802, N4718);
or OR4 (N5544, N5542, N3618, N4811, N147);
buf BUF1 (N5545, N5537);
or OR4 (N5546, N5540, N5179, N1496, N2672);
not NOT1 (N5547, N5541);
xor XOR2 (N5548, N5544, N3449);
nor NOR4 (N5549, N5547, N4055, N2736, N2313);
nand NAND3 (N5550, N5538, N1772, N5481);
buf BUF1 (N5551, N5548);
nor NOR2 (N5552, N5550, N2186);
xor XOR2 (N5553, N5509, N1519);
and AND2 (N5554, N5553, N1528);
buf BUF1 (N5555, N5514);
not NOT1 (N5556, N5549);
xor XOR2 (N5557, N5552, N2729);
buf BUF1 (N5558, N5546);
and AND3 (N5559, N5508, N4013, N4332);
nor NOR2 (N5560, N5543, N4024);
nor NOR3 (N5561, N5560, N2169, N1395);
nand NAND4 (N5562, N5551, N693, N2890, N795);
xor XOR2 (N5563, N5545, N3214);
or OR4 (N5564, N5559, N5348, N1238, N3178);
nand NAND2 (N5565, N5554, N1035);
buf BUF1 (N5566, N5558);
not NOT1 (N5567, N5564);
not NOT1 (N5568, N5563);
nand NAND2 (N5569, N5561, N4685);
nand NAND3 (N5570, N5522, N5073, N2757);
and AND2 (N5571, N5567, N2931);
nor NOR2 (N5572, N5566, N765);
nand NAND4 (N5573, N5568, N5098, N2012, N1523);
xor XOR2 (N5574, N5556, N3576);
buf BUF1 (N5575, N5557);
nor NOR2 (N5576, N5573, N2848);
nor NOR3 (N5577, N5565, N707, N3435);
buf BUF1 (N5578, N5572);
or OR3 (N5579, N5574, N1185, N30);
buf BUF1 (N5580, N5575);
nor NOR4 (N5581, N5578, N2658, N3968, N3764);
not NOT1 (N5582, N5562);
nand NAND3 (N5583, N5571, N4582, N1707);
buf BUF1 (N5584, N5577);
nor NOR4 (N5585, N5584, N3419, N1656, N1209);
not NOT1 (N5586, N5582);
xor XOR2 (N5587, N5583, N5038);
not NOT1 (N5588, N5586);
buf BUF1 (N5589, N5569);
and AND2 (N5590, N5580, N771);
or OR4 (N5591, N5585, N3623, N1769, N1164);
and AND4 (N5592, N5576, N2028, N3117, N4571);
and AND4 (N5593, N5570, N3451, N1771, N223);
xor XOR2 (N5594, N5587, N4802);
nand NAND4 (N5595, N5555, N1936, N1785, N3590);
or OR3 (N5596, N5581, N775, N111);
xor XOR2 (N5597, N5595, N3828);
and AND2 (N5598, N5594, N3600);
not NOT1 (N5599, N5592);
and AND3 (N5600, N5589, N1405, N1199);
or OR4 (N5601, N5599, N3629, N4247, N2647);
nor NOR3 (N5602, N5598, N1113, N2769);
not NOT1 (N5603, N5588);
buf BUF1 (N5604, N5593);
or OR2 (N5605, N5601, N519);
not NOT1 (N5606, N5603);
buf BUF1 (N5607, N5605);
nor NOR4 (N5608, N5600, N546, N3480, N1363);
not NOT1 (N5609, N5604);
not NOT1 (N5610, N5606);
buf BUF1 (N5611, N5602);
nand NAND2 (N5612, N5590, N245);
or OR4 (N5613, N5609, N897, N2822, N5315);
nand NAND4 (N5614, N5591, N244, N101, N3540);
buf BUF1 (N5615, N5610);
nand NAND3 (N5616, N5607, N2709, N1385);
nand NAND4 (N5617, N5579, N3447, N1967, N1820);
and AND3 (N5618, N5614, N1724, N2351);
or OR4 (N5619, N5611, N229, N223, N232);
and AND4 (N5620, N5615, N284, N1958, N2720);
and AND4 (N5621, N5597, N4116, N5467, N3525);
nand NAND4 (N5622, N5613, N5605, N350, N1198);
or OR3 (N5623, N5621, N5109, N4020);
xor XOR2 (N5624, N5620, N616);
and AND3 (N5625, N5623, N4277, N1143);
and AND2 (N5626, N5596, N2874);
nand NAND3 (N5627, N5625, N5335, N5574);
not NOT1 (N5628, N5622);
or OR2 (N5629, N5618, N3511);
not NOT1 (N5630, N5617);
nand NAND2 (N5631, N5612, N3958);
not NOT1 (N5632, N5608);
nor NOR3 (N5633, N5631, N2597, N1355);
xor XOR2 (N5634, N5627, N5254);
not NOT1 (N5635, N5628);
nand NAND4 (N5636, N5633, N2068, N3295, N667);
not NOT1 (N5637, N5626);
nand NAND2 (N5638, N5632, N5044);
nor NOR3 (N5639, N5636, N4622, N3274);
nand NAND2 (N5640, N5629, N1046);
not NOT1 (N5641, N5640);
not NOT1 (N5642, N5619);
and AND2 (N5643, N5638, N26);
not NOT1 (N5644, N5616);
or OR3 (N5645, N5644, N288, N1727);
xor XOR2 (N5646, N5643, N1165);
and AND3 (N5647, N5630, N4541, N115);
buf BUF1 (N5648, N5634);
nand NAND3 (N5649, N5648, N2652, N2269);
buf BUF1 (N5650, N5647);
buf BUF1 (N5651, N5646);
not NOT1 (N5652, N5624);
or OR4 (N5653, N5652, N4458, N3331, N1210);
nor NOR4 (N5654, N5642, N340, N2019, N3977);
and AND2 (N5655, N5649, N3386);
or OR3 (N5656, N5651, N180, N3525);
not NOT1 (N5657, N5639);
xor XOR2 (N5658, N5635, N3000);
nor NOR2 (N5659, N5645, N939);
nor NOR2 (N5660, N5657, N3011);
xor XOR2 (N5661, N5654, N2401);
xor XOR2 (N5662, N5655, N2146);
xor XOR2 (N5663, N5650, N260);
xor XOR2 (N5664, N5659, N183);
not NOT1 (N5665, N5656);
not NOT1 (N5666, N5658);
and AND3 (N5667, N5660, N2784, N2948);
xor XOR2 (N5668, N5666, N325);
or OR4 (N5669, N5637, N4583, N3522, N3306);
nand NAND4 (N5670, N5665, N1882, N4933, N951);
xor XOR2 (N5671, N5667, N887);
not NOT1 (N5672, N5670);
nand NAND3 (N5673, N5661, N2943, N3114);
buf BUF1 (N5674, N5673);
nor NOR4 (N5675, N5662, N250, N5620, N1874);
buf BUF1 (N5676, N5675);
and AND2 (N5677, N5676, N1007);
nand NAND3 (N5678, N5668, N3071, N4001);
and AND3 (N5679, N5663, N3215, N4643);
xor XOR2 (N5680, N5678, N3870);
and AND4 (N5681, N5653, N1230, N2713, N3881);
nand NAND4 (N5682, N5641, N4208, N1733, N5352);
buf BUF1 (N5683, N5669);
not NOT1 (N5684, N5683);
or OR2 (N5685, N5684, N4207);
buf BUF1 (N5686, N5680);
or OR4 (N5687, N5682, N1326, N383, N2604);
buf BUF1 (N5688, N5674);
nand NAND4 (N5689, N5686, N5240, N5549, N3757);
or OR2 (N5690, N5679, N332);
not NOT1 (N5691, N5681);
buf BUF1 (N5692, N5687);
and AND3 (N5693, N5689, N2241, N1877);
not NOT1 (N5694, N5664);
or OR2 (N5695, N5693, N4676);
nand NAND2 (N5696, N5677, N4934);
nand NAND2 (N5697, N5671, N1689);
nor NOR4 (N5698, N5685, N3062, N980, N4747);
and AND3 (N5699, N5697, N2910, N1571);
not NOT1 (N5700, N5692);
xor XOR2 (N5701, N5700, N1467);
and AND2 (N5702, N5701, N3782);
or OR4 (N5703, N5702, N4269, N5251, N629);
or OR4 (N5704, N5691, N2448, N2784, N5370);
nor NOR2 (N5705, N5698, N3076);
and AND2 (N5706, N5688, N4516);
nand NAND4 (N5707, N5695, N941, N1170, N3473);
nand NAND2 (N5708, N5690, N5128);
or OR3 (N5709, N5703, N3901, N5550);
xor XOR2 (N5710, N5672, N3599);
or OR4 (N5711, N5710, N1075, N2606, N916);
buf BUF1 (N5712, N5699);
and AND3 (N5713, N5694, N448, N5099);
nor NOR3 (N5714, N5713, N31, N4649);
and AND3 (N5715, N5712, N3107, N4640);
nand NAND2 (N5716, N5715, N2640);
xor XOR2 (N5717, N5714, N4331);
buf BUF1 (N5718, N5716);
nand NAND2 (N5719, N5718, N1140);
not NOT1 (N5720, N5708);
not NOT1 (N5721, N5709);
buf BUF1 (N5722, N5720);
not NOT1 (N5723, N5696);
xor XOR2 (N5724, N5721, N4908);
not NOT1 (N5725, N5705);
nor NOR2 (N5726, N5711, N5170);
and AND2 (N5727, N5707, N3724);
or OR3 (N5728, N5704, N2781, N99);
nand NAND3 (N5729, N5719, N4507, N3290);
xor XOR2 (N5730, N5706, N1320);
buf BUF1 (N5731, N5722);
not NOT1 (N5732, N5724);
nor NOR3 (N5733, N5729, N48, N2965);
buf BUF1 (N5734, N5731);
nand NAND3 (N5735, N5725, N1794, N3928);
nand NAND2 (N5736, N5727, N4454);
xor XOR2 (N5737, N5726, N2950);
buf BUF1 (N5738, N5735);
xor XOR2 (N5739, N5732, N1074);
and AND3 (N5740, N5733, N3339, N300);
and AND2 (N5741, N5737, N3934);
nand NAND3 (N5742, N5728, N382, N488);
buf BUF1 (N5743, N5742);
buf BUF1 (N5744, N5743);
and AND4 (N5745, N5730, N4797, N1775, N3807);
buf BUF1 (N5746, N5723);
nand NAND3 (N5747, N5741, N2911, N2188);
or OR2 (N5748, N5738, N635);
not NOT1 (N5749, N5748);
or OR2 (N5750, N5739, N3528);
xor XOR2 (N5751, N5736, N3527);
nand NAND3 (N5752, N5734, N1726, N3560);
or OR2 (N5753, N5749, N669);
nand NAND4 (N5754, N5717, N2475, N249, N2849);
and AND4 (N5755, N5753, N239, N3931, N2355);
nand NAND3 (N5756, N5752, N3130, N900);
or OR4 (N5757, N5755, N2830, N4685, N4076);
xor XOR2 (N5758, N5747, N425);
or OR4 (N5759, N5740, N1376, N4, N3216);
xor XOR2 (N5760, N5756, N3425);
nor NOR4 (N5761, N5750, N2232, N3148, N3448);
not NOT1 (N5762, N5745);
and AND2 (N5763, N5761, N4709);
nor NOR3 (N5764, N5746, N5135, N1881);
or OR2 (N5765, N5754, N3841);
or OR4 (N5766, N5758, N4413, N3530, N535);
not NOT1 (N5767, N5764);
not NOT1 (N5768, N5760);
nand NAND2 (N5769, N5762, N3479);
and AND3 (N5770, N5765, N1117, N840);
or OR2 (N5771, N5768, N3293);
and AND2 (N5772, N5766, N87);
nor NOR3 (N5773, N5757, N5646, N3784);
xor XOR2 (N5774, N5770, N2398);
buf BUF1 (N5775, N5759);
and AND2 (N5776, N5767, N809);
and AND2 (N5777, N5774, N578);
xor XOR2 (N5778, N5763, N2057);
nand NAND2 (N5779, N5776, N5183);
xor XOR2 (N5780, N5751, N86);
nand NAND3 (N5781, N5778, N2075, N4209);
and AND4 (N5782, N5780, N3359, N1304, N2308);
and AND3 (N5783, N5772, N1969, N2659);
nor NOR3 (N5784, N5775, N2465, N2867);
nand NAND2 (N5785, N5777, N2811);
nand NAND4 (N5786, N5771, N4099, N3158, N3076);
nor NOR3 (N5787, N5781, N5314, N5024);
nand NAND2 (N5788, N5769, N1478);
xor XOR2 (N5789, N5782, N5034);
not NOT1 (N5790, N5786);
xor XOR2 (N5791, N5784, N3348);
nor NOR2 (N5792, N5790, N4267);
buf BUF1 (N5793, N5788);
xor XOR2 (N5794, N5785, N2734);
nor NOR2 (N5795, N5787, N3462);
xor XOR2 (N5796, N5773, N1257);
not NOT1 (N5797, N5793);
or OR4 (N5798, N5783, N5518, N780, N4707);
nor NOR2 (N5799, N5798, N27);
buf BUF1 (N5800, N5792);
xor XOR2 (N5801, N5744, N1487);
nand NAND2 (N5802, N5779, N5599);
xor XOR2 (N5803, N5791, N1371);
xor XOR2 (N5804, N5796, N3311);
not NOT1 (N5805, N5803);
nand NAND2 (N5806, N5789, N2826);
or OR3 (N5807, N5794, N1693, N503);
buf BUF1 (N5808, N5806);
buf BUF1 (N5809, N5799);
nand NAND4 (N5810, N5807, N2450, N4505, N3293);
nand NAND4 (N5811, N5805, N4026, N750, N2255);
xor XOR2 (N5812, N5802, N4670);
buf BUF1 (N5813, N5809);
buf BUF1 (N5814, N5808);
nand NAND3 (N5815, N5800, N3200, N4739);
nor NOR2 (N5816, N5811, N1739);
xor XOR2 (N5817, N5801, N1427);
nor NOR2 (N5818, N5816, N1766);
not NOT1 (N5819, N5812);
buf BUF1 (N5820, N5815);
nand NAND3 (N5821, N5813, N283, N4109);
not NOT1 (N5822, N5795);
xor XOR2 (N5823, N5817, N2249);
and AND4 (N5824, N5821, N4952, N2208, N4385);
buf BUF1 (N5825, N5824);
xor XOR2 (N5826, N5797, N1676);
buf BUF1 (N5827, N5810);
not NOT1 (N5828, N5827);
or OR2 (N5829, N5820, N4910);
nand NAND4 (N5830, N5822, N1123, N3518, N129);
not NOT1 (N5831, N5814);
xor XOR2 (N5832, N5829, N5324);
and AND3 (N5833, N5831, N2225, N432);
buf BUF1 (N5834, N5825);
and AND3 (N5835, N5819, N1631, N3062);
nand NAND2 (N5836, N5818, N1012);
not NOT1 (N5837, N5836);
nor NOR4 (N5838, N5826, N2061, N710, N4890);
and AND3 (N5839, N5834, N4099, N2676);
not NOT1 (N5840, N5823);
not NOT1 (N5841, N5830);
not NOT1 (N5842, N5828);
and AND2 (N5843, N5840, N3320);
nand NAND3 (N5844, N5842, N2784, N2306);
nor NOR4 (N5845, N5833, N72, N1191, N4820);
xor XOR2 (N5846, N5838, N63);
nand NAND4 (N5847, N5835, N5773, N283, N2604);
xor XOR2 (N5848, N5843, N173);
and AND2 (N5849, N5832, N2175);
and AND3 (N5850, N5841, N5595, N1449);
nor NOR4 (N5851, N5846, N794, N1452, N3045);
xor XOR2 (N5852, N5847, N1547);
not NOT1 (N5853, N5839);
or OR4 (N5854, N5851, N2707, N1214, N3992);
not NOT1 (N5855, N5848);
nand NAND2 (N5856, N5852, N4664);
nand NAND2 (N5857, N5849, N3324);
nor NOR4 (N5858, N5855, N353, N5808, N2444);
xor XOR2 (N5859, N5850, N2035);
nand NAND2 (N5860, N5857, N273);
buf BUF1 (N5861, N5860);
xor XOR2 (N5862, N5861, N828);
or OR3 (N5863, N5858, N4745, N357);
not NOT1 (N5864, N5844);
and AND3 (N5865, N5804, N59, N1432);
nand NAND2 (N5866, N5845, N317);
xor XOR2 (N5867, N5864, N5806);
xor XOR2 (N5868, N5862, N4666);
buf BUF1 (N5869, N5863);
xor XOR2 (N5870, N5856, N5571);
nand NAND2 (N5871, N5869, N5183);
or OR2 (N5872, N5866, N5090);
or OR3 (N5873, N5867, N1850, N4487);
buf BUF1 (N5874, N5853);
not NOT1 (N5875, N5870);
nor NOR4 (N5876, N5875, N4789, N4916, N2176);
buf BUF1 (N5877, N5876);
or OR4 (N5878, N5873, N550, N4330, N4835);
nand NAND3 (N5879, N5854, N2027, N41);
xor XOR2 (N5880, N5879, N5320);
nor NOR4 (N5881, N5877, N1349, N3359, N3758);
or OR3 (N5882, N5878, N5047, N5618);
buf BUF1 (N5883, N5865);
and AND3 (N5884, N5871, N2412, N2261);
not NOT1 (N5885, N5874);
or OR4 (N5886, N5868, N4768, N821, N1416);
or OR3 (N5887, N5882, N2159, N1202);
or OR2 (N5888, N5885, N3974);
or OR3 (N5889, N5881, N5050, N2939);
buf BUF1 (N5890, N5883);
buf BUF1 (N5891, N5889);
nor NOR3 (N5892, N5880, N1972, N109);
nor NOR3 (N5893, N5890, N3814, N5374);
nand NAND4 (N5894, N5887, N2234, N2969, N2144);
nor NOR2 (N5895, N5872, N5625);
or OR2 (N5896, N5891, N4294);
xor XOR2 (N5897, N5859, N5719);
nand NAND2 (N5898, N5895, N2332);
or OR3 (N5899, N5892, N312, N4675);
buf BUF1 (N5900, N5897);
buf BUF1 (N5901, N5894);
not NOT1 (N5902, N5893);
nand NAND2 (N5903, N5901, N778);
and AND2 (N5904, N5837, N2467);
xor XOR2 (N5905, N5898, N2067);
and AND4 (N5906, N5888, N2095, N4828, N221);
not NOT1 (N5907, N5905);
xor XOR2 (N5908, N5900, N3251);
not NOT1 (N5909, N5903);
buf BUF1 (N5910, N5899);
or OR4 (N5911, N5908, N4113, N1973, N395);
buf BUF1 (N5912, N5907);
buf BUF1 (N5913, N5904);
buf BUF1 (N5914, N5906);
not NOT1 (N5915, N5912);
and AND3 (N5916, N5884, N3634, N3521);
nor NOR3 (N5917, N5902, N3826, N1139);
xor XOR2 (N5918, N5910, N1924);
and AND4 (N5919, N5913, N3522, N4330, N5728);
xor XOR2 (N5920, N5918, N810);
and AND4 (N5921, N5911, N3824, N592, N565);
xor XOR2 (N5922, N5916, N5416);
buf BUF1 (N5923, N5896);
xor XOR2 (N5924, N5921, N2482);
nor NOR3 (N5925, N5886, N1940, N1122);
not NOT1 (N5926, N5920);
buf BUF1 (N5927, N5914);
xor XOR2 (N5928, N5927, N5507);
xor XOR2 (N5929, N5926, N388);
not NOT1 (N5930, N5923);
not NOT1 (N5931, N5919);
or OR4 (N5932, N5928, N4819, N2228, N3862);
and AND2 (N5933, N5931, N1897);
or OR3 (N5934, N5909, N355, N2862);
buf BUF1 (N5935, N5930);
not NOT1 (N5936, N5925);
and AND3 (N5937, N5934, N4953, N3472);
nand NAND2 (N5938, N5932, N3942);
xor XOR2 (N5939, N5937, N2578);
xor XOR2 (N5940, N5917, N1807);
or OR3 (N5941, N5933, N5710, N4995);
or OR2 (N5942, N5915, N4321);
nor NOR2 (N5943, N5940, N852);
and AND2 (N5944, N5942, N2183);
buf BUF1 (N5945, N5938);
or OR2 (N5946, N5922, N4799);
and AND4 (N5947, N5944, N3282, N903, N1310);
nor NOR4 (N5948, N5924, N4104, N5017, N5831);
and AND2 (N5949, N5945, N2314);
nor NOR2 (N5950, N5936, N1048);
nor NOR2 (N5951, N5929, N1568);
not NOT1 (N5952, N5950);
not NOT1 (N5953, N5947);
xor XOR2 (N5954, N5951, N3884);
nand NAND2 (N5955, N5948, N4912);
and AND3 (N5956, N5949, N3042, N1917);
or OR2 (N5957, N5941, N4498);
nand NAND3 (N5958, N5957, N5743, N2394);
buf BUF1 (N5959, N5955);
buf BUF1 (N5960, N5939);
and AND2 (N5961, N5943, N1896);
or OR2 (N5962, N5959, N89);
xor XOR2 (N5963, N5958, N3883);
buf BUF1 (N5964, N5962);
nand NAND3 (N5965, N5961, N2630, N4103);
nor NOR4 (N5966, N5965, N972, N4009, N5843);
not NOT1 (N5967, N5963);
nor NOR3 (N5968, N5960, N619, N4805);
not NOT1 (N5969, N5935);
or OR4 (N5970, N5952, N4903, N3912, N1390);
and AND2 (N5971, N5970, N3428);
or OR4 (N5972, N5954, N2410, N5412, N2281);
nand NAND3 (N5973, N5964, N2406, N4184);
or OR4 (N5974, N5953, N5767, N374, N5920);
xor XOR2 (N5975, N5966, N4833);
buf BUF1 (N5976, N5972);
nor NOR3 (N5977, N5969, N2225, N4214);
or OR4 (N5978, N5967, N4494, N4998, N3765);
and AND4 (N5979, N5974, N5159, N3119, N2205);
xor XOR2 (N5980, N5976, N1373);
buf BUF1 (N5981, N5973);
nand NAND4 (N5982, N5980, N5188, N4197, N720);
and AND2 (N5983, N5978, N3195);
xor XOR2 (N5984, N5983, N1468);
and AND3 (N5985, N5984, N5359, N5188);
buf BUF1 (N5986, N5968);
or OR2 (N5987, N5971, N864);
nor NOR2 (N5988, N5946, N4279);
xor XOR2 (N5989, N5977, N5735);
xor XOR2 (N5990, N5956, N2614);
nand NAND3 (N5991, N5986, N202, N2907);
nor NOR4 (N5992, N5989, N4966, N1252, N5061);
xor XOR2 (N5993, N5985, N2189);
xor XOR2 (N5994, N5982, N1187);
not NOT1 (N5995, N5987);
xor XOR2 (N5996, N5991, N5638);
and AND2 (N5997, N5988, N5397);
buf BUF1 (N5998, N5990);
not NOT1 (N5999, N5998);
nand NAND2 (N6000, N5981, N4797);
buf BUF1 (N6001, N5994);
nand NAND3 (N6002, N5996, N4638, N5511);
and AND2 (N6003, N5995, N2543);
xor XOR2 (N6004, N6002, N3349);
or OR4 (N6005, N5975, N1820, N4184, N1783);
buf BUF1 (N6006, N5997);
and AND3 (N6007, N6004, N3346, N4763);
or OR4 (N6008, N5979, N4428, N2531, N1877);
not NOT1 (N6009, N6008);
xor XOR2 (N6010, N6007, N3499);
or OR4 (N6011, N5992, N5850, N2414, N3957);
not NOT1 (N6012, N6000);
xor XOR2 (N6013, N5993, N5044);
or OR3 (N6014, N6006, N1292, N3420);
buf BUF1 (N6015, N6012);
nand NAND4 (N6016, N6011, N838, N4436, N5922);
or OR4 (N6017, N6016, N5090, N3560, N713);
buf BUF1 (N6018, N6015);
xor XOR2 (N6019, N6005, N1774);
xor XOR2 (N6020, N5999, N2068);
nor NOR4 (N6021, N6003, N4952, N3372, N3779);
nand NAND3 (N6022, N6019, N4155, N4271);
buf BUF1 (N6023, N6021);
nor NOR4 (N6024, N6022, N5745, N2340, N4610);
nor NOR3 (N6025, N6013, N5641, N4925);
buf BUF1 (N6026, N6014);
buf BUF1 (N6027, N6025);
and AND2 (N6028, N6026, N1392);
nand NAND3 (N6029, N6028, N4595, N3051);
and AND2 (N6030, N6001, N3511);
not NOT1 (N6031, N6030);
nand NAND2 (N6032, N6018, N3177);
or OR3 (N6033, N6029, N3511, N3201);
buf BUF1 (N6034, N6031);
and AND4 (N6035, N6010, N4208, N1591, N1190);
xor XOR2 (N6036, N6009, N3003);
nor NOR4 (N6037, N6034, N3821, N5091, N4035);
xor XOR2 (N6038, N6035, N4977);
nor NOR4 (N6039, N6033, N1478, N5438, N5295);
xor XOR2 (N6040, N6037, N1347);
nor NOR4 (N6041, N6036, N5354, N5016, N1656);
buf BUF1 (N6042, N6038);
xor XOR2 (N6043, N6024, N5050);
or OR2 (N6044, N6040, N5286);
not NOT1 (N6045, N6032);
buf BUF1 (N6046, N6020);
not NOT1 (N6047, N6023);
xor XOR2 (N6048, N6042, N3650);
xor XOR2 (N6049, N6046, N3941);
xor XOR2 (N6050, N6027, N478);
nand NAND4 (N6051, N6044, N5274, N3944, N3456);
xor XOR2 (N6052, N6039, N111);
or OR2 (N6053, N6051, N2288);
or OR3 (N6054, N6041, N2054, N5225);
xor XOR2 (N6055, N6045, N1288);
nand NAND4 (N6056, N6043, N4270, N3826, N2823);
or OR4 (N6057, N6050, N966, N2622, N4024);
or OR2 (N6058, N6053, N494);
nand NAND2 (N6059, N6049, N3080);
nand NAND4 (N6060, N6057, N4477, N976, N2215);
nand NAND3 (N6061, N6017, N1113, N3802);
nand NAND2 (N6062, N6060, N3152);
or OR4 (N6063, N6061, N2887, N5713, N2033);
xor XOR2 (N6064, N6062, N2237);
not NOT1 (N6065, N6047);
xor XOR2 (N6066, N6065, N1409);
nor NOR2 (N6067, N6052, N2382);
buf BUF1 (N6068, N6048);
or OR2 (N6069, N6066, N2125);
not NOT1 (N6070, N6056);
nor NOR2 (N6071, N6058, N4281);
not NOT1 (N6072, N6069);
buf BUF1 (N6073, N6070);
not NOT1 (N6074, N6059);
buf BUF1 (N6075, N6074);
or OR2 (N6076, N6054, N3266);
or OR2 (N6077, N6075, N4759);
xor XOR2 (N6078, N6071, N5578);
nor NOR4 (N6079, N6063, N3716, N73, N5182);
and AND4 (N6080, N6076, N5899, N899, N3928);
nor NOR3 (N6081, N6072, N5304, N5941);
not NOT1 (N6082, N6068);
xor XOR2 (N6083, N6079, N3657);
and AND4 (N6084, N6078, N568, N3163, N1782);
or OR3 (N6085, N6082, N4782, N5961);
nor NOR4 (N6086, N6081, N5062, N2090, N5427);
nand NAND4 (N6087, N6085, N3580, N864, N1654);
or OR2 (N6088, N6064, N2598);
and AND4 (N6089, N6087, N2272, N4517, N1086);
nor NOR4 (N6090, N6080, N2489, N124, N2614);
and AND3 (N6091, N6077, N5862, N1415);
not NOT1 (N6092, N6073);
and AND2 (N6093, N6088, N3733);
not NOT1 (N6094, N6083);
and AND2 (N6095, N6094, N4408);
xor XOR2 (N6096, N6093, N5961);
nand NAND4 (N6097, N6090, N1206, N5936, N4773);
nand NAND4 (N6098, N6086, N4264, N4862, N3708);
buf BUF1 (N6099, N6097);
not NOT1 (N6100, N6055);
or OR4 (N6101, N6100, N3372, N1914, N3098);
or OR3 (N6102, N6084, N4297, N4427);
not NOT1 (N6103, N6092);
and AND4 (N6104, N6103, N2048, N2361, N5210);
and AND2 (N6105, N6096, N2276);
nand NAND3 (N6106, N6102, N598, N5838);
xor XOR2 (N6107, N6089, N2926);
not NOT1 (N6108, N6101);
nand NAND2 (N6109, N6067, N5288);
and AND3 (N6110, N6091, N2288, N2847);
nand NAND4 (N6111, N6109, N2137, N3919, N220);
or OR2 (N6112, N6110, N3052);
or OR4 (N6113, N6099, N2338, N108, N3659);
nor NOR4 (N6114, N6095, N3826, N4208, N2905);
nor NOR3 (N6115, N6107, N5601, N3939);
xor XOR2 (N6116, N6111, N5065);
and AND4 (N6117, N6104, N4611, N2283, N5929);
nand NAND2 (N6118, N6106, N2703);
or OR4 (N6119, N6113, N1600, N662, N3009);
and AND3 (N6120, N6108, N4977, N626);
buf BUF1 (N6121, N6112);
not NOT1 (N6122, N6120);
nand NAND2 (N6123, N6119, N1784);
nor NOR3 (N6124, N6098, N2194, N2222);
or OR4 (N6125, N6105, N2535, N5004, N4852);
or OR2 (N6126, N6122, N2083);
buf BUF1 (N6127, N6117);
or OR4 (N6128, N6124, N5538, N3711, N5253);
xor XOR2 (N6129, N6128, N1789);
or OR4 (N6130, N6114, N2817, N338, N898);
or OR2 (N6131, N6126, N3311);
and AND4 (N6132, N6118, N1799, N1185, N2781);
nand NAND3 (N6133, N6115, N6071, N1229);
nand NAND2 (N6134, N6123, N5088);
nor NOR2 (N6135, N6129, N4559);
buf BUF1 (N6136, N6131);
buf BUF1 (N6137, N6133);
buf BUF1 (N6138, N6132);
nand NAND3 (N6139, N6130, N2432, N3813);
nand NAND2 (N6140, N6127, N5138);
buf BUF1 (N6141, N6137);
and AND2 (N6142, N6125, N3320);
buf BUF1 (N6143, N6136);
or OR3 (N6144, N6134, N2341, N3832);
xor XOR2 (N6145, N6116, N1216);
and AND2 (N6146, N6135, N4737);
xor XOR2 (N6147, N6140, N6105);
nor NOR2 (N6148, N6145, N5560);
buf BUF1 (N6149, N6143);
nor NOR2 (N6150, N6146, N3888);
xor XOR2 (N6151, N6149, N1916);
not NOT1 (N6152, N6144);
nand NAND3 (N6153, N6150, N5396, N4706);
not NOT1 (N6154, N6151);
and AND4 (N6155, N6153, N287, N1279, N4379);
nor NOR3 (N6156, N6154, N6140, N1678);
xor XOR2 (N6157, N6142, N2257);
xor XOR2 (N6158, N6141, N1010);
and AND3 (N6159, N6158, N4120, N1898);
or OR2 (N6160, N6139, N2781);
or OR4 (N6161, N6160, N2010, N5906, N5650);
xor XOR2 (N6162, N6155, N4937);
buf BUF1 (N6163, N6156);
buf BUF1 (N6164, N6152);
and AND3 (N6165, N6164, N3535, N3680);
buf BUF1 (N6166, N6165);
or OR2 (N6167, N6162, N3646);
not NOT1 (N6168, N6157);
nand NAND4 (N6169, N6148, N5490, N753, N2185);
nor NOR3 (N6170, N6161, N62, N2604);
and AND4 (N6171, N6163, N4584, N1843, N4368);
not NOT1 (N6172, N6167);
xor XOR2 (N6173, N6166, N6162);
xor XOR2 (N6174, N6147, N1058);
and AND4 (N6175, N6168, N2643, N2413, N668);
nand NAND4 (N6176, N6172, N5124, N4448, N502);
nand NAND4 (N6177, N6170, N4856, N517, N2662);
buf BUF1 (N6178, N6159);
buf BUF1 (N6179, N6176);
nand NAND4 (N6180, N6174, N5527, N2056, N3489);
not NOT1 (N6181, N6173);
nand NAND3 (N6182, N6121, N3395, N3596);
nand NAND4 (N6183, N6171, N889, N490, N2413);
nor NOR4 (N6184, N6178, N5625, N3697, N3140);
not NOT1 (N6185, N6179);
buf BUF1 (N6186, N6175);
xor XOR2 (N6187, N6182, N663);
xor XOR2 (N6188, N6186, N3770);
buf BUF1 (N6189, N6185);
nand NAND3 (N6190, N6138, N4735, N3898);
xor XOR2 (N6191, N6190, N5667);
or OR4 (N6192, N6177, N659, N5156, N403);
or OR4 (N6193, N6181, N3122, N4648, N5253);
nand NAND4 (N6194, N6183, N5424, N2289, N2215);
or OR3 (N6195, N6187, N1896, N4380);
not NOT1 (N6196, N6189);
nor NOR2 (N6197, N6180, N2373);
buf BUF1 (N6198, N6197);
not NOT1 (N6199, N6194);
nand NAND3 (N6200, N6193, N3519, N4823);
nor NOR2 (N6201, N6196, N4919);
xor XOR2 (N6202, N6192, N1008);
nand NAND3 (N6203, N6191, N3466, N3229);
or OR2 (N6204, N6202, N1560);
not NOT1 (N6205, N6198);
nand NAND4 (N6206, N6195, N5691, N1457, N1601);
buf BUF1 (N6207, N6204);
or OR2 (N6208, N6205, N3753);
buf BUF1 (N6209, N6184);
not NOT1 (N6210, N6207);
nand NAND4 (N6211, N6209, N824, N1039, N4722);
nand NAND2 (N6212, N6203, N1918);
not NOT1 (N6213, N6200);
nor NOR2 (N6214, N6208, N4057);
and AND4 (N6215, N6188, N530, N1567, N5200);
nand NAND3 (N6216, N6212, N2423, N3762);
xor XOR2 (N6217, N6211, N4540);
nand NAND2 (N6218, N6214, N4376);
not NOT1 (N6219, N6201);
xor XOR2 (N6220, N6216, N6162);
buf BUF1 (N6221, N6215);
nor NOR2 (N6222, N6220, N997);
buf BUF1 (N6223, N6199);
nor NOR4 (N6224, N6213, N1987, N2472, N5216);
nor NOR4 (N6225, N6221, N2647, N95, N5324);
xor XOR2 (N6226, N6222, N4734);
nand NAND3 (N6227, N6226, N4890, N6104);
nor NOR2 (N6228, N6225, N4749);
xor XOR2 (N6229, N6227, N2722);
and AND4 (N6230, N6229, N5803, N3550, N5613);
buf BUF1 (N6231, N6219);
not NOT1 (N6232, N6230);
xor XOR2 (N6233, N6218, N752);
or OR3 (N6234, N6206, N946, N3668);
xor XOR2 (N6235, N6224, N3963);
and AND3 (N6236, N6232, N2346, N2372);
buf BUF1 (N6237, N6231);
nor NOR4 (N6238, N6234, N2911, N3812, N5361);
buf BUF1 (N6239, N6223);
not NOT1 (N6240, N6228);
or OR4 (N6241, N6210, N4763, N2871, N840);
buf BUF1 (N6242, N6217);
nor NOR3 (N6243, N6233, N4759, N2496);
and AND2 (N6244, N6237, N5475);
and AND4 (N6245, N6169, N2792, N5632, N5299);
buf BUF1 (N6246, N6245);
buf BUF1 (N6247, N6238);
and AND2 (N6248, N6236, N4372);
xor XOR2 (N6249, N6244, N4249);
buf BUF1 (N6250, N6247);
buf BUF1 (N6251, N6248);
and AND4 (N6252, N6235, N4689, N2762, N4519);
and AND2 (N6253, N6251, N5023);
nor NOR3 (N6254, N6240, N5950, N4669);
not NOT1 (N6255, N6242);
nor NOR4 (N6256, N6255, N3904, N1487, N1864);
xor XOR2 (N6257, N6254, N242);
buf BUF1 (N6258, N6249);
and AND2 (N6259, N6239, N4413);
or OR2 (N6260, N6243, N3942);
and AND4 (N6261, N6258, N3650, N4586, N153);
and AND3 (N6262, N6260, N1845, N2151);
nor NOR2 (N6263, N6250, N741);
nand NAND2 (N6264, N6241, N5729);
or OR4 (N6265, N6261, N1953, N1356, N4530);
buf BUF1 (N6266, N6257);
buf BUF1 (N6267, N6266);
xor XOR2 (N6268, N6267, N2236);
or OR3 (N6269, N6264, N4460, N4331);
xor XOR2 (N6270, N6265, N3600);
nor NOR3 (N6271, N6270, N282, N4684);
xor XOR2 (N6272, N6263, N2763);
not NOT1 (N6273, N6262);
or OR4 (N6274, N6268, N2236, N2696, N1086);
and AND2 (N6275, N6246, N3761);
or OR4 (N6276, N6256, N4062, N2233, N2283);
or OR3 (N6277, N6276, N5105, N2168);
and AND4 (N6278, N6272, N3438, N3044, N5616);
or OR3 (N6279, N6259, N3733, N2734);
not NOT1 (N6280, N6274);
buf BUF1 (N6281, N6252);
not NOT1 (N6282, N6271);
and AND3 (N6283, N6269, N4208, N3196);
not NOT1 (N6284, N6277);
nor NOR4 (N6285, N6253, N1941, N1063, N2813);
or OR2 (N6286, N6283, N5576);
buf BUF1 (N6287, N6286);
or OR2 (N6288, N6280, N571);
or OR2 (N6289, N6288, N5370);
buf BUF1 (N6290, N6289);
buf BUF1 (N6291, N6290);
or OR3 (N6292, N6285, N811, N2639);
and AND3 (N6293, N6273, N1003, N71);
xor XOR2 (N6294, N6284, N544);
nand NAND3 (N6295, N6292, N1147, N1855);
nand NAND2 (N6296, N6279, N5173);
or OR2 (N6297, N6287, N3609);
not NOT1 (N6298, N6293);
buf BUF1 (N6299, N6291);
not NOT1 (N6300, N6296);
nand NAND2 (N6301, N6295, N550);
and AND4 (N6302, N6299, N2716, N2296, N97);
not NOT1 (N6303, N6300);
buf BUF1 (N6304, N6278);
not NOT1 (N6305, N6302);
xor XOR2 (N6306, N6275, N4058);
buf BUF1 (N6307, N6303);
and AND4 (N6308, N6307, N3723, N1766, N1287);
nor NOR4 (N6309, N6297, N5262, N3720, N2833);
xor XOR2 (N6310, N6304, N5094);
nor NOR4 (N6311, N6305, N2657, N4777, N2509);
nand NAND4 (N6312, N6311, N5081, N4384, N267);
not NOT1 (N6313, N6312);
nor NOR4 (N6314, N6298, N5275, N3533, N653);
xor XOR2 (N6315, N6294, N1494);
or OR4 (N6316, N6309, N5745, N2416, N1651);
not NOT1 (N6317, N6282);
or OR4 (N6318, N6301, N4034, N3442, N3878);
nor NOR4 (N6319, N6318, N1292, N4285, N3916);
or OR2 (N6320, N6308, N2223);
nor NOR2 (N6321, N6310, N36);
nand NAND3 (N6322, N6315, N1275, N4830);
or OR4 (N6323, N6320, N5940, N5754, N3330);
and AND3 (N6324, N6313, N5816, N2788);
nand NAND4 (N6325, N6322, N3598, N2558, N5801);
and AND2 (N6326, N6306, N1828);
buf BUF1 (N6327, N6319);
buf BUF1 (N6328, N6324);
not NOT1 (N6329, N6325);
buf BUF1 (N6330, N6321);
xor XOR2 (N6331, N6330, N305);
not NOT1 (N6332, N6317);
buf BUF1 (N6333, N6327);
nor NOR4 (N6334, N6316, N5824, N4343, N1031);
not NOT1 (N6335, N6314);
nand NAND2 (N6336, N6331, N285);
nand NAND4 (N6337, N6323, N4102, N2908, N918);
or OR4 (N6338, N6334, N569, N3530, N6067);
nand NAND4 (N6339, N6326, N2845, N5570, N3762);
buf BUF1 (N6340, N6339);
buf BUF1 (N6341, N6329);
xor XOR2 (N6342, N6328, N199);
xor XOR2 (N6343, N6333, N2251);
and AND4 (N6344, N6336, N2817, N132, N3273);
not NOT1 (N6345, N6344);
xor XOR2 (N6346, N6340, N3839);
not NOT1 (N6347, N6332);
xor XOR2 (N6348, N6337, N1781);
nor NOR4 (N6349, N6341, N3464, N5284, N1269);
and AND3 (N6350, N6338, N3492, N198);
and AND2 (N6351, N6342, N5287);
xor XOR2 (N6352, N6335, N1795);
nand NAND3 (N6353, N6348, N1289, N6191);
not NOT1 (N6354, N6343);
nand NAND3 (N6355, N6281, N3064, N5580);
not NOT1 (N6356, N6354);
and AND3 (N6357, N6345, N2064, N4343);
or OR2 (N6358, N6350, N3603);
and AND4 (N6359, N6353, N3483, N2384, N4761);
or OR3 (N6360, N6349, N295, N518);
buf BUF1 (N6361, N6359);
buf BUF1 (N6362, N6355);
or OR4 (N6363, N6358, N2663, N1640, N559);
or OR4 (N6364, N6356, N3535, N628, N5453);
and AND2 (N6365, N6346, N3613);
xor XOR2 (N6366, N6351, N1883);
nand NAND2 (N6367, N6347, N797);
or OR2 (N6368, N6361, N74);
not NOT1 (N6369, N6360);
xor XOR2 (N6370, N6357, N2057);
and AND3 (N6371, N6362, N2666, N1592);
xor XOR2 (N6372, N6363, N64);
buf BUF1 (N6373, N6368);
xor XOR2 (N6374, N6369, N118);
and AND3 (N6375, N6372, N2268, N4882);
buf BUF1 (N6376, N6364);
not NOT1 (N6377, N6366);
not NOT1 (N6378, N6370);
buf BUF1 (N6379, N6367);
or OR4 (N6380, N6374, N6193, N4420, N1235);
or OR3 (N6381, N6376, N3833, N4893);
not NOT1 (N6382, N6375);
and AND3 (N6383, N6382, N4053, N4150);
and AND4 (N6384, N6373, N4276, N1383, N4230);
xor XOR2 (N6385, N6352, N3208);
buf BUF1 (N6386, N6385);
nor NOR3 (N6387, N6384, N2477, N1428);
nor NOR3 (N6388, N6381, N271, N6275);
nor NOR4 (N6389, N6365, N3852, N3008, N1958);
or OR3 (N6390, N6383, N539, N215);
xor XOR2 (N6391, N6371, N319);
nand NAND3 (N6392, N6378, N1396, N4546);
xor XOR2 (N6393, N6380, N5033);
and AND3 (N6394, N6388, N4486, N5744);
not NOT1 (N6395, N6392);
not NOT1 (N6396, N6393);
not NOT1 (N6397, N6387);
nor NOR3 (N6398, N6394, N977, N2924);
nand NAND4 (N6399, N6395, N1254, N120, N694);
not NOT1 (N6400, N6377);
not NOT1 (N6401, N6397);
not NOT1 (N6402, N6401);
not NOT1 (N6403, N6379);
nor NOR3 (N6404, N6398, N4408, N715);
buf BUF1 (N6405, N6400);
and AND2 (N6406, N6390, N2281);
nor NOR2 (N6407, N6389, N3615);
nor NOR3 (N6408, N6386, N1889, N675);
or OR4 (N6409, N6399, N3556, N3559, N4780);
and AND2 (N6410, N6407, N5129);
xor XOR2 (N6411, N6404, N291);
nor NOR2 (N6412, N6411, N5040);
or OR2 (N6413, N6391, N2466);
not NOT1 (N6414, N6396);
nand NAND4 (N6415, N6410, N4420, N2401, N4186);
and AND3 (N6416, N6405, N2658, N5934);
nand NAND3 (N6417, N6414, N2588, N4814);
xor XOR2 (N6418, N6412, N3440);
buf BUF1 (N6419, N6406);
or OR4 (N6420, N6402, N917, N4646, N4538);
buf BUF1 (N6421, N6415);
nand NAND4 (N6422, N6418, N6189, N4138, N5728);
not NOT1 (N6423, N6420);
nor NOR4 (N6424, N6403, N2657, N5622, N6376);
and AND2 (N6425, N6416, N4169);
nor NOR3 (N6426, N6413, N594, N2756);
buf BUF1 (N6427, N6417);
xor XOR2 (N6428, N6424, N1416);
nand NAND3 (N6429, N6425, N3446, N2293);
not NOT1 (N6430, N6408);
not NOT1 (N6431, N6430);
xor XOR2 (N6432, N6428, N4517);
nand NAND3 (N6433, N6419, N2211, N2145);
xor XOR2 (N6434, N6429, N208);
buf BUF1 (N6435, N6434);
not NOT1 (N6436, N6423);
nor NOR4 (N6437, N6432, N204, N619, N4872);
not NOT1 (N6438, N6421);
buf BUF1 (N6439, N6436);
not NOT1 (N6440, N6437);
not NOT1 (N6441, N6422);
and AND2 (N6442, N6440, N5224);
xor XOR2 (N6443, N6441, N6152);
xor XOR2 (N6444, N6431, N4563);
or OR3 (N6445, N6444, N4038, N819);
xor XOR2 (N6446, N6439, N76);
not NOT1 (N6447, N6446);
nor NOR2 (N6448, N6438, N876);
xor XOR2 (N6449, N6427, N2400);
buf BUF1 (N6450, N6442);
and AND2 (N6451, N6426, N1515);
buf BUF1 (N6452, N6449);
nor NOR2 (N6453, N6447, N568);
xor XOR2 (N6454, N6450, N3696);
xor XOR2 (N6455, N6435, N2528);
xor XOR2 (N6456, N6448, N389);
buf BUF1 (N6457, N6409);
nand NAND4 (N6458, N6456, N1784, N513, N2284);
not NOT1 (N6459, N6451);
nand NAND4 (N6460, N6452, N4892, N4892, N3037);
nor NOR3 (N6461, N6433, N3142, N1223);
buf BUF1 (N6462, N6443);
or OR4 (N6463, N6461, N2268, N2753, N4444);
xor XOR2 (N6464, N6460, N3395);
not NOT1 (N6465, N6458);
nor NOR4 (N6466, N6464, N6352, N921, N3069);
not NOT1 (N6467, N6455);
and AND4 (N6468, N6467, N3033, N4972, N5233);
xor XOR2 (N6469, N6457, N2472);
and AND3 (N6470, N6453, N2143, N2850);
or OR2 (N6471, N6462, N1681);
or OR2 (N6472, N6463, N5808);
and AND2 (N6473, N6468, N4108);
or OR2 (N6474, N6454, N2925);
and AND3 (N6475, N6445, N1657, N3595);
nand NAND2 (N6476, N6473, N4793);
nor NOR3 (N6477, N6465, N4170, N5752);
nor NOR2 (N6478, N6469, N5550);
buf BUF1 (N6479, N6471);
buf BUF1 (N6480, N6475);
nand NAND3 (N6481, N6476, N4543, N3433);
nor NOR3 (N6482, N6478, N6151, N4563);
nand NAND4 (N6483, N6466, N5913, N3211, N3331);
nand NAND2 (N6484, N6470, N5107);
nand NAND2 (N6485, N6480, N6375);
nand NAND2 (N6486, N6477, N6359);
not NOT1 (N6487, N6486);
nand NAND3 (N6488, N6485, N5672, N3675);
not NOT1 (N6489, N6482);
and AND4 (N6490, N6489, N246, N4268, N224);
xor XOR2 (N6491, N6479, N1714);
nor NOR3 (N6492, N6481, N4450, N2862);
buf BUF1 (N6493, N6492);
and AND2 (N6494, N6484, N4486);
not NOT1 (N6495, N6472);
xor XOR2 (N6496, N6494, N4231);
xor XOR2 (N6497, N6459, N4872);
buf BUF1 (N6498, N6474);
buf BUF1 (N6499, N6496);
nor NOR3 (N6500, N6490, N1970, N2280);
nor NOR4 (N6501, N6495, N5806, N3772, N2860);
and AND4 (N6502, N6498, N1360, N5548, N3153);
buf BUF1 (N6503, N6491);
buf BUF1 (N6504, N6501);
and AND3 (N6505, N6499, N2387, N4386);
and AND3 (N6506, N6504, N1153, N4006);
nand NAND4 (N6507, N6493, N2381, N5883, N5352);
and AND2 (N6508, N6500, N5427);
and AND2 (N6509, N6497, N4218);
not NOT1 (N6510, N6503);
buf BUF1 (N6511, N6487);
and AND2 (N6512, N6502, N3940);
and AND4 (N6513, N6505, N120, N5955, N1741);
or OR4 (N6514, N6512, N5472, N3053, N1405);
nor NOR4 (N6515, N6509, N5519, N4603, N6500);
or OR3 (N6516, N6507, N5321, N5413);
and AND3 (N6517, N6513, N6401, N3635);
not NOT1 (N6518, N6506);
xor XOR2 (N6519, N6517, N2784);
buf BUF1 (N6520, N6515);
nor NOR4 (N6521, N6518, N4294, N2607, N2587);
xor XOR2 (N6522, N6511, N208);
xor XOR2 (N6523, N6519, N2751);
and AND4 (N6524, N6508, N2219, N3571, N4478);
and AND2 (N6525, N6522, N144);
and AND3 (N6526, N6521, N3769, N5456);
buf BUF1 (N6527, N6483);
or OR4 (N6528, N6514, N5383, N2597, N5922);
not NOT1 (N6529, N6528);
and AND2 (N6530, N6527, N6312);
nand NAND4 (N6531, N6523, N3831, N3999, N1074);
and AND3 (N6532, N6516, N3381, N731);
or OR4 (N6533, N6526, N4620, N2885, N938);
nor NOR2 (N6534, N6525, N1110);
nand NAND2 (N6535, N6531, N1706);
and AND3 (N6536, N6524, N4809, N4536);
xor XOR2 (N6537, N6510, N3373);
and AND4 (N6538, N6536, N4822, N3119, N6024);
nor NOR3 (N6539, N6534, N4754, N2098);
buf BUF1 (N6540, N6529);
not NOT1 (N6541, N6532);
or OR3 (N6542, N6520, N6147, N1947);
nand NAND2 (N6543, N6541, N6502);
xor XOR2 (N6544, N6543, N5049);
nand NAND2 (N6545, N6533, N3039);
xor XOR2 (N6546, N6539, N4198);
and AND3 (N6547, N6530, N6346, N2478);
buf BUF1 (N6548, N6547);
nand NAND3 (N6549, N6544, N3135, N4424);
nand NAND3 (N6550, N6545, N3909, N4150);
nor NOR3 (N6551, N6537, N4385, N729);
xor XOR2 (N6552, N6542, N183);
nor NOR2 (N6553, N6550, N652);
xor XOR2 (N6554, N6553, N964);
not NOT1 (N6555, N6540);
nand NAND2 (N6556, N6546, N4596);
not NOT1 (N6557, N6538);
nor NOR2 (N6558, N6535, N5150);
buf BUF1 (N6559, N6558);
and AND2 (N6560, N6549, N2119);
nor NOR4 (N6561, N6551, N5246, N2703, N6323);
nor NOR2 (N6562, N6555, N5688);
nand NAND4 (N6563, N6557, N6484, N3853, N1195);
buf BUF1 (N6564, N6554);
nand NAND3 (N6565, N6560, N3995, N3926);
xor XOR2 (N6566, N6565, N2846);
nor NOR2 (N6567, N6488, N1139);
and AND4 (N6568, N6548, N3754, N6452, N1244);
nor NOR3 (N6569, N6566, N1826, N6350);
xor XOR2 (N6570, N6552, N4477);
nand NAND3 (N6571, N6569, N597, N6446);
and AND3 (N6572, N6567, N2553, N336);
or OR3 (N6573, N6571, N580, N6517);
nor NOR2 (N6574, N6561, N2785);
xor XOR2 (N6575, N6574, N1267);
nor NOR2 (N6576, N6556, N3765);
and AND4 (N6577, N6562, N6083, N1837, N3707);
xor XOR2 (N6578, N6559, N6177);
or OR2 (N6579, N6578, N6467);
xor XOR2 (N6580, N6563, N3213);
nand NAND3 (N6581, N6576, N2092, N6578);
nor NOR4 (N6582, N6570, N6404, N1144, N1081);
not NOT1 (N6583, N6577);
xor XOR2 (N6584, N6575, N3853);
nor NOR4 (N6585, N6572, N1439, N1276, N5373);
or OR3 (N6586, N6582, N1236, N2598);
and AND2 (N6587, N6584, N6523);
buf BUF1 (N6588, N6587);
xor XOR2 (N6589, N6579, N4656);
nor NOR2 (N6590, N6580, N2272);
nand NAND3 (N6591, N6590, N2714, N1102);
xor XOR2 (N6592, N6583, N3957);
or OR2 (N6593, N6581, N5943);
or OR4 (N6594, N6588, N3800, N1154, N4584);
xor XOR2 (N6595, N6586, N3770);
and AND4 (N6596, N6591, N6154, N86, N718);
nor NOR4 (N6597, N6592, N2175, N1248, N2339);
xor XOR2 (N6598, N6585, N5110);
not NOT1 (N6599, N6598);
nand NAND4 (N6600, N6589, N1938, N5401, N6087);
and AND4 (N6601, N6573, N4002, N2268, N6085);
nor NOR4 (N6602, N6599, N6174, N4446, N992);
not NOT1 (N6603, N6568);
buf BUF1 (N6604, N6603);
nor NOR2 (N6605, N6600, N3946);
xor XOR2 (N6606, N6596, N5399);
nand NAND4 (N6607, N6605, N3451, N1949, N2871);
nor NOR2 (N6608, N6597, N4396);
xor XOR2 (N6609, N6608, N4315);
not NOT1 (N6610, N6609);
or OR3 (N6611, N6593, N1617, N6272);
buf BUF1 (N6612, N6602);
or OR4 (N6613, N6595, N92, N4344, N3551);
nand NAND2 (N6614, N6606, N2185);
xor XOR2 (N6615, N6610, N2803);
nor NOR3 (N6616, N6594, N6081, N5869);
nor NOR2 (N6617, N6564, N1878);
and AND2 (N6618, N6613, N1119);
nand NAND2 (N6619, N6604, N2725);
xor XOR2 (N6620, N6614, N1417);
nor NOR2 (N6621, N6607, N3783);
or OR3 (N6622, N6616, N2750, N2035);
and AND2 (N6623, N6617, N5260);
or OR2 (N6624, N6611, N282);
or OR3 (N6625, N6615, N119, N656);
nand NAND3 (N6626, N6622, N365, N2369);
or OR2 (N6627, N6612, N3690);
nor NOR4 (N6628, N6624, N2380, N5280, N3587);
buf BUF1 (N6629, N6621);
and AND3 (N6630, N6628, N2995, N1665);
xor XOR2 (N6631, N6627, N2490);
or OR3 (N6632, N6623, N3419, N3482);
or OR4 (N6633, N6625, N4900, N3762, N3861);
buf BUF1 (N6634, N6626);
not NOT1 (N6635, N6619);
and AND2 (N6636, N6629, N817);
not NOT1 (N6637, N6636);
xor XOR2 (N6638, N6633, N6129);
xor XOR2 (N6639, N6635, N1226);
or OR2 (N6640, N6637, N5920);
nand NAND2 (N6641, N6601, N2268);
nand NAND3 (N6642, N6632, N4479, N5336);
nor NOR4 (N6643, N6630, N2273, N1182, N5027);
or OR2 (N6644, N6643, N2562);
nand NAND4 (N6645, N6631, N539, N2456, N494);
not NOT1 (N6646, N6618);
xor XOR2 (N6647, N6640, N6576);
or OR3 (N6648, N6645, N580, N3961);
nand NAND3 (N6649, N6647, N228, N5335);
and AND3 (N6650, N6620, N5131, N4884);
and AND4 (N6651, N6644, N5926, N4516, N4363);
or OR4 (N6652, N6649, N351, N2055, N1084);
not NOT1 (N6653, N6651);
or OR2 (N6654, N6642, N701);
and AND4 (N6655, N6650, N6330, N3534, N4563);
or OR4 (N6656, N6646, N6049, N64, N6624);
buf BUF1 (N6657, N6654);
nand NAND3 (N6658, N6657, N2697, N3343);
and AND2 (N6659, N6653, N2712);
xor XOR2 (N6660, N6652, N4169);
nand NAND3 (N6661, N6638, N1786, N1635);
not NOT1 (N6662, N6660);
and AND4 (N6663, N6641, N4193, N3549, N3182);
not NOT1 (N6664, N6634);
and AND2 (N6665, N6656, N429);
not NOT1 (N6666, N6655);
or OR4 (N6667, N6659, N5455, N3711, N709);
xor XOR2 (N6668, N6661, N4237);
xor XOR2 (N6669, N6664, N3114);
xor XOR2 (N6670, N6658, N3059);
nor NOR3 (N6671, N6639, N4800, N2478);
or OR3 (N6672, N6670, N1202, N1775);
nand NAND4 (N6673, N6648, N4638, N1112, N3792);
buf BUF1 (N6674, N6667);
and AND3 (N6675, N6674, N3686, N4312);
nand NAND4 (N6676, N6663, N1733, N799, N4017);
xor XOR2 (N6677, N6676, N5700);
nand NAND3 (N6678, N6672, N742, N573);
and AND2 (N6679, N6666, N594);
not NOT1 (N6680, N6673);
and AND4 (N6681, N6662, N6564, N6463, N2909);
nand NAND3 (N6682, N6680, N4006, N3066);
xor XOR2 (N6683, N6682, N1238);
buf BUF1 (N6684, N6669);
buf BUF1 (N6685, N6684);
nor NOR3 (N6686, N6683, N4653, N6065);
buf BUF1 (N6687, N6681);
nand NAND4 (N6688, N6686, N5120, N3330, N5944);
xor XOR2 (N6689, N6668, N1065);
nand NAND4 (N6690, N6687, N3852, N1404, N2157);
nand NAND4 (N6691, N6689, N5352, N2739, N5366);
or OR4 (N6692, N6671, N2588, N3578, N4257);
nand NAND4 (N6693, N6690, N235, N5937, N1045);
nor NOR4 (N6694, N6685, N4754, N1230, N5310);
buf BUF1 (N6695, N6691);
and AND3 (N6696, N6665, N6274, N4787);
nand NAND3 (N6697, N6696, N4210, N2125);
nor NOR4 (N6698, N6688, N2317, N5083, N1748);
not NOT1 (N6699, N6675);
buf BUF1 (N6700, N6679);
and AND4 (N6701, N6695, N4867, N1537, N400);
not NOT1 (N6702, N6693);
xor XOR2 (N6703, N6699, N1045);
buf BUF1 (N6704, N6678);
and AND2 (N6705, N6701, N3768);
not NOT1 (N6706, N6702);
not NOT1 (N6707, N6697);
or OR4 (N6708, N6706, N2281, N1668, N4475);
not NOT1 (N6709, N6677);
and AND2 (N6710, N6694, N4897);
xor XOR2 (N6711, N6707, N5805);
nand NAND4 (N6712, N6709, N3206, N2460, N4817);
xor XOR2 (N6713, N6712, N2530);
xor XOR2 (N6714, N6711, N2776);
not NOT1 (N6715, N6698);
xor XOR2 (N6716, N6705, N3122);
nand NAND3 (N6717, N6703, N2638, N5447);
not NOT1 (N6718, N6717);
xor XOR2 (N6719, N6692, N2601);
nor NOR4 (N6720, N6719, N4768, N5595, N1124);
or OR4 (N6721, N6718, N2178, N1811, N2261);
xor XOR2 (N6722, N6713, N4235);
nand NAND2 (N6723, N6720, N1650);
xor XOR2 (N6724, N6710, N3659);
and AND4 (N6725, N6708, N6203, N2052, N2363);
nor NOR2 (N6726, N6723, N2896);
nand NAND3 (N6727, N6700, N3701, N5414);
xor XOR2 (N6728, N6722, N349);
xor XOR2 (N6729, N6728, N3125);
buf BUF1 (N6730, N6714);
and AND3 (N6731, N6704, N1903, N3090);
or OR4 (N6732, N6715, N3403, N1851, N5175);
not NOT1 (N6733, N6729);
buf BUF1 (N6734, N6733);
or OR4 (N6735, N6732, N3516, N6606, N3626);
and AND2 (N6736, N6726, N4398);
xor XOR2 (N6737, N6735, N2244);
or OR3 (N6738, N6730, N4329, N923);
xor XOR2 (N6739, N6734, N5057);
or OR4 (N6740, N6739, N4938, N5879, N594);
buf BUF1 (N6741, N6731);
xor XOR2 (N6742, N6736, N1258);
or OR3 (N6743, N6742, N6488, N2040);
xor XOR2 (N6744, N6737, N2510);
not NOT1 (N6745, N6721);
xor XOR2 (N6746, N6744, N3848);
not NOT1 (N6747, N6746);
or OR2 (N6748, N6745, N610);
and AND4 (N6749, N6741, N6075, N229, N2533);
nor NOR3 (N6750, N6743, N2996, N2182);
nand NAND3 (N6751, N6725, N1140, N6207);
and AND4 (N6752, N6738, N1941, N197, N2388);
not NOT1 (N6753, N6752);
nor NOR4 (N6754, N6753, N2191, N5802, N2274);
and AND4 (N6755, N6727, N2116, N2155, N2650);
buf BUF1 (N6756, N6749);
nor NOR3 (N6757, N6747, N9, N1793);
xor XOR2 (N6758, N6751, N5411);
buf BUF1 (N6759, N6757);
nand NAND2 (N6760, N6758, N4940);
nand NAND2 (N6761, N6756, N653);
nand NAND2 (N6762, N6759, N403);
xor XOR2 (N6763, N6750, N5174);
buf BUF1 (N6764, N6716);
xor XOR2 (N6765, N6762, N4822);
buf BUF1 (N6766, N6760);
nand NAND3 (N6767, N6724, N4888, N667);
xor XOR2 (N6768, N6765, N5042);
nor NOR2 (N6769, N6748, N5126);
nand NAND2 (N6770, N6764, N5241);
nand NAND2 (N6771, N6769, N5371);
and AND4 (N6772, N6755, N2836, N6350, N4128);
not NOT1 (N6773, N6768);
or OR4 (N6774, N6773, N1855, N6702, N670);
not NOT1 (N6775, N6740);
nand NAND2 (N6776, N6771, N2861);
xor XOR2 (N6777, N6754, N2777);
and AND2 (N6778, N6775, N1988);
xor XOR2 (N6779, N6761, N663);
xor XOR2 (N6780, N6766, N975);
nor NOR2 (N6781, N6774, N2801);
nor NOR4 (N6782, N6781, N2878, N4162, N6402);
and AND3 (N6783, N6763, N1843, N3125);
xor XOR2 (N6784, N6779, N5129);
buf BUF1 (N6785, N6772);
nor NOR2 (N6786, N6785, N322);
nand NAND2 (N6787, N6786, N2924);
or OR4 (N6788, N6783, N2954, N2801, N6398);
nor NOR3 (N6789, N6782, N2494, N5232);
and AND3 (N6790, N6778, N447, N3921);
not NOT1 (N6791, N6767);
not NOT1 (N6792, N6776);
nand NAND2 (N6793, N6791, N3620);
and AND2 (N6794, N6793, N5736);
or OR4 (N6795, N6784, N2190, N3555, N6487);
and AND2 (N6796, N6789, N2420);
buf BUF1 (N6797, N6794);
and AND3 (N6798, N6792, N4211, N3582);
nand NAND4 (N6799, N6770, N2361, N905, N2453);
nor NOR4 (N6800, N6795, N4477, N157, N1861);
or OR2 (N6801, N6777, N2811);
xor XOR2 (N6802, N6797, N1062);
not NOT1 (N6803, N6799);
or OR4 (N6804, N6796, N2350, N1727, N2431);
nand NAND2 (N6805, N6802, N4691);
not NOT1 (N6806, N6788);
or OR3 (N6807, N6801, N3809, N883);
nand NAND2 (N6808, N6804, N1066);
and AND4 (N6809, N6803, N6754, N2305, N4509);
xor XOR2 (N6810, N6790, N2267);
nor NOR2 (N6811, N6807, N498);
xor XOR2 (N6812, N6800, N4660);
not NOT1 (N6813, N6808);
not NOT1 (N6814, N6813);
buf BUF1 (N6815, N6810);
and AND4 (N6816, N6805, N345, N881, N2300);
buf BUF1 (N6817, N6806);
or OR2 (N6818, N6812, N1854);
and AND2 (N6819, N6780, N4347);
nor NOR3 (N6820, N6809, N2981, N3368);
or OR4 (N6821, N6798, N1061, N6252, N4676);
not NOT1 (N6822, N6819);
nor NOR2 (N6823, N6787, N5197);
and AND3 (N6824, N6811, N2797, N366);
xor XOR2 (N6825, N6821, N2915);
nor NOR3 (N6826, N6815, N1129, N1775);
and AND4 (N6827, N6814, N1627, N970, N3452);
or OR4 (N6828, N6824, N5451, N3545, N807);
nor NOR2 (N6829, N6818, N3387);
nand NAND3 (N6830, N6826, N3437, N2950);
and AND2 (N6831, N6817, N5468);
and AND4 (N6832, N6825, N3752, N48, N677);
nand NAND2 (N6833, N6820, N1031);
not NOT1 (N6834, N6829);
nand NAND3 (N6835, N6828, N3844, N3158);
xor XOR2 (N6836, N6831, N2281);
nor NOR4 (N6837, N6823, N3027, N1355, N5221);
nor NOR2 (N6838, N6830, N6393);
nand NAND2 (N6839, N6834, N4826);
xor XOR2 (N6840, N6822, N1649);
xor XOR2 (N6841, N6827, N86);
nor NOR2 (N6842, N6833, N5007);
xor XOR2 (N6843, N6842, N447);
nand NAND2 (N6844, N6843, N3871);
nor NOR4 (N6845, N6837, N4663, N6298, N399);
nor NOR2 (N6846, N6841, N4825);
and AND4 (N6847, N6832, N4749, N5316, N966);
nand NAND3 (N6848, N6847, N6125, N4429);
xor XOR2 (N6849, N6845, N80);
xor XOR2 (N6850, N6839, N3036);
not NOT1 (N6851, N6850);
xor XOR2 (N6852, N6849, N303);
xor XOR2 (N6853, N6851, N2874);
xor XOR2 (N6854, N6835, N5687);
and AND2 (N6855, N6848, N4402);
nand NAND2 (N6856, N6844, N5643);
and AND4 (N6857, N6840, N4784, N3357, N676);
and AND2 (N6858, N6854, N3676);
xor XOR2 (N6859, N6846, N708);
not NOT1 (N6860, N6855);
or OR2 (N6861, N6857, N1361);
or OR2 (N6862, N6838, N5870);
buf BUF1 (N6863, N6860);
buf BUF1 (N6864, N6856);
or OR4 (N6865, N6836, N5265, N1545, N6145);
or OR4 (N6866, N6852, N476, N1537, N3373);
nand NAND3 (N6867, N6864, N6685, N6576);
xor XOR2 (N6868, N6858, N4573);
nand NAND2 (N6869, N6816, N4207);
xor XOR2 (N6870, N6861, N2901);
or OR4 (N6871, N6868, N988, N4720, N638);
or OR4 (N6872, N6869, N5936, N5360, N4014);
or OR2 (N6873, N6865, N4345);
or OR3 (N6874, N6871, N5236, N4881);
nor NOR3 (N6875, N6870, N6236, N5446);
nor NOR4 (N6876, N6872, N5099, N3407, N3716);
and AND3 (N6877, N6866, N1929, N1854);
buf BUF1 (N6878, N6876);
nand NAND2 (N6879, N6878, N4320);
buf BUF1 (N6880, N6879);
and AND4 (N6881, N6853, N1313, N331, N6716);
xor XOR2 (N6882, N6862, N5769);
nor NOR3 (N6883, N6859, N5014, N2228);
nand NAND4 (N6884, N6877, N1626, N427, N6661);
or OR4 (N6885, N6873, N2958, N3831, N6136);
buf BUF1 (N6886, N6883);
not NOT1 (N6887, N6863);
xor XOR2 (N6888, N6886, N1768);
buf BUF1 (N6889, N6882);
nand NAND3 (N6890, N6885, N1669, N601);
nand NAND4 (N6891, N6888, N1455, N1418, N2629);
nor NOR4 (N6892, N6890, N3860, N4794, N4464);
buf BUF1 (N6893, N6867);
not NOT1 (N6894, N6880);
nand NAND2 (N6895, N6891, N5058);
not NOT1 (N6896, N6893);
nor NOR2 (N6897, N6889, N2882);
and AND2 (N6898, N6894, N3680);
buf BUF1 (N6899, N6898);
not NOT1 (N6900, N6884);
buf BUF1 (N6901, N6900);
nand NAND3 (N6902, N6874, N4801, N5111);
nand NAND3 (N6903, N6887, N6221, N673);
xor XOR2 (N6904, N6903, N2361);
and AND3 (N6905, N6895, N5326, N3748);
buf BUF1 (N6906, N6897);
nand NAND2 (N6907, N6902, N5587);
or OR3 (N6908, N6901, N5217, N564);
and AND3 (N6909, N6875, N6493, N3270);
and AND2 (N6910, N6907, N394);
not NOT1 (N6911, N6906);
and AND3 (N6912, N6881, N3826, N4123);
or OR3 (N6913, N6910, N2295, N6255);
nor NOR3 (N6914, N6913, N411, N3457);
or OR2 (N6915, N6911, N3071);
nor NOR4 (N6916, N6899, N809, N744, N3474);
and AND2 (N6917, N6892, N1028);
not NOT1 (N6918, N6896);
xor XOR2 (N6919, N6908, N6574);
buf BUF1 (N6920, N6904);
xor XOR2 (N6921, N6915, N6433);
xor XOR2 (N6922, N6905, N4451);
not NOT1 (N6923, N6916);
buf BUF1 (N6924, N6917);
nand NAND3 (N6925, N6920, N5734, N258);
and AND4 (N6926, N6909, N3558, N6114, N6578);
xor XOR2 (N6927, N6925, N1380);
nand NAND2 (N6928, N6921, N3315);
nand NAND3 (N6929, N6918, N6695, N1454);
xor XOR2 (N6930, N6927, N5504);
xor XOR2 (N6931, N6926, N4428);
nor NOR3 (N6932, N6922, N3240, N6045);
not NOT1 (N6933, N6928);
not NOT1 (N6934, N6924);
or OR2 (N6935, N6912, N2896);
not NOT1 (N6936, N6929);
or OR2 (N6937, N6930, N4285);
xor XOR2 (N6938, N6933, N2095);
or OR2 (N6939, N6935, N2064);
nand NAND3 (N6940, N6932, N1815, N6882);
not NOT1 (N6941, N6939);
buf BUF1 (N6942, N6940);
buf BUF1 (N6943, N6942);
not NOT1 (N6944, N6943);
nand NAND4 (N6945, N6923, N3648, N2648, N165);
buf BUF1 (N6946, N6938);
buf BUF1 (N6947, N6946);
nor NOR4 (N6948, N6936, N4788, N2638, N5239);
or OR4 (N6949, N6937, N5094, N2281, N1427);
xor XOR2 (N6950, N6941, N2175);
or OR4 (N6951, N6944, N6928, N1078, N6473);
xor XOR2 (N6952, N6934, N3932);
and AND4 (N6953, N6914, N5419, N6772, N5037);
not NOT1 (N6954, N6952);
nor NOR2 (N6955, N6949, N3226);
not NOT1 (N6956, N6953);
and AND2 (N6957, N6919, N5427);
and AND2 (N6958, N6947, N1745);
or OR4 (N6959, N6948, N67, N3896, N706);
and AND2 (N6960, N6950, N4994);
nor NOR3 (N6961, N6960, N4993, N1112);
not NOT1 (N6962, N6955);
nor NOR4 (N6963, N6958, N6786, N6372, N3202);
buf BUF1 (N6964, N6957);
or OR2 (N6965, N6959, N5135);
xor XOR2 (N6966, N6962, N2229);
buf BUF1 (N6967, N6954);
nand NAND3 (N6968, N6966, N4690, N6462);
or OR4 (N6969, N6961, N4422, N5212, N1726);
not NOT1 (N6970, N6969);
not NOT1 (N6971, N6963);
nor NOR4 (N6972, N6965, N6176, N3596, N1867);
buf BUF1 (N6973, N6968);
and AND3 (N6974, N6945, N2327, N3859);
not NOT1 (N6975, N6956);
nand NAND4 (N6976, N6964, N4576, N2412, N1606);
nand NAND4 (N6977, N6971, N3155, N4323, N4991);
or OR3 (N6978, N6951, N1387, N3271);
nand NAND4 (N6979, N6967, N5537, N4949, N2268);
and AND3 (N6980, N6970, N446, N3752);
nand NAND3 (N6981, N6973, N6668, N904);
or OR2 (N6982, N6931, N4177);
nand NAND3 (N6983, N6981, N1790, N2079);
nor NOR4 (N6984, N6977, N1234, N4426, N79);
xor XOR2 (N6985, N6972, N3442);
buf BUF1 (N6986, N6974);
and AND2 (N6987, N6975, N4397);
nand NAND2 (N6988, N6983, N5486);
xor XOR2 (N6989, N6978, N6400);
xor XOR2 (N6990, N6986, N1364);
and AND3 (N6991, N6988, N3470, N6);
nor NOR2 (N6992, N6982, N1589);
nand NAND4 (N6993, N6984, N1172, N4417, N5600);
nand NAND4 (N6994, N6980, N3658, N4138, N4101);
nand NAND3 (N6995, N6991, N5739, N5441);
and AND2 (N6996, N6989, N3008);
and AND4 (N6997, N6979, N2458, N1404, N6328);
or OR3 (N6998, N6997, N3969, N315);
buf BUF1 (N6999, N6976);
nor NOR4 (N7000, N6992, N883, N6593, N116);
nor NOR4 (N7001, N7000, N1074, N4895, N6840);
buf BUF1 (N7002, N6987);
and AND2 (N7003, N6993, N4065);
nor NOR4 (N7004, N7001, N383, N6427, N2533);
and AND2 (N7005, N6998, N1812);
nor NOR3 (N7006, N6985, N6281, N2133);
nor NOR3 (N7007, N7003, N4863, N6385);
or OR3 (N7008, N6990, N5080, N2479);
not NOT1 (N7009, N7007);
not NOT1 (N7010, N7002);
buf BUF1 (N7011, N7008);
or OR2 (N7012, N7010, N1022);
or OR2 (N7013, N7011, N5786);
or OR4 (N7014, N7012, N3096, N2558, N3834);
nor NOR2 (N7015, N6999, N2405);
xor XOR2 (N7016, N7009, N3766);
xor XOR2 (N7017, N7016, N6695);
not NOT1 (N7018, N7005);
xor XOR2 (N7019, N7004, N601);
or OR4 (N7020, N6994, N1729, N6069, N1795);
or OR2 (N7021, N7019, N1739);
xor XOR2 (N7022, N6996, N1397);
or OR4 (N7023, N7021, N311, N6542, N1503);
buf BUF1 (N7024, N7006);
not NOT1 (N7025, N7023);
buf BUF1 (N7026, N7018);
xor XOR2 (N7027, N7026, N5834);
and AND2 (N7028, N7014, N5236);
nor NOR4 (N7029, N7027, N3962, N1365, N1339);
or OR4 (N7030, N7022, N6338, N2609, N3507);
not NOT1 (N7031, N6995);
xor XOR2 (N7032, N7025, N2406);
buf BUF1 (N7033, N7031);
xor XOR2 (N7034, N7017, N1940);
or OR2 (N7035, N7024, N6269);
and AND2 (N7036, N7029, N4561);
or OR3 (N7037, N7033, N2416, N666);
nor NOR3 (N7038, N7015, N1496, N6239);
buf BUF1 (N7039, N7036);
not NOT1 (N7040, N7032);
buf BUF1 (N7041, N7038);
nor NOR2 (N7042, N7040, N6496);
buf BUF1 (N7043, N7035);
xor XOR2 (N7044, N7043, N6048);
xor XOR2 (N7045, N7028, N6543);
not NOT1 (N7046, N7034);
xor XOR2 (N7047, N7039, N5411);
and AND4 (N7048, N7030, N5888, N1717, N5166);
buf BUF1 (N7049, N7048);
not NOT1 (N7050, N7045);
not NOT1 (N7051, N7050);
not NOT1 (N7052, N7046);
xor XOR2 (N7053, N7047, N5288);
buf BUF1 (N7054, N7042);
or OR4 (N7055, N7037, N1941, N2648, N5750);
and AND2 (N7056, N7055, N5280);
and AND3 (N7057, N7052, N2722, N2717);
and AND2 (N7058, N7044, N693);
xor XOR2 (N7059, N7049, N1559);
buf BUF1 (N7060, N7041);
nand NAND3 (N7061, N7057, N3403, N3369);
nor NOR3 (N7062, N7061, N6522, N5917);
nand NAND2 (N7063, N7060, N5355);
buf BUF1 (N7064, N7053);
nand NAND2 (N7065, N7054, N4923);
not NOT1 (N7066, N7020);
nand NAND2 (N7067, N7056, N893);
or OR3 (N7068, N7067, N445, N1942);
not NOT1 (N7069, N7013);
and AND4 (N7070, N7058, N385, N5794, N231);
xor XOR2 (N7071, N7070, N2971);
and AND3 (N7072, N7065, N2076, N6214);
buf BUF1 (N7073, N7064);
buf BUF1 (N7074, N7073);
and AND4 (N7075, N7069, N6518, N6712, N1513);
not NOT1 (N7076, N7075);
nor NOR2 (N7077, N7068, N2598);
xor XOR2 (N7078, N7071, N6051);
nand NAND4 (N7079, N7059, N3342, N6852, N20);
xor XOR2 (N7080, N7072, N45);
buf BUF1 (N7081, N7080);
or OR2 (N7082, N7051, N2254);
nand NAND2 (N7083, N7078, N503);
xor XOR2 (N7084, N7062, N3527);
not NOT1 (N7085, N7063);
nand NAND2 (N7086, N7084, N2987);
xor XOR2 (N7087, N7079, N4212);
nand NAND4 (N7088, N7074, N2905, N2492, N4118);
xor XOR2 (N7089, N7081, N3068);
and AND4 (N7090, N7089, N4546, N5418, N1149);
xor XOR2 (N7091, N7086, N6362);
xor XOR2 (N7092, N7087, N3586);
or OR4 (N7093, N7076, N5761, N4654, N5367);
not NOT1 (N7094, N7082);
and AND4 (N7095, N7090, N1640, N4581, N1651);
and AND3 (N7096, N7066, N3088, N921);
xor XOR2 (N7097, N7095, N718);
xor XOR2 (N7098, N7096, N5083);
not NOT1 (N7099, N7077);
nand NAND2 (N7100, N7091, N5151);
or OR3 (N7101, N7083, N4434, N3362);
or OR2 (N7102, N7100, N4947);
xor XOR2 (N7103, N7092, N6912);
buf BUF1 (N7104, N7085);
and AND2 (N7105, N7101, N1327);
xor XOR2 (N7106, N7105, N4665);
nand NAND3 (N7107, N7099, N2942, N4767);
xor XOR2 (N7108, N7098, N1913);
or OR4 (N7109, N7106, N4746, N2914, N2264);
buf BUF1 (N7110, N7093);
not NOT1 (N7111, N7102);
and AND3 (N7112, N7104, N1150, N4310);
and AND2 (N7113, N7107, N6921);
not NOT1 (N7114, N7111);
or OR4 (N7115, N7088, N2352, N3827, N1328);
or OR3 (N7116, N7103, N3143, N955);
xor XOR2 (N7117, N7116, N5677);
nand NAND4 (N7118, N7094, N5113, N3739, N2450);
xor XOR2 (N7119, N7114, N5290);
and AND4 (N7120, N7118, N4513, N838, N5524);
xor XOR2 (N7121, N7119, N1753);
nor NOR3 (N7122, N7109, N2742, N5308);
buf BUF1 (N7123, N7112);
or OR2 (N7124, N7108, N3056);
or OR3 (N7125, N7124, N785, N2458);
nor NOR2 (N7126, N7117, N4043);
not NOT1 (N7127, N7097);
nor NOR4 (N7128, N7126, N3226, N5780, N4697);
and AND3 (N7129, N7115, N182, N6541);
buf BUF1 (N7130, N7110);
xor XOR2 (N7131, N7121, N6076);
buf BUF1 (N7132, N7113);
buf BUF1 (N7133, N7127);
xor XOR2 (N7134, N7120, N3427);
buf BUF1 (N7135, N7123);
and AND2 (N7136, N7135, N2521);
nand NAND4 (N7137, N7128, N5124, N2986, N3607);
and AND2 (N7138, N7122, N1105);
nand NAND4 (N7139, N7129, N6839, N3633, N1199);
not NOT1 (N7140, N7136);
not NOT1 (N7141, N7132);
not NOT1 (N7142, N7125);
nand NAND4 (N7143, N7133, N6203, N3036, N6425);
or OR4 (N7144, N7138, N2466, N42, N1544);
or OR3 (N7145, N7131, N1831, N2141);
nor NOR2 (N7146, N7134, N3666);
or OR4 (N7147, N7143, N4055, N974, N4676);
and AND4 (N7148, N7145, N5130, N4672, N748);
nand NAND4 (N7149, N7137, N1858, N3218, N101);
not NOT1 (N7150, N7130);
or OR4 (N7151, N7150, N1802, N3905, N2830);
and AND3 (N7152, N7148, N5594, N2559);
nand NAND4 (N7153, N7139, N3281, N5230, N3286);
buf BUF1 (N7154, N7149);
or OR2 (N7155, N7141, N4792);
and AND3 (N7156, N7140, N1571, N1991);
xor XOR2 (N7157, N7144, N5204);
xor XOR2 (N7158, N7147, N6249);
buf BUF1 (N7159, N7142);
or OR3 (N7160, N7152, N5847, N415);
nand NAND2 (N7161, N7155, N1911);
buf BUF1 (N7162, N7158);
nor NOR4 (N7163, N7151, N2263, N5210, N5753);
or OR4 (N7164, N7156, N1284, N3620, N1161);
nor NOR2 (N7165, N7161, N4635);
nor NOR4 (N7166, N7164, N430, N5605, N882);
buf BUF1 (N7167, N7165);
nor NOR2 (N7168, N7163, N6812);
buf BUF1 (N7169, N7146);
or OR2 (N7170, N7167, N5895);
not NOT1 (N7171, N7159);
nor NOR4 (N7172, N7160, N6841, N2650, N2421);
buf BUF1 (N7173, N7157);
and AND4 (N7174, N7153, N7053, N1855, N4793);
and AND2 (N7175, N7154, N5179);
buf BUF1 (N7176, N7172);
nand NAND3 (N7177, N7175, N4877, N6949);
xor XOR2 (N7178, N7166, N217);
not NOT1 (N7179, N7176);
and AND3 (N7180, N7169, N2039, N1688);
or OR2 (N7181, N7174, N6305);
not NOT1 (N7182, N7173);
or OR2 (N7183, N7179, N5021);
not NOT1 (N7184, N7181);
nor NOR3 (N7185, N7178, N3497, N4864);
not NOT1 (N7186, N7170);
and AND4 (N7187, N7162, N3213, N4544, N7103);
nand NAND4 (N7188, N7184, N3939, N3675, N2129);
not NOT1 (N7189, N7187);
xor XOR2 (N7190, N7185, N979);
xor XOR2 (N7191, N7180, N2822);
not NOT1 (N7192, N7171);
or OR4 (N7193, N7182, N1477, N4947, N1213);
buf BUF1 (N7194, N7168);
and AND4 (N7195, N7192, N2171, N3799, N6549);
nand NAND2 (N7196, N7191, N2295);
xor XOR2 (N7197, N7190, N643);
and AND3 (N7198, N7186, N2547, N6222);
buf BUF1 (N7199, N7196);
not NOT1 (N7200, N7177);
or OR4 (N7201, N7189, N4378, N5949, N4065);
and AND3 (N7202, N7200, N2066, N4446);
nand NAND4 (N7203, N7202, N797, N662, N523);
xor XOR2 (N7204, N7197, N1484);
not NOT1 (N7205, N7198);
or OR4 (N7206, N7193, N28, N6594, N6044);
buf BUF1 (N7207, N7205);
not NOT1 (N7208, N7188);
not NOT1 (N7209, N7195);
nor NOR4 (N7210, N7209, N2162, N1822, N1001);
xor XOR2 (N7211, N7201, N11);
not NOT1 (N7212, N7206);
or OR3 (N7213, N7183, N6717, N2091);
buf BUF1 (N7214, N7211);
buf BUF1 (N7215, N7199);
buf BUF1 (N7216, N7194);
nor NOR4 (N7217, N7207, N2188, N3992, N2056);
and AND4 (N7218, N7212, N4250, N1879, N5744);
or OR2 (N7219, N7208, N6599);
and AND4 (N7220, N7218, N264, N1339, N937);
nor NOR2 (N7221, N7204, N1078);
nor NOR2 (N7222, N7214, N4772);
buf BUF1 (N7223, N7210);
nand NAND2 (N7224, N7215, N6221);
or OR4 (N7225, N7217, N3307, N2853, N5136);
nand NAND2 (N7226, N7221, N2375);
buf BUF1 (N7227, N7219);
xor XOR2 (N7228, N7216, N5937);
not NOT1 (N7229, N7228);
and AND2 (N7230, N7213, N6478);
or OR3 (N7231, N7229, N186, N5744);
xor XOR2 (N7232, N7227, N1829);
xor XOR2 (N7233, N7220, N2753);
nor NOR3 (N7234, N7231, N1778, N928);
buf BUF1 (N7235, N7230);
nor NOR3 (N7236, N7226, N2376, N5493);
nand NAND4 (N7237, N7236, N6499, N538, N2725);
xor XOR2 (N7238, N7233, N4277);
nor NOR2 (N7239, N7234, N3525);
buf BUF1 (N7240, N7237);
or OR4 (N7241, N7224, N5098, N5701, N6720);
xor XOR2 (N7242, N7222, N2012);
nand NAND3 (N7243, N7242, N7111, N5757);
xor XOR2 (N7244, N7225, N5213);
xor XOR2 (N7245, N7240, N2577);
xor XOR2 (N7246, N7241, N1837);
and AND4 (N7247, N7239, N4633, N992, N3401);
or OR4 (N7248, N7223, N4026, N5029, N6335);
and AND4 (N7249, N7244, N6977, N7158, N6665);
not NOT1 (N7250, N7243);
xor XOR2 (N7251, N7238, N1930);
xor XOR2 (N7252, N7232, N6110);
nand NAND3 (N7253, N7250, N3188, N6797);
buf BUF1 (N7254, N7235);
buf BUF1 (N7255, N7245);
buf BUF1 (N7256, N7248);
xor XOR2 (N7257, N7247, N5474);
nor NOR2 (N7258, N7256, N1983);
and AND2 (N7259, N7252, N872);
and AND4 (N7260, N7257, N6131, N5429, N5047);
buf BUF1 (N7261, N7260);
not NOT1 (N7262, N7255);
not NOT1 (N7263, N7249);
or OR3 (N7264, N7263, N550, N1951);
buf BUF1 (N7265, N7261);
and AND2 (N7266, N7259, N1423);
nand NAND2 (N7267, N7264, N1710);
xor XOR2 (N7268, N7251, N4924);
nor NOR3 (N7269, N7262, N461, N1089);
or OR4 (N7270, N7203, N4078, N6202, N3305);
and AND3 (N7271, N7266, N5360, N2434);
and AND2 (N7272, N7268, N3035);
not NOT1 (N7273, N7272);
or OR2 (N7274, N7267, N4390);
and AND3 (N7275, N7270, N3542, N776);
not NOT1 (N7276, N7254);
nor NOR4 (N7277, N7258, N6320, N6967, N5598);
or OR2 (N7278, N7271, N6338);
xor XOR2 (N7279, N7269, N203);
nand NAND4 (N7280, N7279, N4833, N3327, N3125);
not NOT1 (N7281, N7280);
or OR3 (N7282, N7275, N4016, N2241);
and AND2 (N7283, N7265, N2402);
buf BUF1 (N7284, N7253);
xor XOR2 (N7285, N7283, N5366);
buf BUF1 (N7286, N7281);
xor XOR2 (N7287, N7284, N1838);
and AND3 (N7288, N7276, N3364, N2165);
or OR3 (N7289, N7287, N3810, N2665);
and AND4 (N7290, N7286, N4807, N5189, N4580);
buf BUF1 (N7291, N7274);
nor NOR3 (N7292, N7278, N3480, N3140);
xor XOR2 (N7293, N7246, N1570);
buf BUF1 (N7294, N7282);
or OR2 (N7295, N7291, N165);
xor XOR2 (N7296, N7294, N1394);
and AND3 (N7297, N7289, N6982, N1641);
and AND3 (N7298, N7273, N4575, N374);
buf BUF1 (N7299, N7295);
not NOT1 (N7300, N7298);
buf BUF1 (N7301, N7290);
nand NAND4 (N7302, N7293, N2411, N3236, N3234);
or OR3 (N7303, N7277, N5756, N5081);
nand NAND3 (N7304, N7292, N1948, N4599);
nand NAND4 (N7305, N7304, N6062, N4361, N1758);
or OR2 (N7306, N7303, N5373);
or OR3 (N7307, N7300, N578, N2147);
nand NAND2 (N7308, N7288, N2556);
not NOT1 (N7309, N7299);
not NOT1 (N7310, N7307);
nand NAND3 (N7311, N7302, N2218, N1718);
or OR3 (N7312, N7306, N7044, N1755);
and AND3 (N7313, N7297, N3281, N2426);
not NOT1 (N7314, N7309);
and AND2 (N7315, N7285, N1799);
and AND2 (N7316, N7315, N1914);
or OR3 (N7317, N7312, N3382, N1515);
nand NAND3 (N7318, N7314, N3532, N6588);
not NOT1 (N7319, N7301);
nor NOR3 (N7320, N7313, N2942, N1633);
and AND3 (N7321, N7311, N3998, N5483);
xor XOR2 (N7322, N7296, N3475);
not NOT1 (N7323, N7320);
nand NAND4 (N7324, N7308, N4161, N7000, N1097);
buf BUF1 (N7325, N7305);
nor NOR3 (N7326, N7318, N314, N486);
xor XOR2 (N7327, N7326, N2805);
or OR2 (N7328, N7321, N3458);
nor NOR2 (N7329, N7324, N6722);
or OR2 (N7330, N7310, N3035);
nand NAND4 (N7331, N7319, N1379, N3540, N3138);
nand NAND4 (N7332, N7316, N1437, N3537, N1875);
and AND3 (N7333, N7331, N2779, N4327);
xor XOR2 (N7334, N7317, N4134);
not NOT1 (N7335, N7330);
nor NOR3 (N7336, N7335, N2491, N6542);
and AND3 (N7337, N7332, N2870, N5785);
buf BUF1 (N7338, N7333);
and AND4 (N7339, N7329, N5602, N5902, N6337);
buf BUF1 (N7340, N7328);
buf BUF1 (N7341, N7327);
nor NOR4 (N7342, N7322, N4933, N2339, N1731);
not NOT1 (N7343, N7336);
buf BUF1 (N7344, N7343);
xor XOR2 (N7345, N7337, N237);
nor NOR4 (N7346, N7345, N5620, N3556, N3208);
not NOT1 (N7347, N7339);
nand NAND3 (N7348, N7344, N3237, N4615);
xor XOR2 (N7349, N7348, N6946);
not NOT1 (N7350, N7346);
or OR3 (N7351, N7338, N1561, N5205);
nand NAND4 (N7352, N7347, N5945, N1277, N3365);
not NOT1 (N7353, N7325);
and AND2 (N7354, N7341, N3804);
nor NOR2 (N7355, N7334, N4834);
not NOT1 (N7356, N7323);
nor NOR2 (N7357, N7356, N1234);
not NOT1 (N7358, N7351);
and AND3 (N7359, N7342, N4697, N5744);
nand NAND3 (N7360, N7357, N6342, N3296);
and AND2 (N7361, N7350, N1660);
and AND3 (N7362, N7358, N5935, N7315);
nand NAND3 (N7363, N7355, N5792, N6905);
xor XOR2 (N7364, N7349, N2744);
not NOT1 (N7365, N7359);
nand NAND2 (N7366, N7352, N910);
and AND2 (N7367, N7363, N3410);
or OR2 (N7368, N7361, N752);
buf BUF1 (N7369, N7362);
and AND4 (N7370, N7340, N3102, N4175, N1498);
and AND4 (N7371, N7364, N145, N6912, N5016);
xor XOR2 (N7372, N7370, N1075);
or OR2 (N7373, N7360, N5474);
nor NOR4 (N7374, N7354, N6640, N2356, N829);
nor NOR4 (N7375, N7372, N821, N5796, N3450);
not NOT1 (N7376, N7366);
nor NOR2 (N7377, N7373, N3922);
nor NOR2 (N7378, N7377, N3796);
nor NOR3 (N7379, N7365, N3533, N1665);
or OR4 (N7380, N7376, N551, N1625, N2885);
not NOT1 (N7381, N7353);
and AND2 (N7382, N7374, N3731);
xor XOR2 (N7383, N7375, N2889);
not NOT1 (N7384, N7383);
or OR3 (N7385, N7371, N3881, N1004);
xor XOR2 (N7386, N7382, N3367);
nand NAND4 (N7387, N7378, N579, N1809, N3057);
nor NOR4 (N7388, N7385, N6417, N415, N4931);
and AND3 (N7389, N7386, N5254, N2218);
or OR4 (N7390, N7368, N2908, N3144, N2958);
not NOT1 (N7391, N7381);
and AND3 (N7392, N7387, N5136, N5813);
buf BUF1 (N7393, N7379);
xor XOR2 (N7394, N7392, N2067);
not NOT1 (N7395, N7380);
nand NAND2 (N7396, N7391, N3476);
xor XOR2 (N7397, N7394, N394);
or OR3 (N7398, N7397, N4623, N5049);
nor NOR2 (N7399, N7369, N3764);
not NOT1 (N7400, N7389);
xor XOR2 (N7401, N7390, N6698);
buf BUF1 (N7402, N7384);
nor NOR4 (N7403, N7400, N5727, N4797, N6062);
and AND4 (N7404, N7395, N665, N4466, N3100);
xor XOR2 (N7405, N7393, N3504);
and AND3 (N7406, N7388, N4821, N1117);
not NOT1 (N7407, N7404);
not NOT1 (N7408, N7399);
or OR4 (N7409, N7403, N1035, N3799, N4567);
xor XOR2 (N7410, N7402, N913);
not NOT1 (N7411, N7367);
nor NOR4 (N7412, N7401, N737, N1230, N2161);
xor XOR2 (N7413, N7396, N595);
xor XOR2 (N7414, N7411, N2130);
nor NOR3 (N7415, N7414, N3898, N3368);
nor NOR2 (N7416, N7410, N3969);
and AND4 (N7417, N7405, N7010, N5425, N6666);
buf BUF1 (N7418, N7408);
not NOT1 (N7419, N7398);
or OR4 (N7420, N7416, N3911, N3380, N3100);
or OR4 (N7421, N7418, N278, N1400, N1305);
not NOT1 (N7422, N7409);
and AND2 (N7423, N7413, N3540);
and AND4 (N7424, N7415, N3639, N4726, N1659);
not NOT1 (N7425, N7424);
not NOT1 (N7426, N7407);
nand NAND4 (N7427, N7419, N3446, N7107, N1289);
nor NOR4 (N7428, N7425, N7177, N5334, N2556);
or OR4 (N7429, N7426, N5780, N795, N915);
or OR2 (N7430, N7422, N2836);
or OR4 (N7431, N7412, N42, N5625, N2944);
nor NOR2 (N7432, N7421, N6050);
xor XOR2 (N7433, N7417, N7036);
not NOT1 (N7434, N7420);
or OR3 (N7435, N7423, N5530, N3471);
and AND2 (N7436, N7435, N4680);
nor NOR3 (N7437, N7406, N4990, N1653);
not NOT1 (N7438, N7433);
and AND3 (N7439, N7432, N7236, N1429);
buf BUF1 (N7440, N7439);
buf BUF1 (N7441, N7436);
xor XOR2 (N7442, N7428, N4447);
nand NAND3 (N7443, N7437, N1967, N4295);
or OR4 (N7444, N7438, N3022, N6972, N193);
xor XOR2 (N7445, N7440, N933);
not NOT1 (N7446, N7444);
and AND4 (N7447, N7442, N709, N4965, N5686);
nand NAND4 (N7448, N7446, N103, N5036, N1220);
buf BUF1 (N7449, N7448);
or OR2 (N7450, N7441, N2660);
xor XOR2 (N7451, N7445, N4922);
nor NOR3 (N7452, N7450, N6422, N6938);
nor NOR4 (N7453, N7449, N2524, N225, N6551);
buf BUF1 (N7454, N7453);
and AND3 (N7455, N7434, N6248, N5406);
or OR4 (N7456, N7431, N4132, N4920, N3375);
buf BUF1 (N7457, N7455);
and AND4 (N7458, N7452, N2962, N2216, N1896);
nand NAND3 (N7459, N7458, N6880, N3725);
or OR3 (N7460, N7457, N4708, N2419);
not NOT1 (N7461, N7459);
not NOT1 (N7462, N7429);
xor XOR2 (N7463, N7456, N715);
and AND3 (N7464, N7462, N4254, N4030);
or OR3 (N7465, N7430, N1665, N1760);
and AND4 (N7466, N7463, N3170, N7378, N2944);
and AND2 (N7467, N7427, N7229);
and AND4 (N7468, N7454, N3125, N5735, N2361);
nor NOR4 (N7469, N7466, N1642, N5350, N4960);
nor NOR4 (N7470, N7467, N2675, N1053, N6936);
and AND3 (N7471, N7470, N980, N6642);
not NOT1 (N7472, N7465);
and AND2 (N7473, N7468, N1669);
nor NOR4 (N7474, N7471, N6712, N4341, N6785);
not NOT1 (N7475, N7447);
buf BUF1 (N7476, N7475);
nand NAND3 (N7477, N7451, N4735, N1294);
and AND4 (N7478, N7477, N1000, N1592, N3456);
nor NOR2 (N7479, N7476, N3742);
buf BUF1 (N7480, N7479);
or OR3 (N7481, N7474, N5040, N4354);
and AND3 (N7482, N7461, N5774, N2784);
nand NAND4 (N7483, N7478, N234, N603, N5049);
not NOT1 (N7484, N7480);
nor NOR3 (N7485, N7473, N3473, N2657);
not NOT1 (N7486, N7472);
nor NOR3 (N7487, N7484, N16, N5665);
or OR3 (N7488, N7481, N3829, N4928);
nor NOR2 (N7489, N7469, N6595);
not NOT1 (N7490, N7483);
nor NOR4 (N7491, N7464, N1286, N3205, N1648);
and AND2 (N7492, N7487, N5381);
nor NOR4 (N7493, N7489, N5289, N7083, N3099);
nand NAND2 (N7494, N7485, N1775);
buf BUF1 (N7495, N7493);
nand NAND4 (N7496, N7495, N3312, N7001, N1379);
buf BUF1 (N7497, N7496);
and AND2 (N7498, N7490, N2851);
not NOT1 (N7499, N7482);
and AND3 (N7500, N7443, N7223, N2753);
and AND4 (N7501, N7500, N2744, N4560, N7186);
buf BUF1 (N7502, N7492);
or OR4 (N7503, N7494, N1663, N6539, N3551);
buf BUF1 (N7504, N7503);
buf BUF1 (N7505, N7497);
and AND3 (N7506, N7486, N5629, N3321);
buf BUF1 (N7507, N7504);
nor NOR4 (N7508, N7491, N4419, N5609, N2174);
buf BUF1 (N7509, N7507);
and AND2 (N7510, N7505, N2164);
or OR4 (N7511, N7498, N6179, N7066, N6568);
not NOT1 (N7512, N7488);
buf BUF1 (N7513, N7508);
and AND4 (N7514, N7510, N873, N4033, N784);
nor NOR2 (N7515, N7506, N5032);
nand NAND3 (N7516, N7509, N2028, N5110);
not NOT1 (N7517, N7511);
nand NAND3 (N7518, N7517, N1544, N4989);
nand NAND2 (N7519, N7513, N1721);
buf BUF1 (N7520, N7502);
nand NAND3 (N7521, N7501, N4165, N660);
buf BUF1 (N7522, N7520);
nand NAND3 (N7523, N7499, N752, N2562);
or OR2 (N7524, N7514, N6650);
nand NAND2 (N7525, N7522, N3303);
and AND3 (N7526, N7518, N5272, N2686);
not NOT1 (N7527, N7519);
nor NOR2 (N7528, N7523, N6773);
buf BUF1 (N7529, N7512);
and AND2 (N7530, N7527, N7062);
nor NOR2 (N7531, N7460, N247);
and AND4 (N7532, N7529, N6294, N5817, N4592);
not NOT1 (N7533, N7532);
not NOT1 (N7534, N7531);
xor XOR2 (N7535, N7534, N592);
buf BUF1 (N7536, N7530);
buf BUF1 (N7537, N7526);
buf BUF1 (N7538, N7535);
nand NAND3 (N7539, N7538, N908, N2531);
nand NAND3 (N7540, N7539, N3664, N5814);
buf BUF1 (N7541, N7536);
not NOT1 (N7542, N7533);
xor XOR2 (N7543, N7537, N1462);
and AND2 (N7544, N7521, N886);
buf BUF1 (N7545, N7528);
and AND3 (N7546, N7515, N3561, N6812);
nand NAND2 (N7547, N7546, N870);
nand NAND2 (N7548, N7543, N1111);
not NOT1 (N7549, N7548);
or OR2 (N7550, N7524, N1488);
nand NAND4 (N7551, N7542, N3277, N145, N5941);
xor XOR2 (N7552, N7549, N2798);
and AND3 (N7553, N7544, N1214, N3759);
buf BUF1 (N7554, N7552);
nand NAND2 (N7555, N7540, N1375);
and AND3 (N7556, N7553, N3294, N5575);
buf BUF1 (N7557, N7555);
nor NOR2 (N7558, N7541, N6183);
not NOT1 (N7559, N7554);
and AND3 (N7560, N7525, N2687, N104);
not NOT1 (N7561, N7559);
xor XOR2 (N7562, N7560, N1941);
and AND3 (N7563, N7547, N5349, N3722);
or OR3 (N7564, N7561, N2605, N2554);
nor NOR4 (N7565, N7562, N2538, N1653, N3457);
xor XOR2 (N7566, N7564, N7494);
buf BUF1 (N7567, N7566);
nand NAND2 (N7568, N7516, N3150);
buf BUF1 (N7569, N7558);
buf BUF1 (N7570, N7551);
nor NOR4 (N7571, N7570, N6632, N5438, N6175);
nor NOR3 (N7572, N7568, N449, N6537);
nor NOR3 (N7573, N7557, N1009, N934);
and AND2 (N7574, N7545, N4802);
nor NOR4 (N7575, N7556, N7396, N200, N1867);
buf BUF1 (N7576, N7571);
and AND3 (N7577, N7574, N1221, N4947);
xor XOR2 (N7578, N7550, N2524);
or OR2 (N7579, N7569, N5817);
and AND3 (N7580, N7576, N943, N3576);
xor XOR2 (N7581, N7579, N7546);
nand NAND4 (N7582, N7578, N966, N6511, N2548);
nand NAND3 (N7583, N7575, N4687, N2347);
and AND3 (N7584, N7583, N1702, N1502);
xor XOR2 (N7585, N7577, N6334);
buf BUF1 (N7586, N7585);
buf BUF1 (N7587, N7565);
buf BUF1 (N7588, N7573);
nand NAND3 (N7589, N7572, N3360, N2588);
not NOT1 (N7590, N7584);
nor NOR2 (N7591, N7588, N3798);
not NOT1 (N7592, N7580);
not NOT1 (N7593, N7587);
and AND3 (N7594, N7581, N1459, N88);
or OR3 (N7595, N7563, N3679, N699);
xor XOR2 (N7596, N7567, N2121);
xor XOR2 (N7597, N7590, N2734);
or OR4 (N7598, N7591, N6967, N2980, N1988);
buf BUF1 (N7599, N7597);
and AND3 (N7600, N7596, N5117, N3338);
nand NAND3 (N7601, N7598, N3720, N3347);
buf BUF1 (N7602, N7599);
and AND4 (N7603, N7582, N2762, N474, N1062);
buf BUF1 (N7604, N7592);
xor XOR2 (N7605, N7586, N1629);
buf BUF1 (N7606, N7589);
xor XOR2 (N7607, N7600, N1818);
not NOT1 (N7608, N7595);
nor NOR3 (N7609, N7605, N1933, N1753);
nand NAND2 (N7610, N7608, N6117);
or OR4 (N7611, N7594, N2505, N5796, N5275);
buf BUF1 (N7612, N7602);
or OR3 (N7613, N7606, N3946, N2584);
xor XOR2 (N7614, N7607, N4357);
buf BUF1 (N7615, N7604);
and AND4 (N7616, N7615, N6863, N5301, N7480);
nor NOR2 (N7617, N7609, N665);
nor NOR3 (N7618, N7601, N4020, N2716);
and AND2 (N7619, N7616, N5935);
or OR4 (N7620, N7611, N4756, N2590, N5907);
nor NOR2 (N7621, N7603, N6220);
nor NOR3 (N7622, N7621, N1295, N4717);
nor NOR2 (N7623, N7614, N5705);
and AND3 (N7624, N7618, N683, N3651);
not NOT1 (N7625, N7623);
xor XOR2 (N7626, N7624, N4806);
nor NOR4 (N7627, N7619, N6369, N2369, N2930);
nor NOR3 (N7628, N7626, N4704, N2457);
nand NAND3 (N7629, N7622, N3226, N1496);
buf BUF1 (N7630, N7613);
or OR3 (N7631, N7629, N6760, N4757);
xor XOR2 (N7632, N7627, N1153);
buf BUF1 (N7633, N7628);
nand NAND4 (N7634, N7625, N5232, N2323, N3937);
or OR4 (N7635, N7617, N5875, N2890, N4442);
and AND2 (N7636, N7630, N2847);
buf BUF1 (N7637, N7631);
nor NOR4 (N7638, N7634, N5186, N4552, N5748);
not NOT1 (N7639, N7637);
nor NOR3 (N7640, N7610, N3419, N2732);
buf BUF1 (N7641, N7633);
not NOT1 (N7642, N7635);
or OR3 (N7643, N7639, N3351, N5410);
nand NAND4 (N7644, N7638, N1865, N6948, N3833);
or OR2 (N7645, N7644, N3381);
buf BUF1 (N7646, N7593);
nor NOR2 (N7647, N7632, N50);
buf BUF1 (N7648, N7612);
not NOT1 (N7649, N7648);
not NOT1 (N7650, N7645);
or OR3 (N7651, N7649, N5599, N5355);
not NOT1 (N7652, N7643);
xor XOR2 (N7653, N7620, N3267);
nor NOR4 (N7654, N7652, N3329, N2375, N7456);
nand NAND4 (N7655, N7640, N5375, N5467, N1168);
nand NAND4 (N7656, N7646, N5227, N3322, N2125);
nand NAND3 (N7657, N7636, N2370, N3018);
and AND3 (N7658, N7656, N4930, N2902);
nor NOR2 (N7659, N7642, N31);
not NOT1 (N7660, N7657);
or OR4 (N7661, N7641, N6516, N1842, N1591);
xor XOR2 (N7662, N7660, N6937);
or OR2 (N7663, N7651, N2907);
and AND2 (N7664, N7650, N4696);
xor XOR2 (N7665, N7659, N1003);
not NOT1 (N7666, N7663);
nand NAND4 (N7667, N7662, N1228, N3184, N5248);
buf BUF1 (N7668, N7653);
and AND2 (N7669, N7655, N2672);
buf BUF1 (N7670, N7669);
and AND2 (N7671, N7658, N6621);
and AND3 (N7672, N7670, N2588, N6479);
not NOT1 (N7673, N7654);
or OR2 (N7674, N7668, N238);
xor XOR2 (N7675, N7672, N914);
or OR3 (N7676, N7661, N5184, N2650);
or OR3 (N7677, N7676, N2986, N655);
buf BUF1 (N7678, N7647);
xor XOR2 (N7679, N7677, N6670);
buf BUF1 (N7680, N7667);
xor XOR2 (N7681, N7665, N4946);
not NOT1 (N7682, N7678);
or OR2 (N7683, N7673, N580);
nor NOR2 (N7684, N7680, N7170);
not NOT1 (N7685, N7679);
not NOT1 (N7686, N7666);
xor XOR2 (N7687, N7684, N3297);
and AND3 (N7688, N7686, N2546, N2895);
buf BUF1 (N7689, N7683);
not NOT1 (N7690, N7688);
not NOT1 (N7691, N7689);
nor NOR3 (N7692, N7690, N6117, N5351);
or OR4 (N7693, N7681, N6417, N1963, N5151);
xor XOR2 (N7694, N7692, N5367);
buf BUF1 (N7695, N7693);
and AND3 (N7696, N7674, N7358, N4935);
nor NOR3 (N7697, N7682, N6657, N6678);
and AND2 (N7698, N7694, N3987);
not NOT1 (N7699, N7695);
nor NOR4 (N7700, N7697, N1465, N1819, N6096);
or OR3 (N7701, N7671, N2884, N64);
or OR2 (N7702, N7685, N2793);
xor XOR2 (N7703, N7701, N3936);
and AND2 (N7704, N7696, N4951);
nand NAND3 (N7705, N7704, N659, N1420);
not NOT1 (N7706, N7703);
or OR3 (N7707, N7706, N363, N1117);
buf BUF1 (N7708, N7698);
or OR2 (N7709, N7687, N722);
buf BUF1 (N7710, N7702);
or OR4 (N7711, N7708, N1315, N5466, N4158);
nand NAND3 (N7712, N7709, N6547, N3651);
nor NOR2 (N7713, N7675, N7120);
xor XOR2 (N7714, N7699, N4222);
xor XOR2 (N7715, N7691, N7274);
nor NOR4 (N7716, N7711, N3329, N6046, N3095);
nand NAND2 (N7717, N7714, N991);
or OR3 (N7718, N7710, N5213, N5777);
xor XOR2 (N7719, N7716, N4256);
not NOT1 (N7720, N7719);
not NOT1 (N7721, N7718);
or OR3 (N7722, N7721, N2090, N726);
nand NAND4 (N7723, N7712, N7677, N3029, N5562);
or OR4 (N7724, N7664, N5550, N4313, N5034);
or OR4 (N7725, N7724, N29, N1421, N7067);
nand NAND4 (N7726, N7700, N6045, N7257, N659);
nand NAND3 (N7727, N7715, N1011, N3689);
xor XOR2 (N7728, N7727, N1615);
and AND3 (N7729, N7705, N5613, N3363);
nor NOR2 (N7730, N7729, N6667);
nand NAND4 (N7731, N7717, N3310, N7629, N1833);
xor XOR2 (N7732, N7728, N7233);
buf BUF1 (N7733, N7731);
xor XOR2 (N7734, N7726, N924);
buf BUF1 (N7735, N7733);
xor XOR2 (N7736, N7722, N4316);
nand NAND4 (N7737, N7720, N2165, N1651, N3002);
nand NAND3 (N7738, N7737, N5636, N3622);
xor XOR2 (N7739, N7736, N7446);
nor NOR4 (N7740, N7707, N7267, N4844, N4140);
nor NOR4 (N7741, N7732, N3646, N6397, N5784);
not NOT1 (N7742, N7725);
buf BUF1 (N7743, N7734);
or OR3 (N7744, N7740, N188, N598);
not NOT1 (N7745, N7742);
xor XOR2 (N7746, N7738, N4795);
and AND4 (N7747, N7741, N2239, N7035, N6178);
not NOT1 (N7748, N7745);
xor XOR2 (N7749, N7735, N5886);
nand NAND2 (N7750, N7744, N6948);
nor NOR3 (N7751, N7739, N835, N2555);
nor NOR3 (N7752, N7749, N704, N6767);
nor NOR3 (N7753, N7743, N3385, N5213);
nand NAND4 (N7754, N7746, N7014, N3233, N4294);
and AND3 (N7755, N7751, N7029, N5490);
or OR4 (N7756, N7752, N3233, N5669, N7505);
and AND2 (N7757, N7713, N7498);
nand NAND2 (N7758, N7750, N7456);
buf BUF1 (N7759, N7754);
not NOT1 (N7760, N7755);
nand NAND2 (N7761, N7756, N6757);
nand NAND2 (N7762, N7747, N4455);
not NOT1 (N7763, N7730);
nor NOR4 (N7764, N7753, N5285, N774, N455);
and AND4 (N7765, N7762, N7655, N6625, N2650);
nand NAND3 (N7766, N7761, N6047, N3201);
xor XOR2 (N7767, N7748, N4630);
or OR4 (N7768, N7766, N4330, N7314, N5832);
xor XOR2 (N7769, N7763, N6640);
or OR4 (N7770, N7757, N802, N5072, N7672);
buf BUF1 (N7771, N7769);
or OR4 (N7772, N7759, N4743, N2554, N3860);
or OR4 (N7773, N7760, N1938, N231, N2918);
and AND4 (N7774, N7765, N5336, N1999, N2824);
buf BUF1 (N7775, N7768);
nor NOR4 (N7776, N7764, N1146, N3703, N7298);
and AND3 (N7777, N7776, N2040, N2324);
or OR2 (N7778, N7777, N2692);
nand NAND4 (N7779, N7758, N3654, N7605, N7559);
or OR2 (N7780, N7771, N7103);
xor XOR2 (N7781, N7774, N1383);
xor XOR2 (N7782, N7773, N2276);
xor XOR2 (N7783, N7775, N7598);
xor XOR2 (N7784, N7782, N6225);
xor XOR2 (N7785, N7780, N2941);
buf BUF1 (N7786, N7770);
buf BUF1 (N7787, N7783);
or OR2 (N7788, N7787, N2057);
not NOT1 (N7789, N7788);
xor XOR2 (N7790, N7786, N4296);
and AND4 (N7791, N7778, N3288, N4178, N4827);
xor XOR2 (N7792, N7767, N764);
not NOT1 (N7793, N7789);
or OR2 (N7794, N7779, N2584);
and AND3 (N7795, N7784, N4479, N5388);
and AND3 (N7796, N7790, N4972, N2538);
and AND3 (N7797, N7794, N4875, N1897);
buf BUF1 (N7798, N7795);
or OR4 (N7799, N7772, N4476, N7077, N2599);
buf BUF1 (N7800, N7791);
or OR4 (N7801, N7785, N713, N3695, N6698);
and AND4 (N7802, N7801, N2989, N2850, N4352);
nand NAND3 (N7803, N7793, N4146, N1405);
and AND4 (N7804, N7800, N1815, N5118, N4127);
not NOT1 (N7805, N7803);
and AND3 (N7806, N7798, N903, N3125);
buf BUF1 (N7807, N7796);
not NOT1 (N7808, N7807);
nand NAND4 (N7809, N7799, N2392, N3018, N644);
xor XOR2 (N7810, N7723, N6045);
or OR3 (N7811, N7792, N5059, N3843);
xor XOR2 (N7812, N7797, N839);
buf BUF1 (N7813, N7781);
buf BUF1 (N7814, N7812);
xor XOR2 (N7815, N7806, N7523);
nor NOR4 (N7816, N7805, N1088, N2614, N4590);
not NOT1 (N7817, N7809);
nor NOR2 (N7818, N7813, N5196);
or OR4 (N7819, N7804, N6963, N1783, N5208);
buf BUF1 (N7820, N7816);
nor NOR2 (N7821, N7811, N3152);
nor NOR4 (N7822, N7817, N1185, N246, N6153);
nand NAND4 (N7823, N7810, N4788, N3547, N7635);
nor NOR2 (N7824, N7814, N6992);
buf BUF1 (N7825, N7819);
not NOT1 (N7826, N7822);
or OR4 (N7827, N7820, N4671, N1853, N5180);
not NOT1 (N7828, N7802);
and AND3 (N7829, N7824, N3676, N4636);
and AND3 (N7830, N7808, N5521, N1413);
not NOT1 (N7831, N7828);
not NOT1 (N7832, N7831);
nand NAND3 (N7833, N7829, N2769, N3221);
and AND3 (N7834, N7830, N6249, N2709);
buf BUF1 (N7835, N7826);
and AND3 (N7836, N7821, N837, N5285);
or OR3 (N7837, N7836, N5917, N6034);
or OR4 (N7838, N7823, N201, N6571, N596);
xor XOR2 (N7839, N7827, N3091);
not NOT1 (N7840, N7832);
nor NOR4 (N7841, N7825, N3155, N1238, N2646);
nor NOR2 (N7842, N7837, N4185);
nand NAND4 (N7843, N7835, N2015, N2729, N107);
xor XOR2 (N7844, N7834, N203);
not NOT1 (N7845, N7843);
nand NAND4 (N7846, N7842, N4034, N3029, N5793);
or OR3 (N7847, N7818, N348, N2404);
or OR3 (N7848, N7840, N7043, N6814);
xor XOR2 (N7849, N7848, N7558);
xor XOR2 (N7850, N7815, N5244);
not NOT1 (N7851, N7841);
or OR4 (N7852, N7850, N6051, N179, N3745);
and AND2 (N7853, N7844, N7804);
not NOT1 (N7854, N7851);
or OR3 (N7855, N7853, N7689, N6820);
and AND3 (N7856, N7847, N3094, N6521);
nor NOR3 (N7857, N7855, N5723, N462);
and AND4 (N7858, N7849, N3108, N3393, N2520);
buf BUF1 (N7859, N7845);
nand NAND3 (N7860, N7856, N4048, N6905);
nand NAND4 (N7861, N7857, N5138, N2227, N4190);
xor XOR2 (N7862, N7839, N7018);
not NOT1 (N7863, N7862);
xor XOR2 (N7864, N7838, N7065);
xor XOR2 (N7865, N7863, N1599);
xor XOR2 (N7866, N7854, N1879);
nand NAND2 (N7867, N7859, N647);
nand NAND3 (N7868, N7852, N5998, N3067);
nand NAND3 (N7869, N7858, N7843, N4538);
xor XOR2 (N7870, N7833, N4324);
or OR4 (N7871, N7866, N1287, N1473, N7355);
nand NAND4 (N7872, N7846, N3659, N1383, N4023);
or OR3 (N7873, N7869, N7408, N1877);
nand NAND2 (N7874, N7867, N6064);
not NOT1 (N7875, N7873);
nand NAND3 (N7876, N7875, N6697, N1529);
xor XOR2 (N7877, N7874, N4610);
not NOT1 (N7878, N7871);
and AND3 (N7879, N7876, N4472, N6858);
nand NAND3 (N7880, N7864, N4867, N3984);
nor NOR2 (N7881, N7870, N5380);
not NOT1 (N7882, N7879);
nand NAND3 (N7883, N7865, N6858, N3090);
xor XOR2 (N7884, N7868, N67);
buf BUF1 (N7885, N7877);
or OR4 (N7886, N7880, N4050, N5690, N272);
nand NAND4 (N7887, N7884, N5644, N845, N7013);
xor XOR2 (N7888, N7860, N4634);
xor XOR2 (N7889, N7883, N2338);
and AND3 (N7890, N7882, N3282, N5641);
nand NAND3 (N7891, N7885, N2747, N7218);
not NOT1 (N7892, N7888);
and AND2 (N7893, N7889, N5883);
not NOT1 (N7894, N7886);
not NOT1 (N7895, N7878);
buf BUF1 (N7896, N7881);
not NOT1 (N7897, N7895);
nor NOR2 (N7898, N7896, N1508);
buf BUF1 (N7899, N7892);
buf BUF1 (N7900, N7861);
xor XOR2 (N7901, N7893, N3930);
buf BUF1 (N7902, N7901);
nand NAND4 (N7903, N7887, N1997, N2098, N5068);
not NOT1 (N7904, N7903);
nor NOR2 (N7905, N7891, N2535);
nor NOR2 (N7906, N7894, N282);
and AND3 (N7907, N7906, N3516, N746);
xor XOR2 (N7908, N7905, N6976);
and AND3 (N7909, N7872, N886, N3833);
nand NAND4 (N7910, N7898, N7449, N4487, N6742);
and AND2 (N7911, N7899, N3265);
xor XOR2 (N7912, N7911, N4225);
or OR4 (N7913, N7900, N2652, N1149, N2186);
xor XOR2 (N7914, N7907, N4685);
or OR4 (N7915, N7902, N3096, N6254, N4198);
and AND2 (N7916, N7904, N6083);
xor XOR2 (N7917, N7890, N7274);
and AND4 (N7918, N7915, N1383, N3113, N3328);
or OR3 (N7919, N7916, N7867, N5565);
or OR3 (N7920, N7910, N3586, N2943);
not NOT1 (N7921, N7897);
not NOT1 (N7922, N7912);
not NOT1 (N7923, N7917);
and AND3 (N7924, N7919, N4198, N7613);
and AND4 (N7925, N7908, N585, N4860, N3454);
buf BUF1 (N7926, N7923);
or OR4 (N7927, N7913, N771, N612, N6729);
and AND2 (N7928, N7918, N495);
buf BUF1 (N7929, N7914);
xor XOR2 (N7930, N7909, N4020);
nand NAND2 (N7931, N7925, N7624);
not NOT1 (N7932, N7931);
not NOT1 (N7933, N7920);
nor NOR4 (N7934, N7922, N4478, N4230, N7358);
nor NOR3 (N7935, N7921, N850, N777);
or OR2 (N7936, N7935, N2847);
or OR2 (N7937, N7924, N4761);
xor XOR2 (N7938, N7933, N6923);
nand NAND2 (N7939, N7934, N4450);
or OR4 (N7940, N7926, N2642, N5636, N2346);
nand NAND3 (N7941, N7937, N4349, N6555);
not NOT1 (N7942, N7940);
buf BUF1 (N7943, N7928);
nand NAND4 (N7944, N7943, N6163, N543, N3683);
not NOT1 (N7945, N7941);
or OR3 (N7946, N7938, N3089, N5324);
or OR4 (N7947, N7932, N5825, N4088, N1567);
buf BUF1 (N7948, N7929);
nand NAND4 (N7949, N7939, N5541, N383, N856);
nor NOR3 (N7950, N7947, N7809, N488);
not NOT1 (N7951, N7948);
and AND2 (N7952, N7950, N2767);
nor NOR2 (N7953, N7946, N507);
xor XOR2 (N7954, N7949, N7951);
nor NOR3 (N7955, N4503, N2763, N5096);
buf BUF1 (N7956, N7952);
nand NAND3 (N7957, N7927, N4544, N4469);
and AND2 (N7958, N7936, N1960);
xor XOR2 (N7959, N7958, N941);
buf BUF1 (N7960, N7942);
nand NAND4 (N7961, N7955, N3700, N3307, N6102);
or OR3 (N7962, N7953, N858, N1826);
or OR2 (N7963, N7944, N5659);
buf BUF1 (N7964, N7962);
xor XOR2 (N7965, N7954, N4731);
or OR3 (N7966, N7930, N7086, N4396);
buf BUF1 (N7967, N7963);
buf BUF1 (N7968, N7959);
and AND3 (N7969, N7966, N4329, N4808);
buf BUF1 (N7970, N7969);
nand NAND3 (N7971, N7956, N1339, N5356);
xor XOR2 (N7972, N7971, N7071);
not NOT1 (N7973, N7964);
or OR3 (N7974, N7967, N7057, N5731);
not NOT1 (N7975, N7968);
buf BUF1 (N7976, N7974);
nand NAND3 (N7977, N7976, N7470, N3485);
xor XOR2 (N7978, N7972, N6573);
and AND3 (N7979, N7970, N802, N4058);
and AND4 (N7980, N7973, N2032, N4556, N5286);
nand NAND3 (N7981, N7980, N5496, N7704);
buf BUF1 (N7982, N7975);
or OR3 (N7983, N7981, N2253, N1012);
buf BUF1 (N7984, N7978);
xor XOR2 (N7985, N7960, N7556);
and AND2 (N7986, N7965, N6438);
or OR3 (N7987, N7982, N1282, N3937);
and AND2 (N7988, N7977, N4911);
or OR4 (N7989, N7988, N5176, N2241, N744);
or OR3 (N7990, N7961, N6586, N7788);
buf BUF1 (N7991, N7989);
buf BUF1 (N7992, N7991);
nand NAND4 (N7993, N7986, N7503, N532, N7332);
and AND3 (N7994, N7945, N2995, N1071);
and AND3 (N7995, N7979, N4282, N7050);
and AND2 (N7996, N7983, N7554);
nand NAND3 (N7997, N7993, N5262, N7601);
and AND4 (N7998, N7987, N5204, N1812, N5917);
nand NAND4 (N7999, N7996, N5839, N6086, N4278);
nor NOR3 (N8000, N7999, N5679, N3420);
not NOT1 (N8001, N7957);
or OR4 (N8002, N7994, N5156, N393, N2782);
nor NOR2 (N8003, N7997, N6067);
and AND2 (N8004, N8002, N3391);
or OR2 (N8005, N8000, N7771);
nand NAND2 (N8006, N8001, N6026);
xor XOR2 (N8007, N7998, N2538);
not NOT1 (N8008, N7992);
not NOT1 (N8009, N7984);
xor XOR2 (N8010, N8004, N2979);
nor NOR3 (N8011, N7990, N942, N2033);
not NOT1 (N8012, N8007);
and AND2 (N8013, N8005, N7300);
not NOT1 (N8014, N7995);
not NOT1 (N8015, N8009);
buf BUF1 (N8016, N8013);
xor XOR2 (N8017, N7985, N7231);
nor NOR2 (N8018, N8012, N5284);
buf BUF1 (N8019, N8006);
buf BUF1 (N8020, N8011);
not NOT1 (N8021, N8016);
or OR4 (N8022, N8015, N3685, N7276, N2815);
xor XOR2 (N8023, N8022, N792);
nor NOR4 (N8024, N8003, N327, N1866, N3901);
not NOT1 (N8025, N8010);
nor NOR4 (N8026, N8021, N372, N5770, N315);
or OR3 (N8027, N8017, N2486, N781);
buf BUF1 (N8028, N8014);
or OR2 (N8029, N8026, N7860);
or OR4 (N8030, N8023, N2151, N149, N1518);
and AND4 (N8031, N8020, N2537, N5047, N4837);
nand NAND3 (N8032, N8029, N4174, N2436);
xor XOR2 (N8033, N8030, N1657);
buf BUF1 (N8034, N8028);
and AND2 (N8035, N8031, N7676);
not NOT1 (N8036, N8027);
and AND4 (N8037, N8033, N4928, N4103, N1335);
buf BUF1 (N8038, N8036);
not NOT1 (N8039, N8037);
buf BUF1 (N8040, N8035);
not NOT1 (N8041, N8039);
and AND2 (N8042, N8032, N4865);
nand NAND4 (N8043, N8038, N3142, N1556, N6347);
and AND4 (N8044, N8041, N6671, N4607, N5390);
buf BUF1 (N8045, N8008);
not NOT1 (N8046, N8034);
buf BUF1 (N8047, N8046);
buf BUF1 (N8048, N8019);
or OR4 (N8049, N8048, N3975, N6244, N7583);
xor XOR2 (N8050, N8018, N2415);
xor XOR2 (N8051, N8044, N442);
nand NAND4 (N8052, N8024, N1532, N7068, N3253);
and AND4 (N8053, N8043, N2519, N271, N1742);
not NOT1 (N8054, N8042);
nand NAND2 (N8055, N8045, N5987);
not NOT1 (N8056, N8040);
buf BUF1 (N8057, N8047);
not NOT1 (N8058, N8051);
nor NOR2 (N8059, N8049, N1877);
buf BUF1 (N8060, N8057);
not NOT1 (N8061, N8052);
or OR4 (N8062, N8059, N530, N2259, N1512);
or OR2 (N8063, N8025, N4849);
nor NOR2 (N8064, N8063, N2172);
and AND2 (N8065, N8062, N136);
nand NAND4 (N8066, N8050, N6609, N5875, N3333);
xor XOR2 (N8067, N8055, N710);
nand NAND4 (N8068, N8067, N4625, N1779, N6740);
and AND2 (N8069, N8068, N6093);
nor NOR2 (N8070, N8053, N2610);
nor NOR3 (N8071, N8058, N2516, N5400);
nor NOR3 (N8072, N8056, N6894, N7861);
buf BUF1 (N8073, N8064);
xor XOR2 (N8074, N8065, N5628);
and AND3 (N8075, N8060, N5684, N5780);
xor XOR2 (N8076, N8061, N4245);
xor XOR2 (N8077, N8070, N4608);
nor NOR3 (N8078, N8066, N4908, N2964);
not NOT1 (N8079, N8069);
not NOT1 (N8080, N8074);
and AND2 (N8081, N8073, N5631);
nand NAND3 (N8082, N8079, N1724, N5350);
or OR3 (N8083, N8082, N5153, N637);
nor NOR2 (N8084, N8080, N5325);
nand NAND2 (N8085, N8071, N6451);
nor NOR3 (N8086, N8085, N6762, N1011);
and AND3 (N8087, N8076, N2496, N7558);
nor NOR2 (N8088, N8087, N2135);
and AND2 (N8089, N8083, N6827);
not NOT1 (N8090, N8089);
and AND2 (N8091, N8078, N5078);
not NOT1 (N8092, N8075);
nor NOR2 (N8093, N8086, N5877);
and AND3 (N8094, N8054, N3632, N681);
or OR4 (N8095, N8092, N5296, N6000, N7153);
xor XOR2 (N8096, N8090, N6722);
nand NAND4 (N8097, N8093, N7952, N6556, N6999);
nand NAND4 (N8098, N8077, N5996, N7097, N577);
not NOT1 (N8099, N8095);
and AND2 (N8100, N8081, N6371);
nor NOR4 (N8101, N8088, N250, N5370, N7393);
xor XOR2 (N8102, N8100, N2950);
nor NOR4 (N8103, N8102, N2222, N2013, N6505);
buf BUF1 (N8104, N8096);
or OR2 (N8105, N8103, N3313);
and AND2 (N8106, N8105, N6745);
buf BUF1 (N8107, N8072);
xor XOR2 (N8108, N8107, N7891);
and AND3 (N8109, N8098, N5834, N2548);
not NOT1 (N8110, N8106);
and AND2 (N8111, N8084, N865);
and AND3 (N8112, N8110, N1766, N5445);
nor NOR2 (N8113, N8094, N6885);
nor NOR4 (N8114, N8109, N4237, N5142, N6536);
and AND2 (N8115, N8091, N5450);
or OR3 (N8116, N8114, N2201, N7024);
xor XOR2 (N8117, N8113, N1391);
nor NOR4 (N8118, N8099, N5244, N3009, N5411);
buf BUF1 (N8119, N8116);
not NOT1 (N8120, N8097);
nand NAND4 (N8121, N8104, N6941, N1132, N6344);
or OR4 (N8122, N8111, N5845, N5453, N759);
or OR2 (N8123, N8117, N3259);
buf BUF1 (N8124, N8123);
xor XOR2 (N8125, N8121, N6863);
or OR3 (N8126, N8118, N6824, N6245);
nand NAND3 (N8127, N8108, N4400, N5424);
or OR2 (N8128, N8120, N965);
xor XOR2 (N8129, N8125, N4973);
buf BUF1 (N8130, N8127);
nand NAND2 (N8131, N8122, N2872);
or OR4 (N8132, N8128, N5426, N1660, N4712);
nand NAND4 (N8133, N8112, N3280, N1267, N6919);
xor XOR2 (N8134, N8119, N4975);
or OR2 (N8135, N8131, N1838);
not NOT1 (N8136, N8126);
nor NOR2 (N8137, N8136, N14);
nor NOR4 (N8138, N8130, N4464, N3210, N7390);
buf BUF1 (N8139, N8134);
buf BUF1 (N8140, N8137);
or OR2 (N8141, N8133, N3715);
buf BUF1 (N8142, N8132);
or OR4 (N8143, N8101, N1408, N3499, N5206);
or OR3 (N8144, N8129, N561, N3211);
or OR2 (N8145, N8141, N6541);
or OR2 (N8146, N8142, N3067);
not NOT1 (N8147, N8140);
not NOT1 (N8148, N8143);
not NOT1 (N8149, N8115);
or OR4 (N8150, N8148, N3528, N5244, N6211);
nand NAND3 (N8151, N8147, N4701, N6153);
and AND4 (N8152, N8139, N757, N3446, N7218);
not NOT1 (N8153, N8135);
or OR4 (N8154, N8145, N7975, N7400, N2151);
xor XOR2 (N8155, N8150, N3787);
or OR4 (N8156, N8146, N5385, N2699, N4870);
xor XOR2 (N8157, N8153, N2789);
or OR3 (N8158, N8154, N1889, N3630);
nand NAND2 (N8159, N8149, N662);
nor NOR2 (N8160, N8155, N8005);
xor XOR2 (N8161, N8160, N6300);
nand NAND2 (N8162, N8151, N1757);
and AND2 (N8163, N8159, N6511);
and AND3 (N8164, N8163, N2452, N4288);
nor NOR2 (N8165, N8164, N7907);
buf BUF1 (N8166, N8144);
buf BUF1 (N8167, N8156);
not NOT1 (N8168, N8138);
not NOT1 (N8169, N8165);
or OR4 (N8170, N8162, N96, N6613, N3052);
and AND2 (N8171, N8168, N7668);
not NOT1 (N8172, N8158);
nor NOR3 (N8173, N8167, N3561, N2106);
buf BUF1 (N8174, N8157);
or OR2 (N8175, N8172, N1741);
or OR2 (N8176, N8169, N3904);
nor NOR4 (N8177, N8174, N4325, N7646, N6737);
and AND3 (N8178, N8161, N2392, N701);
nand NAND3 (N8179, N8171, N5138, N2531);
and AND2 (N8180, N8170, N5524);
nand NAND4 (N8181, N8124, N121, N2763, N2843);
xor XOR2 (N8182, N8176, N3216);
or OR2 (N8183, N8179, N3688);
not NOT1 (N8184, N8175);
nand NAND4 (N8185, N8152, N7929, N5214, N4437);
and AND4 (N8186, N8181, N418, N7233, N1263);
xor XOR2 (N8187, N8184, N136);
or OR2 (N8188, N8183, N7068);
nand NAND4 (N8189, N8182, N1330, N6948, N1709);
or OR2 (N8190, N8188, N6708);
buf BUF1 (N8191, N8180);
not NOT1 (N8192, N8178);
not NOT1 (N8193, N8177);
or OR3 (N8194, N8189, N5163, N7026);
buf BUF1 (N8195, N8173);
nand NAND4 (N8196, N8194, N290, N2095, N6038);
not NOT1 (N8197, N8190);
xor XOR2 (N8198, N8191, N7491);
nor NOR2 (N8199, N8192, N1292);
nor NOR2 (N8200, N8198, N1013);
xor XOR2 (N8201, N8195, N5852);
buf BUF1 (N8202, N8187);
nand NAND3 (N8203, N8196, N2051, N26);
or OR4 (N8204, N8193, N5209, N5795, N6819);
not NOT1 (N8205, N8185);
not NOT1 (N8206, N8202);
xor XOR2 (N8207, N8197, N6734);
nand NAND2 (N8208, N8186, N6664);
xor XOR2 (N8209, N8207, N5107);
xor XOR2 (N8210, N8204, N3360);
buf BUF1 (N8211, N8208);
or OR4 (N8212, N8200, N7796, N7319, N6501);
buf BUF1 (N8213, N8210);
and AND2 (N8214, N8205, N586);
not NOT1 (N8215, N8206);
nor NOR3 (N8216, N8213, N1932, N3353);
buf BUF1 (N8217, N8211);
not NOT1 (N8218, N8212);
buf BUF1 (N8219, N8217);
xor XOR2 (N8220, N8214, N4156);
not NOT1 (N8221, N8209);
nand NAND2 (N8222, N8219, N6028);
nor NOR2 (N8223, N8203, N3158);
nand NAND3 (N8224, N8220, N1965, N8079);
or OR2 (N8225, N8222, N710);
buf BUF1 (N8226, N8201);
xor XOR2 (N8227, N8223, N3401);
nand NAND2 (N8228, N8227, N3824);
or OR2 (N8229, N8224, N6852);
xor XOR2 (N8230, N8215, N6001);
not NOT1 (N8231, N8199);
or OR2 (N8232, N8226, N4777);
and AND2 (N8233, N8225, N2822);
nor NOR4 (N8234, N8221, N4583, N5337, N3683);
nand NAND2 (N8235, N8228, N4122);
buf BUF1 (N8236, N8216);
and AND2 (N8237, N8235, N7999);
not NOT1 (N8238, N8166);
xor XOR2 (N8239, N8231, N1188);
nand NAND2 (N8240, N8232, N5014);
buf BUF1 (N8241, N8234);
and AND2 (N8242, N8240, N4178);
buf BUF1 (N8243, N8242);
and AND3 (N8244, N8241, N6986, N4020);
xor XOR2 (N8245, N8244, N4697);
and AND3 (N8246, N8239, N1046, N930);
and AND2 (N8247, N8238, N7837);
and AND4 (N8248, N8236, N4205, N5113, N3629);
nor NOR4 (N8249, N8218, N20, N1067, N7918);
or OR3 (N8250, N8246, N467, N2542);
buf BUF1 (N8251, N8247);
not NOT1 (N8252, N8250);
or OR2 (N8253, N8249, N3497);
and AND2 (N8254, N8243, N1008);
not NOT1 (N8255, N8254);
nor NOR2 (N8256, N8252, N7689);
not NOT1 (N8257, N8248);
nand NAND3 (N8258, N8233, N7123, N2835);
not NOT1 (N8259, N8255);
and AND4 (N8260, N8230, N6051, N6959, N3360);
and AND4 (N8261, N8256, N5740, N3572, N6788);
not NOT1 (N8262, N8245);
or OR4 (N8263, N8237, N3142, N177, N5086);
nor NOR4 (N8264, N8263, N1426, N1450, N1834);
not NOT1 (N8265, N8259);
xor XOR2 (N8266, N8257, N7142);
or OR4 (N8267, N8258, N6780, N6501, N5606);
nor NOR4 (N8268, N8265, N7080, N1151, N8219);
or OR2 (N8269, N8229, N1138);
buf BUF1 (N8270, N8260);
buf BUF1 (N8271, N8251);
nand NAND2 (N8272, N8268, N5536);
and AND4 (N8273, N8261, N2836, N206, N299);
not NOT1 (N8274, N8270);
nor NOR3 (N8275, N8269, N2792, N719);
nand NAND2 (N8276, N8253, N311);
and AND4 (N8277, N8266, N2730, N4194, N6573);
nand NAND4 (N8278, N8271, N5915, N5380, N6012);
not NOT1 (N8279, N8262);
nand NAND3 (N8280, N8272, N7069, N4190);
nor NOR4 (N8281, N8275, N4867, N2036, N2741);
nor NOR3 (N8282, N8281, N641, N8084);
xor XOR2 (N8283, N8267, N1616);
xor XOR2 (N8284, N8279, N6700);
nand NAND4 (N8285, N8284, N6212, N5242, N5581);
buf BUF1 (N8286, N8273);
nor NOR4 (N8287, N8283, N4341, N2310, N8073);
buf BUF1 (N8288, N8274);
xor XOR2 (N8289, N8280, N5832);
buf BUF1 (N8290, N8287);
and AND3 (N8291, N8289, N3948, N3029);
nand NAND4 (N8292, N8264, N7837, N1994, N3608);
nand NAND2 (N8293, N8282, N2021);
not NOT1 (N8294, N8278);
buf BUF1 (N8295, N8276);
xor XOR2 (N8296, N8285, N5828);
nor NOR2 (N8297, N8286, N486);
not NOT1 (N8298, N8294);
or OR4 (N8299, N8292, N561, N2833, N1597);
nor NOR4 (N8300, N8295, N622, N4778, N4360);
or OR3 (N8301, N8300, N4634, N1797);
xor XOR2 (N8302, N8277, N4862);
or OR3 (N8303, N8297, N6298, N1979);
nand NAND2 (N8304, N8303, N5127);
not NOT1 (N8305, N8304);
and AND4 (N8306, N8298, N2058, N6812, N6762);
buf BUF1 (N8307, N8290);
nor NOR3 (N8308, N8305, N5593, N5595);
not NOT1 (N8309, N8306);
buf BUF1 (N8310, N8296);
nand NAND4 (N8311, N8291, N7983, N7563, N5933);
xor XOR2 (N8312, N8301, N7372);
xor XOR2 (N8313, N8312, N3418);
nand NAND2 (N8314, N8311, N938);
not NOT1 (N8315, N8299);
xor XOR2 (N8316, N8288, N5615);
not NOT1 (N8317, N8307);
buf BUF1 (N8318, N8302);
not NOT1 (N8319, N8313);
nor NOR3 (N8320, N8317, N6574, N219);
buf BUF1 (N8321, N8308);
nand NAND2 (N8322, N8314, N873);
nand NAND4 (N8323, N8316, N3567, N2772, N5375);
or OR4 (N8324, N8309, N4843, N2890, N4210);
not NOT1 (N8325, N8315);
nand NAND4 (N8326, N8318, N2408, N235, N5026);
and AND4 (N8327, N8310, N8100, N4672, N5606);
nor NOR3 (N8328, N8327, N7279, N7825);
buf BUF1 (N8329, N8319);
or OR3 (N8330, N8320, N4759, N6327);
nor NOR4 (N8331, N8330, N5685, N8228, N2182);
buf BUF1 (N8332, N8328);
or OR2 (N8333, N8321, N2506);
and AND3 (N8334, N8293, N4197, N358);
buf BUF1 (N8335, N8323);
or OR2 (N8336, N8332, N5481);
buf BUF1 (N8337, N8333);
buf BUF1 (N8338, N8326);
nand NAND2 (N8339, N8329, N996);
or OR4 (N8340, N8338, N3685, N8269, N8178);
and AND2 (N8341, N8324, N5594);
xor XOR2 (N8342, N8325, N2073);
buf BUF1 (N8343, N8337);
not NOT1 (N8344, N8334);
xor XOR2 (N8345, N8336, N5037);
or OR2 (N8346, N8344, N4834);
and AND2 (N8347, N8322, N3792);
and AND4 (N8348, N8340, N6721, N8228, N3459);
nor NOR2 (N8349, N8335, N3320);
nor NOR3 (N8350, N8342, N8217, N32);
or OR2 (N8351, N8339, N4020);
nand NAND3 (N8352, N8343, N5455, N2936);
nand NAND2 (N8353, N8331, N3933);
or OR3 (N8354, N8353, N5125, N1921);
and AND2 (N8355, N8345, N6010);
not NOT1 (N8356, N8350);
and AND2 (N8357, N8348, N7661);
nor NOR3 (N8358, N8346, N1308, N4622);
xor XOR2 (N8359, N8341, N6712);
nand NAND2 (N8360, N8359, N939);
or OR2 (N8361, N8356, N1394);
xor XOR2 (N8362, N8351, N2479);
and AND2 (N8363, N8358, N4335);
nor NOR4 (N8364, N8347, N2724, N1611, N5798);
or OR4 (N8365, N8361, N6137, N8048, N5122);
and AND4 (N8366, N8349, N3272, N2216, N7073);
not NOT1 (N8367, N8357);
nor NOR2 (N8368, N8355, N2098);
xor XOR2 (N8369, N8366, N5770);
buf BUF1 (N8370, N8368);
xor XOR2 (N8371, N8365, N6443);
not NOT1 (N8372, N8364);
buf BUF1 (N8373, N8362);
nand NAND2 (N8374, N8367, N5512);
or OR2 (N8375, N8372, N1484);
xor XOR2 (N8376, N8373, N7472);
and AND2 (N8377, N8363, N1660);
not NOT1 (N8378, N8354);
or OR4 (N8379, N8376, N5192, N1315, N6304);
buf BUF1 (N8380, N8371);
nand NAND2 (N8381, N8369, N4135);
buf BUF1 (N8382, N8352);
buf BUF1 (N8383, N8374);
nand NAND4 (N8384, N8383, N4330, N6299, N3440);
nor NOR4 (N8385, N8382, N7867, N4274, N7053);
xor XOR2 (N8386, N8379, N1060);
nor NOR2 (N8387, N8386, N5422);
nand NAND4 (N8388, N8387, N1863, N4966, N4802);
nor NOR3 (N8389, N8378, N4933, N7269);
and AND3 (N8390, N8388, N6892, N8240);
nand NAND4 (N8391, N8381, N2665, N3556, N5295);
or OR3 (N8392, N8360, N3966, N656);
nor NOR3 (N8393, N8375, N2404, N923);
nor NOR3 (N8394, N8390, N2318, N7802);
and AND3 (N8395, N8385, N3820, N2350);
nand NAND2 (N8396, N8377, N636);
or OR2 (N8397, N8393, N6857);
or OR4 (N8398, N8370, N3517, N1121, N3426);
buf BUF1 (N8399, N8394);
or OR3 (N8400, N8391, N1202, N40);
nor NOR4 (N8401, N8399, N2157, N7241, N5003);
not NOT1 (N8402, N8396);
buf BUF1 (N8403, N8398);
buf BUF1 (N8404, N8403);
and AND4 (N8405, N8384, N7230, N5508, N2513);
xor XOR2 (N8406, N8404, N3997);
or OR4 (N8407, N8395, N2795, N2814, N1845);
buf BUF1 (N8408, N8392);
buf BUF1 (N8409, N8408);
nor NOR3 (N8410, N8402, N3452, N591);
or OR3 (N8411, N8389, N1414, N3703);
and AND2 (N8412, N8409, N1764);
not NOT1 (N8413, N8410);
and AND4 (N8414, N8401, N679, N1191, N5237);
xor XOR2 (N8415, N8380, N5768);
xor XOR2 (N8416, N8397, N5923);
and AND4 (N8417, N8407, N5729, N6722, N5969);
not NOT1 (N8418, N8416);
nand NAND3 (N8419, N8406, N5770, N4903);
xor XOR2 (N8420, N8419, N1897);
nor NOR3 (N8421, N8420, N5484, N4558);
nor NOR4 (N8422, N8405, N3685, N4302, N7517);
buf BUF1 (N8423, N8400);
nor NOR2 (N8424, N8418, N7545);
nor NOR4 (N8425, N8411, N943, N4351, N4883);
and AND2 (N8426, N8413, N4566);
not NOT1 (N8427, N8424);
or OR4 (N8428, N8415, N2952, N3041, N2475);
or OR2 (N8429, N8426, N3190);
nor NOR3 (N8430, N8429, N962, N8191);
buf BUF1 (N8431, N8423);
nor NOR4 (N8432, N8412, N446, N1165, N1037);
and AND3 (N8433, N8427, N263, N623);
and AND2 (N8434, N8422, N3832);
buf BUF1 (N8435, N8428);
not NOT1 (N8436, N8430);
buf BUF1 (N8437, N8432);
nor NOR2 (N8438, N8435, N5488);
nor NOR2 (N8439, N8421, N2967);
or OR3 (N8440, N8431, N4225, N7154);
not NOT1 (N8441, N8440);
not NOT1 (N8442, N8437);
or OR3 (N8443, N8441, N6486, N5809);
xor XOR2 (N8444, N8414, N5835);
xor XOR2 (N8445, N8425, N7537);
or OR2 (N8446, N8445, N5120);
not NOT1 (N8447, N8446);
not NOT1 (N8448, N8443);
or OR2 (N8449, N8447, N134);
nand NAND3 (N8450, N8417, N5073, N4899);
buf BUF1 (N8451, N8450);
xor XOR2 (N8452, N8438, N3032);
not NOT1 (N8453, N8434);
nor NOR3 (N8454, N8448, N4791, N7733);
or OR4 (N8455, N8436, N2807, N1925, N5944);
buf BUF1 (N8456, N8452);
nand NAND3 (N8457, N8439, N4996, N3264);
and AND2 (N8458, N8457, N8046);
and AND4 (N8459, N8456, N3818, N7274, N907);
buf BUF1 (N8460, N8459);
nor NOR4 (N8461, N8444, N4943, N4146, N8147);
nand NAND2 (N8462, N8460, N2519);
xor XOR2 (N8463, N8455, N1993);
not NOT1 (N8464, N8433);
or OR2 (N8465, N8458, N4142);
and AND3 (N8466, N8463, N7497, N7317);
and AND3 (N8467, N8464, N1739, N3082);
or OR2 (N8468, N8454, N4103);
and AND4 (N8469, N8442, N1014, N2889, N4937);
or OR2 (N8470, N8462, N918);
and AND3 (N8471, N8470, N2937, N832);
nand NAND2 (N8472, N8468, N3911);
or OR3 (N8473, N8453, N7738, N2283);
xor XOR2 (N8474, N8466, N4099);
and AND3 (N8475, N8461, N4466, N4907);
and AND2 (N8476, N8471, N3453);
and AND3 (N8477, N8465, N8458, N2687);
nor NOR2 (N8478, N8473, N2217);
buf BUF1 (N8479, N8476);
buf BUF1 (N8480, N8451);
buf BUF1 (N8481, N8480);
not NOT1 (N8482, N8472);
nor NOR2 (N8483, N8449, N473);
xor XOR2 (N8484, N8481, N531);
xor XOR2 (N8485, N8483, N3572);
not NOT1 (N8486, N8477);
not NOT1 (N8487, N8482);
or OR2 (N8488, N8474, N1925);
not NOT1 (N8489, N8469);
nor NOR3 (N8490, N8485, N6936, N7086);
not NOT1 (N8491, N8488);
buf BUF1 (N8492, N8484);
not NOT1 (N8493, N8467);
nor NOR4 (N8494, N8486, N3925, N7369, N2495);
nand NAND2 (N8495, N8491, N4454);
and AND4 (N8496, N8487, N4813, N2230, N3661);
and AND3 (N8497, N8475, N2837, N5548);
not NOT1 (N8498, N8494);
and AND3 (N8499, N8492, N984, N4110);
xor XOR2 (N8500, N8490, N1472);
nor NOR4 (N8501, N8478, N3138, N2052, N7429);
or OR3 (N8502, N8489, N1751, N3921);
nand NAND2 (N8503, N8500, N1330);
nor NOR4 (N8504, N8502, N8266, N4100, N1272);
not NOT1 (N8505, N8496);
and AND3 (N8506, N8499, N7635, N5134);
and AND2 (N8507, N8493, N294);
nor NOR3 (N8508, N8501, N300, N7392);
nor NOR4 (N8509, N8495, N4381, N6006, N4943);
and AND3 (N8510, N8498, N3375, N5661);
xor XOR2 (N8511, N8506, N2953);
or OR2 (N8512, N8510, N5873);
nor NOR2 (N8513, N8511, N5802);
xor XOR2 (N8514, N8505, N6213);
buf BUF1 (N8515, N8513);
nor NOR4 (N8516, N8503, N8039, N6699, N5591);
or OR4 (N8517, N8512, N2728, N5629, N7255);
nand NAND3 (N8518, N8509, N8237, N7217);
nand NAND2 (N8519, N8479, N246);
and AND2 (N8520, N8515, N7161);
nor NOR2 (N8521, N8504, N1674);
not NOT1 (N8522, N8508);
xor XOR2 (N8523, N8507, N6148);
and AND3 (N8524, N8520, N3969, N4718);
and AND3 (N8525, N8523, N5224, N4589);
nand NAND2 (N8526, N8519, N2694);
nand NAND4 (N8527, N8524, N3356, N3869, N129);
and AND3 (N8528, N8521, N2906, N5367);
nor NOR2 (N8529, N8497, N5101);
not NOT1 (N8530, N8526);
not NOT1 (N8531, N8528);
not NOT1 (N8532, N8530);
buf BUF1 (N8533, N8514);
nand NAND4 (N8534, N8517, N6379, N6527, N3254);
nand NAND4 (N8535, N8525, N1721, N4123, N7619);
buf BUF1 (N8536, N8529);
or OR3 (N8537, N8527, N3501, N4153);
not NOT1 (N8538, N8522);
or OR2 (N8539, N8537, N2019);
xor XOR2 (N8540, N8538, N6976);
and AND2 (N8541, N8539, N1833);
not NOT1 (N8542, N8540);
buf BUF1 (N8543, N8531);
nand NAND4 (N8544, N8533, N2169, N1900, N5767);
buf BUF1 (N8545, N8516);
nand NAND3 (N8546, N8542, N392, N6207);
nand NAND4 (N8547, N8536, N7936, N6981, N2007);
and AND3 (N8548, N8541, N5170, N6692);
buf BUF1 (N8549, N8534);
buf BUF1 (N8550, N8544);
not NOT1 (N8551, N8550);
or OR3 (N8552, N8551, N8237, N6924);
not NOT1 (N8553, N8545);
xor XOR2 (N8554, N8553, N5681);
xor XOR2 (N8555, N8535, N6330);
nand NAND4 (N8556, N8518, N717, N6145, N253);
buf BUF1 (N8557, N8543);
xor XOR2 (N8558, N8549, N3699);
or OR2 (N8559, N8547, N3198);
nor NOR3 (N8560, N8548, N7882, N7246);
or OR2 (N8561, N8554, N8141);
xor XOR2 (N8562, N8555, N6843);
buf BUF1 (N8563, N8558);
nor NOR4 (N8564, N8556, N6437, N7772, N1358);
not NOT1 (N8565, N8552);
xor XOR2 (N8566, N8564, N7069);
nand NAND4 (N8567, N8563, N4240, N5500, N7654);
xor XOR2 (N8568, N8546, N1845);
not NOT1 (N8569, N8532);
buf BUF1 (N8570, N8568);
not NOT1 (N8571, N8557);
buf BUF1 (N8572, N8561);
and AND3 (N8573, N8569, N6015, N6367);
or OR3 (N8574, N8572, N2721, N270);
or OR3 (N8575, N8565, N3137, N4011);
nor NOR4 (N8576, N8562, N6733, N4845, N1084);
or OR2 (N8577, N8560, N5631);
nor NOR3 (N8578, N8570, N3983, N4562);
and AND4 (N8579, N8566, N5459, N8197, N2186);
not NOT1 (N8580, N8573);
and AND2 (N8581, N8575, N7787);
not NOT1 (N8582, N8559);
not NOT1 (N8583, N8571);
buf BUF1 (N8584, N8567);
xor XOR2 (N8585, N8574, N6652);
nand NAND4 (N8586, N8576, N7839, N2154, N6779);
nor NOR2 (N8587, N8581, N4482);
nor NOR4 (N8588, N8582, N6858, N3341, N2165);
nor NOR4 (N8589, N8585, N1853, N230, N5867);
or OR4 (N8590, N8577, N7452, N5359, N6288);
nor NOR3 (N8591, N8579, N8182, N4650);
xor XOR2 (N8592, N8587, N7701);
not NOT1 (N8593, N8588);
and AND2 (N8594, N8589, N4438);
and AND3 (N8595, N8593, N4569, N606);
or OR3 (N8596, N8584, N425, N6326);
buf BUF1 (N8597, N8592);
xor XOR2 (N8598, N8580, N4497);
nand NAND2 (N8599, N8596, N1088);
nor NOR4 (N8600, N8595, N964, N7528, N1695);
xor XOR2 (N8601, N8590, N7581);
not NOT1 (N8602, N8598);
buf BUF1 (N8603, N8597);
not NOT1 (N8604, N8603);
or OR3 (N8605, N8604, N6216, N492);
or OR3 (N8606, N8578, N1440, N194);
and AND2 (N8607, N8606, N8218);
buf BUF1 (N8608, N8601);
not NOT1 (N8609, N8583);
buf BUF1 (N8610, N8609);
and AND4 (N8611, N8608, N7908, N6913, N4915);
nand NAND3 (N8612, N8600, N728, N4841);
buf BUF1 (N8613, N8586);
nor NOR4 (N8614, N8610, N3241, N5997, N4134);
buf BUF1 (N8615, N8612);
xor XOR2 (N8616, N8591, N6310);
xor XOR2 (N8617, N8594, N3626);
or OR4 (N8618, N8615, N252, N7177, N5824);
nor NOR3 (N8619, N8613, N3577, N4125);
xor XOR2 (N8620, N8617, N7946);
nand NAND4 (N8621, N8607, N4130, N1508, N8357);
not NOT1 (N8622, N8616);
and AND3 (N8623, N8605, N2176, N382);
or OR2 (N8624, N8602, N8432);
or OR4 (N8625, N8618, N1462, N2126, N4943);
nor NOR3 (N8626, N8623, N6361, N2929);
not NOT1 (N8627, N8625);
and AND4 (N8628, N8614, N4632, N1190, N6752);
xor XOR2 (N8629, N8624, N3132);
nand NAND2 (N8630, N8629, N6546);
and AND4 (N8631, N8627, N4641, N714, N3667);
xor XOR2 (N8632, N8626, N1296);
nand NAND4 (N8633, N8631, N4576, N8243, N920);
not NOT1 (N8634, N8632);
xor XOR2 (N8635, N8633, N442);
and AND3 (N8636, N8622, N7718, N6165);
or OR4 (N8637, N8599, N2743, N980, N1434);
and AND4 (N8638, N8619, N7074, N346, N356);
not NOT1 (N8639, N8628);
not NOT1 (N8640, N8611);
not NOT1 (N8641, N8630);
buf BUF1 (N8642, N8639);
and AND3 (N8643, N8620, N2353, N423);
and AND3 (N8644, N8642, N1083, N6167);
buf BUF1 (N8645, N8636);
nand NAND2 (N8646, N8641, N8497);
not NOT1 (N8647, N8635);
nand NAND3 (N8648, N8621, N1531, N8285);
xor XOR2 (N8649, N8638, N3626);
not NOT1 (N8650, N8643);
nor NOR2 (N8651, N8649, N7012);
buf BUF1 (N8652, N8648);
xor XOR2 (N8653, N8650, N349);
buf BUF1 (N8654, N8645);
xor XOR2 (N8655, N8647, N3720);
buf BUF1 (N8656, N8653);
or OR4 (N8657, N8646, N3949, N1914, N1875);
xor XOR2 (N8658, N8657, N7612);
not NOT1 (N8659, N8640);
not NOT1 (N8660, N8656);
nand NAND4 (N8661, N8652, N2739, N5767, N2104);
buf BUF1 (N8662, N8661);
xor XOR2 (N8663, N8654, N4029);
not NOT1 (N8664, N8634);
buf BUF1 (N8665, N8660);
not NOT1 (N8666, N8651);
not NOT1 (N8667, N8659);
or OR3 (N8668, N8644, N4501, N7039);
and AND4 (N8669, N8658, N122, N2989, N8300);
and AND2 (N8670, N8668, N5194);
buf BUF1 (N8671, N8667);
xor XOR2 (N8672, N8665, N6701);
or OR3 (N8673, N8671, N4510, N6611);
xor XOR2 (N8674, N8666, N7385);
buf BUF1 (N8675, N8669);
not NOT1 (N8676, N8674);
nor NOR2 (N8677, N8664, N967);
not NOT1 (N8678, N8673);
or OR2 (N8679, N8663, N6451);
or OR2 (N8680, N8670, N240);
or OR4 (N8681, N8680, N5422, N3443, N3971);
not NOT1 (N8682, N8637);
xor XOR2 (N8683, N8677, N5715);
nor NOR4 (N8684, N8672, N6148, N419, N4217);
buf BUF1 (N8685, N8676);
and AND3 (N8686, N8683, N4831, N3824);
nand NAND3 (N8687, N8681, N8006, N3205);
and AND2 (N8688, N8685, N838);
nor NOR2 (N8689, N8682, N2265);
buf BUF1 (N8690, N8662);
nor NOR4 (N8691, N8686, N5279, N4018, N8509);
buf BUF1 (N8692, N8690);
nand NAND4 (N8693, N8692, N8442, N4238, N3443);
xor XOR2 (N8694, N8691, N2157);
and AND2 (N8695, N8689, N6914);
and AND3 (N8696, N8695, N2171, N5172);
nor NOR3 (N8697, N8694, N8472, N5471);
nand NAND2 (N8698, N8687, N2776);
nand NAND4 (N8699, N8675, N1982, N4304, N2464);
nor NOR3 (N8700, N8684, N6714, N1615);
nor NOR2 (N8701, N8688, N4041);
nand NAND4 (N8702, N8679, N2099, N7768, N1559);
xor XOR2 (N8703, N8655, N7352);
or OR3 (N8704, N8702, N5888, N2969);
nand NAND2 (N8705, N8698, N4667);
xor XOR2 (N8706, N8704, N8629);
nor NOR3 (N8707, N8705, N1828, N8395);
buf BUF1 (N8708, N8699);
buf BUF1 (N8709, N8707);
and AND2 (N8710, N8701, N5028);
and AND3 (N8711, N8708, N37, N241);
nor NOR3 (N8712, N8700, N3186, N3758);
and AND4 (N8713, N8697, N3375, N3652, N4706);
not NOT1 (N8714, N8693);
and AND4 (N8715, N8710, N3058, N5970, N3883);
or OR2 (N8716, N8713, N8656);
buf BUF1 (N8717, N8714);
and AND4 (N8718, N8706, N837, N5759, N3332);
not NOT1 (N8719, N8678);
xor XOR2 (N8720, N8717, N6281);
xor XOR2 (N8721, N8703, N5327);
nor NOR3 (N8722, N8712, N3451, N4506);
xor XOR2 (N8723, N8720, N817);
xor XOR2 (N8724, N8722, N7699);
buf BUF1 (N8725, N8696);
nand NAND3 (N8726, N8716, N2613, N4640);
xor XOR2 (N8727, N8718, N7576);
or OR4 (N8728, N8715, N5577, N145, N6333);
and AND4 (N8729, N8711, N7680, N6027, N6312);
or OR3 (N8730, N8719, N5066, N2380);
nor NOR4 (N8731, N8728, N691, N2475, N180);
xor XOR2 (N8732, N8729, N4217);
nand NAND2 (N8733, N8724, N7269);
xor XOR2 (N8734, N8731, N2228);
not NOT1 (N8735, N8732);
or OR4 (N8736, N8723, N3790, N5152, N4742);
nor NOR2 (N8737, N8736, N4438);
buf BUF1 (N8738, N8721);
xor XOR2 (N8739, N8725, N2092);
and AND2 (N8740, N8733, N2226);
or OR2 (N8741, N8730, N2170);
and AND2 (N8742, N8734, N6389);
nand NAND3 (N8743, N8726, N8148, N7956);
buf BUF1 (N8744, N8737);
or OR3 (N8745, N8742, N4186, N1095);
xor XOR2 (N8746, N8740, N2426);
xor XOR2 (N8747, N8741, N6293);
and AND4 (N8748, N8709, N2292, N2865, N4159);
or OR3 (N8749, N8735, N8140, N8058);
nor NOR3 (N8750, N8747, N3419, N5749);
nand NAND4 (N8751, N8748, N8053, N2023, N4701);
xor XOR2 (N8752, N8743, N1666);
buf BUF1 (N8753, N8746);
and AND4 (N8754, N8749, N667, N2452, N6136);
nor NOR2 (N8755, N8727, N8249);
xor XOR2 (N8756, N8745, N2762);
buf BUF1 (N8757, N8753);
and AND3 (N8758, N8755, N133, N3512);
not NOT1 (N8759, N8738);
xor XOR2 (N8760, N8739, N5954);
or OR2 (N8761, N8751, N7915);
buf BUF1 (N8762, N8759);
not NOT1 (N8763, N8756);
nor NOR2 (N8764, N8763, N3101);
nand NAND4 (N8765, N8758, N6254, N7406, N2420);
and AND3 (N8766, N8757, N2933, N3383);
buf BUF1 (N8767, N8754);
not NOT1 (N8768, N8750);
or OR3 (N8769, N8744, N8301, N3977);
nand NAND4 (N8770, N8761, N6247, N7861, N3990);
buf BUF1 (N8771, N8764);
xor XOR2 (N8772, N8760, N5338);
nor NOR4 (N8773, N8752, N573, N1758, N5625);
not NOT1 (N8774, N8769);
nor NOR4 (N8775, N8773, N8506, N7238, N2956);
nor NOR2 (N8776, N8768, N8122);
nor NOR4 (N8777, N8776, N1397, N8454, N2474);
buf BUF1 (N8778, N8772);
and AND4 (N8779, N8775, N970, N4349, N2176);
and AND2 (N8780, N8766, N3123);
not NOT1 (N8781, N8778);
or OR2 (N8782, N8780, N6529);
not NOT1 (N8783, N8765);
not NOT1 (N8784, N8782);
buf BUF1 (N8785, N8784);
not NOT1 (N8786, N8785);
nand NAND2 (N8787, N8781, N327);
or OR3 (N8788, N8787, N7967, N3710);
nand NAND4 (N8789, N8786, N7827, N1511, N318);
nand NAND2 (N8790, N8762, N8137);
or OR2 (N8791, N8777, N3247);
xor XOR2 (N8792, N8790, N3522);
nand NAND4 (N8793, N8771, N5083, N6499, N7835);
nand NAND2 (N8794, N8770, N367);
and AND2 (N8795, N8794, N3819);
not NOT1 (N8796, N8792);
nor NOR4 (N8797, N8791, N7398, N8755, N6684);
buf BUF1 (N8798, N8788);
not NOT1 (N8799, N8783);
nor NOR3 (N8800, N8795, N1065, N6460);
nand NAND2 (N8801, N8796, N4646);
nand NAND3 (N8802, N8800, N8417, N2068);
xor XOR2 (N8803, N8801, N8058);
nor NOR4 (N8804, N8793, N1934, N6592, N7635);
and AND4 (N8805, N8799, N4676, N8054, N6446);
or OR2 (N8806, N8802, N7278);
xor XOR2 (N8807, N8774, N8697);
nand NAND2 (N8808, N8804, N4088);
nor NOR4 (N8809, N8805, N1921, N3785, N3373);
and AND3 (N8810, N8789, N4170, N2384);
xor XOR2 (N8811, N8806, N2784);
xor XOR2 (N8812, N8811, N8011);
nor NOR4 (N8813, N8809, N1145, N1295, N6260);
nor NOR2 (N8814, N8767, N7529);
xor XOR2 (N8815, N8798, N7052);
buf BUF1 (N8816, N8803);
and AND3 (N8817, N8797, N5470, N8434);
xor XOR2 (N8818, N8812, N4281);
buf BUF1 (N8819, N8815);
and AND2 (N8820, N8810, N5790);
nor NOR3 (N8821, N8808, N7707, N3273);
or OR3 (N8822, N8779, N6609, N1575);
and AND2 (N8823, N8822, N3138);
or OR4 (N8824, N8807, N3048, N1525, N8522);
not NOT1 (N8825, N8823);
buf BUF1 (N8826, N8825);
nand NAND2 (N8827, N8819, N4500);
or OR3 (N8828, N8824, N633, N944);
xor XOR2 (N8829, N8827, N5114);
buf BUF1 (N8830, N8829);
or OR2 (N8831, N8830, N7587);
nand NAND3 (N8832, N8820, N5776, N7017);
xor XOR2 (N8833, N8832, N5532);
not NOT1 (N8834, N8826);
or OR3 (N8835, N8828, N8707, N2064);
not NOT1 (N8836, N8813);
or OR4 (N8837, N8821, N3060, N2689, N982);
buf BUF1 (N8838, N8817);
and AND2 (N8839, N8816, N4027);
and AND4 (N8840, N8833, N1706, N8299, N1995);
nand NAND3 (N8841, N8835, N8633, N7964);
xor XOR2 (N8842, N8834, N293);
nand NAND4 (N8843, N8814, N7688, N8138, N8687);
or OR4 (N8844, N8831, N6352, N1082, N8136);
xor XOR2 (N8845, N8836, N1038);
nor NOR4 (N8846, N8840, N6438, N5231, N6553);
and AND2 (N8847, N8844, N5866);
and AND2 (N8848, N8818, N6466);
xor XOR2 (N8849, N8841, N167);
nor NOR3 (N8850, N8837, N2295, N2644);
and AND2 (N8851, N8845, N4162);
and AND2 (N8852, N8850, N696);
not NOT1 (N8853, N8847);
xor XOR2 (N8854, N8843, N1820);
or OR4 (N8855, N8842, N2979, N2455, N7732);
buf BUF1 (N8856, N8846);
buf BUF1 (N8857, N8854);
nand NAND4 (N8858, N8851, N6527, N4977, N1349);
buf BUF1 (N8859, N8839);
nand NAND2 (N8860, N8852, N4975);
not NOT1 (N8861, N8855);
nand NAND4 (N8862, N8859, N7168, N4873, N6688);
xor XOR2 (N8863, N8848, N385);
or OR2 (N8864, N8863, N6259);
buf BUF1 (N8865, N8860);
and AND4 (N8866, N8853, N8523, N2706, N6882);
and AND4 (N8867, N8858, N4255, N5846, N3408);
or OR4 (N8868, N8857, N8709, N7237, N2913);
nand NAND2 (N8869, N8865, N4985);
xor XOR2 (N8870, N8867, N393);
and AND2 (N8871, N8870, N1025);
nor NOR4 (N8872, N8864, N5927, N7869, N4596);
xor XOR2 (N8873, N8862, N2487);
nand NAND2 (N8874, N8869, N6872);
nand NAND3 (N8875, N8838, N820, N2455);
xor XOR2 (N8876, N8873, N8835);
buf BUF1 (N8877, N8872);
and AND2 (N8878, N8849, N6998);
xor XOR2 (N8879, N8868, N5609);
buf BUF1 (N8880, N8866);
and AND2 (N8881, N8875, N4398);
not NOT1 (N8882, N8856);
not NOT1 (N8883, N8881);
nand NAND4 (N8884, N8877, N5368, N2392, N3094);
nand NAND4 (N8885, N8884, N385, N718, N3349);
nor NOR4 (N8886, N8880, N1475, N6843, N581);
nor NOR3 (N8887, N8883, N4772, N6474);
buf BUF1 (N8888, N8887);
not NOT1 (N8889, N8882);
nand NAND3 (N8890, N8885, N7283, N1814);
or OR3 (N8891, N8861, N4071, N6072);
nor NOR4 (N8892, N8891, N2862, N1912, N1417);
nor NOR4 (N8893, N8879, N6885, N2785, N3578);
xor XOR2 (N8894, N8893, N6206);
or OR4 (N8895, N8894, N1402, N8256, N1492);
nand NAND4 (N8896, N8890, N2249, N1103, N1208);
nor NOR3 (N8897, N8889, N2192, N2532);
buf BUF1 (N8898, N8892);
nand NAND4 (N8899, N8886, N3532, N6309, N1782);
nand NAND3 (N8900, N8899, N1045, N6652);
or OR3 (N8901, N8871, N1998, N1152);
xor XOR2 (N8902, N8888, N420);
xor XOR2 (N8903, N8878, N2924);
xor XOR2 (N8904, N8895, N3643);
not NOT1 (N8905, N8901);
not NOT1 (N8906, N8874);
nor NOR3 (N8907, N8902, N330, N8515);
buf BUF1 (N8908, N8876);
and AND4 (N8909, N8896, N4815, N755, N2989);
or OR2 (N8910, N8904, N3530);
buf BUF1 (N8911, N8909);
and AND3 (N8912, N8903, N8783, N3660);
or OR2 (N8913, N8910, N569);
nand NAND3 (N8914, N8897, N7542, N2502);
not NOT1 (N8915, N8914);
buf BUF1 (N8916, N8907);
or OR2 (N8917, N8900, N4954);
buf BUF1 (N8918, N8906);
or OR2 (N8919, N8918, N7606);
or OR3 (N8920, N8917, N3543, N5528);
buf BUF1 (N8921, N8920);
nand NAND4 (N8922, N8908, N5287, N1775, N2537);
nand NAND2 (N8923, N8898, N5912);
buf BUF1 (N8924, N8921);
xor XOR2 (N8925, N8912, N464);
xor XOR2 (N8926, N8911, N4256);
nor NOR2 (N8927, N8922, N1062);
and AND2 (N8928, N8926, N4433);
xor XOR2 (N8929, N8913, N3388);
xor XOR2 (N8930, N8924, N5861);
not NOT1 (N8931, N8905);
buf BUF1 (N8932, N8919);
and AND2 (N8933, N8923, N1147);
xor XOR2 (N8934, N8916, N127);
not NOT1 (N8935, N8934);
xor XOR2 (N8936, N8927, N3147);
nand NAND2 (N8937, N8936, N4225);
xor XOR2 (N8938, N8937, N203);
buf BUF1 (N8939, N8931);
or OR2 (N8940, N8938, N6566);
nand NAND3 (N8941, N8930, N120, N5577);
nor NOR4 (N8942, N8940, N6278, N7229, N7923);
nand NAND3 (N8943, N8932, N8029, N2585);
not NOT1 (N8944, N8943);
nor NOR3 (N8945, N8942, N7173, N8519);
buf BUF1 (N8946, N8935);
xor XOR2 (N8947, N8929, N1331);
nand NAND4 (N8948, N8947, N1555, N1036, N1068);
or OR4 (N8949, N8933, N16, N5091, N2152);
and AND3 (N8950, N8948, N7570, N6130);
or OR4 (N8951, N8949, N8200, N7174, N7506);
nand NAND4 (N8952, N8946, N7870, N2921, N878);
not NOT1 (N8953, N8925);
buf BUF1 (N8954, N8950);
nor NOR3 (N8955, N8952, N968, N2274);
xor XOR2 (N8956, N8939, N6709);
nor NOR3 (N8957, N8944, N325, N4856);
or OR4 (N8958, N8928, N1037, N8117, N286);
xor XOR2 (N8959, N8915, N6913);
nor NOR3 (N8960, N8953, N7693, N3780);
not NOT1 (N8961, N8960);
not NOT1 (N8962, N8954);
nand NAND3 (N8963, N8961, N6629, N7913);
xor XOR2 (N8964, N8962, N4380);
or OR3 (N8965, N8958, N4892, N1539);
buf BUF1 (N8966, N8945);
and AND3 (N8967, N8956, N8008, N5749);
buf BUF1 (N8968, N8965);
not NOT1 (N8969, N8968);
xor XOR2 (N8970, N8941, N2982);
nor NOR3 (N8971, N8967, N2879, N2935);
not NOT1 (N8972, N8959);
nor NOR3 (N8973, N8969, N7909, N4748);
not NOT1 (N8974, N8972);
and AND2 (N8975, N8963, N3363);
nand NAND4 (N8976, N8971, N723, N260, N8542);
buf BUF1 (N8977, N8973);
nand NAND2 (N8978, N8970, N2906);
buf BUF1 (N8979, N8976);
nor NOR3 (N8980, N8951, N8783, N1812);
nor NOR3 (N8981, N8979, N6040, N8166);
xor XOR2 (N8982, N8977, N906);
and AND4 (N8983, N8957, N3727, N1269, N1013);
not NOT1 (N8984, N8978);
nor NOR3 (N8985, N8980, N8663, N3639);
nor NOR4 (N8986, N8974, N5932, N8947, N1017);
xor XOR2 (N8987, N8982, N3104);
xor XOR2 (N8988, N8986, N6363);
nor NOR4 (N8989, N8984, N6933, N7842, N7619);
nand NAND4 (N8990, N8983, N4340, N2275, N722);
xor XOR2 (N8991, N8990, N4159);
nor NOR4 (N8992, N8981, N3603, N4048, N6784);
not NOT1 (N8993, N8964);
not NOT1 (N8994, N8992);
xor XOR2 (N8995, N8966, N3181);
and AND3 (N8996, N8975, N5020, N4330);
nor NOR2 (N8997, N8955, N5744);
not NOT1 (N8998, N8989);
or OR4 (N8999, N8993, N1710, N8456, N4977);
buf BUF1 (N9000, N8999);
buf BUF1 (N9001, N8995);
nor NOR4 (N9002, N8991, N236, N1652, N576);
not NOT1 (N9003, N9001);
nor NOR3 (N9004, N8994, N2195, N1899);
nor NOR3 (N9005, N8998, N231, N4437);
and AND4 (N9006, N8988, N4219, N1187, N8710);
not NOT1 (N9007, N9004);
not NOT1 (N9008, N8997);
not NOT1 (N9009, N9007);
nand NAND3 (N9010, N9005, N3406, N3298);
or OR2 (N9011, N9000, N2091);
nor NOR2 (N9012, N9002, N506);
xor XOR2 (N9013, N9010, N7706);
nor NOR3 (N9014, N9008, N6085, N8941);
xor XOR2 (N9015, N9006, N4506);
or OR3 (N9016, N9011, N3454, N2617);
buf BUF1 (N9017, N8996);
nand NAND2 (N9018, N9014, N4946);
xor XOR2 (N9019, N9016, N1961);
not NOT1 (N9020, N9015);
xor XOR2 (N9021, N9003, N8672);
and AND2 (N9022, N9019, N733);
buf BUF1 (N9023, N9017);
or OR2 (N9024, N9012, N464);
xor XOR2 (N9025, N8987, N5248);
or OR3 (N9026, N9018, N8066, N1248);
and AND4 (N9027, N9021, N581, N1425, N1889);
xor XOR2 (N9028, N9022, N277);
and AND2 (N9029, N9013, N1497);
nor NOR4 (N9030, N9027, N3139, N1372, N7363);
nor NOR3 (N9031, N9020, N6709, N7772);
and AND3 (N9032, N9031, N2756, N4246);
and AND2 (N9033, N9023, N4136);
nor NOR4 (N9034, N9028, N626, N1920, N6166);
nor NOR3 (N9035, N9030, N2443, N1657);
or OR3 (N9036, N9033, N909, N9007);
and AND3 (N9037, N9026, N764, N3720);
and AND4 (N9038, N9035, N1101, N585, N4162);
or OR4 (N9039, N9009, N3485, N6921, N3720);
xor XOR2 (N9040, N9025, N3702);
xor XOR2 (N9041, N9036, N243);
and AND2 (N9042, N9032, N526);
not NOT1 (N9043, N8985);
not NOT1 (N9044, N9029);
and AND2 (N9045, N9043, N2174);
nor NOR4 (N9046, N9040, N3262, N747, N2984);
or OR3 (N9047, N9042, N3927, N7836);
not NOT1 (N9048, N9041);
not NOT1 (N9049, N9039);
and AND3 (N9050, N9034, N2574, N8305);
not NOT1 (N9051, N9037);
and AND3 (N9052, N9044, N480, N3770);
buf BUF1 (N9053, N9024);
nand NAND3 (N9054, N9049, N2978, N6229);
xor XOR2 (N9055, N9045, N4068);
xor XOR2 (N9056, N9053, N8627);
or OR3 (N9057, N9052, N599, N7640);
nand NAND4 (N9058, N9054, N3343, N1157, N984);
and AND4 (N9059, N9047, N8886, N643, N4736);
nand NAND4 (N9060, N9056, N8953, N3558, N2001);
not NOT1 (N9061, N9048);
and AND3 (N9062, N9061, N3425, N8551);
xor XOR2 (N9063, N9055, N264);
nor NOR4 (N9064, N9046, N4489, N5934, N2626);
buf BUF1 (N9065, N9062);
nand NAND4 (N9066, N9058, N3769, N5867, N4250);
and AND2 (N9067, N9038, N4955);
nand NAND4 (N9068, N9063, N6310, N3346, N8073);
buf BUF1 (N9069, N9065);
not NOT1 (N9070, N9057);
nand NAND4 (N9071, N9067, N3253, N1929, N3659);
nand NAND2 (N9072, N9070, N3848);
nand NAND3 (N9073, N9060, N8336, N4942);
nor NOR2 (N9074, N9050, N1797);
and AND2 (N9075, N9059, N2721);
not NOT1 (N9076, N9075);
xor XOR2 (N9077, N9066, N6289);
not NOT1 (N9078, N9074);
not NOT1 (N9079, N9076);
buf BUF1 (N9080, N9064);
and AND2 (N9081, N9071, N4957);
and AND3 (N9082, N9073, N6882, N3794);
buf BUF1 (N9083, N9079);
buf BUF1 (N9084, N9081);
or OR3 (N9085, N9072, N4333, N6126);
nand NAND2 (N9086, N9085, N2892);
not NOT1 (N9087, N9069);
nand NAND2 (N9088, N9082, N770);
xor XOR2 (N9089, N9088, N176);
buf BUF1 (N9090, N9084);
nor NOR4 (N9091, N9051, N1376, N6431, N4531);
xor XOR2 (N9092, N9086, N5315);
nor NOR2 (N9093, N9083, N7809);
nand NAND4 (N9094, N9078, N4797, N5484, N6671);
nand NAND3 (N9095, N9094, N7827, N3877);
buf BUF1 (N9096, N9090);
and AND2 (N9097, N9092, N5790);
and AND2 (N9098, N9089, N7852);
not NOT1 (N9099, N9097);
and AND4 (N9100, N9087, N6468, N5390, N5354);
nand NAND4 (N9101, N9098, N7222, N1963, N8295);
buf BUF1 (N9102, N9091);
xor XOR2 (N9103, N9099, N2396);
xor XOR2 (N9104, N9096, N8080);
nor NOR3 (N9105, N9100, N536, N8100);
nor NOR3 (N9106, N9095, N8827, N7068);
nor NOR4 (N9107, N9104, N5122, N6686, N896);
buf BUF1 (N9108, N9107);
xor XOR2 (N9109, N9080, N1440);
or OR2 (N9110, N9093, N4057);
xor XOR2 (N9111, N9110, N1255);
nand NAND4 (N9112, N9068, N6198, N2091, N5100);
nand NAND3 (N9113, N9106, N6177, N6931);
and AND4 (N9114, N9108, N7862, N3039, N293);
and AND3 (N9115, N9113, N7327, N3009);
not NOT1 (N9116, N9101);
nor NOR4 (N9117, N9105, N1667, N5180, N3995);
nor NOR4 (N9118, N9109, N1253, N3344, N4007);
xor XOR2 (N9119, N9115, N4425);
xor XOR2 (N9120, N9103, N2476);
nor NOR3 (N9121, N9118, N687, N1415);
or OR3 (N9122, N9077, N1373, N6454);
buf BUF1 (N9123, N9112);
or OR3 (N9124, N9114, N1494, N2059);
nand NAND3 (N9125, N9116, N6451, N7339);
nand NAND4 (N9126, N9120, N7048, N8402, N2763);
buf BUF1 (N9127, N9126);
not NOT1 (N9128, N9127);
xor XOR2 (N9129, N9117, N6886);
nand NAND3 (N9130, N9122, N2019, N7412);
or OR2 (N9131, N9125, N1038);
or OR2 (N9132, N9111, N6845);
nand NAND4 (N9133, N9123, N5231, N3093, N3488);
or OR2 (N9134, N9124, N7370);
buf BUF1 (N9135, N9131);
nand NAND3 (N9136, N9130, N4482, N9058);
buf BUF1 (N9137, N9136);
buf BUF1 (N9138, N9129);
nor NOR4 (N9139, N9119, N3321, N1346, N5706);
nor NOR2 (N9140, N9135, N6878);
nand NAND3 (N9141, N9138, N1110, N3084);
xor XOR2 (N9142, N9132, N4950);
not NOT1 (N9143, N9121);
nor NOR4 (N9144, N9128, N7271, N4283, N2143);
and AND4 (N9145, N9143, N6065, N5611, N4461);
not NOT1 (N9146, N9139);
not NOT1 (N9147, N9137);
nor NOR2 (N9148, N9142, N8771);
not NOT1 (N9149, N9146);
and AND4 (N9150, N9141, N7812, N6600, N2572);
xor XOR2 (N9151, N9102, N5511);
buf BUF1 (N9152, N9133);
nor NOR3 (N9153, N9150, N2220, N3244);
not NOT1 (N9154, N9134);
and AND3 (N9155, N9154, N8906, N505);
and AND4 (N9156, N9145, N5614, N4782, N257);
and AND3 (N9157, N9153, N755, N8190);
or OR4 (N9158, N9156, N5250, N1490, N4831);
and AND4 (N9159, N9155, N8473, N9010, N3288);
nor NOR4 (N9160, N9149, N7978, N1421, N9101);
nor NOR2 (N9161, N9158, N1863);
buf BUF1 (N9162, N9152);
buf BUF1 (N9163, N9160);
buf BUF1 (N9164, N9162);
not NOT1 (N9165, N9161);
and AND3 (N9166, N9159, N4713, N8281);
or OR4 (N9167, N9165, N5923, N5453, N1638);
nor NOR3 (N9168, N9167, N7793, N3723);
nor NOR3 (N9169, N9163, N3961, N5547);
nand NAND4 (N9170, N9140, N7117, N4258, N7063);
xor XOR2 (N9171, N9164, N2920);
buf BUF1 (N9172, N9157);
buf BUF1 (N9173, N9168);
nor NOR2 (N9174, N9173, N4806);
xor XOR2 (N9175, N9147, N7768);
and AND2 (N9176, N9175, N6582);
or OR3 (N9177, N9169, N1011, N4066);
nor NOR2 (N9178, N9171, N3811);
buf BUF1 (N9179, N9148);
nor NOR3 (N9180, N9166, N7896, N5053);
or OR3 (N9181, N9176, N4463, N4671);
xor XOR2 (N9182, N9178, N3258);
nand NAND2 (N9183, N9179, N73);
or OR2 (N9184, N9172, N1057);
nand NAND3 (N9185, N9177, N7422, N4315);
nor NOR4 (N9186, N9181, N2012, N4363, N312);
not NOT1 (N9187, N9151);
nor NOR2 (N9188, N9180, N5167);
buf BUF1 (N9189, N9187);
and AND2 (N9190, N9183, N3171);
and AND4 (N9191, N9144, N621, N4157, N3827);
and AND3 (N9192, N9174, N3735, N1457);
not NOT1 (N9193, N9190);
xor XOR2 (N9194, N9184, N5011);
or OR3 (N9195, N9189, N51, N5932);
not NOT1 (N9196, N9186);
not NOT1 (N9197, N9191);
or OR2 (N9198, N9194, N344);
nor NOR4 (N9199, N9185, N2290, N7708, N2927);
buf BUF1 (N9200, N9170);
nor NOR2 (N9201, N9182, N1302);
buf BUF1 (N9202, N9197);
buf BUF1 (N9203, N9198);
nor NOR3 (N9204, N9203, N7433, N197);
buf BUF1 (N9205, N9202);
and AND3 (N9206, N9204, N9098, N334);
xor XOR2 (N9207, N9201, N5753);
or OR3 (N9208, N9196, N8064, N8606);
not NOT1 (N9209, N9207);
nor NOR4 (N9210, N9199, N3943, N933, N5549);
and AND3 (N9211, N9188, N4508, N2789);
buf BUF1 (N9212, N9209);
xor XOR2 (N9213, N9193, N9096);
not NOT1 (N9214, N9192);
nand NAND3 (N9215, N9211, N5471, N3063);
not NOT1 (N9216, N9210);
and AND2 (N9217, N9200, N4734);
nand NAND2 (N9218, N9206, N2018);
buf BUF1 (N9219, N9213);
nand NAND2 (N9220, N9214, N1421);
buf BUF1 (N9221, N9219);
not NOT1 (N9222, N9220);
or OR2 (N9223, N9221, N6235);
buf BUF1 (N9224, N9208);
and AND4 (N9225, N9216, N1140, N213, N1268);
buf BUF1 (N9226, N9223);
and AND2 (N9227, N9222, N1834);
not NOT1 (N9228, N9227);
xor XOR2 (N9229, N9226, N3392);
buf BUF1 (N9230, N9225);
nor NOR2 (N9231, N9230, N7075);
buf BUF1 (N9232, N9231);
nor NOR2 (N9233, N9212, N2655);
xor XOR2 (N9234, N9232, N6137);
nand NAND3 (N9235, N9233, N6862, N3376);
and AND2 (N9236, N9218, N2032);
nand NAND3 (N9237, N9228, N1325, N5892);
or OR2 (N9238, N9235, N2592);
or OR3 (N9239, N9217, N6926, N8106);
or OR3 (N9240, N9205, N4653, N8910);
xor XOR2 (N9241, N9234, N8559);
nor NOR2 (N9242, N9215, N6621);
nand NAND3 (N9243, N9224, N717, N1260);
or OR4 (N9244, N9240, N7906, N5576, N4551);
nor NOR3 (N9245, N9195, N409, N473);
not NOT1 (N9246, N9245);
buf BUF1 (N9247, N9244);
nand NAND2 (N9248, N9239, N5809);
or OR3 (N9249, N9238, N5160, N7547);
not NOT1 (N9250, N9249);
nor NOR4 (N9251, N9229, N7036, N1490, N1403);
not NOT1 (N9252, N9251);
not NOT1 (N9253, N9252);
or OR2 (N9254, N9237, N1450);
not NOT1 (N9255, N9253);
nor NOR2 (N9256, N9246, N9002);
or OR2 (N9257, N9255, N2426);
nand NAND3 (N9258, N9250, N7093, N1161);
or OR4 (N9259, N9247, N2306, N5414, N6736);
buf BUF1 (N9260, N9258);
or OR3 (N9261, N9248, N3512, N3135);
buf BUF1 (N9262, N9261);
buf BUF1 (N9263, N9257);
buf BUF1 (N9264, N9243);
xor XOR2 (N9265, N9260, N3262);
nor NOR4 (N9266, N9259, N5686, N1683, N6062);
or OR3 (N9267, N9264, N2577, N4950);
nor NOR2 (N9268, N9262, N1729);
xor XOR2 (N9269, N9263, N4093);
nor NOR4 (N9270, N9265, N5445, N2466, N8037);
nor NOR2 (N9271, N9241, N7705);
nor NOR2 (N9272, N9271, N427);
nand NAND2 (N9273, N9270, N8366);
nand NAND2 (N9274, N9267, N8963);
nor NOR2 (N9275, N9256, N6220);
buf BUF1 (N9276, N9266);
not NOT1 (N9277, N9242);
buf BUF1 (N9278, N9269);
nor NOR3 (N9279, N9277, N4993, N3553);
and AND3 (N9280, N9274, N301, N6091);
nor NOR4 (N9281, N9278, N524, N2109, N5559);
nand NAND2 (N9282, N9272, N8424);
nand NAND2 (N9283, N9236, N6054);
not NOT1 (N9284, N9280);
nand NAND3 (N9285, N9268, N7912, N8882);
nand NAND4 (N9286, N9275, N5708, N6851, N4249);
or OR2 (N9287, N9284, N729);
nor NOR3 (N9288, N9281, N262, N8529);
nand NAND2 (N9289, N9254, N3834);
buf BUF1 (N9290, N9282);
or OR4 (N9291, N9279, N7413, N1340, N252);
buf BUF1 (N9292, N9287);
xor XOR2 (N9293, N9292, N5185);
and AND2 (N9294, N9291, N6107);
nor NOR4 (N9295, N9276, N8966, N2063, N8082);
not NOT1 (N9296, N9283);
not NOT1 (N9297, N9273);
or OR4 (N9298, N9290, N5320, N6630, N2687);
and AND4 (N9299, N9294, N595, N407, N6234);
nand NAND4 (N9300, N9296, N8662, N2784, N8813);
nor NOR2 (N9301, N9297, N6919);
or OR3 (N9302, N9301, N4744, N6061);
nand NAND4 (N9303, N9295, N6360, N2355, N7173);
nand NAND2 (N9304, N9289, N1043);
buf BUF1 (N9305, N9300);
not NOT1 (N9306, N9298);
buf BUF1 (N9307, N9305);
buf BUF1 (N9308, N9286);
buf BUF1 (N9309, N9293);
xor XOR2 (N9310, N9302, N1501);
and AND4 (N9311, N9310, N1541, N7088, N544);
xor XOR2 (N9312, N9303, N8034);
xor XOR2 (N9313, N9309, N916);
nor NOR3 (N9314, N9299, N5068, N3976);
and AND2 (N9315, N9313, N2317);
and AND3 (N9316, N9308, N4412, N2447);
nor NOR2 (N9317, N9316, N6977);
or OR2 (N9318, N9312, N2590);
nor NOR4 (N9319, N9318, N7784, N4002, N6959);
nor NOR2 (N9320, N9285, N9103);
and AND2 (N9321, N9317, N7507);
nor NOR4 (N9322, N9311, N7996, N321, N7887);
nand NAND2 (N9323, N9320, N7802);
nand NAND4 (N9324, N9323, N8629, N690, N338);
nand NAND4 (N9325, N9315, N680, N2182, N2743);
buf BUF1 (N9326, N9307);
xor XOR2 (N9327, N9322, N2679);
not NOT1 (N9328, N9326);
and AND2 (N9329, N9321, N8505);
nor NOR4 (N9330, N9314, N8682, N4354, N2688);
not NOT1 (N9331, N9330);
buf BUF1 (N9332, N9306);
buf BUF1 (N9333, N9325);
or OR4 (N9334, N9324, N5651, N3567, N8377);
nor NOR2 (N9335, N9288, N3677);
and AND2 (N9336, N9329, N1412);
not NOT1 (N9337, N9304);
not NOT1 (N9338, N9336);
or OR4 (N9339, N9319, N3379, N2451, N7793);
and AND4 (N9340, N9335, N3756, N2865, N7931);
or OR3 (N9341, N9338, N4000, N2315);
or OR2 (N9342, N9337, N1447);
and AND3 (N9343, N9339, N2369, N795);
nand NAND3 (N9344, N9332, N2400, N8098);
buf BUF1 (N9345, N9328);
and AND3 (N9346, N9342, N740, N4854);
not NOT1 (N9347, N9334);
nand NAND3 (N9348, N9327, N6287, N3879);
and AND3 (N9349, N9344, N4456, N8434);
or OR4 (N9350, N9349, N325, N7509, N4716);
buf BUF1 (N9351, N9340);
and AND4 (N9352, N9345, N7255, N8997, N8294);
not NOT1 (N9353, N9352);
or OR2 (N9354, N9350, N1800);
and AND4 (N9355, N9347, N8472, N1505, N2236);
and AND3 (N9356, N9354, N7575, N9143);
nand NAND2 (N9357, N9346, N403);
not NOT1 (N9358, N9341);
nor NOR3 (N9359, N9333, N890, N4904);
buf BUF1 (N9360, N9356);
and AND3 (N9361, N9358, N4840, N1999);
xor XOR2 (N9362, N9359, N1100);
xor XOR2 (N9363, N9343, N6305);
nor NOR4 (N9364, N9357, N2209, N5870, N3273);
and AND2 (N9365, N9361, N6045);
nand NAND3 (N9366, N9362, N1886, N6721);
nor NOR3 (N9367, N9365, N5095, N7438);
buf BUF1 (N9368, N9351);
xor XOR2 (N9369, N9367, N4588);
buf BUF1 (N9370, N9368);
nand NAND4 (N9371, N9363, N9077, N5498, N3089);
not NOT1 (N9372, N9371);
nand NAND3 (N9373, N9369, N9207, N5314);
nor NOR4 (N9374, N9360, N1003, N4104, N3127);
or OR3 (N9375, N9373, N9315, N471);
buf BUF1 (N9376, N9353);
and AND4 (N9377, N9374, N1927, N820, N7164);
nand NAND3 (N9378, N9377, N5019, N1324);
nor NOR2 (N9379, N9348, N3794);
nor NOR4 (N9380, N9331, N629, N2913, N1905);
nand NAND4 (N9381, N9378, N7507, N2698, N5305);
buf BUF1 (N9382, N9375);
nor NOR3 (N9383, N9380, N8563, N2828);
or OR3 (N9384, N9366, N3879, N3932);
not NOT1 (N9385, N9379);
xor XOR2 (N9386, N9384, N2455);
nor NOR3 (N9387, N9355, N1163, N4601);
and AND4 (N9388, N9385, N5503, N5334, N1538);
and AND4 (N9389, N9376, N1300, N9264, N6517);
and AND4 (N9390, N9389, N4210, N6285, N6205);
nor NOR3 (N9391, N9388, N5059, N1806);
not NOT1 (N9392, N9370);
or OR3 (N9393, N9387, N6674, N9214);
and AND4 (N9394, N9383, N7756, N751, N1942);
xor XOR2 (N9395, N9390, N8299);
nand NAND3 (N9396, N9372, N4675, N386);
nor NOR3 (N9397, N9393, N3525, N3272);
or OR2 (N9398, N9391, N2799);
xor XOR2 (N9399, N9364, N8632);
xor XOR2 (N9400, N9395, N8172);
and AND4 (N9401, N9394, N2687, N8964, N2463);
and AND4 (N9402, N9382, N9192, N798, N200);
nor NOR4 (N9403, N9398, N5176, N110, N335);
nand NAND4 (N9404, N9381, N4177, N6537, N7440);
nand NAND3 (N9405, N9397, N8933, N867);
not NOT1 (N9406, N9404);
xor XOR2 (N9407, N9392, N6656);
not NOT1 (N9408, N9396);
not NOT1 (N9409, N9403);
xor XOR2 (N9410, N9400, N8100);
nand NAND3 (N9411, N9401, N1439, N2291);
and AND4 (N9412, N9399, N5876, N2012, N5508);
or OR4 (N9413, N9407, N4106, N7110, N9211);
or OR2 (N9414, N9408, N1217);
buf BUF1 (N9415, N9386);
not NOT1 (N9416, N9414);
nor NOR2 (N9417, N9402, N783);
buf BUF1 (N9418, N9406);
xor XOR2 (N9419, N9410, N4473);
not NOT1 (N9420, N9405);
buf BUF1 (N9421, N9419);
and AND2 (N9422, N9411, N9034);
nor NOR4 (N9423, N9418, N6268, N8645, N867);
or OR2 (N9424, N9417, N6111);
nor NOR2 (N9425, N9423, N1390);
nor NOR2 (N9426, N9415, N42);
nor NOR2 (N9427, N9409, N659);
nor NOR3 (N9428, N9422, N3508, N5711);
and AND3 (N9429, N9420, N7638, N3809);
nor NOR2 (N9430, N9428, N7924);
or OR3 (N9431, N9424, N1651, N6577);
not NOT1 (N9432, N9426);
and AND3 (N9433, N9427, N7599, N7657);
nand NAND3 (N9434, N9413, N8903, N7026);
nand NAND2 (N9435, N9412, N2898);
nand NAND3 (N9436, N9433, N7075, N8939);
buf BUF1 (N9437, N9425);
buf BUF1 (N9438, N9416);
nand NAND4 (N9439, N9437, N5660, N5284, N7239);
nand NAND3 (N9440, N9434, N1708, N3356);
buf BUF1 (N9441, N9436);
and AND3 (N9442, N9421, N849, N6079);
xor XOR2 (N9443, N9439, N5408);
and AND2 (N9444, N9429, N5336);
xor XOR2 (N9445, N9444, N1061);
and AND2 (N9446, N9443, N7751);
nor NOR2 (N9447, N9435, N3591);
nor NOR3 (N9448, N9441, N7547, N3563);
or OR2 (N9449, N9432, N2117);
nand NAND2 (N9450, N9442, N6746);
or OR3 (N9451, N9447, N3460, N8796);
or OR2 (N9452, N9431, N7023);
xor XOR2 (N9453, N9452, N1799);
buf BUF1 (N9454, N9446);
and AND2 (N9455, N9430, N7569);
nor NOR4 (N9456, N9448, N7096, N2093, N3003);
and AND4 (N9457, N9445, N128, N7137, N2503);
nand NAND2 (N9458, N9457, N87);
xor XOR2 (N9459, N9455, N8038);
not NOT1 (N9460, N9458);
and AND3 (N9461, N9453, N7988, N8422);
or OR4 (N9462, N9451, N8915, N8492, N1910);
nand NAND3 (N9463, N9454, N7771, N2119);
and AND4 (N9464, N9463, N4524, N5148, N2702);
xor XOR2 (N9465, N9438, N6794);
and AND3 (N9466, N9450, N4869, N3491);
nand NAND4 (N9467, N9461, N113, N9254, N4999);
buf BUF1 (N9468, N9456);
nor NOR4 (N9469, N9465, N6689, N887, N6838);
and AND3 (N9470, N9469, N6130, N993);
nor NOR3 (N9471, N9440, N2212, N6391);
nor NOR3 (N9472, N9467, N3894, N5932);
xor XOR2 (N9473, N9460, N4999);
xor XOR2 (N9474, N9471, N9284);
xor XOR2 (N9475, N9466, N5841);
nor NOR4 (N9476, N9449, N8301, N5290, N3976);
buf BUF1 (N9477, N9474);
xor XOR2 (N9478, N9464, N8835);
not NOT1 (N9479, N9462);
xor XOR2 (N9480, N9470, N2679);
and AND4 (N9481, N9475, N5829, N5824, N2383);
xor XOR2 (N9482, N9481, N6709);
and AND2 (N9483, N9479, N2749);
xor XOR2 (N9484, N9468, N2669);
not NOT1 (N9485, N9477);
nor NOR2 (N9486, N9484, N200);
xor XOR2 (N9487, N9478, N2081);
buf BUF1 (N9488, N9482);
not NOT1 (N9489, N9473);
or OR3 (N9490, N9486, N1980, N8528);
not NOT1 (N9491, N9485);
nor NOR4 (N9492, N9483, N1668, N30, N7503);
nor NOR4 (N9493, N9488, N1509, N2821, N1065);
and AND3 (N9494, N9491, N2503, N2228);
nand NAND3 (N9495, N9459, N2594, N2287);
or OR4 (N9496, N9487, N3411, N8389, N8506);
nand NAND2 (N9497, N9496, N1856);
nor NOR3 (N9498, N9490, N2624, N5770);
xor XOR2 (N9499, N9495, N9303);
xor XOR2 (N9500, N9493, N3317);
and AND2 (N9501, N9498, N3497);
buf BUF1 (N9502, N9500);
or OR2 (N9503, N9501, N1227);
not NOT1 (N9504, N9489);
nand NAND4 (N9505, N9503, N2673, N4469, N2466);
nand NAND3 (N9506, N9494, N3613, N3803);
not NOT1 (N9507, N9472);
and AND4 (N9508, N9499, N5590, N8297, N8179);
or OR3 (N9509, N9492, N827, N3555);
nor NOR2 (N9510, N9504, N4377);
and AND4 (N9511, N9506, N4886, N7039, N8117);
xor XOR2 (N9512, N9480, N6155);
nor NOR4 (N9513, N9476, N8316, N3627, N6685);
nand NAND2 (N9514, N9511, N6737);
or OR3 (N9515, N9497, N9500, N5397);
buf BUF1 (N9516, N9515);
xor XOR2 (N9517, N9510, N1917);
and AND2 (N9518, N9516, N2590);
nor NOR2 (N9519, N9513, N2514);
buf BUF1 (N9520, N9512);
or OR3 (N9521, N9517, N4512, N7752);
nand NAND2 (N9522, N9521, N6349);
xor XOR2 (N9523, N9522, N4747);
not NOT1 (N9524, N9518);
not NOT1 (N9525, N9507);
nor NOR3 (N9526, N9505, N5109, N7464);
buf BUF1 (N9527, N9519);
not NOT1 (N9528, N9527);
or OR4 (N9529, N9526, N6690, N8720, N6294);
nand NAND3 (N9530, N9529, N6148, N9465);
and AND3 (N9531, N9509, N6638, N9207);
nand NAND2 (N9532, N9528, N1831);
not NOT1 (N9533, N9525);
nor NOR2 (N9534, N9502, N6790);
xor XOR2 (N9535, N9534, N4403);
xor XOR2 (N9536, N9524, N9085);
buf BUF1 (N9537, N9532);
nand NAND4 (N9538, N9530, N1325, N2273, N7382);
nand NAND2 (N9539, N9535, N5005);
or OR2 (N9540, N9539, N5195);
nand NAND2 (N9541, N9520, N895);
nor NOR2 (N9542, N9508, N2437);
and AND4 (N9543, N9538, N1161, N8986, N6360);
buf BUF1 (N9544, N9542);
or OR4 (N9545, N9543, N1840, N567, N4199);
nor NOR3 (N9546, N9544, N5033, N3982);
nand NAND4 (N9547, N9537, N5709, N7840, N398);
nand NAND2 (N9548, N9523, N5632);
or OR3 (N9549, N9546, N2256, N2323);
buf BUF1 (N9550, N9536);
and AND4 (N9551, N9514, N8698, N2249, N4807);
or OR3 (N9552, N9550, N8886, N5366);
buf BUF1 (N9553, N9531);
and AND2 (N9554, N9549, N3542);
nor NOR2 (N9555, N9554, N4544);
xor XOR2 (N9556, N9555, N3058);
nor NOR4 (N9557, N9533, N573, N6404, N2281);
or OR3 (N9558, N9548, N1981, N1476);
nand NAND3 (N9559, N9545, N4256, N6895);
xor XOR2 (N9560, N9559, N9281);
or OR4 (N9561, N9541, N8475, N3460, N1067);
and AND4 (N9562, N9561, N5732, N4150, N2911);
nand NAND2 (N9563, N9556, N7266);
not NOT1 (N9564, N9558);
and AND2 (N9565, N9564, N1836);
nor NOR2 (N9566, N9565, N3337);
and AND3 (N9567, N9566, N5755, N8951);
or OR3 (N9568, N9562, N267, N2767);
or OR4 (N9569, N9540, N5169, N3672, N4514);
nand NAND4 (N9570, N9567, N3432, N1734, N7103);
and AND3 (N9571, N9569, N2572, N4731);
nor NOR3 (N9572, N9568, N8533, N4785);
not NOT1 (N9573, N9551);
xor XOR2 (N9574, N9570, N1660);
buf BUF1 (N9575, N9552);
buf BUF1 (N9576, N9557);
xor XOR2 (N9577, N9573, N2807);
and AND3 (N9578, N9576, N6866, N1629);
not NOT1 (N9579, N9577);
and AND4 (N9580, N9579, N175, N8962, N7500);
nor NOR4 (N9581, N9574, N6299, N8869, N1972);
nand NAND4 (N9582, N9578, N4005, N7655, N227);
not NOT1 (N9583, N9582);
not NOT1 (N9584, N9572);
nor NOR3 (N9585, N9584, N7190, N1136);
or OR2 (N9586, N9553, N7212);
nor NOR2 (N9587, N9581, N2412);
xor XOR2 (N9588, N9547, N5883);
and AND3 (N9589, N9563, N1261, N1395);
not NOT1 (N9590, N9588);
or OR2 (N9591, N9571, N8310);
and AND3 (N9592, N9587, N3174, N2099);
buf BUF1 (N9593, N9575);
not NOT1 (N9594, N9560);
nor NOR2 (N9595, N9593, N9202);
buf BUF1 (N9596, N9594);
buf BUF1 (N9597, N9592);
buf BUF1 (N9598, N9583);
not NOT1 (N9599, N9595);
nor NOR4 (N9600, N9597, N5181, N9596, N9075);
nor NOR4 (N9601, N5962, N1745, N8005, N5953);
and AND4 (N9602, N9601, N3710, N9294, N1787);
nor NOR3 (N9603, N9591, N5712, N1960);
not NOT1 (N9604, N9585);
nand NAND2 (N9605, N9589, N4541);
not NOT1 (N9606, N9590);
nand NAND4 (N9607, N9603, N6470, N3836, N6217);
not NOT1 (N9608, N9580);
buf BUF1 (N9609, N9600);
and AND3 (N9610, N9606, N9519, N8576);
or OR4 (N9611, N9607, N7696, N7356, N2883);
or OR4 (N9612, N9586, N8327, N6093, N1140);
buf BUF1 (N9613, N9612);
nand NAND4 (N9614, N9613, N8902, N1760, N2992);
nor NOR3 (N9615, N9599, N4908, N6365);
xor XOR2 (N9616, N9605, N1264);
buf BUF1 (N9617, N9608);
nor NOR3 (N9618, N9602, N816, N3765);
xor XOR2 (N9619, N9617, N5850);
not NOT1 (N9620, N9610);
and AND4 (N9621, N9615, N3233, N487, N9126);
xor XOR2 (N9622, N9604, N6605);
or OR2 (N9623, N9616, N1420);
buf BUF1 (N9624, N9620);
not NOT1 (N9625, N9609);
buf BUF1 (N9626, N9625);
or OR4 (N9627, N9621, N6167, N1182, N7951);
or OR4 (N9628, N9622, N1322, N4370, N6669);
not NOT1 (N9629, N9611);
nand NAND4 (N9630, N9628, N1020, N8512, N5015);
nand NAND3 (N9631, N9598, N5738, N7012);
or OR2 (N9632, N9626, N2214);
nand NAND4 (N9633, N9632, N8062, N3106, N6546);
nand NAND4 (N9634, N9618, N444, N4325, N5335);
and AND3 (N9635, N9627, N4129, N4233);
or OR4 (N9636, N9630, N2537, N7380, N7791);
or OR4 (N9637, N9633, N7924, N4233, N7495);
or OR4 (N9638, N9624, N7251, N5739, N5258);
buf BUF1 (N9639, N9638);
buf BUF1 (N9640, N9639);
nor NOR3 (N9641, N9637, N6520, N2635);
not NOT1 (N9642, N9629);
xor XOR2 (N9643, N9642, N2667);
nand NAND3 (N9644, N9640, N9263, N6195);
buf BUF1 (N9645, N9644);
xor XOR2 (N9646, N9645, N6219);
nor NOR2 (N9647, N9619, N3496);
nor NOR2 (N9648, N9636, N7388);
nor NOR2 (N9649, N9643, N3202);
nor NOR2 (N9650, N9648, N2141);
not NOT1 (N9651, N9623);
or OR3 (N9652, N9631, N158, N6824);
not NOT1 (N9653, N9649);
nor NOR3 (N9654, N9653, N5720, N940);
buf BUF1 (N9655, N9652);
buf BUF1 (N9656, N9646);
xor XOR2 (N9657, N9655, N5427);
nor NOR4 (N9658, N9647, N1438, N4126, N12);
not NOT1 (N9659, N9641);
not NOT1 (N9660, N9656);
nand NAND3 (N9661, N9650, N2345, N553);
and AND3 (N9662, N9635, N697, N4009);
nor NOR2 (N9663, N9658, N6419);
buf BUF1 (N9664, N9663);
and AND2 (N9665, N9662, N8620);
or OR4 (N9666, N9661, N3410, N3169, N3755);
buf BUF1 (N9667, N9666);
or OR4 (N9668, N9614, N1841, N2014, N6907);
nand NAND2 (N9669, N9659, N46);
or OR4 (N9670, N9669, N9231, N8354, N3089);
not NOT1 (N9671, N9654);
or OR2 (N9672, N9665, N4188);
nand NAND4 (N9673, N9634, N2880, N9151, N3572);
xor XOR2 (N9674, N9664, N1885);
nor NOR4 (N9675, N9670, N3414, N7320, N848);
buf BUF1 (N9676, N9674);
nor NOR4 (N9677, N9676, N8562, N8957, N1605);
nand NAND2 (N9678, N9677, N8157);
not NOT1 (N9679, N9673);
not NOT1 (N9680, N9660);
buf BUF1 (N9681, N9680);
or OR2 (N9682, N9675, N95);
nand NAND2 (N9683, N9671, N1505);
and AND3 (N9684, N9651, N538, N984);
buf BUF1 (N9685, N9679);
or OR3 (N9686, N9682, N3732, N8214);
nor NOR4 (N9687, N9672, N3362, N9129, N3037);
buf BUF1 (N9688, N9687);
nor NOR2 (N9689, N9657, N3254);
buf BUF1 (N9690, N9667);
and AND4 (N9691, N9688, N5842, N8943, N6642);
buf BUF1 (N9692, N9684);
not NOT1 (N9693, N9690);
buf BUF1 (N9694, N9683);
nand NAND4 (N9695, N9681, N5154, N2396, N6304);
xor XOR2 (N9696, N9691, N9536);
nand NAND2 (N9697, N9692, N5377);
nor NOR3 (N9698, N9668, N469, N7244);
and AND3 (N9699, N9696, N6471, N4338);
xor XOR2 (N9700, N9678, N3301);
xor XOR2 (N9701, N9695, N7076);
and AND4 (N9702, N9700, N2998, N1555, N4250);
xor XOR2 (N9703, N9694, N1480);
xor XOR2 (N9704, N9697, N7885);
buf BUF1 (N9705, N9699);
nand NAND4 (N9706, N9705, N4033, N3228, N588);
nor NOR4 (N9707, N9686, N6803, N1004, N3934);
or OR2 (N9708, N9701, N3149);
not NOT1 (N9709, N9707);
not NOT1 (N9710, N9708);
not NOT1 (N9711, N9698);
buf BUF1 (N9712, N9704);
xor XOR2 (N9713, N9702, N2647);
buf BUF1 (N9714, N9713);
and AND3 (N9715, N9709, N3699, N1126);
buf BUF1 (N9716, N9711);
xor XOR2 (N9717, N9710, N7193);
nand NAND2 (N9718, N9717, N2032);
and AND4 (N9719, N9715, N4554, N8956, N1549);
nor NOR3 (N9720, N9706, N6243, N8380);
and AND4 (N9721, N9685, N4090, N8960, N2519);
nand NAND3 (N9722, N9720, N4421, N3271);
or OR2 (N9723, N9721, N8741);
nor NOR3 (N9724, N9723, N7087, N9160);
buf BUF1 (N9725, N9703);
buf BUF1 (N9726, N9722);
nor NOR2 (N9727, N9718, N4569);
or OR4 (N9728, N9719, N379, N691, N1721);
buf BUF1 (N9729, N9726);
nor NOR3 (N9730, N9725, N2765, N5516);
or OR3 (N9731, N9727, N7146, N1567);
nand NAND4 (N9732, N9729, N5643, N166, N6477);
nand NAND2 (N9733, N9730, N5805);
and AND4 (N9734, N9693, N5986, N8952, N8690);
or OR4 (N9735, N9714, N3991, N3962, N2133);
nand NAND2 (N9736, N9734, N4148);
nand NAND2 (N9737, N9724, N7909);
nand NAND3 (N9738, N9728, N5719, N6993);
not NOT1 (N9739, N9716);
xor XOR2 (N9740, N9689, N240);
nor NOR2 (N9741, N9739, N9085);
buf BUF1 (N9742, N9741);
and AND4 (N9743, N9731, N6250, N8342, N4215);
nor NOR2 (N9744, N9735, N8351);
nand NAND2 (N9745, N9743, N4354);
not NOT1 (N9746, N9742);
xor XOR2 (N9747, N9740, N8768);
or OR2 (N9748, N9738, N3905);
xor XOR2 (N9749, N9732, N3127);
buf BUF1 (N9750, N9745);
and AND2 (N9751, N9748, N7078);
nand NAND3 (N9752, N9733, N5351, N4522);
buf BUF1 (N9753, N9749);
and AND4 (N9754, N9712, N3771, N434, N4867);
nor NOR3 (N9755, N9736, N5804, N4628);
buf BUF1 (N9756, N9744);
and AND2 (N9757, N9753, N381);
xor XOR2 (N9758, N9751, N6554);
or OR4 (N9759, N9737, N4772, N5247, N5033);
and AND4 (N9760, N9754, N5018, N948, N488);
or OR4 (N9761, N9760, N3072, N7096, N4019);
not NOT1 (N9762, N9752);
not NOT1 (N9763, N9762);
and AND2 (N9764, N9746, N9227);
and AND4 (N9765, N9761, N3523, N556, N7587);
not NOT1 (N9766, N9756);
or OR3 (N9767, N9758, N3543, N4231);
buf BUF1 (N9768, N9755);
or OR3 (N9769, N9767, N2357, N5092);
not NOT1 (N9770, N9769);
nor NOR3 (N9771, N9747, N8203, N2277);
nand NAND3 (N9772, N9759, N3614, N4838);
xor XOR2 (N9773, N9772, N2248);
not NOT1 (N9774, N9771);
not NOT1 (N9775, N9770);
nand NAND3 (N9776, N9766, N1896, N4122);
not NOT1 (N9777, N9765);
or OR2 (N9778, N9750, N5528);
nor NOR2 (N9779, N9777, N7944);
nand NAND2 (N9780, N9768, N1633);
or OR3 (N9781, N9776, N8729, N5177);
nor NOR3 (N9782, N9781, N7231, N5523);
nand NAND4 (N9783, N9778, N9713, N8598, N5742);
and AND3 (N9784, N9780, N6053, N2017);
xor XOR2 (N9785, N9757, N52);
or OR3 (N9786, N9782, N7161, N5300);
or OR4 (N9787, N9786, N574, N980, N4806);
nand NAND3 (N9788, N9784, N7689, N5875);
xor XOR2 (N9789, N9785, N7350);
and AND2 (N9790, N9789, N6464);
not NOT1 (N9791, N9764);
not NOT1 (N9792, N9763);
nand NAND3 (N9793, N9787, N8220, N3227);
and AND2 (N9794, N9788, N2980);
buf BUF1 (N9795, N9792);
or OR4 (N9796, N9774, N4442, N5926, N530);
buf BUF1 (N9797, N9783);
nand NAND3 (N9798, N9794, N8716, N551);
not NOT1 (N9799, N9798);
nand NAND3 (N9800, N9799, N1516, N1247);
nor NOR3 (N9801, N9791, N4919, N8291);
or OR4 (N9802, N9779, N7457, N163, N6553);
xor XOR2 (N9803, N9802, N7953);
not NOT1 (N9804, N9773);
nor NOR2 (N9805, N9800, N1284);
not NOT1 (N9806, N9775);
buf BUF1 (N9807, N9796);
nor NOR4 (N9808, N9805, N7452, N2785, N2671);
xor XOR2 (N9809, N9806, N3617);
and AND2 (N9810, N9801, N4737);
nor NOR2 (N9811, N9808, N9265);
buf BUF1 (N9812, N9793);
nor NOR2 (N9813, N9807, N8701);
or OR3 (N9814, N9810, N8009, N2737);
not NOT1 (N9815, N9811);
or OR4 (N9816, N9790, N1958, N5414, N7453);
nand NAND3 (N9817, N9814, N6458, N826);
nand NAND4 (N9818, N9809, N8997, N5132, N2344);
nand NAND4 (N9819, N9803, N984, N7149, N186);
or OR2 (N9820, N9817, N9664);
xor XOR2 (N9821, N9816, N2627);
xor XOR2 (N9822, N9795, N7264);
xor XOR2 (N9823, N9812, N7413);
xor XOR2 (N9824, N9813, N9440);
nor NOR2 (N9825, N9820, N3458);
and AND4 (N9826, N9821, N8892, N857, N4769);
buf BUF1 (N9827, N9797);
buf BUF1 (N9828, N9827);
buf BUF1 (N9829, N9828);
nor NOR4 (N9830, N9825, N5392, N2891, N9073);
and AND2 (N9831, N9819, N4944);
and AND2 (N9832, N9815, N5202);
and AND2 (N9833, N9832, N8383);
buf BUF1 (N9834, N9823);
not NOT1 (N9835, N9834);
xor XOR2 (N9836, N9833, N1997);
nand NAND4 (N9837, N9818, N1058, N6064, N8039);
xor XOR2 (N9838, N9836, N875);
buf BUF1 (N9839, N9824);
xor XOR2 (N9840, N9838, N5828);
xor XOR2 (N9841, N9822, N3950);
not NOT1 (N9842, N9830);
nand NAND4 (N9843, N9837, N1112, N2987, N5793);
not NOT1 (N9844, N9826);
not NOT1 (N9845, N9842);
nand NAND4 (N9846, N9835, N4777, N1258, N2184);
and AND2 (N9847, N9840, N3854);
xor XOR2 (N9848, N9845, N9462);
and AND3 (N9849, N9829, N4310, N462);
nor NOR4 (N9850, N9849, N7900, N5061, N8454);
not NOT1 (N9851, N9844);
xor XOR2 (N9852, N9846, N5471);
and AND4 (N9853, N9847, N3612, N7009, N3898);
buf BUF1 (N9854, N9850);
xor XOR2 (N9855, N9804, N6757);
not NOT1 (N9856, N9841);
xor XOR2 (N9857, N9854, N8381);
xor XOR2 (N9858, N9852, N7835);
nand NAND3 (N9859, N9843, N9681, N7399);
not NOT1 (N9860, N9858);
buf BUF1 (N9861, N9857);
nor NOR4 (N9862, N9859, N5171, N7263, N5586);
xor XOR2 (N9863, N9860, N4178);
or OR2 (N9864, N9851, N8134);
xor XOR2 (N9865, N9863, N292);
buf BUF1 (N9866, N9864);
nor NOR3 (N9867, N9856, N7136, N6198);
buf BUF1 (N9868, N9861);
buf BUF1 (N9869, N9855);
nand NAND3 (N9870, N9866, N1533, N2560);
not NOT1 (N9871, N9853);
nand NAND4 (N9872, N9865, N4609, N9369, N1327);
nor NOR2 (N9873, N9862, N9279);
or OR3 (N9874, N9867, N5660, N8718);
xor XOR2 (N9875, N9871, N864);
nor NOR3 (N9876, N9870, N202, N7017);
and AND3 (N9877, N9872, N7555, N328);
not NOT1 (N9878, N9876);
buf BUF1 (N9879, N9868);
and AND4 (N9880, N9874, N6738, N9779, N1400);
buf BUF1 (N9881, N9877);
buf BUF1 (N9882, N9848);
not NOT1 (N9883, N9873);
not NOT1 (N9884, N9869);
nor NOR3 (N9885, N9881, N229, N7912);
nand NAND3 (N9886, N9878, N8683, N5652);
or OR2 (N9887, N9839, N5417);
buf BUF1 (N9888, N9880);
buf BUF1 (N9889, N9887);
not NOT1 (N9890, N9888);
or OR3 (N9891, N9875, N8533, N350);
xor XOR2 (N9892, N9879, N5581);
or OR3 (N9893, N9882, N2720, N2279);
nand NAND4 (N9894, N9884, N1956, N3262, N5103);
nor NOR2 (N9895, N9886, N3824);
and AND3 (N9896, N9885, N6862, N8955);
not NOT1 (N9897, N9892);
and AND4 (N9898, N9891, N3639, N8549, N5455);
nor NOR4 (N9899, N9890, N5279, N9038, N4940);
or OR4 (N9900, N9894, N7604, N1173, N787);
nand NAND2 (N9901, N9883, N4563);
or OR2 (N9902, N9831, N9113);
nor NOR3 (N9903, N9896, N2701, N5793);
or OR3 (N9904, N9902, N4883, N1619);
buf BUF1 (N9905, N9897);
nand NAND4 (N9906, N9905, N3148, N9108, N2497);
xor XOR2 (N9907, N9898, N3414);
and AND2 (N9908, N9901, N6985);
not NOT1 (N9909, N9907);
or OR2 (N9910, N9889, N1743);
not NOT1 (N9911, N9908);
nor NOR2 (N9912, N9893, N6623);
or OR3 (N9913, N9900, N1851, N9052);
nand NAND3 (N9914, N9912, N1742, N4321);
nand NAND2 (N9915, N9914, N9354);
buf BUF1 (N9916, N9913);
nor NOR3 (N9917, N9909, N7382, N2168);
buf BUF1 (N9918, N9904);
nand NAND2 (N9919, N9915, N1047);
nand NAND4 (N9920, N9911, N7619, N3752, N4944);
or OR4 (N9921, N9895, N7672, N1523, N2655);
nand NAND4 (N9922, N9918, N4981, N3418, N4270);
not NOT1 (N9923, N9899);
and AND3 (N9924, N9916, N7536, N3060);
nor NOR3 (N9925, N9920, N6579, N5647);
buf BUF1 (N9926, N9924);
and AND4 (N9927, N9903, N954, N5570, N8617);
not NOT1 (N9928, N9926);
nor NOR2 (N9929, N9928, N1380);
or OR3 (N9930, N9919, N3507, N6722);
nand NAND2 (N9931, N9910, N8760);
xor XOR2 (N9932, N9929, N7532);
xor XOR2 (N9933, N9932, N4297);
nor NOR4 (N9934, N9930, N183, N5682, N7851);
not NOT1 (N9935, N9933);
xor XOR2 (N9936, N9922, N8076);
xor XOR2 (N9937, N9935, N6197);
and AND4 (N9938, N9917, N8156, N8126, N8788);
nand NAND4 (N9939, N9936, N55, N9705, N3419);
and AND2 (N9940, N9906, N5568);
xor XOR2 (N9941, N9939, N4765);
buf BUF1 (N9942, N9923);
nor NOR3 (N9943, N9940, N2845, N6531);
and AND2 (N9944, N9943, N3438);
or OR2 (N9945, N9937, N4734);
nor NOR4 (N9946, N9944, N8994, N4338, N1985);
nor NOR4 (N9947, N9925, N8374, N7945, N2096);
xor XOR2 (N9948, N9921, N2078);
or OR2 (N9949, N9938, N2394);
nor NOR4 (N9950, N9945, N2356, N6476, N1545);
buf BUF1 (N9951, N9931);
nor NOR3 (N9952, N9949, N8520, N8162);
nand NAND4 (N9953, N9948, N2348, N8238, N5306);
and AND4 (N9954, N9946, N982, N7428, N4476);
nand NAND4 (N9955, N9950, N8728, N9488, N8141);
not NOT1 (N9956, N9955);
and AND2 (N9957, N9942, N5344);
nand NAND3 (N9958, N9941, N5828, N9099);
xor XOR2 (N9959, N9927, N3347);
or OR3 (N9960, N9954, N2350, N511);
or OR3 (N9961, N9952, N2902, N2488);
xor XOR2 (N9962, N9953, N9237);
not NOT1 (N9963, N9958);
buf BUF1 (N9964, N9960);
xor XOR2 (N9965, N9959, N5575);
and AND3 (N9966, N9934, N2030, N186);
and AND2 (N9967, N9966, N649);
or OR4 (N9968, N9965, N3901, N3886, N222);
nand NAND2 (N9969, N9967, N4380);
or OR4 (N9970, N9964, N6700, N3015, N9756);
nor NOR3 (N9971, N9961, N9097, N8991);
not NOT1 (N9972, N9968);
or OR2 (N9973, N9972, N8785);
or OR4 (N9974, N9973, N4815, N9199, N4565);
not NOT1 (N9975, N9971);
nand NAND2 (N9976, N9963, N748);
nor NOR4 (N9977, N9975, N1815, N8896, N2065);
buf BUF1 (N9978, N9956);
buf BUF1 (N9979, N9951);
buf BUF1 (N9980, N9977);
xor XOR2 (N9981, N9969, N4486);
xor XOR2 (N9982, N9957, N6055);
not NOT1 (N9983, N9981);
or OR3 (N9984, N9947, N2918, N6269);
not NOT1 (N9985, N9970);
nand NAND4 (N9986, N9984, N1236, N9259, N7501);
buf BUF1 (N9987, N9962);
xor XOR2 (N9988, N9983, N7174);
nand NAND4 (N9989, N9986, N6008, N7707, N9873);
nand NAND3 (N9990, N9976, N6274, N8082);
buf BUF1 (N9991, N9989);
and AND2 (N9992, N9987, N8491);
nor NOR3 (N9993, N9979, N4970, N7452);
not NOT1 (N9994, N9991);
nor NOR4 (N9995, N9980, N7319, N9553, N1160);
nand NAND4 (N9996, N9974, N2467, N7043, N5808);
not NOT1 (N9997, N9996);
nand NAND4 (N9998, N9978, N8194, N4172, N9854);
nor NOR2 (N9999, N9998, N1186);
nand NAND2 (N10000, N9994, N444);
xor XOR2 (N10001, N9992, N3695);
nor NOR3 (N10002, N9999, N7980, N2876);
nand NAND3 (N10003, N10001, N5239, N4821);
buf BUF1 (N10004, N9995);
not NOT1 (N10005, N9997);
nor NOR2 (N10006, N9982, N3485);
and AND3 (N10007, N10000, N3874, N1322);
or OR2 (N10008, N10002, N6308);
not NOT1 (N10009, N10006);
nor NOR3 (N10010, N9988, N3524, N8380);
xor XOR2 (N10011, N10007, N8592);
nor NOR4 (N10012, N9993, N4948, N9936, N7329);
xor XOR2 (N10013, N9990, N6622);
buf BUF1 (N10014, N10013);
nand NAND3 (N10015, N10003, N5068, N8959);
nor NOR4 (N10016, N10009, N2489, N4555, N2713);
nand NAND2 (N10017, N10008, N3465);
not NOT1 (N10018, N10015);
and AND3 (N10019, N10005, N2460, N7823);
and AND2 (N10020, N10014, N4648);
buf BUF1 (N10021, N10011);
or OR2 (N10022, N10019, N7145);
nand NAND2 (N10023, N10017, N2798);
nand NAND2 (N10024, N9985, N2497);
nand NAND3 (N10025, N10024, N3163, N9419);
not NOT1 (N10026, N10010);
xor XOR2 (N10027, N10016, N7272);
and AND3 (N10028, N10020, N5421, N4765);
or OR4 (N10029, N10027, N5283, N5326, N6333);
xor XOR2 (N10030, N10026, N5013);
nor NOR2 (N10031, N10018, N923);
xor XOR2 (N10032, N10029, N8037);
or OR2 (N10033, N10028, N3455);
not NOT1 (N10034, N10025);
not NOT1 (N10035, N10022);
xor XOR2 (N10036, N10034, N2489);
or OR3 (N10037, N10035, N4672, N6762);
buf BUF1 (N10038, N10031);
xor XOR2 (N10039, N10030, N7362);
and AND4 (N10040, N10036, N4656, N580, N5875);
or OR2 (N10041, N10039, N4060);
not NOT1 (N10042, N10041);
buf BUF1 (N10043, N10037);
not NOT1 (N10044, N10040);
buf BUF1 (N10045, N10042);
nor NOR4 (N10046, N10012, N2285, N7872, N2467);
nor NOR3 (N10047, N10004, N3993, N503);
not NOT1 (N10048, N10038);
nand NAND2 (N10049, N10033, N4953);
and AND2 (N10050, N10045, N2787);
not NOT1 (N10051, N10049);
nand NAND3 (N10052, N10050, N1134, N779);
and AND2 (N10053, N10052, N7632);
not NOT1 (N10054, N10048);
nor NOR4 (N10055, N10043, N8410, N3019, N676);
buf BUF1 (N10056, N10023);
buf BUF1 (N10057, N10021);
not NOT1 (N10058, N10046);
nor NOR2 (N10059, N10054, N1790);
not NOT1 (N10060, N10056);
buf BUF1 (N10061, N10053);
nor NOR2 (N10062, N10051, N9814);
and AND3 (N10063, N10059, N3002, N4685);
or OR3 (N10064, N10057, N8769, N6853);
and AND2 (N10065, N10063, N5909);
buf BUF1 (N10066, N10062);
and AND4 (N10067, N10064, N5724, N7711, N6221);
nor NOR2 (N10068, N10066, N2379);
nor NOR3 (N10069, N10061, N6574, N5966);
not NOT1 (N10070, N10055);
or OR2 (N10071, N10060, N2019);
xor XOR2 (N10072, N10071, N6100);
or OR4 (N10073, N10032, N1449, N7012, N4681);
xor XOR2 (N10074, N10068, N4832);
xor XOR2 (N10075, N10047, N4328);
nand NAND4 (N10076, N10073, N1664, N5271, N634);
nand NAND2 (N10077, N10044, N6281);
buf BUF1 (N10078, N10072);
nand NAND3 (N10079, N10077, N5685, N5746);
not NOT1 (N10080, N10058);
buf BUF1 (N10081, N10074);
buf BUF1 (N10082, N10076);
buf BUF1 (N10083, N10082);
and AND3 (N10084, N10069, N4401, N1609);
nand NAND3 (N10085, N10083, N1828, N5286);
nor NOR3 (N10086, N10079, N4626, N6014);
xor XOR2 (N10087, N10065, N5158);
nand NAND4 (N10088, N10084, N5893, N3001, N1057);
or OR4 (N10089, N10088, N3130, N4819, N266);
not NOT1 (N10090, N10078);
not NOT1 (N10091, N10080);
buf BUF1 (N10092, N10081);
or OR2 (N10093, N10092, N6300);
or OR4 (N10094, N10070, N6907, N6477, N3685);
and AND4 (N10095, N10086, N3556, N8173, N1391);
nor NOR2 (N10096, N10093, N6690);
not NOT1 (N10097, N10095);
not NOT1 (N10098, N10090);
xor XOR2 (N10099, N10089, N7969);
buf BUF1 (N10100, N10067);
xor XOR2 (N10101, N10097, N2157);
not NOT1 (N10102, N10075);
xor XOR2 (N10103, N10094, N8278);
and AND2 (N10104, N10098, N5085);
xor XOR2 (N10105, N10104, N5056);
buf BUF1 (N10106, N10105);
xor XOR2 (N10107, N10102, N166);
nor NOR2 (N10108, N10100, N3441);
buf BUF1 (N10109, N10101);
not NOT1 (N10110, N10107);
nand NAND2 (N10111, N10109, N7854);
nor NOR4 (N10112, N10103, N5414, N4636, N1948);
nand NAND4 (N10113, N10110, N4358, N4362, N7284);
and AND3 (N10114, N10091, N4766, N8327);
and AND2 (N10115, N10099, N8636);
nand NAND2 (N10116, N10096, N5108);
nand NAND4 (N10117, N10085, N7477, N3212, N5335);
and AND3 (N10118, N10106, N9213, N2411);
nor NOR2 (N10119, N10118, N3220);
not NOT1 (N10120, N10111);
nor NOR4 (N10121, N10115, N966, N1038, N6311);
buf BUF1 (N10122, N10119);
and AND3 (N10123, N10117, N4171, N7637);
and AND3 (N10124, N10120, N6282, N6314);
nor NOR3 (N10125, N10112, N6327, N9193);
nand NAND2 (N10126, N10114, N5717);
or OR2 (N10127, N10121, N3360);
or OR3 (N10128, N10113, N4971, N2154);
and AND4 (N10129, N10108, N5386, N8140, N3536);
or OR4 (N10130, N10124, N1316, N4404, N3716);
not NOT1 (N10131, N10125);
not NOT1 (N10132, N10116);
not NOT1 (N10133, N10130);
buf BUF1 (N10134, N10127);
buf BUF1 (N10135, N10132);
buf BUF1 (N10136, N10087);
xor XOR2 (N10137, N10131, N591);
not NOT1 (N10138, N10129);
or OR2 (N10139, N10134, N8984);
not NOT1 (N10140, N10137);
and AND3 (N10141, N10138, N8720, N4721);
or OR4 (N10142, N10135, N7497, N9429, N9277);
or OR4 (N10143, N10122, N1465, N9013, N2839);
xor XOR2 (N10144, N10133, N5187);
buf BUF1 (N10145, N10123);
nand NAND2 (N10146, N10145, N1846);
buf BUF1 (N10147, N10140);
nand NAND3 (N10148, N10146, N4803, N3960);
nor NOR2 (N10149, N10141, N9863);
xor XOR2 (N10150, N10147, N2259);
buf BUF1 (N10151, N10126);
buf BUF1 (N10152, N10128);
and AND2 (N10153, N10152, N1870);
buf BUF1 (N10154, N10144);
buf BUF1 (N10155, N10154);
nor NOR4 (N10156, N10155, N2769, N8948, N6570);
nor NOR3 (N10157, N10156, N7449, N278);
or OR4 (N10158, N10143, N8309, N8670, N802);
nor NOR4 (N10159, N10149, N8074, N7922, N4923);
nor NOR2 (N10160, N10139, N190);
nand NAND3 (N10161, N10160, N6935, N218);
xor XOR2 (N10162, N10151, N7221);
not NOT1 (N10163, N10157);
nand NAND3 (N10164, N10158, N5487, N9678);
nor NOR2 (N10165, N10148, N2994);
nor NOR2 (N10166, N10153, N3287);
and AND3 (N10167, N10150, N2220, N645);
not NOT1 (N10168, N10166);
buf BUF1 (N10169, N10163);
xor XOR2 (N10170, N10167, N2605);
and AND4 (N10171, N10165, N7823, N8726, N5296);
nor NOR2 (N10172, N10169, N7812);
xor XOR2 (N10173, N10159, N2806);
or OR3 (N10174, N10172, N8128, N1970);
not NOT1 (N10175, N10170);
not NOT1 (N10176, N10136);
xor XOR2 (N10177, N10162, N1354);
xor XOR2 (N10178, N10168, N9530);
xor XOR2 (N10179, N10177, N8061);
nand NAND3 (N10180, N10175, N4715, N2775);
buf BUF1 (N10181, N10176);
xor XOR2 (N10182, N10174, N4139);
or OR3 (N10183, N10142, N6945, N6418);
not NOT1 (N10184, N10182);
and AND2 (N10185, N10179, N7104);
or OR4 (N10186, N10161, N7425, N930, N10117);
and AND3 (N10187, N10180, N8608, N4168);
nor NOR4 (N10188, N10178, N7970, N5551, N6139);
buf BUF1 (N10189, N10184);
buf BUF1 (N10190, N10187);
or OR3 (N10191, N10188, N4341, N6596);
nor NOR4 (N10192, N10190, N2611, N348, N8268);
nand NAND3 (N10193, N10183, N2708, N9474);
xor XOR2 (N10194, N10181, N6117);
nor NOR4 (N10195, N10164, N9410, N22, N3007);
buf BUF1 (N10196, N10193);
and AND2 (N10197, N10194, N3719);
or OR3 (N10198, N10186, N8128, N7814);
not NOT1 (N10199, N10185);
or OR2 (N10200, N10189, N2030);
nand NAND4 (N10201, N10198, N1041, N6398, N1459);
nand NAND3 (N10202, N10197, N5083, N4598);
or OR4 (N10203, N10192, N2975, N5106, N1203);
nor NOR3 (N10204, N10203, N1915, N8539);
buf BUF1 (N10205, N10200);
xor XOR2 (N10206, N10199, N5399);
and AND3 (N10207, N10202, N2364, N1236);
nand NAND2 (N10208, N10171, N9969);
buf BUF1 (N10209, N10201);
nor NOR4 (N10210, N10195, N7987, N536, N8754);
nand NAND4 (N10211, N10206, N6878, N4680, N4228);
and AND3 (N10212, N10173, N2677, N4886);
xor XOR2 (N10213, N10196, N3221);
or OR3 (N10214, N10191, N1135, N8304);
buf BUF1 (N10215, N10213);
nor NOR4 (N10216, N10210, N1820, N2253, N9244);
nor NOR4 (N10217, N10212, N2587, N3054, N8710);
nand NAND2 (N10218, N10204, N4047);
xor XOR2 (N10219, N10215, N4811);
nand NAND3 (N10220, N10207, N3810, N1063);
xor XOR2 (N10221, N10216, N4594);
nor NOR4 (N10222, N10209, N9458, N1741, N1614);
or OR4 (N10223, N10220, N1091, N5028, N6356);
not NOT1 (N10224, N10211);
not NOT1 (N10225, N10217);
nand NAND2 (N10226, N10222, N240);
nand NAND3 (N10227, N10218, N1215, N4647);
and AND3 (N10228, N10208, N9291, N5689);
or OR2 (N10229, N10205, N7409);
xor XOR2 (N10230, N10225, N566);
nor NOR3 (N10231, N10221, N1540, N5788);
or OR4 (N10232, N10229, N7028, N9425, N9853);
buf BUF1 (N10233, N10226);
not NOT1 (N10234, N10230);
nand NAND4 (N10235, N10227, N6566, N6734, N575);
nand NAND4 (N10236, N10214, N8482, N1260, N1803);
and AND3 (N10237, N10224, N5590, N10050);
xor XOR2 (N10238, N10232, N7378);
or OR4 (N10239, N10228, N255, N2517, N4771);
not NOT1 (N10240, N10233);
buf BUF1 (N10241, N10238);
nand NAND2 (N10242, N10240, N2665);
and AND3 (N10243, N10219, N3070, N9265);
and AND4 (N10244, N10241, N879, N2713, N8103);
xor XOR2 (N10245, N10236, N7876);
or OR3 (N10246, N10223, N9813, N7108);
or OR3 (N10247, N10235, N8414, N2337);
and AND4 (N10248, N10246, N6094, N3060, N4171);
not NOT1 (N10249, N10234);
or OR4 (N10250, N10249, N7892, N5017, N4808);
nand NAND4 (N10251, N10239, N6078, N2280, N9624);
or OR3 (N10252, N10244, N7058, N7742);
nor NOR4 (N10253, N10251, N2849, N6883, N3687);
nor NOR3 (N10254, N10248, N1324, N8482);
and AND4 (N10255, N10242, N2367, N7683, N1197);
and AND4 (N10256, N10237, N7068, N4100, N7019);
nand NAND4 (N10257, N10253, N3101, N1095, N5132);
xor XOR2 (N10258, N10243, N5297);
buf BUF1 (N10259, N10256);
not NOT1 (N10260, N10255);
nor NOR4 (N10261, N10259, N7739, N9121, N1065);
or OR2 (N10262, N10260, N7328);
not NOT1 (N10263, N10262);
nand NAND2 (N10264, N10250, N6902);
or OR4 (N10265, N10263, N9975, N7618, N8545);
not NOT1 (N10266, N10264);
xor XOR2 (N10267, N10231, N10117);
or OR3 (N10268, N10258, N5818, N9749);
and AND2 (N10269, N10261, N3147);
and AND2 (N10270, N10252, N2309);
nand NAND4 (N10271, N10265, N1385, N4401, N6840);
not NOT1 (N10272, N10254);
xor XOR2 (N10273, N10271, N7421);
nor NOR3 (N10274, N10269, N6416, N4463);
nand NAND3 (N10275, N10247, N8792, N3390);
and AND4 (N10276, N10245, N6747, N2928, N1675);
nor NOR2 (N10277, N10270, N5363);
nand NAND4 (N10278, N10267, N5423, N7728, N7981);
not NOT1 (N10279, N10268);
xor XOR2 (N10280, N10276, N8310);
nor NOR4 (N10281, N10266, N3266, N6179, N5680);
nor NOR2 (N10282, N10274, N2608);
xor XOR2 (N10283, N10280, N1198);
or OR4 (N10284, N10257, N230, N3839, N4395);
and AND2 (N10285, N10284, N3746);
buf BUF1 (N10286, N10272);
nand NAND4 (N10287, N10283, N5448, N112, N5781);
or OR2 (N10288, N10287, N7237);
or OR2 (N10289, N10285, N2426);
and AND4 (N10290, N10278, N2635, N7273, N1450);
and AND3 (N10291, N10273, N765, N10265);
buf BUF1 (N10292, N10286);
xor XOR2 (N10293, N10282, N7293);
not NOT1 (N10294, N10291);
not NOT1 (N10295, N10292);
and AND2 (N10296, N10290, N6221);
nor NOR2 (N10297, N10275, N5742);
or OR2 (N10298, N10279, N2348);
nor NOR4 (N10299, N10297, N9445, N4604, N3745);
or OR3 (N10300, N10296, N10180, N10098);
or OR3 (N10301, N10299, N9214, N5178);
nand NAND4 (N10302, N10289, N3272, N577, N8926);
nand NAND2 (N10303, N10302, N4561);
xor XOR2 (N10304, N10294, N1627);
or OR3 (N10305, N10300, N7143, N252);
xor XOR2 (N10306, N10298, N6867);
buf BUF1 (N10307, N10277);
buf BUF1 (N10308, N10301);
and AND2 (N10309, N10281, N2386);
not NOT1 (N10310, N10304);
nand NAND4 (N10311, N10307, N6674, N1120, N582);
or OR3 (N10312, N10288, N6402, N8714);
nand NAND2 (N10313, N10305, N1750);
buf BUF1 (N10314, N10309);
or OR4 (N10315, N10293, N7999, N8040, N1364);
xor XOR2 (N10316, N10311, N4777);
not NOT1 (N10317, N10316);
not NOT1 (N10318, N10313);
or OR3 (N10319, N10306, N8638, N9569);
xor XOR2 (N10320, N10318, N6099);
nand NAND2 (N10321, N10303, N699);
nand NAND2 (N10322, N10320, N957);
and AND4 (N10323, N10322, N9399, N9046, N8166);
nand NAND2 (N10324, N10315, N3306);
and AND3 (N10325, N10310, N4780, N856);
or OR3 (N10326, N10314, N2285, N1689);
buf BUF1 (N10327, N10312);
and AND4 (N10328, N10319, N5164, N4715, N2801);
not NOT1 (N10329, N10295);
and AND3 (N10330, N10329, N4562, N2710);
buf BUF1 (N10331, N10328);
xor XOR2 (N10332, N10330, N5464);
nor NOR3 (N10333, N10326, N9218, N429);
buf BUF1 (N10334, N10333);
or OR2 (N10335, N10308, N7813);
buf BUF1 (N10336, N10325);
and AND3 (N10337, N10321, N5142, N5254);
nor NOR3 (N10338, N10332, N2789, N9203);
not NOT1 (N10339, N10324);
xor XOR2 (N10340, N10317, N8238);
and AND4 (N10341, N10338, N9836, N6160, N2601);
nor NOR4 (N10342, N10336, N10003, N8547, N1588);
nand NAND2 (N10343, N10323, N7359);
nor NOR3 (N10344, N10327, N10142, N22);
and AND3 (N10345, N10341, N9798, N5307);
or OR4 (N10346, N10334, N3201, N4128, N8279);
nor NOR4 (N10347, N10345, N9553, N24, N7459);
not NOT1 (N10348, N10340);
nand NAND2 (N10349, N10344, N9016);
buf BUF1 (N10350, N10335);
and AND3 (N10351, N10343, N9332, N9724);
not NOT1 (N10352, N10331);
xor XOR2 (N10353, N10347, N9819);
xor XOR2 (N10354, N10353, N5915);
and AND4 (N10355, N10352, N9417, N1954, N5376);
or OR4 (N10356, N10342, N8444, N4392, N1552);
buf BUF1 (N10357, N10339);
nand NAND4 (N10358, N10348, N6248, N4417, N6616);
buf BUF1 (N10359, N10355);
xor XOR2 (N10360, N10351, N5055);
or OR4 (N10361, N10357, N2574, N3612, N8471);
or OR2 (N10362, N10346, N2847);
buf BUF1 (N10363, N10358);
or OR4 (N10364, N10363, N6657, N8029, N2863);
or OR4 (N10365, N10350, N2328, N2821, N2733);
or OR2 (N10366, N10361, N2126);
or OR2 (N10367, N10366, N5680);
or OR3 (N10368, N10337, N8059, N4368);
and AND4 (N10369, N10359, N4439, N1654, N9623);
nand NAND4 (N10370, N10364, N9132, N304, N9695);
and AND4 (N10371, N10354, N3037, N6349, N2746);
buf BUF1 (N10372, N10360);
nand NAND3 (N10373, N10349, N5410, N4061);
not NOT1 (N10374, N10362);
buf BUF1 (N10375, N10365);
not NOT1 (N10376, N10371);
and AND2 (N10377, N10372, N4371);
buf BUF1 (N10378, N10374);
xor XOR2 (N10379, N10367, N7302);
and AND2 (N10380, N10379, N169);
buf BUF1 (N10381, N10356);
nor NOR4 (N10382, N10373, N734, N7486, N1775);
nor NOR4 (N10383, N10381, N1552, N7303, N7431);
xor XOR2 (N10384, N10382, N10327);
buf BUF1 (N10385, N10376);
nand NAND3 (N10386, N10378, N2726, N1221);
nand NAND2 (N10387, N10369, N4963);
not NOT1 (N10388, N10368);
not NOT1 (N10389, N10375);
and AND2 (N10390, N10389, N210);
or OR4 (N10391, N10377, N6804, N3618, N53);
and AND3 (N10392, N10380, N6496, N9862);
or OR4 (N10393, N10387, N4803, N6323, N3763);
not NOT1 (N10394, N10383);
nor NOR2 (N10395, N10388, N3269);
xor XOR2 (N10396, N10390, N8296);
xor XOR2 (N10397, N10396, N5864);
xor XOR2 (N10398, N10370, N758);
xor XOR2 (N10399, N10391, N10099);
nor NOR3 (N10400, N10397, N9967, N4998);
nor NOR2 (N10401, N10386, N4356);
xor XOR2 (N10402, N10385, N9363);
and AND2 (N10403, N10401, N3281);
or OR4 (N10404, N10399, N8849, N7347, N8398);
buf BUF1 (N10405, N10395);
nand NAND4 (N10406, N10403, N6617, N380, N1731);
nor NOR2 (N10407, N10402, N4565);
nor NOR2 (N10408, N10400, N960);
buf BUF1 (N10409, N10398);
nor NOR2 (N10410, N10404, N1789);
and AND3 (N10411, N10409, N3471, N4943);
and AND4 (N10412, N10392, N10018, N5863, N10025);
not NOT1 (N10413, N10384);
nor NOR2 (N10414, N10413, N2220);
nor NOR2 (N10415, N10410, N7198);
not NOT1 (N10416, N10412);
or OR4 (N10417, N10405, N8821, N7610, N8208);
xor XOR2 (N10418, N10414, N9946);
or OR3 (N10419, N10417, N6941, N7927);
and AND3 (N10420, N10415, N3788, N435);
and AND4 (N10421, N10418, N9259, N4952, N10025);
xor XOR2 (N10422, N10411, N3448);
nor NOR4 (N10423, N10419, N5795, N884, N201);
xor XOR2 (N10424, N10416, N1454);
or OR4 (N10425, N10423, N8176, N3198, N8536);
or OR4 (N10426, N10421, N625, N1215, N1664);
not NOT1 (N10427, N10420);
xor XOR2 (N10428, N10393, N3035);
xor XOR2 (N10429, N10407, N7344);
not NOT1 (N10430, N10429);
or OR4 (N10431, N10406, N6853, N2964, N949);
and AND4 (N10432, N10426, N9017, N1035, N5395);
nor NOR4 (N10433, N10432, N8528, N6905, N8844);
or OR4 (N10434, N10408, N7693, N1406, N2077);
nand NAND4 (N10435, N10427, N10134, N1886, N7653);
and AND2 (N10436, N10435, N6697);
xor XOR2 (N10437, N10434, N5916);
nor NOR2 (N10438, N10437, N7378);
or OR4 (N10439, N10394, N8354, N9446, N3155);
xor XOR2 (N10440, N10433, N9308);
not NOT1 (N10441, N10440);
or OR4 (N10442, N10430, N5689, N3148, N8051);
not NOT1 (N10443, N10439);
not NOT1 (N10444, N10428);
nor NOR2 (N10445, N10425, N4060);
not NOT1 (N10446, N10422);
or OR3 (N10447, N10442, N9287, N1476);
and AND2 (N10448, N10447, N2880);
or OR2 (N10449, N10443, N8216);
nor NOR2 (N10450, N10438, N7825);
and AND3 (N10451, N10424, N4481, N1542);
xor XOR2 (N10452, N10450, N1579);
not NOT1 (N10453, N10446);
buf BUF1 (N10454, N10444);
not NOT1 (N10455, N10441);
nand NAND3 (N10456, N10445, N6539, N5113);
or OR3 (N10457, N10453, N9217, N3900);
not NOT1 (N10458, N10451);
and AND4 (N10459, N10457, N5856, N8428, N9039);
buf BUF1 (N10460, N10449);
nor NOR2 (N10461, N10436, N5306);
nor NOR4 (N10462, N10461, N3592, N8362, N7437);
nor NOR2 (N10463, N10456, N8143);
nor NOR2 (N10464, N10459, N9945);
xor XOR2 (N10465, N10454, N10399);
xor XOR2 (N10466, N10431, N7149);
nor NOR2 (N10467, N10452, N1955);
and AND2 (N10468, N10466, N2804);
nor NOR3 (N10469, N10467, N8319, N2044);
xor XOR2 (N10470, N10460, N1275);
not NOT1 (N10471, N10448);
or OR3 (N10472, N10468, N5323, N2832);
xor XOR2 (N10473, N10472, N9711);
and AND3 (N10474, N10463, N9571, N2534);
xor XOR2 (N10475, N10455, N6207);
nor NOR2 (N10476, N10473, N7028);
nand NAND3 (N10477, N10469, N1210, N4671);
and AND3 (N10478, N10476, N2698, N2832);
xor XOR2 (N10479, N10470, N6416);
buf BUF1 (N10480, N10462);
and AND3 (N10481, N10464, N2620, N399);
not NOT1 (N10482, N10480);
xor XOR2 (N10483, N10477, N4579);
not NOT1 (N10484, N10458);
or OR3 (N10485, N10484, N7656, N5607);
xor XOR2 (N10486, N10482, N5950);
nor NOR3 (N10487, N10483, N9084, N8311);
not NOT1 (N10488, N10487);
not NOT1 (N10489, N10481);
not NOT1 (N10490, N10478);
nand NAND4 (N10491, N10479, N1628, N9264, N2933);
buf BUF1 (N10492, N10474);
and AND3 (N10493, N10471, N7774, N10205);
or OR3 (N10494, N10488, N2556, N7281);
and AND4 (N10495, N10475, N5758, N372, N2848);
buf BUF1 (N10496, N10490);
not NOT1 (N10497, N10493);
not NOT1 (N10498, N10489);
buf BUF1 (N10499, N10485);
xor XOR2 (N10500, N10491, N3343);
or OR2 (N10501, N10496, N2988);
nand NAND2 (N10502, N10465, N6799);
and AND4 (N10503, N10500, N3671, N6324, N309);
and AND3 (N10504, N10498, N3328, N7774);
buf BUF1 (N10505, N10503);
or OR2 (N10506, N10505, N8336);
buf BUF1 (N10507, N10494);
nand NAND2 (N10508, N10497, N2602);
xor XOR2 (N10509, N10495, N6654);
nor NOR2 (N10510, N10509, N6640);
nor NOR3 (N10511, N10492, N1394, N4136);
xor XOR2 (N10512, N10507, N2943);
nor NOR4 (N10513, N10512, N172, N9079, N7252);
nand NAND3 (N10514, N10513, N2116, N1800);
and AND3 (N10515, N10511, N9510, N5760);
buf BUF1 (N10516, N10508);
not NOT1 (N10517, N10506);
nor NOR2 (N10518, N10517, N4753);
xor XOR2 (N10519, N10501, N1350);
xor XOR2 (N10520, N10519, N3606);
nor NOR2 (N10521, N10510, N4907);
xor XOR2 (N10522, N10504, N6944);
nand NAND2 (N10523, N10502, N1032);
nor NOR3 (N10524, N10499, N7691, N4602);
nand NAND4 (N10525, N10518, N5916, N8854, N1028);
xor XOR2 (N10526, N10520, N3330);
buf BUF1 (N10527, N10514);
buf BUF1 (N10528, N10516);
nor NOR2 (N10529, N10524, N7692);
or OR2 (N10530, N10486, N9204);
nand NAND4 (N10531, N10527, N58, N7871, N438);
xor XOR2 (N10532, N10530, N3446);
nand NAND3 (N10533, N10515, N3905, N10047);
not NOT1 (N10534, N10528);
nor NOR3 (N10535, N10521, N9794, N517);
buf BUF1 (N10536, N10532);
nor NOR4 (N10537, N10522, N6552, N8142, N7651);
not NOT1 (N10538, N10529);
nor NOR4 (N10539, N10534, N3406, N10497, N8451);
not NOT1 (N10540, N10533);
and AND4 (N10541, N10526, N8381, N9361, N6663);
not NOT1 (N10542, N10535);
buf BUF1 (N10543, N10537);
nor NOR3 (N10544, N10531, N6736, N1106);
xor XOR2 (N10545, N10543, N3633);
and AND2 (N10546, N10541, N2507);
nand NAND4 (N10547, N10545, N6927, N6463, N233);
xor XOR2 (N10548, N10539, N1042);
nand NAND4 (N10549, N10540, N10469, N7366, N4093);
xor XOR2 (N10550, N10544, N7537);
and AND4 (N10551, N10550, N1723, N3049, N5475);
not NOT1 (N10552, N10551);
nand NAND3 (N10553, N10536, N1016, N1504);
not NOT1 (N10554, N10546);
not NOT1 (N10555, N10542);
or OR2 (N10556, N10553, N8557);
and AND4 (N10557, N10555, N4238, N2923, N5810);
nor NOR3 (N10558, N10554, N6194, N4351);
xor XOR2 (N10559, N10548, N818);
nor NOR3 (N10560, N10538, N200, N4222);
xor XOR2 (N10561, N10556, N5449);
or OR3 (N10562, N10552, N1526, N8039);
xor XOR2 (N10563, N10562, N2768);
buf BUF1 (N10564, N10523);
and AND2 (N10565, N10564, N8457);
or OR4 (N10566, N10558, N5937, N6514, N898);
and AND4 (N10567, N10561, N8141, N243, N2050);
buf BUF1 (N10568, N10566);
not NOT1 (N10569, N10557);
buf BUF1 (N10570, N10525);
xor XOR2 (N10571, N10569, N2383);
not NOT1 (N10572, N10547);
nand NAND3 (N10573, N10559, N249, N2902);
or OR4 (N10574, N10571, N3875, N1414, N3771);
buf BUF1 (N10575, N10573);
buf BUF1 (N10576, N10568);
buf BUF1 (N10577, N10574);
not NOT1 (N10578, N10567);
or OR2 (N10579, N10563, N10184);
or OR3 (N10580, N10572, N4746, N6857);
and AND3 (N10581, N10549, N225, N8889);
buf BUF1 (N10582, N10575);
nor NOR4 (N10583, N10582, N5530, N2162, N3501);
and AND2 (N10584, N10580, N4045);
nand NAND3 (N10585, N10577, N613, N3842);
or OR4 (N10586, N10578, N8363, N181, N1008);
nor NOR4 (N10587, N10581, N8598, N7394, N6089);
nor NOR2 (N10588, N10576, N8359);
nand NAND3 (N10589, N10587, N4131, N6671);
or OR3 (N10590, N10579, N5591, N8194);
nand NAND2 (N10591, N10584, N1416);
xor XOR2 (N10592, N10565, N2554);
not NOT1 (N10593, N10570);
buf BUF1 (N10594, N10593);
nor NOR2 (N10595, N10585, N2382);
xor XOR2 (N10596, N10586, N8041);
buf BUF1 (N10597, N10589);
buf BUF1 (N10598, N10560);
buf BUF1 (N10599, N10588);
nor NOR2 (N10600, N10598, N4524);
not NOT1 (N10601, N10596);
nand NAND2 (N10602, N10599, N6009);
xor XOR2 (N10603, N10592, N12);
and AND2 (N10604, N10583, N6285);
or OR3 (N10605, N10604, N3164, N1531);
buf BUF1 (N10606, N10601);
xor XOR2 (N10607, N10591, N2436);
and AND4 (N10608, N10606, N3810, N5455, N2400);
and AND4 (N10609, N10597, N907, N7558, N9004);
not NOT1 (N10610, N10600);
nand NAND2 (N10611, N10590, N10226);
or OR4 (N10612, N10607, N5479, N961, N10402);
or OR2 (N10613, N10608, N9135);
and AND4 (N10614, N10609, N2200, N7224, N3055);
nor NOR3 (N10615, N10611, N707, N8406);
or OR4 (N10616, N10610, N9072, N7056, N7404);
not NOT1 (N10617, N10612);
nor NOR3 (N10618, N10617, N9454, N5046);
nor NOR4 (N10619, N10613, N8613, N6104, N10614);
and AND4 (N10620, N8903, N8091, N8994, N4921);
or OR4 (N10621, N10619, N4484, N7409, N6631);
and AND3 (N10622, N10616, N2665, N2183);
or OR3 (N10623, N10615, N1945, N2581);
and AND4 (N10624, N10623, N7497, N2260, N2447);
xor XOR2 (N10625, N10624, N6720);
and AND3 (N10626, N10595, N6199, N795);
xor XOR2 (N10627, N10603, N5211);
and AND4 (N10628, N10621, N1579, N6601, N6198);
and AND3 (N10629, N10625, N1532, N1118);
xor XOR2 (N10630, N10620, N4536);
and AND2 (N10631, N10630, N698);
nand NAND3 (N10632, N10605, N2129, N7435);
buf BUF1 (N10633, N10627);
or OR3 (N10634, N10602, N6133, N639);
xor XOR2 (N10635, N10633, N3980);
nor NOR3 (N10636, N10635, N6942, N6662);
not NOT1 (N10637, N10632);
and AND3 (N10638, N10594, N1237, N6577);
buf BUF1 (N10639, N10631);
buf BUF1 (N10640, N10636);
or OR4 (N10641, N10628, N1783, N3191, N8078);
and AND4 (N10642, N10629, N7373, N8395, N6328);
xor XOR2 (N10643, N10642, N8685);
nor NOR3 (N10644, N10634, N3392, N9935);
or OR3 (N10645, N10637, N1622, N9443);
or OR4 (N10646, N10645, N7944, N2554, N8691);
or OR3 (N10647, N10644, N2315, N3978);
xor XOR2 (N10648, N10641, N4601);
and AND2 (N10649, N10648, N9787);
nor NOR2 (N10650, N10618, N6871);
buf BUF1 (N10651, N10638);
xor XOR2 (N10652, N10639, N6243);
and AND2 (N10653, N10640, N1138);
and AND3 (N10654, N10649, N3084, N277);
or OR2 (N10655, N10650, N2854);
nor NOR4 (N10656, N10646, N3600, N10081, N4531);
and AND2 (N10657, N10652, N3877);
nor NOR4 (N10658, N10653, N9904, N3713, N4255);
nand NAND2 (N10659, N10622, N5774);
xor XOR2 (N10660, N10655, N9829);
nand NAND2 (N10661, N10654, N8422);
nand NAND3 (N10662, N10660, N10172, N174);
xor XOR2 (N10663, N10647, N3644);
not NOT1 (N10664, N10626);
not NOT1 (N10665, N10663);
xor XOR2 (N10666, N10661, N83);
nor NOR4 (N10667, N10659, N10227, N985, N6610);
or OR2 (N10668, N10662, N1393);
or OR3 (N10669, N10668, N6655, N568);
and AND3 (N10670, N10643, N9590, N901);
xor XOR2 (N10671, N10667, N6863);
xor XOR2 (N10672, N10656, N10129);
xor XOR2 (N10673, N10672, N8460);
nor NOR2 (N10674, N10666, N5594);
or OR3 (N10675, N10657, N7766, N5406);
or OR4 (N10676, N10658, N7438, N9020, N6757);
and AND3 (N10677, N10670, N4518, N9083);
xor XOR2 (N10678, N10673, N9172);
buf BUF1 (N10679, N10664);
xor XOR2 (N10680, N10677, N8683);
not NOT1 (N10681, N10671);
nor NOR3 (N10682, N10680, N4948, N10674);
buf BUF1 (N10683, N5401);
or OR3 (N10684, N10681, N3221, N7214);
or OR4 (N10685, N10684, N862, N602, N2106);
or OR2 (N10686, N10679, N8034);
and AND3 (N10687, N10675, N457, N9830);
buf BUF1 (N10688, N10665);
and AND4 (N10689, N10683, N3923, N6500, N158);
not NOT1 (N10690, N10669);
and AND3 (N10691, N10676, N6545, N4194);
and AND4 (N10692, N10689, N3173, N9842, N6185);
buf BUF1 (N10693, N10691);
xor XOR2 (N10694, N10690, N9718);
and AND2 (N10695, N10692, N10606);
nand NAND4 (N10696, N10687, N512, N8676, N1361);
nor NOR2 (N10697, N10651, N2169);
nor NOR4 (N10698, N10686, N5140, N2750, N962);
nor NOR3 (N10699, N10682, N1121, N7122);
nand NAND4 (N10700, N10695, N363, N5369, N8701);
nand NAND2 (N10701, N10685, N590);
not NOT1 (N10702, N10698);
xor XOR2 (N10703, N10697, N6692);
xor XOR2 (N10704, N10688, N3018);
buf BUF1 (N10705, N10702);
nand NAND4 (N10706, N10701, N5993, N6072, N9084);
nand NAND2 (N10707, N10704, N751);
not NOT1 (N10708, N10705);
nand NAND3 (N10709, N10706, N599, N6042);
not NOT1 (N10710, N10708);
nor NOR2 (N10711, N10707, N6228);
or OR4 (N10712, N10711, N8628, N10030, N7691);
nor NOR3 (N10713, N10703, N2995, N7966);
and AND2 (N10714, N10712, N4587);
or OR3 (N10715, N10714, N9043, N972);
and AND2 (N10716, N10694, N3506);
buf BUF1 (N10717, N10678);
buf BUF1 (N10718, N10709);
buf BUF1 (N10719, N10713);
or OR4 (N10720, N10719, N7375, N9672, N850);
buf BUF1 (N10721, N10699);
xor XOR2 (N10722, N10693, N6995);
nor NOR2 (N10723, N10722, N2779);
or OR3 (N10724, N10716, N5103, N9087);
and AND4 (N10725, N10710, N9706, N7191, N9065);
not NOT1 (N10726, N10725);
nand NAND2 (N10727, N10726, N7006);
xor XOR2 (N10728, N10715, N5705);
nand NAND3 (N10729, N10720, N9525, N8363);
or OR3 (N10730, N10696, N3297, N3530);
not NOT1 (N10731, N10729);
nor NOR3 (N10732, N10721, N6730, N2941);
and AND4 (N10733, N10731, N4321, N9870, N8453);
nor NOR4 (N10734, N10724, N4040, N338, N10388);
not NOT1 (N10735, N10723);
nand NAND4 (N10736, N10734, N9615, N3460, N6892);
xor XOR2 (N10737, N10732, N1841);
buf BUF1 (N10738, N10733);
and AND4 (N10739, N10700, N4080, N938, N2864);
or OR2 (N10740, N10738, N8437);
xor XOR2 (N10741, N10730, N4153);
not NOT1 (N10742, N10737);
xor XOR2 (N10743, N10735, N2254);
and AND3 (N10744, N10718, N10539, N4646);
nor NOR2 (N10745, N10742, N6496);
not NOT1 (N10746, N10727);
or OR3 (N10747, N10741, N5147, N7472);
not NOT1 (N10748, N10739);
not NOT1 (N10749, N10746);
nand NAND4 (N10750, N10748, N7960, N60, N2209);
nand NAND4 (N10751, N10717, N9000, N4590, N7440);
or OR4 (N10752, N10743, N8781, N6540, N9163);
and AND2 (N10753, N10750, N1462);
nand NAND4 (N10754, N10751, N3729, N6894, N1921);
or OR3 (N10755, N10728, N10442, N7152);
xor XOR2 (N10756, N10754, N10744);
not NOT1 (N10757, N8332);
or OR4 (N10758, N10757, N4650, N5745, N1883);
not NOT1 (N10759, N10758);
or OR3 (N10760, N10753, N2113, N8341);
nor NOR2 (N10761, N10756, N3280);
not NOT1 (N10762, N10740);
xor XOR2 (N10763, N10760, N9690);
nand NAND4 (N10764, N10747, N9610, N8478, N5651);
and AND3 (N10765, N10759, N6554, N10413);
nor NOR4 (N10766, N10762, N5413, N10656, N8310);
buf BUF1 (N10767, N10749);
xor XOR2 (N10768, N10752, N6433);
or OR2 (N10769, N10736, N8008);
and AND4 (N10770, N10766, N3250, N1308, N1972);
or OR4 (N10771, N10770, N8745, N10660, N3763);
not NOT1 (N10772, N10767);
not NOT1 (N10773, N10763);
and AND2 (N10774, N10755, N6360);
not NOT1 (N10775, N10765);
buf BUF1 (N10776, N10768);
buf BUF1 (N10777, N10771);
nor NOR2 (N10778, N10774, N1233);
and AND2 (N10779, N10764, N6129);
buf BUF1 (N10780, N10772);
nor NOR2 (N10781, N10776, N2748);
nor NOR3 (N10782, N10780, N5255, N10165);
nor NOR3 (N10783, N10761, N481, N2242);
or OR2 (N10784, N10745, N8355);
not NOT1 (N10785, N10777);
or OR3 (N10786, N10782, N7969, N8647);
or OR4 (N10787, N10785, N5686, N8270, N7467);
buf BUF1 (N10788, N10773);
not NOT1 (N10789, N10784);
not NOT1 (N10790, N10778);
or OR3 (N10791, N10783, N8452, N8284);
nand NAND4 (N10792, N10791, N159, N83, N274);
nand NAND4 (N10793, N10792, N9017, N9865, N4709);
not NOT1 (N10794, N10781);
nor NOR4 (N10795, N10779, N3055, N3647, N3437);
or OR4 (N10796, N10787, N4445, N1417, N334);
nand NAND3 (N10797, N10786, N7032, N1890);
not NOT1 (N10798, N10790);
nor NOR3 (N10799, N10789, N1071, N5748);
and AND4 (N10800, N10769, N4308, N9528, N5385);
not NOT1 (N10801, N10799);
or OR3 (N10802, N10788, N7605, N10214);
or OR2 (N10803, N10801, N6708);
nand NAND2 (N10804, N10802, N9156);
not NOT1 (N10805, N10795);
or OR3 (N10806, N10793, N1800, N2992);
and AND3 (N10807, N10805, N7809, N3867);
or OR3 (N10808, N10796, N1541, N5125);
xor XOR2 (N10809, N10800, N1291);
buf BUF1 (N10810, N10797);
and AND3 (N10811, N10807, N7122, N8048);
buf BUF1 (N10812, N10804);
or OR2 (N10813, N10794, N753);
xor XOR2 (N10814, N10812, N188);
nand NAND2 (N10815, N10811, N2309);
or OR3 (N10816, N10815, N6937, N9401);
xor XOR2 (N10817, N10816, N4556);
not NOT1 (N10818, N10775);
and AND2 (N10819, N10814, N134);
and AND4 (N10820, N10809, N3887, N9518, N515);
xor XOR2 (N10821, N10813, N4755);
and AND2 (N10822, N10818, N4827);
nor NOR3 (N10823, N10810, N1959, N1803);
buf BUF1 (N10824, N10823);
nand NAND2 (N10825, N10822, N4180);
xor XOR2 (N10826, N10798, N3330);
or OR4 (N10827, N10808, N4128, N8150, N2385);
buf BUF1 (N10828, N10803);
xor XOR2 (N10829, N10825, N3073);
not NOT1 (N10830, N10806);
nor NOR3 (N10831, N10830, N910, N6872);
xor XOR2 (N10832, N10819, N8246);
not NOT1 (N10833, N10831);
buf BUF1 (N10834, N10827);
xor XOR2 (N10835, N10832, N9467);
nand NAND4 (N10836, N10835, N883, N2871, N8684);
xor XOR2 (N10837, N10828, N4102);
and AND3 (N10838, N10826, N1592, N4599);
or OR4 (N10839, N10833, N9096, N7940, N5910);
xor XOR2 (N10840, N10836, N1776);
nor NOR3 (N10841, N10824, N8969, N8188);
xor XOR2 (N10842, N10841, N230);
xor XOR2 (N10843, N10834, N8800);
nor NOR3 (N10844, N10842, N2347, N6277);
not NOT1 (N10845, N10840);
buf BUF1 (N10846, N10817);
nand NAND3 (N10847, N10820, N8418, N6860);
not NOT1 (N10848, N10837);
nand NAND3 (N10849, N10838, N3397, N1364);
or OR4 (N10850, N10844, N1004, N8730, N9577);
buf BUF1 (N10851, N10847);
xor XOR2 (N10852, N10845, N7491);
nand NAND3 (N10853, N10851, N1958, N6698);
xor XOR2 (N10854, N10853, N1783);
and AND4 (N10855, N10846, N3408, N1630, N2696);
or OR4 (N10856, N10850, N2709, N3273, N10469);
buf BUF1 (N10857, N10849);
nand NAND3 (N10858, N10854, N4762, N7410);
and AND3 (N10859, N10858, N3131, N45);
and AND3 (N10860, N10839, N1891, N3183);
nand NAND4 (N10861, N10860, N6074, N1868, N3055);
not NOT1 (N10862, N10859);
nand NAND3 (N10863, N10862, N7886, N2816);
buf BUF1 (N10864, N10857);
buf BUF1 (N10865, N10852);
and AND2 (N10866, N10848, N2791);
nand NAND2 (N10867, N10829, N1373);
xor XOR2 (N10868, N10855, N5850);
and AND3 (N10869, N10861, N3047, N4622);
not NOT1 (N10870, N10868);
xor XOR2 (N10871, N10870, N2191);
nand NAND3 (N10872, N10843, N6110, N8847);
not NOT1 (N10873, N10872);
xor XOR2 (N10874, N10856, N7977);
and AND3 (N10875, N10866, N8193, N10543);
nand NAND4 (N10876, N10871, N10066, N10599, N6125);
buf BUF1 (N10877, N10865);
nor NOR2 (N10878, N10876, N9641);
or OR3 (N10879, N10864, N956, N10040);
or OR2 (N10880, N10875, N2186);
nand NAND3 (N10881, N10821, N9087, N2665);
nand NAND2 (N10882, N10869, N10773);
not NOT1 (N10883, N10878);
or OR3 (N10884, N10879, N3430, N2992);
nor NOR2 (N10885, N10884, N444);
or OR3 (N10886, N10877, N9615, N4065);
buf BUF1 (N10887, N10874);
nor NOR4 (N10888, N10886, N9374, N1304, N9890);
nor NOR4 (N10889, N10883, N5146, N8865, N4602);
nor NOR2 (N10890, N10887, N10108);
nand NAND2 (N10891, N10863, N2795);
buf BUF1 (N10892, N10867);
or OR3 (N10893, N10890, N4683, N2987);
not NOT1 (N10894, N10880);
or OR3 (N10895, N10888, N7573, N2170);
and AND2 (N10896, N10873, N6099);
and AND3 (N10897, N10895, N3324, N4061);
buf BUF1 (N10898, N10897);
nor NOR2 (N10899, N10882, N9559);
or OR2 (N10900, N10892, N9189);
xor XOR2 (N10901, N10899, N124);
buf BUF1 (N10902, N10891);
or OR3 (N10903, N10901, N4378, N1337);
buf BUF1 (N10904, N10881);
nand NAND4 (N10905, N10896, N3865, N3421, N1855);
buf BUF1 (N10906, N10905);
not NOT1 (N10907, N10906);
xor XOR2 (N10908, N10893, N1459);
nor NOR4 (N10909, N10898, N6010, N4145, N10873);
not NOT1 (N10910, N10908);
and AND4 (N10911, N10894, N2145, N6336, N7080);
nand NAND4 (N10912, N10903, N7807, N349, N9160);
xor XOR2 (N10913, N10910, N2105);
and AND4 (N10914, N10900, N9231, N6691, N3999);
xor XOR2 (N10915, N10913, N5327);
nor NOR4 (N10916, N10911, N4025, N9907, N7351);
and AND4 (N10917, N10912, N8401, N2844, N5318);
and AND3 (N10918, N10904, N6472, N9875);
buf BUF1 (N10919, N10885);
nand NAND3 (N10920, N10909, N5861, N91);
or OR4 (N10921, N10915, N10490, N4562, N6708);
and AND3 (N10922, N10920, N4124, N6589);
buf BUF1 (N10923, N10919);
nand NAND4 (N10924, N10914, N3659, N9005, N5885);
and AND3 (N10925, N10922, N4684, N2965);
buf BUF1 (N10926, N10907);
buf BUF1 (N10927, N10902);
xor XOR2 (N10928, N10927, N8181);
and AND3 (N10929, N10918, N635, N7664);
buf BUF1 (N10930, N10923);
and AND2 (N10931, N10924, N2151);
and AND2 (N10932, N10931, N4037);
and AND2 (N10933, N10930, N9151);
and AND4 (N10934, N10925, N7697, N1852, N567);
not NOT1 (N10935, N10934);
nor NOR3 (N10936, N10926, N2622, N4666);
buf BUF1 (N10937, N10921);
or OR4 (N10938, N10932, N7682, N3944, N2098);
nor NOR4 (N10939, N10889, N6802, N8658, N4778);
nand NAND3 (N10940, N10916, N5129, N4407);
not NOT1 (N10941, N10939);
nor NOR2 (N10942, N10941, N9187);
and AND3 (N10943, N10936, N503, N7403);
not NOT1 (N10944, N10937);
xor XOR2 (N10945, N10942, N8252);
or OR2 (N10946, N10917, N7474);
buf BUF1 (N10947, N10946);
not NOT1 (N10948, N10929);
not NOT1 (N10949, N10947);
nor NOR4 (N10950, N10944, N252, N4671, N4276);
buf BUF1 (N10951, N10943);
or OR4 (N10952, N10933, N59, N6098, N1521);
xor XOR2 (N10953, N10940, N7737);
nor NOR4 (N10954, N10953, N7686, N514, N2070);
not NOT1 (N10955, N10928);
not NOT1 (N10956, N10952);
not NOT1 (N10957, N10945);
nand NAND4 (N10958, N10948, N9476, N3154, N8091);
nand NAND3 (N10959, N10951, N4886, N2981);
buf BUF1 (N10960, N10954);
not NOT1 (N10961, N10959);
not NOT1 (N10962, N10955);
not NOT1 (N10963, N10956);
buf BUF1 (N10964, N10962);
or OR2 (N10965, N10960, N8900);
not NOT1 (N10966, N10965);
and AND3 (N10967, N10964, N7327, N6854);
buf BUF1 (N10968, N10938);
and AND3 (N10969, N10958, N3660, N4549);
or OR3 (N10970, N10969, N2175, N10033);
nand NAND4 (N10971, N10961, N1291, N8963, N7348);
not NOT1 (N10972, N10935);
buf BUF1 (N10973, N10972);
nand NAND4 (N10974, N10950, N3358, N10850, N3179);
or OR4 (N10975, N10966, N5735, N5212, N10131);
nor NOR2 (N10976, N10975, N5045);
and AND3 (N10977, N10976, N4689, N1357);
or OR2 (N10978, N10963, N5241);
or OR4 (N10979, N10974, N7393, N1527, N35);
buf BUF1 (N10980, N10971);
not NOT1 (N10981, N10977);
or OR3 (N10982, N10978, N4361, N7951);
nor NOR2 (N10983, N10970, N5071);
nor NOR4 (N10984, N10957, N703, N3840, N796);
nand NAND2 (N10985, N10973, N140);
nor NOR3 (N10986, N10982, N9894, N4230);
nor NOR3 (N10987, N10985, N264, N6076);
nand NAND4 (N10988, N10987, N2010, N8667, N3354);
or OR3 (N10989, N10980, N6455, N2859);
not NOT1 (N10990, N10981);
buf BUF1 (N10991, N10988);
or OR3 (N10992, N10979, N1098, N8941);
not NOT1 (N10993, N10990);
nor NOR2 (N10994, N10984, N3255);
nor NOR3 (N10995, N10967, N7842, N2021);
not NOT1 (N10996, N10991);
not NOT1 (N10997, N10986);
xor XOR2 (N10998, N10995, N5228);
buf BUF1 (N10999, N10949);
not NOT1 (N11000, N10994);
not NOT1 (N11001, N10996);
and AND2 (N11002, N10998, N8552);
and AND4 (N11003, N10997, N2580, N1609, N10032);
nor NOR4 (N11004, N11000, N7352, N4422, N1418);
xor XOR2 (N11005, N10989, N6536);
nor NOR2 (N11006, N11002, N3036);
nand NAND3 (N11007, N11005, N2169, N3920);
or OR3 (N11008, N11003, N1373, N10510);
nand NAND4 (N11009, N10992, N3245, N10675, N4373);
xor XOR2 (N11010, N11009, N4482);
buf BUF1 (N11011, N11010);
and AND3 (N11012, N10983, N5350, N8416);
xor XOR2 (N11013, N11007, N10816);
buf BUF1 (N11014, N11013);
and AND3 (N11015, N11011, N5671, N3371);
buf BUF1 (N11016, N11015);
nand NAND3 (N11017, N11016, N1515, N700);
not NOT1 (N11018, N11001);
xor XOR2 (N11019, N11018, N5311);
xor XOR2 (N11020, N10968, N3260);
xor XOR2 (N11021, N10999, N1803);
buf BUF1 (N11022, N11012);
buf BUF1 (N11023, N11017);
and AND4 (N11024, N11022, N8855, N4513, N8845);
and AND4 (N11025, N11023, N10553, N6392, N1360);
or OR3 (N11026, N11019, N2518, N9132);
not NOT1 (N11027, N11006);
and AND4 (N11028, N11024, N6791, N6043, N6946);
buf BUF1 (N11029, N11014);
buf BUF1 (N11030, N11028);
buf BUF1 (N11031, N11027);
nand NAND3 (N11032, N11021, N4728, N7337);
not NOT1 (N11033, N11032);
and AND2 (N11034, N11025, N1288);
and AND2 (N11035, N11004, N1264);
not NOT1 (N11036, N11031);
and AND3 (N11037, N11026, N6359, N10062);
and AND4 (N11038, N11037, N7302, N6698, N6818);
nand NAND4 (N11039, N11020, N1837, N3133, N216);
nand NAND3 (N11040, N11030, N7132, N6256);
xor XOR2 (N11041, N11029, N7418);
or OR3 (N11042, N11041, N9982, N4843);
nor NOR4 (N11043, N11008, N528, N10337, N4854);
or OR3 (N11044, N11042, N6628, N8126);
xor XOR2 (N11045, N11038, N3645);
xor XOR2 (N11046, N11045, N10446);
nor NOR4 (N11047, N11046, N1265, N3320, N4270);
buf BUF1 (N11048, N11036);
and AND3 (N11049, N11039, N9560, N4642);
xor XOR2 (N11050, N11043, N3985);
not NOT1 (N11051, N10993);
nand NAND2 (N11052, N11049, N1867);
nand NAND4 (N11053, N11048, N2705, N8107, N572);
buf BUF1 (N11054, N11033);
nor NOR3 (N11055, N11040, N4120, N6613);
and AND3 (N11056, N11055, N2316, N2278);
buf BUF1 (N11057, N11051);
not NOT1 (N11058, N11052);
buf BUF1 (N11059, N11054);
not NOT1 (N11060, N11035);
or OR2 (N11061, N11034, N10793);
and AND4 (N11062, N11061, N3420, N9052, N7567);
not NOT1 (N11063, N11057);
and AND3 (N11064, N11047, N9209, N2229);
nand NAND2 (N11065, N11064, N6520);
buf BUF1 (N11066, N11050);
or OR4 (N11067, N11053, N8975, N4162, N6241);
nor NOR3 (N11068, N11059, N3140, N6125);
buf BUF1 (N11069, N11044);
nand NAND3 (N11070, N11069, N9382, N8504);
buf BUF1 (N11071, N11058);
or OR4 (N11072, N11063, N8521, N5287, N9050);
or OR4 (N11073, N11068, N377, N1573, N7656);
xor XOR2 (N11074, N11071, N11009);
and AND3 (N11075, N11066, N5858, N8786);
or OR3 (N11076, N11075, N8558, N2448);
xor XOR2 (N11077, N11070, N953);
or OR4 (N11078, N11072, N8659, N10292, N2425);
nand NAND2 (N11079, N11065, N7613);
or OR4 (N11080, N11074, N7184, N5674, N1453);
not NOT1 (N11081, N11076);
or OR4 (N11082, N11077, N10204, N1233, N5064);
nor NOR3 (N11083, N11056, N6728, N3457);
xor XOR2 (N11084, N11079, N8366);
and AND3 (N11085, N11060, N2658, N8524);
buf BUF1 (N11086, N11078);
and AND4 (N11087, N11073, N7679, N6850, N4378);
buf BUF1 (N11088, N11082);
or OR2 (N11089, N11081, N8229);
xor XOR2 (N11090, N11080, N2044);
nand NAND4 (N11091, N11085, N3683, N5155, N2600);
nand NAND3 (N11092, N11062, N8482, N7814);
not NOT1 (N11093, N11083);
and AND2 (N11094, N11087, N840);
buf BUF1 (N11095, N11088);
nand NAND3 (N11096, N11091, N3583, N9583);
xor XOR2 (N11097, N11067, N1895);
xor XOR2 (N11098, N11097, N10954);
not NOT1 (N11099, N11098);
and AND3 (N11100, N11086, N1297, N300);
not NOT1 (N11101, N11095);
nand NAND4 (N11102, N11089, N6560, N9164, N1016);
and AND3 (N11103, N11090, N7852, N4867);
nand NAND2 (N11104, N11096, N1991);
buf BUF1 (N11105, N11099);
nand NAND3 (N11106, N11102, N2794, N5699);
nor NOR3 (N11107, N11092, N10097, N2203);
nand NAND2 (N11108, N11104, N4111);
buf BUF1 (N11109, N11100);
nand NAND3 (N11110, N11093, N2736, N2222);
xor XOR2 (N11111, N11101, N6335);
xor XOR2 (N11112, N11109, N3582);
not NOT1 (N11113, N11106);
not NOT1 (N11114, N11111);
nand NAND2 (N11115, N11108, N3232);
nand NAND2 (N11116, N11084, N8252);
nor NOR4 (N11117, N11115, N1611, N5490, N3939);
and AND4 (N11118, N11094, N10471, N903, N7101);
or OR4 (N11119, N11114, N10557, N9282, N10409);
not NOT1 (N11120, N11107);
and AND2 (N11121, N11105, N9179);
xor XOR2 (N11122, N11119, N5337);
buf BUF1 (N11123, N11110);
nor NOR2 (N11124, N11123, N4218);
nand NAND4 (N11125, N11112, N276, N6973, N5673);
nor NOR4 (N11126, N11121, N4804, N482, N3038);
xor XOR2 (N11127, N11103, N7029);
nand NAND2 (N11128, N11118, N9803);
and AND2 (N11129, N11128, N9397);
and AND2 (N11130, N11116, N3610);
not NOT1 (N11131, N11130);
and AND4 (N11132, N11117, N2575, N889, N221);
and AND3 (N11133, N11113, N706, N3579);
buf BUF1 (N11134, N11131);
xor XOR2 (N11135, N11133, N5553);
nand NAND2 (N11136, N11125, N2144);
xor XOR2 (N11137, N11120, N505);
nand NAND2 (N11138, N11122, N1807);
and AND2 (N11139, N11132, N328);
nor NOR3 (N11140, N11124, N5791, N7763);
not NOT1 (N11141, N11129);
not NOT1 (N11142, N11138);
not NOT1 (N11143, N11127);
buf BUF1 (N11144, N11139);
buf BUF1 (N11145, N11143);
nand NAND2 (N11146, N11137, N89);
not NOT1 (N11147, N11126);
and AND3 (N11148, N11136, N3388, N8713);
nand NAND3 (N11149, N11144, N590, N7566);
not NOT1 (N11150, N11141);
and AND3 (N11151, N11135, N722, N7093);
not NOT1 (N11152, N11147);
or OR4 (N11153, N11146, N5216, N1801, N10792);
xor XOR2 (N11154, N11152, N9197);
nand NAND4 (N11155, N11134, N3460, N4007, N94);
or OR2 (N11156, N11151, N5804);
nand NAND2 (N11157, N11156, N3533);
and AND3 (N11158, N11148, N7999, N2427);
nor NOR4 (N11159, N11157, N4508, N4048, N2662);
xor XOR2 (N11160, N11140, N5797);
nor NOR4 (N11161, N11145, N3032, N9192, N8582);
not NOT1 (N11162, N11158);
nor NOR2 (N11163, N11154, N3572);
xor XOR2 (N11164, N11155, N5007);
nand NAND2 (N11165, N11162, N7284);
nor NOR4 (N11166, N11159, N2145, N7867, N8188);
buf BUF1 (N11167, N11142);
not NOT1 (N11168, N11150);
nor NOR4 (N11169, N11167, N3115, N9110, N9281);
buf BUF1 (N11170, N11149);
nor NOR2 (N11171, N11160, N2512);
buf BUF1 (N11172, N11166);
and AND2 (N11173, N11171, N8653);
not NOT1 (N11174, N11164);
nand NAND2 (N11175, N11161, N3551);
or OR2 (N11176, N11174, N6286);
nor NOR3 (N11177, N11172, N8079, N581);
nor NOR2 (N11178, N11165, N8861);
and AND4 (N11179, N11178, N9466, N5365, N4114);
nand NAND4 (N11180, N11175, N6265, N6735, N9398);
nand NAND4 (N11181, N11168, N5495, N3653, N8664);
nand NAND4 (N11182, N11177, N8569, N9769, N4344);
buf BUF1 (N11183, N11169);
not NOT1 (N11184, N11170);
buf BUF1 (N11185, N11153);
or OR2 (N11186, N11163, N7398);
xor XOR2 (N11187, N11176, N7616);
buf BUF1 (N11188, N11186);
not NOT1 (N11189, N11182);
or OR2 (N11190, N11185, N6818);
xor XOR2 (N11191, N11183, N8408);
buf BUF1 (N11192, N11191);
buf BUF1 (N11193, N11181);
nor NOR4 (N11194, N11180, N9059, N7430, N5286);
not NOT1 (N11195, N11194);
and AND2 (N11196, N11188, N2998);
and AND2 (N11197, N11184, N3866);
nor NOR3 (N11198, N11195, N7426, N7176);
not NOT1 (N11199, N11189);
nor NOR2 (N11200, N11190, N7929);
buf BUF1 (N11201, N11198);
nor NOR4 (N11202, N11179, N2200, N10358, N9983);
or OR4 (N11203, N11202, N7985, N5785, N2805);
nand NAND2 (N11204, N11173, N4552);
not NOT1 (N11205, N11193);
nand NAND4 (N11206, N11196, N2714, N3812, N8177);
nand NAND2 (N11207, N11204, N10994);
nor NOR2 (N11208, N11187, N6762);
not NOT1 (N11209, N11208);
xor XOR2 (N11210, N11197, N4189);
nor NOR4 (N11211, N11210, N9124, N6566, N4080);
nor NOR3 (N11212, N11201, N8638, N1730);
and AND2 (N11213, N11200, N1604);
and AND4 (N11214, N11207, N8116, N9701, N9703);
or OR3 (N11215, N11214, N6646, N2629);
and AND2 (N11216, N11213, N3969);
buf BUF1 (N11217, N11216);
and AND4 (N11218, N11203, N824, N1915, N103);
nand NAND2 (N11219, N11217, N1992);
nor NOR4 (N11220, N11215, N1850, N7749, N8409);
buf BUF1 (N11221, N11212);
nand NAND2 (N11222, N11199, N8386);
and AND3 (N11223, N11211, N7849, N10326);
or OR2 (N11224, N11218, N4040);
not NOT1 (N11225, N11206);
nand NAND4 (N11226, N11220, N2952, N4862, N6451);
and AND2 (N11227, N11192, N5545);
and AND2 (N11228, N11227, N7849);
or OR3 (N11229, N11226, N914, N5071);
nand NAND4 (N11230, N11228, N602, N1205, N9278);
or OR2 (N11231, N11230, N5453);
or OR4 (N11232, N11223, N10878, N50, N1038);
buf BUF1 (N11233, N11222);
not NOT1 (N11234, N11225);
and AND4 (N11235, N11221, N8932, N4881, N8861);
or OR2 (N11236, N11232, N8418);
not NOT1 (N11237, N11233);
not NOT1 (N11238, N11205);
buf BUF1 (N11239, N11219);
or OR2 (N11240, N11224, N1188);
not NOT1 (N11241, N11236);
xor XOR2 (N11242, N11235, N10058);
nand NAND3 (N11243, N11234, N5782, N9819);
or OR2 (N11244, N11238, N10681);
and AND3 (N11245, N11209, N4314, N9220);
nand NAND4 (N11246, N11242, N5355, N7961, N1792);
xor XOR2 (N11247, N11237, N3829);
buf BUF1 (N11248, N11245);
buf BUF1 (N11249, N11246);
not NOT1 (N11250, N11247);
or OR4 (N11251, N11239, N9158, N138, N6272);
not NOT1 (N11252, N11229);
buf BUF1 (N11253, N11248);
nand NAND3 (N11254, N11253, N5055, N5778);
nor NOR2 (N11255, N11231, N10041);
or OR4 (N11256, N11250, N10579, N4067, N6136);
not NOT1 (N11257, N11249);
not NOT1 (N11258, N11252);
nor NOR2 (N11259, N11254, N5886);
nor NOR4 (N11260, N11256, N3578, N5179, N2587);
nand NAND4 (N11261, N11240, N2792, N10581, N3346);
nand NAND2 (N11262, N11241, N8411);
nand NAND2 (N11263, N11258, N10392);
or OR4 (N11264, N11257, N4690, N1855, N7525);
nand NAND3 (N11265, N11264, N3900, N3932);
or OR4 (N11266, N11243, N6229, N633, N3411);
nor NOR4 (N11267, N11259, N11138, N2346, N796);
and AND2 (N11268, N11266, N498);
nor NOR2 (N11269, N11265, N9571);
not NOT1 (N11270, N11260);
xor XOR2 (N11271, N11261, N5268);
or OR3 (N11272, N11270, N5950, N1774);
not NOT1 (N11273, N11251);
xor XOR2 (N11274, N11268, N7636);
buf BUF1 (N11275, N11262);
or OR4 (N11276, N11275, N4449, N8975, N137);
or OR3 (N11277, N11255, N8362, N7119);
and AND3 (N11278, N11277, N8665, N8226);
and AND4 (N11279, N11276, N4635, N11073, N4325);
xor XOR2 (N11280, N11278, N679);
or OR4 (N11281, N11279, N1828, N8914, N5798);
nor NOR4 (N11282, N11280, N1194, N3247, N10323);
xor XOR2 (N11283, N11273, N2975);
nand NAND2 (N11284, N11267, N5617);
or OR4 (N11285, N11284, N9051, N6791, N10702);
buf BUF1 (N11286, N11282);
nand NAND4 (N11287, N11274, N1683, N10935, N7370);
and AND2 (N11288, N11287, N1591);
not NOT1 (N11289, N11286);
buf BUF1 (N11290, N11271);
xor XOR2 (N11291, N11263, N9086);
buf BUF1 (N11292, N11291);
and AND4 (N11293, N11289, N4119, N7057, N7135);
buf BUF1 (N11294, N11283);
xor XOR2 (N11295, N11290, N1909);
not NOT1 (N11296, N11288);
nor NOR3 (N11297, N11281, N2006, N344);
nor NOR3 (N11298, N11293, N10256, N1441);
xor XOR2 (N11299, N11269, N10842);
xor XOR2 (N11300, N11295, N5930);
not NOT1 (N11301, N11298);
xor XOR2 (N11302, N11299, N7771);
buf BUF1 (N11303, N11302);
xor XOR2 (N11304, N11301, N5810);
or OR2 (N11305, N11272, N297);
nand NAND4 (N11306, N11300, N2381, N3869, N4204);
nand NAND2 (N11307, N11297, N7459);
nand NAND2 (N11308, N11305, N83);
nor NOR4 (N11309, N11306, N8462, N4831, N3251);
and AND2 (N11310, N11296, N2585);
or OR4 (N11311, N11303, N336, N9151, N8138);
or OR3 (N11312, N11294, N3068, N3723);
or OR2 (N11313, N11309, N8710);
buf BUF1 (N11314, N11310);
or OR4 (N11315, N11307, N9098, N4532, N9592);
xor XOR2 (N11316, N11314, N8266);
nor NOR4 (N11317, N11244, N9024, N2125, N4099);
xor XOR2 (N11318, N11316, N880);
or OR3 (N11319, N11315, N7836, N87);
not NOT1 (N11320, N11313);
or OR2 (N11321, N11312, N6344);
not NOT1 (N11322, N11317);
nor NOR4 (N11323, N11322, N6850, N2120, N5270);
buf BUF1 (N11324, N11323);
or OR2 (N11325, N11311, N10370);
xor XOR2 (N11326, N11318, N4799);
nor NOR2 (N11327, N11304, N3449);
buf BUF1 (N11328, N11308);
xor XOR2 (N11329, N11321, N4110);
or OR2 (N11330, N11285, N5645);
or OR3 (N11331, N11330, N5385, N6188);
nand NAND3 (N11332, N11326, N11121, N2410);
not NOT1 (N11333, N11292);
and AND2 (N11334, N11320, N3748);
buf BUF1 (N11335, N11325);
nand NAND3 (N11336, N11329, N6508, N8232);
and AND2 (N11337, N11332, N4342);
buf BUF1 (N11338, N11333);
not NOT1 (N11339, N11327);
nand NAND4 (N11340, N11336, N10583, N633, N5271);
not NOT1 (N11341, N11331);
nor NOR4 (N11342, N11339, N581, N10799, N11158);
or OR4 (N11343, N11340, N9717, N4661, N1632);
not NOT1 (N11344, N11341);
nor NOR3 (N11345, N11319, N4395, N10579);
not NOT1 (N11346, N11335);
buf BUF1 (N11347, N11346);
or OR4 (N11348, N11338, N2232, N4750, N10290);
buf BUF1 (N11349, N11342);
xor XOR2 (N11350, N11343, N8868);
not NOT1 (N11351, N11349);
or OR4 (N11352, N11348, N9768, N7213, N10105);
xor XOR2 (N11353, N11334, N982);
not NOT1 (N11354, N11350);
buf BUF1 (N11355, N11354);
not NOT1 (N11356, N11353);
nor NOR4 (N11357, N11324, N9998, N5269, N10526);
and AND3 (N11358, N11351, N9946, N5301);
xor XOR2 (N11359, N11328, N189);
buf BUF1 (N11360, N11359);
or OR4 (N11361, N11356, N8768, N829, N10868);
not NOT1 (N11362, N11360);
and AND2 (N11363, N11358, N6616);
or OR4 (N11364, N11355, N9918, N11064, N3191);
or OR4 (N11365, N11337, N3316, N7341, N5237);
nor NOR3 (N11366, N11364, N6527, N6814);
nor NOR2 (N11367, N11357, N1479);
not NOT1 (N11368, N11367);
buf BUF1 (N11369, N11362);
nor NOR2 (N11370, N11347, N10352);
xor XOR2 (N11371, N11369, N6194);
or OR4 (N11372, N11365, N8324, N8813, N6146);
xor XOR2 (N11373, N11352, N1469);
nor NOR4 (N11374, N11372, N1964, N2178, N7495);
nor NOR2 (N11375, N11363, N10342);
not NOT1 (N11376, N11345);
not NOT1 (N11377, N11366);
nand NAND2 (N11378, N11374, N9689);
buf BUF1 (N11379, N11344);
xor XOR2 (N11380, N11373, N7542);
and AND4 (N11381, N11368, N5332, N6032, N4122);
or OR3 (N11382, N11371, N5379, N9976);
xor XOR2 (N11383, N11370, N9062);
nand NAND4 (N11384, N11383, N10765, N11243, N819);
xor XOR2 (N11385, N11376, N10890);
xor XOR2 (N11386, N11380, N7220);
not NOT1 (N11387, N11381);
xor XOR2 (N11388, N11387, N2469);
xor XOR2 (N11389, N11375, N2606);
nand NAND2 (N11390, N11386, N3208);
or OR3 (N11391, N11389, N1475, N4929);
or OR3 (N11392, N11361, N11153, N2994);
or OR4 (N11393, N11384, N3774, N2694, N3550);
not NOT1 (N11394, N11382);
nand NAND4 (N11395, N11392, N497, N698, N1446);
xor XOR2 (N11396, N11385, N2387);
buf BUF1 (N11397, N11390);
or OR3 (N11398, N11377, N6438, N5224);
nor NOR2 (N11399, N11378, N3058);
or OR4 (N11400, N11379, N9736, N9990, N3709);
buf BUF1 (N11401, N11391);
not NOT1 (N11402, N11398);
xor XOR2 (N11403, N11396, N710);
nor NOR2 (N11404, N11394, N4250);
nor NOR2 (N11405, N11395, N6945);
xor XOR2 (N11406, N11404, N706);
not NOT1 (N11407, N11401);
xor XOR2 (N11408, N11406, N2720);
xor XOR2 (N11409, N11407, N6329);
nor NOR2 (N11410, N11399, N2558);
nor NOR4 (N11411, N11408, N1510, N8212, N6410);
buf BUF1 (N11412, N11388);
buf BUF1 (N11413, N11400);
nor NOR4 (N11414, N11409, N3464, N4280, N10365);
not NOT1 (N11415, N11403);
not NOT1 (N11416, N11414);
xor XOR2 (N11417, N11415, N7656);
nor NOR4 (N11418, N11416, N10305, N10074, N5461);
nor NOR4 (N11419, N11397, N380, N1699, N3569);
and AND4 (N11420, N11410, N6576, N3362, N9907);
and AND3 (N11421, N11412, N9364, N10419);
xor XOR2 (N11422, N11405, N10110);
nand NAND2 (N11423, N11413, N6602);
or OR3 (N11424, N11421, N8454, N7812);
or OR2 (N11425, N11411, N5692);
and AND3 (N11426, N11425, N5989, N11020);
xor XOR2 (N11427, N11417, N6440);
and AND2 (N11428, N11426, N8887);
buf BUF1 (N11429, N11428);
not NOT1 (N11430, N11420);
buf BUF1 (N11431, N11429);
xor XOR2 (N11432, N11419, N7826);
and AND4 (N11433, N11431, N9505, N6269, N8737);
xor XOR2 (N11434, N11433, N10553);
buf BUF1 (N11435, N11424);
nor NOR2 (N11436, N11430, N11207);
not NOT1 (N11437, N11422);
and AND2 (N11438, N11436, N9022);
buf BUF1 (N11439, N11402);
or OR3 (N11440, N11435, N84, N4754);
or OR3 (N11441, N11438, N8377, N4318);
xor XOR2 (N11442, N11432, N1774);
nor NOR3 (N11443, N11440, N4264, N9647);
nor NOR2 (N11444, N11442, N5360);
nand NAND3 (N11445, N11439, N9890, N1583);
nor NOR4 (N11446, N11443, N3986, N2993, N2635);
xor XOR2 (N11447, N11445, N2253);
nand NAND3 (N11448, N11418, N5016, N5437);
and AND3 (N11449, N11441, N7689, N6856);
nor NOR2 (N11450, N11448, N1638);
nand NAND4 (N11451, N11423, N8624, N3748, N10754);
or OR2 (N11452, N11393, N3029);
and AND3 (N11453, N11451, N9338, N5725);
buf BUF1 (N11454, N11446);
buf BUF1 (N11455, N11452);
and AND4 (N11456, N11434, N8605, N6702, N10718);
nand NAND4 (N11457, N11437, N8549, N10610, N9020);
not NOT1 (N11458, N11444);
not NOT1 (N11459, N11454);
xor XOR2 (N11460, N11458, N9555);
and AND4 (N11461, N11453, N1925, N6655, N3754);
nand NAND2 (N11462, N11450, N5918);
not NOT1 (N11463, N11427);
buf BUF1 (N11464, N11461);
or OR3 (N11465, N11462, N7483, N9441);
and AND4 (N11466, N11449, N10257, N767, N6706);
xor XOR2 (N11467, N11457, N9145);
xor XOR2 (N11468, N11464, N9163);
nor NOR3 (N11469, N11460, N6983, N7495);
nor NOR2 (N11470, N11468, N9199);
xor XOR2 (N11471, N11447, N1399);
xor XOR2 (N11472, N11455, N6147);
not NOT1 (N11473, N11470);
nand NAND2 (N11474, N11465, N1529);
buf BUF1 (N11475, N11456);
not NOT1 (N11476, N11475);
not NOT1 (N11477, N11459);
xor XOR2 (N11478, N11463, N3842);
buf BUF1 (N11479, N11478);
buf BUF1 (N11480, N11471);
and AND4 (N11481, N11473, N1241, N8743, N6460);
nand NAND2 (N11482, N11481, N8776);
not NOT1 (N11483, N11466);
nand NAND2 (N11484, N11483, N1864);
not NOT1 (N11485, N11480);
nand NAND3 (N11486, N11469, N2517, N5963);
nor NOR2 (N11487, N11485, N7923);
xor XOR2 (N11488, N11476, N6787);
or OR3 (N11489, N11488, N3310, N10260);
nand NAND4 (N11490, N11467, N2223, N6031, N4328);
nand NAND3 (N11491, N11489, N3163, N3085);
not NOT1 (N11492, N11479);
and AND4 (N11493, N11472, N10394, N9481, N1105);
nor NOR4 (N11494, N11490, N8725, N10556, N39);
and AND3 (N11495, N11487, N3027, N11071);
or OR4 (N11496, N11474, N11332, N8282, N1369);
and AND4 (N11497, N11486, N5732, N8631, N5160);
nor NOR4 (N11498, N11477, N6033, N2744, N10148);
or OR2 (N11499, N11491, N4724);
nor NOR3 (N11500, N11499, N8353, N6733);
nand NAND2 (N11501, N11496, N10735);
xor XOR2 (N11502, N11482, N9106);
nand NAND2 (N11503, N11494, N2975);
nor NOR2 (N11504, N11495, N9728);
and AND2 (N11505, N11493, N1261);
not NOT1 (N11506, N11505);
buf BUF1 (N11507, N11484);
nand NAND3 (N11508, N11506, N1620, N3636);
xor XOR2 (N11509, N11497, N9997);
nand NAND3 (N11510, N11502, N5589, N4526);
xor XOR2 (N11511, N11498, N10286);
xor XOR2 (N11512, N11504, N409);
nor NOR2 (N11513, N11507, N3740);
and AND2 (N11514, N11508, N9335);
nor NOR4 (N11515, N11512, N9594, N5970, N3143);
not NOT1 (N11516, N11513);
nand NAND3 (N11517, N11514, N10024, N6514);
xor XOR2 (N11518, N11509, N2169);
and AND3 (N11519, N11503, N1646, N10523);
nand NAND4 (N11520, N11518, N2163, N10656, N2056);
nor NOR2 (N11521, N11492, N10001);
xor XOR2 (N11522, N11517, N4037);
not NOT1 (N11523, N11515);
nand NAND4 (N11524, N11521, N153, N4406, N4894);
xor XOR2 (N11525, N11511, N2028);
nand NAND3 (N11526, N11500, N2569, N7630);
xor XOR2 (N11527, N11526, N1294);
and AND3 (N11528, N11501, N3799, N7402);
and AND2 (N11529, N11519, N1713);
xor XOR2 (N11530, N11510, N259);
or OR4 (N11531, N11516, N6971, N7297, N212);
nand NAND2 (N11532, N11531, N1624);
or OR2 (N11533, N11529, N6016);
or OR4 (N11534, N11520, N2228, N352, N1724);
xor XOR2 (N11535, N11522, N4340);
xor XOR2 (N11536, N11528, N7133);
not NOT1 (N11537, N11534);
buf BUF1 (N11538, N11537);
or OR4 (N11539, N11524, N10447, N10170, N6971);
nor NOR3 (N11540, N11539, N7623, N5519);
and AND2 (N11541, N11525, N7923);
nand NAND2 (N11542, N11538, N10527);
or OR2 (N11543, N11535, N4423);
buf BUF1 (N11544, N11523);
or OR2 (N11545, N11543, N2886);
xor XOR2 (N11546, N11542, N10216);
and AND3 (N11547, N11536, N7888, N5153);
not NOT1 (N11548, N11544);
xor XOR2 (N11549, N11527, N8246);
nor NOR2 (N11550, N11530, N2714);
nand NAND4 (N11551, N11545, N7152, N751, N4363);
xor XOR2 (N11552, N11540, N5757);
not NOT1 (N11553, N11533);
not NOT1 (N11554, N11546);
or OR4 (N11555, N11551, N11232, N446, N3393);
or OR4 (N11556, N11541, N6751, N9190, N4814);
xor XOR2 (N11557, N11550, N2030);
and AND2 (N11558, N11554, N10083);
and AND2 (N11559, N11558, N7267);
not NOT1 (N11560, N11559);
nor NOR2 (N11561, N11549, N1514);
not NOT1 (N11562, N11532);
nor NOR4 (N11563, N11553, N10774, N3293, N10721);
buf BUF1 (N11564, N11563);
or OR2 (N11565, N11552, N7728);
nand NAND3 (N11566, N11548, N3478, N10924);
xor XOR2 (N11567, N11561, N6665);
nand NAND3 (N11568, N11556, N2507, N2335);
not NOT1 (N11569, N11562);
nor NOR3 (N11570, N11547, N9046, N4305);
nand NAND2 (N11571, N11568, N8963);
or OR2 (N11572, N11560, N3205);
nor NOR3 (N11573, N11571, N4720, N4685);
nand NAND2 (N11574, N11573, N3379);
nor NOR2 (N11575, N11555, N3350);
buf BUF1 (N11576, N11567);
buf BUF1 (N11577, N11575);
buf BUF1 (N11578, N11566);
xor XOR2 (N11579, N11569, N9426);
not NOT1 (N11580, N11574);
not NOT1 (N11581, N11579);
or OR2 (N11582, N11581, N10486);
not NOT1 (N11583, N11577);
nand NAND2 (N11584, N11578, N52);
not NOT1 (N11585, N11580);
nand NAND4 (N11586, N11585, N11299, N2621, N9894);
nor NOR3 (N11587, N11570, N9742, N3896);
and AND4 (N11588, N11582, N4628, N4947, N7401);
not NOT1 (N11589, N11572);
xor XOR2 (N11590, N11586, N9790);
nor NOR2 (N11591, N11587, N4264);
and AND2 (N11592, N11591, N4994);
not NOT1 (N11593, N11557);
nor NOR2 (N11594, N11592, N2466);
buf BUF1 (N11595, N11594);
nand NAND3 (N11596, N11583, N266, N11582);
nand NAND3 (N11597, N11565, N9548, N1290);
nor NOR4 (N11598, N11590, N8338, N8040, N3256);
nand NAND2 (N11599, N11595, N6529);
and AND2 (N11600, N11589, N1281);
buf BUF1 (N11601, N11593);
or OR4 (N11602, N11588, N9325, N6077, N3402);
nor NOR2 (N11603, N11597, N5469);
xor XOR2 (N11604, N11602, N3880);
nor NOR3 (N11605, N11598, N2666, N1738);
not NOT1 (N11606, N11604);
xor XOR2 (N11607, N11576, N6238);
nor NOR2 (N11608, N11603, N939);
xor XOR2 (N11609, N11606, N848);
and AND2 (N11610, N11608, N9703);
nor NOR4 (N11611, N11607, N11238, N5970, N10584);
and AND2 (N11612, N11610, N3722);
nor NOR4 (N11613, N11599, N7094, N7204, N9124);
buf BUF1 (N11614, N11612);
nor NOR3 (N11615, N11614, N2889, N11445);
and AND3 (N11616, N11615, N2620, N6846);
nand NAND3 (N11617, N11605, N3424, N5582);
buf BUF1 (N11618, N11584);
or OR2 (N11619, N11611, N4676);
xor XOR2 (N11620, N11619, N4199);
nand NAND2 (N11621, N11609, N3293);
xor XOR2 (N11622, N11600, N2321);
not NOT1 (N11623, N11613);
xor XOR2 (N11624, N11564, N9381);
and AND2 (N11625, N11596, N3079);
not NOT1 (N11626, N11616);
nor NOR4 (N11627, N11621, N8252, N3982, N624);
or OR2 (N11628, N11625, N8346);
buf BUF1 (N11629, N11618);
not NOT1 (N11630, N11624);
or OR4 (N11631, N11620, N9846, N3776, N2001);
or OR3 (N11632, N11601, N2512, N8954);
or OR3 (N11633, N11623, N8797, N4610);
nor NOR4 (N11634, N11630, N1197, N825, N1354);
or OR4 (N11635, N11634, N10567, N6302, N9888);
nor NOR3 (N11636, N11632, N10149, N1533);
not NOT1 (N11637, N11627);
buf BUF1 (N11638, N11617);
and AND2 (N11639, N11636, N937);
and AND2 (N11640, N11628, N9491);
nor NOR3 (N11641, N11622, N3341, N8777);
or OR2 (N11642, N11629, N8085);
xor XOR2 (N11643, N11637, N11504);
or OR4 (N11644, N11635, N8317, N2238, N2890);
nor NOR3 (N11645, N11644, N7848, N8354);
xor XOR2 (N11646, N11639, N11100);
xor XOR2 (N11647, N11646, N6142);
nand NAND2 (N11648, N11640, N8308);
and AND2 (N11649, N11643, N6101);
and AND2 (N11650, N11649, N1530);
xor XOR2 (N11651, N11641, N2557);
nor NOR2 (N11652, N11626, N5662);
not NOT1 (N11653, N11638);
or OR4 (N11654, N11633, N7209, N6714, N580);
and AND3 (N11655, N11651, N8960, N9727);
or OR2 (N11656, N11653, N10745);
and AND2 (N11657, N11655, N2224);
and AND3 (N11658, N11656, N9732, N9407);
buf BUF1 (N11659, N11652);
and AND4 (N11660, N11657, N9235, N2695, N8595);
not NOT1 (N11661, N11660);
xor XOR2 (N11662, N11654, N9969);
and AND2 (N11663, N11647, N10011);
buf BUF1 (N11664, N11642);
nand NAND4 (N11665, N11658, N3639, N340, N5414);
nand NAND4 (N11666, N11645, N5545, N7713, N4115);
xor XOR2 (N11667, N11664, N9442);
or OR4 (N11668, N11659, N3386, N8629, N1019);
xor XOR2 (N11669, N11665, N11375);
not NOT1 (N11670, N11666);
nand NAND2 (N11671, N11631, N622);
or OR3 (N11672, N11671, N5011, N8224);
nand NAND2 (N11673, N11648, N8675);
and AND4 (N11674, N11663, N5794, N2437, N3773);
and AND4 (N11675, N11668, N9785, N8203, N8776);
and AND2 (N11676, N11674, N4981);
xor XOR2 (N11677, N11670, N7033);
buf BUF1 (N11678, N11673);
or OR4 (N11679, N11677, N2028, N6872, N9897);
nor NOR4 (N11680, N11667, N10013, N3990, N11321);
nor NOR3 (N11681, N11669, N3338, N6448);
nand NAND3 (N11682, N11672, N894, N3462);
and AND4 (N11683, N11661, N4846, N5518, N6563);
xor XOR2 (N11684, N11662, N1981);
nor NOR3 (N11685, N11682, N8384, N2855);
and AND2 (N11686, N11684, N10943);
and AND2 (N11687, N11675, N403);
not NOT1 (N11688, N11679);
xor XOR2 (N11689, N11681, N10040);
xor XOR2 (N11690, N11683, N58);
or OR2 (N11691, N11678, N2961);
and AND4 (N11692, N11688, N1618, N3144, N2821);
and AND4 (N11693, N11676, N4487, N9678, N2659);
buf BUF1 (N11694, N11680);
nand NAND4 (N11695, N11693, N11276, N10379, N4574);
nand NAND2 (N11696, N11695, N2619);
or OR3 (N11697, N11696, N7587, N3967);
not NOT1 (N11698, N11697);
buf BUF1 (N11699, N11692);
buf BUF1 (N11700, N11690);
buf BUF1 (N11701, N11689);
nand NAND2 (N11702, N11686, N3522);
or OR2 (N11703, N11691, N11348);
nand NAND2 (N11704, N11687, N11068);
buf BUF1 (N11705, N11701);
xor XOR2 (N11706, N11694, N11646);
and AND4 (N11707, N11706, N4508, N820, N11691);
nand NAND4 (N11708, N11707, N10435, N6437, N9136);
xor XOR2 (N11709, N11702, N5737);
or OR2 (N11710, N11650, N831);
xor XOR2 (N11711, N11703, N3369);
nand NAND4 (N11712, N11711, N1258, N11309, N5555);
and AND2 (N11713, N11710, N11320);
nand NAND4 (N11714, N11708, N5592, N3526, N9658);
buf BUF1 (N11715, N11714);
not NOT1 (N11716, N11700);
xor XOR2 (N11717, N11712, N7675);
and AND4 (N11718, N11715, N8953, N5919, N7071);
and AND2 (N11719, N11698, N6755);
and AND3 (N11720, N11699, N9548, N11114);
or OR4 (N11721, N11720, N5536, N3824, N3649);
buf BUF1 (N11722, N11721);
nor NOR4 (N11723, N11705, N4027, N8686, N10305);
and AND2 (N11724, N11713, N9854);
nand NAND4 (N11725, N11704, N6124, N279, N6514);
and AND2 (N11726, N11725, N7219);
nand NAND4 (N11727, N11723, N8116, N4914, N4389);
buf BUF1 (N11728, N11718);
xor XOR2 (N11729, N11717, N10250);
and AND3 (N11730, N11716, N10667, N5135);
buf BUF1 (N11731, N11722);
and AND4 (N11732, N11728, N412, N6256, N6694);
xor XOR2 (N11733, N11726, N8330);
xor XOR2 (N11734, N11724, N4967);
xor XOR2 (N11735, N11734, N8485);
nand NAND4 (N11736, N11733, N10879, N10820, N3140);
buf BUF1 (N11737, N11709);
xor XOR2 (N11738, N11727, N8923);
and AND3 (N11739, N11729, N685, N69);
not NOT1 (N11740, N11731);
or OR4 (N11741, N11736, N10134, N8211, N8131);
or OR4 (N11742, N11685, N3183, N5491, N3817);
not NOT1 (N11743, N11741);
not NOT1 (N11744, N11739);
and AND4 (N11745, N11738, N5189, N8379, N5135);
buf BUF1 (N11746, N11730);
xor XOR2 (N11747, N11746, N5792);
or OR3 (N11748, N11719, N8963, N3742);
buf BUF1 (N11749, N11743);
nor NOR2 (N11750, N11749, N10442);
buf BUF1 (N11751, N11735);
nor NOR4 (N11752, N11732, N1969, N11201, N5052);
or OR2 (N11753, N11742, N8852);
not NOT1 (N11754, N11737);
nor NOR3 (N11755, N11745, N11354, N1354);
or OR4 (N11756, N11755, N4489, N7933, N6916);
xor XOR2 (N11757, N11747, N2897);
or OR3 (N11758, N11751, N3470, N11083);
not NOT1 (N11759, N11752);
nor NOR2 (N11760, N11758, N4301);
buf BUF1 (N11761, N11753);
and AND2 (N11762, N11761, N6655);
buf BUF1 (N11763, N11748);
xor XOR2 (N11764, N11750, N8852);
not NOT1 (N11765, N11763);
buf BUF1 (N11766, N11759);
xor XOR2 (N11767, N11744, N2933);
nor NOR4 (N11768, N11757, N7719, N11658, N2163);
nor NOR2 (N11769, N11760, N3254);
not NOT1 (N11770, N11767);
xor XOR2 (N11771, N11768, N6412);
or OR4 (N11772, N11756, N7612, N1575, N9076);
nor NOR3 (N11773, N11740, N9233, N2331);
not NOT1 (N11774, N11762);
nor NOR3 (N11775, N11771, N11414, N3679);
and AND3 (N11776, N11772, N10937, N7863);
not NOT1 (N11777, N11754);
xor XOR2 (N11778, N11770, N10593);
or OR2 (N11779, N11765, N4378);
not NOT1 (N11780, N11778);
buf BUF1 (N11781, N11769);
xor XOR2 (N11782, N11764, N11465);
buf BUF1 (N11783, N11782);
not NOT1 (N11784, N11776);
and AND4 (N11785, N11779, N8441, N4894, N7389);
not NOT1 (N11786, N11773);
or OR4 (N11787, N11777, N2075, N4444, N4522);
nor NOR4 (N11788, N11775, N5711, N9973, N8550);
nor NOR3 (N11789, N11787, N2199, N10544);
not NOT1 (N11790, N11766);
or OR2 (N11791, N11789, N8977);
buf BUF1 (N11792, N11791);
nand NAND4 (N11793, N11783, N2537, N10604, N7898);
and AND3 (N11794, N11792, N4519, N4454);
nor NOR4 (N11795, N11784, N4928, N1569, N4849);
nand NAND2 (N11796, N11781, N9999);
and AND4 (N11797, N11790, N596, N7385, N4580);
xor XOR2 (N11798, N11794, N1402);
nor NOR2 (N11799, N11796, N5778);
not NOT1 (N11800, N11797);
or OR2 (N11801, N11786, N2445);
or OR2 (N11802, N11798, N9921);
nand NAND4 (N11803, N11801, N5819, N3834, N11691);
and AND2 (N11804, N11788, N6993);
nand NAND4 (N11805, N11804, N1150, N8866, N5705);
buf BUF1 (N11806, N11793);
nor NOR3 (N11807, N11805, N5660, N1135);
buf BUF1 (N11808, N11807);
and AND2 (N11809, N11785, N7718);
not NOT1 (N11810, N11774);
nor NOR4 (N11811, N11808, N5064, N9149, N6024);
nand NAND3 (N11812, N11811, N8957, N1486);
xor XOR2 (N11813, N11780, N9520);
nand NAND2 (N11814, N11812, N10920);
or OR4 (N11815, N11813, N9810, N11123, N5584);
xor XOR2 (N11816, N11803, N7393);
nand NAND3 (N11817, N11810, N353, N2267);
nor NOR3 (N11818, N11800, N4327, N8572);
buf BUF1 (N11819, N11799);
nor NOR3 (N11820, N11816, N7560, N11453);
buf BUF1 (N11821, N11814);
nand NAND2 (N11822, N11820, N5226);
and AND2 (N11823, N11809, N35);
xor XOR2 (N11824, N11818, N8444);
xor XOR2 (N11825, N11817, N9474);
nand NAND2 (N11826, N11823, N10138);
and AND3 (N11827, N11825, N2788, N1092);
nor NOR2 (N11828, N11795, N7732);
or OR3 (N11829, N11819, N3669, N7875);
and AND3 (N11830, N11829, N5776, N8083);
not NOT1 (N11831, N11822);
or OR4 (N11832, N11828, N1887, N1434, N9235);
buf BUF1 (N11833, N11824);
or OR3 (N11834, N11815, N8459, N6574);
buf BUF1 (N11835, N11833);
buf BUF1 (N11836, N11826);
buf BUF1 (N11837, N11835);
or OR3 (N11838, N11836, N9694, N8605);
not NOT1 (N11839, N11806);
buf BUF1 (N11840, N11839);
xor XOR2 (N11841, N11802, N3575);
or OR3 (N11842, N11834, N3953, N3067);
nand NAND3 (N11843, N11841, N3946, N1644);
xor XOR2 (N11844, N11831, N574);
not NOT1 (N11845, N11827);
nor NOR3 (N11846, N11845, N2847, N11559);
buf BUF1 (N11847, N11821);
not NOT1 (N11848, N11832);
xor XOR2 (N11849, N11830, N5040);
nand NAND4 (N11850, N11842, N10490, N4096, N8577);
buf BUF1 (N11851, N11846);
and AND4 (N11852, N11847, N1714, N8569, N8652);
xor XOR2 (N11853, N11851, N10925);
or OR4 (N11854, N11837, N3531, N7853, N725);
and AND2 (N11855, N11848, N4919);
buf BUF1 (N11856, N11840);
and AND3 (N11857, N11853, N9281, N8127);
nand NAND4 (N11858, N11843, N8638, N6027, N8657);
not NOT1 (N11859, N11844);
or OR2 (N11860, N11849, N7109);
or OR3 (N11861, N11854, N6504, N7869);
or OR3 (N11862, N11856, N8017, N11814);
not NOT1 (N11863, N11858);
or OR3 (N11864, N11862, N661, N3242);
nand NAND4 (N11865, N11863, N9217, N10915, N5318);
nand NAND2 (N11866, N11865, N4512);
buf BUF1 (N11867, N11864);
not NOT1 (N11868, N11861);
xor XOR2 (N11869, N11860, N1734);
buf BUF1 (N11870, N11859);
xor XOR2 (N11871, N11866, N8560);
xor XOR2 (N11872, N11869, N6607);
buf BUF1 (N11873, N11838);
buf BUF1 (N11874, N11868);
or OR2 (N11875, N11857, N11493);
nor NOR2 (N11876, N11852, N9798);
not NOT1 (N11877, N11867);
or OR2 (N11878, N11870, N6116);
buf BUF1 (N11879, N11877);
or OR3 (N11880, N11879, N11606, N8735);
or OR4 (N11881, N11855, N9524, N11595, N10517);
and AND2 (N11882, N11876, N6285);
and AND3 (N11883, N11881, N5037, N1701);
or OR4 (N11884, N11850, N10700, N8417, N11012);
not NOT1 (N11885, N11880);
xor XOR2 (N11886, N11878, N335);
or OR4 (N11887, N11871, N1620, N7995, N11836);
and AND2 (N11888, N11884, N298);
and AND3 (N11889, N11887, N1422, N5674);
or OR2 (N11890, N11882, N2179);
buf BUF1 (N11891, N11890);
nand NAND4 (N11892, N11885, N2691, N5588, N9444);
xor XOR2 (N11893, N11872, N9437);
nor NOR4 (N11894, N11889, N800, N4708, N6431);
buf BUF1 (N11895, N11894);
not NOT1 (N11896, N11875);
nand NAND2 (N11897, N11892, N9779);
and AND3 (N11898, N11888, N6390, N10889);
and AND2 (N11899, N11893, N10931);
or OR2 (N11900, N11895, N5425);
buf BUF1 (N11901, N11874);
nor NOR4 (N11902, N11900, N2730, N6639, N5516);
and AND3 (N11903, N11896, N4426, N11257);
nand NAND4 (N11904, N11902, N5311, N6131, N3790);
and AND4 (N11905, N11873, N8837, N2130, N9922);
and AND4 (N11906, N11886, N9037, N8542, N3299);
and AND3 (N11907, N11904, N3232, N7792);
not NOT1 (N11908, N11883);
not NOT1 (N11909, N11899);
buf BUF1 (N11910, N11897);
and AND2 (N11911, N11903, N7274);
or OR3 (N11912, N11906, N265, N5334);
xor XOR2 (N11913, N11910, N7857);
and AND4 (N11914, N11898, N7822, N6340, N6283);
xor XOR2 (N11915, N11901, N6982);
buf BUF1 (N11916, N11912);
nor NOR4 (N11917, N11914, N7580, N3261, N10252);
xor XOR2 (N11918, N11915, N10263);
nor NOR2 (N11919, N11916, N4753);
or OR3 (N11920, N11909, N5733, N11719);
nor NOR4 (N11921, N11911, N5424, N1075, N11413);
buf BUF1 (N11922, N11905);
nor NOR2 (N11923, N11920, N1327);
or OR2 (N11924, N11891, N8354);
buf BUF1 (N11925, N11908);
or OR4 (N11926, N11921, N6432, N8191, N22);
buf BUF1 (N11927, N11925);
or OR2 (N11928, N11918, N10432);
nand NAND4 (N11929, N11924, N10269, N6623, N2226);
nand NAND4 (N11930, N11919, N9232, N4507, N1976);
xor XOR2 (N11931, N11907, N8744);
or OR3 (N11932, N11926, N3400, N9425);
and AND3 (N11933, N11928, N2503, N514);
or OR4 (N11934, N11923, N6509, N1490, N9287);
buf BUF1 (N11935, N11930);
xor XOR2 (N11936, N11931, N4468);
buf BUF1 (N11937, N11933);
not NOT1 (N11938, N11913);
nor NOR2 (N11939, N11937, N3341);
and AND2 (N11940, N11938, N7728);
and AND2 (N11941, N11939, N7223);
buf BUF1 (N11942, N11941);
nand NAND3 (N11943, N11917, N9078, N11633);
and AND3 (N11944, N11934, N3514, N2464);
or OR4 (N11945, N11936, N3064, N3866, N8450);
and AND3 (N11946, N11945, N4798, N1187);
not NOT1 (N11947, N11944);
nand NAND4 (N11948, N11946, N6650, N7200, N5035);
nand NAND2 (N11949, N11948, N7787);
nand NAND4 (N11950, N11947, N6078, N6146, N9482);
not NOT1 (N11951, N11929);
nor NOR3 (N11952, N11940, N1685, N1618);
buf BUF1 (N11953, N11922);
or OR3 (N11954, N11932, N3063, N985);
buf BUF1 (N11955, N11949);
nand NAND4 (N11956, N11943, N3297, N1731, N6039);
nor NOR2 (N11957, N11951, N6277);
nand NAND4 (N11958, N11956, N11252, N2588, N5583);
or OR2 (N11959, N11950, N7188);
buf BUF1 (N11960, N11942);
nand NAND2 (N11961, N11952, N9974);
nand NAND4 (N11962, N11957, N8483, N6164, N6518);
nand NAND3 (N11963, N11954, N11785, N5476);
and AND3 (N11964, N11961, N7245, N2516);
xor XOR2 (N11965, N11962, N1677);
or OR2 (N11966, N11963, N2574);
xor XOR2 (N11967, N11935, N4219);
nand NAND4 (N11968, N11958, N3686, N10132, N4209);
buf BUF1 (N11969, N11960);
or OR2 (N11970, N11964, N11518);
buf BUF1 (N11971, N11965);
or OR4 (N11972, N11955, N11942, N9669, N1736);
not NOT1 (N11973, N11967);
and AND3 (N11974, N11959, N1025, N4970);
xor XOR2 (N11975, N11973, N5671);
nor NOR4 (N11976, N11971, N7025, N9062, N10337);
not NOT1 (N11977, N11966);
not NOT1 (N11978, N11968);
xor XOR2 (N11979, N11953, N98);
and AND4 (N11980, N11976, N38, N6834, N11492);
and AND3 (N11981, N11970, N11497, N7816);
not NOT1 (N11982, N11969);
xor XOR2 (N11983, N11981, N876);
not NOT1 (N11984, N11975);
buf BUF1 (N11985, N11979);
and AND4 (N11986, N11972, N6398, N626, N10839);
xor XOR2 (N11987, N11983, N5422);
nand NAND3 (N11988, N11977, N1341, N7986);
nor NOR3 (N11989, N11980, N11795, N141);
or OR4 (N11990, N11989, N6578, N9037, N1561);
nor NOR2 (N11991, N11984, N1);
or OR2 (N11992, N11974, N4725);
buf BUF1 (N11993, N11986);
xor XOR2 (N11994, N11927, N1707);
nand NAND4 (N11995, N11993, N2976, N7048, N10540);
and AND4 (N11996, N11978, N8341, N8107, N4575);
and AND2 (N11997, N11994, N6682);
not NOT1 (N11998, N11996);
or OR2 (N11999, N11985, N5940);
buf BUF1 (N12000, N11999);
not NOT1 (N12001, N11988);
xor XOR2 (N12002, N11991, N9075);
buf BUF1 (N12003, N12002);
or OR2 (N12004, N11995, N8290);
buf BUF1 (N12005, N11998);
and AND2 (N12006, N12001, N6969);
xor XOR2 (N12007, N11997, N11495);
xor XOR2 (N12008, N11990, N8696);
buf BUF1 (N12009, N12005);
buf BUF1 (N12010, N12000);
buf BUF1 (N12011, N11992);
nor NOR2 (N12012, N11982, N3911);
not NOT1 (N12013, N12012);
not NOT1 (N12014, N12007);
nor NOR2 (N12015, N12003, N9541);
and AND2 (N12016, N12011, N4857);
not NOT1 (N12017, N12014);
buf BUF1 (N12018, N12009);
nor NOR2 (N12019, N12008, N10015);
nor NOR4 (N12020, N12019, N10216, N2694, N8280);
nand NAND3 (N12021, N12013, N8532, N11478);
or OR4 (N12022, N12010, N6508, N1607, N8421);
and AND2 (N12023, N12017, N7594);
xor XOR2 (N12024, N12016, N1397);
buf BUF1 (N12025, N11987);
or OR4 (N12026, N12023, N7292, N627, N4493);
buf BUF1 (N12027, N12026);
xor XOR2 (N12028, N12027, N9553);
nand NAND4 (N12029, N12004, N10733, N10407, N1973);
or OR3 (N12030, N12020, N1525, N2687);
or OR3 (N12031, N12024, N9341, N1392);
and AND2 (N12032, N12021, N7614);
nand NAND4 (N12033, N12006, N2634, N8049, N6771);
or OR3 (N12034, N12033, N8433, N1926);
nor NOR4 (N12035, N12034, N11717, N7118, N237);
or OR2 (N12036, N12031, N4557);
nand NAND2 (N12037, N12035, N486);
and AND2 (N12038, N12037, N5146);
xor XOR2 (N12039, N12028, N11005);
and AND4 (N12040, N12022, N6294, N8757, N9160);
and AND3 (N12041, N12036, N2776, N4387);
xor XOR2 (N12042, N12040, N8572);
xor XOR2 (N12043, N12018, N2957);
not NOT1 (N12044, N12041);
buf BUF1 (N12045, N12042);
or OR2 (N12046, N12045, N932);
nand NAND2 (N12047, N12038, N9632);
or OR2 (N12048, N12015, N3155);
buf BUF1 (N12049, N12048);
or OR3 (N12050, N12043, N10556, N3417);
nor NOR4 (N12051, N12032, N1823, N6718, N840);
nand NAND2 (N12052, N12025, N6957);
buf BUF1 (N12053, N12047);
and AND2 (N12054, N12049, N5627);
not NOT1 (N12055, N12044);
not NOT1 (N12056, N12050);
nand NAND4 (N12057, N12054, N3060, N3582, N9483);
nor NOR2 (N12058, N12057, N4931);
or OR3 (N12059, N12055, N8966, N554);
or OR4 (N12060, N12058, N8313, N7523, N4159);
buf BUF1 (N12061, N12059);
and AND3 (N12062, N12039, N664, N8837);
nand NAND4 (N12063, N12060, N7412, N4861, N3644);
and AND2 (N12064, N12053, N934);
and AND4 (N12065, N12064, N6833, N11349, N3849);
or OR2 (N12066, N12056, N2501);
buf BUF1 (N12067, N12030);
xor XOR2 (N12068, N12046, N9412);
buf BUF1 (N12069, N12065);
or OR4 (N12070, N12063, N8144, N6623, N3998);
xor XOR2 (N12071, N12062, N7410);
buf BUF1 (N12072, N12029);
not NOT1 (N12073, N12052);
or OR2 (N12074, N12073, N9908);
buf BUF1 (N12075, N12067);
or OR4 (N12076, N12070, N3832, N7410, N2854);
and AND3 (N12077, N12074, N11845, N5692);
buf BUF1 (N12078, N12069);
and AND3 (N12079, N12072, N6267, N5160);
xor XOR2 (N12080, N12078, N5071);
buf BUF1 (N12081, N12071);
buf BUF1 (N12082, N12061);
nor NOR2 (N12083, N12077, N5577);
not NOT1 (N12084, N12066);
or OR4 (N12085, N12075, N6744, N4436, N9656);
xor XOR2 (N12086, N12080, N7315);
nand NAND2 (N12087, N12068, N6476);
and AND2 (N12088, N12083, N330);
or OR4 (N12089, N12084, N11559, N7555, N1547);
nand NAND3 (N12090, N12085, N8353, N8122);
not NOT1 (N12091, N12089);
and AND4 (N12092, N12090, N1886, N930, N8016);
and AND4 (N12093, N12092, N2289, N8798, N529);
xor XOR2 (N12094, N12087, N4585);
nor NOR3 (N12095, N12051, N1558, N8566);
nand NAND2 (N12096, N12086, N6304);
nand NAND2 (N12097, N12079, N11922);
and AND4 (N12098, N12095, N3538, N10454, N7129);
nand NAND4 (N12099, N12094, N4218, N1099, N11473);
or OR4 (N12100, N12097, N10676, N4746, N3532);
buf BUF1 (N12101, N12091);
buf BUF1 (N12102, N12100);
and AND2 (N12103, N12099, N7450);
nand NAND4 (N12104, N12081, N3875, N10746, N10176);
and AND4 (N12105, N12101, N2178, N7558, N4597);
buf BUF1 (N12106, N12104);
xor XOR2 (N12107, N12103, N10097);
nor NOR3 (N12108, N12076, N8204, N3245);
xor XOR2 (N12109, N12106, N5200);
and AND2 (N12110, N12096, N6592);
not NOT1 (N12111, N12109);
buf BUF1 (N12112, N12105);
buf BUF1 (N12113, N12082);
or OR2 (N12114, N12088, N10791);
xor XOR2 (N12115, N12113, N11781);
and AND3 (N12116, N12115, N6315, N11113);
nor NOR2 (N12117, N12098, N6104);
not NOT1 (N12118, N12114);
nor NOR3 (N12119, N12110, N3720, N10673);
not NOT1 (N12120, N12108);
nor NOR4 (N12121, N12111, N8329, N9942, N2905);
or OR3 (N12122, N12112, N9058, N5775);
or OR2 (N12123, N12121, N10605);
not NOT1 (N12124, N12118);
not NOT1 (N12125, N12122);
nand NAND2 (N12126, N12119, N5232);
nand NAND2 (N12127, N12116, N1672);
not NOT1 (N12128, N12117);
buf BUF1 (N12129, N12102);
nor NOR3 (N12130, N12127, N7500, N449);
not NOT1 (N12131, N12093);
nor NOR4 (N12132, N12123, N2210, N4621, N9217);
and AND2 (N12133, N12124, N5705);
buf BUF1 (N12134, N12133);
buf BUF1 (N12135, N12120);
not NOT1 (N12136, N12130);
and AND3 (N12137, N12129, N6759, N6711);
or OR3 (N12138, N12126, N3876, N8530);
nor NOR2 (N12139, N12128, N433);
and AND2 (N12140, N12135, N11764);
or OR4 (N12141, N12107, N8102, N1733, N8704);
nor NOR3 (N12142, N12141, N1195, N3432);
buf BUF1 (N12143, N12139);
or OR3 (N12144, N12132, N8708, N10078);
nor NOR2 (N12145, N12140, N12138);
nor NOR2 (N12146, N9513, N5693);
or OR3 (N12147, N12144, N1611, N6513);
and AND2 (N12148, N12146, N2543);
or OR3 (N12149, N12145, N11165, N3217);
nand NAND4 (N12150, N12148, N3218, N9027, N11854);
not NOT1 (N12151, N12149);
buf BUF1 (N12152, N12151);
buf BUF1 (N12153, N12142);
nor NOR3 (N12154, N12147, N226, N656);
or OR3 (N12155, N12125, N3841, N1165);
or OR3 (N12156, N12154, N5405, N5246);
and AND2 (N12157, N12153, N3961);
and AND4 (N12158, N12137, N4569, N1370, N11743);
nor NOR2 (N12159, N12158, N10166);
and AND3 (N12160, N12152, N2122, N7005);
nand NAND4 (N12161, N12155, N6645, N7443, N10269);
nand NAND2 (N12162, N12161, N819);
nand NAND4 (N12163, N12159, N1239, N2386, N11890);
nor NOR2 (N12164, N12163, N1220);
nand NAND3 (N12165, N12131, N4590, N6602);
nor NOR3 (N12166, N12136, N1141, N6464);
not NOT1 (N12167, N12162);
not NOT1 (N12168, N12165);
or OR3 (N12169, N12166, N10940, N6736);
buf BUF1 (N12170, N12156);
not NOT1 (N12171, N12167);
and AND2 (N12172, N12168, N10109);
or OR4 (N12173, N12134, N5537, N2207, N5465);
nor NOR2 (N12174, N12169, N2568);
and AND2 (N12175, N12173, N1081);
nor NOR2 (N12176, N12171, N11900);
nor NOR2 (N12177, N12174, N2029);
or OR2 (N12178, N12170, N5597);
xor XOR2 (N12179, N12150, N169);
buf BUF1 (N12180, N12175);
not NOT1 (N12181, N12172);
nor NOR3 (N12182, N12181, N3398, N937);
or OR3 (N12183, N12177, N7870, N6516);
or OR4 (N12184, N12176, N5895, N9781, N10315);
buf BUF1 (N12185, N12143);
buf BUF1 (N12186, N12185);
or OR4 (N12187, N12186, N10452, N1827, N7223);
not NOT1 (N12188, N12182);
and AND4 (N12189, N12187, N3510, N7017, N4510);
buf BUF1 (N12190, N12180);
nand NAND2 (N12191, N12189, N422);
not NOT1 (N12192, N12179);
xor XOR2 (N12193, N12157, N11407);
nor NOR4 (N12194, N12192, N10586, N10131, N2519);
and AND4 (N12195, N12194, N11890, N9283, N2258);
and AND4 (N12196, N12188, N1107, N10177, N7818);
or OR4 (N12197, N12193, N6235, N10314, N3900);
or OR4 (N12198, N12184, N9779, N569, N5550);
or OR4 (N12199, N12196, N4360, N2246, N1826);
xor XOR2 (N12200, N12197, N5624);
or OR3 (N12201, N12199, N10719, N7917);
not NOT1 (N12202, N12164);
nor NOR4 (N12203, N12202, N8929, N11421, N9709);
and AND3 (N12204, N12200, N6273, N12125);
nand NAND2 (N12205, N12160, N9128);
and AND4 (N12206, N12198, N287, N5246, N3646);
nand NAND4 (N12207, N12205, N3921, N9907, N11720);
xor XOR2 (N12208, N12201, N5750);
and AND2 (N12209, N12190, N7309);
xor XOR2 (N12210, N12208, N8469);
nor NOR4 (N12211, N12183, N7171, N9828, N2278);
xor XOR2 (N12212, N12203, N1501);
and AND3 (N12213, N12209, N975, N11217);
buf BUF1 (N12214, N12195);
nand NAND4 (N12215, N12178, N3445, N3827, N1342);
buf BUF1 (N12216, N12215);
nand NAND2 (N12217, N12206, N10604);
or OR4 (N12218, N12204, N9517, N3970, N1336);
nand NAND3 (N12219, N12191, N7978, N3081);
or OR4 (N12220, N12218, N3295, N7622, N537);
xor XOR2 (N12221, N12207, N10870);
or OR3 (N12222, N12214, N2573, N5637);
nor NOR3 (N12223, N12216, N8490, N9591);
xor XOR2 (N12224, N12211, N4829);
and AND2 (N12225, N12220, N10777);
and AND2 (N12226, N12221, N1026);
not NOT1 (N12227, N12217);
or OR3 (N12228, N12224, N6628, N9599);
or OR4 (N12229, N12225, N6032, N5374, N5765);
buf BUF1 (N12230, N12223);
not NOT1 (N12231, N12227);
buf BUF1 (N12232, N12222);
and AND4 (N12233, N12212, N10806, N10586, N10164);
xor XOR2 (N12234, N12213, N9261);
nand NAND3 (N12235, N12231, N4596, N4355);
xor XOR2 (N12236, N12229, N2261);
not NOT1 (N12237, N12234);
nand NAND2 (N12238, N12233, N4511);
not NOT1 (N12239, N12226);
or OR3 (N12240, N12210, N566, N1893);
not NOT1 (N12241, N12230);
nand NAND4 (N12242, N12237, N3855, N8637, N7074);
buf BUF1 (N12243, N12236);
not NOT1 (N12244, N12232);
xor XOR2 (N12245, N12228, N1079);
nor NOR3 (N12246, N12245, N5136, N6006);
nor NOR2 (N12247, N12219, N909);
nand NAND3 (N12248, N12247, N6886, N4045);
nand NAND4 (N12249, N12243, N6239, N7189, N11620);
buf BUF1 (N12250, N12248);
nor NOR2 (N12251, N12238, N11998);
buf BUF1 (N12252, N12239);
xor XOR2 (N12253, N12252, N2115);
and AND2 (N12254, N12251, N9766);
and AND2 (N12255, N12249, N1059);
or OR4 (N12256, N12242, N8260, N3662, N7426);
or OR4 (N12257, N12254, N8450, N9914, N1394);
buf BUF1 (N12258, N12240);
not NOT1 (N12259, N12241);
and AND2 (N12260, N12256, N12239);
buf BUF1 (N12261, N12260);
or OR2 (N12262, N12246, N2471);
and AND2 (N12263, N12235, N326);
and AND3 (N12264, N12258, N7876, N8179);
or OR3 (N12265, N12259, N4874, N11888);
nand NAND4 (N12266, N12261, N2624, N11760, N414);
nand NAND3 (N12267, N12263, N11422, N6299);
nand NAND3 (N12268, N12265, N8085, N1795);
xor XOR2 (N12269, N12257, N11722);
not NOT1 (N12270, N12253);
not NOT1 (N12271, N12268);
nor NOR3 (N12272, N12244, N7790, N4195);
nand NAND4 (N12273, N12264, N11977, N4463, N7689);
and AND3 (N12274, N12262, N80, N8239);
xor XOR2 (N12275, N12267, N7035);
nor NOR2 (N12276, N12274, N8145);
nor NOR3 (N12277, N12269, N8216, N10627);
nor NOR2 (N12278, N12277, N821);
and AND3 (N12279, N12276, N2981, N12244);
xor XOR2 (N12280, N12255, N4683);
or OR3 (N12281, N12279, N11183, N10819);
nor NOR4 (N12282, N12266, N8661, N3681, N6068);
and AND3 (N12283, N12278, N9362, N1726);
nand NAND2 (N12284, N12280, N4381);
not NOT1 (N12285, N12270);
buf BUF1 (N12286, N12285);
or OR2 (N12287, N12275, N9362);
nor NOR3 (N12288, N12271, N2118, N10109);
nor NOR2 (N12289, N12286, N350);
buf BUF1 (N12290, N12284);
not NOT1 (N12291, N12250);
nand NAND3 (N12292, N12272, N357, N11094);
xor XOR2 (N12293, N12288, N7193);
or OR2 (N12294, N12287, N4425);
xor XOR2 (N12295, N12289, N1047);
and AND4 (N12296, N12281, N2420, N8697, N4116);
not NOT1 (N12297, N12290);
not NOT1 (N12298, N12291);
buf BUF1 (N12299, N12283);
not NOT1 (N12300, N12273);
xor XOR2 (N12301, N12296, N3379);
buf BUF1 (N12302, N12294);
buf BUF1 (N12303, N12297);
buf BUF1 (N12304, N12302);
and AND2 (N12305, N12301, N6064);
nor NOR4 (N12306, N12299, N1658, N6885, N529);
xor XOR2 (N12307, N12303, N7604);
not NOT1 (N12308, N12292);
and AND2 (N12309, N12308, N3796);
nand NAND3 (N12310, N12298, N1734, N10706);
nand NAND4 (N12311, N12300, N2955, N8300, N10129);
not NOT1 (N12312, N12310);
nor NOR2 (N12313, N12304, N7036);
and AND4 (N12314, N12282, N5777, N9310, N9176);
nand NAND3 (N12315, N12311, N372, N2507);
or OR2 (N12316, N12307, N2226);
xor XOR2 (N12317, N12306, N1597);
or OR4 (N12318, N12314, N5567, N1228, N2388);
xor XOR2 (N12319, N12312, N7858);
nand NAND4 (N12320, N12316, N2917, N1250, N343);
nand NAND3 (N12321, N12309, N4420, N4554);
nand NAND3 (N12322, N12305, N2648, N7074);
not NOT1 (N12323, N12321);
or OR2 (N12324, N12323, N1853);
nor NOR2 (N12325, N12315, N3986);
or OR2 (N12326, N12318, N1673);
nor NOR4 (N12327, N12325, N2177, N3214, N10824);
or OR4 (N12328, N12293, N9178, N2940, N7324);
and AND3 (N12329, N12328, N2780, N10770);
not NOT1 (N12330, N12324);
nand NAND3 (N12331, N12313, N9209, N9748);
and AND3 (N12332, N12319, N11756, N3033);
xor XOR2 (N12333, N12322, N10999);
nand NAND2 (N12334, N12326, N9774);
not NOT1 (N12335, N12332);
and AND3 (N12336, N12327, N5168, N12052);
nor NOR3 (N12337, N12317, N5581, N3668);
nor NOR3 (N12338, N12295, N3304, N8518);
xor XOR2 (N12339, N12320, N1887);
not NOT1 (N12340, N12335);
not NOT1 (N12341, N12331);
buf BUF1 (N12342, N12337);
or OR4 (N12343, N12330, N7991, N5262, N5527);
buf BUF1 (N12344, N12340);
not NOT1 (N12345, N12339);
and AND3 (N12346, N12343, N6690, N4150);
buf BUF1 (N12347, N12336);
xor XOR2 (N12348, N12334, N4120);
nand NAND2 (N12349, N12347, N6265);
nand NAND4 (N12350, N12338, N2261, N11617, N7190);
nor NOR3 (N12351, N12344, N4885, N9066);
and AND3 (N12352, N12348, N4808, N6661);
xor XOR2 (N12353, N12346, N683);
not NOT1 (N12354, N12350);
not NOT1 (N12355, N12341);
and AND4 (N12356, N12333, N991, N9717, N8985);
xor XOR2 (N12357, N12353, N890);
nor NOR4 (N12358, N12342, N5743, N2901, N6196);
buf BUF1 (N12359, N12354);
xor XOR2 (N12360, N12351, N8051);
xor XOR2 (N12361, N12352, N223);
or OR3 (N12362, N12329, N11230, N4192);
nor NOR3 (N12363, N12356, N9853, N2232);
or OR3 (N12364, N12358, N4765, N7468);
nand NAND2 (N12365, N12361, N6743);
nor NOR4 (N12366, N12365, N10507, N1117, N20);
nor NOR3 (N12367, N12357, N2352, N291);
or OR2 (N12368, N12360, N11125);
or OR4 (N12369, N12363, N9913, N8261, N9433);
nand NAND2 (N12370, N12355, N8324);
nand NAND2 (N12371, N12369, N2407);
not NOT1 (N12372, N12368);
nor NOR2 (N12373, N12364, N320);
nor NOR3 (N12374, N12372, N6705, N11329);
or OR4 (N12375, N12370, N152, N4383, N8503);
or OR4 (N12376, N12349, N10690, N10369, N9115);
buf BUF1 (N12377, N12373);
not NOT1 (N12378, N12362);
nor NOR3 (N12379, N12378, N1025, N11122);
nand NAND2 (N12380, N12367, N6910);
or OR4 (N12381, N12376, N439, N156, N3189);
nor NOR2 (N12382, N12366, N10360);
and AND3 (N12383, N12380, N8083, N5568);
or OR4 (N12384, N12377, N8251, N1087, N5751);
and AND4 (N12385, N12345, N5405, N8033, N10773);
buf BUF1 (N12386, N12381);
xor XOR2 (N12387, N12375, N5171);
or OR3 (N12388, N12379, N10869, N2930);
nand NAND3 (N12389, N12383, N12028, N8793);
nor NOR2 (N12390, N12374, N11192);
nand NAND2 (N12391, N12388, N6783);
buf BUF1 (N12392, N12386);
nand NAND3 (N12393, N12387, N7698, N7705);
or OR4 (N12394, N12391, N7293, N4330, N12336);
nand NAND2 (N12395, N12390, N2895);
buf BUF1 (N12396, N12371);
or OR2 (N12397, N12389, N6105);
not NOT1 (N12398, N12385);
nor NOR3 (N12399, N12359, N3907, N12030);
and AND4 (N12400, N12384, N1407, N2006, N2680);
or OR4 (N12401, N12400, N11574, N9384, N10852);
nor NOR4 (N12402, N12394, N5847, N699, N6997);
xor XOR2 (N12403, N12393, N9039);
not NOT1 (N12404, N12399);
and AND2 (N12405, N12392, N11810);
xor XOR2 (N12406, N12401, N12022);
or OR4 (N12407, N12398, N11769, N7486, N9705);
buf BUF1 (N12408, N12395);
or OR2 (N12409, N12397, N1816);
not NOT1 (N12410, N12404);
and AND4 (N12411, N12405, N1567, N1054, N5654);
nor NOR3 (N12412, N12402, N173, N3057);
or OR3 (N12413, N12382, N1100, N4746);
or OR2 (N12414, N12408, N6375);
nor NOR4 (N12415, N12413, N5048, N8128, N12118);
or OR2 (N12416, N12412, N2402);
nor NOR4 (N12417, N12409, N482, N10725, N6796);
and AND2 (N12418, N12410, N6482);
and AND4 (N12419, N12396, N2927, N10201, N2735);
xor XOR2 (N12420, N12416, N6030);
nand NAND4 (N12421, N12403, N7919, N11727, N4277);
and AND4 (N12422, N12411, N5461, N5887, N5942);
or OR2 (N12423, N12419, N195);
nor NOR4 (N12424, N12417, N7857, N4886, N3910);
buf BUF1 (N12425, N12420);
xor XOR2 (N12426, N12423, N9504);
or OR2 (N12427, N12421, N11209);
and AND4 (N12428, N12415, N6252, N8765, N5776);
xor XOR2 (N12429, N12427, N9153);
or OR3 (N12430, N12418, N10561, N7166);
and AND2 (N12431, N12428, N8317);
not NOT1 (N12432, N12430);
nand NAND4 (N12433, N12407, N10576, N4744, N1514);
and AND3 (N12434, N12406, N7177, N7552);
and AND4 (N12435, N12431, N3263, N11373, N9134);
not NOT1 (N12436, N12433);
and AND3 (N12437, N12414, N11445, N526);
not NOT1 (N12438, N12422);
nor NOR2 (N12439, N12432, N4083);
nor NOR4 (N12440, N12429, N812, N9669, N1139);
xor XOR2 (N12441, N12436, N3684);
or OR2 (N12442, N12439, N891);
buf BUF1 (N12443, N12437);
or OR2 (N12444, N12435, N1143);
and AND3 (N12445, N12444, N1937, N8512);
nand NAND3 (N12446, N12424, N7257, N9163);
xor XOR2 (N12447, N12441, N6368);
or OR4 (N12448, N12447, N12028, N11807, N6362);
or OR4 (N12449, N12442, N2921, N2094, N6516);
not NOT1 (N12450, N12443);
or OR3 (N12451, N12434, N8188, N11623);
or OR2 (N12452, N12445, N4292);
or OR2 (N12453, N12451, N4559);
not NOT1 (N12454, N12425);
nor NOR4 (N12455, N12450, N5421, N11321, N5484);
and AND2 (N12456, N12454, N6536);
or OR3 (N12457, N12455, N4824, N7623);
buf BUF1 (N12458, N12449);
not NOT1 (N12459, N12426);
and AND2 (N12460, N12448, N11495);
and AND2 (N12461, N12452, N11970);
buf BUF1 (N12462, N12461);
and AND3 (N12463, N12457, N10893, N6149);
nor NOR4 (N12464, N12440, N6141, N2355, N9940);
or OR4 (N12465, N12458, N7228, N12332, N5970);
nor NOR2 (N12466, N12456, N8403);
and AND4 (N12467, N12466, N2448, N8331, N9372);
not NOT1 (N12468, N12459);
nand NAND3 (N12469, N12453, N10690, N4286);
nand NAND3 (N12470, N12446, N10481, N7067);
not NOT1 (N12471, N12438);
not NOT1 (N12472, N12471);
nand NAND4 (N12473, N12469, N2005, N2814, N11221);
buf BUF1 (N12474, N12473);
nand NAND4 (N12475, N12470, N8767, N6324, N11214);
or OR2 (N12476, N12475, N5927);
xor XOR2 (N12477, N12463, N5079);
nor NOR3 (N12478, N12465, N1901, N3135);
nand NAND4 (N12479, N12460, N3783, N9804, N3471);
or OR4 (N12480, N12472, N769, N4103, N10025);
and AND4 (N12481, N12468, N5847, N4884, N547);
xor XOR2 (N12482, N12474, N9286);
nand NAND4 (N12483, N12481, N10352, N2661, N3960);
xor XOR2 (N12484, N12479, N839);
or OR2 (N12485, N12482, N209);
nor NOR4 (N12486, N12485, N5036, N9142, N2993);
or OR4 (N12487, N12477, N10395, N5927, N358);
nand NAND3 (N12488, N12476, N7923, N1630);
nor NOR2 (N12489, N12487, N2069);
not NOT1 (N12490, N12488);
buf BUF1 (N12491, N12462);
xor XOR2 (N12492, N12464, N4491);
nand NAND4 (N12493, N12467, N8578, N6398, N10001);
nor NOR4 (N12494, N12491, N4447, N1605, N2445);
nand NAND4 (N12495, N12492, N4800, N4832, N11487);
buf BUF1 (N12496, N12484);
nand NAND4 (N12497, N12486, N7504, N9940, N5248);
nor NOR3 (N12498, N12495, N4575, N964);
or OR3 (N12499, N12494, N11921, N9691);
and AND3 (N12500, N12498, N8459, N8964);
nand NAND4 (N12501, N12493, N937, N3657, N3235);
nand NAND4 (N12502, N12480, N5644, N4617, N9026);
xor XOR2 (N12503, N12489, N794);
not NOT1 (N12504, N12500);
or OR2 (N12505, N12497, N3739);
or OR4 (N12506, N12504, N7869, N5828, N2891);
buf BUF1 (N12507, N12499);
xor XOR2 (N12508, N12502, N102);
xor XOR2 (N12509, N12483, N2676);
nor NOR3 (N12510, N12501, N2881, N9429);
buf BUF1 (N12511, N12506);
not NOT1 (N12512, N12490);
buf BUF1 (N12513, N12505);
not NOT1 (N12514, N12509);
buf BUF1 (N12515, N12503);
and AND3 (N12516, N12478, N2340, N446);
or OR4 (N12517, N12511, N9667, N9705, N3471);
nor NOR2 (N12518, N12516, N12457);
nor NOR3 (N12519, N12517, N1518, N10281);
nor NOR2 (N12520, N12518, N3272);
buf BUF1 (N12521, N12515);
nand NAND4 (N12522, N12513, N4032, N7422, N3759);
not NOT1 (N12523, N12521);
and AND3 (N12524, N12510, N7477, N4806);
or OR4 (N12525, N12523, N7464, N1013, N6793);
buf BUF1 (N12526, N12524);
and AND4 (N12527, N12507, N9755, N1168, N9392);
buf BUF1 (N12528, N12512);
or OR4 (N12529, N12526, N1645, N9403, N5265);
or OR4 (N12530, N12508, N1839, N7585, N5966);
nand NAND3 (N12531, N12514, N2768, N5239);
nor NOR2 (N12532, N12531, N5735);
or OR3 (N12533, N12496, N10062, N11543);
nor NOR2 (N12534, N12527, N2892);
not NOT1 (N12535, N12532);
not NOT1 (N12536, N12533);
nand NAND4 (N12537, N12529, N4887, N1179, N1710);
nor NOR3 (N12538, N12530, N2212, N5473);
or OR3 (N12539, N12528, N10219, N9913);
nor NOR4 (N12540, N12525, N5913, N1142, N5355);
not NOT1 (N12541, N12522);
and AND3 (N12542, N12538, N696, N12125);
buf BUF1 (N12543, N12541);
nor NOR2 (N12544, N12542, N8739);
buf BUF1 (N12545, N12535);
nor NOR3 (N12546, N12520, N10096, N4031);
xor XOR2 (N12547, N12546, N2586);
xor XOR2 (N12548, N12539, N9638);
not NOT1 (N12549, N12519);
or OR2 (N12550, N12536, N9690);
nor NOR3 (N12551, N12543, N6361, N10616);
nand NAND2 (N12552, N12550, N9790);
or OR4 (N12553, N12552, N12515, N10875, N12439);
xor XOR2 (N12554, N12551, N1805);
buf BUF1 (N12555, N12540);
nand NAND2 (N12556, N12548, N5194);
xor XOR2 (N12557, N12554, N11690);
buf BUF1 (N12558, N12537);
and AND4 (N12559, N12555, N8290, N10464, N11375);
nand NAND4 (N12560, N12559, N10420, N1068, N12481);
xor XOR2 (N12561, N12545, N10916);
nor NOR3 (N12562, N12560, N3217, N5940);
and AND4 (N12563, N12558, N2728, N2142, N7231);
xor XOR2 (N12564, N12547, N4314);
nor NOR3 (N12565, N12562, N11453, N1833);
not NOT1 (N12566, N12553);
nand NAND4 (N12567, N12566, N7726, N1790, N1535);
nand NAND4 (N12568, N12564, N8548, N5710, N2700);
or OR2 (N12569, N12534, N10639);
not NOT1 (N12570, N12565);
or OR3 (N12571, N12567, N9626, N5873);
and AND3 (N12572, N12557, N3811, N9761);
nor NOR3 (N12573, N12572, N7059, N9394);
buf BUF1 (N12574, N12570);
nor NOR2 (N12575, N12568, N8295);
or OR2 (N12576, N12574, N287);
nor NOR3 (N12577, N12569, N5781, N4318);
and AND4 (N12578, N12576, N2581, N9629, N4737);
nor NOR4 (N12579, N12563, N8163, N573, N457);
nor NOR3 (N12580, N12549, N5474, N11976);
nand NAND3 (N12581, N12579, N8866, N8603);
buf BUF1 (N12582, N12577);
or OR3 (N12583, N12580, N668, N8939);
nand NAND3 (N12584, N12571, N2380, N3722);
nor NOR2 (N12585, N12583, N6409);
not NOT1 (N12586, N12573);
or OR4 (N12587, N12582, N12250, N5882, N7737);
or OR4 (N12588, N12587, N6254, N8658, N3101);
or OR3 (N12589, N12578, N8837, N12378);
not NOT1 (N12590, N12586);
nand NAND2 (N12591, N12590, N7937);
and AND3 (N12592, N12589, N7839, N12266);
buf BUF1 (N12593, N12592);
xor XOR2 (N12594, N12591, N6968);
or OR2 (N12595, N12544, N4814);
or OR2 (N12596, N12561, N6133);
and AND2 (N12597, N12595, N1486);
buf BUF1 (N12598, N12575);
nand NAND3 (N12599, N12588, N6908, N4475);
or OR3 (N12600, N12598, N1006, N2957);
not NOT1 (N12601, N12594);
not NOT1 (N12602, N12585);
or OR4 (N12603, N12599, N6355, N3911, N4551);
xor XOR2 (N12604, N12593, N4151);
buf BUF1 (N12605, N12584);
buf BUF1 (N12606, N12581);
buf BUF1 (N12607, N12556);
buf BUF1 (N12608, N12600);
xor XOR2 (N12609, N12606, N11505);
or OR2 (N12610, N12609, N5147);
nand NAND2 (N12611, N12601, N1327);
or OR2 (N12612, N12604, N6242);
not NOT1 (N12613, N12610);
or OR4 (N12614, N12597, N12154, N8188, N10274);
and AND3 (N12615, N12602, N12575, N4355);
not NOT1 (N12616, N12613);
nor NOR4 (N12617, N12607, N12066, N3645, N6192);
or OR2 (N12618, N12605, N10578);
not NOT1 (N12619, N12616);
or OR3 (N12620, N12603, N9102, N7567);
nor NOR2 (N12621, N12617, N9212);
nor NOR4 (N12622, N12618, N7373, N7874, N9901);
and AND3 (N12623, N12614, N11652, N1530);
xor XOR2 (N12624, N12611, N1254);
not NOT1 (N12625, N12621);
not NOT1 (N12626, N12596);
or OR3 (N12627, N12615, N3429, N7152);
and AND2 (N12628, N12620, N2496);
or OR3 (N12629, N12623, N11612, N12179);
and AND3 (N12630, N12612, N935, N6807);
nand NAND4 (N12631, N12627, N2310, N296, N5);
not NOT1 (N12632, N12622);
buf BUF1 (N12633, N12630);
or OR3 (N12634, N12625, N7680, N6733);
not NOT1 (N12635, N12634);
nor NOR3 (N12636, N12629, N1961, N6994);
buf BUF1 (N12637, N12626);
or OR3 (N12638, N12633, N1497, N7040);
xor XOR2 (N12639, N12624, N10888);
nand NAND3 (N12640, N12638, N8802, N3459);
not NOT1 (N12641, N12636);
not NOT1 (N12642, N12608);
and AND2 (N12643, N12637, N10687);
or OR3 (N12644, N12619, N1984, N4913);
nor NOR4 (N12645, N12635, N3294, N9430, N6649);
xor XOR2 (N12646, N12642, N8671);
buf BUF1 (N12647, N12632);
and AND4 (N12648, N12639, N8824, N9165, N6755);
xor XOR2 (N12649, N12647, N10606);
or OR2 (N12650, N12643, N9675);
not NOT1 (N12651, N12644);
nand NAND4 (N12652, N12641, N9764, N980, N4538);
buf BUF1 (N12653, N12646);
buf BUF1 (N12654, N12650);
nor NOR3 (N12655, N12640, N11763, N7586);
nand NAND2 (N12656, N12653, N2394);
or OR2 (N12657, N12628, N5718);
buf BUF1 (N12658, N12656);
not NOT1 (N12659, N12645);
buf BUF1 (N12660, N12659);
or OR4 (N12661, N12657, N9372, N4920, N6521);
or OR4 (N12662, N12654, N3535, N6007, N6332);
not NOT1 (N12663, N12660);
and AND3 (N12664, N12648, N6735, N4518);
and AND2 (N12665, N12663, N9127);
nor NOR3 (N12666, N12631, N11992, N49);
and AND4 (N12667, N12664, N10257, N2327, N493);
xor XOR2 (N12668, N12655, N7454);
and AND3 (N12669, N12661, N12386, N9793);
nor NOR3 (N12670, N12668, N2218, N1690);
buf BUF1 (N12671, N12669);
xor XOR2 (N12672, N12666, N4654);
nor NOR4 (N12673, N12651, N1784, N10887, N3924);
xor XOR2 (N12674, N12658, N3998);
nand NAND3 (N12675, N12649, N5639, N6354);
buf BUF1 (N12676, N12674);
buf BUF1 (N12677, N12676);
buf BUF1 (N12678, N12667);
and AND3 (N12679, N12673, N5780, N11416);
or OR4 (N12680, N12678, N652, N1343, N7249);
nor NOR2 (N12681, N12665, N3700);
xor XOR2 (N12682, N12671, N2517);
not NOT1 (N12683, N12652);
nand NAND4 (N12684, N12662, N3797, N6845, N3207);
or OR2 (N12685, N12670, N1023);
or OR4 (N12686, N12684, N11988, N31, N9412);
not NOT1 (N12687, N12681);
or OR3 (N12688, N12687, N5683, N5234);
xor XOR2 (N12689, N12686, N1608);
buf BUF1 (N12690, N12682);
buf BUF1 (N12691, N12680);
nand NAND2 (N12692, N12672, N6702);
nor NOR3 (N12693, N12690, N729, N6329);
not NOT1 (N12694, N12688);
xor XOR2 (N12695, N12675, N2561);
or OR3 (N12696, N12677, N120, N2309);
buf BUF1 (N12697, N12679);
buf BUF1 (N12698, N12689);
xor XOR2 (N12699, N12695, N2222);
or OR3 (N12700, N12691, N6110, N2108);
nand NAND3 (N12701, N12697, N10631, N3761);
nor NOR3 (N12702, N12683, N7016, N2696);
xor XOR2 (N12703, N12696, N8564);
or OR3 (N12704, N12701, N8724, N4841);
nand NAND3 (N12705, N12698, N3237, N3107);
or OR2 (N12706, N12685, N3120);
or OR3 (N12707, N12694, N2181, N11381);
and AND4 (N12708, N12703, N4069, N12111, N8649);
buf BUF1 (N12709, N12706);
xor XOR2 (N12710, N12692, N7810);
xor XOR2 (N12711, N12700, N2908);
and AND4 (N12712, N12702, N7490, N5238, N5840);
or OR4 (N12713, N12707, N12236, N2009, N8451);
and AND3 (N12714, N12693, N5839, N3418);
buf BUF1 (N12715, N12704);
nor NOR3 (N12716, N12712, N8654, N12112);
and AND4 (N12717, N12711, N5021, N7932, N3622);
and AND4 (N12718, N12713, N2126, N1900, N1934);
nor NOR3 (N12719, N12716, N9919, N4482);
buf BUF1 (N12720, N12717);
not NOT1 (N12721, N12714);
nor NOR4 (N12722, N12708, N9354, N11299, N96);
and AND2 (N12723, N12709, N10546);
nor NOR3 (N12724, N12718, N10573, N1682);
or OR3 (N12725, N12721, N12013, N2496);
not NOT1 (N12726, N12720);
xor XOR2 (N12727, N12719, N7637);
buf BUF1 (N12728, N12726);
nor NOR4 (N12729, N12715, N12532, N12602, N8190);
buf BUF1 (N12730, N12710);
nor NOR2 (N12731, N12722, N6052);
not NOT1 (N12732, N12727);
xor XOR2 (N12733, N12731, N5233);
buf BUF1 (N12734, N12730);
not NOT1 (N12735, N12732);
not NOT1 (N12736, N12725);
buf BUF1 (N12737, N12723);
buf BUF1 (N12738, N12733);
buf BUF1 (N12739, N12734);
xor XOR2 (N12740, N12736, N5694);
nor NOR3 (N12741, N12735, N7421, N4290);
nand NAND3 (N12742, N12737, N8075, N4343);
and AND3 (N12743, N12740, N1282, N7815);
buf BUF1 (N12744, N12741);
xor XOR2 (N12745, N12743, N12596);
nor NOR3 (N12746, N12729, N11215, N3512);
nor NOR2 (N12747, N12724, N11589);
nand NAND3 (N12748, N12744, N12744, N3022);
not NOT1 (N12749, N12699);
or OR2 (N12750, N12745, N4134);
or OR3 (N12751, N12748, N11881, N2704);
buf BUF1 (N12752, N12738);
nand NAND2 (N12753, N12739, N858);
or OR2 (N12754, N12742, N9582);
nor NOR3 (N12755, N12749, N10572, N12222);
or OR2 (N12756, N12751, N4533);
and AND4 (N12757, N12747, N2464, N4735, N4025);
xor XOR2 (N12758, N12753, N50);
or OR4 (N12759, N12752, N4602, N12299, N10013);
nand NAND3 (N12760, N12759, N3990, N9876);
not NOT1 (N12761, N12750);
and AND3 (N12762, N12728, N7870, N4741);
and AND2 (N12763, N12760, N4775);
nand NAND4 (N12764, N12756, N4159, N823, N4842);
not NOT1 (N12765, N12764);
nor NOR4 (N12766, N12758, N12538, N1352, N7798);
xor XOR2 (N12767, N12754, N6040);
nor NOR3 (N12768, N12761, N4169, N10618);
xor XOR2 (N12769, N12765, N9964);
buf BUF1 (N12770, N12705);
and AND2 (N12771, N12767, N2799);
or OR3 (N12772, N12762, N1228, N1271);
xor XOR2 (N12773, N12769, N5582);
and AND4 (N12774, N12771, N10906, N10267, N2985);
and AND2 (N12775, N12774, N6888);
or OR4 (N12776, N12763, N6062, N6842, N2895);
buf BUF1 (N12777, N12757);
or OR2 (N12778, N12766, N665);
nand NAND4 (N12779, N12775, N6937, N1004, N10806);
buf BUF1 (N12780, N12779);
buf BUF1 (N12781, N12776);
nor NOR2 (N12782, N12772, N4566);
nor NOR2 (N12783, N12746, N8650);
buf BUF1 (N12784, N12780);
xor XOR2 (N12785, N12782, N5407);
and AND2 (N12786, N12785, N6235);
not NOT1 (N12787, N12786);
nor NOR2 (N12788, N12783, N11568);
or OR3 (N12789, N12770, N827, N8561);
nor NOR3 (N12790, N12755, N6935, N9913);
nand NAND4 (N12791, N12789, N1805, N11161, N539);
nand NAND3 (N12792, N12791, N12575, N7964);
nor NOR4 (N12793, N12784, N7811, N4049, N340);
and AND2 (N12794, N12792, N11010);
or OR2 (N12795, N12768, N9285);
or OR2 (N12796, N12794, N1260);
nor NOR4 (N12797, N12773, N4823, N5149, N10369);
or OR2 (N12798, N12795, N6676);
or OR2 (N12799, N12797, N1949);
buf BUF1 (N12800, N12777);
nor NOR4 (N12801, N12798, N3674, N10079, N4315);
buf BUF1 (N12802, N12799);
buf BUF1 (N12803, N12788);
or OR2 (N12804, N12793, N6950);
or OR4 (N12805, N12778, N7972, N1352, N2171);
or OR2 (N12806, N12805, N10483);
nor NOR2 (N12807, N12803, N2780);
buf BUF1 (N12808, N12801);
and AND4 (N12809, N12806, N2878, N9770, N2147);
xor XOR2 (N12810, N12802, N10307);
and AND3 (N12811, N12796, N299, N11991);
or OR4 (N12812, N12811, N8488, N4188, N2247);
not NOT1 (N12813, N12808);
nor NOR2 (N12814, N12810, N7344);
buf BUF1 (N12815, N12807);
nand NAND2 (N12816, N12814, N7837);
endmodule