// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N6405,N6414,N6416,N6406,N6418,N6420,N6409,N6419,N6412,N6421;

not NOT1 (N22, N14);
and AND2 (N23, N17, N13);
nand NAND3 (N24, N13, N4, N13);
buf BUF1 (N25, N9);
nor NOR3 (N26, N7, N1, N20);
and AND3 (N27, N6, N9, N25);
xor XOR2 (N28, N9, N5);
or OR2 (N29, N22, N16);
nor NOR2 (N30, N20, N2);
buf BUF1 (N31, N4);
buf BUF1 (N32, N6);
buf BUF1 (N33, N25);
or OR4 (N34, N32, N2, N18, N21);
nor NOR4 (N35, N27, N10, N30, N3);
nor NOR3 (N36, N32, N29, N13);
and AND2 (N37, N15, N24);
nand NAND3 (N38, N4, N35, N1);
or OR4 (N39, N22, N25, N3, N20);
xor XOR2 (N40, N31, N4);
and AND4 (N41, N39, N27, N14, N4);
or OR4 (N42, N41, N20, N35, N41);
not NOT1 (N43, N42);
nor NOR2 (N44, N43, N26);
not NOT1 (N45, N7);
or OR2 (N46, N23, N3);
xor XOR2 (N47, N36, N27);
buf BUF1 (N48, N28);
nand NAND3 (N49, N38, N33, N13);
nor NOR4 (N50, N22, N18, N37, N25);
buf BUF1 (N51, N43);
nor NOR4 (N52, N40, N9, N31, N5);
not NOT1 (N53, N49);
nor NOR3 (N54, N45, N5, N47);
nand NAND3 (N55, N32, N40, N27);
nor NOR2 (N56, N34, N6);
not NOT1 (N57, N52);
xor XOR2 (N58, N55, N50);
not NOT1 (N59, N25);
nor NOR4 (N60, N48, N46, N28, N21);
xor XOR2 (N61, N4, N26);
xor XOR2 (N62, N51, N6);
nand NAND3 (N63, N62, N31, N6);
and AND4 (N64, N53, N62, N57, N62);
buf BUF1 (N65, N61);
nor NOR2 (N66, N29, N4);
nand NAND3 (N67, N44, N10, N6);
buf BUF1 (N68, N63);
xor XOR2 (N69, N68, N51);
nand NAND2 (N70, N67, N33);
nor NOR4 (N71, N59, N58, N42, N56);
not NOT1 (N72, N60);
buf BUF1 (N73, N28);
xor XOR2 (N74, N5, N51);
xor XOR2 (N75, N74, N37);
or OR3 (N76, N65, N7, N17);
nand NAND4 (N77, N70, N15, N36, N17);
not NOT1 (N78, N76);
xor XOR2 (N79, N77, N51);
buf BUF1 (N80, N75);
nand NAND4 (N81, N73, N70, N54, N33);
nor NOR2 (N82, N56, N57);
nand NAND2 (N83, N69, N77);
nor NOR3 (N84, N83, N35, N28);
nand NAND4 (N85, N72, N73, N69, N31);
nand NAND4 (N86, N82, N57, N4, N74);
nand NAND3 (N87, N84, N39, N36);
not NOT1 (N88, N80);
xor XOR2 (N89, N87, N53);
nor NOR4 (N90, N85, N44, N84, N8);
nor NOR2 (N91, N64, N15);
nand NAND2 (N92, N88, N2);
or OR3 (N93, N71, N22, N5);
or OR4 (N94, N89, N38, N37, N90);
nand NAND4 (N95, N22, N40, N21, N32);
nor NOR2 (N96, N94, N37);
nor NOR4 (N97, N79, N92, N35, N34);
and AND4 (N98, N79, N53, N12, N44);
nand NAND3 (N99, N86, N95, N55);
nand NAND4 (N100, N32, N74, N42, N7);
not NOT1 (N101, N66);
buf BUF1 (N102, N91);
and AND2 (N103, N100, N70);
or OR3 (N104, N96, N101, N42);
or OR4 (N105, N56, N29, N104, N52);
buf BUF1 (N106, N53);
xor XOR2 (N107, N93, N38);
buf BUF1 (N108, N103);
not NOT1 (N109, N99);
nor NOR3 (N110, N102, N22, N22);
or OR4 (N111, N105, N69, N2, N83);
or OR2 (N112, N98, N7);
xor XOR2 (N113, N110, N111);
nand NAND4 (N114, N106, N12, N76, N37);
and AND4 (N115, N52, N92, N42, N41);
not NOT1 (N116, N78);
and AND2 (N117, N115, N15);
buf BUF1 (N118, N108);
nand NAND3 (N119, N81, N32, N12);
buf BUF1 (N120, N113);
not NOT1 (N121, N116);
xor XOR2 (N122, N114, N107);
not NOT1 (N123, N90);
xor XOR2 (N124, N117, N26);
and AND3 (N125, N97, N5, N30);
and AND2 (N126, N124, N35);
buf BUF1 (N127, N126);
or OR2 (N128, N112, N6);
nand NAND2 (N129, N123, N38);
nand NAND2 (N130, N122, N79);
nand NAND3 (N131, N120, N106, N66);
xor XOR2 (N132, N109, N30);
nand NAND3 (N133, N132, N63, N4);
buf BUF1 (N134, N130);
buf BUF1 (N135, N133);
not NOT1 (N136, N135);
nor NOR2 (N137, N134, N96);
not NOT1 (N138, N118);
buf BUF1 (N139, N131);
not NOT1 (N140, N139);
nor NOR2 (N141, N121, N137);
nor NOR2 (N142, N6, N128);
nand NAND4 (N143, N20, N53, N134, N125);
buf BUF1 (N144, N56);
and AND3 (N145, N127, N120, N31);
xor XOR2 (N146, N141, N19);
or OR3 (N147, N146, N126, N116);
buf BUF1 (N148, N138);
nand NAND3 (N149, N129, N132, N99);
nor NOR2 (N150, N145, N43);
and AND4 (N151, N140, N139, N19, N134);
not NOT1 (N152, N136);
xor XOR2 (N153, N152, N81);
and AND2 (N154, N144, N67);
nand NAND2 (N155, N153, N123);
nor NOR2 (N156, N143, N80);
nand NAND2 (N157, N119, N137);
buf BUF1 (N158, N150);
nor NOR2 (N159, N155, N116);
xor XOR2 (N160, N149, N88);
nand NAND3 (N161, N160, N72, N93);
or OR4 (N162, N159, N90, N72, N37);
nand NAND2 (N163, N147, N124);
buf BUF1 (N164, N157);
buf BUF1 (N165, N161);
and AND2 (N166, N158, N19);
nor NOR4 (N167, N154, N44, N131, N53);
not NOT1 (N168, N164);
or OR2 (N169, N162, N105);
and AND3 (N170, N166, N104, N140);
or OR2 (N171, N163, N162);
not NOT1 (N172, N167);
xor XOR2 (N173, N156, N151);
xor XOR2 (N174, N123, N43);
nor NOR4 (N175, N172, N19, N117, N104);
nand NAND2 (N176, N170, N130);
not NOT1 (N177, N169);
nand NAND3 (N178, N175, N169, N70);
xor XOR2 (N179, N173, N168);
buf BUF1 (N180, N89);
not NOT1 (N181, N171);
xor XOR2 (N182, N165, N97);
xor XOR2 (N183, N181, N14);
and AND2 (N184, N174, N17);
or OR3 (N185, N179, N17, N113);
nor NOR2 (N186, N183, N72);
xor XOR2 (N187, N180, N151);
and AND3 (N188, N182, N100, N62);
or OR2 (N189, N178, N164);
or OR4 (N190, N189, N82, N13, N23);
nand NAND2 (N191, N142, N8);
buf BUF1 (N192, N177);
and AND4 (N193, N191, N89, N176, N101);
buf BUF1 (N194, N137);
nor NOR3 (N195, N193, N49, N130);
nand NAND2 (N196, N190, N145);
and AND3 (N197, N185, N144, N124);
and AND3 (N198, N184, N43, N12);
or OR4 (N199, N196, N159, N142, N110);
not NOT1 (N200, N188);
and AND3 (N201, N194, N66, N104);
and AND4 (N202, N148, N125, N100, N163);
not NOT1 (N203, N187);
xor XOR2 (N204, N202, N55);
or OR3 (N205, N204, N19, N106);
xor XOR2 (N206, N186, N171);
nand NAND2 (N207, N203, N184);
buf BUF1 (N208, N195);
or OR2 (N209, N208, N143);
not NOT1 (N210, N197);
nand NAND4 (N211, N200, N175, N101, N168);
xor XOR2 (N212, N192, N13);
and AND4 (N213, N205, N8, N37, N139);
or OR2 (N214, N211, N92);
xor XOR2 (N215, N210, N6);
or OR2 (N216, N206, N107);
nand NAND2 (N217, N207, N120);
and AND2 (N218, N212, N3);
and AND4 (N219, N213, N208, N150, N130);
buf BUF1 (N220, N216);
not NOT1 (N221, N209);
not NOT1 (N222, N198);
xor XOR2 (N223, N222, N136);
and AND2 (N224, N201, N57);
nor NOR2 (N225, N223, N74);
and AND3 (N226, N215, N214, N92);
buf BUF1 (N227, N83);
nor NOR2 (N228, N225, N52);
not NOT1 (N229, N221);
nand NAND3 (N230, N218, N98, N170);
and AND3 (N231, N199, N9, N209);
and AND4 (N232, N217, N84, N164, N26);
nor NOR3 (N233, N230, N140, N92);
nor NOR3 (N234, N227, N91, N19);
nand NAND4 (N235, N224, N73, N38, N215);
or OR2 (N236, N232, N42);
not NOT1 (N237, N235);
xor XOR2 (N238, N220, N235);
or OR2 (N239, N219, N194);
nand NAND3 (N240, N238, N148, N115);
nor NOR2 (N241, N240, N93);
or OR4 (N242, N228, N62, N48, N187);
xor XOR2 (N243, N234, N186);
or OR4 (N244, N233, N112, N68, N4);
xor XOR2 (N245, N231, N242);
or OR3 (N246, N92, N76, N9);
nand NAND4 (N247, N229, N33, N167, N104);
nand NAND2 (N248, N237, N237);
xor XOR2 (N249, N246, N86);
nor NOR4 (N250, N236, N20, N29, N141);
not NOT1 (N251, N249);
not NOT1 (N252, N243);
or OR4 (N253, N247, N242, N228, N141);
not NOT1 (N254, N252);
xor XOR2 (N255, N241, N219);
nand NAND3 (N256, N226, N179, N220);
not NOT1 (N257, N248);
and AND4 (N258, N253, N177, N254, N47);
xor XOR2 (N259, N251, N82);
not NOT1 (N260, N227);
buf BUF1 (N261, N245);
or OR4 (N262, N258, N119, N7, N194);
nor NOR3 (N263, N261, N197, N130);
nor NOR3 (N264, N263, N112, N51);
nand NAND3 (N265, N259, N230, N100);
nand NAND2 (N266, N264, N68);
or OR2 (N267, N260, N248);
buf BUF1 (N268, N250);
not NOT1 (N269, N265);
and AND2 (N270, N256, N169);
nor NOR4 (N271, N268, N97, N54, N103);
nor NOR3 (N272, N266, N36, N196);
not NOT1 (N273, N272);
nor NOR3 (N274, N255, N227, N217);
buf BUF1 (N275, N244);
and AND3 (N276, N267, N223, N177);
nand NAND2 (N277, N270, N272);
buf BUF1 (N278, N277);
or OR4 (N279, N274, N178, N163, N107);
xor XOR2 (N280, N262, N147);
nor NOR3 (N281, N269, N190, N129);
and AND2 (N282, N257, N62);
buf BUF1 (N283, N282);
buf BUF1 (N284, N283);
nor NOR4 (N285, N271, N277, N107, N71);
or OR4 (N286, N285, N209, N207, N251);
nand NAND2 (N287, N280, N279);
or OR2 (N288, N62, N25);
nand NAND3 (N289, N287, N26, N73);
not NOT1 (N290, N276);
not NOT1 (N291, N289);
xor XOR2 (N292, N278, N224);
or OR3 (N293, N290, N134, N66);
or OR2 (N294, N291, N11);
or OR2 (N295, N292, N261);
not NOT1 (N296, N239);
xor XOR2 (N297, N281, N96);
or OR3 (N298, N297, N219, N293);
buf BUF1 (N299, N42);
and AND3 (N300, N299, N199, N163);
xor XOR2 (N301, N273, N64);
nand NAND4 (N302, N288, N210, N37, N218);
nor NOR2 (N303, N301, N256);
or OR4 (N304, N296, N108, N149, N38);
not NOT1 (N305, N284);
xor XOR2 (N306, N300, N134);
and AND3 (N307, N305, N3, N89);
or OR4 (N308, N286, N77, N221, N267);
nand NAND2 (N309, N306, N68);
nor NOR2 (N310, N294, N284);
buf BUF1 (N311, N307);
nor NOR4 (N312, N302, N242, N42, N31);
nand NAND3 (N313, N308, N111, N79);
or OR3 (N314, N295, N238, N116);
not NOT1 (N315, N312);
nor NOR4 (N316, N310, N291, N270, N128);
or OR3 (N317, N315, N285, N32);
xor XOR2 (N318, N311, N228);
and AND2 (N319, N316, N63);
xor XOR2 (N320, N309, N304);
or OR2 (N321, N296, N195);
nand NAND3 (N322, N318, N33, N180);
xor XOR2 (N323, N321, N202);
buf BUF1 (N324, N317);
or OR2 (N325, N314, N281);
or OR4 (N326, N325, N2, N307, N145);
buf BUF1 (N327, N275);
nor NOR2 (N328, N322, N197);
nor NOR2 (N329, N303, N154);
nand NAND3 (N330, N323, N116, N199);
and AND3 (N331, N320, N132, N34);
xor XOR2 (N332, N331, N204);
not NOT1 (N333, N330);
and AND2 (N334, N326, N205);
xor XOR2 (N335, N327, N300);
nand NAND3 (N336, N329, N9, N318);
nand NAND2 (N337, N313, N168);
nand NAND4 (N338, N319, N22, N167, N284);
and AND3 (N339, N334, N263, N129);
and AND2 (N340, N333, N223);
not NOT1 (N341, N298);
nand NAND4 (N342, N332, N147, N144, N223);
buf BUF1 (N343, N335);
or OR4 (N344, N324, N283, N151, N49);
or OR2 (N345, N338, N337);
or OR3 (N346, N278, N183, N250);
nor NOR2 (N347, N342, N44);
not NOT1 (N348, N345);
nand NAND3 (N349, N328, N189, N63);
or OR3 (N350, N339, N65, N316);
xor XOR2 (N351, N341, N178);
buf BUF1 (N352, N351);
nor NOR2 (N353, N336, N11);
nor NOR4 (N354, N349, N258, N203, N255);
nand NAND4 (N355, N344, N311, N220, N298);
buf BUF1 (N356, N343);
not NOT1 (N357, N355);
nor NOR2 (N358, N350, N79);
and AND3 (N359, N354, N90, N170);
nand NAND4 (N360, N357, N154, N36, N82);
buf BUF1 (N361, N352);
nor NOR4 (N362, N340, N5, N278, N216);
nand NAND2 (N363, N356, N80);
buf BUF1 (N364, N346);
nor NOR4 (N365, N347, N103, N316, N56);
nor NOR3 (N366, N348, N245, N155);
nand NAND4 (N367, N353, N178, N161, N175);
or OR4 (N368, N367, N228, N178, N6);
buf BUF1 (N369, N358);
or OR3 (N370, N361, N278, N139);
nor NOR3 (N371, N370, N242, N255);
nand NAND4 (N372, N371, N355, N202, N265);
nand NAND2 (N373, N372, N12);
or OR3 (N374, N366, N151, N125);
nor NOR2 (N375, N369, N314);
xor XOR2 (N376, N360, N373);
nor NOR3 (N377, N335, N249, N372);
and AND4 (N378, N377, N154, N169, N254);
buf BUF1 (N379, N378);
not NOT1 (N380, N359);
or OR3 (N381, N379, N312, N13);
not NOT1 (N382, N376);
nor NOR3 (N383, N363, N86, N37);
not NOT1 (N384, N375);
and AND3 (N385, N368, N121, N263);
buf BUF1 (N386, N380);
xor XOR2 (N387, N382, N162);
buf BUF1 (N388, N364);
or OR3 (N389, N383, N8, N2);
nand NAND3 (N390, N388, N298, N262);
and AND2 (N391, N387, N390);
buf BUF1 (N392, N118);
or OR2 (N393, N374, N144);
not NOT1 (N394, N392);
nand NAND4 (N395, N384, N270, N379, N3);
nor NOR4 (N396, N362, N227, N281, N295);
not NOT1 (N397, N365);
or OR3 (N398, N385, N267, N128);
not NOT1 (N399, N398);
not NOT1 (N400, N396);
nand NAND2 (N401, N399, N394);
and AND4 (N402, N165, N196, N250, N347);
or OR4 (N403, N386, N54, N74, N402);
nor NOR2 (N404, N219, N264);
not NOT1 (N405, N397);
or OR4 (N406, N401, N165, N271, N97);
xor XOR2 (N407, N381, N58);
or OR3 (N408, N405, N236, N233);
not NOT1 (N409, N403);
nand NAND4 (N410, N400, N15, N219, N349);
buf BUF1 (N411, N408);
not NOT1 (N412, N391);
xor XOR2 (N413, N407, N390);
nand NAND3 (N414, N395, N47, N49);
and AND4 (N415, N413, N240, N109, N161);
nor NOR3 (N416, N410, N34, N91);
nor NOR2 (N417, N411, N164);
nor NOR3 (N418, N389, N162, N50);
buf BUF1 (N419, N409);
nand NAND4 (N420, N415, N216, N28, N167);
buf BUF1 (N421, N419);
nand NAND4 (N422, N420, N283, N187, N61);
xor XOR2 (N423, N422, N308);
or OR2 (N424, N421, N331);
not NOT1 (N425, N416);
xor XOR2 (N426, N418, N323);
nand NAND2 (N427, N425, N64);
nor NOR4 (N428, N417, N262, N322, N85);
xor XOR2 (N429, N414, N302);
buf BUF1 (N430, N412);
buf BUF1 (N431, N430);
buf BUF1 (N432, N427);
not NOT1 (N433, N424);
not NOT1 (N434, N432);
buf BUF1 (N435, N429);
buf BUF1 (N436, N393);
nand NAND3 (N437, N436, N81, N33);
nand NAND4 (N438, N435, N276, N23, N431);
and AND3 (N439, N328, N19, N365);
or OR4 (N440, N428, N425, N219, N68);
and AND4 (N441, N440, N137, N7, N360);
buf BUF1 (N442, N438);
and AND2 (N443, N439, N102);
xor XOR2 (N444, N441, N198);
and AND4 (N445, N442, N335, N7, N175);
nand NAND3 (N446, N434, N352, N278);
xor XOR2 (N447, N437, N39);
and AND3 (N448, N404, N89, N302);
nor NOR3 (N449, N448, N213, N318);
or OR2 (N450, N423, N3);
xor XOR2 (N451, N445, N95);
or OR3 (N452, N446, N196, N337);
not NOT1 (N453, N451);
nand NAND2 (N454, N444, N318);
nand NAND2 (N455, N452, N305);
and AND2 (N456, N426, N171);
xor XOR2 (N457, N433, N34);
xor XOR2 (N458, N406, N359);
xor XOR2 (N459, N455, N371);
and AND3 (N460, N443, N305, N99);
buf BUF1 (N461, N458);
not NOT1 (N462, N461);
xor XOR2 (N463, N460, N285);
not NOT1 (N464, N447);
not NOT1 (N465, N450);
nor NOR3 (N466, N453, N10, N25);
and AND3 (N467, N463, N377, N51);
not NOT1 (N468, N466);
and AND2 (N469, N465, N119);
or OR4 (N470, N468, N56, N406, N401);
not NOT1 (N471, N449);
and AND4 (N472, N467, N392, N216, N146);
nand NAND3 (N473, N454, N156, N299);
nand NAND3 (N474, N456, N189, N218);
not NOT1 (N475, N457);
nand NAND3 (N476, N475, N31, N275);
nor NOR3 (N477, N470, N170, N45);
nand NAND4 (N478, N476, N120, N140, N29);
nand NAND3 (N479, N471, N183, N412);
nand NAND2 (N480, N478, N262);
nand NAND2 (N481, N469, N266);
not NOT1 (N482, N462);
buf BUF1 (N483, N472);
nand NAND4 (N484, N479, N420, N94, N233);
or OR2 (N485, N473, N246);
nand NAND3 (N486, N483, N311, N87);
nor NOR3 (N487, N481, N137, N286);
and AND3 (N488, N474, N91, N171);
and AND4 (N489, N464, N20, N416, N450);
nor NOR3 (N490, N477, N447, N47);
nand NAND4 (N491, N489, N360, N46, N54);
nor NOR2 (N492, N488, N272);
nand NAND4 (N493, N485, N174, N132, N351);
nand NAND4 (N494, N492, N122, N35, N486);
and AND2 (N495, N88, N209);
buf BUF1 (N496, N490);
or OR2 (N497, N484, N445);
buf BUF1 (N498, N494);
xor XOR2 (N499, N495, N383);
or OR2 (N500, N487, N393);
buf BUF1 (N501, N497);
xor XOR2 (N502, N493, N434);
xor XOR2 (N503, N500, N9);
nand NAND3 (N504, N459, N113, N296);
xor XOR2 (N505, N499, N149);
buf BUF1 (N506, N504);
nand NAND2 (N507, N496, N242);
xor XOR2 (N508, N498, N1);
xor XOR2 (N509, N503, N94);
nand NAND3 (N510, N505, N480, N47);
xor XOR2 (N511, N338, N428);
xor XOR2 (N512, N482, N93);
or OR4 (N513, N509, N361, N198, N64);
buf BUF1 (N514, N513);
not NOT1 (N515, N507);
xor XOR2 (N516, N491, N204);
buf BUF1 (N517, N514);
not NOT1 (N518, N506);
and AND4 (N519, N502, N383, N341, N190);
nand NAND3 (N520, N515, N451, N13);
or OR2 (N521, N517, N172);
nor NOR2 (N522, N516, N19);
buf BUF1 (N523, N510);
not NOT1 (N524, N512);
xor XOR2 (N525, N520, N351);
and AND2 (N526, N511, N498);
not NOT1 (N527, N519);
or OR3 (N528, N518, N369, N367);
and AND4 (N529, N522, N465, N517, N463);
nor NOR2 (N530, N526, N322);
not NOT1 (N531, N508);
nand NAND4 (N532, N530, N201, N485, N304);
xor XOR2 (N533, N524, N28);
xor XOR2 (N534, N533, N87);
buf BUF1 (N535, N532);
nor NOR3 (N536, N534, N53, N3);
and AND3 (N537, N501, N73, N493);
nand NAND2 (N538, N529, N272);
and AND3 (N539, N538, N311, N157);
buf BUF1 (N540, N535);
and AND2 (N541, N527, N31);
or OR4 (N542, N525, N95, N275, N432);
and AND2 (N543, N521, N127);
buf BUF1 (N544, N542);
not NOT1 (N545, N523);
buf BUF1 (N546, N545);
xor XOR2 (N547, N531, N183);
nand NAND2 (N548, N528, N80);
or OR2 (N549, N543, N269);
nand NAND4 (N550, N546, N340, N464, N153);
not NOT1 (N551, N536);
or OR2 (N552, N551, N329);
xor XOR2 (N553, N540, N55);
buf BUF1 (N554, N550);
not NOT1 (N555, N552);
not NOT1 (N556, N548);
xor XOR2 (N557, N555, N76);
buf BUF1 (N558, N541);
not NOT1 (N559, N554);
buf BUF1 (N560, N553);
buf BUF1 (N561, N544);
nor NOR2 (N562, N556, N34);
not NOT1 (N563, N558);
or OR4 (N564, N562, N188, N385, N548);
not NOT1 (N565, N564);
buf BUF1 (N566, N565);
nor NOR2 (N567, N549, N193);
xor XOR2 (N568, N560, N341);
not NOT1 (N569, N547);
nand NAND4 (N570, N557, N505, N316, N520);
not NOT1 (N571, N561);
buf BUF1 (N572, N571);
nand NAND2 (N573, N566, N555);
and AND4 (N574, N570, N369, N95, N405);
xor XOR2 (N575, N573, N562);
nor NOR3 (N576, N537, N118, N60);
nand NAND4 (N577, N575, N496, N56, N419);
not NOT1 (N578, N574);
not NOT1 (N579, N563);
and AND4 (N580, N572, N2, N368, N341);
nor NOR2 (N581, N539, N15);
nand NAND2 (N582, N568, N328);
nand NAND4 (N583, N567, N233, N324, N358);
or OR3 (N584, N577, N460, N569);
or OR2 (N585, N564, N215);
and AND3 (N586, N582, N143, N377);
and AND2 (N587, N576, N439);
buf BUF1 (N588, N581);
not NOT1 (N589, N583);
nand NAND4 (N590, N585, N135, N100, N5);
xor XOR2 (N591, N559, N218);
nand NAND3 (N592, N587, N319, N91);
xor XOR2 (N593, N584, N6);
xor XOR2 (N594, N591, N203);
not NOT1 (N595, N590);
buf BUF1 (N596, N593);
or OR3 (N597, N592, N108, N28);
not NOT1 (N598, N596);
nor NOR4 (N599, N595, N483, N155, N394);
buf BUF1 (N600, N580);
or OR4 (N601, N578, N228, N127, N56);
xor XOR2 (N602, N598, N343);
xor XOR2 (N603, N594, N228);
buf BUF1 (N604, N586);
not NOT1 (N605, N603);
and AND3 (N606, N605, N531, N605);
buf BUF1 (N607, N589);
not NOT1 (N608, N602);
not NOT1 (N609, N606);
and AND4 (N610, N600, N594, N514, N330);
and AND4 (N611, N609, N7, N98, N110);
buf BUF1 (N612, N607);
or OR4 (N613, N599, N450, N473, N73);
buf BUF1 (N614, N588);
nand NAND3 (N615, N612, N554, N475);
nand NAND4 (N616, N579, N499, N237, N55);
buf BUF1 (N617, N610);
nand NAND3 (N618, N613, N178, N309);
nor NOR3 (N619, N616, N265, N44);
and AND4 (N620, N601, N347, N426, N54);
nand NAND3 (N621, N604, N329, N371);
and AND4 (N622, N617, N27, N201, N615);
xor XOR2 (N623, N162, N565);
not NOT1 (N624, N622);
nand NAND2 (N625, N619, N5);
buf BUF1 (N626, N623);
xor XOR2 (N627, N597, N95);
and AND4 (N628, N627, N8, N543, N311);
and AND2 (N629, N626, N389);
xor XOR2 (N630, N614, N370);
buf BUF1 (N631, N624);
nor NOR2 (N632, N630, N127);
buf BUF1 (N633, N629);
not NOT1 (N634, N631);
xor XOR2 (N635, N620, N458);
nand NAND4 (N636, N625, N159, N435, N321);
and AND3 (N637, N628, N494, N71);
nor NOR4 (N638, N611, N217, N131, N226);
not NOT1 (N639, N632);
or OR3 (N640, N634, N86, N626);
or OR4 (N641, N638, N46, N52, N457);
buf BUF1 (N642, N621);
xor XOR2 (N643, N639, N116);
and AND2 (N644, N635, N634);
nor NOR3 (N645, N641, N285, N339);
xor XOR2 (N646, N636, N111);
nand NAND4 (N647, N618, N255, N615, N398);
xor XOR2 (N648, N640, N458);
buf BUF1 (N649, N648);
nand NAND4 (N650, N633, N439, N102, N10);
nand NAND4 (N651, N644, N241, N106, N604);
buf BUF1 (N652, N650);
not NOT1 (N653, N651);
nand NAND4 (N654, N649, N204, N432, N136);
or OR3 (N655, N646, N444, N338);
nor NOR3 (N656, N643, N84, N118);
xor XOR2 (N657, N642, N174);
xor XOR2 (N658, N653, N57);
or OR4 (N659, N658, N222, N432, N155);
or OR2 (N660, N647, N67);
nand NAND2 (N661, N608, N334);
nor NOR4 (N662, N660, N587, N354, N73);
not NOT1 (N663, N654);
or OR2 (N664, N645, N611);
nor NOR2 (N665, N652, N443);
nand NAND3 (N666, N663, N244, N6);
nand NAND3 (N667, N661, N528, N279);
or OR2 (N668, N637, N95);
and AND3 (N669, N664, N395, N377);
buf BUF1 (N670, N666);
or OR2 (N671, N670, N212);
nand NAND3 (N672, N667, N242, N466);
nand NAND3 (N673, N669, N661, N344);
or OR2 (N674, N672, N404);
nand NAND4 (N675, N656, N308, N58, N437);
and AND3 (N676, N675, N67, N385);
nor NOR4 (N677, N657, N91, N405, N539);
buf BUF1 (N678, N673);
nand NAND2 (N679, N674, N371);
not NOT1 (N680, N668);
buf BUF1 (N681, N677);
nor NOR3 (N682, N681, N475, N45);
or OR4 (N683, N659, N470, N410, N345);
buf BUF1 (N684, N680);
and AND2 (N685, N678, N456);
or OR2 (N686, N662, N597);
not NOT1 (N687, N684);
not NOT1 (N688, N686);
xor XOR2 (N689, N682, N279);
not NOT1 (N690, N665);
not NOT1 (N691, N671);
nor NOR4 (N692, N691, N532, N663, N608);
nand NAND4 (N693, N655, N305, N552, N27);
and AND2 (N694, N688, N646);
and AND4 (N695, N693, N684, N342, N31);
buf BUF1 (N696, N689);
xor XOR2 (N697, N687, N445);
not NOT1 (N698, N676);
or OR4 (N699, N683, N183, N158, N636);
or OR4 (N700, N695, N681, N268, N438);
nand NAND3 (N701, N698, N394, N408);
nand NAND2 (N702, N701, N62);
nor NOR4 (N703, N690, N690, N481, N41);
and AND2 (N704, N685, N181);
buf BUF1 (N705, N679);
nand NAND4 (N706, N702, N481, N540, N444);
or OR2 (N707, N699, N251);
and AND3 (N708, N704, N586, N217);
or OR4 (N709, N696, N183, N200, N530);
or OR4 (N710, N697, N68, N170, N525);
or OR4 (N711, N703, N85, N171, N132);
xor XOR2 (N712, N694, N592);
nor NOR2 (N713, N709, N397);
or OR2 (N714, N708, N308);
nor NOR4 (N715, N711, N704, N191, N479);
and AND4 (N716, N712, N142, N620, N74);
buf BUF1 (N717, N710);
xor XOR2 (N718, N713, N279);
nor NOR3 (N719, N692, N122, N355);
buf BUF1 (N720, N719);
nor NOR4 (N721, N716, N163, N177, N254);
buf BUF1 (N722, N700);
xor XOR2 (N723, N715, N616);
and AND4 (N724, N722, N700, N163, N542);
buf BUF1 (N725, N720);
or OR2 (N726, N706, N245);
buf BUF1 (N727, N726);
or OR2 (N728, N717, N259);
and AND3 (N729, N728, N20, N628);
and AND4 (N730, N725, N301, N392, N317);
buf BUF1 (N731, N707);
buf BUF1 (N732, N730);
nand NAND3 (N733, N727, N545, N550);
nand NAND3 (N734, N714, N264, N358);
not NOT1 (N735, N721);
not NOT1 (N736, N724);
xor XOR2 (N737, N735, N227);
nor NOR3 (N738, N729, N662, N697);
nor NOR3 (N739, N705, N226, N666);
not NOT1 (N740, N737);
or OR2 (N741, N718, N78);
or OR2 (N742, N734, N327);
nand NAND3 (N743, N736, N656, N580);
or OR3 (N744, N743, N626, N564);
not NOT1 (N745, N740);
and AND4 (N746, N738, N98, N185, N148);
or OR2 (N747, N739, N298);
not NOT1 (N748, N744);
nor NOR2 (N749, N742, N569);
not NOT1 (N750, N733);
and AND4 (N751, N750, N637, N610, N568);
nor NOR3 (N752, N723, N333, N514);
xor XOR2 (N753, N746, N583);
nand NAND4 (N754, N741, N145, N357, N381);
or OR3 (N755, N751, N351, N591);
nand NAND2 (N756, N755, N540);
buf BUF1 (N757, N731);
buf BUF1 (N758, N747);
not NOT1 (N759, N748);
nand NAND2 (N760, N757, N533);
nor NOR3 (N761, N759, N394, N356);
xor XOR2 (N762, N754, N589);
or OR2 (N763, N749, N136);
buf BUF1 (N764, N756);
or OR3 (N765, N764, N42, N274);
not NOT1 (N766, N762);
or OR4 (N767, N760, N197, N562, N134);
nor NOR4 (N768, N761, N530, N220, N366);
xor XOR2 (N769, N753, N409);
nor NOR3 (N770, N766, N698, N119);
xor XOR2 (N771, N763, N359);
and AND4 (N772, N768, N532, N703, N426);
and AND3 (N773, N765, N376, N674);
nor NOR3 (N774, N769, N66, N368);
and AND4 (N775, N752, N272, N525, N22);
nor NOR4 (N776, N775, N702, N629, N90);
not NOT1 (N777, N732);
and AND2 (N778, N767, N437);
buf BUF1 (N779, N758);
nor NOR3 (N780, N745, N731, N233);
not NOT1 (N781, N778);
xor XOR2 (N782, N781, N633);
buf BUF1 (N783, N780);
xor XOR2 (N784, N776, N608);
nor NOR3 (N785, N771, N89, N646);
and AND3 (N786, N770, N215, N575);
nor NOR2 (N787, N786, N695);
nor NOR2 (N788, N784, N365);
nand NAND3 (N789, N772, N436, N34);
nand NAND2 (N790, N774, N380);
nor NOR3 (N791, N773, N789, N571);
xor XOR2 (N792, N428, N617);
not NOT1 (N793, N777);
buf BUF1 (N794, N793);
buf BUF1 (N795, N787);
buf BUF1 (N796, N779);
not NOT1 (N797, N792);
nand NAND4 (N798, N783, N613, N168, N319);
not NOT1 (N799, N791);
xor XOR2 (N800, N794, N572);
not NOT1 (N801, N785);
and AND3 (N802, N798, N299, N735);
or OR3 (N803, N790, N301, N401);
nor NOR2 (N804, N803, N164);
not NOT1 (N805, N802);
and AND3 (N806, N795, N619, N679);
nand NAND3 (N807, N801, N501, N532);
or OR2 (N808, N804, N461);
xor XOR2 (N809, N806, N209);
nor NOR2 (N810, N788, N705);
and AND2 (N811, N799, N699);
buf BUF1 (N812, N807);
nand NAND3 (N813, N812, N371, N273);
nand NAND4 (N814, N811, N805, N495, N145);
or OR4 (N815, N680, N151, N365, N481);
nor NOR2 (N816, N810, N594);
nand NAND2 (N817, N813, N4);
and AND2 (N818, N815, N673);
xor XOR2 (N819, N818, N221);
and AND2 (N820, N797, N349);
and AND4 (N821, N816, N311, N484, N302);
not NOT1 (N822, N808);
and AND3 (N823, N809, N230, N370);
nand NAND2 (N824, N823, N165);
and AND3 (N825, N821, N262, N128);
nor NOR4 (N826, N824, N501, N589, N553);
nor NOR4 (N827, N826, N246, N291, N222);
xor XOR2 (N828, N825, N638);
and AND3 (N829, N800, N104, N498);
or OR2 (N830, N782, N586);
not NOT1 (N831, N814);
or OR4 (N832, N828, N594, N198, N572);
not NOT1 (N833, N817);
nor NOR4 (N834, N833, N405, N761, N363);
nand NAND4 (N835, N829, N15, N215, N394);
and AND4 (N836, N820, N270, N578, N793);
xor XOR2 (N837, N832, N718);
xor XOR2 (N838, N827, N41);
nor NOR2 (N839, N796, N47);
or OR2 (N840, N831, N315);
nor NOR3 (N841, N838, N504, N683);
and AND2 (N842, N840, N4);
xor XOR2 (N843, N822, N206);
nand NAND4 (N844, N843, N415, N200, N18);
nand NAND3 (N845, N841, N507, N59);
buf BUF1 (N846, N830);
not NOT1 (N847, N819);
and AND2 (N848, N844, N44);
xor XOR2 (N849, N836, N403);
nor NOR3 (N850, N846, N47, N441);
not NOT1 (N851, N847);
nor NOR4 (N852, N839, N335, N768, N593);
nand NAND4 (N853, N850, N375, N602, N815);
xor XOR2 (N854, N842, N586);
nor NOR2 (N855, N848, N369);
buf BUF1 (N856, N849);
or OR4 (N857, N854, N347, N35, N95);
and AND4 (N858, N853, N278, N465, N244);
xor XOR2 (N859, N858, N414);
xor XOR2 (N860, N851, N783);
or OR4 (N861, N845, N680, N298, N640);
nand NAND2 (N862, N859, N554);
buf BUF1 (N863, N852);
buf BUF1 (N864, N860);
not NOT1 (N865, N861);
xor XOR2 (N866, N856, N337);
xor XOR2 (N867, N835, N513);
xor XOR2 (N868, N867, N653);
xor XOR2 (N869, N865, N765);
not NOT1 (N870, N864);
or OR4 (N871, N866, N150, N85, N627);
not NOT1 (N872, N834);
or OR3 (N873, N869, N428, N459);
not NOT1 (N874, N837);
or OR3 (N875, N863, N554, N410);
buf BUF1 (N876, N868);
buf BUF1 (N877, N872);
not NOT1 (N878, N870);
or OR4 (N879, N878, N179, N796, N400);
or OR2 (N880, N855, N428);
and AND4 (N881, N857, N655, N505, N428);
buf BUF1 (N882, N877);
not NOT1 (N883, N874);
nand NAND2 (N884, N875, N448);
nor NOR2 (N885, N883, N227);
nand NAND4 (N886, N871, N679, N557, N250);
nand NAND4 (N887, N881, N573, N327, N830);
and AND3 (N888, N873, N424, N50);
xor XOR2 (N889, N880, N635);
and AND2 (N890, N886, N448);
buf BUF1 (N891, N889);
and AND3 (N892, N885, N694, N465);
and AND4 (N893, N891, N142, N523, N107);
nand NAND4 (N894, N888, N598, N601, N176);
buf BUF1 (N895, N876);
not NOT1 (N896, N879);
buf BUF1 (N897, N895);
and AND3 (N898, N893, N440, N760);
or OR4 (N899, N890, N265, N552, N89);
nand NAND4 (N900, N897, N567, N507, N67);
nand NAND2 (N901, N898, N714);
and AND4 (N902, N901, N519, N44, N472);
buf BUF1 (N903, N899);
or OR3 (N904, N887, N519, N568);
nand NAND2 (N905, N882, N224);
and AND3 (N906, N903, N700, N147);
nand NAND3 (N907, N884, N327, N690);
and AND4 (N908, N896, N411, N818, N439);
buf BUF1 (N909, N894);
and AND4 (N910, N904, N544, N614, N891);
not NOT1 (N911, N900);
nand NAND2 (N912, N910, N161);
buf BUF1 (N913, N909);
buf BUF1 (N914, N907);
nor NOR2 (N915, N913, N271);
xor XOR2 (N916, N911, N825);
not NOT1 (N917, N912);
not NOT1 (N918, N906);
nor NOR4 (N919, N916, N747, N804, N494);
not NOT1 (N920, N902);
or OR4 (N921, N915, N531, N147, N101);
nand NAND4 (N922, N918, N447, N918, N806);
buf BUF1 (N923, N908);
nand NAND2 (N924, N914, N42);
nor NOR3 (N925, N924, N462, N209);
nand NAND2 (N926, N925, N394);
nand NAND2 (N927, N917, N795);
not NOT1 (N928, N926);
not NOT1 (N929, N919);
nor NOR2 (N930, N892, N718);
and AND2 (N931, N928, N252);
or OR3 (N932, N920, N188, N529);
nor NOR4 (N933, N932, N838, N811, N806);
not NOT1 (N934, N927);
nand NAND2 (N935, N921, N359);
not NOT1 (N936, N931);
not NOT1 (N937, N905);
and AND4 (N938, N922, N35, N223, N269);
and AND4 (N939, N934, N461, N689, N364);
or OR2 (N940, N939, N25);
xor XOR2 (N941, N862, N67);
buf BUF1 (N942, N935);
nand NAND4 (N943, N930, N178, N320, N310);
not NOT1 (N944, N929);
not NOT1 (N945, N944);
and AND4 (N946, N933, N161, N143, N367);
and AND2 (N947, N936, N13);
not NOT1 (N948, N923);
buf BUF1 (N949, N947);
or OR4 (N950, N937, N372, N517, N675);
buf BUF1 (N951, N938);
or OR3 (N952, N951, N56, N374);
nor NOR3 (N953, N950, N108, N144);
or OR4 (N954, N946, N874, N775, N475);
nand NAND2 (N955, N952, N645);
nor NOR3 (N956, N949, N719, N345);
buf BUF1 (N957, N956);
nand NAND3 (N958, N945, N912, N808);
or OR2 (N959, N958, N539);
and AND4 (N960, N955, N289, N699, N222);
xor XOR2 (N961, N957, N254);
not NOT1 (N962, N959);
nor NOR4 (N963, N960, N30, N873, N906);
buf BUF1 (N964, N962);
and AND3 (N965, N954, N711, N505);
not NOT1 (N966, N964);
or OR2 (N967, N965, N127);
and AND4 (N968, N940, N272, N625, N19);
and AND2 (N969, N961, N923);
xor XOR2 (N970, N943, N312);
or OR3 (N971, N953, N155, N869);
xor XOR2 (N972, N948, N668);
and AND3 (N973, N972, N364, N891);
and AND3 (N974, N973, N296, N124);
and AND3 (N975, N969, N525, N880);
and AND2 (N976, N942, N891);
nor NOR2 (N977, N975, N936);
not NOT1 (N978, N974);
not NOT1 (N979, N941);
not NOT1 (N980, N979);
nor NOR4 (N981, N963, N456, N675, N73);
not NOT1 (N982, N980);
buf BUF1 (N983, N982);
or OR3 (N984, N977, N633, N126);
and AND3 (N985, N967, N723, N827);
buf BUF1 (N986, N971);
or OR4 (N987, N986, N885, N278, N123);
nand NAND2 (N988, N981, N381);
or OR2 (N989, N976, N576);
and AND3 (N990, N983, N510, N10);
buf BUF1 (N991, N985);
nand NAND2 (N992, N966, N822);
not NOT1 (N993, N992);
nor NOR2 (N994, N993, N796);
buf BUF1 (N995, N989);
buf BUF1 (N996, N987);
nor NOR3 (N997, N988, N405, N493);
xor XOR2 (N998, N995, N121);
xor XOR2 (N999, N996, N659);
not NOT1 (N1000, N998);
or OR2 (N1001, N994, N498);
nand NAND4 (N1002, N997, N865, N842, N172);
nand NAND2 (N1003, N990, N574);
buf BUF1 (N1004, N1003);
and AND2 (N1005, N1001, N977);
xor XOR2 (N1006, N968, N542);
or OR4 (N1007, N970, N207, N817, N599);
nor NOR3 (N1008, N984, N10, N1002);
buf BUF1 (N1009, N76);
xor XOR2 (N1010, N1009, N568);
nor NOR2 (N1011, N1008, N814);
xor XOR2 (N1012, N1010, N822);
not NOT1 (N1013, N999);
or OR3 (N1014, N991, N795, N979);
and AND3 (N1015, N1011, N701, N388);
nor NOR2 (N1016, N1015, N341);
or OR3 (N1017, N1000, N163, N692);
xor XOR2 (N1018, N1007, N316);
nor NOR4 (N1019, N1004, N532, N574, N427);
buf BUF1 (N1020, N1019);
or OR2 (N1021, N1012, N945);
xor XOR2 (N1022, N1016, N455);
buf BUF1 (N1023, N1021);
and AND4 (N1024, N1018, N965, N774, N85);
nor NOR4 (N1025, N1020, N222, N838, N317);
or OR2 (N1026, N1005, N390);
buf BUF1 (N1027, N1025);
buf BUF1 (N1028, N1006);
or OR3 (N1029, N1023, N552, N207);
or OR4 (N1030, N1028, N410, N792, N1);
or OR3 (N1031, N1030, N686, N343);
or OR4 (N1032, N1027, N676, N9, N544);
or OR4 (N1033, N1029, N396, N237, N377);
xor XOR2 (N1034, N1017, N654);
nand NAND2 (N1035, N1034, N581);
not NOT1 (N1036, N1022);
xor XOR2 (N1037, N978, N988);
nand NAND3 (N1038, N1033, N589, N71);
buf BUF1 (N1039, N1026);
buf BUF1 (N1040, N1031);
nor NOR4 (N1041, N1040, N957, N375, N526);
xor XOR2 (N1042, N1013, N355);
not NOT1 (N1043, N1037);
and AND3 (N1044, N1036, N317, N462);
buf BUF1 (N1045, N1038);
and AND4 (N1046, N1044, N199, N512, N49);
not NOT1 (N1047, N1043);
nor NOR4 (N1048, N1024, N617, N458, N286);
xor XOR2 (N1049, N1041, N776);
nor NOR4 (N1050, N1048, N635, N264, N688);
nand NAND4 (N1051, N1045, N625, N379, N110);
nor NOR4 (N1052, N1051, N1001, N767, N818);
buf BUF1 (N1053, N1032);
nand NAND2 (N1054, N1035, N54);
nand NAND4 (N1055, N1014, N441, N103, N295);
buf BUF1 (N1056, N1050);
xor XOR2 (N1057, N1055, N250);
not NOT1 (N1058, N1047);
buf BUF1 (N1059, N1046);
not NOT1 (N1060, N1052);
and AND4 (N1061, N1042, N602, N270, N305);
nor NOR2 (N1062, N1060, N362);
nand NAND2 (N1063, N1039, N74);
nor NOR4 (N1064, N1063, N781, N327, N410);
not NOT1 (N1065, N1059);
nor NOR3 (N1066, N1054, N512, N394);
buf BUF1 (N1067, N1066);
not NOT1 (N1068, N1049);
buf BUF1 (N1069, N1065);
buf BUF1 (N1070, N1068);
nand NAND2 (N1071, N1058, N265);
buf BUF1 (N1072, N1069);
xor XOR2 (N1073, N1071, N983);
nor NOR4 (N1074, N1073, N717, N139, N679);
nand NAND3 (N1075, N1053, N436, N755);
nand NAND2 (N1076, N1072, N769);
xor XOR2 (N1077, N1057, N526);
nor NOR4 (N1078, N1067, N552, N426, N48);
buf BUF1 (N1079, N1056);
buf BUF1 (N1080, N1074);
nand NAND3 (N1081, N1070, N841, N400);
xor XOR2 (N1082, N1075, N822);
or OR4 (N1083, N1076, N280, N364, N303);
and AND4 (N1084, N1083, N289, N821, N464);
nor NOR3 (N1085, N1081, N859, N418);
nor NOR4 (N1086, N1061, N296, N217, N332);
nand NAND3 (N1087, N1062, N573, N271);
or OR3 (N1088, N1064, N648, N766);
nor NOR3 (N1089, N1086, N684, N361);
buf BUF1 (N1090, N1087);
xor XOR2 (N1091, N1088, N941);
nor NOR3 (N1092, N1079, N57, N68);
nor NOR4 (N1093, N1084, N977, N875, N338);
buf BUF1 (N1094, N1092);
not NOT1 (N1095, N1093);
xor XOR2 (N1096, N1090, N122);
not NOT1 (N1097, N1095);
nand NAND2 (N1098, N1078, N444);
nand NAND2 (N1099, N1091, N602);
buf BUF1 (N1100, N1089);
buf BUF1 (N1101, N1098);
nor NOR3 (N1102, N1085, N186, N442);
xor XOR2 (N1103, N1080, N483);
buf BUF1 (N1104, N1094);
buf BUF1 (N1105, N1100);
xor XOR2 (N1106, N1101, N399);
xor XOR2 (N1107, N1077, N804);
or OR3 (N1108, N1105, N313, N565);
nor NOR4 (N1109, N1102, N600, N947, N926);
buf BUF1 (N1110, N1106);
xor XOR2 (N1111, N1108, N837);
and AND3 (N1112, N1107, N1045, N146);
nand NAND2 (N1113, N1111, N177);
not NOT1 (N1114, N1110);
buf BUF1 (N1115, N1103);
nand NAND2 (N1116, N1096, N779);
and AND3 (N1117, N1097, N57, N323);
and AND3 (N1118, N1109, N413, N849);
not NOT1 (N1119, N1113);
and AND2 (N1120, N1115, N789);
buf BUF1 (N1121, N1119);
buf BUF1 (N1122, N1120);
nor NOR4 (N1123, N1116, N635, N620, N856);
xor XOR2 (N1124, N1112, N744);
not NOT1 (N1125, N1122);
nor NOR4 (N1126, N1114, N650, N915, N1085);
not NOT1 (N1127, N1118);
xor XOR2 (N1128, N1127, N1125);
not NOT1 (N1129, N950);
or OR2 (N1130, N1124, N566);
nor NOR3 (N1131, N1126, N543, N367);
or OR2 (N1132, N1128, N1025);
and AND3 (N1133, N1082, N762, N140);
not NOT1 (N1134, N1099);
nor NOR4 (N1135, N1134, N239, N522, N690);
not NOT1 (N1136, N1104);
or OR4 (N1137, N1135, N250, N1057, N926);
or OR3 (N1138, N1137, N1034, N741);
buf BUF1 (N1139, N1131);
nand NAND3 (N1140, N1136, N747, N514);
and AND3 (N1141, N1139, N638, N1049);
and AND4 (N1142, N1129, N882, N332, N778);
buf BUF1 (N1143, N1123);
nor NOR2 (N1144, N1141, N533);
or OR2 (N1145, N1121, N762);
or OR2 (N1146, N1143, N671);
and AND3 (N1147, N1133, N506, N108);
buf BUF1 (N1148, N1138);
buf BUF1 (N1149, N1145);
nor NOR4 (N1150, N1117, N1114, N293, N693);
buf BUF1 (N1151, N1132);
not NOT1 (N1152, N1148);
xor XOR2 (N1153, N1152, N1045);
xor XOR2 (N1154, N1151, N301);
and AND4 (N1155, N1153, N758, N85, N565);
nand NAND4 (N1156, N1147, N376, N1058, N587);
nor NOR3 (N1157, N1144, N352, N1099);
not NOT1 (N1158, N1142);
xor XOR2 (N1159, N1154, N749);
and AND3 (N1160, N1140, N513, N95);
nand NAND3 (N1161, N1155, N751, N286);
or OR4 (N1162, N1161, N449, N834, N364);
xor XOR2 (N1163, N1149, N1060);
buf BUF1 (N1164, N1162);
and AND2 (N1165, N1160, N837);
nand NAND4 (N1166, N1158, N640, N741, N221);
and AND4 (N1167, N1164, N127, N552, N179);
not NOT1 (N1168, N1150);
and AND4 (N1169, N1157, N699, N666, N878);
or OR4 (N1170, N1156, N54, N873, N1052);
xor XOR2 (N1171, N1159, N377);
not NOT1 (N1172, N1165);
not NOT1 (N1173, N1168);
nand NAND3 (N1174, N1171, N774, N853);
nor NOR4 (N1175, N1130, N382, N554, N282);
and AND4 (N1176, N1167, N857, N1011, N1136);
buf BUF1 (N1177, N1170);
nor NOR4 (N1178, N1176, N1022, N686, N879);
or OR4 (N1179, N1172, N1131, N241, N609);
nand NAND2 (N1180, N1163, N393);
and AND4 (N1181, N1175, N1136, N568, N31);
xor XOR2 (N1182, N1146, N656);
nor NOR3 (N1183, N1169, N917, N318);
xor XOR2 (N1184, N1177, N445);
buf BUF1 (N1185, N1180);
nor NOR3 (N1186, N1173, N857, N1023);
and AND3 (N1187, N1174, N1185, N561);
xor XOR2 (N1188, N134, N530);
and AND2 (N1189, N1178, N54);
nand NAND2 (N1190, N1182, N568);
buf BUF1 (N1191, N1186);
and AND3 (N1192, N1190, N655, N709);
not NOT1 (N1193, N1184);
xor XOR2 (N1194, N1188, N285);
xor XOR2 (N1195, N1192, N112);
and AND3 (N1196, N1189, N264, N530);
not NOT1 (N1197, N1195);
or OR2 (N1198, N1197, N1150);
not NOT1 (N1199, N1194);
xor XOR2 (N1200, N1191, N713);
not NOT1 (N1201, N1198);
or OR3 (N1202, N1183, N273, N1110);
buf BUF1 (N1203, N1187);
nand NAND4 (N1204, N1199, N309, N1116, N192);
or OR2 (N1205, N1203, N303);
and AND4 (N1206, N1202, N1088, N611, N804);
and AND2 (N1207, N1204, N257);
nand NAND4 (N1208, N1201, N439, N1039, N1171);
or OR4 (N1209, N1166, N677, N1050, N946);
or OR2 (N1210, N1207, N102);
buf BUF1 (N1211, N1181);
nor NOR2 (N1212, N1196, N262);
nor NOR4 (N1213, N1209, N17, N906, N835);
and AND4 (N1214, N1200, N547, N280, N747);
not NOT1 (N1215, N1214);
and AND2 (N1216, N1193, N868);
or OR3 (N1217, N1212, N324, N861);
and AND3 (N1218, N1210, N180, N132);
or OR3 (N1219, N1179, N1170, N400);
nor NOR2 (N1220, N1216, N922);
xor XOR2 (N1221, N1219, N417);
buf BUF1 (N1222, N1217);
or OR3 (N1223, N1218, N226, N217);
not NOT1 (N1224, N1208);
xor XOR2 (N1225, N1224, N207);
buf BUF1 (N1226, N1221);
not NOT1 (N1227, N1211);
nand NAND4 (N1228, N1206, N1038, N1128, N945);
nand NAND4 (N1229, N1223, N1062, N1210, N286);
nor NOR3 (N1230, N1220, N29, N1127);
xor XOR2 (N1231, N1227, N217);
or OR2 (N1232, N1213, N602);
xor XOR2 (N1233, N1230, N1014);
buf BUF1 (N1234, N1215);
or OR3 (N1235, N1234, N85, N328);
not NOT1 (N1236, N1225);
and AND2 (N1237, N1235, N500);
not NOT1 (N1238, N1222);
nand NAND4 (N1239, N1233, N1011, N586, N566);
not NOT1 (N1240, N1238);
or OR3 (N1241, N1231, N825, N465);
nor NOR4 (N1242, N1205, N902, N551, N482);
or OR4 (N1243, N1229, N986, N46, N352);
or OR2 (N1244, N1237, N1064);
and AND4 (N1245, N1232, N346, N95, N937);
or OR3 (N1246, N1243, N874, N168);
or OR3 (N1247, N1228, N76, N276);
not NOT1 (N1248, N1247);
or OR4 (N1249, N1240, N107, N395, N1183);
or OR2 (N1250, N1241, N350);
nand NAND4 (N1251, N1226, N1130, N282, N923);
xor XOR2 (N1252, N1244, N426);
nand NAND4 (N1253, N1242, N34, N466, N119);
xor XOR2 (N1254, N1248, N78);
xor XOR2 (N1255, N1239, N198);
not NOT1 (N1256, N1245);
and AND2 (N1257, N1246, N1256);
nor NOR3 (N1258, N739, N2, N196);
not NOT1 (N1259, N1254);
and AND4 (N1260, N1258, N1079, N372, N887);
and AND2 (N1261, N1252, N798);
buf BUF1 (N1262, N1251);
buf BUF1 (N1263, N1261);
or OR4 (N1264, N1260, N564, N394, N479);
nand NAND4 (N1265, N1250, N419, N664, N711);
nand NAND4 (N1266, N1263, N1215, N310, N745);
nand NAND3 (N1267, N1255, N57, N1129);
or OR2 (N1268, N1265, N507);
xor XOR2 (N1269, N1249, N1254);
nor NOR3 (N1270, N1253, N1224, N1192);
nor NOR4 (N1271, N1267, N1081, N292, N809);
not NOT1 (N1272, N1269);
and AND4 (N1273, N1268, N1261, N323, N1252);
nor NOR3 (N1274, N1257, N770, N925);
not NOT1 (N1275, N1264);
nand NAND3 (N1276, N1274, N670, N997);
or OR2 (N1277, N1271, N823);
and AND2 (N1278, N1270, N229);
xor XOR2 (N1279, N1278, N1217);
buf BUF1 (N1280, N1275);
nor NOR4 (N1281, N1262, N797, N402, N1234);
or OR2 (N1282, N1259, N225);
buf BUF1 (N1283, N1282);
and AND4 (N1284, N1273, N136, N441, N172);
or OR4 (N1285, N1284, N1161, N382, N217);
not NOT1 (N1286, N1279);
nor NOR2 (N1287, N1280, N310);
nor NOR2 (N1288, N1272, N422);
or OR3 (N1289, N1277, N314, N1238);
nor NOR2 (N1290, N1281, N1098);
and AND3 (N1291, N1287, N491, N622);
nand NAND3 (N1292, N1286, N695, N147);
and AND4 (N1293, N1290, N659, N1247, N819);
xor XOR2 (N1294, N1289, N1090);
xor XOR2 (N1295, N1283, N401);
nor NOR3 (N1296, N1236, N650, N272);
xor XOR2 (N1297, N1293, N147);
buf BUF1 (N1298, N1297);
buf BUF1 (N1299, N1291);
xor XOR2 (N1300, N1292, N363);
nor NOR4 (N1301, N1298, N1000, N871, N492);
xor XOR2 (N1302, N1295, N326);
nor NOR2 (N1303, N1301, N379);
and AND4 (N1304, N1299, N1043, N465, N743);
buf BUF1 (N1305, N1294);
nand NAND2 (N1306, N1303, N926);
not NOT1 (N1307, N1305);
or OR3 (N1308, N1302, N1187, N833);
nand NAND2 (N1309, N1288, N1013);
not NOT1 (N1310, N1309);
not NOT1 (N1311, N1276);
nand NAND2 (N1312, N1304, N1237);
buf BUF1 (N1313, N1296);
nor NOR3 (N1314, N1312, N967, N398);
buf BUF1 (N1315, N1310);
nand NAND2 (N1316, N1285, N1212);
nor NOR4 (N1317, N1315, N1180, N736, N232);
nand NAND2 (N1318, N1313, N542);
buf BUF1 (N1319, N1300);
and AND2 (N1320, N1316, N1009);
xor XOR2 (N1321, N1266, N852);
not NOT1 (N1322, N1318);
and AND4 (N1323, N1317, N875, N375, N968);
nor NOR2 (N1324, N1308, N1186);
nand NAND3 (N1325, N1319, N1088, N1222);
not NOT1 (N1326, N1314);
nand NAND2 (N1327, N1326, N168);
or OR3 (N1328, N1306, N845, N675);
nor NOR3 (N1329, N1307, N790, N157);
not NOT1 (N1330, N1325);
or OR2 (N1331, N1328, N1115);
buf BUF1 (N1332, N1331);
nand NAND3 (N1333, N1330, N560, N834);
not NOT1 (N1334, N1332);
nor NOR2 (N1335, N1322, N301);
nand NAND2 (N1336, N1320, N120);
and AND3 (N1337, N1336, N1289, N490);
nand NAND3 (N1338, N1323, N198, N742);
and AND4 (N1339, N1327, N385, N663, N751);
nor NOR3 (N1340, N1339, N1326, N1184);
nor NOR4 (N1341, N1311, N1003, N829, N636);
nand NAND2 (N1342, N1329, N1215);
and AND3 (N1343, N1338, N701, N456);
nand NAND3 (N1344, N1340, N838, N258);
nand NAND3 (N1345, N1343, N484, N909);
nor NOR4 (N1346, N1341, N92, N932, N719);
xor XOR2 (N1347, N1335, N269);
and AND3 (N1348, N1345, N714, N1319);
or OR4 (N1349, N1347, N872, N528, N903);
xor XOR2 (N1350, N1321, N1052);
or OR3 (N1351, N1342, N733, N1009);
nor NOR2 (N1352, N1351, N1095);
nand NAND2 (N1353, N1333, N1294);
or OR2 (N1354, N1349, N21);
buf BUF1 (N1355, N1348);
or OR2 (N1356, N1337, N608);
not NOT1 (N1357, N1344);
xor XOR2 (N1358, N1346, N1203);
and AND2 (N1359, N1357, N988);
buf BUF1 (N1360, N1359);
not NOT1 (N1361, N1324);
or OR4 (N1362, N1354, N1285, N201, N492);
nor NOR3 (N1363, N1352, N150, N731);
or OR2 (N1364, N1361, N427);
not NOT1 (N1365, N1334);
not NOT1 (N1366, N1353);
not NOT1 (N1367, N1360);
xor XOR2 (N1368, N1363, N206);
nor NOR2 (N1369, N1367, N1115);
or OR4 (N1370, N1368, N560, N486, N1033);
xor XOR2 (N1371, N1350, N601);
buf BUF1 (N1372, N1362);
xor XOR2 (N1373, N1372, N834);
buf BUF1 (N1374, N1365);
or OR3 (N1375, N1371, N17, N269);
and AND4 (N1376, N1366, N1040, N442, N25);
not NOT1 (N1377, N1370);
or OR3 (N1378, N1376, N112, N547);
not NOT1 (N1379, N1377);
buf BUF1 (N1380, N1364);
nand NAND2 (N1381, N1373, N829);
and AND3 (N1382, N1369, N358, N1025);
not NOT1 (N1383, N1358);
or OR2 (N1384, N1383, N896);
and AND3 (N1385, N1382, N128, N819);
nor NOR3 (N1386, N1356, N275, N196);
and AND4 (N1387, N1385, N558, N1365, N491);
nor NOR2 (N1388, N1379, N1233);
xor XOR2 (N1389, N1387, N208);
or OR3 (N1390, N1381, N1016, N778);
xor XOR2 (N1391, N1375, N181);
nand NAND3 (N1392, N1374, N748, N897);
xor XOR2 (N1393, N1355, N866);
nand NAND4 (N1394, N1389, N779, N377, N745);
not NOT1 (N1395, N1393);
not NOT1 (N1396, N1390);
or OR2 (N1397, N1396, N29);
nor NOR2 (N1398, N1397, N879);
nor NOR4 (N1399, N1388, N618, N701, N1054);
or OR3 (N1400, N1380, N884, N214);
nor NOR4 (N1401, N1394, N406, N353, N1124);
nand NAND3 (N1402, N1399, N1128, N57);
nor NOR4 (N1403, N1402, N1225, N1117, N239);
or OR2 (N1404, N1400, N922);
xor XOR2 (N1405, N1391, N1217);
nor NOR4 (N1406, N1392, N493, N215, N933);
xor XOR2 (N1407, N1403, N748);
buf BUF1 (N1408, N1395);
not NOT1 (N1409, N1398);
buf BUF1 (N1410, N1409);
and AND4 (N1411, N1410, N494, N251, N1101);
or OR3 (N1412, N1378, N173, N394);
nand NAND2 (N1413, N1411, N411);
nand NAND3 (N1414, N1407, N111, N645);
and AND3 (N1415, N1412, N1356, N206);
and AND4 (N1416, N1413, N14, N462, N736);
buf BUF1 (N1417, N1404);
nand NAND2 (N1418, N1384, N1065);
not NOT1 (N1419, N1405);
or OR2 (N1420, N1401, N494);
xor XOR2 (N1421, N1386, N424);
and AND2 (N1422, N1417, N1171);
buf BUF1 (N1423, N1408);
nand NAND4 (N1424, N1422, N1041, N266, N53);
nand NAND3 (N1425, N1418, N751, N296);
or OR4 (N1426, N1425, N1351, N1359, N702);
xor XOR2 (N1427, N1414, N778);
and AND4 (N1428, N1426, N955, N424, N907);
or OR2 (N1429, N1424, N603);
nand NAND2 (N1430, N1420, N654);
nor NOR2 (N1431, N1428, N1160);
nand NAND4 (N1432, N1429, N183, N678, N1216);
nand NAND3 (N1433, N1423, N663, N1335);
not NOT1 (N1434, N1432);
or OR3 (N1435, N1406, N605, N1291);
nor NOR3 (N1436, N1415, N253, N1173);
buf BUF1 (N1437, N1431);
and AND4 (N1438, N1434, N1145, N1208, N1403);
xor XOR2 (N1439, N1419, N1079);
nor NOR2 (N1440, N1416, N771);
nor NOR4 (N1441, N1421, N1327, N1310, N1028);
xor XOR2 (N1442, N1441, N966);
xor XOR2 (N1443, N1442, N13);
nor NOR4 (N1444, N1440, N370, N984, N437);
xor XOR2 (N1445, N1430, N575);
not NOT1 (N1446, N1435);
nand NAND3 (N1447, N1437, N294, N818);
nand NAND3 (N1448, N1436, N222, N555);
and AND4 (N1449, N1446, N1145, N1344, N927);
xor XOR2 (N1450, N1449, N35);
nor NOR4 (N1451, N1448, N267, N1071, N205);
nor NOR3 (N1452, N1444, N199, N384);
or OR4 (N1453, N1443, N948, N1139, N253);
not NOT1 (N1454, N1452);
or OR2 (N1455, N1454, N301);
nor NOR3 (N1456, N1451, N5, N1003);
buf BUF1 (N1457, N1427);
xor XOR2 (N1458, N1433, N1313);
nor NOR2 (N1459, N1453, N845);
and AND4 (N1460, N1439, N1250, N1077, N1250);
nor NOR3 (N1461, N1460, N510, N120);
nand NAND2 (N1462, N1457, N941);
buf BUF1 (N1463, N1445);
nor NOR2 (N1464, N1461, N8);
or OR3 (N1465, N1464, N471, N1398);
not NOT1 (N1466, N1455);
nor NOR2 (N1467, N1465, N1023);
and AND3 (N1468, N1458, N442, N1178);
or OR3 (N1469, N1467, N951, N1323);
or OR4 (N1470, N1447, N131, N228, N578);
not NOT1 (N1471, N1468);
or OR4 (N1472, N1450, N1174, N1423, N742);
nand NAND4 (N1473, N1471, N1248, N644, N107);
xor XOR2 (N1474, N1470, N1336);
or OR4 (N1475, N1438, N32, N1286, N651);
nand NAND2 (N1476, N1456, N538);
buf BUF1 (N1477, N1473);
or OR3 (N1478, N1469, N602, N181);
not NOT1 (N1479, N1477);
nor NOR3 (N1480, N1466, N1210, N49);
nand NAND3 (N1481, N1478, N605, N32);
xor XOR2 (N1482, N1474, N258);
or OR4 (N1483, N1462, N595, N891, N200);
buf BUF1 (N1484, N1483);
nand NAND4 (N1485, N1459, N1033, N913, N78);
buf BUF1 (N1486, N1481);
buf BUF1 (N1487, N1486);
nor NOR3 (N1488, N1487, N804, N1296);
xor XOR2 (N1489, N1488, N1254);
xor XOR2 (N1490, N1480, N887);
buf BUF1 (N1491, N1489);
nor NOR4 (N1492, N1490, N704, N502, N30);
not NOT1 (N1493, N1492);
not NOT1 (N1494, N1484);
nand NAND2 (N1495, N1476, N777);
nor NOR4 (N1496, N1472, N280, N1207, N799);
or OR2 (N1497, N1463, N124);
not NOT1 (N1498, N1493);
nand NAND3 (N1499, N1495, N217, N1298);
buf BUF1 (N1500, N1498);
xor XOR2 (N1501, N1482, N852);
nor NOR3 (N1502, N1497, N339, N191);
nor NOR2 (N1503, N1501, N32);
xor XOR2 (N1504, N1503, N990);
nor NOR2 (N1505, N1500, N734);
nand NAND2 (N1506, N1494, N1439);
nand NAND3 (N1507, N1502, N915, N241);
and AND4 (N1508, N1507, N544, N993, N233);
not NOT1 (N1509, N1475);
xor XOR2 (N1510, N1485, N587);
xor XOR2 (N1511, N1496, N1077);
nand NAND3 (N1512, N1508, N958, N1508);
not NOT1 (N1513, N1479);
xor XOR2 (N1514, N1510, N738);
or OR2 (N1515, N1505, N662);
and AND4 (N1516, N1514, N446, N672, N1487);
xor XOR2 (N1517, N1506, N932);
buf BUF1 (N1518, N1499);
buf BUF1 (N1519, N1512);
buf BUF1 (N1520, N1491);
nand NAND4 (N1521, N1518, N1403, N948, N1242);
not NOT1 (N1522, N1521);
not NOT1 (N1523, N1515);
nor NOR2 (N1524, N1513, N234);
not NOT1 (N1525, N1509);
buf BUF1 (N1526, N1517);
not NOT1 (N1527, N1504);
xor XOR2 (N1528, N1525, N688);
nand NAND3 (N1529, N1519, N1371, N795);
nand NAND4 (N1530, N1528, N946, N1052, N596);
xor XOR2 (N1531, N1527, N857);
and AND2 (N1532, N1524, N1324);
nor NOR4 (N1533, N1522, N608, N1451, N654);
nor NOR3 (N1534, N1531, N728, N1431);
buf BUF1 (N1535, N1530);
or OR3 (N1536, N1520, N1080, N886);
and AND2 (N1537, N1536, N690);
nor NOR4 (N1538, N1535, N857, N580, N605);
xor XOR2 (N1539, N1523, N863);
buf BUF1 (N1540, N1516);
or OR4 (N1541, N1529, N69, N514, N1250);
or OR2 (N1542, N1511, N600);
not NOT1 (N1543, N1541);
xor XOR2 (N1544, N1542, N1510);
nand NAND2 (N1545, N1533, N51);
not NOT1 (N1546, N1537);
buf BUF1 (N1547, N1545);
and AND2 (N1548, N1540, N266);
nor NOR2 (N1549, N1532, N867);
not NOT1 (N1550, N1539);
nor NOR2 (N1551, N1544, N117);
xor XOR2 (N1552, N1549, N391);
buf BUF1 (N1553, N1551);
nand NAND4 (N1554, N1534, N152, N1171, N274);
not NOT1 (N1555, N1552);
nand NAND3 (N1556, N1543, N357, N471);
buf BUF1 (N1557, N1550);
not NOT1 (N1558, N1555);
or OR3 (N1559, N1538, N278, N522);
nand NAND2 (N1560, N1554, N13);
xor XOR2 (N1561, N1559, N1338);
or OR2 (N1562, N1553, N555);
buf BUF1 (N1563, N1556);
buf BUF1 (N1564, N1561);
buf BUF1 (N1565, N1558);
not NOT1 (N1566, N1547);
nand NAND4 (N1567, N1557, N1428, N484, N351);
nand NAND4 (N1568, N1566, N1151, N682, N1034);
nor NOR4 (N1569, N1564, N730, N457, N991);
nand NAND3 (N1570, N1546, N842, N728);
buf BUF1 (N1571, N1560);
xor XOR2 (N1572, N1567, N1473);
and AND2 (N1573, N1562, N1148);
nor NOR4 (N1574, N1569, N971, N979, N871);
or OR4 (N1575, N1563, N263, N1120, N948);
not NOT1 (N1576, N1572);
or OR4 (N1577, N1574, N182, N161, N1346);
buf BUF1 (N1578, N1573);
or OR2 (N1579, N1575, N610);
nor NOR3 (N1580, N1579, N446, N981);
nor NOR3 (N1581, N1548, N1309, N1123);
nand NAND3 (N1582, N1565, N692, N908);
buf BUF1 (N1583, N1578);
and AND4 (N1584, N1581, N601, N53, N1213);
or OR2 (N1585, N1580, N1464);
buf BUF1 (N1586, N1570);
and AND4 (N1587, N1577, N657, N394, N97);
not NOT1 (N1588, N1571);
xor XOR2 (N1589, N1576, N180);
nor NOR4 (N1590, N1589, N1310, N734, N85);
nand NAND2 (N1591, N1584, N270);
not NOT1 (N1592, N1591);
nor NOR3 (N1593, N1582, N132, N1559);
nor NOR2 (N1594, N1568, N927);
or OR4 (N1595, N1592, N1111, N1176, N466);
nand NAND3 (N1596, N1588, N1208, N67);
or OR3 (N1597, N1596, N838, N1096);
and AND4 (N1598, N1526, N1039, N712, N1116);
nand NAND2 (N1599, N1597, N708);
buf BUF1 (N1600, N1586);
nor NOR4 (N1601, N1590, N1216, N210, N615);
nand NAND2 (N1602, N1594, N86);
not NOT1 (N1603, N1593);
not NOT1 (N1604, N1598);
and AND4 (N1605, N1604, N725, N925, N71);
xor XOR2 (N1606, N1583, N1313);
buf BUF1 (N1607, N1606);
not NOT1 (N1608, N1585);
buf BUF1 (N1609, N1608);
buf BUF1 (N1610, N1595);
xor XOR2 (N1611, N1607, N960);
buf BUF1 (N1612, N1605);
nand NAND4 (N1613, N1612, N576, N888, N982);
nand NAND3 (N1614, N1613, N332, N1157);
and AND4 (N1615, N1587, N414, N109, N858);
or OR2 (N1616, N1601, N1443);
or OR3 (N1617, N1610, N1593, N198);
nand NAND2 (N1618, N1600, N895);
or OR3 (N1619, N1599, N1208, N415);
xor XOR2 (N1620, N1611, N446);
and AND4 (N1621, N1619, N1004, N1001, N1170);
nand NAND3 (N1622, N1609, N1506, N1502);
nor NOR2 (N1623, N1614, N1167);
not NOT1 (N1624, N1602);
and AND2 (N1625, N1624, N1250);
nor NOR2 (N1626, N1622, N396);
xor XOR2 (N1627, N1623, N1423);
nand NAND2 (N1628, N1603, N1060);
buf BUF1 (N1629, N1626);
nor NOR2 (N1630, N1615, N1134);
not NOT1 (N1631, N1620);
and AND4 (N1632, N1617, N1173, N505, N1112);
nand NAND4 (N1633, N1625, N640, N1386, N1235);
xor XOR2 (N1634, N1628, N1559);
or OR2 (N1635, N1618, N880);
and AND2 (N1636, N1634, N695);
xor XOR2 (N1637, N1633, N1469);
or OR3 (N1638, N1631, N1312, N1344);
not NOT1 (N1639, N1629);
buf BUF1 (N1640, N1639);
xor XOR2 (N1641, N1621, N625);
or OR2 (N1642, N1630, N886);
not NOT1 (N1643, N1636);
or OR4 (N1644, N1637, N350, N1470, N734);
or OR3 (N1645, N1616, N1306, N548);
nor NOR2 (N1646, N1645, N466);
or OR2 (N1647, N1627, N588);
nand NAND3 (N1648, N1643, N1201, N1318);
and AND4 (N1649, N1632, N49, N929, N233);
xor XOR2 (N1650, N1641, N146);
nand NAND4 (N1651, N1640, N414, N376, N1111);
xor XOR2 (N1652, N1649, N117);
xor XOR2 (N1653, N1648, N555);
not NOT1 (N1654, N1646);
or OR4 (N1655, N1638, N1056, N255, N324);
nand NAND4 (N1656, N1647, N1260, N432, N1370);
or OR4 (N1657, N1642, N22, N128, N101);
not NOT1 (N1658, N1657);
nand NAND3 (N1659, N1654, N792, N1247);
nor NOR3 (N1660, N1652, N273, N444);
and AND3 (N1661, N1653, N1625, N1247);
or OR3 (N1662, N1661, N398, N217);
not NOT1 (N1663, N1650);
nand NAND4 (N1664, N1659, N954, N365, N588);
nor NOR2 (N1665, N1663, N549);
and AND3 (N1666, N1651, N1521, N1432);
or OR3 (N1667, N1660, N1415, N542);
buf BUF1 (N1668, N1665);
nand NAND2 (N1669, N1664, N496);
xor XOR2 (N1670, N1668, N1052);
buf BUF1 (N1671, N1662);
nand NAND4 (N1672, N1658, N1605, N936, N1393);
or OR3 (N1673, N1671, N1130, N789);
xor XOR2 (N1674, N1655, N962);
xor XOR2 (N1675, N1673, N1043);
or OR4 (N1676, N1635, N606, N1614, N978);
and AND3 (N1677, N1672, N1638, N1555);
nand NAND4 (N1678, N1676, N829, N920, N982);
buf BUF1 (N1679, N1644);
buf BUF1 (N1680, N1674);
buf BUF1 (N1681, N1666);
not NOT1 (N1682, N1679);
nand NAND4 (N1683, N1670, N1050, N1237, N833);
or OR2 (N1684, N1675, N44);
not NOT1 (N1685, N1678);
and AND3 (N1686, N1669, N1295, N404);
nand NAND3 (N1687, N1682, N32, N863);
nand NAND4 (N1688, N1683, N1517, N1584, N775);
buf BUF1 (N1689, N1685);
or OR2 (N1690, N1687, N1573);
or OR3 (N1691, N1667, N724, N1614);
buf BUF1 (N1692, N1684);
nor NOR2 (N1693, N1680, N23);
buf BUF1 (N1694, N1693);
or OR2 (N1695, N1677, N546);
xor XOR2 (N1696, N1686, N1115);
nor NOR3 (N1697, N1694, N545, N222);
or OR4 (N1698, N1681, N1362, N507, N574);
nor NOR2 (N1699, N1656, N1478);
buf BUF1 (N1700, N1692);
not NOT1 (N1701, N1691);
nand NAND3 (N1702, N1688, N1022, N1247);
nand NAND4 (N1703, N1700, N1177, N215, N832);
nand NAND4 (N1704, N1699, N1682, N583, N1493);
nand NAND3 (N1705, N1702, N920, N1484);
or OR4 (N1706, N1696, N684, N769, N344);
or OR4 (N1707, N1701, N727, N640, N646);
xor XOR2 (N1708, N1690, N1083);
nor NOR3 (N1709, N1706, N1477, N1560);
and AND2 (N1710, N1689, N1620);
and AND3 (N1711, N1710, N744, N1256);
xor XOR2 (N1712, N1707, N1435);
not NOT1 (N1713, N1703);
not NOT1 (N1714, N1709);
or OR3 (N1715, N1698, N1530, N1505);
or OR2 (N1716, N1715, N437);
or OR2 (N1717, N1697, N531);
buf BUF1 (N1718, N1717);
nand NAND3 (N1719, N1712, N534, N1616);
or OR2 (N1720, N1714, N1681);
xor XOR2 (N1721, N1716, N1059);
and AND2 (N1722, N1720, N1482);
nand NAND3 (N1723, N1719, N793, N340);
and AND3 (N1724, N1705, N739, N1555);
nand NAND3 (N1725, N1713, N403, N1427);
or OR4 (N1726, N1724, N123, N1271, N479);
buf BUF1 (N1727, N1723);
buf BUF1 (N1728, N1721);
or OR3 (N1729, N1718, N1669, N1083);
not NOT1 (N1730, N1729);
not NOT1 (N1731, N1725);
and AND4 (N1732, N1704, N1212, N1187, N511);
xor XOR2 (N1733, N1730, N1084);
buf BUF1 (N1734, N1733);
xor XOR2 (N1735, N1695, N1673);
not NOT1 (N1736, N1727);
not NOT1 (N1737, N1734);
or OR2 (N1738, N1735, N84);
not NOT1 (N1739, N1728);
xor XOR2 (N1740, N1736, N661);
xor XOR2 (N1741, N1722, N431);
buf BUF1 (N1742, N1739);
buf BUF1 (N1743, N1737);
and AND3 (N1744, N1731, N138, N831);
nand NAND2 (N1745, N1711, N1314);
and AND3 (N1746, N1744, N263, N468);
nand NAND4 (N1747, N1743, N1523, N1647, N1344);
nor NOR3 (N1748, N1732, N1655, N315);
not NOT1 (N1749, N1745);
not NOT1 (N1750, N1742);
buf BUF1 (N1751, N1738);
and AND2 (N1752, N1740, N1534);
not NOT1 (N1753, N1750);
not NOT1 (N1754, N1748);
buf BUF1 (N1755, N1726);
nor NOR2 (N1756, N1755, N277);
not NOT1 (N1757, N1708);
nor NOR4 (N1758, N1754, N598, N1119, N415);
xor XOR2 (N1759, N1751, N1040);
xor XOR2 (N1760, N1747, N261);
not NOT1 (N1761, N1758);
xor XOR2 (N1762, N1749, N903);
and AND2 (N1763, N1753, N1442);
buf BUF1 (N1764, N1741);
buf BUF1 (N1765, N1762);
or OR4 (N1766, N1746, N833, N1674, N365);
nor NOR2 (N1767, N1764, N1685);
buf BUF1 (N1768, N1765);
nand NAND4 (N1769, N1752, N668, N1677, N529);
nand NAND2 (N1770, N1767, N140);
nor NOR4 (N1771, N1760, N1493, N213, N506);
nor NOR4 (N1772, N1771, N1473, N1592, N590);
or OR2 (N1773, N1759, N1453);
nor NOR4 (N1774, N1768, N1103, N269, N517);
not NOT1 (N1775, N1756);
and AND4 (N1776, N1757, N1510, N1699, N184);
and AND2 (N1777, N1773, N739);
buf BUF1 (N1778, N1761);
nor NOR2 (N1779, N1763, N512);
buf BUF1 (N1780, N1774);
nor NOR2 (N1781, N1770, N805);
or OR2 (N1782, N1776, N324);
nand NAND3 (N1783, N1780, N757, N36);
nand NAND3 (N1784, N1777, N782, N759);
xor XOR2 (N1785, N1769, N1546);
or OR4 (N1786, N1782, N953, N1186, N1551);
and AND4 (N1787, N1781, N190, N1564, N687);
and AND3 (N1788, N1766, N793, N1359);
or OR3 (N1789, N1785, N1543, N973);
xor XOR2 (N1790, N1775, N1159);
xor XOR2 (N1791, N1779, N1721);
or OR3 (N1792, N1790, N947, N570);
buf BUF1 (N1793, N1772);
or OR3 (N1794, N1786, N970, N855);
nor NOR3 (N1795, N1794, N1153, N1458);
nand NAND2 (N1796, N1795, N622);
not NOT1 (N1797, N1787);
and AND2 (N1798, N1791, N1223);
or OR4 (N1799, N1784, N1377, N1147, N897);
buf BUF1 (N1800, N1798);
and AND3 (N1801, N1793, N1229, N1756);
xor XOR2 (N1802, N1800, N1414);
not NOT1 (N1803, N1796);
buf BUF1 (N1804, N1783);
nor NOR3 (N1805, N1789, N784, N797);
and AND3 (N1806, N1799, N968, N960);
nor NOR3 (N1807, N1804, N421, N953);
and AND2 (N1808, N1797, N793);
or OR2 (N1809, N1778, N1309);
not NOT1 (N1810, N1792);
not NOT1 (N1811, N1802);
and AND3 (N1812, N1808, N108, N426);
or OR4 (N1813, N1805, N865, N71, N387);
or OR2 (N1814, N1807, N1479);
nor NOR4 (N1815, N1810, N911, N1507, N1522);
nor NOR3 (N1816, N1811, N828, N1139);
buf BUF1 (N1817, N1815);
nand NAND4 (N1818, N1812, N834, N1678, N1120);
or OR4 (N1819, N1801, N525, N1426, N589);
buf BUF1 (N1820, N1809);
nand NAND3 (N1821, N1816, N111, N822);
xor XOR2 (N1822, N1803, N1073);
nand NAND3 (N1823, N1817, N698, N288);
nor NOR4 (N1824, N1814, N1128, N1048, N1330);
nand NAND4 (N1825, N1818, N1161, N826, N1822);
buf BUF1 (N1826, N1597);
not NOT1 (N1827, N1819);
xor XOR2 (N1828, N1823, N1781);
nand NAND4 (N1829, N1806, N1787, N424, N746);
not NOT1 (N1830, N1813);
nor NOR4 (N1831, N1821, N1747, N1483, N1100);
buf BUF1 (N1832, N1828);
nor NOR4 (N1833, N1827, N591, N121, N1424);
nand NAND3 (N1834, N1832, N132, N324);
or OR3 (N1835, N1830, N293, N58);
not NOT1 (N1836, N1835);
buf BUF1 (N1837, N1826);
and AND4 (N1838, N1834, N529, N979, N812);
buf BUF1 (N1839, N1831);
buf BUF1 (N1840, N1837);
nor NOR2 (N1841, N1833, N835);
buf BUF1 (N1842, N1788);
xor XOR2 (N1843, N1839, N401);
nand NAND2 (N1844, N1838, N409);
nand NAND4 (N1845, N1843, N1161, N1450, N1188);
not NOT1 (N1846, N1820);
nand NAND4 (N1847, N1825, N765, N130, N1368);
nor NOR3 (N1848, N1842, N619, N239);
or OR2 (N1849, N1840, N392);
and AND4 (N1850, N1844, N1029, N782, N643);
nor NOR2 (N1851, N1841, N1701);
nor NOR2 (N1852, N1824, N477);
and AND4 (N1853, N1849, N1213, N172, N692);
not NOT1 (N1854, N1851);
nor NOR2 (N1855, N1853, N520);
not NOT1 (N1856, N1850);
nor NOR3 (N1857, N1845, N1662, N1577);
xor XOR2 (N1858, N1846, N944);
nand NAND2 (N1859, N1856, N1643);
buf BUF1 (N1860, N1855);
nand NAND4 (N1861, N1848, N1146, N1328, N1663);
xor XOR2 (N1862, N1861, N1433);
or OR2 (N1863, N1860, N947);
nand NAND4 (N1864, N1863, N341, N759, N1437);
xor XOR2 (N1865, N1847, N888);
and AND4 (N1866, N1854, N356, N1449, N201);
xor XOR2 (N1867, N1857, N287);
nand NAND2 (N1868, N1867, N128);
or OR4 (N1869, N1836, N874, N227, N703);
nor NOR2 (N1870, N1852, N852);
not NOT1 (N1871, N1868);
nand NAND3 (N1872, N1864, N158, N1074);
nor NOR2 (N1873, N1866, N1834);
nor NOR2 (N1874, N1858, N1037);
or OR4 (N1875, N1869, N196, N1666, N736);
not NOT1 (N1876, N1862);
xor XOR2 (N1877, N1874, N710);
not NOT1 (N1878, N1871);
nor NOR3 (N1879, N1875, N392, N596);
nand NAND4 (N1880, N1879, N506, N947, N743);
xor XOR2 (N1881, N1876, N881);
and AND3 (N1882, N1870, N1462, N1367);
nor NOR2 (N1883, N1882, N1112);
not NOT1 (N1884, N1878);
or OR3 (N1885, N1883, N675, N1527);
nand NAND2 (N1886, N1865, N307);
not NOT1 (N1887, N1872);
nor NOR2 (N1888, N1886, N1885);
nand NAND3 (N1889, N69, N784, N496);
buf BUF1 (N1890, N1877);
not NOT1 (N1891, N1884);
nand NAND3 (N1892, N1891, N1742, N1610);
xor XOR2 (N1893, N1881, N1473);
nand NAND4 (N1894, N1890, N1193, N616, N423);
nand NAND4 (N1895, N1887, N1291, N301, N684);
nor NOR4 (N1896, N1880, N1388, N1736, N1071);
nand NAND4 (N1897, N1893, N683, N1533, N789);
or OR4 (N1898, N1895, N1023, N371, N395);
and AND2 (N1899, N1898, N771);
or OR4 (N1900, N1897, N1604, N380, N884);
or OR4 (N1901, N1859, N727, N1686, N1495);
and AND2 (N1902, N1894, N1847);
buf BUF1 (N1903, N1829);
nor NOR2 (N1904, N1888, N1770);
and AND4 (N1905, N1901, N1285, N1333, N1751);
and AND2 (N1906, N1889, N1353);
nand NAND4 (N1907, N1902, N1278, N750, N1029);
or OR2 (N1908, N1896, N1149);
or OR2 (N1909, N1907, N810);
nor NOR3 (N1910, N1903, N1261, N1425);
buf BUF1 (N1911, N1909);
xor XOR2 (N1912, N1910, N1116);
buf BUF1 (N1913, N1904);
not NOT1 (N1914, N1892);
and AND3 (N1915, N1899, N1453, N1486);
buf BUF1 (N1916, N1908);
or OR3 (N1917, N1916, N615, N433);
xor XOR2 (N1918, N1906, N750);
and AND2 (N1919, N1913, N425);
and AND2 (N1920, N1915, N969);
nand NAND3 (N1921, N1911, N812, N1057);
or OR4 (N1922, N1900, N1341, N1210, N1573);
and AND4 (N1923, N1873, N1661, N220, N726);
buf BUF1 (N1924, N1918);
not NOT1 (N1925, N1919);
and AND4 (N1926, N1912, N68, N120, N1197);
nand NAND3 (N1927, N1905, N769, N320);
or OR2 (N1928, N1921, N616);
nand NAND4 (N1929, N1923, N720, N137, N685);
not NOT1 (N1930, N1924);
not NOT1 (N1931, N1925);
nor NOR2 (N1932, N1920, N1876);
xor XOR2 (N1933, N1932, N34);
nor NOR3 (N1934, N1927, N1724, N1196);
or OR4 (N1935, N1929, N696, N1044, N1055);
not NOT1 (N1936, N1934);
nor NOR3 (N1937, N1914, N772, N1319);
nand NAND4 (N1938, N1935, N1283, N1668, N1011);
and AND4 (N1939, N1938, N64, N1897, N1398);
or OR3 (N1940, N1936, N317, N162);
and AND3 (N1941, N1917, N1364, N159);
xor XOR2 (N1942, N1931, N431);
and AND4 (N1943, N1922, N143, N1733, N95);
nand NAND4 (N1944, N1942, N1941, N688, N1603);
and AND4 (N1945, N1037, N305, N416, N1869);
and AND3 (N1946, N1945, N396, N1403);
nand NAND4 (N1947, N1944, N1464, N1465, N1896);
buf BUF1 (N1948, N1939);
nand NAND4 (N1949, N1948, N1446, N1763, N224);
nand NAND3 (N1950, N1937, N817, N149);
nand NAND2 (N1951, N1950, N816);
buf BUF1 (N1952, N1951);
nor NOR2 (N1953, N1943, N1653);
nand NAND4 (N1954, N1940, N1467, N751, N1441);
xor XOR2 (N1955, N1933, N946);
xor XOR2 (N1956, N1952, N821);
and AND3 (N1957, N1947, N202, N1418);
not NOT1 (N1958, N1956);
xor XOR2 (N1959, N1957, N958);
nand NAND4 (N1960, N1953, N1379, N32, N1596);
nor NOR2 (N1961, N1955, N1657);
nor NOR2 (N1962, N1961, N35);
xor XOR2 (N1963, N1959, N897);
or OR4 (N1964, N1930, N63, N1167, N1334);
and AND3 (N1965, N1960, N249, N198);
xor XOR2 (N1966, N1964, N1165);
nor NOR3 (N1967, N1954, N947, N1306);
nand NAND4 (N1968, N1958, N1841, N928, N859);
nor NOR2 (N1969, N1967, N636);
nand NAND2 (N1970, N1965, N31);
xor XOR2 (N1971, N1949, N1122);
xor XOR2 (N1972, N1969, N1635);
buf BUF1 (N1973, N1971);
buf BUF1 (N1974, N1966);
not NOT1 (N1975, N1972);
or OR2 (N1976, N1973, N527);
xor XOR2 (N1977, N1974, N185);
or OR3 (N1978, N1975, N19, N758);
or OR3 (N1979, N1978, N1790, N1899);
nand NAND4 (N1980, N1979, N964, N1818, N105);
xor XOR2 (N1981, N1946, N671);
buf BUF1 (N1982, N1981);
and AND2 (N1983, N1982, N380);
xor XOR2 (N1984, N1968, N858);
and AND3 (N1985, N1980, N531, N657);
nor NOR3 (N1986, N1976, N197, N540);
xor XOR2 (N1987, N1928, N575);
not NOT1 (N1988, N1987);
not NOT1 (N1989, N1988);
nand NAND3 (N1990, N1983, N1450, N191);
buf BUF1 (N1991, N1984);
nor NOR4 (N1992, N1962, N618, N1218, N1267);
and AND4 (N1993, N1963, N1246, N284, N62);
and AND2 (N1994, N1989, N1022);
and AND3 (N1995, N1990, N957, N1555);
buf BUF1 (N1996, N1994);
or OR2 (N1997, N1993, N1069);
buf BUF1 (N1998, N1985);
nor NOR4 (N1999, N1970, N160, N294, N147);
and AND3 (N2000, N1995, N575, N1534);
and AND3 (N2001, N1997, N1403, N497);
nor NOR3 (N2002, N2000, N703, N1769);
xor XOR2 (N2003, N1991, N7);
nand NAND4 (N2004, N1992, N1243, N1433, N43);
buf BUF1 (N2005, N2002);
nor NOR2 (N2006, N1977, N1450);
and AND2 (N2007, N2003, N705);
xor XOR2 (N2008, N2005, N1364);
nand NAND3 (N2009, N1996, N1030, N1000);
nand NAND2 (N2010, N2008, N1777);
nor NOR4 (N2011, N1926, N508, N1820, N1953);
nor NOR3 (N2012, N1998, N1428, N823);
nand NAND3 (N2013, N2011, N1621, N1641);
buf BUF1 (N2014, N2006);
buf BUF1 (N2015, N2004);
not NOT1 (N2016, N2015);
nand NAND3 (N2017, N2012, N1123, N1955);
or OR2 (N2018, N1986, N412);
nand NAND4 (N2019, N2013, N1309, N563, N1123);
nor NOR2 (N2020, N2001, N1237);
buf BUF1 (N2021, N1999);
nor NOR3 (N2022, N2017, N200, N1822);
not NOT1 (N2023, N2009);
and AND2 (N2024, N2007, N712);
not NOT1 (N2025, N2014);
xor XOR2 (N2026, N2022, N2025);
nand NAND2 (N2027, N2015, N1560);
nor NOR3 (N2028, N2026, N102, N1296);
and AND2 (N2029, N2016, N1199);
nor NOR3 (N2030, N2019, N1776, N1300);
xor XOR2 (N2031, N2029, N46);
nand NAND2 (N2032, N2023, N1312);
or OR3 (N2033, N2018, N1788, N1245);
and AND4 (N2034, N2020, N1120, N1327, N333);
and AND2 (N2035, N2010, N1739);
nor NOR3 (N2036, N2021, N682, N190);
buf BUF1 (N2037, N2028);
nand NAND2 (N2038, N2034, N1647);
buf BUF1 (N2039, N2033);
and AND3 (N2040, N2039, N1273, N1847);
nand NAND2 (N2041, N2035, N200);
xor XOR2 (N2042, N2041, N698);
not NOT1 (N2043, N2040);
not NOT1 (N2044, N2038);
not NOT1 (N2045, N2042);
and AND2 (N2046, N2031, N257);
buf BUF1 (N2047, N2024);
xor XOR2 (N2048, N2027, N1460);
and AND2 (N2049, N2032, N1025);
and AND4 (N2050, N2036, N1087, N224, N1483);
or OR3 (N2051, N2048, N12, N795);
nand NAND3 (N2052, N2050, N579, N629);
xor XOR2 (N2053, N2045, N1344);
and AND2 (N2054, N2049, N270);
nor NOR2 (N2055, N2053, N724);
xor XOR2 (N2056, N2047, N1799);
nor NOR4 (N2057, N2055, N884, N1239, N1270);
and AND2 (N2058, N2037, N531);
nand NAND2 (N2059, N2058, N738);
nor NOR2 (N2060, N2052, N181);
nor NOR2 (N2061, N2044, N1451);
or OR3 (N2062, N2060, N1442, N1716);
not NOT1 (N2063, N2057);
xor XOR2 (N2064, N2030, N1948);
nor NOR4 (N2065, N2043, N1558, N709, N255);
buf BUF1 (N2066, N2054);
or OR4 (N2067, N2062, N18, N529, N873);
not NOT1 (N2068, N2063);
nor NOR2 (N2069, N2064, N1335);
nand NAND4 (N2070, N2051, N916, N1221, N772);
and AND2 (N2071, N2065, N1909);
nand NAND2 (N2072, N2068, N1931);
nand NAND2 (N2073, N2059, N1366);
not NOT1 (N2074, N2061);
or OR2 (N2075, N2072, N762);
and AND4 (N2076, N2073, N1451, N1744, N1940);
buf BUF1 (N2077, N2070);
nand NAND2 (N2078, N2071, N1347);
xor XOR2 (N2079, N2067, N1318);
or OR4 (N2080, N2078, N2056, N439, N820);
xor XOR2 (N2081, N585, N1386);
or OR2 (N2082, N2080, N1325);
xor XOR2 (N2083, N2075, N264);
nor NOR4 (N2084, N2046, N2000, N843, N1542);
or OR3 (N2085, N2076, N363, N503);
buf BUF1 (N2086, N2085);
nor NOR3 (N2087, N2066, N727, N1192);
nand NAND3 (N2088, N2086, N390, N1144);
xor XOR2 (N2089, N2069, N1890);
xor XOR2 (N2090, N2074, N1336);
nand NAND3 (N2091, N2088, N365, N883);
not NOT1 (N2092, N2084);
nand NAND3 (N2093, N2079, N1481, N1162);
buf BUF1 (N2094, N2092);
or OR4 (N2095, N2082, N1225, N1639, N64);
and AND3 (N2096, N2094, N1490, N139);
buf BUF1 (N2097, N2077);
and AND3 (N2098, N2083, N1462, N1219);
or OR2 (N2099, N2089, N1891);
buf BUF1 (N2100, N2095);
buf BUF1 (N2101, N2087);
nor NOR2 (N2102, N2097, N714);
not NOT1 (N2103, N2081);
not NOT1 (N2104, N2100);
nand NAND3 (N2105, N2091, N1501, N834);
nand NAND4 (N2106, N2093, N1261, N352, N511);
buf BUF1 (N2107, N2103);
nand NAND3 (N2108, N2104, N1624, N1151);
or OR3 (N2109, N2106, N1267, N359);
nand NAND3 (N2110, N2105, N658, N154);
nor NOR4 (N2111, N2101, N583, N636, N931);
and AND2 (N2112, N2108, N1974);
nor NOR3 (N2113, N2109, N448, N1331);
nand NAND3 (N2114, N2111, N67, N311);
buf BUF1 (N2115, N2102);
buf BUF1 (N2116, N2110);
not NOT1 (N2117, N2090);
and AND4 (N2118, N2107, N949, N553, N232);
buf BUF1 (N2119, N2112);
nand NAND4 (N2120, N2116, N1936, N167, N653);
and AND3 (N2121, N2098, N1221, N1938);
not NOT1 (N2122, N2119);
xor XOR2 (N2123, N2122, N908);
or OR4 (N2124, N2096, N500, N2050, N2074);
and AND4 (N2125, N2099, N720, N1588, N433);
not NOT1 (N2126, N2115);
xor XOR2 (N2127, N2126, N719);
not NOT1 (N2128, N2123);
buf BUF1 (N2129, N2121);
buf BUF1 (N2130, N2113);
or OR4 (N2131, N2129, N1553, N1095, N1015);
nor NOR2 (N2132, N2131, N1739);
xor XOR2 (N2133, N2127, N946);
nand NAND3 (N2134, N2120, N253, N2048);
and AND2 (N2135, N2128, N343);
xor XOR2 (N2136, N2133, N2021);
or OR4 (N2137, N2114, N1551, N1941, N1870);
buf BUF1 (N2138, N2130);
nor NOR3 (N2139, N2134, N1068, N1518);
nand NAND2 (N2140, N2136, N512);
nor NOR3 (N2141, N2117, N80, N1962);
buf BUF1 (N2142, N2138);
not NOT1 (N2143, N2141);
nand NAND2 (N2144, N2135, N1885);
nand NAND4 (N2145, N2124, N2141, N263, N1696);
nand NAND4 (N2146, N2125, N2134, N881, N1328);
nor NOR4 (N2147, N2142, N325, N900, N1061);
nand NAND3 (N2148, N2140, N586, N1060);
not NOT1 (N2149, N2146);
nor NOR2 (N2150, N2148, N141);
nand NAND2 (N2151, N2137, N23);
nand NAND4 (N2152, N2118, N1547, N1053, N560);
nor NOR2 (N2153, N2143, N691);
nand NAND4 (N2154, N2147, N1053, N1002, N1808);
buf BUF1 (N2155, N2150);
not NOT1 (N2156, N2153);
and AND4 (N2157, N2152, N1164, N46, N432);
not NOT1 (N2158, N2132);
xor XOR2 (N2159, N2154, N160);
xor XOR2 (N2160, N2156, N2065);
buf BUF1 (N2161, N2139);
or OR3 (N2162, N2161, N2151, N1048);
nand NAND2 (N2163, N486, N21);
buf BUF1 (N2164, N2160);
not NOT1 (N2165, N2149);
and AND3 (N2166, N2163, N583, N348);
and AND2 (N2167, N2164, N630);
xor XOR2 (N2168, N2162, N691);
nand NAND3 (N2169, N2157, N2006, N1637);
buf BUF1 (N2170, N2166);
not NOT1 (N2171, N2169);
xor XOR2 (N2172, N2170, N635);
or OR4 (N2173, N2165, N894, N1244, N25);
buf BUF1 (N2174, N2173);
buf BUF1 (N2175, N2168);
nand NAND2 (N2176, N2158, N1822);
or OR3 (N2177, N2145, N1286, N258);
nor NOR4 (N2178, N2177, N573, N1672, N2144);
not NOT1 (N2179, N330);
buf BUF1 (N2180, N2175);
or OR4 (N2181, N2159, N2067, N1177, N1945);
xor XOR2 (N2182, N2179, N644);
buf BUF1 (N2183, N2167);
or OR3 (N2184, N2182, N1038, N959);
nor NOR4 (N2185, N2183, N841, N529, N672);
buf BUF1 (N2186, N2185);
not NOT1 (N2187, N2172);
nor NOR4 (N2188, N2186, N459, N1487, N9);
nand NAND4 (N2189, N2176, N58, N1643, N1154);
or OR2 (N2190, N2155, N779);
nand NAND2 (N2191, N2171, N664);
buf BUF1 (N2192, N2178);
xor XOR2 (N2193, N2174, N598);
or OR2 (N2194, N2187, N1946);
and AND2 (N2195, N2190, N965);
or OR3 (N2196, N2188, N128, N138);
or OR3 (N2197, N2180, N582, N2077);
or OR4 (N2198, N2196, N535, N2113, N1475);
nand NAND3 (N2199, N2197, N14, N1690);
xor XOR2 (N2200, N2191, N170);
not NOT1 (N2201, N2189);
xor XOR2 (N2202, N2199, N1714);
nand NAND4 (N2203, N2193, N1511, N450, N1032);
xor XOR2 (N2204, N2181, N2077);
nor NOR4 (N2205, N2200, N730, N1088, N792);
buf BUF1 (N2206, N2195);
or OR3 (N2207, N2206, N629, N263);
nor NOR3 (N2208, N2198, N2144, N38);
not NOT1 (N2209, N2184);
nand NAND4 (N2210, N2207, N1513, N570, N1544);
buf BUF1 (N2211, N2203);
and AND3 (N2212, N2204, N1772, N839);
and AND3 (N2213, N2201, N2142, N690);
and AND4 (N2214, N2210, N1281, N1052, N924);
nor NOR2 (N2215, N2205, N1481);
or OR3 (N2216, N2209, N123, N2004);
buf BUF1 (N2217, N2215);
and AND3 (N2218, N2213, N407, N503);
xor XOR2 (N2219, N2217, N1080);
or OR3 (N2220, N2208, N432, N1555);
and AND4 (N2221, N2211, N424, N1856, N1610);
and AND2 (N2222, N2218, N1163);
xor XOR2 (N2223, N2219, N1949);
or OR4 (N2224, N2202, N945, N611, N689);
and AND2 (N2225, N2220, N436);
nor NOR2 (N2226, N2223, N400);
nor NOR4 (N2227, N2194, N1978, N1622, N420);
and AND4 (N2228, N2222, N748, N103, N1238);
buf BUF1 (N2229, N2192);
not NOT1 (N2230, N2216);
nor NOR2 (N2231, N2214, N2034);
xor XOR2 (N2232, N2228, N1758);
and AND2 (N2233, N2229, N2151);
xor XOR2 (N2234, N2212, N1473);
nor NOR2 (N2235, N2226, N412);
buf BUF1 (N2236, N2235);
nand NAND2 (N2237, N2234, N799);
not NOT1 (N2238, N2236);
xor XOR2 (N2239, N2238, N609);
nor NOR3 (N2240, N2224, N743, N586);
nand NAND3 (N2241, N2225, N1120, N271);
or OR4 (N2242, N2232, N1820, N1380, N1198);
not NOT1 (N2243, N2241);
nand NAND2 (N2244, N2221, N1406);
and AND4 (N2245, N2233, N352, N234, N2073);
nor NOR2 (N2246, N2239, N1112);
nor NOR2 (N2247, N2230, N2103);
buf BUF1 (N2248, N2242);
nand NAND4 (N2249, N2245, N242, N167, N276);
and AND2 (N2250, N2237, N508);
nand NAND2 (N2251, N2240, N1287);
or OR2 (N2252, N2251, N773);
nor NOR3 (N2253, N2243, N393, N737);
buf BUF1 (N2254, N2227);
not NOT1 (N2255, N2248);
xor XOR2 (N2256, N2247, N812);
nor NOR2 (N2257, N2254, N902);
not NOT1 (N2258, N2255);
nor NOR2 (N2259, N2231, N169);
or OR3 (N2260, N2258, N2052, N2026);
not NOT1 (N2261, N2253);
or OR4 (N2262, N2252, N1637, N591, N145);
not NOT1 (N2263, N2256);
xor XOR2 (N2264, N2257, N303);
buf BUF1 (N2265, N2262);
xor XOR2 (N2266, N2244, N1322);
not NOT1 (N2267, N2259);
xor XOR2 (N2268, N2266, N688);
nor NOR2 (N2269, N2268, N443);
not NOT1 (N2270, N2250);
nor NOR4 (N2271, N2270, N556, N481, N1718);
buf BUF1 (N2272, N2260);
nand NAND3 (N2273, N2263, N1993, N974);
xor XOR2 (N2274, N2265, N1260);
nor NOR3 (N2275, N2249, N555, N1033);
buf BUF1 (N2276, N2273);
nor NOR4 (N2277, N2246, N646, N800, N2085);
xor XOR2 (N2278, N2269, N531);
and AND3 (N2279, N2276, N196, N1962);
nand NAND4 (N2280, N2278, N1990, N2124, N1989);
not NOT1 (N2281, N2275);
nand NAND2 (N2282, N2280, N769);
or OR3 (N2283, N2279, N1188, N1542);
buf BUF1 (N2284, N2264);
nor NOR2 (N2285, N2271, N308);
or OR2 (N2286, N2283, N738);
nand NAND3 (N2287, N2286, N85, N2102);
xor XOR2 (N2288, N2284, N1489);
nor NOR3 (N2289, N2287, N384, N1377);
buf BUF1 (N2290, N2288);
buf BUF1 (N2291, N2281);
or OR2 (N2292, N2289, N1238);
not NOT1 (N2293, N2282);
and AND4 (N2294, N2267, N1106, N1009, N17);
or OR2 (N2295, N2291, N1169);
or OR3 (N2296, N2294, N1947, N1968);
not NOT1 (N2297, N2285);
buf BUF1 (N2298, N2296);
and AND2 (N2299, N2295, N1754);
nor NOR2 (N2300, N2292, N694);
not NOT1 (N2301, N2300);
and AND2 (N2302, N2299, N151);
buf BUF1 (N2303, N2302);
nand NAND4 (N2304, N2290, N2214, N1868, N1181);
nand NAND2 (N2305, N2277, N431);
xor XOR2 (N2306, N2297, N1524);
buf BUF1 (N2307, N2293);
nand NAND3 (N2308, N2305, N212, N88);
and AND2 (N2309, N2261, N186);
xor XOR2 (N2310, N2309, N1840);
xor XOR2 (N2311, N2303, N278);
buf BUF1 (N2312, N2274);
nor NOR4 (N2313, N2308, N341, N1086, N192);
buf BUF1 (N2314, N2301);
buf BUF1 (N2315, N2311);
buf BUF1 (N2316, N2307);
buf BUF1 (N2317, N2315);
or OR3 (N2318, N2298, N433, N2260);
nand NAND4 (N2319, N2304, N1558, N1558, N9);
xor XOR2 (N2320, N2313, N894);
buf BUF1 (N2321, N2314);
and AND3 (N2322, N2320, N2206, N2214);
nand NAND2 (N2323, N2321, N789);
and AND4 (N2324, N2316, N1699, N2095, N1437);
nand NAND3 (N2325, N2322, N1571, N62);
or OR2 (N2326, N2318, N1606);
buf BUF1 (N2327, N2317);
not NOT1 (N2328, N2319);
buf BUF1 (N2329, N2325);
nor NOR4 (N2330, N2326, N1954, N671, N79);
nand NAND3 (N2331, N2330, N932, N451);
xor XOR2 (N2332, N2324, N259);
or OR3 (N2333, N2331, N1853, N48);
buf BUF1 (N2334, N2328);
not NOT1 (N2335, N2333);
buf BUF1 (N2336, N2306);
nand NAND4 (N2337, N2310, N20, N2098, N925);
xor XOR2 (N2338, N2329, N220);
and AND4 (N2339, N2338, N1676, N1692, N2114);
and AND2 (N2340, N2312, N450);
nand NAND4 (N2341, N2340, N2080, N2124, N2272);
nand NAND4 (N2342, N1148, N437, N1442, N395);
buf BUF1 (N2343, N2341);
xor XOR2 (N2344, N2343, N212);
and AND4 (N2345, N2332, N834, N1002, N1566);
buf BUF1 (N2346, N2344);
or OR4 (N2347, N2335, N919, N2268, N338);
xor XOR2 (N2348, N2327, N2130);
and AND3 (N2349, N2346, N121, N883);
nor NOR3 (N2350, N2345, N833, N1552);
buf BUF1 (N2351, N2347);
xor XOR2 (N2352, N2350, N1652);
xor XOR2 (N2353, N2323, N441);
buf BUF1 (N2354, N2351);
or OR3 (N2355, N2353, N814, N2035);
xor XOR2 (N2356, N2336, N808);
not NOT1 (N2357, N2334);
nor NOR2 (N2358, N2337, N316);
not NOT1 (N2359, N2349);
not NOT1 (N2360, N2356);
and AND4 (N2361, N2352, N1720, N2090, N1036);
not NOT1 (N2362, N2342);
or OR3 (N2363, N2354, N259, N525);
not NOT1 (N2364, N2361);
nand NAND3 (N2365, N2363, N1041, N2148);
nand NAND2 (N2366, N2364, N2056);
or OR2 (N2367, N2339, N369);
xor XOR2 (N2368, N2348, N346);
buf BUF1 (N2369, N2366);
not NOT1 (N2370, N2357);
nor NOR3 (N2371, N2365, N1716, N1429);
xor XOR2 (N2372, N2368, N742);
nor NOR4 (N2373, N2358, N35, N1045, N2251);
xor XOR2 (N2374, N2355, N75);
buf BUF1 (N2375, N2367);
buf BUF1 (N2376, N2373);
not NOT1 (N2377, N2375);
nor NOR2 (N2378, N2372, N2299);
xor XOR2 (N2379, N2362, N1227);
xor XOR2 (N2380, N2370, N483);
nor NOR3 (N2381, N2376, N55, N1846);
not NOT1 (N2382, N2360);
xor XOR2 (N2383, N2382, N540);
and AND2 (N2384, N2374, N1863);
xor XOR2 (N2385, N2377, N797);
nor NOR2 (N2386, N2380, N1263);
not NOT1 (N2387, N2371);
nor NOR4 (N2388, N2359, N944, N202, N43);
nand NAND4 (N2389, N2385, N2285, N1337, N2083);
and AND2 (N2390, N2386, N1104);
not NOT1 (N2391, N2384);
nor NOR2 (N2392, N2383, N570);
buf BUF1 (N2393, N2379);
nand NAND4 (N2394, N2393, N1542, N1522, N1946);
not NOT1 (N2395, N2387);
xor XOR2 (N2396, N2378, N1191);
buf BUF1 (N2397, N2394);
buf BUF1 (N2398, N2388);
and AND4 (N2399, N2398, N1014, N1329, N190);
buf BUF1 (N2400, N2369);
not NOT1 (N2401, N2399);
nand NAND2 (N2402, N2389, N68);
or OR3 (N2403, N2391, N116, N1664);
and AND4 (N2404, N2390, N1898, N1978, N2246);
xor XOR2 (N2405, N2395, N1107);
nand NAND4 (N2406, N2396, N728, N958, N1260);
not NOT1 (N2407, N2400);
and AND4 (N2408, N2392, N1464, N1173, N2330);
xor XOR2 (N2409, N2402, N1040);
and AND3 (N2410, N2408, N849, N2132);
or OR3 (N2411, N2406, N2101, N117);
nor NOR4 (N2412, N2403, N889, N512, N1160);
nand NAND2 (N2413, N2397, N2372);
xor XOR2 (N2414, N2412, N465);
and AND4 (N2415, N2413, N730, N1495, N100);
not NOT1 (N2416, N2414);
not NOT1 (N2417, N2401);
xor XOR2 (N2418, N2409, N324);
or OR2 (N2419, N2418, N1529);
and AND2 (N2420, N2415, N143);
nor NOR3 (N2421, N2416, N464, N1761);
and AND4 (N2422, N2417, N1397, N964, N1898);
and AND2 (N2423, N2421, N1414);
buf BUF1 (N2424, N2405);
or OR2 (N2425, N2423, N1524);
nand NAND3 (N2426, N2381, N1141, N2072);
or OR4 (N2427, N2407, N1038, N1401, N549);
not NOT1 (N2428, N2422);
nor NOR4 (N2429, N2404, N1194, N1415, N1169);
or OR2 (N2430, N2420, N1580);
nand NAND4 (N2431, N2411, N143, N1278, N2062);
buf BUF1 (N2432, N2419);
xor XOR2 (N2433, N2425, N896);
not NOT1 (N2434, N2429);
nor NOR4 (N2435, N2434, N1668, N2263, N2363);
or OR4 (N2436, N2432, N1148, N806, N644);
buf BUF1 (N2437, N2431);
xor XOR2 (N2438, N2424, N340);
buf BUF1 (N2439, N2427);
not NOT1 (N2440, N2430);
nor NOR4 (N2441, N2426, N1275, N692, N308);
nand NAND4 (N2442, N2437, N895, N1486, N1753);
nand NAND4 (N2443, N2441, N994, N2066, N67);
nand NAND2 (N2444, N2435, N11);
xor XOR2 (N2445, N2444, N593);
nand NAND2 (N2446, N2428, N2046);
buf BUF1 (N2447, N2439);
xor XOR2 (N2448, N2433, N2419);
or OR4 (N2449, N2436, N1831, N455, N2375);
buf BUF1 (N2450, N2438);
nor NOR4 (N2451, N2442, N498, N832, N846);
buf BUF1 (N2452, N2410);
xor XOR2 (N2453, N2445, N372);
nor NOR3 (N2454, N2451, N220, N949);
nand NAND4 (N2455, N2446, N1832, N401, N1366);
not NOT1 (N2456, N2452);
nor NOR2 (N2457, N2448, N248);
nor NOR4 (N2458, N2457, N1078, N1882, N783);
and AND2 (N2459, N2455, N1947);
nor NOR2 (N2460, N2456, N1943);
nor NOR4 (N2461, N2453, N1777, N1260, N1330);
or OR3 (N2462, N2447, N733, N919);
nand NAND3 (N2463, N2462, N1386, N2098);
xor XOR2 (N2464, N2463, N1679);
nor NOR2 (N2465, N2443, N1931);
or OR4 (N2466, N2449, N1628, N827, N262);
and AND2 (N2467, N2465, N1400);
nor NOR2 (N2468, N2459, N1089);
nand NAND3 (N2469, N2458, N7, N14);
xor XOR2 (N2470, N2464, N1698);
nor NOR2 (N2471, N2466, N701);
nor NOR2 (N2472, N2450, N37);
and AND4 (N2473, N2440, N344, N429, N878);
buf BUF1 (N2474, N2467);
nor NOR3 (N2475, N2471, N2165, N1916);
nor NOR3 (N2476, N2468, N1893, N659);
buf BUF1 (N2477, N2475);
not NOT1 (N2478, N2454);
not NOT1 (N2479, N2460);
nor NOR3 (N2480, N2478, N845, N555);
buf BUF1 (N2481, N2474);
xor XOR2 (N2482, N2469, N241);
and AND2 (N2483, N2479, N131);
and AND2 (N2484, N2476, N842);
xor XOR2 (N2485, N2473, N2402);
buf BUF1 (N2486, N2483);
not NOT1 (N2487, N2484);
buf BUF1 (N2488, N2477);
nor NOR3 (N2489, N2486, N260, N676);
xor XOR2 (N2490, N2461, N593);
and AND4 (N2491, N2472, N1135, N188, N891);
nor NOR4 (N2492, N2470, N1079, N207, N343);
buf BUF1 (N2493, N2490);
xor XOR2 (N2494, N2492, N879);
buf BUF1 (N2495, N2485);
or OR3 (N2496, N2489, N1134, N867);
or OR2 (N2497, N2494, N600);
xor XOR2 (N2498, N2491, N603);
nor NOR3 (N2499, N2493, N178, N1772);
not NOT1 (N2500, N2495);
xor XOR2 (N2501, N2498, N2330);
nand NAND4 (N2502, N2487, N1827, N1672, N127);
buf BUF1 (N2503, N2501);
not NOT1 (N2504, N2502);
xor XOR2 (N2505, N2488, N724);
or OR4 (N2506, N2503, N1501, N903, N138);
or OR2 (N2507, N2506, N426);
not NOT1 (N2508, N2507);
buf BUF1 (N2509, N2481);
not NOT1 (N2510, N2499);
and AND3 (N2511, N2482, N1477, N666);
nor NOR2 (N2512, N2509, N646);
or OR3 (N2513, N2511, N814, N2459);
or OR2 (N2514, N2512, N338);
or OR3 (N2515, N2504, N2410, N2021);
or OR4 (N2516, N2505, N2098, N1757, N2106);
buf BUF1 (N2517, N2514);
not NOT1 (N2518, N2497);
buf BUF1 (N2519, N2518);
not NOT1 (N2520, N2496);
or OR3 (N2521, N2513, N394, N26);
xor XOR2 (N2522, N2521, N2100);
nor NOR3 (N2523, N2522, N229, N1623);
nor NOR3 (N2524, N2516, N1026, N1774);
nor NOR3 (N2525, N2524, N1667, N2090);
xor XOR2 (N2526, N2517, N712);
xor XOR2 (N2527, N2515, N683);
nor NOR2 (N2528, N2526, N391);
nor NOR4 (N2529, N2527, N2099, N2136, N1731);
nand NAND4 (N2530, N2519, N280, N1161, N2311);
or OR4 (N2531, N2523, N2009, N975, N2026);
not NOT1 (N2532, N2528);
and AND4 (N2533, N2532, N1531, N520, N2128);
buf BUF1 (N2534, N2508);
buf BUF1 (N2535, N2510);
nand NAND4 (N2536, N2534, N1189, N2247, N348);
buf BUF1 (N2537, N2533);
and AND3 (N2538, N2525, N976, N2063);
or OR3 (N2539, N2520, N1275, N1620);
nand NAND3 (N2540, N2500, N1196, N1135);
or OR4 (N2541, N2531, N1693, N463, N1492);
not NOT1 (N2542, N2540);
nor NOR4 (N2543, N2530, N787, N1291, N2489);
not NOT1 (N2544, N2536);
nand NAND2 (N2545, N2542, N542);
or OR3 (N2546, N2537, N1087, N2242);
not NOT1 (N2547, N2480);
nor NOR2 (N2548, N2529, N1020);
nor NOR3 (N2549, N2538, N1989, N292);
nor NOR2 (N2550, N2544, N473);
or OR4 (N2551, N2547, N582, N1182, N1567);
and AND2 (N2552, N2543, N1721);
not NOT1 (N2553, N2541);
or OR2 (N2554, N2551, N596);
xor XOR2 (N2555, N2546, N349);
nand NAND2 (N2556, N2548, N1569);
xor XOR2 (N2557, N2549, N1409);
and AND3 (N2558, N2545, N1722, N1873);
nor NOR2 (N2559, N2557, N1941);
xor XOR2 (N2560, N2555, N1746);
not NOT1 (N2561, N2553);
nor NOR3 (N2562, N2561, N1286, N1546);
nand NAND3 (N2563, N2562, N1232, N2002);
nand NAND3 (N2564, N2539, N2093, N1836);
nand NAND2 (N2565, N2563, N533);
nand NAND4 (N2566, N2554, N111, N680, N2295);
not NOT1 (N2567, N2550);
or OR2 (N2568, N2558, N2396);
nor NOR4 (N2569, N2567, N1105, N949, N756);
nand NAND4 (N2570, N2566, N1046, N2297, N1201);
nor NOR2 (N2571, N2559, N1369);
nor NOR4 (N2572, N2569, N858, N1366, N2389);
not NOT1 (N2573, N2570);
xor XOR2 (N2574, N2565, N329);
buf BUF1 (N2575, N2573);
nor NOR4 (N2576, N2568, N832, N752, N2240);
buf BUF1 (N2577, N2575);
or OR4 (N2578, N2571, N1495, N454, N2256);
and AND3 (N2579, N2556, N2260, N1160);
xor XOR2 (N2580, N2578, N1070);
xor XOR2 (N2581, N2572, N447);
or OR3 (N2582, N2574, N316, N1917);
buf BUF1 (N2583, N2564);
xor XOR2 (N2584, N2552, N763);
nor NOR2 (N2585, N2580, N273);
nor NOR3 (N2586, N2584, N67, N2288);
nand NAND4 (N2587, N2582, N2504, N1146, N979);
nand NAND3 (N2588, N2577, N129, N1002);
buf BUF1 (N2589, N2588);
buf BUF1 (N2590, N2587);
xor XOR2 (N2591, N2581, N690);
nor NOR4 (N2592, N2591, N901, N2126, N2468);
nor NOR2 (N2593, N2585, N1404);
or OR2 (N2594, N2586, N1587);
or OR4 (N2595, N2579, N2583, N2256, N2035);
buf BUF1 (N2596, N1460);
nor NOR3 (N2597, N2560, N796, N317);
nor NOR4 (N2598, N2535, N298, N923, N2285);
xor XOR2 (N2599, N2590, N2522);
not NOT1 (N2600, N2576);
nor NOR2 (N2601, N2597, N2296);
nand NAND3 (N2602, N2592, N1844, N1582);
buf BUF1 (N2603, N2596);
and AND4 (N2604, N2600, N816, N428, N2480);
xor XOR2 (N2605, N2602, N1488);
xor XOR2 (N2606, N2589, N1307);
not NOT1 (N2607, N2601);
or OR3 (N2608, N2606, N750, N239);
xor XOR2 (N2609, N2608, N649);
xor XOR2 (N2610, N2603, N2589);
and AND2 (N2611, N2604, N284);
or OR2 (N2612, N2593, N2275);
or OR3 (N2613, N2611, N156, N2107);
nand NAND3 (N2614, N2598, N2249, N2072);
nor NOR2 (N2615, N2610, N1719);
and AND2 (N2616, N2607, N271);
or OR2 (N2617, N2612, N12);
nor NOR2 (N2618, N2614, N1109);
nand NAND4 (N2619, N2594, N1562, N635, N1252);
and AND4 (N2620, N2615, N312, N821, N255);
and AND4 (N2621, N2609, N189, N509, N2097);
xor XOR2 (N2622, N2616, N872);
not NOT1 (N2623, N2617);
or OR2 (N2624, N2623, N904);
nor NOR3 (N2625, N2622, N168, N1965);
nor NOR3 (N2626, N2621, N1782, N335);
buf BUF1 (N2627, N2618);
not NOT1 (N2628, N2605);
nor NOR2 (N2629, N2624, N2049);
nor NOR3 (N2630, N2595, N1501, N1879);
buf BUF1 (N2631, N2619);
not NOT1 (N2632, N2629);
not NOT1 (N2633, N2628);
not NOT1 (N2634, N2620);
and AND4 (N2635, N2634, N90, N2436, N253);
not NOT1 (N2636, N2633);
not NOT1 (N2637, N2625);
nor NOR3 (N2638, N2632, N93, N367);
nor NOR2 (N2639, N2638, N2295);
or OR4 (N2640, N2599, N2577, N2161, N2472);
and AND3 (N2641, N2639, N845, N1146);
and AND4 (N2642, N2631, N898, N546, N2072);
not NOT1 (N2643, N2641);
and AND2 (N2644, N2635, N400);
buf BUF1 (N2645, N2637);
nor NOR2 (N2646, N2627, N2573);
nand NAND4 (N2647, N2613, N132, N686, N2117);
nand NAND2 (N2648, N2644, N768);
and AND2 (N2649, N2647, N1366);
nor NOR2 (N2650, N2649, N2335);
and AND4 (N2651, N2630, N591, N2370, N327);
nand NAND4 (N2652, N2651, N2434, N1000, N1481);
nor NOR2 (N2653, N2643, N2321);
not NOT1 (N2654, N2653);
and AND3 (N2655, N2646, N2191, N2460);
buf BUF1 (N2656, N2636);
xor XOR2 (N2657, N2655, N354);
nor NOR4 (N2658, N2654, N1230, N1210, N1388);
not NOT1 (N2659, N2626);
nand NAND4 (N2660, N2656, N237, N719, N2342);
nand NAND4 (N2661, N2657, N1313, N1827, N2403);
nor NOR4 (N2662, N2660, N1247, N607, N2128);
xor XOR2 (N2663, N2658, N1608);
and AND4 (N2664, N2661, N2427, N94, N327);
nor NOR2 (N2665, N2652, N1744);
nand NAND2 (N2666, N2650, N664);
or OR4 (N2667, N2640, N766, N1338, N333);
buf BUF1 (N2668, N2659);
and AND2 (N2669, N2668, N864);
xor XOR2 (N2670, N2669, N2156);
and AND2 (N2671, N2666, N2277);
xor XOR2 (N2672, N2664, N274);
or OR2 (N2673, N2665, N1871);
and AND4 (N2674, N2667, N686, N839, N498);
nand NAND2 (N2675, N2645, N952);
nand NAND4 (N2676, N2671, N1220, N2292, N1065);
not NOT1 (N2677, N2673);
or OR4 (N2678, N2663, N515, N1329, N1043);
xor XOR2 (N2679, N2678, N2237);
xor XOR2 (N2680, N2662, N977);
xor XOR2 (N2681, N2674, N877);
xor XOR2 (N2682, N2675, N2311);
nor NOR4 (N2683, N2672, N2207, N2637, N2498);
nor NOR2 (N2684, N2642, N1638);
and AND2 (N2685, N2684, N2346);
or OR3 (N2686, N2681, N1744, N81);
nand NAND3 (N2687, N2670, N1030, N1628);
or OR2 (N2688, N2683, N375);
not NOT1 (N2689, N2680);
and AND4 (N2690, N2648, N589, N1843, N2030);
not NOT1 (N2691, N2690);
not NOT1 (N2692, N2691);
or OR4 (N2693, N2689, N710, N1330, N1673);
xor XOR2 (N2694, N2676, N482);
buf BUF1 (N2695, N2685);
not NOT1 (N2696, N2687);
not NOT1 (N2697, N2696);
nand NAND3 (N2698, N2679, N2680, N2434);
nor NOR4 (N2699, N2693, N1515, N1858, N2196);
or OR3 (N2700, N2694, N1124, N1749);
nand NAND4 (N2701, N2682, N1565, N775, N947);
nor NOR3 (N2702, N2695, N776, N1878);
and AND3 (N2703, N2677, N871, N1507);
not NOT1 (N2704, N2697);
nand NAND3 (N2705, N2686, N750, N708);
not NOT1 (N2706, N2702);
nand NAND2 (N2707, N2701, N2074);
nor NOR2 (N2708, N2704, N2199);
nor NOR2 (N2709, N2698, N30);
nor NOR3 (N2710, N2700, N361, N1715);
or OR4 (N2711, N2708, N958, N1460, N1733);
buf BUF1 (N2712, N2703);
buf BUF1 (N2713, N2712);
or OR2 (N2714, N2706, N2473);
nand NAND4 (N2715, N2713, N1102, N2210, N2664);
or OR2 (N2716, N2699, N2565);
and AND4 (N2717, N2711, N1061, N224, N2386);
or OR2 (N2718, N2692, N2226);
xor XOR2 (N2719, N2709, N861);
or OR2 (N2720, N2717, N1927);
nor NOR3 (N2721, N2707, N1060, N1493);
xor XOR2 (N2722, N2718, N2289);
or OR3 (N2723, N2721, N2409, N1955);
nand NAND4 (N2724, N2716, N925, N662, N353);
nand NAND2 (N2725, N2719, N2641);
and AND3 (N2726, N2725, N472, N2069);
buf BUF1 (N2727, N2722);
buf BUF1 (N2728, N2688);
not NOT1 (N2729, N2714);
or OR3 (N2730, N2720, N1153, N2434);
not NOT1 (N2731, N2724);
buf BUF1 (N2732, N2715);
not NOT1 (N2733, N2730);
or OR3 (N2734, N2726, N177, N1735);
nand NAND2 (N2735, N2732, N300);
and AND3 (N2736, N2727, N219, N2046);
and AND3 (N2737, N2731, N12, N2447);
buf BUF1 (N2738, N2737);
nand NAND2 (N2739, N2728, N108);
xor XOR2 (N2740, N2736, N1319);
nor NOR3 (N2741, N2729, N1104, N610);
and AND4 (N2742, N2733, N1776, N2369, N2177);
and AND2 (N2743, N2705, N444);
buf BUF1 (N2744, N2723);
nand NAND2 (N2745, N2740, N2109);
or OR3 (N2746, N2741, N1133, N853);
or OR2 (N2747, N2735, N1976);
and AND4 (N2748, N2743, N2639, N543, N1660);
and AND4 (N2749, N2739, N1267, N2333, N649);
nand NAND2 (N2750, N2745, N428);
nand NAND2 (N2751, N2734, N973);
or OR3 (N2752, N2742, N2213, N596);
or OR2 (N2753, N2747, N452);
xor XOR2 (N2754, N2750, N2545);
or OR4 (N2755, N2748, N2563, N1691, N845);
nand NAND3 (N2756, N2710, N403, N2272);
nand NAND2 (N2757, N2755, N603);
xor XOR2 (N2758, N2749, N1161);
nand NAND3 (N2759, N2754, N1243, N727);
nand NAND4 (N2760, N2758, N1980, N2540, N1781);
and AND4 (N2761, N2756, N1437, N668, N2067);
buf BUF1 (N2762, N2761);
and AND2 (N2763, N2759, N2442);
or OR2 (N2764, N2751, N858);
nand NAND2 (N2765, N2757, N431);
and AND2 (N2766, N2746, N1384);
nor NOR2 (N2767, N2766, N2278);
buf BUF1 (N2768, N2764);
xor XOR2 (N2769, N2760, N693);
xor XOR2 (N2770, N2768, N1056);
and AND3 (N2771, N2752, N577, N397);
nand NAND2 (N2772, N2767, N2404);
not NOT1 (N2773, N2753);
nor NOR2 (N2774, N2769, N1598);
not NOT1 (N2775, N2774);
not NOT1 (N2776, N2744);
nor NOR4 (N2777, N2776, N626, N2295, N2235);
xor XOR2 (N2778, N2771, N2057);
buf BUF1 (N2779, N2738);
nand NAND4 (N2780, N2763, N2640, N2510, N1900);
not NOT1 (N2781, N2779);
xor XOR2 (N2782, N2781, N2104);
buf BUF1 (N2783, N2765);
nor NOR3 (N2784, N2773, N636, N2165);
buf BUF1 (N2785, N2775);
or OR2 (N2786, N2770, N135);
and AND3 (N2787, N2785, N2756, N1070);
nand NAND4 (N2788, N2783, N1392, N437, N2273);
and AND3 (N2789, N2788, N1411, N1968);
xor XOR2 (N2790, N2789, N425);
and AND4 (N2791, N2787, N299, N1879, N1245);
nand NAND4 (N2792, N2762, N1946, N1995, N2200);
or OR4 (N2793, N2792, N309, N327, N842);
or OR3 (N2794, N2786, N1935, N1056);
and AND3 (N2795, N2777, N2460, N993);
nor NOR4 (N2796, N2778, N1432, N2329, N818);
buf BUF1 (N2797, N2784);
or OR3 (N2798, N2796, N157, N291);
xor XOR2 (N2799, N2780, N960);
nand NAND3 (N2800, N2798, N732, N1563);
nand NAND2 (N2801, N2797, N1541);
or OR4 (N2802, N2793, N714, N1370, N1151);
or OR4 (N2803, N2799, N428, N2482, N620);
xor XOR2 (N2804, N2794, N55);
buf BUF1 (N2805, N2795);
not NOT1 (N2806, N2772);
nand NAND3 (N2807, N2800, N1393, N1553);
buf BUF1 (N2808, N2807);
buf BUF1 (N2809, N2782);
and AND3 (N2810, N2809, N1863, N1713);
nor NOR4 (N2811, N2810, N2286, N358, N1556);
buf BUF1 (N2812, N2801);
nor NOR3 (N2813, N2811, N709, N731);
not NOT1 (N2814, N2791);
buf BUF1 (N2815, N2802);
buf BUF1 (N2816, N2804);
or OR2 (N2817, N2806, N61);
nand NAND3 (N2818, N2805, N1815, N1319);
nand NAND2 (N2819, N2812, N1425);
not NOT1 (N2820, N2815);
xor XOR2 (N2821, N2817, N1614);
xor XOR2 (N2822, N2819, N1897);
nor NOR3 (N2823, N2813, N1618, N1878);
not NOT1 (N2824, N2822);
not NOT1 (N2825, N2814);
xor XOR2 (N2826, N2821, N2614);
nor NOR3 (N2827, N2808, N408, N867);
nor NOR3 (N2828, N2825, N63, N1626);
buf BUF1 (N2829, N2828);
nand NAND3 (N2830, N2827, N1836, N1484);
buf BUF1 (N2831, N2830);
nor NOR2 (N2832, N2823, N52);
or OR2 (N2833, N2803, N2022);
not NOT1 (N2834, N2818);
nor NOR3 (N2835, N2824, N948, N413);
buf BUF1 (N2836, N2832);
and AND2 (N2837, N2836, N2716);
and AND2 (N2838, N2829, N2180);
nand NAND2 (N2839, N2790, N1597);
xor XOR2 (N2840, N2833, N2093);
buf BUF1 (N2841, N2831);
or OR3 (N2842, N2837, N2226, N2665);
buf BUF1 (N2843, N2839);
and AND2 (N2844, N2826, N36);
nor NOR2 (N2845, N2816, N1463);
not NOT1 (N2846, N2838);
xor XOR2 (N2847, N2844, N136);
nor NOR3 (N2848, N2845, N2386, N2414);
buf BUF1 (N2849, N2835);
xor XOR2 (N2850, N2847, N1981);
and AND3 (N2851, N2846, N127, N2713);
and AND2 (N2852, N2834, N1286);
nor NOR3 (N2853, N2849, N2331, N2847);
nand NAND3 (N2854, N2820, N2259, N2105);
xor XOR2 (N2855, N2841, N2811);
nor NOR2 (N2856, N2843, N1636);
nand NAND2 (N2857, N2840, N1796);
or OR3 (N2858, N2851, N1411, N2020);
nor NOR4 (N2859, N2842, N2627, N817, N671);
xor XOR2 (N2860, N2857, N2674);
or OR3 (N2861, N2854, N2565, N1799);
and AND2 (N2862, N2859, N641);
and AND4 (N2863, N2862, N1135, N2184, N1969);
and AND3 (N2864, N2863, N1766, N2297);
xor XOR2 (N2865, N2856, N1044);
not NOT1 (N2866, N2850);
buf BUF1 (N2867, N2855);
xor XOR2 (N2868, N2865, N2040);
xor XOR2 (N2869, N2867, N2417);
xor XOR2 (N2870, N2848, N1643);
buf BUF1 (N2871, N2866);
buf BUF1 (N2872, N2852);
or OR4 (N2873, N2864, N1498, N2374, N958);
nor NOR4 (N2874, N2868, N790, N1237, N362);
nand NAND3 (N2875, N2869, N1154, N545);
not NOT1 (N2876, N2860);
not NOT1 (N2877, N2861);
and AND2 (N2878, N2853, N1233);
nand NAND2 (N2879, N2876, N158);
or OR2 (N2880, N2874, N1531);
nand NAND4 (N2881, N2871, N1069, N1981, N1202);
xor XOR2 (N2882, N2877, N977);
xor XOR2 (N2883, N2880, N763);
or OR2 (N2884, N2872, N66);
or OR2 (N2885, N2881, N239);
xor XOR2 (N2886, N2884, N2765);
nor NOR3 (N2887, N2858, N1539, N818);
buf BUF1 (N2888, N2878);
nand NAND2 (N2889, N2888, N2688);
nand NAND4 (N2890, N2879, N1175, N867, N1099);
or OR3 (N2891, N2890, N601, N508);
nand NAND2 (N2892, N2875, N2657);
and AND4 (N2893, N2883, N2412, N2095, N326);
buf BUF1 (N2894, N2882);
and AND4 (N2895, N2870, N1461, N406, N1791);
xor XOR2 (N2896, N2885, N349);
xor XOR2 (N2897, N2896, N2365);
nor NOR3 (N2898, N2873, N1410, N258);
xor XOR2 (N2899, N2891, N1708);
not NOT1 (N2900, N2899);
nor NOR3 (N2901, N2895, N1115, N2852);
nor NOR3 (N2902, N2901, N110, N2007);
and AND4 (N2903, N2894, N1472, N2577, N2054);
buf BUF1 (N2904, N2892);
buf BUF1 (N2905, N2893);
and AND3 (N2906, N2887, N620, N1197);
and AND2 (N2907, N2889, N2112);
not NOT1 (N2908, N2900);
not NOT1 (N2909, N2897);
buf BUF1 (N2910, N2908);
and AND4 (N2911, N2903, N764, N1747, N314);
or OR2 (N2912, N2906, N2097);
nor NOR3 (N2913, N2898, N2221, N1792);
nor NOR2 (N2914, N2902, N369);
xor XOR2 (N2915, N2909, N851);
buf BUF1 (N2916, N2904);
or OR3 (N2917, N2886, N571, N2741);
or OR2 (N2918, N2905, N2190);
buf BUF1 (N2919, N2907);
nand NAND3 (N2920, N2913, N1990, N1714);
or OR4 (N2921, N2915, N57, N2722, N2494);
buf BUF1 (N2922, N2911);
buf BUF1 (N2923, N2922);
or OR4 (N2924, N2921, N2795, N1156, N2275);
nand NAND4 (N2925, N2923, N374, N2413, N1651);
xor XOR2 (N2926, N2925, N2675);
not NOT1 (N2927, N2912);
nor NOR4 (N2928, N2910, N2604, N73, N326);
nor NOR3 (N2929, N2918, N2220, N1439);
and AND2 (N2930, N2920, N2322);
buf BUF1 (N2931, N2924);
and AND4 (N2932, N2916, N2520, N2, N1342);
buf BUF1 (N2933, N2927);
nand NAND3 (N2934, N2928, N1724, N1393);
nand NAND3 (N2935, N2917, N209, N780);
or OR2 (N2936, N2919, N2675);
not NOT1 (N2937, N2930);
nor NOR3 (N2938, N2936, N1204, N1237);
buf BUF1 (N2939, N2935);
nor NOR2 (N2940, N2926, N2808);
nor NOR2 (N2941, N2939, N2066);
nand NAND4 (N2942, N2933, N1902, N2923, N494);
xor XOR2 (N2943, N2934, N445);
xor XOR2 (N2944, N2937, N1624);
not NOT1 (N2945, N2940);
or OR4 (N2946, N2943, N1820, N2691, N213);
or OR4 (N2947, N2942, N1485, N719, N2353);
nor NOR3 (N2948, N2947, N1343, N1067);
not NOT1 (N2949, N2914);
nand NAND2 (N2950, N2932, N569);
nor NOR3 (N2951, N2944, N2189, N1231);
not NOT1 (N2952, N2951);
not NOT1 (N2953, N2941);
nand NAND3 (N2954, N2945, N1104, N1437);
or OR2 (N2955, N2952, N796);
or OR3 (N2956, N2946, N864, N1417);
buf BUF1 (N2957, N2948);
nand NAND4 (N2958, N2931, N879, N2078, N1145);
or OR3 (N2959, N2957, N2352, N517);
or OR2 (N2960, N2955, N2152);
nand NAND4 (N2961, N2938, N2441, N737, N2118);
buf BUF1 (N2962, N2950);
not NOT1 (N2963, N2949);
xor XOR2 (N2964, N2962, N640);
nand NAND3 (N2965, N2960, N1964, N1515);
not NOT1 (N2966, N2961);
xor XOR2 (N2967, N2964, N790);
not NOT1 (N2968, N2966);
or OR4 (N2969, N2963, N2867, N2019, N1572);
not NOT1 (N2970, N2953);
not NOT1 (N2971, N2969);
buf BUF1 (N2972, N2968);
nor NOR2 (N2973, N2970, N1364);
not NOT1 (N2974, N2959);
nor NOR4 (N2975, N2956, N524, N2920, N1195);
not NOT1 (N2976, N2958);
xor XOR2 (N2977, N2972, N467);
and AND4 (N2978, N2974, N100, N905, N1305);
or OR2 (N2979, N2977, N763);
nand NAND4 (N2980, N2978, N2946, N1673, N1940);
nand NAND4 (N2981, N2954, N2824, N1113, N769);
and AND4 (N2982, N2981, N79, N2308, N258);
not NOT1 (N2983, N2979);
not NOT1 (N2984, N2965);
and AND3 (N2985, N2973, N716, N1322);
nor NOR2 (N2986, N2929, N732);
xor XOR2 (N2987, N2984, N2466);
xor XOR2 (N2988, N2967, N2330);
nor NOR3 (N2989, N2986, N2433, N580);
nor NOR2 (N2990, N2985, N2614);
nor NOR2 (N2991, N2976, N650);
nor NOR4 (N2992, N2989, N2455, N1407, N2731);
nor NOR4 (N2993, N2987, N2562, N1988, N1506);
xor XOR2 (N2994, N2982, N756);
or OR3 (N2995, N2975, N165, N783);
xor XOR2 (N2996, N2994, N12);
nor NOR3 (N2997, N2980, N1681, N1779);
buf BUF1 (N2998, N2993);
buf BUF1 (N2999, N2971);
nand NAND3 (N3000, N2988, N1320, N1190);
and AND3 (N3001, N2998, N181, N1532);
nor NOR4 (N3002, N2992, N2951, N1189, N2424);
nor NOR2 (N3003, N2999, N559);
xor XOR2 (N3004, N2983, N2633);
or OR3 (N3005, N3004, N202, N1223);
or OR4 (N3006, N2991, N1414, N742, N121);
or OR4 (N3007, N3005, N556, N1290, N867);
and AND4 (N3008, N2996, N397, N620, N2622);
xor XOR2 (N3009, N3006, N1979);
not NOT1 (N3010, N3001);
or OR2 (N3011, N2995, N713);
or OR4 (N3012, N3011, N2702, N2619, N419);
and AND3 (N3013, N3010, N2909, N1480);
not NOT1 (N3014, N3009);
nand NAND3 (N3015, N3007, N107, N735);
nand NAND3 (N3016, N3012, N2891, N470);
nor NOR2 (N3017, N3002, N2386);
buf BUF1 (N3018, N3014);
nor NOR3 (N3019, N3018, N1050, N355);
buf BUF1 (N3020, N2997);
not NOT1 (N3021, N3008);
and AND2 (N3022, N3015, N2504);
nor NOR4 (N3023, N3003, N778, N1884, N2050);
or OR4 (N3024, N3021, N2421, N453, N851);
nor NOR2 (N3025, N3019, N1648);
or OR4 (N3026, N3017, N36, N2420, N2838);
not NOT1 (N3027, N2990);
nand NAND4 (N3028, N3020, N119, N2410, N671);
nor NOR2 (N3029, N3013, N2252);
xor XOR2 (N3030, N3027, N2238);
or OR2 (N3031, N3024, N2296);
nor NOR3 (N3032, N3028, N1592, N2276);
not NOT1 (N3033, N3023);
buf BUF1 (N3034, N3031);
xor XOR2 (N3035, N3000, N1501);
xor XOR2 (N3036, N3029, N2679);
xor XOR2 (N3037, N3030, N2292);
or OR2 (N3038, N3022, N295);
and AND3 (N3039, N3016, N1881, N2189);
xor XOR2 (N3040, N3036, N480);
nand NAND3 (N3041, N3032, N1663, N1397);
nor NOR3 (N3042, N3039, N637, N1427);
and AND2 (N3043, N3042, N2534);
nor NOR4 (N3044, N3025, N1862, N83, N500);
and AND4 (N3045, N3041, N2440, N1972, N1080);
nand NAND2 (N3046, N3035, N1509);
not NOT1 (N3047, N3026);
xor XOR2 (N3048, N3038, N2376);
buf BUF1 (N3049, N3047);
or OR4 (N3050, N3046, N1939, N385, N1106);
buf BUF1 (N3051, N3037);
xor XOR2 (N3052, N3044, N2148);
not NOT1 (N3053, N3050);
nand NAND4 (N3054, N3045, N2414, N435, N1010);
xor XOR2 (N3055, N3049, N240);
not NOT1 (N3056, N3053);
nand NAND2 (N3057, N3055, N1963);
buf BUF1 (N3058, N3052);
nand NAND3 (N3059, N3034, N631, N162);
not NOT1 (N3060, N3043);
or OR4 (N3061, N3056, N1656, N2432, N2087);
buf BUF1 (N3062, N3059);
and AND2 (N3063, N3048, N784);
nand NAND3 (N3064, N3061, N2788, N2057);
nor NOR3 (N3065, N3054, N161, N1813);
buf BUF1 (N3066, N3057);
nor NOR3 (N3067, N3040, N373, N1043);
or OR3 (N3068, N3058, N2989, N2264);
nand NAND4 (N3069, N3065, N2194, N1832, N1176);
xor XOR2 (N3070, N3060, N663);
or OR4 (N3071, N3062, N2259, N1512, N1165);
buf BUF1 (N3072, N3063);
not NOT1 (N3073, N3067);
not NOT1 (N3074, N3064);
or OR3 (N3075, N3071, N286, N1953);
nor NOR2 (N3076, N3075, N382);
and AND4 (N3077, N3072, N1222, N1139, N1444);
nor NOR3 (N3078, N3077, N925, N523);
nand NAND2 (N3079, N3070, N2311);
or OR2 (N3080, N3079, N743);
or OR4 (N3081, N3076, N2957, N2975, N528);
not NOT1 (N3082, N3080);
and AND3 (N3083, N3068, N2509, N619);
nor NOR4 (N3084, N3083, N2043, N2625, N2416);
not NOT1 (N3085, N3081);
not NOT1 (N3086, N3069);
or OR3 (N3087, N3033, N2407, N2208);
or OR2 (N3088, N3085, N2182);
or OR4 (N3089, N3082, N617, N300, N1012);
and AND4 (N3090, N3086, N414, N58, N975);
or OR2 (N3091, N3066, N2243);
buf BUF1 (N3092, N3074);
nand NAND3 (N3093, N3078, N1707, N2807);
buf BUF1 (N3094, N3089);
buf BUF1 (N3095, N3051);
nand NAND4 (N3096, N3094, N1086, N923, N1018);
nand NAND4 (N3097, N3093, N1682, N3029, N688);
or OR4 (N3098, N3088, N2407, N2124, N1324);
not NOT1 (N3099, N3096);
xor XOR2 (N3100, N3090, N1403);
xor XOR2 (N3101, N3097, N2988);
not NOT1 (N3102, N3084);
or OR4 (N3103, N3087, N2430, N2974, N193);
or OR2 (N3104, N3100, N1007);
and AND2 (N3105, N3101, N2141);
xor XOR2 (N3106, N3099, N2178);
and AND4 (N3107, N3106, N1063, N1073, N1807);
and AND3 (N3108, N3104, N861, N1322);
or OR4 (N3109, N3103, N2543, N397, N2758);
nor NOR2 (N3110, N3107, N1972);
xor XOR2 (N3111, N3102, N508);
buf BUF1 (N3112, N3111);
nor NOR3 (N3113, N3091, N1279, N2495);
not NOT1 (N3114, N3113);
nand NAND4 (N3115, N3073, N2133, N1317, N1233);
xor XOR2 (N3116, N3112, N1330);
nor NOR3 (N3117, N3115, N644, N3047);
or OR3 (N3118, N3117, N516, N1615);
nor NOR4 (N3119, N3092, N2161, N2512, N1451);
nor NOR2 (N3120, N3119, N1043);
or OR3 (N3121, N3116, N2641, N3103);
xor XOR2 (N3122, N3110, N2033);
not NOT1 (N3123, N3120);
buf BUF1 (N3124, N3105);
nor NOR3 (N3125, N3098, N908, N1162);
nor NOR2 (N3126, N3118, N725);
and AND4 (N3127, N3124, N329, N2750, N3025);
not NOT1 (N3128, N3126);
not NOT1 (N3129, N3108);
nor NOR4 (N3130, N3122, N717, N479, N1212);
nor NOR4 (N3131, N3109, N58, N16, N1195);
or OR4 (N3132, N3121, N1499, N1009, N2590);
and AND4 (N3133, N3128, N1505, N3046, N2534);
nor NOR3 (N3134, N3131, N1568, N799);
not NOT1 (N3135, N3129);
not NOT1 (N3136, N3133);
nor NOR4 (N3137, N3132, N3073, N2492, N233);
xor XOR2 (N3138, N3135, N3100);
nand NAND4 (N3139, N3114, N3027, N531, N2724);
nor NOR2 (N3140, N3134, N2527);
nor NOR2 (N3141, N3138, N1716);
xor XOR2 (N3142, N3140, N1140);
not NOT1 (N3143, N3095);
or OR4 (N3144, N3136, N1956, N1359, N1450);
and AND3 (N3145, N3143, N1741, N2946);
buf BUF1 (N3146, N3139);
buf BUF1 (N3147, N3144);
nor NOR4 (N3148, N3125, N1849, N1312, N1389);
buf BUF1 (N3149, N3123);
buf BUF1 (N3150, N3130);
nand NAND3 (N3151, N3147, N581, N1113);
not NOT1 (N3152, N3149);
nor NOR4 (N3153, N3127, N1459, N1228, N1448);
nand NAND3 (N3154, N3146, N570, N3096);
nand NAND2 (N3155, N3152, N780);
xor XOR2 (N3156, N3148, N390);
nand NAND2 (N3157, N3151, N3040);
nor NOR4 (N3158, N3154, N3051, N383, N1211);
buf BUF1 (N3159, N3142);
buf BUF1 (N3160, N3153);
buf BUF1 (N3161, N3141);
buf BUF1 (N3162, N3159);
buf BUF1 (N3163, N3161);
or OR3 (N3164, N3156, N375, N2733);
and AND2 (N3165, N3155, N2964);
nor NOR2 (N3166, N3160, N1956);
nor NOR3 (N3167, N3164, N1914, N1391);
nor NOR2 (N3168, N3163, N403);
nand NAND3 (N3169, N3157, N2759, N2547);
and AND3 (N3170, N3158, N918, N1527);
nand NAND4 (N3171, N3170, N2126, N93, N1956);
buf BUF1 (N3172, N3167);
or OR3 (N3173, N3172, N2382, N3159);
buf BUF1 (N3174, N3173);
and AND3 (N3175, N3171, N2300, N101);
xor XOR2 (N3176, N3165, N2111);
xor XOR2 (N3177, N3166, N2706);
nor NOR2 (N3178, N3176, N878);
or OR4 (N3179, N3177, N403, N2851, N904);
xor XOR2 (N3180, N3179, N1833);
buf BUF1 (N3181, N3162);
buf BUF1 (N3182, N3178);
and AND3 (N3183, N3181, N1719, N3118);
and AND4 (N3184, N3137, N2520, N2412, N1143);
nand NAND4 (N3185, N3150, N2760, N1813, N908);
xor XOR2 (N3186, N3183, N1094);
nand NAND4 (N3187, N3174, N3091, N2370, N865);
buf BUF1 (N3188, N3185);
xor XOR2 (N3189, N3145, N3051);
xor XOR2 (N3190, N3186, N687);
nand NAND2 (N3191, N3180, N1483);
nand NAND4 (N3192, N3191, N44, N2226, N2312);
and AND2 (N3193, N3169, N1028);
nand NAND4 (N3194, N3190, N2529, N2871, N227);
or OR3 (N3195, N3184, N1744, N18);
buf BUF1 (N3196, N3195);
or OR3 (N3197, N3168, N847, N3116);
nand NAND2 (N3198, N3189, N2824);
not NOT1 (N3199, N3182);
xor XOR2 (N3200, N3194, N141);
or OR3 (N3201, N3187, N1396, N2576);
and AND3 (N3202, N3188, N127, N2780);
or OR2 (N3203, N3196, N1646);
and AND2 (N3204, N3192, N2786);
and AND4 (N3205, N3203, N1921, N996, N3180);
not NOT1 (N3206, N3175);
nand NAND3 (N3207, N3201, N1548, N207);
xor XOR2 (N3208, N3193, N972);
nand NAND3 (N3209, N3199, N1901, N2556);
buf BUF1 (N3210, N3197);
xor XOR2 (N3211, N3210, N517);
or OR3 (N3212, N3208, N1931, N1492);
xor XOR2 (N3213, N3206, N1607);
not NOT1 (N3214, N3200);
nand NAND2 (N3215, N3207, N2979);
and AND3 (N3216, N3202, N1803, N1672);
or OR2 (N3217, N3213, N2897);
and AND4 (N3218, N3216, N3144, N989, N2014);
not NOT1 (N3219, N3205);
buf BUF1 (N3220, N3204);
nor NOR3 (N3221, N3217, N144, N2353);
not NOT1 (N3222, N3214);
not NOT1 (N3223, N3218);
buf BUF1 (N3224, N3211);
or OR2 (N3225, N3224, N2735);
buf BUF1 (N3226, N3215);
nand NAND3 (N3227, N3220, N857, N1175);
nand NAND2 (N3228, N3221, N2859);
nor NOR3 (N3229, N3227, N249, N496);
not NOT1 (N3230, N3219);
buf BUF1 (N3231, N3225);
and AND2 (N3232, N3226, N171);
or OR3 (N3233, N3209, N2394, N2669);
xor XOR2 (N3234, N3228, N531);
not NOT1 (N3235, N3234);
buf BUF1 (N3236, N3235);
xor XOR2 (N3237, N3212, N941);
or OR2 (N3238, N3229, N2301);
or OR3 (N3239, N3238, N660, N1038);
not NOT1 (N3240, N3198);
nor NOR3 (N3241, N3236, N1045, N2969);
nor NOR4 (N3242, N3222, N346, N2330, N3);
and AND3 (N3243, N3232, N603, N56);
and AND3 (N3244, N3231, N2803, N1016);
not NOT1 (N3245, N3230);
xor XOR2 (N3246, N3243, N1270);
or OR4 (N3247, N3244, N2709, N2117, N2638);
or OR2 (N3248, N3240, N1450);
not NOT1 (N3249, N3241);
nor NOR4 (N3250, N3242, N2712, N1232, N424);
nor NOR4 (N3251, N3245, N2618, N1872, N2974);
buf BUF1 (N3252, N3251);
buf BUF1 (N3253, N3233);
buf BUF1 (N3254, N3252);
nand NAND4 (N3255, N3249, N2613, N3092, N1184);
nand NAND4 (N3256, N3247, N2872, N3190, N2041);
nand NAND2 (N3257, N3255, N1653);
and AND4 (N3258, N3257, N620, N555, N778);
not NOT1 (N3259, N3239);
and AND2 (N3260, N3259, N770);
nand NAND3 (N3261, N3253, N2759, N2382);
not NOT1 (N3262, N3248);
xor XOR2 (N3263, N3254, N2227);
nor NOR4 (N3264, N3261, N148, N3245, N708);
or OR2 (N3265, N3237, N2931);
buf BUF1 (N3266, N3223);
and AND2 (N3267, N3263, N1736);
not NOT1 (N3268, N3265);
nand NAND2 (N3269, N3262, N2185);
or OR4 (N3270, N3266, N1880, N2169, N2209);
not NOT1 (N3271, N3269);
and AND2 (N3272, N3250, N1441);
xor XOR2 (N3273, N3272, N1609);
not NOT1 (N3274, N3258);
xor XOR2 (N3275, N3264, N1388);
not NOT1 (N3276, N3267);
not NOT1 (N3277, N3276);
and AND2 (N3278, N3273, N2007);
buf BUF1 (N3279, N3256);
nor NOR4 (N3280, N3278, N1384, N911, N1705);
and AND4 (N3281, N3274, N2579, N321, N254);
not NOT1 (N3282, N3277);
not NOT1 (N3283, N3281);
or OR4 (N3284, N3283, N2468, N703, N2183);
buf BUF1 (N3285, N3271);
xor XOR2 (N3286, N3279, N2);
nor NOR3 (N3287, N3260, N1285, N2204);
and AND3 (N3288, N3282, N557, N1403);
xor XOR2 (N3289, N3246, N128);
buf BUF1 (N3290, N3289);
nor NOR2 (N3291, N3268, N777);
buf BUF1 (N3292, N3288);
nor NOR4 (N3293, N3280, N2801, N2386, N2750);
buf BUF1 (N3294, N3287);
and AND2 (N3295, N3285, N2845);
and AND4 (N3296, N3275, N2347, N3010, N558);
nand NAND2 (N3297, N3286, N462);
nand NAND3 (N3298, N3284, N288, N1609);
nor NOR4 (N3299, N3291, N4, N3175, N2501);
nor NOR2 (N3300, N3299, N1930);
buf BUF1 (N3301, N3298);
xor XOR2 (N3302, N3292, N1759);
and AND3 (N3303, N3301, N461, N2158);
nand NAND2 (N3304, N3303, N1679);
buf BUF1 (N3305, N3290);
and AND4 (N3306, N3305, N1267, N3040, N1047);
not NOT1 (N3307, N3294);
not NOT1 (N3308, N3300);
and AND4 (N3309, N3297, N3229, N2761, N558);
nor NOR3 (N3310, N3308, N1664, N1318);
buf BUF1 (N3311, N3310);
and AND4 (N3312, N3296, N620, N777, N2979);
nor NOR3 (N3313, N3306, N1493, N763);
not NOT1 (N3314, N3302);
or OR3 (N3315, N3304, N404, N752);
and AND2 (N3316, N3270, N2585);
or OR4 (N3317, N3316, N462, N3098, N1311);
xor XOR2 (N3318, N3293, N2933);
nor NOR2 (N3319, N3318, N882);
nor NOR2 (N3320, N3307, N459);
not NOT1 (N3321, N3313);
nor NOR4 (N3322, N3309, N1538, N2559, N1026);
nand NAND2 (N3323, N3314, N886);
and AND2 (N3324, N3312, N610);
or OR3 (N3325, N3317, N2413, N2114);
not NOT1 (N3326, N3311);
not NOT1 (N3327, N3324);
buf BUF1 (N3328, N3327);
and AND3 (N3329, N3319, N3185, N330);
and AND2 (N3330, N3295, N1799);
or OR2 (N3331, N3328, N1453);
buf BUF1 (N3332, N3321);
nor NOR4 (N3333, N3331, N2014, N2330, N1284);
buf BUF1 (N3334, N3320);
not NOT1 (N3335, N3323);
nand NAND3 (N3336, N3334, N2148, N1381);
nor NOR4 (N3337, N3332, N1044, N141, N2777);
nand NAND4 (N3338, N3337, N2627, N26, N1898);
not NOT1 (N3339, N3336);
and AND4 (N3340, N3315, N1128, N2361, N867);
or OR3 (N3341, N3340, N63, N692);
xor XOR2 (N3342, N3341, N1977);
and AND3 (N3343, N3339, N2093, N2563);
and AND4 (N3344, N3342, N123, N2019, N847);
and AND2 (N3345, N3343, N1253);
and AND3 (N3346, N3326, N1124, N1395);
or OR4 (N3347, N3325, N989, N1147, N3155);
not NOT1 (N3348, N3346);
and AND4 (N3349, N3329, N3317, N3277, N1616);
xor XOR2 (N3350, N3335, N1919);
or OR2 (N3351, N3344, N1049);
not NOT1 (N3352, N3350);
not NOT1 (N3353, N3352);
nand NAND4 (N3354, N3333, N603, N3149, N2453);
nor NOR4 (N3355, N3347, N985, N2471, N3053);
not NOT1 (N3356, N3338);
or OR2 (N3357, N3330, N1713);
nand NAND4 (N3358, N3351, N2962, N43, N1285);
and AND4 (N3359, N3322, N2136, N2458, N3254);
buf BUF1 (N3360, N3355);
nor NOR4 (N3361, N3348, N1572, N3097, N1513);
xor XOR2 (N3362, N3359, N1080);
nor NOR4 (N3363, N3361, N495, N759, N870);
nor NOR2 (N3364, N3345, N1176);
nand NAND2 (N3365, N3349, N1448);
nand NAND4 (N3366, N3360, N1366, N2882, N1840);
nand NAND3 (N3367, N3365, N3269, N1566);
nor NOR3 (N3368, N3357, N2238, N3141);
nor NOR3 (N3369, N3368, N299, N3272);
nor NOR4 (N3370, N3362, N2344, N57, N1223);
not NOT1 (N3371, N3364);
not NOT1 (N3372, N3356);
xor XOR2 (N3373, N3371, N2376);
and AND3 (N3374, N3370, N2453, N1726);
and AND4 (N3375, N3353, N1150, N904, N1726);
and AND3 (N3376, N3372, N854, N1311);
xor XOR2 (N3377, N3354, N3337);
and AND4 (N3378, N3376, N116, N726, N761);
and AND2 (N3379, N3374, N3165);
not NOT1 (N3380, N3373);
xor XOR2 (N3381, N3366, N1111);
nand NAND3 (N3382, N3378, N2979, N1683);
buf BUF1 (N3383, N3369);
and AND4 (N3384, N3381, N2131, N2219, N2296);
or OR3 (N3385, N3383, N2959, N5);
buf BUF1 (N3386, N3363);
xor XOR2 (N3387, N3377, N2669);
nand NAND4 (N3388, N3367, N1504, N3342, N1930);
not NOT1 (N3389, N3380);
buf BUF1 (N3390, N3384);
not NOT1 (N3391, N3389);
xor XOR2 (N3392, N3375, N1920);
nor NOR3 (N3393, N3382, N2613, N674);
or OR4 (N3394, N3358, N1054, N270, N701);
not NOT1 (N3395, N3379);
nor NOR3 (N3396, N3390, N1910, N1192);
buf BUF1 (N3397, N3393);
nand NAND2 (N3398, N3388, N2479);
buf BUF1 (N3399, N3396);
nor NOR2 (N3400, N3397, N3376);
and AND2 (N3401, N3385, N3047);
nor NOR3 (N3402, N3398, N1643, N953);
and AND3 (N3403, N3392, N1964, N3396);
not NOT1 (N3404, N3395);
and AND2 (N3405, N3404, N1433);
and AND4 (N3406, N3401, N210, N2434, N2407);
nand NAND2 (N3407, N3403, N2380);
not NOT1 (N3408, N3402);
and AND2 (N3409, N3387, N2782);
xor XOR2 (N3410, N3394, N711);
not NOT1 (N3411, N3410);
and AND2 (N3412, N3407, N3312);
buf BUF1 (N3413, N3412);
or OR2 (N3414, N3405, N2260);
not NOT1 (N3415, N3391);
nand NAND2 (N3416, N3386, N342);
not NOT1 (N3417, N3415);
xor XOR2 (N3418, N3416, N907);
buf BUF1 (N3419, N3414);
not NOT1 (N3420, N3417);
xor XOR2 (N3421, N3420, N1246);
nor NOR2 (N3422, N3400, N266);
nand NAND2 (N3423, N3418, N421);
buf BUF1 (N3424, N3422);
nor NOR4 (N3425, N3419, N3178, N581, N1272);
not NOT1 (N3426, N3411);
buf BUF1 (N3427, N3399);
or OR3 (N3428, N3408, N307, N2457);
nand NAND4 (N3429, N3428, N2909, N610, N371);
nor NOR2 (N3430, N3425, N2938);
nor NOR2 (N3431, N3423, N2211);
nor NOR2 (N3432, N3429, N2646);
xor XOR2 (N3433, N3406, N745);
or OR4 (N3434, N3424, N94, N2623, N3094);
not NOT1 (N3435, N3432);
not NOT1 (N3436, N3431);
or OR3 (N3437, N3427, N2949, N1583);
nand NAND4 (N3438, N3436, N2686, N2058, N1232);
nand NAND3 (N3439, N3426, N1030, N3232);
nor NOR3 (N3440, N3430, N609, N51);
nor NOR3 (N3441, N3438, N1758, N488);
buf BUF1 (N3442, N3409);
nand NAND3 (N3443, N3439, N2101, N226);
not NOT1 (N3444, N3434);
buf BUF1 (N3445, N3433);
and AND3 (N3446, N3437, N1325, N1898);
or OR3 (N3447, N3442, N1567, N509);
not NOT1 (N3448, N3435);
buf BUF1 (N3449, N3441);
nand NAND3 (N3450, N3443, N2111, N1222);
or OR3 (N3451, N3450, N867, N775);
or OR3 (N3452, N3449, N1460, N2270);
nor NOR4 (N3453, N3445, N2629, N2164, N3017);
xor XOR2 (N3454, N3447, N645);
nor NOR2 (N3455, N3421, N927);
and AND4 (N3456, N3453, N2523, N1126, N3127);
nor NOR4 (N3457, N3454, N37, N77, N1920);
and AND2 (N3458, N3440, N2331);
not NOT1 (N3459, N3446);
not NOT1 (N3460, N3459);
not NOT1 (N3461, N3448);
buf BUF1 (N3462, N3444);
not NOT1 (N3463, N3461);
xor XOR2 (N3464, N3460, N2620);
nand NAND2 (N3465, N3463, N291);
nor NOR2 (N3466, N3455, N2517);
not NOT1 (N3467, N3458);
xor XOR2 (N3468, N3451, N1336);
xor XOR2 (N3469, N3462, N1817);
nand NAND4 (N3470, N3464, N182, N1462, N2334);
or OR3 (N3471, N3469, N2099, N2047);
buf BUF1 (N3472, N3466);
xor XOR2 (N3473, N3452, N393);
xor XOR2 (N3474, N3471, N2218);
nor NOR4 (N3475, N3457, N580, N1344, N2124);
or OR2 (N3476, N3472, N866);
nor NOR2 (N3477, N3467, N1262);
xor XOR2 (N3478, N3477, N2404);
and AND2 (N3479, N3476, N1348);
xor XOR2 (N3480, N3474, N198);
nand NAND3 (N3481, N3456, N2394, N381);
and AND4 (N3482, N3480, N3415, N525, N894);
xor XOR2 (N3483, N3473, N2147);
and AND4 (N3484, N3468, N2311, N2153, N2529);
not NOT1 (N3485, N3470);
nor NOR4 (N3486, N3484, N2275, N2420, N1733);
nor NOR4 (N3487, N3479, N668, N1371, N619);
or OR2 (N3488, N3481, N2634);
xor XOR2 (N3489, N3465, N1891);
xor XOR2 (N3490, N3489, N460);
nand NAND3 (N3491, N3482, N2608, N1690);
buf BUF1 (N3492, N3478);
and AND3 (N3493, N3492, N2298, N455);
or OR3 (N3494, N3488, N1710, N1344);
or OR4 (N3495, N3490, N1248, N1039, N2170);
and AND3 (N3496, N3491, N992, N815);
nand NAND2 (N3497, N3486, N2482);
buf BUF1 (N3498, N3475);
or OR3 (N3499, N3494, N2084, N2411);
nand NAND2 (N3500, N3487, N2391);
nand NAND4 (N3501, N3485, N2334, N259, N207);
nor NOR2 (N3502, N3493, N384);
nor NOR3 (N3503, N3413, N2571, N2022);
nor NOR2 (N3504, N3502, N12);
xor XOR2 (N3505, N3501, N670);
not NOT1 (N3506, N3504);
xor XOR2 (N3507, N3495, N2413);
nand NAND2 (N3508, N3499, N816);
buf BUF1 (N3509, N3498);
not NOT1 (N3510, N3506);
not NOT1 (N3511, N3500);
nor NOR2 (N3512, N3503, N3022);
and AND4 (N3513, N3496, N2166, N1108, N1042);
xor XOR2 (N3514, N3513, N158);
nor NOR2 (N3515, N3514, N1580);
buf BUF1 (N3516, N3512);
or OR3 (N3517, N3508, N389, N2170);
nor NOR2 (N3518, N3510, N2938);
not NOT1 (N3519, N3497);
xor XOR2 (N3520, N3518, N243);
and AND4 (N3521, N3520, N93, N2622, N1766);
nand NAND3 (N3522, N3516, N2983, N1585);
xor XOR2 (N3523, N3519, N1214);
xor XOR2 (N3524, N3509, N1651);
xor XOR2 (N3525, N3507, N1092);
nand NAND4 (N3526, N3523, N492, N2016, N2087);
nand NAND4 (N3527, N3483, N1133, N2248, N1413);
and AND2 (N3528, N3521, N691);
nand NAND3 (N3529, N3517, N131, N1814);
nand NAND4 (N3530, N3522, N2720, N28, N2499);
buf BUF1 (N3531, N3525);
nor NOR3 (N3532, N3531, N1773, N2805);
xor XOR2 (N3533, N3532, N1240);
or OR4 (N3534, N3511, N765, N529, N3342);
xor XOR2 (N3535, N3530, N1809);
xor XOR2 (N3536, N3524, N3116);
buf BUF1 (N3537, N3515);
and AND2 (N3538, N3533, N257);
nor NOR3 (N3539, N3527, N1735, N3284);
and AND3 (N3540, N3537, N801, N1111);
buf BUF1 (N3541, N3529);
buf BUF1 (N3542, N3534);
nor NOR2 (N3543, N3528, N3147);
not NOT1 (N3544, N3538);
not NOT1 (N3545, N3535);
not NOT1 (N3546, N3540);
nor NOR3 (N3547, N3539, N1004, N1609);
buf BUF1 (N3548, N3544);
buf BUF1 (N3549, N3547);
nor NOR3 (N3550, N3545, N420, N2245);
buf BUF1 (N3551, N3550);
nand NAND3 (N3552, N3549, N2395, N2929);
buf BUF1 (N3553, N3552);
and AND3 (N3554, N3553, N2974, N1737);
nor NOR4 (N3555, N3543, N403, N984, N1089);
not NOT1 (N3556, N3541);
and AND2 (N3557, N3546, N185);
xor XOR2 (N3558, N3556, N1021);
or OR2 (N3559, N3554, N2311);
nor NOR2 (N3560, N3557, N742);
nor NOR3 (N3561, N3558, N3453, N3108);
nor NOR2 (N3562, N3559, N1687);
or OR3 (N3563, N3562, N143, N1826);
xor XOR2 (N3564, N3548, N2443);
or OR2 (N3565, N3563, N1268);
and AND3 (N3566, N3561, N1948, N764);
not NOT1 (N3567, N3526);
xor XOR2 (N3568, N3560, N980);
not NOT1 (N3569, N3564);
nand NAND2 (N3570, N3551, N1056);
xor XOR2 (N3571, N3568, N1113);
nor NOR4 (N3572, N3505, N2867, N312, N277);
or OR2 (N3573, N3555, N1609);
and AND3 (N3574, N3570, N1787, N3055);
nor NOR2 (N3575, N3572, N2936);
or OR4 (N3576, N3575, N1176, N3384, N1300);
not NOT1 (N3577, N3542);
and AND4 (N3578, N3573, N2963, N3227, N2215);
xor XOR2 (N3579, N3567, N991);
buf BUF1 (N3580, N3578);
nand NAND3 (N3581, N3565, N1299, N3053);
and AND3 (N3582, N3581, N2303, N391);
or OR3 (N3583, N3574, N3125, N120);
xor XOR2 (N3584, N3577, N1731);
or OR3 (N3585, N3571, N2443, N1967);
and AND3 (N3586, N3585, N3582, N433);
nor NOR2 (N3587, N3358, N2580);
buf BUF1 (N3588, N3566);
or OR4 (N3589, N3536, N448, N3571, N1404);
and AND2 (N3590, N3569, N3372);
or OR2 (N3591, N3589, N3209);
or OR4 (N3592, N3588, N2753, N864, N1235);
or OR2 (N3593, N3590, N2055);
or OR2 (N3594, N3593, N3441);
buf BUF1 (N3595, N3579);
and AND2 (N3596, N3594, N2703);
and AND2 (N3597, N3583, N775);
buf BUF1 (N3598, N3591);
buf BUF1 (N3599, N3587);
nor NOR3 (N3600, N3599, N3201, N797);
nand NAND4 (N3601, N3592, N3235, N1656, N2332);
nor NOR3 (N3602, N3595, N2045, N108);
nand NAND3 (N3603, N3586, N247, N707);
nand NAND3 (N3604, N3596, N817, N1244);
and AND3 (N3605, N3597, N3342, N3206);
or OR4 (N3606, N3603, N2863, N46, N3252);
not NOT1 (N3607, N3584);
buf BUF1 (N3608, N3607);
and AND4 (N3609, N3606, N2885, N286, N1169);
buf BUF1 (N3610, N3605);
nand NAND4 (N3611, N3601, N455, N3049, N180);
nand NAND2 (N3612, N3600, N91);
xor XOR2 (N3613, N3598, N558);
or OR4 (N3614, N3609, N392, N3291, N1037);
nor NOR2 (N3615, N3612, N1308);
nor NOR3 (N3616, N3580, N2142, N3064);
nor NOR4 (N3617, N3615, N3490, N2572, N2636);
or OR2 (N3618, N3604, N2988);
not NOT1 (N3619, N3610);
xor XOR2 (N3620, N3614, N260);
and AND2 (N3621, N3602, N756);
nor NOR2 (N3622, N3616, N435);
and AND2 (N3623, N3608, N2772);
nor NOR4 (N3624, N3619, N924, N744, N1072);
nand NAND3 (N3625, N3611, N2624, N3138);
buf BUF1 (N3626, N3618);
not NOT1 (N3627, N3613);
nand NAND3 (N3628, N3624, N1008, N267);
not NOT1 (N3629, N3576);
or OR3 (N3630, N3625, N103, N1823);
buf BUF1 (N3631, N3617);
or OR2 (N3632, N3623, N2587);
not NOT1 (N3633, N3628);
or OR4 (N3634, N3631, N124, N993, N3206);
buf BUF1 (N3635, N3629);
xor XOR2 (N3636, N3626, N2448);
buf BUF1 (N3637, N3627);
and AND3 (N3638, N3637, N3002, N3618);
xor XOR2 (N3639, N3622, N1290);
nor NOR3 (N3640, N3633, N3425, N3540);
buf BUF1 (N3641, N3638);
xor XOR2 (N3642, N3621, N368);
and AND2 (N3643, N3636, N1758);
xor XOR2 (N3644, N3639, N3246);
and AND3 (N3645, N3640, N2082, N1354);
and AND4 (N3646, N3635, N2513, N3516, N2069);
and AND2 (N3647, N3620, N1895);
and AND3 (N3648, N3646, N1930, N575);
and AND4 (N3649, N3634, N3589, N1412, N12);
and AND3 (N3650, N3645, N3009, N3208);
and AND3 (N3651, N3642, N2112, N3115);
or OR3 (N3652, N3651, N1130, N1220);
xor XOR2 (N3653, N3650, N689);
nand NAND2 (N3654, N3632, N786);
buf BUF1 (N3655, N3654);
or OR4 (N3656, N3655, N2368, N65, N1173);
nand NAND2 (N3657, N3653, N1192);
nand NAND3 (N3658, N3652, N1938, N3329);
not NOT1 (N3659, N3644);
nor NOR4 (N3660, N3630, N1286, N2502, N1583);
nor NOR2 (N3661, N3643, N1560);
nor NOR3 (N3662, N3660, N506, N2209);
buf BUF1 (N3663, N3662);
buf BUF1 (N3664, N3656);
and AND3 (N3665, N3649, N2537, N2590);
or OR3 (N3666, N3648, N710, N994);
not NOT1 (N3667, N3663);
nand NAND4 (N3668, N3657, N163, N1239, N1969);
nand NAND3 (N3669, N3666, N961, N905);
and AND4 (N3670, N3668, N376, N2933, N2274);
xor XOR2 (N3671, N3659, N2100);
nor NOR3 (N3672, N3671, N2577, N154);
xor XOR2 (N3673, N3672, N2717);
xor XOR2 (N3674, N3658, N2480);
not NOT1 (N3675, N3661);
buf BUF1 (N3676, N3674);
nand NAND3 (N3677, N3647, N78, N1466);
or OR2 (N3678, N3677, N2034);
xor XOR2 (N3679, N3675, N1647);
and AND3 (N3680, N3667, N2868, N1726);
buf BUF1 (N3681, N3678);
xor XOR2 (N3682, N3670, N1587);
nor NOR4 (N3683, N3669, N1445, N885, N2188);
buf BUF1 (N3684, N3680);
nor NOR4 (N3685, N3684, N2101, N921, N3551);
xor XOR2 (N3686, N3664, N994);
nor NOR4 (N3687, N3685, N126, N1878, N537);
nand NAND4 (N3688, N3681, N835, N3490, N2988);
buf BUF1 (N3689, N3686);
or OR3 (N3690, N3641, N3647, N2348);
and AND3 (N3691, N3683, N1706, N1235);
not NOT1 (N3692, N3690);
or OR2 (N3693, N3673, N2389);
xor XOR2 (N3694, N3687, N2084);
or OR4 (N3695, N3689, N3566, N163, N2989);
nor NOR3 (N3696, N3679, N806, N1982);
nor NOR4 (N3697, N3696, N1607, N834, N135);
buf BUF1 (N3698, N3692);
nand NAND4 (N3699, N3693, N3271, N1504, N1161);
xor XOR2 (N3700, N3695, N802);
nand NAND3 (N3701, N3682, N856, N645);
nand NAND4 (N3702, N3676, N3330, N2749, N1926);
xor XOR2 (N3703, N3699, N861);
or OR4 (N3704, N3703, N453, N2802, N107);
nand NAND2 (N3705, N3691, N92);
nor NOR3 (N3706, N3688, N2300, N87);
xor XOR2 (N3707, N3706, N2873);
nor NOR4 (N3708, N3700, N414, N2490, N2833);
nand NAND2 (N3709, N3702, N1647);
nor NOR2 (N3710, N3697, N1990);
nand NAND4 (N3711, N3698, N2812, N687, N3465);
xor XOR2 (N3712, N3711, N2133);
and AND3 (N3713, N3705, N3451, N3482);
nand NAND2 (N3714, N3710, N1799);
nor NOR4 (N3715, N3704, N2007, N3497, N3303);
not NOT1 (N3716, N3694);
buf BUF1 (N3717, N3708);
nor NOR2 (N3718, N3715, N2192);
not NOT1 (N3719, N3707);
nor NOR4 (N3720, N3709, N2019, N1938, N2895);
nor NOR4 (N3721, N3665, N2000, N2152, N2463);
or OR4 (N3722, N3716, N3652, N1238, N786);
or OR2 (N3723, N3720, N1906);
buf BUF1 (N3724, N3723);
nor NOR3 (N3725, N3721, N2515, N1985);
buf BUF1 (N3726, N3718);
or OR2 (N3727, N3724, N305);
xor XOR2 (N3728, N3712, N188);
buf BUF1 (N3729, N3719);
xor XOR2 (N3730, N3725, N1665);
not NOT1 (N3731, N3730);
nand NAND2 (N3732, N3713, N3480);
and AND3 (N3733, N3701, N787, N2655);
nor NOR3 (N3734, N3727, N1277, N1826);
or OR4 (N3735, N3717, N3291, N1351, N822);
xor XOR2 (N3736, N3735, N3064);
or OR2 (N3737, N3734, N173);
nand NAND2 (N3738, N3714, N98);
buf BUF1 (N3739, N3733);
nor NOR3 (N3740, N3737, N738, N1604);
or OR2 (N3741, N3729, N2122);
not NOT1 (N3742, N3731);
not NOT1 (N3743, N3739);
nand NAND2 (N3744, N3741, N3481);
nand NAND3 (N3745, N3732, N1178, N1550);
and AND4 (N3746, N3743, N2226, N3180, N3248);
or OR4 (N3747, N3744, N2907, N406, N58);
buf BUF1 (N3748, N3736);
and AND3 (N3749, N3747, N1641, N2724);
xor XOR2 (N3750, N3746, N1584);
buf BUF1 (N3751, N3722);
or OR4 (N3752, N3748, N1329, N2705, N2969);
xor XOR2 (N3753, N3745, N1129);
not NOT1 (N3754, N3750);
or OR4 (N3755, N3749, N1105, N3524, N3005);
not NOT1 (N3756, N3754);
xor XOR2 (N3757, N3740, N229);
and AND3 (N3758, N3757, N2648, N2086);
nor NOR4 (N3759, N3752, N3681, N2136, N679);
or OR3 (N3760, N3753, N3000, N864);
not NOT1 (N3761, N3728);
or OR2 (N3762, N3756, N2677);
and AND3 (N3763, N3759, N2939, N1366);
or OR4 (N3764, N3755, N1208, N1569, N3005);
xor XOR2 (N3765, N3758, N3623);
not NOT1 (N3766, N3765);
and AND2 (N3767, N3766, N3414);
or OR2 (N3768, N3751, N1773);
and AND3 (N3769, N3768, N2304, N1113);
nor NOR4 (N3770, N3764, N672, N3439, N293);
buf BUF1 (N3771, N3767);
and AND2 (N3772, N3738, N2932);
not NOT1 (N3773, N3769);
nand NAND4 (N3774, N3772, N2413, N3177, N935);
nor NOR3 (N3775, N3761, N3592, N2658);
and AND2 (N3776, N3760, N1304);
buf BUF1 (N3777, N3774);
and AND4 (N3778, N3762, N2821, N2361, N1942);
or OR2 (N3779, N3771, N1034);
xor XOR2 (N3780, N3726, N1981);
and AND2 (N3781, N3770, N1255);
buf BUF1 (N3782, N3778);
not NOT1 (N3783, N3775);
nor NOR4 (N3784, N3783, N565, N1176, N1322);
xor XOR2 (N3785, N3742, N2819);
not NOT1 (N3786, N3784);
nand NAND2 (N3787, N3785, N1377);
not NOT1 (N3788, N3773);
and AND2 (N3789, N3777, N2749);
and AND3 (N3790, N3781, N3658, N1041);
or OR3 (N3791, N3763, N1566, N792);
not NOT1 (N3792, N3779);
or OR3 (N3793, N3782, N3091, N2903);
and AND3 (N3794, N3776, N1963, N2363);
nand NAND3 (N3795, N3780, N1629, N3390);
and AND3 (N3796, N3788, N2004, N3027);
xor XOR2 (N3797, N3786, N804);
buf BUF1 (N3798, N3787);
nor NOR4 (N3799, N3794, N3249, N3783, N1233);
xor XOR2 (N3800, N3797, N1712);
nor NOR3 (N3801, N3789, N1825, N794);
xor XOR2 (N3802, N3799, N2705);
or OR2 (N3803, N3798, N1463);
nand NAND4 (N3804, N3793, N697, N2105, N3620);
not NOT1 (N3805, N3791);
nand NAND2 (N3806, N3795, N836);
nor NOR4 (N3807, N3796, N3316, N1102, N3791);
nor NOR3 (N3808, N3803, N2092, N2955);
xor XOR2 (N3809, N3802, N1187);
nor NOR4 (N3810, N3804, N463, N1629, N2479);
nor NOR4 (N3811, N3790, N2653, N1175, N2207);
not NOT1 (N3812, N3811);
nor NOR4 (N3813, N3809, N674, N67, N1022);
and AND4 (N3814, N3806, N2702, N2436, N3305);
or OR4 (N3815, N3792, N2787, N324, N1244);
nor NOR2 (N3816, N3812, N99);
nor NOR4 (N3817, N3816, N488, N3736, N508);
xor XOR2 (N3818, N3808, N1037);
nand NAND2 (N3819, N3814, N1562);
buf BUF1 (N3820, N3818);
or OR2 (N3821, N3801, N1220);
or OR3 (N3822, N3810, N2550, N3376);
not NOT1 (N3823, N3820);
or OR2 (N3824, N3805, N2571);
not NOT1 (N3825, N3819);
and AND4 (N3826, N3800, N2861, N2431, N2014);
or OR4 (N3827, N3821, N2221, N2257, N67);
nor NOR3 (N3828, N3815, N1277, N3156);
buf BUF1 (N3829, N3823);
nand NAND4 (N3830, N3813, N3218, N1929, N2513);
not NOT1 (N3831, N3807);
and AND3 (N3832, N3831, N1404, N2665);
buf BUF1 (N3833, N3832);
xor XOR2 (N3834, N3824, N1827);
nor NOR3 (N3835, N3829, N2483, N3102);
nor NOR3 (N3836, N3828, N3462, N3425);
and AND3 (N3837, N3822, N1858, N1785);
xor XOR2 (N3838, N3833, N2272);
buf BUF1 (N3839, N3830);
not NOT1 (N3840, N3817);
nor NOR4 (N3841, N3840, N3244, N2477, N2566);
nand NAND2 (N3842, N3839, N132);
buf BUF1 (N3843, N3825);
buf BUF1 (N3844, N3835);
nor NOR3 (N3845, N3838, N3753, N1714);
and AND4 (N3846, N3842, N3449, N1540, N2463);
xor XOR2 (N3847, N3834, N3307);
and AND3 (N3848, N3841, N980, N1760);
and AND4 (N3849, N3846, N656, N559, N1085);
xor XOR2 (N3850, N3827, N2505);
buf BUF1 (N3851, N3845);
or OR4 (N3852, N3836, N2554, N13, N650);
xor XOR2 (N3853, N3849, N857);
not NOT1 (N3854, N3853);
or OR2 (N3855, N3848, N2222);
or OR3 (N3856, N3843, N2141, N2971);
and AND2 (N3857, N3847, N1957);
nor NOR2 (N3858, N3854, N426);
buf BUF1 (N3859, N3850);
nor NOR2 (N3860, N3858, N3634);
nor NOR2 (N3861, N3844, N2112);
or OR3 (N3862, N3856, N2983, N2537);
xor XOR2 (N3863, N3851, N2957);
or OR2 (N3864, N3859, N3773);
xor XOR2 (N3865, N3860, N3763);
and AND3 (N3866, N3826, N2765, N1100);
xor XOR2 (N3867, N3864, N2506);
nand NAND4 (N3868, N3852, N2266, N2777, N2541);
and AND3 (N3869, N3861, N3356, N2011);
nor NOR3 (N3870, N3862, N3663, N1306);
nor NOR4 (N3871, N3868, N3652, N789, N301);
and AND2 (N3872, N3869, N3353);
or OR4 (N3873, N3870, N2046, N742, N1498);
or OR2 (N3874, N3873, N1368);
not NOT1 (N3875, N3855);
buf BUF1 (N3876, N3872);
nor NOR4 (N3877, N3875, N884, N942, N135);
xor XOR2 (N3878, N3837, N91);
and AND3 (N3879, N3867, N2090, N2584);
and AND4 (N3880, N3874, N1025, N814, N2771);
nand NAND3 (N3881, N3880, N2294, N989);
nor NOR3 (N3882, N3863, N3726, N2963);
nor NOR2 (N3883, N3877, N1720);
nand NAND4 (N3884, N3876, N3615, N3357, N1308);
xor XOR2 (N3885, N3865, N1014);
nand NAND3 (N3886, N3866, N3514, N3835);
nor NOR3 (N3887, N3884, N703, N590);
buf BUF1 (N3888, N3882);
nor NOR2 (N3889, N3883, N2949);
nand NAND4 (N3890, N3857, N2319, N1399, N3069);
nor NOR3 (N3891, N3887, N335, N532);
and AND4 (N3892, N3878, N2842, N3665, N2744);
not NOT1 (N3893, N3885);
nand NAND4 (N3894, N3871, N813, N3574, N1313);
or OR3 (N3895, N3889, N1858, N374);
nand NAND2 (N3896, N3890, N319);
nor NOR4 (N3897, N3886, N3749, N2725, N3487);
buf BUF1 (N3898, N3888);
or OR4 (N3899, N3896, N2333, N2682, N1209);
and AND4 (N3900, N3894, N201, N2289, N1052);
or OR4 (N3901, N3899, N928, N249, N651);
nor NOR2 (N3902, N3898, N1351);
nand NAND2 (N3903, N3891, N3668);
nand NAND3 (N3904, N3895, N2301, N323);
nand NAND3 (N3905, N3893, N2453, N3323);
or OR4 (N3906, N3901, N1725, N2528, N3323);
or OR3 (N3907, N3879, N383, N357);
and AND2 (N3908, N3907, N3266);
nor NOR2 (N3909, N3897, N2334);
nor NOR2 (N3910, N3904, N699);
buf BUF1 (N3911, N3905);
nand NAND4 (N3912, N3909, N1366, N2066, N1377);
and AND2 (N3913, N3900, N922);
not NOT1 (N3914, N3892);
nor NOR4 (N3915, N3912, N1789, N1911, N3680);
or OR3 (N3916, N3902, N3361, N3695);
or OR4 (N3917, N3908, N3597, N1475, N1880);
nor NOR2 (N3918, N3913, N2758);
and AND4 (N3919, N3917, N1295, N3914, N3101);
buf BUF1 (N3920, N2566);
nand NAND3 (N3921, N3911, N1054, N2093);
buf BUF1 (N3922, N3881);
nor NOR4 (N3923, N3906, N2353, N3803, N2823);
and AND3 (N3924, N3903, N2986, N3825);
nand NAND2 (N3925, N3918, N1272);
and AND2 (N3926, N3919, N1757);
and AND4 (N3927, N3910, N3776, N595, N1148);
not NOT1 (N3928, N3925);
and AND3 (N3929, N3928, N1651, N254);
buf BUF1 (N3930, N3923);
not NOT1 (N3931, N3922);
not NOT1 (N3932, N3931);
not NOT1 (N3933, N3927);
buf BUF1 (N3934, N3932);
or OR4 (N3935, N3926, N3303, N2540, N3292);
nand NAND4 (N3936, N3935, N2412, N1576, N2725);
or OR2 (N3937, N3921, N3030);
not NOT1 (N3938, N3936);
and AND4 (N3939, N3916, N2019, N237, N1240);
nor NOR2 (N3940, N3915, N293);
or OR2 (N3941, N3939, N844);
buf BUF1 (N3942, N3933);
nor NOR4 (N3943, N3924, N3796, N1983, N1137);
xor XOR2 (N3944, N3942, N3933);
and AND3 (N3945, N3943, N998, N3346);
buf BUF1 (N3946, N3944);
and AND3 (N3947, N3930, N1605, N1748);
or OR3 (N3948, N3946, N2797, N1654);
not NOT1 (N3949, N3920);
or OR2 (N3950, N3934, N197);
buf BUF1 (N3951, N3937);
not NOT1 (N3952, N3945);
xor XOR2 (N3953, N3941, N909);
nor NOR4 (N3954, N3953, N3596, N3830, N676);
nand NAND4 (N3955, N3938, N279, N353, N43);
xor XOR2 (N3956, N3948, N1296);
and AND4 (N3957, N3947, N1216, N3853, N1601);
buf BUF1 (N3958, N3940);
nand NAND4 (N3959, N3950, N955, N2403, N3011);
or OR4 (N3960, N3952, N1223, N2489, N2853);
and AND3 (N3961, N3958, N1449, N3611);
not NOT1 (N3962, N3929);
and AND2 (N3963, N3954, N248);
nor NOR4 (N3964, N3956, N1862, N630, N3520);
nand NAND2 (N3965, N3949, N2938);
not NOT1 (N3966, N3960);
xor XOR2 (N3967, N3951, N24);
or OR3 (N3968, N3959, N2038, N2870);
or OR3 (N3969, N3962, N3612, N2888);
or OR4 (N3970, N3969, N1865, N1510, N2214);
nor NOR4 (N3971, N3957, N3375, N2570, N1300);
or OR2 (N3972, N3967, N3958);
not NOT1 (N3973, N3964);
nand NAND2 (N3974, N3971, N225);
nor NOR4 (N3975, N3955, N2471, N720, N1841);
nand NAND2 (N3976, N3968, N947);
xor XOR2 (N3977, N3965, N2139);
buf BUF1 (N3978, N3963);
buf BUF1 (N3979, N3975);
nand NAND4 (N3980, N3966, N639, N2866, N1316);
xor XOR2 (N3981, N3978, N1984);
or OR2 (N3982, N3977, N903);
nor NOR4 (N3983, N3981, N203, N3271, N3509);
and AND2 (N3984, N3982, N2629);
xor XOR2 (N3985, N3961, N2722);
buf BUF1 (N3986, N3973);
buf BUF1 (N3987, N3985);
nor NOR3 (N3988, N3972, N1599, N1421);
not NOT1 (N3989, N3984);
or OR4 (N3990, N3986, N1235, N2078, N241);
or OR2 (N3991, N3987, N1393);
nand NAND2 (N3992, N3983, N1354);
nor NOR3 (N3993, N3988, N2150, N3783);
xor XOR2 (N3994, N3992, N2664);
nor NOR3 (N3995, N3976, N2947, N2753);
xor XOR2 (N3996, N3991, N1932);
nor NOR4 (N3997, N3990, N2586, N86, N198);
buf BUF1 (N3998, N3995);
and AND2 (N3999, N3974, N2568);
and AND4 (N4000, N3998, N3960, N3140, N3369);
xor XOR2 (N4001, N3997, N2849);
or OR3 (N4002, N3999, N3039, N542);
buf BUF1 (N4003, N3979);
xor XOR2 (N4004, N3994, N2150);
and AND2 (N4005, N3993, N1172);
nand NAND4 (N4006, N4002, N2186, N629, N2133);
buf BUF1 (N4007, N3970);
and AND3 (N4008, N4001, N1565, N3897);
nand NAND4 (N4009, N3996, N305, N1443, N279);
nand NAND2 (N4010, N4009, N105);
not NOT1 (N4011, N4000);
or OR3 (N4012, N4010, N1948, N2060);
nand NAND2 (N4013, N4005, N2692);
nand NAND4 (N4014, N4008, N2512, N3217, N2699);
not NOT1 (N4015, N3989);
not NOT1 (N4016, N4004);
and AND4 (N4017, N4011, N1769, N391, N1532);
or OR3 (N4018, N3980, N221, N2436);
and AND3 (N4019, N4012, N1889, N2232);
nand NAND4 (N4020, N4019, N1754, N2869, N2793);
nor NOR3 (N4021, N4016, N74, N2209);
and AND4 (N4022, N4006, N3857, N488, N585);
buf BUF1 (N4023, N4013);
not NOT1 (N4024, N4014);
nand NAND2 (N4025, N4017, N1148);
and AND3 (N4026, N4021, N1076, N800);
nor NOR4 (N4027, N4018, N778, N2824, N2885);
nand NAND2 (N4028, N4015, N4018);
or OR3 (N4029, N4026, N233, N3057);
not NOT1 (N4030, N4020);
buf BUF1 (N4031, N4024);
buf BUF1 (N4032, N4031);
or OR2 (N4033, N4028, N1057);
nand NAND3 (N4034, N4033, N3810, N1744);
buf BUF1 (N4035, N4023);
and AND3 (N4036, N4032, N2868, N747);
and AND3 (N4037, N4007, N3182, N2428);
xor XOR2 (N4038, N4035, N1184);
nand NAND4 (N4039, N4037, N965, N3809, N3478);
nor NOR4 (N4040, N4003, N1663, N3005, N1833);
xor XOR2 (N4041, N4038, N1138);
or OR3 (N4042, N4041, N1281, N2291);
nor NOR4 (N4043, N4029, N597, N3202, N381);
nor NOR4 (N4044, N4022, N1853, N1525, N1541);
or OR2 (N4045, N4040, N142);
and AND3 (N4046, N4044, N3304, N3941);
nand NAND4 (N4047, N4034, N1542, N2731, N1060);
and AND2 (N4048, N4039, N3706);
xor XOR2 (N4049, N4030, N1215);
nand NAND3 (N4050, N4036, N2294, N2617);
not NOT1 (N4051, N4046);
nand NAND4 (N4052, N4027, N507, N3983, N1077);
nor NOR4 (N4053, N4051, N113, N1567, N745);
xor XOR2 (N4054, N4053, N3918);
xor XOR2 (N4055, N4050, N3180);
not NOT1 (N4056, N4047);
and AND4 (N4057, N4045, N3238, N1085, N2684);
and AND2 (N4058, N4043, N2896);
xor XOR2 (N4059, N4056, N2211);
not NOT1 (N4060, N4052);
and AND4 (N4061, N4058, N2283, N2134, N453);
or OR4 (N4062, N4025, N3675, N806, N1589);
and AND4 (N4063, N4054, N492, N805, N981);
nand NAND3 (N4064, N4059, N3099, N904);
buf BUF1 (N4065, N4048);
or OR4 (N4066, N4061, N3591, N3597, N2306);
buf BUF1 (N4067, N4062);
or OR2 (N4068, N4065, N2269);
nor NOR4 (N4069, N4063, N706, N3514, N2202);
and AND2 (N4070, N4064, N2839);
nor NOR3 (N4071, N4060, N1196, N2552);
xor XOR2 (N4072, N4057, N3546);
and AND3 (N4073, N4071, N198, N1253);
buf BUF1 (N4074, N4049);
or OR4 (N4075, N4069, N648, N2467, N2955);
not NOT1 (N4076, N4074);
nor NOR4 (N4077, N4066, N3234, N148, N931);
nor NOR4 (N4078, N4076, N2432, N985, N1934);
xor XOR2 (N4079, N4075, N3168);
xor XOR2 (N4080, N4072, N3904);
nand NAND4 (N4081, N4079, N6, N3180, N1533);
nand NAND3 (N4082, N4070, N2172, N1803);
or OR2 (N4083, N4082, N646);
and AND3 (N4084, N4081, N441, N3228);
not NOT1 (N4085, N4083);
and AND4 (N4086, N4055, N202, N1100, N3013);
not NOT1 (N4087, N4080);
nand NAND4 (N4088, N4086, N3326, N3446, N3599);
not NOT1 (N4089, N4068);
xor XOR2 (N4090, N4084, N1081);
and AND2 (N4091, N4078, N2753);
buf BUF1 (N4092, N4090);
or OR3 (N4093, N4092, N2839, N443);
nor NOR2 (N4094, N4067, N384);
buf BUF1 (N4095, N4089);
nand NAND2 (N4096, N4087, N1008);
nor NOR2 (N4097, N4073, N3373);
nand NAND2 (N4098, N4096, N3132);
and AND4 (N4099, N4093, N3809, N1100, N3894);
xor XOR2 (N4100, N4098, N478);
xor XOR2 (N4101, N4094, N1509);
nand NAND2 (N4102, N4085, N498);
or OR3 (N4103, N4095, N1361, N3133);
buf BUF1 (N4104, N4097);
buf BUF1 (N4105, N4091);
xor XOR2 (N4106, N4104, N2881);
buf BUF1 (N4107, N4105);
not NOT1 (N4108, N4103);
nor NOR3 (N4109, N4099, N3394, N294);
or OR4 (N4110, N4088, N1219, N3496, N1568);
and AND2 (N4111, N4100, N850);
and AND4 (N4112, N4077, N3123, N1742, N2388);
nand NAND2 (N4113, N4106, N2447);
nand NAND4 (N4114, N4101, N2223, N725, N3890);
nand NAND2 (N4115, N4109, N2750);
nor NOR4 (N4116, N4110, N1218, N700, N2269);
xor XOR2 (N4117, N4114, N65);
xor XOR2 (N4118, N4117, N1987);
and AND2 (N4119, N4042, N1761);
nand NAND2 (N4120, N4119, N223);
xor XOR2 (N4121, N4116, N1204);
nor NOR4 (N4122, N4113, N2726, N3881, N1132);
buf BUF1 (N4123, N4102);
xor XOR2 (N4124, N4111, N95);
and AND3 (N4125, N4107, N3571, N2245);
not NOT1 (N4126, N4120);
nand NAND2 (N4127, N4112, N2232);
xor XOR2 (N4128, N4125, N1571);
nor NOR3 (N4129, N4127, N2404, N3449);
nand NAND4 (N4130, N4123, N3842, N627, N120);
buf BUF1 (N4131, N4129);
nor NOR4 (N4132, N4128, N1990, N2465, N3302);
xor XOR2 (N4133, N4121, N3572);
nand NAND2 (N4134, N4118, N978);
not NOT1 (N4135, N4115);
nor NOR3 (N4136, N4134, N3519, N2954);
not NOT1 (N4137, N4122);
nor NOR4 (N4138, N4135, N3348, N1972, N2261);
nor NOR2 (N4139, N4133, N736);
not NOT1 (N4140, N4126);
or OR4 (N4141, N4130, N2845, N2394, N396);
or OR2 (N4142, N4139, N1785);
buf BUF1 (N4143, N4132);
not NOT1 (N4144, N4142);
nor NOR2 (N4145, N4143, N775);
and AND2 (N4146, N4141, N2383);
xor XOR2 (N4147, N4140, N4012);
and AND4 (N4148, N4138, N1798, N1061, N1725);
and AND3 (N4149, N4146, N1402, N3537);
not NOT1 (N4150, N4137);
and AND2 (N4151, N4150, N1265);
buf BUF1 (N4152, N4145);
nand NAND2 (N4153, N4144, N3387);
xor XOR2 (N4154, N4152, N3229);
nor NOR4 (N4155, N4153, N2342, N2384, N2357);
buf BUF1 (N4156, N4155);
nor NOR2 (N4157, N4108, N3724);
nor NOR2 (N4158, N4149, N51);
or OR2 (N4159, N4124, N1146);
xor XOR2 (N4160, N4158, N3675);
or OR4 (N4161, N4159, N3146, N3311, N3852);
or OR4 (N4162, N4161, N500, N3253, N1797);
and AND3 (N4163, N4148, N2896, N165);
nor NOR3 (N4164, N4156, N1373, N1215);
xor XOR2 (N4165, N4154, N2063);
buf BUF1 (N4166, N4165);
nor NOR2 (N4167, N4163, N3034);
and AND2 (N4168, N4151, N3501);
buf BUF1 (N4169, N4167);
nor NOR4 (N4170, N4169, N3262, N2357, N4115);
nor NOR3 (N4171, N4147, N727, N3481);
or OR4 (N4172, N4171, N888, N3564, N2988);
not NOT1 (N4173, N4162);
not NOT1 (N4174, N4166);
xor XOR2 (N4175, N4174, N1218);
buf BUF1 (N4176, N4175);
nand NAND3 (N4177, N4176, N1565, N3596);
xor XOR2 (N4178, N4168, N1915);
buf BUF1 (N4179, N4178);
nor NOR4 (N4180, N4136, N3218, N3211, N1757);
xor XOR2 (N4181, N4177, N319);
buf BUF1 (N4182, N4180);
or OR3 (N4183, N4170, N3239, N1504);
nor NOR2 (N4184, N4172, N710);
and AND3 (N4185, N4181, N1321, N1824);
xor XOR2 (N4186, N4131, N3125);
xor XOR2 (N4187, N4182, N3303);
not NOT1 (N4188, N4164);
not NOT1 (N4189, N4160);
nand NAND4 (N4190, N4188, N3796, N3847, N3462);
xor XOR2 (N4191, N4189, N1716);
and AND2 (N4192, N4185, N3192);
nand NAND3 (N4193, N4190, N204, N2949);
or OR2 (N4194, N4186, N2747);
not NOT1 (N4195, N4183);
nor NOR2 (N4196, N4194, N1585);
not NOT1 (N4197, N4193);
nand NAND4 (N4198, N4195, N3293, N4176, N3984);
xor XOR2 (N4199, N4179, N2962);
nor NOR4 (N4200, N4196, N4093, N322, N4190);
and AND2 (N4201, N4187, N3986);
nor NOR4 (N4202, N4198, N1378, N2495, N3578);
nor NOR2 (N4203, N4202, N2608);
and AND4 (N4204, N4201, N3957, N3143, N2067);
or OR2 (N4205, N4157, N2231);
or OR2 (N4206, N4205, N1030);
not NOT1 (N4207, N4173);
xor XOR2 (N4208, N4197, N2549);
and AND3 (N4209, N4203, N1056, N1546);
nand NAND3 (N4210, N4204, N2497, N3093);
xor XOR2 (N4211, N4191, N3839);
nand NAND2 (N4212, N4199, N2386);
and AND2 (N4213, N4211, N4187);
nor NOR3 (N4214, N4207, N429, N1754);
and AND3 (N4215, N4200, N3004, N1090);
nand NAND2 (N4216, N4210, N1394);
and AND4 (N4217, N4216, N1012, N2757, N2443);
xor XOR2 (N4218, N4184, N973);
nor NOR4 (N4219, N4218, N1677, N3293, N3031);
buf BUF1 (N4220, N4192);
and AND4 (N4221, N4209, N2732, N1246, N479);
and AND4 (N4222, N4214, N3472, N3553, N1024);
and AND4 (N4223, N4215, N1099, N2710, N3353);
nand NAND2 (N4224, N4223, N3450);
xor XOR2 (N4225, N4208, N2810);
nand NAND4 (N4226, N4225, N2601, N3711, N2164);
and AND3 (N4227, N4212, N25, N3271);
or OR2 (N4228, N4222, N275);
and AND4 (N4229, N4217, N2102, N3191, N3353);
and AND2 (N4230, N4220, N4026);
or OR2 (N4231, N4219, N3841);
nand NAND3 (N4232, N4230, N2028, N3070);
or OR2 (N4233, N4231, N1461);
xor XOR2 (N4234, N4224, N3680);
not NOT1 (N4235, N4234);
and AND2 (N4236, N4206, N760);
and AND3 (N4237, N4226, N147, N475);
xor XOR2 (N4238, N4221, N1561);
or OR2 (N4239, N4213, N2026);
nand NAND3 (N4240, N4228, N3457, N1458);
nor NOR2 (N4241, N4240, N357);
or OR2 (N4242, N4237, N1506);
nor NOR2 (N4243, N4242, N3512);
or OR3 (N4244, N4243, N2812, N3679);
or OR4 (N4245, N4236, N1869, N309, N2834);
nor NOR2 (N4246, N4239, N3976);
not NOT1 (N4247, N4235);
xor XOR2 (N4248, N4229, N2319);
or OR2 (N4249, N4247, N550);
not NOT1 (N4250, N4249);
or OR2 (N4251, N4248, N243);
xor XOR2 (N4252, N4246, N3167);
and AND2 (N4253, N4250, N3960);
and AND2 (N4254, N4253, N3276);
and AND3 (N4255, N4251, N2924, N492);
nor NOR2 (N4256, N4252, N3741);
buf BUF1 (N4257, N4238);
nor NOR3 (N4258, N4241, N2042, N3042);
not NOT1 (N4259, N4257);
or OR2 (N4260, N4258, N1611);
nand NAND2 (N4261, N4254, N1358);
buf BUF1 (N4262, N4255);
nor NOR3 (N4263, N4232, N4162, N2077);
nor NOR3 (N4264, N4262, N2461, N1956);
buf BUF1 (N4265, N4259);
or OR4 (N4266, N4245, N1698, N1017, N435);
buf BUF1 (N4267, N4266);
buf BUF1 (N4268, N4227);
nor NOR4 (N4269, N4265, N3107, N537, N1332);
not NOT1 (N4270, N4268);
xor XOR2 (N4271, N4264, N3310);
nand NAND2 (N4272, N4261, N1991);
nand NAND2 (N4273, N4260, N1899);
or OR4 (N4274, N4267, N1664, N2959, N2040);
or OR4 (N4275, N4244, N554, N3907, N2790);
and AND3 (N4276, N4271, N2190, N833);
or OR2 (N4277, N4256, N2384);
xor XOR2 (N4278, N4269, N1907);
buf BUF1 (N4279, N4278);
xor XOR2 (N4280, N4273, N387);
buf BUF1 (N4281, N4279);
nand NAND2 (N4282, N4275, N2296);
or OR2 (N4283, N4282, N911);
or OR4 (N4284, N4280, N2767, N1049, N219);
or OR2 (N4285, N4281, N3589);
and AND3 (N4286, N4284, N729, N2953);
buf BUF1 (N4287, N4233);
nand NAND3 (N4288, N4272, N1628, N2530);
xor XOR2 (N4289, N4263, N4106);
and AND3 (N4290, N4288, N3248, N4132);
and AND4 (N4291, N4274, N1932, N941, N3586);
nand NAND2 (N4292, N4289, N1184);
not NOT1 (N4293, N4286);
not NOT1 (N4294, N4292);
or OR4 (N4295, N4285, N4176, N1916, N57);
and AND3 (N4296, N4293, N784, N2972);
buf BUF1 (N4297, N4283);
and AND2 (N4298, N4277, N4225);
and AND4 (N4299, N4298, N896, N1692, N73);
nor NOR4 (N4300, N4270, N1874, N1569, N2753);
not NOT1 (N4301, N4296);
nand NAND3 (N4302, N4299, N1209, N4012);
not NOT1 (N4303, N4300);
and AND4 (N4304, N4297, N1910, N1567, N1597);
or OR4 (N4305, N4304, N320, N407, N2851);
or OR3 (N4306, N4303, N3380, N3186);
nor NOR3 (N4307, N4301, N2907, N2760);
buf BUF1 (N4308, N4306);
nand NAND3 (N4309, N4291, N2144, N536);
or OR3 (N4310, N4308, N3071, N2394);
buf BUF1 (N4311, N4310);
not NOT1 (N4312, N4276);
or OR4 (N4313, N4290, N2531, N2644, N2463);
nand NAND3 (N4314, N4295, N3110, N1604);
xor XOR2 (N4315, N4302, N1295);
and AND3 (N4316, N4309, N3151, N4256);
buf BUF1 (N4317, N4313);
xor XOR2 (N4318, N4314, N1);
and AND2 (N4319, N4311, N4091);
xor XOR2 (N4320, N4319, N1967);
or OR2 (N4321, N4305, N3679);
xor XOR2 (N4322, N4315, N2398);
not NOT1 (N4323, N4321);
xor XOR2 (N4324, N4287, N3957);
nor NOR2 (N4325, N4322, N2159);
xor XOR2 (N4326, N4320, N2105);
and AND4 (N4327, N4294, N1854, N1132, N1315);
nand NAND3 (N4328, N4317, N837, N3330);
nand NAND4 (N4329, N4316, N3605, N1968, N2843);
xor XOR2 (N4330, N4324, N1527);
or OR2 (N4331, N4328, N2396);
or OR4 (N4332, N4318, N2371, N1172, N938);
buf BUF1 (N4333, N4325);
and AND4 (N4334, N4326, N3782, N322, N3045);
nor NOR2 (N4335, N4329, N4030);
buf BUF1 (N4336, N4334);
xor XOR2 (N4337, N4332, N4091);
xor XOR2 (N4338, N4331, N1977);
or OR4 (N4339, N4338, N944, N3648, N3642);
or OR2 (N4340, N4339, N324);
and AND4 (N4341, N4335, N454, N1257, N2388);
nor NOR4 (N4342, N4337, N517, N984, N83);
and AND2 (N4343, N4333, N840);
nor NOR2 (N4344, N4307, N683);
not NOT1 (N4345, N4327);
and AND3 (N4346, N4342, N3179, N3440);
or OR4 (N4347, N4340, N1050, N3352, N2900);
and AND2 (N4348, N4330, N2794);
and AND4 (N4349, N4341, N164, N1705, N3968);
buf BUF1 (N4350, N4312);
nor NOR2 (N4351, N4345, N3014);
not NOT1 (N4352, N4349);
not NOT1 (N4353, N4336);
not NOT1 (N4354, N4347);
or OR3 (N4355, N4353, N878, N714);
or OR3 (N4356, N4346, N3649, N1766);
buf BUF1 (N4357, N4352);
nand NAND2 (N4358, N4351, N2080);
nand NAND3 (N4359, N4323, N1773, N3985);
and AND2 (N4360, N4344, N988);
and AND4 (N4361, N4343, N4277, N1243, N2092);
not NOT1 (N4362, N4356);
buf BUF1 (N4363, N4362);
not NOT1 (N4364, N4357);
nor NOR2 (N4365, N4348, N507);
nor NOR3 (N4366, N4359, N1114, N1135);
xor XOR2 (N4367, N4364, N3456);
buf BUF1 (N4368, N4354);
and AND2 (N4369, N4350, N2748);
not NOT1 (N4370, N4355);
nor NOR4 (N4371, N4358, N4213, N580, N1584);
and AND3 (N4372, N4361, N2919, N3607);
or OR4 (N4373, N4360, N4213, N4128, N3995);
not NOT1 (N4374, N4371);
or OR3 (N4375, N4366, N70, N2281);
or OR4 (N4376, N4373, N677, N316, N1363);
and AND4 (N4377, N4367, N1107, N575, N3120);
nand NAND3 (N4378, N4365, N2228, N1654);
xor XOR2 (N4379, N4370, N1367);
and AND2 (N4380, N4376, N3661);
xor XOR2 (N4381, N4378, N3692);
xor XOR2 (N4382, N4381, N2055);
nand NAND4 (N4383, N4375, N3626, N3930, N3816);
or OR4 (N4384, N4368, N2429, N1643, N3460);
or OR2 (N4385, N4380, N3847);
buf BUF1 (N4386, N4382);
not NOT1 (N4387, N4383);
nand NAND3 (N4388, N4384, N2388, N742);
buf BUF1 (N4389, N4386);
nand NAND4 (N4390, N4387, N1263, N4262, N255);
or OR4 (N4391, N4363, N788, N2184, N3554);
nor NOR4 (N4392, N4385, N485, N1162, N527);
and AND2 (N4393, N4389, N2837);
and AND2 (N4394, N4391, N2317);
buf BUF1 (N4395, N4374);
xor XOR2 (N4396, N4377, N600);
buf BUF1 (N4397, N4392);
and AND3 (N4398, N4394, N3237, N2633);
or OR3 (N4399, N4397, N2847, N3997);
or OR4 (N4400, N4395, N81, N4044, N3769);
nand NAND2 (N4401, N4399, N2054);
or OR3 (N4402, N4390, N1840, N2137);
not NOT1 (N4403, N4396);
not NOT1 (N4404, N4388);
nor NOR3 (N4405, N4369, N1406, N1741);
or OR2 (N4406, N4400, N3187);
buf BUF1 (N4407, N4379);
and AND2 (N4408, N4372, N1976);
nor NOR2 (N4409, N4406, N301);
and AND3 (N4410, N4393, N1610, N898);
and AND4 (N4411, N4410, N2474, N1658, N3196);
or OR3 (N4412, N4407, N928, N757);
not NOT1 (N4413, N4404);
nand NAND2 (N4414, N4412, N1966);
not NOT1 (N4415, N4413);
xor XOR2 (N4416, N4403, N1830);
nor NOR3 (N4417, N4409, N3080, N2802);
buf BUF1 (N4418, N4411);
nand NAND2 (N4419, N4418, N879);
nor NOR2 (N4420, N4402, N3196);
buf BUF1 (N4421, N4405);
nor NOR4 (N4422, N4421, N2385, N3576, N4206);
xor XOR2 (N4423, N4408, N2229);
and AND3 (N4424, N4398, N551, N2438);
buf BUF1 (N4425, N4422);
not NOT1 (N4426, N4416);
and AND4 (N4427, N4425, N4054, N2982, N407);
or OR3 (N4428, N4419, N4332, N1125);
buf BUF1 (N4429, N4417);
and AND4 (N4430, N4415, N2934, N459, N3287);
and AND2 (N4431, N4414, N2437);
xor XOR2 (N4432, N4420, N1745);
not NOT1 (N4433, N4427);
and AND2 (N4434, N4424, N4413);
or OR4 (N4435, N4401, N2716, N2869, N3824);
and AND3 (N4436, N4435, N875, N4014);
nor NOR4 (N4437, N4436, N2963, N2617, N4043);
not NOT1 (N4438, N4423);
xor XOR2 (N4439, N4431, N3226);
or OR2 (N4440, N4429, N2674);
xor XOR2 (N4441, N4428, N3598);
nand NAND2 (N4442, N4438, N1524);
buf BUF1 (N4443, N4434);
and AND3 (N4444, N4441, N914, N534);
not NOT1 (N4445, N4440);
and AND2 (N4446, N4443, N2168);
nor NOR3 (N4447, N4426, N3566, N2698);
or OR4 (N4448, N4447, N2391, N1408, N729);
not NOT1 (N4449, N4442);
or OR4 (N4450, N4430, N2071, N540, N626);
buf BUF1 (N4451, N4433);
buf BUF1 (N4452, N4439);
or OR3 (N4453, N4432, N681, N2431);
xor XOR2 (N4454, N4445, N3590);
not NOT1 (N4455, N4452);
not NOT1 (N4456, N4448);
xor XOR2 (N4457, N4444, N1667);
or OR4 (N4458, N4437, N3164, N2150, N3989);
xor XOR2 (N4459, N4454, N3579);
or OR3 (N4460, N4458, N1881, N433);
nor NOR3 (N4461, N4453, N2833, N4443);
xor XOR2 (N4462, N4450, N3963);
and AND4 (N4463, N4455, N2043, N3458, N3315);
or OR3 (N4464, N4451, N4151, N3296);
or OR3 (N4465, N4462, N724, N1028);
and AND2 (N4466, N4446, N533);
and AND3 (N4467, N4459, N1346, N4109);
not NOT1 (N4468, N4465);
nand NAND4 (N4469, N4466, N34, N1763, N2169);
xor XOR2 (N4470, N4460, N2116);
and AND4 (N4471, N4469, N2092, N307, N2177);
nand NAND2 (N4472, N4471, N2216);
or OR3 (N4473, N4461, N2697, N296);
or OR3 (N4474, N4467, N955, N4191);
nor NOR2 (N4475, N4470, N4417);
xor XOR2 (N4476, N4464, N1812);
or OR2 (N4477, N4463, N4390);
buf BUF1 (N4478, N4472);
nor NOR2 (N4479, N4475, N1129);
nand NAND4 (N4480, N4476, N1162, N2156, N510);
xor XOR2 (N4481, N4474, N3649);
not NOT1 (N4482, N4477);
or OR3 (N4483, N4456, N162, N2765);
nor NOR4 (N4484, N4473, N2100, N2077, N2696);
not NOT1 (N4485, N4468);
not NOT1 (N4486, N4478);
and AND2 (N4487, N4449, N4072);
not NOT1 (N4488, N4485);
xor XOR2 (N4489, N4488, N831);
nor NOR4 (N4490, N4484, N1787, N870, N405);
not NOT1 (N4491, N4486);
and AND2 (N4492, N4480, N2159);
xor XOR2 (N4493, N4479, N1309);
xor XOR2 (N4494, N4492, N1676);
xor XOR2 (N4495, N4481, N2643);
and AND2 (N4496, N4483, N1578);
xor XOR2 (N4497, N4495, N3309);
xor XOR2 (N4498, N4496, N1538);
xor XOR2 (N4499, N4482, N3325);
and AND3 (N4500, N4489, N904, N2402);
nor NOR3 (N4501, N4487, N1723, N1343);
and AND4 (N4502, N4500, N3925, N2405, N62);
or OR4 (N4503, N4498, N2386, N3220, N4492);
nand NAND3 (N4504, N4499, N3790, N791);
buf BUF1 (N4505, N4501);
or OR4 (N4506, N4502, N3088, N2706, N3487);
nor NOR3 (N4507, N4457, N377, N3324);
nor NOR2 (N4508, N4497, N1514);
and AND3 (N4509, N4493, N1580, N1975);
nor NOR2 (N4510, N4505, N3209);
or OR3 (N4511, N4508, N2975, N3153);
not NOT1 (N4512, N4511);
buf BUF1 (N4513, N4494);
buf BUF1 (N4514, N4491);
nor NOR3 (N4515, N4513, N3386, N348);
buf BUF1 (N4516, N4515);
and AND3 (N4517, N4490, N3435, N452);
buf BUF1 (N4518, N4516);
buf BUF1 (N4519, N4509);
xor XOR2 (N4520, N4514, N2506);
nand NAND3 (N4521, N4503, N1012, N1834);
and AND2 (N4522, N4506, N3547);
buf BUF1 (N4523, N4518);
buf BUF1 (N4524, N4510);
buf BUF1 (N4525, N4523);
not NOT1 (N4526, N4507);
nor NOR2 (N4527, N4524, N3131);
not NOT1 (N4528, N4526);
nand NAND3 (N4529, N4528, N687, N2642);
not NOT1 (N4530, N4521);
not NOT1 (N4531, N4520);
not NOT1 (N4532, N4517);
buf BUF1 (N4533, N4532);
xor XOR2 (N4534, N4512, N4067);
nor NOR3 (N4535, N4504, N376, N2827);
xor XOR2 (N4536, N4535, N1949);
nand NAND3 (N4537, N4536, N810, N1248);
buf BUF1 (N4538, N4537);
and AND4 (N4539, N4530, N2845, N1931, N2167);
or OR2 (N4540, N4539, N3280);
and AND4 (N4541, N4527, N132, N501, N2590);
buf BUF1 (N4542, N4533);
or OR2 (N4543, N4540, N4036);
not NOT1 (N4544, N4538);
buf BUF1 (N4545, N4543);
buf BUF1 (N4546, N4534);
buf BUF1 (N4547, N4531);
not NOT1 (N4548, N4546);
nor NOR2 (N4549, N4544, N3248);
or OR3 (N4550, N4547, N4510, N1863);
nor NOR2 (N4551, N4522, N4197);
xor XOR2 (N4552, N4548, N1550);
and AND2 (N4553, N4529, N1008);
or OR4 (N4554, N4553, N1339, N1753, N552);
xor XOR2 (N4555, N4541, N3167);
and AND2 (N4556, N4525, N2422);
buf BUF1 (N4557, N4551);
and AND4 (N4558, N4552, N1436, N3328, N59);
not NOT1 (N4559, N4550);
nor NOR3 (N4560, N4545, N2503, N3987);
buf BUF1 (N4561, N4560);
nand NAND3 (N4562, N4561, N1220, N1364);
nand NAND2 (N4563, N4555, N2176);
nand NAND2 (N4564, N4556, N4351);
or OR4 (N4565, N4519, N1601, N4470, N1208);
nand NAND2 (N4566, N4554, N1422);
not NOT1 (N4567, N4563);
nand NAND2 (N4568, N4565, N1469);
xor XOR2 (N4569, N4559, N4180);
and AND4 (N4570, N4542, N1730, N1686, N552);
nand NAND2 (N4571, N4557, N2633);
buf BUF1 (N4572, N4564);
and AND3 (N4573, N4558, N2365, N1699);
xor XOR2 (N4574, N4566, N1187);
and AND3 (N4575, N4568, N118, N3902);
nand NAND4 (N4576, N4549, N1011, N3382, N1647);
nand NAND4 (N4577, N4575, N4386, N2501, N2535);
buf BUF1 (N4578, N4567);
nand NAND3 (N4579, N4578, N4540, N385);
xor XOR2 (N4580, N4573, N2468);
not NOT1 (N4581, N4570);
and AND4 (N4582, N4574, N3086, N387, N2438);
buf BUF1 (N4583, N4572);
nor NOR4 (N4584, N4562, N777, N2790, N2605);
and AND2 (N4585, N4571, N3793);
nand NAND4 (N4586, N4577, N4052, N4463, N2284);
buf BUF1 (N4587, N4579);
not NOT1 (N4588, N4587);
xor XOR2 (N4589, N4580, N1641);
and AND4 (N4590, N4583, N3801, N2506, N2932);
nor NOR2 (N4591, N4590, N3521);
buf BUF1 (N4592, N4582);
nand NAND3 (N4593, N4569, N241, N3172);
and AND4 (N4594, N4589, N1324, N3758, N1103);
nor NOR2 (N4595, N4584, N1338);
and AND3 (N4596, N4591, N3519, N2439);
and AND3 (N4597, N4594, N1031, N1416);
xor XOR2 (N4598, N4576, N1467);
or OR3 (N4599, N4597, N2701, N3182);
not NOT1 (N4600, N4599);
and AND2 (N4601, N4588, N3394);
not NOT1 (N4602, N4595);
not NOT1 (N4603, N4592);
nor NOR4 (N4604, N4586, N2701, N3953, N3028);
xor XOR2 (N4605, N4600, N667);
buf BUF1 (N4606, N4596);
not NOT1 (N4607, N4606);
not NOT1 (N4608, N4585);
and AND4 (N4609, N4607, N202, N4165, N3748);
nand NAND3 (N4610, N4593, N3121, N1586);
not NOT1 (N4611, N4610);
or OR2 (N4612, N4603, N4118);
and AND4 (N4613, N4608, N2351, N4425, N4187);
not NOT1 (N4614, N4609);
buf BUF1 (N4615, N4598);
nor NOR3 (N4616, N4581, N4219, N4000);
nor NOR2 (N4617, N4614, N558);
buf BUF1 (N4618, N4605);
buf BUF1 (N4619, N4601);
or OR4 (N4620, N4604, N4482, N1089, N1108);
buf BUF1 (N4621, N4612);
buf BUF1 (N4622, N4619);
nand NAND3 (N4623, N4615, N7, N2605);
not NOT1 (N4624, N4617);
xor XOR2 (N4625, N4623, N2951);
xor XOR2 (N4626, N4622, N4475);
nor NOR3 (N4627, N4625, N2775, N1751);
and AND2 (N4628, N4616, N3090);
buf BUF1 (N4629, N4618);
nand NAND3 (N4630, N4611, N163, N2047);
and AND4 (N4631, N4626, N3038, N890, N2602);
xor XOR2 (N4632, N4602, N3023);
nand NAND2 (N4633, N4627, N3944);
buf BUF1 (N4634, N4632);
xor XOR2 (N4635, N4613, N866);
nor NOR4 (N4636, N4631, N2548, N79, N2612);
nor NOR4 (N4637, N4628, N900, N2034, N4154);
nand NAND4 (N4638, N4637, N1406, N2194, N428);
nor NOR3 (N4639, N4620, N2004, N1241);
nand NAND3 (N4640, N4621, N1413, N3759);
buf BUF1 (N4641, N4640);
xor XOR2 (N4642, N4629, N792);
not NOT1 (N4643, N4624);
nand NAND4 (N4644, N4643, N197, N1301, N3562);
nand NAND3 (N4645, N4644, N2802, N2975);
and AND3 (N4646, N4638, N309, N2135);
and AND4 (N4647, N4634, N1521, N1856, N585);
nand NAND4 (N4648, N4645, N373, N3865, N1895);
nor NOR4 (N4649, N4648, N2899, N2877, N4273);
not NOT1 (N4650, N4641);
buf BUF1 (N4651, N4649);
not NOT1 (N4652, N4650);
nand NAND4 (N4653, N4630, N88, N4161, N1707);
and AND2 (N4654, N4647, N3760);
buf BUF1 (N4655, N4636);
nor NOR3 (N4656, N4642, N1612, N4166);
nand NAND3 (N4657, N4654, N988, N3662);
buf BUF1 (N4658, N4633);
buf BUF1 (N4659, N4656);
buf BUF1 (N4660, N4635);
xor XOR2 (N4661, N4653, N1724);
and AND2 (N4662, N4646, N2419);
and AND4 (N4663, N4655, N4310, N3539, N4050);
nor NOR3 (N4664, N4660, N4102, N3888);
nand NAND3 (N4665, N4661, N1071, N1402);
xor XOR2 (N4666, N4639, N4378);
and AND2 (N4667, N4659, N298);
xor XOR2 (N4668, N4651, N3307);
buf BUF1 (N4669, N4658);
or OR2 (N4670, N4668, N2598);
or OR2 (N4671, N4662, N3836);
nor NOR4 (N4672, N4671, N3939, N637, N4441);
buf BUF1 (N4673, N4672);
and AND3 (N4674, N4673, N3717, N1230);
nor NOR4 (N4675, N4667, N1560, N694, N1641);
and AND4 (N4676, N4670, N219, N1724, N3411);
nor NOR4 (N4677, N4669, N1323, N3504, N1501);
nand NAND4 (N4678, N4657, N2597, N2418, N2625);
and AND2 (N4679, N4676, N3170);
not NOT1 (N4680, N4679);
not NOT1 (N4681, N4665);
nor NOR4 (N4682, N4680, N582, N968, N1789);
xor XOR2 (N4683, N4652, N755);
buf BUF1 (N4684, N4666);
buf BUF1 (N4685, N4678);
nor NOR2 (N4686, N4682, N1936);
nor NOR4 (N4687, N4685, N2906, N1718, N7);
nand NAND3 (N4688, N4686, N2121, N171);
nand NAND3 (N4689, N4683, N507, N518);
nand NAND2 (N4690, N4687, N3159);
xor XOR2 (N4691, N4674, N3816);
xor XOR2 (N4692, N4689, N963);
nor NOR2 (N4693, N4681, N2108);
not NOT1 (N4694, N4675);
xor XOR2 (N4695, N4692, N1195);
and AND3 (N4696, N4664, N4240, N135);
nor NOR3 (N4697, N4693, N590, N84);
not NOT1 (N4698, N4691);
not NOT1 (N4699, N4684);
nor NOR4 (N4700, N4695, N1454, N546, N1267);
or OR3 (N4701, N4697, N2686, N3754);
nor NOR4 (N4702, N4701, N1613, N2473, N2801);
nand NAND4 (N4703, N4663, N1419, N876, N2216);
buf BUF1 (N4704, N4688);
nor NOR4 (N4705, N4703, N1664, N3494, N2854);
nor NOR4 (N4706, N4696, N3658, N1724, N515);
xor XOR2 (N4707, N4699, N225);
buf BUF1 (N4708, N4704);
nand NAND3 (N4709, N4698, N4510, N3748);
and AND3 (N4710, N4708, N141, N2112);
xor XOR2 (N4711, N4700, N1267);
nor NOR4 (N4712, N4677, N2494, N4225, N46);
xor XOR2 (N4713, N4707, N4078);
buf BUF1 (N4714, N4711);
buf BUF1 (N4715, N4690);
buf BUF1 (N4716, N4712);
nor NOR4 (N4717, N4716, N2163, N825, N1487);
nand NAND3 (N4718, N4710, N2272, N2336);
not NOT1 (N4719, N4702);
xor XOR2 (N4720, N4715, N4511);
or OR3 (N4721, N4709, N3558, N4545);
not NOT1 (N4722, N4706);
not NOT1 (N4723, N4717);
and AND2 (N4724, N4694, N4487);
nor NOR2 (N4725, N4705, N3094);
or OR4 (N4726, N4725, N143, N1819, N3209);
not NOT1 (N4727, N4721);
nor NOR3 (N4728, N4718, N773, N3031);
buf BUF1 (N4729, N4714);
nand NAND3 (N4730, N4722, N3110, N623);
not NOT1 (N4731, N4720);
nor NOR4 (N4732, N4731, N664, N2920, N3717);
and AND4 (N4733, N4719, N2451, N4687, N1519);
or OR4 (N4734, N4733, N1652, N1704, N3589);
or OR2 (N4735, N4734, N3952);
nor NOR4 (N4736, N4728, N1221, N4105, N241);
buf BUF1 (N4737, N4726);
not NOT1 (N4738, N4737);
not NOT1 (N4739, N4713);
nand NAND4 (N4740, N4729, N4491, N4187, N4548);
and AND3 (N4741, N4730, N3739, N2464);
buf BUF1 (N4742, N4727);
buf BUF1 (N4743, N4724);
buf BUF1 (N4744, N4741);
or OR4 (N4745, N4740, N2329, N3756, N3857);
not NOT1 (N4746, N4742);
not NOT1 (N4747, N4744);
nand NAND2 (N4748, N4723, N2780);
xor XOR2 (N4749, N4739, N1817);
and AND4 (N4750, N4743, N4472, N406, N731);
and AND4 (N4751, N4748, N1744, N1994, N163);
not NOT1 (N4752, N4732);
buf BUF1 (N4753, N4746);
not NOT1 (N4754, N4745);
xor XOR2 (N4755, N4736, N1298);
not NOT1 (N4756, N4752);
nand NAND3 (N4757, N4755, N1322, N2197);
nand NAND4 (N4758, N4747, N3295, N1190, N4542);
nor NOR4 (N4759, N4749, N3483, N688, N3214);
and AND3 (N4760, N4753, N39, N2987);
and AND4 (N4761, N4756, N1273, N4666, N4155);
and AND3 (N4762, N4760, N1511, N3298);
nor NOR2 (N4763, N4735, N2516);
xor XOR2 (N4764, N4738, N1763);
and AND3 (N4765, N4754, N2636, N3630);
not NOT1 (N4766, N4762);
nor NOR2 (N4767, N4763, N1124);
and AND3 (N4768, N4757, N55, N2042);
or OR4 (N4769, N4761, N2365, N1886, N3134);
nor NOR2 (N4770, N4768, N2555);
buf BUF1 (N4771, N4769);
xor XOR2 (N4772, N4770, N3445);
not NOT1 (N4773, N4765);
nand NAND2 (N4774, N4766, N3502);
and AND4 (N4775, N4751, N3090, N2156, N3964);
nor NOR4 (N4776, N4759, N2071, N1240, N531);
not NOT1 (N4777, N4776);
or OR4 (N4778, N4775, N2095, N4661, N420);
nand NAND4 (N4779, N4773, N598, N1545, N2977);
buf BUF1 (N4780, N4767);
buf BUF1 (N4781, N4774);
nand NAND2 (N4782, N4772, N653);
buf BUF1 (N4783, N4781);
not NOT1 (N4784, N4783);
and AND3 (N4785, N4784, N4293, N4774);
nand NAND3 (N4786, N4782, N3590, N1143);
buf BUF1 (N4787, N4779);
xor XOR2 (N4788, N4778, N2595);
xor XOR2 (N4789, N4764, N1544);
not NOT1 (N4790, N4785);
xor XOR2 (N4791, N4758, N1085);
or OR3 (N4792, N4777, N4599, N3967);
and AND2 (N4793, N4787, N983);
or OR2 (N4794, N4771, N118);
xor XOR2 (N4795, N4792, N2071);
nand NAND2 (N4796, N4788, N4694);
not NOT1 (N4797, N4796);
buf BUF1 (N4798, N4791);
and AND3 (N4799, N4780, N2742, N4134);
nor NOR3 (N4800, N4789, N2547, N3815);
nand NAND4 (N4801, N4798, N1605, N4658, N4202);
nand NAND3 (N4802, N4793, N1570, N533);
buf BUF1 (N4803, N4797);
buf BUF1 (N4804, N4803);
buf BUF1 (N4805, N4799);
or OR2 (N4806, N4794, N3736);
buf BUF1 (N4807, N4806);
nor NOR4 (N4808, N4786, N2038, N1797, N3152);
nand NAND4 (N4809, N4750, N1362, N394, N4117);
buf BUF1 (N4810, N4801);
or OR2 (N4811, N4802, N144);
buf BUF1 (N4812, N4805);
and AND4 (N4813, N4804, N2362, N3969, N260);
and AND3 (N4814, N4812, N2477, N3023);
not NOT1 (N4815, N4813);
not NOT1 (N4816, N4810);
buf BUF1 (N4817, N4795);
nor NOR4 (N4818, N4807, N2215, N1624, N4816);
nor NOR4 (N4819, N700, N3880, N4585, N743);
buf BUF1 (N4820, N4817);
or OR4 (N4821, N4820, N1137, N2786, N3236);
nor NOR4 (N4822, N4808, N771, N3870, N3591);
buf BUF1 (N4823, N4811);
and AND4 (N4824, N4818, N965, N2779, N3539);
nand NAND2 (N4825, N4819, N3966);
nor NOR4 (N4826, N4790, N566, N2361, N1348);
nand NAND4 (N4827, N4821, N4400, N3258, N4059);
xor XOR2 (N4828, N4815, N4044);
xor XOR2 (N4829, N4814, N4631);
and AND3 (N4830, N4827, N4493, N1578);
and AND4 (N4831, N4809, N4136, N792, N1311);
nor NOR3 (N4832, N4826, N621, N1152);
nand NAND3 (N4833, N4830, N1898, N3694);
and AND4 (N4834, N4824, N460, N3881, N4117);
and AND3 (N4835, N4825, N3868, N1551);
xor XOR2 (N4836, N4800, N3967);
buf BUF1 (N4837, N4829);
or OR2 (N4838, N4835, N2655);
nor NOR4 (N4839, N4822, N517, N1612, N612);
not NOT1 (N4840, N4839);
not NOT1 (N4841, N4838);
not NOT1 (N4842, N4832);
xor XOR2 (N4843, N4823, N3593);
not NOT1 (N4844, N4842);
buf BUF1 (N4845, N4844);
nor NOR2 (N4846, N4843, N2951);
nor NOR3 (N4847, N4840, N2546, N4425);
nor NOR3 (N4848, N4841, N2103, N3664);
and AND3 (N4849, N4828, N4292, N266);
or OR3 (N4850, N4833, N3965, N1312);
nor NOR2 (N4851, N4850, N812);
and AND4 (N4852, N4836, N1057, N4677, N2595);
buf BUF1 (N4853, N4847);
nand NAND3 (N4854, N4831, N1791, N1537);
buf BUF1 (N4855, N4851);
not NOT1 (N4856, N4848);
or OR2 (N4857, N4834, N3574);
nor NOR3 (N4858, N4857, N2360, N4314);
and AND3 (N4859, N4854, N4065, N1953);
nor NOR4 (N4860, N4846, N4435, N1408, N4028);
or OR4 (N4861, N4845, N3421, N3208, N782);
nor NOR2 (N4862, N4856, N3197);
or OR2 (N4863, N4837, N4447);
and AND4 (N4864, N4852, N3947, N499, N4588);
nand NAND3 (N4865, N4855, N1391, N4700);
nor NOR3 (N4866, N4849, N813, N2099);
or OR2 (N4867, N4862, N3898);
nor NOR3 (N4868, N4861, N2400, N1723);
nand NAND3 (N4869, N4859, N1438, N563);
nand NAND2 (N4870, N4860, N2732);
and AND4 (N4871, N4853, N2365, N3172, N3598);
nand NAND3 (N4872, N4864, N4444, N3279);
nand NAND3 (N4873, N4871, N4233, N777);
and AND4 (N4874, N4867, N2541, N2956, N1690);
buf BUF1 (N4875, N4858);
buf BUF1 (N4876, N4863);
nand NAND2 (N4877, N4870, N1270);
nand NAND3 (N4878, N4875, N1571, N69);
xor XOR2 (N4879, N4869, N3199);
xor XOR2 (N4880, N4879, N2353);
and AND2 (N4881, N4876, N1178);
or OR2 (N4882, N4880, N2861);
xor XOR2 (N4883, N4873, N2623);
nor NOR4 (N4884, N4872, N252, N2534, N4664);
buf BUF1 (N4885, N4866);
xor XOR2 (N4886, N4883, N1669);
or OR4 (N4887, N4881, N3362, N653, N2146);
or OR3 (N4888, N4887, N284, N4311);
or OR4 (N4889, N4888, N853, N2357, N3451);
nor NOR2 (N4890, N4886, N1488);
and AND2 (N4891, N4865, N2229);
or OR3 (N4892, N4889, N4748, N4265);
and AND4 (N4893, N4892, N4127, N1115, N3869);
nor NOR4 (N4894, N4893, N4083, N558, N4016);
or OR3 (N4895, N4874, N2438, N4818);
nand NAND4 (N4896, N4890, N1432, N1343, N2634);
not NOT1 (N4897, N4868);
xor XOR2 (N4898, N4894, N377);
buf BUF1 (N4899, N4878);
nor NOR3 (N4900, N4895, N3116, N4848);
buf BUF1 (N4901, N4891);
buf BUF1 (N4902, N4885);
or OR4 (N4903, N4901, N4393, N1373, N3395);
not NOT1 (N4904, N4902);
not NOT1 (N4905, N4900);
nand NAND2 (N4906, N4904, N4536);
or OR2 (N4907, N4906, N2373);
and AND3 (N4908, N4896, N2607, N1113);
or OR3 (N4909, N4907, N2929, N3629);
xor XOR2 (N4910, N4905, N938);
nor NOR4 (N4911, N4908, N807, N3036, N3366);
xor XOR2 (N4912, N4911, N3197);
not NOT1 (N4913, N4877);
not NOT1 (N4914, N4898);
buf BUF1 (N4915, N4912);
xor XOR2 (N4916, N4910, N229);
nand NAND3 (N4917, N4915, N752, N3318);
nand NAND3 (N4918, N4903, N916, N114);
buf BUF1 (N4919, N4914);
not NOT1 (N4920, N4882);
not NOT1 (N4921, N4909);
or OR4 (N4922, N4884, N4370, N874, N4417);
or OR2 (N4923, N4922, N4413);
buf BUF1 (N4924, N4919);
nor NOR3 (N4925, N4918, N1571, N2230);
and AND4 (N4926, N4923, N568, N3696, N279);
nor NOR2 (N4927, N4897, N874);
not NOT1 (N4928, N4913);
not NOT1 (N4929, N4917);
buf BUF1 (N4930, N4916);
or OR3 (N4931, N4899, N2057, N4189);
not NOT1 (N4932, N4928);
and AND4 (N4933, N4925, N2256, N1572, N4015);
nor NOR3 (N4934, N4927, N2579, N4630);
and AND2 (N4935, N4931, N802);
or OR4 (N4936, N4926, N3912, N1903, N2);
and AND2 (N4937, N4920, N934);
and AND4 (N4938, N4929, N63, N3228, N61);
or OR2 (N4939, N4930, N3163);
not NOT1 (N4940, N4937);
nor NOR2 (N4941, N4938, N3045);
or OR4 (N4942, N4934, N2247, N2841, N3274);
not NOT1 (N4943, N4932);
or OR2 (N4944, N4936, N1752);
nor NOR4 (N4945, N4933, N2794, N794, N4552);
or OR4 (N4946, N4935, N141, N1670, N221);
or OR3 (N4947, N4924, N2266, N2497);
or OR3 (N4948, N4942, N2507, N4236);
xor XOR2 (N4949, N4948, N4612);
or OR3 (N4950, N4946, N2416, N205);
xor XOR2 (N4951, N4947, N838);
or OR2 (N4952, N4940, N2790);
nor NOR3 (N4953, N4949, N1807, N3046);
nand NAND4 (N4954, N4951, N3483, N4265, N2171);
nand NAND2 (N4955, N4943, N3839);
nor NOR4 (N4956, N4939, N2978, N3799, N1310);
xor XOR2 (N4957, N4952, N4898);
and AND2 (N4958, N4950, N2214);
not NOT1 (N4959, N4953);
not NOT1 (N4960, N4957);
buf BUF1 (N4961, N4956);
nand NAND3 (N4962, N4960, N2318, N4617);
nand NAND3 (N4963, N4945, N707, N680);
nand NAND3 (N4964, N4958, N1599, N4397);
and AND3 (N4965, N4944, N4077, N2569);
nand NAND3 (N4966, N4964, N4345, N135);
or OR4 (N4967, N4966, N3772, N1321, N3819);
and AND3 (N4968, N4954, N3036, N2246);
buf BUF1 (N4969, N4963);
nand NAND4 (N4970, N4959, N3479, N182, N3149);
buf BUF1 (N4971, N4962);
nand NAND2 (N4972, N4968, N3910);
nand NAND3 (N4973, N4941, N4036, N2110);
xor XOR2 (N4974, N4973, N2439);
nand NAND3 (N4975, N4921, N4110, N56);
not NOT1 (N4976, N4974);
nand NAND2 (N4977, N4965, N1518);
xor XOR2 (N4978, N4969, N484);
or OR4 (N4979, N4961, N2169, N1679, N1932);
buf BUF1 (N4980, N4975);
not NOT1 (N4981, N4978);
not NOT1 (N4982, N4979);
and AND3 (N4983, N4976, N372, N1384);
and AND4 (N4984, N4955, N3431, N1320, N3620);
and AND3 (N4985, N4970, N661, N4184);
xor XOR2 (N4986, N4977, N180);
buf BUF1 (N4987, N4983);
nand NAND2 (N4988, N4981, N1943);
and AND2 (N4989, N4971, N1680);
buf BUF1 (N4990, N4984);
or OR3 (N4991, N4967, N2675, N998);
nand NAND2 (N4992, N4987, N3263);
nor NOR4 (N4993, N4986, N557, N1820, N1899);
nand NAND4 (N4994, N4990, N2707, N1575, N2710);
nor NOR3 (N4995, N4985, N4850, N3405);
or OR4 (N4996, N4991, N4233, N2725, N4342);
xor XOR2 (N4997, N4972, N1826);
buf BUF1 (N4998, N4988);
xor XOR2 (N4999, N4992, N4675);
buf BUF1 (N5000, N4980);
or OR2 (N5001, N5000, N4002);
nor NOR4 (N5002, N4994, N3663, N1619, N4702);
nand NAND4 (N5003, N5002, N3740, N1412, N2030);
or OR3 (N5004, N5003, N1108, N3352);
and AND2 (N5005, N4982, N1588);
and AND2 (N5006, N4995, N4016);
and AND3 (N5007, N4996, N143, N3844);
not NOT1 (N5008, N5004);
and AND4 (N5009, N5005, N3469, N4975, N1801);
buf BUF1 (N5010, N5009);
not NOT1 (N5011, N5008);
buf BUF1 (N5012, N4997);
and AND4 (N5013, N5001, N3920, N1923, N2273);
and AND3 (N5014, N4998, N3003, N1402);
nand NAND2 (N5015, N4989, N3035);
xor XOR2 (N5016, N4993, N450);
and AND4 (N5017, N5006, N1062, N53, N2012);
xor XOR2 (N5018, N5013, N2823);
nand NAND4 (N5019, N4999, N4211, N1097, N1009);
buf BUF1 (N5020, N5015);
nand NAND3 (N5021, N5007, N2227, N2423);
nor NOR4 (N5022, N5021, N903, N4376, N4930);
buf BUF1 (N5023, N5014);
buf BUF1 (N5024, N5022);
and AND3 (N5025, N5020, N4617, N757);
xor XOR2 (N5026, N5023, N2126);
or OR2 (N5027, N5025, N946);
not NOT1 (N5028, N5012);
xor XOR2 (N5029, N5026, N864);
xor XOR2 (N5030, N5018, N551);
buf BUF1 (N5031, N5030);
or OR4 (N5032, N5010, N1037, N3085, N2130);
xor XOR2 (N5033, N5024, N140);
and AND3 (N5034, N5031, N3584, N1679);
or OR4 (N5035, N5016, N2882, N4442, N4979);
and AND4 (N5036, N5019, N2747, N2734, N4717);
nor NOR3 (N5037, N5033, N1589, N3771);
buf BUF1 (N5038, N5017);
xor XOR2 (N5039, N5036, N888);
and AND3 (N5040, N5035, N3792, N2811);
or OR2 (N5041, N5037, N4561);
buf BUF1 (N5042, N5032);
xor XOR2 (N5043, N5034, N4357);
xor XOR2 (N5044, N5039, N2413);
and AND2 (N5045, N5011, N4846);
nand NAND4 (N5046, N5040, N1235, N2015, N2084);
nand NAND4 (N5047, N5028, N4350, N2065, N3259);
buf BUF1 (N5048, N5042);
buf BUF1 (N5049, N5043);
or OR4 (N5050, N5047, N25, N5024, N4971);
or OR3 (N5051, N5045, N614, N4727);
or OR2 (N5052, N5049, N3984);
buf BUF1 (N5053, N5048);
xor XOR2 (N5054, N5052, N2276);
not NOT1 (N5055, N5027);
nor NOR3 (N5056, N5029, N4752, N2337);
nor NOR2 (N5057, N5053, N4755);
nand NAND4 (N5058, N5056, N4650, N3266, N654);
and AND3 (N5059, N5041, N3546, N3685);
xor XOR2 (N5060, N5057, N4702);
xor XOR2 (N5061, N5051, N4118);
and AND4 (N5062, N5044, N3395, N3855, N3521);
buf BUF1 (N5063, N5062);
and AND2 (N5064, N5058, N4391);
nor NOR4 (N5065, N5063, N2980, N459, N1584);
nor NOR2 (N5066, N5060, N1732);
or OR4 (N5067, N5054, N1254, N3767, N4383);
xor XOR2 (N5068, N5065, N1786);
or OR4 (N5069, N5067, N1986, N127, N4074);
xor XOR2 (N5070, N5055, N4159);
nor NOR2 (N5071, N5068, N1064);
not NOT1 (N5072, N5066);
nor NOR3 (N5073, N5046, N4291, N304);
buf BUF1 (N5074, N5072);
nor NOR2 (N5075, N5050, N2406);
nor NOR2 (N5076, N5074, N4138);
buf BUF1 (N5077, N5070);
buf BUF1 (N5078, N5064);
buf BUF1 (N5079, N5078);
nor NOR4 (N5080, N5075, N3492, N2470, N3424);
nand NAND4 (N5081, N5077, N4906, N1583, N417);
or OR4 (N5082, N5080, N3145, N1167, N1181);
buf BUF1 (N5083, N5071);
buf BUF1 (N5084, N5076);
nor NOR4 (N5085, N5069, N170, N998, N4379);
not NOT1 (N5086, N5085);
and AND4 (N5087, N5084, N4219, N1129, N4093);
nand NAND2 (N5088, N5086, N526);
nand NAND4 (N5089, N5038, N4454, N5054, N4017);
not NOT1 (N5090, N5082);
xor XOR2 (N5091, N5089, N4684);
buf BUF1 (N5092, N5088);
buf BUF1 (N5093, N5092);
xor XOR2 (N5094, N5079, N387);
or OR3 (N5095, N5061, N3778, N838);
nand NAND3 (N5096, N5087, N1834, N1462);
nand NAND4 (N5097, N5090, N375, N1614, N2836);
buf BUF1 (N5098, N5095);
xor XOR2 (N5099, N5091, N2502);
nand NAND3 (N5100, N5096, N4605, N2565);
nor NOR3 (N5101, N5093, N2456, N4230);
not NOT1 (N5102, N5097);
nor NOR4 (N5103, N5100, N4301, N676, N3365);
nor NOR4 (N5104, N5098, N4830, N2999, N4520);
xor XOR2 (N5105, N5073, N4144);
or OR4 (N5106, N5083, N705, N3636, N2092);
not NOT1 (N5107, N5081);
and AND3 (N5108, N5106, N1328, N3942);
nor NOR4 (N5109, N5107, N2012, N4006, N2370);
xor XOR2 (N5110, N5108, N2761);
buf BUF1 (N5111, N5103);
not NOT1 (N5112, N5059);
or OR4 (N5113, N5101, N3556, N2462, N2280);
nand NAND3 (N5114, N5099, N4641, N2106);
buf BUF1 (N5115, N5113);
not NOT1 (N5116, N5094);
nor NOR3 (N5117, N5105, N1047, N2323);
nand NAND4 (N5118, N5111, N2487, N4306, N2956);
xor XOR2 (N5119, N5104, N4828);
not NOT1 (N5120, N5118);
not NOT1 (N5121, N5102);
nor NOR2 (N5122, N5109, N5090);
not NOT1 (N5123, N5112);
not NOT1 (N5124, N5110);
buf BUF1 (N5125, N5119);
nand NAND3 (N5126, N5122, N1702, N1834);
buf BUF1 (N5127, N5121);
and AND2 (N5128, N5116, N3860);
buf BUF1 (N5129, N5124);
nand NAND3 (N5130, N5129, N3242, N3859);
buf BUF1 (N5131, N5120);
and AND4 (N5132, N5123, N4710, N2678, N1048);
nor NOR3 (N5133, N5131, N406, N3230);
not NOT1 (N5134, N5128);
buf BUF1 (N5135, N5132);
nand NAND4 (N5136, N5130, N5068, N4563, N3354);
or OR2 (N5137, N5114, N1062);
nand NAND3 (N5138, N5135, N3102, N175);
and AND3 (N5139, N5126, N1682, N200);
and AND4 (N5140, N5134, N4787, N1457, N3568);
xor XOR2 (N5141, N5136, N2224);
or OR2 (N5142, N5127, N825);
nor NOR4 (N5143, N5115, N4545, N2366, N281);
buf BUF1 (N5144, N5138);
buf BUF1 (N5145, N5139);
xor XOR2 (N5146, N5137, N3008);
xor XOR2 (N5147, N5125, N4217);
or OR2 (N5148, N5117, N3521);
nor NOR2 (N5149, N5133, N1778);
buf BUF1 (N5150, N5147);
nand NAND2 (N5151, N5150, N2816);
and AND4 (N5152, N5148, N2524, N3085, N989);
nor NOR4 (N5153, N5145, N3759, N4783, N1829);
buf BUF1 (N5154, N5141);
nor NOR2 (N5155, N5149, N998);
and AND3 (N5156, N5151, N4252, N1070);
and AND4 (N5157, N5146, N1351, N5153, N209);
xor XOR2 (N5158, N4158, N4072);
buf BUF1 (N5159, N5158);
nand NAND3 (N5160, N5144, N510, N799);
xor XOR2 (N5161, N5156, N865);
nand NAND3 (N5162, N5152, N148, N738);
nor NOR2 (N5163, N5159, N3704);
nand NAND4 (N5164, N5143, N1219, N4443, N3943);
or OR3 (N5165, N5142, N3833, N2792);
or OR4 (N5166, N5140, N1672, N1140, N1445);
or OR3 (N5167, N5157, N2731, N1544);
xor XOR2 (N5168, N5155, N3081);
xor XOR2 (N5169, N5165, N3806);
and AND2 (N5170, N5164, N1121);
not NOT1 (N5171, N5167);
or OR4 (N5172, N5171, N264, N3918, N1412);
buf BUF1 (N5173, N5169);
and AND4 (N5174, N5170, N1581, N3152, N4147);
buf BUF1 (N5175, N5168);
not NOT1 (N5176, N5173);
buf BUF1 (N5177, N5174);
nand NAND4 (N5178, N5176, N2001, N2762, N4510);
not NOT1 (N5179, N5161);
xor XOR2 (N5180, N5163, N1619);
nand NAND3 (N5181, N5177, N4985, N1166);
nor NOR4 (N5182, N5172, N4540, N810, N4584);
nor NOR3 (N5183, N5166, N1433, N2688);
nor NOR3 (N5184, N5183, N2889, N740);
buf BUF1 (N5185, N5184);
nor NOR2 (N5186, N5154, N224);
nor NOR2 (N5187, N5160, N4474);
or OR3 (N5188, N5180, N2791, N2346);
buf BUF1 (N5189, N5187);
or OR2 (N5190, N5181, N1160);
xor XOR2 (N5191, N5179, N2852);
or OR3 (N5192, N5182, N2268, N1687);
xor XOR2 (N5193, N5185, N1262);
nand NAND3 (N5194, N5186, N444, N2622);
and AND3 (N5195, N5178, N2667, N2902);
not NOT1 (N5196, N5191);
or OR4 (N5197, N5162, N1519, N4888, N1985);
or OR4 (N5198, N5196, N3794, N3032, N3708);
and AND4 (N5199, N5189, N4169, N3527, N1113);
buf BUF1 (N5200, N5199);
not NOT1 (N5201, N5200);
and AND3 (N5202, N5188, N3985, N4745);
nand NAND2 (N5203, N5193, N2915);
nor NOR3 (N5204, N5198, N1734, N1517);
and AND4 (N5205, N5175, N2200, N4380, N550);
or OR3 (N5206, N5201, N4698, N321);
nand NAND3 (N5207, N5202, N5030, N4631);
buf BUF1 (N5208, N5190);
or OR4 (N5209, N5207, N3005, N2039, N412);
and AND2 (N5210, N5206, N3453);
xor XOR2 (N5211, N5205, N1244);
xor XOR2 (N5212, N5203, N3349);
and AND3 (N5213, N5211, N1690, N3973);
xor XOR2 (N5214, N5212, N1418);
nor NOR2 (N5215, N5210, N457);
and AND4 (N5216, N5194, N2486, N854, N3865);
buf BUF1 (N5217, N5215);
buf BUF1 (N5218, N5213);
xor XOR2 (N5219, N5214, N1281);
not NOT1 (N5220, N5216);
and AND3 (N5221, N5218, N2379, N627);
nand NAND3 (N5222, N5219, N1178, N2589);
buf BUF1 (N5223, N5221);
xor XOR2 (N5224, N5197, N208);
buf BUF1 (N5225, N5209);
or OR2 (N5226, N5222, N2842);
nand NAND2 (N5227, N5225, N5005);
nor NOR4 (N5228, N5217, N5032, N974, N159);
xor XOR2 (N5229, N5220, N1169);
nor NOR4 (N5230, N5224, N17, N4070, N2868);
xor XOR2 (N5231, N5192, N2232);
buf BUF1 (N5232, N5195);
or OR3 (N5233, N5226, N1858, N1941);
nand NAND2 (N5234, N5233, N3477);
nand NAND2 (N5235, N5223, N622);
or OR3 (N5236, N5231, N2686, N5147);
nor NOR3 (N5237, N5227, N2780, N3052);
not NOT1 (N5238, N5228);
nor NOR2 (N5239, N5229, N574);
xor XOR2 (N5240, N5235, N2777);
and AND4 (N5241, N5236, N1138, N25, N2995);
nand NAND4 (N5242, N5237, N3555, N870, N862);
nor NOR3 (N5243, N5239, N1356, N394);
buf BUF1 (N5244, N5204);
xor XOR2 (N5245, N5241, N5223);
not NOT1 (N5246, N5245);
xor XOR2 (N5247, N5238, N3604);
nand NAND3 (N5248, N5230, N5120, N2075);
nor NOR2 (N5249, N5208, N3700);
nand NAND2 (N5250, N5246, N2142);
and AND2 (N5251, N5234, N1899);
and AND4 (N5252, N5242, N1285, N2710, N4730);
buf BUF1 (N5253, N5244);
not NOT1 (N5254, N5240);
and AND3 (N5255, N5252, N4337, N3642);
and AND3 (N5256, N5232, N2912, N4484);
or OR2 (N5257, N5253, N586);
and AND2 (N5258, N5243, N5132);
nor NOR2 (N5259, N5254, N4574);
or OR4 (N5260, N5256, N4753, N5163, N315);
nand NAND2 (N5261, N5260, N1471);
and AND4 (N5262, N5250, N3951, N3813, N4328);
nand NAND2 (N5263, N5262, N3201);
nand NAND4 (N5264, N5248, N2491, N1537, N1205);
and AND3 (N5265, N5259, N3119, N678);
nand NAND2 (N5266, N5261, N1522);
and AND4 (N5267, N5249, N1473, N4201, N1201);
not NOT1 (N5268, N5266);
not NOT1 (N5269, N5257);
xor XOR2 (N5270, N5269, N3829);
nor NOR4 (N5271, N5258, N5077, N2066, N3231);
nor NOR2 (N5272, N5267, N1843);
buf BUF1 (N5273, N5271);
not NOT1 (N5274, N5273);
buf BUF1 (N5275, N5247);
not NOT1 (N5276, N5274);
nor NOR2 (N5277, N5276, N3074);
not NOT1 (N5278, N5268);
or OR4 (N5279, N5275, N1478, N4694, N2125);
xor XOR2 (N5280, N5272, N4608);
nor NOR3 (N5281, N5280, N4898, N2637);
buf BUF1 (N5282, N5255);
nand NAND4 (N5283, N5270, N4881, N3091, N3354);
and AND4 (N5284, N5278, N7, N3464, N2076);
nand NAND2 (N5285, N5264, N939);
not NOT1 (N5286, N5282);
not NOT1 (N5287, N5251);
not NOT1 (N5288, N5287);
or OR4 (N5289, N5263, N1939, N4032, N5061);
or OR4 (N5290, N5283, N941, N3073, N4214);
and AND2 (N5291, N5279, N3393);
nand NAND4 (N5292, N5277, N1846, N3995, N5019);
or OR2 (N5293, N5290, N3718);
xor XOR2 (N5294, N5286, N3193);
or OR3 (N5295, N5294, N2744, N258);
and AND4 (N5296, N5288, N3709, N2659, N4191);
nand NAND3 (N5297, N5296, N2646, N5211);
or OR4 (N5298, N5291, N1389, N2763, N1698);
nand NAND2 (N5299, N5298, N576);
nor NOR3 (N5300, N5295, N193, N3555);
and AND4 (N5301, N5281, N2097, N491, N4533);
and AND3 (N5302, N5293, N1637, N3975);
and AND4 (N5303, N5292, N531, N2880, N3214);
or OR4 (N5304, N5289, N2138, N2963, N3622);
xor XOR2 (N5305, N5284, N670);
and AND4 (N5306, N5301, N3293, N2687, N1111);
buf BUF1 (N5307, N5306);
nor NOR2 (N5308, N5299, N3567);
nor NOR2 (N5309, N5302, N2425);
and AND4 (N5310, N5309, N1847, N2888, N1750);
nand NAND3 (N5311, N5285, N220, N2112);
not NOT1 (N5312, N5297);
xor XOR2 (N5313, N5310, N2548);
buf BUF1 (N5314, N5308);
or OR2 (N5315, N5312, N4585);
nor NOR3 (N5316, N5303, N3722, N2895);
nor NOR4 (N5317, N5313, N4719, N82, N4432);
nand NAND3 (N5318, N5316, N3192, N4146);
xor XOR2 (N5319, N5304, N56);
xor XOR2 (N5320, N5265, N3288);
buf BUF1 (N5321, N5317);
and AND2 (N5322, N5314, N359);
nand NAND3 (N5323, N5315, N2363, N4501);
nor NOR3 (N5324, N5307, N2592, N1680);
nand NAND4 (N5325, N5300, N723, N573, N1745);
buf BUF1 (N5326, N5311);
nand NAND4 (N5327, N5321, N4467, N3609, N757);
nor NOR2 (N5328, N5324, N4522);
and AND4 (N5329, N5326, N4172, N2628, N2681);
xor XOR2 (N5330, N5329, N596);
not NOT1 (N5331, N5325);
not NOT1 (N5332, N5319);
buf BUF1 (N5333, N5323);
or OR4 (N5334, N5331, N2340, N3170, N3840);
nor NOR4 (N5335, N5332, N3960, N4256, N4314);
or OR2 (N5336, N5327, N2215);
buf BUF1 (N5337, N5334);
nor NOR3 (N5338, N5333, N225, N2726);
buf BUF1 (N5339, N5330);
and AND2 (N5340, N5305, N1087);
nand NAND3 (N5341, N5340, N184, N3864);
nor NOR2 (N5342, N5341, N3857);
buf BUF1 (N5343, N5328);
not NOT1 (N5344, N5335);
not NOT1 (N5345, N5338);
nor NOR3 (N5346, N5322, N2688, N1924);
xor XOR2 (N5347, N5346, N2433);
buf BUF1 (N5348, N5320);
not NOT1 (N5349, N5318);
or OR2 (N5350, N5349, N534);
not NOT1 (N5351, N5342);
nand NAND2 (N5352, N5343, N112);
or OR2 (N5353, N5347, N1338);
not NOT1 (N5354, N5350);
xor XOR2 (N5355, N5339, N3660);
not NOT1 (N5356, N5354);
xor XOR2 (N5357, N5353, N1789);
buf BUF1 (N5358, N5357);
nand NAND2 (N5359, N5356, N685);
xor XOR2 (N5360, N5351, N800);
not NOT1 (N5361, N5355);
xor XOR2 (N5362, N5360, N725);
not NOT1 (N5363, N5348);
and AND4 (N5364, N5352, N2672, N1015, N4018);
and AND2 (N5365, N5363, N3202);
xor XOR2 (N5366, N5364, N398);
or OR4 (N5367, N5359, N2550, N1126, N4177);
or OR3 (N5368, N5367, N4960, N3241);
buf BUF1 (N5369, N5358);
nand NAND2 (N5370, N5337, N1486);
or OR3 (N5371, N5368, N3050, N4379);
or OR3 (N5372, N5365, N5240, N4926);
nand NAND3 (N5373, N5369, N2662, N5067);
not NOT1 (N5374, N5361);
xor XOR2 (N5375, N5372, N186);
nor NOR2 (N5376, N5374, N79);
or OR4 (N5377, N5373, N1888, N275, N262);
and AND3 (N5378, N5362, N3309, N2914);
nand NAND4 (N5379, N5345, N2785, N5170, N4352);
or OR3 (N5380, N5370, N1378, N4266);
buf BUF1 (N5381, N5379);
or OR2 (N5382, N5381, N3789);
buf BUF1 (N5383, N5344);
not NOT1 (N5384, N5377);
and AND3 (N5385, N5376, N137, N1686);
or OR2 (N5386, N5371, N2381);
or OR3 (N5387, N5383, N3192, N4083);
or OR4 (N5388, N5366, N3137, N4607, N464);
xor XOR2 (N5389, N5375, N3441);
and AND3 (N5390, N5388, N3578, N267);
xor XOR2 (N5391, N5387, N1028);
nand NAND3 (N5392, N5382, N3064, N1712);
nor NOR3 (N5393, N5390, N3624, N4052);
nand NAND3 (N5394, N5378, N947, N2128);
and AND3 (N5395, N5336, N3868, N3802);
nor NOR2 (N5396, N5394, N119);
not NOT1 (N5397, N5380);
or OR3 (N5398, N5389, N5353, N501);
nand NAND4 (N5399, N5385, N171, N2265, N1130);
not NOT1 (N5400, N5399);
buf BUF1 (N5401, N5397);
and AND3 (N5402, N5401, N2248, N2944);
or OR2 (N5403, N5392, N2333);
and AND2 (N5404, N5386, N3171);
buf BUF1 (N5405, N5393);
nand NAND4 (N5406, N5403, N4024, N5059, N2854);
or OR2 (N5407, N5400, N4043);
and AND4 (N5408, N5407, N1422, N4801, N661);
buf BUF1 (N5409, N5406);
xor XOR2 (N5410, N5405, N3113);
and AND3 (N5411, N5396, N3949, N1709);
nor NOR4 (N5412, N5395, N3137, N2130, N3352);
xor XOR2 (N5413, N5410, N4466);
xor XOR2 (N5414, N5408, N488);
nand NAND4 (N5415, N5413, N5156, N4070, N2056);
or OR2 (N5416, N5411, N2462);
buf BUF1 (N5417, N5414);
and AND2 (N5418, N5391, N3963);
or OR4 (N5419, N5402, N4937, N1754, N4536);
nand NAND3 (N5420, N5409, N1802, N938);
xor XOR2 (N5421, N5420, N3790);
buf BUF1 (N5422, N5415);
nor NOR3 (N5423, N5421, N1267, N1240);
xor XOR2 (N5424, N5422, N442);
buf BUF1 (N5425, N5404);
not NOT1 (N5426, N5416);
buf BUF1 (N5427, N5424);
xor XOR2 (N5428, N5418, N35);
and AND2 (N5429, N5426, N1230);
or OR4 (N5430, N5423, N3746, N1796, N1027);
and AND2 (N5431, N5419, N1638);
or OR4 (N5432, N5431, N4049, N1425, N2704);
and AND4 (N5433, N5384, N3234, N3458, N4292);
and AND4 (N5434, N5425, N4921, N697, N1585);
buf BUF1 (N5435, N5412);
or OR2 (N5436, N5398, N2827);
nor NOR2 (N5437, N5429, N1628);
buf BUF1 (N5438, N5432);
buf BUF1 (N5439, N5434);
or OR2 (N5440, N5436, N337);
nor NOR4 (N5441, N5435, N158, N1971, N1916);
nor NOR4 (N5442, N5439, N335, N415, N5315);
buf BUF1 (N5443, N5442);
not NOT1 (N5444, N5433);
not NOT1 (N5445, N5438);
buf BUF1 (N5446, N5445);
or OR2 (N5447, N5443, N3286);
nand NAND2 (N5448, N5430, N1031);
xor XOR2 (N5449, N5437, N682);
nand NAND4 (N5450, N5428, N838, N1587, N3574);
and AND2 (N5451, N5444, N2880);
nor NOR2 (N5452, N5417, N3662);
nand NAND4 (N5453, N5441, N4637, N210, N3363);
not NOT1 (N5454, N5453);
or OR4 (N5455, N5427, N1836, N4552, N4736);
and AND2 (N5456, N5455, N4597);
and AND2 (N5457, N5449, N1196);
nor NOR4 (N5458, N5451, N2323, N3888, N1607);
buf BUF1 (N5459, N5456);
nand NAND3 (N5460, N5446, N2542, N1039);
or OR2 (N5461, N5458, N1270);
or OR4 (N5462, N5460, N226, N549, N585);
not NOT1 (N5463, N5450);
nor NOR4 (N5464, N5457, N3944, N5152, N2899);
or OR2 (N5465, N5452, N1199);
not NOT1 (N5466, N5459);
xor XOR2 (N5467, N5461, N1975);
buf BUF1 (N5468, N5462);
xor XOR2 (N5469, N5465, N876);
not NOT1 (N5470, N5466);
not NOT1 (N5471, N5440);
nor NOR4 (N5472, N5463, N4662, N531, N1053);
nor NOR3 (N5473, N5468, N3743, N4243);
nor NOR3 (N5474, N5467, N5368, N2387);
nand NAND4 (N5475, N5448, N4964, N3735, N3442);
not NOT1 (N5476, N5470);
xor XOR2 (N5477, N5475, N412);
xor XOR2 (N5478, N5477, N822);
not NOT1 (N5479, N5447);
buf BUF1 (N5480, N5474);
or OR2 (N5481, N5472, N3984);
nor NOR3 (N5482, N5480, N5417, N3142);
not NOT1 (N5483, N5464);
not NOT1 (N5484, N5483);
nand NAND4 (N5485, N5481, N133, N4807, N4891);
not NOT1 (N5486, N5485);
xor XOR2 (N5487, N5454, N4966);
buf BUF1 (N5488, N5486);
xor XOR2 (N5489, N5488, N3275);
buf BUF1 (N5490, N5487);
xor XOR2 (N5491, N5479, N3348);
xor XOR2 (N5492, N5491, N2474);
nand NAND4 (N5493, N5484, N1351, N4443, N359);
nor NOR3 (N5494, N5476, N175, N1214);
nand NAND3 (N5495, N5489, N3488, N3136);
or OR3 (N5496, N5494, N4282, N2598);
or OR4 (N5497, N5490, N82, N1140, N2672);
buf BUF1 (N5498, N5473);
xor XOR2 (N5499, N5496, N135);
nor NOR4 (N5500, N5498, N2040, N668, N1610);
nand NAND4 (N5501, N5492, N3567, N4922, N3081);
and AND2 (N5502, N5478, N2730);
or OR3 (N5503, N5482, N591, N297);
buf BUF1 (N5504, N5497);
buf BUF1 (N5505, N5501);
nor NOR4 (N5506, N5504, N3779, N3726, N5336);
or OR2 (N5507, N5503, N4984);
and AND2 (N5508, N5500, N1784);
and AND2 (N5509, N5499, N1648);
nand NAND2 (N5510, N5506, N3083);
buf BUF1 (N5511, N5471);
and AND4 (N5512, N5495, N4962, N2696, N2475);
or OR3 (N5513, N5493, N1932, N3192);
nand NAND3 (N5514, N5505, N2790, N2665);
nor NOR4 (N5515, N5513, N3812, N3647, N3650);
nor NOR4 (N5516, N5515, N4912, N1310, N90);
nor NOR2 (N5517, N5511, N2087);
and AND3 (N5518, N5510, N5486, N1277);
buf BUF1 (N5519, N5518);
and AND2 (N5520, N5508, N4879);
and AND4 (N5521, N5512, N3446, N1326, N3976);
or OR4 (N5522, N5507, N3704, N4522, N4051);
buf BUF1 (N5523, N5519);
buf BUF1 (N5524, N5521);
and AND4 (N5525, N5524, N3022, N522, N509);
buf BUF1 (N5526, N5502);
buf BUF1 (N5527, N5523);
and AND2 (N5528, N5509, N5504);
or OR4 (N5529, N5517, N284, N4684, N2641);
nand NAND2 (N5530, N5529, N668);
or OR4 (N5531, N5530, N2212, N160, N2172);
and AND3 (N5532, N5516, N2215, N4630);
nor NOR4 (N5533, N5532, N974, N1542, N1910);
not NOT1 (N5534, N5526);
buf BUF1 (N5535, N5522);
not NOT1 (N5536, N5520);
nand NAND4 (N5537, N5536, N90, N2159, N2794);
buf BUF1 (N5538, N5469);
not NOT1 (N5539, N5538);
or OR2 (N5540, N5535, N2837);
xor XOR2 (N5541, N5534, N4963);
nand NAND3 (N5542, N5527, N4801, N423);
buf BUF1 (N5543, N5537);
xor XOR2 (N5544, N5542, N3380);
not NOT1 (N5545, N5533);
nor NOR4 (N5546, N5528, N1935, N4272, N5476);
or OR3 (N5547, N5540, N4120, N2826);
xor XOR2 (N5548, N5546, N612);
nor NOR2 (N5549, N5544, N1708);
not NOT1 (N5550, N5549);
or OR2 (N5551, N5531, N5260);
nand NAND3 (N5552, N5543, N868, N2187);
nor NOR4 (N5553, N5552, N4037, N5233, N257);
or OR2 (N5554, N5545, N4926);
xor XOR2 (N5555, N5539, N408);
buf BUF1 (N5556, N5514);
nor NOR3 (N5557, N5525, N4353, N2993);
xor XOR2 (N5558, N5555, N2327);
or OR3 (N5559, N5550, N4019, N1527);
buf BUF1 (N5560, N5559);
or OR4 (N5561, N5560, N5508, N1021, N1597);
and AND3 (N5562, N5547, N3089, N5234);
nand NAND4 (N5563, N5557, N4395, N1528, N2895);
not NOT1 (N5564, N5554);
and AND3 (N5565, N5564, N5357, N3422);
nor NOR3 (N5566, N5565, N4809, N4741);
not NOT1 (N5567, N5558);
xor XOR2 (N5568, N5551, N3737);
or OR3 (N5569, N5568, N5531, N1026);
nand NAND4 (N5570, N5563, N2263, N4582, N5521);
not NOT1 (N5571, N5541);
buf BUF1 (N5572, N5566);
nor NOR2 (N5573, N5567, N4866);
nand NAND2 (N5574, N5570, N4085);
or OR4 (N5575, N5569, N57, N3231, N5223);
nand NAND2 (N5576, N5548, N2677);
nor NOR3 (N5577, N5562, N3858, N3150);
xor XOR2 (N5578, N5561, N2114);
not NOT1 (N5579, N5553);
or OR4 (N5580, N5556, N3238, N3338, N1562);
xor XOR2 (N5581, N5580, N3860);
nand NAND2 (N5582, N5578, N2250);
not NOT1 (N5583, N5572);
nand NAND3 (N5584, N5574, N2378, N813);
not NOT1 (N5585, N5576);
or OR2 (N5586, N5571, N5310);
nand NAND4 (N5587, N5575, N3021, N4532, N3168);
xor XOR2 (N5588, N5587, N4361);
buf BUF1 (N5589, N5577);
xor XOR2 (N5590, N5589, N3718);
xor XOR2 (N5591, N5582, N3458);
nor NOR2 (N5592, N5585, N1508);
nor NOR3 (N5593, N5581, N2721, N2710);
nor NOR3 (N5594, N5573, N3562, N4129);
and AND4 (N5595, N5588, N727, N499, N4643);
nor NOR3 (N5596, N5583, N356, N583);
nor NOR4 (N5597, N5594, N2771, N4181, N2141);
and AND3 (N5598, N5596, N392, N4242);
xor XOR2 (N5599, N5593, N2764);
nor NOR3 (N5600, N5584, N3821, N3497);
xor XOR2 (N5601, N5599, N781);
xor XOR2 (N5602, N5595, N3474);
not NOT1 (N5603, N5597);
buf BUF1 (N5604, N5591);
nand NAND2 (N5605, N5590, N3533);
buf BUF1 (N5606, N5598);
not NOT1 (N5607, N5579);
or OR2 (N5608, N5602, N1618);
nor NOR4 (N5609, N5608, N2405, N1886, N3545);
nor NOR3 (N5610, N5607, N1389, N3391);
nand NAND3 (N5611, N5604, N4953, N3911);
nor NOR2 (N5612, N5592, N4185);
and AND2 (N5613, N5601, N1714);
or OR3 (N5614, N5610, N4429, N4625);
xor XOR2 (N5615, N5614, N4036);
buf BUF1 (N5616, N5603);
xor XOR2 (N5617, N5612, N4067);
buf BUF1 (N5618, N5605);
xor XOR2 (N5619, N5609, N5554);
and AND2 (N5620, N5617, N3385);
nand NAND4 (N5621, N5586, N1180, N1427, N4978);
xor XOR2 (N5622, N5616, N3612);
not NOT1 (N5623, N5600);
buf BUF1 (N5624, N5615);
nor NOR4 (N5625, N5622, N782, N4456, N933);
and AND2 (N5626, N5625, N3466);
xor XOR2 (N5627, N5620, N2887);
and AND3 (N5628, N5618, N2808, N5081);
and AND4 (N5629, N5611, N3512, N2326, N215);
or OR2 (N5630, N5623, N4624);
xor XOR2 (N5631, N5627, N2565);
or OR3 (N5632, N5629, N3312, N1509);
buf BUF1 (N5633, N5631);
buf BUF1 (N5634, N5606);
nor NOR2 (N5635, N5630, N2231);
xor XOR2 (N5636, N5633, N226);
and AND2 (N5637, N5626, N3642);
buf BUF1 (N5638, N5621);
xor XOR2 (N5639, N5635, N4243);
nand NAND2 (N5640, N5637, N3804);
not NOT1 (N5641, N5640);
not NOT1 (N5642, N5619);
nand NAND4 (N5643, N5639, N691, N4571, N1454);
not NOT1 (N5644, N5613);
nor NOR3 (N5645, N5628, N819, N4685);
and AND3 (N5646, N5645, N5050, N683);
nand NAND4 (N5647, N5642, N621, N1240, N2222);
and AND4 (N5648, N5624, N3762, N4388, N91);
nor NOR3 (N5649, N5634, N1014, N1684);
buf BUF1 (N5650, N5638);
not NOT1 (N5651, N5632);
buf BUF1 (N5652, N5649);
xor XOR2 (N5653, N5647, N870);
xor XOR2 (N5654, N5648, N3107);
nand NAND2 (N5655, N5636, N1776);
not NOT1 (N5656, N5646);
buf BUF1 (N5657, N5652);
or OR2 (N5658, N5656, N4993);
buf BUF1 (N5659, N5658);
and AND3 (N5660, N5659, N4730, N3099);
buf BUF1 (N5661, N5641);
nor NOR3 (N5662, N5643, N4425, N5615);
nor NOR2 (N5663, N5662, N1257);
buf BUF1 (N5664, N5655);
buf BUF1 (N5665, N5663);
or OR3 (N5666, N5664, N4268, N2117);
buf BUF1 (N5667, N5660);
xor XOR2 (N5668, N5644, N2234);
nand NAND2 (N5669, N5668, N4551);
buf BUF1 (N5670, N5661);
and AND2 (N5671, N5670, N2614);
and AND3 (N5672, N5651, N2476, N2886);
nand NAND3 (N5673, N5657, N5298, N452);
nor NOR2 (N5674, N5653, N377);
or OR3 (N5675, N5650, N1607, N3243);
nand NAND2 (N5676, N5666, N5525);
buf BUF1 (N5677, N5673);
buf BUF1 (N5678, N5674);
or OR4 (N5679, N5676, N1051, N4810, N2873);
or OR4 (N5680, N5667, N5358, N5226, N3393);
nand NAND3 (N5681, N5675, N2213, N1296);
or OR3 (N5682, N5680, N736, N3114);
nand NAND3 (N5683, N5678, N1064, N2916);
xor XOR2 (N5684, N5682, N2891);
or OR2 (N5685, N5669, N4463);
nand NAND2 (N5686, N5671, N695);
nand NAND2 (N5687, N5679, N2063);
nor NOR3 (N5688, N5687, N3277, N814);
buf BUF1 (N5689, N5684);
nand NAND2 (N5690, N5689, N2959);
nor NOR3 (N5691, N5672, N2662, N1127);
nand NAND3 (N5692, N5677, N2650, N3033);
nand NAND3 (N5693, N5681, N3003, N2145);
or OR2 (N5694, N5692, N1737);
nor NOR2 (N5695, N5690, N888);
not NOT1 (N5696, N5665);
not NOT1 (N5697, N5694);
and AND4 (N5698, N5683, N154, N1216, N5071);
nand NAND4 (N5699, N5685, N774, N2062, N3040);
nor NOR3 (N5700, N5686, N261, N1374);
not NOT1 (N5701, N5699);
xor XOR2 (N5702, N5701, N700);
xor XOR2 (N5703, N5702, N2770);
nor NOR3 (N5704, N5654, N4244, N1063);
xor XOR2 (N5705, N5697, N5637);
xor XOR2 (N5706, N5704, N3847);
not NOT1 (N5707, N5705);
and AND4 (N5708, N5698, N2012, N4409, N5634);
not NOT1 (N5709, N5707);
nand NAND2 (N5710, N5708, N3180);
not NOT1 (N5711, N5695);
and AND4 (N5712, N5711, N5008, N1861, N3149);
and AND4 (N5713, N5693, N847, N2114, N1813);
or OR3 (N5714, N5713, N3801, N805);
and AND4 (N5715, N5712, N2197, N4050, N5694);
nand NAND3 (N5716, N5691, N5516, N2773);
buf BUF1 (N5717, N5714);
and AND3 (N5718, N5710, N2975, N4247);
nand NAND2 (N5719, N5696, N9);
and AND4 (N5720, N5703, N450, N3244, N4114);
buf BUF1 (N5721, N5715);
or OR3 (N5722, N5706, N1287, N1080);
or OR3 (N5723, N5709, N445, N2558);
nand NAND2 (N5724, N5721, N4301);
nor NOR4 (N5725, N5700, N3588, N3487, N3101);
not NOT1 (N5726, N5718);
not NOT1 (N5727, N5726);
and AND4 (N5728, N5688, N4262, N4448, N2875);
nand NAND4 (N5729, N5720, N2925, N467, N3339);
or OR2 (N5730, N5724, N3013);
xor XOR2 (N5731, N5722, N4787);
nor NOR4 (N5732, N5731, N2572, N4178, N5643);
nor NOR2 (N5733, N5727, N4155);
not NOT1 (N5734, N5723);
nand NAND3 (N5735, N5734, N1301, N3021);
or OR2 (N5736, N5717, N3256);
not NOT1 (N5737, N5728);
not NOT1 (N5738, N5737);
or OR4 (N5739, N5716, N4075, N2627, N2291);
or OR2 (N5740, N5736, N440);
nand NAND2 (N5741, N5735, N5716);
and AND2 (N5742, N5725, N529);
nand NAND2 (N5743, N5740, N205);
nor NOR4 (N5744, N5742, N5545, N319, N636);
nor NOR2 (N5745, N5729, N5549);
xor XOR2 (N5746, N5741, N1641);
and AND3 (N5747, N5732, N3230, N2283);
nor NOR3 (N5748, N5739, N2501, N808);
xor XOR2 (N5749, N5745, N273);
or OR4 (N5750, N5744, N894, N4728, N2377);
xor XOR2 (N5751, N5748, N80);
and AND3 (N5752, N5749, N3767, N3480);
not NOT1 (N5753, N5747);
and AND4 (N5754, N5730, N1486, N3698, N4076);
nor NOR4 (N5755, N5743, N1278, N5449, N4496);
nor NOR3 (N5756, N5755, N4752, N362);
or OR3 (N5757, N5754, N4347, N3938);
nor NOR3 (N5758, N5733, N3459, N3626);
buf BUF1 (N5759, N5738);
nor NOR2 (N5760, N5758, N3752);
not NOT1 (N5761, N5750);
xor XOR2 (N5762, N5761, N782);
buf BUF1 (N5763, N5719);
not NOT1 (N5764, N5753);
or OR3 (N5765, N5752, N1520, N3795);
xor XOR2 (N5766, N5762, N2680);
nand NAND3 (N5767, N5757, N4070, N4683);
and AND2 (N5768, N5751, N3166);
or OR4 (N5769, N5764, N2891, N2173, N4669);
nand NAND3 (N5770, N5768, N3128, N913);
or OR2 (N5771, N5765, N1069);
nor NOR4 (N5772, N5759, N2030, N2557, N1993);
and AND2 (N5773, N5746, N1178);
and AND4 (N5774, N5770, N2447, N3116, N1575);
or OR4 (N5775, N5766, N876, N5698, N739);
buf BUF1 (N5776, N5774);
xor XOR2 (N5777, N5756, N2368);
nor NOR2 (N5778, N5777, N4896);
xor XOR2 (N5779, N5775, N453);
buf BUF1 (N5780, N5772);
xor XOR2 (N5781, N5780, N4374);
nand NAND3 (N5782, N5767, N1613, N1900);
nor NOR3 (N5783, N5773, N3947, N5519);
not NOT1 (N5784, N5781);
or OR4 (N5785, N5763, N479, N4683, N5510);
nand NAND3 (N5786, N5776, N1930, N626);
not NOT1 (N5787, N5760);
or OR3 (N5788, N5786, N444, N292);
or OR3 (N5789, N5788, N751, N131);
buf BUF1 (N5790, N5782);
not NOT1 (N5791, N5769);
and AND4 (N5792, N5779, N2005, N1134, N2020);
and AND2 (N5793, N5789, N3252);
or OR3 (N5794, N5784, N1428, N1175);
buf BUF1 (N5795, N5794);
or OR3 (N5796, N5783, N1104, N2484);
nor NOR2 (N5797, N5785, N183);
not NOT1 (N5798, N5797);
xor XOR2 (N5799, N5795, N4666);
buf BUF1 (N5800, N5778);
not NOT1 (N5801, N5798);
nand NAND3 (N5802, N5801, N1354, N208);
buf BUF1 (N5803, N5800);
not NOT1 (N5804, N5802);
buf BUF1 (N5805, N5793);
xor XOR2 (N5806, N5803, N5663);
and AND3 (N5807, N5787, N4250, N1992);
buf BUF1 (N5808, N5796);
nand NAND4 (N5809, N5771, N290, N5093, N4375);
nor NOR3 (N5810, N5799, N5711, N502);
nor NOR4 (N5811, N5807, N2056, N2740, N4903);
buf BUF1 (N5812, N5792);
nor NOR4 (N5813, N5810, N668, N3916, N3911);
nand NAND4 (N5814, N5811, N1319, N3641, N3421);
xor XOR2 (N5815, N5814, N3601);
nand NAND4 (N5816, N5808, N146, N2288, N2538);
not NOT1 (N5817, N5791);
nand NAND4 (N5818, N5816, N4143, N3900, N5696);
not NOT1 (N5819, N5790);
or OR4 (N5820, N5817, N5508, N4738, N2029);
or OR2 (N5821, N5812, N3637);
or OR4 (N5822, N5818, N5463, N3402, N2667);
nor NOR2 (N5823, N5806, N4306);
not NOT1 (N5824, N5805);
and AND2 (N5825, N5821, N1619);
buf BUF1 (N5826, N5809);
not NOT1 (N5827, N5813);
buf BUF1 (N5828, N5827);
nor NOR3 (N5829, N5815, N3095, N5232);
nand NAND2 (N5830, N5828, N1920);
buf BUF1 (N5831, N5825);
buf BUF1 (N5832, N5804);
nand NAND3 (N5833, N5826, N1375, N5282);
and AND4 (N5834, N5822, N4707, N3629, N408);
and AND2 (N5835, N5833, N599);
buf BUF1 (N5836, N5829);
nand NAND3 (N5837, N5820, N26, N3867);
nand NAND3 (N5838, N5836, N3384, N3487);
buf BUF1 (N5839, N5838);
not NOT1 (N5840, N5837);
xor XOR2 (N5841, N5831, N2225);
or OR4 (N5842, N5840, N4394, N5293, N4693);
not NOT1 (N5843, N5839);
buf BUF1 (N5844, N5824);
nor NOR3 (N5845, N5823, N4849, N1227);
nor NOR2 (N5846, N5835, N4257);
not NOT1 (N5847, N5834);
nand NAND3 (N5848, N5841, N1720, N4282);
or OR4 (N5849, N5847, N3069, N4277, N5037);
not NOT1 (N5850, N5845);
xor XOR2 (N5851, N5819, N2937);
not NOT1 (N5852, N5846);
nand NAND3 (N5853, N5844, N4146, N4041);
nor NOR4 (N5854, N5832, N446, N4661, N2420);
xor XOR2 (N5855, N5848, N88);
and AND4 (N5856, N5853, N3437, N5127, N4721);
buf BUF1 (N5857, N5852);
buf BUF1 (N5858, N5856);
or OR4 (N5859, N5858, N5649, N1687, N787);
or OR2 (N5860, N5854, N3155);
or OR4 (N5861, N5842, N2864, N2038, N5698);
and AND2 (N5862, N5849, N4390);
not NOT1 (N5863, N5830);
and AND2 (N5864, N5843, N1869);
or OR4 (N5865, N5863, N2039, N3879, N1878);
xor XOR2 (N5866, N5851, N4596);
nor NOR3 (N5867, N5864, N2848, N841);
xor XOR2 (N5868, N5855, N4165);
and AND2 (N5869, N5861, N2607);
and AND2 (N5870, N5850, N5164);
buf BUF1 (N5871, N5869);
and AND3 (N5872, N5865, N16, N847);
buf BUF1 (N5873, N5859);
not NOT1 (N5874, N5872);
not NOT1 (N5875, N5868);
buf BUF1 (N5876, N5873);
xor XOR2 (N5877, N5867, N3375);
not NOT1 (N5878, N5866);
xor XOR2 (N5879, N5857, N935);
nand NAND3 (N5880, N5862, N4829, N3400);
xor XOR2 (N5881, N5880, N1511);
and AND4 (N5882, N5871, N4548, N1947, N3084);
or OR2 (N5883, N5878, N4813);
buf BUF1 (N5884, N5881);
not NOT1 (N5885, N5860);
nand NAND3 (N5886, N5884, N73, N2922);
xor XOR2 (N5887, N5879, N2471);
buf BUF1 (N5888, N5870);
buf BUF1 (N5889, N5874);
xor XOR2 (N5890, N5887, N1621);
or OR3 (N5891, N5886, N3572, N4793);
nand NAND3 (N5892, N5885, N5398, N3695);
nand NAND3 (N5893, N5890, N3737, N81);
and AND2 (N5894, N5888, N5206);
and AND2 (N5895, N5889, N5557);
or OR3 (N5896, N5892, N3466, N3388);
not NOT1 (N5897, N5891);
and AND4 (N5898, N5895, N2278, N1481, N5850);
buf BUF1 (N5899, N5897);
not NOT1 (N5900, N5894);
or OR2 (N5901, N5899, N5847);
not NOT1 (N5902, N5900);
nor NOR3 (N5903, N5896, N903, N2916);
and AND4 (N5904, N5898, N4140, N3551, N2106);
or OR4 (N5905, N5882, N520, N368, N4176);
not NOT1 (N5906, N5905);
not NOT1 (N5907, N5903);
nor NOR4 (N5908, N5904, N777, N185, N4152);
and AND2 (N5909, N5893, N2740);
and AND3 (N5910, N5883, N4062, N917);
or OR2 (N5911, N5875, N2205);
xor XOR2 (N5912, N5909, N796);
and AND4 (N5913, N5907, N5139, N1051, N4679);
xor XOR2 (N5914, N5910, N936);
nor NOR4 (N5915, N5913, N4940, N5448, N855);
xor XOR2 (N5916, N5912, N122);
buf BUF1 (N5917, N5908);
not NOT1 (N5918, N5916);
buf BUF1 (N5919, N5902);
xor XOR2 (N5920, N5918, N651);
buf BUF1 (N5921, N5919);
xor XOR2 (N5922, N5915, N2012);
xor XOR2 (N5923, N5901, N2007);
xor XOR2 (N5924, N5920, N2068);
buf BUF1 (N5925, N5911);
buf BUF1 (N5926, N5923);
nand NAND2 (N5927, N5924, N5693);
and AND4 (N5928, N5927, N472, N5492, N1769);
and AND4 (N5929, N5921, N5308, N3752, N5552);
nor NOR2 (N5930, N5906, N858);
xor XOR2 (N5931, N5926, N4798);
nor NOR2 (N5932, N5930, N2792);
nor NOR4 (N5933, N5931, N2676, N285, N5158);
or OR4 (N5934, N5877, N5812, N2649, N1278);
nand NAND4 (N5935, N5932, N4699, N1780, N5750);
xor XOR2 (N5936, N5928, N4482);
or OR4 (N5937, N5929, N734, N4627, N3499);
or OR3 (N5938, N5914, N583, N677);
buf BUF1 (N5939, N5934);
not NOT1 (N5940, N5939);
nor NOR4 (N5941, N5925, N4051, N4758, N3131);
xor XOR2 (N5942, N5941, N1750);
nor NOR3 (N5943, N5937, N5131, N1684);
xor XOR2 (N5944, N5876, N1179);
or OR4 (N5945, N5917, N1141, N3861, N1937);
buf BUF1 (N5946, N5942);
buf BUF1 (N5947, N5938);
or OR2 (N5948, N5933, N2983);
xor XOR2 (N5949, N5946, N5674);
not NOT1 (N5950, N5944);
nand NAND4 (N5951, N5949, N5628, N237, N361);
buf BUF1 (N5952, N5947);
or OR3 (N5953, N5952, N1898, N1815);
xor XOR2 (N5954, N5951, N2520);
nor NOR2 (N5955, N5936, N5762);
nand NAND4 (N5956, N5948, N2952, N3433, N2072);
and AND4 (N5957, N5922, N1471, N2303, N3844);
nor NOR3 (N5958, N5956, N5385, N3737);
buf BUF1 (N5959, N5957);
or OR3 (N5960, N5945, N4941, N5730);
xor XOR2 (N5961, N5959, N491);
or OR4 (N5962, N5961, N293, N1508, N3093);
not NOT1 (N5963, N5962);
nand NAND2 (N5964, N5963, N2658);
or OR2 (N5965, N5953, N2874);
or OR3 (N5966, N5954, N2535, N1289);
or OR2 (N5967, N5935, N5148);
and AND4 (N5968, N5943, N3253, N5180, N3819);
not NOT1 (N5969, N5958);
nor NOR2 (N5970, N5940, N888);
or OR3 (N5971, N5969, N2785, N4496);
xor XOR2 (N5972, N5971, N1760);
xor XOR2 (N5973, N5964, N5798);
not NOT1 (N5974, N5973);
xor XOR2 (N5975, N5966, N5308);
and AND4 (N5976, N5974, N4574, N1810, N3361);
and AND4 (N5977, N5972, N4434, N149, N313);
buf BUF1 (N5978, N5955);
or OR2 (N5979, N5965, N5425);
and AND3 (N5980, N5978, N5361, N3499);
xor XOR2 (N5981, N5968, N965);
nor NOR3 (N5982, N5979, N5206, N3486);
and AND3 (N5983, N5982, N2302, N144);
not NOT1 (N5984, N5970);
not NOT1 (N5985, N5981);
not NOT1 (N5986, N5983);
and AND2 (N5987, N5986, N91);
nand NAND2 (N5988, N5984, N2787);
buf BUF1 (N5989, N5960);
nor NOR4 (N5990, N5977, N3342, N3983, N1361);
buf BUF1 (N5991, N5976);
nor NOR4 (N5992, N5950, N349, N739, N5229);
and AND3 (N5993, N5967, N1941, N5220);
and AND4 (N5994, N5985, N5020, N1057, N849);
buf BUF1 (N5995, N5987);
nor NOR2 (N5996, N5975, N290);
not NOT1 (N5997, N5994);
or OR3 (N5998, N5990, N4412, N2627);
and AND3 (N5999, N5993, N4890, N4144);
buf BUF1 (N6000, N5991);
buf BUF1 (N6001, N5997);
not NOT1 (N6002, N5995);
nor NOR3 (N6003, N5996, N2442, N1267);
and AND2 (N6004, N5988, N4261);
not NOT1 (N6005, N5989);
xor XOR2 (N6006, N6000, N468);
not NOT1 (N6007, N5999);
buf BUF1 (N6008, N6005);
nor NOR2 (N6009, N5980, N5613);
or OR2 (N6010, N6001, N3622);
xor XOR2 (N6011, N6007, N4881);
or OR3 (N6012, N5992, N1640, N3478);
buf BUF1 (N6013, N6009);
nor NOR2 (N6014, N6008, N2182);
or OR4 (N6015, N6004, N5134, N3941, N15);
xor XOR2 (N6016, N6003, N1123);
not NOT1 (N6017, N6014);
nor NOR2 (N6018, N6016, N5827);
nand NAND2 (N6019, N6012, N5895);
and AND2 (N6020, N6015, N1265);
not NOT1 (N6021, N5998);
buf BUF1 (N6022, N6013);
nand NAND4 (N6023, N6011, N5038, N3727, N2995);
and AND2 (N6024, N6020, N2439);
buf BUF1 (N6025, N6024);
xor XOR2 (N6026, N6017, N4585);
not NOT1 (N6027, N6002);
or OR2 (N6028, N6026, N5821);
and AND2 (N6029, N6019, N5274);
or OR4 (N6030, N6029, N3982, N2826, N5719);
nand NAND4 (N6031, N6022, N1137, N4467, N5565);
nor NOR3 (N6032, N6028, N3743, N3661);
buf BUF1 (N6033, N6030);
buf BUF1 (N6034, N6025);
nor NOR4 (N6035, N6033, N1724, N1630, N802);
or OR3 (N6036, N6034, N695, N5214);
and AND3 (N6037, N6018, N935, N800);
nor NOR2 (N6038, N6010, N5646);
buf BUF1 (N6039, N6035);
xor XOR2 (N6040, N6039, N1087);
nor NOR3 (N6041, N6032, N3494, N3679);
or OR4 (N6042, N6031, N1671, N1830, N3815);
xor XOR2 (N6043, N6042, N5823);
and AND2 (N6044, N6027, N3168);
buf BUF1 (N6045, N6036);
xor XOR2 (N6046, N6023, N5345);
buf BUF1 (N6047, N6043);
nand NAND2 (N6048, N6021, N3143);
xor XOR2 (N6049, N6006, N2423);
and AND2 (N6050, N6048, N851);
xor XOR2 (N6051, N6040, N3541);
nor NOR3 (N6052, N6049, N2833, N5699);
or OR2 (N6053, N6047, N469);
not NOT1 (N6054, N6041);
nand NAND2 (N6055, N6046, N844);
or OR3 (N6056, N6054, N5355, N1462);
nand NAND3 (N6057, N6050, N4774, N4554);
not NOT1 (N6058, N6051);
not NOT1 (N6059, N6057);
not NOT1 (N6060, N6056);
nand NAND3 (N6061, N6037, N5089, N3273);
buf BUF1 (N6062, N6060);
buf BUF1 (N6063, N6052);
xor XOR2 (N6064, N6055, N1246);
xor XOR2 (N6065, N6044, N5204);
or OR3 (N6066, N6038, N3243, N2143);
not NOT1 (N6067, N6066);
nand NAND4 (N6068, N6067, N667, N1339, N4021);
xor XOR2 (N6069, N6045, N4734);
or OR4 (N6070, N6063, N1355, N230, N4700);
nor NOR4 (N6071, N6064, N2316, N1674, N1937);
xor XOR2 (N6072, N6062, N4148);
or OR2 (N6073, N6058, N1460);
and AND2 (N6074, N6053, N4748);
nand NAND4 (N6075, N6059, N3489, N1954, N3994);
and AND4 (N6076, N6074, N402, N1031, N58);
xor XOR2 (N6077, N6070, N2827);
nor NOR2 (N6078, N6071, N3654);
or OR2 (N6079, N6068, N4818);
and AND4 (N6080, N6061, N198, N5980, N3642);
or OR4 (N6081, N6065, N6055, N4259, N4987);
buf BUF1 (N6082, N6079);
not NOT1 (N6083, N6082);
and AND3 (N6084, N6083, N898, N3192);
buf BUF1 (N6085, N6075);
not NOT1 (N6086, N6072);
nor NOR3 (N6087, N6085, N4337, N216);
nor NOR3 (N6088, N6069, N4760, N4723);
and AND4 (N6089, N6081, N1587, N3723, N611);
nor NOR3 (N6090, N6080, N5267, N4995);
and AND2 (N6091, N6090, N4312);
xor XOR2 (N6092, N6078, N5793);
and AND4 (N6093, N6087, N2409, N1623, N4947);
buf BUF1 (N6094, N6093);
and AND2 (N6095, N6089, N1384);
not NOT1 (N6096, N6086);
not NOT1 (N6097, N6084);
buf BUF1 (N6098, N6077);
nand NAND2 (N6099, N6098, N1612);
and AND2 (N6100, N6092, N2599);
nor NOR2 (N6101, N6091, N783);
not NOT1 (N6102, N6101);
nand NAND2 (N6103, N6097, N6056);
nand NAND3 (N6104, N6103, N319, N519);
xor XOR2 (N6105, N6095, N4882);
buf BUF1 (N6106, N6104);
nand NAND4 (N6107, N6100, N3158, N1997, N719);
and AND2 (N6108, N6076, N2224);
nand NAND3 (N6109, N6106, N5302, N3904);
not NOT1 (N6110, N6094);
and AND3 (N6111, N6102, N3058, N4933);
nor NOR3 (N6112, N6107, N2642, N5129);
buf BUF1 (N6113, N6108);
nand NAND4 (N6114, N6109, N2416, N510, N434);
and AND4 (N6115, N6099, N5588, N5883, N3155);
xor XOR2 (N6116, N6112, N3326);
or OR4 (N6117, N6113, N400, N4180, N1400);
xor XOR2 (N6118, N6110, N3146);
nor NOR2 (N6119, N6073, N5980);
not NOT1 (N6120, N6088);
or OR2 (N6121, N6111, N1353);
nand NAND2 (N6122, N6114, N4841);
or OR2 (N6123, N6122, N5750);
nor NOR4 (N6124, N6118, N3427, N325, N5299);
or OR3 (N6125, N6116, N3297, N529);
xor XOR2 (N6126, N6117, N3464);
nor NOR4 (N6127, N6124, N5770, N4659, N2738);
not NOT1 (N6128, N6105);
or OR4 (N6129, N6123, N853, N140, N2737);
xor XOR2 (N6130, N6096, N1185);
and AND3 (N6131, N6120, N3380, N4669);
not NOT1 (N6132, N6119);
buf BUF1 (N6133, N6126);
nand NAND3 (N6134, N6132, N3059, N1997);
and AND3 (N6135, N6128, N3379, N9);
buf BUF1 (N6136, N6125);
xor XOR2 (N6137, N6115, N1260);
not NOT1 (N6138, N6135);
xor XOR2 (N6139, N6133, N3512);
xor XOR2 (N6140, N6136, N162);
xor XOR2 (N6141, N6139, N892);
nor NOR2 (N6142, N6141, N1737);
xor XOR2 (N6143, N6138, N2480);
or OR4 (N6144, N6134, N1906, N2386, N4284);
nand NAND2 (N6145, N6144, N3492);
buf BUF1 (N6146, N6129);
or OR3 (N6147, N6146, N4426, N1285);
or OR2 (N6148, N6145, N2552);
or OR3 (N6149, N6147, N5030, N3822);
nand NAND3 (N6150, N6140, N1789, N2232);
not NOT1 (N6151, N6130);
and AND2 (N6152, N6143, N416);
not NOT1 (N6153, N6148);
and AND2 (N6154, N6131, N4459);
or OR3 (N6155, N6149, N5230, N2179);
nor NOR2 (N6156, N6137, N5163);
not NOT1 (N6157, N6156);
or OR2 (N6158, N6157, N5019);
xor XOR2 (N6159, N6121, N597);
or OR3 (N6160, N6142, N5611, N691);
nand NAND2 (N6161, N6155, N1808);
buf BUF1 (N6162, N6153);
xor XOR2 (N6163, N6150, N914);
buf BUF1 (N6164, N6161);
or OR3 (N6165, N6152, N5489, N3037);
xor XOR2 (N6166, N6165, N4842);
and AND4 (N6167, N6158, N3729, N2889, N220);
xor XOR2 (N6168, N6166, N511);
or OR2 (N6169, N6167, N6069);
or OR2 (N6170, N6154, N5527);
nor NOR3 (N6171, N6163, N3882, N2545);
not NOT1 (N6172, N6159);
and AND3 (N6173, N6171, N568, N5190);
not NOT1 (N6174, N6169);
and AND3 (N6175, N6162, N5062, N3373);
nor NOR2 (N6176, N6151, N4785);
and AND2 (N6177, N6127, N1737);
not NOT1 (N6178, N6170);
or OR4 (N6179, N6178, N4354, N5801, N6022);
not NOT1 (N6180, N6177);
and AND4 (N6181, N6179, N6170, N3481, N4914);
buf BUF1 (N6182, N6173);
and AND2 (N6183, N6172, N5610);
or OR2 (N6184, N6183, N1401);
buf BUF1 (N6185, N6182);
nand NAND2 (N6186, N6168, N2710);
and AND4 (N6187, N6164, N98, N3265, N820);
nand NAND2 (N6188, N6185, N6177);
not NOT1 (N6189, N6186);
not NOT1 (N6190, N6189);
buf BUF1 (N6191, N6160);
or OR4 (N6192, N6180, N1370, N1836, N5823);
xor XOR2 (N6193, N6191, N2402);
not NOT1 (N6194, N6174);
nand NAND3 (N6195, N6188, N5499, N609);
nand NAND2 (N6196, N6175, N5522);
or OR4 (N6197, N6192, N5975, N2706, N705);
buf BUF1 (N6198, N6193);
or OR2 (N6199, N6197, N5566);
nand NAND2 (N6200, N6176, N1050);
or OR3 (N6201, N6184, N4050, N719);
buf BUF1 (N6202, N6199);
and AND3 (N6203, N6187, N3474, N5774);
or OR3 (N6204, N6195, N554, N1139);
or OR3 (N6205, N6200, N5527, N2180);
nor NOR2 (N6206, N6203, N321);
buf BUF1 (N6207, N6196);
nor NOR2 (N6208, N6202, N3820);
xor XOR2 (N6209, N6190, N74);
xor XOR2 (N6210, N6209, N76);
and AND4 (N6211, N6207, N1644, N1961, N1961);
not NOT1 (N6212, N6211);
and AND4 (N6213, N6210, N2703, N5015, N3972);
nor NOR4 (N6214, N6205, N5150, N2356, N860);
xor XOR2 (N6215, N6214, N5868);
not NOT1 (N6216, N6181);
nand NAND2 (N6217, N6213, N3216);
buf BUF1 (N6218, N6212);
xor XOR2 (N6219, N6216, N3430);
or OR4 (N6220, N6217, N5855, N3141, N63);
nand NAND3 (N6221, N6208, N5409, N5974);
not NOT1 (N6222, N6194);
buf BUF1 (N6223, N6215);
nand NAND3 (N6224, N6221, N2641, N2241);
buf BUF1 (N6225, N6204);
or OR3 (N6226, N6222, N725, N615);
xor XOR2 (N6227, N6201, N2190);
nand NAND2 (N6228, N6223, N1879);
xor XOR2 (N6229, N6226, N1272);
and AND3 (N6230, N6229, N4798, N4053);
nor NOR2 (N6231, N6206, N1159);
or OR3 (N6232, N6219, N2550, N2936);
nand NAND2 (N6233, N6218, N3426);
not NOT1 (N6234, N6232);
buf BUF1 (N6235, N6227);
nor NOR3 (N6236, N6224, N1216, N4773);
or OR2 (N6237, N6230, N1099);
buf BUF1 (N6238, N6198);
and AND3 (N6239, N6228, N2069, N2288);
buf BUF1 (N6240, N6225);
xor XOR2 (N6241, N6238, N2650);
not NOT1 (N6242, N6240);
not NOT1 (N6243, N6241);
xor XOR2 (N6244, N6236, N5553);
buf BUF1 (N6245, N6244);
and AND2 (N6246, N6234, N580);
not NOT1 (N6247, N6246);
not NOT1 (N6248, N6231);
or OR4 (N6249, N6220, N3906, N328, N2776);
not NOT1 (N6250, N6243);
xor XOR2 (N6251, N6248, N4046);
or OR4 (N6252, N6239, N886, N634, N5773);
nand NAND4 (N6253, N6237, N1798, N1420, N13);
xor XOR2 (N6254, N6252, N3326);
not NOT1 (N6255, N6247);
buf BUF1 (N6256, N6251);
and AND2 (N6257, N6235, N3066);
or OR2 (N6258, N6233, N1782);
nor NOR2 (N6259, N6258, N2420);
xor XOR2 (N6260, N6254, N4649);
nor NOR4 (N6261, N6253, N1165, N4768, N4693);
not NOT1 (N6262, N6261);
not NOT1 (N6263, N6255);
nand NAND2 (N6264, N6256, N198);
nor NOR4 (N6265, N6257, N2367, N68, N2111);
or OR2 (N6266, N6265, N5899);
and AND4 (N6267, N6266, N944, N3178, N2258);
xor XOR2 (N6268, N6259, N4295);
not NOT1 (N6269, N6262);
not NOT1 (N6270, N6268);
nand NAND3 (N6271, N6269, N5168, N5245);
nor NOR3 (N6272, N6245, N2018, N4778);
not NOT1 (N6273, N6263);
not NOT1 (N6274, N6267);
not NOT1 (N6275, N6271);
not NOT1 (N6276, N6272);
xor XOR2 (N6277, N6270, N3044);
nand NAND2 (N6278, N6249, N4727);
and AND3 (N6279, N6274, N4707, N2351);
nand NAND3 (N6280, N6264, N3080, N4556);
or OR3 (N6281, N6277, N4541, N5431);
nand NAND3 (N6282, N6276, N4969, N4886);
buf BUF1 (N6283, N6280);
buf BUF1 (N6284, N6279);
nand NAND2 (N6285, N6283, N1308);
xor XOR2 (N6286, N6281, N1478);
nor NOR4 (N6287, N6282, N1056, N4151, N2227);
and AND4 (N6288, N6284, N5405, N5350, N3071);
nor NOR2 (N6289, N6287, N2771);
xor XOR2 (N6290, N6275, N5516);
nor NOR4 (N6291, N6290, N3759, N3448, N3331);
nor NOR2 (N6292, N6242, N3547);
nor NOR4 (N6293, N6292, N2781, N2056, N3602);
or OR3 (N6294, N6285, N2868, N3302);
buf BUF1 (N6295, N6286);
not NOT1 (N6296, N6250);
nand NAND4 (N6297, N6260, N3588, N1256, N4586);
nand NAND4 (N6298, N6295, N3823, N5573, N1456);
xor XOR2 (N6299, N6297, N4226);
xor XOR2 (N6300, N6299, N5214);
nand NAND2 (N6301, N6298, N3452);
buf BUF1 (N6302, N6288);
and AND4 (N6303, N6296, N4027, N1355, N1957);
nor NOR2 (N6304, N6289, N4706);
not NOT1 (N6305, N6293);
xor XOR2 (N6306, N6304, N2238);
buf BUF1 (N6307, N6303);
buf BUF1 (N6308, N6291);
nand NAND2 (N6309, N6294, N1363);
and AND2 (N6310, N6302, N2677);
not NOT1 (N6311, N6310);
not NOT1 (N6312, N6306);
nand NAND4 (N6313, N6300, N3717, N5331, N2030);
nand NAND3 (N6314, N6308, N934, N2930);
not NOT1 (N6315, N6305);
nand NAND3 (N6316, N6312, N277, N3502);
and AND4 (N6317, N6273, N4058, N1960, N4223);
or OR2 (N6318, N6278, N3747);
xor XOR2 (N6319, N6315, N1738);
not NOT1 (N6320, N6317);
nor NOR2 (N6321, N6313, N3986);
nand NAND4 (N6322, N6316, N5042, N879, N1980);
not NOT1 (N6323, N6311);
nand NAND3 (N6324, N6314, N4335, N3497);
buf BUF1 (N6325, N6321);
buf BUF1 (N6326, N6318);
not NOT1 (N6327, N6323);
xor XOR2 (N6328, N6307, N6149);
xor XOR2 (N6329, N6324, N6246);
nand NAND3 (N6330, N6322, N4667, N1584);
nor NOR2 (N6331, N6330, N4885);
nor NOR4 (N6332, N6309, N3234, N248, N2920);
xor XOR2 (N6333, N6332, N5320);
nor NOR2 (N6334, N6328, N3062);
buf BUF1 (N6335, N6326);
or OR2 (N6336, N6335, N4962);
buf BUF1 (N6337, N6301);
nor NOR3 (N6338, N6336, N4002, N180);
buf BUF1 (N6339, N6334);
and AND4 (N6340, N6329, N5640, N3083, N5916);
buf BUF1 (N6341, N6337);
or OR3 (N6342, N6325, N567, N701);
and AND2 (N6343, N6341, N2811);
not NOT1 (N6344, N6342);
or OR4 (N6345, N6319, N4612, N3113, N2888);
and AND3 (N6346, N6320, N1976, N3125);
buf BUF1 (N6347, N6339);
nand NAND4 (N6348, N6346, N1610, N2906, N32);
buf BUF1 (N6349, N6347);
nand NAND3 (N6350, N6333, N6239, N2941);
buf BUF1 (N6351, N6340);
and AND2 (N6352, N6343, N438);
buf BUF1 (N6353, N6327);
not NOT1 (N6354, N6348);
not NOT1 (N6355, N6353);
and AND3 (N6356, N6352, N727, N3254);
or OR2 (N6357, N6345, N16);
not NOT1 (N6358, N6350);
not NOT1 (N6359, N6354);
buf BUF1 (N6360, N6359);
xor XOR2 (N6361, N6357, N2515);
not NOT1 (N6362, N6361);
not NOT1 (N6363, N6360);
xor XOR2 (N6364, N6356, N5451);
not NOT1 (N6365, N6364);
not NOT1 (N6366, N6362);
nor NOR3 (N6367, N6366, N6216, N2968);
and AND3 (N6368, N6363, N639, N4550);
and AND2 (N6369, N6367, N1191);
xor XOR2 (N6370, N6368, N4904);
or OR2 (N6371, N6349, N2276);
buf BUF1 (N6372, N6338);
xor XOR2 (N6373, N6371, N2633);
and AND4 (N6374, N6344, N5842, N2062, N427);
xor XOR2 (N6375, N6369, N205);
or OR2 (N6376, N6373, N4517);
xor XOR2 (N6377, N6355, N365);
or OR3 (N6378, N6372, N5055, N4984);
nand NAND4 (N6379, N6378, N6311, N5778, N3847);
xor XOR2 (N6380, N6375, N5250);
nand NAND2 (N6381, N6377, N4300);
nor NOR4 (N6382, N6381, N555, N177, N2848);
or OR2 (N6383, N6351, N5644);
and AND4 (N6384, N6358, N6254, N1965, N5341);
buf BUF1 (N6385, N6370);
xor XOR2 (N6386, N6384, N1246);
nor NOR2 (N6387, N6379, N2852);
or OR4 (N6388, N6382, N5319, N5600, N6125);
not NOT1 (N6389, N6387);
not NOT1 (N6390, N6388);
not NOT1 (N6391, N6389);
and AND2 (N6392, N6365, N4276);
nor NOR4 (N6393, N6380, N5029, N1676, N3302);
or OR4 (N6394, N6385, N3663, N6184, N950);
or OR4 (N6395, N6374, N4187, N4459, N498);
xor XOR2 (N6396, N6376, N2572);
buf BUF1 (N6397, N6391);
nor NOR2 (N6398, N6386, N3759);
or OR2 (N6399, N6390, N5445);
not NOT1 (N6400, N6398);
xor XOR2 (N6401, N6331, N4385);
and AND3 (N6402, N6394, N2266, N4624);
buf BUF1 (N6403, N6395);
nand NAND2 (N6404, N6393, N3346);
nand NAND2 (N6405, N6402, N3587);
not NOT1 (N6406, N6396);
nor NOR3 (N6407, N6404, N5841, N2291);
or OR2 (N6408, N6397, N4435);
or OR3 (N6409, N6392, N2118, N2288);
and AND3 (N6410, N6408, N5774, N5546);
or OR4 (N6411, N6407, N3209, N5303, N1976);
or OR4 (N6412, N6400, N507, N487, N2323);
nor NOR4 (N6413, N6411, N1630, N4880, N4027);
nor NOR4 (N6414, N6383, N556, N88, N291);
xor XOR2 (N6415, N6413, N4349);
not NOT1 (N6416, N6410);
nand NAND3 (N6417, N6399, N4354, N217);
or OR3 (N6418, N6403, N2078, N6350);
nor NOR4 (N6419, N6401, N2074, N949, N1198);
xor XOR2 (N6420, N6415, N1834);
nand NAND4 (N6421, N6417, N5493, N2928, N2148);
endmodule