// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N2010,N2007,N2003,N2012,N1989,N2006,N2011,N2000,N2009,N2013;

buf BUF1 (N14, N6);
xor XOR2 (N15, N6, N6);
nor NOR3 (N16, N11, N14, N3);
not NOT1 (N17, N10);
and AND4 (N18, N3, N2, N11, N13);
nor NOR2 (N19, N7, N2);
buf BUF1 (N20, N5);
buf BUF1 (N21, N7);
or OR3 (N22, N6, N8, N21);
or OR4 (N23, N1, N4, N17, N9);
or OR2 (N24, N15, N4);
and AND4 (N25, N18, N4, N24, N20);
xor XOR2 (N26, N12, N16);
or OR2 (N27, N19, N2);
nor NOR3 (N28, N10, N27, N23);
and AND3 (N29, N11, N27, N4);
xor XOR2 (N30, N9, N10);
and AND4 (N31, N9, N27, N6, N22);
nor NOR2 (N32, N11, N17);
xor XOR2 (N33, N17, N9);
nand NAND3 (N34, N15, N12, N15);
nor NOR4 (N35, N32, N16, N6, N9);
nand NAND4 (N36, N12, N13, N26, N8);
nand NAND4 (N37, N16, N29, N26, N13);
nand NAND3 (N38, N5, N14, N30);
not NOT1 (N39, N32);
buf BUF1 (N40, N33);
nand NAND4 (N41, N40, N33, N21, N20);
and AND3 (N42, N41, N20, N21);
xor XOR2 (N43, N37, N39);
xor XOR2 (N44, N8, N41);
nand NAND4 (N45, N34, N3, N30, N4);
nor NOR2 (N46, N36, N18);
or OR4 (N47, N43, N37, N10, N41);
xor XOR2 (N48, N42, N5);
buf BUF1 (N49, N31);
and AND2 (N50, N47, N34);
and AND4 (N51, N35, N24, N33, N28);
nand NAND4 (N52, N15, N34, N30, N19);
xor XOR2 (N53, N51, N33);
xor XOR2 (N54, N49, N40);
not NOT1 (N55, N45);
not NOT1 (N56, N55);
and AND4 (N57, N56, N13, N54, N32);
or OR4 (N58, N6, N31, N30, N22);
nor NOR4 (N59, N38, N2, N47, N39);
xor XOR2 (N60, N59, N1);
nand NAND3 (N61, N50, N16, N1);
not NOT1 (N62, N46);
and AND4 (N63, N48, N17, N41, N14);
xor XOR2 (N64, N61, N29);
nor NOR2 (N65, N44, N28);
not NOT1 (N66, N62);
buf BUF1 (N67, N66);
and AND2 (N68, N58, N7);
buf BUF1 (N69, N57);
nor NOR2 (N70, N65, N56);
nor NOR2 (N71, N68, N63);
buf BUF1 (N72, N17);
nand NAND3 (N73, N71, N23, N19);
buf BUF1 (N74, N25);
and AND4 (N75, N52, N34, N28, N72);
xor XOR2 (N76, N1, N22);
nand NAND4 (N77, N75, N53, N23, N56);
not NOT1 (N78, N55);
nand NAND3 (N79, N70, N39, N56);
not NOT1 (N80, N74);
or OR4 (N81, N79, N52, N18, N7);
nand NAND2 (N82, N80, N12);
nand NAND4 (N83, N82, N2, N44, N43);
nand NAND3 (N84, N64, N57, N55);
not NOT1 (N85, N60);
buf BUF1 (N86, N73);
or OR3 (N87, N76, N31, N40);
and AND4 (N88, N78, N39, N65, N69);
or OR4 (N89, N40, N21, N4, N26);
xor XOR2 (N90, N81, N60);
or OR3 (N91, N85, N74, N23);
buf BUF1 (N92, N91);
xor XOR2 (N93, N77, N91);
not NOT1 (N94, N89);
xor XOR2 (N95, N84, N20);
nor NOR2 (N96, N67, N82);
or OR3 (N97, N83, N37, N16);
nor NOR3 (N98, N96, N8, N29);
or OR3 (N99, N98, N24, N4);
xor XOR2 (N100, N87, N45);
nand NAND4 (N101, N90, N8, N9, N13);
not NOT1 (N102, N86);
nand NAND3 (N103, N88, N101, N98);
nand NAND3 (N104, N39, N32, N40);
not NOT1 (N105, N94);
nor NOR2 (N106, N100, N35);
xor XOR2 (N107, N99, N20);
nor NOR3 (N108, N92, N7, N65);
xor XOR2 (N109, N102, N45);
nand NAND2 (N110, N103, N56);
nand NAND2 (N111, N107, N44);
nor NOR2 (N112, N104, N90);
and AND4 (N113, N93, N59, N95, N50);
xor XOR2 (N114, N110, N23);
nand NAND4 (N115, N60, N30, N54, N83);
buf BUF1 (N116, N97);
nor NOR4 (N117, N111, N71, N50, N94);
and AND2 (N118, N109, N100);
and AND4 (N119, N106, N64, N32, N29);
nand NAND2 (N120, N115, N87);
buf BUF1 (N121, N116);
not NOT1 (N122, N105);
and AND4 (N123, N119, N40, N16, N108);
buf BUF1 (N124, N22);
not NOT1 (N125, N117);
nor NOR3 (N126, N113, N19, N114);
xor XOR2 (N127, N35, N35);
or OR4 (N128, N125, N45, N119, N102);
xor XOR2 (N129, N122, N68);
buf BUF1 (N130, N127);
buf BUF1 (N131, N130);
or OR3 (N132, N118, N17, N32);
nand NAND3 (N133, N129, N9, N61);
xor XOR2 (N134, N124, N67);
and AND2 (N135, N134, N50);
or OR3 (N136, N120, N5, N83);
not NOT1 (N137, N112);
and AND4 (N138, N135, N81, N22, N66);
not NOT1 (N139, N131);
not NOT1 (N140, N121);
not NOT1 (N141, N123);
and AND4 (N142, N126, N88, N74, N87);
or OR2 (N143, N141, N76);
buf BUF1 (N144, N139);
nand NAND3 (N145, N132, N75, N57);
not NOT1 (N146, N133);
xor XOR2 (N147, N138, N45);
or OR3 (N148, N140, N90, N79);
not NOT1 (N149, N137);
and AND3 (N150, N142, N132, N89);
buf BUF1 (N151, N146);
nand NAND4 (N152, N128, N26, N103, N3);
and AND3 (N153, N149, N101, N124);
not NOT1 (N154, N147);
or OR2 (N155, N145, N97);
buf BUF1 (N156, N154);
buf BUF1 (N157, N143);
nor NOR4 (N158, N157, N79, N101, N65);
buf BUF1 (N159, N150);
nand NAND4 (N160, N156, N104, N117, N113);
or OR2 (N161, N151, N135);
nor NOR3 (N162, N161, N72, N11);
nor NOR2 (N163, N152, N144);
nor NOR3 (N164, N91, N80, N62);
buf BUF1 (N165, N153);
nor NOR2 (N166, N165, N120);
buf BUF1 (N167, N162);
nand NAND2 (N168, N136, N35);
xor XOR2 (N169, N166, N17);
or OR4 (N170, N168, N106, N91, N61);
not NOT1 (N171, N160);
xor XOR2 (N172, N169, N57);
or OR4 (N173, N167, N164, N16, N100);
buf BUF1 (N174, N127);
or OR3 (N175, N173, N105, N117);
nand NAND2 (N176, N163, N116);
nor NOR3 (N177, N159, N76, N141);
xor XOR2 (N178, N172, N64);
not NOT1 (N179, N148);
or OR2 (N180, N177, N20);
not NOT1 (N181, N176);
or OR3 (N182, N180, N154, N168);
xor XOR2 (N183, N181, N143);
nor NOR3 (N184, N158, N108, N10);
buf BUF1 (N185, N155);
or OR2 (N186, N182, N113);
and AND3 (N187, N184, N17, N140);
nand NAND2 (N188, N174, N4);
or OR3 (N189, N188, N7, N16);
nand NAND4 (N190, N175, N154, N115, N138);
nor NOR2 (N191, N187, N81);
nand NAND2 (N192, N186, N59);
nor NOR3 (N193, N185, N157, N143);
not NOT1 (N194, N178);
xor XOR2 (N195, N191, N21);
buf BUF1 (N196, N195);
buf BUF1 (N197, N183);
buf BUF1 (N198, N170);
nand NAND3 (N199, N196, N159, N130);
buf BUF1 (N200, N197);
nand NAND3 (N201, N189, N19, N168);
or OR2 (N202, N190, N58);
xor XOR2 (N203, N202, N13);
or OR2 (N204, N192, N194);
not NOT1 (N205, N133);
or OR4 (N206, N193, N117, N56, N7);
or OR3 (N207, N203, N166, N152);
and AND4 (N208, N205, N121, N52, N120);
nor NOR3 (N209, N198, N123, N146);
nand NAND2 (N210, N179, N76);
xor XOR2 (N211, N171, N40);
not NOT1 (N212, N204);
buf BUF1 (N213, N201);
and AND4 (N214, N209, N61, N87, N141);
buf BUF1 (N215, N212);
nand NAND3 (N216, N200, N175, N72);
not NOT1 (N217, N207);
nor NOR3 (N218, N208, N8, N133);
xor XOR2 (N219, N218, N158);
not NOT1 (N220, N216);
not NOT1 (N221, N215);
nand NAND2 (N222, N211, N68);
or OR4 (N223, N222, N1, N40, N24);
xor XOR2 (N224, N221, N195);
and AND3 (N225, N213, N8, N95);
xor XOR2 (N226, N219, N96);
or OR4 (N227, N223, N111, N184, N51);
nand NAND2 (N228, N225, N10);
nand NAND4 (N229, N206, N45, N177, N49);
or OR2 (N230, N210, N13);
nand NAND3 (N231, N227, N52, N59);
nor NOR4 (N232, N230, N116, N216, N152);
not NOT1 (N233, N217);
and AND4 (N234, N199, N60, N171, N192);
xor XOR2 (N235, N214, N90);
or OR3 (N236, N228, N207, N57);
and AND3 (N237, N224, N173, N189);
buf BUF1 (N238, N236);
or OR3 (N239, N237, N159, N211);
or OR4 (N240, N233, N186, N92, N55);
nand NAND4 (N241, N226, N57, N16, N16);
nor NOR2 (N242, N229, N11);
buf BUF1 (N243, N239);
buf BUF1 (N244, N242);
xor XOR2 (N245, N238, N114);
not NOT1 (N246, N243);
not NOT1 (N247, N245);
or OR3 (N248, N220, N247, N32);
buf BUF1 (N249, N122);
and AND4 (N250, N235, N8, N240, N73);
not NOT1 (N251, N212);
buf BUF1 (N252, N249);
nor NOR3 (N253, N244, N183, N83);
xor XOR2 (N254, N253, N7);
and AND3 (N255, N232, N224, N113);
or OR2 (N256, N231, N189);
and AND3 (N257, N252, N137, N33);
nor NOR3 (N258, N257, N6, N143);
or OR2 (N259, N250, N197);
xor XOR2 (N260, N258, N21);
nor NOR4 (N261, N234, N84, N155, N137);
nand NAND3 (N262, N260, N151, N102);
buf BUF1 (N263, N256);
nand NAND2 (N264, N259, N225);
not NOT1 (N265, N246);
nor NOR3 (N266, N248, N181, N112);
nor NOR3 (N267, N265, N101, N165);
nand NAND3 (N268, N266, N131, N262);
buf BUF1 (N269, N220);
nor NOR2 (N270, N263, N99);
nor NOR4 (N271, N268, N76, N125, N168);
nand NAND4 (N272, N264, N245, N154, N192);
buf BUF1 (N273, N254);
nor NOR4 (N274, N269, N91, N39, N205);
or OR2 (N275, N271, N126);
nor NOR2 (N276, N241, N57);
nand NAND3 (N277, N261, N172, N102);
not NOT1 (N278, N267);
and AND3 (N279, N251, N62, N247);
xor XOR2 (N280, N277, N153);
and AND4 (N281, N276, N3, N265, N87);
nor NOR2 (N282, N279, N79);
nand NAND2 (N283, N278, N229);
buf BUF1 (N284, N275);
or OR4 (N285, N274, N143, N219, N161);
and AND4 (N286, N283, N49, N156, N251);
or OR3 (N287, N272, N247, N148);
nor NOR2 (N288, N284, N148);
nor NOR3 (N289, N255, N244, N198);
nor NOR2 (N290, N281, N254);
and AND2 (N291, N282, N109);
nand NAND4 (N292, N291, N12, N66, N3);
nand NAND4 (N293, N288, N117, N198, N287);
xor XOR2 (N294, N282, N277);
nor NOR4 (N295, N290, N276, N242, N129);
buf BUF1 (N296, N293);
nand NAND4 (N297, N296, N31, N258, N117);
buf BUF1 (N298, N297);
nor NOR2 (N299, N295, N85);
nor NOR4 (N300, N292, N235, N52, N54);
and AND4 (N301, N298, N290, N67, N274);
buf BUF1 (N302, N299);
nor NOR2 (N303, N273, N62);
nand NAND3 (N304, N300, N219, N82);
nor NOR3 (N305, N285, N181, N113);
buf BUF1 (N306, N303);
nor NOR4 (N307, N306, N269, N102, N242);
and AND4 (N308, N270, N127, N10, N306);
xor XOR2 (N309, N286, N100);
buf BUF1 (N310, N302);
or OR4 (N311, N280, N32, N9, N294);
nand NAND2 (N312, N91, N127);
buf BUF1 (N313, N304);
nand NAND2 (N314, N308, N150);
nand NAND4 (N315, N314, N232, N174, N308);
not NOT1 (N316, N313);
xor XOR2 (N317, N289, N254);
or OR3 (N318, N305, N231, N226);
or OR4 (N319, N310, N40, N317, N110);
and AND4 (N320, N230, N290, N248, N313);
nand NAND4 (N321, N315, N122, N60, N307);
nand NAND3 (N322, N155, N116, N276);
nand NAND3 (N323, N318, N81, N297);
nor NOR3 (N324, N321, N71, N281);
nand NAND4 (N325, N320, N52, N76, N251);
nor NOR2 (N326, N325, N12);
nand NAND2 (N327, N316, N8);
xor XOR2 (N328, N324, N216);
not NOT1 (N329, N322);
and AND3 (N330, N312, N126, N109);
buf BUF1 (N331, N311);
xor XOR2 (N332, N301, N7);
nand NAND2 (N333, N331, N254);
or OR2 (N334, N329, N32);
nor NOR2 (N335, N332, N52);
and AND2 (N336, N333, N163);
nor NOR2 (N337, N328, N277);
and AND3 (N338, N309, N280, N272);
nor NOR3 (N339, N338, N136, N38);
buf BUF1 (N340, N330);
nand NAND3 (N341, N337, N145, N237);
or OR4 (N342, N336, N105, N174, N177);
xor XOR2 (N343, N341, N323);
buf BUF1 (N344, N316);
nand NAND2 (N345, N340, N218);
not NOT1 (N346, N343);
or OR3 (N347, N326, N195, N208);
xor XOR2 (N348, N342, N289);
nand NAND2 (N349, N345, N213);
buf BUF1 (N350, N347);
not NOT1 (N351, N348);
not NOT1 (N352, N349);
nor NOR3 (N353, N346, N161, N263);
nand NAND3 (N354, N335, N247, N9);
buf BUF1 (N355, N353);
nand NAND2 (N356, N355, N326);
or OR3 (N357, N334, N57, N235);
xor XOR2 (N358, N351, N164);
nand NAND2 (N359, N356, N155);
not NOT1 (N360, N327);
not NOT1 (N361, N339);
nor NOR3 (N362, N319, N194, N34);
and AND4 (N363, N361, N362, N68, N56);
and AND3 (N364, N349, N27, N53);
buf BUF1 (N365, N363);
nor NOR2 (N366, N352, N177);
nor NOR2 (N367, N357, N269);
not NOT1 (N368, N359);
nand NAND4 (N369, N350, N232, N217, N156);
buf BUF1 (N370, N360);
buf BUF1 (N371, N368);
xor XOR2 (N372, N344, N37);
xor XOR2 (N373, N354, N66);
nand NAND4 (N374, N369, N100, N236, N176);
nor NOR2 (N375, N372, N1);
nor NOR4 (N376, N371, N292, N133, N306);
xor XOR2 (N377, N375, N40);
xor XOR2 (N378, N358, N369);
not NOT1 (N379, N370);
not NOT1 (N380, N373);
or OR3 (N381, N380, N220, N252);
and AND3 (N382, N365, N118, N160);
nand NAND4 (N383, N377, N221, N272, N32);
or OR4 (N384, N378, N34, N224, N346);
xor XOR2 (N385, N384, N167);
not NOT1 (N386, N367);
nor NOR3 (N387, N381, N249, N119);
or OR3 (N388, N383, N365, N253);
buf BUF1 (N389, N382);
and AND4 (N390, N364, N277, N28, N169);
and AND4 (N391, N388, N332, N179, N186);
and AND3 (N392, N387, N201, N343);
and AND4 (N393, N385, N123, N296, N342);
xor XOR2 (N394, N389, N30);
not NOT1 (N395, N379);
or OR3 (N396, N390, N5, N283);
not NOT1 (N397, N394);
xor XOR2 (N398, N386, N128);
or OR4 (N399, N398, N217, N290, N36);
buf BUF1 (N400, N392);
and AND3 (N401, N399, N278, N244);
xor XOR2 (N402, N400, N314);
nor NOR2 (N403, N391, N374);
and AND4 (N404, N180, N130, N167, N275);
nor NOR2 (N405, N397, N165);
nand NAND3 (N406, N393, N40, N227);
xor XOR2 (N407, N404, N209);
buf BUF1 (N408, N405);
or OR4 (N409, N401, N325, N350, N196);
not NOT1 (N410, N406);
nor NOR4 (N411, N409, N82, N180, N174);
or OR2 (N412, N403, N314);
nor NOR4 (N413, N395, N147, N155, N125);
and AND3 (N414, N408, N16, N27);
and AND2 (N415, N407, N34);
and AND4 (N416, N402, N144, N176, N119);
and AND2 (N417, N413, N219);
or OR4 (N418, N396, N282, N192, N320);
buf BUF1 (N419, N416);
nand NAND3 (N420, N366, N354, N303);
and AND2 (N421, N412, N165);
not NOT1 (N422, N417);
nand NAND4 (N423, N376, N333, N223, N291);
or OR3 (N424, N422, N227, N351);
nor NOR3 (N425, N424, N301, N73);
nor NOR3 (N426, N411, N124, N135);
or OR2 (N427, N423, N409);
xor XOR2 (N428, N415, N190);
and AND3 (N429, N410, N327, N227);
xor XOR2 (N430, N414, N157);
nor NOR4 (N431, N418, N225, N295, N240);
nand NAND3 (N432, N425, N59, N340);
nor NOR3 (N433, N428, N138, N289);
not NOT1 (N434, N426);
buf BUF1 (N435, N421);
and AND3 (N436, N420, N425, N71);
buf BUF1 (N437, N430);
and AND3 (N438, N436, N125, N62);
or OR3 (N439, N431, N45, N296);
xor XOR2 (N440, N435, N112);
and AND2 (N441, N438, N242);
xor XOR2 (N442, N441, N26);
xor XOR2 (N443, N439, N323);
or OR4 (N444, N442, N155, N382, N233);
xor XOR2 (N445, N437, N227);
buf BUF1 (N446, N429);
nor NOR4 (N447, N434, N218, N374, N328);
buf BUF1 (N448, N419);
xor XOR2 (N449, N445, N22);
and AND4 (N450, N433, N84, N278, N229);
nand NAND3 (N451, N449, N365, N83);
and AND2 (N452, N427, N203);
nand NAND3 (N453, N440, N372, N400);
and AND4 (N454, N451, N385, N161, N180);
buf BUF1 (N455, N454);
buf BUF1 (N456, N455);
nor NOR2 (N457, N432, N156);
nand NAND4 (N458, N457, N162, N7, N245);
buf BUF1 (N459, N447);
xor XOR2 (N460, N458, N94);
nand NAND4 (N461, N460, N355, N83, N347);
nor NOR3 (N462, N443, N144, N207);
or OR3 (N463, N444, N216, N8);
buf BUF1 (N464, N452);
and AND2 (N465, N453, N327);
nor NOR2 (N466, N450, N22);
nand NAND2 (N467, N456, N54);
and AND2 (N468, N461, N181);
and AND4 (N469, N459, N426, N237, N185);
nand NAND2 (N470, N465, N120);
nor NOR4 (N471, N468, N315, N428, N221);
nor NOR3 (N472, N469, N32, N169);
xor XOR2 (N473, N470, N114);
or OR3 (N474, N472, N183, N274);
nor NOR2 (N475, N467, N181);
not NOT1 (N476, N446);
and AND2 (N477, N448, N234);
nand NAND3 (N478, N475, N1, N223);
nor NOR2 (N479, N471, N365);
not NOT1 (N480, N466);
not NOT1 (N481, N479);
buf BUF1 (N482, N476);
or OR2 (N483, N462, N451);
xor XOR2 (N484, N480, N248);
nand NAND2 (N485, N483, N191);
nor NOR4 (N486, N484, N45, N70, N240);
nand NAND2 (N487, N477, N33);
and AND3 (N488, N482, N164, N362);
and AND4 (N489, N486, N281, N193, N356);
or OR2 (N490, N488, N446);
not NOT1 (N491, N489);
nand NAND4 (N492, N485, N476, N238, N387);
xor XOR2 (N493, N473, N248);
or OR3 (N494, N490, N108, N91);
nor NOR2 (N495, N474, N144);
buf BUF1 (N496, N481);
and AND4 (N497, N464, N387, N377, N449);
or OR2 (N498, N492, N283);
and AND3 (N499, N498, N306, N470);
and AND4 (N500, N496, N401, N453, N304);
xor XOR2 (N501, N500, N66);
buf BUF1 (N502, N493);
buf BUF1 (N503, N494);
xor XOR2 (N504, N502, N238);
buf BUF1 (N505, N487);
xor XOR2 (N506, N491, N23);
xor XOR2 (N507, N478, N450);
buf BUF1 (N508, N506);
not NOT1 (N509, N508);
nor NOR3 (N510, N499, N247, N300);
or OR2 (N511, N509, N48);
or OR3 (N512, N507, N23, N499);
buf BUF1 (N513, N510);
xor XOR2 (N514, N503, N396);
buf BUF1 (N515, N495);
nand NAND4 (N516, N515, N437, N229, N174);
and AND2 (N517, N516, N490);
and AND4 (N518, N511, N419, N491, N204);
nand NAND2 (N519, N501, N412);
buf BUF1 (N520, N504);
not NOT1 (N521, N463);
xor XOR2 (N522, N513, N142);
and AND3 (N523, N518, N427, N323);
not NOT1 (N524, N512);
xor XOR2 (N525, N522, N338);
buf BUF1 (N526, N523);
buf BUF1 (N527, N505);
nand NAND2 (N528, N497, N75);
nor NOR3 (N529, N526, N486, N81);
nand NAND2 (N530, N527, N106);
and AND4 (N531, N524, N342, N438, N126);
nor NOR4 (N532, N521, N473, N412, N393);
buf BUF1 (N533, N528);
not NOT1 (N534, N532);
nand NAND3 (N535, N534, N43, N232);
or OR2 (N536, N525, N463);
xor XOR2 (N537, N535, N471);
nand NAND2 (N538, N533, N344);
not NOT1 (N539, N538);
nor NOR2 (N540, N536, N165);
not NOT1 (N541, N520);
and AND2 (N542, N519, N218);
nor NOR2 (N543, N514, N379);
buf BUF1 (N544, N537);
and AND2 (N545, N531, N92);
buf BUF1 (N546, N542);
or OR4 (N547, N517, N443, N157, N543);
xor XOR2 (N548, N539, N485);
nand NAND2 (N549, N170, N295);
nand NAND2 (N550, N544, N448);
or OR2 (N551, N529, N32);
nor NOR3 (N552, N547, N53, N18);
xor XOR2 (N553, N541, N334);
not NOT1 (N554, N549);
not NOT1 (N555, N530);
xor XOR2 (N556, N546, N480);
and AND2 (N557, N550, N316);
xor XOR2 (N558, N551, N413);
or OR4 (N559, N554, N282, N147, N173);
nand NAND3 (N560, N557, N291, N460);
or OR2 (N561, N556, N298);
and AND4 (N562, N540, N260, N354, N365);
xor XOR2 (N563, N555, N291);
buf BUF1 (N564, N563);
nor NOR2 (N565, N561, N53);
xor XOR2 (N566, N560, N337);
and AND3 (N567, N564, N283, N170);
xor XOR2 (N568, N558, N100);
not NOT1 (N569, N553);
and AND4 (N570, N559, N220, N108, N7);
xor XOR2 (N571, N568, N271);
or OR2 (N572, N567, N353);
and AND3 (N573, N565, N387, N129);
and AND2 (N574, N552, N317);
buf BUF1 (N575, N545);
xor XOR2 (N576, N569, N9);
buf BUF1 (N577, N572);
xor XOR2 (N578, N566, N451);
buf BUF1 (N579, N571);
or OR3 (N580, N578, N50, N473);
not NOT1 (N581, N575);
nand NAND3 (N582, N580, N561, N259);
nor NOR4 (N583, N581, N499, N491, N322);
nor NOR2 (N584, N579, N489);
buf BUF1 (N585, N582);
nor NOR4 (N586, N573, N350, N133, N42);
nor NOR2 (N587, N585, N439);
buf BUF1 (N588, N570);
nand NAND2 (N589, N588, N403);
xor XOR2 (N590, N589, N192);
buf BUF1 (N591, N562);
xor XOR2 (N592, N576, N191);
not NOT1 (N593, N590);
buf BUF1 (N594, N583);
not NOT1 (N595, N587);
buf BUF1 (N596, N594);
buf BUF1 (N597, N574);
not NOT1 (N598, N548);
xor XOR2 (N599, N595, N4);
xor XOR2 (N600, N584, N578);
buf BUF1 (N601, N593);
nand NAND2 (N602, N577, N373);
nor NOR2 (N603, N601, N369);
xor XOR2 (N604, N597, N274);
xor XOR2 (N605, N596, N416);
nor NOR2 (N606, N586, N150);
or OR3 (N607, N604, N57, N122);
and AND2 (N608, N607, N535);
nand NAND2 (N609, N602, N415);
buf BUF1 (N610, N609);
nand NAND2 (N611, N591, N378);
xor XOR2 (N612, N605, N440);
buf BUF1 (N613, N610);
xor XOR2 (N614, N608, N103);
and AND2 (N615, N613, N57);
xor XOR2 (N616, N606, N68);
buf BUF1 (N617, N614);
buf BUF1 (N618, N598);
or OR2 (N619, N603, N379);
or OR2 (N620, N616, N442);
nand NAND2 (N621, N617, N25);
nand NAND2 (N622, N620, N595);
xor XOR2 (N623, N621, N338);
not NOT1 (N624, N611);
buf BUF1 (N625, N612);
nor NOR2 (N626, N619, N470);
not NOT1 (N627, N600);
buf BUF1 (N628, N626);
xor XOR2 (N629, N622, N98);
nand NAND4 (N630, N624, N593, N52, N431);
and AND3 (N631, N628, N72, N407);
xor XOR2 (N632, N599, N530);
buf BUF1 (N633, N632);
and AND4 (N634, N627, N616, N600, N12);
not NOT1 (N635, N625);
buf BUF1 (N636, N631);
xor XOR2 (N637, N615, N158);
buf BUF1 (N638, N634);
buf BUF1 (N639, N637);
and AND2 (N640, N629, N509);
or OR3 (N641, N633, N11, N494);
nor NOR4 (N642, N592, N434, N440, N34);
or OR4 (N643, N638, N34, N321, N223);
not NOT1 (N644, N641);
buf BUF1 (N645, N635);
nand NAND4 (N646, N640, N499, N23, N473);
and AND4 (N647, N643, N562, N55, N230);
nand NAND2 (N648, N645, N405);
or OR4 (N649, N630, N589, N308, N224);
nand NAND2 (N650, N649, N300);
nor NOR2 (N651, N636, N338);
nor NOR2 (N652, N648, N389);
xor XOR2 (N653, N644, N433);
xor XOR2 (N654, N652, N616);
not NOT1 (N655, N653);
xor XOR2 (N656, N647, N187);
xor XOR2 (N657, N639, N67);
and AND3 (N658, N642, N406, N100);
xor XOR2 (N659, N655, N139);
not NOT1 (N660, N656);
nor NOR2 (N661, N654, N336);
or OR4 (N662, N658, N53, N346, N434);
and AND4 (N663, N646, N580, N442, N240);
not NOT1 (N664, N661);
not NOT1 (N665, N623);
or OR2 (N666, N665, N39);
xor XOR2 (N667, N650, N317);
and AND4 (N668, N657, N345, N492, N421);
or OR3 (N669, N668, N308, N452);
nor NOR3 (N670, N669, N311, N510);
not NOT1 (N671, N666);
nor NOR2 (N672, N651, N548);
and AND4 (N673, N672, N21, N414, N279);
nor NOR4 (N674, N660, N55, N83, N660);
and AND4 (N675, N663, N228, N259, N514);
and AND3 (N676, N674, N129, N186);
buf BUF1 (N677, N671);
nor NOR2 (N678, N667, N134);
or OR2 (N679, N664, N106);
buf BUF1 (N680, N618);
xor XOR2 (N681, N678, N132);
nand NAND3 (N682, N659, N445, N404);
not NOT1 (N683, N670);
and AND4 (N684, N681, N565, N430, N211);
or OR4 (N685, N677, N197, N427, N611);
nand NAND3 (N686, N680, N159, N272);
not NOT1 (N687, N676);
buf BUF1 (N688, N686);
and AND4 (N689, N679, N97, N332, N8);
and AND2 (N690, N688, N499);
nand NAND4 (N691, N687, N330, N434, N173);
nand NAND3 (N692, N689, N429, N551);
nand NAND2 (N693, N684, N141);
not NOT1 (N694, N683);
xor XOR2 (N695, N662, N558);
nor NOR4 (N696, N673, N571, N629, N490);
and AND4 (N697, N695, N20, N130, N137);
nand NAND4 (N698, N675, N544, N468, N423);
nor NOR2 (N699, N682, N449);
nor NOR4 (N700, N699, N220, N95, N515);
or OR2 (N701, N690, N147);
or OR3 (N702, N697, N577, N204);
nand NAND2 (N703, N691, N660);
buf BUF1 (N704, N692);
or OR4 (N705, N693, N210, N166, N149);
or OR3 (N706, N703, N673, N154);
and AND2 (N707, N701, N123);
xor XOR2 (N708, N705, N191);
xor XOR2 (N709, N707, N601);
or OR4 (N710, N696, N185, N373, N488);
nand NAND4 (N711, N700, N184, N162, N223);
buf BUF1 (N712, N704);
buf BUF1 (N713, N694);
nor NOR4 (N714, N698, N270, N418, N74);
not NOT1 (N715, N685);
xor XOR2 (N716, N708, N432);
buf BUF1 (N717, N716);
xor XOR2 (N718, N711, N58);
buf BUF1 (N719, N713);
nand NAND3 (N720, N702, N15, N643);
nor NOR3 (N721, N714, N331, N36);
or OR4 (N722, N718, N283, N373, N623);
buf BUF1 (N723, N721);
and AND2 (N724, N709, N640);
xor XOR2 (N725, N723, N659);
or OR4 (N726, N717, N714, N531, N47);
buf BUF1 (N727, N725);
xor XOR2 (N728, N726, N516);
nor NOR3 (N729, N727, N516, N448);
buf BUF1 (N730, N722);
nor NOR3 (N731, N730, N383, N474);
buf BUF1 (N732, N724);
nand NAND4 (N733, N715, N116, N287, N606);
or OR2 (N734, N706, N676);
nand NAND2 (N735, N712, N262);
buf BUF1 (N736, N735);
not NOT1 (N737, N733);
nand NAND3 (N738, N737, N656, N167);
nor NOR2 (N739, N731, N651);
nor NOR4 (N740, N738, N267, N409, N8);
xor XOR2 (N741, N728, N576);
or OR2 (N742, N740, N412);
not NOT1 (N743, N719);
nand NAND2 (N744, N742, N103);
nand NAND2 (N745, N710, N96);
and AND4 (N746, N732, N566, N342, N518);
and AND2 (N747, N729, N476);
nor NOR3 (N748, N744, N233, N319);
nand NAND2 (N749, N734, N673);
nor NOR3 (N750, N743, N551, N441);
not NOT1 (N751, N750);
nand NAND2 (N752, N746, N17);
and AND4 (N753, N752, N464, N290, N667);
and AND2 (N754, N739, N595);
nor NOR2 (N755, N751, N382);
nand NAND2 (N756, N748, N615);
not NOT1 (N757, N720);
not NOT1 (N758, N747);
xor XOR2 (N759, N757, N119);
nand NAND3 (N760, N759, N396, N555);
buf BUF1 (N761, N749);
buf BUF1 (N762, N760);
and AND3 (N763, N761, N253, N695);
nand NAND4 (N764, N741, N367, N517, N479);
or OR2 (N765, N764, N518);
nor NOR4 (N766, N755, N684, N410, N514);
not NOT1 (N767, N754);
buf BUF1 (N768, N762);
and AND2 (N769, N756, N669);
and AND3 (N770, N745, N692, N732);
nor NOR3 (N771, N758, N313, N751);
nor NOR4 (N772, N770, N311, N144, N256);
xor XOR2 (N773, N763, N714);
xor XOR2 (N774, N768, N84);
not NOT1 (N775, N767);
nand NAND3 (N776, N771, N137, N105);
and AND4 (N777, N773, N331, N356, N617);
or OR4 (N778, N772, N95, N244, N415);
nor NOR2 (N779, N774, N778);
nand NAND2 (N780, N399, N514);
or OR4 (N781, N776, N138, N605, N124);
not NOT1 (N782, N753);
nor NOR4 (N783, N765, N716, N433, N663);
and AND4 (N784, N736, N508, N326, N180);
not NOT1 (N785, N784);
or OR4 (N786, N769, N559, N41, N345);
nor NOR4 (N787, N777, N19, N532, N398);
xor XOR2 (N788, N781, N246);
xor XOR2 (N789, N780, N325);
nor NOR3 (N790, N789, N335, N48);
xor XOR2 (N791, N786, N551);
xor XOR2 (N792, N791, N195);
buf BUF1 (N793, N787);
xor XOR2 (N794, N779, N606);
xor XOR2 (N795, N782, N525);
and AND3 (N796, N790, N792, N688);
and AND4 (N797, N71, N684, N764, N281);
xor XOR2 (N798, N793, N700);
xor XOR2 (N799, N797, N797);
not NOT1 (N800, N783);
xor XOR2 (N801, N794, N733);
and AND2 (N802, N788, N409);
and AND4 (N803, N801, N793, N174, N430);
nand NAND4 (N804, N785, N441, N788, N362);
nor NOR2 (N805, N796, N353);
nand NAND2 (N806, N798, N360);
and AND3 (N807, N805, N242, N15);
and AND2 (N808, N799, N273);
or OR4 (N809, N775, N214, N668, N100);
not NOT1 (N810, N807);
xor XOR2 (N811, N806, N620);
buf BUF1 (N812, N802);
nand NAND4 (N813, N811, N385, N227, N773);
buf BUF1 (N814, N804);
not NOT1 (N815, N803);
buf BUF1 (N816, N809);
or OR2 (N817, N810, N401);
or OR4 (N818, N817, N311, N208, N607);
or OR4 (N819, N816, N104, N739, N729);
not NOT1 (N820, N814);
buf BUF1 (N821, N818);
not NOT1 (N822, N821);
buf BUF1 (N823, N800);
buf BUF1 (N824, N819);
nor NOR3 (N825, N812, N695, N159);
or OR4 (N826, N820, N706, N664, N289);
nand NAND4 (N827, N823, N296, N752, N447);
and AND2 (N828, N766, N645);
and AND3 (N829, N828, N633, N460);
nand NAND2 (N830, N825, N369);
buf BUF1 (N831, N813);
nor NOR2 (N832, N830, N239);
or OR3 (N833, N822, N41, N208);
or OR4 (N834, N808, N71, N266, N833);
buf BUF1 (N835, N104);
or OR3 (N836, N824, N420, N95);
nand NAND2 (N837, N795, N537);
and AND2 (N838, N827, N479);
nor NOR4 (N839, N829, N415, N671, N457);
buf BUF1 (N840, N836);
nor NOR3 (N841, N834, N573, N608);
nand NAND2 (N842, N826, N431);
and AND4 (N843, N839, N674, N578, N448);
nor NOR3 (N844, N840, N494, N524);
and AND3 (N845, N838, N240, N623);
not NOT1 (N846, N815);
not NOT1 (N847, N846);
and AND2 (N848, N845, N31);
and AND4 (N849, N841, N567, N501, N715);
nand NAND4 (N850, N848, N8, N357, N570);
nand NAND3 (N851, N850, N320, N802);
not NOT1 (N852, N849);
nand NAND4 (N853, N847, N49, N205, N760);
or OR4 (N854, N852, N806, N313, N349);
xor XOR2 (N855, N854, N29);
buf BUF1 (N856, N837);
nor NOR3 (N857, N832, N664, N690);
not NOT1 (N858, N853);
buf BUF1 (N859, N835);
xor XOR2 (N860, N858, N775);
buf BUF1 (N861, N859);
or OR4 (N862, N860, N405, N124, N325);
and AND4 (N863, N856, N144, N206, N670);
and AND4 (N864, N844, N760, N6, N460);
not NOT1 (N865, N843);
nor NOR2 (N866, N855, N834);
or OR4 (N867, N863, N534, N258, N436);
not NOT1 (N868, N864);
not NOT1 (N869, N842);
not NOT1 (N870, N869);
and AND3 (N871, N831, N641, N396);
or OR4 (N872, N857, N50, N786, N570);
buf BUF1 (N873, N872);
xor XOR2 (N874, N870, N243);
or OR4 (N875, N874, N75, N218, N226);
nand NAND2 (N876, N873, N182);
and AND2 (N877, N851, N274);
nand NAND4 (N878, N876, N574, N254, N209);
and AND4 (N879, N878, N526, N795, N823);
or OR4 (N880, N879, N861, N474, N19);
not NOT1 (N881, N457);
xor XOR2 (N882, N877, N272);
xor XOR2 (N883, N871, N867);
nand NAND2 (N884, N804, N745);
and AND4 (N885, N880, N516, N166, N498);
nand NAND4 (N886, N882, N230, N30, N332);
not NOT1 (N887, N862);
and AND4 (N888, N887, N596, N809, N51);
or OR4 (N889, N886, N350, N591, N395);
nor NOR3 (N890, N884, N55, N44);
nor NOR3 (N891, N868, N223, N41);
not NOT1 (N892, N875);
nand NAND4 (N893, N866, N761, N405, N492);
and AND3 (N894, N865, N679, N591);
nand NAND4 (N895, N893, N653, N700, N197);
nand NAND4 (N896, N890, N86, N546, N272);
not NOT1 (N897, N883);
not NOT1 (N898, N888);
buf BUF1 (N899, N896);
nor NOR3 (N900, N892, N413, N477);
buf BUF1 (N901, N900);
nand NAND2 (N902, N901, N885);
and AND4 (N903, N575, N683, N590, N435);
nand NAND3 (N904, N894, N692, N195);
or OR2 (N905, N891, N603);
and AND4 (N906, N898, N235, N133, N20);
and AND4 (N907, N906, N248, N106, N856);
nand NAND3 (N908, N903, N639, N831);
nor NOR2 (N909, N895, N215);
xor XOR2 (N910, N905, N442);
nor NOR3 (N911, N889, N336, N700);
and AND4 (N912, N899, N273, N389, N181);
buf BUF1 (N913, N911);
and AND2 (N914, N907, N869);
buf BUF1 (N915, N910);
xor XOR2 (N916, N912, N232);
or OR4 (N917, N902, N434, N602, N699);
buf BUF1 (N918, N917);
buf BUF1 (N919, N916);
nor NOR4 (N920, N918, N854, N860, N887);
nand NAND4 (N921, N913, N616, N841, N638);
buf BUF1 (N922, N921);
xor XOR2 (N923, N897, N656);
and AND3 (N924, N923, N859, N439);
nor NOR4 (N925, N908, N339, N317, N435);
buf BUF1 (N926, N914);
nor NOR4 (N927, N922, N867, N71, N440);
not NOT1 (N928, N904);
and AND4 (N929, N928, N664, N523, N923);
xor XOR2 (N930, N909, N27);
or OR2 (N931, N881, N368);
not NOT1 (N932, N924);
and AND2 (N933, N915, N443);
nor NOR3 (N934, N927, N172, N365);
buf BUF1 (N935, N932);
or OR3 (N936, N925, N705, N651);
buf BUF1 (N937, N936);
or OR3 (N938, N926, N745, N477);
or OR2 (N939, N934, N718);
nand NAND2 (N940, N919, N597);
buf BUF1 (N941, N920);
nor NOR2 (N942, N935, N626);
or OR3 (N943, N930, N835, N820);
nand NAND3 (N944, N942, N488, N70);
xor XOR2 (N945, N931, N667);
xor XOR2 (N946, N944, N529);
nor NOR3 (N947, N938, N552, N901);
buf BUF1 (N948, N939);
nor NOR3 (N949, N946, N806, N347);
buf BUF1 (N950, N943);
nand NAND3 (N951, N945, N536, N680);
and AND3 (N952, N948, N936, N584);
nor NOR4 (N953, N950, N870, N479, N556);
xor XOR2 (N954, N933, N746);
not NOT1 (N955, N952);
not NOT1 (N956, N955);
or OR4 (N957, N951, N231, N777, N313);
nand NAND2 (N958, N929, N533);
or OR4 (N959, N940, N749, N617, N703);
xor XOR2 (N960, N941, N151);
nor NOR4 (N961, N947, N851, N388, N776);
xor XOR2 (N962, N956, N491);
buf BUF1 (N963, N953);
not NOT1 (N964, N961);
not NOT1 (N965, N949);
nor NOR4 (N966, N958, N186, N109, N537);
buf BUF1 (N967, N966);
or OR2 (N968, N963, N120);
buf BUF1 (N969, N937);
nand NAND2 (N970, N967, N143);
and AND3 (N971, N964, N513, N319);
or OR4 (N972, N968, N801, N470, N841);
and AND4 (N973, N957, N835, N271, N852);
buf BUF1 (N974, N971);
and AND2 (N975, N954, N185);
and AND4 (N976, N974, N119, N236, N10);
not NOT1 (N977, N962);
nand NAND2 (N978, N977, N316);
not NOT1 (N979, N972);
xor XOR2 (N980, N978, N527);
xor XOR2 (N981, N969, N415);
not NOT1 (N982, N965);
xor XOR2 (N983, N959, N79);
nand NAND3 (N984, N960, N632, N412);
and AND4 (N985, N983, N673, N948, N70);
xor XOR2 (N986, N970, N852);
not NOT1 (N987, N976);
nand NAND2 (N988, N987, N800);
nor NOR3 (N989, N986, N219, N964);
or OR2 (N990, N979, N277);
buf BUF1 (N991, N984);
or OR3 (N992, N990, N470, N296);
nor NOR4 (N993, N980, N672, N129, N367);
xor XOR2 (N994, N988, N871);
and AND2 (N995, N985, N486);
nor NOR3 (N996, N975, N517, N894);
nor NOR4 (N997, N993, N207, N982, N246);
nand NAND3 (N998, N475, N604, N488);
and AND2 (N999, N995, N68);
not NOT1 (N1000, N991);
buf BUF1 (N1001, N997);
buf BUF1 (N1002, N1001);
xor XOR2 (N1003, N996, N524);
buf BUF1 (N1004, N1003);
and AND3 (N1005, N989, N136, N110);
and AND4 (N1006, N994, N126, N682, N659);
xor XOR2 (N1007, N1000, N277);
buf BUF1 (N1008, N1002);
nand NAND3 (N1009, N999, N755, N340);
nor NOR4 (N1010, N1008, N85, N755, N691);
buf BUF1 (N1011, N1006);
nand NAND3 (N1012, N1004, N911, N196);
nor NOR4 (N1013, N973, N465, N729, N642);
xor XOR2 (N1014, N992, N820);
and AND2 (N1015, N998, N508);
and AND2 (N1016, N981, N913);
and AND3 (N1017, N1013, N1001, N402);
buf BUF1 (N1018, N1016);
nand NAND2 (N1019, N1009, N470);
not NOT1 (N1020, N1014);
nor NOR4 (N1021, N1015, N858, N713, N259);
or OR2 (N1022, N1012, N582);
and AND4 (N1023, N1018, N483, N795, N507);
and AND3 (N1024, N1019, N79, N336);
not NOT1 (N1025, N1022);
and AND4 (N1026, N1020, N816, N49, N626);
buf BUF1 (N1027, N1021);
or OR2 (N1028, N1017, N488);
buf BUF1 (N1029, N1010);
buf BUF1 (N1030, N1007);
xor XOR2 (N1031, N1025, N138);
or OR2 (N1032, N1011, N734);
nor NOR2 (N1033, N1030, N650);
nor NOR4 (N1034, N1027, N303, N71, N802);
nand NAND4 (N1035, N1032, N134, N1031, N691);
and AND3 (N1036, N240, N649, N771);
not NOT1 (N1037, N1029);
xor XOR2 (N1038, N1028, N715);
and AND2 (N1039, N1005, N846);
nand NAND2 (N1040, N1024, N159);
buf BUF1 (N1041, N1040);
and AND4 (N1042, N1041, N933, N991, N709);
nand NAND2 (N1043, N1038, N35);
or OR4 (N1044, N1034, N515, N319, N82);
buf BUF1 (N1045, N1035);
nand NAND3 (N1046, N1036, N912, N798);
and AND3 (N1047, N1039, N273, N222);
nand NAND2 (N1048, N1047, N820);
xor XOR2 (N1049, N1023, N157);
nor NOR4 (N1050, N1044, N646, N539, N760);
nor NOR3 (N1051, N1042, N985, N277);
not NOT1 (N1052, N1045);
nand NAND3 (N1053, N1050, N276, N872);
buf BUF1 (N1054, N1026);
nand NAND4 (N1055, N1053, N456, N81, N1004);
nor NOR4 (N1056, N1046, N229, N540, N234);
or OR2 (N1057, N1055, N312);
and AND2 (N1058, N1056, N697);
or OR4 (N1059, N1048, N641, N300, N79);
buf BUF1 (N1060, N1059);
nor NOR4 (N1061, N1054, N6, N109, N197);
buf BUF1 (N1062, N1051);
xor XOR2 (N1063, N1061, N255);
and AND3 (N1064, N1058, N408, N276);
buf BUF1 (N1065, N1064);
or OR4 (N1066, N1052, N1022, N319, N110);
nor NOR3 (N1067, N1057, N44, N100);
not NOT1 (N1068, N1066);
nor NOR4 (N1069, N1033, N73, N499, N189);
buf BUF1 (N1070, N1062);
and AND3 (N1071, N1060, N700, N578);
and AND4 (N1072, N1063, N598, N1036, N139);
nand NAND4 (N1073, N1071, N39, N272, N320);
or OR4 (N1074, N1070, N569, N867, N846);
and AND2 (N1075, N1073, N170);
buf BUF1 (N1076, N1072);
and AND2 (N1077, N1075, N666);
not NOT1 (N1078, N1077);
and AND3 (N1079, N1078, N379, N399);
nor NOR2 (N1080, N1069, N680);
nor NOR2 (N1081, N1049, N92);
nand NAND2 (N1082, N1079, N809);
buf BUF1 (N1083, N1080);
buf BUF1 (N1084, N1043);
buf BUF1 (N1085, N1082);
nand NAND2 (N1086, N1065, N112);
not NOT1 (N1087, N1076);
or OR2 (N1088, N1067, N394);
xor XOR2 (N1089, N1088, N364);
nor NOR3 (N1090, N1074, N490, N485);
xor XOR2 (N1091, N1085, N427);
not NOT1 (N1092, N1037);
nand NAND2 (N1093, N1090, N147);
xor XOR2 (N1094, N1091, N475);
not NOT1 (N1095, N1089);
nand NAND3 (N1096, N1093, N138, N979);
buf BUF1 (N1097, N1094);
and AND2 (N1098, N1081, N709);
xor XOR2 (N1099, N1084, N798);
not NOT1 (N1100, N1099);
buf BUF1 (N1101, N1098);
buf BUF1 (N1102, N1101);
buf BUF1 (N1103, N1092);
and AND2 (N1104, N1083, N596);
nand NAND2 (N1105, N1097, N100);
buf BUF1 (N1106, N1068);
and AND4 (N1107, N1095, N1100, N912, N759);
xor XOR2 (N1108, N1071, N232);
nand NAND3 (N1109, N1104, N1024, N841);
nor NOR4 (N1110, N1107, N985, N81, N40);
xor XOR2 (N1111, N1109, N796);
or OR4 (N1112, N1086, N1095, N244, N867);
nor NOR3 (N1113, N1103, N907, N638);
and AND4 (N1114, N1113, N55, N315, N1096);
buf BUF1 (N1115, N835);
or OR3 (N1116, N1112, N118, N691);
xor XOR2 (N1117, N1114, N432);
or OR3 (N1118, N1105, N718, N409);
nor NOR3 (N1119, N1106, N609, N501);
nor NOR4 (N1120, N1102, N934, N413, N600);
not NOT1 (N1121, N1119);
nand NAND3 (N1122, N1108, N334, N504);
xor XOR2 (N1123, N1111, N413);
or OR2 (N1124, N1122, N710);
or OR3 (N1125, N1087, N261, N158);
xor XOR2 (N1126, N1125, N14);
xor XOR2 (N1127, N1124, N424);
xor XOR2 (N1128, N1121, N146);
or OR2 (N1129, N1126, N619);
and AND2 (N1130, N1127, N323);
buf BUF1 (N1131, N1110);
not NOT1 (N1132, N1130);
buf BUF1 (N1133, N1131);
xor XOR2 (N1134, N1116, N887);
buf BUF1 (N1135, N1115);
xor XOR2 (N1136, N1128, N507);
nor NOR4 (N1137, N1129, N1029, N1112, N448);
buf BUF1 (N1138, N1135);
not NOT1 (N1139, N1117);
and AND3 (N1140, N1132, N323, N119);
nor NOR2 (N1141, N1120, N250);
not NOT1 (N1142, N1137);
and AND2 (N1143, N1123, N214);
or OR4 (N1144, N1136, N74, N61, N549);
or OR3 (N1145, N1139, N975, N1021);
or OR2 (N1146, N1144, N602);
nor NOR4 (N1147, N1146, N349, N118, N865);
nand NAND2 (N1148, N1147, N137);
xor XOR2 (N1149, N1145, N449);
nor NOR3 (N1150, N1118, N959, N1024);
not NOT1 (N1151, N1148);
not NOT1 (N1152, N1134);
xor XOR2 (N1153, N1142, N56);
buf BUF1 (N1154, N1153);
and AND3 (N1155, N1141, N175, N839);
xor XOR2 (N1156, N1143, N386);
nor NOR3 (N1157, N1154, N948, N599);
not NOT1 (N1158, N1151);
xor XOR2 (N1159, N1156, N47);
xor XOR2 (N1160, N1149, N724);
or OR3 (N1161, N1140, N975, N894);
buf BUF1 (N1162, N1158);
nand NAND4 (N1163, N1133, N723, N819, N849);
nand NAND2 (N1164, N1155, N692);
nor NOR4 (N1165, N1138, N952, N362, N563);
xor XOR2 (N1166, N1164, N325);
nand NAND2 (N1167, N1162, N911);
xor XOR2 (N1168, N1166, N568);
and AND2 (N1169, N1163, N659);
nor NOR2 (N1170, N1165, N197);
nor NOR3 (N1171, N1169, N1025, N829);
not NOT1 (N1172, N1161);
and AND4 (N1173, N1168, N46, N390, N51);
and AND2 (N1174, N1171, N1163);
buf BUF1 (N1175, N1157);
not NOT1 (N1176, N1173);
not NOT1 (N1177, N1167);
or OR2 (N1178, N1172, N962);
nand NAND3 (N1179, N1177, N146, N288);
nor NOR4 (N1180, N1179, N923, N713, N166);
nand NAND2 (N1181, N1159, N350);
nor NOR3 (N1182, N1176, N116, N692);
or OR2 (N1183, N1160, N674);
buf BUF1 (N1184, N1170);
and AND2 (N1185, N1181, N362);
nor NOR4 (N1186, N1178, N1161, N473, N716);
and AND3 (N1187, N1185, N990, N1185);
buf BUF1 (N1188, N1150);
nand NAND4 (N1189, N1186, N991, N1173, N282);
not NOT1 (N1190, N1174);
nand NAND4 (N1191, N1180, N528, N491, N775);
not NOT1 (N1192, N1182);
xor XOR2 (N1193, N1192, N695);
buf BUF1 (N1194, N1188);
not NOT1 (N1195, N1152);
and AND2 (N1196, N1190, N574);
buf BUF1 (N1197, N1194);
not NOT1 (N1198, N1193);
xor XOR2 (N1199, N1195, N71);
and AND3 (N1200, N1183, N499, N946);
not NOT1 (N1201, N1184);
nor NOR4 (N1202, N1200, N542, N1159, N1193);
or OR2 (N1203, N1199, N1082);
nand NAND3 (N1204, N1197, N533, N771);
xor XOR2 (N1205, N1196, N1029);
not NOT1 (N1206, N1189);
and AND2 (N1207, N1206, N263);
buf BUF1 (N1208, N1201);
nand NAND3 (N1209, N1202, N818, N659);
and AND2 (N1210, N1205, N601);
and AND2 (N1211, N1203, N745);
nor NOR3 (N1212, N1187, N943, N512);
nand NAND3 (N1213, N1211, N819, N1180);
or OR4 (N1214, N1212, N87, N344, N216);
or OR4 (N1215, N1208, N777, N185, N529);
and AND3 (N1216, N1210, N807, N1127);
buf BUF1 (N1217, N1198);
buf BUF1 (N1218, N1214);
buf BUF1 (N1219, N1218);
and AND2 (N1220, N1207, N621);
nand NAND2 (N1221, N1215, N729);
nor NOR4 (N1222, N1217, N763, N809, N1200);
and AND3 (N1223, N1220, N1012, N366);
not NOT1 (N1224, N1175);
and AND4 (N1225, N1221, N1156, N529, N689);
and AND2 (N1226, N1222, N701);
nor NOR4 (N1227, N1223, N326, N1150, N819);
not NOT1 (N1228, N1209);
nor NOR4 (N1229, N1191, N1035, N351, N606);
and AND4 (N1230, N1216, N447, N108, N895);
or OR2 (N1231, N1219, N1080);
nor NOR2 (N1232, N1225, N707);
xor XOR2 (N1233, N1226, N390);
and AND3 (N1234, N1229, N139, N1053);
buf BUF1 (N1235, N1213);
nor NOR3 (N1236, N1204, N492, N1138);
and AND3 (N1237, N1224, N361, N1023);
buf BUF1 (N1238, N1234);
not NOT1 (N1239, N1228);
nor NOR2 (N1240, N1237, N244);
nor NOR3 (N1241, N1230, N661, N123);
nor NOR2 (N1242, N1235, N952);
or OR4 (N1243, N1239, N988, N414, N736);
nand NAND3 (N1244, N1240, N1002, N985);
nor NOR2 (N1245, N1243, N514);
and AND4 (N1246, N1227, N894, N319, N453);
not NOT1 (N1247, N1236);
nand NAND3 (N1248, N1232, N1148, N1193);
nand NAND3 (N1249, N1246, N207, N624);
or OR3 (N1250, N1233, N651, N390);
buf BUF1 (N1251, N1238);
or OR3 (N1252, N1250, N514, N646);
and AND2 (N1253, N1252, N302);
and AND3 (N1254, N1253, N613, N248);
xor XOR2 (N1255, N1251, N617);
nand NAND2 (N1256, N1248, N525);
and AND2 (N1257, N1255, N515);
xor XOR2 (N1258, N1241, N226);
and AND2 (N1259, N1244, N485);
buf BUF1 (N1260, N1249);
buf BUF1 (N1261, N1256);
and AND3 (N1262, N1247, N380, N627);
nor NOR3 (N1263, N1231, N1005, N1001);
nand NAND2 (N1264, N1261, N220);
nand NAND3 (N1265, N1242, N79, N1257);
or OR2 (N1266, N350, N80);
nand NAND3 (N1267, N1262, N584, N765);
nand NAND3 (N1268, N1266, N307, N1054);
or OR2 (N1269, N1268, N11);
and AND4 (N1270, N1264, N1237, N767, N715);
and AND2 (N1271, N1259, N181);
not NOT1 (N1272, N1265);
not NOT1 (N1273, N1272);
and AND2 (N1274, N1271, N436);
nor NOR3 (N1275, N1260, N1137, N476);
not NOT1 (N1276, N1275);
xor XOR2 (N1277, N1267, N260);
nand NAND3 (N1278, N1273, N1238, N1073);
nor NOR3 (N1279, N1269, N938, N696);
xor XOR2 (N1280, N1254, N425);
xor XOR2 (N1281, N1270, N966);
nor NOR3 (N1282, N1276, N1212, N796);
not NOT1 (N1283, N1263);
or OR4 (N1284, N1274, N512, N847, N170);
nand NAND2 (N1285, N1277, N1165);
nand NAND2 (N1286, N1281, N247);
and AND4 (N1287, N1286, N1226, N186, N35);
and AND3 (N1288, N1283, N1225, N576);
or OR2 (N1289, N1284, N596);
not NOT1 (N1290, N1245);
xor XOR2 (N1291, N1282, N1242);
nand NAND4 (N1292, N1287, N1004, N1254, N1180);
xor XOR2 (N1293, N1289, N609);
xor XOR2 (N1294, N1288, N718);
nor NOR2 (N1295, N1292, N1253);
xor XOR2 (N1296, N1258, N434);
and AND4 (N1297, N1294, N176, N1130, N79);
xor XOR2 (N1298, N1291, N986);
nand NAND3 (N1299, N1290, N449, N193);
not NOT1 (N1300, N1278);
or OR2 (N1301, N1297, N1300);
and AND4 (N1302, N110, N572, N1292, N854);
or OR4 (N1303, N1280, N46, N238, N363);
and AND3 (N1304, N1285, N787, N989);
nor NOR4 (N1305, N1279, N1011, N1200, N989);
not NOT1 (N1306, N1302);
buf BUF1 (N1307, N1295);
not NOT1 (N1308, N1293);
nand NAND3 (N1309, N1303, N201, N798);
buf BUF1 (N1310, N1309);
or OR3 (N1311, N1310, N47, N1131);
nor NOR3 (N1312, N1296, N765, N151);
xor XOR2 (N1313, N1312, N349);
or OR4 (N1314, N1311, N19, N488, N640);
nand NAND2 (N1315, N1298, N211);
not NOT1 (N1316, N1299);
not NOT1 (N1317, N1314);
nor NOR4 (N1318, N1313, N892, N5, N301);
nand NAND3 (N1319, N1316, N1281, N141);
buf BUF1 (N1320, N1318);
nor NOR2 (N1321, N1308, N673);
nor NOR3 (N1322, N1305, N881, N293);
and AND2 (N1323, N1307, N911);
not NOT1 (N1324, N1320);
not NOT1 (N1325, N1321);
or OR2 (N1326, N1319, N190);
nor NOR4 (N1327, N1324, N191, N334, N540);
nor NOR2 (N1328, N1304, N645);
not NOT1 (N1329, N1317);
xor XOR2 (N1330, N1323, N1201);
and AND2 (N1331, N1325, N1292);
xor XOR2 (N1332, N1306, N1324);
buf BUF1 (N1333, N1327);
nand NAND2 (N1334, N1326, N942);
not NOT1 (N1335, N1330);
or OR3 (N1336, N1333, N777, N906);
or OR2 (N1337, N1336, N295);
or OR2 (N1338, N1301, N1270);
and AND3 (N1339, N1334, N949, N474);
and AND4 (N1340, N1329, N1308, N1337, N82);
and AND3 (N1341, N463, N86, N1249);
not NOT1 (N1342, N1331);
nor NOR3 (N1343, N1315, N252, N474);
or OR2 (N1344, N1328, N297);
xor XOR2 (N1345, N1343, N1332);
not NOT1 (N1346, N777);
xor XOR2 (N1347, N1341, N1211);
or OR3 (N1348, N1345, N823, N837);
or OR3 (N1349, N1347, N333, N686);
nand NAND3 (N1350, N1322, N994, N642);
nor NOR3 (N1351, N1340, N887, N829);
xor XOR2 (N1352, N1346, N141);
buf BUF1 (N1353, N1352);
not NOT1 (N1354, N1344);
and AND2 (N1355, N1338, N1068);
buf BUF1 (N1356, N1355);
or OR2 (N1357, N1339, N387);
or OR3 (N1358, N1351, N1238, N67);
buf BUF1 (N1359, N1353);
or OR3 (N1360, N1335, N401, N1113);
nor NOR4 (N1361, N1359, N286, N1201, N657);
xor XOR2 (N1362, N1361, N191);
buf BUF1 (N1363, N1348);
nand NAND2 (N1364, N1362, N958);
buf BUF1 (N1365, N1364);
or OR2 (N1366, N1349, N1360);
not NOT1 (N1367, N97);
nor NOR3 (N1368, N1365, N69, N1138);
buf BUF1 (N1369, N1358);
buf BUF1 (N1370, N1354);
xor XOR2 (N1371, N1357, N453);
not NOT1 (N1372, N1366);
nand NAND4 (N1373, N1370, N129, N382, N999);
or OR2 (N1374, N1356, N318);
xor XOR2 (N1375, N1372, N24);
nor NOR3 (N1376, N1373, N250, N154);
xor XOR2 (N1377, N1369, N498);
or OR2 (N1378, N1342, N752);
not NOT1 (N1379, N1377);
nor NOR4 (N1380, N1374, N649, N33, N187);
nor NOR4 (N1381, N1379, N1000, N726, N194);
buf BUF1 (N1382, N1381);
or OR3 (N1383, N1378, N59, N1194);
buf BUF1 (N1384, N1376);
xor XOR2 (N1385, N1368, N1224);
and AND3 (N1386, N1380, N246, N1084);
xor XOR2 (N1387, N1350, N524);
xor XOR2 (N1388, N1375, N674);
not NOT1 (N1389, N1387);
nor NOR4 (N1390, N1386, N344, N179, N493);
not NOT1 (N1391, N1367);
buf BUF1 (N1392, N1385);
not NOT1 (N1393, N1371);
nand NAND2 (N1394, N1383, N605);
or OR2 (N1395, N1363, N866);
nor NOR3 (N1396, N1393, N1235, N968);
and AND3 (N1397, N1384, N645, N1142);
or OR4 (N1398, N1389, N1056, N332, N1101);
buf BUF1 (N1399, N1394);
nor NOR4 (N1400, N1396, N14, N1050, N857);
or OR4 (N1401, N1400, N666, N1059, N242);
nor NOR4 (N1402, N1395, N152, N273, N1096);
and AND2 (N1403, N1397, N1322);
not NOT1 (N1404, N1401);
or OR3 (N1405, N1398, N177, N510);
or OR3 (N1406, N1390, N708, N1);
or OR3 (N1407, N1399, N1145, N320);
and AND3 (N1408, N1392, N897, N613);
xor XOR2 (N1409, N1406, N978);
xor XOR2 (N1410, N1407, N382);
not NOT1 (N1411, N1408);
nand NAND3 (N1412, N1402, N927, N232);
and AND4 (N1413, N1405, N563, N321, N131);
nand NAND3 (N1414, N1409, N647, N1273);
nor NOR2 (N1415, N1411, N281);
nand NAND2 (N1416, N1403, N560);
and AND3 (N1417, N1382, N871, N6);
buf BUF1 (N1418, N1391);
not NOT1 (N1419, N1413);
nand NAND4 (N1420, N1415, N1352, N589, N1077);
xor XOR2 (N1421, N1419, N211);
not NOT1 (N1422, N1418);
not NOT1 (N1423, N1412);
nand NAND3 (N1424, N1414, N156, N922);
nand NAND3 (N1425, N1417, N1243, N235);
nor NOR4 (N1426, N1421, N1035, N1291, N186);
and AND3 (N1427, N1388, N611, N1270);
nand NAND3 (N1428, N1426, N478, N38);
xor XOR2 (N1429, N1404, N414);
and AND2 (N1430, N1429, N599);
and AND4 (N1431, N1427, N134, N1397, N547);
nor NOR3 (N1432, N1420, N923, N663);
buf BUF1 (N1433, N1428);
nand NAND3 (N1434, N1410, N814, N710);
not NOT1 (N1435, N1432);
nand NAND2 (N1436, N1416, N1335);
nor NOR2 (N1437, N1431, N346);
xor XOR2 (N1438, N1437, N101);
xor XOR2 (N1439, N1424, N806);
buf BUF1 (N1440, N1434);
nand NAND2 (N1441, N1438, N433);
not NOT1 (N1442, N1439);
not NOT1 (N1443, N1442);
nor NOR4 (N1444, N1425, N1008, N458, N605);
nor NOR4 (N1445, N1444, N91, N898, N1335);
buf BUF1 (N1446, N1436);
or OR4 (N1447, N1441, N945, N1034, N224);
not NOT1 (N1448, N1446);
or OR3 (N1449, N1422, N934, N265);
buf BUF1 (N1450, N1423);
xor XOR2 (N1451, N1448, N835);
or OR4 (N1452, N1450, N267, N225, N289);
nor NOR3 (N1453, N1443, N347, N196);
nand NAND4 (N1454, N1433, N643, N545, N874);
or OR2 (N1455, N1452, N1018);
and AND4 (N1456, N1440, N668, N889, N1439);
or OR4 (N1457, N1451, N471, N1154, N340);
and AND3 (N1458, N1453, N1154, N362);
not NOT1 (N1459, N1430);
buf BUF1 (N1460, N1454);
not NOT1 (N1461, N1455);
xor XOR2 (N1462, N1445, N776);
xor XOR2 (N1463, N1456, N208);
nand NAND3 (N1464, N1463, N589, N578);
and AND4 (N1465, N1460, N14, N304, N962);
nor NOR4 (N1466, N1459, N334, N846, N1285);
nor NOR2 (N1467, N1465, N1351);
buf BUF1 (N1468, N1466);
buf BUF1 (N1469, N1435);
and AND3 (N1470, N1462, N385, N1156);
nor NOR4 (N1471, N1457, N805, N557, N1135);
not NOT1 (N1472, N1461);
nor NOR2 (N1473, N1471, N574);
or OR4 (N1474, N1449, N813, N1198, N497);
xor XOR2 (N1475, N1472, N1094);
nor NOR2 (N1476, N1468, N220);
xor XOR2 (N1477, N1469, N909);
buf BUF1 (N1478, N1477);
xor XOR2 (N1479, N1474, N492);
nor NOR2 (N1480, N1458, N190);
xor XOR2 (N1481, N1475, N882);
xor XOR2 (N1482, N1478, N218);
or OR3 (N1483, N1473, N686, N658);
xor XOR2 (N1484, N1447, N1298);
not NOT1 (N1485, N1481);
and AND3 (N1486, N1464, N1348, N953);
xor XOR2 (N1487, N1484, N1325);
or OR2 (N1488, N1476, N335);
and AND4 (N1489, N1467, N171, N909, N1232);
or OR2 (N1490, N1488, N110);
nand NAND4 (N1491, N1482, N555, N97, N537);
nor NOR3 (N1492, N1486, N790, N683);
nor NOR4 (N1493, N1492, N1366, N749, N1231);
and AND2 (N1494, N1489, N260);
xor XOR2 (N1495, N1490, N1313);
nand NAND4 (N1496, N1479, N1113, N658, N909);
not NOT1 (N1497, N1491);
nor NOR2 (N1498, N1483, N371);
and AND2 (N1499, N1495, N1296);
buf BUF1 (N1500, N1497);
and AND3 (N1501, N1499, N200, N861);
not NOT1 (N1502, N1487);
and AND3 (N1503, N1485, N874, N1116);
not NOT1 (N1504, N1496);
xor XOR2 (N1505, N1493, N900);
nand NAND3 (N1506, N1503, N1215, N1311);
xor XOR2 (N1507, N1504, N1176);
nand NAND3 (N1508, N1470, N1249, N1127);
nor NOR4 (N1509, N1505, N1278, N672, N881);
not NOT1 (N1510, N1480);
or OR2 (N1511, N1501, N1377);
and AND3 (N1512, N1509, N370, N1115);
nor NOR2 (N1513, N1507, N1507);
not NOT1 (N1514, N1513);
nor NOR2 (N1515, N1500, N579);
nand NAND2 (N1516, N1514, N137);
nor NOR3 (N1517, N1506, N50, N481);
or OR2 (N1518, N1511, N1015);
nand NAND2 (N1519, N1515, N306);
and AND2 (N1520, N1518, N197);
xor XOR2 (N1521, N1510, N573);
buf BUF1 (N1522, N1498);
xor XOR2 (N1523, N1520, N447);
nor NOR2 (N1524, N1517, N922);
nor NOR3 (N1525, N1502, N188, N448);
or OR2 (N1526, N1519, N839);
not NOT1 (N1527, N1525);
and AND2 (N1528, N1508, N52);
buf BUF1 (N1529, N1522);
not NOT1 (N1530, N1529);
xor XOR2 (N1531, N1528, N1366);
or OR3 (N1532, N1512, N538, N407);
nand NAND3 (N1533, N1521, N1331, N805);
xor XOR2 (N1534, N1530, N1465);
nor NOR2 (N1535, N1531, N1262);
and AND2 (N1536, N1523, N1477);
nand NAND4 (N1537, N1533, N454, N1441, N916);
not NOT1 (N1538, N1536);
and AND4 (N1539, N1538, N306, N516, N31);
buf BUF1 (N1540, N1526);
buf BUF1 (N1541, N1524);
not NOT1 (N1542, N1537);
not NOT1 (N1543, N1527);
nand NAND2 (N1544, N1542, N562);
nand NAND4 (N1545, N1535, N1232, N368, N1364);
and AND2 (N1546, N1541, N960);
and AND3 (N1547, N1494, N1070, N645);
and AND2 (N1548, N1546, N1248);
nor NOR3 (N1549, N1545, N506, N1129);
buf BUF1 (N1550, N1539);
and AND2 (N1551, N1550, N1254);
nor NOR3 (N1552, N1551, N534, N1082);
nor NOR2 (N1553, N1540, N651);
nand NAND3 (N1554, N1516, N283, N500);
not NOT1 (N1555, N1532);
or OR2 (N1556, N1534, N192);
nand NAND4 (N1557, N1547, N162, N631, N466);
nand NAND2 (N1558, N1554, N91);
or OR2 (N1559, N1549, N411);
buf BUF1 (N1560, N1557);
buf BUF1 (N1561, N1553);
nor NOR2 (N1562, N1552, N447);
xor XOR2 (N1563, N1562, N587);
nor NOR4 (N1564, N1559, N1497, N195, N968);
xor XOR2 (N1565, N1563, N526);
xor XOR2 (N1566, N1543, N1058);
not NOT1 (N1567, N1544);
and AND2 (N1568, N1564, N21);
or OR4 (N1569, N1561, N632, N1270, N499);
xor XOR2 (N1570, N1555, N52);
not NOT1 (N1571, N1560);
nand NAND4 (N1572, N1570, N766, N233, N1061);
nand NAND2 (N1573, N1567, N1275);
or OR2 (N1574, N1572, N87);
xor XOR2 (N1575, N1568, N637);
not NOT1 (N1576, N1566);
not NOT1 (N1577, N1574);
or OR4 (N1578, N1558, N686, N1479, N908);
or OR2 (N1579, N1565, N1083);
xor XOR2 (N1580, N1556, N747);
buf BUF1 (N1581, N1571);
nor NOR4 (N1582, N1576, N57, N675, N485);
nor NOR4 (N1583, N1575, N1219, N810, N1011);
not NOT1 (N1584, N1580);
nand NAND3 (N1585, N1584, N259, N1583);
buf BUF1 (N1586, N1406);
xor XOR2 (N1587, N1579, N860);
nor NOR2 (N1588, N1577, N923);
nor NOR2 (N1589, N1581, N790);
buf BUF1 (N1590, N1573);
nand NAND3 (N1591, N1569, N1372, N765);
nor NOR3 (N1592, N1582, N712, N1426);
not NOT1 (N1593, N1587);
xor XOR2 (N1594, N1589, N1476);
or OR4 (N1595, N1592, N1110, N175, N635);
nand NAND3 (N1596, N1594, N6, N867);
and AND3 (N1597, N1585, N1501, N825);
nand NAND4 (N1598, N1590, N1164, N1390, N136);
or OR4 (N1599, N1586, N362, N1427, N270);
nor NOR2 (N1600, N1596, N1172);
and AND3 (N1601, N1593, N49, N1530);
nand NAND3 (N1602, N1598, N342, N373);
buf BUF1 (N1603, N1588);
or OR3 (N1604, N1548, N1009, N820);
and AND3 (N1605, N1602, N1126, N1430);
xor XOR2 (N1606, N1600, N224);
and AND3 (N1607, N1597, N91, N195);
xor XOR2 (N1608, N1607, N1071);
nor NOR2 (N1609, N1604, N517);
buf BUF1 (N1610, N1606);
nor NOR2 (N1611, N1591, N962);
nor NOR2 (N1612, N1601, N497);
nand NAND4 (N1613, N1595, N59, N999, N395);
nor NOR3 (N1614, N1609, N812, N1385);
xor XOR2 (N1615, N1599, N1298);
and AND2 (N1616, N1578, N1577);
nand NAND3 (N1617, N1614, N954, N123);
or OR2 (N1618, N1605, N1037);
and AND3 (N1619, N1610, N710, N581);
nand NAND3 (N1620, N1619, N1542, N235);
nor NOR4 (N1621, N1613, N681, N516, N45);
nor NOR2 (N1622, N1611, N237);
buf BUF1 (N1623, N1612);
nor NOR3 (N1624, N1618, N16, N205);
not NOT1 (N1625, N1608);
nor NOR2 (N1626, N1617, N1148);
nor NOR4 (N1627, N1625, N1375, N575, N651);
nand NAND4 (N1628, N1621, N1061, N610, N1013);
nor NOR3 (N1629, N1628, N1237, N366);
and AND3 (N1630, N1620, N1011, N1503);
or OR3 (N1631, N1627, N617, N1497);
nor NOR4 (N1632, N1626, N1461, N25, N157);
or OR3 (N1633, N1632, N1239, N891);
or OR3 (N1634, N1615, N439, N320);
xor XOR2 (N1635, N1633, N1390);
or OR2 (N1636, N1622, N372);
nand NAND4 (N1637, N1623, N250, N1569, N306);
buf BUF1 (N1638, N1635);
xor XOR2 (N1639, N1637, N1184);
or OR4 (N1640, N1639, N1604, N409, N1490);
nor NOR2 (N1641, N1640, N820);
nor NOR4 (N1642, N1636, N1278, N749, N1489);
or OR2 (N1643, N1616, N1021);
and AND3 (N1644, N1603, N277, N1371);
buf BUF1 (N1645, N1624);
not NOT1 (N1646, N1634);
buf BUF1 (N1647, N1642);
not NOT1 (N1648, N1630);
buf BUF1 (N1649, N1641);
nand NAND4 (N1650, N1646, N578, N1215, N561);
or OR3 (N1651, N1649, N743, N307);
nand NAND4 (N1652, N1644, N1372, N125, N941);
and AND2 (N1653, N1648, N468);
buf BUF1 (N1654, N1647);
not NOT1 (N1655, N1653);
or OR2 (N1656, N1643, N1344);
and AND3 (N1657, N1631, N1339, N907);
not NOT1 (N1658, N1657);
buf BUF1 (N1659, N1652);
nor NOR3 (N1660, N1655, N645, N644);
and AND2 (N1661, N1638, N606);
nor NOR2 (N1662, N1654, N895);
nand NAND4 (N1663, N1629, N636, N506, N1150);
and AND2 (N1664, N1660, N826);
nand NAND3 (N1665, N1664, N125, N1420);
and AND4 (N1666, N1650, N1225, N1386, N1253);
nand NAND4 (N1667, N1658, N1356, N470, N538);
buf BUF1 (N1668, N1659);
xor XOR2 (N1669, N1656, N1336);
buf BUF1 (N1670, N1645);
xor XOR2 (N1671, N1663, N1415);
not NOT1 (N1672, N1671);
nand NAND4 (N1673, N1661, N400, N955, N711);
buf BUF1 (N1674, N1672);
and AND3 (N1675, N1674, N1466, N1373);
nand NAND4 (N1676, N1662, N373, N1365, N1387);
and AND3 (N1677, N1665, N189, N1030);
nor NOR4 (N1678, N1670, N247, N1641, N740);
not NOT1 (N1679, N1675);
xor XOR2 (N1680, N1666, N1087);
nand NAND4 (N1681, N1673, N214, N1076, N1538);
or OR4 (N1682, N1677, N658, N1520, N204);
not NOT1 (N1683, N1679);
and AND4 (N1684, N1669, N1554, N711, N359);
not NOT1 (N1685, N1684);
nor NOR3 (N1686, N1682, N264, N1291);
nand NAND4 (N1687, N1685, N408, N819, N641);
nor NOR3 (N1688, N1667, N929, N724);
xor XOR2 (N1689, N1683, N738);
xor XOR2 (N1690, N1676, N105);
xor XOR2 (N1691, N1680, N275);
nor NOR4 (N1692, N1689, N582, N1648, N570);
buf BUF1 (N1693, N1668);
or OR3 (N1694, N1690, N685, N886);
not NOT1 (N1695, N1686);
not NOT1 (N1696, N1694);
nor NOR3 (N1697, N1695, N1601, N339);
nor NOR2 (N1698, N1692, N872);
xor XOR2 (N1699, N1698, N1644);
nor NOR2 (N1700, N1687, N1135);
or OR3 (N1701, N1651, N803, N1153);
not NOT1 (N1702, N1701);
and AND2 (N1703, N1681, N730);
nand NAND4 (N1704, N1699, N1029, N1089, N863);
xor XOR2 (N1705, N1678, N519);
or OR4 (N1706, N1688, N1395, N1521, N1004);
not NOT1 (N1707, N1697);
xor XOR2 (N1708, N1703, N106);
not NOT1 (N1709, N1706);
not NOT1 (N1710, N1700);
and AND4 (N1711, N1705, N642, N1266, N1092);
not NOT1 (N1712, N1693);
nand NAND4 (N1713, N1708, N1608, N821, N445);
and AND4 (N1714, N1691, N203, N1396, N840);
nand NAND3 (N1715, N1707, N527, N532);
xor XOR2 (N1716, N1713, N595);
nor NOR3 (N1717, N1704, N1674, N1482);
nor NOR3 (N1718, N1711, N102, N336);
xor XOR2 (N1719, N1702, N886);
nor NOR2 (N1720, N1716, N463);
xor XOR2 (N1721, N1709, N1463);
not NOT1 (N1722, N1712);
xor XOR2 (N1723, N1720, N767);
nor NOR4 (N1724, N1721, N117, N1145, N974);
buf BUF1 (N1725, N1724);
not NOT1 (N1726, N1710);
or OR3 (N1727, N1725, N977, N739);
nand NAND4 (N1728, N1714, N1144, N855, N1397);
not NOT1 (N1729, N1717);
or OR3 (N1730, N1715, N230, N275);
or OR2 (N1731, N1723, N511);
xor XOR2 (N1732, N1731, N424);
xor XOR2 (N1733, N1718, N968);
xor XOR2 (N1734, N1733, N1239);
not NOT1 (N1735, N1729);
not NOT1 (N1736, N1726);
and AND2 (N1737, N1735, N493);
buf BUF1 (N1738, N1734);
nor NOR4 (N1739, N1730, N974, N1196, N536);
or OR2 (N1740, N1732, N138);
nand NAND2 (N1741, N1736, N1363);
and AND2 (N1742, N1719, N1001);
or OR3 (N1743, N1738, N902, N1030);
xor XOR2 (N1744, N1722, N1361);
buf BUF1 (N1745, N1740);
xor XOR2 (N1746, N1739, N570);
or OR3 (N1747, N1696, N193, N973);
and AND4 (N1748, N1747, N603, N235, N1487);
and AND4 (N1749, N1742, N1127, N1384, N1563);
buf BUF1 (N1750, N1741);
or OR3 (N1751, N1743, N1268, N999);
and AND2 (N1752, N1737, N776);
xor XOR2 (N1753, N1728, N732);
nand NAND4 (N1754, N1748, N518, N1251, N1009);
nor NOR4 (N1755, N1746, N850, N541, N1542);
nand NAND3 (N1756, N1752, N1502, N1584);
nand NAND2 (N1757, N1755, N45);
nor NOR3 (N1758, N1749, N1098, N739);
or OR4 (N1759, N1757, N583, N1679, N186);
and AND4 (N1760, N1745, N230, N843, N1669);
nor NOR3 (N1761, N1759, N1538, N1693);
or OR2 (N1762, N1753, N451);
buf BUF1 (N1763, N1758);
nor NOR4 (N1764, N1750, N194, N307, N1521);
not NOT1 (N1765, N1762);
and AND3 (N1766, N1727, N206, N1560);
not NOT1 (N1767, N1760);
nand NAND2 (N1768, N1767, N1517);
xor XOR2 (N1769, N1754, N1290);
and AND2 (N1770, N1769, N493);
xor XOR2 (N1771, N1766, N1693);
nand NAND2 (N1772, N1771, N504);
nor NOR3 (N1773, N1756, N1340, N677);
nor NOR4 (N1774, N1772, N1321, N1695, N989);
and AND2 (N1775, N1774, N1004);
buf BUF1 (N1776, N1775);
nand NAND3 (N1777, N1770, N1387, N1489);
or OR4 (N1778, N1765, N588, N720, N506);
not NOT1 (N1779, N1764);
buf BUF1 (N1780, N1751);
or OR3 (N1781, N1744, N301, N1257);
and AND2 (N1782, N1763, N125);
nor NOR2 (N1783, N1777, N1251);
xor XOR2 (N1784, N1761, N1610);
buf BUF1 (N1785, N1780);
xor XOR2 (N1786, N1784, N1503);
not NOT1 (N1787, N1785);
nor NOR3 (N1788, N1782, N603, N228);
buf BUF1 (N1789, N1768);
buf BUF1 (N1790, N1773);
not NOT1 (N1791, N1783);
xor XOR2 (N1792, N1788, N659);
xor XOR2 (N1793, N1779, N21);
nand NAND2 (N1794, N1793, N132);
or OR3 (N1795, N1776, N1506, N1614);
buf BUF1 (N1796, N1791);
buf BUF1 (N1797, N1789);
nand NAND2 (N1798, N1790, N1059);
or OR3 (N1799, N1795, N1139, N1093);
nor NOR2 (N1800, N1781, N1623);
or OR3 (N1801, N1786, N1637, N1080);
buf BUF1 (N1802, N1800);
or OR3 (N1803, N1802, N1205, N228);
nand NAND4 (N1804, N1797, N1259, N12, N230);
nor NOR3 (N1805, N1804, N416, N1307);
nand NAND2 (N1806, N1805, N1173);
or OR3 (N1807, N1803, N1065, N1160);
not NOT1 (N1808, N1792);
not NOT1 (N1809, N1808);
and AND4 (N1810, N1807, N363, N305, N760);
not NOT1 (N1811, N1810);
buf BUF1 (N1812, N1799);
not NOT1 (N1813, N1801);
or OR3 (N1814, N1811, N1139, N1110);
and AND2 (N1815, N1812, N1702);
xor XOR2 (N1816, N1778, N1748);
buf BUF1 (N1817, N1814);
or OR4 (N1818, N1816, N1210, N600, N1482);
nand NAND2 (N1819, N1815, N722);
and AND4 (N1820, N1809, N245, N631, N49);
or OR2 (N1821, N1806, N1371);
not NOT1 (N1822, N1820);
and AND4 (N1823, N1819, N862, N316, N11);
and AND3 (N1824, N1813, N301, N692);
not NOT1 (N1825, N1798);
not NOT1 (N1826, N1787);
and AND2 (N1827, N1821, N1543);
or OR4 (N1828, N1822, N495, N547, N620);
xor XOR2 (N1829, N1826, N1659);
xor XOR2 (N1830, N1794, N1259);
nor NOR2 (N1831, N1817, N360);
and AND4 (N1832, N1829, N1021, N1791, N1357);
or OR2 (N1833, N1825, N1115);
and AND2 (N1834, N1796, N811);
or OR2 (N1835, N1823, N694);
nor NOR4 (N1836, N1830, N1746, N1774, N1650);
and AND4 (N1837, N1828, N953, N329, N267);
nor NOR3 (N1838, N1837, N8, N697);
buf BUF1 (N1839, N1831);
xor XOR2 (N1840, N1832, N533);
nor NOR3 (N1841, N1818, N1603, N1321);
buf BUF1 (N1842, N1834);
or OR3 (N1843, N1838, N207, N558);
and AND3 (N1844, N1842, N1715, N616);
xor XOR2 (N1845, N1835, N145);
xor XOR2 (N1846, N1824, N701);
xor XOR2 (N1847, N1840, N1385);
not NOT1 (N1848, N1836);
nand NAND2 (N1849, N1847, N189);
nand NAND3 (N1850, N1848, N1305, N1046);
and AND3 (N1851, N1846, N150, N661);
xor XOR2 (N1852, N1843, N798);
buf BUF1 (N1853, N1833);
not NOT1 (N1854, N1841);
and AND2 (N1855, N1827, N1554);
buf BUF1 (N1856, N1855);
buf BUF1 (N1857, N1850);
not NOT1 (N1858, N1854);
not NOT1 (N1859, N1851);
xor XOR2 (N1860, N1857, N1394);
and AND2 (N1861, N1839, N1527);
and AND3 (N1862, N1858, N1756, N943);
buf BUF1 (N1863, N1849);
nor NOR2 (N1864, N1860, N450);
not NOT1 (N1865, N1852);
nor NOR2 (N1866, N1856, N770);
and AND4 (N1867, N1866, N1368, N31, N288);
not NOT1 (N1868, N1867);
xor XOR2 (N1869, N1853, N1133);
and AND2 (N1870, N1865, N1708);
or OR3 (N1871, N1845, N758, N1308);
xor XOR2 (N1872, N1859, N1227);
and AND2 (N1873, N1868, N1477);
nand NAND2 (N1874, N1863, N1554);
or OR2 (N1875, N1873, N148);
or OR3 (N1876, N1844, N1812, N1344);
and AND2 (N1877, N1874, N702);
nand NAND4 (N1878, N1864, N1085, N117, N609);
nor NOR2 (N1879, N1875, N883);
or OR2 (N1880, N1869, N1590);
nand NAND2 (N1881, N1870, N1590);
buf BUF1 (N1882, N1880);
nor NOR4 (N1883, N1861, N1105, N212, N1494);
not NOT1 (N1884, N1862);
or OR3 (N1885, N1871, N1088, N1297);
not NOT1 (N1886, N1872);
and AND2 (N1887, N1886, N621);
xor XOR2 (N1888, N1878, N1150);
or OR3 (N1889, N1882, N1832, N1751);
and AND4 (N1890, N1877, N227, N201, N1111);
nand NAND2 (N1891, N1890, N761);
or OR2 (N1892, N1888, N617);
or OR2 (N1893, N1883, N141);
nand NAND3 (N1894, N1887, N1494, N251);
xor XOR2 (N1895, N1884, N1865);
xor XOR2 (N1896, N1893, N280);
and AND4 (N1897, N1876, N1419, N1116, N510);
not NOT1 (N1898, N1879);
not NOT1 (N1899, N1896);
nor NOR2 (N1900, N1881, N1720);
xor XOR2 (N1901, N1892, N898);
or OR2 (N1902, N1899, N1626);
xor XOR2 (N1903, N1900, N1220);
or OR2 (N1904, N1898, N1753);
nand NAND3 (N1905, N1891, N1193, N1762);
or OR3 (N1906, N1897, N11, N1552);
nand NAND2 (N1907, N1894, N1296);
nor NOR3 (N1908, N1904, N688, N966);
xor XOR2 (N1909, N1908, N1246);
and AND2 (N1910, N1889, N828);
not NOT1 (N1911, N1906);
nand NAND2 (N1912, N1907, N1714);
not NOT1 (N1913, N1902);
not NOT1 (N1914, N1913);
nand NAND3 (N1915, N1885, N825, N603);
not NOT1 (N1916, N1914);
not NOT1 (N1917, N1912);
nand NAND3 (N1918, N1916, N926, N1643);
buf BUF1 (N1919, N1918);
buf BUF1 (N1920, N1919);
nand NAND4 (N1921, N1911, N629, N895, N649);
buf BUF1 (N1922, N1901);
and AND2 (N1923, N1903, N173);
xor XOR2 (N1924, N1921, N1196);
buf BUF1 (N1925, N1895);
nand NAND3 (N1926, N1905, N636, N1631);
buf BUF1 (N1927, N1910);
and AND2 (N1928, N1917, N1475);
or OR3 (N1929, N1926, N886, N1434);
nand NAND3 (N1930, N1920, N1, N666);
and AND4 (N1931, N1927, N830, N714, N802);
nand NAND4 (N1932, N1931, N1725, N1777, N398);
nor NOR2 (N1933, N1925, N750);
nor NOR4 (N1934, N1923, N661, N1286, N468);
not NOT1 (N1935, N1934);
not NOT1 (N1936, N1915);
or OR2 (N1937, N1928, N988);
xor XOR2 (N1938, N1924, N144);
and AND3 (N1939, N1935, N1643, N819);
or OR3 (N1940, N1936, N750, N1625);
nor NOR2 (N1941, N1930, N1806);
or OR4 (N1942, N1941, N1771, N804, N1036);
and AND2 (N1943, N1940, N647);
xor XOR2 (N1944, N1937, N1941);
nand NAND2 (N1945, N1929, N860);
or OR3 (N1946, N1943, N736, N1194);
nor NOR4 (N1947, N1942, N630, N980, N736);
nand NAND2 (N1948, N1947, N235);
or OR4 (N1949, N1945, N1876, N695, N955);
xor XOR2 (N1950, N1946, N48);
not NOT1 (N1951, N1909);
and AND2 (N1952, N1950, N1592);
not NOT1 (N1953, N1951);
buf BUF1 (N1954, N1948);
xor XOR2 (N1955, N1922, N280);
buf BUF1 (N1956, N1952);
nand NAND3 (N1957, N1932, N1348, N1597);
nand NAND3 (N1958, N1954, N404, N1135);
nor NOR3 (N1959, N1933, N1077, N1678);
and AND2 (N1960, N1959, N645);
xor XOR2 (N1961, N1938, N83);
nor NOR3 (N1962, N1939, N1575, N600);
buf BUF1 (N1963, N1962);
buf BUF1 (N1964, N1949);
or OR3 (N1965, N1944, N615, N828);
and AND3 (N1966, N1961, N1937, N245);
buf BUF1 (N1967, N1965);
nor NOR3 (N1968, N1963, N1499, N752);
or OR2 (N1969, N1968, N1038);
buf BUF1 (N1970, N1956);
nor NOR4 (N1971, N1957, N1095, N1856, N1969);
nor NOR3 (N1972, N1221, N772, N699);
buf BUF1 (N1973, N1972);
and AND3 (N1974, N1960, N1865, N65);
xor XOR2 (N1975, N1966, N493);
nand NAND4 (N1976, N1974, N337, N1438, N981);
xor XOR2 (N1977, N1975, N856);
xor XOR2 (N1978, N1953, N842);
not NOT1 (N1979, N1976);
buf BUF1 (N1980, N1973);
not NOT1 (N1981, N1955);
and AND4 (N1982, N1977, N114, N1336, N482);
and AND4 (N1983, N1979, N427, N858, N717);
not NOT1 (N1984, N1958);
nand NAND4 (N1985, N1982, N1061, N1650, N1841);
nor NOR4 (N1986, N1983, N1513, N1269, N55);
or OR2 (N1987, N1970, N50);
buf BUF1 (N1988, N1985);
and AND4 (N1989, N1986, N1170, N549, N683);
not NOT1 (N1990, N1971);
buf BUF1 (N1991, N1987);
and AND2 (N1992, N1988, N238);
nor NOR4 (N1993, N1992, N1327, N236, N1746);
xor XOR2 (N1994, N1967, N424);
xor XOR2 (N1995, N1993, N1100);
not NOT1 (N1996, N1964);
buf BUF1 (N1997, N1994);
nor NOR2 (N1998, N1991, N1928);
buf BUF1 (N1999, N1990);
buf BUF1 (N2000, N1980);
nor NOR4 (N2001, N1996, N1364, N356, N1475);
nor NOR2 (N2002, N1984, N808);
and AND2 (N2003, N1995, N136);
xor XOR2 (N2004, N1978, N1494);
xor XOR2 (N2005, N2004, N791);
nand NAND4 (N2006, N1981, N898, N1320, N1086);
nor NOR3 (N2007, N2001, N632, N1984);
nand NAND4 (N2008, N1999, N843, N293, N1979);
not NOT1 (N2009, N2002);
nor NOR3 (N2010, N1997, N213, N1005);
buf BUF1 (N2011, N2008);
nor NOR2 (N2012, N2005, N169);
and AND4 (N2013, N1998, N1702, N1951, N1742);
endmodule