// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N4010,N4011,N3997,N4009,N3994,N3979,N4007,N4004,N4006,N4012;

not NOT1 (N13, N2);
xor XOR2 (N14, N7, N7);
xor XOR2 (N15, N14, N9);
or OR2 (N16, N13, N2);
buf BUF1 (N17, N5);
xor XOR2 (N18, N7, N6);
or OR3 (N19, N12, N17, N14);
and AND3 (N20, N1, N7, N8);
and AND2 (N21, N18, N14);
xor XOR2 (N22, N20, N17);
nor NOR3 (N23, N22, N7, N18);
and AND3 (N24, N5, N4, N4);
nand NAND2 (N25, N5, N23);
or OR4 (N26, N3, N19, N25, N23);
and AND3 (N27, N2, N22, N24);
nor NOR2 (N28, N14, N4);
or OR2 (N29, N12, N23);
nand NAND4 (N30, N29, N6, N20, N29);
buf BUF1 (N31, N23);
xor XOR2 (N32, N20, N3);
and AND4 (N33, N24, N23, N32, N24);
and AND3 (N34, N31, N15, N6);
or OR4 (N35, N14, N24, N11, N11);
or OR3 (N36, N10, N6, N17);
xor XOR2 (N37, N33, N27);
nand NAND2 (N38, N9, N1);
or OR3 (N39, N21, N28, N34);
buf BUF1 (N40, N35);
buf BUF1 (N41, N37);
and AND4 (N42, N19, N3, N13, N35);
not NOT1 (N43, N24);
or OR4 (N44, N42, N16, N37, N35);
buf BUF1 (N45, N8);
nor NOR4 (N46, N36, N10, N7, N17);
nand NAND3 (N47, N44, N17, N21);
buf BUF1 (N48, N43);
xor XOR2 (N49, N46, N1);
or OR4 (N50, N30, N41, N1, N37);
not NOT1 (N51, N20);
xor XOR2 (N52, N47, N8);
xor XOR2 (N53, N48, N31);
buf BUF1 (N54, N53);
xor XOR2 (N55, N51, N22);
buf BUF1 (N56, N45);
or OR2 (N57, N50, N32);
not NOT1 (N58, N54);
nor NOR2 (N59, N49, N27);
not NOT1 (N60, N39);
xor XOR2 (N61, N26, N43);
buf BUF1 (N62, N38);
nand NAND4 (N63, N59, N48, N27, N54);
or OR3 (N64, N40, N56, N12);
or OR3 (N65, N31, N35, N3);
buf BUF1 (N66, N58);
not NOT1 (N67, N61);
nand NAND4 (N68, N66, N16, N20, N23);
and AND3 (N69, N65, N62, N13);
or OR4 (N70, N67, N22, N63, N2);
xor XOR2 (N71, N30, N4);
nor NOR2 (N72, N58, N52);
nor NOR4 (N73, N6, N20, N43, N63);
nor NOR2 (N74, N57, N65);
nor NOR3 (N75, N72, N58, N7);
nand NAND2 (N76, N74, N44);
nand NAND4 (N77, N73, N40, N68, N2);
nand NAND3 (N78, N71, N70, N4);
buf BUF1 (N79, N25);
xor XOR2 (N80, N35, N19);
and AND4 (N81, N75, N61, N60, N5);
not NOT1 (N82, N39);
xor XOR2 (N83, N79, N82);
xor XOR2 (N84, N38, N61);
or OR4 (N85, N80, N25, N81, N65);
xor XOR2 (N86, N48, N69);
not NOT1 (N87, N34);
buf BUF1 (N88, N55);
nor NOR2 (N89, N86, N80);
and AND2 (N90, N76, N68);
xor XOR2 (N91, N78, N71);
buf BUF1 (N92, N77);
xor XOR2 (N93, N90, N64);
and AND3 (N94, N7, N28, N3);
buf BUF1 (N95, N93);
buf BUF1 (N96, N91);
not NOT1 (N97, N94);
nor NOR2 (N98, N83, N2);
xor XOR2 (N99, N87, N80);
nor NOR4 (N100, N98, N73, N30, N10);
and AND2 (N101, N100, N71);
or OR3 (N102, N97, N89, N63);
nand NAND4 (N103, N40, N24, N42, N78);
xor XOR2 (N104, N96, N78);
nand NAND4 (N105, N99, N83, N38, N56);
nor NOR4 (N106, N103, N99, N5, N70);
buf BUF1 (N107, N92);
nand NAND3 (N108, N88, N19, N25);
nand NAND2 (N109, N108, N96);
nor NOR2 (N110, N107, N94);
not NOT1 (N111, N84);
and AND2 (N112, N95, N64);
nand NAND3 (N113, N109, N49, N17);
not NOT1 (N114, N113);
and AND3 (N115, N114, N75, N82);
or OR4 (N116, N115, N53, N21, N104);
nor NOR4 (N117, N35, N65, N72, N67);
nand NAND3 (N118, N111, N39, N35);
xor XOR2 (N119, N105, N69);
and AND4 (N120, N101, N34, N54, N80);
xor XOR2 (N121, N110, N11);
buf BUF1 (N122, N116);
not NOT1 (N123, N119);
nand NAND2 (N124, N118, N35);
nor NOR4 (N125, N124, N4, N14, N76);
xor XOR2 (N126, N121, N121);
nor NOR4 (N127, N123, N16, N49, N11);
or OR2 (N128, N126, N37);
buf BUF1 (N129, N127);
xor XOR2 (N130, N106, N101);
or OR4 (N131, N102, N15, N81, N29);
or OR4 (N132, N122, N39, N99, N96);
nor NOR2 (N133, N125, N12);
nand NAND2 (N134, N130, N11);
nor NOR2 (N135, N85, N14);
not NOT1 (N136, N134);
not NOT1 (N137, N129);
or OR3 (N138, N133, N122, N57);
nand NAND4 (N139, N117, N69, N100, N92);
xor XOR2 (N140, N128, N133);
or OR4 (N141, N137, N69, N17, N1);
or OR3 (N142, N138, N65, N91);
not NOT1 (N143, N141);
xor XOR2 (N144, N120, N56);
not NOT1 (N145, N136);
xor XOR2 (N146, N112, N71);
or OR2 (N147, N132, N123);
xor XOR2 (N148, N139, N68);
not NOT1 (N149, N142);
or OR3 (N150, N148, N59, N53);
xor XOR2 (N151, N147, N6);
not NOT1 (N152, N144);
or OR4 (N153, N152, N115, N74, N95);
or OR3 (N154, N149, N70, N137);
buf BUF1 (N155, N143);
nor NOR2 (N156, N135, N23);
buf BUF1 (N157, N151);
nand NAND4 (N158, N157, N14, N66, N115);
buf BUF1 (N159, N153);
or OR3 (N160, N159, N39, N34);
or OR4 (N161, N146, N113, N33, N145);
not NOT1 (N162, N55);
and AND4 (N163, N158, N23, N97, N114);
xor XOR2 (N164, N160, N32);
or OR3 (N165, N155, N126, N29);
or OR4 (N166, N165, N73, N50, N146);
buf BUF1 (N167, N166);
nand NAND4 (N168, N156, N51, N2, N116);
not NOT1 (N169, N140);
buf BUF1 (N170, N162);
nor NOR4 (N171, N168, N86, N87, N2);
not NOT1 (N172, N163);
nor NOR3 (N173, N171, N46, N141);
buf BUF1 (N174, N161);
nand NAND3 (N175, N167, N131, N169);
nand NAND4 (N176, N161, N51, N60, N159);
xor XOR2 (N177, N75, N47);
and AND3 (N178, N154, N29, N168);
xor XOR2 (N179, N173, N18);
nor NOR4 (N180, N170, N86, N110, N17);
xor XOR2 (N181, N177, N11);
buf BUF1 (N182, N172);
buf BUF1 (N183, N178);
nand NAND2 (N184, N180, N143);
not NOT1 (N185, N181);
nand NAND2 (N186, N150, N59);
xor XOR2 (N187, N183, N153);
not NOT1 (N188, N175);
and AND3 (N189, N185, N82, N144);
buf BUF1 (N190, N176);
or OR2 (N191, N188, N168);
xor XOR2 (N192, N164, N102);
buf BUF1 (N193, N179);
and AND3 (N194, N191, N14, N179);
nand NAND4 (N195, N174, N29, N71, N32);
and AND4 (N196, N187, N78, N62, N25);
buf BUF1 (N197, N190);
nor NOR2 (N198, N192, N69);
nand NAND4 (N199, N197, N83, N92, N48);
nand NAND4 (N200, N193, N196, N150, N90);
xor XOR2 (N201, N158, N5);
and AND4 (N202, N195, N42, N144, N196);
nand NAND2 (N203, N202, N89);
not NOT1 (N204, N194);
and AND2 (N205, N186, N100);
not NOT1 (N206, N203);
buf BUF1 (N207, N198);
not NOT1 (N208, N184);
and AND3 (N209, N189, N79, N69);
and AND2 (N210, N205, N185);
nand NAND3 (N211, N199, N3, N195);
xor XOR2 (N212, N182, N101);
and AND4 (N213, N200, N137, N212, N92);
nand NAND3 (N214, N86, N192, N142);
nor NOR4 (N215, N213, N204, N10, N32);
and AND2 (N216, N28, N20);
nand NAND2 (N217, N201, N47);
not NOT1 (N218, N214);
nand NAND4 (N219, N215, N96, N188, N183);
or OR4 (N220, N209, N124, N172, N213);
not NOT1 (N221, N217);
nand NAND4 (N222, N211, N55, N5, N42);
not NOT1 (N223, N221);
and AND2 (N224, N208, N202);
or OR2 (N225, N224, N93);
xor XOR2 (N226, N220, N93);
xor XOR2 (N227, N206, N179);
nand NAND2 (N228, N216, N202);
and AND2 (N229, N223, N82);
nand NAND4 (N230, N225, N164, N172, N143);
and AND4 (N231, N222, N182, N130, N152);
and AND2 (N232, N229, N64);
nand NAND3 (N233, N230, N96, N176);
buf BUF1 (N234, N210);
buf BUF1 (N235, N232);
xor XOR2 (N236, N218, N158);
buf BUF1 (N237, N228);
nor NOR2 (N238, N207, N175);
nand NAND3 (N239, N227, N203, N215);
xor XOR2 (N240, N235, N89);
xor XOR2 (N241, N234, N182);
buf BUF1 (N242, N226);
and AND4 (N243, N238, N41, N88, N242);
not NOT1 (N244, N48);
and AND2 (N245, N231, N131);
or OR3 (N246, N245, N101, N240);
or OR2 (N247, N194, N174);
or OR4 (N248, N241, N22, N90, N185);
not NOT1 (N249, N219);
or OR2 (N250, N237, N112);
nor NOR3 (N251, N246, N163, N21);
and AND4 (N252, N248, N83, N97, N34);
not NOT1 (N253, N233);
buf BUF1 (N254, N244);
or OR2 (N255, N254, N244);
not NOT1 (N256, N251);
or OR2 (N257, N247, N141);
xor XOR2 (N258, N249, N95);
not NOT1 (N259, N243);
or OR3 (N260, N252, N102, N142);
buf BUF1 (N261, N236);
and AND4 (N262, N239, N182, N84, N204);
nand NAND4 (N263, N253, N40, N119, N109);
buf BUF1 (N264, N260);
nand NAND3 (N265, N263, N97, N237);
buf BUF1 (N266, N261);
buf BUF1 (N267, N255);
nand NAND2 (N268, N264, N45);
xor XOR2 (N269, N257, N36);
nand NAND3 (N270, N265, N49, N202);
and AND4 (N271, N259, N153, N41, N211);
and AND4 (N272, N271, N13, N67, N110);
and AND2 (N273, N269, N28);
nor NOR4 (N274, N272, N42, N4, N227);
not NOT1 (N275, N268);
not NOT1 (N276, N266);
buf BUF1 (N277, N267);
and AND3 (N278, N275, N90, N31);
or OR4 (N279, N276, N212, N254, N42);
not NOT1 (N280, N250);
and AND3 (N281, N258, N55, N78);
not NOT1 (N282, N277);
nand NAND3 (N283, N274, N115, N216);
nand NAND4 (N284, N270, N160, N61, N58);
nor NOR3 (N285, N262, N204, N230);
not NOT1 (N286, N284);
and AND2 (N287, N282, N119);
nor NOR2 (N288, N278, N195);
and AND3 (N289, N287, N97, N5);
and AND3 (N290, N283, N181, N162);
and AND2 (N291, N280, N285);
not NOT1 (N292, N216);
nand NAND3 (N293, N288, N99, N179);
not NOT1 (N294, N273);
xor XOR2 (N295, N290, N170);
or OR4 (N296, N295, N155, N167, N248);
and AND4 (N297, N296, N104, N233, N194);
xor XOR2 (N298, N279, N183);
and AND3 (N299, N291, N121, N57);
xor XOR2 (N300, N299, N132);
and AND4 (N301, N298, N54, N298, N11);
xor XOR2 (N302, N286, N118);
or OR3 (N303, N289, N244, N299);
not NOT1 (N304, N297);
nand NAND4 (N305, N301, N137, N14, N121);
and AND2 (N306, N256, N242);
or OR3 (N307, N281, N31, N34);
buf BUF1 (N308, N293);
nor NOR3 (N309, N294, N154, N76);
not NOT1 (N310, N292);
or OR2 (N311, N305, N187);
and AND4 (N312, N304, N220, N295, N39);
nor NOR2 (N313, N307, N309);
not NOT1 (N314, N256);
or OR3 (N315, N312, N264, N159);
xor XOR2 (N316, N303, N299);
not NOT1 (N317, N300);
not NOT1 (N318, N311);
and AND4 (N319, N306, N174, N52, N250);
nand NAND4 (N320, N314, N197, N134, N256);
xor XOR2 (N321, N316, N198);
or OR4 (N322, N315, N56, N300, N49);
nand NAND4 (N323, N322, N95, N312, N28);
nand NAND2 (N324, N302, N322);
nand NAND3 (N325, N321, N140, N31);
nor NOR3 (N326, N324, N315, N141);
and AND4 (N327, N318, N263, N30, N89);
not NOT1 (N328, N325);
not NOT1 (N329, N317);
nor NOR2 (N330, N313, N325);
nand NAND2 (N331, N310, N95);
not NOT1 (N332, N327);
nand NAND2 (N333, N331, N50);
nor NOR3 (N334, N326, N307, N252);
and AND2 (N335, N329, N220);
or OR4 (N336, N328, N240, N285, N84);
nor NOR4 (N337, N323, N325, N295, N193);
nor NOR4 (N338, N337, N268, N288, N114);
or OR2 (N339, N319, N126);
nor NOR2 (N340, N339, N317);
or OR4 (N341, N333, N171, N65, N14);
or OR2 (N342, N332, N326);
nand NAND2 (N343, N330, N21);
or OR4 (N344, N336, N293, N285, N193);
not NOT1 (N345, N338);
nor NOR2 (N346, N335, N81);
xor XOR2 (N347, N334, N314);
nor NOR2 (N348, N341, N133);
xor XOR2 (N349, N320, N221);
not NOT1 (N350, N348);
or OR4 (N351, N344, N284, N281, N313);
buf BUF1 (N352, N351);
and AND3 (N353, N342, N218, N75);
xor XOR2 (N354, N353, N140);
and AND3 (N355, N350, N41, N22);
and AND2 (N356, N355, N130);
and AND4 (N357, N349, N173, N288, N86);
nor NOR3 (N358, N340, N233, N214);
not NOT1 (N359, N352);
not NOT1 (N360, N358);
buf BUF1 (N361, N359);
not NOT1 (N362, N357);
and AND4 (N363, N356, N210, N74, N268);
nand NAND2 (N364, N308, N101);
and AND4 (N365, N363, N237, N301, N105);
nand NAND3 (N366, N343, N262, N50);
not NOT1 (N367, N366);
nand NAND4 (N368, N347, N273, N344, N224);
not NOT1 (N369, N367);
nand NAND4 (N370, N369, N26, N278, N200);
not NOT1 (N371, N368);
buf BUF1 (N372, N361);
and AND4 (N373, N345, N247, N68, N47);
nand NAND2 (N374, N362, N188);
nor NOR3 (N375, N372, N8, N317);
and AND4 (N376, N346, N315, N335, N311);
xor XOR2 (N377, N375, N257);
buf BUF1 (N378, N376);
nor NOR2 (N379, N373, N127);
nand NAND2 (N380, N360, N354);
not NOT1 (N381, N132);
nor NOR3 (N382, N371, N73, N46);
nor NOR2 (N383, N379, N204);
nand NAND2 (N384, N378, N239);
nand NAND4 (N385, N382, N243, N89, N112);
nor NOR4 (N386, N370, N139, N204, N314);
xor XOR2 (N387, N386, N299);
xor XOR2 (N388, N384, N281);
xor XOR2 (N389, N377, N181);
nor NOR4 (N390, N385, N382, N337, N161);
xor XOR2 (N391, N390, N76);
nand NAND2 (N392, N374, N258);
xor XOR2 (N393, N389, N172);
xor XOR2 (N394, N381, N229);
or OR2 (N395, N383, N151);
not NOT1 (N396, N391);
buf BUF1 (N397, N395);
xor XOR2 (N398, N388, N189);
buf BUF1 (N399, N393);
or OR4 (N400, N365, N215, N341, N50);
and AND2 (N401, N392, N157);
nand NAND4 (N402, N401, N348, N285, N22);
nor NOR4 (N403, N402, N43, N236, N297);
and AND4 (N404, N397, N217, N316, N18);
nand NAND3 (N405, N404, N138, N56);
or OR4 (N406, N364, N129, N293, N227);
nand NAND4 (N407, N405, N394, N354, N272);
nand NAND4 (N408, N401, N301, N28, N18);
and AND2 (N409, N398, N25);
nor NOR4 (N410, N406, N2, N12, N123);
nand NAND3 (N411, N380, N380, N253);
and AND2 (N412, N396, N273);
and AND3 (N413, N408, N410, N221);
and AND2 (N414, N373, N10);
and AND3 (N415, N413, N182, N171);
and AND3 (N416, N403, N127, N175);
or OR4 (N417, N387, N205, N53, N171);
nand NAND2 (N418, N414, N289);
not NOT1 (N419, N400);
or OR4 (N420, N409, N379, N23, N283);
or OR3 (N421, N418, N107, N208);
buf BUF1 (N422, N415);
nor NOR2 (N423, N417, N36);
nand NAND3 (N424, N423, N141, N165);
nand NAND2 (N425, N416, N281);
and AND3 (N426, N424, N265, N274);
xor XOR2 (N427, N411, N324);
nor NOR3 (N428, N422, N50, N300);
not NOT1 (N429, N428);
xor XOR2 (N430, N425, N344);
or OR4 (N431, N429, N277, N203, N264);
nor NOR3 (N432, N430, N351, N165);
nand NAND2 (N433, N427, N432);
nor NOR2 (N434, N204, N270);
and AND2 (N435, N421, N30);
buf BUF1 (N436, N407);
nor NOR3 (N437, N399, N270, N411);
not NOT1 (N438, N431);
nand NAND4 (N439, N436, N294, N160, N430);
nor NOR3 (N440, N412, N376, N269);
and AND3 (N441, N426, N408, N102);
not NOT1 (N442, N439);
and AND4 (N443, N420, N404, N277, N210);
nand NAND4 (N444, N433, N323, N329, N167);
not NOT1 (N445, N438);
buf BUF1 (N446, N440);
nor NOR2 (N447, N446, N394);
nand NAND3 (N448, N444, N267, N81);
xor XOR2 (N449, N419, N169);
nand NAND2 (N450, N437, N429);
and AND2 (N451, N443, N361);
and AND4 (N452, N441, N251, N26, N270);
xor XOR2 (N453, N445, N23);
nor NOR3 (N454, N453, N54, N315);
nand NAND3 (N455, N448, N306, N85);
nand NAND2 (N456, N455, N61);
or OR2 (N457, N434, N76);
buf BUF1 (N458, N450);
and AND3 (N459, N451, N439, N55);
or OR3 (N460, N447, N77, N305);
nand NAND2 (N461, N457, N320);
buf BUF1 (N462, N452);
and AND4 (N463, N461, N14, N383, N198);
nand NAND2 (N464, N435, N275);
and AND4 (N465, N456, N428, N212, N142);
nor NOR4 (N466, N458, N43, N286, N204);
nand NAND2 (N467, N465, N149);
not NOT1 (N468, N462);
or OR4 (N469, N467, N358, N292, N253);
nand NAND3 (N470, N464, N319, N282);
buf BUF1 (N471, N469);
nor NOR2 (N472, N463, N160);
or OR3 (N473, N459, N336, N341);
nor NOR2 (N474, N460, N406);
xor XOR2 (N475, N471, N62);
nor NOR4 (N476, N449, N221, N95, N451);
xor XOR2 (N477, N470, N350);
not NOT1 (N478, N454);
or OR4 (N479, N475, N416, N99, N463);
buf BUF1 (N480, N473);
buf BUF1 (N481, N474);
buf BUF1 (N482, N480);
and AND4 (N483, N468, N138, N349, N410);
nand NAND2 (N484, N483, N80);
nor NOR4 (N485, N484, N333, N278, N52);
or OR2 (N486, N476, N393);
not NOT1 (N487, N482);
buf BUF1 (N488, N481);
buf BUF1 (N489, N488);
xor XOR2 (N490, N478, N377);
not NOT1 (N491, N479);
and AND4 (N492, N491, N431, N337, N49);
buf BUF1 (N493, N485);
buf BUF1 (N494, N477);
and AND3 (N495, N489, N362, N361);
nand NAND3 (N496, N490, N76, N1);
and AND4 (N497, N486, N488, N47, N261);
xor XOR2 (N498, N487, N476);
and AND3 (N499, N498, N476, N400);
nor NOR4 (N500, N442, N376, N413, N310);
or OR3 (N501, N492, N290, N351);
not NOT1 (N502, N500);
or OR2 (N503, N496, N155);
not NOT1 (N504, N499);
nor NOR3 (N505, N502, N145, N325);
and AND3 (N506, N504, N220, N358);
nor NOR4 (N507, N497, N268, N247, N197);
xor XOR2 (N508, N466, N216);
or OR2 (N509, N503, N292);
xor XOR2 (N510, N472, N425);
and AND3 (N511, N508, N331, N489);
buf BUF1 (N512, N495);
not NOT1 (N513, N493);
nor NOR2 (N514, N510, N311);
not NOT1 (N515, N512);
nor NOR3 (N516, N507, N440, N382);
nor NOR4 (N517, N514, N332, N219, N19);
nand NAND4 (N518, N509, N194, N186, N315);
and AND2 (N519, N511, N317);
and AND3 (N520, N513, N502, N117);
or OR3 (N521, N494, N93, N359);
nor NOR2 (N522, N519, N313);
and AND2 (N523, N516, N28);
xor XOR2 (N524, N523, N521);
and AND4 (N525, N271, N393, N289, N104);
or OR2 (N526, N520, N439);
nor NOR3 (N527, N522, N5, N477);
nor NOR4 (N528, N526, N177, N108, N342);
nand NAND4 (N529, N518, N516, N342, N230);
nand NAND3 (N530, N515, N277, N358);
nand NAND3 (N531, N530, N420, N346);
nand NAND3 (N532, N524, N469, N398);
not NOT1 (N533, N527);
not NOT1 (N534, N532);
nor NOR2 (N535, N534, N474);
nand NAND3 (N536, N501, N441, N191);
xor XOR2 (N537, N506, N353);
not NOT1 (N538, N505);
buf BUF1 (N539, N538);
not NOT1 (N540, N528);
nor NOR3 (N541, N517, N307, N183);
and AND4 (N542, N536, N359, N347, N382);
not NOT1 (N543, N525);
or OR4 (N544, N531, N23, N347, N386);
not NOT1 (N545, N533);
nor NOR4 (N546, N544, N211, N48, N195);
or OR2 (N547, N543, N284);
and AND2 (N548, N537, N172);
nand NAND3 (N549, N540, N103, N535);
not NOT1 (N550, N180);
nand NAND4 (N551, N529, N427, N217, N484);
buf BUF1 (N552, N545);
nand NAND2 (N553, N549, N418);
buf BUF1 (N554, N552);
nor NOR2 (N555, N551, N413);
buf BUF1 (N556, N554);
xor XOR2 (N557, N539, N111);
not NOT1 (N558, N541);
nand NAND2 (N559, N550, N386);
nor NOR4 (N560, N547, N435, N123, N467);
and AND3 (N561, N555, N522, N466);
not NOT1 (N562, N553);
xor XOR2 (N563, N556, N182);
xor XOR2 (N564, N562, N25);
buf BUF1 (N565, N560);
buf BUF1 (N566, N542);
not NOT1 (N567, N559);
or OR2 (N568, N557, N175);
xor XOR2 (N569, N561, N513);
or OR3 (N570, N566, N76, N430);
or OR3 (N571, N570, N136, N456);
nand NAND3 (N572, N565, N117, N99);
not NOT1 (N573, N568);
and AND3 (N574, N567, N501, N299);
nand NAND4 (N575, N558, N28, N37, N522);
not NOT1 (N576, N574);
nand NAND4 (N577, N546, N94, N379, N94);
or OR2 (N578, N577, N237);
nor NOR4 (N579, N571, N275, N90, N313);
nand NAND4 (N580, N563, N52, N500, N312);
and AND2 (N581, N578, N383);
nand NAND3 (N582, N569, N124, N91);
nand NAND3 (N583, N575, N390, N252);
or OR2 (N584, N582, N494);
nand NAND3 (N585, N572, N512, N489);
and AND2 (N586, N580, N117);
and AND4 (N587, N584, N531, N306, N429);
and AND3 (N588, N548, N553, N255);
xor XOR2 (N589, N581, N193);
and AND4 (N590, N579, N322, N149, N379);
xor XOR2 (N591, N576, N285);
xor XOR2 (N592, N585, N521);
nand NAND4 (N593, N592, N502, N249, N213);
nand NAND4 (N594, N564, N384, N167, N314);
nand NAND3 (N595, N593, N111, N350);
nand NAND4 (N596, N591, N391, N444, N578);
or OR3 (N597, N594, N363, N268);
nor NOR3 (N598, N586, N236, N542);
xor XOR2 (N599, N595, N126);
xor XOR2 (N600, N583, N277);
xor XOR2 (N601, N598, N512);
buf BUF1 (N602, N589);
buf BUF1 (N603, N602);
nand NAND4 (N604, N590, N37, N454, N505);
nand NAND2 (N605, N573, N160);
not NOT1 (N606, N587);
nor NOR2 (N607, N596, N124);
nand NAND4 (N608, N607, N197, N552, N445);
nand NAND3 (N609, N603, N31, N212);
nand NAND3 (N610, N604, N473, N231);
buf BUF1 (N611, N599);
nand NAND4 (N612, N600, N449, N213, N26);
nor NOR2 (N613, N601, N425);
buf BUF1 (N614, N611);
nand NAND4 (N615, N606, N87, N63, N327);
xor XOR2 (N616, N612, N462);
buf BUF1 (N617, N609);
nor NOR4 (N618, N588, N104, N443, N511);
and AND2 (N619, N618, N589);
not NOT1 (N620, N610);
not NOT1 (N621, N613);
and AND2 (N622, N614, N49);
buf BUF1 (N623, N605);
and AND3 (N624, N620, N317, N15);
buf BUF1 (N625, N617);
nand NAND2 (N626, N619, N585);
buf BUF1 (N627, N626);
xor XOR2 (N628, N622, N38);
or OR2 (N629, N623, N350);
nor NOR4 (N630, N629, N515, N295, N5);
nor NOR4 (N631, N597, N439, N33, N415);
xor XOR2 (N632, N621, N433);
nor NOR4 (N633, N625, N197, N506, N31);
nor NOR4 (N634, N631, N262, N206, N384);
buf BUF1 (N635, N624);
not NOT1 (N636, N635);
nor NOR2 (N637, N627, N176);
nor NOR2 (N638, N628, N502);
buf BUF1 (N639, N615);
buf BUF1 (N640, N637);
nor NOR3 (N641, N633, N37, N145);
buf BUF1 (N642, N636);
nand NAND2 (N643, N608, N36);
buf BUF1 (N644, N642);
buf BUF1 (N645, N632);
and AND3 (N646, N616, N562, N162);
xor XOR2 (N647, N638, N149);
not NOT1 (N648, N645);
buf BUF1 (N649, N646);
or OR4 (N650, N647, N526, N347, N251);
nor NOR3 (N651, N630, N380, N104);
nor NOR3 (N652, N643, N426, N401);
nand NAND3 (N653, N651, N507, N582);
not NOT1 (N654, N641);
nor NOR4 (N655, N644, N188, N96, N385);
nor NOR3 (N656, N648, N112, N286);
not NOT1 (N657, N654);
xor XOR2 (N658, N655, N148);
nand NAND2 (N659, N650, N293);
nand NAND4 (N660, N656, N167, N527, N530);
nor NOR3 (N661, N657, N266, N242);
nor NOR4 (N662, N640, N551, N608, N30);
xor XOR2 (N663, N639, N325);
nand NAND4 (N664, N662, N515, N48, N32);
nand NAND3 (N665, N649, N575, N601);
and AND2 (N666, N663, N28);
nor NOR3 (N667, N634, N247, N361);
or OR3 (N668, N666, N160, N610);
nand NAND3 (N669, N652, N598, N56);
and AND3 (N670, N659, N235, N44);
and AND2 (N671, N658, N160);
nand NAND4 (N672, N668, N297, N417, N594);
buf BUF1 (N673, N653);
and AND4 (N674, N669, N483, N160, N446);
nand NAND3 (N675, N665, N283, N582);
nor NOR2 (N676, N674, N152);
or OR4 (N677, N671, N659, N116, N673);
nand NAND3 (N678, N171, N398, N635);
not NOT1 (N679, N676);
and AND4 (N680, N664, N72, N178, N353);
buf BUF1 (N681, N670);
or OR2 (N682, N672, N307);
nor NOR2 (N683, N677, N437);
nor NOR2 (N684, N681, N666);
buf BUF1 (N685, N667);
buf BUF1 (N686, N682);
or OR3 (N687, N686, N38, N233);
xor XOR2 (N688, N678, N362);
not NOT1 (N689, N683);
buf BUF1 (N690, N660);
or OR2 (N691, N687, N332);
and AND4 (N692, N688, N453, N491, N575);
not NOT1 (N693, N692);
nor NOR4 (N694, N680, N7, N323, N109);
and AND4 (N695, N690, N165, N637, N178);
not NOT1 (N696, N675);
not NOT1 (N697, N684);
xor XOR2 (N698, N697, N328);
nor NOR4 (N699, N696, N229, N539, N546);
nor NOR2 (N700, N685, N309);
buf BUF1 (N701, N698);
nor NOR4 (N702, N693, N312, N474, N269);
not NOT1 (N703, N689);
xor XOR2 (N704, N691, N210);
nand NAND2 (N705, N679, N607);
and AND2 (N706, N701, N179);
xor XOR2 (N707, N700, N95);
and AND4 (N708, N702, N688, N149, N247);
and AND4 (N709, N661, N676, N455, N584);
buf BUF1 (N710, N709);
and AND3 (N711, N694, N125, N195);
xor XOR2 (N712, N708, N288);
not NOT1 (N713, N707);
not NOT1 (N714, N705);
nor NOR2 (N715, N712, N523);
xor XOR2 (N716, N704, N309);
xor XOR2 (N717, N699, N380);
and AND3 (N718, N711, N204, N449);
xor XOR2 (N719, N703, N382);
or OR4 (N720, N695, N244, N109, N423);
or OR3 (N721, N719, N316, N76);
xor XOR2 (N722, N710, N78);
xor XOR2 (N723, N706, N252);
and AND4 (N724, N722, N531, N342, N519);
or OR3 (N725, N717, N31, N11);
and AND2 (N726, N720, N66);
buf BUF1 (N727, N715);
nor NOR2 (N728, N713, N209);
nand NAND3 (N729, N716, N434, N619);
nor NOR4 (N730, N728, N459, N650, N40);
xor XOR2 (N731, N725, N388);
nor NOR2 (N732, N721, N22);
and AND2 (N733, N714, N118);
xor XOR2 (N734, N727, N502);
nand NAND4 (N735, N718, N311, N92, N578);
nor NOR3 (N736, N723, N365, N670);
xor XOR2 (N737, N734, N244);
nor NOR2 (N738, N736, N244);
xor XOR2 (N739, N729, N111);
xor XOR2 (N740, N730, N101);
and AND3 (N741, N737, N457, N534);
or OR2 (N742, N738, N691);
or OR3 (N743, N726, N590, N58);
nor NOR4 (N744, N743, N10, N404, N90);
nand NAND2 (N745, N744, N327);
xor XOR2 (N746, N739, N219);
nor NOR3 (N747, N745, N108, N577);
nand NAND4 (N748, N742, N39, N270, N240);
not NOT1 (N749, N746);
nand NAND2 (N750, N747, N134);
or OR2 (N751, N733, N3);
not NOT1 (N752, N751);
or OR2 (N753, N740, N565);
not NOT1 (N754, N748);
and AND3 (N755, N724, N544, N745);
or OR2 (N756, N735, N582);
xor XOR2 (N757, N752, N273);
not NOT1 (N758, N755);
nor NOR2 (N759, N749, N559);
xor XOR2 (N760, N759, N148);
nand NAND2 (N761, N731, N626);
or OR4 (N762, N758, N595, N544, N661);
and AND4 (N763, N757, N752, N216, N514);
buf BUF1 (N764, N753);
or OR2 (N765, N762, N715);
xor XOR2 (N766, N741, N315);
xor XOR2 (N767, N754, N479);
or OR3 (N768, N760, N621, N552);
nor NOR3 (N769, N767, N392, N671);
nand NAND4 (N770, N766, N345, N441, N26);
buf BUF1 (N771, N769);
nor NOR4 (N772, N763, N656, N643, N685);
xor XOR2 (N773, N772, N561);
xor XOR2 (N774, N765, N370);
nor NOR2 (N775, N773, N760);
not NOT1 (N776, N756);
xor XOR2 (N777, N761, N399);
not NOT1 (N778, N777);
nor NOR4 (N779, N764, N710, N690, N146);
or OR2 (N780, N779, N455);
nand NAND3 (N781, N776, N217, N513);
not NOT1 (N782, N778);
nand NAND3 (N783, N732, N776, N103);
nor NOR2 (N784, N770, N240);
and AND4 (N785, N768, N762, N335, N673);
and AND3 (N786, N771, N147, N662);
xor XOR2 (N787, N774, N272);
xor XOR2 (N788, N781, N633);
not NOT1 (N789, N780);
nor NOR4 (N790, N775, N265, N243, N476);
buf BUF1 (N791, N750);
or OR4 (N792, N784, N382, N737, N153);
and AND2 (N793, N782, N525);
and AND3 (N794, N789, N54, N772);
and AND3 (N795, N791, N68, N770);
not NOT1 (N796, N785);
and AND3 (N797, N795, N278, N309);
buf BUF1 (N798, N790);
not NOT1 (N799, N786);
buf BUF1 (N800, N796);
nand NAND2 (N801, N797, N330);
not NOT1 (N802, N800);
nand NAND4 (N803, N801, N756, N256, N736);
buf BUF1 (N804, N799);
xor XOR2 (N805, N787, N13);
not NOT1 (N806, N783);
or OR4 (N807, N805, N176, N602, N532);
or OR2 (N808, N793, N211);
and AND2 (N809, N788, N39);
buf BUF1 (N810, N794);
nand NAND2 (N811, N792, N42);
nand NAND3 (N812, N798, N217, N140);
or OR3 (N813, N804, N726, N650);
xor XOR2 (N814, N811, N145);
and AND3 (N815, N807, N293, N243);
not NOT1 (N816, N803);
buf BUF1 (N817, N806);
and AND3 (N818, N815, N195, N287);
nor NOR3 (N819, N802, N630, N148);
not NOT1 (N820, N817);
and AND2 (N821, N809, N160);
nand NAND2 (N822, N816, N281);
buf BUF1 (N823, N810);
not NOT1 (N824, N814);
or OR2 (N825, N824, N69);
nand NAND2 (N826, N822, N208);
xor XOR2 (N827, N821, N680);
nor NOR3 (N828, N826, N87, N511);
nand NAND2 (N829, N808, N646);
xor XOR2 (N830, N823, N218);
buf BUF1 (N831, N830);
buf BUF1 (N832, N812);
nor NOR3 (N833, N832, N675, N231);
not NOT1 (N834, N831);
xor XOR2 (N835, N827, N750);
or OR2 (N836, N835, N762);
or OR2 (N837, N813, N433);
nor NOR4 (N838, N834, N763, N763, N207);
nand NAND3 (N839, N828, N338, N758);
nand NAND4 (N840, N825, N592, N65, N494);
nor NOR2 (N841, N829, N397);
not NOT1 (N842, N837);
not NOT1 (N843, N833);
or OR4 (N844, N818, N627, N357, N807);
xor XOR2 (N845, N836, N474);
buf BUF1 (N846, N845);
buf BUF1 (N847, N844);
xor XOR2 (N848, N847, N503);
nor NOR3 (N849, N841, N122, N530);
or OR4 (N850, N839, N816, N91, N407);
or OR3 (N851, N838, N462, N239);
or OR4 (N852, N840, N760, N437, N578);
or OR2 (N853, N848, N410);
nor NOR2 (N854, N846, N651);
not NOT1 (N855, N820);
nor NOR2 (N856, N850, N595);
buf BUF1 (N857, N849);
not NOT1 (N858, N842);
buf BUF1 (N859, N851);
nand NAND3 (N860, N852, N509, N719);
nor NOR2 (N861, N856, N355);
nor NOR3 (N862, N843, N770, N843);
buf BUF1 (N863, N819);
or OR3 (N864, N860, N181, N378);
not NOT1 (N865, N859);
nor NOR2 (N866, N863, N524);
nand NAND3 (N867, N862, N133, N755);
buf BUF1 (N868, N865);
and AND4 (N869, N868, N669, N29, N64);
or OR2 (N870, N857, N167);
nor NOR4 (N871, N861, N751, N338, N155);
xor XOR2 (N872, N858, N850);
or OR2 (N873, N867, N692);
nand NAND3 (N874, N866, N382, N74);
xor XOR2 (N875, N873, N298);
nand NAND4 (N876, N869, N846, N789, N621);
or OR3 (N877, N876, N737, N738);
not NOT1 (N878, N874);
nor NOR4 (N879, N875, N570, N810, N859);
or OR3 (N880, N871, N250, N543);
and AND3 (N881, N877, N235, N453);
buf BUF1 (N882, N855);
nor NOR2 (N883, N854, N116);
nand NAND4 (N884, N880, N595, N689, N466);
and AND4 (N885, N883, N722, N475, N558);
buf BUF1 (N886, N882);
buf BUF1 (N887, N881);
and AND2 (N888, N878, N575);
nand NAND2 (N889, N870, N99);
buf BUF1 (N890, N888);
nand NAND4 (N891, N879, N483, N401, N341);
buf BUF1 (N892, N885);
buf BUF1 (N893, N892);
and AND2 (N894, N891, N563);
not NOT1 (N895, N886);
not NOT1 (N896, N864);
not NOT1 (N897, N895);
nor NOR3 (N898, N896, N790, N802);
nor NOR3 (N899, N893, N389, N598);
nand NAND2 (N900, N872, N580);
and AND4 (N901, N890, N604, N654, N308);
buf BUF1 (N902, N894);
xor XOR2 (N903, N897, N433);
or OR4 (N904, N898, N611, N103, N57);
and AND3 (N905, N904, N674, N445);
nand NAND2 (N906, N901, N707);
nand NAND4 (N907, N853, N206, N418, N267);
nor NOR3 (N908, N884, N806, N13);
xor XOR2 (N909, N889, N478);
or OR4 (N910, N899, N329, N644, N98);
nand NAND3 (N911, N905, N282, N800);
and AND4 (N912, N908, N227, N463, N616);
or OR3 (N913, N912, N781, N610);
buf BUF1 (N914, N911);
not NOT1 (N915, N910);
buf BUF1 (N916, N887);
xor XOR2 (N917, N907, N47);
nor NOR2 (N918, N915, N155);
or OR2 (N919, N916, N531);
nor NOR4 (N920, N919, N164, N220, N156);
xor XOR2 (N921, N902, N210);
not NOT1 (N922, N906);
or OR4 (N923, N909, N569, N693, N496);
buf BUF1 (N924, N917);
buf BUF1 (N925, N924);
buf BUF1 (N926, N922);
xor XOR2 (N927, N903, N419);
or OR2 (N928, N923, N836);
or OR4 (N929, N926, N659, N742, N199);
nor NOR4 (N930, N928, N350, N471, N161);
or OR2 (N931, N913, N924);
buf BUF1 (N932, N930);
or OR2 (N933, N929, N557);
or OR2 (N934, N920, N492);
buf BUF1 (N935, N900);
buf BUF1 (N936, N934);
not NOT1 (N937, N932);
xor XOR2 (N938, N918, N39);
buf BUF1 (N939, N931);
or OR3 (N940, N937, N552, N730);
nand NAND4 (N941, N935, N600, N819, N323);
xor XOR2 (N942, N933, N861);
not NOT1 (N943, N927);
not NOT1 (N944, N925);
buf BUF1 (N945, N944);
and AND3 (N946, N942, N60, N760);
buf BUF1 (N947, N943);
nor NOR3 (N948, N938, N469, N139);
nor NOR3 (N949, N939, N492, N706);
nand NAND3 (N950, N936, N738, N168);
or OR3 (N951, N948, N445, N139);
or OR4 (N952, N940, N49, N635, N460);
xor XOR2 (N953, N921, N435);
xor XOR2 (N954, N941, N260);
nor NOR4 (N955, N954, N668, N114, N82);
buf BUF1 (N956, N945);
and AND2 (N957, N950, N452);
nand NAND2 (N958, N955, N868);
buf BUF1 (N959, N956);
xor XOR2 (N960, N958, N280);
nand NAND4 (N961, N951, N846, N563, N210);
buf BUF1 (N962, N959);
not NOT1 (N963, N960);
not NOT1 (N964, N962);
xor XOR2 (N965, N961, N740);
buf BUF1 (N966, N964);
and AND3 (N967, N952, N676, N948);
not NOT1 (N968, N946);
buf BUF1 (N969, N947);
nand NAND2 (N970, N963, N222);
buf BUF1 (N971, N968);
and AND3 (N972, N957, N208, N755);
and AND4 (N973, N914, N579, N456, N45);
or OR3 (N974, N969, N193, N654);
buf BUF1 (N975, N973);
nand NAND2 (N976, N970, N513);
xor XOR2 (N977, N953, N384);
xor XOR2 (N978, N974, N444);
nor NOR4 (N979, N966, N968, N297, N351);
and AND4 (N980, N976, N324, N867, N533);
nor NOR4 (N981, N971, N850, N373, N755);
buf BUF1 (N982, N975);
and AND2 (N983, N977, N562);
and AND4 (N984, N980, N856, N423, N154);
and AND2 (N985, N979, N660);
not NOT1 (N986, N985);
buf BUF1 (N987, N978);
xor XOR2 (N988, N967, N687);
xor XOR2 (N989, N981, N557);
nor NOR2 (N990, N949, N125);
nand NAND3 (N991, N982, N971, N457);
not NOT1 (N992, N989);
buf BUF1 (N993, N990);
xor XOR2 (N994, N991, N660);
buf BUF1 (N995, N984);
xor XOR2 (N996, N988, N524);
and AND2 (N997, N986, N963);
nor NOR3 (N998, N996, N431, N802);
nand NAND4 (N999, N995, N138, N309, N430);
nand NAND4 (N1000, N998, N569, N414, N168);
nand NAND2 (N1001, N992, N943);
or OR4 (N1002, N1000, N63, N547, N236);
and AND4 (N1003, N999, N967, N91, N978);
and AND3 (N1004, N965, N607, N61);
or OR3 (N1005, N1001, N65, N691);
nand NAND4 (N1006, N1004, N360, N534, N568);
nor NOR2 (N1007, N997, N266);
nand NAND2 (N1008, N987, N685);
and AND3 (N1009, N1003, N869, N462);
or OR4 (N1010, N1006, N241, N128, N327);
nand NAND4 (N1011, N1002, N63, N313, N970);
or OR2 (N1012, N1009, N931);
nor NOR3 (N1013, N993, N752, N67);
nand NAND3 (N1014, N1011, N681, N170);
not NOT1 (N1015, N1012);
nor NOR4 (N1016, N972, N986, N277, N433);
or OR3 (N1017, N1016, N592, N326);
nand NAND2 (N1018, N1014, N364);
and AND4 (N1019, N1013, N456, N556, N285);
xor XOR2 (N1020, N1017, N813);
not NOT1 (N1021, N1019);
not NOT1 (N1022, N1020);
nand NAND3 (N1023, N1008, N128, N696);
or OR3 (N1024, N1005, N224, N474);
or OR3 (N1025, N1023, N855, N79);
not NOT1 (N1026, N1021);
buf BUF1 (N1027, N1018);
buf BUF1 (N1028, N1022);
xor XOR2 (N1029, N994, N387);
or OR2 (N1030, N1007, N630);
and AND3 (N1031, N1026, N472, N423);
xor XOR2 (N1032, N1010, N50);
nor NOR2 (N1033, N983, N1027);
nor NOR3 (N1034, N465, N409, N515);
and AND3 (N1035, N1032, N501, N914);
xor XOR2 (N1036, N1015, N80);
nor NOR4 (N1037, N1024, N726, N110, N831);
or OR4 (N1038, N1034, N1026, N918, N818);
or OR4 (N1039, N1037, N152, N914, N978);
and AND2 (N1040, N1028, N578);
and AND4 (N1041, N1029, N720, N283, N960);
or OR2 (N1042, N1041, N303);
buf BUF1 (N1043, N1042);
buf BUF1 (N1044, N1031);
nand NAND4 (N1045, N1025, N381, N852, N284);
and AND3 (N1046, N1035, N37, N457);
and AND3 (N1047, N1045, N79, N798);
not NOT1 (N1048, N1030);
nor NOR2 (N1049, N1046, N714);
not NOT1 (N1050, N1040);
or OR3 (N1051, N1038, N654, N983);
nand NAND4 (N1052, N1036, N785, N17, N778);
xor XOR2 (N1053, N1043, N176);
not NOT1 (N1054, N1050);
buf BUF1 (N1055, N1039);
and AND2 (N1056, N1051, N1049);
and AND2 (N1057, N114, N946);
xor XOR2 (N1058, N1048, N536);
or OR2 (N1059, N1053, N6);
buf BUF1 (N1060, N1047);
nand NAND2 (N1061, N1054, N619);
xor XOR2 (N1062, N1059, N776);
nand NAND4 (N1063, N1057, N232, N683, N959);
and AND2 (N1064, N1061, N161);
or OR3 (N1065, N1044, N789, N1031);
nand NAND4 (N1066, N1064, N879, N122, N941);
and AND3 (N1067, N1065, N578, N243);
not NOT1 (N1068, N1063);
xor XOR2 (N1069, N1052, N728);
buf BUF1 (N1070, N1069);
xor XOR2 (N1071, N1066, N518);
nand NAND2 (N1072, N1062, N679);
nand NAND4 (N1073, N1058, N566, N862, N152);
nand NAND3 (N1074, N1068, N833, N954);
and AND4 (N1075, N1073, N886, N924, N826);
or OR4 (N1076, N1071, N822, N571, N224);
and AND3 (N1077, N1070, N1035, N26);
buf BUF1 (N1078, N1055);
nor NOR2 (N1079, N1060, N1075);
buf BUF1 (N1080, N639);
and AND2 (N1081, N1076, N105);
nor NOR4 (N1082, N1077, N589, N40, N642);
xor XOR2 (N1083, N1033, N60);
buf BUF1 (N1084, N1072);
buf BUF1 (N1085, N1082);
not NOT1 (N1086, N1083);
not NOT1 (N1087, N1084);
not NOT1 (N1088, N1078);
nand NAND3 (N1089, N1086, N1, N275);
not NOT1 (N1090, N1080);
xor XOR2 (N1091, N1074, N280);
not NOT1 (N1092, N1087);
not NOT1 (N1093, N1091);
and AND4 (N1094, N1090, N1052, N492, N177);
and AND2 (N1095, N1089, N8);
or OR3 (N1096, N1093, N967, N983);
or OR2 (N1097, N1079, N556);
nor NOR3 (N1098, N1097, N156, N137);
and AND2 (N1099, N1067, N58);
buf BUF1 (N1100, N1094);
nand NAND2 (N1101, N1099, N662);
nor NOR2 (N1102, N1101, N642);
and AND4 (N1103, N1098, N767, N62, N1083);
nor NOR3 (N1104, N1095, N871, N633);
nor NOR3 (N1105, N1088, N480, N191);
buf BUF1 (N1106, N1105);
not NOT1 (N1107, N1100);
and AND4 (N1108, N1081, N981, N959, N324);
and AND4 (N1109, N1104, N614, N25, N426);
not NOT1 (N1110, N1096);
buf BUF1 (N1111, N1085);
or OR3 (N1112, N1107, N106, N1055);
nor NOR3 (N1113, N1102, N362, N75);
xor XOR2 (N1114, N1111, N732);
and AND2 (N1115, N1114, N1050);
buf BUF1 (N1116, N1056);
nand NAND2 (N1117, N1113, N538);
nor NOR3 (N1118, N1115, N945, N771);
and AND2 (N1119, N1117, N766);
nor NOR3 (N1120, N1108, N315, N930);
xor XOR2 (N1121, N1106, N32);
and AND3 (N1122, N1110, N892, N126);
nor NOR4 (N1123, N1118, N284, N503, N836);
nor NOR3 (N1124, N1116, N723, N577);
or OR2 (N1125, N1109, N783);
and AND4 (N1126, N1121, N673, N620, N1038);
or OR4 (N1127, N1119, N757, N13, N940);
buf BUF1 (N1128, N1103);
nor NOR3 (N1129, N1123, N354, N827);
or OR2 (N1130, N1120, N817);
nand NAND3 (N1131, N1092, N412, N383);
not NOT1 (N1132, N1130);
and AND3 (N1133, N1128, N39, N217);
buf BUF1 (N1134, N1129);
buf BUF1 (N1135, N1124);
nor NOR4 (N1136, N1126, N955, N1019, N732);
nor NOR2 (N1137, N1112, N199);
not NOT1 (N1138, N1134);
or OR2 (N1139, N1122, N527);
and AND3 (N1140, N1136, N1139, N970);
or OR3 (N1141, N933, N317, N438);
or OR4 (N1142, N1137, N513, N976, N302);
nor NOR4 (N1143, N1142, N29, N455, N831);
and AND4 (N1144, N1141, N504, N895, N252);
xor XOR2 (N1145, N1127, N751);
and AND3 (N1146, N1145, N891, N109);
xor XOR2 (N1147, N1140, N1101);
not NOT1 (N1148, N1144);
not NOT1 (N1149, N1132);
xor XOR2 (N1150, N1133, N37);
nor NOR3 (N1151, N1147, N912, N958);
xor XOR2 (N1152, N1125, N946);
not NOT1 (N1153, N1146);
not NOT1 (N1154, N1153);
and AND3 (N1155, N1152, N606, N592);
buf BUF1 (N1156, N1138);
nor NOR4 (N1157, N1150, N941, N982, N931);
nand NAND3 (N1158, N1149, N1082, N978);
nand NAND4 (N1159, N1151, N706, N179, N524);
xor XOR2 (N1160, N1157, N891);
nand NAND4 (N1161, N1148, N703, N43, N139);
buf BUF1 (N1162, N1158);
or OR2 (N1163, N1161, N177);
and AND3 (N1164, N1154, N1025, N448);
and AND2 (N1165, N1156, N766);
xor XOR2 (N1166, N1164, N904);
and AND4 (N1167, N1135, N850, N569, N281);
nor NOR2 (N1168, N1143, N130);
xor XOR2 (N1169, N1155, N809);
and AND4 (N1170, N1131, N682, N840, N765);
not NOT1 (N1171, N1160);
and AND2 (N1172, N1169, N777);
xor XOR2 (N1173, N1163, N524);
and AND3 (N1174, N1173, N102, N967);
not NOT1 (N1175, N1171);
not NOT1 (N1176, N1168);
xor XOR2 (N1177, N1176, N246);
nor NOR3 (N1178, N1170, N652, N686);
and AND2 (N1179, N1162, N694);
nand NAND4 (N1180, N1165, N750, N544, N599);
not NOT1 (N1181, N1167);
nand NAND3 (N1182, N1175, N10, N534);
and AND4 (N1183, N1178, N1056, N599, N938);
nand NAND2 (N1184, N1174, N251);
xor XOR2 (N1185, N1180, N474);
nor NOR2 (N1186, N1181, N257);
and AND2 (N1187, N1177, N1152);
not NOT1 (N1188, N1187);
or OR4 (N1189, N1188, N719, N619, N828);
xor XOR2 (N1190, N1182, N108);
nand NAND4 (N1191, N1190, N816, N940, N315);
buf BUF1 (N1192, N1183);
xor XOR2 (N1193, N1185, N1095);
nand NAND2 (N1194, N1186, N396);
not NOT1 (N1195, N1166);
buf BUF1 (N1196, N1179);
buf BUF1 (N1197, N1192);
nand NAND4 (N1198, N1197, N1096, N231, N736);
and AND3 (N1199, N1184, N203, N653);
or OR3 (N1200, N1195, N250, N492);
xor XOR2 (N1201, N1191, N805);
and AND2 (N1202, N1198, N290);
xor XOR2 (N1203, N1189, N417);
nor NOR4 (N1204, N1159, N25, N707, N77);
or OR3 (N1205, N1196, N979, N547);
not NOT1 (N1206, N1202);
not NOT1 (N1207, N1199);
not NOT1 (N1208, N1193);
nand NAND3 (N1209, N1172, N919, N715);
and AND4 (N1210, N1207, N462, N357, N363);
and AND4 (N1211, N1208, N270, N908, N555);
or OR3 (N1212, N1206, N941, N79);
xor XOR2 (N1213, N1200, N407);
and AND2 (N1214, N1203, N631);
and AND3 (N1215, N1213, N440, N698);
buf BUF1 (N1216, N1212);
buf BUF1 (N1217, N1216);
not NOT1 (N1218, N1194);
not NOT1 (N1219, N1217);
and AND2 (N1220, N1214, N964);
or OR2 (N1221, N1209, N647);
and AND4 (N1222, N1205, N425, N904, N860);
nor NOR2 (N1223, N1222, N356);
nor NOR3 (N1224, N1201, N850, N898);
buf BUF1 (N1225, N1215);
nor NOR3 (N1226, N1204, N32, N587);
nor NOR2 (N1227, N1221, N1087);
nand NAND4 (N1228, N1223, N145, N1144, N1219);
and AND3 (N1229, N687, N574, N1047);
not NOT1 (N1230, N1224);
nor NOR2 (N1231, N1228, N303);
or OR3 (N1232, N1211, N982, N925);
or OR4 (N1233, N1210, N312, N235, N191);
nand NAND4 (N1234, N1229, N481, N1029, N819);
and AND2 (N1235, N1233, N821);
and AND4 (N1236, N1235, N1156, N886, N71);
xor XOR2 (N1237, N1220, N615);
or OR4 (N1238, N1218, N341, N996, N930);
xor XOR2 (N1239, N1230, N1141);
or OR3 (N1240, N1232, N615, N808);
nand NAND2 (N1241, N1239, N1128);
nand NAND2 (N1242, N1236, N649);
or OR2 (N1243, N1227, N478);
and AND3 (N1244, N1237, N116, N646);
not NOT1 (N1245, N1241);
or OR4 (N1246, N1240, N275, N451, N981);
nand NAND3 (N1247, N1238, N144, N593);
nand NAND2 (N1248, N1247, N348);
nor NOR3 (N1249, N1244, N121, N1193);
xor XOR2 (N1250, N1245, N1225);
not NOT1 (N1251, N389);
nand NAND3 (N1252, N1246, N367, N303);
not NOT1 (N1253, N1231);
xor XOR2 (N1254, N1234, N262);
not NOT1 (N1255, N1248);
and AND4 (N1256, N1249, N665, N963, N195);
and AND3 (N1257, N1254, N305, N255);
nor NOR4 (N1258, N1253, N429, N98, N274);
xor XOR2 (N1259, N1250, N589);
nand NAND2 (N1260, N1259, N1008);
not NOT1 (N1261, N1257);
not NOT1 (N1262, N1242);
or OR4 (N1263, N1262, N1204, N557, N675);
and AND4 (N1264, N1263, N316, N800, N210);
not NOT1 (N1265, N1260);
xor XOR2 (N1266, N1261, N1057);
buf BUF1 (N1267, N1256);
nor NOR4 (N1268, N1267, N1266, N1061, N1246);
not NOT1 (N1269, N140);
buf BUF1 (N1270, N1255);
nor NOR2 (N1271, N1270, N1094);
nor NOR3 (N1272, N1226, N887, N570);
buf BUF1 (N1273, N1272);
or OR2 (N1274, N1258, N544);
and AND3 (N1275, N1274, N1254, N7);
nand NAND4 (N1276, N1273, N192, N537, N1066);
and AND4 (N1277, N1251, N888, N820, N29);
buf BUF1 (N1278, N1276);
xor XOR2 (N1279, N1265, N1162);
not NOT1 (N1280, N1264);
or OR2 (N1281, N1252, N347);
not NOT1 (N1282, N1243);
nor NOR4 (N1283, N1278, N476, N1057, N402);
not NOT1 (N1284, N1281);
and AND2 (N1285, N1277, N1024);
nand NAND3 (N1286, N1285, N407, N322);
and AND4 (N1287, N1271, N606, N8, N771);
xor XOR2 (N1288, N1284, N1236);
nor NOR4 (N1289, N1286, N859, N682, N1105);
or OR4 (N1290, N1288, N57, N1167, N1185);
and AND2 (N1291, N1289, N838);
xor XOR2 (N1292, N1280, N918);
nand NAND3 (N1293, N1291, N358, N237);
xor XOR2 (N1294, N1290, N25);
nor NOR2 (N1295, N1287, N853);
or OR4 (N1296, N1279, N519, N1152, N537);
or OR4 (N1297, N1294, N861, N1240, N22);
xor XOR2 (N1298, N1295, N1009);
or OR3 (N1299, N1282, N693, N648);
not NOT1 (N1300, N1268);
nor NOR3 (N1301, N1300, N31, N892);
buf BUF1 (N1302, N1293);
nor NOR3 (N1303, N1298, N1128, N41);
and AND2 (N1304, N1299, N1194);
nand NAND2 (N1305, N1304, N824);
and AND3 (N1306, N1283, N1168, N1204);
and AND3 (N1307, N1303, N1298, N110);
not NOT1 (N1308, N1296);
not NOT1 (N1309, N1292);
or OR4 (N1310, N1307, N444, N467, N439);
xor XOR2 (N1311, N1302, N1170);
or OR2 (N1312, N1275, N401);
or OR3 (N1313, N1310, N607, N266);
or OR4 (N1314, N1309, N1235, N630, N391);
buf BUF1 (N1315, N1305);
nor NOR4 (N1316, N1301, N908, N137, N23);
or OR2 (N1317, N1316, N347);
nor NOR2 (N1318, N1314, N252);
or OR2 (N1319, N1318, N663);
buf BUF1 (N1320, N1297);
or OR4 (N1321, N1313, N650, N1282, N527);
buf BUF1 (N1322, N1319);
and AND3 (N1323, N1320, N473, N406);
buf BUF1 (N1324, N1317);
and AND2 (N1325, N1306, N129);
and AND2 (N1326, N1323, N728);
nor NOR2 (N1327, N1324, N1260);
not NOT1 (N1328, N1315);
buf BUF1 (N1329, N1312);
xor XOR2 (N1330, N1311, N551);
or OR4 (N1331, N1328, N950, N686, N757);
nand NAND4 (N1332, N1325, N71, N683, N1251);
or OR3 (N1333, N1326, N701, N187);
xor XOR2 (N1334, N1269, N31);
or OR4 (N1335, N1322, N1245, N445, N404);
buf BUF1 (N1336, N1308);
nand NAND3 (N1337, N1334, N936, N466);
nand NAND3 (N1338, N1327, N649, N1232);
or OR2 (N1339, N1338, N208);
nand NAND2 (N1340, N1335, N1104);
nand NAND4 (N1341, N1330, N263, N303, N1327);
not NOT1 (N1342, N1329);
and AND4 (N1343, N1321, N10, N38, N218);
or OR2 (N1344, N1341, N468);
xor XOR2 (N1345, N1337, N1296);
and AND2 (N1346, N1339, N893);
and AND4 (N1347, N1336, N57, N105, N714);
not NOT1 (N1348, N1332);
buf BUF1 (N1349, N1343);
nor NOR3 (N1350, N1348, N41, N355);
and AND2 (N1351, N1331, N1321);
and AND3 (N1352, N1347, N1104, N314);
buf BUF1 (N1353, N1340);
not NOT1 (N1354, N1349);
buf BUF1 (N1355, N1346);
nor NOR4 (N1356, N1351, N1185, N377, N120);
nand NAND3 (N1357, N1353, N940, N200);
buf BUF1 (N1358, N1342);
buf BUF1 (N1359, N1333);
nor NOR3 (N1360, N1352, N267, N1212);
nand NAND3 (N1361, N1354, N1347, N44);
buf BUF1 (N1362, N1361);
or OR2 (N1363, N1357, N331);
or OR2 (N1364, N1345, N716);
buf BUF1 (N1365, N1350);
or OR4 (N1366, N1362, N655, N714, N527);
nand NAND4 (N1367, N1364, N465, N1232, N577);
nor NOR2 (N1368, N1366, N1344);
or OR4 (N1369, N1340, N1332, N63, N338);
nand NAND3 (N1370, N1365, N1175, N182);
or OR3 (N1371, N1359, N276, N1264);
and AND3 (N1372, N1370, N1252, N636);
nand NAND3 (N1373, N1358, N1334, N934);
buf BUF1 (N1374, N1356);
buf BUF1 (N1375, N1369);
not NOT1 (N1376, N1363);
not NOT1 (N1377, N1368);
nand NAND4 (N1378, N1372, N529, N1300, N940);
nand NAND4 (N1379, N1374, N179, N31, N1333);
buf BUF1 (N1380, N1367);
nand NAND2 (N1381, N1360, N333);
nand NAND2 (N1382, N1375, N1222);
not NOT1 (N1383, N1379);
nand NAND4 (N1384, N1381, N1201, N528, N176);
not NOT1 (N1385, N1380);
not NOT1 (N1386, N1376);
buf BUF1 (N1387, N1385);
nor NOR2 (N1388, N1382, N1360);
not NOT1 (N1389, N1378);
not NOT1 (N1390, N1373);
not NOT1 (N1391, N1389);
or OR3 (N1392, N1388, N45, N891);
or OR2 (N1393, N1386, N179);
nor NOR3 (N1394, N1392, N640, N330);
xor XOR2 (N1395, N1355, N1349);
and AND3 (N1396, N1391, N649, N883);
or OR3 (N1397, N1377, N51, N1324);
nand NAND3 (N1398, N1384, N1335, N755);
and AND3 (N1399, N1396, N430, N1398);
or OR3 (N1400, N277, N1297, N1268);
or OR4 (N1401, N1393, N247, N563, N547);
and AND3 (N1402, N1387, N676, N677);
buf BUF1 (N1403, N1397);
and AND4 (N1404, N1400, N930, N44, N838);
nand NAND3 (N1405, N1395, N145, N1204);
and AND4 (N1406, N1402, N79, N1042, N733);
nor NOR4 (N1407, N1406, N78, N1337, N385);
nor NOR4 (N1408, N1390, N215, N1348, N1379);
buf BUF1 (N1409, N1405);
not NOT1 (N1410, N1408);
or OR3 (N1411, N1403, N132, N659);
nor NOR3 (N1412, N1410, N903, N1409);
nand NAND4 (N1413, N516, N983, N229, N67);
not NOT1 (N1414, N1401);
and AND2 (N1415, N1394, N1155);
or OR2 (N1416, N1412, N407);
nor NOR3 (N1417, N1411, N1327, N226);
or OR4 (N1418, N1404, N179, N92, N631);
not NOT1 (N1419, N1416);
and AND4 (N1420, N1417, N307, N426, N1368);
not NOT1 (N1421, N1371);
nor NOR2 (N1422, N1383, N152);
xor XOR2 (N1423, N1421, N1106);
xor XOR2 (N1424, N1423, N204);
xor XOR2 (N1425, N1407, N161);
xor XOR2 (N1426, N1422, N1315);
or OR3 (N1427, N1415, N287, N303);
buf BUF1 (N1428, N1419);
or OR3 (N1429, N1399, N37, N905);
xor XOR2 (N1430, N1428, N529);
nand NAND3 (N1431, N1425, N598, N915);
and AND3 (N1432, N1426, N1351, N865);
nand NAND2 (N1433, N1431, N459);
not NOT1 (N1434, N1418);
or OR2 (N1435, N1413, N846);
not NOT1 (N1436, N1420);
buf BUF1 (N1437, N1429);
nor NOR2 (N1438, N1434, N304);
buf BUF1 (N1439, N1424);
or OR2 (N1440, N1438, N931);
not NOT1 (N1441, N1439);
nor NOR4 (N1442, N1440, N1248, N254, N58);
and AND2 (N1443, N1432, N663);
nor NOR4 (N1444, N1414, N345, N721, N672);
buf BUF1 (N1445, N1444);
and AND2 (N1446, N1435, N1279);
nor NOR4 (N1447, N1433, N968, N1387, N372);
xor XOR2 (N1448, N1447, N95);
nand NAND2 (N1449, N1448, N1039);
and AND2 (N1450, N1449, N143);
nand NAND3 (N1451, N1445, N195, N807);
or OR3 (N1452, N1442, N1446, N276);
nor NOR2 (N1453, N43, N561);
nand NAND3 (N1454, N1443, N532, N1245);
xor XOR2 (N1455, N1453, N599);
xor XOR2 (N1456, N1450, N459);
or OR4 (N1457, N1436, N482, N613, N316);
and AND3 (N1458, N1427, N1033, N386);
xor XOR2 (N1459, N1441, N1399);
not NOT1 (N1460, N1430);
not NOT1 (N1461, N1437);
nor NOR2 (N1462, N1451, N517);
not NOT1 (N1463, N1459);
not NOT1 (N1464, N1455);
xor XOR2 (N1465, N1460, N777);
buf BUF1 (N1466, N1461);
not NOT1 (N1467, N1466);
nand NAND4 (N1468, N1458, N1160, N162, N1321);
not NOT1 (N1469, N1462);
buf BUF1 (N1470, N1469);
nand NAND2 (N1471, N1463, N1222);
xor XOR2 (N1472, N1454, N339);
nor NOR3 (N1473, N1464, N1266, N175);
not NOT1 (N1474, N1472);
nand NAND2 (N1475, N1474, N784);
nor NOR2 (N1476, N1452, N137);
not NOT1 (N1477, N1465);
nand NAND4 (N1478, N1468, N3, N345, N518);
or OR2 (N1479, N1477, N448);
not NOT1 (N1480, N1467);
nand NAND4 (N1481, N1480, N1335, N441, N234);
and AND2 (N1482, N1481, N1365);
xor XOR2 (N1483, N1470, N1087);
and AND2 (N1484, N1478, N983);
not NOT1 (N1485, N1479);
buf BUF1 (N1486, N1475);
xor XOR2 (N1487, N1484, N184);
or OR2 (N1488, N1483, N264);
nor NOR3 (N1489, N1471, N91, N1311);
or OR2 (N1490, N1485, N216);
buf BUF1 (N1491, N1457);
nand NAND3 (N1492, N1489, N1271, N1264);
xor XOR2 (N1493, N1491, N274);
or OR4 (N1494, N1486, N32, N651, N683);
or OR3 (N1495, N1473, N952, N1067);
not NOT1 (N1496, N1482);
or OR2 (N1497, N1495, N371);
buf BUF1 (N1498, N1490);
xor XOR2 (N1499, N1456, N788);
nand NAND4 (N1500, N1488, N633, N867, N767);
nand NAND2 (N1501, N1492, N15);
buf BUF1 (N1502, N1494);
nand NAND2 (N1503, N1496, N592);
and AND3 (N1504, N1476, N585, N757);
and AND3 (N1505, N1487, N68, N73);
buf BUF1 (N1506, N1493);
not NOT1 (N1507, N1501);
xor XOR2 (N1508, N1503, N241);
xor XOR2 (N1509, N1507, N376);
not NOT1 (N1510, N1509);
not NOT1 (N1511, N1504);
buf BUF1 (N1512, N1497);
buf BUF1 (N1513, N1505);
or OR4 (N1514, N1506, N341, N817, N1223);
nand NAND4 (N1515, N1511, N506, N108, N1367);
nand NAND2 (N1516, N1513, N242);
nand NAND4 (N1517, N1512, N116, N692, N331);
xor XOR2 (N1518, N1499, N533);
nor NOR4 (N1519, N1515, N1061, N1473, N49);
buf BUF1 (N1520, N1516);
not NOT1 (N1521, N1518);
nor NOR3 (N1522, N1498, N929, N663);
nor NOR2 (N1523, N1522, N138);
nand NAND2 (N1524, N1508, N812);
nor NOR4 (N1525, N1524, N1336, N1193, N1518);
or OR4 (N1526, N1521, N839, N1114, N1523);
nand NAND3 (N1527, N482, N159, N960);
buf BUF1 (N1528, N1520);
xor XOR2 (N1529, N1514, N1137);
nor NOR2 (N1530, N1510, N391);
nor NOR3 (N1531, N1529, N402, N1232);
not NOT1 (N1532, N1519);
nand NAND2 (N1533, N1500, N520);
nand NAND2 (N1534, N1517, N1249);
buf BUF1 (N1535, N1502);
or OR2 (N1536, N1526, N1202);
nor NOR2 (N1537, N1531, N470);
buf BUF1 (N1538, N1532);
or OR3 (N1539, N1530, N39, N1133);
xor XOR2 (N1540, N1527, N969);
or OR3 (N1541, N1538, N560, N1338);
not NOT1 (N1542, N1525);
nand NAND4 (N1543, N1542, N1025, N863, N961);
buf BUF1 (N1544, N1533);
or OR2 (N1545, N1536, N1377);
not NOT1 (N1546, N1543);
xor XOR2 (N1547, N1541, N1313);
not NOT1 (N1548, N1545);
nand NAND3 (N1549, N1546, N636, N979);
and AND2 (N1550, N1548, N121);
buf BUF1 (N1551, N1539);
not NOT1 (N1552, N1540);
buf BUF1 (N1553, N1552);
or OR2 (N1554, N1544, N300);
nand NAND2 (N1555, N1537, N721);
buf BUF1 (N1556, N1550);
xor XOR2 (N1557, N1547, N389);
not NOT1 (N1558, N1555);
or OR3 (N1559, N1528, N1020, N1518);
not NOT1 (N1560, N1556);
and AND4 (N1561, N1535, N1005, N387, N290);
or OR2 (N1562, N1553, N359);
nand NAND2 (N1563, N1554, N362);
buf BUF1 (N1564, N1557);
or OR2 (N1565, N1563, N1534);
nor NOR4 (N1566, N692, N90, N1307, N528);
nor NOR3 (N1567, N1558, N9, N1311);
not NOT1 (N1568, N1566);
xor XOR2 (N1569, N1562, N627);
and AND3 (N1570, N1559, N424, N1387);
nand NAND2 (N1571, N1549, N1217);
buf BUF1 (N1572, N1565);
or OR4 (N1573, N1569, N1165, N1006, N99);
xor XOR2 (N1574, N1572, N173);
buf BUF1 (N1575, N1573);
not NOT1 (N1576, N1575);
nor NOR2 (N1577, N1574, N1135);
nor NOR3 (N1578, N1571, N892, N310);
buf BUF1 (N1579, N1578);
nand NAND4 (N1580, N1564, N1271, N829, N662);
or OR4 (N1581, N1568, N325, N428, N1242);
nor NOR3 (N1582, N1576, N1395, N1345);
nor NOR4 (N1583, N1577, N727, N1242, N1392);
xor XOR2 (N1584, N1583, N890);
nor NOR2 (N1585, N1561, N88);
xor XOR2 (N1586, N1585, N1009);
and AND2 (N1587, N1580, N1307);
buf BUF1 (N1588, N1567);
nand NAND2 (N1589, N1570, N418);
nand NAND2 (N1590, N1560, N1410);
and AND3 (N1591, N1587, N110, N352);
xor XOR2 (N1592, N1589, N598);
and AND3 (N1593, N1551, N1193, N176);
or OR3 (N1594, N1582, N198, N675);
or OR4 (N1595, N1584, N121, N1156, N669);
or OR4 (N1596, N1593, N1116, N628, N1264);
nand NAND3 (N1597, N1588, N839, N313);
xor XOR2 (N1598, N1594, N1474);
not NOT1 (N1599, N1595);
nor NOR3 (N1600, N1586, N1107, N305);
buf BUF1 (N1601, N1581);
and AND3 (N1602, N1579, N1393, N1356);
or OR3 (N1603, N1601, N228, N74);
nand NAND2 (N1604, N1596, N890);
buf BUF1 (N1605, N1602);
buf BUF1 (N1606, N1590);
buf BUF1 (N1607, N1592);
buf BUF1 (N1608, N1600);
and AND3 (N1609, N1603, N1339, N691);
buf BUF1 (N1610, N1597);
nor NOR2 (N1611, N1591, N825);
nand NAND2 (N1612, N1599, N939);
xor XOR2 (N1613, N1605, N1352);
buf BUF1 (N1614, N1609);
nand NAND2 (N1615, N1612, N410);
buf BUF1 (N1616, N1606);
xor XOR2 (N1617, N1616, N974);
nand NAND2 (N1618, N1614, N1331);
buf BUF1 (N1619, N1618);
nand NAND2 (N1620, N1611, N556);
and AND4 (N1621, N1604, N21, N493, N303);
and AND4 (N1622, N1621, N1084, N1272, N1113);
and AND3 (N1623, N1607, N1012, N1564);
xor XOR2 (N1624, N1598, N332);
nand NAND2 (N1625, N1622, N545);
or OR4 (N1626, N1625, N1408, N979, N85);
or OR4 (N1627, N1610, N314, N1257, N1388);
nand NAND2 (N1628, N1613, N310);
or OR3 (N1629, N1620, N129, N817);
or OR4 (N1630, N1617, N163, N890, N645);
buf BUF1 (N1631, N1626);
or OR2 (N1632, N1631, N242);
not NOT1 (N1633, N1608);
or OR2 (N1634, N1619, N502);
not NOT1 (N1635, N1623);
and AND3 (N1636, N1633, N417, N5);
nand NAND3 (N1637, N1634, N1265, N809);
or OR4 (N1638, N1627, N1578, N671, N636);
nor NOR4 (N1639, N1637, N595, N1508, N474);
not NOT1 (N1640, N1624);
and AND4 (N1641, N1638, N461, N377, N720);
nand NAND4 (N1642, N1640, N1552, N798, N967);
or OR4 (N1643, N1628, N1099, N123, N65);
xor XOR2 (N1644, N1641, N77);
buf BUF1 (N1645, N1632);
buf BUF1 (N1646, N1635);
or OR2 (N1647, N1645, N699);
or OR2 (N1648, N1643, N1380);
or OR3 (N1649, N1648, N1364, N735);
nand NAND3 (N1650, N1644, N626, N931);
not NOT1 (N1651, N1646);
nand NAND2 (N1652, N1630, N241);
or OR4 (N1653, N1636, N1198, N114, N95);
xor XOR2 (N1654, N1642, N827);
buf BUF1 (N1655, N1650);
or OR3 (N1656, N1655, N1047, N1139);
buf BUF1 (N1657, N1656);
and AND2 (N1658, N1629, N1531);
xor XOR2 (N1659, N1647, N573);
not NOT1 (N1660, N1654);
nand NAND2 (N1661, N1659, N80);
buf BUF1 (N1662, N1653);
xor XOR2 (N1663, N1661, N482);
nor NOR2 (N1664, N1652, N1435);
nor NOR2 (N1665, N1658, N163);
or OR2 (N1666, N1662, N286);
and AND2 (N1667, N1657, N620);
nor NOR4 (N1668, N1660, N1214, N751, N500);
not NOT1 (N1669, N1615);
not NOT1 (N1670, N1649);
not NOT1 (N1671, N1663);
nand NAND2 (N1672, N1668, N171);
xor XOR2 (N1673, N1667, N224);
or OR3 (N1674, N1672, N1447, N283);
buf BUF1 (N1675, N1666);
and AND3 (N1676, N1674, N13, N1015);
nand NAND2 (N1677, N1651, N908);
nand NAND3 (N1678, N1673, N1295, N612);
nor NOR3 (N1679, N1677, N508, N1031);
not NOT1 (N1680, N1665);
not NOT1 (N1681, N1676);
buf BUF1 (N1682, N1681);
nand NAND2 (N1683, N1670, N552);
buf BUF1 (N1684, N1664);
and AND3 (N1685, N1675, N113, N1394);
not NOT1 (N1686, N1679);
not NOT1 (N1687, N1639);
and AND4 (N1688, N1680, N1112, N279, N673);
or OR3 (N1689, N1688, N887, N678);
not NOT1 (N1690, N1683);
nand NAND3 (N1691, N1678, N1515, N601);
nor NOR4 (N1692, N1685, N1596, N1367, N145);
not NOT1 (N1693, N1671);
xor XOR2 (N1694, N1690, N463);
nor NOR3 (N1695, N1689, N933, N864);
xor XOR2 (N1696, N1682, N1542);
and AND2 (N1697, N1686, N407);
buf BUF1 (N1698, N1691);
or OR2 (N1699, N1694, N471);
or OR2 (N1700, N1687, N543);
nor NOR3 (N1701, N1695, N614, N536);
xor XOR2 (N1702, N1693, N1072);
nor NOR2 (N1703, N1701, N791);
xor XOR2 (N1704, N1669, N1604);
not NOT1 (N1705, N1697);
not NOT1 (N1706, N1692);
xor XOR2 (N1707, N1699, N22);
and AND3 (N1708, N1696, N1189, N484);
xor XOR2 (N1709, N1706, N1508);
and AND3 (N1710, N1704, N192, N27);
not NOT1 (N1711, N1710);
buf BUF1 (N1712, N1711);
nor NOR3 (N1713, N1698, N836, N1611);
and AND3 (N1714, N1702, N611, N1567);
and AND2 (N1715, N1707, N228);
buf BUF1 (N1716, N1700);
not NOT1 (N1717, N1708);
not NOT1 (N1718, N1703);
or OR3 (N1719, N1713, N746, N1230);
not NOT1 (N1720, N1712);
buf BUF1 (N1721, N1718);
or OR3 (N1722, N1714, N941, N676);
xor XOR2 (N1723, N1717, N396);
or OR3 (N1724, N1716, N209, N1456);
buf BUF1 (N1725, N1705);
not NOT1 (N1726, N1725);
nand NAND3 (N1727, N1723, N1188, N1581);
not NOT1 (N1728, N1722);
and AND2 (N1729, N1724, N407);
nand NAND2 (N1730, N1728, N919);
xor XOR2 (N1731, N1720, N440);
or OR2 (N1732, N1709, N270);
xor XOR2 (N1733, N1684, N869);
buf BUF1 (N1734, N1715);
nand NAND2 (N1735, N1721, N176);
and AND3 (N1736, N1733, N663, N1222);
nor NOR2 (N1737, N1731, N180);
nand NAND3 (N1738, N1730, N192, N1704);
nor NOR2 (N1739, N1737, N159);
nor NOR2 (N1740, N1736, N107);
or OR3 (N1741, N1729, N781, N1727);
not NOT1 (N1742, N134);
buf BUF1 (N1743, N1719);
xor XOR2 (N1744, N1734, N1115);
buf BUF1 (N1745, N1740);
not NOT1 (N1746, N1739);
buf BUF1 (N1747, N1732);
xor XOR2 (N1748, N1726, N197);
not NOT1 (N1749, N1735);
nand NAND3 (N1750, N1745, N1233, N1105);
or OR3 (N1751, N1748, N1382, N1255);
nand NAND4 (N1752, N1742, N483, N831, N1680);
nand NAND2 (N1753, N1751, N224);
and AND2 (N1754, N1738, N39);
not NOT1 (N1755, N1752);
xor XOR2 (N1756, N1750, N364);
buf BUF1 (N1757, N1749);
and AND3 (N1758, N1757, N1554, N117);
not NOT1 (N1759, N1754);
nand NAND4 (N1760, N1741, N1275, N1579, N553);
and AND4 (N1761, N1760, N614, N1568, N106);
nand NAND3 (N1762, N1758, N1157, N127);
xor XOR2 (N1763, N1759, N851);
xor XOR2 (N1764, N1763, N448);
nor NOR2 (N1765, N1743, N1702);
nand NAND3 (N1766, N1761, N936, N549);
or OR3 (N1767, N1764, N1217, N79);
buf BUF1 (N1768, N1747);
not NOT1 (N1769, N1766);
or OR4 (N1770, N1746, N1751, N1528, N65);
buf BUF1 (N1771, N1769);
and AND2 (N1772, N1753, N820);
or OR3 (N1773, N1767, N221, N1468);
xor XOR2 (N1774, N1771, N564);
or OR2 (N1775, N1765, N678);
xor XOR2 (N1776, N1773, N1245);
buf BUF1 (N1777, N1776);
and AND3 (N1778, N1744, N76, N1669);
or OR3 (N1779, N1770, N1437, N1215);
not NOT1 (N1780, N1778);
nand NAND3 (N1781, N1774, N780, N700);
nor NOR2 (N1782, N1781, N258);
and AND3 (N1783, N1782, N1305, N581);
buf BUF1 (N1784, N1772);
not NOT1 (N1785, N1783);
nand NAND2 (N1786, N1755, N682);
nand NAND4 (N1787, N1786, N518, N279, N226);
buf BUF1 (N1788, N1768);
not NOT1 (N1789, N1787);
and AND4 (N1790, N1775, N1218, N762, N911);
and AND3 (N1791, N1789, N748, N1602);
xor XOR2 (N1792, N1779, N627);
and AND2 (N1793, N1792, N478);
or OR4 (N1794, N1790, N1502, N1426, N1490);
xor XOR2 (N1795, N1780, N1343);
nand NAND4 (N1796, N1784, N174, N920, N105);
nand NAND2 (N1797, N1756, N132);
nor NOR2 (N1798, N1788, N623);
nor NOR3 (N1799, N1785, N1583, N966);
buf BUF1 (N1800, N1777);
or OR2 (N1801, N1795, N1167);
or OR4 (N1802, N1793, N1534, N261, N742);
xor XOR2 (N1803, N1800, N1431);
xor XOR2 (N1804, N1802, N1103);
nand NAND4 (N1805, N1798, N405, N1618, N374);
and AND2 (N1806, N1799, N1666);
nand NAND2 (N1807, N1762, N1767);
buf BUF1 (N1808, N1796);
and AND4 (N1809, N1806, N635, N840, N794);
nor NOR2 (N1810, N1809, N942);
not NOT1 (N1811, N1810);
nor NOR3 (N1812, N1791, N404, N884);
or OR2 (N1813, N1812, N306);
or OR2 (N1814, N1804, N998);
nand NAND4 (N1815, N1807, N1288, N562, N770);
nand NAND4 (N1816, N1803, N356, N745, N1525);
xor XOR2 (N1817, N1814, N266);
nand NAND2 (N1818, N1811, N1771);
or OR4 (N1819, N1815, N1063, N979, N769);
and AND4 (N1820, N1818, N989, N720, N63);
xor XOR2 (N1821, N1797, N581);
nand NAND4 (N1822, N1816, N1657, N1473, N611);
xor XOR2 (N1823, N1817, N1159);
xor XOR2 (N1824, N1823, N1674);
not NOT1 (N1825, N1821);
nand NAND3 (N1826, N1801, N1522, N1726);
not NOT1 (N1827, N1805);
nor NOR4 (N1828, N1808, N98, N1095, N326);
nor NOR2 (N1829, N1827, N538);
nor NOR3 (N1830, N1813, N466, N643);
and AND2 (N1831, N1830, N831);
not NOT1 (N1832, N1819);
xor XOR2 (N1833, N1825, N1635);
and AND4 (N1834, N1826, N224, N1430, N1055);
buf BUF1 (N1835, N1820);
buf BUF1 (N1836, N1832);
nor NOR3 (N1837, N1831, N549, N430);
nor NOR3 (N1838, N1836, N236, N433);
nor NOR2 (N1839, N1794, N1480);
not NOT1 (N1840, N1829);
nand NAND4 (N1841, N1840, N1207, N1316, N1650);
and AND3 (N1842, N1822, N442, N1387);
buf BUF1 (N1843, N1828);
xor XOR2 (N1844, N1824, N1026);
nor NOR2 (N1845, N1838, N66);
not NOT1 (N1846, N1841);
or OR2 (N1847, N1845, N260);
and AND2 (N1848, N1839, N584);
nand NAND3 (N1849, N1848, N1031, N384);
nand NAND3 (N1850, N1849, N562, N1144);
nand NAND3 (N1851, N1842, N766, N90);
xor XOR2 (N1852, N1846, N890);
xor XOR2 (N1853, N1844, N137);
or OR4 (N1854, N1837, N527, N977, N1785);
and AND3 (N1855, N1833, N289, N1758);
nor NOR4 (N1856, N1855, N300, N907, N1080);
and AND3 (N1857, N1854, N1697, N762);
nor NOR2 (N1858, N1835, N1476);
xor XOR2 (N1859, N1853, N498);
nor NOR2 (N1860, N1852, N1270);
nand NAND4 (N1861, N1850, N986, N383, N195);
not NOT1 (N1862, N1860);
xor XOR2 (N1863, N1851, N1528);
buf BUF1 (N1864, N1859);
nand NAND3 (N1865, N1863, N1177, N565);
nand NAND4 (N1866, N1847, N1122, N1219, N711);
xor XOR2 (N1867, N1858, N768);
not NOT1 (N1868, N1862);
and AND4 (N1869, N1866, N286, N1859, N520);
nor NOR2 (N1870, N1857, N573);
buf BUF1 (N1871, N1861);
nor NOR2 (N1872, N1868, N793);
not NOT1 (N1873, N1870);
nor NOR4 (N1874, N1856, N536, N160, N1612);
nand NAND3 (N1875, N1843, N745, N297);
and AND3 (N1876, N1871, N1421, N1005);
and AND2 (N1877, N1876, N389);
or OR2 (N1878, N1877, N1337);
buf BUF1 (N1879, N1873);
not NOT1 (N1880, N1864);
not NOT1 (N1881, N1875);
or OR3 (N1882, N1880, N395, N1104);
or OR2 (N1883, N1867, N710);
or OR3 (N1884, N1869, N1437, N1465);
xor XOR2 (N1885, N1865, N815);
nand NAND2 (N1886, N1884, N1168);
not NOT1 (N1887, N1879);
not NOT1 (N1888, N1872);
not NOT1 (N1889, N1887);
buf BUF1 (N1890, N1882);
nor NOR3 (N1891, N1888, N945, N1611);
buf BUF1 (N1892, N1883);
buf BUF1 (N1893, N1886);
nand NAND3 (N1894, N1881, N98, N1031);
and AND2 (N1895, N1892, N50);
not NOT1 (N1896, N1874);
nor NOR4 (N1897, N1885, N1718, N1424, N1125);
or OR4 (N1898, N1834, N1766, N1490, N103);
and AND3 (N1899, N1897, N1615, N1808);
xor XOR2 (N1900, N1893, N1276);
or OR2 (N1901, N1890, N743);
and AND3 (N1902, N1896, N952, N1594);
and AND4 (N1903, N1895, N521, N901, N853);
xor XOR2 (N1904, N1891, N668);
or OR2 (N1905, N1898, N1521);
buf BUF1 (N1906, N1903);
buf BUF1 (N1907, N1889);
not NOT1 (N1908, N1894);
buf BUF1 (N1909, N1905);
not NOT1 (N1910, N1909);
nand NAND3 (N1911, N1900, N1884, N1644);
not NOT1 (N1912, N1907);
nand NAND2 (N1913, N1904, N1544);
nor NOR2 (N1914, N1910, N1293);
or OR2 (N1915, N1901, N443);
buf BUF1 (N1916, N1911);
nand NAND3 (N1917, N1916, N1512, N362);
and AND4 (N1918, N1899, N1819, N1764, N161);
nand NAND2 (N1919, N1878, N646);
or OR2 (N1920, N1918, N1449);
buf BUF1 (N1921, N1906);
xor XOR2 (N1922, N1921, N34);
and AND3 (N1923, N1908, N531, N1909);
and AND2 (N1924, N1917, N1776);
not NOT1 (N1925, N1913);
not NOT1 (N1926, N1915);
and AND2 (N1927, N1902, N922);
nand NAND3 (N1928, N1926, N294, N747);
and AND2 (N1929, N1928, N1300);
and AND3 (N1930, N1924, N1352, N995);
buf BUF1 (N1931, N1919);
and AND3 (N1932, N1920, N1064, N529);
or OR2 (N1933, N1925, N1335);
and AND3 (N1934, N1912, N1478, N1323);
nor NOR4 (N1935, N1922, N1500, N35, N329);
and AND4 (N1936, N1933, N391, N1791, N763);
nand NAND2 (N1937, N1935, N1005);
xor XOR2 (N1938, N1931, N52);
xor XOR2 (N1939, N1932, N334);
and AND3 (N1940, N1929, N27, N913);
nor NOR2 (N1941, N1930, N1175);
nor NOR2 (N1942, N1936, N1416);
or OR3 (N1943, N1934, N327, N1038);
xor XOR2 (N1944, N1943, N1162);
buf BUF1 (N1945, N1941);
not NOT1 (N1946, N1944);
nor NOR3 (N1947, N1938, N475, N1110);
xor XOR2 (N1948, N1939, N244);
and AND2 (N1949, N1948, N373);
not NOT1 (N1950, N1949);
nand NAND4 (N1951, N1914, N89, N578, N1808);
xor XOR2 (N1952, N1937, N208);
and AND3 (N1953, N1951, N1475, N1091);
nor NOR2 (N1954, N1947, N766);
and AND2 (N1955, N1950, N849);
xor XOR2 (N1956, N1952, N1392);
and AND4 (N1957, N1953, N362, N1196, N1822);
and AND3 (N1958, N1955, N1048, N825);
not NOT1 (N1959, N1957);
not NOT1 (N1960, N1942);
nand NAND3 (N1961, N1960, N102, N1696);
or OR3 (N1962, N1954, N687, N97);
xor XOR2 (N1963, N1958, N1440);
not NOT1 (N1964, N1940);
nand NAND3 (N1965, N1956, N181, N925);
nand NAND3 (N1966, N1923, N125, N284);
or OR2 (N1967, N1959, N277);
nor NOR2 (N1968, N1961, N503);
xor XOR2 (N1969, N1945, N1198);
not NOT1 (N1970, N1927);
and AND4 (N1971, N1966, N363, N1876, N685);
nand NAND3 (N1972, N1971, N1545, N987);
xor XOR2 (N1973, N1972, N721);
nor NOR3 (N1974, N1970, N1586, N1754);
nor NOR3 (N1975, N1968, N1541, N1973);
nor NOR3 (N1976, N61, N571, N1491);
and AND2 (N1977, N1967, N149);
not NOT1 (N1978, N1976);
not NOT1 (N1979, N1974);
not NOT1 (N1980, N1975);
xor XOR2 (N1981, N1964, N264);
nand NAND2 (N1982, N1963, N1162);
not NOT1 (N1983, N1977);
not NOT1 (N1984, N1982);
nand NAND4 (N1985, N1978, N483, N871, N1103);
buf BUF1 (N1986, N1981);
nor NOR3 (N1987, N1969, N330, N508);
and AND3 (N1988, N1984, N1014, N775);
xor XOR2 (N1989, N1979, N1935);
nor NOR2 (N1990, N1946, N1546);
and AND4 (N1991, N1986, N681, N57, N975);
or OR4 (N1992, N1990, N1959, N1971, N1497);
not NOT1 (N1993, N1989);
nand NAND3 (N1994, N1965, N487, N586);
nor NOR4 (N1995, N1987, N44, N1495, N300);
and AND4 (N1996, N1980, N1854, N1238, N1869);
nand NAND3 (N1997, N1996, N594, N960);
nand NAND3 (N1998, N1995, N875, N916);
buf BUF1 (N1999, N1997);
nand NAND2 (N2000, N1993, N1197);
not NOT1 (N2001, N1994);
nor NOR2 (N2002, N1991, N528);
and AND2 (N2003, N1985, N78);
nand NAND3 (N2004, N1988, N690, N515);
or OR3 (N2005, N1992, N485, N1334);
buf BUF1 (N2006, N1962);
buf BUF1 (N2007, N2006);
nand NAND3 (N2008, N2007, N17, N1204);
nor NOR2 (N2009, N2002, N777);
or OR2 (N2010, N2000, N868);
and AND2 (N2011, N2004, N1035);
xor XOR2 (N2012, N2001, N802);
nand NAND2 (N2013, N1999, N1090);
or OR4 (N2014, N2003, N1927, N1884, N1384);
not NOT1 (N2015, N1983);
or OR2 (N2016, N2013, N1681);
buf BUF1 (N2017, N2012);
nor NOR3 (N2018, N2005, N251, N857);
nand NAND2 (N2019, N2014, N1079);
buf BUF1 (N2020, N2009);
or OR4 (N2021, N2019, N933, N812, N61);
nor NOR4 (N2022, N1998, N1125, N585, N912);
and AND3 (N2023, N2010, N1075, N989);
or OR4 (N2024, N2008, N181, N1789, N37);
nand NAND2 (N2025, N2023, N1041);
not NOT1 (N2026, N2016);
nor NOR2 (N2027, N2026, N1929);
or OR3 (N2028, N2018, N5, N1410);
nor NOR2 (N2029, N2028, N364);
nand NAND3 (N2030, N2020, N1359, N1926);
nand NAND2 (N2031, N2022, N1889);
not NOT1 (N2032, N2031);
buf BUF1 (N2033, N2015);
xor XOR2 (N2034, N2024, N234);
nand NAND2 (N2035, N2033, N157);
xor XOR2 (N2036, N2034, N875);
and AND3 (N2037, N2011, N1233, N411);
not NOT1 (N2038, N2030);
nor NOR4 (N2039, N2027, N1960, N779, N583);
and AND2 (N2040, N2035, N623);
nor NOR3 (N2041, N2040, N1965, N595);
or OR2 (N2042, N2017, N507);
xor XOR2 (N2043, N2021, N1429);
not NOT1 (N2044, N2029);
nor NOR4 (N2045, N2042, N691, N1599, N1702);
buf BUF1 (N2046, N2025);
nor NOR2 (N2047, N2037, N857);
and AND2 (N2048, N2045, N1121);
nor NOR4 (N2049, N2046, N933, N1351, N443);
nor NOR4 (N2050, N2049, N1697, N712, N1113);
and AND3 (N2051, N2048, N472, N1066);
buf BUF1 (N2052, N2038);
and AND2 (N2053, N2032, N562);
buf BUF1 (N2054, N2044);
not NOT1 (N2055, N2050);
or OR3 (N2056, N2036, N592, N244);
buf BUF1 (N2057, N2039);
nor NOR4 (N2058, N2056, N1855, N1425, N1489);
not NOT1 (N2059, N2058);
and AND4 (N2060, N2057, N908, N1982, N1882);
and AND3 (N2061, N2053, N2051, N666);
or OR4 (N2062, N1059, N808, N285, N38);
xor XOR2 (N2063, N2052, N1624);
or OR3 (N2064, N2063, N1971, N913);
not NOT1 (N2065, N2054);
xor XOR2 (N2066, N2047, N406);
nor NOR2 (N2067, N2062, N1178);
nor NOR3 (N2068, N2064, N863, N1584);
not NOT1 (N2069, N2041);
not NOT1 (N2070, N2069);
xor XOR2 (N2071, N2061, N883);
and AND4 (N2072, N2043, N512, N1621, N1166);
buf BUF1 (N2073, N2072);
not NOT1 (N2074, N2071);
nand NAND2 (N2075, N2067, N1390);
and AND3 (N2076, N2074, N1705, N37);
nor NOR2 (N2077, N2070, N1481);
and AND2 (N2078, N2066, N815);
buf BUF1 (N2079, N2068);
nor NOR4 (N2080, N2059, N654, N1958, N314);
and AND3 (N2081, N2077, N543, N802);
and AND4 (N2082, N2073, N1199, N995, N205);
nand NAND2 (N2083, N2055, N1692);
not NOT1 (N2084, N2076);
or OR3 (N2085, N2082, N905, N68);
nand NAND3 (N2086, N2075, N601, N649);
xor XOR2 (N2087, N2083, N1034);
buf BUF1 (N2088, N2078);
nand NAND2 (N2089, N2079, N363);
nor NOR3 (N2090, N2087, N227, N964);
and AND3 (N2091, N2086, N1642, N534);
or OR3 (N2092, N2060, N1935, N1033);
nor NOR3 (N2093, N2091, N1944, N1801);
and AND3 (N2094, N2092, N1307, N1673);
and AND2 (N2095, N2088, N1050);
or OR3 (N2096, N2094, N1964, N1435);
and AND3 (N2097, N2090, N452, N952);
nand NAND2 (N2098, N2096, N1639);
or OR3 (N2099, N2065, N1857, N670);
buf BUF1 (N2100, N2080);
or OR3 (N2101, N2097, N2011, N323);
buf BUF1 (N2102, N2101);
nand NAND4 (N2103, N2085, N280, N832, N2044);
and AND2 (N2104, N2099, N730);
not NOT1 (N2105, N2100);
or OR2 (N2106, N2089, N996);
not NOT1 (N2107, N2095);
nand NAND3 (N2108, N2081, N1833, N1668);
nand NAND2 (N2109, N2105, N41);
xor XOR2 (N2110, N2107, N1881);
nand NAND3 (N2111, N2108, N471, N979);
buf BUF1 (N2112, N2098);
and AND4 (N2113, N2104, N1664, N1535, N130);
nand NAND4 (N2114, N2093, N1729, N994, N1352);
not NOT1 (N2115, N2102);
nor NOR2 (N2116, N2114, N1835);
nand NAND3 (N2117, N2113, N993, N925);
nor NOR3 (N2118, N2084, N851, N1993);
buf BUF1 (N2119, N2111);
nor NOR4 (N2120, N2116, N1381, N645, N1186);
nor NOR2 (N2121, N2112, N576);
buf BUF1 (N2122, N2117);
xor XOR2 (N2123, N2109, N1097);
not NOT1 (N2124, N2103);
and AND2 (N2125, N2120, N2013);
xor XOR2 (N2126, N2115, N827);
or OR2 (N2127, N2125, N737);
xor XOR2 (N2128, N2123, N1479);
nand NAND3 (N2129, N2124, N806, N1560);
and AND3 (N2130, N2119, N314, N221);
xor XOR2 (N2131, N2122, N2020);
buf BUF1 (N2132, N2106);
nor NOR2 (N2133, N2118, N394);
xor XOR2 (N2134, N2132, N1888);
xor XOR2 (N2135, N2129, N1301);
and AND2 (N2136, N2135, N1867);
nand NAND2 (N2137, N2121, N1586);
xor XOR2 (N2138, N2128, N352);
nor NOR3 (N2139, N2133, N1785, N2054);
nor NOR3 (N2140, N2130, N2133, N1939);
nand NAND2 (N2141, N2127, N263);
xor XOR2 (N2142, N2137, N2082);
not NOT1 (N2143, N2140);
not NOT1 (N2144, N2141);
buf BUF1 (N2145, N2126);
buf BUF1 (N2146, N2142);
or OR3 (N2147, N2110, N2032, N1995);
not NOT1 (N2148, N2134);
xor XOR2 (N2149, N2148, N119);
nand NAND4 (N2150, N2145, N1932, N7, N1380);
and AND3 (N2151, N2150, N233, N419);
buf BUF1 (N2152, N2147);
not NOT1 (N2153, N2149);
or OR4 (N2154, N2143, N729, N1035, N1912);
nor NOR4 (N2155, N2136, N199, N657, N264);
or OR4 (N2156, N2131, N1514, N744, N741);
nand NAND2 (N2157, N2138, N498);
and AND2 (N2158, N2144, N192);
buf BUF1 (N2159, N2154);
or OR2 (N2160, N2139, N1522);
and AND2 (N2161, N2152, N1186);
and AND2 (N2162, N2156, N433);
and AND4 (N2163, N2151, N1215, N1213, N493);
buf BUF1 (N2164, N2163);
or OR3 (N2165, N2158, N114, N2153);
not NOT1 (N2166, N1520);
nand NAND2 (N2167, N2165, N995);
nand NAND2 (N2168, N2160, N1303);
nor NOR3 (N2169, N2159, N1812, N1924);
nor NOR3 (N2170, N2162, N442, N1420);
buf BUF1 (N2171, N2168);
buf BUF1 (N2172, N2164);
buf BUF1 (N2173, N2169);
or OR4 (N2174, N2155, N1979, N14, N396);
buf BUF1 (N2175, N2157);
nor NOR4 (N2176, N2174, N1957, N1525, N1004);
nand NAND2 (N2177, N2171, N971);
xor XOR2 (N2178, N2167, N1955);
not NOT1 (N2179, N2177);
nand NAND4 (N2180, N2172, N1461, N1099, N177);
xor XOR2 (N2181, N2178, N862);
or OR3 (N2182, N2180, N753, N1175);
nand NAND3 (N2183, N2181, N1448, N1509);
not NOT1 (N2184, N2182);
buf BUF1 (N2185, N2184);
or OR3 (N2186, N2176, N1199, N132);
buf BUF1 (N2187, N2170);
buf BUF1 (N2188, N2183);
and AND4 (N2189, N2179, N1204, N700, N1266);
or OR3 (N2190, N2146, N1001, N408);
not NOT1 (N2191, N2187);
not NOT1 (N2192, N2191);
buf BUF1 (N2193, N2161);
nand NAND3 (N2194, N2189, N1286, N1351);
or OR2 (N2195, N2185, N876);
buf BUF1 (N2196, N2173);
buf BUF1 (N2197, N2196);
nand NAND2 (N2198, N2190, N1780);
buf BUF1 (N2199, N2194);
not NOT1 (N2200, N2186);
not NOT1 (N2201, N2200);
nand NAND2 (N2202, N2201, N807);
buf BUF1 (N2203, N2166);
nor NOR3 (N2204, N2203, N1880, N2008);
nand NAND2 (N2205, N2195, N706);
or OR4 (N2206, N2192, N1463, N2035, N701);
not NOT1 (N2207, N2205);
xor XOR2 (N2208, N2193, N7);
xor XOR2 (N2209, N2207, N1214);
nor NOR4 (N2210, N2175, N601, N327, N1922);
or OR2 (N2211, N2209, N340);
buf BUF1 (N2212, N2198);
xor XOR2 (N2213, N2202, N1178);
nor NOR4 (N2214, N2204, N1916, N658, N2165);
or OR4 (N2215, N2199, N1700, N411, N2018);
buf BUF1 (N2216, N2206);
nor NOR4 (N2217, N2210, N1311, N1925, N1758);
and AND3 (N2218, N2215, N135, N449);
xor XOR2 (N2219, N2188, N1547);
and AND2 (N2220, N2216, N237);
nor NOR3 (N2221, N2197, N71, N665);
nand NAND2 (N2222, N2220, N162);
nor NOR4 (N2223, N2221, N530, N1199, N1995);
or OR2 (N2224, N2214, N1392);
buf BUF1 (N2225, N2212);
nand NAND2 (N2226, N2213, N2097);
buf BUF1 (N2227, N2218);
xor XOR2 (N2228, N2223, N261);
not NOT1 (N2229, N2224);
or OR3 (N2230, N2228, N1458, N384);
not NOT1 (N2231, N2211);
nand NAND3 (N2232, N2226, N712, N2174);
or OR3 (N2233, N2217, N1223, N1563);
or OR2 (N2234, N2222, N1234);
not NOT1 (N2235, N2230);
xor XOR2 (N2236, N2232, N1262);
nand NAND4 (N2237, N2233, N597, N531, N403);
buf BUF1 (N2238, N2225);
buf BUF1 (N2239, N2231);
nor NOR2 (N2240, N2234, N393);
and AND2 (N2241, N2227, N297);
nor NOR3 (N2242, N2241, N960, N760);
and AND3 (N2243, N2240, N1376, N715);
not NOT1 (N2244, N2235);
nand NAND3 (N2245, N2236, N155, N455);
nor NOR3 (N2246, N2238, N643, N639);
and AND4 (N2247, N2239, N1968, N250, N1307);
and AND4 (N2248, N2208, N1072, N2171, N254);
nand NAND2 (N2249, N2243, N1056);
nand NAND2 (N2250, N2249, N2159);
nor NOR2 (N2251, N2245, N505);
or OR2 (N2252, N2247, N703);
buf BUF1 (N2253, N2250);
xor XOR2 (N2254, N2248, N1981);
buf BUF1 (N2255, N2237);
nor NOR4 (N2256, N2252, N1493, N1579, N1076);
buf BUF1 (N2257, N2242);
nor NOR2 (N2258, N2251, N767);
and AND3 (N2259, N2256, N930, N685);
nor NOR3 (N2260, N2244, N826, N587);
buf BUF1 (N2261, N2219);
not NOT1 (N2262, N2261);
not NOT1 (N2263, N2255);
nor NOR3 (N2264, N2259, N317, N633);
xor XOR2 (N2265, N2253, N797);
xor XOR2 (N2266, N2229, N2018);
xor XOR2 (N2267, N2246, N518);
nor NOR2 (N2268, N2258, N1325);
not NOT1 (N2269, N2262);
nor NOR3 (N2270, N2268, N425, N532);
buf BUF1 (N2271, N2265);
nor NOR3 (N2272, N2270, N1431, N1415);
nand NAND3 (N2273, N2260, N1992, N1590);
buf BUF1 (N2274, N2267);
and AND4 (N2275, N2257, N88, N252, N1684);
and AND4 (N2276, N2272, N623, N1377, N1219);
and AND4 (N2277, N2264, N1228, N811, N2171);
and AND3 (N2278, N2269, N96, N1017);
not NOT1 (N2279, N2266);
nor NOR2 (N2280, N2275, N1949);
buf BUF1 (N2281, N2276);
not NOT1 (N2282, N2280);
nand NAND3 (N2283, N2281, N1408, N1083);
and AND2 (N2284, N2263, N188);
nand NAND3 (N2285, N2277, N1761, N1943);
nand NAND3 (N2286, N2282, N173, N1427);
nand NAND2 (N2287, N2283, N784);
or OR4 (N2288, N2254, N1803, N1958, N1505);
xor XOR2 (N2289, N2278, N1953);
nor NOR2 (N2290, N2279, N851);
nand NAND2 (N2291, N2287, N1225);
buf BUF1 (N2292, N2271);
buf BUF1 (N2293, N2289);
nor NOR3 (N2294, N2286, N1284, N1448);
xor XOR2 (N2295, N2285, N1840);
buf BUF1 (N2296, N2291);
nand NAND3 (N2297, N2284, N1653, N495);
and AND4 (N2298, N2295, N1672, N686, N2288);
or OR4 (N2299, N548, N460, N884, N237);
nand NAND2 (N2300, N2294, N1391);
or OR3 (N2301, N2273, N1562, N917);
buf BUF1 (N2302, N2300);
nand NAND4 (N2303, N2298, N465, N1418, N320);
not NOT1 (N2304, N2303);
not NOT1 (N2305, N2304);
and AND3 (N2306, N2296, N201, N106);
and AND3 (N2307, N2306, N1785, N1612);
and AND2 (N2308, N2301, N1835);
buf BUF1 (N2309, N2297);
not NOT1 (N2310, N2290);
and AND2 (N2311, N2307, N989);
xor XOR2 (N2312, N2309, N242);
not NOT1 (N2313, N2293);
xor XOR2 (N2314, N2312, N393);
or OR4 (N2315, N2274, N921, N2123, N1391);
nand NAND4 (N2316, N2308, N2297, N2299, N543);
not NOT1 (N2317, N56);
nand NAND2 (N2318, N2311, N258);
nor NOR2 (N2319, N2302, N412);
buf BUF1 (N2320, N2292);
nor NOR3 (N2321, N2305, N1711, N1552);
or OR2 (N2322, N2316, N1786);
nor NOR4 (N2323, N2314, N1781, N1280, N722);
not NOT1 (N2324, N2321);
not NOT1 (N2325, N2318);
nor NOR4 (N2326, N2315, N2092, N1943, N461);
nor NOR3 (N2327, N2322, N2131, N122);
buf BUF1 (N2328, N2327);
buf BUF1 (N2329, N2324);
buf BUF1 (N2330, N2328);
or OR3 (N2331, N2326, N482, N1189);
nand NAND3 (N2332, N2317, N885, N153);
not NOT1 (N2333, N2329);
or OR3 (N2334, N2333, N993, N285);
buf BUF1 (N2335, N2319);
and AND2 (N2336, N2323, N1278);
not NOT1 (N2337, N2335);
not NOT1 (N2338, N2336);
buf BUF1 (N2339, N2334);
nor NOR3 (N2340, N2313, N1090, N814);
and AND3 (N2341, N2340, N189, N756);
or OR2 (N2342, N2320, N1073);
or OR2 (N2343, N2339, N2204);
xor XOR2 (N2344, N2341, N2178);
buf BUF1 (N2345, N2338);
nor NOR4 (N2346, N2344, N407, N824, N695);
nand NAND4 (N2347, N2346, N1608, N1149, N1002);
nand NAND3 (N2348, N2330, N976, N704);
or OR2 (N2349, N2343, N941);
nand NAND4 (N2350, N2342, N1970, N783, N2233);
not NOT1 (N2351, N2337);
xor XOR2 (N2352, N2325, N1434);
nor NOR2 (N2353, N2348, N873);
buf BUF1 (N2354, N2347);
nand NAND3 (N2355, N2350, N2265, N2062);
or OR3 (N2356, N2332, N178, N275);
not NOT1 (N2357, N2349);
buf BUF1 (N2358, N2345);
nand NAND2 (N2359, N2356, N1488);
buf BUF1 (N2360, N2357);
buf BUF1 (N2361, N2354);
or OR4 (N2362, N2361, N1952, N857, N903);
nor NOR2 (N2363, N2355, N2117);
and AND4 (N2364, N2363, N261, N970, N949);
nand NAND3 (N2365, N2353, N521, N638);
and AND2 (N2366, N2310, N699);
nand NAND2 (N2367, N2351, N592);
not NOT1 (N2368, N2362);
and AND3 (N2369, N2364, N2193, N179);
nand NAND3 (N2370, N2358, N821, N207);
not NOT1 (N2371, N2359);
and AND3 (N2372, N2369, N2211, N1966);
not NOT1 (N2373, N2372);
xor XOR2 (N2374, N2371, N1583);
nand NAND2 (N2375, N2331, N300);
or OR2 (N2376, N2366, N1270);
not NOT1 (N2377, N2373);
not NOT1 (N2378, N2367);
buf BUF1 (N2379, N2375);
and AND2 (N2380, N2378, N2365);
or OR4 (N2381, N1109, N1230, N1319, N1428);
or OR2 (N2382, N2370, N1468);
nor NOR4 (N2383, N2360, N1651, N340, N566);
nand NAND2 (N2384, N2382, N1492);
nor NOR4 (N2385, N2379, N1715, N1781, N2136);
not NOT1 (N2386, N2352);
buf BUF1 (N2387, N2381);
nor NOR2 (N2388, N2376, N1728);
or OR3 (N2389, N2377, N1429, N2090);
nor NOR3 (N2390, N2383, N882, N1983);
not NOT1 (N2391, N2388);
or OR4 (N2392, N2391, N804, N827, N1806);
or OR2 (N2393, N2380, N843);
buf BUF1 (N2394, N2389);
nor NOR3 (N2395, N2390, N1270, N267);
xor XOR2 (N2396, N2395, N1579);
or OR3 (N2397, N2385, N1574, N723);
nand NAND3 (N2398, N2393, N1442, N1405);
or OR2 (N2399, N2397, N1953);
nor NOR2 (N2400, N2394, N1324);
or OR2 (N2401, N2398, N2370);
or OR2 (N2402, N2396, N1441);
and AND3 (N2403, N2401, N1439, N1793);
xor XOR2 (N2404, N2384, N2103);
nand NAND2 (N2405, N2403, N1976);
not NOT1 (N2406, N2400);
nor NOR3 (N2407, N2402, N1553, N837);
nand NAND2 (N2408, N2407, N703);
nand NAND4 (N2409, N2405, N892, N423, N1157);
buf BUF1 (N2410, N2374);
nand NAND2 (N2411, N2404, N1165);
not NOT1 (N2412, N2399);
not NOT1 (N2413, N2412);
nor NOR3 (N2414, N2387, N1783, N1739);
not NOT1 (N2415, N2409);
xor XOR2 (N2416, N2411, N50);
nand NAND3 (N2417, N2410, N1446, N815);
xor XOR2 (N2418, N2386, N140);
xor XOR2 (N2419, N2418, N850);
or OR3 (N2420, N2408, N1935, N934);
buf BUF1 (N2421, N2415);
buf BUF1 (N2422, N2413);
buf BUF1 (N2423, N2392);
not NOT1 (N2424, N2368);
buf BUF1 (N2425, N2421);
and AND4 (N2426, N2416, N2312, N1035, N255);
or OR3 (N2427, N2419, N2257, N1099);
buf BUF1 (N2428, N2417);
xor XOR2 (N2429, N2414, N204);
or OR3 (N2430, N2422, N628, N466);
nand NAND4 (N2431, N2427, N1068, N2327, N978);
or OR4 (N2432, N2429, N2287, N487, N1219);
nor NOR2 (N2433, N2428, N219);
nand NAND3 (N2434, N2425, N1214, N529);
xor XOR2 (N2435, N2424, N1218);
or OR2 (N2436, N2430, N2212);
not NOT1 (N2437, N2433);
and AND3 (N2438, N2420, N2222, N2345);
nor NOR2 (N2439, N2423, N504);
nor NOR4 (N2440, N2406, N732, N1976, N1732);
nand NAND3 (N2441, N2436, N935, N1586);
buf BUF1 (N2442, N2435);
and AND3 (N2443, N2440, N951, N1188);
and AND3 (N2444, N2441, N731, N616);
nand NAND2 (N2445, N2432, N450);
nand NAND3 (N2446, N2437, N62, N126);
nand NAND2 (N2447, N2445, N947);
nor NOR3 (N2448, N2426, N1995, N2256);
nand NAND3 (N2449, N2446, N1657, N642);
buf BUF1 (N2450, N2439);
buf BUF1 (N2451, N2443);
not NOT1 (N2452, N2449);
or OR4 (N2453, N2447, N723, N66, N1941);
nor NOR2 (N2454, N2452, N1020);
xor XOR2 (N2455, N2431, N2149);
buf BUF1 (N2456, N2442);
not NOT1 (N2457, N2451);
buf BUF1 (N2458, N2455);
not NOT1 (N2459, N2450);
nor NOR2 (N2460, N2457, N2155);
or OR4 (N2461, N2438, N920, N2066, N1501);
not NOT1 (N2462, N2456);
or OR2 (N2463, N2434, N1262);
not NOT1 (N2464, N2463);
or OR4 (N2465, N2464, N1497, N1046, N735);
not NOT1 (N2466, N2460);
xor XOR2 (N2467, N2454, N802);
buf BUF1 (N2468, N2462);
or OR3 (N2469, N2461, N1544, N37);
xor XOR2 (N2470, N2444, N662);
nand NAND2 (N2471, N2459, N964);
and AND2 (N2472, N2466, N2231);
buf BUF1 (N2473, N2469);
or OR3 (N2474, N2468, N540, N2344);
and AND2 (N2475, N2453, N1036);
nand NAND3 (N2476, N2471, N13, N2282);
not NOT1 (N2477, N2467);
xor XOR2 (N2478, N2470, N2116);
buf BUF1 (N2479, N2473);
not NOT1 (N2480, N2472);
and AND2 (N2481, N2474, N1941);
or OR2 (N2482, N2477, N1971);
buf BUF1 (N2483, N2480);
nor NOR4 (N2484, N2448, N1260, N1682, N2063);
nand NAND2 (N2485, N2483, N3);
or OR4 (N2486, N2485, N1346, N813, N1920);
or OR4 (N2487, N2458, N732, N1768, N960);
nor NOR4 (N2488, N2484, N1481, N353, N2144);
not NOT1 (N2489, N2475);
not NOT1 (N2490, N2476);
buf BUF1 (N2491, N2481);
xor XOR2 (N2492, N2488, N2028);
or OR2 (N2493, N2489, N1272);
or OR3 (N2494, N2486, N1368, N426);
and AND2 (N2495, N2493, N1295);
xor XOR2 (N2496, N2490, N801);
and AND4 (N2497, N2496, N2022, N1171, N2325);
not NOT1 (N2498, N2465);
xor XOR2 (N2499, N2497, N572);
nor NOR3 (N2500, N2494, N1196, N2404);
nor NOR4 (N2501, N2479, N479, N456, N1768);
nand NAND2 (N2502, N2498, N1542);
nand NAND3 (N2503, N2501, N1194, N815);
not NOT1 (N2504, N2482);
not NOT1 (N2505, N2487);
buf BUF1 (N2506, N2495);
nor NOR4 (N2507, N2505, N1440, N771, N1372);
and AND3 (N2508, N2503, N1866, N1447);
xor XOR2 (N2509, N2506, N261);
or OR2 (N2510, N2502, N1233);
nand NAND3 (N2511, N2478, N669, N1994);
nand NAND3 (N2512, N2511, N1592, N1868);
nor NOR2 (N2513, N2491, N1107);
nor NOR2 (N2514, N2507, N1515);
and AND2 (N2515, N2492, N2212);
not NOT1 (N2516, N2509);
not NOT1 (N2517, N2512);
nand NAND3 (N2518, N2504, N1090, N1120);
xor XOR2 (N2519, N2510, N2504);
and AND2 (N2520, N2515, N243);
not NOT1 (N2521, N2517);
not NOT1 (N2522, N2520);
nor NOR2 (N2523, N2500, N598);
xor XOR2 (N2524, N2508, N2389);
or OR2 (N2525, N2522, N2432);
nor NOR3 (N2526, N2523, N424, N2094);
nand NAND3 (N2527, N2526, N2380, N2222);
nand NAND4 (N2528, N2519, N295, N361, N272);
nor NOR3 (N2529, N2514, N383, N1205);
buf BUF1 (N2530, N2521);
xor XOR2 (N2531, N2525, N1966);
and AND4 (N2532, N2529, N1807, N100, N2441);
xor XOR2 (N2533, N2531, N1218);
nand NAND3 (N2534, N2513, N2520, N136);
and AND2 (N2535, N2516, N2159);
nand NAND3 (N2536, N2528, N37, N682);
and AND2 (N2537, N2533, N2295);
nor NOR2 (N2538, N2534, N1572);
not NOT1 (N2539, N2499);
and AND2 (N2540, N2537, N1900);
not NOT1 (N2541, N2532);
buf BUF1 (N2542, N2530);
and AND4 (N2543, N2527, N2096, N2429, N837);
nor NOR3 (N2544, N2524, N559, N1805);
not NOT1 (N2545, N2518);
and AND2 (N2546, N2540, N548);
and AND3 (N2547, N2538, N842, N478);
buf BUF1 (N2548, N2546);
or OR2 (N2549, N2542, N2094);
nand NAND3 (N2550, N2536, N772, N98);
and AND2 (N2551, N2544, N2037);
not NOT1 (N2552, N2551);
and AND2 (N2553, N2547, N2466);
not NOT1 (N2554, N2553);
not NOT1 (N2555, N2550);
not NOT1 (N2556, N2549);
nand NAND4 (N2557, N2556, N29, N49, N1405);
buf BUF1 (N2558, N2543);
nor NOR4 (N2559, N2545, N473, N643, N898);
not NOT1 (N2560, N2535);
not NOT1 (N2561, N2559);
and AND2 (N2562, N2548, N1370);
not NOT1 (N2563, N2552);
or OR3 (N2564, N2561, N815, N1311);
not NOT1 (N2565, N2564);
nor NOR4 (N2566, N2563, N1682, N2417, N1904);
not NOT1 (N2567, N2566);
nand NAND2 (N2568, N2555, N411);
not NOT1 (N2569, N2567);
not NOT1 (N2570, N2541);
nand NAND4 (N2571, N2560, N2506, N935, N1510);
buf BUF1 (N2572, N2569);
buf BUF1 (N2573, N2570);
xor XOR2 (N2574, N2568, N1355);
and AND2 (N2575, N2539, N2343);
and AND2 (N2576, N2557, N1791);
buf BUF1 (N2577, N2558);
xor XOR2 (N2578, N2554, N346);
not NOT1 (N2579, N2571);
or OR4 (N2580, N2576, N2405, N1891, N1465);
buf BUF1 (N2581, N2574);
nor NOR4 (N2582, N2578, N1307, N1090, N2536);
buf BUF1 (N2583, N2565);
nand NAND3 (N2584, N2575, N484, N537);
not NOT1 (N2585, N2580);
nor NOR4 (N2586, N2572, N1947, N2456, N1340);
or OR3 (N2587, N2573, N672, N2019);
and AND3 (N2588, N2583, N987, N1485);
and AND4 (N2589, N2586, N1322, N2351, N2256);
nand NAND2 (N2590, N2589, N2581);
or OR3 (N2591, N817, N300, N269);
nor NOR2 (N2592, N2585, N783);
nor NOR4 (N2593, N2590, N2274, N193, N238);
and AND3 (N2594, N2588, N238, N822);
not NOT1 (N2595, N2594);
nand NAND2 (N2596, N2579, N1535);
nor NOR3 (N2597, N2595, N2338, N2153);
nor NOR3 (N2598, N2597, N1691, N1953);
not NOT1 (N2599, N2577);
nand NAND2 (N2600, N2591, N777);
nand NAND3 (N2601, N2593, N555, N2506);
xor XOR2 (N2602, N2562, N1550);
not NOT1 (N2603, N2598);
or OR2 (N2604, N2599, N362);
buf BUF1 (N2605, N2600);
nand NAND4 (N2606, N2605, N1836, N92, N1309);
or OR3 (N2607, N2596, N1655, N1360);
not NOT1 (N2608, N2604);
or OR4 (N2609, N2584, N1830, N2558, N364);
buf BUF1 (N2610, N2602);
buf BUF1 (N2611, N2587);
and AND3 (N2612, N2592, N2009, N2110);
xor XOR2 (N2613, N2610, N646);
nor NOR3 (N2614, N2608, N1554, N239);
or OR2 (N2615, N2603, N381);
xor XOR2 (N2616, N2611, N2091);
not NOT1 (N2617, N2612);
and AND2 (N2618, N2617, N1094);
nor NOR2 (N2619, N2613, N245);
nand NAND4 (N2620, N2582, N1789, N794, N2340);
nor NOR3 (N2621, N2618, N809, N2594);
not NOT1 (N2622, N2606);
buf BUF1 (N2623, N2601);
buf BUF1 (N2624, N2607);
and AND2 (N2625, N2620, N1200);
or OR3 (N2626, N2625, N1790, N1229);
not NOT1 (N2627, N2616);
not NOT1 (N2628, N2609);
buf BUF1 (N2629, N2619);
nor NOR4 (N2630, N2627, N627, N1888, N2298);
and AND3 (N2631, N2630, N481, N352);
buf BUF1 (N2632, N2624);
xor XOR2 (N2633, N2626, N584);
not NOT1 (N2634, N2622);
xor XOR2 (N2635, N2615, N616);
and AND2 (N2636, N2634, N2372);
and AND2 (N2637, N2628, N1052);
not NOT1 (N2638, N2637);
buf BUF1 (N2639, N2614);
not NOT1 (N2640, N2635);
nor NOR4 (N2641, N2621, N1943, N2303, N835);
xor XOR2 (N2642, N2631, N1478);
not NOT1 (N2643, N2633);
not NOT1 (N2644, N2629);
nor NOR4 (N2645, N2636, N1139, N1206, N706);
buf BUF1 (N2646, N2632);
nor NOR2 (N2647, N2640, N739);
or OR2 (N2648, N2646, N422);
nor NOR3 (N2649, N2645, N1494, N395);
not NOT1 (N2650, N2647);
nand NAND2 (N2651, N2638, N308);
nor NOR2 (N2652, N2641, N754);
or OR4 (N2653, N2642, N1629, N547, N247);
xor XOR2 (N2654, N2644, N2274);
or OR2 (N2655, N2653, N37);
xor XOR2 (N2656, N2639, N2014);
or OR4 (N2657, N2652, N1503, N299, N1539);
not NOT1 (N2658, N2643);
xor XOR2 (N2659, N2648, N570);
nand NAND4 (N2660, N2623, N1414, N2193, N170);
nand NAND2 (N2661, N2657, N1330);
or OR4 (N2662, N2661, N2597, N774, N2461);
or OR4 (N2663, N2656, N554, N316, N1);
nand NAND2 (N2664, N2655, N2474);
xor XOR2 (N2665, N2660, N2518);
not NOT1 (N2666, N2651);
xor XOR2 (N2667, N2666, N517);
nor NOR4 (N2668, N2654, N1965, N1535, N1586);
nor NOR2 (N2669, N2658, N2597);
buf BUF1 (N2670, N2669);
not NOT1 (N2671, N2659);
nand NAND4 (N2672, N2667, N1276, N2349, N606);
and AND4 (N2673, N2663, N369, N2128, N167);
nand NAND3 (N2674, N2670, N2258, N256);
buf BUF1 (N2675, N2668);
or OR2 (N2676, N2675, N1960);
nand NAND4 (N2677, N2650, N2351, N2585, N2258);
not NOT1 (N2678, N2677);
xor XOR2 (N2679, N2678, N874);
xor XOR2 (N2680, N2676, N1032);
and AND3 (N2681, N2649, N57, N1885);
xor XOR2 (N2682, N2672, N1474);
not NOT1 (N2683, N2662);
not NOT1 (N2684, N2673);
nor NOR2 (N2685, N2665, N522);
or OR2 (N2686, N2671, N2276);
nand NAND4 (N2687, N2686, N961, N2590, N2153);
or OR3 (N2688, N2687, N744, N2433);
nor NOR3 (N2689, N2688, N1940, N576);
nor NOR4 (N2690, N2679, N839, N1250, N2393);
xor XOR2 (N2691, N2682, N608);
nand NAND4 (N2692, N2691, N2295, N342, N1063);
nand NAND4 (N2693, N2684, N1255, N1767, N1178);
or OR2 (N2694, N2681, N1888);
nand NAND2 (N2695, N2674, N2081);
nor NOR3 (N2696, N2683, N2418, N1941);
and AND4 (N2697, N2692, N67, N563, N553);
or OR2 (N2698, N2689, N744);
or OR4 (N2699, N2693, N1100, N2464, N304);
not NOT1 (N2700, N2680);
and AND2 (N2701, N2685, N2278);
nor NOR2 (N2702, N2699, N658);
and AND3 (N2703, N2700, N1126, N84);
not NOT1 (N2704, N2664);
not NOT1 (N2705, N2697);
or OR4 (N2706, N2694, N1687, N610, N1908);
buf BUF1 (N2707, N2704);
xor XOR2 (N2708, N2706, N2455);
nand NAND4 (N2709, N2698, N582, N2138, N243);
not NOT1 (N2710, N2707);
buf BUF1 (N2711, N2705);
buf BUF1 (N2712, N2709);
nor NOR2 (N2713, N2701, N1678);
nor NOR2 (N2714, N2690, N137);
xor XOR2 (N2715, N2714, N340);
xor XOR2 (N2716, N2711, N581);
not NOT1 (N2717, N2713);
nor NOR2 (N2718, N2703, N1143);
xor XOR2 (N2719, N2708, N776);
nor NOR4 (N2720, N2716, N506, N979, N68);
buf BUF1 (N2721, N2720);
and AND2 (N2722, N2710, N2136);
or OR3 (N2723, N2702, N1787, N1592);
or OR2 (N2724, N2721, N250);
nand NAND2 (N2725, N2719, N1492);
xor XOR2 (N2726, N2723, N1434);
nand NAND2 (N2727, N2717, N608);
and AND4 (N2728, N2696, N1067, N648, N1290);
not NOT1 (N2729, N2712);
xor XOR2 (N2730, N2722, N378);
and AND2 (N2731, N2725, N814);
and AND3 (N2732, N2731, N1460, N2658);
not NOT1 (N2733, N2727);
or OR3 (N2734, N2732, N332, N2536);
and AND4 (N2735, N2729, N2193, N1210, N1109);
and AND2 (N2736, N2730, N408);
not NOT1 (N2737, N2724);
nor NOR2 (N2738, N2733, N1333);
and AND2 (N2739, N2726, N890);
and AND4 (N2740, N2739, N1951, N236, N1706);
or OR2 (N2741, N2736, N100);
and AND4 (N2742, N2728, N1143, N1973, N1057);
buf BUF1 (N2743, N2695);
buf BUF1 (N2744, N2718);
or OR3 (N2745, N2715, N934, N157);
nand NAND2 (N2746, N2744, N1584);
not NOT1 (N2747, N2742);
nand NAND4 (N2748, N2747, N505, N2357, N2423);
or OR2 (N2749, N2734, N1683);
xor XOR2 (N2750, N2749, N624);
not NOT1 (N2751, N2746);
xor XOR2 (N2752, N2748, N37);
xor XOR2 (N2753, N2735, N1031);
and AND2 (N2754, N2738, N1337);
buf BUF1 (N2755, N2737);
or OR4 (N2756, N2751, N1964, N809, N2299);
nand NAND2 (N2757, N2756, N2107);
nand NAND2 (N2758, N2741, N548);
xor XOR2 (N2759, N2745, N1810);
nand NAND2 (N2760, N2752, N2414);
nor NOR3 (N2761, N2740, N1371, N2230);
nand NAND3 (N2762, N2755, N463, N172);
and AND2 (N2763, N2757, N1722);
nand NAND4 (N2764, N2762, N1050, N1714, N2634);
nor NOR3 (N2765, N2759, N1427, N1300);
nand NAND3 (N2766, N2765, N1668, N158);
xor XOR2 (N2767, N2758, N2137);
nand NAND2 (N2768, N2766, N155);
buf BUF1 (N2769, N2743);
and AND4 (N2770, N2753, N1153, N712, N64);
not NOT1 (N2771, N2770);
buf BUF1 (N2772, N2750);
and AND2 (N2773, N2767, N2285);
or OR4 (N2774, N2764, N2741, N1323, N1579);
or OR2 (N2775, N2768, N1629);
nand NAND3 (N2776, N2760, N85, N2286);
not NOT1 (N2777, N2771);
buf BUF1 (N2778, N2761);
nand NAND2 (N2779, N2772, N13);
nand NAND3 (N2780, N2774, N335, N2456);
not NOT1 (N2781, N2775);
buf BUF1 (N2782, N2763);
not NOT1 (N2783, N2781);
not NOT1 (N2784, N2782);
xor XOR2 (N2785, N2754, N2710);
xor XOR2 (N2786, N2778, N1394);
nor NOR3 (N2787, N2784, N945, N332);
nand NAND4 (N2788, N2785, N1063, N1872, N2076);
or OR3 (N2789, N2779, N1829, N717);
buf BUF1 (N2790, N2787);
xor XOR2 (N2791, N2788, N2306);
nor NOR4 (N2792, N2790, N989, N1412, N392);
buf BUF1 (N2793, N2786);
and AND2 (N2794, N2773, N1990);
nor NOR3 (N2795, N2783, N725, N2446);
nor NOR4 (N2796, N2792, N1008, N1042, N109);
nand NAND2 (N2797, N2780, N2495);
buf BUF1 (N2798, N2769);
nand NAND3 (N2799, N2795, N2513, N385);
not NOT1 (N2800, N2791);
xor XOR2 (N2801, N2794, N893);
and AND3 (N2802, N2776, N2161, N2557);
not NOT1 (N2803, N2798);
and AND3 (N2804, N2801, N1677, N1977);
xor XOR2 (N2805, N2796, N2622);
and AND3 (N2806, N2804, N1551, N2231);
nand NAND4 (N2807, N2793, N1985, N2480, N1224);
and AND3 (N2808, N2807, N2756, N414);
xor XOR2 (N2809, N2803, N5);
xor XOR2 (N2810, N2802, N2543);
nand NAND3 (N2811, N2809, N2127, N2760);
nor NOR4 (N2812, N2811, N1402, N126, N42);
xor XOR2 (N2813, N2805, N459);
and AND4 (N2814, N2813, N1316, N1984, N2805);
xor XOR2 (N2815, N2800, N188);
and AND2 (N2816, N2789, N1763);
xor XOR2 (N2817, N2799, N1985);
nand NAND3 (N2818, N2817, N108, N2743);
or OR3 (N2819, N2797, N2714, N2548);
xor XOR2 (N2820, N2812, N141);
or OR2 (N2821, N2777, N1294);
not NOT1 (N2822, N2818);
buf BUF1 (N2823, N2808);
not NOT1 (N2824, N2821);
and AND3 (N2825, N2816, N1988, N777);
and AND3 (N2826, N2806, N1317, N2766);
not NOT1 (N2827, N2824);
and AND2 (N2828, N2823, N1054);
and AND4 (N2829, N2814, N1968, N1669, N515);
or OR4 (N2830, N2826, N1892, N1066, N1050);
buf BUF1 (N2831, N2822);
not NOT1 (N2832, N2831);
nand NAND3 (N2833, N2819, N101, N2299);
not NOT1 (N2834, N2829);
xor XOR2 (N2835, N2828, N1070);
or OR3 (N2836, N2832, N2734, N526);
buf BUF1 (N2837, N2825);
and AND4 (N2838, N2830, N951, N216, N660);
buf BUF1 (N2839, N2815);
nor NOR4 (N2840, N2810, N2829, N121, N2796);
nand NAND3 (N2841, N2820, N2196, N2143);
nand NAND3 (N2842, N2833, N2027, N1439);
nor NOR3 (N2843, N2840, N1264, N138);
nor NOR3 (N2844, N2837, N430, N1053);
nor NOR2 (N2845, N2836, N386);
or OR4 (N2846, N2838, N2124, N2626, N1359);
and AND4 (N2847, N2844, N1736, N2756, N1111);
and AND3 (N2848, N2835, N1720, N1777);
xor XOR2 (N2849, N2846, N51);
nor NOR4 (N2850, N2839, N898, N320, N1779);
and AND3 (N2851, N2834, N2057, N2542);
nor NOR2 (N2852, N2841, N1112);
nor NOR2 (N2853, N2850, N416);
nand NAND2 (N2854, N2827, N1875);
and AND3 (N2855, N2843, N308, N1602);
nor NOR4 (N2856, N2854, N2293, N1819, N454);
nor NOR4 (N2857, N2842, N2315, N1126, N1500);
nand NAND2 (N2858, N2848, N1526);
not NOT1 (N2859, N2858);
buf BUF1 (N2860, N2847);
nand NAND3 (N2861, N2851, N1031, N195);
or OR4 (N2862, N2857, N891, N1635, N2006);
or OR3 (N2863, N2855, N2327, N270);
buf BUF1 (N2864, N2849);
or OR4 (N2865, N2856, N1123, N1038, N913);
not NOT1 (N2866, N2864);
and AND4 (N2867, N2865, N1963, N1468, N855);
or OR2 (N2868, N2866, N1985);
or OR3 (N2869, N2853, N1406, N1842);
or OR2 (N2870, N2867, N2319);
xor XOR2 (N2871, N2845, N1122);
buf BUF1 (N2872, N2868);
not NOT1 (N2873, N2863);
not NOT1 (N2874, N2859);
nand NAND2 (N2875, N2873, N2554);
or OR4 (N2876, N2875, N372, N1827, N2236);
not NOT1 (N2877, N2870);
nor NOR3 (N2878, N2877, N2719, N2690);
xor XOR2 (N2879, N2878, N192);
and AND2 (N2880, N2861, N2177);
or OR4 (N2881, N2872, N582, N102, N1618);
or OR2 (N2882, N2869, N2109);
or OR2 (N2883, N2871, N361);
or OR2 (N2884, N2879, N1408);
nand NAND2 (N2885, N2874, N2212);
or OR2 (N2886, N2881, N2659);
nor NOR4 (N2887, N2883, N1668, N2841, N104);
nor NOR4 (N2888, N2860, N1021, N748, N654);
nand NAND2 (N2889, N2885, N2266);
buf BUF1 (N2890, N2876);
not NOT1 (N2891, N2882);
xor XOR2 (N2892, N2888, N1776);
not NOT1 (N2893, N2862);
and AND4 (N2894, N2852, N2831, N2296, N255);
nor NOR4 (N2895, N2892, N2842, N1254, N830);
or OR4 (N2896, N2891, N2530, N929, N559);
xor XOR2 (N2897, N2894, N849);
not NOT1 (N2898, N2896);
xor XOR2 (N2899, N2884, N2721);
or OR4 (N2900, N2887, N2469, N1604, N1015);
nand NAND2 (N2901, N2895, N2649);
nor NOR2 (N2902, N2893, N351);
xor XOR2 (N2903, N2900, N2224);
or OR4 (N2904, N2902, N2755, N2879, N2177);
buf BUF1 (N2905, N2897);
not NOT1 (N2906, N2901);
nand NAND2 (N2907, N2899, N972);
nand NAND2 (N2908, N2903, N1273);
nor NOR2 (N2909, N2905, N589);
not NOT1 (N2910, N2889);
and AND4 (N2911, N2880, N2560, N2632, N127);
not NOT1 (N2912, N2886);
not NOT1 (N2913, N2908);
and AND4 (N2914, N2890, N1453, N64, N387);
or OR4 (N2915, N2909, N1377, N2470, N766);
not NOT1 (N2916, N2898);
xor XOR2 (N2917, N2910, N1569);
nand NAND4 (N2918, N2906, N2895, N2235, N882);
xor XOR2 (N2919, N2907, N773);
buf BUF1 (N2920, N2917);
nand NAND4 (N2921, N2914, N1043, N2201, N1306);
nand NAND4 (N2922, N2918, N1578, N2335, N2230);
not NOT1 (N2923, N2921);
nand NAND4 (N2924, N2913, N1808, N2848, N2817);
not NOT1 (N2925, N2916);
or OR2 (N2926, N2924, N1419);
not NOT1 (N2927, N2920);
buf BUF1 (N2928, N2904);
nand NAND4 (N2929, N2927, N1118, N2120, N928);
not NOT1 (N2930, N2915);
buf BUF1 (N2931, N2925);
not NOT1 (N2932, N2930);
buf BUF1 (N2933, N2922);
not NOT1 (N2934, N2932);
buf BUF1 (N2935, N2926);
xor XOR2 (N2936, N2931, N2444);
nand NAND3 (N2937, N2919, N2170, N1038);
nand NAND3 (N2938, N2911, N591, N472);
not NOT1 (N2939, N2928);
xor XOR2 (N2940, N2937, N1616);
nand NAND4 (N2941, N2935, N1266, N2285, N238);
not NOT1 (N2942, N2934);
nor NOR3 (N2943, N2938, N2699, N864);
xor XOR2 (N2944, N2929, N1206);
or OR4 (N2945, N2941, N1525, N2041, N1936);
buf BUF1 (N2946, N2945);
and AND3 (N2947, N2946, N699, N1251);
buf BUF1 (N2948, N2936);
xor XOR2 (N2949, N2942, N1187);
or OR2 (N2950, N2948, N681);
and AND3 (N2951, N2940, N2823, N1267);
nand NAND2 (N2952, N2950, N2435);
not NOT1 (N2953, N2951);
not NOT1 (N2954, N2947);
not NOT1 (N2955, N2944);
nor NOR4 (N2956, N2933, N1543, N628, N2115);
and AND4 (N2957, N2939, N2164, N710, N2873);
nand NAND4 (N2958, N2956, N390, N925, N1475);
nand NAND4 (N2959, N2949, N2910, N1445, N350);
xor XOR2 (N2960, N2943, N51);
nor NOR3 (N2961, N2952, N2288, N1223);
buf BUF1 (N2962, N2923);
not NOT1 (N2963, N2958);
not NOT1 (N2964, N2957);
xor XOR2 (N2965, N2962, N1425);
xor XOR2 (N2966, N2960, N2333);
nor NOR3 (N2967, N2966, N470, N2686);
nand NAND3 (N2968, N2963, N2745, N2025);
and AND2 (N2969, N2964, N1301);
or OR2 (N2970, N2912, N1134);
or OR3 (N2971, N2953, N1651, N2707);
buf BUF1 (N2972, N2959);
xor XOR2 (N2973, N2955, N1148);
and AND4 (N2974, N2970, N625, N1641, N2084);
nor NOR4 (N2975, N2974, N1797, N1183, N2869);
xor XOR2 (N2976, N2961, N1932);
xor XOR2 (N2977, N2968, N1434);
xor XOR2 (N2978, N2971, N2710);
xor XOR2 (N2979, N2978, N1310);
or OR3 (N2980, N2973, N1184, N2144);
or OR4 (N2981, N2979, N300, N1914, N1396);
or OR3 (N2982, N2977, N1455, N2005);
buf BUF1 (N2983, N2967);
or OR2 (N2984, N2976, N1668);
buf BUF1 (N2985, N2983);
or OR2 (N2986, N2982, N1139);
buf BUF1 (N2987, N2984);
and AND2 (N2988, N2954, N807);
xor XOR2 (N2989, N2981, N66);
nand NAND2 (N2990, N2989, N952);
and AND3 (N2991, N2975, N1839, N463);
xor XOR2 (N2992, N2986, N1295);
or OR3 (N2993, N2969, N2991, N2286);
not NOT1 (N2994, N2952);
not NOT1 (N2995, N2972);
not NOT1 (N2996, N2985);
buf BUF1 (N2997, N2992);
buf BUF1 (N2998, N2995);
not NOT1 (N2999, N2994);
nor NOR2 (N3000, N2965, N157);
or OR2 (N3001, N2999, N1607);
not NOT1 (N3002, N2990);
nand NAND4 (N3003, N3001, N906, N417, N1858);
buf BUF1 (N3004, N3000);
and AND3 (N3005, N2998, N985, N412);
not NOT1 (N3006, N3005);
buf BUF1 (N3007, N3003);
and AND3 (N3008, N2996, N1751, N1532);
nor NOR4 (N3009, N3006, N657, N173, N1020);
nand NAND2 (N3010, N3009, N954);
nand NAND3 (N3011, N2993, N2266, N2417);
not NOT1 (N3012, N3011);
buf BUF1 (N3013, N3008);
xor XOR2 (N3014, N3012, N510);
nor NOR3 (N3015, N3002, N2951, N2017);
nor NOR4 (N3016, N3004, N213, N2290, N2327);
not NOT1 (N3017, N3015);
nand NAND2 (N3018, N3013, N1025);
and AND2 (N3019, N2988, N2071);
buf BUF1 (N3020, N2980);
or OR3 (N3021, N3017, N2212, N1742);
buf BUF1 (N3022, N3014);
xor XOR2 (N3023, N3020, N1510);
not NOT1 (N3024, N2987);
not NOT1 (N3025, N3023);
xor XOR2 (N3026, N3022, N2758);
or OR4 (N3027, N3026, N757, N806, N749);
buf BUF1 (N3028, N3007);
xor XOR2 (N3029, N3028, N2579);
nand NAND2 (N3030, N3024, N464);
and AND3 (N3031, N3030, N25, N282);
not NOT1 (N3032, N2997);
or OR2 (N3033, N3019, N592);
not NOT1 (N3034, N3010);
or OR3 (N3035, N3034, N2438, N357);
buf BUF1 (N3036, N3016);
or OR2 (N3037, N3031, N2919);
buf BUF1 (N3038, N3029);
buf BUF1 (N3039, N3025);
xor XOR2 (N3040, N3035, N2313);
buf BUF1 (N3041, N3036);
buf BUF1 (N3042, N3021);
xor XOR2 (N3043, N3037, N2728);
nand NAND3 (N3044, N3038, N2928, N611);
not NOT1 (N3045, N3042);
xor XOR2 (N3046, N3032, N2925);
nand NAND2 (N3047, N3041, N198);
xor XOR2 (N3048, N3018, N1954);
xor XOR2 (N3049, N3044, N1383);
nand NAND3 (N3050, N3033, N2442, N1935);
or OR3 (N3051, N3047, N467, N1588);
nand NAND4 (N3052, N3049, N2386, N97, N2606);
not NOT1 (N3053, N3046);
or OR3 (N3054, N3027, N1232, N266);
xor XOR2 (N3055, N3052, N1762);
not NOT1 (N3056, N3045);
xor XOR2 (N3057, N3056, N1529);
not NOT1 (N3058, N3040);
not NOT1 (N3059, N3048);
not NOT1 (N3060, N3057);
nor NOR4 (N3061, N3051, N892, N707, N1318);
not NOT1 (N3062, N3039);
not NOT1 (N3063, N3053);
or OR3 (N3064, N3063, N1316, N520);
nand NAND3 (N3065, N3064, N2827, N2587);
and AND2 (N3066, N3062, N796);
not NOT1 (N3067, N3058);
buf BUF1 (N3068, N3059);
nor NOR3 (N3069, N3067, N1604, N1842);
nor NOR3 (N3070, N3065, N2202, N929);
or OR3 (N3071, N3043, N2245, N2091);
not NOT1 (N3072, N3068);
nand NAND4 (N3073, N3060, N1454, N2366, N440);
nor NOR2 (N3074, N3050, N737);
nor NOR4 (N3075, N3066, N2138, N2276, N2947);
buf BUF1 (N3076, N3055);
not NOT1 (N3077, N3070);
buf BUF1 (N3078, N3072);
not NOT1 (N3079, N3071);
buf BUF1 (N3080, N3079);
xor XOR2 (N3081, N3061, N825);
buf BUF1 (N3082, N3069);
buf BUF1 (N3083, N3074);
nand NAND3 (N3084, N3054, N2011, N1915);
or OR4 (N3085, N3081, N1441, N1559, N1832);
nor NOR2 (N3086, N3084, N1322);
nand NAND2 (N3087, N3086, N351);
not NOT1 (N3088, N3085);
nor NOR2 (N3089, N3078, N92);
nor NOR3 (N3090, N3089, N149, N1364);
and AND3 (N3091, N3087, N34, N1079);
and AND4 (N3092, N3083, N2641, N290, N3020);
not NOT1 (N3093, N3073);
buf BUF1 (N3094, N3092);
nor NOR4 (N3095, N3088, N1178, N77, N1490);
buf BUF1 (N3096, N3076);
or OR3 (N3097, N3095, N2609, N676);
buf BUF1 (N3098, N3094);
nor NOR2 (N3099, N3075, N1042);
and AND2 (N3100, N3082, N260);
not NOT1 (N3101, N3080);
and AND2 (N3102, N3100, N2503);
xor XOR2 (N3103, N3101, N200);
or OR2 (N3104, N3077, N946);
nand NAND4 (N3105, N3096, N743, N1168, N2606);
buf BUF1 (N3106, N3102);
nor NOR2 (N3107, N3097, N464);
and AND4 (N3108, N3107, N823, N2882, N1030);
buf BUF1 (N3109, N3098);
not NOT1 (N3110, N3091);
xor XOR2 (N3111, N3110, N1816);
nor NOR2 (N3112, N3090, N2993);
nor NOR3 (N3113, N3108, N76, N2096);
nand NAND2 (N3114, N3103, N2227);
nand NAND4 (N3115, N3111, N36, N1069, N1443);
buf BUF1 (N3116, N3106);
xor XOR2 (N3117, N3112, N1174);
xor XOR2 (N3118, N3115, N864);
nand NAND3 (N3119, N3116, N932, N621);
not NOT1 (N3120, N3117);
and AND3 (N3121, N3120, N2496, N493);
not NOT1 (N3122, N3104);
nor NOR2 (N3123, N3121, N47);
xor XOR2 (N3124, N3114, N3084);
not NOT1 (N3125, N3119);
nand NAND3 (N3126, N3099, N1693, N2533);
or OR4 (N3127, N3125, N646, N140, N602);
nand NAND2 (N3128, N3122, N1516);
or OR4 (N3129, N3124, N1872, N1543, N861);
nand NAND2 (N3130, N3129, N178);
buf BUF1 (N3131, N3105);
xor XOR2 (N3132, N3118, N1831);
buf BUF1 (N3133, N3131);
nand NAND3 (N3134, N3127, N1255, N1613);
nor NOR2 (N3135, N3132, N284);
buf BUF1 (N3136, N3135);
buf BUF1 (N3137, N3130);
or OR3 (N3138, N3123, N2269, N783);
not NOT1 (N3139, N3137);
nor NOR2 (N3140, N3126, N2650);
or OR2 (N3141, N3128, N1112);
buf BUF1 (N3142, N3113);
buf BUF1 (N3143, N3093);
xor XOR2 (N3144, N3109, N438);
buf BUF1 (N3145, N3144);
buf BUF1 (N3146, N3138);
or OR4 (N3147, N3140, N2257, N393, N21);
and AND3 (N3148, N3141, N1679, N2248);
or OR2 (N3149, N3136, N2980);
xor XOR2 (N3150, N3146, N466);
not NOT1 (N3151, N3143);
buf BUF1 (N3152, N3147);
and AND3 (N3153, N3148, N1885, N1412);
xor XOR2 (N3154, N3142, N662);
and AND2 (N3155, N3149, N503);
xor XOR2 (N3156, N3152, N2938);
nor NOR4 (N3157, N3153, N717, N2375, N593);
not NOT1 (N3158, N3139);
nor NOR4 (N3159, N3133, N2991, N693, N14);
or OR3 (N3160, N3155, N942, N2511);
buf BUF1 (N3161, N3160);
nor NOR2 (N3162, N3158, N1764);
not NOT1 (N3163, N3156);
nor NOR3 (N3164, N3134, N58, N2513);
not NOT1 (N3165, N3159);
and AND2 (N3166, N3161, N803);
not NOT1 (N3167, N3164);
nand NAND2 (N3168, N3162, N1650);
and AND3 (N3169, N3166, N2856, N2134);
or OR3 (N3170, N3163, N1632, N1369);
nor NOR3 (N3171, N3145, N2186, N2670);
or OR3 (N3172, N3169, N2054, N1678);
nor NOR2 (N3173, N3154, N1844);
nor NOR2 (N3174, N3157, N2485);
not NOT1 (N3175, N3151);
nor NOR4 (N3176, N3170, N1692, N1208, N2394);
or OR2 (N3177, N3171, N1748);
and AND3 (N3178, N3174, N2350, N1161);
xor XOR2 (N3179, N3178, N954);
and AND3 (N3180, N3167, N2709, N2889);
buf BUF1 (N3181, N3179);
or OR3 (N3182, N3165, N693, N801);
nand NAND3 (N3183, N3180, N1892, N700);
buf BUF1 (N3184, N3172);
not NOT1 (N3185, N3175);
and AND3 (N3186, N3181, N874, N1519);
not NOT1 (N3187, N3176);
buf BUF1 (N3188, N3150);
buf BUF1 (N3189, N3182);
or OR3 (N3190, N3185, N1010, N2816);
or OR3 (N3191, N3177, N135, N2031);
and AND2 (N3192, N3173, N696);
buf BUF1 (N3193, N3187);
not NOT1 (N3194, N3193);
nand NAND3 (N3195, N3183, N1721, N2806);
not NOT1 (N3196, N3189);
or OR4 (N3197, N3190, N2618, N3058, N2211);
not NOT1 (N3198, N3192);
xor XOR2 (N3199, N3186, N1411);
nand NAND3 (N3200, N3194, N332, N890);
nand NAND2 (N3201, N3184, N3028);
and AND2 (N3202, N3195, N976);
xor XOR2 (N3203, N3188, N174);
or OR4 (N3204, N3200, N2585, N1300, N672);
or OR2 (N3205, N3204, N3070);
nand NAND4 (N3206, N3203, N729, N2898, N449);
buf BUF1 (N3207, N3198);
nand NAND4 (N3208, N3191, N2311, N2513, N1312);
or OR4 (N3209, N3202, N3016, N812, N620);
nor NOR2 (N3210, N3168, N2960);
xor XOR2 (N3211, N3196, N1887);
or OR3 (N3212, N3197, N291, N1145);
buf BUF1 (N3213, N3208);
nand NAND4 (N3214, N3212, N621, N1626, N2998);
xor XOR2 (N3215, N3209, N907);
not NOT1 (N3216, N3211);
not NOT1 (N3217, N3205);
or OR4 (N3218, N3217, N2104, N321, N1179);
not NOT1 (N3219, N3214);
not NOT1 (N3220, N3213);
nand NAND2 (N3221, N3220, N348);
not NOT1 (N3222, N3201);
buf BUF1 (N3223, N3222);
or OR3 (N3224, N3210, N1541, N844);
xor XOR2 (N3225, N3199, N1277);
nand NAND4 (N3226, N3224, N3043, N3179, N530);
not NOT1 (N3227, N3206);
or OR4 (N3228, N3219, N1059, N1162, N33);
nand NAND4 (N3229, N3223, N2351, N227, N2002);
buf BUF1 (N3230, N3215);
not NOT1 (N3231, N3216);
xor XOR2 (N3232, N3228, N3115);
xor XOR2 (N3233, N3227, N2771);
nor NOR3 (N3234, N3226, N998, N1034);
or OR3 (N3235, N3234, N2651, N2634);
not NOT1 (N3236, N3218);
nand NAND4 (N3237, N3221, N423, N1132, N1716);
xor XOR2 (N3238, N3232, N2776);
xor XOR2 (N3239, N3233, N2420);
or OR4 (N3240, N3229, N783, N2388, N1036);
not NOT1 (N3241, N3207);
buf BUF1 (N3242, N3231);
nor NOR2 (N3243, N3242, N2142);
nor NOR3 (N3244, N3237, N2367, N2882);
or OR2 (N3245, N3225, N1757);
nand NAND2 (N3246, N3244, N1627);
nand NAND4 (N3247, N3240, N1316, N1597, N1693);
xor XOR2 (N3248, N3241, N3034);
xor XOR2 (N3249, N3248, N1084);
nor NOR3 (N3250, N3245, N785, N2975);
xor XOR2 (N3251, N3239, N253);
and AND3 (N3252, N3230, N2535, N2801);
and AND2 (N3253, N3247, N1774);
xor XOR2 (N3254, N3249, N1196);
not NOT1 (N3255, N3252);
not NOT1 (N3256, N3255);
xor XOR2 (N3257, N3235, N1501);
xor XOR2 (N3258, N3251, N226);
nor NOR2 (N3259, N3246, N197);
buf BUF1 (N3260, N3257);
or OR3 (N3261, N3260, N764, N1981);
nand NAND3 (N3262, N3253, N3072, N2414);
xor XOR2 (N3263, N3256, N2085);
and AND3 (N3264, N3254, N570, N1596);
buf BUF1 (N3265, N3236);
nand NAND3 (N3266, N3243, N1731, N1387);
nor NOR4 (N3267, N3264, N875, N2926, N585);
xor XOR2 (N3268, N3238, N2724);
buf BUF1 (N3269, N3263);
not NOT1 (N3270, N3259);
or OR4 (N3271, N3265, N3063, N2523, N2327);
nand NAND4 (N3272, N3269, N101, N24, N2541);
nand NAND4 (N3273, N3266, N356, N723, N1607);
buf BUF1 (N3274, N3268);
and AND2 (N3275, N3267, N2792);
xor XOR2 (N3276, N3270, N1518);
xor XOR2 (N3277, N3250, N2929);
nor NOR4 (N3278, N3272, N1310, N242, N471);
buf BUF1 (N3279, N3276);
nand NAND2 (N3280, N3261, N344);
or OR2 (N3281, N3278, N2613);
not NOT1 (N3282, N3277);
and AND4 (N3283, N3271, N67, N1561, N432);
not NOT1 (N3284, N3275);
xor XOR2 (N3285, N3282, N2852);
xor XOR2 (N3286, N3280, N2357);
xor XOR2 (N3287, N3258, N2562);
buf BUF1 (N3288, N3285);
or OR3 (N3289, N3279, N862, N2112);
nor NOR2 (N3290, N3289, N1534);
or OR3 (N3291, N3274, N483, N2760);
not NOT1 (N3292, N3262);
and AND2 (N3293, N3273, N2892);
xor XOR2 (N3294, N3293, N1621);
nand NAND3 (N3295, N3290, N2212, N3191);
not NOT1 (N3296, N3292);
and AND4 (N3297, N3281, N2721, N589, N1967);
nor NOR4 (N3298, N3291, N1928, N1421, N2741);
nor NOR4 (N3299, N3296, N2265, N600, N3161);
not NOT1 (N3300, N3298);
nor NOR2 (N3301, N3288, N1801);
not NOT1 (N3302, N3300);
not NOT1 (N3303, N3295);
nor NOR2 (N3304, N3286, N586);
not NOT1 (N3305, N3297);
not NOT1 (N3306, N3299);
or OR4 (N3307, N3304, N1117, N867, N807);
xor XOR2 (N3308, N3307, N515);
nand NAND4 (N3309, N3283, N1367, N2562, N940);
or OR4 (N3310, N3306, N2405, N1730, N1189);
or OR3 (N3311, N3303, N1908, N1909);
or OR3 (N3312, N3294, N1776, N1641);
xor XOR2 (N3313, N3287, N145);
or OR2 (N3314, N3309, N3242);
not NOT1 (N3315, N3301);
not NOT1 (N3316, N3284);
buf BUF1 (N3317, N3311);
or OR2 (N3318, N3313, N1518);
and AND3 (N3319, N3318, N1664, N275);
or OR3 (N3320, N3310, N1156, N791);
buf BUF1 (N3321, N3314);
and AND2 (N3322, N3302, N2944);
xor XOR2 (N3323, N3312, N1912);
nor NOR3 (N3324, N3317, N2222, N1567);
and AND4 (N3325, N3324, N1453, N3290, N2636);
not NOT1 (N3326, N3315);
or OR2 (N3327, N3326, N509);
xor XOR2 (N3328, N3320, N2387);
or OR3 (N3329, N3322, N1584, N2732);
nor NOR2 (N3330, N3323, N2779);
and AND3 (N3331, N3327, N2699, N2668);
nand NAND4 (N3332, N3319, N1417, N2483, N448);
buf BUF1 (N3333, N3305);
and AND3 (N3334, N3330, N2906, N1503);
nand NAND3 (N3335, N3321, N1360, N711);
or OR4 (N3336, N3332, N3136, N1636, N486);
nand NAND2 (N3337, N3325, N3112);
nand NAND3 (N3338, N3331, N100, N3311);
nand NAND4 (N3339, N3328, N883, N812, N725);
nand NAND3 (N3340, N3333, N355, N574);
or OR3 (N3341, N3308, N2021, N2968);
xor XOR2 (N3342, N3339, N2125);
not NOT1 (N3343, N3316);
xor XOR2 (N3344, N3336, N2722);
nand NAND4 (N3345, N3338, N2802, N2370, N578);
and AND2 (N3346, N3342, N2707);
nand NAND4 (N3347, N3340, N1053, N1443, N469);
or OR4 (N3348, N3346, N1944, N2904, N3279);
nor NOR3 (N3349, N3348, N686, N1385);
not NOT1 (N3350, N3343);
nor NOR4 (N3351, N3350, N335, N3156, N2176);
buf BUF1 (N3352, N3344);
not NOT1 (N3353, N3345);
nand NAND4 (N3354, N3352, N2509, N2616, N2502);
buf BUF1 (N3355, N3347);
buf BUF1 (N3356, N3351);
not NOT1 (N3357, N3334);
not NOT1 (N3358, N3335);
and AND2 (N3359, N3341, N1297);
buf BUF1 (N3360, N3349);
not NOT1 (N3361, N3337);
not NOT1 (N3362, N3359);
buf BUF1 (N3363, N3358);
nor NOR2 (N3364, N3362, N3344);
buf BUF1 (N3365, N3353);
xor XOR2 (N3366, N3356, N2593);
or OR2 (N3367, N3363, N2115);
and AND2 (N3368, N3354, N2121);
and AND3 (N3369, N3329, N308, N3286);
nand NAND3 (N3370, N3369, N174, N1037);
nand NAND2 (N3371, N3367, N1289);
nor NOR4 (N3372, N3366, N2148, N1746, N1478);
nor NOR4 (N3373, N3365, N1263, N1876, N3225);
and AND4 (N3374, N3368, N875, N707, N2214);
and AND3 (N3375, N3360, N29, N1967);
nand NAND3 (N3376, N3370, N2301, N524);
or OR2 (N3377, N3364, N2466);
xor XOR2 (N3378, N3373, N337);
nand NAND2 (N3379, N3374, N2674);
buf BUF1 (N3380, N3361);
and AND3 (N3381, N3379, N1794, N1547);
and AND4 (N3382, N3381, N3121, N967, N1239);
nand NAND3 (N3383, N3355, N1866, N2344);
xor XOR2 (N3384, N3372, N734);
buf BUF1 (N3385, N3378);
and AND3 (N3386, N3357, N45, N2802);
and AND3 (N3387, N3385, N1253, N911);
and AND3 (N3388, N3387, N1298, N978);
or OR2 (N3389, N3382, N2556);
not NOT1 (N3390, N3371);
xor XOR2 (N3391, N3376, N529);
nor NOR4 (N3392, N3375, N2459, N793, N2712);
buf BUF1 (N3393, N3377);
not NOT1 (N3394, N3392);
or OR4 (N3395, N3390, N953, N3159, N2131);
nand NAND3 (N3396, N3380, N3092, N1810);
and AND2 (N3397, N3386, N2735);
xor XOR2 (N3398, N3396, N2180);
xor XOR2 (N3399, N3389, N1915);
nand NAND4 (N3400, N3384, N2899, N1845, N1529);
buf BUF1 (N3401, N3383);
nand NAND2 (N3402, N3400, N2918);
not NOT1 (N3403, N3398);
and AND3 (N3404, N3395, N2895, N407);
and AND3 (N3405, N3397, N2716, N518);
not NOT1 (N3406, N3391);
or OR3 (N3407, N3394, N2354, N332);
buf BUF1 (N3408, N3402);
buf BUF1 (N3409, N3388);
nand NAND3 (N3410, N3409, N2685, N3185);
nand NAND2 (N3411, N3407, N1923);
not NOT1 (N3412, N3404);
xor XOR2 (N3413, N3393, N2325);
or OR3 (N3414, N3405, N2355, N3316);
or OR2 (N3415, N3401, N2765);
or OR4 (N3416, N3403, N1372, N3377, N2339);
nor NOR4 (N3417, N3399, N1992, N3114, N508);
not NOT1 (N3418, N3414);
and AND2 (N3419, N3411, N1907);
not NOT1 (N3420, N3406);
not NOT1 (N3421, N3410);
buf BUF1 (N3422, N3418);
xor XOR2 (N3423, N3417, N2940);
nand NAND2 (N3424, N3408, N2760);
and AND2 (N3425, N3422, N2626);
xor XOR2 (N3426, N3416, N775);
or OR2 (N3427, N3420, N2660);
and AND2 (N3428, N3419, N3273);
xor XOR2 (N3429, N3413, N2926);
nand NAND2 (N3430, N3429, N2370);
xor XOR2 (N3431, N3412, N772);
xor XOR2 (N3432, N3427, N2102);
nor NOR2 (N3433, N3428, N2732);
and AND3 (N3434, N3433, N2044, N431);
buf BUF1 (N3435, N3423);
nand NAND3 (N3436, N3432, N2237, N2087);
xor XOR2 (N3437, N3425, N1646);
buf BUF1 (N3438, N3421);
and AND3 (N3439, N3434, N1361, N2177);
nor NOR3 (N3440, N3424, N1249, N926);
nand NAND3 (N3441, N3431, N2140, N377);
buf BUF1 (N3442, N3437);
xor XOR2 (N3443, N3439, N1161);
nor NOR2 (N3444, N3426, N1813);
buf BUF1 (N3445, N3440);
nand NAND2 (N3446, N3436, N209);
buf BUF1 (N3447, N3435);
buf BUF1 (N3448, N3443);
nand NAND4 (N3449, N3448, N19, N538, N1004);
and AND3 (N3450, N3415, N409, N1946);
and AND4 (N3451, N3441, N1675, N3181, N1769);
and AND3 (N3452, N3445, N428, N3369);
buf BUF1 (N3453, N3442);
or OR4 (N3454, N3430, N2636, N2030, N1921);
buf BUF1 (N3455, N3450);
xor XOR2 (N3456, N3447, N1532);
nand NAND2 (N3457, N3452, N3365);
and AND4 (N3458, N3456, N100, N1278, N1892);
nand NAND3 (N3459, N3454, N2577, N775);
and AND2 (N3460, N3451, N1849);
and AND4 (N3461, N3460, N1261, N3417, N850);
or OR3 (N3462, N3459, N1992, N2494);
buf BUF1 (N3463, N3462);
and AND3 (N3464, N3453, N1205, N1080);
or OR4 (N3465, N3458, N3241, N1919, N68);
buf BUF1 (N3466, N3446);
buf BUF1 (N3467, N3444);
buf BUF1 (N3468, N3457);
nand NAND3 (N3469, N3465, N2692, N423);
or OR4 (N3470, N3464, N1355, N2794, N1917);
buf BUF1 (N3471, N3449);
nand NAND3 (N3472, N3463, N862, N1034);
nand NAND3 (N3473, N3438, N1932, N1497);
buf BUF1 (N3474, N3472);
nand NAND3 (N3475, N3467, N11, N46);
not NOT1 (N3476, N3461);
buf BUF1 (N3477, N3470);
nor NOR3 (N3478, N3466, N919, N1299);
and AND4 (N3479, N3469, N2126, N1327, N1449);
xor XOR2 (N3480, N3479, N1067);
nor NOR2 (N3481, N3478, N2114);
nand NAND2 (N3482, N3475, N2186);
or OR2 (N3483, N3474, N2578);
buf BUF1 (N3484, N3480);
nor NOR3 (N3485, N3468, N2560, N650);
nor NOR2 (N3486, N3483, N3327);
and AND4 (N3487, N3455, N1376, N2205, N2023);
nor NOR3 (N3488, N3486, N504, N1287);
nand NAND2 (N3489, N3485, N450);
or OR3 (N3490, N3488, N1356, N288);
not NOT1 (N3491, N3482);
buf BUF1 (N3492, N3489);
xor XOR2 (N3493, N3471, N3003);
xor XOR2 (N3494, N3476, N1975);
nand NAND2 (N3495, N3477, N1876);
nor NOR4 (N3496, N3490, N1783, N92, N2212);
buf BUF1 (N3497, N3496);
or OR4 (N3498, N3497, N3124, N3051, N1069);
nor NOR2 (N3499, N3481, N2);
or OR4 (N3500, N3484, N3023, N641, N2892);
not NOT1 (N3501, N3491);
nand NAND3 (N3502, N3487, N791, N110);
nor NOR4 (N3503, N3494, N1874, N1615, N2035);
buf BUF1 (N3504, N3501);
not NOT1 (N3505, N3473);
nor NOR3 (N3506, N3500, N2312, N2684);
nor NOR4 (N3507, N3503, N2532, N2294, N1040);
and AND3 (N3508, N3492, N1723, N2789);
not NOT1 (N3509, N3502);
not NOT1 (N3510, N3504);
nand NAND2 (N3511, N3498, N2627);
not NOT1 (N3512, N3508);
nor NOR4 (N3513, N3493, N1867, N2030, N3038);
nor NOR4 (N3514, N3513, N1472, N1990, N3123);
nor NOR4 (N3515, N3512, N3081, N3132, N1058);
xor XOR2 (N3516, N3510, N3455);
buf BUF1 (N3517, N3499);
nand NAND3 (N3518, N3516, N3030, N1512);
buf BUF1 (N3519, N3495);
or OR3 (N3520, N3515, N1120, N968);
or OR4 (N3521, N3505, N1725, N2789, N1303);
buf BUF1 (N3522, N3506);
and AND2 (N3523, N3509, N143);
xor XOR2 (N3524, N3520, N2090);
nor NOR4 (N3525, N3519, N2710, N1888, N3424);
nor NOR2 (N3526, N3514, N1148);
nor NOR2 (N3527, N3525, N3267);
nor NOR4 (N3528, N3518, N1654, N2845, N812);
xor XOR2 (N3529, N3511, N676);
nor NOR2 (N3530, N3526, N1818);
buf BUF1 (N3531, N3521);
nor NOR2 (N3532, N3524, N1472);
xor XOR2 (N3533, N3517, N2885);
nand NAND2 (N3534, N3531, N2139);
nand NAND2 (N3535, N3530, N1313);
or OR4 (N3536, N3507, N1770, N2844, N851);
and AND4 (N3537, N3534, N2980, N978, N2494);
not NOT1 (N3538, N3532);
buf BUF1 (N3539, N3537);
nand NAND4 (N3540, N3522, N3000, N726, N1711);
nor NOR4 (N3541, N3528, N801, N269, N1199);
xor XOR2 (N3542, N3523, N1766);
nand NAND4 (N3543, N3541, N3180, N824, N2018);
not NOT1 (N3544, N3538);
xor XOR2 (N3545, N3540, N2158);
and AND2 (N3546, N3527, N2434);
and AND2 (N3547, N3535, N3121);
nand NAND3 (N3548, N3545, N2553, N1603);
or OR2 (N3549, N3529, N2522);
or OR2 (N3550, N3536, N1378);
or OR2 (N3551, N3533, N2697);
nand NAND2 (N3552, N3549, N2783);
nor NOR3 (N3553, N3539, N2806, N1579);
or OR2 (N3554, N3542, N3208);
buf BUF1 (N3555, N3550);
buf BUF1 (N3556, N3555);
nor NOR3 (N3557, N3543, N15, N2195);
not NOT1 (N3558, N3551);
nor NOR3 (N3559, N3547, N1314, N2653);
buf BUF1 (N3560, N3546);
or OR4 (N3561, N3553, N2309, N928, N2998);
nand NAND4 (N3562, N3552, N737, N2862, N181);
nor NOR2 (N3563, N3557, N2449);
or OR3 (N3564, N3548, N3327, N3071);
buf BUF1 (N3565, N3556);
or OR3 (N3566, N3563, N3129, N221);
buf BUF1 (N3567, N3560);
nor NOR4 (N3568, N3562, N3399, N1760, N1398);
nand NAND2 (N3569, N3558, N1685);
and AND3 (N3570, N3565, N2349, N2459);
and AND3 (N3571, N3566, N617, N1510);
xor XOR2 (N3572, N3571, N1679);
nand NAND4 (N3573, N3570, N3562, N2731, N801);
or OR2 (N3574, N3559, N364);
xor XOR2 (N3575, N3572, N1274);
not NOT1 (N3576, N3561);
and AND3 (N3577, N3568, N2873, N2015);
nand NAND4 (N3578, N3554, N2261, N2061, N2593);
not NOT1 (N3579, N3576);
nor NOR3 (N3580, N3569, N1623, N1585);
xor XOR2 (N3581, N3544, N1136);
buf BUF1 (N3582, N3577);
nand NAND4 (N3583, N3580, N572, N1528, N2161);
xor XOR2 (N3584, N3579, N2765);
xor XOR2 (N3585, N3581, N3467);
xor XOR2 (N3586, N3567, N767);
xor XOR2 (N3587, N3585, N1282);
or OR2 (N3588, N3582, N2255);
xor XOR2 (N3589, N3564, N676);
and AND2 (N3590, N3588, N3101);
nor NOR3 (N3591, N3586, N3430, N357);
buf BUF1 (N3592, N3583);
nand NAND3 (N3593, N3592, N1655, N3050);
nor NOR2 (N3594, N3573, N1394);
and AND4 (N3595, N3590, N1103, N2582, N2258);
or OR2 (N3596, N3575, N306);
xor XOR2 (N3597, N3587, N3497);
xor XOR2 (N3598, N3594, N3363);
nand NAND2 (N3599, N3578, N2102);
nor NOR4 (N3600, N3599, N1070, N3, N3513);
nand NAND2 (N3601, N3589, N2494);
or OR2 (N3602, N3601, N1998);
or OR2 (N3603, N3597, N2501);
or OR2 (N3604, N3591, N386);
nand NAND4 (N3605, N3574, N1016, N2724, N2187);
not NOT1 (N3606, N3605);
or OR3 (N3607, N3593, N1578, N477);
not NOT1 (N3608, N3596);
xor XOR2 (N3609, N3608, N251);
not NOT1 (N3610, N3602);
or OR3 (N3611, N3584, N377, N1684);
not NOT1 (N3612, N3611);
xor XOR2 (N3613, N3606, N2874);
nor NOR4 (N3614, N3612, N389, N2788, N1445);
or OR4 (N3615, N3604, N2597, N1045, N1293);
xor XOR2 (N3616, N3598, N14);
buf BUF1 (N3617, N3609);
or OR3 (N3618, N3613, N454, N1548);
or OR2 (N3619, N3614, N2898);
or OR3 (N3620, N3615, N1346, N3010);
nor NOR2 (N3621, N3619, N533);
nand NAND4 (N3622, N3616, N313, N787, N2898);
xor XOR2 (N3623, N3618, N3272);
buf BUF1 (N3624, N3607);
nand NAND2 (N3625, N3603, N1519);
nand NAND3 (N3626, N3624, N1711, N3605);
not NOT1 (N3627, N3623);
nand NAND3 (N3628, N3627, N1969, N2049);
nor NOR4 (N3629, N3625, N2947, N3366, N143);
or OR2 (N3630, N3629, N2552);
not NOT1 (N3631, N3617);
nor NOR2 (N3632, N3631, N2432);
xor XOR2 (N3633, N3610, N2721);
or OR3 (N3634, N3630, N1546, N1335);
not NOT1 (N3635, N3600);
and AND2 (N3636, N3632, N1039);
nand NAND3 (N3637, N3628, N121, N2030);
not NOT1 (N3638, N3633);
nand NAND3 (N3639, N3637, N3633, N894);
and AND2 (N3640, N3626, N1655);
xor XOR2 (N3641, N3620, N942);
nor NOR3 (N3642, N3595, N1106, N1067);
buf BUF1 (N3643, N3641);
buf BUF1 (N3644, N3640);
nand NAND3 (N3645, N3639, N3517, N2137);
or OR3 (N3646, N3635, N2327, N295);
not NOT1 (N3647, N3645);
not NOT1 (N3648, N3622);
or OR3 (N3649, N3648, N621, N2675);
nor NOR2 (N3650, N3634, N2789);
nand NAND2 (N3651, N3642, N1314);
nor NOR3 (N3652, N3651, N32, N1590);
or OR2 (N3653, N3621, N739);
nor NOR3 (N3654, N3650, N2800, N1966);
and AND2 (N3655, N3653, N7);
and AND4 (N3656, N3647, N723, N3616, N3624);
nand NAND4 (N3657, N3652, N3341, N2151, N287);
or OR3 (N3658, N3657, N449, N2901);
nand NAND4 (N3659, N3643, N391, N1974, N1552);
or OR4 (N3660, N3656, N196, N2520, N1994);
nand NAND4 (N3661, N3659, N3316, N528, N22);
buf BUF1 (N3662, N3655);
nand NAND3 (N3663, N3646, N1385, N1475);
xor XOR2 (N3664, N3658, N1076);
xor XOR2 (N3665, N3661, N1403);
nor NOR2 (N3666, N3654, N1405);
nand NAND3 (N3667, N3664, N2116, N3010);
xor XOR2 (N3668, N3660, N1034);
or OR4 (N3669, N3636, N497, N2091, N598);
nor NOR2 (N3670, N3663, N3279);
nand NAND2 (N3671, N3667, N1254);
xor XOR2 (N3672, N3665, N2797);
xor XOR2 (N3673, N3666, N2381);
and AND2 (N3674, N3649, N3355);
or OR3 (N3675, N3644, N477, N2164);
buf BUF1 (N3676, N3671);
not NOT1 (N3677, N3669);
nor NOR2 (N3678, N3674, N2529);
not NOT1 (N3679, N3638);
xor XOR2 (N3680, N3678, N3041);
buf BUF1 (N3681, N3676);
not NOT1 (N3682, N3677);
and AND4 (N3683, N3675, N40, N1876, N2740);
and AND4 (N3684, N3673, N2101, N552, N2460);
not NOT1 (N3685, N3679);
or OR2 (N3686, N3680, N3319);
nand NAND4 (N3687, N3683, N2488, N2895, N2585);
xor XOR2 (N3688, N3668, N2042);
or OR2 (N3689, N3672, N2076);
nand NAND2 (N3690, N3687, N1865);
nor NOR3 (N3691, N3685, N2652, N3084);
or OR2 (N3692, N3688, N196);
nor NOR3 (N3693, N3689, N579, N3397);
and AND2 (N3694, N3681, N439);
not NOT1 (N3695, N3684);
not NOT1 (N3696, N3690);
nor NOR3 (N3697, N3696, N110, N178);
xor XOR2 (N3698, N3694, N2915);
not NOT1 (N3699, N3697);
nand NAND2 (N3700, N3662, N3361);
buf BUF1 (N3701, N3670);
nor NOR2 (N3702, N3695, N3614);
buf BUF1 (N3703, N3700);
and AND3 (N3704, N3701, N2298, N2749);
xor XOR2 (N3705, N3698, N3496);
and AND4 (N3706, N3686, N1323, N3399, N2913);
buf BUF1 (N3707, N3699);
nor NOR3 (N3708, N3692, N1153, N647);
not NOT1 (N3709, N3693);
buf BUF1 (N3710, N3691);
buf BUF1 (N3711, N3705);
buf BUF1 (N3712, N3709);
nor NOR3 (N3713, N3712, N1536, N1562);
buf BUF1 (N3714, N3707);
xor XOR2 (N3715, N3682, N1512);
or OR2 (N3716, N3713, N2636);
xor XOR2 (N3717, N3708, N911);
not NOT1 (N3718, N3704);
and AND2 (N3719, N3717, N1098);
buf BUF1 (N3720, N3718);
or OR2 (N3721, N3703, N3295);
and AND4 (N3722, N3719, N3028, N79, N149);
buf BUF1 (N3723, N3716);
nor NOR2 (N3724, N3715, N950);
xor XOR2 (N3725, N3706, N720);
buf BUF1 (N3726, N3722);
and AND2 (N3727, N3725, N2870);
nand NAND3 (N3728, N3727, N2671, N1653);
or OR3 (N3729, N3721, N921, N399);
nand NAND2 (N3730, N3726, N1943);
or OR3 (N3731, N3723, N3700, N128);
or OR3 (N3732, N3728, N738, N3518);
nand NAND3 (N3733, N3731, N2230, N3036);
or OR4 (N3734, N3729, N2280, N604, N2664);
xor XOR2 (N3735, N3711, N1496);
nor NOR3 (N3736, N3734, N709, N746);
nand NAND3 (N3737, N3702, N2845, N1285);
buf BUF1 (N3738, N3732);
xor XOR2 (N3739, N3724, N1991);
nor NOR4 (N3740, N3735, N3286, N3172, N3490);
not NOT1 (N3741, N3733);
and AND3 (N3742, N3720, N1028, N257);
buf BUF1 (N3743, N3738);
nand NAND3 (N3744, N3742, N2450, N1557);
nand NAND4 (N3745, N3714, N2481, N2787, N3087);
not NOT1 (N3746, N3730);
nor NOR4 (N3747, N3737, N1514, N2467, N247);
not NOT1 (N3748, N3740);
nand NAND3 (N3749, N3741, N3074, N1043);
nand NAND4 (N3750, N3746, N1266, N1775, N2734);
buf BUF1 (N3751, N3736);
not NOT1 (N3752, N3750);
buf BUF1 (N3753, N3739);
and AND4 (N3754, N3751, N2195, N2418, N1478);
nand NAND3 (N3755, N3748, N2816, N2526);
buf BUF1 (N3756, N3755);
or OR2 (N3757, N3744, N759);
buf BUF1 (N3758, N3756);
nor NOR3 (N3759, N3758, N3646, N890);
buf BUF1 (N3760, N3743);
not NOT1 (N3761, N3710);
xor XOR2 (N3762, N3752, N3400);
nand NAND3 (N3763, N3761, N2999, N1226);
or OR3 (N3764, N3763, N505, N3628);
xor XOR2 (N3765, N3747, N3567);
xor XOR2 (N3766, N3764, N249);
nand NAND3 (N3767, N3765, N3553, N1426);
nor NOR2 (N3768, N3757, N521);
not NOT1 (N3769, N3745);
or OR3 (N3770, N3759, N2459, N675);
buf BUF1 (N3771, N3767);
or OR4 (N3772, N3749, N6, N2347, N2081);
not NOT1 (N3773, N3754);
nor NOR2 (N3774, N3772, N159);
and AND4 (N3775, N3762, N3000, N2309, N3375);
buf BUF1 (N3776, N3773);
and AND2 (N3777, N3753, N1360);
xor XOR2 (N3778, N3770, N925);
and AND4 (N3779, N3766, N2947, N230, N2645);
not NOT1 (N3780, N3760);
nand NAND4 (N3781, N3778, N2560, N1746, N3655);
nand NAND3 (N3782, N3777, N1111, N3366);
xor XOR2 (N3783, N3781, N53);
or OR4 (N3784, N3771, N2934, N3577, N129);
buf BUF1 (N3785, N3784);
or OR2 (N3786, N3779, N3444);
and AND4 (N3787, N3774, N3320, N1115, N2926);
xor XOR2 (N3788, N3776, N1092);
nor NOR4 (N3789, N3787, N1104, N2416, N2217);
nor NOR3 (N3790, N3782, N251, N3047);
nor NOR4 (N3791, N3775, N295, N1417, N3250);
or OR3 (N3792, N3783, N792, N202);
not NOT1 (N3793, N3786);
not NOT1 (N3794, N3789);
nor NOR2 (N3795, N3785, N3580);
not NOT1 (N3796, N3788);
and AND4 (N3797, N3796, N347, N2745, N529);
not NOT1 (N3798, N3791);
and AND4 (N3799, N3798, N2598, N2873, N2949);
and AND2 (N3800, N3795, N440);
xor XOR2 (N3801, N3793, N452);
nor NOR4 (N3802, N3769, N1281, N2949, N1380);
and AND2 (N3803, N3790, N1230);
not NOT1 (N3804, N3794);
buf BUF1 (N3805, N3804);
buf BUF1 (N3806, N3799);
not NOT1 (N3807, N3802);
xor XOR2 (N3808, N3768, N1168);
xor XOR2 (N3809, N3800, N3571);
and AND2 (N3810, N3809, N665);
nor NOR4 (N3811, N3807, N1093, N1574, N722);
and AND3 (N3812, N3803, N3578, N319);
nor NOR2 (N3813, N3810, N1211);
nand NAND2 (N3814, N3812, N400);
nand NAND3 (N3815, N3813, N3338, N1299);
nand NAND2 (N3816, N3806, N2681);
and AND3 (N3817, N3808, N2172, N899);
nor NOR2 (N3818, N3816, N913);
nand NAND3 (N3819, N3780, N2932, N2267);
buf BUF1 (N3820, N3814);
nand NAND2 (N3821, N3820, N1759);
and AND3 (N3822, N3815, N1943, N924);
or OR2 (N3823, N3805, N182);
not NOT1 (N3824, N3822);
not NOT1 (N3825, N3792);
buf BUF1 (N3826, N3801);
not NOT1 (N3827, N3821);
nand NAND4 (N3828, N3824, N2785, N3407, N2157);
not NOT1 (N3829, N3825);
buf BUF1 (N3830, N3817);
and AND2 (N3831, N3819, N3781);
nand NAND2 (N3832, N3826, N3718);
nor NOR2 (N3833, N3829, N2503);
buf BUF1 (N3834, N3827);
and AND3 (N3835, N3797, N2744, N3766);
and AND3 (N3836, N3823, N2021, N2037);
not NOT1 (N3837, N3833);
nor NOR4 (N3838, N3832, N173, N871, N1944);
or OR2 (N3839, N3834, N42);
xor XOR2 (N3840, N3818, N574);
or OR3 (N3841, N3840, N975, N2256);
xor XOR2 (N3842, N3830, N3116);
or OR4 (N3843, N3811, N2850, N3092, N1339);
nand NAND2 (N3844, N3828, N3151);
buf BUF1 (N3845, N3842);
nor NOR4 (N3846, N3838, N1293, N3427, N3556);
not NOT1 (N3847, N3831);
buf BUF1 (N3848, N3845);
not NOT1 (N3849, N3843);
nand NAND3 (N3850, N3839, N2957, N748);
not NOT1 (N3851, N3836);
nand NAND3 (N3852, N3844, N622, N2017);
or OR3 (N3853, N3849, N2008, N2707);
nor NOR4 (N3854, N3841, N3721, N3608, N968);
or OR3 (N3855, N3846, N3413, N264);
or OR4 (N3856, N3853, N1450, N2237, N3311);
nor NOR4 (N3857, N3855, N2203, N3554, N866);
xor XOR2 (N3858, N3857, N1091);
or OR4 (N3859, N3854, N2768, N3265, N3155);
and AND2 (N3860, N3859, N3459);
or OR4 (N3861, N3848, N3375, N957, N56);
nand NAND2 (N3862, N3850, N1297);
nand NAND3 (N3863, N3861, N664, N28);
and AND3 (N3864, N3835, N1674, N2736);
and AND3 (N3865, N3862, N2800, N554);
nor NOR4 (N3866, N3864, N2279, N370, N2167);
nor NOR3 (N3867, N3866, N2099, N1254);
nor NOR2 (N3868, N3858, N3257);
nor NOR4 (N3869, N3865, N1131, N1492, N368);
nand NAND2 (N3870, N3868, N1016);
nand NAND4 (N3871, N3867, N1264, N1195, N3337);
or OR2 (N3872, N3852, N3086);
nor NOR2 (N3873, N3860, N2690);
and AND2 (N3874, N3851, N771);
buf BUF1 (N3875, N3872);
buf BUF1 (N3876, N3873);
nand NAND2 (N3877, N3871, N2946);
not NOT1 (N3878, N3847);
nor NOR2 (N3879, N3870, N615);
nand NAND4 (N3880, N3877, N2702, N2912, N2918);
nand NAND3 (N3881, N3869, N2462, N1633);
buf BUF1 (N3882, N3881);
xor XOR2 (N3883, N3882, N1034);
not NOT1 (N3884, N3837);
and AND4 (N3885, N3874, N2301, N2819, N2183);
nor NOR2 (N3886, N3875, N3045);
nor NOR4 (N3887, N3863, N931, N3735, N2668);
nor NOR4 (N3888, N3885, N966, N1834, N688);
xor XOR2 (N3889, N3879, N1876);
not NOT1 (N3890, N3878);
not NOT1 (N3891, N3888);
nor NOR2 (N3892, N3889, N2776);
not NOT1 (N3893, N3883);
nand NAND3 (N3894, N3856, N2400, N2807);
or OR2 (N3895, N3886, N2943);
or OR4 (N3896, N3887, N1935, N2116, N1442);
or OR2 (N3897, N3890, N1140);
buf BUF1 (N3898, N3894);
or OR2 (N3899, N3896, N2485);
nand NAND4 (N3900, N3892, N300, N325, N221);
xor XOR2 (N3901, N3895, N2067);
not NOT1 (N3902, N3900);
not NOT1 (N3903, N3902);
nor NOR4 (N3904, N3893, N2603, N110, N1728);
xor XOR2 (N3905, N3898, N1513);
nand NAND2 (N3906, N3905, N1473);
nor NOR2 (N3907, N3901, N2486);
xor XOR2 (N3908, N3891, N991);
nor NOR2 (N3909, N3906, N2736);
xor XOR2 (N3910, N3907, N3282);
nand NAND2 (N3911, N3899, N3270);
nor NOR4 (N3912, N3903, N1801, N780, N2551);
nor NOR3 (N3913, N3904, N3473, N1120);
and AND3 (N3914, N3884, N2619, N43);
and AND4 (N3915, N3908, N1402, N1891, N1310);
nand NAND2 (N3916, N3880, N1434);
buf BUF1 (N3917, N3914);
xor XOR2 (N3918, N3912, N3492);
and AND3 (N3919, N3876, N2022, N1354);
buf BUF1 (N3920, N3917);
buf BUF1 (N3921, N3897);
nand NAND2 (N3922, N3911, N841);
and AND3 (N3923, N3913, N2521, N3559);
nand NAND4 (N3924, N3915, N2187, N2445, N1214);
not NOT1 (N3925, N3909);
xor XOR2 (N3926, N3925, N1209);
xor XOR2 (N3927, N3920, N3059);
buf BUF1 (N3928, N3916);
xor XOR2 (N3929, N3923, N511);
xor XOR2 (N3930, N3910, N3655);
nand NAND4 (N3931, N3930, N647, N1505, N1209);
xor XOR2 (N3932, N3928, N3620);
not NOT1 (N3933, N3921);
nand NAND3 (N3934, N3931, N160, N2821);
nand NAND4 (N3935, N3926, N2385, N1512, N2780);
or OR3 (N3936, N3924, N805, N3431);
buf BUF1 (N3937, N3929);
or OR2 (N3938, N3935, N189);
nand NAND2 (N3939, N3938, N216);
not NOT1 (N3940, N3937);
xor XOR2 (N3941, N3932, N2676);
nor NOR3 (N3942, N3936, N188, N3513);
and AND3 (N3943, N3940, N2033, N2733);
xor XOR2 (N3944, N3943, N139);
not NOT1 (N3945, N3934);
nor NOR3 (N3946, N3933, N1564, N674);
xor XOR2 (N3947, N3939, N2540);
or OR2 (N3948, N3919, N581);
or OR3 (N3949, N3942, N385, N705);
or OR3 (N3950, N3946, N573, N3604);
buf BUF1 (N3951, N3944);
nor NOR2 (N3952, N3922, N3510);
xor XOR2 (N3953, N3918, N2589);
nand NAND4 (N3954, N3947, N1579, N3297, N3046);
buf BUF1 (N3955, N3945);
not NOT1 (N3956, N3951);
or OR2 (N3957, N3954, N3668);
buf BUF1 (N3958, N3927);
buf BUF1 (N3959, N3948);
nor NOR3 (N3960, N3955, N1914, N3775);
nor NOR2 (N3961, N3956, N1831);
not NOT1 (N3962, N3941);
xor XOR2 (N3963, N3959, N2777);
and AND3 (N3964, N3960, N2504, N1078);
not NOT1 (N3965, N3957);
not NOT1 (N3966, N3963);
xor XOR2 (N3967, N3958, N1884);
nand NAND2 (N3968, N3965, N722);
not NOT1 (N3969, N3961);
xor XOR2 (N3970, N3969, N3381);
xor XOR2 (N3971, N3949, N2811);
xor XOR2 (N3972, N3967, N564);
and AND2 (N3973, N3971, N665);
nand NAND2 (N3974, N3970, N3837);
or OR2 (N3975, N3950, N148);
xor XOR2 (N3976, N3966, N3512);
nand NAND4 (N3977, N3974, N3540, N1844, N1352);
nand NAND2 (N3978, N3972, N2099);
not NOT1 (N3979, N3976);
xor XOR2 (N3980, N3952, N1590);
nand NAND3 (N3981, N3953, N3451, N2945);
xor XOR2 (N3982, N3980, N1777);
nor NOR4 (N3983, N3982, N2145, N1814, N526);
nand NAND2 (N3984, N3978, N2554);
and AND2 (N3985, N3975, N3440);
nor NOR4 (N3986, N3984, N3384, N1014, N2568);
or OR4 (N3987, N3981, N2697, N3698, N1663);
not NOT1 (N3988, N3977);
nand NAND3 (N3989, N3986, N2905, N2571);
or OR3 (N3990, N3968, N2, N1736);
and AND4 (N3991, N3987, N2615, N1448, N2179);
not NOT1 (N3992, N3989);
and AND4 (N3993, N3973, N2511, N2726, N1844);
not NOT1 (N3994, N3991);
xor XOR2 (N3995, N3964, N3407);
or OR2 (N3996, N3990, N3163);
xor XOR2 (N3997, N3962, N378);
and AND4 (N3998, N3988, N3919, N3957, N1988);
buf BUF1 (N3999, N3996);
nand NAND2 (N4000, N3992, N3611);
nand NAND2 (N4001, N3993, N1097);
nand NAND4 (N4002, N3985, N3803, N971, N1957);
not NOT1 (N4003, N4002);
nand NAND4 (N4004, N3983, N3458, N1379, N1724);
xor XOR2 (N4005, N4000, N1190);
xor XOR2 (N4006, N4001, N1472);
nand NAND3 (N4007, N3998, N776, N424);
buf BUF1 (N4008, N3999);
not NOT1 (N4009, N4003);
nor NOR3 (N4010, N4008, N708, N2442);
or OR4 (N4011, N4005, N190, N2786, N2315);
and AND2 (N4012, N3995, N2418);
endmodule