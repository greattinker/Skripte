// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N3202,N3213,N3211,N3190,N3216,N3199,N3208,N3212,N3197,N3218;

nor NOR2 (N19, N13, N4);
or OR3 (N20, N15, N11, N19);
nor NOR4 (N21, N12, N11, N1, N19);
xor XOR2 (N22, N4, N12);
nand NAND2 (N23, N9, N4);
xor XOR2 (N24, N23, N1);
nand NAND3 (N25, N17, N10, N1);
and AND4 (N26, N12, N2, N14, N19);
nor NOR2 (N27, N8, N4);
buf BUF1 (N28, N22);
nor NOR2 (N29, N10, N23);
or OR4 (N30, N10, N10, N1, N10);
nor NOR2 (N31, N2, N19);
nor NOR3 (N32, N25, N18, N15);
and AND2 (N33, N29, N6);
or OR4 (N34, N20, N11, N26, N33);
or OR3 (N35, N19, N18, N3);
nor NOR3 (N36, N7, N4, N4);
or OR4 (N37, N32, N5, N26, N34);
or OR2 (N38, N4, N17);
not NOT1 (N39, N21);
nand NAND2 (N40, N31, N1);
buf BUF1 (N41, N39);
nor NOR3 (N42, N27, N10, N10);
and AND4 (N43, N28, N37, N27, N24);
nand NAND4 (N44, N19, N42, N9, N37);
xor XOR2 (N45, N11, N44);
or OR2 (N46, N14, N12);
xor XOR2 (N47, N9, N28);
or OR3 (N48, N47, N16, N24);
or OR2 (N49, N41, N1);
buf BUF1 (N50, N49);
not NOT1 (N51, N45);
nand NAND2 (N52, N35, N17);
nand NAND2 (N53, N50, N49);
and AND2 (N54, N38, N19);
and AND2 (N55, N53, N41);
not NOT1 (N56, N52);
not NOT1 (N57, N30);
not NOT1 (N58, N46);
and AND3 (N59, N55, N47, N2);
nor NOR2 (N60, N36, N8);
not NOT1 (N61, N56);
nor NOR2 (N62, N40, N23);
and AND4 (N63, N59, N16, N55, N33);
xor XOR2 (N64, N58, N13);
buf BUF1 (N65, N51);
buf BUF1 (N66, N57);
not NOT1 (N67, N65);
buf BUF1 (N68, N67);
buf BUF1 (N69, N61);
nor NOR4 (N70, N48, N5, N59, N23);
buf BUF1 (N71, N69);
buf BUF1 (N72, N54);
not NOT1 (N73, N63);
and AND4 (N74, N70, N12, N71, N66);
and AND2 (N75, N38, N31);
nand NAND4 (N76, N19, N32, N44, N70);
nand NAND2 (N77, N64, N49);
and AND2 (N78, N43, N46);
nand NAND3 (N79, N60, N24, N50);
xor XOR2 (N80, N74, N53);
nor NOR4 (N81, N68, N16, N32, N46);
not NOT1 (N82, N78);
or OR4 (N83, N82, N17, N29, N27);
xor XOR2 (N84, N76, N19);
not NOT1 (N85, N83);
not NOT1 (N86, N84);
or OR4 (N87, N79, N10, N40, N62);
or OR2 (N88, N15, N9);
xor XOR2 (N89, N80, N31);
nand NAND4 (N90, N77, N86, N49, N75);
xor XOR2 (N91, N68, N48);
nor NOR3 (N92, N50, N83, N80);
and AND2 (N93, N73, N43);
buf BUF1 (N94, N89);
xor XOR2 (N95, N90, N41);
or OR4 (N96, N95, N40, N63, N48);
buf BUF1 (N97, N94);
nor NOR2 (N98, N85, N5);
and AND2 (N99, N72, N83);
nor NOR3 (N100, N96, N32, N26);
or OR2 (N101, N91, N74);
nand NAND3 (N102, N100, N50, N6);
and AND3 (N103, N98, N2, N95);
xor XOR2 (N104, N87, N75);
and AND3 (N105, N92, N89, N33);
xor XOR2 (N106, N104, N102);
nand NAND4 (N107, N44, N51, N92, N27);
buf BUF1 (N108, N106);
and AND4 (N109, N105, N17, N26, N74);
nand NAND2 (N110, N103, N35);
and AND4 (N111, N81, N110, N50, N103);
xor XOR2 (N112, N90, N60);
or OR4 (N113, N107, N94, N31, N68);
not NOT1 (N114, N99);
or OR4 (N115, N97, N60, N69, N10);
and AND4 (N116, N113, N35, N53, N82);
xor XOR2 (N117, N116, N77);
xor XOR2 (N118, N101, N9);
and AND2 (N119, N108, N45);
buf BUF1 (N120, N117);
and AND3 (N121, N119, N54, N107);
nor NOR4 (N122, N121, N16, N114, N118);
not NOT1 (N123, N79);
xor XOR2 (N124, N1, N28);
and AND2 (N125, N109, N36);
or OR2 (N126, N123, N24);
buf BUF1 (N127, N93);
or OR2 (N128, N124, N12);
nand NAND3 (N129, N125, N74, N71);
nor NOR3 (N130, N115, N41, N77);
buf BUF1 (N131, N126);
buf BUF1 (N132, N127);
or OR2 (N133, N112, N30);
not NOT1 (N134, N133);
not NOT1 (N135, N122);
or OR4 (N136, N130, N55, N29, N119);
xor XOR2 (N137, N129, N37);
nor NOR4 (N138, N136, N95, N124, N78);
xor XOR2 (N139, N135, N6);
not NOT1 (N140, N88);
nor NOR4 (N141, N132, N1, N28, N104);
not NOT1 (N142, N131);
and AND3 (N143, N141, N76, N135);
nor NOR3 (N144, N143, N33, N55);
not NOT1 (N145, N134);
or OR3 (N146, N142, N127, N64);
xor XOR2 (N147, N120, N10);
not NOT1 (N148, N139);
not NOT1 (N149, N146);
not NOT1 (N150, N144);
buf BUF1 (N151, N138);
xor XOR2 (N152, N147, N20);
nand NAND2 (N153, N140, N150);
or OR2 (N154, N3, N26);
and AND2 (N155, N149, N53);
nand NAND3 (N156, N151, N75, N121);
buf BUF1 (N157, N137);
not NOT1 (N158, N156);
and AND2 (N159, N154, N11);
nand NAND3 (N160, N128, N115, N86);
not NOT1 (N161, N158);
nor NOR4 (N162, N148, N84, N29, N160);
or OR4 (N163, N91, N154, N38, N159);
nor NOR2 (N164, N98, N154);
and AND3 (N165, N153, N117, N15);
not NOT1 (N166, N165);
and AND3 (N167, N161, N143, N42);
buf BUF1 (N168, N167);
and AND4 (N169, N168, N71, N38, N23);
nand NAND2 (N170, N169, N106);
buf BUF1 (N171, N157);
nand NAND4 (N172, N145, N24, N34, N25);
or OR2 (N173, N111, N80);
and AND3 (N174, N155, N115, N97);
nor NOR4 (N175, N173, N149, N105, N102);
nand NAND3 (N176, N174, N133, N145);
not NOT1 (N177, N176);
nor NOR2 (N178, N163, N85);
xor XOR2 (N179, N172, N127);
not NOT1 (N180, N178);
xor XOR2 (N181, N177, N156);
nor NOR4 (N182, N181, N161, N15, N151);
or OR4 (N183, N170, N93, N52, N114);
buf BUF1 (N184, N171);
buf BUF1 (N185, N162);
not NOT1 (N186, N184);
and AND2 (N187, N180, N67);
and AND2 (N188, N186, N96);
and AND2 (N189, N175, N150);
not NOT1 (N190, N183);
nor NOR2 (N191, N187, N30);
xor XOR2 (N192, N191, N163);
and AND4 (N193, N166, N165, N89, N53);
nand NAND2 (N194, N182, N190);
not NOT1 (N195, N7);
and AND2 (N196, N193, N186);
and AND2 (N197, N195, N42);
nand NAND3 (N198, N164, N90, N183);
or OR2 (N199, N188, N99);
nor NOR2 (N200, N197, N71);
and AND3 (N201, N152, N104, N183);
nor NOR3 (N202, N194, N151, N180);
and AND2 (N203, N192, N32);
and AND3 (N204, N199, N14, N40);
nor NOR4 (N205, N204, N99, N80, N104);
or OR4 (N206, N205, N75, N133, N9);
not NOT1 (N207, N198);
nand NAND3 (N208, N185, N3, N132);
or OR3 (N209, N200, N110, N166);
and AND3 (N210, N179, N133, N118);
and AND3 (N211, N189, N99, N51);
buf BUF1 (N212, N208);
buf BUF1 (N213, N212);
buf BUF1 (N214, N207);
xor XOR2 (N215, N213, N82);
nor NOR3 (N216, N196, N62, N79);
and AND2 (N217, N206, N63);
not NOT1 (N218, N216);
not NOT1 (N219, N217);
buf BUF1 (N220, N211);
nand NAND2 (N221, N202, N8);
xor XOR2 (N222, N203, N79);
nor NOR2 (N223, N209, N179);
nor NOR2 (N224, N220, N162);
xor XOR2 (N225, N222, N97);
buf BUF1 (N226, N201);
or OR3 (N227, N223, N140, N62);
nand NAND3 (N228, N225, N129, N190);
nand NAND2 (N229, N226, N173);
or OR4 (N230, N210, N190, N224, N142);
xor XOR2 (N231, N145, N128);
xor XOR2 (N232, N221, N19);
not NOT1 (N233, N219);
and AND2 (N234, N228, N77);
nor NOR3 (N235, N234, N56, N202);
xor XOR2 (N236, N233, N5);
not NOT1 (N237, N230);
xor XOR2 (N238, N215, N99);
or OR3 (N239, N235, N194, N66);
nand NAND4 (N240, N218, N52, N86, N38);
buf BUF1 (N241, N229);
nand NAND3 (N242, N241, N63, N72);
xor XOR2 (N243, N214, N200);
buf BUF1 (N244, N240);
buf BUF1 (N245, N236);
and AND3 (N246, N231, N27, N157);
nor NOR3 (N247, N227, N214, N21);
and AND4 (N248, N246, N244, N68, N121);
buf BUF1 (N249, N198);
xor XOR2 (N250, N238, N237);
xor XOR2 (N251, N228, N1);
nor NOR2 (N252, N249, N211);
not NOT1 (N253, N252);
xor XOR2 (N254, N245, N51);
and AND3 (N255, N253, N48, N204);
or OR2 (N256, N242, N252);
buf BUF1 (N257, N232);
xor XOR2 (N258, N248, N76);
or OR3 (N259, N250, N209, N211);
or OR3 (N260, N247, N83, N189);
not NOT1 (N261, N260);
xor XOR2 (N262, N254, N113);
nor NOR3 (N263, N239, N195, N111);
or OR4 (N264, N262, N183, N189, N113);
xor XOR2 (N265, N243, N208);
not NOT1 (N266, N257);
xor XOR2 (N267, N265, N168);
not NOT1 (N268, N267);
and AND2 (N269, N264, N228);
nor NOR2 (N270, N251, N92);
or OR3 (N271, N266, N18, N249);
not NOT1 (N272, N263);
nor NOR2 (N273, N261, N234);
nand NAND4 (N274, N259, N160, N127, N243);
buf BUF1 (N275, N274);
not NOT1 (N276, N256);
buf BUF1 (N277, N273);
nor NOR4 (N278, N277, N15, N105, N52);
and AND4 (N279, N278, N155, N235, N36);
or OR2 (N280, N276, N91);
buf BUF1 (N281, N280);
not NOT1 (N282, N269);
or OR3 (N283, N268, N24, N86);
and AND3 (N284, N271, N137, N95);
and AND4 (N285, N272, N36, N273, N272);
nor NOR3 (N286, N283, N185, N2);
not NOT1 (N287, N279);
xor XOR2 (N288, N285, N226);
xor XOR2 (N289, N284, N88);
xor XOR2 (N290, N281, N8);
xor XOR2 (N291, N287, N184);
and AND3 (N292, N286, N99, N97);
and AND4 (N293, N291, N147, N215, N69);
not NOT1 (N294, N270);
buf BUF1 (N295, N293);
or OR3 (N296, N288, N202, N118);
buf BUF1 (N297, N292);
nand NAND2 (N298, N295, N278);
not NOT1 (N299, N258);
nor NOR4 (N300, N294, N213, N295, N250);
and AND4 (N301, N255, N80, N210, N273);
not NOT1 (N302, N275);
nand NAND2 (N303, N297, N230);
xor XOR2 (N304, N282, N256);
nor NOR4 (N305, N299, N70, N157, N99);
nand NAND4 (N306, N298, N250, N193, N34);
buf BUF1 (N307, N289);
nor NOR3 (N308, N305, N67, N111);
buf BUF1 (N309, N301);
xor XOR2 (N310, N306, N253);
or OR4 (N311, N303, N21, N134, N96);
not NOT1 (N312, N290);
buf BUF1 (N313, N309);
nor NOR4 (N314, N311, N129, N36, N134);
nor NOR4 (N315, N313, N11, N31, N4);
xor XOR2 (N316, N296, N145);
nor NOR3 (N317, N310, N107, N219);
buf BUF1 (N318, N316);
nor NOR3 (N319, N307, N248, N49);
not NOT1 (N320, N302);
not NOT1 (N321, N317);
and AND4 (N322, N320, N122, N20, N17);
nand NAND3 (N323, N304, N159, N218);
not NOT1 (N324, N315);
nor NOR3 (N325, N323, N11, N87);
buf BUF1 (N326, N322);
xor XOR2 (N327, N321, N315);
or OR2 (N328, N319, N258);
nor NOR2 (N329, N328, N239);
xor XOR2 (N330, N324, N102);
nand NAND2 (N331, N329, N4);
and AND3 (N332, N318, N99, N303);
nor NOR3 (N333, N314, N166, N21);
nor NOR3 (N334, N330, N70, N270);
nand NAND3 (N335, N325, N233, N101);
xor XOR2 (N336, N300, N52);
nor NOR2 (N337, N336, N220);
and AND2 (N338, N333, N87);
and AND3 (N339, N335, N16, N182);
xor XOR2 (N340, N308, N286);
and AND2 (N341, N331, N172);
buf BUF1 (N342, N339);
nor NOR3 (N343, N327, N313, N261);
or OR4 (N344, N343, N341, N309, N144);
and AND2 (N345, N203, N57);
xor XOR2 (N346, N345, N167);
not NOT1 (N347, N346);
and AND4 (N348, N312, N155, N106, N142);
nand NAND2 (N349, N338, N232);
nor NOR3 (N350, N334, N62, N271);
and AND4 (N351, N326, N243, N310, N102);
or OR3 (N352, N344, N78, N198);
buf BUF1 (N353, N349);
buf BUF1 (N354, N353);
not NOT1 (N355, N348);
xor XOR2 (N356, N337, N19);
buf BUF1 (N357, N356);
not NOT1 (N358, N342);
not NOT1 (N359, N355);
buf BUF1 (N360, N332);
and AND3 (N361, N358, N251, N343);
nor NOR2 (N362, N357, N115);
nor NOR4 (N363, N362, N203, N238, N6);
buf BUF1 (N364, N352);
not NOT1 (N365, N354);
or OR3 (N366, N347, N344, N347);
not NOT1 (N367, N363);
not NOT1 (N368, N366);
and AND2 (N369, N351, N307);
not NOT1 (N370, N361);
buf BUF1 (N371, N368);
nor NOR4 (N372, N365, N184, N94, N371);
xor XOR2 (N373, N260, N202);
buf BUF1 (N374, N372);
and AND4 (N375, N364, N7, N288, N342);
nand NAND4 (N376, N350, N85, N50, N76);
xor XOR2 (N377, N367, N16);
buf BUF1 (N378, N373);
and AND4 (N379, N370, N364, N92, N44);
nand NAND2 (N380, N340, N223);
not NOT1 (N381, N375);
buf BUF1 (N382, N359);
xor XOR2 (N383, N381, N173);
or OR3 (N384, N380, N134, N31);
not NOT1 (N385, N369);
nor NOR3 (N386, N376, N296, N18);
buf BUF1 (N387, N385);
and AND3 (N388, N383, N246, N373);
not NOT1 (N389, N379);
or OR2 (N390, N387, N55);
xor XOR2 (N391, N390, N377);
not NOT1 (N392, N128);
not NOT1 (N393, N389);
or OR2 (N394, N386, N359);
xor XOR2 (N395, N391, N203);
buf BUF1 (N396, N393);
or OR3 (N397, N382, N385, N93);
or OR2 (N398, N395, N310);
nor NOR3 (N399, N378, N294, N310);
and AND3 (N400, N397, N284, N293);
nor NOR4 (N401, N398, N226, N227, N384);
and AND4 (N402, N277, N384, N52, N46);
xor XOR2 (N403, N392, N210);
not NOT1 (N404, N374);
nor NOR2 (N405, N388, N55);
not NOT1 (N406, N360);
nand NAND4 (N407, N399, N253, N154, N202);
nor NOR2 (N408, N404, N138);
nor NOR4 (N409, N406, N37, N358, N127);
not NOT1 (N410, N403);
buf BUF1 (N411, N402);
not NOT1 (N412, N401);
and AND2 (N413, N410, N45);
and AND3 (N414, N407, N412, N43);
nor NOR3 (N415, N213, N307, N170);
buf BUF1 (N416, N396);
and AND4 (N417, N415, N99, N199, N287);
not NOT1 (N418, N400);
nand NAND4 (N419, N405, N247, N7, N347);
or OR2 (N420, N418, N14);
xor XOR2 (N421, N414, N412);
not NOT1 (N422, N411);
nor NOR4 (N423, N394, N44, N29, N220);
and AND2 (N424, N413, N375);
buf BUF1 (N425, N420);
not NOT1 (N426, N425);
nor NOR3 (N427, N424, N292, N137);
or OR3 (N428, N427, N11, N54);
not NOT1 (N429, N409);
xor XOR2 (N430, N416, N161);
nand NAND3 (N431, N422, N70, N335);
nor NOR3 (N432, N419, N227, N253);
or OR3 (N433, N431, N229, N11);
nand NAND2 (N434, N423, N395);
not NOT1 (N435, N429);
not NOT1 (N436, N434);
nor NOR2 (N437, N417, N91);
and AND3 (N438, N436, N29, N24);
nor NOR2 (N439, N435, N73);
xor XOR2 (N440, N421, N245);
or OR4 (N441, N428, N202, N96, N128);
nand NAND2 (N442, N441, N152);
or OR2 (N443, N437, N320);
and AND2 (N444, N442, N132);
buf BUF1 (N445, N438);
xor XOR2 (N446, N439, N112);
and AND3 (N447, N426, N72, N215);
xor XOR2 (N448, N408, N152);
or OR2 (N449, N433, N332);
xor XOR2 (N450, N432, N169);
xor XOR2 (N451, N449, N99);
and AND2 (N452, N440, N181);
not NOT1 (N453, N444);
nand NAND3 (N454, N445, N132, N156);
xor XOR2 (N455, N451, N391);
or OR2 (N456, N453, N210);
nor NOR4 (N457, N456, N380, N290, N404);
not NOT1 (N458, N443);
not NOT1 (N459, N446);
xor XOR2 (N460, N448, N32);
xor XOR2 (N461, N447, N137);
nand NAND4 (N462, N450, N272, N208, N105);
nor NOR3 (N463, N430, N13, N3);
xor XOR2 (N464, N463, N11);
or OR4 (N465, N458, N342, N231, N278);
buf BUF1 (N466, N454);
buf BUF1 (N467, N452);
not NOT1 (N468, N461);
xor XOR2 (N469, N455, N183);
not NOT1 (N470, N464);
and AND4 (N471, N470, N36, N397, N448);
not NOT1 (N472, N460);
xor XOR2 (N473, N462, N467);
buf BUF1 (N474, N152);
or OR2 (N475, N471, N446);
nand NAND3 (N476, N459, N127, N118);
nor NOR4 (N477, N466, N322, N346, N339);
nor NOR4 (N478, N468, N170, N441, N188);
and AND2 (N479, N457, N417);
nor NOR4 (N480, N479, N371, N21, N359);
xor XOR2 (N481, N474, N468);
or OR2 (N482, N478, N451);
buf BUF1 (N483, N480);
or OR2 (N484, N475, N223);
nor NOR3 (N485, N472, N77, N69);
buf BUF1 (N486, N477);
not NOT1 (N487, N482);
and AND2 (N488, N486, N451);
nand NAND2 (N489, N488, N327);
or OR4 (N490, N487, N183, N160, N158);
and AND2 (N491, N490, N196);
or OR3 (N492, N469, N106, N246);
nand NAND4 (N493, N491, N374, N276, N278);
not NOT1 (N494, N485);
xor XOR2 (N495, N492, N290);
not NOT1 (N496, N465);
buf BUF1 (N497, N481);
nor NOR2 (N498, N473, N92);
buf BUF1 (N499, N498);
and AND3 (N500, N484, N74, N487);
xor XOR2 (N501, N495, N190);
not NOT1 (N502, N476);
nand NAND3 (N503, N489, N164, N105);
not NOT1 (N504, N497);
nand NAND2 (N505, N494, N223);
and AND3 (N506, N504, N278, N471);
and AND4 (N507, N499, N487, N284, N481);
nand NAND2 (N508, N506, N484);
not NOT1 (N509, N500);
nor NOR4 (N510, N496, N85, N233, N151);
nor NOR4 (N511, N502, N87, N499, N166);
nor NOR2 (N512, N510, N134);
nand NAND3 (N513, N512, N54, N300);
xor XOR2 (N514, N503, N258);
not NOT1 (N515, N507);
xor XOR2 (N516, N514, N455);
not NOT1 (N517, N516);
nor NOR3 (N518, N483, N385, N361);
and AND4 (N519, N518, N97, N82, N289);
nand NAND3 (N520, N501, N172, N467);
not NOT1 (N521, N509);
and AND3 (N522, N508, N178, N155);
or OR3 (N523, N505, N40, N484);
buf BUF1 (N524, N517);
nand NAND4 (N525, N515, N23, N305, N114);
and AND2 (N526, N493, N313);
nand NAND3 (N527, N524, N163, N35);
or OR2 (N528, N511, N318);
xor XOR2 (N529, N519, N452);
not NOT1 (N530, N526);
xor XOR2 (N531, N525, N64);
not NOT1 (N532, N521);
xor XOR2 (N533, N527, N169);
and AND2 (N534, N523, N170);
nor NOR2 (N535, N534, N149);
nand NAND4 (N536, N529, N414, N86, N482);
and AND2 (N537, N532, N352);
buf BUF1 (N538, N530);
not NOT1 (N539, N528);
or OR4 (N540, N539, N174, N538, N518);
or OR4 (N541, N248, N316, N409, N103);
not NOT1 (N542, N536);
buf BUF1 (N543, N542);
nand NAND4 (N544, N535, N367, N478, N94);
xor XOR2 (N545, N522, N208);
not NOT1 (N546, N533);
or OR4 (N547, N546, N171, N512, N524);
nor NOR3 (N548, N544, N474, N106);
xor XOR2 (N549, N547, N226);
buf BUF1 (N550, N543);
nor NOR4 (N551, N541, N103, N116, N479);
not NOT1 (N552, N540);
not NOT1 (N553, N552);
nor NOR3 (N554, N537, N16, N78);
and AND2 (N555, N550, N518);
nand NAND3 (N556, N531, N476, N174);
or OR4 (N557, N556, N189, N457, N410);
nor NOR3 (N558, N513, N334, N272);
and AND4 (N559, N548, N324, N115, N97);
not NOT1 (N560, N558);
buf BUF1 (N561, N557);
and AND4 (N562, N545, N172, N385, N49);
and AND3 (N563, N554, N292, N467);
nand NAND4 (N564, N520, N540, N534, N406);
buf BUF1 (N565, N555);
nand NAND4 (N566, N553, N324, N61, N317);
and AND2 (N567, N563, N532);
and AND3 (N568, N559, N564, N202);
xor XOR2 (N569, N243, N459);
nand NAND2 (N570, N561, N477);
nand NAND2 (N571, N551, N566);
buf BUF1 (N572, N388);
nand NAND2 (N573, N560, N382);
and AND2 (N574, N573, N107);
or OR3 (N575, N572, N559, N109);
not NOT1 (N576, N569);
nor NOR2 (N577, N571, N47);
nand NAND4 (N578, N568, N260, N161, N68);
and AND4 (N579, N570, N474, N195, N476);
or OR4 (N580, N577, N147, N190, N488);
nor NOR4 (N581, N549, N334, N529, N388);
nor NOR2 (N582, N562, N369);
or OR4 (N583, N580, N202, N132, N551);
nor NOR4 (N584, N575, N446, N94, N518);
not NOT1 (N585, N574);
nand NAND2 (N586, N581, N149);
or OR2 (N587, N582, N361);
nand NAND2 (N588, N576, N465);
xor XOR2 (N589, N588, N575);
or OR2 (N590, N586, N504);
or OR3 (N591, N583, N516, N424);
buf BUF1 (N592, N579);
xor XOR2 (N593, N591, N290);
and AND2 (N594, N578, N82);
nor NOR4 (N595, N594, N442, N208, N17);
nand NAND2 (N596, N567, N259);
xor XOR2 (N597, N585, N554);
nand NAND3 (N598, N592, N437, N60);
nand NAND3 (N599, N598, N598, N411);
buf BUF1 (N600, N584);
xor XOR2 (N601, N595, N190);
nor NOR4 (N602, N601, N99, N131, N315);
and AND4 (N603, N587, N292, N402, N473);
buf BUF1 (N604, N603);
not NOT1 (N605, N589);
xor XOR2 (N606, N565, N133);
buf BUF1 (N607, N606);
nand NAND4 (N608, N597, N595, N408, N257);
nand NAND2 (N609, N596, N443);
buf BUF1 (N610, N590);
nor NOR4 (N611, N600, N169, N596, N495);
nand NAND2 (N612, N593, N499);
or OR4 (N613, N612, N547, N349, N5);
nand NAND4 (N614, N610, N35, N507, N235);
nand NAND3 (N615, N604, N346, N4);
not NOT1 (N616, N614);
buf BUF1 (N617, N599);
and AND4 (N618, N617, N185, N211, N370);
and AND2 (N619, N613, N352);
buf BUF1 (N620, N605);
not NOT1 (N621, N620);
nand NAND4 (N622, N615, N370, N157, N554);
xor XOR2 (N623, N621, N328);
nor NOR4 (N624, N607, N314, N149, N578);
or OR4 (N625, N618, N372, N501, N94);
or OR2 (N626, N611, N605);
buf BUF1 (N627, N616);
buf BUF1 (N628, N623);
or OR3 (N629, N619, N381, N588);
and AND2 (N630, N629, N224);
not NOT1 (N631, N627);
nor NOR3 (N632, N631, N262, N273);
nand NAND3 (N633, N624, N381, N235);
buf BUF1 (N634, N622);
and AND4 (N635, N634, N345, N172, N174);
or OR2 (N636, N632, N428);
nand NAND2 (N637, N608, N78);
not NOT1 (N638, N636);
xor XOR2 (N639, N625, N350);
nor NOR3 (N640, N637, N153, N607);
or OR4 (N641, N602, N329, N265, N161);
buf BUF1 (N642, N641);
nand NAND2 (N643, N633, N542);
nor NOR3 (N644, N643, N376, N301);
buf BUF1 (N645, N626);
nor NOR3 (N646, N630, N326, N308);
xor XOR2 (N647, N635, N201);
buf BUF1 (N648, N642);
and AND4 (N649, N638, N127, N267, N488);
xor XOR2 (N650, N645, N90);
and AND2 (N651, N646, N647);
buf BUF1 (N652, N200);
xor XOR2 (N653, N650, N45);
nor NOR4 (N654, N644, N499, N560, N73);
not NOT1 (N655, N609);
xor XOR2 (N656, N640, N465);
nor NOR2 (N657, N655, N2);
nand NAND2 (N658, N652, N570);
nor NOR2 (N659, N656, N487);
not NOT1 (N660, N639);
nor NOR3 (N661, N649, N335, N520);
not NOT1 (N662, N628);
nor NOR2 (N663, N651, N30);
not NOT1 (N664, N654);
and AND2 (N665, N662, N275);
buf BUF1 (N666, N657);
or OR3 (N667, N661, N38, N284);
nor NOR2 (N668, N659, N119);
not NOT1 (N669, N666);
nand NAND2 (N670, N658, N309);
xor XOR2 (N671, N665, N320);
or OR3 (N672, N671, N522, N392);
not NOT1 (N673, N660);
or OR3 (N674, N672, N585, N453);
or OR4 (N675, N663, N617, N571, N655);
xor XOR2 (N676, N668, N237);
nor NOR3 (N677, N676, N3, N288);
not NOT1 (N678, N677);
and AND2 (N679, N667, N537);
nor NOR3 (N680, N653, N270, N231);
or OR3 (N681, N674, N458, N380);
not NOT1 (N682, N680);
nor NOR4 (N683, N681, N240, N445, N405);
nor NOR3 (N684, N673, N473, N172);
and AND3 (N685, N684, N180, N407);
nor NOR3 (N686, N669, N594, N66);
nand NAND2 (N687, N686, N469);
not NOT1 (N688, N648);
or OR2 (N689, N688, N557);
nand NAND3 (N690, N685, N139, N173);
buf BUF1 (N691, N679);
nand NAND3 (N692, N690, N139, N167);
and AND3 (N693, N670, N167, N557);
nand NAND3 (N694, N664, N194, N615);
buf BUF1 (N695, N693);
buf BUF1 (N696, N682);
nor NOR4 (N697, N678, N249, N540, N637);
and AND2 (N698, N675, N525);
nand NAND4 (N699, N692, N397, N151, N81);
nor NOR2 (N700, N699, N254);
buf BUF1 (N701, N696);
nand NAND2 (N702, N701, N90);
and AND2 (N703, N687, N366);
xor XOR2 (N704, N689, N168);
buf BUF1 (N705, N683);
or OR3 (N706, N703, N522, N588);
buf BUF1 (N707, N700);
xor XOR2 (N708, N706, N295);
xor XOR2 (N709, N698, N62);
and AND3 (N710, N691, N629, N182);
buf BUF1 (N711, N709);
nor NOR3 (N712, N702, N121, N301);
buf BUF1 (N713, N697);
or OR3 (N714, N707, N294, N349);
xor XOR2 (N715, N708, N553);
nand NAND3 (N716, N713, N476, N248);
or OR2 (N717, N694, N309);
not NOT1 (N718, N715);
nor NOR4 (N719, N717, N424, N687, N206);
nor NOR2 (N720, N705, N667);
or OR2 (N721, N718, N617);
buf BUF1 (N722, N714);
or OR3 (N723, N710, N602, N123);
buf BUF1 (N724, N719);
or OR2 (N725, N704, N212);
and AND3 (N726, N712, N436, N43);
xor XOR2 (N727, N721, N723);
not NOT1 (N728, N200);
nand NAND2 (N729, N726, N66);
nor NOR2 (N730, N722, N656);
not NOT1 (N731, N728);
or OR3 (N732, N725, N253, N512);
buf BUF1 (N733, N724);
xor XOR2 (N734, N720, N60);
buf BUF1 (N735, N732);
or OR4 (N736, N711, N609, N613, N128);
or OR4 (N737, N695, N566, N372, N663);
nor NOR4 (N738, N730, N657, N4, N76);
not NOT1 (N739, N734);
or OR3 (N740, N736, N432, N452);
not NOT1 (N741, N739);
buf BUF1 (N742, N738);
nand NAND3 (N743, N716, N351, N121);
and AND4 (N744, N735, N632, N589, N595);
or OR3 (N745, N729, N66, N491);
xor XOR2 (N746, N733, N270);
buf BUF1 (N747, N737);
nand NAND4 (N748, N741, N478, N635, N418);
nor NOR3 (N749, N746, N8, N495);
not NOT1 (N750, N727);
nor NOR2 (N751, N747, N368);
buf BUF1 (N752, N745);
buf BUF1 (N753, N740);
nand NAND2 (N754, N752, N71);
xor XOR2 (N755, N750, N5);
or OR3 (N756, N749, N167, N558);
nand NAND4 (N757, N751, N192, N297, N182);
nor NOR2 (N758, N743, N174);
xor XOR2 (N759, N754, N258);
nor NOR4 (N760, N756, N65, N743, N16);
nor NOR2 (N761, N759, N2);
not NOT1 (N762, N742);
nand NAND4 (N763, N755, N447, N377, N644);
nand NAND3 (N764, N753, N49, N658);
xor XOR2 (N765, N748, N740);
and AND3 (N766, N758, N622, N683);
or OR3 (N767, N764, N595, N692);
buf BUF1 (N768, N763);
not NOT1 (N769, N761);
or OR2 (N770, N765, N54);
buf BUF1 (N771, N766);
xor XOR2 (N772, N731, N147);
or OR2 (N773, N762, N250);
nand NAND4 (N774, N771, N473, N53, N566);
and AND3 (N775, N768, N50, N283);
xor XOR2 (N776, N773, N406);
nand NAND4 (N777, N775, N573, N591, N430);
nand NAND2 (N778, N767, N84);
not NOT1 (N779, N778);
nor NOR4 (N780, N757, N716, N462, N489);
nor NOR3 (N781, N770, N603, N159);
xor XOR2 (N782, N760, N113);
and AND3 (N783, N744, N625, N111);
nand NAND2 (N784, N782, N176);
buf BUF1 (N785, N769);
nor NOR2 (N786, N780, N502);
or OR2 (N787, N776, N303);
nand NAND3 (N788, N787, N750, N385);
not NOT1 (N789, N788);
and AND3 (N790, N789, N732, N407);
not NOT1 (N791, N779);
buf BUF1 (N792, N785);
or OR4 (N793, N781, N725, N650, N171);
or OR2 (N794, N792, N161);
nand NAND2 (N795, N790, N35);
or OR4 (N796, N794, N486, N791, N706);
not NOT1 (N797, N49);
not NOT1 (N798, N795);
or OR3 (N799, N796, N298, N523);
or OR3 (N800, N799, N215, N680);
nor NOR3 (N801, N772, N414, N764);
or OR2 (N802, N777, N144);
nand NAND3 (N803, N801, N20, N463);
nand NAND2 (N804, N784, N119);
or OR2 (N805, N798, N718);
xor XOR2 (N806, N800, N83);
or OR3 (N807, N806, N300, N269);
xor XOR2 (N808, N783, N348);
or OR4 (N809, N786, N337, N67, N261);
nor NOR4 (N810, N793, N635, N113, N582);
buf BUF1 (N811, N810);
not NOT1 (N812, N807);
not NOT1 (N813, N804);
nand NAND4 (N814, N803, N694, N318, N259);
nor NOR2 (N815, N802, N48);
not NOT1 (N816, N815);
nor NOR4 (N817, N809, N417, N126, N271);
nor NOR4 (N818, N817, N627, N178, N746);
not NOT1 (N819, N811);
nand NAND2 (N820, N774, N560);
nand NAND4 (N821, N812, N201, N286, N621);
nor NOR3 (N822, N821, N702, N616);
not NOT1 (N823, N814);
not NOT1 (N824, N820);
xor XOR2 (N825, N797, N689);
nand NAND2 (N826, N823, N19);
not NOT1 (N827, N808);
or OR2 (N828, N822, N566);
not NOT1 (N829, N816);
nor NOR2 (N830, N818, N2);
not NOT1 (N831, N805);
and AND3 (N832, N830, N548, N610);
and AND2 (N833, N829, N50);
buf BUF1 (N834, N831);
or OR4 (N835, N819, N351, N471, N131);
nor NOR4 (N836, N832, N440, N229, N427);
and AND2 (N837, N826, N95);
nor NOR4 (N838, N813, N256, N101, N561);
or OR4 (N839, N827, N101, N83, N55);
xor XOR2 (N840, N825, N443);
and AND3 (N841, N837, N290, N822);
not NOT1 (N842, N824);
nor NOR3 (N843, N836, N254, N441);
buf BUF1 (N844, N839);
nor NOR4 (N845, N841, N740, N365, N752);
xor XOR2 (N846, N834, N159);
or OR2 (N847, N845, N812);
not NOT1 (N848, N847);
buf BUF1 (N849, N840);
xor XOR2 (N850, N846, N58);
nand NAND3 (N851, N848, N133, N35);
nor NOR4 (N852, N844, N613, N403, N363);
nand NAND4 (N853, N828, N235, N627, N135);
and AND3 (N854, N842, N161, N531);
not NOT1 (N855, N852);
nand NAND4 (N856, N833, N399, N491, N544);
nand NAND2 (N857, N850, N829);
and AND3 (N858, N849, N176, N155);
and AND2 (N859, N855, N160);
or OR3 (N860, N843, N412, N33);
and AND3 (N861, N853, N210, N57);
and AND3 (N862, N857, N389, N742);
or OR2 (N863, N854, N810);
xor XOR2 (N864, N860, N648);
not NOT1 (N865, N856);
not NOT1 (N866, N865);
nand NAND2 (N867, N859, N443);
and AND2 (N868, N863, N867);
nor NOR4 (N869, N389, N696, N401, N80);
xor XOR2 (N870, N835, N654);
not NOT1 (N871, N858);
or OR3 (N872, N868, N836, N846);
or OR2 (N873, N838, N157);
buf BUF1 (N874, N864);
and AND3 (N875, N862, N689, N587);
nand NAND2 (N876, N873, N541);
xor XOR2 (N877, N866, N377);
nand NAND2 (N878, N869, N108);
not NOT1 (N879, N871);
not NOT1 (N880, N870);
buf BUF1 (N881, N872);
or OR2 (N882, N875, N801);
not NOT1 (N883, N876);
xor XOR2 (N884, N861, N147);
nand NAND2 (N885, N878, N860);
and AND4 (N886, N877, N28, N478, N141);
not NOT1 (N887, N881);
and AND3 (N888, N887, N743, N481);
or OR2 (N889, N888, N17);
not NOT1 (N890, N879);
nor NOR4 (N891, N883, N127, N812, N238);
xor XOR2 (N892, N885, N592);
or OR3 (N893, N890, N290, N514);
and AND3 (N894, N892, N429, N65);
not NOT1 (N895, N884);
xor XOR2 (N896, N889, N612);
and AND2 (N897, N886, N308);
nor NOR4 (N898, N882, N496, N883, N1);
and AND4 (N899, N893, N330, N492, N200);
and AND3 (N900, N851, N220, N173);
buf BUF1 (N901, N897);
not NOT1 (N902, N880);
nor NOR3 (N903, N902, N863, N331);
and AND4 (N904, N896, N6, N306, N740);
xor XOR2 (N905, N874, N473);
nand NAND2 (N906, N891, N742);
xor XOR2 (N907, N898, N461);
and AND3 (N908, N904, N105, N852);
nor NOR2 (N909, N908, N447);
and AND4 (N910, N906, N814, N731, N399);
or OR2 (N911, N905, N601);
not NOT1 (N912, N907);
not NOT1 (N913, N901);
buf BUF1 (N914, N900);
and AND4 (N915, N909, N427, N691, N813);
buf BUF1 (N916, N913);
nand NAND4 (N917, N914, N797, N777, N386);
xor XOR2 (N918, N911, N186);
and AND3 (N919, N899, N51, N205);
nor NOR2 (N920, N894, N915);
or OR4 (N921, N703, N811, N405, N132);
nor NOR2 (N922, N919, N812);
not NOT1 (N923, N922);
nor NOR3 (N924, N895, N170, N449);
nor NOR2 (N925, N918, N780);
xor XOR2 (N926, N917, N741);
xor XOR2 (N927, N921, N424);
xor XOR2 (N928, N923, N728);
not NOT1 (N929, N925);
not NOT1 (N930, N920);
buf BUF1 (N931, N924);
xor XOR2 (N932, N928, N253);
or OR4 (N933, N929, N144, N554, N181);
xor XOR2 (N934, N916, N429);
nor NOR4 (N935, N933, N873, N631, N359);
xor XOR2 (N936, N926, N429);
nor NOR4 (N937, N935, N138, N141, N649);
or OR3 (N938, N910, N846, N60);
nor NOR3 (N939, N927, N731, N92);
not NOT1 (N940, N937);
nand NAND2 (N941, N938, N885);
or OR4 (N942, N930, N855, N616, N822);
nor NOR2 (N943, N940, N86);
xor XOR2 (N944, N934, N696);
nand NAND2 (N945, N903, N776);
nor NOR3 (N946, N939, N453, N922);
or OR4 (N947, N936, N831, N680, N713);
nor NOR4 (N948, N947, N750, N278, N649);
buf BUF1 (N949, N944);
and AND4 (N950, N912, N591, N719, N63);
or OR3 (N951, N945, N287, N545);
xor XOR2 (N952, N942, N836);
not NOT1 (N953, N950);
xor XOR2 (N954, N948, N298);
xor XOR2 (N955, N941, N59);
not NOT1 (N956, N953);
buf BUF1 (N957, N943);
and AND3 (N958, N946, N460, N282);
or OR2 (N959, N932, N921);
and AND3 (N960, N956, N217, N17);
nand NAND2 (N961, N954, N110);
or OR2 (N962, N951, N279);
nand NAND3 (N963, N931, N175, N904);
nand NAND4 (N964, N957, N516, N140, N534);
nand NAND4 (N965, N964, N316, N698, N181);
xor XOR2 (N966, N949, N23);
nor NOR2 (N967, N961, N511);
or OR4 (N968, N960, N706, N92, N821);
nor NOR2 (N969, N955, N84);
buf BUF1 (N970, N966);
or OR2 (N971, N969, N924);
nor NOR4 (N972, N965, N966, N398, N184);
or OR3 (N973, N971, N958, N824);
or OR3 (N974, N263, N895, N677);
and AND2 (N975, N970, N742);
or OR2 (N976, N972, N149);
buf BUF1 (N977, N968);
nor NOR4 (N978, N973, N533, N551, N114);
not NOT1 (N979, N977);
xor XOR2 (N980, N974, N138);
and AND2 (N981, N975, N810);
nand NAND3 (N982, N979, N625, N610);
buf BUF1 (N983, N962);
nor NOR3 (N984, N976, N35, N520);
and AND4 (N985, N952, N561, N294, N367);
or OR4 (N986, N982, N625, N18, N859);
and AND2 (N987, N985, N533);
xor XOR2 (N988, N984, N368);
or OR4 (N989, N981, N300, N19, N987);
buf BUF1 (N990, N752);
or OR3 (N991, N980, N416, N189);
buf BUF1 (N992, N978);
not NOT1 (N993, N992);
buf BUF1 (N994, N988);
xor XOR2 (N995, N983, N228);
buf BUF1 (N996, N995);
nand NAND2 (N997, N994, N871);
or OR4 (N998, N989, N729, N707, N180);
or OR3 (N999, N996, N347, N535);
and AND4 (N1000, N997, N677, N90, N526);
and AND4 (N1001, N990, N67, N461, N104);
xor XOR2 (N1002, N1000, N8);
not NOT1 (N1003, N999);
not NOT1 (N1004, N959);
nor NOR4 (N1005, N963, N580, N879, N605);
or OR3 (N1006, N993, N78, N49);
xor XOR2 (N1007, N991, N932);
or OR4 (N1008, N1004, N612, N937, N986);
xor XOR2 (N1009, N253, N647);
or OR2 (N1010, N1003, N692);
not NOT1 (N1011, N1002);
xor XOR2 (N1012, N1011, N332);
nand NAND3 (N1013, N1006, N996, N17);
buf BUF1 (N1014, N1010);
nand NAND2 (N1015, N998, N241);
or OR4 (N1016, N1012, N370, N146, N870);
not NOT1 (N1017, N1015);
xor XOR2 (N1018, N1016, N804);
xor XOR2 (N1019, N1018, N15);
not NOT1 (N1020, N1009);
nor NOR4 (N1021, N1020, N721, N855, N111);
not NOT1 (N1022, N1008);
buf BUF1 (N1023, N1021);
not NOT1 (N1024, N1007);
nand NAND3 (N1025, N1017, N378, N355);
and AND2 (N1026, N1025, N320);
xor XOR2 (N1027, N1023, N583);
nor NOR3 (N1028, N967, N994, N611);
or OR4 (N1029, N1024, N937, N809, N421);
or OR4 (N1030, N1028, N979, N909, N447);
buf BUF1 (N1031, N1014);
buf BUF1 (N1032, N1001);
and AND3 (N1033, N1019, N429, N290);
nor NOR2 (N1034, N1005, N419);
or OR2 (N1035, N1033, N731);
and AND4 (N1036, N1035, N712, N334, N424);
or OR2 (N1037, N1027, N960);
nand NAND3 (N1038, N1036, N43, N760);
or OR2 (N1039, N1034, N867);
not NOT1 (N1040, N1038);
nor NOR2 (N1041, N1029, N905);
not NOT1 (N1042, N1013);
xor XOR2 (N1043, N1031, N264);
xor XOR2 (N1044, N1040, N651);
not NOT1 (N1045, N1032);
or OR2 (N1046, N1022, N106);
nand NAND2 (N1047, N1046, N332);
nor NOR4 (N1048, N1037, N154, N959, N628);
not NOT1 (N1049, N1042);
not NOT1 (N1050, N1030);
and AND3 (N1051, N1039, N313, N758);
and AND3 (N1052, N1050, N123, N174);
xor XOR2 (N1053, N1045, N6);
xor XOR2 (N1054, N1052, N138);
nor NOR4 (N1055, N1053, N127, N5, N565);
nor NOR2 (N1056, N1044, N992);
xor XOR2 (N1057, N1054, N278);
and AND4 (N1058, N1051, N122, N686, N1004);
buf BUF1 (N1059, N1058);
nor NOR4 (N1060, N1041, N929, N1054, N816);
not NOT1 (N1061, N1026);
buf BUF1 (N1062, N1048);
xor XOR2 (N1063, N1049, N149);
nand NAND4 (N1064, N1047, N338, N102, N935);
or OR2 (N1065, N1059, N603);
xor XOR2 (N1066, N1062, N489);
or OR2 (N1067, N1065, N770);
nor NOR2 (N1068, N1043, N419);
nand NAND2 (N1069, N1067, N768);
nor NOR3 (N1070, N1056, N141, N362);
and AND2 (N1071, N1064, N831);
or OR4 (N1072, N1070, N944, N42, N450);
buf BUF1 (N1073, N1061);
xor XOR2 (N1074, N1060, N585);
or OR4 (N1075, N1071, N956, N172, N817);
buf BUF1 (N1076, N1063);
buf BUF1 (N1077, N1074);
xor XOR2 (N1078, N1072, N888);
xor XOR2 (N1079, N1077, N575);
nor NOR2 (N1080, N1078, N647);
nand NAND4 (N1081, N1076, N23, N277, N580);
nor NOR2 (N1082, N1075, N194);
buf BUF1 (N1083, N1069);
nand NAND2 (N1084, N1079, N57);
and AND2 (N1085, N1057, N508);
not NOT1 (N1086, N1083);
not NOT1 (N1087, N1055);
nand NAND4 (N1088, N1084, N775, N513, N716);
not NOT1 (N1089, N1068);
nor NOR3 (N1090, N1089, N774, N256);
nand NAND4 (N1091, N1066, N261, N983, N418);
xor XOR2 (N1092, N1090, N826);
buf BUF1 (N1093, N1087);
xor XOR2 (N1094, N1085, N213);
buf BUF1 (N1095, N1092);
and AND4 (N1096, N1081, N303, N1074, N88);
nand NAND3 (N1097, N1093, N1046, N813);
and AND3 (N1098, N1086, N797, N947);
and AND4 (N1099, N1097, N292, N679, N516);
not NOT1 (N1100, N1099);
and AND4 (N1101, N1080, N699, N614, N298);
nand NAND2 (N1102, N1091, N669);
and AND2 (N1103, N1073, N568);
xor XOR2 (N1104, N1098, N29);
and AND4 (N1105, N1102, N403, N67, N486);
nor NOR3 (N1106, N1095, N224, N1050);
nor NOR2 (N1107, N1101, N192);
not NOT1 (N1108, N1106);
or OR3 (N1109, N1082, N214, N200);
and AND2 (N1110, N1104, N738);
nand NAND3 (N1111, N1108, N1066, N523);
or OR3 (N1112, N1109, N657, N783);
buf BUF1 (N1113, N1105);
xor XOR2 (N1114, N1100, N918);
and AND4 (N1115, N1088, N610, N186, N1066);
or OR4 (N1116, N1115, N151, N377, N925);
or OR3 (N1117, N1116, N914, N521);
and AND3 (N1118, N1111, N722, N907);
and AND2 (N1119, N1110, N956);
nand NAND3 (N1120, N1096, N150, N323);
not NOT1 (N1121, N1094);
buf BUF1 (N1122, N1113);
nand NAND2 (N1123, N1118, N915);
nor NOR2 (N1124, N1122, N844);
xor XOR2 (N1125, N1103, N1010);
not NOT1 (N1126, N1112);
nor NOR2 (N1127, N1123, N647);
or OR2 (N1128, N1124, N681);
not NOT1 (N1129, N1128);
xor XOR2 (N1130, N1117, N726);
nor NOR3 (N1131, N1120, N230, N558);
xor XOR2 (N1132, N1114, N275);
nor NOR3 (N1133, N1126, N9, N457);
nor NOR4 (N1134, N1133, N331, N686, N1071);
buf BUF1 (N1135, N1119);
buf BUF1 (N1136, N1135);
nand NAND3 (N1137, N1129, N974, N806);
not NOT1 (N1138, N1131);
nor NOR2 (N1139, N1127, N348);
xor XOR2 (N1140, N1130, N707);
and AND3 (N1141, N1121, N811, N398);
and AND2 (N1142, N1134, N538);
xor XOR2 (N1143, N1140, N40);
nand NAND3 (N1144, N1138, N142, N429);
nor NOR4 (N1145, N1125, N113, N1061, N381);
not NOT1 (N1146, N1141);
not NOT1 (N1147, N1136);
not NOT1 (N1148, N1132);
and AND3 (N1149, N1148, N1035, N260);
nand NAND4 (N1150, N1147, N752, N512, N232);
and AND3 (N1151, N1149, N113, N834);
nand NAND2 (N1152, N1137, N973);
nor NOR3 (N1153, N1143, N654, N137);
and AND4 (N1154, N1151, N888, N704, N830);
and AND3 (N1155, N1142, N809, N128);
xor XOR2 (N1156, N1139, N660);
or OR3 (N1157, N1144, N638, N663);
buf BUF1 (N1158, N1152);
nor NOR4 (N1159, N1158, N1095, N1122, N639);
or OR2 (N1160, N1145, N15);
or OR3 (N1161, N1160, N96, N611);
or OR4 (N1162, N1153, N523, N1154, N225);
nor NOR3 (N1163, N389, N73, N1005);
nor NOR2 (N1164, N1159, N137);
buf BUF1 (N1165, N1156);
and AND4 (N1166, N1155, N1031, N1050, N1134);
nor NOR4 (N1167, N1150, N1065, N880, N297);
nand NAND3 (N1168, N1167, N446, N198);
nor NOR3 (N1169, N1164, N135, N892);
and AND3 (N1170, N1168, N1156, N84);
xor XOR2 (N1171, N1146, N560);
or OR3 (N1172, N1165, N30, N404);
or OR3 (N1173, N1166, N22, N155);
nand NAND2 (N1174, N1169, N336);
and AND2 (N1175, N1170, N739);
xor XOR2 (N1176, N1163, N1033);
not NOT1 (N1177, N1162);
nand NAND4 (N1178, N1176, N626, N69, N1121);
and AND2 (N1179, N1174, N610);
nor NOR2 (N1180, N1107, N454);
nand NAND3 (N1181, N1180, N667, N317);
or OR4 (N1182, N1171, N296, N1129, N148);
not NOT1 (N1183, N1182);
buf BUF1 (N1184, N1161);
and AND3 (N1185, N1157, N1082, N191);
nand NAND4 (N1186, N1179, N801, N415, N311);
buf BUF1 (N1187, N1185);
or OR2 (N1188, N1184, N1183);
nor NOR4 (N1189, N438, N488, N1119, N639);
or OR4 (N1190, N1173, N612, N337, N369);
or OR2 (N1191, N1178, N379);
xor XOR2 (N1192, N1186, N126);
buf BUF1 (N1193, N1187);
buf BUF1 (N1194, N1172);
buf BUF1 (N1195, N1192);
nor NOR3 (N1196, N1194, N1170, N903);
nor NOR3 (N1197, N1188, N705, N320);
xor XOR2 (N1198, N1189, N186);
or OR4 (N1199, N1197, N1169, N636, N1134);
and AND3 (N1200, N1199, N2, N983);
buf BUF1 (N1201, N1177);
nand NAND4 (N1202, N1201, N116, N1073, N1161);
nor NOR2 (N1203, N1196, N986);
buf BUF1 (N1204, N1198);
xor XOR2 (N1205, N1195, N608);
not NOT1 (N1206, N1202);
nand NAND4 (N1207, N1175, N449, N1002, N610);
or OR3 (N1208, N1191, N1037, N1165);
nand NAND2 (N1209, N1190, N1142);
or OR4 (N1210, N1193, N690, N167, N228);
and AND3 (N1211, N1206, N439, N50);
xor XOR2 (N1212, N1200, N815);
or OR2 (N1213, N1207, N1206);
xor XOR2 (N1214, N1208, N1125);
buf BUF1 (N1215, N1211);
nand NAND2 (N1216, N1205, N74);
buf BUF1 (N1217, N1215);
nand NAND4 (N1218, N1210, N1141, N966, N1102);
nand NAND2 (N1219, N1217, N749);
xor XOR2 (N1220, N1214, N461);
xor XOR2 (N1221, N1218, N762);
nand NAND2 (N1222, N1204, N923);
buf BUF1 (N1223, N1212);
and AND2 (N1224, N1203, N693);
nor NOR2 (N1225, N1219, N1064);
nand NAND2 (N1226, N1213, N673);
nor NOR4 (N1227, N1216, N583, N1088, N1219);
buf BUF1 (N1228, N1227);
or OR2 (N1229, N1224, N174);
buf BUF1 (N1230, N1209);
and AND4 (N1231, N1225, N1034, N433, N825);
xor XOR2 (N1232, N1228, N667);
buf BUF1 (N1233, N1221);
xor XOR2 (N1234, N1230, N1053);
buf BUF1 (N1235, N1222);
nand NAND3 (N1236, N1231, N997, N5);
or OR3 (N1237, N1234, N785, N432);
not NOT1 (N1238, N1233);
or OR2 (N1239, N1235, N1057);
buf BUF1 (N1240, N1226);
nor NOR2 (N1241, N1236, N575);
or OR4 (N1242, N1229, N682, N989, N1136);
and AND4 (N1243, N1239, N113, N215, N920);
and AND4 (N1244, N1232, N555, N1154, N47);
buf BUF1 (N1245, N1241);
or OR4 (N1246, N1223, N628, N144, N380);
and AND2 (N1247, N1242, N581);
and AND3 (N1248, N1245, N1208, N43);
not NOT1 (N1249, N1240);
nor NOR3 (N1250, N1246, N480, N60);
or OR2 (N1251, N1181, N1247);
xor XOR2 (N1252, N1003, N944);
or OR3 (N1253, N1244, N1223, N255);
xor XOR2 (N1254, N1252, N634);
nand NAND3 (N1255, N1248, N250, N843);
and AND3 (N1256, N1254, N193, N464);
xor XOR2 (N1257, N1256, N1234);
and AND4 (N1258, N1253, N562, N959, N1257);
and AND3 (N1259, N186, N738, N1150);
nand NAND3 (N1260, N1258, N839, N24);
and AND3 (N1261, N1259, N66, N87);
nand NAND3 (N1262, N1260, N497, N847);
xor XOR2 (N1263, N1251, N958);
xor XOR2 (N1264, N1249, N253);
buf BUF1 (N1265, N1264);
buf BUF1 (N1266, N1237);
buf BUF1 (N1267, N1255);
buf BUF1 (N1268, N1261);
nor NOR3 (N1269, N1262, N805, N1079);
nor NOR2 (N1270, N1243, N1079);
not NOT1 (N1271, N1238);
xor XOR2 (N1272, N1263, N1024);
buf BUF1 (N1273, N1266);
and AND4 (N1274, N1267, N1167, N286, N978);
not NOT1 (N1275, N1220);
nor NOR4 (N1276, N1271, N294, N85, N299);
not NOT1 (N1277, N1269);
buf BUF1 (N1278, N1274);
and AND2 (N1279, N1277, N124);
xor XOR2 (N1280, N1265, N1014);
and AND4 (N1281, N1250, N459, N281, N283);
and AND2 (N1282, N1276, N1242);
xor XOR2 (N1283, N1282, N118);
nor NOR4 (N1284, N1279, N337, N1081, N870);
and AND3 (N1285, N1284, N1008, N1282);
and AND2 (N1286, N1278, N167);
not NOT1 (N1287, N1275);
xor XOR2 (N1288, N1268, N16);
xor XOR2 (N1289, N1273, N872);
not NOT1 (N1290, N1288);
xor XOR2 (N1291, N1287, N625);
not NOT1 (N1292, N1289);
buf BUF1 (N1293, N1286);
buf BUF1 (N1294, N1293);
and AND3 (N1295, N1285, N902, N979);
buf BUF1 (N1296, N1283);
nor NOR2 (N1297, N1295, N178);
buf BUF1 (N1298, N1297);
or OR3 (N1299, N1270, N743, N1298);
nor NOR3 (N1300, N908, N280, N433);
buf BUF1 (N1301, N1290);
xor XOR2 (N1302, N1291, N1166);
buf BUF1 (N1303, N1296);
nor NOR4 (N1304, N1294, N1161, N774, N60);
not NOT1 (N1305, N1292);
not NOT1 (N1306, N1301);
not NOT1 (N1307, N1305);
nor NOR4 (N1308, N1272, N453, N1242, N253);
nand NAND3 (N1309, N1302, N397, N582);
nand NAND2 (N1310, N1300, N1153);
not NOT1 (N1311, N1310);
xor XOR2 (N1312, N1307, N990);
or OR4 (N1313, N1306, N18, N846, N759);
not NOT1 (N1314, N1313);
not NOT1 (N1315, N1299);
not NOT1 (N1316, N1314);
nor NOR3 (N1317, N1315, N518, N1103);
not NOT1 (N1318, N1316);
nor NOR3 (N1319, N1312, N387, N530);
or OR3 (N1320, N1318, N756, N1094);
not NOT1 (N1321, N1320);
xor XOR2 (N1322, N1281, N318);
or OR3 (N1323, N1317, N20, N795);
or OR3 (N1324, N1319, N230, N1120);
buf BUF1 (N1325, N1308);
not NOT1 (N1326, N1311);
xor XOR2 (N1327, N1309, N548);
not NOT1 (N1328, N1326);
xor XOR2 (N1329, N1321, N1204);
not NOT1 (N1330, N1280);
nor NOR4 (N1331, N1324, N1285, N455, N650);
and AND4 (N1332, N1331, N7, N1031, N335);
not NOT1 (N1333, N1329);
not NOT1 (N1334, N1327);
nand NAND3 (N1335, N1325, N1219, N878);
nor NOR2 (N1336, N1332, N1247);
and AND3 (N1337, N1330, N1223, N890);
or OR3 (N1338, N1322, N166, N855);
not NOT1 (N1339, N1333);
nor NOR3 (N1340, N1303, N1334, N912);
or OR2 (N1341, N747, N988);
buf BUF1 (N1342, N1337);
nand NAND2 (N1343, N1336, N499);
not NOT1 (N1344, N1335);
buf BUF1 (N1345, N1342);
and AND4 (N1346, N1344, N882, N1275, N681);
nand NAND3 (N1347, N1339, N944, N764);
or OR3 (N1348, N1338, N1282, N1203);
or OR2 (N1349, N1304, N336);
xor XOR2 (N1350, N1345, N142);
nor NOR4 (N1351, N1350, N33, N858, N836);
not NOT1 (N1352, N1347);
nor NOR4 (N1353, N1340, N1044, N527, N588);
not NOT1 (N1354, N1353);
buf BUF1 (N1355, N1346);
nor NOR2 (N1356, N1343, N723);
not NOT1 (N1357, N1355);
nand NAND2 (N1358, N1341, N879);
buf BUF1 (N1359, N1348);
nand NAND4 (N1360, N1356, N1133, N517, N153);
xor XOR2 (N1361, N1328, N547);
buf BUF1 (N1362, N1357);
xor XOR2 (N1363, N1359, N112);
xor XOR2 (N1364, N1360, N301);
xor XOR2 (N1365, N1352, N141);
nand NAND2 (N1366, N1349, N1182);
not NOT1 (N1367, N1361);
or OR3 (N1368, N1367, N254, N1132);
not NOT1 (N1369, N1366);
xor XOR2 (N1370, N1323, N268);
nor NOR4 (N1371, N1369, N27, N243, N311);
nor NOR3 (N1372, N1351, N524, N872);
not NOT1 (N1373, N1358);
buf BUF1 (N1374, N1373);
not NOT1 (N1375, N1363);
xor XOR2 (N1376, N1354, N488);
nand NAND2 (N1377, N1371, N448);
nor NOR3 (N1378, N1374, N956, N1136);
buf BUF1 (N1379, N1375);
nor NOR4 (N1380, N1368, N244, N893, N755);
not NOT1 (N1381, N1379);
nor NOR3 (N1382, N1365, N727, N428);
xor XOR2 (N1383, N1381, N1250);
buf BUF1 (N1384, N1378);
or OR4 (N1385, N1362, N93, N15, N688);
buf BUF1 (N1386, N1364);
nand NAND4 (N1387, N1382, N632, N630, N529);
or OR4 (N1388, N1383, N1291, N196, N627);
nor NOR3 (N1389, N1388, N277, N1303);
xor XOR2 (N1390, N1389, N573);
nand NAND4 (N1391, N1386, N824, N401, N632);
nand NAND3 (N1392, N1376, N116, N1311);
nor NOR4 (N1393, N1384, N475, N976, N261);
nor NOR2 (N1394, N1392, N494);
nor NOR3 (N1395, N1370, N652, N950);
not NOT1 (N1396, N1380);
not NOT1 (N1397, N1393);
not NOT1 (N1398, N1390);
or OR2 (N1399, N1398, N793);
and AND3 (N1400, N1395, N1357, N535);
xor XOR2 (N1401, N1391, N1002);
nand NAND2 (N1402, N1397, N270);
nand NAND4 (N1403, N1402, N854, N203, N560);
buf BUF1 (N1404, N1385);
nor NOR4 (N1405, N1399, N882, N681, N642);
nand NAND3 (N1406, N1403, N859, N731);
nand NAND4 (N1407, N1404, N135, N7, N811);
nand NAND3 (N1408, N1372, N1072, N1162);
nand NAND4 (N1409, N1408, N1059, N1400, N509);
or OR3 (N1410, N930, N231, N510);
nor NOR2 (N1411, N1377, N706);
not NOT1 (N1412, N1410);
not NOT1 (N1413, N1409);
buf BUF1 (N1414, N1412);
not NOT1 (N1415, N1396);
buf BUF1 (N1416, N1415);
nor NOR3 (N1417, N1407, N1355, N1201);
nor NOR2 (N1418, N1414, N905);
nor NOR3 (N1419, N1406, N774, N399);
or OR4 (N1420, N1394, N115, N760, N316);
xor XOR2 (N1421, N1411, N864);
and AND3 (N1422, N1405, N162, N535);
nand NAND2 (N1423, N1422, N1341);
nand NAND4 (N1424, N1419, N838, N511, N354);
buf BUF1 (N1425, N1416);
not NOT1 (N1426, N1424);
not NOT1 (N1427, N1387);
and AND4 (N1428, N1418, N85, N1250, N382);
xor XOR2 (N1429, N1401, N1277);
buf BUF1 (N1430, N1423);
or OR3 (N1431, N1427, N1177, N821);
and AND4 (N1432, N1430, N1264, N454, N581);
nor NOR3 (N1433, N1428, N325, N1329);
xor XOR2 (N1434, N1417, N1059);
and AND2 (N1435, N1434, N1209);
nand NAND3 (N1436, N1435, N371, N1276);
and AND2 (N1437, N1429, N436);
not NOT1 (N1438, N1433);
nand NAND3 (N1439, N1425, N148, N126);
nand NAND2 (N1440, N1413, N978);
or OR4 (N1441, N1431, N1025, N1437, N473);
nor NOR3 (N1442, N1361, N271, N68);
or OR4 (N1443, N1426, N758, N1040, N586);
and AND3 (N1444, N1442, N860, N375);
or OR4 (N1445, N1443, N889, N105, N1186);
nor NOR4 (N1446, N1436, N434, N1408, N1288);
xor XOR2 (N1447, N1446, N777);
not NOT1 (N1448, N1420);
nand NAND4 (N1449, N1440, N336, N1203, N708);
nor NOR3 (N1450, N1421, N513, N574);
xor XOR2 (N1451, N1445, N794);
or OR4 (N1452, N1438, N1289, N563, N330);
or OR3 (N1453, N1441, N1214, N574);
not NOT1 (N1454, N1449);
nand NAND4 (N1455, N1439, N156, N177, N802);
buf BUF1 (N1456, N1454);
or OR4 (N1457, N1450, N575, N1106, N1336);
and AND4 (N1458, N1432, N577, N1187, N961);
nor NOR2 (N1459, N1451, N919);
and AND3 (N1460, N1453, N736, N1179);
not NOT1 (N1461, N1447);
buf BUF1 (N1462, N1452);
not NOT1 (N1463, N1461);
nand NAND3 (N1464, N1462, N162, N80);
and AND4 (N1465, N1460, N1069, N431, N859);
buf BUF1 (N1466, N1463);
not NOT1 (N1467, N1466);
xor XOR2 (N1468, N1467, N1061);
buf BUF1 (N1469, N1458);
and AND3 (N1470, N1469, N1284, N811);
nor NOR3 (N1471, N1456, N1256, N146);
not NOT1 (N1472, N1468);
nand NAND2 (N1473, N1464, N1392);
nor NOR3 (N1474, N1465, N704, N1189);
or OR2 (N1475, N1444, N302);
or OR4 (N1476, N1471, N468, N384, N47);
buf BUF1 (N1477, N1459);
xor XOR2 (N1478, N1470, N47);
nand NAND4 (N1479, N1477, N229, N385, N1326);
or OR3 (N1480, N1448, N1261, N1033);
not NOT1 (N1481, N1476);
not NOT1 (N1482, N1472);
xor XOR2 (N1483, N1478, N676);
xor XOR2 (N1484, N1482, N608);
buf BUF1 (N1485, N1483);
buf BUF1 (N1486, N1475);
nor NOR3 (N1487, N1481, N923, N1028);
not NOT1 (N1488, N1474);
nor NOR3 (N1489, N1479, N787, N1013);
not NOT1 (N1490, N1488);
not NOT1 (N1491, N1486);
nand NAND4 (N1492, N1480, N1187, N636, N781);
not NOT1 (N1493, N1489);
and AND4 (N1494, N1457, N78, N750, N246);
xor XOR2 (N1495, N1473, N222);
xor XOR2 (N1496, N1490, N979);
nand NAND4 (N1497, N1491, N1071, N997, N954);
nor NOR2 (N1498, N1487, N1336);
not NOT1 (N1499, N1485);
xor XOR2 (N1500, N1492, N555);
or OR3 (N1501, N1496, N1348, N615);
nor NOR4 (N1502, N1494, N1013, N1078, N513);
xor XOR2 (N1503, N1502, N1016);
xor XOR2 (N1504, N1455, N1308);
and AND3 (N1505, N1504, N516, N776);
nor NOR4 (N1506, N1500, N309, N190, N293);
not NOT1 (N1507, N1498);
buf BUF1 (N1508, N1499);
xor XOR2 (N1509, N1503, N830);
xor XOR2 (N1510, N1484, N968);
not NOT1 (N1511, N1510);
not NOT1 (N1512, N1511);
and AND4 (N1513, N1508, N769, N1198, N604);
nor NOR3 (N1514, N1497, N78, N415);
not NOT1 (N1515, N1501);
buf BUF1 (N1516, N1495);
not NOT1 (N1517, N1514);
buf BUF1 (N1518, N1493);
xor XOR2 (N1519, N1513, N1389);
nor NOR2 (N1520, N1509, N300);
and AND3 (N1521, N1519, N28, N1282);
xor XOR2 (N1522, N1515, N1362);
xor XOR2 (N1523, N1505, N791);
or OR3 (N1524, N1518, N1155, N785);
not NOT1 (N1525, N1522);
buf BUF1 (N1526, N1521);
nand NAND4 (N1527, N1507, N1193, N1431, N982);
not NOT1 (N1528, N1523);
nand NAND4 (N1529, N1506, N1045, N680, N34);
or OR3 (N1530, N1517, N431, N1191);
and AND4 (N1531, N1524, N163, N1092, N42);
not NOT1 (N1532, N1516);
nor NOR2 (N1533, N1525, N581);
or OR3 (N1534, N1520, N1298, N809);
or OR3 (N1535, N1532, N1045, N1403);
nor NOR4 (N1536, N1530, N1306, N813, N927);
not NOT1 (N1537, N1534);
xor XOR2 (N1538, N1531, N604);
not NOT1 (N1539, N1528);
xor XOR2 (N1540, N1536, N856);
buf BUF1 (N1541, N1527);
nor NOR2 (N1542, N1529, N623);
nand NAND3 (N1543, N1538, N514, N741);
nor NOR4 (N1544, N1512, N289, N1267, N58);
and AND4 (N1545, N1543, N777, N372, N21);
not NOT1 (N1546, N1535);
not NOT1 (N1547, N1546);
xor XOR2 (N1548, N1544, N304);
not NOT1 (N1549, N1547);
nor NOR2 (N1550, N1549, N1016);
nor NOR2 (N1551, N1526, N1040);
nand NAND2 (N1552, N1551, N460);
nor NOR3 (N1553, N1548, N134, N927);
nand NAND4 (N1554, N1533, N329, N1546, N1465);
nand NAND4 (N1555, N1554, N1072, N1317, N633);
xor XOR2 (N1556, N1542, N1257);
buf BUF1 (N1557, N1552);
or OR2 (N1558, N1553, N422);
or OR4 (N1559, N1537, N57, N1358, N1290);
xor XOR2 (N1560, N1558, N1186);
nand NAND4 (N1561, N1556, N1426, N751, N1086);
xor XOR2 (N1562, N1561, N18);
buf BUF1 (N1563, N1555);
nand NAND2 (N1564, N1550, N359);
or OR4 (N1565, N1560, N1447, N656, N879);
or OR3 (N1566, N1565, N1542, N622);
and AND4 (N1567, N1563, N179, N262, N433);
xor XOR2 (N1568, N1567, N1278);
nor NOR2 (N1569, N1545, N1176);
or OR2 (N1570, N1568, N79);
nand NAND3 (N1571, N1564, N932, N725);
or OR3 (N1572, N1540, N599, N1128);
or OR2 (N1573, N1571, N1399);
buf BUF1 (N1574, N1557);
and AND2 (N1575, N1562, N577);
and AND4 (N1576, N1566, N1396, N463, N1100);
nand NAND4 (N1577, N1559, N360, N929, N289);
and AND4 (N1578, N1577, N402, N1325, N1295);
nand NAND2 (N1579, N1541, N1187);
buf BUF1 (N1580, N1578);
and AND3 (N1581, N1539, N644, N789);
not NOT1 (N1582, N1574);
and AND3 (N1583, N1576, N558, N281);
or OR3 (N1584, N1570, N1452, N1275);
nand NAND2 (N1585, N1569, N207);
nor NOR2 (N1586, N1581, N77);
buf BUF1 (N1587, N1575);
buf BUF1 (N1588, N1583);
and AND3 (N1589, N1587, N506, N779);
buf BUF1 (N1590, N1589);
or OR3 (N1591, N1590, N628, N1343);
buf BUF1 (N1592, N1579);
nor NOR2 (N1593, N1572, N966);
nand NAND4 (N1594, N1592, N644, N1030, N1534);
not NOT1 (N1595, N1584);
or OR3 (N1596, N1588, N138, N747);
or OR3 (N1597, N1594, N1377, N240);
and AND2 (N1598, N1596, N747);
xor XOR2 (N1599, N1591, N1159);
not NOT1 (N1600, N1593);
and AND2 (N1601, N1600, N1156);
xor XOR2 (N1602, N1595, N912);
not NOT1 (N1603, N1573);
nor NOR3 (N1604, N1586, N240, N1380);
nand NAND2 (N1605, N1603, N555);
buf BUF1 (N1606, N1602);
nand NAND4 (N1607, N1582, N75, N1285, N567);
and AND2 (N1608, N1606, N1375);
or OR3 (N1609, N1580, N45, N1492);
buf BUF1 (N1610, N1604);
or OR3 (N1611, N1608, N730, N978);
buf BUF1 (N1612, N1609);
and AND3 (N1613, N1597, N1004, N1201);
nor NOR3 (N1614, N1599, N1483, N1247);
nor NOR3 (N1615, N1601, N735, N835);
not NOT1 (N1616, N1612);
xor XOR2 (N1617, N1611, N820);
or OR2 (N1618, N1610, N1095);
nand NAND4 (N1619, N1617, N140, N289, N778);
nand NAND4 (N1620, N1614, N406, N1576, N1371);
or OR3 (N1621, N1598, N1127, N318);
or OR3 (N1622, N1619, N1256, N1612);
buf BUF1 (N1623, N1585);
xor XOR2 (N1624, N1607, N1015);
xor XOR2 (N1625, N1605, N334);
nor NOR2 (N1626, N1622, N1617);
nor NOR4 (N1627, N1626, N1134, N319, N559);
nor NOR4 (N1628, N1625, N1450, N5, N233);
or OR4 (N1629, N1624, N560, N587, N1377);
nor NOR2 (N1630, N1629, N209);
nand NAND4 (N1631, N1615, N1565, N1376, N156);
buf BUF1 (N1632, N1623);
or OR2 (N1633, N1618, N1507);
and AND2 (N1634, N1631, N1113);
nor NOR4 (N1635, N1627, N804, N1628, N139);
nand NAND3 (N1636, N600, N127, N163);
and AND3 (N1637, N1633, N1407, N723);
xor XOR2 (N1638, N1637, N314);
nand NAND2 (N1639, N1613, N218);
or OR3 (N1640, N1638, N1126, N474);
or OR3 (N1641, N1635, N539, N433);
nand NAND2 (N1642, N1630, N1393);
xor XOR2 (N1643, N1642, N805);
xor XOR2 (N1644, N1643, N368);
buf BUF1 (N1645, N1641);
or OR3 (N1646, N1621, N122, N1330);
and AND2 (N1647, N1645, N156);
buf BUF1 (N1648, N1646);
or OR3 (N1649, N1648, N98, N1329);
xor XOR2 (N1650, N1640, N869);
buf BUF1 (N1651, N1634);
nand NAND3 (N1652, N1650, N821, N529);
xor XOR2 (N1653, N1616, N190);
nand NAND2 (N1654, N1649, N512);
nor NOR2 (N1655, N1653, N936);
nor NOR4 (N1656, N1652, N1621, N1646, N1327);
and AND2 (N1657, N1639, N630);
xor XOR2 (N1658, N1656, N811);
and AND2 (N1659, N1657, N1551);
not NOT1 (N1660, N1620);
buf BUF1 (N1661, N1654);
xor XOR2 (N1662, N1632, N1463);
xor XOR2 (N1663, N1644, N1279);
not NOT1 (N1664, N1651);
not NOT1 (N1665, N1636);
buf BUF1 (N1666, N1658);
or OR2 (N1667, N1660, N461);
not NOT1 (N1668, N1647);
xor XOR2 (N1669, N1659, N925);
not NOT1 (N1670, N1669);
not NOT1 (N1671, N1670);
nor NOR4 (N1672, N1662, N1448, N1451, N188);
and AND4 (N1673, N1664, N1544, N1234, N1423);
nand NAND4 (N1674, N1673, N917, N412, N237);
or OR2 (N1675, N1667, N1172);
xor XOR2 (N1676, N1655, N78);
and AND4 (N1677, N1661, N41, N159, N509);
not NOT1 (N1678, N1666);
xor XOR2 (N1679, N1674, N764);
and AND2 (N1680, N1678, N1325);
xor XOR2 (N1681, N1675, N132);
and AND4 (N1682, N1676, N1500, N1435, N1011);
nor NOR3 (N1683, N1680, N353, N1554);
or OR3 (N1684, N1681, N659, N1114);
xor XOR2 (N1685, N1677, N1638);
or OR4 (N1686, N1685, N1630, N1278, N929);
nor NOR4 (N1687, N1679, N107, N175, N317);
xor XOR2 (N1688, N1682, N1620);
nor NOR2 (N1689, N1687, N261);
xor XOR2 (N1690, N1686, N1028);
or OR4 (N1691, N1684, N1327, N1025, N1538);
buf BUF1 (N1692, N1665);
and AND3 (N1693, N1663, N282, N530);
xor XOR2 (N1694, N1671, N1616);
xor XOR2 (N1695, N1668, N1536);
or OR4 (N1696, N1683, N1305, N108, N985);
not NOT1 (N1697, N1690);
xor XOR2 (N1698, N1697, N340);
buf BUF1 (N1699, N1688);
nand NAND2 (N1700, N1692, N725);
nand NAND4 (N1701, N1693, N1179, N609, N302);
nand NAND3 (N1702, N1691, N1664, N500);
and AND2 (N1703, N1672, N334);
nor NOR4 (N1704, N1701, N1001, N1269, N1377);
or OR4 (N1705, N1694, N1152, N1649, N559);
and AND3 (N1706, N1702, N615, N739);
nor NOR3 (N1707, N1705, N1287, N764);
xor XOR2 (N1708, N1700, N1558);
buf BUF1 (N1709, N1704);
nor NOR3 (N1710, N1695, N1342, N32);
buf BUF1 (N1711, N1710);
and AND3 (N1712, N1698, N566, N904);
or OR3 (N1713, N1706, N1556, N1707);
nand NAND2 (N1714, N968, N1052);
or OR2 (N1715, N1711, N996);
buf BUF1 (N1716, N1708);
nor NOR4 (N1717, N1716, N576, N433, N1348);
nor NOR2 (N1718, N1712, N1624);
and AND4 (N1719, N1696, N1582, N104, N187);
and AND2 (N1720, N1709, N1076);
xor XOR2 (N1721, N1699, N1234);
buf BUF1 (N1722, N1703);
or OR2 (N1723, N1719, N877);
or OR3 (N1724, N1722, N388, N995);
nor NOR2 (N1725, N1714, N234);
nand NAND3 (N1726, N1725, N645, N1176);
not NOT1 (N1727, N1718);
buf BUF1 (N1728, N1715);
nor NOR2 (N1729, N1713, N17);
buf BUF1 (N1730, N1729);
and AND3 (N1731, N1726, N1226, N1297);
not NOT1 (N1732, N1689);
nand NAND3 (N1733, N1720, N1437, N926);
xor XOR2 (N1734, N1731, N1500);
xor XOR2 (N1735, N1721, N1709);
and AND4 (N1736, N1724, N1016, N1027, N1574);
not NOT1 (N1737, N1733);
nor NOR4 (N1738, N1732, N528, N497, N1197);
and AND4 (N1739, N1730, N1321, N1595, N304);
buf BUF1 (N1740, N1739);
or OR4 (N1741, N1738, N1560, N1130, N210);
or OR2 (N1742, N1727, N1391);
xor XOR2 (N1743, N1742, N1408);
xor XOR2 (N1744, N1741, N178);
nand NAND3 (N1745, N1734, N354, N829);
xor XOR2 (N1746, N1723, N1446);
not NOT1 (N1747, N1737);
buf BUF1 (N1748, N1747);
nand NAND2 (N1749, N1735, N459);
not NOT1 (N1750, N1717);
xor XOR2 (N1751, N1745, N295);
nor NOR2 (N1752, N1746, N1501);
and AND2 (N1753, N1728, N1376);
and AND4 (N1754, N1751, N1205, N674, N1679);
nand NAND3 (N1755, N1744, N536, N1742);
or OR3 (N1756, N1753, N283, N10);
xor XOR2 (N1757, N1740, N741);
or OR2 (N1758, N1754, N155);
buf BUF1 (N1759, N1757);
nor NOR2 (N1760, N1755, N1532);
or OR3 (N1761, N1758, N1247, N1324);
buf BUF1 (N1762, N1743);
and AND2 (N1763, N1760, N1663);
buf BUF1 (N1764, N1748);
buf BUF1 (N1765, N1762);
nor NOR3 (N1766, N1752, N881, N1143);
xor XOR2 (N1767, N1750, N1204);
buf BUF1 (N1768, N1761);
xor XOR2 (N1769, N1756, N1203);
nor NOR3 (N1770, N1764, N1005, N1469);
or OR2 (N1771, N1766, N1111);
buf BUF1 (N1772, N1767);
buf BUF1 (N1773, N1770);
or OR2 (N1774, N1765, N1109);
or OR4 (N1775, N1771, N1183, N23, N605);
nor NOR2 (N1776, N1769, N516);
or OR4 (N1777, N1759, N1753, N1287, N456);
nor NOR3 (N1778, N1772, N779, N1720);
xor XOR2 (N1779, N1768, N123);
or OR2 (N1780, N1736, N1713);
xor XOR2 (N1781, N1779, N24);
and AND2 (N1782, N1776, N968);
buf BUF1 (N1783, N1749);
buf BUF1 (N1784, N1783);
buf BUF1 (N1785, N1775);
or OR2 (N1786, N1763, N903);
not NOT1 (N1787, N1784);
nand NAND2 (N1788, N1774, N1097);
and AND2 (N1789, N1777, N943);
or OR4 (N1790, N1787, N673, N795, N1207);
not NOT1 (N1791, N1789);
or OR4 (N1792, N1790, N1039, N560, N811);
nand NAND3 (N1793, N1781, N1277, N341);
buf BUF1 (N1794, N1785);
buf BUF1 (N1795, N1780);
nor NOR2 (N1796, N1791, N869);
not NOT1 (N1797, N1792);
not NOT1 (N1798, N1795);
nand NAND4 (N1799, N1773, N761, N1636, N826);
xor XOR2 (N1800, N1782, N1103);
nor NOR3 (N1801, N1799, N1598, N1294);
xor XOR2 (N1802, N1796, N1487);
xor XOR2 (N1803, N1800, N1517);
nor NOR3 (N1804, N1802, N1027, N338);
and AND4 (N1805, N1794, N1772, N454, N1158);
or OR2 (N1806, N1805, N778);
nand NAND2 (N1807, N1788, N91);
xor XOR2 (N1808, N1778, N75);
buf BUF1 (N1809, N1808);
xor XOR2 (N1810, N1804, N1290);
nor NOR4 (N1811, N1798, N290, N1625, N1148);
not NOT1 (N1812, N1793);
nand NAND3 (N1813, N1801, N256, N1429);
buf BUF1 (N1814, N1806);
and AND3 (N1815, N1813, N1606, N306);
or OR4 (N1816, N1812, N79, N846, N381);
or OR3 (N1817, N1786, N559, N233);
or OR4 (N1818, N1816, N1301, N1207, N1162);
nor NOR3 (N1819, N1817, N1678, N573);
nand NAND2 (N1820, N1814, N482);
or OR2 (N1821, N1807, N869);
nor NOR2 (N1822, N1819, N804);
and AND4 (N1823, N1810, N817, N1320, N1678);
or OR4 (N1824, N1803, N977, N443, N298);
or OR4 (N1825, N1821, N1501, N30, N773);
nor NOR3 (N1826, N1815, N1452, N805);
not NOT1 (N1827, N1797);
and AND2 (N1828, N1826, N12);
nor NOR2 (N1829, N1818, N1100);
or OR4 (N1830, N1828, N1802, N663, N1667);
and AND2 (N1831, N1827, N361);
xor XOR2 (N1832, N1811, N1172);
xor XOR2 (N1833, N1831, N1344);
xor XOR2 (N1834, N1829, N499);
nand NAND2 (N1835, N1809, N219);
nand NAND3 (N1836, N1822, N685, N228);
nor NOR4 (N1837, N1825, N1110, N1157, N1116);
or OR4 (N1838, N1830, N90, N94, N1216);
or OR2 (N1839, N1836, N622);
xor XOR2 (N1840, N1837, N747);
xor XOR2 (N1841, N1833, N841);
nand NAND4 (N1842, N1823, N724, N1396, N1030);
and AND2 (N1843, N1842, N1658);
not NOT1 (N1844, N1838);
nor NOR4 (N1845, N1841, N1740, N471, N21);
xor XOR2 (N1846, N1845, N10);
or OR3 (N1847, N1840, N178, N1364);
nor NOR4 (N1848, N1835, N13, N924, N1730);
buf BUF1 (N1849, N1834);
xor XOR2 (N1850, N1839, N1125);
nor NOR4 (N1851, N1824, N608, N1550, N1657);
nand NAND3 (N1852, N1851, N780, N46);
or OR3 (N1853, N1846, N872, N731);
buf BUF1 (N1854, N1843);
nor NOR3 (N1855, N1853, N1390, N813);
and AND4 (N1856, N1832, N1470, N917, N484);
buf BUF1 (N1857, N1844);
xor XOR2 (N1858, N1856, N1512);
not NOT1 (N1859, N1820);
nand NAND4 (N1860, N1850, N718, N1622, N813);
nand NAND3 (N1861, N1858, N91, N1029);
xor XOR2 (N1862, N1854, N74);
xor XOR2 (N1863, N1860, N1204);
buf BUF1 (N1864, N1847);
not NOT1 (N1865, N1848);
nand NAND3 (N1866, N1852, N1790, N1674);
or OR3 (N1867, N1861, N428, N90);
or OR2 (N1868, N1864, N231);
buf BUF1 (N1869, N1849);
not NOT1 (N1870, N1866);
xor XOR2 (N1871, N1857, N1120);
or OR3 (N1872, N1863, N1526, N1800);
and AND4 (N1873, N1870, N1828, N1592, N377);
nor NOR3 (N1874, N1865, N420, N1019);
and AND4 (N1875, N1855, N120, N368, N609);
xor XOR2 (N1876, N1871, N1056);
not NOT1 (N1877, N1867);
buf BUF1 (N1878, N1875);
nor NOR3 (N1879, N1878, N1645, N653);
nand NAND4 (N1880, N1873, N290, N1364, N1151);
nor NOR4 (N1881, N1859, N5, N695, N1424);
or OR3 (N1882, N1879, N224, N1780);
nor NOR3 (N1883, N1877, N8, N756);
and AND2 (N1884, N1862, N1768);
or OR4 (N1885, N1876, N1218, N1587, N1082);
or OR4 (N1886, N1874, N1132, N1136, N1882);
or OR2 (N1887, N515, N660);
not NOT1 (N1888, N1880);
nor NOR3 (N1889, N1869, N793, N1319);
buf BUF1 (N1890, N1868);
nand NAND3 (N1891, N1885, N1170, N1099);
nor NOR3 (N1892, N1886, N1729, N369);
buf BUF1 (N1893, N1884);
and AND2 (N1894, N1892, N295);
buf BUF1 (N1895, N1887);
buf BUF1 (N1896, N1891);
not NOT1 (N1897, N1872);
buf BUF1 (N1898, N1889);
buf BUF1 (N1899, N1881);
or OR2 (N1900, N1883, N348);
and AND2 (N1901, N1894, N1102);
nand NAND4 (N1902, N1893, N1814, N164, N284);
and AND4 (N1903, N1902, N1305, N1538, N846);
and AND2 (N1904, N1890, N1550);
nand NAND3 (N1905, N1897, N103, N1391);
and AND3 (N1906, N1905, N1828, N760);
or OR4 (N1907, N1898, N1491, N788, N818);
nand NAND2 (N1908, N1907, N533);
buf BUF1 (N1909, N1896);
or OR4 (N1910, N1904, N1266, N1338, N327);
or OR2 (N1911, N1909, N124);
nor NOR3 (N1912, N1911, N1614, N1167);
xor XOR2 (N1913, N1895, N1705);
buf BUF1 (N1914, N1910);
xor XOR2 (N1915, N1906, N1550);
nor NOR2 (N1916, N1899, N765);
or OR3 (N1917, N1916, N319, N1649);
or OR2 (N1918, N1901, N1883);
buf BUF1 (N1919, N1913);
or OR2 (N1920, N1915, N1368);
buf BUF1 (N1921, N1900);
xor XOR2 (N1922, N1917, N128);
xor XOR2 (N1923, N1908, N658);
buf BUF1 (N1924, N1923);
not NOT1 (N1925, N1912);
not NOT1 (N1926, N1918);
not NOT1 (N1927, N1920);
nor NOR2 (N1928, N1924, N1431);
or OR3 (N1929, N1925, N1157, N914);
or OR3 (N1930, N1919, N664, N1745);
not NOT1 (N1931, N1903);
or OR2 (N1932, N1888, N531);
and AND4 (N1933, N1932, N1044, N772, N1673);
or OR4 (N1934, N1921, N1354, N1007, N264);
buf BUF1 (N1935, N1914);
and AND2 (N1936, N1935, N270);
nor NOR3 (N1937, N1931, N297, N586);
or OR4 (N1938, N1927, N86, N1766, N1269);
nor NOR3 (N1939, N1922, N1437, N325);
buf BUF1 (N1940, N1926);
buf BUF1 (N1941, N1937);
and AND3 (N1942, N1936, N912, N1507);
not NOT1 (N1943, N1940);
buf BUF1 (N1944, N1928);
xor XOR2 (N1945, N1941, N1509);
xor XOR2 (N1946, N1939, N932);
not NOT1 (N1947, N1929);
nand NAND4 (N1948, N1934, N875, N990, N878);
nand NAND3 (N1949, N1944, N282, N1817);
not NOT1 (N1950, N1943);
or OR3 (N1951, N1942, N1557, N1329);
xor XOR2 (N1952, N1949, N1119);
nand NAND4 (N1953, N1951, N1871, N1661, N1520);
xor XOR2 (N1954, N1933, N1124);
buf BUF1 (N1955, N1938);
nor NOR3 (N1956, N1954, N1832, N1021);
nand NAND4 (N1957, N1955, N858, N1329, N164);
xor XOR2 (N1958, N1957, N1700);
xor XOR2 (N1959, N1948, N983);
nand NAND3 (N1960, N1952, N838, N989);
buf BUF1 (N1961, N1947);
nor NOR2 (N1962, N1950, N1231);
xor XOR2 (N1963, N1946, N1407);
buf BUF1 (N1964, N1963);
or OR4 (N1965, N1964, N435, N1562, N138);
nor NOR2 (N1966, N1959, N1820);
nand NAND3 (N1967, N1965, N1873, N596);
or OR3 (N1968, N1966, N1785, N50);
nor NOR4 (N1969, N1967, N23, N1304, N81);
nand NAND3 (N1970, N1945, N1547, N1150);
buf BUF1 (N1971, N1962);
buf BUF1 (N1972, N1971);
not NOT1 (N1973, N1969);
and AND3 (N1974, N1958, N1586, N1676);
nand NAND4 (N1975, N1960, N1922, N431, N109);
xor XOR2 (N1976, N1975, N1249);
xor XOR2 (N1977, N1953, N1098);
and AND3 (N1978, N1976, N1200, N94);
xor XOR2 (N1979, N1961, N1107);
or OR2 (N1980, N1979, N171);
not NOT1 (N1981, N1930);
xor XOR2 (N1982, N1956, N1030);
nand NAND2 (N1983, N1977, N1568);
or OR4 (N1984, N1972, N727, N449, N363);
nand NAND3 (N1985, N1983, N594, N823);
and AND2 (N1986, N1973, N519);
nand NAND3 (N1987, N1974, N684, N64);
or OR2 (N1988, N1985, N1144);
xor XOR2 (N1989, N1978, N417);
and AND4 (N1990, N1986, N337, N1637, N146);
or OR3 (N1991, N1989, N1959, N139);
and AND3 (N1992, N1987, N1816, N527);
or OR4 (N1993, N1981, N981, N883, N844);
not NOT1 (N1994, N1993);
or OR3 (N1995, N1984, N1112, N1316);
buf BUF1 (N1996, N1970);
and AND4 (N1997, N1992, N1762, N1156, N1054);
xor XOR2 (N1998, N1968, N1868);
not NOT1 (N1999, N1990);
not NOT1 (N2000, N1997);
or OR3 (N2001, N1991, N1309, N1380);
nor NOR4 (N2002, N1988, N1383, N256, N1866);
buf BUF1 (N2003, N1996);
nand NAND3 (N2004, N1980, N94, N1642);
and AND3 (N2005, N1998, N1316, N700);
nor NOR3 (N2006, N2002, N726, N862);
buf BUF1 (N2007, N1995);
not NOT1 (N2008, N2001);
or OR3 (N2009, N2006, N503, N1938);
nor NOR3 (N2010, N2000, N931, N1027);
nor NOR2 (N2011, N2003, N1490);
xor XOR2 (N2012, N2007, N310);
xor XOR2 (N2013, N2012, N622);
nor NOR3 (N2014, N1999, N272, N344);
or OR3 (N2015, N2014, N469, N2000);
or OR4 (N2016, N2015, N1357, N649, N356);
nor NOR4 (N2017, N1982, N1319, N1685, N1615);
or OR4 (N2018, N2013, N560, N1093, N1176);
xor XOR2 (N2019, N2017, N1364);
and AND2 (N2020, N2019, N632);
nor NOR3 (N2021, N2004, N1931, N2005);
and AND2 (N2022, N1524, N537);
and AND4 (N2023, N2009, N172, N1639, N849);
nor NOR4 (N2024, N2016, N442, N341, N1949);
and AND2 (N2025, N1994, N998);
nand NAND2 (N2026, N2011, N675);
and AND3 (N2027, N2023, N1016, N382);
xor XOR2 (N2028, N2025, N1220);
buf BUF1 (N2029, N2022);
or OR2 (N2030, N2026, N1237);
and AND2 (N2031, N2010, N517);
nor NOR2 (N2032, N2024, N44);
xor XOR2 (N2033, N2018, N910);
xor XOR2 (N2034, N2029, N603);
not NOT1 (N2035, N2008);
and AND4 (N2036, N2030, N1424, N667, N208);
nand NAND2 (N2037, N2035, N1485);
not NOT1 (N2038, N2034);
xor XOR2 (N2039, N2033, N1698);
nor NOR2 (N2040, N2028, N976);
nand NAND2 (N2041, N2032, N615);
nand NAND3 (N2042, N2040, N1020, N769);
xor XOR2 (N2043, N2021, N1827);
nand NAND4 (N2044, N2041, N2016, N135, N1781);
buf BUF1 (N2045, N2037);
nor NOR4 (N2046, N2031, N1130, N1204, N325);
xor XOR2 (N2047, N2027, N790);
and AND3 (N2048, N2036, N456, N467);
buf BUF1 (N2049, N2047);
buf BUF1 (N2050, N2038);
not NOT1 (N2051, N2046);
nand NAND3 (N2052, N2050, N92, N1532);
nor NOR2 (N2053, N2020, N1463);
not NOT1 (N2054, N2051);
or OR4 (N2055, N2045, N987, N635, N1084);
xor XOR2 (N2056, N2053, N679);
not NOT1 (N2057, N2043);
not NOT1 (N2058, N2048);
xor XOR2 (N2059, N2039, N1029);
xor XOR2 (N2060, N2042, N1595);
buf BUF1 (N2061, N2059);
not NOT1 (N2062, N2060);
and AND2 (N2063, N2056, N1463);
not NOT1 (N2064, N2054);
buf BUF1 (N2065, N2052);
buf BUF1 (N2066, N2062);
or OR2 (N2067, N2063, N2032);
nor NOR3 (N2068, N2058, N872, N1774);
buf BUF1 (N2069, N2044);
or OR4 (N2070, N2068, N904, N498, N1462);
or OR2 (N2071, N2064, N1668);
buf BUF1 (N2072, N2070);
and AND4 (N2073, N2057, N7, N990, N1509);
buf BUF1 (N2074, N2055);
xor XOR2 (N2075, N2065, N406);
nor NOR3 (N2076, N2075, N1941, N1108);
xor XOR2 (N2077, N2061, N1369);
nor NOR2 (N2078, N2069, N1572);
buf BUF1 (N2079, N2072);
and AND3 (N2080, N2049, N884, N1033);
or OR4 (N2081, N2074, N1256, N712, N267);
nor NOR4 (N2082, N2079, N225, N342, N457);
buf BUF1 (N2083, N2077);
nand NAND2 (N2084, N2076, N1709);
and AND2 (N2085, N2081, N730);
nand NAND2 (N2086, N2085, N2028);
not NOT1 (N2087, N2083);
or OR2 (N2088, N2071, N2000);
not NOT1 (N2089, N2087);
buf BUF1 (N2090, N2088);
nor NOR4 (N2091, N2067, N1531, N1555, N267);
and AND2 (N2092, N2091, N929);
xor XOR2 (N2093, N2089, N704);
or OR4 (N2094, N2092, N1156, N1780, N485);
xor XOR2 (N2095, N2066, N520);
nor NOR3 (N2096, N2090, N765, N290);
buf BUF1 (N2097, N2082);
xor XOR2 (N2098, N2084, N504);
buf BUF1 (N2099, N2078);
nand NAND3 (N2100, N2080, N86, N1340);
buf BUF1 (N2101, N2099);
and AND3 (N2102, N2101, N2033, N1940);
nor NOR3 (N2103, N2073, N302, N1248);
buf BUF1 (N2104, N2103);
nand NAND3 (N2105, N2100, N1162, N662);
or OR4 (N2106, N2098, N587, N832, N408);
or OR4 (N2107, N2097, N1548, N151, N1822);
nor NOR3 (N2108, N2095, N2059, N978);
xor XOR2 (N2109, N2107, N2088);
nand NAND3 (N2110, N2105, N417, N639);
and AND2 (N2111, N2096, N518);
xor XOR2 (N2112, N2110, N187);
xor XOR2 (N2113, N2111, N76);
nor NOR2 (N2114, N2113, N1050);
not NOT1 (N2115, N2109);
not NOT1 (N2116, N2106);
nand NAND2 (N2117, N2102, N1470);
xor XOR2 (N2118, N2093, N924);
nor NOR2 (N2119, N2112, N161);
and AND3 (N2120, N2108, N1571, N1512);
not NOT1 (N2121, N2119);
xor XOR2 (N2122, N2114, N1652);
or OR2 (N2123, N2094, N1525);
not NOT1 (N2124, N2118);
buf BUF1 (N2125, N2123);
and AND2 (N2126, N2125, N1683);
or OR2 (N2127, N2086, N1606);
nor NOR4 (N2128, N2126, N1540, N1943, N332);
not NOT1 (N2129, N2117);
and AND3 (N2130, N2115, N1829, N636);
not NOT1 (N2131, N2122);
buf BUF1 (N2132, N2120);
not NOT1 (N2133, N2127);
nand NAND2 (N2134, N2104, N1438);
buf BUF1 (N2135, N2133);
not NOT1 (N2136, N2128);
xor XOR2 (N2137, N2131, N1030);
nor NOR4 (N2138, N2132, N1932, N1324, N1792);
buf BUF1 (N2139, N2134);
xor XOR2 (N2140, N2124, N516);
nand NAND4 (N2141, N2136, N2023, N1793, N1870);
or OR4 (N2142, N2141, N169, N535, N769);
and AND3 (N2143, N2116, N576, N924);
buf BUF1 (N2144, N2142);
not NOT1 (N2145, N2135);
or OR4 (N2146, N2129, N633, N1277, N1722);
or OR2 (N2147, N2140, N464);
or OR4 (N2148, N2137, N1508, N1684, N422);
and AND3 (N2149, N2148, N2075, N1769);
nand NAND4 (N2150, N2149, N233, N195, N1410);
buf BUF1 (N2151, N2150);
nor NOR3 (N2152, N2144, N481, N774);
xor XOR2 (N2153, N2130, N671);
or OR3 (N2154, N2121, N1602, N715);
xor XOR2 (N2155, N2147, N640);
buf BUF1 (N2156, N2155);
buf BUF1 (N2157, N2153);
buf BUF1 (N2158, N2151);
or OR2 (N2159, N2157, N470);
not NOT1 (N2160, N2156);
and AND3 (N2161, N2159, N587, N78);
buf BUF1 (N2162, N2145);
not NOT1 (N2163, N2158);
or OR3 (N2164, N2154, N1957, N27);
xor XOR2 (N2165, N2164, N1100);
or OR4 (N2166, N2139, N80, N1930, N203);
xor XOR2 (N2167, N2146, N792);
nor NOR3 (N2168, N2161, N2070, N1061);
xor XOR2 (N2169, N2165, N731);
nor NOR2 (N2170, N2168, N257);
nor NOR2 (N2171, N2143, N1202);
or OR4 (N2172, N2171, N1164, N73, N1520);
nor NOR3 (N2173, N2162, N147, N216);
nor NOR3 (N2174, N2152, N1498, N62);
buf BUF1 (N2175, N2166);
nor NOR4 (N2176, N2173, N382, N1230, N777);
and AND3 (N2177, N2138, N396, N42);
not NOT1 (N2178, N2163);
and AND2 (N2179, N2160, N1387);
buf BUF1 (N2180, N2179);
or OR2 (N2181, N2175, N860);
buf BUF1 (N2182, N2178);
not NOT1 (N2183, N2170);
xor XOR2 (N2184, N2182, N1756);
nand NAND2 (N2185, N2184, N1159);
buf BUF1 (N2186, N2169);
and AND3 (N2187, N2167, N1380, N1475);
and AND3 (N2188, N2177, N1451, N1326);
or OR3 (N2189, N2180, N290, N1505);
xor XOR2 (N2190, N2183, N559);
and AND3 (N2191, N2187, N1487, N283);
buf BUF1 (N2192, N2172);
xor XOR2 (N2193, N2176, N954);
xor XOR2 (N2194, N2188, N1013);
nand NAND4 (N2195, N2174, N1304, N1218, N230);
buf BUF1 (N2196, N2189);
buf BUF1 (N2197, N2196);
nand NAND2 (N2198, N2195, N2065);
xor XOR2 (N2199, N2181, N595);
and AND2 (N2200, N2197, N322);
not NOT1 (N2201, N2191);
nand NAND2 (N2202, N2185, N339);
buf BUF1 (N2203, N2200);
or OR3 (N2204, N2193, N1629, N935);
nor NOR3 (N2205, N2190, N1538, N76);
xor XOR2 (N2206, N2199, N537);
nor NOR2 (N2207, N2206, N1045);
or OR4 (N2208, N2186, N594, N1259, N1367);
xor XOR2 (N2209, N2204, N1622);
buf BUF1 (N2210, N2208);
or OR3 (N2211, N2202, N997, N719);
or OR4 (N2212, N2209, N308, N1801, N1782);
or OR2 (N2213, N2207, N261);
or OR3 (N2214, N2194, N671, N1756);
nand NAND2 (N2215, N2203, N2038);
nand NAND3 (N2216, N2215, N1792, N1776);
and AND3 (N2217, N2192, N1179, N285);
nor NOR2 (N2218, N2214, N450);
buf BUF1 (N2219, N2210);
or OR2 (N2220, N2205, N474);
xor XOR2 (N2221, N2212, N717);
not NOT1 (N2222, N2217);
nand NAND2 (N2223, N2219, N2116);
nand NAND2 (N2224, N2221, N364);
and AND2 (N2225, N2224, N449);
xor XOR2 (N2226, N2201, N1005);
and AND2 (N2227, N2222, N125);
and AND3 (N2228, N2213, N2144, N499);
xor XOR2 (N2229, N2227, N1054);
nand NAND4 (N2230, N2216, N936, N1268, N2122);
nand NAND3 (N2231, N2218, N1785, N646);
and AND2 (N2232, N2229, N872);
buf BUF1 (N2233, N2198);
nand NAND3 (N2234, N2226, N1850, N311);
nand NAND3 (N2235, N2228, N781, N2127);
not NOT1 (N2236, N2231);
xor XOR2 (N2237, N2235, N961);
nor NOR2 (N2238, N2233, N1516);
xor XOR2 (N2239, N2232, N920);
not NOT1 (N2240, N2239);
nor NOR3 (N2241, N2237, N843, N1171);
xor XOR2 (N2242, N2225, N2145);
nor NOR3 (N2243, N2241, N600, N1628);
xor XOR2 (N2244, N2223, N2046);
nor NOR2 (N2245, N2243, N476);
nand NAND3 (N2246, N2220, N1442, N1252);
buf BUF1 (N2247, N2234);
buf BUF1 (N2248, N2236);
buf BUF1 (N2249, N2211);
or OR4 (N2250, N2230, N46, N1571, N429);
xor XOR2 (N2251, N2245, N421);
buf BUF1 (N2252, N2240);
nor NOR3 (N2253, N2238, N471, N1952);
xor XOR2 (N2254, N2250, N1614);
buf BUF1 (N2255, N2254);
nor NOR3 (N2256, N2251, N827, N1150);
not NOT1 (N2257, N2253);
xor XOR2 (N2258, N2244, N383);
buf BUF1 (N2259, N2248);
nand NAND2 (N2260, N2258, N491);
or OR4 (N2261, N2249, N833, N907, N89);
nor NOR2 (N2262, N2256, N1876);
and AND3 (N2263, N2246, N575, N2053);
nand NAND2 (N2264, N2259, N1867);
and AND3 (N2265, N2263, N191, N971);
not NOT1 (N2266, N2257);
not NOT1 (N2267, N2264);
nor NOR4 (N2268, N2262, N928, N6, N1701);
not NOT1 (N2269, N2242);
nor NOR3 (N2270, N2269, N667, N1706);
not NOT1 (N2271, N2268);
and AND3 (N2272, N2270, N1113, N1931);
or OR2 (N2273, N2260, N398);
and AND3 (N2274, N2252, N1398, N386);
and AND4 (N2275, N2272, N1590, N2076, N968);
and AND3 (N2276, N2266, N842, N980);
nor NOR4 (N2277, N2265, N480, N1704, N868);
nand NAND2 (N2278, N2255, N764);
and AND3 (N2279, N2261, N1371, N1586);
nor NOR4 (N2280, N2273, N951, N1819, N524);
nand NAND3 (N2281, N2275, N485, N175);
buf BUF1 (N2282, N2279);
xor XOR2 (N2283, N2267, N1832);
nor NOR3 (N2284, N2280, N1544, N1502);
buf BUF1 (N2285, N2283);
xor XOR2 (N2286, N2281, N949);
xor XOR2 (N2287, N2274, N1111);
nand NAND2 (N2288, N2278, N58);
or OR4 (N2289, N2282, N2125, N837, N5);
buf BUF1 (N2290, N2289);
and AND4 (N2291, N2287, N1777, N1863, N105);
not NOT1 (N2292, N2247);
xor XOR2 (N2293, N2286, N1490);
xor XOR2 (N2294, N2293, N795);
nand NAND2 (N2295, N2288, N258);
nor NOR2 (N2296, N2292, N1013);
nand NAND2 (N2297, N2285, N784);
or OR2 (N2298, N2295, N531);
or OR3 (N2299, N2277, N888, N1089);
and AND4 (N2300, N2297, N2003, N1109, N1667);
nand NAND2 (N2301, N2294, N1322);
buf BUF1 (N2302, N2276);
and AND2 (N2303, N2291, N525);
not NOT1 (N2304, N2271);
not NOT1 (N2305, N2296);
or OR4 (N2306, N2302, N2255, N1455, N596);
or OR4 (N2307, N2290, N1765, N2068, N300);
not NOT1 (N2308, N2303);
nand NAND2 (N2309, N2301, N1698);
not NOT1 (N2310, N2305);
nand NAND3 (N2311, N2299, N471, N1276);
not NOT1 (N2312, N2304);
and AND2 (N2313, N2308, N588);
nand NAND4 (N2314, N2298, N1971, N97, N1113);
not NOT1 (N2315, N2284);
xor XOR2 (N2316, N2306, N1000);
xor XOR2 (N2317, N2316, N2086);
nand NAND4 (N2318, N2307, N1636, N883, N347);
nor NOR2 (N2319, N2311, N21);
nor NOR4 (N2320, N2309, N2221, N2008, N933);
buf BUF1 (N2321, N2315);
buf BUF1 (N2322, N2321);
not NOT1 (N2323, N2320);
nand NAND2 (N2324, N2310, N1284);
not NOT1 (N2325, N2319);
or OR4 (N2326, N2325, N29, N466, N991);
nor NOR2 (N2327, N2318, N99);
or OR3 (N2328, N2314, N2054, N1290);
xor XOR2 (N2329, N2324, N2304);
nand NAND3 (N2330, N2327, N2251, N2270);
not NOT1 (N2331, N2312);
not NOT1 (N2332, N2300);
buf BUF1 (N2333, N2331);
nand NAND3 (N2334, N2332, N1185, N490);
buf BUF1 (N2335, N2328);
not NOT1 (N2336, N2335);
and AND3 (N2337, N2333, N1092, N1895);
not NOT1 (N2338, N2322);
nand NAND3 (N2339, N2323, N2196, N1220);
not NOT1 (N2340, N2339);
nor NOR3 (N2341, N2330, N612, N831);
not NOT1 (N2342, N2329);
buf BUF1 (N2343, N2337);
buf BUF1 (N2344, N2338);
or OR3 (N2345, N2344, N1117, N95);
not NOT1 (N2346, N2341);
nor NOR4 (N2347, N2336, N1947, N837, N939);
not NOT1 (N2348, N2342);
and AND2 (N2349, N2340, N2182);
nor NOR4 (N2350, N2317, N818, N606, N1827);
nor NOR4 (N2351, N2346, N769, N2145, N794);
and AND3 (N2352, N2326, N1289, N1553);
nand NAND4 (N2353, N2334, N622, N1348, N59);
and AND2 (N2354, N2313, N2042);
buf BUF1 (N2355, N2348);
buf BUF1 (N2356, N2349);
xor XOR2 (N2357, N2351, N1002);
xor XOR2 (N2358, N2345, N365);
and AND2 (N2359, N2356, N1836);
nand NAND4 (N2360, N2359, N978, N1263, N2226);
not NOT1 (N2361, N2354);
and AND4 (N2362, N2358, N528, N773, N705);
buf BUF1 (N2363, N2352);
nand NAND3 (N2364, N2347, N2205, N89);
and AND3 (N2365, N2350, N1748, N1839);
not NOT1 (N2366, N2363);
nor NOR3 (N2367, N2353, N288, N782);
or OR2 (N2368, N2361, N897);
not NOT1 (N2369, N2355);
nand NAND4 (N2370, N2365, N2038, N2066, N2067);
xor XOR2 (N2371, N2368, N414);
nand NAND2 (N2372, N2366, N1573);
or OR2 (N2373, N2357, N2051);
not NOT1 (N2374, N2343);
nand NAND2 (N2375, N2367, N297);
xor XOR2 (N2376, N2362, N192);
not NOT1 (N2377, N2376);
nand NAND2 (N2378, N2360, N1193);
xor XOR2 (N2379, N2375, N604);
xor XOR2 (N2380, N2370, N83);
and AND2 (N2381, N2374, N2317);
buf BUF1 (N2382, N2378);
or OR3 (N2383, N2379, N1324, N1528);
nor NOR3 (N2384, N2369, N1658, N1121);
nor NOR2 (N2385, N2384, N2082);
and AND3 (N2386, N2381, N1094, N1339);
nor NOR3 (N2387, N2377, N367, N1328);
and AND3 (N2388, N2383, N1529, N844);
nor NOR2 (N2389, N2380, N1596);
nor NOR3 (N2390, N2385, N498, N3);
or OR4 (N2391, N2387, N1137, N261, N478);
nand NAND2 (N2392, N2388, N27);
xor XOR2 (N2393, N2391, N729);
buf BUF1 (N2394, N2389);
buf BUF1 (N2395, N2393);
or OR3 (N2396, N2371, N2071, N1143);
not NOT1 (N2397, N2372);
and AND2 (N2398, N2373, N1358);
nor NOR4 (N2399, N2398, N1709, N552, N1590);
nand NAND4 (N2400, N2364, N1121, N2086, N136);
or OR2 (N2401, N2396, N983);
or OR4 (N2402, N2397, N2075, N2264, N2241);
not NOT1 (N2403, N2395);
nand NAND2 (N2404, N2402, N2372);
not NOT1 (N2405, N2401);
nand NAND4 (N2406, N2382, N372, N2378, N1759);
xor XOR2 (N2407, N2406, N1039);
not NOT1 (N2408, N2405);
not NOT1 (N2409, N2400);
not NOT1 (N2410, N2386);
buf BUF1 (N2411, N2409);
buf BUF1 (N2412, N2407);
nor NOR4 (N2413, N2412, N785, N325, N411);
or OR4 (N2414, N2411, N1019, N1126, N621);
or OR4 (N2415, N2410, N1028, N2110, N1372);
not NOT1 (N2416, N2415);
and AND2 (N2417, N2399, N1321);
xor XOR2 (N2418, N2417, N1283);
and AND2 (N2419, N2413, N1235);
xor XOR2 (N2420, N2394, N268);
buf BUF1 (N2421, N2419);
xor XOR2 (N2422, N2414, N2217);
or OR4 (N2423, N2390, N954, N1983, N2343);
buf BUF1 (N2424, N2420);
nand NAND4 (N2425, N2392, N162, N1302, N2407);
nor NOR2 (N2426, N2408, N2389);
nor NOR4 (N2427, N2421, N663, N1192, N1765);
buf BUF1 (N2428, N2427);
and AND4 (N2429, N2422, N1775, N93, N880);
xor XOR2 (N2430, N2403, N2256);
nand NAND2 (N2431, N2429, N2100);
buf BUF1 (N2432, N2431);
or OR2 (N2433, N2418, N1076);
nor NOR2 (N2434, N2425, N2071);
nand NAND2 (N2435, N2430, N815);
and AND3 (N2436, N2426, N1501, N1383);
nor NOR3 (N2437, N2404, N1420, N1387);
nor NOR4 (N2438, N2428, N978, N806, N1005);
and AND2 (N2439, N2435, N420);
not NOT1 (N2440, N2436);
buf BUF1 (N2441, N2424);
buf BUF1 (N2442, N2416);
or OR2 (N2443, N2423, N629);
or OR3 (N2444, N2442, N1432, N901);
or OR3 (N2445, N2444, N509, N2401);
nand NAND3 (N2446, N2434, N492, N1053);
xor XOR2 (N2447, N2432, N700);
and AND3 (N2448, N2433, N2400, N2297);
not NOT1 (N2449, N2441);
nand NAND4 (N2450, N2438, N956, N1132, N892);
not NOT1 (N2451, N2450);
xor XOR2 (N2452, N2446, N517);
nor NOR4 (N2453, N2448, N892, N707, N228);
not NOT1 (N2454, N2440);
nor NOR3 (N2455, N2449, N1779, N2005);
and AND4 (N2456, N2452, N239, N908, N502);
xor XOR2 (N2457, N2453, N1327);
xor XOR2 (N2458, N2445, N1386);
xor XOR2 (N2459, N2447, N883);
xor XOR2 (N2460, N2458, N742);
and AND2 (N2461, N2455, N546);
buf BUF1 (N2462, N2439);
nor NOR3 (N2463, N2457, N1439, N804);
nor NOR4 (N2464, N2459, N504, N299, N524);
not NOT1 (N2465, N2461);
nand NAND3 (N2466, N2456, N182, N504);
or OR4 (N2467, N2462, N267, N841, N1867);
and AND3 (N2468, N2460, N2434, N1416);
nand NAND2 (N2469, N2451, N2463);
or OR2 (N2470, N2457, N2333);
and AND4 (N2471, N2469, N1237, N291, N2102);
nand NAND3 (N2472, N2454, N1473, N1212);
nand NAND4 (N2473, N2464, N197, N1586, N1860);
buf BUF1 (N2474, N2472);
nand NAND2 (N2475, N2443, N1626);
or OR3 (N2476, N2467, N2443, N640);
nor NOR2 (N2477, N2470, N859);
xor XOR2 (N2478, N2474, N1382);
buf BUF1 (N2479, N2437);
not NOT1 (N2480, N2473);
nand NAND2 (N2481, N2478, N853);
buf BUF1 (N2482, N2477);
nand NAND4 (N2483, N2475, N1816, N182, N246);
buf BUF1 (N2484, N2479);
and AND4 (N2485, N2481, N1892, N201, N1669);
not NOT1 (N2486, N2468);
or OR3 (N2487, N2465, N2399, N1155);
and AND4 (N2488, N2487, N1027, N1737, N1142);
not NOT1 (N2489, N2486);
xor XOR2 (N2490, N2485, N165);
and AND2 (N2491, N2484, N434);
xor XOR2 (N2492, N2490, N2221);
nor NOR2 (N2493, N2476, N1267);
and AND2 (N2494, N2493, N1762);
nand NAND2 (N2495, N2482, N1194);
or OR4 (N2496, N2466, N1709, N16, N1085);
and AND2 (N2497, N2496, N265);
nor NOR3 (N2498, N2491, N322, N1461);
not NOT1 (N2499, N2480);
or OR4 (N2500, N2489, N1819, N573, N2230);
xor XOR2 (N2501, N2499, N139);
buf BUF1 (N2502, N2494);
nor NOR4 (N2503, N2497, N1779, N1218, N2327);
nand NAND4 (N2504, N2503, N1057, N991, N1360);
nand NAND3 (N2505, N2488, N747, N2137);
nand NAND3 (N2506, N2504, N1142, N2444);
nor NOR3 (N2507, N2505, N2116, N316);
or OR2 (N2508, N2501, N1600);
nor NOR3 (N2509, N2508, N315, N86);
or OR2 (N2510, N2500, N2225);
nand NAND4 (N2511, N2506, N2263, N1215, N1613);
nand NAND3 (N2512, N2492, N1742, N916);
not NOT1 (N2513, N2510);
nor NOR4 (N2514, N2509, N850, N1364, N454);
nor NOR3 (N2515, N2471, N159, N1103);
not NOT1 (N2516, N2495);
not NOT1 (N2517, N2516);
not NOT1 (N2518, N2514);
nand NAND4 (N2519, N2511, N2109, N2109, N55);
xor XOR2 (N2520, N2515, N934);
buf BUF1 (N2521, N2513);
xor XOR2 (N2522, N2517, N1334);
or OR2 (N2523, N2518, N250);
or OR4 (N2524, N2512, N360, N1842, N751);
and AND2 (N2525, N2483, N733);
nand NAND2 (N2526, N2522, N2308);
nor NOR3 (N2527, N2519, N2390, N1047);
nand NAND4 (N2528, N2525, N235, N1131, N2392);
nor NOR2 (N2529, N2521, N557);
buf BUF1 (N2530, N2507);
xor XOR2 (N2531, N2502, N1098);
and AND2 (N2532, N2524, N1096);
and AND3 (N2533, N2526, N669, N463);
not NOT1 (N2534, N2530);
or OR3 (N2535, N2498, N375, N1981);
not NOT1 (N2536, N2531);
and AND3 (N2537, N2527, N2134, N1383);
nand NAND4 (N2538, N2535, N1955, N166, N434);
and AND3 (N2539, N2534, N1989, N1527);
nand NAND2 (N2540, N2536, N1963);
or OR3 (N2541, N2523, N918, N2359);
or OR2 (N2542, N2541, N1530);
xor XOR2 (N2543, N2520, N1714);
nand NAND2 (N2544, N2540, N1882);
or OR4 (N2545, N2537, N2056, N846, N1355);
not NOT1 (N2546, N2528);
or OR4 (N2547, N2545, N543, N2027, N988);
and AND4 (N2548, N2538, N854, N2460, N1351);
nor NOR3 (N2549, N2547, N353, N1275);
or OR3 (N2550, N2532, N905, N2444);
nor NOR2 (N2551, N2550, N1290);
nor NOR4 (N2552, N2544, N1756, N295, N693);
buf BUF1 (N2553, N2543);
nor NOR2 (N2554, N2552, N808);
nor NOR2 (N2555, N2553, N650);
nand NAND3 (N2556, N2554, N2367, N835);
xor XOR2 (N2557, N2533, N1759);
nand NAND2 (N2558, N2542, N1664);
xor XOR2 (N2559, N2557, N985);
buf BUF1 (N2560, N2539);
nor NOR3 (N2561, N2548, N2355, N98);
nand NAND4 (N2562, N2560, N1828, N480, N341);
nand NAND2 (N2563, N2546, N2305);
or OR3 (N2564, N2562, N500, N52);
xor XOR2 (N2565, N2556, N2148);
not NOT1 (N2566, N2551);
nor NOR3 (N2567, N2529, N495, N831);
buf BUF1 (N2568, N2558);
or OR3 (N2569, N2566, N623, N2421);
and AND4 (N2570, N2568, N743, N1076, N2264);
xor XOR2 (N2571, N2565, N1129);
not NOT1 (N2572, N2567);
nand NAND2 (N2573, N2572, N1510);
xor XOR2 (N2574, N2559, N1431);
nor NOR2 (N2575, N2570, N966);
buf BUF1 (N2576, N2549);
not NOT1 (N2577, N2564);
not NOT1 (N2578, N2577);
not NOT1 (N2579, N2561);
xor XOR2 (N2580, N2555, N1938);
and AND3 (N2581, N2576, N2390, N589);
and AND3 (N2582, N2569, N591, N180);
not NOT1 (N2583, N2563);
and AND4 (N2584, N2579, N659, N617, N421);
and AND4 (N2585, N2580, N54, N93, N1710);
buf BUF1 (N2586, N2584);
or OR4 (N2587, N2578, N2214, N556, N355);
xor XOR2 (N2588, N2581, N1172);
or OR3 (N2589, N2586, N534, N1461);
and AND3 (N2590, N2573, N564, N530);
nor NOR3 (N2591, N2575, N720, N737);
xor XOR2 (N2592, N2571, N704);
and AND3 (N2593, N2588, N221, N1359);
and AND3 (N2594, N2592, N2198, N1809);
not NOT1 (N2595, N2583);
and AND3 (N2596, N2595, N1232, N1414);
buf BUF1 (N2597, N2574);
and AND2 (N2598, N2590, N525);
not NOT1 (N2599, N2589);
nand NAND4 (N2600, N2596, N867, N1790, N2567);
not NOT1 (N2601, N2582);
buf BUF1 (N2602, N2594);
buf BUF1 (N2603, N2587);
xor XOR2 (N2604, N2603, N952);
not NOT1 (N2605, N2598);
nor NOR3 (N2606, N2585, N1228, N272);
or OR2 (N2607, N2606, N298);
and AND3 (N2608, N2597, N1082, N2017);
and AND3 (N2609, N2605, N1366, N2339);
nand NAND3 (N2610, N2601, N491, N2511);
nor NOR2 (N2611, N2600, N2340);
and AND2 (N2612, N2604, N75);
nor NOR3 (N2613, N2609, N814, N1012);
or OR3 (N2614, N2591, N1203, N2552);
xor XOR2 (N2615, N2607, N1319);
nand NAND3 (N2616, N2599, N926, N261);
nor NOR4 (N2617, N2602, N148, N1811, N168);
not NOT1 (N2618, N2610);
buf BUF1 (N2619, N2616);
and AND3 (N2620, N2593, N319, N1607);
or OR2 (N2621, N2612, N495);
or OR3 (N2622, N2615, N960, N1227);
or OR2 (N2623, N2613, N323);
not NOT1 (N2624, N2621);
nor NOR3 (N2625, N2611, N776, N2569);
nor NOR4 (N2626, N2618, N1803, N2066, N515);
and AND3 (N2627, N2625, N1314, N310);
nor NOR3 (N2628, N2627, N2420, N331);
and AND3 (N2629, N2622, N1234, N2474);
nand NAND3 (N2630, N2629, N2405, N2361);
nand NAND3 (N2631, N2617, N1033, N551);
xor XOR2 (N2632, N2614, N2030);
nor NOR4 (N2633, N2626, N1410, N1342, N1821);
nand NAND3 (N2634, N2608, N2188, N769);
not NOT1 (N2635, N2633);
buf BUF1 (N2636, N2620);
not NOT1 (N2637, N2630);
or OR3 (N2638, N2632, N1246, N671);
and AND4 (N2639, N2636, N37, N2458, N1011);
not NOT1 (N2640, N2639);
nand NAND4 (N2641, N2631, N602, N20, N468);
nand NAND4 (N2642, N2634, N1712, N1335, N1606);
and AND3 (N2643, N2635, N528, N509);
nand NAND3 (N2644, N2637, N2426, N968);
not NOT1 (N2645, N2638);
nand NAND2 (N2646, N2641, N1013);
nor NOR2 (N2647, N2623, N174);
nand NAND3 (N2648, N2624, N534, N1107);
nor NOR4 (N2649, N2644, N500, N159, N2195);
nand NAND2 (N2650, N2646, N964);
and AND3 (N2651, N2640, N1615, N275);
nor NOR3 (N2652, N2642, N162, N460);
not NOT1 (N2653, N2628);
or OR2 (N2654, N2651, N1366);
or OR2 (N2655, N2619, N2541);
xor XOR2 (N2656, N2643, N700);
not NOT1 (N2657, N2653);
nor NOR2 (N2658, N2648, N37);
nor NOR4 (N2659, N2657, N2231, N2603, N2130);
not NOT1 (N2660, N2658);
buf BUF1 (N2661, N2650);
and AND4 (N2662, N2652, N2078, N1149, N684);
nor NOR2 (N2663, N2661, N585);
nand NAND4 (N2664, N2655, N186, N2640, N2370);
nand NAND2 (N2665, N2654, N303);
nand NAND2 (N2666, N2647, N180);
not NOT1 (N2667, N2659);
nor NOR3 (N2668, N2649, N215, N1561);
and AND2 (N2669, N2662, N2109);
and AND4 (N2670, N2660, N740, N1425, N2537);
nor NOR3 (N2671, N2670, N1531, N496);
nor NOR2 (N2672, N2667, N865);
nand NAND2 (N2673, N2668, N455);
nand NAND2 (N2674, N2665, N811);
nor NOR2 (N2675, N2673, N1650);
nor NOR2 (N2676, N2672, N867);
not NOT1 (N2677, N2664);
xor XOR2 (N2678, N2656, N207);
not NOT1 (N2679, N2669);
or OR2 (N2680, N2674, N2635);
xor XOR2 (N2681, N2676, N1664);
buf BUF1 (N2682, N2681);
or OR4 (N2683, N2675, N2099, N850, N1658);
nand NAND2 (N2684, N2679, N887);
not NOT1 (N2685, N2678);
buf BUF1 (N2686, N2684);
not NOT1 (N2687, N2671);
and AND3 (N2688, N2687, N1145, N67);
nor NOR3 (N2689, N2682, N1845, N720);
not NOT1 (N2690, N2680);
and AND3 (N2691, N2645, N820, N185);
and AND2 (N2692, N2686, N2089);
xor XOR2 (N2693, N2688, N885);
nor NOR3 (N2694, N2689, N1297, N1983);
nor NOR3 (N2695, N2694, N2588, N1198);
and AND2 (N2696, N2677, N405);
or OR2 (N2697, N2683, N1730);
not NOT1 (N2698, N2693);
nor NOR3 (N2699, N2696, N1111, N2083);
not NOT1 (N2700, N2697);
nand NAND2 (N2701, N2695, N362);
or OR3 (N2702, N2691, N2469, N1358);
buf BUF1 (N2703, N2666);
xor XOR2 (N2704, N2685, N2126);
or OR2 (N2705, N2702, N1677);
nand NAND4 (N2706, N2703, N913, N2652, N2049);
or OR2 (N2707, N2699, N1877);
and AND4 (N2708, N2707, N601, N464, N1300);
buf BUF1 (N2709, N2705);
not NOT1 (N2710, N2709);
and AND3 (N2711, N2690, N2300, N1599);
or OR2 (N2712, N2663, N1042);
not NOT1 (N2713, N2706);
nor NOR4 (N2714, N2692, N474, N2208, N2120);
and AND2 (N2715, N2698, N2648);
nand NAND2 (N2716, N2714, N114);
nand NAND2 (N2717, N2713, N1559);
or OR3 (N2718, N2716, N2259, N850);
xor XOR2 (N2719, N2718, N407);
nor NOR2 (N2720, N2708, N1312);
not NOT1 (N2721, N2704);
buf BUF1 (N2722, N2710);
and AND4 (N2723, N2719, N43, N1031, N2111);
nand NAND4 (N2724, N2700, N2082, N499, N246);
or OR3 (N2725, N2722, N287, N1496);
or OR2 (N2726, N2712, N2389);
xor XOR2 (N2727, N2720, N2262);
buf BUF1 (N2728, N2724);
nor NOR2 (N2729, N2701, N174);
buf BUF1 (N2730, N2727);
not NOT1 (N2731, N2730);
buf BUF1 (N2732, N2728);
or OR3 (N2733, N2721, N641, N1333);
nand NAND2 (N2734, N2711, N2467);
not NOT1 (N2735, N2731);
nand NAND4 (N2736, N2734, N599, N1550, N637);
buf BUF1 (N2737, N2717);
nor NOR4 (N2738, N2726, N1432, N275, N497);
nor NOR3 (N2739, N2733, N2052, N688);
buf BUF1 (N2740, N2729);
nor NOR3 (N2741, N2736, N663, N16);
not NOT1 (N2742, N2732);
nor NOR2 (N2743, N2742, N1798);
not NOT1 (N2744, N2743);
not NOT1 (N2745, N2740);
and AND3 (N2746, N2741, N2048, N1791);
nor NOR2 (N2747, N2745, N2552);
and AND4 (N2748, N2746, N1046, N1469, N594);
not NOT1 (N2749, N2738);
nand NAND3 (N2750, N2725, N1465, N140);
nand NAND4 (N2751, N2739, N1086, N2340, N2189);
buf BUF1 (N2752, N2750);
not NOT1 (N2753, N2748);
and AND2 (N2754, N2749, N1944);
not NOT1 (N2755, N2737);
and AND3 (N2756, N2747, N875, N1279);
buf BUF1 (N2757, N2751);
nor NOR4 (N2758, N2756, N2037, N2592, N1715);
nand NAND4 (N2759, N2754, N2250, N2607, N897);
xor XOR2 (N2760, N2753, N2394);
nor NOR4 (N2761, N2752, N1701, N2604, N2261);
nor NOR4 (N2762, N2723, N1723, N596, N2396);
nor NOR3 (N2763, N2759, N1993, N1860);
xor XOR2 (N2764, N2755, N2701);
buf BUF1 (N2765, N2760);
buf BUF1 (N2766, N2761);
not NOT1 (N2767, N2765);
xor XOR2 (N2768, N2735, N2252);
nand NAND2 (N2769, N2763, N2090);
and AND2 (N2770, N2715, N36);
and AND3 (N2771, N2770, N1606, N846);
buf BUF1 (N2772, N2762);
or OR2 (N2773, N2764, N935);
nor NOR2 (N2774, N2771, N2573);
and AND3 (N2775, N2744, N2415, N2138);
and AND2 (N2776, N2767, N2386);
nand NAND3 (N2777, N2766, N1228, N662);
not NOT1 (N2778, N2758);
buf BUF1 (N2779, N2757);
or OR2 (N2780, N2776, N1224);
nand NAND3 (N2781, N2779, N1582, N88);
xor XOR2 (N2782, N2773, N256);
not NOT1 (N2783, N2774);
buf BUF1 (N2784, N2782);
or OR2 (N2785, N2781, N1005);
buf BUF1 (N2786, N2775);
and AND3 (N2787, N2778, N789, N2284);
nand NAND4 (N2788, N2786, N928, N1042, N2251);
xor XOR2 (N2789, N2769, N1165);
nand NAND2 (N2790, N2788, N1249);
buf BUF1 (N2791, N2784);
and AND4 (N2792, N2787, N36, N1806, N262);
and AND3 (N2793, N2791, N41, N1726);
and AND4 (N2794, N2785, N1515, N2722, N1673);
xor XOR2 (N2795, N2783, N816);
xor XOR2 (N2796, N2792, N1029);
xor XOR2 (N2797, N2772, N246);
not NOT1 (N2798, N2789);
and AND2 (N2799, N2790, N1899);
xor XOR2 (N2800, N2777, N1046);
nor NOR2 (N2801, N2800, N276);
xor XOR2 (N2802, N2797, N592);
xor XOR2 (N2803, N2798, N1208);
or OR2 (N2804, N2780, N970);
xor XOR2 (N2805, N2795, N2010);
buf BUF1 (N2806, N2802);
xor XOR2 (N2807, N2806, N2197);
nand NAND3 (N2808, N2803, N539, N2166);
and AND2 (N2809, N2799, N141);
and AND3 (N2810, N2793, N2416, N2536);
nor NOR4 (N2811, N2805, N1597, N2658, N2687);
nor NOR2 (N2812, N2801, N2472);
xor XOR2 (N2813, N2796, N2300);
xor XOR2 (N2814, N2810, N1246);
not NOT1 (N2815, N2807);
not NOT1 (N2816, N2804);
not NOT1 (N2817, N2811);
or OR3 (N2818, N2817, N201, N2133);
and AND3 (N2819, N2808, N2436, N2000);
nand NAND3 (N2820, N2815, N1927, N102);
xor XOR2 (N2821, N2809, N1841);
nor NOR4 (N2822, N2768, N767, N1666, N2540);
xor XOR2 (N2823, N2821, N1168);
and AND2 (N2824, N2816, N2566);
nor NOR3 (N2825, N2812, N74, N1052);
nand NAND4 (N2826, N2820, N2379, N1876, N877);
or OR4 (N2827, N2826, N841, N1778, N1229);
nand NAND4 (N2828, N2824, N1048, N351, N893);
nand NAND2 (N2829, N2825, N2281);
buf BUF1 (N2830, N2822);
buf BUF1 (N2831, N2814);
nor NOR3 (N2832, N2828, N2299, N2358);
nor NOR3 (N2833, N2794, N671, N1196);
nor NOR4 (N2834, N2819, N551, N1252, N1952);
not NOT1 (N2835, N2818);
buf BUF1 (N2836, N2829);
and AND2 (N2837, N2831, N1396);
nor NOR3 (N2838, N2823, N1430, N1267);
buf BUF1 (N2839, N2813);
or OR3 (N2840, N2834, N1406, N2029);
xor XOR2 (N2841, N2827, N1741);
buf BUF1 (N2842, N2835);
nor NOR3 (N2843, N2842, N696, N473);
not NOT1 (N2844, N2836);
nor NOR4 (N2845, N2839, N1412, N674, N632);
or OR3 (N2846, N2843, N318, N1133);
nand NAND4 (N2847, N2830, N1690, N724, N1072);
nand NAND2 (N2848, N2837, N365);
nand NAND2 (N2849, N2847, N1087);
or OR4 (N2850, N2833, N2146, N12, N2193);
or OR3 (N2851, N2846, N1910, N2785);
buf BUF1 (N2852, N2851);
or OR2 (N2853, N2845, N2181);
not NOT1 (N2854, N2832);
and AND4 (N2855, N2841, N675, N970, N2217);
xor XOR2 (N2856, N2853, N1419);
xor XOR2 (N2857, N2849, N2613);
buf BUF1 (N2858, N2857);
buf BUF1 (N2859, N2838);
and AND4 (N2860, N2854, N929, N2415, N417);
nor NOR2 (N2861, N2850, N2789);
not NOT1 (N2862, N2858);
not NOT1 (N2863, N2840);
xor XOR2 (N2864, N2848, N2128);
not NOT1 (N2865, N2852);
not NOT1 (N2866, N2855);
and AND3 (N2867, N2864, N144, N2457);
xor XOR2 (N2868, N2861, N1506);
nand NAND3 (N2869, N2859, N1813, N2594);
and AND4 (N2870, N2865, N422, N2860, N180);
or OR2 (N2871, N2642, N2566);
buf BUF1 (N2872, N2863);
buf BUF1 (N2873, N2872);
nor NOR4 (N2874, N2856, N2483, N2295, N316);
not NOT1 (N2875, N2874);
buf BUF1 (N2876, N2869);
not NOT1 (N2877, N2873);
xor XOR2 (N2878, N2876, N553);
or OR2 (N2879, N2868, N658);
or OR2 (N2880, N2866, N2000);
nor NOR4 (N2881, N2867, N1546, N864, N1438);
nor NOR3 (N2882, N2879, N548, N2543);
buf BUF1 (N2883, N2877);
and AND3 (N2884, N2844, N300, N2845);
and AND3 (N2885, N2875, N1158, N260);
nor NOR3 (N2886, N2882, N1941, N714);
not NOT1 (N2887, N2886);
nor NOR3 (N2888, N2871, N2525, N1906);
or OR2 (N2889, N2870, N2713);
nand NAND4 (N2890, N2878, N1328, N1116, N1232);
not NOT1 (N2891, N2881);
buf BUF1 (N2892, N2884);
or OR2 (N2893, N2889, N2114);
xor XOR2 (N2894, N2893, N967);
nand NAND2 (N2895, N2880, N1342);
xor XOR2 (N2896, N2888, N1888);
nor NOR2 (N2897, N2894, N560);
nand NAND3 (N2898, N2896, N317, N1990);
or OR3 (N2899, N2885, N2206, N2700);
and AND4 (N2900, N2890, N335, N2612, N2893);
nand NAND2 (N2901, N2891, N102);
buf BUF1 (N2902, N2901);
nor NOR4 (N2903, N2902, N1625, N1678, N289);
xor XOR2 (N2904, N2903, N1317);
nand NAND2 (N2905, N2895, N2857);
or OR3 (N2906, N2897, N2417, N510);
nand NAND4 (N2907, N2904, N484, N1076, N1726);
nand NAND2 (N2908, N2905, N1864);
nor NOR2 (N2909, N2908, N2500);
buf BUF1 (N2910, N2909);
or OR2 (N2911, N2862, N93);
xor XOR2 (N2912, N2906, N1986);
not NOT1 (N2913, N2898);
buf BUF1 (N2914, N2892);
nand NAND3 (N2915, N2910, N2362, N1430);
and AND4 (N2916, N2887, N1655, N701, N1066);
nor NOR3 (N2917, N2912, N2824, N2089);
nor NOR3 (N2918, N2900, N2042, N741);
xor XOR2 (N2919, N2914, N2133);
and AND3 (N2920, N2899, N2034, N1837);
not NOT1 (N2921, N2916);
nand NAND2 (N2922, N2919, N2347);
nor NOR3 (N2923, N2918, N1316, N2118);
buf BUF1 (N2924, N2907);
buf BUF1 (N2925, N2920);
or OR3 (N2926, N2921, N232, N2743);
buf BUF1 (N2927, N2883);
nor NOR4 (N2928, N2927, N1472, N874, N1396);
buf BUF1 (N2929, N2923);
nand NAND3 (N2930, N2928, N1717, N1348);
nand NAND3 (N2931, N2917, N763, N2248);
nand NAND4 (N2932, N2930, N2569, N711, N2697);
not NOT1 (N2933, N2924);
buf BUF1 (N2934, N2915);
buf BUF1 (N2935, N2913);
xor XOR2 (N2936, N2922, N1771);
nor NOR3 (N2937, N2934, N2121, N1845);
nand NAND4 (N2938, N2926, N537, N2222, N48);
not NOT1 (N2939, N2932);
nor NOR4 (N2940, N2911, N1349, N147, N2617);
not NOT1 (N2941, N2931);
or OR3 (N2942, N2936, N2923, N614);
buf BUF1 (N2943, N2942);
nor NOR2 (N2944, N2937, N2276);
or OR2 (N2945, N2943, N950);
nor NOR2 (N2946, N2933, N1883);
xor XOR2 (N2947, N2944, N465);
not NOT1 (N2948, N2940);
nor NOR4 (N2949, N2939, N1529, N932, N1125);
buf BUF1 (N2950, N2948);
nor NOR3 (N2951, N2938, N1929, N233);
or OR3 (N2952, N2949, N800, N759);
or OR2 (N2953, N2935, N432);
nor NOR4 (N2954, N2952, N810, N2005, N2068);
and AND2 (N2955, N2951, N2079);
or OR3 (N2956, N2950, N351, N557);
xor XOR2 (N2957, N2956, N1804);
xor XOR2 (N2958, N2945, N127);
and AND2 (N2959, N2957, N1181);
nand NAND2 (N2960, N2929, N1699);
not NOT1 (N2961, N2954);
buf BUF1 (N2962, N2955);
or OR2 (N2963, N2953, N459);
xor XOR2 (N2964, N2961, N2698);
xor XOR2 (N2965, N2959, N2843);
and AND2 (N2966, N2925, N1347);
and AND2 (N2967, N2966, N254);
and AND4 (N2968, N2941, N2475, N426, N418);
not NOT1 (N2969, N2946);
nand NAND3 (N2970, N2965, N539, N1948);
or OR2 (N2971, N2963, N1587);
and AND2 (N2972, N2958, N6);
xor XOR2 (N2973, N2964, N928);
nor NOR2 (N2974, N2947, N2864);
or OR3 (N2975, N2960, N11, N223);
nand NAND3 (N2976, N2970, N1302, N1311);
xor XOR2 (N2977, N2973, N1403);
nand NAND4 (N2978, N2968, N2409, N712, N522);
not NOT1 (N2979, N2971);
nor NOR3 (N2980, N2976, N955, N503);
and AND3 (N2981, N2978, N2805, N1966);
not NOT1 (N2982, N2981);
nand NAND2 (N2983, N2969, N2299);
not NOT1 (N2984, N2975);
and AND2 (N2985, N2974, N762);
not NOT1 (N2986, N2977);
nor NOR4 (N2987, N2986, N1069, N457, N611);
nor NOR2 (N2988, N2982, N2942);
or OR4 (N2989, N2979, N2858, N86, N2088);
buf BUF1 (N2990, N2967);
buf BUF1 (N2991, N2985);
buf BUF1 (N2992, N2991);
buf BUF1 (N2993, N2992);
or OR2 (N2994, N2984, N2286);
not NOT1 (N2995, N2962);
nand NAND2 (N2996, N2995, N984);
nor NOR3 (N2997, N2990, N2275, N2111);
and AND4 (N2998, N2989, N1520, N1542, N448);
or OR2 (N2999, N2997, N239);
nor NOR2 (N3000, N2987, N1721);
nand NAND2 (N3001, N2983, N666);
not NOT1 (N3002, N2996);
and AND3 (N3003, N3000, N42, N56);
or OR3 (N3004, N2972, N1249, N416);
not NOT1 (N3005, N2993);
not NOT1 (N3006, N2988);
not NOT1 (N3007, N3002);
nor NOR3 (N3008, N3004, N2956, N2470);
nand NAND2 (N3009, N3006, N574);
nor NOR2 (N3010, N3008, N2233);
nand NAND4 (N3011, N2999, N1211, N2783, N1768);
buf BUF1 (N3012, N2998);
xor XOR2 (N3013, N3009, N2189);
and AND3 (N3014, N3007, N373, N490);
xor XOR2 (N3015, N3005, N324);
nor NOR4 (N3016, N2980, N630, N1383, N2000);
not NOT1 (N3017, N2994);
buf BUF1 (N3018, N3017);
or OR4 (N3019, N3018, N445, N1848, N2234);
or OR4 (N3020, N3015, N2116, N2425, N2091);
not NOT1 (N3021, N3013);
nor NOR3 (N3022, N3014, N2545, N1668);
not NOT1 (N3023, N3001);
or OR4 (N3024, N3023, N1699, N1251, N727);
buf BUF1 (N3025, N3020);
nand NAND4 (N3026, N3024, N1353, N1019, N2550);
and AND4 (N3027, N3011, N1486, N677, N1373);
nand NAND3 (N3028, N3012, N1298, N1875);
nand NAND2 (N3029, N3021, N1246);
nand NAND3 (N3030, N3019, N1718, N1208);
or OR3 (N3031, N3028, N494, N69);
buf BUF1 (N3032, N3029);
not NOT1 (N3033, N3003);
nand NAND3 (N3034, N3027, N2581, N636);
or OR3 (N3035, N3033, N2271, N2057);
nor NOR3 (N3036, N3031, N1081, N1830);
nor NOR2 (N3037, N3036, N375);
or OR4 (N3038, N3010, N2303, N1717, N2418);
buf BUF1 (N3039, N3034);
not NOT1 (N3040, N3022);
nand NAND2 (N3041, N3032, N2349);
nand NAND2 (N3042, N3025, N2111);
not NOT1 (N3043, N3041);
not NOT1 (N3044, N3043);
xor XOR2 (N3045, N3030, N1059);
not NOT1 (N3046, N3035);
nor NOR3 (N3047, N3039, N1675, N712);
xor XOR2 (N3048, N3044, N2580);
and AND2 (N3049, N3048, N1724);
xor XOR2 (N3050, N3045, N2450);
nand NAND4 (N3051, N3046, N1637, N1070, N498);
nand NAND4 (N3052, N3038, N2744, N2248, N2770);
nor NOR4 (N3053, N3037, N2977, N1896, N871);
not NOT1 (N3054, N3052);
buf BUF1 (N3055, N3047);
or OR2 (N3056, N3049, N2148);
not NOT1 (N3057, N3040);
not NOT1 (N3058, N3016);
nor NOR4 (N3059, N3055, N362, N2719, N884);
or OR4 (N3060, N3054, N2529, N2389, N594);
or OR4 (N3061, N3059, N2930, N874, N1774);
not NOT1 (N3062, N3050);
nand NAND4 (N3063, N3058, N2357, N1413, N523);
xor XOR2 (N3064, N3051, N1938);
buf BUF1 (N3065, N3062);
nor NOR2 (N3066, N3064, N1187);
buf BUF1 (N3067, N3053);
xor XOR2 (N3068, N3057, N2083);
or OR4 (N3069, N3042, N2882, N1883, N524);
or OR2 (N3070, N3056, N1243);
buf BUF1 (N3071, N3026);
and AND2 (N3072, N3061, N2765);
and AND3 (N3073, N3070, N1856, N2320);
nor NOR3 (N3074, N3067, N90, N990);
xor XOR2 (N3075, N3065, N2648);
nor NOR3 (N3076, N3069, N1619, N1378);
nand NAND3 (N3077, N3068, N1043, N2825);
nand NAND2 (N3078, N3063, N1051);
buf BUF1 (N3079, N3060);
and AND3 (N3080, N3077, N163, N111);
nor NOR3 (N3081, N3072, N116, N419);
nor NOR3 (N3082, N3074, N2068, N3019);
nor NOR4 (N3083, N3082, N174, N2553, N980);
or OR3 (N3084, N3078, N1784, N1780);
nor NOR4 (N3085, N3076, N1251, N1286, N1542);
and AND2 (N3086, N3073, N2716);
nand NAND3 (N3087, N3081, N989, N966);
xor XOR2 (N3088, N3075, N2555);
xor XOR2 (N3089, N3086, N2952);
not NOT1 (N3090, N3080);
or OR2 (N3091, N3087, N2419);
xor XOR2 (N3092, N3089, N1138);
buf BUF1 (N3093, N3066);
nor NOR2 (N3094, N3071, N692);
or OR2 (N3095, N3088, N955);
not NOT1 (N3096, N3094);
or OR3 (N3097, N3083, N65, N2904);
nor NOR4 (N3098, N3090, N1758, N3060, N857);
nand NAND4 (N3099, N3097, N188, N999, N2988);
xor XOR2 (N3100, N3095, N574);
or OR3 (N3101, N3084, N51, N2897);
not NOT1 (N3102, N3092);
and AND2 (N3103, N3101, N1517);
not NOT1 (N3104, N3100);
and AND4 (N3105, N3103, N221, N2105, N3041);
nor NOR3 (N3106, N3091, N981, N411);
nand NAND4 (N3107, N3105, N1925, N900, N343);
buf BUF1 (N3108, N3093);
not NOT1 (N3109, N3079);
nand NAND4 (N3110, N3102, N456, N1191, N748);
nor NOR3 (N3111, N3110, N714, N2758);
or OR4 (N3112, N3096, N1594, N15, N68);
not NOT1 (N3113, N3108);
xor XOR2 (N3114, N3099, N231);
nand NAND4 (N3115, N3085, N996, N1856, N52);
xor XOR2 (N3116, N3111, N2901);
nor NOR3 (N3117, N3104, N1259, N2433);
and AND4 (N3118, N3115, N2956, N2942, N2554);
not NOT1 (N3119, N3117);
nand NAND2 (N3120, N3112, N213);
nor NOR2 (N3121, N3098, N2381);
and AND4 (N3122, N3118, N3010, N1362, N1835);
xor XOR2 (N3123, N3114, N1070);
nor NOR3 (N3124, N3116, N1138, N2841);
or OR4 (N3125, N3121, N1821, N1500, N2023);
xor XOR2 (N3126, N3120, N1285);
xor XOR2 (N3127, N3122, N2114);
buf BUF1 (N3128, N3125);
nor NOR3 (N3129, N3119, N886, N1539);
xor XOR2 (N3130, N3124, N2733);
buf BUF1 (N3131, N3106);
xor XOR2 (N3132, N3126, N1140);
or OR2 (N3133, N3129, N385);
xor XOR2 (N3134, N3128, N1952);
buf BUF1 (N3135, N3130);
and AND4 (N3136, N3127, N228, N853, N1944);
and AND4 (N3137, N3132, N2581, N1456, N1463);
buf BUF1 (N3138, N3109);
and AND4 (N3139, N3123, N1545, N259, N905);
nor NOR2 (N3140, N3139, N1941);
nor NOR3 (N3141, N3135, N2892, N621);
buf BUF1 (N3142, N3137);
buf BUF1 (N3143, N3133);
buf BUF1 (N3144, N3141);
nand NAND2 (N3145, N3136, N411);
buf BUF1 (N3146, N3138);
nand NAND3 (N3147, N3113, N2158, N1965);
or OR4 (N3148, N3140, N704, N2322, N797);
not NOT1 (N3149, N3148);
nand NAND2 (N3150, N3143, N1447);
buf BUF1 (N3151, N3142);
nor NOR4 (N3152, N3151, N64, N1805, N1263);
nor NOR2 (N3153, N3134, N1599);
xor XOR2 (N3154, N3146, N684);
nand NAND2 (N3155, N3150, N385);
or OR3 (N3156, N3147, N1127, N2902);
xor XOR2 (N3157, N3156, N22);
nand NAND3 (N3158, N3149, N2917, N1832);
or OR4 (N3159, N3153, N1012, N871, N1645);
nand NAND3 (N3160, N3154, N853, N910);
and AND3 (N3161, N3159, N1732, N2356);
or OR3 (N3162, N3155, N2241, N795);
not NOT1 (N3163, N3160);
buf BUF1 (N3164, N3131);
not NOT1 (N3165, N3152);
and AND2 (N3166, N3161, N992);
and AND3 (N3167, N3107, N1881, N1366);
nor NOR2 (N3168, N3165, N863);
nor NOR2 (N3169, N3162, N2604);
xor XOR2 (N3170, N3166, N1457);
not NOT1 (N3171, N3158);
nand NAND2 (N3172, N3157, N3106);
buf BUF1 (N3173, N3171);
xor XOR2 (N3174, N3164, N573);
buf BUF1 (N3175, N3168);
or OR4 (N3176, N3170, N2325, N808, N534);
xor XOR2 (N3177, N3167, N1403);
or OR4 (N3178, N3169, N3099, N979, N2855);
buf BUF1 (N3179, N3144);
buf BUF1 (N3180, N3175);
and AND4 (N3181, N3180, N2021, N1477, N2522);
nand NAND3 (N3182, N3173, N1932, N939);
buf BUF1 (N3183, N3145);
nor NOR3 (N3184, N3183, N3137, N1847);
xor XOR2 (N3185, N3176, N1897);
nand NAND4 (N3186, N3179, N822, N2255, N1699);
buf BUF1 (N3187, N3186);
xor XOR2 (N3188, N3163, N186);
nand NAND3 (N3189, N3178, N2522, N207);
buf BUF1 (N3190, N3177);
and AND4 (N3191, N3172, N81, N1291, N2422);
buf BUF1 (N3192, N3187);
xor XOR2 (N3193, N3192, N2836);
not NOT1 (N3194, N3182);
xor XOR2 (N3195, N3185, N1536);
nand NAND2 (N3196, N3188, N2832);
not NOT1 (N3197, N3184);
or OR2 (N3198, N3191, N340);
nor NOR2 (N3199, N3174, N721);
nor NOR2 (N3200, N3198, N596);
nand NAND4 (N3201, N3196, N1067, N1020, N3122);
or OR2 (N3202, N3194, N3035);
or OR3 (N3203, N3189, N1647, N2613);
nor NOR3 (N3204, N3195, N3043, N2267);
nand NAND2 (N3205, N3193, N1819);
and AND2 (N3206, N3203, N1921);
not NOT1 (N3207, N3205);
nor NOR4 (N3208, N3201, N955, N2771, N874);
buf BUF1 (N3209, N3204);
nand NAND4 (N3210, N3181, N1232, N2829, N2058);
xor XOR2 (N3211, N3210, N3125);
xor XOR2 (N3212, N3200, N1331);
buf BUF1 (N3213, N3207);
buf BUF1 (N3214, N3209);
nand NAND2 (N3215, N3214, N2356);
nand NAND4 (N3216, N3206, N948, N1835, N2640);
nor NOR4 (N3217, N3215, N785, N2772, N291);
and AND3 (N3218, N3217, N3144, N1329);
endmodule