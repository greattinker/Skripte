// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;

output N708,N692,N697,N676,N710,N707,N709,N705,N704,N711;

nor NOR3 (N12, N9, N5, N3);
not NOT1 (N13, N10);
nand NAND4 (N14, N3, N7, N6, N11);
or OR4 (N15, N13, N10, N13, N1);
or OR3 (N16, N10, N1, N6);
or OR2 (N17, N9, N3);
nand NAND2 (N18, N1, N17);
or OR2 (N19, N17, N7);
nand NAND2 (N20, N19, N11);
nand NAND3 (N21, N11, N20, N20);
or OR4 (N22, N11, N9, N20, N15);
and AND4 (N23, N7, N9, N18, N13);
not NOT1 (N24, N3);
nor NOR4 (N25, N8, N2, N7, N8);
not NOT1 (N26, N23);
nor NOR4 (N27, N7, N6, N23, N20);
buf BUF1 (N28, N14);
nand NAND3 (N29, N22, N2, N6);
or OR4 (N30, N24, N13, N5, N11);
and AND2 (N31, N5, N15);
not NOT1 (N32, N16);
nand NAND4 (N33, N21, N27, N5, N16);
and AND3 (N34, N13, N16, N7);
or OR2 (N35, N30, N5);
buf BUF1 (N36, N12);
or OR2 (N37, N32, N3);
and AND3 (N38, N36, N35, N14);
buf BUF1 (N39, N10);
nor NOR4 (N40, N25, N12, N4, N21);
nor NOR2 (N41, N38, N3);
nor NOR4 (N42, N41, N16, N8, N23);
xor XOR2 (N43, N31, N28);
xor XOR2 (N44, N32, N12);
and AND3 (N45, N37, N13, N42);
buf BUF1 (N46, N41);
buf BUF1 (N47, N29);
xor XOR2 (N48, N44, N2);
buf BUF1 (N49, N48);
or OR3 (N50, N49, N23, N18);
nand NAND4 (N51, N47, N42, N42, N37);
xor XOR2 (N52, N46, N27);
or OR4 (N53, N39, N4, N20, N26);
buf BUF1 (N54, N37);
or OR3 (N55, N43, N27, N53);
not NOT1 (N56, N51);
and AND2 (N57, N35, N10);
buf BUF1 (N58, N33);
and AND4 (N59, N45, N45, N20, N20);
xor XOR2 (N60, N56, N59);
not NOT1 (N61, N33);
buf BUF1 (N62, N61);
xor XOR2 (N63, N50, N44);
buf BUF1 (N64, N62);
nor NOR4 (N65, N60, N15, N21, N20);
or OR4 (N66, N57, N52, N34, N19);
buf BUF1 (N67, N18);
nand NAND3 (N68, N23, N22, N28);
nor NOR2 (N69, N65, N28);
nand NAND4 (N70, N58, N49, N63, N13);
and AND2 (N71, N43, N48);
nand NAND4 (N72, N68, N53, N60, N29);
or OR3 (N73, N67, N51, N42);
nand NAND3 (N74, N40, N21, N70);
and AND4 (N75, N48, N66, N46, N54);
nand NAND3 (N76, N49, N11, N21);
nand NAND4 (N77, N63, N48, N28, N31);
not NOT1 (N78, N55);
nor NOR3 (N79, N75, N41, N8);
xor XOR2 (N80, N64, N5);
not NOT1 (N81, N71);
nand NAND2 (N82, N81, N77);
nor NOR4 (N83, N16, N37, N39, N19);
not NOT1 (N84, N82);
nand NAND2 (N85, N83, N83);
and AND3 (N86, N69, N82, N77);
buf BUF1 (N87, N73);
or OR2 (N88, N80, N82);
xor XOR2 (N89, N76, N47);
or OR3 (N90, N86, N78, N23);
nor NOR3 (N91, N3, N18, N10);
xor XOR2 (N92, N87, N45);
nor NOR4 (N93, N85, N9, N66, N62);
buf BUF1 (N94, N79);
nand NAND2 (N95, N84, N43);
and AND3 (N96, N88, N46, N16);
buf BUF1 (N97, N72);
or OR2 (N98, N97, N5);
not NOT1 (N99, N98);
nand NAND3 (N100, N92, N17, N71);
nor NOR3 (N101, N74, N23, N60);
or OR4 (N102, N93, N58, N49, N92);
or OR4 (N103, N99, N100, N37, N16);
nand NAND2 (N104, N37, N50);
nand NAND3 (N105, N102, N20, N64);
not NOT1 (N106, N90);
not NOT1 (N107, N95);
xor XOR2 (N108, N103, N86);
not NOT1 (N109, N101);
buf BUF1 (N110, N108);
nand NAND2 (N111, N91, N24);
buf BUF1 (N112, N96);
nand NAND3 (N113, N94, N3, N28);
and AND2 (N114, N106, N12);
xor XOR2 (N115, N113, N80);
nand NAND3 (N116, N111, N8, N81);
not NOT1 (N117, N114);
xor XOR2 (N118, N112, N78);
buf BUF1 (N119, N109);
buf BUF1 (N120, N107);
nor NOR3 (N121, N105, N73, N48);
not NOT1 (N122, N117);
nand NAND4 (N123, N110, N110, N58, N88);
or OR4 (N124, N118, N17, N98, N85);
or OR2 (N125, N104, N15);
and AND4 (N126, N120, N109, N78, N71);
buf BUF1 (N127, N121);
buf BUF1 (N128, N89);
buf BUF1 (N129, N116);
and AND2 (N130, N122, N33);
nand NAND4 (N131, N129, N21, N34, N119);
not NOT1 (N132, N105);
nand NAND4 (N133, N131, N95, N51, N52);
and AND3 (N134, N130, N101, N81);
nand NAND3 (N135, N125, N87, N3);
buf BUF1 (N136, N135);
xor XOR2 (N137, N128, N21);
xor XOR2 (N138, N127, N92);
buf BUF1 (N139, N124);
not NOT1 (N140, N126);
buf BUF1 (N141, N136);
buf BUF1 (N142, N137);
xor XOR2 (N143, N139, N84);
buf BUF1 (N144, N132);
nor NOR2 (N145, N144, N59);
not NOT1 (N146, N138);
nor NOR3 (N147, N123, N139, N51);
nor NOR4 (N148, N145, N72, N124, N95);
buf BUF1 (N149, N147);
nand NAND4 (N150, N115, N47, N94, N98);
buf BUF1 (N151, N148);
not NOT1 (N152, N134);
nand NAND2 (N153, N150, N38);
or OR3 (N154, N142, N49, N127);
nand NAND2 (N155, N153, N62);
not NOT1 (N156, N154);
nand NAND2 (N157, N152, N99);
nor NOR3 (N158, N157, N52, N33);
not NOT1 (N159, N141);
nor NOR4 (N160, N155, N16, N15, N55);
xor XOR2 (N161, N146, N39);
not NOT1 (N162, N143);
or OR3 (N163, N161, N130, N52);
xor XOR2 (N164, N140, N44);
not NOT1 (N165, N156);
nand NAND3 (N166, N159, N43, N66);
buf BUF1 (N167, N164);
nand NAND4 (N168, N151, N48, N161, N35);
nor NOR3 (N169, N160, N105, N10);
or OR2 (N170, N169, N71);
or OR3 (N171, N158, N45, N84);
and AND2 (N172, N162, N22);
not NOT1 (N173, N168);
and AND3 (N174, N163, N123, N52);
and AND2 (N175, N170, N119);
or OR2 (N176, N166, N148);
not NOT1 (N177, N165);
nor NOR4 (N178, N173, N29, N142, N30);
buf BUF1 (N179, N167);
and AND3 (N180, N171, N38, N158);
buf BUF1 (N181, N172);
xor XOR2 (N182, N174, N155);
or OR2 (N183, N181, N165);
not NOT1 (N184, N180);
and AND2 (N185, N133, N172);
nor NOR4 (N186, N179, N157, N113, N147);
and AND4 (N187, N176, N67, N32, N97);
or OR3 (N188, N185, N181, N37);
buf BUF1 (N189, N182);
xor XOR2 (N190, N184, N148);
or OR3 (N191, N177, N186, N46);
or OR3 (N192, N79, N27, N5);
and AND3 (N193, N190, N187, N143);
not NOT1 (N194, N113);
not NOT1 (N195, N175);
xor XOR2 (N196, N178, N35);
nor NOR2 (N197, N191, N3);
nand NAND4 (N198, N195, N104, N3, N38);
not NOT1 (N199, N183);
or OR4 (N200, N189, N158, N177, N174);
xor XOR2 (N201, N149, N1);
nor NOR3 (N202, N199, N50, N47);
or OR3 (N203, N192, N5, N184);
xor XOR2 (N204, N196, N107);
buf BUF1 (N205, N202);
nor NOR2 (N206, N201, N70);
or OR2 (N207, N205, N126);
or OR2 (N208, N198, N137);
not NOT1 (N209, N208);
or OR2 (N210, N188, N107);
nand NAND2 (N211, N200, N16);
and AND4 (N212, N210, N150, N19, N178);
xor XOR2 (N213, N204, N124);
and AND3 (N214, N193, N147, N166);
or OR2 (N215, N211, N107);
and AND3 (N216, N194, N137, N32);
buf BUF1 (N217, N197);
buf BUF1 (N218, N214);
nor NOR3 (N219, N216, N2, N20);
not NOT1 (N220, N215);
nor NOR4 (N221, N218, N166, N220, N158);
buf BUF1 (N222, N171);
or OR4 (N223, N212, N97, N166, N63);
nand NAND4 (N224, N219, N103, N59, N36);
and AND4 (N225, N221, N32, N121, N21);
xor XOR2 (N226, N213, N102);
buf BUF1 (N227, N217);
nand NAND4 (N228, N209, N53, N110, N182);
nor NOR2 (N229, N223, N137);
or OR4 (N230, N203, N32, N87, N136);
and AND2 (N231, N222, N191);
not NOT1 (N232, N229);
nor NOR2 (N233, N225, N220);
or OR2 (N234, N228, N156);
and AND2 (N235, N224, N11);
nor NOR3 (N236, N234, N165, N84);
nand NAND2 (N237, N233, N68);
xor XOR2 (N238, N206, N94);
and AND2 (N239, N231, N71);
and AND4 (N240, N237, N123, N108, N212);
buf BUF1 (N241, N230);
nor NOR2 (N242, N235, N143);
not NOT1 (N243, N241);
and AND3 (N244, N207, N20, N226);
buf BUF1 (N245, N41);
not NOT1 (N246, N238);
buf BUF1 (N247, N239);
xor XOR2 (N248, N242, N189);
buf BUF1 (N249, N248);
not NOT1 (N250, N236);
or OR3 (N251, N232, N150, N131);
not NOT1 (N252, N243);
and AND3 (N253, N247, N24, N152);
and AND2 (N254, N240, N29);
xor XOR2 (N255, N245, N20);
and AND3 (N256, N251, N159, N131);
and AND3 (N257, N227, N179, N96);
nor NOR3 (N258, N257, N2, N173);
buf BUF1 (N259, N249);
nand NAND3 (N260, N255, N9, N99);
nand NAND2 (N261, N258, N148);
nand NAND4 (N262, N253, N145, N121, N66);
xor XOR2 (N263, N254, N172);
buf BUF1 (N264, N263);
or OR4 (N265, N264, N150, N157, N31);
or OR3 (N266, N262, N126, N207);
or OR3 (N267, N261, N102, N6);
or OR2 (N268, N246, N85);
or OR2 (N269, N252, N203);
nor NOR4 (N270, N256, N10, N55, N183);
not NOT1 (N271, N268);
xor XOR2 (N272, N269, N252);
not NOT1 (N273, N250);
buf BUF1 (N274, N265);
buf BUF1 (N275, N273);
and AND3 (N276, N274, N152, N268);
and AND2 (N277, N276, N80);
or OR4 (N278, N271, N190, N195, N49);
nor NOR3 (N279, N267, N89, N10);
not NOT1 (N280, N278);
or OR2 (N281, N275, N118);
and AND3 (N282, N280, N71, N214);
xor XOR2 (N283, N259, N271);
not NOT1 (N284, N244);
xor XOR2 (N285, N279, N53);
and AND2 (N286, N272, N41);
nand NAND3 (N287, N281, N122, N41);
and AND2 (N288, N266, N37);
xor XOR2 (N289, N285, N236);
buf BUF1 (N290, N270);
nor NOR4 (N291, N286, N137, N150, N232);
not NOT1 (N292, N277);
nand NAND2 (N293, N283, N260);
and AND3 (N294, N27, N210, N133);
and AND4 (N295, N289, N111, N188, N3);
and AND4 (N296, N294, N106, N96, N273);
xor XOR2 (N297, N295, N20);
nand NAND4 (N298, N290, N102, N115, N162);
or OR2 (N299, N288, N290);
nor NOR3 (N300, N287, N267, N267);
nor NOR2 (N301, N297, N248);
or OR3 (N302, N300, N167, N7);
or OR4 (N303, N282, N262, N246, N33);
not NOT1 (N304, N284);
nand NAND4 (N305, N292, N243, N280, N107);
nand NAND4 (N306, N298, N232, N164, N175);
and AND4 (N307, N306, N215, N293, N24);
nand NAND3 (N308, N114, N21, N21);
or OR4 (N309, N304, N183, N173, N11);
nor NOR2 (N310, N303, N187);
xor XOR2 (N311, N291, N76);
and AND4 (N312, N301, N117, N264, N34);
nor NOR3 (N313, N302, N86, N60);
not NOT1 (N314, N305);
not NOT1 (N315, N310);
and AND2 (N316, N296, N69);
and AND3 (N317, N308, N91, N153);
buf BUF1 (N318, N307);
or OR4 (N319, N316, N5, N136, N54);
not NOT1 (N320, N317);
nand NAND3 (N321, N314, N127, N87);
nor NOR2 (N322, N312, N307);
nand NAND2 (N323, N315, N240);
xor XOR2 (N324, N318, N225);
nand NAND4 (N325, N309, N197, N195, N235);
nor NOR4 (N326, N321, N77, N273, N167);
and AND2 (N327, N324, N72);
nand NAND4 (N328, N299, N277, N76, N168);
not NOT1 (N329, N325);
buf BUF1 (N330, N319);
buf BUF1 (N331, N329);
nand NAND4 (N332, N322, N230, N247, N296);
xor XOR2 (N333, N311, N293);
and AND3 (N334, N333, N26, N327);
not NOT1 (N335, N145);
buf BUF1 (N336, N320);
nand NAND2 (N337, N326, N158);
not NOT1 (N338, N336);
nor NOR2 (N339, N328, N107);
xor XOR2 (N340, N337, N168);
and AND3 (N341, N313, N191, N36);
nor NOR4 (N342, N335, N263, N259, N262);
buf BUF1 (N343, N334);
or OR4 (N344, N339, N203, N202, N224);
or OR3 (N345, N342, N288, N282);
and AND3 (N346, N340, N49, N211);
buf BUF1 (N347, N330);
not NOT1 (N348, N343);
or OR4 (N349, N338, N135, N275, N98);
and AND4 (N350, N344, N206, N253, N29);
or OR2 (N351, N345, N213);
or OR3 (N352, N348, N126, N146);
and AND3 (N353, N349, N7, N228);
nor NOR3 (N354, N347, N345, N158);
not NOT1 (N355, N350);
not NOT1 (N356, N323);
nand NAND2 (N357, N354, N114);
nand NAND2 (N358, N331, N334);
not NOT1 (N359, N332);
buf BUF1 (N360, N352);
or OR2 (N361, N358, N297);
xor XOR2 (N362, N360, N296);
not NOT1 (N363, N359);
nor NOR4 (N364, N351, N341, N86, N161);
xor XOR2 (N365, N136, N88);
or OR4 (N366, N356, N93, N52, N267);
nand NAND2 (N367, N363, N254);
buf BUF1 (N368, N364);
and AND3 (N369, N357, N101, N10);
not NOT1 (N370, N361);
buf BUF1 (N371, N370);
nand NAND2 (N372, N368, N91);
not NOT1 (N373, N371);
and AND3 (N374, N365, N278, N342);
nor NOR4 (N375, N353, N318, N117, N245);
and AND2 (N376, N367, N311);
nand NAND4 (N377, N366, N184, N279, N22);
nand NAND3 (N378, N372, N112, N297);
or OR4 (N379, N374, N319, N360, N33);
and AND2 (N380, N379, N73);
nor NOR4 (N381, N375, N225, N18, N371);
or OR4 (N382, N380, N56, N376, N85);
nand NAND3 (N383, N173, N71, N49);
or OR2 (N384, N346, N67);
and AND3 (N385, N377, N9, N196);
not NOT1 (N386, N373);
nand NAND2 (N387, N381, N217);
not NOT1 (N388, N369);
nor NOR2 (N389, N362, N29);
xor XOR2 (N390, N378, N156);
nor NOR2 (N391, N389, N214);
nand NAND2 (N392, N382, N388);
nor NOR3 (N393, N74, N142, N372);
xor XOR2 (N394, N355, N309);
and AND3 (N395, N384, N138, N314);
buf BUF1 (N396, N393);
and AND2 (N397, N387, N320);
nand NAND2 (N398, N394, N120);
nand NAND3 (N399, N391, N208, N304);
and AND4 (N400, N385, N352, N344, N216);
or OR4 (N401, N392, N125, N60, N137);
and AND4 (N402, N390, N363, N244, N340);
nand NAND3 (N403, N383, N108, N182);
or OR3 (N404, N403, N194, N176);
buf BUF1 (N405, N398);
and AND3 (N406, N400, N227, N11);
nor NOR3 (N407, N397, N49, N208);
xor XOR2 (N408, N401, N129);
or OR3 (N409, N405, N139, N322);
buf BUF1 (N410, N409);
or OR3 (N411, N404, N99, N365);
buf BUF1 (N412, N396);
nand NAND2 (N413, N399, N75);
buf BUF1 (N414, N408);
not NOT1 (N415, N411);
buf BUF1 (N416, N413);
nor NOR4 (N417, N407, N198, N157, N202);
not NOT1 (N418, N416);
not NOT1 (N419, N410);
nor NOR4 (N420, N419, N103, N271, N235);
nand NAND2 (N421, N386, N272);
xor XOR2 (N422, N421, N18);
and AND3 (N423, N417, N43, N286);
and AND3 (N424, N423, N381, N201);
and AND3 (N425, N395, N286, N5);
or OR4 (N426, N420, N201, N170, N147);
not NOT1 (N427, N426);
buf BUF1 (N428, N415);
or OR2 (N429, N414, N32);
xor XOR2 (N430, N427, N412);
buf BUF1 (N431, N20);
nand NAND2 (N432, N422, N395);
nand NAND2 (N433, N428, N168);
and AND3 (N434, N429, N177, N119);
or OR4 (N435, N425, N387, N166, N399);
not NOT1 (N436, N431);
nand NAND3 (N437, N402, N24, N274);
buf BUF1 (N438, N434);
nand NAND4 (N439, N436, N82, N28, N126);
or OR3 (N440, N433, N413, N167);
or OR2 (N441, N418, N97);
or OR4 (N442, N437, N438, N201, N428);
xor XOR2 (N443, N116, N126);
and AND4 (N444, N442, N423, N219, N113);
xor XOR2 (N445, N439, N187);
nand NAND3 (N446, N435, N115, N22);
or OR2 (N447, N406, N425);
not NOT1 (N448, N441);
nor NOR3 (N449, N432, N418, N264);
xor XOR2 (N450, N447, N424);
and AND2 (N451, N373, N54);
nor NOR4 (N452, N444, N169, N395, N202);
nand NAND3 (N453, N452, N346, N185);
or OR3 (N454, N430, N268, N8);
nand NAND4 (N455, N448, N94, N44, N400);
nand NAND2 (N456, N443, N414);
nor NOR2 (N457, N453, N325);
nand NAND2 (N458, N446, N25);
nor NOR2 (N459, N454, N267);
xor XOR2 (N460, N457, N38);
or OR3 (N461, N445, N199, N357);
or OR4 (N462, N456, N155, N157, N76);
not NOT1 (N463, N458);
nor NOR4 (N464, N459, N252, N425, N353);
and AND4 (N465, N440, N308, N459, N218);
and AND2 (N466, N460, N306);
buf BUF1 (N467, N455);
not NOT1 (N468, N451);
or OR4 (N469, N463, N438, N198, N310);
nand NAND2 (N470, N467, N265);
buf BUF1 (N471, N461);
buf BUF1 (N472, N469);
nor NOR4 (N473, N468, N378, N222, N191);
not NOT1 (N474, N466);
nor NOR4 (N475, N470, N324, N443, N283);
buf BUF1 (N476, N464);
nand NAND4 (N477, N462, N173, N271, N282);
nor NOR3 (N478, N476, N362, N339);
buf BUF1 (N479, N465);
not NOT1 (N480, N471);
nand NAND4 (N481, N477, N205, N221, N370);
nor NOR2 (N482, N475, N444);
nor NOR4 (N483, N479, N198, N113, N208);
or OR4 (N484, N450, N161, N143, N289);
or OR2 (N485, N480, N258);
not NOT1 (N486, N481);
xor XOR2 (N487, N482, N361);
not NOT1 (N488, N486);
or OR3 (N489, N474, N375, N341);
nor NOR2 (N490, N483, N372);
and AND4 (N491, N473, N77, N13, N274);
nand NAND3 (N492, N484, N243, N375);
buf BUF1 (N493, N487);
nor NOR4 (N494, N493, N452, N54, N27);
nand NAND3 (N495, N472, N91, N410);
not NOT1 (N496, N491);
nor NOR3 (N497, N492, N169, N444);
xor XOR2 (N498, N478, N446);
or OR4 (N499, N497, N22, N25, N44);
not NOT1 (N500, N485);
buf BUF1 (N501, N499);
not NOT1 (N502, N489);
or OR4 (N503, N496, N459, N322, N292);
not NOT1 (N504, N495);
and AND4 (N505, N504, N463, N401, N489);
not NOT1 (N506, N449);
nand NAND2 (N507, N505, N341);
buf BUF1 (N508, N488);
nand NAND4 (N509, N508, N437, N285, N10);
nor NOR3 (N510, N501, N505, N405);
nor NOR2 (N511, N490, N450);
nor NOR2 (N512, N502, N207);
or OR3 (N513, N503, N120, N58);
nor NOR3 (N514, N507, N273, N66);
nor NOR3 (N515, N506, N417, N274);
not NOT1 (N516, N500);
nand NAND4 (N517, N498, N473, N307, N54);
buf BUF1 (N518, N514);
not NOT1 (N519, N510);
nor NOR2 (N520, N511, N467);
nand NAND3 (N521, N512, N249, N143);
nor NOR4 (N522, N519, N386, N329, N402);
nand NAND4 (N523, N509, N360, N105, N457);
not NOT1 (N524, N515);
and AND3 (N525, N521, N394, N23);
xor XOR2 (N526, N524, N66);
nor NOR3 (N527, N518, N9, N226);
nor NOR2 (N528, N513, N349);
nand NAND4 (N529, N525, N55, N108, N62);
nand NAND4 (N530, N517, N295, N177, N197);
xor XOR2 (N531, N520, N232);
xor XOR2 (N532, N516, N380);
and AND3 (N533, N526, N273, N405);
not NOT1 (N534, N530);
nor NOR4 (N535, N534, N93, N342, N273);
or OR4 (N536, N535, N412, N133, N498);
nor NOR3 (N537, N533, N377, N184);
or OR2 (N538, N529, N175);
not NOT1 (N539, N532);
buf BUF1 (N540, N537);
and AND2 (N541, N540, N467);
nor NOR4 (N542, N527, N48, N411, N310);
xor XOR2 (N543, N536, N116);
not NOT1 (N544, N528);
not NOT1 (N545, N544);
buf BUF1 (N546, N531);
not NOT1 (N547, N543);
or OR4 (N548, N542, N335, N61, N251);
and AND3 (N549, N539, N376, N10);
nor NOR2 (N550, N546, N190);
buf BUF1 (N551, N538);
buf BUF1 (N552, N550);
not NOT1 (N553, N522);
nand NAND4 (N554, N523, N87, N544, N10);
nand NAND3 (N555, N541, N241, N22);
buf BUF1 (N556, N548);
not NOT1 (N557, N549);
nand NAND4 (N558, N547, N422, N552, N252);
nand NAND3 (N559, N300, N470, N474);
not NOT1 (N560, N558);
nand NAND3 (N561, N560, N348, N507);
or OR2 (N562, N494, N485);
nor NOR2 (N563, N562, N249);
or OR4 (N564, N563, N505, N168, N394);
xor XOR2 (N565, N553, N335);
nand NAND2 (N566, N565, N323);
buf BUF1 (N567, N561);
or OR4 (N568, N557, N113, N433, N428);
or OR4 (N569, N556, N3, N278, N509);
buf BUF1 (N570, N567);
buf BUF1 (N571, N545);
nand NAND3 (N572, N570, N540, N161);
nor NOR3 (N573, N572, N332, N319);
or OR2 (N574, N564, N537);
nor NOR3 (N575, N551, N144, N377);
xor XOR2 (N576, N559, N87);
nand NAND4 (N577, N566, N210, N176, N372);
and AND3 (N578, N575, N32, N130);
not NOT1 (N579, N576);
buf BUF1 (N580, N579);
or OR2 (N581, N577, N440);
nor NOR4 (N582, N571, N294, N352, N116);
nand NAND4 (N583, N568, N98, N268, N21);
not NOT1 (N584, N573);
not NOT1 (N585, N578);
or OR3 (N586, N584, N546, N508);
nand NAND2 (N587, N585, N179);
not NOT1 (N588, N580);
not NOT1 (N589, N581);
not NOT1 (N590, N582);
nand NAND2 (N591, N589, N387);
or OR2 (N592, N587, N407);
xor XOR2 (N593, N554, N28);
or OR2 (N594, N586, N371);
xor XOR2 (N595, N593, N581);
nand NAND2 (N596, N591, N249);
not NOT1 (N597, N596);
or OR3 (N598, N590, N180, N273);
nor NOR2 (N599, N598, N95);
or OR3 (N600, N594, N355, N257);
buf BUF1 (N601, N595);
not NOT1 (N602, N599);
nand NAND3 (N603, N592, N580, N25);
and AND2 (N604, N583, N1);
nor NOR4 (N605, N588, N83, N63, N536);
xor XOR2 (N606, N574, N434);
buf BUF1 (N607, N604);
and AND2 (N608, N603, N205);
xor XOR2 (N609, N555, N603);
buf BUF1 (N610, N605);
not NOT1 (N611, N601);
nand NAND2 (N612, N609, N504);
and AND4 (N613, N602, N226, N190, N135);
nand NAND3 (N614, N600, N275, N584);
not NOT1 (N615, N606);
and AND4 (N616, N612, N256, N465, N342);
nor NOR2 (N617, N569, N572);
and AND2 (N618, N608, N492);
not NOT1 (N619, N597);
nand NAND3 (N620, N610, N181, N433);
nand NAND3 (N621, N618, N117, N7);
and AND4 (N622, N614, N364, N396, N300);
xor XOR2 (N623, N620, N297);
xor XOR2 (N624, N611, N492);
nor NOR3 (N625, N619, N80, N46);
xor XOR2 (N626, N621, N137);
not NOT1 (N627, N624);
and AND4 (N628, N623, N425, N428, N53);
xor XOR2 (N629, N617, N244);
xor XOR2 (N630, N622, N526);
buf BUF1 (N631, N616);
nand NAND3 (N632, N625, N66, N545);
xor XOR2 (N633, N628, N542);
not NOT1 (N634, N630);
or OR3 (N635, N615, N165, N59);
nand NAND4 (N636, N631, N17, N351, N194);
and AND4 (N637, N633, N326, N426, N510);
nor NOR4 (N638, N626, N220, N496, N49);
not NOT1 (N639, N634);
not NOT1 (N640, N607);
nor NOR4 (N641, N639, N560, N281, N416);
nor NOR2 (N642, N635, N140);
or OR2 (N643, N638, N39);
nor NOR3 (N644, N632, N72, N27);
and AND2 (N645, N643, N295);
and AND2 (N646, N629, N512);
buf BUF1 (N647, N644);
and AND4 (N648, N637, N477, N558, N172);
xor XOR2 (N649, N640, N109);
nor NOR3 (N650, N646, N575, N303);
nand NAND2 (N651, N648, N136);
nand NAND4 (N652, N627, N425, N142, N153);
nand NAND3 (N653, N641, N230, N28);
xor XOR2 (N654, N652, N171);
nor NOR2 (N655, N649, N125);
xor XOR2 (N656, N651, N48);
buf BUF1 (N657, N653);
xor XOR2 (N658, N642, N92);
buf BUF1 (N659, N636);
nand NAND3 (N660, N645, N584, N86);
not NOT1 (N661, N656);
or OR4 (N662, N659, N433, N368, N543);
nand NAND4 (N663, N650, N15, N572, N469);
and AND2 (N664, N661, N469);
xor XOR2 (N665, N658, N63);
buf BUF1 (N666, N663);
nand NAND4 (N667, N655, N429, N55, N32);
and AND4 (N668, N613, N58, N234, N107);
nand NAND2 (N669, N667, N230);
nor NOR3 (N670, N657, N534, N454);
or OR2 (N671, N660, N347);
xor XOR2 (N672, N669, N385);
nand NAND3 (N673, N670, N261, N231);
or OR2 (N674, N666, N624);
xor XOR2 (N675, N662, N351);
not NOT1 (N676, N675);
nor NOR2 (N677, N673, N431);
and AND3 (N678, N647, N390, N217);
and AND4 (N679, N664, N279, N381, N124);
and AND4 (N680, N665, N312, N514, N647);
xor XOR2 (N681, N654, N55);
buf BUF1 (N682, N679);
xor XOR2 (N683, N682, N451);
nand NAND4 (N684, N681, N476, N352, N347);
xor XOR2 (N685, N678, N298);
buf BUF1 (N686, N683);
xor XOR2 (N687, N668, N555);
nor NOR4 (N688, N687, N681, N87, N425);
not NOT1 (N689, N684);
xor XOR2 (N690, N674, N220);
not NOT1 (N691, N690);
xor XOR2 (N692, N688, N598);
nor NOR4 (N693, N685, N330, N562, N220);
nand NAND2 (N694, N677, N631);
or OR4 (N695, N694, N245, N100, N465);
nor NOR3 (N696, N686, N32, N332);
nand NAND2 (N697, N672, N357);
xor XOR2 (N698, N689, N526);
nor NOR2 (N699, N691, N211);
nand NAND2 (N700, N698, N37);
and AND4 (N701, N699, N267, N688, N415);
and AND2 (N702, N680, N6);
not NOT1 (N703, N702);
nand NAND4 (N704, N700, N7, N420, N79);
nor NOR3 (N705, N696, N145, N273);
and AND3 (N706, N701, N66, N2);
not NOT1 (N707, N693);
buf BUF1 (N708, N671);
and AND3 (N709, N703, N127, N15);
and AND3 (N710, N706, N310, N221);
buf BUF1 (N711, N695);
endmodule