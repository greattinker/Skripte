// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N795,N804,N805,N798,N809,N815,N785,N813,N796,N816;

and AND4 (N17, N15, N6, N11, N11);
nor NOR2 (N18, N15, N14);
not NOT1 (N19, N3);
or OR2 (N20, N1, N7);
or OR4 (N21, N12, N2, N10, N8);
or OR4 (N22, N9, N6, N10, N15);
nor NOR3 (N23, N20, N14, N8);
buf BUF1 (N24, N3);
and AND3 (N25, N10, N23, N1);
and AND3 (N26, N15, N20, N14);
nand NAND3 (N27, N11, N1, N24);
nand NAND3 (N28, N19, N13, N23);
nand NAND2 (N29, N19, N9);
xor XOR2 (N30, N27, N7);
or OR3 (N31, N5, N17, N27);
xor XOR2 (N32, N18, N25);
and AND2 (N33, N18, N26);
buf BUF1 (N34, N24);
or OR4 (N35, N21, N29, N2, N21);
and AND3 (N36, N9, N18, N22);
buf BUF1 (N37, N29);
not NOT1 (N38, N25);
or OR4 (N39, N38, N29, N37, N18);
xor XOR2 (N40, N22, N6);
not NOT1 (N41, N34);
buf BUF1 (N42, N41);
or OR3 (N43, N35, N37, N39);
or OR3 (N44, N25, N19, N19);
not NOT1 (N45, N43);
nor NOR4 (N46, N33, N35, N12, N38);
buf BUF1 (N47, N45);
xor XOR2 (N48, N47, N4);
and AND3 (N49, N40, N1, N35);
buf BUF1 (N50, N48);
nand NAND2 (N51, N46, N11);
and AND4 (N52, N31, N35, N34, N33);
buf BUF1 (N53, N36);
xor XOR2 (N54, N50, N28);
not NOT1 (N55, N16);
nor NOR4 (N56, N51, N5, N15, N33);
not NOT1 (N57, N55);
nor NOR3 (N58, N53, N47, N42);
buf BUF1 (N59, N58);
or OR2 (N60, N37, N19);
not NOT1 (N61, N44);
xor XOR2 (N62, N61, N47);
and AND2 (N63, N62, N41);
nor NOR3 (N64, N59, N25, N14);
nand NAND3 (N65, N56, N56, N37);
buf BUF1 (N66, N54);
xor XOR2 (N67, N57, N44);
and AND4 (N68, N63, N56, N4, N60);
nand NAND2 (N69, N34, N16);
nor NOR4 (N70, N64, N61, N36, N29);
buf BUF1 (N71, N65);
xor XOR2 (N72, N71, N64);
and AND3 (N73, N70, N65, N51);
and AND4 (N74, N30, N35, N10, N47);
nand NAND2 (N75, N73, N63);
not NOT1 (N76, N52);
buf BUF1 (N77, N72);
not NOT1 (N78, N77);
nor NOR2 (N79, N66, N35);
nor NOR3 (N80, N75, N67, N64);
not NOT1 (N81, N61);
nor NOR2 (N82, N49, N62);
and AND2 (N83, N68, N76);
buf BUF1 (N84, N82);
and AND4 (N85, N80, N64, N21, N29);
nand NAND4 (N86, N41, N10, N34, N65);
buf BUF1 (N87, N78);
not NOT1 (N88, N69);
not NOT1 (N89, N85);
not NOT1 (N90, N74);
and AND4 (N91, N86, N70, N50, N53);
not NOT1 (N92, N91);
not NOT1 (N93, N89);
xor XOR2 (N94, N87, N62);
xor XOR2 (N95, N83, N78);
buf BUF1 (N96, N90);
buf BUF1 (N97, N84);
buf BUF1 (N98, N96);
buf BUF1 (N99, N32);
nor NOR3 (N100, N95, N26, N96);
not NOT1 (N101, N98);
not NOT1 (N102, N97);
xor XOR2 (N103, N94, N80);
xor XOR2 (N104, N81, N47);
buf BUF1 (N105, N104);
nor NOR2 (N106, N101, N65);
or OR3 (N107, N79, N78, N74);
nand NAND3 (N108, N105, N49, N45);
not NOT1 (N109, N103);
nand NAND3 (N110, N102, N103, N26);
and AND3 (N111, N110, N102, N99);
buf BUF1 (N112, N111);
nor NOR4 (N113, N35, N93, N52, N37);
buf BUF1 (N114, N26);
nand NAND2 (N115, N92, N36);
not NOT1 (N116, N108);
not NOT1 (N117, N116);
nor NOR2 (N118, N113, N50);
xor XOR2 (N119, N115, N103);
buf BUF1 (N120, N112);
nand NAND2 (N121, N100, N59);
xor XOR2 (N122, N118, N26);
or OR3 (N123, N114, N82, N108);
nor NOR4 (N124, N120, N100, N51, N4);
not NOT1 (N125, N106);
nor NOR4 (N126, N107, N72, N117, N118);
nand NAND2 (N127, N93, N15);
and AND2 (N128, N123, N18);
nand NAND3 (N129, N124, N95, N65);
buf BUF1 (N130, N119);
or OR4 (N131, N109, N27, N67, N86);
nand NAND3 (N132, N126, N16, N81);
nor NOR4 (N133, N125, N129, N75, N7);
buf BUF1 (N134, N96);
not NOT1 (N135, N133);
buf BUF1 (N136, N134);
and AND4 (N137, N131, N69, N132, N92);
nor NOR3 (N138, N28, N94, N43);
nor NOR2 (N139, N136, N40);
nand NAND2 (N140, N130, N115);
and AND3 (N141, N135, N23, N130);
or OR3 (N142, N140, N127, N53);
nand NAND4 (N143, N103, N48, N98, N47);
or OR3 (N144, N143, N100, N4);
or OR3 (N145, N137, N129, N58);
and AND2 (N146, N139, N69);
not NOT1 (N147, N145);
buf BUF1 (N148, N121);
xor XOR2 (N149, N128, N134);
nor NOR3 (N150, N138, N27, N17);
xor XOR2 (N151, N88, N1);
nand NAND4 (N152, N150, N115, N79, N24);
nor NOR3 (N153, N141, N143, N135);
and AND4 (N154, N153, N59, N62, N51);
xor XOR2 (N155, N149, N27);
and AND4 (N156, N147, N75, N15, N1);
nor NOR3 (N157, N146, N95, N136);
xor XOR2 (N158, N156, N117);
nand NAND2 (N159, N155, N31);
nor NOR4 (N160, N148, N88, N85, N134);
xor XOR2 (N161, N152, N49);
not NOT1 (N162, N144);
not NOT1 (N163, N158);
nor NOR4 (N164, N122, N100, N3, N120);
and AND2 (N165, N142, N6);
and AND4 (N166, N154, N157, N138, N75);
buf BUF1 (N167, N73);
nor NOR2 (N168, N161, N46);
and AND4 (N169, N167, N96, N21, N58);
nor NOR4 (N170, N169, N138, N26, N88);
nor NOR4 (N171, N165, N136, N138, N164);
nor NOR2 (N172, N7, N34);
xor XOR2 (N173, N170, N146);
xor XOR2 (N174, N151, N163);
or OR4 (N175, N69, N172, N146, N123);
buf BUF1 (N176, N169);
buf BUF1 (N177, N176);
or OR2 (N178, N162, N109);
or OR2 (N179, N174, N51);
not NOT1 (N180, N171);
nor NOR4 (N181, N177, N138, N42, N170);
nand NAND4 (N182, N159, N157, N38, N134);
not NOT1 (N183, N178);
not NOT1 (N184, N179);
and AND2 (N185, N180, N87);
nor NOR3 (N186, N185, N33, N183);
buf BUF1 (N187, N90);
or OR3 (N188, N184, N81, N94);
nor NOR2 (N189, N188, N182);
or OR2 (N190, N181, N76);
nand NAND3 (N191, N117, N151, N31);
nor NOR4 (N192, N160, N188, N164, N38);
buf BUF1 (N193, N192);
and AND3 (N194, N175, N84, N132);
nor NOR3 (N195, N189, N102, N32);
or OR3 (N196, N186, N174, N185);
and AND4 (N197, N173, N66, N181, N53);
and AND3 (N198, N190, N17, N85);
and AND4 (N199, N198, N39, N36, N192);
and AND4 (N200, N196, N54, N196, N94);
or OR3 (N201, N191, N162, N72);
nand NAND3 (N202, N168, N62, N130);
nand NAND3 (N203, N166, N87, N190);
xor XOR2 (N204, N202, N21);
not NOT1 (N205, N197);
buf BUF1 (N206, N203);
and AND3 (N207, N201, N172, N70);
buf BUF1 (N208, N205);
nand NAND3 (N209, N194, N205, N66);
or OR4 (N210, N204, N136, N48, N84);
buf BUF1 (N211, N209);
nand NAND2 (N212, N193, N176);
not NOT1 (N213, N195);
not NOT1 (N214, N206);
and AND4 (N215, N207, N155, N190, N26);
not NOT1 (N216, N214);
xor XOR2 (N217, N210, N167);
nand NAND2 (N218, N213, N110);
buf BUF1 (N219, N187);
or OR2 (N220, N212, N176);
nand NAND3 (N221, N219, N130, N106);
or OR4 (N222, N217, N153, N55, N20);
not NOT1 (N223, N222);
or OR4 (N224, N223, N82, N21, N12);
buf BUF1 (N225, N224);
not NOT1 (N226, N200);
not NOT1 (N227, N208);
nand NAND2 (N228, N220, N207);
nor NOR2 (N229, N226, N5);
xor XOR2 (N230, N218, N114);
and AND2 (N231, N227, N223);
not NOT1 (N232, N230);
buf BUF1 (N233, N211);
buf BUF1 (N234, N229);
buf BUF1 (N235, N228);
nand NAND4 (N236, N199, N139, N34, N191);
and AND3 (N237, N215, N213, N135);
nor NOR2 (N238, N232, N3);
and AND3 (N239, N225, N84, N18);
not NOT1 (N240, N237);
buf BUF1 (N241, N236);
not NOT1 (N242, N235);
or OR4 (N243, N240, N55, N141, N182);
nor NOR2 (N244, N238, N41);
buf BUF1 (N245, N242);
not NOT1 (N246, N239);
and AND4 (N247, N234, N99, N192, N85);
buf BUF1 (N248, N246);
not NOT1 (N249, N241);
buf BUF1 (N250, N248);
or OR2 (N251, N231, N15);
not NOT1 (N252, N233);
or OR4 (N253, N250, N82, N215, N238);
and AND3 (N254, N216, N124, N66);
nor NOR4 (N255, N244, N232, N234, N125);
xor XOR2 (N256, N221, N242);
and AND3 (N257, N243, N174, N147);
and AND2 (N258, N247, N50);
and AND4 (N259, N255, N213, N202, N121);
and AND3 (N260, N256, N86, N163);
nor NOR2 (N261, N249, N160);
or OR3 (N262, N245, N7, N16);
not NOT1 (N263, N251);
nand NAND3 (N264, N263, N203, N48);
not NOT1 (N265, N264);
not NOT1 (N266, N252);
and AND2 (N267, N262, N8);
buf BUF1 (N268, N267);
or OR2 (N269, N265, N88);
nor NOR2 (N270, N254, N222);
xor XOR2 (N271, N266, N48);
xor XOR2 (N272, N269, N226);
or OR4 (N273, N258, N267, N5, N89);
not NOT1 (N274, N273);
xor XOR2 (N275, N257, N144);
or OR2 (N276, N259, N262);
buf BUF1 (N277, N274);
xor XOR2 (N278, N276, N235);
not NOT1 (N279, N278);
buf BUF1 (N280, N272);
nand NAND4 (N281, N260, N193, N191, N89);
or OR2 (N282, N271, N125);
nor NOR3 (N283, N280, N67, N212);
not NOT1 (N284, N283);
not NOT1 (N285, N284);
not NOT1 (N286, N281);
xor XOR2 (N287, N261, N177);
and AND3 (N288, N285, N36, N20);
nor NOR2 (N289, N275, N288);
and AND3 (N290, N263, N116, N65);
or OR3 (N291, N282, N270, N205);
xor XOR2 (N292, N195, N241);
xor XOR2 (N293, N279, N49);
buf BUF1 (N294, N286);
buf BUF1 (N295, N268);
buf BUF1 (N296, N289);
not NOT1 (N297, N287);
buf BUF1 (N298, N296);
not NOT1 (N299, N292);
and AND4 (N300, N298, N102, N26, N162);
not NOT1 (N301, N295);
buf BUF1 (N302, N277);
or OR2 (N303, N290, N100);
not NOT1 (N304, N253);
and AND4 (N305, N303, N183, N285, N218);
and AND2 (N306, N299, N191);
xor XOR2 (N307, N293, N84);
nor NOR2 (N308, N291, N216);
xor XOR2 (N309, N304, N7);
and AND4 (N310, N300, N309, N118, N180);
and AND3 (N311, N275, N15, N46);
xor XOR2 (N312, N305, N193);
not NOT1 (N313, N302);
not NOT1 (N314, N312);
nand NAND4 (N315, N313, N266, N114, N204);
nand NAND2 (N316, N308, N142);
not NOT1 (N317, N311);
buf BUF1 (N318, N315);
buf BUF1 (N319, N314);
buf BUF1 (N320, N319);
not NOT1 (N321, N318);
not NOT1 (N322, N307);
not NOT1 (N323, N316);
buf BUF1 (N324, N306);
and AND2 (N325, N317, N200);
buf BUF1 (N326, N323);
not NOT1 (N327, N301);
buf BUF1 (N328, N326);
nand NAND3 (N329, N328, N27, N311);
or OR3 (N330, N325, N269, N82);
and AND2 (N331, N321, N16);
nand NAND2 (N332, N330, N297);
or OR2 (N333, N196, N322);
nand NAND4 (N334, N281, N178, N127, N144);
nor NOR4 (N335, N327, N121, N193, N319);
xor XOR2 (N336, N332, N111);
and AND2 (N337, N335, N230);
nand NAND2 (N338, N336, N214);
xor XOR2 (N339, N333, N195);
xor XOR2 (N340, N310, N231);
not NOT1 (N341, N337);
xor XOR2 (N342, N331, N338);
nor NOR2 (N343, N45, N122);
buf BUF1 (N344, N342);
and AND3 (N345, N344, N151, N178);
xor XOR2 (N346, N334, N319);
nand NAND2 (N347, N324, N327);
nand NAND4 (N348, N320, N259, N113, N109);
buf BUF1 (N349, N346);
not NOT1 (N350, N347);
and AND3 (N351, N341, N259, N175);
nor NOR4 (N352, N349, N273, N12, N268);
nand NAND4 (N353, N343, N219, N69, N89);
nor NOR3 (N354, N294, N85, N307);
nor NOR3 (N355, N350, N181, N243);
xor XOR2 (N356, N345, N294);
xor XOR2 (N357, N339, N224);
or OR2 (N358, N329, N100);
nand NAND2 (N359, N355, N2);
and AND2 (N360, N340, N354);
nand NAND3 (N361, N104, N174, N93);
buf BUF1 (N362, N358);
nor NOR3 (N363, N361, N53, N153);
xor XOR2 (N364, N348, N63);
not NOT1 (N365, N363);
nor NOR2 (N366, N356, N9);
and AND3 (N367, N365, N163, N80);
not NOT1 (N368, N364);
not NOT1 (N369, N368);
not NOT1 (N370, N351);
not NOT1 (N371, N352);
or OR2 (N372, N357, N298);
or OR2 (N373, N369, N207);
nor NOR3 (N374, N373, N66, N217);
nor NOR4 (N375, N370, N103, N337, N198);
nand NAND4 (N376, N375, N346, N74, N147);
and AND3 (N377, N374, N155, N149);
nand NAND2 (N378, N367, N322);
not NOT1 (N379, N362);
nor NOR3 (N380, N360, N81, N256);
nand NAND4 (N381, N378, N115, N327, N87);
nor NOR3 (N382, N359, N99, N99);
and AND3 (N383, N380, N187, N240);
not NOT1 (N384, N377);
buf BUF1 (N385, N382);
buf BUF1 (N386, N376);
nor NOR4 (N387, N386, N317, N48, N313);
and AND4 (N388, N383, N100, N86, N227);
nand NAND3 (N389, N385, N181, N309);
nand NAND2 (N390, N379, N169);
nand NAND4 (N391, N390, N319, N116, N244);
nor NOR2 (N392, N387, N40);
nand NAND2 (N393, N391, N140);
nor NOR2 (N394, N353, N264);
not NOT1 (N395, N388);
buf BUF1 (N396, N384);
nand NAND3 (N397, N389, N20, N138);
buf BUF1 (N398, N381);
nand NAND3 (N399, N393, N51, N292);
xor XOR2 (N400, N399, N339);
nor NOR2 (N401, N398, N82);
not NOT1 (N402, N396);
or OR3 (N403, N394, N172, N350);
not NOT1 (N404, N372);
or OR4 (N405, N404, N164, N33, N112);
nand NAND3 (N406, N401, N360, N197);
not NOT1 (N407, N395);
nor NOR3 (N408, N397, N399, N285);
nor NOR4 (N409, N408, N167, N28, N162);
buf BUF1 (N410, N407);
and AND2 (N411, N392, N263);
or OR4 (N412, N400, N132, N250, N243);
xor XOR2 (N413, N412, N88);
nand NAND3 (N414, N403, N383, N137);
xor XOR2 (N415, N411, N295);
or OR2 (N416, N410, N9);
nand NAND4 (N417, N414, N416, N140, N307);
and AND4 (N418, N197, N100, N17, N211);
or OR4 (N419, N413, N398, N200, N96);
buf BUF1 (N420, N417);
and AND4 (N421, N406, N276, N416, N36);
nand NAND4 (N422, N366, N20, N298, N336);
buf BUF1 (N423, N422);
or OR3 (N424, N409, N160, N29);
buf BUF1 (N425, N415);
and AND2 (N426, N423, N352);
and AND4 (N427, N418, N338, N111, N245);
not NOT1 (N428, N426);
not NOT1 (N429, N419);
xor XOR2 (N430, N425, N280);
xor XOR2 (N431, N430, N415);
nand NAND4 (N432, N405, N254, N195, N253);
xor XOR2 (N433, N429, N195);
or OR2 (N434, N402, N4);
and AND4 (N435, N371, N353, N312, N341);
xor XOR2 (N436, N420, N127);
not NOT1 (N437, N421);
xor XOR2 (N438, N424, N398);
nand NAND2 (N439, N434, N98);
xor XOR2 (N440, N428, N193);
or OR2 (N441, N431, N225);
and AND3 (N442, N439, N327, N32);
not NOT1 (N443, N438);
nor NOR2 (N444, N440, N84);
and AND2 (N445, N441, N125);
not NOT1 (N446, N445);
not NOT1 (N447, N444);
nand NAND3 (N448, N432, N110, N237);
and AND3 (N449, N436, N306, N362);
and AND3 (N450, N427, N363, N172);
or OR3 (N451, N443, N368, N175);
and AND4 (N452, N435, N204, N93, N78);
nor NOR2 (N453, N446, N389);
or OR4 (N454, N447, N289, N443, N401);
or OR2 (N455, N449, N346);
not NOT1 (N456, N448);
nor NOR4 (N457, N452, N294, N86, N142);
nand NAND2 (N458, N437, N67);
xor XOR2 (N459, N451, N199);
nor NOR2 (N460, N433, N301);
and AND4 (N461, N454, N225, N20, N449);
or OR4 (N462, N455, N345, N430, N311);
not NOT1 (N463, N459);
or OR3 (N464, N461, N103, N72);
nor NOR2 (N465, N457, N144);
buf BUF1 (N466, N450);
and AND4 (N467, N458, N102, N299, N156);
buf BUF1 (N468, N463);
not NOT1 (N469, N468);
or OR2 (N470, N466, N78);
and AND2 (N471, N464, N393);
not NOT1 (N472, N469);
not NOT1 (N473, N472);
and AND4 (N474, N471, N231, N347, N149);
and AND3 (N475, N453, N75, N117);
nand NAND2 (N476, N460, N168);
xor XOR2 (N477, N456, N95);
buf BUF1 (N478, N473);
nand NAND4 (N479, N477, N109, N45, N43);
xor XOR2 (N480, N475, N133);
xor XOR2 (N481, N442, N84);
buf BUF1 (N482, N478);
or OR2 (N483, N470, N402);
and AND4 (N484, N474, N140, N275, N376);
nor NOR4 (N485, N484, N426, N261, N219);
nor NOR3 (N486, N462, N441, N298);
and AND4 (N487, N482, N181, N352, N409);
not NOT1 (N488, N487);
not NOT1 (N489, N488);
and AND3 (N490, N465, N469, N272);
not NOT1 (N491, N483);
and AND3 (N492, N489, N457, N384);
and AND4 (N493, N491, N82, N147, N265);
or OR4 (N494, N485, N72, N169, N344);
nor NOR2 (N495, N476, N258);
xor XOR2 (N496, N479, N317);
buf BUF1 (N497, N481);
nand NAND2 (N498, N480, N169);
or OR2 (N499, N495, N433);
xor XOR2 (N500, N499, N245);
nand NAND3 (N501, N496, N500, N37);
not NOT1 (N502, N132);
or OR3 (N503, N493, N402, N340);
buf BUF1 (N504, N502);
nand NAND2 (N505, N490, N79);
nor NOR2 (N506, N498, N462);
not NOT1 (N507, N506);
and AND2 (N508, N497, N25);
xor XOR2 (N509, N503, N336);
buf BUF1 (N510, N492);
nand NAND4 (N511, N501, N79, N124, N159);
or OR4 (N512, N507, N260, N480, N252);
nand NAND2 (N513, N509, N121);
or OR4 (N514, N510, N297, N235, N170);
nand NAND3 (N515, N513, N430, N108);
and AND4 (N516, N511, N172, N350, N294);
or OR2 (N517, N516, N382);
not NOT1 (N518, N517);
not NOT1 (N519, N486);
buf BUF1 (N520, N518);
nand NAND4 (N521, N504, N463, N392, N119);
buf BUF1 (N522, N514);
not NOT1 (N523, N467);
or OR3 (N524, N522, N3, N364);
nand NAND4 (N525, N521, N137, N189, N71);
nor NOR2 (N526, N515, N167);
not NOT1 (N527, N525);
or OR3 (N528, N523, N47, N357);
buf BUF1 (N529, N519);
and AND4 (N530, N508, N124, N40, N502);
nand NAND2 (N531, N527, N125);
nand NAND4 (N532, N531, N378, N253, N429);
or OR3 (N533, N530, N71, N453);
and AND2 (N534, N505, N220);
nand NAND3 (N535, N529, N408, N182);
and AND4 (N536, N512, N37, N90, N454);
nor NOR4 (N537, N528, N442, N88, N217);
nand NAND2 (N538, N534, N220);
or OR4 (N539, N532, N75, N448, N119);
or OR4 (N540, N494, N474, N296, N482);
xor XOR2 (N541, N533, N352);
nand NAND4 (N542, N524, N457, N232, N126);
xor XOR2 (N543, N535, N209);
xor XOR2 (N544, N543, N364);
xor XOR2 (N545, N536, N115);
buf BUF1 (N546, N544);
nand NAND3 (N547, N540, N145, N375);
nand NAND2 (N548, N539, N509);
or OR2 (N549, N545, N83);
and AND3 (N550, N538, N474, N535);
nand NAND3 (N551, N520, N38, N525);
not NOT1 (N552, N537);
nor NOR2 (N553, N548, N503);
and AND3 (N554, N547, N150, N545);
nand NAND4 (N555, N551, N127, N518, N177);
nand NAND2 (N556, N549, N548);
nor NOR2 (N557, N554, N490);
buf BUF1 (N558, N541);
buf BUF1 (N559, N557);
xor XOR2 (N560, N546, N204);
or OR3 (N561, N553, N278, N544);
nand NAND3 (N562, N542, N168, N465);
nor NOR4 (N563, N562, N36, N468, N110);
and AND4 (N564, N561, N126, N169, N506);
and AND4 (N565, N555, N259, N8, N66);
or OR2 (N566, N564, N243);
not NOT1 (N567, N550);
not NOT1 (N568, N556);
nand NAND4 (N569, N552, N5, N63, N321);
or OR2 (N570, N526, N321);
xor XOR2 (N571, N558, N43);
xor XOR2 (N572, N570, N254);
not NOT1 (N573, N566);
not NOT1 (N574, N563);
buf BUF1 (N575, N571);
nand NAND4 (N576, N559, N543, N122, N444);
nor NOR2 (N577, N572, N203);
and AND3 (N578, N560, N122, N291);
and AND2 (N579, N575, N571);
and AND4 (N580, N574, N478, N565, N224);
nand NAND3 (N581, N387, N438, N186);
xor XOR2 (N582, N580, N153);
or OR4 (N583, N579, N406, N122, N574);
not NOT1 (N584, N573);
nor NOR3 (N585, N583, N228, N143);
buf BUF1 (N586, N581);
and AND4 (N587, N567, N494, N486, N468);
nand NAND3 (N588, N585, N293, N278);
and AND2 (N589, N584, N169);
and AND2 (N590, N568, N571);
xor XOR2 (N591, N589, N194);
buf BUF1 (N592, N588);
buf BUF1 (N593, N591);
and AND4 (N594, N590, N592, N533, N559);
and AND3 (N595, N146, N350, N475);
xor XOR2 (N596, N586, N422);
buf BUF1 (N597, N569);
or OR3 (N598, N594, N55, N550);
or OR3 (N599, N595, N111, N495);
and AND3 (N600, N576, N514, N474);
nand NAND4 (N601, N598, N518, N411, N235);
nand NAND2 (N602, N582, N68);
or OR2 (N603, N587, N145);
not NOT1 (N604, N600);
buf BUF1 (N605, N599);
nand NAND3 (N606, N601, N505, N274);
not NOT1 (N607, N602);
nand NAND4 (N608, N596, N523, N375, N331);
not NOT1 (N609, N608);
xor XOR2 (N610, N605, N105);
xor XOR2 (N611, N610, N226);
xor XOR2 (N612, N577, N391);
xor XOR2 (N613, N609, N296);
nor NOR4 (N614, N613, N228, N38, N41);
nor NOR2 (N615, N578, N139);
not NOT1 (N616, N612);
buf BUF1 (N617, N616);
nand NAND4 (N618, N611, N289, N236, N315);
not NOT1 (N619, N614);
buf BUF1 (N620, N603);
nand NAND4 (N621, N615, N213, N619, N116);
nand NAND4 (N622, N10, N431, N256, N547);
xor XOR2 (N623, N607, N225);
and AND4 (N624, N622, N176, N92, N490);
xor XOR2 (N625, N593, N119);
not NOT1 (N626, N620);
or OR2 (N627, N618, N272);
xor XOR2 (N628, N621, N607);
and AND4 (N629, N624, N9, N272, N4);
buf BUF1 (N630, N627);
and AND2 (N631, N630, N571);
or OR4 (N632, N628, N229, N33, N88);
not NOT1 (N633, N625);
buf BUF1 (N634, N617);
not NOT1 (N635, N606);
not NOT1 (N636, N604);
not NOT1 (N637, N633);
not NOT1 (N638, N631);
xor XOR2 (N639, N635, N435);
or OR2 (N640, N629, N635);
xor XOR2 (N641, N638, N36);
nand NAND3 (N642, N634, N501, N47);
buf BUF1 (N643, N626);
not NOT1 (N644, N623);
nand NAND2 (N645, N644, N580);
not NOT1 (N646, N636);
nor NOR3 (N647, N643, N225, N633);
xor XOR2 (N648, N641, N421);
nand NAND3 (N649, N642, N70, N278);
and AND4 (N650, N640, N448, N562, N354);
and AND4 (N651, N639, N56, N319, N540);
xor XOR2 (N652, N648, N238);
nand NAND3 (N653, N645, N350, N205);
not NOT1 (N654, N647);
or OR3 (N655, N653, N57, N596);
and AND2 (N656, N649, N130);
nand NAND2 (N657, N655, N290);
or OR4 (N658, N657, N368, N428, N436);
not NOT1 (N659, N652);
not NOT1 (N660, N637);
buf BUF1 (N661, N650);
and AND4 (N662, N654, N481, N380, N645);
nand NAND3 (N663, N658, N404, N310);
xor XOR2 (N664, N646, N498);
buf BUF1 (N665, N664);
buf BUF1 (N666, N660);
and AND4 (N667, N656, N485, N276, N274);
and AND3 (N668, N665, N353, N47);
and AND3 (N669, N663, N394, N629);
and AND3 (N670, N667, N659, N70);
buf BUF1 (N671, N63);
nand NAND3 (N672, N597, N39, N301);
not NOT1 (N673, N670);
nand NAND3 (N674, N632, N491, N488);
nand NAND3 (N675, N669, N638, N237);
and AND3 (N676, N651, N620, N202);
or OR3 (N677, N661, N4, N351);
nor NOR2 (N678, N674, N152);
nand NAND3 (N679, N668, N605, N48);
nand NAND4 (N680, N677, N399, N393, N618);
xor XOR2 (N681, N666, N257);
xor XOR2 (N682, N673, N487);
nand NAND3 (N683, N672, N589, N576);
nand NAND4 (N684, N676, N656, N276, N606);
and AND2 (N685, N678, N284);
buf BUF1 (N686, N685);
xor XOR2 (N687, N682, N402);
nor NOR3 (N688, N684, N199, N372);
and AND3 (N689, N671, N422, N46);
or OR3 (N690, N687, N107, N9);
not NOT1 (N691, N690);
xor XOR2 (N692, N680, N301);
or OR4 (N693, N686, N250, N40, N117);
nor NOR3 (N694, N679, N148, N416);
xor XOR2 (N695, N689, N233);
and AND2 (N696, N675, N338);
and AND3 (N697, N694, N252, N269);
buf BUF1 (N698, N688);
not NOT1 (N699, N693);
or OR3 (N700, N692, N601, N360);
xor XOR2 (N701, N697, N322);
nor NOR3 (N702, N695, N511, N387);
and AND4 (N703, N681, N303, N372, N517);
nor NOR2 (N704, N699, N517);
and AND4 (N705, N691, N280, N217, N512);
xor XOR2 (N706, N698, N121);
xor XOR2 (N707, N683, N231);
not NOT1 (N708, N702);
and AND4 (N709, N696, N578, N527, N707);
buf BUF1 (N710, N2);
nand NAND3 (N711, N703, N619, N423);
xor XOR2 (N712, N701, N59);
buf BUF1 (N713, N712);
buf BUF1 (N714, N710);
or OR2 (N715, N704, N681);
not NOT1 (N716, N708);
and AND2 (N717, N713, N180);
and AND3 (N718, N706, N635, N225);
not NOT1 (N719, N705);
or OR4 (N720, N662, N116, N585, N671);
buf BUF1 (N721, N714);
not NOT1 (N722, N719);
or OR4 (N723, N700, N37, N395, N405);
or OR2 (N724, N711, N652);
nor NOR2 (N725, N715, N141);
not NOT1 (N726, N718);
nor NOR4 (N727, N726, N95, N324, N302);
and AND3 (N728, N727, N530, N574);
and AND4 (N729, N725, N646, N674, N690);
nor NOR3 (N730, N723, N180, N211);
nand NAND3 (N731, N722, N408, N571);
and AND2 (N732, N731, N261);
nand NAND4 (N733, N716, N350, N645, N25);
nand NAND2 (N734, N720, N109);
buf BUF1 (N735, N733);
not NOT1 (N736, N721);
nor NOR4 (N737, N730, N445, N544, N49);
nand NAND3 (N738, N735, N467, N406);
or OR2 (N739, N738, N135);
not NOT1 (N740, N734);
buf BUF1 (N741, N717);
buf BUF1 (N742, N724);
not NOT1 (N743, N742);
nand NAND4 (N744, N709, N107, N181, N515);
buf BUF1 (N745, N732);
nand NAND4 (N746, N745, N185, N588, N180);
and AND3 (N747, N741, N394, N345);
and AND3 (N748, N747, N83, N170);
nor NOR3 (N749, N739, N159, N180);
buf BUF1 (N750, N737);
nor NOR4 (N751, N729, N288, N552, N491);
not NOT1 (N752, N740);
nor NOR2 (N753, N751, N551);
nor NOR2 (N754, N728, N597);
or OR4 (N755, N744, N492, N208, N712);
xor XOR2 (N756, N746, N510);
and AND2 (N757, N736, N654);
and AND3 (N758, N748, N528, N459);
xor XOR2 (N759, N752, N618);
or OR4 (N760, N755, N385, N559, N374);
nor NOR2 (N761, N750, N315);
and AND2 (N762, N754, N624);
not NOT1 (N763, N743);
nor NOR2 (N764, N759, N174);
xor XOR2 (N765, N757, N453);
or OR4 (N766, N764, N417, N219, N564);
or OR4 (N767, N749, N432, N422, N57);
xor XOR2 (N768, N761, N81);
nand NAND2 (N769, N765, N642);
and AND2 (N770, N767, N312);
buf BUF1 (N771, N770);
not NOT1 (N772, N762);
nor NOR3 (N773, N772, N763, N584);
xor XOR2 (N774, N216, N600);
nor NOR3 (N775, N771, N350, N219);
xor XOR2 (N776, N775, N417);
nor NOR2 (N777, N766, N516);
or OR4 (N778, N769, N733, N556, N166);
or OR4 (N779, N773, N188, N139, N296);
buf BUF1 (N780, N774);
nor NOR4 (N781, N776, N205, N42, N140);
buf BUF1 (N782, N760);
nand NAND4 (N783, N753, N111, N455, N684);
not NOT1 (N784, N780);
and AND4 (N785, N758, N686, N467, N218);
or OR4 (N786, N783, N701, N648, N753);
and AND3 (N787, N779, N221, N478);
not NOT1 (N788, N781);
xor XOR2 (N789, N782, N118);
buf BUF1 (N790, N786);
xor XOR2 (N791, N788, N725);
nand NAND3 (N792, N787, N236, N721);
nor NOR4 (N793, N756, N268, N456, N731);
xor XOR2 (N794, N790, N222);
buf BUF1 (N795, N793);
not NOT1 (N796, N792);
nor NOR4 (N797, N784, N778, N338, N330);
and AND2 (N798, N430, N20);
not NOT1 (N799, N789);
and AND3 (N800, N791, N65, N415);
nor NOR3 (N801, N768, N750, N294);
buf BUF1 (N802, N799);
nor NOR3 (N803, N797, N48, N123);
or OR3 (N804, N802, N590, N472);
xor XOR2 (N805, N777, N323);
or OR2 (N806, N801, N41);
buf BUF1 (N807, N803);
and AND2 (N808, N806, N578);
and AND4 (N809, N807, N279, N218, N68);
or OR3 (N810, N808, N122, N732);
buf BUF1 (N811, N794);
nor NOR2 (N812, N810, N222);
nor NOR3 (N813, N811, N230, N741);
nand NAND3 (N814, N812, N378, N661);
xor XOR2 (N815, N800, N390);
nand NAND3 (N816, N814, N358, N226);
endmodule