// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N1490,N1505,N1503,N1506,N1495,N1494,N1509,N1501,N1508,N1510;

and AND2 (N11, N1, N4);
and AND4 (N12, N11, N10, N3, N3);
xor XOR2 (N13, N9, N4);
or OR4 (N14, N1, N11, N12, N13);
and AND4 (N15, N14, N5, N13, N6);
nor NOR3 (N16, N15, N1, N6);
nor NOR4 (N17, N2, N4, N5, N12);
nor NOR3 (N18, N4, N14, N10);
nor NOR2 (N19, N2, N8);
nand NAND2 (N20, N2, N8);
xor XOR2 (N21, N1, N7);
not NOT1 (N22, N9);
and AND4 (N23, N2, N19, N18, N12);
or OR2 (N24, N9, N20);
buf BUF1 (N25, N7);
nor NOR4 (N26, N17, N16, N22, N9);
xor XOR2 (N27, N21, N23);
nor NOR3 (N28, N21, N12, N17);
or OR2 (N29, N9, N19);
and AND3 (N30, N7, N18, N17);
xor XOR2 (N31, N1, N13);
nand NAND2 (N32, N12, N14);
xor XOR2 (N33, N13, N14);
nand NAND2 (N34, N30, N16);
xor XOR2 (N35, N31, N20);
and AND3 (N36, N24, N31, N14);
buf BUF1 (N37, N29);
nor NOR3 (N38, N26, N25, N6);
not NOT1 (N39, N6);
or OR2 (N40, N28, N20);
xor XOR2 (N41, N38, N31);
or OR3 (N42, N41, N5, N34);
not NOT1 (N43, N9);
xor XOR2 (N44, N43, N6);
or OR2 (N45, N27, N25);
nor NOR3 (N46, N37, N45, N15);
buf BUF1 (N47, N42);
not NOT1 (N48, N10);
buf BUF1 (N49, N46);
xor XOR2 (N50, N35, N29);
nand NAND4 (N51, N36, N7, N14, N27);
buf BUF1 (N52, N32);
not NOT1 (N53, N44);
nor NOR3 (N54, N53, N37, N8);
nor NOR4 (N55, N40, N10, N8, N11);
or OR2 (N56, N48, N25);
or OR3 (N57, N55, N27, N46);
or OR3 (N58, N51, N13, N37);
or OR4 (N59, N56, N21, N51, N24);
buf BUF1 (N60, N58);
nor NOR2 (N61, N59, N7);
buf BUF1 (N62, N61);
not NOT1 (N63, N39);
and AND2 (N64, N57, N14);
nand NAND3 (N65, N54, N2, N14);
nand NAND4 (N66, N62, N61, N12, N6);
not NOT1 (N67, N47);
xor XOR2 (N68, N33, N4);
xor XOR2 (N69, N60, N53);
buf BUF1 (N70, N66);
not NOT1 (N71, N68);
not NOT1 (N72, N50);
and AND3 (N73, N64, N50, N13);
nor NOR2 (N74, N70, N49);
nand NAND2 (N75, N44, N61);
nand NAND3 (N76, N65, N66, N16);
buf BUF1 (N77, N63);
nor NOR2 (N78, N77, N69);
and AND2 (N79, N37, N22);
nor NOR2 (N80, N75, N52);
buf BUF1 (N81, N57);
and AND3 (N82, N74, N7, N62);
or OR3 (N83, N82, N74, N77);
xor XOR2 (N84, N79, N41);
nand NAND3 (N85, N67, N5, N23);
nor NOR2 (N86, N84, N53);
and AND4 (N87, N71, N64, N4, N56);
not NOT1 (N88, N78);
not NOT1 (N89, N81);
xor XOR2 (N90, N73, N32);
nand NAND3 (N91, N85, N37, N62);
xor XOR2 (N92, N80, N70);
buf BUF1 (N93, N72);
not NOT1 (N94, N88);
or OR3 (N95, N83, N49, N48);
nor NOR3 (N96, N86, N32, N95);
nand NAND4 (N97, N2, N10, N34, N20);
nand NAND4 (N98, N92, N42, N47, N47);
xor XOR2 (N99, N91, N7);
nand NAND2 (N100, N94, N44);
nor NOR3 (N101, N93, N10, N68);
nand NAND2 (N102, N97, N17);
xor XOR2 (N103, N96, N25);
or OR4 (N104, N87, N58, N75, N1);
nand NAND4 (N105, N99, N56, N36, N57);
nand NAND3 (N106, N89, N72, N101);
xor XOR2 (N107, N30, N101);
or OR3 (N108, N100, N13, N27);
and AND3 (N109, N98, N83, N75);
and AND4 (N110, N109, N44, N19, N87);
nand NAND2 (N111, N102, N57);
nand NAND4 (N112, N111, N102, N76, N109);
buf BUF1 (N113, N82);
and AND3 (N114, N107, N17, N105);
nor NOR4 (N115, N99, N104, N99, N32);
and AND4 (N116, N95, N9, N99, N110);
nor NOR3 (N117, N52, N42, N102);
xor XOR2 (N118, N117, N25);
or OR2 (N119, N106, N40);
nor NOR4 (N120, N119, N76, N22, N21);
nor NOR2 (N121, N90, N86);
nor NOR3 (N122, N115, N64, N16);
not NOT1 (N123, N113);
not NOT1 (N124, N121);
and AND2 (N125, N114, N107);
buf BUF1 (N126, N123);
nor NOR3 (N127, N120, N100, N70);
not NOT1 (N128, N122);
buf BUF1 (N129, N128);
not NOT1 (N130, N129);
xor XOR2 (N131, N125, N12);
not NOT1 (N132, N124);
or OR3 (N133, N132, N88, N17);
or OR4 (N134, N103, N28, N78, N6);
xor XOR2 (N135, N131, N37);
xor XOR2 (N136, N118, N62);
nand NAND4 (N137, N134, N64, N43, N99);
nor NOR2 (N138, N133, N67);
and AND2 (N139, N135, N47);
and AND4 (N140, N138, N41, N135, N100);
xor XOR2 (N141, N116, N119);
not NOT1 (N142, N141);
buf BUF1 (N143, N136);
not NOT1 (N144, N127);
not NOT1 (N145, N130);
or OR2 (N146, N126, N73);
xor XOR2 (N147, N139, N52);
nor NOR2 (N148, N147, N38);
not NOT1 (N149, N108);
buf BUF1 (N150, N140);
buf BUF1 (N151, N144);
nor NOR2 (N152, N145, N145);
buf BUF1 (N153, N148);
nand NAND4 (N154, N142, N114, N116, N8);
xor XOR2 (N155, N154, N71);
and AND4 (N156, N155, N29, N116, N35);
nand NAND4 (N157, N151, N2, N114, N22);
not NOT1 (N158, N156);
nor NOR2 (N159, N112, N47);
and AND3 (N160, N150, N120, N35);
or OR2 (N161, N152, N55);
nand NAND4 (N162, N153, N2, N100, N65);
xor XOR2 (N163, N157, N107);
nor NOR4 (N164, N149, N129, N61, N13);
and AND4 (N165, N137, N63, N133, N81);
nand NAND2 (N166, N146, N4);
not NOT1 (N167, N166);
and AND2 (N168, N163, N124);
buf BUF1 (N169, N160);
or OR3 (N170, N159, N69, N44);
and AND3 (N171, N143, N79, N133);
buf BUF1 (N172, N171);
or OR3 (N173, N172, N77, N70);
nor NOR2 (N174, N161, N31);
nand NAND3 (N175, N169, N12, N16);
or OR2 (N176, N162, N60);
xor XOR2 (N177, N175, N35);
nand NAND3 (N178, N173, N102, N111);
or OR3 (N179, N177, N126, N23);
and AND2 (N180, N168, N138);
xor XOR2 (N181, N164, N82);
and AND3 (N182, N158, N43, N78);
not NOT1 (N183, N179);
or OR3 (N184, N181, N109, N38);
buf BUF1 (N185, N178);
nand NAND2 (N186, N184, N180);
and AND3 (N187, N141, N173, N149);
or OR4 (N188, N165, N50, N27, N110);
xor XOR2 (N189, N188, N125);
nand NAND4 (N190, N170, N171, N97, N58);
nand NAND4 (N191, N189, N134, N71, N124);
nor NOR3 (N192, N185, N76, N38);
xor XOR2 (N193, N192, N187);
xor XOR2 (N194, N127, N178);
nor NOR2 (N195, N183, N139);
or OR4 (N196, N182, N145, N67, N40);
nor NOR2 (N197, N176, N194);
nand NAND2 (N198, N25, N175);
and AND2 (N199, N186, N139);
buf BUF1 (N200, N167);
not NOT1 (N201, N195);
nor NOR3 (N202, N191, N58, N192);
or OR4 (N203, N202, N91, N19, N60);
and AND2 (N204, N190, N101);
buf BUF1 (N205, N200);
buf BUF1 (N206, N198);
nand NAND3 (N207, N206, N17, N179);
not NOT1 (N208, N207);
nand NAND3 (N209, N174, N161, N160);
buf BUF1 (N210, N204);
nor NOR4 (N211, N208, N70, N24, N200);
and AND4 (N212, N205, N176, N48, N113);
buf BUF1 (N213, N203);
buf BUF1 (N214, N199);
nor NOR2 (N215, N193, N178);
nor NOR3 (N216, N213, N126, N94);
nor NOR2 (N217, N209, N5);
not NOT1 (N218, N215);
buf BUF1 (N219, N217);
not NOT1 (N220, N210);
buf BUF1 (N221, N219);
and AND3 (N222, N221, N48, N13);
xor XOR2 (N223, N197, N198);
nand NAND3 (N224, N218, N122, N151);
xor XOR2 (N225, N201, N39);
and AND2 (N226, N223, N19);
and AND2 (N227, N216, N60);
xor XOR2 (N228, N224, N46);
nor NOR4 (N229, N196, N222, N130, N3);
not NOT1 (N230, N2);
xor XOR2 (N231, N229, N121);
nor NOR3 (N232, N227, N137, N213);
or OR2 (N233, N230, N164);
nor NOR4 (N234, N232, N168, N158, N174);
or OR4 (N235, N231, N100, N202, N6);
and AND4 (N236, N212, N115, N25, N183);
buf BUF1 (N237, N226);
and AND3 (N238, N237, N202, N203);
or OR3 (N239, N220, N21, N172);
buf BUF1 (N240, N239);
nand NAND2 (N241, N211, N223);
nor NOR4 (N242, N236, N123, N67, N6);
and AND3 (N243, N235, N162, N232);
and AND4 (N244, N214, N229, N21, N160);
buf BUF1 (N245, N225);
xor XOR2 (N246, N245, N227);
or OR3 (N247, N244, N207, N109);
nor NOR3 (N248, N234, N172, N163);
or OR4 (N249, N242, N239, N70, N11);
and AND2 (N250, N241, N41);
nor NOR3 (N251, N246, N155, N118);
nand NAND2 (N252, N248, N234);
not NOT1 (N253, N233);
not NOT1 (N254, N238);
xor XOR2 (N255, N249, N16);
buf BUF1 (N256, N243);
nor NOR2 (N257, N252, N202);
not NOT1 (N258, N256);
nor NOR2 (N259, N257, N167);
nand NAND2 (N260, N253, N94);
xor XOR2 (N261, N240, N91);
nand NAND3 (N262, N254, N14, N35);
or OR3 (N263, N251, N83, N203);
xor XOR2 (N264, N255, N88);
not NOT1 (N265, N261);
nor NOR3 (N266, N259, N85, N179);
xor XOR2 (N267, N247, N14);
nor NOR2 (N268, N265, N66);
or OR4 (N269, N267, N117, N212, N44);
or OR4 (N270, N268, N244, N216, N251);
buf BUF1 (N271, N258);
nand NAND3 (N272, N260, N200, N200);
not NOT1 (N273, N271);
nand NAND2 (N274, N270, N120);
not NOT1 (N275, N264);
not NOT1 (N276, N228);
buf BUF1 (N277, N276);
buf BUF1 (N278, N275);
nand NAND2 (N279, N263, N203);
nand NAND3 (N280, N272, N248, N202);
nor NOR3 (N281, N274, N179, N38);
nand NAND2 (N282, N262, N172);
nor NOR2 (N283, N266, N271);
and AND4 (N284, N273, N29, N193, N73);
buf BUF1 (N285, N282);
xor XOR2 (N286, N283, N10);
nand NAND3 (N287, N286, N139, N202);
buf BUF1 (N288, N280);
not NOT1 (N289, N281);
xor XOR2 (N290, N277, N247);
or OR2 (N291, N284, N62);
nand NAND3 (N292, N290, N169, N46);
and AND4 (N293, N288, N211, N22, N276);
and AND2 (N294, N250, N84);
xor XOR2 (N295, N289, N200);
buf BUF1 (N296, N287);
or OR4 (N297, N294, N72, N130, N153);
buf BUF1 (N298, N293);
and AND4 (N299, N269, N75, N178, N252);
nor NOR4 (N300, N285, N147, N162, N122);
and AND2 (N301, N297, N104);
xor XOR2 (N302, N296, N85);
and AND3 (N303, N301, N225, N75);
and AND4 (N304, N299, N198, N300, N186);
xor XOR2 (N305, N61, N294);
xor XOR2 (N306, N305, N96);
or OR2 (N307, N302, N17);
or OR3 (N308, N298, N217, N30);
and AND4 (N309, N306, N39, N279, N179);
nor NOR4 (N310, N25, N176, N133, N30);
and AND2 (N311, N309, N119);
nor NOR3 (N312, N292, N151, N225);
and AND2 (N313, N308, N280);
and AND2 (N314, N291, N56);
buf BUF1 (N315, N312);
and AND4 (N316, N307, N184, N226, N313);
and AND4 (N317, N191, N17, N285, N285);
not NOT1 (N318, N278);
and AND2 (N319, N304, N259);
xor XOR2 (N320, N317, N42);
buf BUF1 (N321, N320);
nand NAND2 (N322, N316, N258);
nor NOR2 (N323, N315, N208);
xor XOR2 (N324, N295, N30);
not NOT1 (N325, N311);
nor NOR4 (N326, N323, N152, N107, N27);
nor NOR4 (N327, N314, N171, N149, N18);
xor XOR2 (N328, N322, N311);
nand NAND4 (N329, N318, N302, N78, N169);
not NOT1 (N330, N324);
buf BUF1 (N331, N327);
nor NOR3 (N332, N303, N146, N37);
not NOT1 (N333, N330);
and AND4 (N334, N329, N274, N320, N160);
not NOT1 (N335, N326);
and AND2 (N336, N325, N335);
xor XOR2 (N337, N95, N203);
buf BUF1 (N338, N337);
nand NAND2 (N339, N336, N245);
and AND2 (N340, N338, N44);
nor NOR4 (N341, N339, N168, N245, N76);
and AND4 (N342, N328, N164, N203, N199);
nor NOR2 (N343, N310, N179);
or OR3 (N344, N332, N281, N121);
or OR2 (N345, N343, N46);
not NOT1 (N346, N331);
or OR2 (N347, N334, N346);
or OR2 (N348, N66, N19);
and AND3 (N349, N347, N121, N199);
buf BUF1 (N350, N340);
buf BUF1 (N351, N319);
xor XOR2 (N352, N341, N17);
not NOT1 (N353, N342);
not NOT1 (N354, N353);
or OR4 (N355, N350, N329, N219, N258);
xor XOR2 (N356, N333, N104);
nand NAND4 (N357, N344, N128, N175, N103);
or OR4 (N358, N345, N333, N10, N112);
or OR4 (N359, N349, N246, N235, N300);
or OR4 (N360, N321, N292, N260, N175);
xor XOR2 (N361, N352, N322);
not NOT1 (N362, N351);
buf BUF1 (N363, N354);
or OR4 (N364, N360, N226, N119, N282);
or OR3 (N365, N356, N77, N104);
not NOT1 (N366, N355);
or OR3 (N367, N361, N276, N70);
nor NOR4 (N368, N364, N239, N11, N1);
nand NAND4 (N369, N365, N92, N199, N169);
and AND3 (N370, N362, N28, N229);
nand NAND3 (N371, N370, N370, N64);
xor XOR2 (N372, N363, N120);
or OR2 (N373, N359, N367);
nand NAND3 (N374, N179, N185, N223);
not NOT1 (N375, N368);
buf BUF1 (N376, N374);
or OR4 (N377, N375, N218, N223, N370);
nand NAND2 (N378, N371, N363);
not NOT1 (N379, N348);
nor NOR3 (N380, N376, N248, N210);
buf BUF1 (N381, N378);
or OR3 (N382, N369, N378, N114);
and AND2 (N383, N377, N43);
nor NOR2 (N384, N372, N186);
and AND3 (N385, N384, N332, N185);
xor XOR2 (N386, N385, N57);
nand NAND3 (N387, N357, N376, N237);
xor XOR2 (N388, N380, N47);
buf BUF1 (N389, N381);
nand NAND2 (N390, N379, N175);
not NOT1 (N391, N389);
buf BUF1 (N392, N366);
not NOT1 (N393, N392);
and AND4 (N394, N373, N241, N201, N302);
nand NAND2 (N395, N388, N108);
nor NOR2 (N396, N358, N389);
nand NAND3 (N397, N394, N351, N70);
not NOT1 (N398, N382);
and AND4 (N399, N395, N277, N242, N333);
not NOT1 (N400, N398);
or OR3 (N401, N396, N269, N204);
buf BUF1 (N402, N393);
xor XOR2 (N403, N399, N249);
and AND3 (N404, N390, N370, N34);
or OR2 (N405, N397, N327);
xor XOR2 (N406, N391, N379);
or OR2 (N407, N403, N270);
nand NAND3 (N408, N404, N386, N123);
buf BUF1 (N409, N76);
nand NAND2 (N410, N387, N364);
not NOT1 (N411, N402);
not NOT1 (N412, N401);
nand NAND3 (N413, N412, N72, N14);
xor XOR2 (N414, N400, N311);
xor XOR2 (N415, N411, N91);
and AND2 (N416, N413, N92);
xor XOR2 (N417, N383, N90);
or OR4 (N418, N416, N386, N13, N28);
not NOT1 (N419, N405);
not NOT1 (N420, N414);
or OR3 (N421, N407, N93, N226);
or OR4 (N422, N410, N360, N183, N229);
xor XOR2 (N423, N418, N22);
nor NOR2 (N424, N421, N80);
not NOT1 (N425, N406);
or OR3 (N426, N419, N417, N2);
not NOT1 (N427, N346);
nor NOR3 (N428, N427, N292, N105);
not NOT1 (N429, N424);
and AND3 (N430, N423, N39, N51);
nand NAND2 (N431, N429, N348);
xor XOR2 (N432, N415, N60);
nor NOR4 (N433, N430, N241, N194, N419);
nand NAND3 (N434, N408, N188, N42);
and AND4 (N435, N433, N204, N319, N394);
buf BUF1 (N436, N432);
or OR2 (N437, N409, N118);
or OR2 (N438, N437, N405);
or OR4 (N439, N434, N143, N436, N187);
xor XOR2 (N440, N72, N276);
or OR4 (N441, N428, N235, N204, N44);
not NOT1 (N442, N426);
xor XOR2 (N443, N440, N387);
nand NAND4 (N444, N442, N305, N394, N54);
and AND3 (N445, N425, N256, N399);
or OR4 (N446, N445, N392, N7, N18);
nor NOR4 (N447, N443, N287, N409, N112);
nand NAND3 (N448, N438, N270, N86);
nor NOR2 (N449, N431, N365);
or OR3 (N450, N422, N330, N24);
buf BUF1 (N451, N439);
buf BUF1 (N452, N451);
xor XOR2 (N453, N446, N131);
xor XOR2 (N454, N449, N395);
not NOT1 (N455, N435);
xor XOR2 (N456, N448, N377);
or OR4 (N457, N450, N444, N456, N174);
nand NAND4 (N458, N159, N157, N167, N439);
and AND2 (N459, N13, N81);
or OR3 (N460, N441, N33, N239);
and AND3 (N461, N452, N22, N262);
not NOT1 (N462, N459);
buf BUF1 (N463, N447);
xor XOR2 (N464, N458, N312);
xor XOR2 (N465, N454, N193);
xor XOR2 (N466, N455, N212);
or OR4 (N467, N460, N233, N267, N397);
not NOT1 (N468, N465);
or OR3 (N469, N420, N273, N312);
nand NAND3 (N470, N467, N9, N132);
nor NOR2 (N471, N466, N26);
nand NAND2 (N472, N463, N109);
buf BUF1 (N473, N453);
nor NOR2 (N474, N461, N366);
nor NOR2 (N475, N468, N417);
or OR3 (N476, N470, N37, N214);
not NOT1 (N477, N462);
not NOT1 (N478, N472);
and AND2 (N479, N469, N5);
buf BUF1 (N480, N476);
nor NOR3 (N481, N473, N253, N331);
and AND3 (N482, N464, N388, N204);
or OR3 (N483, N479, N191, N87);
not NOT1 (N484, N471);
xor XOR2 (N485, N483, N202);
nor NOR4 (N486, N480, N416, N479, N165);
nor NOR3 (N487, N484, N142, N134);
nand NAND4 (N488, N478, N181, N450, N164);
or OR4 (N489, N482, N162, N218, N104);
buf BUF1 (N490, N488);
xor XOR2 (N491, N485, N33);
xor XOR2 (N492, N489, N491);
and AND4 (N493, N95, N362, N375, N464);
buf BUF1 (N494, N487);
nor NOR2 (N495, N494, N69);
nand NAND4 (N496, N492, N449, N187, N114);
or OR3 (N497, N490, N280, N89);
nor NOR3 (N498, N477, N378, N118);
nand NAND4 (N499, N495, N186, N199, N469);
not NOT1 (N500, N475);
nor NOR2 (N501, N496, N240);
xor XOR2 (N502, N457, N467);
and AND2 (N503, N474, N46);
and AND3 (N504, N486, N192, N451);
xor XOR2 (N505, N493, N463);
nor NOR3 (N506, N502, N139, N72);
buf BUF1 (N507, N504);
nor NOR3 (N508, N505, N142, N323);
not NOT1 (N509, N500);
xor XOR2 (N510, N506, N393);
xor XOR2 (N511, N509, N478);
xor XOR2 (N512, N481, N257);
nand NAND2 (N513, N510, N504);
or OR3 (N514, N499, N347, N398);
not NOT1 (N515, N508);
nor NOR2 (N516, N503, N448);
xor XOR2 (N517, N513, N272);
not NOT1 (N518, N501);
and AND2 (N519, N512, N1);
nor NOR3 (N520, N518, N58, N514);
nand NAND3 (N521, N199, N269, N283);
buf BUF1 (N522, N521);
nand NAND4 (N523, N507, N424, N239, N412);
not NOT1 (N524, N515);
nand NAND4 (N525, N520, N239, N350, N238);
nand NAND4 (N526, N498, N163, N424, N448);
or OR4 (N527, N516, N32, N216, N520);
not NOT1 (N528, N526);
and AND4 (N529, N519, N17, N486, N501);
nor NOR3 (N530, N528, N384, N309);
not NOT1 (N531, N523);
or OR4 (N532, N522, N497, N439, N507);
buf BUF1 (N533, N193);
nand NAND4 (N534, N511, N514, N468, N60);
and AND4 (N535, N529, N68, N447, N456);
or OR4 (N536, N534, N295, N412, N305);
nor NOR2 (N537, N535, N154);
nand NAND4 (N538, N536, N137, N425, N177);
and AND4 (N539, N537, N268, N141, N326);
nor NOR4 (N540, N539, N271, N443, N203);
nand NAND4 (N541, N533, N411, N110, N225);
buf BUF1 (N542, N540);
or OR4 (N543, N531, N457, N525, N427);
nor NOR3 (N544, N500, N381, N175);
xor XOR2 (N545, N538, N544);
xor XOR2 (N546, N389, N162);
nand NAND2 (N547, N541, N29);
buf BUF1 (N548, N545);
or OR3 (N549, N530, N346, N528);
not NOT1 (N550, N517);
and AND4 (N551, N524, N509, N250, N478);
and AND3 (N552, N550, N318, N217);
nor NOR4 (N553, N543, N92, N66, N289);
xor XOR2 (N554, N546, N40);
nand NAND4 (N555, N554, N27, N364, N56);
buf BUF1 (N556, N542);
not NOT1 (N557, N552);
or OR2 (N558, N553, N125);
nor NOR3 (N559, N557, N81, N517);
nand NAND4 (N560, N549, N132, N520, N522);
nor NOR2 (N561, N551, N200);
or OR4 (N562, N548, N523, N6, N102);
nor NOR2 (N563, N547, N238);
or OR4 (N564, N563, N289, N269, N489);
nand NAND3 (N565, N564, N430, N441);
buf BUF1 (N566, N556);
nand NAND3 (N567, N560, N257, N383);
not NOT1 (N568, N562);
or OR3 (N569, N532, N402, N489);
and AND4 (N570, N561, N154, N317, N190);
nor NOR4 (N571, N558, N527, N352, N164);
nor NOR2 (N572, N407, N146);
xor XOR2 (N573, N565, N473);
buf BUF1 (N574, N566);
buf BUF1 (N575, N573);
not NOT1 (N576, N570);
buf BUF1 (N577, N568);
buf BUF1 (N578, N571);
nor NOR3 (N579, N555, N213, N508);
nand NAND3 (N580, N567, N422, N12);
not NOT1 (N581, N569);
xor XOR2 (N582, N559, N451);
nand NAND2 (N583, N577, N312);
nor NOR4 (N584, N574, N267, N327, N128);
nor NOR3 (N585, N581, N410, N462);
nand NAND4 (N586, N578, N413, N550, N581);
nor NOR3 (N587, N572, N140, N190);
buf BUF1 (N588, N585);
and AND4 (N589, N586, N453, N574, N576);
xor XOR2 (N590, N332, N451);
buf BUF1 (N591, N575);
or OR4 (N592, N580, N473, N529, N568);
nor NOR2 (N593, N584, N64);
or OR2 (N594, N582, N435);
nand NAND4 (N595, N583, N545, N376, N98);
and AND2 (N596, N588, N27);
and AND3 (N597, N592, N390, N581);
not NOT1 (N598, N595);
buf BUF1 (N599, N597);
buf BUF1 (N600, N599);
or OR4 (N601, N600, N344, N135, N384);
nor NOR4 (N602, N601, N122, N291, N400);
nor NOR2 (N603, N587, N18);
nor NOR4 (N604, N579, N302, N147, N50);
buf BUF1 (N605, N589);
buf BUF1 (N606, N593);
not NOT1 (N607, N591);
and AND3 (N608, N594, N303, N358);
nand NAND2 (N609, N596, N149);
or OR3 (N610, N604, N535, N14);
buf BUF1 (N611, N602);
not NOT1 (N612, N605);
not NOT1 (N613, N606);
not NOT1 (N614, N609);
buf BUF1 (N615, N590);
nor NOR2 (N616, N613, N417);
nor NOR2 (N617, N603, N52);
not NOT1 (N618, N616);
nor NOR2 (N619, N608, N61);
and AND4 (N620, N614, N289, N270, N336);
nor NOR3 (N621, N615, N217, N45);
not NOT1 (N622, N620);
buf BUF1 (N623, N617);
or OR4 (N624, N607, N228, N191, N460);
nand NAND2 (N625, N619, N195);
and AND4 (N626, N625, N354, N107, N573);
nand NAND3 (N627, N621, N333, N235);
or OR3 (N628, N623, N565, N141);
nor NOR3 (N629, N611, N67, N228);
xor XOR2 (N630, N627, N407);
buf BUF1 (N631, N630);
xor XOR2 (N632, N618, N491);
nand NAND3 (N633, N624, N70, N37);
and AND3 (N634, N598, N494, N503);
xor XOR2 (N635, N610, N197);
not NOT1 (N636, N622);
xor XOR2 (N637, N632, N46);
nand NAND4 (N638, N629, N497, N582, N253);
nand NAND4 (N639, N634, N17, N303, N360);
or OR2 (N640, N638, N558);
not NOT1 (N641, N640);
nand NAND3 (N642, N628, N114, N295);
nand NAND3 (N643, N642, N140, N134);
nor NOR2 (N644, N626, N73);
or OR4 (N645, N644, N8, N294, N574);
nor NOR3 (N646, N639, N23, N621);
and AND3 (N647, N631, N61, N628);
or OR3 (N648, N647, N481, N150);
nor NOR4 (N649, N648, N430, N104, N165);
not NOT1 (N650, N636);
buf BUF1 (N651, N645);
or OR3 (N652, N612, N573, N320);
or OR4 (N653, N649, N140, N407, N229);
or OR2 (N654, N643, N96);
buf BUF1 (N655, N646);
buf BUF1 (N656, N635);
not NOT1 (N657, N655);
or OR4 (N658, N637, N644, N5, N404);
not NOT1 (N659, N652);
buf BUF1 (N660, N656);
or OR2 (N661, N651, N480);
or OR4 (N662, N641, N641, N428, N245);
buf BUF1 (N663, N662);
and AND3 (N664, N658, N143, N291);
and AND3 (N665, N660, N531, N11);
not NOT1 (N666, N661);
buf BUF1 (N667, N633);
or OR2 (N668, N663, N630);
nand NAND4 (N669, N659, N443, N197, N231);
or OR4 (N670, N657, N144, N102, N569);
xor XOR2 (N671, N653, N270);
not NOT1 (N672, N666);
buf BUF1 (N673, N665);
nand NAND4 (N674, N664, N351, N317, N415);
or OR4 (N675, N650, N174, N48, N425);
xor XOR2 (N676, N673, N467);
or OR3 (N677, N675, N110, N67);
nand NAND2 (N678, N672, N645);
and AND4 (N679, N670, N279, N403, N74);
nand NAND2 (N680, N669, N137);
or OR3 (N681, N668, N462, N211);
not NOT1 (N682, N667);
buf BUF1 (N683, N677);
not NOT1 (N684, N680);
nand NAND4 (N685, N684, N243, N523, N133);
buf BUF1 (N686, N682);
and AND4 (N687, N681, N611, N597, N645);
nand NAND3 (N688, N654, N51, N151);
and AND3 (N689, N688, N37, N600);
and AND2 (N690, N674, N168);
xor XOR2 (N691, N671, N203);
not NOT1 (N692, N687);
not NOT1 (N693, N690);
or OR4 (N694, N692, N650, N141, N579);
nand NAND3 (N695, N689, N648, N579);
nand NAND4 (N696, N683, N495, N615, N564);
nand NAND2 (N697, N693, N475);
not NOT1 (N698, N678);
nand NAND3 (N699, N696, N446, N697);
not NOT1 (N700, N228);
nand NAND2 (N701, N700, N6);
nor NOR3 (N702, N685, N107, N300);
xor XOR2 (N703, N679, N605);
nor NOR3 (N704, N676, N662, N84);
nand NAND3 (N705, N694, N284, N562);
or OR2 (N706, N704, N339);
nor NOR3 (N707, N686, N186, N347);
and AND4 (N708, N698, N618, N9, N15);
or OR4 (N709, N705, N66, N437, N648);
nor NOR4 (N710, N701, N328, N465, N465);
nor NOR4 (N711, N708, N565, N366, N584);
or OR2 (N712, N709, N339);
or OR2 (N713, N712, N427);
or OR4 (N714, N702, N534, N356, N372);
and AND3 (N715, N703, N702, N312);
not NOT1 (N716, N715);
buf BUF1 (N717, N711);
or OR3 (N718, N717, N12, N206);
buf BUF1 (N719, N713);
buf BUF1 (N720, N710);
or OR3 (N721, N718, N556, N132);
nor NOR3 (N722, N716, N466, N281);
or OR3 (N723, N706, N471, N108);
xor XOR2 (N724, N714, N406);
xor XOR2 (N725, N722, N499);
nand NAND2 (N726, N719, N366);
nand NAND2 (N727, N695, N721);
nand NAND4 (N728, N569, N343, N103, N591);
and AND3 (N729, N727, N570, N456);
nor NOR3 (N730, N724, N563, N448);
or OR4 (N731, N728, N44, N672, N3);
not NOT1 (N732, N707);
or OR3 (N733, N726, N426, N239);
nand NAND3 (N734, N732, N333, N464);
nand NAND3 (N735, N723, N141, N711);
xor XOR2 (N736, N691, N602);
nand NAND2 (N737, N720, N636);
and AND3 (N738, N736, N734, N213);
buf BUF1 (N739, N477);
not NOT1 (N740, N737);
or OR2 (N741, N735, N404);
buf BUF1 (N742, N730);
buf BUF1 (N743, N731);
or OR3 (N744, N740, N153, N424);
and AND4 (N745, N729, N64, N495, N56);
nand NAND4 (N746, N733, N350, N211, N606);
nand NAND2 (N747, N746, N214);
not NOT1 (N748, N741);
not NOT1 (N749, N748);
not NOT1 (N750, N738);
xor XOR2 (N751, N739, N166);
or OR4 (N752, N751, N392, N360, N381);
or OR3 (N753, N750, N638, N735);
not NOT1 (N754, N725);
buf BUF1 (N755, N754);
nand NAND3 (N756, N753, N609, N636);
or OR4 (N757, N744, N131, N352, N123);
buf BUF1 (N758, N742);
xor XOR2 (N759, N699, N356);
buf BUF1 (N760, N749);
and AND2 (N761, N759, N646);
not NOT1 (N762, N756);
nand NAND3 (N763, N762, N43, N571);
not NOT1 (N764, N758);
nand NAND2 (N765, N763, N397);
not NOT1 (N766, N761);
not NOT1 (N767, N757);
nor NOR2 (N768, N760, N545);
xor XOR2 (N769, N767, N570);
buf BUF1 (N770, N745);
not NOT1 (N771, N766);
buf BUF1 (N772, N752);
xor XOR2 (N773, N769, N666);
and AND4 (N774, N764, N580, N609, N667);
xor XOR2 (N775, N768, N578);
buf BUF1 (N776, N775);
nor NOR2 (N777, N776, N402);
or OR2 (N778, N777, N733);
not NOT1 (N779, N774);
and AND2 (N780, N778, N450);
xor XOR2 (N781, N780, N97);
not NOT1 (N782, N765);
xor XOR2 (N783, N781, N303);
buf BUF1 (N784, N772);
not NOT1 (N785, N773);
nand NAND2 (N786, N747, N659);
nor NOR4 (N787, N785, N228, N748, N135);
not NOT1 (N788, N787);
buf BUF1 (N789, N779);
or OR4 (N790, N788, N714, N345, N177);
or OR2 (N791, N790, N289);
not NOT1 (N792, N786);
xor XOR2 (N793, N791, N28);
nand NAND2 (N794, N789, N298);
nor NOR2 (N795, N792, N397);
not NOT1 (N796, N782);
nand NAND3 (N797, N796, N580, N549);
or OR3 (N798, N793, N355, N426);
not NOT1 (N799, N794);
and AND2 (N800, N795, N709);
xor XOR2 (N801, N783, N381);
and AND3 (N802, N800, N761, N571);
xor XOR2 (N803, N802, N456);
buf BUF1 (N804, N784);
and AND3 (N805, N799, N700, N163);
or OR2 (N806, N804, N88);
nor NOR3 (N807, N743, N778, N289);
xor XOR2 (N808, N798, N479);
nor NOR3 (N809, N803, N287, N199);
buf BUF1 (N810, N755);
buf BUF1 (N811, N771);
nor NOR3 (N812, N770, N25, N25);
or OR3 (N813, N806, N135, N729);
nor NOR3 (N814, N797, N378, N584);
buf BUF1 (N815, N809);
xor XOR2 (N816, N805, N197);
and AND3 (N817, N810, N329, N399);
not NOT1 (N818, N813);
nand NAND4 (N819, N817, N653, N41, N209);
nor NOR2 (N820, N812, N306);
nand NAND2 (N821, N816, N523);
and AND4 (N822, N807, N546, N37, N361);
and AND3 (N823, N819, N122, N698);
and AND4 (N824, N808, N311, N678, N738);
or OR4 (N825, N824, N698, N412, N206);
nor NOR3 (N826, N815, N345, N321);
nor NOR4 (N827, N801, N300, N64, N404);
and AND3 (N828, N822, N503, N651);
not NOT1 (N829, N823);
xor XOR2 (N830, N821, N218);
xor XOR2 (N831, N826, N413);
buf BUF1 (N832, N820);
or OR2 (N833, N830, N641);
not NOT1 (N834, N829);
and AND3 (N835, N818, N119, N298);
buf BUF1 (N836, N814);
or OR4 (N837, N825, N299, N439, N650);
xor XOR2 (N838, N832, N38);
and AND3 (N839, N811, N784, N781);
nand NAND3 (N840, N836, N12, N400);
or OR3 (N841, N828, N242, N349);
not NOT1 (N842, N833);
nor NOR4 (N843, N835, N511, N181, N726);
not NOT1 (N844, N843);
or OR2 (N845, N844, N714);
nor NOR4 (N846, N845, N337, N695, N554);
nand NAND4 (N847, N841, N467, N425, N292);
buf BUF1 (N848, N838);
nand NAND4 (N849, N846, N792, N366, N737);
buf BUF1 (N850, N831);
nand NAND4 (N851, N827, N227, N710, N313);
not NOT1 (N852, N849);
not NOT1 (N853, N842);
not NOT1 (N854, N848);
xor XOR2 (N855, N853, N480);
nor NOR3 (N856, N847, N678, N292);
or OR4 (N857, N851, N4, N292, N500);
nand NAND4 (N858, N839, N375, N164, N101);
not NOT1 (N859, N858);
buf BUF1 (N860, N837);
and AND4 (N861, N857, N504, N99, N610);
not NOT1 (N862, N859);
nor NOR2 (N863, N852, N517);
xor XOR2 (N864, N856, N596);
nor NOR2 (N865, N860, N366);
nor NOR3 (N866, N863, N433, N28);
xor XOR2 (N867, N864, N144);
nor NOR4 (N868, N854, N638, N541, N201);
buf BUF1 (N869, N840);
nor NOR4 (N870, N865, N666, N515, N852);
nor NOR4 (N871, N862, N679, N58, N30);
buf BUF1 (N872, N855);
and AND3 (N873, N834, N148, N441);
and AND2 (N874, N870, N775);
nand NAND2 (N875, N850, N244);
not NOT1 (N876, N871);
and AND2 (N877, N876, N641);
nand NAND4 (N878, N861, N240, N316, N511);
xor XOR2 (N879, N866, N515);
and AND4 (N880, N878, N505, N441, N816);
xor XOR2 (N881, N869, N346);
nand NAND3 (N882, N875, N219, N564);
xor XOR2 (N883, N881, N123);
nand NAND2 (N884, N873, N304);
and AND4 (N885, N877, N131, N442, N869);
or OR2 (N886, N885, N86);
buf BUF1 (N887, N867);
or OR2 (N888, N879, N677);
not NOT1 (N889, N872);
or OR4 (N890, N889, N306, N215, N414);
not NOT1 (N891, N868);
nor NOR4 (N892, N882, N742, N416, N431);
not NOT1 (N893, N884);
and AND3 (N894, N880, N594, N358);
not NOT1 (N895, N890);
nand NAND3 (N896, N892, N57, N618);
nand NAND2 (N897, N883, N6);
nor NOR4 (N898, N895, N289, N267, N634);
and AND2 (N899, N888, N485);
and AND4 (N900, N886, N311, N390, N633);
and AND3 (N901, N898, N473, N165);
and AND4 (N902, N893, N850, N131, N129);
buf BUF1 (N903, N901);
xor XOR2 (N904, N887, N502);
or OR4 (N905, N874, N420, N374, N479);
or OR2 (N906, N891, N343);
nor NOR4 (N907, N897, N754, N723, N304);
nor NOR2 (N908, N902, N853);
or OR4 (N909, N900, N686, N468, N52);
nand NAND2 (N910, N905, N293);
and AND2 (N911, N909, N48);
not NOT1 (N912, N911);
nand NAND2 (N913, N903, N628);
xor XOR2 (N914, N910, N682);
or OR2 (N915, N913, N430);
xor XOR2 (N916, N899, N705);
nor NOR4 (N917, N908, N302, N594, N537);
nor NOR4 (N918, N916, N44, N107, N886);
not NOT1 (N919, N914);
nand NAND2 (N920, N896, N797);
nor NOR4 (N921, N920, N790, N324, N899);
nor NOR3 (N922, N906, N504, N84);
nor NOR2 (N923, N907, N652);
not NOT1 (N924, N894);
nand NAND2 (N925, N924, N401);
not NOT1 (N926, N922);
nand NAND4 (N927, N926, N58, N556, N376);
xor XOR2 (N928, N925, N426);
nor NOR4 (N929, N919, N109, N293, N408);
buf BUF1 (N930, N928);
nand NAND2 (N931, N923, N199);
not NOT1 (N932, N917);
nand NAND3 (N933, N931, N663, N890);
buf BUF1 (N934, N904);
nor NOR3 (N935, N912, N36, N325);
nand NAND4 (N936, N927, N766, N881, N7);
buf BUF1 (N937, N935);
and AND4 (N938, N932, N248, N345, N430);
nand NAND3 (N939, N918, N272, N97);
and AND4 (N940, N933, N166, N14, N87);
xor XOR2 (N941, N929, N675);
not NOT1 (N942, N940);
or OR2 (N943, N934, N71);
buf BUF1 (N944, N942);
or OR3 (N945, N938, N548, N934);
and AND4 (N946, N943, N532, N391, N641);
nor NOR4 (N947, N945, N909, N271, N222);
and AND4 (N948, N947, N786, N325, N118);
xor XOR2 (N949, N937, N454);
xor XOR2 (N950, N936, N846);
nor NOR3 (N951, N915, N201, N679);
nor NOR2 (N952, N950, N209);
xor XOR2 (N953, N921, N251);
nor NOR3 (N954, N939, N676, N730);
or OR3 (N955, N944, N311, N560);
not NOT1 (N956, N953);
or OR4 (N957, N951, N141, N533, N945);
or OR2 (N958, N956, N783);
and AND3 (N959, N941, N740, N224);
nor NOR2 (N960, N958, N403);
buf BUF1 (N961, N946);
xor XOR2 (N962, N930, N226);
and AND2 (N963, N960, N776);
nor NOR3 (N964, N955, N234, N208);
nor NOR3 (N965, N948, N570, N399);
not NOT1 (N966, N963);
and AND4 (N967, N962, N655, N758, N874);
buf BUF1 (N968, N965);
or OR2 (N969, N949, N844);
xor XOR2 (N970, N967, N394);
xor XOR2 (N971, N961, N47);
buf BUF1 (N972, N968);
nand NAND2 (N973, N959, N496);
xor XOR2 (N974, N969, N829);
buf BUF1 (N975, N952);
xor XOR2 (N976, N975, N396);
nor NOR4 (N977, N974, N938, N329, N900);
not NOT1 (N978, N957);
xor XOR2 (N979, N964, N343);
xor XOR2 (N980, N976, N46);
or OR3 (N981, N979, N928, N507);
xor XOR2 (N982, N978, N25);
or OR3 (N983, N971, N288, N749);
nand NAND4 (N984, N983, N941, N837, N458);
nand NAND3 (N985, N973, N133, N279);
nand NAND2 (N986, N966, N336);
or OR2 (N987, N984, N508);
and AND4 (N988, N981, N49, N966, N285);
nor NOR2 (N989, N988, N548);
or OR3 (N990, N986, N984, N113);
or OR3 (N991, N985, N584, N759);
not NOT1 (N992, N980);
xor XOR2 (N993, N977, N51);
nor NOR3 (N994, N982, N456, N401);
nand NAND3 (N995, N994, N621, N684);
nor NOR4 (N996, N991, N69, N718, N19);
xor XOR2 (N997, N954, N944);
nand NAND4 (N998, N996, N987, N602, N975);
or OR4 (N999, N773, N813, N447, N671);
not NOT1 (N1000, N995);
nor NOR3 (N1001, N999, N928, N213);
buf BUF1 (N1002, N990);
nor NOR3 (N1003, N993, N322, N969);
xor XOR2 (N1004, N1003, N263);
or OR4 (N1005, N998, N473, N680, N687);
or OR3 (N1006, N970, N207, N562);
nor NOR2 (N1007, N1006, N111);
nand NAND3 (N1008, N972, N859, N462);
nor NOR4 (N1009, N997, N782, N761, N244);
buf BUF1 (N1010, N1005);
and AND4 (N1011, N1000, N934, N611, N827);
or OR2 (N1012, N1011, N71);
or OR4 (N1013, N1002, N105, N939, N115);
not NOT1 (N1014, N1008);
nand NAND3 (N1015, N1009, N139, N312);
buf BUF1 (N1016, N992);
or OR4 (N1017, N1004, N782, N860, N629);
not NOT1 (N1018, N1001);
and AND3 (N1019, N1012, N781, N170);
buf BUF1 (N1020, N1019);
nor NOR2 (N1021, N989, N513);
or OR2 (N1022, N1017, N973);
or OR4 (N1023, N1021, N231, N119, N887);
and AND2 (N1024, N1015, N72);
nand NAND4 (N1025, N1007, N133, N600, N7);
xor XOR2 (N1026, N1020, N275);
nand NAND3 (N1027, N1025, N591, N219);
buf BUF1 (N1028, N1022);
nor NOR2 (N1029, N1014, N62);
buf BUF1 (N1030, N1026);
buf BUF1 (N1031, N1023);
nor NOR3 (N1032, N1018, N128, N875);
nor NOR4 (N1033, N1010, N1016, N337, N764);
xor XOR2 (N1034, N751, N287);
nand NAND3 (N1035, N1031, N923, N458);
xor XOR2 (N1036, N1024, N996);
not NOT1 (N1037, N1027);
not NOT1 (N1038, N1036);
xor XOR2 (N1039, N1013, N882);
nor NOR4 (N1040, N1039, N725, N610, N369);
and AND2 (N1041, N1030, N249);
xor XOR2 (N1042, N1032, N116);
not NOT1 (N1043, N1033);
buf BUF1 (N1044, N1034);
and AND2 (N1045, N1043, N1000);
nand NAND4 (N1046, N1045, N649, N819, N238);
and AND4 (N1047, N1037, N837, N15, N752);
xor XOR2 (N1048, N1040, N988);
not NOT1 (N1049, N1047);
or OR2 (N1050, N1042, N1012);
buf BUF1 (N1051, N1029);
buf BUF1 (N1052, N1046);
xor XOR2 (N1053, N1049, N935);
xor XOR2 (N1054, N1041, N99);
xor XOR2 (N1055, N1038, N667);
nor NOR2 (N1056, N1055, N801);
nor NOR4 (N1057, N1051, N386, N882, N924);
buf BUF1 (N1058, N1053);
buf BUF1 (N1059, N1054);
or OR2 (N1060, N1050, N884);
not NOT1 (N1061, N1060);
nand NAND3 (N1062, N1044, N254, N116);
nand NAND3 (N1063, N1048, N658, N12);
xor XOR2 (N1064, N1059, N522);
not NOT1 (N1065, N1062);
and AND4 (N1066, N1058, N1036, N165, N785);
buf BUF1 (N1067, N1028);
nand NAND4 (N1068, N1056, N794, N520, N893);
nand NAND2 (N1069, N1061, N553);
not NOT1 (N1070, N1068);
or OR2 (N1071, N1035, N712);
or OR2 (N1072, N1070, N538);
xor XOR2 (N1073, N1064, N319);
buf BUF1 (N1074, N1052);
nor NOR4 (N1075, N1074, N147, N1016, N138);
nand NAND3 (N1076, N1067, N1010, N788);
and AND3 (N1077, N1071, N713, N244);
nand NAND4 (N1078, N1057, N796, N339, N648);
not NOT1 (N1079, N1077);
and AND2 (N1080, N1073, N346);
nor NOR2 (N1081, N1080, N633);
or OR3 (N1082, N1069, N532, N821);
and AND4 (N1083, N1065, N189, N550, N983);
or OR3 (N1084, N1076, N204, N18);
xor XOR2 (N1085, N1081, N1066);
xor XOR2 (N1086, N865, N770);
nand NAND4 (N1087, N1085, N483, N718, N825);
not NOT1 (N1088, N1063);
nor NOR2 (N1089, N1086, N708);
buf BUF1 (N1090, N1083);
buf BUF1 (N1091, N1075);
nor NOR2 (N1092, N1090, N42);
and AND2 (N1093, N1088, N794);
nand NAND4 (N1094, N1093, N398, N944, N858);
nand NAND2 (N1095, N1091, N217);
nand NAND3 (N1096, N1087, N883, N955);
xor XOR2 (N1097, N1078, N418);
and AND2 (N1098, N1084, N525);
nand NAND2 (N1099, N1095, N671);
nor NOR3 (N1100, N1097, N340, N38);
and AND2 (N1101, N1082, N524);
or OR3 (N1102, N1101, N1089, N459);
or OR2 (N1103, N445, N167);
and AND4 (N1104, N1079, N514, N979, N470);
nor NOR3 (N1105, N1096, N878, N42);
and AND4 (N1106, N1100, N256, N81, N892);
nor NOR2 (N1107, N1105, N308);
xor XOR2 (N1108, N1104, N832);
nand NAND2 (N1109, N1092, N1075);
xor XOR2 (N1110, N1107, N43);
and AND3 (N1111, N1099, N73, N643);
nand NAND3 (N1112, N1109, N493, N1076);
not NOT1 (N1113, N1102);
nor NOR2 (N1114, N1111, N1067);
nand NAND3 (N1115, N1098, N752, N747);
xor XOR2 (N1116, N1110, N541);
not NOT1 (N1117, N1112);
nor NOR2 (N1118, N1094, N136);
not NOT1 (N1119, N1115);
nor NOR3 (N1120, N1108, N653, N341);
not NOT1 (N1121, N1113);
xor XOR2 (N1122, N1120, N422);
or OR2 (N1123, N1114, N309);
nor NOR2 (N1124, N1072, N758);
nor NOR4 (N1125, N1106, N793, N931, N197);
not NOT1 (N1126, N1118);
xor XOR2 (N1127, N1126, N285);
or OR4 (N1128, N1123, N786, N173, N779);
not NOT1 (N1129, N1127);
xor XOR2 (N1130, N1125, N172);
or OR2 (N1131, N1121, N508);
nor NOR2 (N1132, N1131, N728);
not NOT1 (N1133, N1128);
xor XOR2 (N1134, N1133, N664);
nor NOR4 (N1135, N1130, N318, N1116, N337);
xor XOR2 (N1136, N606, N384);
buf BUF1 (N1137, N1135);
and AND3 (N1138, N1117, N953, N11);
buf BUF1 (N1139, N1103);
or OR4 (N1140, N1138, N909, N66, N457);
or OR3 (N1141, N1139, N809, N208);
not NOT1 (N1142, N1134);
not NOT1 (N1143, N1140);
and AND2 (N1144, N1143, N961);
not NOT1 (N1145, N1142);
not NOT1 (N1146, N1124);
not NOT1 (N1147, N1136);
or OR3 (N1148, N1141, N391, N458);
or OR3 (N1149, N1122, N498, N169);
xor XOR2 (N1150, N1147, N927);
buf BUF1 (N1151, N1148);
xor XOR2 (N1152, N1137, N1013);
and AND4 (N1153, N1146, N523, N769, N543);
nor NOR3 (N1154, N1119, N520, N457);
or OR4 (N1155, N1153, N22, N1123, N557);
not NOT1 (N1156, N1132);
not NOT1 (N1157, N1156);
buf BUF1 (N1158, N1129);
nand NAND4 (N1159, N1145, N126, N500, N395);
and AND2 (N1160, N1144, N996);
nand NAND2 (N1161, N1149, N169);
nand NAND4 (N1162, N1150, N634, N367, N478);
not NOT1 (N1163, N1159);
nand NAND4 (N1164, N1158, N459, N595, N937);
or OR2 (N1165, N1162, N20);
not NOT1 (N1166, N1163);
and AND3 (N1167, N1151, N357, N804);
or OR3 (N1168, N1167, N416, N813);
xor XOR2 (N1169, N1157, N779);
xor XOR2 (N1170, N1166, N766);
not NOT1 (N1171, N1160);
buf BUF1 (N1172, N1152);
nand NAND3 (N1173, N1171, N1022, N480);
buf BUF1 (N1174, N1165);
not NOT1 (N1175, N1154);
buf BUF1 (N1176, N1168);
buf BUF1 (N1177, N1173);
or OR3 (N1178, N1170, N606, N1107);
buf BUF1 (N1179, N1175);
nand NAND3 (N1180, N1177, N1162, N819);
xor XOR2 (N1181, N1164, N383);
buf BUF1 (N1182, N1176);
not NOT1 (N1183, N1182);
or OR2 (N1184, N1180, N131);
nor NOR2 (N1185, N1174, N518);
or OR3 (N1186, N1181, N949, N106);
or OR4 (N1187, N1179, N958, N450, N383);
or OR4 (N1188, N1178, N974, N379, N566);
xor XOR2 (N1189, N1187, N888);
nor NOR3 (N1190, N1183, N374, N493);
not NOT1 (N1191, N1186);
nand NAND2 (N1192, N1190, N501);
buf BUF1 (N1193, N1184);
xor XOR2 (N1194, N1155, N378);
nor NOR3 (N1195, N1192, N224, N422);
or OR4 (N1196, N1191, N751, N812, N578);
and AND4 (N1197, N1172, N3, N532, N19);
nand NAND3 (N1198, N1169, N915, N1048);
buf BUF1 (N1199, N1193);
and AND3 (N1200, N1161, N776, N1024);
and AND2 (N1201, N1194, N944);
nor NOR2 (N1202, N1195, N1043);
or OR3 (N1203, N1198, N525, N221);
nand NAND4 (N1204, N1196, N1109, N1113, N1045);
not NOT1 (N1205, N1189);
nor NOR4 (N1206, N1199, N1121, N956, N100);
buf BUF1 (N1207, N1205);
buf BUF1 (N1208, N1185);
not NOT1 (N1209, N1202);
buf BUF1 (N1210, N1201);
nand NAND4 (N1211, N1206, N373, N911, N35);
or OR2 (N1212, N1210, N930);
or OR4 (N1213, N1209, N1195, N747, N347);
buf BUF1 (N1214, N1213);
or OR3 (N1215, N1203, N80, N781);
or OR2 (N1216, N1200, N834);
and AND3 (N1217, N1215, N748, N813);
and AND2 (N1218, N1197, N35);
nand NAND4 (N1219, N1218, N306, N995, N957);
and AND4 (N1220, N1208, N113, N87, N288);
nor NOR3 (N1221, N1211, N345, N289);
nand NAND2 (N1222, N1217, N254);
buf BUF1 (N1223, N1221);
not NOT1 (N1224, N1204);
nand NAND4 (N1225, N1188, N191, N707, N397);
xor XOR2 (N1226, N1224, N997);
buf BUF1 (N1227, N1207);
or OR2 (N1228, N1219, N203);
and AND4 (N1229, N1214, N663, N580, N248);
xor XOR2 (N1230, N1223, N1119);
not NOT1 (N1231, N1230);
and AND2 (N1232, N1220, N374);
or OR4 (N1233, N1222, N116, N705, N63);
or OR2 (N1234, N1226, N717);
nand NAND3 (N1235, N1234, N889, N115);
not NOT1 (N1236, N1233);
xor XOR2 (N1237, N1236, N542);
or OR3 (N1238, N1228, N547, N522);
nand NAND2 (N1239, N1232, N1021);
or OR2 (N1240, N1237, N1173);
nand NAND4 (N1241, N1229, N976, N503, N463);
and AND2 (N1242, N1238, N1177);
or OR2 (N1243, N1225, N311);
or OR3 (N1244, N1240, N127, N775);
or OR4 (N1245, N1242, N149, N280, N981);
not NOT1 (N1246, N1243);
not NOT1 (N1247, N1245);
or OR3 (N1248, N1246, N211, N504);
xor XOR2 (N1249, N1212, N627);
buf BUF1 (N1250, N1231);
buf BUF1 (N1251, N1250);
not NOT1 (N1252, N1251);
and AND2 (N1253, N1227, N1012);
or OR3 (N1254, N1247, N986, N968);
buf BUF1 (N1255, N1254);
nor NOR2 (N1256, N1235, N893);
and AND4 (N1257, N1252, N1134, N528, N98);
nand NAND3 (N1258, N1244, N614, N675);
not NOT1 (N1259, N1255);
nor NOR4 (N1260, N1249, N1225, N887, N309);
nor NOR4 (N1261, N1239, N938, N1145, N70);
buf BUF1 (N1262, N1241);
buf BUF1 (N1263, N1256);
and AND3 (N1264, N1257, N531, N1083);
nand NAND2 (N1265, N1264, N725);
not NOT1 (N1266, N1216);
not NOT1 (N1267, N1266);
or OR3 (N1268, N1260, N1174, N371);
not NOT1 (N1269, N1261);
nor NOR2 (N1270, N1268, N473);
nor NOR4 (N1271, N1270, N211, N235, N1162);
or OR4 (N1272, N1253, N110, N364, N1158);
not NOT1 (N1273, N1259);
and AND3 (N1274, N1265, N899, N1079);
nor NOR2 (N1275, N1269, N537);
nand NAND4 (N1276, N1248, N195, N464, N140);
xor XOR2 (N1277, N1267, N378);
and AND4 (N1278, N1263, N931, N1104, N540);
nand NAND3 (N1279, N1278, N912, N978);
xor XOR2 (N1280, N1272, N1117);
nand NAND3 (N1281, N1275, N147, N144);
xor XOR2 (N1282, N1277, N1136);
nor NOR2 (N1283, N1276, N983);
or OR3 (N1284, N1258, N740, N117);
or OR2 (N1285, N1271, N997);
nand NAND4 (N1286, N1285, N1087, N688, N1238);
nand NAND4 (N1287, N1283, N409, N726, N786);
nor NOR4 (N1288, N1279, N113, N540, N1140);
nand NAND3 (N1289, N1287, N305, N143);
and AND4 (N1290, N1286, N17, N782, N903);
xor XOR2 (N1291, N1262, N615);
or OR3 (N1292, N1274, N710, N1109);
xor XOR2 (N1293, N1282, N171);
nor NOR2 (N1294, N1281, N792);
nor NOR4 (N1295, N1280, N690, N533, N359);
or OR2 (N1296, N1293, N974);
not NOT1 (N1297, N1273);
or OR2 (N1298, N1294, N1074);
nor NOR3 (N1299, N1289, N999, N106);
not NOT1 (N1300, N1288);
buf BUF1 (N1301, N1284);
nand NAND3 (N1302, N1296, N96, N355);
not NOT1 (N1303, N1290);
and AND4 (N1304, N1299, N578, N819, N484);
buf BUF1 (N1305, N1291);
xor XOR2 (N1306, N1301, N713);
buf BUF1 (N1307, N1295);
or OR4 (N1308, N1307, N24, N734, N73);
or OR4 (N1309, N1300, N1185, N81, N902);
nor NOR3 (N1310, N1298, N955, N665);
and AND2 (N1311, N1303, N537);
buf BUF1 (N1312, N1306);
and AND4 (N1313, N1292, N1278, N867, N149);
not NOT1 (N1314, N1308);
nand NAND2 (N1315, N1302, N32);
and AND4 (N1316, N1312, N109, N774, N758);
or OR2 (N1317, N1305, N867);
and AND2 (N1318, N1310, N1209);
not NOT1 (N1319, N1315);
buf BUF1 (N1320, N1309);
or OR4 (N1321, N1313, N465, N892, N926);
nor NOR4 (N1322, N1311, N735, N1043, N942);
not NOT1 (N1323, N1317);
and AND2 (N1324, N1319, N444);
and AND3 (N1325, N1314, N644, N936);
nor NOR4 (N1326, N1320, N529, N388, N427);
or OR4 (N1327, N1325, N103, N92, N690);
nor NOR4 (N1328, N1304, N211, N1039, N1316);
nand NAND3 (N1329, N642, N235, N979);
xor XOR2 (N1330, N1324, N199);
buf BUF1 (N1331, N1330);
or OR2 (N1332, N1331, N761);
xor XOR2 (N1333, N1326, N1220);
nand NAND2 (N1334, N1323, N1266);
nand NAND4 (N1335, N1328, N559, N285, N709);
and AND4 (N1336, N1297, N761, N44, N1314);
xor XOR2 (N1337, N1329, N1241);
and AND3 (N1338, N1336, N588, N1071);
and AND2 (N1339, N1322, N123);
nand NAND2 (N1340, N1333, N1248);
nand NAND4 (N1341, N1327, N64, N508, N915);
and AND4 (N1342, N1341, N632, N108, N524);
xor XOR2 (N1343, N1340, N122);
buf BUF1 (N1344, N1335);
or OR3 (N1345, N1344, N1276, N1102);
nand NAND4 (N1346, N1343, N377, N759, N998);
not NOT1 (N1347, N1346);
nor NOR3 (N1348, N1334, N601, N1030);
or OR3 (N1349, N1345, N1266, N1093);
and AND4 (N1350, N1337, N809, N879, N208);
xor XOR2 (N1351, N1347, N421);
xor XOR2 (N1352, N1349, N678);
and AND3 (N1353, N1352, N795, N106);
nand NAND2 (N1354, N1332, N308);
or OR4 (N1355, N1318, N705, N372, N914);
and AND2 (N1356, N1339, N1129);
and AND2 (N1357, N1350, N359);
buf BUF1 (N1358, N1321);
or OR2 (N1359, N1356, N449);
and AND4 (N1360, N1351, N818, N22, N1260);
nand NAND2 (N1361, N1357, N1121);
or OR3 (N1362, N1348, N132, N1266);
not NOT1 (N1363, N1353);
nand NAND4 (N1364, N1342, N735, N1255, N666);
not NOT1 (N1365, N1363);
not NOT1 (N1366, N1361);
or OR4 (N1367, N1365, N13, N1322, N290);
or OR2 (N1368, N1338, N347);
nor NOR3 (N1369, N1364, N1259, N200);
nand NAND2 (N1370, N1368, N249);
nor NOR3 (N1371, N1359, N155, N814);
and AND3 (N1372, N1354, N1283, N1016);
or OR2 (N1373, N1367, N1149);
buf BUF1 (N1374, N1373);
and AND2 (N1375, N1362, N644);
nor NOR2 (N1376, N1355, N295);
xor XOR2 (N1377, N1358, N61);
nor NOR3 (N1378, N1376, N947, N1227);
not NOT1 (N1379, N1372);
buf BUF1 (N1380, N1360);
buf BUF1 (N1381, N1375);
xor XOR2 (N1382, N1366, N746);
or OR2 (N1383, N1381, N276);
not NOT1 (N1384, N1370);
buf BUF1 (N1385, N1378);
nand NAND4 (N1386, N1374, N185, N360, N774);
buf BUF1 (N1387, N1386);
buf BUF1 (N1388, N1383);
not NOT1 (N1389, N1385);
or OR2 (N1390, N1377, N1105);
buf BUF1 (N1391, N1384);
or OR2 (N1392, N1382, N917);
and AND3 (N1393, N1369, N71, N352);
buf BUF1 (N1394, N1371);
or OR3 (N1395, N1392, N762, N1343);
nand NAND4 (N1396, N1393, N12, N806, N784);
nor NOR4 (N1397, N1394, N1103, N851, N1250);
nand NAND4 (N1398, N1396, N1119, N797, N887);
buf BUF1 (N1399, N1387);
nand NAND2 (N1400, N1391, N596);
nand NAND3 (N1401, N1400, N242, N647);
not NOT1 (N1402, N1390);
and AND3 (N1403, N1380, N426, N1044);
xor XOR2 (N1404, N1389, N114);
and AND3 (N1405, N1379, N1167, N1139);
xor XOR2 (N1406, N1401, N913);
or OR4 (N1407, N1406, N1226, N156, N883);
buf BUF1 (N1408, N1398);
and AND2 (N1409, N1408, N64);
not NOT1 (N1410, N1403);
not NOT1 (N1411, N1402);
not NOT1 (N1412, N1411);
xor XOR2 (N1413, N1410, N449);
nand NAND4 (N1414, N1412, N810, N537, N801);
or OR2 (N1415, N1407, N373);
xor XOR2 (N1416, N1409, N322);
and AND2 (N1417, N1388, N1302);
not NOT1 (N1418, N1397);
buf BUF1 (N1419, N1414);
buf BUF1 (N1420, N1417);
or OR4 (N1421, N1420, N628, N734, N787);
and AND3 (N1422, N1416, N126, N63);
and AND2 (N1423, N1395, N993);
xor XOR2 (N1424, N1405, N748);
xor XOR2 (N1425, N1413, N1226);
buf BUF1 (N1426, N1421);
buf BUF1 (N1427, N1425);
nor NOR3 (N1428, N1427, N198, N755);
nand NAND3 (N1429, N1418, N1138, N8);
xor XOR2 (N1430, N1424, N411);
xor XOR2 (N1431, N1428, N1164);
or OR3 (N1432, N1423, N1021, N218);
buf BUF1 (N1433, N1415);
not NOT1 (N1434, N1422);
nor NOR2 (N1435, N1432, N138);
not NOT1 (N1436, N1430);
nor NOR2 (N1437, N1399, N1429);
and AND4 (N1438, N30, N1018, N1322, N739);
buf BUF1 (N1439, N1436);
not NOT1 (N1440, N1438);
nor NOR3 (N1441, N1434, N18, N1155);
or OR3 (N1442, N1433, N428, N154);
buf BUF1 (N1443, N1439);
or OR3 (N1444, N1440, N768, N440);
buf BUF1 (N1445, N1404);
nand NAND3 (N1446, N1437, N997, N71);
not NOT1 (N1447, N1441);
nand NAND3 (N1448, N1419, N1275, N67);
not NOT1 (N1449, N1444);
nor NOR4 (N1450, N1447, N969, N909, N471);
or OR3 (N1451, N1445, N411, N1414);
and AND2 (N1452, N1450, N320);
or OR3 (N1453, N1448, N1203, N460);
nor NOR3 (N1454, N1435, N167, N958);
xor XOR2 (N1455, N1443, N1192);
not NOT1 (N1456, N1446);
nand NAND2 (N1457, N1456, N199);
nand NAND3 (N1458, N1442, N1408, N624);
or OR3 (N1459, N1455, N720, N484);
nor NOR4 (N1460, N1431, N1188, N878, N1345);
nand NAND2 (N1461, N1460, N939);
not NOT1 (N1462, N1452);
or OR3 (N1463, N1459, N978, N833);
xor XOR2 (N1464, N1451, N501);
nor NOR3 (N1465, N1462, N288, N656);
xor XOR2 (N1466, N1454, N1292);
nand NAND4 (N1467, N1449, N1244, N487, N822);
or OR4 (N1468, N1458, N437, N1401, N1365);
buf BUF1 (N1469, N1466);
nand NAND3 (N1470, N1426, N337, N591);
buf BUF1 (N1471, N1464);
nand NAND2 (N1472, N1471, N233);
or OR2 (N1473, N1453, N666);
or OR2 (N1474, N1465, N403);
not NOT1 (N1475, N1467);
buf BUF1 (N1476, N1470);
nand NAND2 (N1477, N1469, N49);
not NOT1 (N1478, N1474);
xor XOR2 (N1479, N1476, N290);
buf BUF1 (N1480, N1457);
nand NAND3 (N1481, N1461, N413, N227);
nand NAND2 (N1482, N1463, N210);
nand NAND2 (N1483, N1481, N1057);
buf BUF1 (N1484, N1473);
nand NAND3 (N1485, N1478, N102, N70);
not NOT1 (N1486, N1479);
nor NOR2 (N1487, N1475, N386);
xor XOR2 (N1488, N1483, N1345);
nor NOR2 (N1489, N1477, N889);
nor NOR4 (N1490, N1482, N320, N1118, N1223);
nand NAND2 (N1491, N1468, N1386);
nand NAND3 (N1492, N1486, N901, N1241);
nand NAND2 (N1493, N1472, N956);
and AND3 (N1494, N1480, N1065, N1140);
or OR2 (N1495, N1492, N43);
xor XOR2 (N1496, N1485, N882);
nand NAND3 (N1497, N1487, N1355, N1480);
or OR3 (N1498, N1496, N444, N1097);
nor NOR3 (N1499, N1489, N674, N1245);
or OR2 (N1500, N1493, N55);
and AND3 (N1501, N1484, N735, N1234);
nand NAND4 (N1502, N1488, N821, N701, N884);
nand NAND2 (N1503, N1491, N494);
not NOT1 (N1504, N1500);
and AND4 (N1505, N1504, N1448, N622, N963);
xor XOR2 (N1506, N1502, N653);
or OR3 (N1507, N1499, N1110, N1294);
xor XOR2 (N1508, N1507, N1418);
or OR4 (N1509, N1497, N1234, N626, N863);
not NOT1 (N1510, N1498);
endmodule