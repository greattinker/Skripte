// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N3523,N3515,N3519,N3513,N3503,N3521,N3514,N3491,N3518,N3524;

nand NAND3 (N25, N22, N21, N3);
nand NAND2 (N26, N11, N25);
not NOT1 (N27, N12);
or OR3 (N28, N13, N3, N5);
nor NOR2 (N29, N5, N13);
nor NOR3 (N30, N9, N3, N7);
nand NAND3 (N31, N21, N24, N19);
xor XOR2 (N32, N14, N22);
nor NOR3 (N33, N14, N16, N7);
buf BUF1 (N34, N19);
and AND4 (N35, N15, N31, N13, N5);
or OR2 (N36, N20, N7);
buf BUF1 (N37, N26);
nand NAND3 (N38, N29, N22, N31);
not NOT1 (N39, N27);
nor NOR3 (N40, N36, N28, N28);
nor NOR2 (N41, N17, N34);
and AND4 (N42, N28, N23, N19, N30);
and AND4 (N43, N13, N7, N23, N33);
nor NOR4 (N44, N2, N22, N5, N28);
xor XOR2 (N45, N44, N22);
nor NOR2 (N46, N40, N9);
not NOT1 (N47, N41);
nand NAND3 (N48, N32, N44, N7);
or OR4 (N49, N45, N15, N26, N19);
and AND4 (N50, N48, N11, N10, N30);
xor XOR2 (N51, N38, N26);
nor NOR3 (N52, N50, N51, N50);
buf BUF1 (N53, N51);
and AND4 (N54, N43, N5, N42, N21);
not NOT1 (N55, N26);
nor NOR2 (N56, N54, N1);
nand NAND3 (N57, N46, N42, N34);
nor NOR2 (N58, N53, N17);
xor XOR2 (N59, N47, N11);
and AND2 (N60, N59, N33);
buf BUF1 (N61, N55);
or OR2 (N62, N60, N36);
buf BUF1 (N63, N39);
xor XOR2 (N64, N49, N12);
nor NOR4 (N65, N61, N10, N49, N34);
not NOT1 (N66, N52);
buf BUF1 (N67, N56);
xor XOR2 (N68, N65, N6);
not NOT1 (N69, N37);
buf BUF1 (N70, N57);
not NOT1 (N71, N64);
and AND2 (N72, N71, N45);
or OR4 (N73, N58, N64, N34, N50);
not NOT1 (N74, N66);
buf BUF1 (N75, N63);
xor XOR2 (N76, N62, N12);
buf BUF1 (N77, N73);
xor XOR2 (N78, N75, N33);
or OR3 (N79, N78, N51, N40);
nand NAND3 (N80, N72, N6, N30);
or OR3 (N81, N35, N72, N73);
or OR3 (N82, N80, N26, N23);
and AND2 (N83, N67, N72);
xor XOR2 (N84, N74, N36);
or OR3 (N85, N83, N68, N26);
not NOT1 (N86, N77);
not NOT1 (N87, N38);
xor XOR2 (N88, N70, N21);
buf BUF1 (N89, N82);
nor NOR2 (N90, N86, N59);
and AND2 (N91, N69, N20);
and AND3 (N92, N90, N45, N46);
and AND4 (N93, N91, N38, N55, N70);
buf BUF1 (N94, N92);
or OR2 (N95, N76, N50);
xor XOR2 (N96, N89, N72);
nor NOR4 (N97, N79, N34, N48, N52);
nor NOR2 (N98, N97, N14);
nor NOR3 (N99, N81, N21, N51);
not NOT1 (N100, N96);
nand NAND4 (N101, N100, N25, N47, N64);
buf BUF1 (N102, N84);
and AND2 (N103, N88, N62);
and AND4 (N104, N98, N23, N92, N56);
nand NAND2 (N105, N104, N27);
and AND2 (N106, N105, N23);
not NOT1 (N107, N93);
not NOT1 (N108, N85);
nor NOR2 (N109, N108, N46);
or OR4 (N110, N106, N63, N10, N2);
xor XOR2 (N111, N102, N48);
nor NOR2 (N112, N87, N26);
buf BUF1 (N113, N94);
xor XOR2 (N114, N110, N113);
not NOT1 (N115, N20);
nor NOR2 (N116, N101, N3);
buf BUF1 (N117, N111);
and AND3 (N118, N117, N31, N60);
nor NOR3 (N119, N112, N48, N108);
nand NAND2 (N120, N118, N37);
nand NAND4 (N121, N109, N84, N22, N24);
not NOT1 (N122, N116);
not NOT1 (N123, N121);
buf BUF1 (N124, N123);
xor XOR2 (N125, N119, N54);
buf BUF1 (N126, N124);
buf BUF1 (N127, N126);
nand NAND2 (N128, N115, N63);
not NOT1 (N129, N114);
nor NOR3 (N130, N95, N102, N124);
buf BUF1 (N131, N130);
nand NAND2 (N132, N122, N51);
buf BUF1 (N133, N132);
and AND2 (N134, N107, N63);
nor NOR2 (N135, N127, N57);
nor NOR2 (N136, N128, N74);
nand NAND3 (N137, N120, N34, N111);
buf BUF1 (N138, N103);
nor NOR2 (N139, N134, N128);
buf BUF1 (N140, N136);
not NOT1 (N141, N133);
or OR3 (N142, N138, N84, N124);
nand NAND3 (N143, N137, N4, N72);
buf BUF1 (N144, N139);
nor NOR3 (N145, N141, N72, N23);
not NOT1 (N146, N99);
not NOT1 (N147, N135);
and AND4 (N148, N145, N38, N87, N108);
not NOT1 (N149, N143);
xor XOR2 (N150, N142, N36);
and AND2 (N151, N149, N37);
or OR2 (N152, N150, N73);
xor XOR2 (N153, N147, N5);
nor NOR4 (N154, N153, N93, N138, N99);
and AND3 (N155, N125, N144, N84);
nor NOR3 (N156, N21, N88, N19);
not NOT1 (N157, N152);
and AND4 (N158, N151, N23, N142, N47);
buf BUF1 (N159, N155);
xor XOR2 (N160, N140, N56);
and AND2 (N161, N129, N11);
buf BUF1 (N162, N156);
xor XOR2 (N163, N160, N49);
nand NAND3 (N164, N161, N25, N24);
not NOT1 (N165, N159);
nand NAND2 (N166, N148, N65);
buf BUF1 (N167, N157);
xor XOR2 (N168, N164, N151);
nand NAND4 (N169, N163, N123, N151, N15);
and AND2 (N170, N167, N82);
nand NAND4 (N171, N170, N110, N56, N15);
xor XOR2 (N172, N165, N83);
xor XOR2 (N173, N162, N38);
nor NOR4 (N174, N172, N90, N117, N70);
nor NOR4 (N175, N158, N47, N144, N138);
nor NOR3 (N176, N171, N19, N46);
or OR4 (N177, N168, N65, N89, N171);
xor XOR2 (N178, N174, N142);
buf BUF1 (N179, N166);
not NOT1 (N180, N169);
not NOT1 (N181, N146);
not NOT1 (N182, N178);
or OR4 (N183, N173, N107, N31, N84);
not NOT1 (N184, N179);
not NOT1 (N185, N175);
not NOT1 (N186, N177);
xor XOR2 (N187, N184, N69);
and AND2 (N188, N187, N183);
xor XOR2 (N189, N26, N146);
not NOT1 (N190, N176);
nor NOR4 (N191, N131, N91, N72, N12);
and AND4 (N192, N186, N143, N140, N94);
and AND3 (N193, N154, N16, N140);
xor XOR2 (N194, N188, N7);
buf BUF1 (N195, N182);
nor NOR3 (N196, N185, N158, N71);
nor NOR3 (N197, N180, N43, N89);
not NOT1 (N198, N191);
and AND3 (N199, N193, N145, N101);
xor XOR2 (N200, N199, N147);
nor NOR2 (N201, N200, N130);
and AND4 (N202, N189, N69, N87, N163);
buf BUF1 (N203, N181);
xor XOR2 (N204, N195, N69);
nand NAND2 (N205, N192, N61);
nand NAND3 (N206, N203, N137, N55);
not NOT1 (N207, N198);
xor XOR2 (N208, N204, N109);
buf BUF1 (N209, N197);
or OR4 (N210, N201, N152, N61, N139);
and AND2 (N211, N206, N196);
buf BUF1 (N212, N74);
buf BUF1 (N213, N210);
and AND4 (N214, N213, N95, N174, N23);
nand NAND3 (N215, N214, N73, N206);
buf BUF1 (N216, N208);
or OR2 (N217, N209, N169);
xor XOR2 (N218, N215, N148);
buf BUF1 (N219, N190);
buf BUF1 (N220, N219);
nand NAND3 (N221, N220, N31, N218);
and AND4 (N222, N10, N71, N197, N40);
not NOT1 (N223, N205);
or OR3 (N224, N223, N38, N24);
buf BUF1 (N225, N212);
buf BUF1 (N226, N194);
buf BUF1 (N227, N225);
buf BUF1 (N228, N207);
buf BUF1 (N229, N221);
and AND4 (N230, N216, N51, N114, N63);
and AND2 (N231, N222, N66);
nand NAND4 (N232, N227, N58, N211, N22);
not NOT1 (N233, N215);
buf BUF1 (N234, N202);
xor XOR2 (N235, N226, N231);
nand NAND4 (N236, N12, N82, N136, N23);
xor XOR2 (N237, N217, N22);
and AND3 (N238, N235, N103, N28);
not NOT1 (N239, N232);
nand NAND4 (N240, N224, N179, N142, N228);
nor NOR2 (N241, N116, N198);
buf BUF1 (N242, N239);
xor XOR2 (N243, N236, N183);
nor NOR2 (N244, N230, N25);
buf BUF1 (N245, N234);
xor XOR2 (N246, N245, N133);
or OR4 (N247, N244, N45, N73, N206);
and AND2 (N248, N233, N20);
and AND3 (N249, N243, N174, N128);
or OR4 (N250, N247, N120, N37, N239);
not NOT1 (N251, N248);
nor NOR3 (N252, N250, N153, N195);
nand NAND3 (N253, N237, N2, N71);
xor XOR2 (N254, N229, N250);
or OR3 (N255, N249, N107, N203);
nor NOR2 (N256, N238, N105);
and AND3 (N257, N242, N49, N109);
nand NAND3 (N258, N246, N16, N43);
not NOT1 (N259, N253);
not NOT1 (N260, N256);
and AND2 (N261, N259, N176);
or OR3 (N262, N257, N99, N176);
not NOT1 (N263, N254);
xor XOR2 (N264, N251, N54);
xor XOR2 (N265, N258, N66);
xor XOR2 (N266, N263, N158);
buf BUF1 (N267, N265);
and AND2 (N268, N267, N67);
or OR2 (N269, N262, N132);
buf BUF1 (N270, N261);
xor XOR2 (N271, N266, N14);
or OR3 (N272, N264, N35, N258);
buf BUF1 (N273, N255);
nor NOR4 (N274, N271, N271, N104, N46);
not NOT1 (N275, N252);
not NOT1 (N276, N241);
xor XOR2 (N277, N270, N43);
not NOT1 (N278, N277);
not NOT1 (N279, N260);
buf BUF1 (N280, N275);
or OR4 (N281, N280, N214, N123, N123);
and AND4 (N282, N240, N218, N49, N7);
xor XOR2 (N283, N268, N19);
or OR4 (N284, N283, N135, N51, N266);
xor XOR2 (N285, N273, N225);
or OR3 (N286, N272, N31, N227);
not NOT1 (N287, N269);
xor XOR2 (N288, N281, N269);
nor NOR4 (N289, N284, N39, N71, N7);
or OR4 (N290, N286, N128, N280, N24);
or OR4 (N291, N287, N108, N60, N99);
and AND2 (N292, N291, N163);
nor NOR2 (N293, N279, N31);
buf BUF1 (N294, N293);
not NOT1 (N295, N292);
nor NOR4 (N296, N295, N138, N124, N169);
xor XOR2 (N297, N278, N144);
nand NAND2 (N298, N282, N61);
nor NOR2 (N299, N294, N133);
and AND3 (N300, N299, N254, N21);
xor XOR2 (N301, N290, N221);
and AND2 (N302, N298, N197);
nor NOR4 (N303, N288, N150, N90, N267);
not NOT1 (N304, N303);
nor NOR4 (N305, N297, N244, N237, N182);
not NOT1 (N306, N285);
buf BUF1 (N307, N302);
not NOT1 (N308, N305);
xor XOR2 (N309, N307, N103);
or OR2 (N310, N276, N263);
buf BUF1 (N311, N289);
nand NAND4 (N312, N311, N263, N232, N236);
xor XOR2 (N313, N309, N75);
nor NOR3 (N314, N300, N299, N187);
buf BUF1 (N315, N310);
buf BUF1 (N316, N301);
or OR4 (N317, N296, N261, N13, N250);
nor NOR4 (N318, N316, N158, N269, N200);
nor NOR2 (N319, N315, N80);
buf BUF1 (N320, N317);
nand NAND4 (N321, N318, N306, N108, N88);
or OR4 (N322, N283, N229, N310, N125);
xor XOR2 (N323, N321, N87);
buf BUF1 (N324, N314);
not NOT1 (N325, N324);
not NOT1 (N326, N313);
and AND4 (N327, N312, N153, N98, N222);
not NOT1 (N328, N322);
buf BUF1 (N329, N328);
buf BUF1 (N330, N320);
and AND4 (N331, N325, N292, N72, N157);
and AND4 (N332, N323, N12, N208, N82);
xor XOR2 (N333, N332, N281);
xor XOR2 (N334, N331, N91);
xor XOR2 (N335, N334, N271);
and AND3 (N336, N333, N211, N210);
and AND4 (N337, N330, N302, N198, N162);
and AND4 (N338, N274, N89, N284, N114);
not NOT1 (N339, N338);
nor NOR2 (N340, N339, N13);
buf BUF1 (N341, N308);
xor XOR2 (N342, N327, N41);
and AND2 (N343, N326, N93);
buf BUF1 (N344, N336);
and AND2 (N345, N337, N69);
nor NOR3 (N346, N343, N332, N76);
and AND2 (N347, N329, N341);
xor XOR2 (N348, N53, N203);
buf BUF1 (N349, N304);
not NOT1 (N350, N335);
nor NOR4 (N351, N346, N280, N269, N144);
or OR4 (N352, N350, N79, N108, N195);
and AND3 (N353, N351, N91, N244);
xor XOR2 (N354, N345, N154);
nand NAND2 (N355, N342, N66);
nor NOR4 (N356, N352, N124, N164, N36);
not NOT1 (N357, N340);
not NOT1 (N358, N357);
not NOT1 (N359, N353);
and AND4 (N360, N344, N265, N15, N45);
nand NAND2 (N361, N348, N108);
and AND4 (N362, N359, N359, N219, N57);
not NOT1 (N363, N356);
buf BUF1 (N364, N358);
buf BUF1 (N365, N347);
nand NAND2 (N366, N365, N47);
buf BUF1 (N367, N361);
xor XOR2 (N368, N366, N244);
nand NAND2 (N369, N364, N312);
and AND4 (N370, N355, N173, N141, N78);
nand NAND3 (N371, N354, N43, N50);
nor NOR2 (N372, N371, N370);
not NOT1 (N373, N268);
nand NAND2 (N374, N349, N132);
not NOT1 (N375, N374);
not NOT1 (N376, N368);
nand NAND4 (N377, N362, N76, N105, N167);
nand NAND4 (N378, N376, N180, N103, N92);
and AND2 (N379, N372, N238);
buf BUF1 (N380, N378);
nand NAND3 (N381, N367, N145, N23);
xor XOR2 (N382, N369, N130);
and AND3 (N383, N380, N129, N316);
not NOT1 (N384, N381);
xor XOR2 (N385, N383, N177);
nand NAND3 (N386, N363, N119, N322);
nor NOR3 (N387, N386, N34, N251);
xor XOR2 (N388, N379, N138);
xor XOR2 (N389, N388, N311);
buf BUF1 (N390, N384);
xor XOR2 (N391, N390, N341);
or OR2 (N392, N391, N154);
nor NOR2 (N393, N377, N10);
xor XOR2 (N394, N382, N175);
and AND3 (N395, N375, N365, N182);
nor NOR3 (N396, N395, N252, N383);
or OR2 (N397, N394, N112);
nor NOR4 (N398, N385, N261, N206, N10);
xor XOR2 (N399, N398, N102);
buf BUF1 (N400, N397);
xor XOR2 (N401, N373, N33);
or OR3 (N402, N396, N139, N279);
nand NAND2 (N403, N392, N370);
nor NOR2 (N404, N387, N111);
not NOT1 (N405, N404);
or OR4 (N406, N393, N144, N342, N380);
and AND3 (N407, N401, N388, N193);
nand NAND2 (N408, N399, N256);
not NOT1 (N409, N360);
or OR3 (N410, N409, N238, N223);
nor NOR4 (N411, N407, N245, N62, N290);
xor XOR2 (N412, N411, N109);
buf BUF1 (N413, N319);
and AND3 (N414, N402, N216, N128);
or OR4 (N415, N405, N174, N183, N339);
buf BUF1 (N416, N406);
nor NOR2 (N417, N415, N393);
not NOT1 (N418, N412);
xor XOR2 (N419, N389, N115);
or OR4 (N420, N408, N86, N222, N309);
xor XOR2 (N421, N420, N176);
or OR2 (N422, N413, N209);
and AND2 (N423, N421, N292);
nand NAND4 (N424, N414, N80, N174, N402);
not NOT1 (N425, N410);
nor NOR2 (N426, N417, N416);
and AND3 (N427, N160, N238, N163);
xor XOR2 (N428, N427, N405);
nand NAND2 (N429, N422, N48);
and AND4 (N430, N428, N14, N206, N295);
or OR4 (N431, N426, N393, N282, N382);
buf BUF1 (N432, N400);
buf BUF1 (N433, N423);
nor NOR3 (N434, N429, N84, N425);
xor XOR2 (N435, N425, N223);
xor XOR2 (N436, N432, N183);
buf BUF1 (N437, N430);
nor NOR3 (N438, N433, N48, N261);
and AND4 (N439, N419, N120, N429, N355);
or OR4 (N440, N439, N283, N261, N68);
xor XOR2 (N441, N424, N52);
nand NAND3 (N442, N441, N74, N79);
buf BUF1 (N443, N436);
and AND4 (N444, N418, N30, N231, N358);
not NOT1 (N445, N438);
and AND2 (N446, N443, N197);
nor NOR3 (N447, N445, N27, N183);
nor NOR2 (N448, N437, N161);
nand NAND2 (N449, N434, N164);
nand NAND2 (N450, N448, N271);
xor XOR2 (N451, N431, N116);
nand NAND4 (N452, N442, N234, N75, N125);
and AND4 (N453, N449, N92, N373, N234);
nor NOR3 (N454, N447, N277, N227);
not NOT1 (N455, N452);
or OR4 (N456, N453, N326, N428, N26);
and AND3 (N457, N455, N293, N282);
buf BUF1 (N458, N440);
not NOT1 (N459, N451);
nand NAND4 (N460, N446, N225, N365, N98);
buf BUF1 (N461, N444);
buf BUF1 (N462, N435);
and AND4 (N463, N462, N111, N274, N18);
nand NAND2 (N464, N459, N323);
xor XOR2 (N465, N456, N101);
nor NOR2 (N466, N460, N362);
not NOT1 (N467, N465);
or OR3 (N468, N454, N382, N140);
or OR3 (N469, N464, N441, N112);
or OR3 (N470, N458, N168, N259);
buf BUF1 (N471, N470);
buf BUF1 (N472, N403);
not NOT1 (N473, N469);
and AND3 (N474, N457, N258, N206);
and AND3 (N475, N450, N129, N266);
xor XOR2 (N476, N466, N243);
nor NOR2 (N477, N461, N445);
not NOT1 (N478, N476);
or OR3 (N479, N472, N294, N472);
xor XOR2 (N480, N474, N212);
xor XOR2 (N481, N463, N124);
or OR3 (N482, N478, N47, N299);
buf BUF1 (N483, N482);
or OR2 (N484, N473, N261);
xor XOR2 (N485, N484, N106);
nor NOR2 (N486, N480, N478);
xor XOR2 (N487, N471, N175);
buf BUF1 (N488, N481);
xor XOR2 (N489, N467, N200);
or OR4 (N490, N477, N8, N195, N181);
nor NOR3 (N491, N488, N116, N101);
buf BUF1 (N492, N479);
xor XOR2 (N493, N490, N149);
buf BUF1 (N494, N493);
not NOT1 (N495, N492);
nor NOR4 (N496, N495, N337, N375, N295);
nand NAND2 (N497, N496, N351);
or OR4 (N498, N468, N379, N351, N146);
nor NOR3 (N499, N491, N183, N393);
buf BUF1 (N500, N498);
not NOT1 (N501, N500);
nand NAND4 (N502, N475, N122, N132, N202);
nor NOR3 (N503, N485, N361, N451);
nand NAND2 (N504, N487, N53);
nand NAND2 (N505, N483, N31);
nor NOR4 (N506, N503, N190, N28, N109);
nor NOR4 (N507, N497, N83, N319, N415);
and AND4 (N508, N494, N271, N214, N269);
and AND3 (N509, N501, N3, N503);
xor XOR2 (N510, N486, N59);
or OR2 (N511, N510, N454);
or OR3 (N512, N505, N474, N50);
xor XOR2 (N513, N512, N406);
buf BUF1 (N514, N507);
buf BUF1 (N515, N499);
and AND2 (N516, N509, N515);
xor XOR2 (N517, N446, N198);
not NOT1 (N518, N513);
nor NOR2 (N519, N489, N269);
or OR3 (N520, N516, N291, N77);
xor XOR2 (N521, N517, N291);
buf BUF1 (N522, N521);
nand NAND2 (N523, N502, N320);
nor NOR3 (N524, N508, N336, N240);
buf BUF1 (N525, N518);
xor XOR2 (N526, N514, N179);
not NOT1 (N527, N519);
xor XOR2 (N528, N511, N14);
xor XOR2 (N529, N522, N62);
nand NAND4 (N530, N529, N346, N347, N3);
xor XOR2 (N531, N520, N97);
nor NOR3 (N532, N524, N157, N260);
and AND2 (N533, N525, N339);
nand NAND3 (N534, N526, N158, N347);
and AND3 (N535, N504, N457, N353);
and AND3 (N536, N527, N98, N114);
and AND3 (N537, N506, N28, N99);
and AND2 (N538, N533, N307);
nand NAND4 (N539, N534, N261, N380, N127);
not NOT1 (N540, N532);
xor XOR2 (N541, N537, N361);
nor NOR3 (N542, N540, N386, N276);
and AND2 (N543, N541, N234);
xor XOR2 (N544, N531, N241);
nand NAND3 (N545, N528, N322, N255);
nand NAND2 (N546, N539, N158);
nor NOR3 (N547, N544, N464, N280);
or OR4 (N548, N545, N215, N55, N514);
buf BUF1 (N549, N523);
and AND3 (N550, N536, N211, N530);
or OR2 (N551, N40, N125);
nor NOR3 (N552, N543, N472, N216);
xor XOR2 (N553, N546, N509);
not NOT1 (N554, N542);
nand NAND2 (N555, N552, N468);
or OR2 (N556, N553, N340);
nor NOR3 (N557, N538, N553, N183);
or OR2 (N558, N548, N331);
buf BUF1 (N559, N558);
nand NAND2 (N560, N551, N207);
buf BUF1 (N561, N549);
nand NAND2 (N562, N556, N493);
not NOT1 (N563, N561);
buf BUF1 (N564, N555);
nand NAND2 (N565, N563, N315);
nor NOR3 (N566, N535, N173, N52);
or OR3 (N567, N557, N59, N208);
or OR3 (N568, N554, N203, N461);
and AND2 (N569, N550, N267);
nor NOR4 (N570, N569, N172, N389, N170);
nor NOR3 (N571, N560, N447, N269);
or OR3 (N572, N559, N368, N537);
not NOT1 (N573, N571);
nor NOR2 (N574, N547, N402);
xor XOR2 (N575, N568, N324);
nor NOR4 (N576, N566, N195, N437, N78);
nand NAND3 (N577, N573, N500, N328);
not NOT1 (N578, N570);
nand NAND3 (N579, N567, N379, N402);
xor XOR2 (N580, N564, N161);
nor NOR2 (N581, N576, N421);
nor NOR2 (N582, N577, N374);
not NOT1 (N583, N575);
and AND2 (N584, N574, N282);
not NOT1 (N585, N578);
buf BUF1 (N586, N582);
and AND3 (N587, N581, N247, N159);
buf BUF1 (N588, N586);
nand NAND4 (N589, N572, N475, N265, N152);
nand NAND2 (N590, N565, N343);
not NOT1 (N591, N588);
buf BUF1 (N592, N583);
nand NAND4 (N593, N585, N285, N111, N15);
not NOT1 (N594, N592);
xor XOR2 (N595, N584, N568);
nand NAND4 (N596, N590, N484, N567, N161);
not NOT1 (N597, N587);
not NOT1 (N598, N595);
buf BUF1 (N599, N591);
or OR4 (N600, N579, N79, N89, N305);
xor XOR2 (N601, N594, N598);
nand NAND2 (N602, N226, N104);
nand NAND4 (N603, N596, N351, N216, N303);
and AND2 (N604, N601, N112);
not NOT1 (N605, N602);
buf BUF1 (N606, N593);
or OR3 (N607, N603, N521, N270);
and AND2 (N608, N580, N530);
not NOT1 (N609, N608);
xor XOR2 (N610, N606, N601);
nor NOR2 (N611, N609, N330);
nor NOR4 (N612, N611, N89, N440, N45);
nand NAND3 (N613, N600, N34, N465);
nor NOR2 (N614, N607, N255);
nor NOR3 (N615, N604, N62, N490);
nand NAND3 (N616, N599, N406, N498);
xor XOR2 (N617, N613, N378);
nand NAND2 (N618, N616, N227);
buf BUF1 (N619, N562);
nand NAND3 (N620, N612, N285, N398);
nand NAND2 (N621, N619, N393);
buf BUF1 (N622, N617);
nand NAND2 (N623, N618, N524);
and AND2 (N624, N615, N322);
nand NAND3 (N625, N622, N533, N465);
xor XOR2 (N626, N597, N559);
and AND4 (N627, N614, N262, N548, N287);
not NOT1 (N628, N626);
buf BUF1 (N629, N620);
buf BUF1 (N630, N621);
and AND2 (N631, N605, N306);
xor XOR2 (N632, N625, N464);
or OR3 (N633, N629, N420, N339);
and AND2 (N634, N628, N150);
nor NOR3 (N635, N631, N593, N77);
buf BUF1 (N636, N624);
nor NOR3 (N637, N610, N413, N236);
xor XOR2 (N638, N632, N38);
xor XOR2 (N639, N635, N164);
or OR4 (N640, N637, N133, N133, N226);
not NOT1 (N641, N633);
nor NOR4 (N642, N634, N53, N294, N514);
nand NAND3 (N643, N589, N222, N65);
nor NOR2 (N644, N642, N241);
xor XOR2 (N645, N641, N570);
and AND2 (N646, N630, N443);
xor XOR2 (N647, N645, N290);
buf BUF1 (N648, N623);
nor NOR2 (N649, N643, N306);
nor NOR4 (N650, N639, N477, N573, N253);
or OR2 (N651, N638, N231);
buf BUF1 (N652, N640);
and AND4 (N653, N651, N609, N175, N131);
nand NAND3 (N654, N652, N427, N239);
nand NAND2 (N655, N653, N276);
xor XOR2 (N656, N655, N70);
or OR2 (N657, N648, N237);
not NOT1 (N658, N647);
nor NOR4 (N659, N650, N414, N35, N334);
nand NAND4 (N660, N659, N380, N437, N530);
buf BUF1 (N661, N627);
nor NOR3 (N662, N658, N525, N45);
buf BUF1 (N663, N649);
or OR2 (N664, N657, N197);
nor NOR4 (N665, N644, N16, N245, N133);
buf BUF1 (N666, N661);
not NOT1 (N667, N666);
nand NAND3 (N668, N636, N260, N344);
xor XOR2 (N669, N646, N127);
or OR3 (N670, N662, N374, N477);
buf BUF1 (N671, N665);
and AND4 (N672, N670, N33, N79, N273);
or OR2 (N673, N664, N654);
nor NOR4 (N674, N287, N580, N104, N29);
nand NAND4 (N675, N660, N503, N234, N216);
or OR4 (N676, N673, N40, N543, N273);
or OR3 (N677, N675, N398, N338);
not NOT1 (N678, N677);
buf BUF1 (N679, N663);
and AND2 (N680, N678, N228);
or OR3 (N681, N679, N322, N487);
xor XOR2 (N682, N669, N400);
and AND2 (N683, N681, N154);
buf BUF1 (N684, N674);
buf BUF1 (N685, N667);
nor NOR3 (N686, N672, N563, N103);
and AND2 (N687, N682, N370);
nand NAND4 (N688, N684, N534, N151, N230);
and AND4 (N689, N685, N440, N348, N24);
not NOT1 (N690, N676);
not NOT1 (N691, N687);
xor XOR2 (N692, N668, N233);
nor NOR3 (N693, N690, N478, N178);
nor NOR4 (N694, N680, N260, N44, N281);
and AND4 (N695, N694, N533, N462, N576);
nand NAND2 (N696, N671, N107);
and AND2 (N697, N686, N169);
xor XOR2 (N698, N693, N512);
or OR4 (N699, N696, N659, N357, N71);
or OR4 (N700, N683, N40, N598, N413);
or OR3 (N701, N695, N153, N415);
nor NOR3 (N702, N697, N467, N420);
nor NOR4 (N703, N701, N230, N611, N360);
not NOT1 (N704, N702);
and AND4 (N705, N704, N688, N388, N116);
xor XOR2 (N706, N591, N289);
buf BUF1 (N707, N700);
not NOT1 (N708, N706);
buf BUF1 (N709, N703);
buf BUF1 (N710, N707);
xor XOR2 (N711, N699, N342);
buf BUF1 (N712, N709);
or OR4 (N713, N692, N203, N89, N617);
nand NAND4 (N714, N656, N556, N68, N698);
nor NOR3 (N715, N199, N9, N368);
buf BUF1 (N716, N710);
and AND4 (N717, N691, N490, N10, N495);
or OR2 (N718, N705, N82);
nand NAND3 (N719, N712, N475, N87);
xor XOR2 (N720, N711, N81);
not NOT1 (N721, N715);
not NOT1 (N722, N714);
or OR4 (N723, N722, N212, N145, N543);
buf BUF1 (N724, N719);
not NOT1 (N725, N717);
or OR4 (N726, N716, N104, N720, N494);
buf BUF1 (N727, N674);
not NOT1 (N728, N718);
nor NOR3 (N729, N726, N417, N364);
xor XOR2 (N730, N727, N195);
and AND2 (N731, N730, N530);
xor XOR2 (N732, N708, N616);
buf BUF1 (N733, N732);
nand NAND2 (N734, N721, N369);
nand NAND2 (N735, N728, N588);
not NOT1 (N736, N723);
nor NOR4 (N737, N736, N365, N687, N155);
not NOT1 (N738, N734);
and AND2 (N739, N689, N9);
buf BUF1 (N740, N724);
nor NOR3 (N741, N738, N423, N402);
and AND3 (N742, N737, N19, N538);
not NOT1 (N743, N731);
nand NAND4 (N744, N713, N363, N550, N300);
xor XOR2 (N745, N725, N708);
nand NAND2 (N746, N745, N544);
not NOT1 (N747, N735);
or OR2 (N748, N741, N73);
not NOT1 (N749, N739);
nand NAND2 (N750, N748, N301);
not NOT1 (N751, N747);
not NOT1 (N752, N742);
or OR4 (N753, N751, N303, N286, N177);
nor NOR2 (N754, N743, N248);
nor NOR4 (N755, N752, N380, N706, N532);
buf BUF1 (N756, N740);
buf BUF1 (N757, N744);
and AND4 (N758, N749, N266, N230, N321);
buf BUF1 (N759, N756);
nor NOR2 (N760, N729, N431);
not NOT1 (N761, N750);
buf BUF1 (N762, N753);
not NOT1 (N763, N760);
nor NOR4 (N764, N754, N625, N338, N85);
nand NAND4 (N765, N746, N140, N645, N495);
nor NOR2 (N766, N761, N477);
nand NAND3 (N767, N758, N702, N655);
nand NAND4 (N768, N763, N99, N94, N234);
not NOT1 (N769, N762);
buf BUF1 (N770, N768);
xor XOR2 (N771, N766, N727);
xor XOR2 (N772, N759, N682);
nor NOR2 (N773, N757, N500);
buf BUF1 (N774, N755);
buf BUF1 (N775, N771);
not NOT1 (N776, N765);
and AND3 (N777, N773, N679, N186);
xor XOR2 (N778, N776, N350);
or OR2 (N779, N777, N151);
nand NAND2 (N780, N767, N15);
and AND3 (N781, N774, N717, N429);
or OR4 (N782, N772, N665, N578, N606);
nand NAND4 (N783, N775, N498, N775, N289);
not NOT1 (N784, N779);
buf BUF1 (N785, N780);
not NOT1 (N786, N781);
nand NAND2 (N787, N770, N772);
or OR3 (N788, N784, N662, N338);
and AND4 (N789, N733, N569, N692, N675);
nor NOR3 (N790, N787, N447, N290);
buf BUF1 (N791, N783);
buf BUF1 (N792, N788);
nor NOR3 (N793, N792, N216, N449);
not NOT1 (N794, N791);
and AND3 (N795, N790, N391, N364);
and AND2 (N796, N785, N288);
and AND4 (N797, N786, N762, N780, N592);
nor NOR4 (N798, N769, N78, N179, N595);
nand NAND2 (N799, N794, N6);
not NOT1 (N800, N795);
not NOT1 (N801, N764);
nor NOR3 (N802, N796, N686, N251);
and AND3 (N803, N778, N534, N410);
nor NOR2 (N804, N800, N771);
nor NOR2 (N805, N793, N296);
and AND3 (N806, N803, N727, N296);
or OR4 (N807, N804, N386, N794, N67);
and AND4 (N808, N789, N773, N612, N562);
nand NAND2 (N809, N806, N383);
or OR4 (N810, N799, N434, N121, N366);
not NOT1 (N811, N802);
or OR2 (N812, N798, N140);
xor XOR2 (N813, N812, N169);
nand NAND3 (N814, N809, N48, N222);
buf BUF1 (N815, N813);
buf BUF1 (N816, N807);
xor XOR2 (N817, N815, N284);
buf BUF1 (N818, N782);
and AND3 (N819, N818, N627, N605);
and AND3 (N820, N819, N614, N111);
nor NOR2 (N821, N805, N670);
nor NOR2 (N822, N811, N560);
xor XOR2 (N823, N797, N711);
nand NAND3 (N824, N801, N610, N239);
xor XOR2 (N825, N821, N778);
buf BUF1 (N826, N820);
nor NOR2 (N827, N810, N333);
and AND3 (N828, N824, N140, N498);
or OR4 (N829, N823, N28, N392, N689);
not NOT1 (N830, N808);
nand NAND3 (N831, N825, N530, N345);
and AND2 (N832, N822, N208);
or OR4 (N833, N814, N646, N273, N728);
and AND4 (N834, N827, N290, N798, N127);
not NOT1 (N835, N817);
xor XOR2 (N836, N835, N473);
and AND4 (N837, N828, N139, N664, N671);
not NOT1 (N838, N832);
or OR2 (N839, N826, N577);
not NOT1 (N840, N837);
not NOT1 (N841, N840);
nand NAND4 (N842, N838, N206, N584, N480);
nor NOR4 (N843, N833, N791, N776, N644);
not NOT1 (N844, N829);
buf BUF1 (N845, N844);
xor XOR2 (N846, N842, N598);
and AND4 (N847, N816, N100, N191, N220);
nand NAND2 (N848, N847, N538);
and AND3 (N849, N831, N338, N236);
buf BUF1 (N850, N849);
not NOT1 (N851, N830);
not NOT1 (N852, N836);
or OR2 (N853, N841, N799);
nor NOR2 (N854, N848, N806);
and AND4 (N855, N850, N20, N196, N312);
or OR3 (N856, N843, N410, N134);
or OR3 (N857, N845, N527, N527);
xor XOR2 (N858, N854, N494);
and AND4 (N859, N856, N258, N722, N251);
xor XOR2 (N860, N857, N361);
not NOT1 (N861, N855);
xor XOR2 (N862, N846, N777);
nand NAND2 (N863, N852, N845);
nand NAND3 (N864, N858, N515, N736);
buf BUF1 (N865, N864);
buf BUF1 (N866, N862);
nor NOR3 (N867, N860, N301, N210);
or OR3 (N868, N834, N344, N9);
nand NAND3 (N869, N863, N758, N112);
not NOT1 (N870, N866);
xor XOR2 (N871, N869, N493);
and AND2 (N872, N861, N540);
nor NOR3 (N873, N853, N397, N204);
or OR4 (N874, N870, N206, N153, N560);
nor NOR4 (N875, N839, N440, N806, N699);
xor XOR2 (N876, N872, N182);
and AND3 (N877, N867, N601, N612);
xor XOR2 (N878, N876, N286);
xor XOR2 (N879, N859, N209);
not NOT1 (N880, N865);
xor XOR2 (N881, N874, N490);
or OR3 (N882, N877, N538, N66);
and AND3 (N883, N871, N172, N463);
nor NOR3 (N884, N875, N78, N596);
buf BUF1 (N885, N879);
or OR3 (N886, N883, N757, N514);
or OR3 (N887, N880, N99, N586);
xor XOR2 (N888, N881, N459);
nor NOR3 (N889, N851, N412, N67);
and AND3 (N890, N885, N462, N134);
buf BUF1 (N891, N886);
nand NAND2 (N892, N888, N532);
nor NOR4 (N893, N889, N124, N833, N117);
not NOT1 (N894, N873);
and AND4 (N895, N893, N710, N290, N217);
or OR3 (N896, N895, N889, N428);
nand NAND3 (N897, N891, N684, N247);
buf BUF1 (N898, N892);
buf BUF1 (N899, N890);
xor XOR2 (N900, N899, N528);
not NOT1 (N901, N878);
and AND3 (N902, N898, N177, N525);
or OR4 (N903, N900, N273, N685, N442);
xor XOR2 (N904, N901, N434);
not NOT1 (N905, N897);
and AND3 (N906, N884, N290, N830);
and AND3 (N907, N902, N371, N330);
nor NOR3 (N908, N906, N221, N262);
not NOT1 (N909, N882);
buf BUF1 (N910, N905);
nand NAND4 (N911, N903, N422, N207, N21);
or OR3 (N912, N908, N602, N803);
or OR3 (N913, N894, N48, N269);
or OR4 (N914, N912, N867, N844, N39);
not NOT1 (N915, N904);
or OR4 (N916, N887, N589, N798, N611);
or OR2 (N917, N868, N5);
or OR4 (N918, N909, N24, N659, N535);
not NOT1 (N919, N907);
not NOT1 (N920, N911);
not NOT1 (N921, N914);
nand NAND3 (N922, N919, N136, N433);
nand NAND4 (N923, N896, N616, N444, N848);
not NOT1 (N924, N917);
not NOT1 (N925, N921);
nor NOR2 (N926, N920, N766);
nor NOR3 (N927, N925, N277, N53);
nand NAND2 (N928, N923, N333);
and AND2 (N929, N926, N278);
and AND2 (N930, N915, N575);
nor NOR2 (N931, N916, N131);
or OR4 (N932, N928, N603, N259, N76);
buf BUF1 (N933, N924);
not NOT1 (N934, N922);
and AND4 (N935, N934, N602, N368, N147);
buf BUF1 (N936, N933);
nor NOR3 (N937, N930, N440, N251);
not NOT1 (N938, N929);
nand NAND3 (N939, N932, N524, N798);
and AND4 (N940, N939, N220, N801, N448);
and AND3 (N941, N910, N446, N760);
xor XOR2 (N942, N913, N879);
buf BUF1 (N943, N941);
or OR4 (N944, N943, N403, N463, N824);
nor NOR3 (N945, N918, N354, N376);
not NOT1 (N946, N931);
nand NAND4 (N947, N927, N188, N665, N69);
not NOT1 (N948, N938);
nand NAND3 (N949, N944, N83, N637);
nor NOR4 (N950, N940, N319, N353, N789);
nor NOR4 (N951, N946, N111, N241, N549);
buf BUF1 (N952, N945);
or OR4 (N953, N948, N793, N724, N404);
nor NOR2 (N954, N953, N197);
not NOT1 (N955, N952);
xor XOR2 (N956, N936, N414);
nand NAND2 (N957, N942, N493);
xor XOR2 (N958, N950, N591);
and AND2 (N959, N956, N861);
buf BUF1 (N960, N955);
nor NOR4 (N961, N959, N712, N44, N902);
not NOT1 (N962, N949);
xor XOR2 (N963, N937, N570);
and AND3 (N964, N963, N142, N638);
xor XOR2 (N965, N951, N103);
not NOT1 (N966, N957);
xor XOR2 (N967, N958, N27);
nor NOR4 (N968, N962, N95, N670, N432);
nor NOR2 (N969, N964, N12);
nand NAND2 (N970, N965, N287);
xor XOR2 (N971, N969, N911);
buf BUF1 (N972, N947);
nand NAND4 (N973, N972, N89, N581, N464);
and AND2 (N974, N971, N763);
xor XOR2 (N975, N960, N532);
xor XOR2 (N976, N954, N370);
buf BUF1 (N977, N967);
and AND4 (N978, N976, N433, N939, N220);
not NOT1 (N979, N975);
buf BUF1 (N980, N968);
xor XOR2 (N981, N978, N466);
nor NOR4 (N982, N966, N798, N602, N791);
nor NOR2 (N983, N979, N708);
nor NOR2 (N984, N970, N22);
buf BUF1 (N985, N980);
not NOT1 (N986, N973);
nand NAND3 (N987, N974, N827, N108);
nand NAND2 (N988, N982, N394);
buf BUF1 (N989, N977);
nor NOR2 (N990, N981, N148);
nand NAND2 (N991, N987, N173);
buf BUF1 (N992, N988);
buf BUF1 (N993, N990);
nand NAND4 (N994, N983, N906, N139, N96);
and AND3 (N995, N992, N410, N828);
nand NAND2 (N996, N993, N778);
xor XOR2 (N997, N989, N835);
buf BUF1 (N998, N985);
nand NAND2 (N999, N986, N599);
buf BUF1 (N1000, N997);
nor NOR2 (N1001, N1000, N816);
and AND4 (N1002, N998, N281, N390, N863);
or OR2 (N1003, N961, N76);
xor XOR2 (N1004, N1002, N748);
or OR2 (N1005, N1004, N493);
or OR4 (N1006, N995, N386, N943, N161);
and AND4 (N1007, N935, N952, N757, N114);
xor XOR2 (N1008, N994, N735);
nor NOR2 (N1009, N1008, N740);
not NOT1 (N1010, N996);
and AND2 (N1011, N1010, N371);
or OR3 (N1012, N1001, N522, N242);
and AND4 (N1013, N1006, N557, N672, N553);
and AND3 (N1014, N1012, N95, N258);
not NOT1 (N1015, N984);
buf BUF1 (N1016, N1007);
nand NAND2 (N1017, N1005, N346);
nand NAND4 (N1018, N1013, N581, N505, N689);
or OR4 (N1019, N1014, N37, N922, N654);
nor NOR4 (N1020, N1003, N794, N976, N68);
nor NOR4 (N1021, N1011, N921, N267, N591);
buf BUF1 (N1022, N1020);
nor NOR2 (N1023, N1015, N207);
nor NOR3 (N1024, N1019, N402, N472);
or OR2 (N1025, N1022, N121);
or OR4 (N1026, N1025, N366, N298, N15);
not NOT1 (N1027, N1021);
not NOT1 (N1028, N1024);
or OR2 (N1029, N1009, N802);
nand NAND3 (N1030, N1026, N169, N502);
or OR2 (N1031, N1028, N713);
and AND2 (N1032, N991, N1014);
nand NAND4 (N1033, N1029, N20, N869, N511);
nand NAND3 (N1034, N1032, N42, N838);
and AND4 (N1035, N1031, N555, N866, N954);
nor NOR3 (N1036, N1030, N476, N953);
nand NAND4 (N1037, N1017, N991, N1024, N904);
xor XOR2 (N1038, N1035, N242);
not NOT1 (N1039, N1018);
nand NAND2 (N1040, N1033, N876);
not NOT1 (N1041, N1036);
or OR2 (N1042, N1023, N153);
not NOT1 (N1043, N1027);
xor XOR2 (N1044, N1016, N100);
not NOT1 (N1045, N1041);
and AND4 (N1046, N1045, N497, N64, N749);
xor XOR2 (N1047, N1040, N504);
or OR3 (N1048, N999, N454, N863);
nand NAND3 (N1049, N1037, N297, N288);
nand NAND3 (N1050, N1038, N212, N782);
nor NOR3 (N1051, N1043, N164, N396);
not NOT1 (N1052, N1051);
nand NAND4 (N1053, N1048, N127, N909, N874);
nand NAND2 (N1054, N1046, N764);
and AND4 (N1055, N1050, N899, N573, N417);
nand NAND2 (N1056, N1034, N752);
buf BUF1 (N1057, N1054);
and AND2 (N1058, N1053, N145);
xor XOR2 (N1059, N1058, N832);
xor XOR2 (N1060, N1044, N294);
nand NAND4 (N1061, N1039, N201, N577, N402);
and AND4 (N1062, N1047, N570, N646, N322);
nor NOR2 (N1063, N1052, N832);
or OR3 (N1064, N1063, N381, N692);
not NOT1 (N1065, N1060);
not NOT1 (N1066, N1056);
and AND4 (N1067, N1062, N982, N532, N920);
nor NOR3 (N1068, N1057, N614, N1017);
xor XOR2 (N1069, N1059, N558);
nand NAND4 (N1070, N1065, N319, N711, N107);
nor NOR3 (N1071, N1066, N616, N114);
xor XOR2 (N1072, N1068, N664);
nand NAND4 (N1073, N1067, N150, N443, N627);
buf BUF1 (N1074, N1070);
not NOT1 (N1075, N1073);
and AND2 (N1076, N1072, N3);
not NOT1 (N1077, N1069);
and AND4 (N1078, N1074, N266, N907, N177);
not NOT1 (N1079, N1075);
or OR4 (N1080, N1077, N3, N277, N798);
not NOT1 (N1081, N1061);
or OR2 (N1082, N1080, N493);
not NOT1 (N1083, N1079);
and AND2 (N1084, N1071, N19);
buf BUF1 (N1085, N1083);
xor XOR2 (N1086, N1076, N30);
nand NAND4 (N1087, N1085, N625, N207, N601);
or OR4 (N1088, N1082, N425, N735, N226);
or OR2 (N1089, N1086, N175);
not NOT1 (N1090, N1088);
buf BUF1 (N1091, N1049);
buf BUF1 (N1092, N1091);
nand NAND3 (N1093, N1092, N804, N935);
nand NAND3 (N1094, N1042, N213, N74);
nand NAND3 (N1095, N1093, N82, N248);
and AND2 (N1096, N1087, N948);
buf BUF1 (N1097, N1095);
nand NAND4 (N1098, N1081, N233, N425, N214);
not NOT1 (N1099, N1089);
buf BUF1 (N1100, N1055);
and AND3 (N1101, N1096, N582, N1004);
not NOT1 (N1102, N1100);
nand NAND3 (N1103, N1098, N337, N344);
and AND2 (N1104, N1101, N985);
or OR3 (N1105, N1090, N499, N460);
and AND3 (N1106, N1097, N918, N589);
nand NAND3 (N1107, N1064, N778, N688);
xor XOR2 (N1108, N1104, N892);
nand NAND4 (N1109, N1103, N542, N361, N321);
xor XOR2 (N1110, N1109, N219);
or OR3 (N1111, N1099, N536, N4);
nor NOR3 (N1112, N1105, N531, N1018);
nor NOR3 (N1113, N1094, N291, N836);
not NOT1 (N1114, N1113);
nand NAND4 (N1115, N1084, N527, N180, N773);
buf BUF1 (N1116, N1115);
not NOT1 (N1117, N1078);
and AND2 (N1118, N1107, N874);
xor XOR2 (N1119, N1116, N1074);
not NOT1 (N1120, N1118);
buf BUF1 (N1121, N1117);
xor XOR2 (N1122, N1119, N1028);
nand NAND3 (N1123, N1110, N764, N451);
and AND3 (N1124, N1120, N406, N105);
not NOT1 (N1125, N1102);
and AND2 (N1126, N1112, N895);
and AND4 (N1127, N1108, N246, N282, N1032);
and AND4 (N1128, N1106, N706, N512, N994);
xor XOR2 (N1129, N1111, N298);
or OR2 (N1130, N1126, N636);
not NOT1 (N1131, N1123);
xor XOR2 (N1132, N1124, N119);
nor NOR3 (N1133, N1122, N152, N683);
nand NAND3 (N1134, N1131, N991, N536);
and AND4 (N1135, N1132, N741, N1115, N1057);
nor NOR3 (N1136, N1129, N219, N181);
and AND4 (N1137, N1136, N784, N174, N1040);
or OR3 (N1138, N1121, N898, N591);
xor XOR2 (N1139, N1130, N236);
and AND4 (N1140, N1135, N90, N299, N264);
or OR4 (N1141, N1139, N639, N162, N527);
xor XOR2 (N1142, N1140, N727);
not NOT1 (N1143, N1138);
xor XOR2 (N1144, N1125, N693);
nand NAND3 (N1145, N1127, N389, N237);
nand NAND4 (N1146, N1143, N488, N902, N505);
nand NAND2 (N1147, N1142, N601);
buf BUF1 (N1148, N1147);
or OR4 (N1149, N1134, N135, N614, N273);
nor NOR2 (N1150, N1133, N281);
nor NOR3 (N1151, N1145, N687, N721);
and AND2 (N1152, N1150, N135);
not NOT1 (N1153, N1144);
nor NOR4 (N1154, N1146, N662, N532, N840);
or OR2 (N1155, N1137, N896);
nor NOR2 (N1156, N1148, N187);
nand NAND3 (N1157, N1155, N763, N364);
or OR4 (N1158, N1153, N32, N921, N339);
nor NOR2 (N1159, N1152, N858);
xor XOR2 (N1160, N1128, N599);
nor NOR3 (N1161, N1160, N488, N1009);
and AND3 (N1162, N1151, N802, N871);
not NOT1 (N1163, N1114);
xor XOR2 (N1164, N1156, N621);
not NOT1 (N1165, N1141);
and AND2 (N1166, N1159, N228);
nor NOR4 (N1167, N1164, N671, N364, N519);
and AND3 (N1168, N1167, N448, N356);
nand NAND2 (N1169, N1157, N1051);
and AND4 (N1170, N1165, N411, N988, N1088);
nand NAND2 (N1171, N1163, N991);
not NOT1 (N1172, N1154);
buf BUF1 (N1173, N1161);
nand NAND4 (N1174, N1149, N585, N730, N400);
nor NOR4 (N1175, N1166, N962, N758, N621);
nor NOR3 (N1176, N1171, N340, N941);
and AND3 (N1177, N1174, N244, N1090);
or OR4 (N1178, N1176, N908, N426, N240);
and AND2 (N1179, N1175, N53);
xor XOR2 (N1180, N1168, N678);
nand NAND4 (N1181, N1169, N230, N496, N1141);
and AND2 (N1182, N1158, N418);
not NOT1 (N1183, N1162);
buf BUF1 (N1184, N1170);
nand NAND2 (N1185, N1173, N921);
nand NAND4 (N1186, N1185, N161, N548, N218);
xor XOR2 (N1187, N1177, N257);
or OR3 (N1188, N1178, N212, N527);
nand NAND4 (N1189, N1172, N932, N492, N512);
or OR3 (N1190, N1189, N996, N851);
or OR4 (N1191, N1181, N1074, N5, N274);
or OR2 (N1192, N1188, N465);
nand NAND3 (N1193, N1190, N1187, N361);
buf BUF1 (N1194, N890);
and AND2 (N1195, N1191, N11);
buf BUF1 (N1196, N1192);
nand NAND3 (N1197, N1196, N347, N123);
not NOT1 (N1198, N1194);
buf BUF1 (N1199, N1193);
and AND4 (N1200, N1195, N244, N359, N542);
nor NOR2 (N1201, N1180, N711);
and AND3 (N1202, N1182, N811, N1142);
xor XOR2 (N1203, N1200, N282);
nor NOR3 (N1204, N1183, N1153, N386);
and AND3 (N1205, N1203, N172, N461);
buf BUF1 (N1206, N1201);
or OR4 (N1207, N1186, N696, N1027, N483);
and AND2 (N1208, N1184, N822);
and AND2 (N1209, N1202, N777);
nor NOR4 (N1210, N1207, N125, N646, N1048);
or OR3 (N1211, N1197, N789, N144);
not NOT1 (N1212, N1208);
xor XOR2 (N1213, N1209, N580);
or OR4 (N1214, N1213, N993, N482, N922);
xor XOR2 (N1215, N1212, N878);
not NOT1 (N1216, N1205);
nand NAND4 (N1217, N1214, N552, N405, N1018);
buf BUF1 (N1218, N1211);
xor XOR2 (N1219, N1217, N441);
and AND3 (N1220, N1206, N1090, N11);
and AND4 (N1221, N1198, N82, N180, N1062);
or OR3 (N1222, N1216, N153, N623);
nand NAND2 (N1223, N1219, N809);
and AND4 (N1224, N1215, N991, N1035, N272);
nor NOR3 (N1225, N1179, N1149, N67);
not NOT1 (N1226, N1224);
or OR3 (N1227, N1222, N109, N593);
buf BUF1 (N1228, N1223);
nand NAND2 (N1229, N1221, N121);
nor NOR4 (N1230, N1226, N98, N772, N328);
or OR2 (N1231, N1204, N396);
not NOT1 (N1232, N1220);
nor NOR4 (N1233, N1229, N474, N662, N1056);
buf BUF1 (N1234, N1225);
buf BUF1 (N1235, N1228);
not NOT1 (N1236, N1199);
and AND2 (N1237, N1227, N1063);
xor XOR2 (N1238, N1230, N288);
or OR3 (N1239, N1237, N1117, N951);
nor NOR2 (N1240, N1238, N623);
nor NOR3 (N1241, N1235, N783, N624);
and AND3 (N1242, N1232, N346, N363);
xor XOR2 (N1243, N1236, N68);
nand NAND2 (N1244, N1218, N541);
buf BUF1 (N1245, N1239);
not NOT1 (N1246, N1233);
or OR3 (N1247, N1243, N14, N209);
nand NAND3 (N1248, N1246, N694, N1139);
not NOT1 (N1249, N1247);
not NOT1 (N1250, N1231);
not NOT1 (N1251, N1234);
nor NOR3 (N1252, N1251, N421, N87);
and AND3 (N1253, N1248, N635, N286);
and AND3 (N1254, N1242, N755, N703);
xor XOR2 (N1255, N1210, N152);
and AND4 (N1256, N1240, N87, N676, N311);
or OR4 (N1257, N1254, N1081, N569, N111);
xor XOR2 (N1258, N1241, N1043);
xor XOR2 (N1259, N1256, N110);
nand NAND2 (N1260, N1244, N1127);
or OR2 (N1261, N1245, N526);
or OR2 (N1262, N1252, N1222);
buf BUF1 (N1263, N1253);
buf BUF1 (N1264, N1261);
buf BUF1 (N1265, N1255);
and AND3 (N1266, N1259, N290, N840);
nand NAND2 (N1267, N1258, N564);
buf BUF1 (N1268, N1250);
not NOT1 (N1269, N1267);
nand NAND4 (N1270, N1265, N619, N650, N1202);
not NOT1 (N1271, N1270);
and AND3 (N1272, N1260, N662, N593);
xor XOR2 (N1273, N1268, N1265);
not NOT1 (N1274, N1264);
nor NOR4 (N1275, N1271, N227, N77, N640);
nand NAND3 (N1276, N1263, N696, N501);
and AND3 (N1277, N1274, N165, N1267);
nor NOR2 (N1278, N1257, N1237);
nor NOR4 (N1279, N1273, N932, N722, N1136);
xor XOR2 (N1280, N1279, N480);
and AND2 (N1281, N1266, N576);
nor NOR4 (N1282, N1262, N330, N712, N200);
and AND2 (N1283, N1249, N120);
not NOT1 (N1284, N1272);
nand NAND3 (N1285, N1276, N454, N342);
buf BUF1 (N1286, N1277);
buf BUF1 (N1287, N1280);
nor NOR4 (N1288, N1283, N593, N1149, N504);
not NOT1 (N1289, N1288);
not NOT1 (N1290, N1289);
or OR2 (N1291, N1285, N1032);
nand NAND4 (N1292, N1291, N83, N956, N489);
nor NOR4 (N1293, N1290, N456, N1283, N802);
or OR4 (N1294, N1293, N563, N27, N455);
and AND3 (N1295, N1282, N1274, N170);
not NOT1 (N1296, N1294);
xor XOR2 (N1297, N1281, N453);
buf BUF1 (N1298, N1292);
buf BUF1 (N1299, N1284);
not NOT1 (N1300, N1286);
or OR4 (N1301, N1287, N194, N802, N973);
buf BUF1 (N1302, N1278);
and AND2 (N1303, N1296, N155);
nor NOR3 (N1304, N1269, N726, N1291);
not NOT1 (N1305, N1300);
buf BUF1 (N1306, N1298);
or OR4 (N1307, N1306, N450, N1151, N1126);
nand NAND3 (N1308, N1297, N220, N770);
nand NAND3 (N1309, N1308, N658, N238);
xor XOR2 (N1310, N1295, N1191);
nand NAND4 (N1311, N1301, N157, N499, N785);
xor XOR2 (N1312, N1305, N160);
and AND4 (N1313, N1302, N341, N827, N135);
and AND3 (N1314, N1312, N1024, N113);
not NOT1 (N1315, N1313);
not NOT1 (N1316, N1275);
or OR3 (N1317, N1316, N922, N749);
not NOT1 (N1318, N1311);
xor XOR2 (N1319, N1315, N1016);
and AND3 (N1320, N1307, N722, N1217);
not NOT1 (N1321, N1319);
xor XOR2 (N1322, N1310, N879);
or OR4 (N1323, N1322, N369, N1258, N335);
or OR2 (N1324, N1318, N42);
buf BUF1 (N1325, N1324);
nand NAND4 (N1326, N1314, N403, N897, N1140);
buf BUF1 (N1327, N1326);
buf BUF1 (N1328, N1320);
not NOT1 (N1329, N1309);
nor NOR2 (N1330, N1317, N79);
and AND3 (N1331, N1330, N573, N502);
not NOT1 (N1332, N1304);
nand NAND4 (N1333, N1299, N1319, N1303, N1136);
and AND2 (N1334, N429, N947);
nand NAND2 (N1335, N1333, N567);
nand NAND2 (N1336, N1328, N80);
nor NOR2 (N1337, N1331, N831);
not NOT1 (N1338, N1323);
nor NOR2 (N1339, N1321, N1166);
and AND4 (N1340, N1336, N664, N189, N760);
nor NOR4 (N1341, N1327, N331, N1282, N379);
nand NAND2 (N1342, N1337, N1187);
or OR2 (N1343, N1340, N603);
or OR2 (N1344, N1334, N363);
and AND3 (N1345, N1325, N300, N655);
buf BUF1 (N1346, N1343);
or OR4 (N1347, N1342, N665, N822, N118);
xor XOR2 (N1348, N1329, N647);
and AND3 (N1349, N1341, N461, N460);
or OR2 (N1350, N1345, N789);
and AND2 (N1351, N1344, N248);
buf BUF1 (N1352, N1351);
xor XOR2 (N1353, N1350, N1271);
not NOT1 (N1354, N1346);
and AND2 (N1355, N1338, N651);
nor NOR2 (N1356, N1339, N621);
or OR3 (N1357, N1356, N48, N710);
and AND2 (N1358, N1332, N483);
buf BUF1 (N1359, N1352);
and AND4 (N1360, N1357, N512, N1257, N1254);
buf BUF1 (N1361, N1358);
and AND4 (N1362, N1348, N634, N1348, N524);
not NOT1 (N1363, N1347);
xor XOR2 (N1364, N1361, N712);
and AND4 (N1365, N1335, N324, N1309, N216);
and AND2 (N1366, N1360, N862);
nand NAND4 (N1367, N1354, N4, N483, N886);
nor NOR4 (N1368, N1359, N250, N677, N288);
xor XOR2 (N1369, N1368, N667);
xor XOR2 (N1370, N1362, N1020);
buf BUF1 (N1371, N1365);
and AND2 (N1372, N1367, N632);
xor XOR2 (N1373, N1363, N25);
or OR2 (N1374, N1353, N214);
nor NOR4 (N1375, N1364, N703, N192, N437);
or OR4 (N1376, N1371, N1238, N631, N994);
nor NOR2 (N1377, N1374, N678);
not NOT1 (N1378, N1355);
xor XOR2 (N1379, N1378, N79);
xor XOR2 (N1380, N1376, N131);
and AND2 (N1381, N1372, N801);
nand NAND3 (N1382, N1349, N722, N760);
or OR4 (N1383, N1382, N875, N244, N1303);
or OR4 (N1384, N1375, N824, N1347, N906);
and AND4 (N1385, N1384, N139, N321, N1080);
or OR4 (N1386, N1379, N673, N16, N235);
nor NOR3 (N1387, N1366, N862, N1012);
nor NOR4 (N1388, N1373, N978, N381, N933);
not NOT1 (N1389, N1380);
and AND2 (N1390, N1381, N425);
and AND4 (N1391, N1388, N898, N762, N1237);
and AND4 (N1392, N1387, N510, N505, N1388);
not NOT1 (N1393, N1390);
nand NAND3 (N1394, N1393, N824, N840);
xor XOR2 (N1395, N1383, N1372);
nand NAND4 (N1396, N1391, N1253, N50, N542);
nand NAND3 (N1397, N1389, N1373, N1055);
nor NOR4 (N1398, N1385, N58, N119, N437);
nor NOR2 (N1399, N1369, N1366);
nand NAND4 (N1400, N1395, N483, N462, N471);
buf BUF1 (N1401, N1394);
xor XOR2 (N1402, N1396, N286);
xor XOR2 (N1403, N1402, N615);
and AND2 (N1404, N1401, N257);
not NOT1 (N1405, N1386);
nor NOR3 (N1406, N1370, N1005, N527);
and AND4 (N1407, N1406, N1331, N710, N971);
buf BUF1 (N1408, N1397);
buf BUF1 (N1409, N1377);
not NOT1 (N1410, N1392);
or OR2 (N1411, N1404, N1014);
nor NOR2 (N1412, N1410, N441);
nor NOR2 (N1413, N1405, N1410);
buf BUF1 (N1414, N1411);
or OR4 (N1415, N1403, N1134, N1202, N139);
nor NOR2 (N1416, N1398, N430);
not NOT1 (N1417, N1413);
not NOT1 (N1418, N1412);
buf BUF1 (N1419, N1408);
xor XOR2 (N1420, N1415, N1363);
xor XOR2 (N1421, N1407, N1215);
not NOT1 (N1422, N1409);
or OR2 (N1423, N1422, N487);
not NOT1 (N1424, N1419);
buf BUF1 (N1425, N1416);
or OR3 (N1426, N1424, N1399, N594);
or OR3 (N1427, N1351, N1238, N332);
and AND2 (N1428, N1421, N1123);
nor NOR4 (N1429, N1426, N621, N893, N510);
nor NOR3 (N1430, N1427, N1241, N25);
nor NOR3 (N1431, N1429, N194, N658);
buf BUF1 (N1432, N1423);
nand NAND4 (N1433, N1430, N634, N1246, N536);
nor NOR2 (N1434, N1425, N1179);
xor XOR2 (N1435, N1434, N21);
and AND2 (N1436, N1414, N866);
nor NOR4 (N1437, N1417, N468, N1199, N98);
not NOT1 (N1438, N1433);
nor NOR3 (N1439, N1431, N939, N160);
not NOT1 (N1440, N1435);
xor XOR2 (N1441, N1439, N558);
buf BUF1 (N1442, N1440);
nand NAND2 (N1443, N1437, N1306);
buf BUF1 (N1444, N1436);
xor XOR2 (N1445, N1438, N260);
nor NOR3 (N1446, N1420, N198, N1071);
nor NOR2 (N1447, N1432, N752);
or OR4 (N1448, N1447, N836, N286, N1349);
nor NOR4 (N1449, N1446, N424, N1207, N1252);
and AND3 (N1450, N1445, N766, N397);
not NOT1 (N1451, N1441);
buf BUF1 (N1452, N1428);
nand NAND4 (N1453, N1448, N1060, N1190, N382);
not NOT1 (N1454, N1453);
nor NOR3 (N1455, N1444, N591, N230);
nand NAND3 (N1456, N1443, N1151, N622);
buf BUF1 (N1457, N1456);
nor NOR4 (N1458, N1449, N805, N411, N778);
and AND4 (N1459, N1457, N344, N376, N574);
not NOT1 (N1460, N1450);
buf BUF1 (N1461, N1454);
nor NOR3 (N1462, N1460, N742, N1078);
buf BUF1 (N1463, N1459);
and AND2 (N1464, N1451, N475);
and AND3 (N1465, N1452, N1362, N252);
not NOT1 (N1466, N1461);
nand NAND2 (N1467, N1458, N2);
and AND3 (N1468, N1455, N1160, N778);
not NOT1 (N1469, N1464);
or OR4 (N1470, N1468, N617, N229, N175);
not NOT1 (N1471, N1418);
nor NOR4 (N1472, N1463, N640, N1412, N639);
buf BUF1 (N1473, N1400);
or OR2 (N1474, N1467, N264);
nor NOR2 (N1475, N1466, N1118);
and AND3 (N1476, N1474, N129, N25);
buf BUF1 (N1477, N1470);
or OR4 (N1478, N1476, N992, N309, N1171);
nor NOR4 (N1479, N1478, N1446, N783, N334);
not NOT1 (N1480, N1475);
buf BUF1 (N1481, N1465);
not NOT1 (N1482, N1442);
nand NAND3 (N1483, N1481, N640, N487);
not NOT1 (N1484, N1472);
nand NAND4 (N1485, N1473, N531, N1369, N1387);
nor NOR3 (N1486, N1477, N467, N945);
nand NAND3 (N1487, N1462, N688, N1030);
nor NOR2 (N1488, N1483, N943);
xor XOR2 (N1489, N1487, N1135);
nor NOR2 (N1490, N1471, N451);
buf BUF1 (N1491, N1488);
xor XOR2 (N1492, N1479, N1239);
buf BUF1 (N1493, N1480);
buf BUF1 (N1494, N1486);
nor NOR3 (N1495, N1484, N22, N725);
not NOT1 (N1496, N1469);
nand NAND4 (N1497, N1495, N1342, N839, N162);
nor NOR3 (N1498, N1491, N193, N1343);
nand NAND3 (N1499, N1498, N974, N1197);
or OR3 (N1500, N1482, N1112, N443);
not NOT1 (N1501, N1499);
nor NOR4 (N1502, N1496, N133, N352, N539);
not NOT1 (N1503, N1500);
nand NAND3 (N1504, N1501, N542, N395);
buf BUF1 (N1505, N1497);
nand NAND2 (N1506, N1502, N703);
buf BUF1 (N1507, N1505);
buf BUF1 (N1508, N1494);
not NOT1 (N1509, N1489);
nand NAND2 (N1510, N1492, N1341);
nand NAND2 (N1511, N1485, N583);
nor NOR2 (N1512, N1506, N953);
nor NOR3 (N1513, N1493, N399, N165);
nor NOR3 (N1514, N1508, N1445, N1020);
nor NOR4 (N1515, N1504, N856, N416, N825);
nand NAND2 (N1516, N1514, N126);
xor XOR2 (N1517, N1507, N1383);
xor XOR2 (N1518, N1515, N1489);
nand NAND4 (N1519, N1510, N419, N1054, N373);
and AND2 (N1520, N1511, N168);
or OR2 (N1521, N1503, N980);
nor NOR3 (N1522, N1520, N1265, N486);
not NOT1 (N1523, N1490);
xor XOR2 (N1524, N1516, N882);
xor XOR2 (N1525, N1517, N792);
xor XOR2 (N1526, N1518, N857);
xor XOR2 (N1527, N1521, N1270);
nand NAND4 (N1528, N1523, N1380, N220, N471);
and AND4 (N1529, N1527, N818, N61, N728);
buf BUF1 (N1530, N1513);
buf BUF1 (N1531, N1526);
nand NAND4 (N1532, N1530, N567, N818, N1026);
buf BUF1 (N1533, N1509);
not NOT1 (N1534, N1529);
nand NAND2 (N1535, N1532, N80);
nor NOR3 (N1536, N1535, N553, N668);
and AND4 (N1537, N1524, N182, N1258, N1067);
not NOT1 (N1538, N1537);
nand NAND2 (N1539, N1512, N166);
xor XOR2 (N1540, N1519, N853);
not NOT1 (N1541, N1531);
nand NAND2 (N1542, N1534, N1439);
not NOT1 (N1543, N1536);
buf BUF1 (N1544, N1542);
xor XOR2 (N1545, N1533, N1159);
or OR2 (N1546, N1528, N60);
nor NOR4 (N1547, N1543, N181, N242, N1178);
nand NAND2 (N1548, N1540, N238);
buf BUF1 (N1549, N1538);
buf BUF1 (N1550, N1541);
nor NOR4 (N1551, N1548, N394, N1426, N950);
not NOT1 (N1552, N1545);
or OR2 (N1553, N1549, N640);
nor NOR4 (N1554, N1553, N77, N466, N58);
xor XOR2 (N1555, N1522, N1052);
or OR3 (N1556, N1554, N79, N261);
and AND2 (N1557, N1547, N871);
nand NAND4 (N1558, N1557, N1077, N426, N756);
or OR4 (N1559, N1552, N1403, N204, N404);
not NOT1 (N1560, N1525);
buf BUF1 (N1561, N1546);
and AND2 (N1562, N1559, N590);
xor XOR2 (N1563, N1561, N267);
xor XOR2 (N1564, N1558, N105);
nand NAND4 (N1565, N1551, N1525, N444, N258);
nor NOR2 (N1566, N1564, N886);
xor XOR2 (N1567, N1565, N664);
or OR3 (N1568, N1544, N699, N367);
not NOT1 (N1569, N1568);
or OR4 (N1570, N1550, N735, N791, N1042);
xor XOR2 (N1571, N1570, N94);
xor XOR2 (N1572, N1556, N1446);
nand NAND2 (N1573, N1572, N377);
xor XOR2 (N1574, N1555, N867);
or OR2 (N1575, N1567, N949);
buf BUF1 (N1576, N1569);
buf BUF1 (N1577, N1539);
buf BUF1 (N1578, N1575);
xor XOR2 (N1579, N1578, N1518);
nand NAND3 (N1580, N1571, N248, N42);
not NOT1 (N1581, N1576);
nor NOR3 (N1582, N1562, N293, N748);
xor XOR2 (N1583, N1573, N29);
or OR2 (N1584, N1560, N482);
nand NAND2 (N1585, N1577, N1052);
nand NAND3 (N1586, N1582, N1198, N435);
nand NAND3 (N1587, N1585, N1183, N944);
or OR3 (N1588, N1587, N725, N483);
buf BUF1 (N1589, N1574);
not NOT1 (N1590, N1580);
nand NAND3 (N1591, N1586, N198, N53);
nand NAND3 (N1592, N1566, N1043, N406);
xor XOR2 (N1593, N1592, N608);
xor XOR2 (N1594, N1583, N1473);
nand NAND2 (N1595, N1581, N609);
nor NOR3 (N1596, N1595, N57, N93);
nand NAND4 (N1597, N1591, N1069, N439, N340);
nand NAND4 (N1598, N1563, N1575, N538, N188);
or OR4 (N1599, N1588, N799, N274, N675);
or OR4 (N1600, N1594, N658, N1244, N1128);
and AND3 (N1601, N1598, N159, N665);
nand NAND2 (N1602, N1579, N538);
xor XOR2 (N1603, N1599, N167);
nor NOR3 (N1604, N1584, N242, N1527);
or OR3 (N1605, N1600, N695, N1507);
xor XOR2 (N1606, N1597, N101);
buf BUF1 (N1607, N1590);
nor NOR2 (N1608, N1604, N268);
xor XOR2 (N1609, N1606, N66);
buf BUF1 (N1610, N1607);
nand NAND2 (N1611, N1589, N168);
nor NOR4 (N1612, N1602, N1280, N240, N1366);
not NOT1 (N1613, N1608);
xor XOR2 (N1614, N1596, N552);
buf BUF1 (N1615, N1593);
and AND3 (N1616, N1612, N1433, N875);
not NOT1 (N1617, N1611);
xor XOR2 (N1618, N1605, N1520);
buf BUF1 (N1619, N1616);
xor XOR2 (N1620, N1603, N409);
nor NOR3 (N1621, N1620, N419, N311);
and AND2 (N1622, N1613, N1463);
or OR3 (N1623, N1617, N568, N654);
or OR3 (N1624, N1619, N799, N1428);
not NOT1 (N1625, N1614);
xor XOR2 (N1626, N1621, N787);
and AND4 (N1627, N1601, N192, N133, N93);
nor NOR3 (N1628, N1627, N875, N241);
and AND3 (N1629, N1628, N860, N77);
or OR4 (N1630, N1624, N852, N317, N1581);
nor NOR2 (N1631, N1618, N562);
and AND4 (N1632, N1622, N870, N593, N1356);
xor XOR2 (N1633, N1630, N717);
not NOT1 (N1634, N1633);
not NOT1 (N1635, N1629);
buf BUF1 (N1636, N1610);
and AND3 (N1637, N1625, N411, N694);
and AND3 (N1638, N1637, N1606, N1060);
not NOT1 (N1639, N1631);
nor NOR2 (N1640, N1634, N755);
not NOT1 (N1641, N1623);
buf BUF1 (N1642, N1626);
or OR2 (N1643, N1638, N218);
buf BUF1 (N1644, N1636);
buf BUF1 (N1645, N1640);
and AND3 (N1646, N1641, N872, N642);
and AND2 (N1647, N1645, N447);
not NOT1 (N1648, N1632);
and AND4 (N1649, N1639, N1611, N1431, N18);
nand NAND3 (N1650, N1615, N1199, N1179);
nand NAND2 (N1651, N1642, N598);
buf BUF1 (N1652, N1649);
not NOT1 (N1653, N1647);
nand NAND4 (N1654, N1609, N1454, N1181, N894);
xor XOR2 (N1655, N1652, N29);
and AND2 (N1656, N1648, N330);
nand NAND3 (N1657, N1643, N480, N1127);
and AND3 (N1658, N1651, N1641, N293);
and AND3 (N1659, N1657, N404, N1537);
not NOT1 (N1660, N1635);
buf BUF1 (N1661, N1650);
xor XOR2 (N1662, N1653, N405);
xor XOR2 (N1663, N1644, N165);
and AND4 (N1664, N1659, N1659, N88, N1323);
buf BUF1 (N1665, N1655);
and AND2 (N1666, N1654, N1110);
buf BUF1 (N1667, N1656);
nor NOR4 (N1668, N1666, N420, N503, N1178);
buf BUF1 (N1669, N1667);
buf BUF1 (N1670, N1669);
and AND3 (N1671, N1665, N1426, N415);
nand NAND2 (N1672, N1664, N1561);
nor NOR3 (N1673, N1658, N10, N57);
buf BUF1 (N1674, N1673);
xor XOR2 (N1675, N1661, N855);
and AND4 (N1676, N1668, N1032, N69, N351);
or OR3 (N1677, N1670, N260, N1139);
nand NAND2 (N1678, N1662, N704);
nand NAND4 (N1679, N1646, N1368, N1518, N40);
nor NOR2 (N1680, N1677, N933);
nand NAND4 (N1681, N1660, N1267, N1467, N381);
and AND4 (N1682, N1663, N726, N1074, N466);
or OR4 (N1683, N1674, N817, N89, N887);
or OR2 (N1684, N1678, N172);
buf BUF1 (N1685, N1683);
not NOT1 (N1686, N1680);
nor NOR4 (N1687, N1682, N753, N865, N490);
nand NAND3 (N1688, N1681, N1227, N815);
nand NAND2 (N1689, N1687, N1222);
buf BUF1 (N1690, N1675);
not NOT1 (N1691, N1688);
not NOT1 (N1692, N1671);
buf BUF1 (N1693, N1692);
nor NOR4 (N1694, N1690, N144, N64, N704);
nand NAND4 (N1695, N1685, N1081, N239, N1576);
not NOT1 (N1696, N1689);
nand NAND4 (N1697, N1684, N75, N1040, N510);
xor XOR2 (N1698, N1686, N1445);
or OR2 (N1699, N1691, N1338);
and AND2 (N1700, N1696, N1055);
buf BUF1 (N1701, N1672);
and AND4 (N1702, N1693, N364, N1499, N1642);
xor XOR2 (N1703, N1679, N1216);
nand NAND2 (N1704, N1703, N894);
xor XOR2 (N1705, N1697, N1185);
nand NAND4 (N1706, N1701, N125, N991, N1064);
not NOT1 (N1707, N1699);
or OR3 (N1708, N1705, N894, N1151);
nor NOR2 (N1709, N1704, N1262);
not NOT1 (N1710, N1707);
and AND3 (N1711, N1698, N1157, N1154);
and AND2 (N1712, N1706, N1664);
nand NAND3 (N1713, N1695, N1139, N138);
or OR2 (N1714, N1676, N596);
nor NOR2 (N1715, N1712, N1391);
and AND3 (N1716, N1713, N1304, N230);
not NOT1 (N1717, N1700);
and AND2 (N1718, N1715, N1480);
buf BUF1 (N1719, N1709);
xor XOR2 (N1720, N1708, N1352);
xor XOR2 (N1721, N1694, N288);
nor NOR4 (N1722, N1719, N1063, N1021, N1197);
not NOT1 (N1723, N1717);
nand NAND2 (N1724, N1722, N1613);
or OR3 (N1725, N1710, N1579, N882);
and AND2 (N1726, N1721, N970);
buf BUF1 (N1727, N1725);
nand NAND4 (N1728, N1718, N906, N1102, N231);
not NOT1 (N1729, N1728);
and AND3 (N1730, N1723, N345, N1153);
buf BUF1 (N1731, N1702);
and AND2 (N1732, N1714, N371);
xor XOR2 (N1733, N1732, N736);
and AND4 (N1734, N1730, N690, N583, N1014);
xor XOR2 (N1735, N1731, N1148);
buf BUF1 (N1736, N1716);
xor XOR2 (N1737, N1724, N1192);
xor XOR2 (N1738, N1736, N357);
and AND4 (N1739, N1738, N1455, N1646, N953);
xor XOR2 (N1740, N1734, N1693);
buf BUF1 (N1741, N1729);
and AND4 (N1742, N1733, N669, N1600, N1055);
or OR2 (N1743, N1720, N638);
buf BUF1 (N1744, N1727);
not NOT1 (N1745, N1742);
nor NOR4 (N1746, N1726, N743, N1041, N1441);
nand NAND2 (N1747, N1737, N739);
and AND4 (N1748, N1735, N1134, N271, N1113);
buf BUF1 (N1749, N1743);
and AND2 (N1750, N1744, N539);
nand NAND3 (N1751, N1745, N378, N1373);
buf BUF1 (N1752, N1750);
buf BUF1 (N1753, N1748);
not NOT1 (N1754, N1739);
or OR2 (N1755, N1711, N1053);
xor XOR2 (N1756, N1741, N1499);
not NOT1 (N1757, N1756);
xor XOR2 (N1758, N1740, N33);
buf BUF1 (N1759, N1746);
xor XOR2 (N1760, N1747, N752);
or OR4 (N1761, N1755, N1213, N1230, N1726);
and AND2 (N1762, N1751, N255);
or OR2 (N1763, N1753, N680);
not NOT1 (N1764, N1754);
nor NOR2 (N1765, N1761, N1374);
or OR4 (N1766, N1762, N48, N181, N651);
nand NAND4 (N1767, N1765, N540, N461, N591);
buf BUF1 (N1768, N1757);
nand NAND4 (N1769, N1749, N1342, N221, N1168);
or OR4 (N1770, N1769, N687, N785, N522);
and AND3 (N1771, N1752, N1269, N1475);
or OR2 (N1772, N1763, N662);
xor XOR2 (N1773, N1759, N522);
and AND4 (N1774, N1772, N1224, N1394, N1759);
xor XOR2 (N1775, N1770, N1715);
xor XOR2 (N1776, N1758, N110);
not NOT1 (N1777, N1760);
nor NOR4 (N1778, N1768, N1735, N1296, N510);
and AND2 (N1779, N1764, N9);
not NOT1 (N1780, N1771);
buf BUF1 (N1781, N1780);
not NOT1 (N1782, N1774);
nor NOR4 (N1783, N1779, N477, N1088, N1250);
xor XOR2 (N1784, N1783, N682);
nor NOR4 (N1785, N1773, N440, N598, N834);
not NOT1 (N1786, N1766);
buf BUF1 (N1787, N1785);
nor NOR4 (N1788, N1781, N1197, N945, N1765);
or OR3 (N1789, N1787, N1427, N502);
or OR4 (N1790, N1788, N276, N1245, N227);
and AND4 (N1791, N1777, N191, N1192, N246);
nor NOR3 (N1792, N1767, N1690, N876);
nand NAND4 (N1793, N1791, N557, N553, N691);
and AND4 (N1794, N1782, N753, N1637, N699);
nor NOR4 (N1795, N1775, N424, N417, N814);
xor XOR2 (N1796, N1784, N1604);
nand NAND4 (N1797, N1796, N964, N1013, N713);
nand NAND2 (N1798, N1793, N1770);
or OR2 (N1799, N1794, N1011);
xor XOR2 (N1800, N1776, N1636);
not NOT1 (N1801, N1797);
not NOT1 (N1802, N1799);
or OR3 (N1803, N1802, N442, N1085);
buf BUF1 (N1804, N1803);
and AND2 (N1805, N1800, N949);
not NOT1 (N1806, N1804);
buf BUF1 (N1807, N1778);
xor XOR2 (N1808, N1786, N904);
nand NAND4 (N1809, N1801, N666, N648, N328);
not NOT1 (N1810, N1807);
or OR3 (N1811, N1795, N1341, N964);
and AND3 (N1812, N1810, N1053, N922);
and AND3 (N1813, N1805, N199, N66);
buf BUF1 (N1814, N1811);
nor NOR2 (N1815, N1806, N1710);
nor NOR4 (N1816, N1815, N1253, N233, N1741);
xor XOR2 (N1817, N1816, N1376);
and AND3 (N1818, N1808, N699, N1379);
xor XOR2 (N1819, N1814, N1696);
and AND2 (N1820, N1809, N709);
nor NOR4 (N1821, N1817, N1047, N325, N709);
nor NOR2 (N1822, N1798, N655);
nand NAND3 (N1823, N1820, N1719, N925);
xor XOR2 (N1824, N1789, N520);
not NOT1 (N1825, N1813);
and AND3 (N1826, N1818, N299, N811);
nand NAND2 (N1827, N1790, N929);
nand NAND3 (N1828, N1819, N1729, N231);
xor XOR2 (N1829, N1824, N1372);
nor NOR4 (N1830, N1825, N546, N317, N584);
nor NOR2 (N1831, N1822, N25);
not NOT1 (N1832, N1829);
or OR3 (N1833, N1812, N1717, N1239);
not NOT1 (N1834, N1827);
buf BUF1 (N1835, N1826);
and AND2 (N1836, N1821, N530);
and AND2 (N1837, N1830, N1633);
nor NOR4 (N1838, N1837, N96, N1721, N1464);
nor NOR3 (N1839, N1832, N472, N1445);
and AND4 (N1840, N1838, N835, N781, N640);
and AND3 (N1841, N1835, N1813, N691);
or OR4 (N1842, N1833, N1069, N494, N385);
nand NAND2 (N1843, N1841, N1036);
buf BUF1 (N1844, N1823);
nor NOR2 (N1845, N1840, N229);
and AND4 (N1846, N1844, N1298, N942, N112);
nor NOR4 (N1847, N1842, N1061, N1572, N1637);
not NOT1 (N1848, N1847);
buf BUF1 (N1849, N1792);
nor NOR3 (N1850, N1834, N1266, N1170);
nand NAND4 (N1851, N1828, N497, N1186, N1298);
nand NAND3 (N1852, N1839, N829, N1181);
not NOT1 (N1853, N1843);
not NOT1 (N1854, N1836);
nand NAND3 (N1855, N1831, N1445, N395);
nand NAND3 (N1856, N1853, N484, N49);
nand NAND4 (N1857, N1856, N7, N1567, N668);
not NOT1 (N1858, N1845);
nor NOR4 (N1859, N1855, N1123, N513, N916);
xor XOR2 (N1860, N1850, N1842);
xor XOR2 (N1861, N1860, N1040);
xor XOR2 (N1862, N1846, N51);
or OR4 (N1863, N1859, N378, N1296, N1370);
or OR2 (N1864, N1863, N31);
and AND2 (N1865, N1858, N1844);
and AND3 (N1866, N1854, N1591, N1002);
not NOT1 (N1867, N1865);
nand NAND4 (N1868, N1862, N137, N507, N1763);
nand NAND4 (N1869, N1868, N1803, N65, N825);
nand NAND2 (N1870, N1849, N1104);
or OR3 (N1871, N1851, N29, N356);
or OR2 (N1872, N1870, N575);
and AND2 (N1873, N1861, N1183);
not NOT1 (N1874, N1869);
and AND3 (N1875, N1867, N1350, N1812);
nor NOR3 (N1876, N1873, N1857, N1207);
buf BUF1 (N1877, N914);
xor XOR2 (N1878, N1866, N818);
or OR3 (N1879, N1878, N1081, N987);
buf BUF1 (N1880, N1872);
buf BUF1 (N1881, N1876);
buf BUF1 (N1882, N1874);
and AND2 (N1883, N1882, N666);
and AND2 (N1884, N1864, N1741);
xor XOR2 (N1885, N1879, N1403);
nand NAND2 (N1886, N1848, N1867);
or OR2 (N1887, N1881, N54);
nor NOR4 (N1888, N1877, N755, N1210, N768);
nand NAND2 (N1889, N1852, N797);
nor NOR3 (N1890, N1884, N991, N1757);
xor XOR2 (N1891, N1875, N400);
not NOT1 (N1892, N1891);
nor NOR3 (N1893, N1889, N928, N1877);
nand NAND3 (N1894, N1885, N45, N525);
not NOT1 (N1895, N1880);
buf BUF1 (N1896, N1895);
and AND4 (N1897, N1886, N1866, N373, N1683);
xor XOR2 (N1898, N1888, N858);
buf BUF1 (N1899, N1871);
buf BUF1 (N1900, N1896);
buf BUF1 (N1901, N1898);
buf BUF1 (N1902, N1883);
not NOT1 (N1903, N1890);
buf BUF1 (N1904, N1892);
nand NAND2 (N1905, N1887, N330);
not NOT1 (N1906, N1893);
or OR3 (N1907, N1905, N1373, N601);
and AND2 (N1908, N1903, N476);
or OR3 (N1909, N1900, N60, N1052);
nor NOR2 (N1910, N1897, N912);
and AND2 (N1911, N1894, N1472);
not NOT1 (N1912, N1901);
not NOT1 (N1913, N1906);
nand NAND3 (N1914, N1912, N1178, N611);
and AND2 (N1915, N1899, N61);
buf BUF1 (N1916, N1914);
nand NAND4 (N1917, N1913, N1910, N1505, N865);
nor NOR3 (N1918, N766, N634, N433);
not NOT1 (N1919, N1907);
xor XOR2 (N1920, N1902, N502);
nand NAND2 (N1921, N1915, N174);
and AND2 (N1922, N1917, N1869);
xor XOR2 (N1923, N1904, N1620);
nor NOR3 (N1924, N1920, N1390, N1698);
buf BUF1 (N1925, N1921);
nor NOR4 (N1926, N1918, N804, N1085, N1516);
nand NAND2 (N1927, N1916, N1777);
xor XOR2 (N1928, N1909, N870);
and AND2 (N1929, N1928, N1107);
nor NOR4 (N1930, N1926, N851, N1232, N41);
buf BUF1 (N1931, N1927);
and AND4 (N1932, N1931, N1844, N1077, N1207);
not NOT1 (N1933, N1922);
or OR4 (N1934, N1925, N1651, N923, N312);
or OR2 (N1935, N1930, N1560);
nor NOR3 (N1936, N1908, N1857, N282);
nand NAND3 (N1937, N1919, N1451, N450);
and AND3 (N1938, N1936, N1527, N445);
nand NAND4 (N1939, N1935, N1465, N694, N188);
xor XOR2 (N1940, N1938, N1521);
xor XOR2 (N1941, N1940, N587);
buf BUF1 (N1942, N1929);
nor NOR4 (N1943, N1939, N1096, N564, N258);
buf BUF1 (N1944, N1942);
nand NAND2 (N1945, N1933, N1713);
or OR3 (N1946, N1932, N718, N1250);
nand NAND3 (N1947, N1944, N245, N117);
not NOT1 (N1948, N1924);
buf BUF1 (N1949, N1948);
and AND3 (N1950, N1943, N1339, N937);
nor NOR2 (N1951, N1947, N658);
or OR4 (N1952, N1951, N1021, N1226, N33);
or OR4 (N1953, N1941, N1104, N1666, N719);
or OR4 (N1954, N1946, N673, N32, N58);
or OR2 (N1955, N1949, N829);
not NOT1 (N1956, N1952);
xor XOR2 (N1957, N1954, N1591);
buf BUF1 (N1958, N1956);
not NOT1 (N1959, N1950);
nor NOR3 (N1960, N1934, N1109, N1586);
nand NAND4 (N1961, N1923, N1622, N136, N709);
not NOT1 (N1962, N1945);
or OR2 (N1963, N1957, N750);
xor XOR2 (N1964, N1962, N790);
buf BUF1 (N1965, N1964);
nand NAND2 (N1966, N1959, N748);
nor NOR3 (N1967, N1965, N96, N615);
nand NAND3 (N1968, N1963, N850, N1538);
xor XOR2 (N1969, N1961, N239);
and AND4 (N1970, N1966, N620, N1065, N655);
nand NAND4 (N1971, N1969, N873, N539, N1697);
nor NOR3 (N1972, N1911, N1508, N491);
nand NAND4 (N1973, N1967, N807, N762, N1413);
xor XOR2 (N1974, N1972, N1937);
not NOT1 (N1975, N1142);
or OR3 (N1976, N1968, N1374, N212);
buf BUF1 (N1977, N1958);
buf BUF1 (N1978, N1953);
nand NAND4 (N1979, N1973, N9, N1538, N1392);
nand NAND4 (N1980, N1976, N554, N1565, N218);
nand NAND3 (N1981, N1960, N285, N335);
not NOT1 (N1982, N1977);
not NOT1 (N1983, N1980);
not NOT1 (N1984, N1955);
buf BUF1 (N1985, N1983);
nor NOR2 (N1986, N1981, N10);
and AND2 (N1987, N1984, N986);
nor NOR4 (N1988, N1978, N399, N1454, N820);
or OR2 (N1989, N1970, N1607);
nand NAND4 (N1990, N1985, N1927, N647, N1448);
and AND4 (N1991, N1982, N1105, N1198, N444);
not NOT1 (N1992, N1988);
buf BUF1 (N1993, N1992);
not NOT1 (N1994, N1987);
nand NAND4 (N1995, N1991, N911, N1645, N14);
and AND3 (N1996, N1986, N1422, N1270);
and AND3 (N1997, N1996, N1705, N1096);
or OR3 (N1998, N1993, N1661, N468);
buf BUF1 (N1999, N1998);
buf BUF1 (N2000, N1974);
or OR2 (N2001, N1997, N1245);
and AND2 (N2002, N2000, N833);
xor XOR2 (N2003, N1989, N970);
nor NOR3 (N2004, N1971, N778, N1427);
not NOT1 (N2005, N2001);
nand NAND4 (N2006, N1979, N1438, N908, N1858);
and AND3 (N2007, N2006, N558, N35);
not NOT1 (N2008, N1999);
not NOT1 (N2009, N2004);
nand NAND2 (N2010, N1990, N1705);
nand NAND2 (N2011, N2003, N1345);
xor XOR2 (N2012, N1975, N1807);
not NOT1 (N2013, N1995);
or OR2 (N2014, N2007, N949);
nand NAND3 (N2015, N2014, N494, N1126);
and AND3 (N2016, N2002, N1926, N1247);
and AND2 (N2017, N2009, N190);
not NOT1 (N2018, N2011);
and AND3 (N2019, N2018, N1646, N211);
nor NOR4 (N2020, N2016, N889, N197, N1129);
or OR2 (N2021, N1994, N1628);
and AND3 (N2022, N2015, N1977, N37);
buf BUF1 (N2023, N2017);
nor NOR3 (N2024, N2022, N444, N1320);
nor NOR4 (N2025, N2005, N823, N598, N1345);
not NOT1 (N2026, N2010);
buf BUF1 (N2027, N2008);
nand NAND4 (N2028, N2027, N1085, N1783, N1468);
and AND2 (N2029, N2020, N157);
or OR4 (N2030, N2028, N122, N1263, N573);
nor NOR3 (N2031, N2013, N902, N1130);
xor XOR2 (N2032, N2026, N1075);
buf BUF1 (N2033, N2032);
and AND3 (N2034, N2024, N1885, N1668);
and AND4 (N2035, N2030, N393, N495, N1108);
or OR2 (N2036, N2023, N30);
and AND4 (N2037, N2025, N1871, N607, N584);
xor XOR2 (N2038, N2029, N1154);
and AND2 (N2039, N2036, N631);
nor NOR2 (N2040, N2019, N226);
not NOT1 (N2041, N2040);
nand NAND3 (N2042, N2012, N1047, N510);
xor XOR2 (N2043, N2031, N1147);
and AND4 (N2044, N2041, N931, N1254, N63);
not NOT1 (N2045, N2044);
and AND2 (N2046, N2043, N1030);
buf BUF1 (N2047, N2045);
and AND4 (N2048, N2035, N994, N35, N1152);
and AND4 (N2049, N2038, N1517, N323, N528);
and AND4 (N2050, N2037, N837, N1800, N43);
nand NAND2 (N2051, N2033, N1555);
xor XOR2 (N2052, N2048, N1148);
buf BUF1 (N2053, N2050);
buf BUF1 (N2054, N2052);
not NOT1 (N2055, N2051);
nand NAND2 (N2056, N2042, N966);
not NOT1 (N2057, N2055);
buf BUF1 (N2058, N2021);
nor NOR3 (N2059, N2057, N1560, N1661);
and AND4 (N2060, N2056, N451, N1894, N602);
xor XOR2 (N2061, N2039, N1770);
not NOT1 (N2062, N2054);
and AND4 (N2063, N2053, N448, N1862, N1824);
nor NOR2 (N2064, N2063, N416);
and AND4 (N2065, N2062, N191, N935, N592);
nand NAND2 (N2066, N2046, N308);
nand NAND4 (N2067, N2064, N55, N1453, N1822);
or OR3 (N2068, N2059, N588, N1101);
buf BUF1 (N2069, N2058);
and AND4 (N2070, N2061, N418, N29, N1546);
not NOT1 (N2071, N2066);
buf BUF1 (N2072, N2067);
not NOT1 (N2073, N2034);
or OR3 (N2074, N2069, N1158, N1700);
buf BUF1 (N2075, N2074);
or OR2 (N2076, N2060, N1937);
buf BUF1 (N2077, N2073);
xor XOR2 (N2078, N2076, N1632);
nand NAND3 (N2079, N2071, N1285, N1393);
nand NAND3 (N2080, N2068, N145, N100);
or OR4 (N2081, N2047, N879, N891, N835);
not NOT1 (N2082, N2077);
buf BUF1 (N2083, N2072);
buf BUF1 (N2084, N2078);
nand NAND3 (N2085, N2070, N158, N728);
xor XOR2 (N2086, N2065, N245);
xor XOR2 (N2087, N2079, N924);
nand NAND3 (N2088, N2087, N935, N1322);
xor XOR2 (N2089, N2088, N643);
nand NAND4 (N2090, N2049, N1815, N775, N341);
xor XOR2 (N2091, N2080, N500);
or OR3 (N2092, N2083, N1124, N387);
buf BUF1 (N2093, N2089);
or OR4 (N2094, N2092, N961, N276, N585);
buf BUF1 (N2095, N2091);
nand NAND4 (N2096, N2093, N1917, N1740, N1576);
or OR2 (N2097, N2081, N456);
nand NAND4 (N2098, N2082, N1608, N1131, N1163);
not NOT1 (N2099, N2094);
nor NOR4 (N2100, N2086, N1566, N406, N1795);
nor NOR2 (N2101, N2098, N1968);
nor NOR4 (N2102, N2084, N733, N503, N668);
or OR4 (N2103, N2097, N1839, N1531, N2006);
and AND3 (N2104, N2096, N6, N1514);
xor XOR2 (N2105, N2085, N900);
or OR2 (N2106, N2101, N833);
not NOT1 (N2107, N2075);
or OR3 (N2108, N2104, N123, N2100);
and AND4 (N2109, N816, N684, N1128, N1417);
not NOT1 (N2110, N2099);
nand NAND4 (N2111, N2103, N1124, N891, N1951);
xor XOR2 (N2112, N2109, N1237);
nand NAND2 (N2113, N2110, N857);
or OR2 (N2114, N2090, N288);
and AND4 (N2115, N2113, N1705, N765, N206);
or OR4 (N2116, N2106, N2066, N540, N1966);
xor XOR2 (N2117, N2114, N531);
nor NOR2 (N2118, N2095, N250);
and AND2 (N2119, N2105, N1253);
buf BUF1 (N2120, N2112);
or OR4 (N2121, N2120, N1277, N1989, N679);
and AND3 (N2122, N2107, N703, N699);
not NOT1 (N2123, N2116);
or OR3 (N2124, N2123, N2098, N1359);
or OR2 (N2125, N2122, N1849);
buf BUF1 (N2126, N2111);
or OR2 (N2127, N2115, N213);
not NOT1 (N2128, N2124);
nand NAND3 (N2129, N2118, N761, N1070);
nand NAND4 (N2130, N2108, N332, N1690, N405);
not NOT1 (N2131, N2126);
nand NAND4 (N2132, N2121, N1193, N2083, N1087);
and AND4 (N2133, N2132, N1393, N2066, N690);
buf BUF1 (N2134, N2133);
nor NOR3 (N2135, N2131, N795, N1417);
not NOT1 (N2136, N2119);
or OR2 (N2137, N2127, N2010);
and AND4 (N2138, N2102, N2057, N968, N1935);
not NOT1 (N2139, N2125);
or OR3 (N2140, N2139, N1691, N1115);
or OR2 (N2141, N2128, N1289);
buf BUF1 (N2142, N2137);
and AND3 (N2143, N2135, N1793, N1089);
and AND3 (N2144, N2130, N970, N2102);
and AND4 (N2145, N2144, N363, N1261, N424);
or OR4 (N2146, N2136, N240, N1990, N1597);
and AND2 (N2147, N2117, N743);
buf BUF1 (N2148, N2134);
or OR2 (N2149, N2148, N1121);
nor NOR2 (N2150, N2141, N564);
buf BUF1 (N2151, N2150);
nand NAND4 (N2152, N2138, N722, N1469, N608);
buf BUF1 (N2153, N2129);
not NOT1 (N2154, N2152);
not NOT1 (N2155, N2147);
not NOT1 (N2156, N2154);
nor NOR4 (N2157, N2146, N1848, N732, N1805);
and AND3 (N2158, N2143, N150, N1460);
and AND2 (N2159, N2153, N766);
not NOT1 (N2160, N2151);
buf BUF1 (N2161, N2160);
or OR2 (N2162, N2158, N1872);
buf BUF1 (N2163, N2157);
buf BUF1 (N2164, N2140);
or OR3 (N2165, N2164, N118, N486);
nor NOR4 (N2166, N2162, N812, N1599, N1435);
or OR4 (N2167, N2165, N1690, N1771, N1035);
or OR3 (N2168, N2145, N440, N28);
and AND4 (N2169, N2155, N1917, N234, N1820);
not NOT1 (N2170, N2159);
nand NAND4 (N2171, N2169, N1796, N2018, N2004);
not NOT1 (N2172, N2161);
and AND3 (N2173, N2163, N1833, N1936);
nor NOR2 (N2174, N2166, N569);
and AND4 (N2175, N2174, N641, N510, N1720);
nand NAND3 (N2176, N2172, N1807, N1923);
and AND2 (N2177, N2173, N1892);
nand NAND3 (N2178, N2171, N17, N249);
or OR3 (N2179, N2175, N606, N1074);
or OR3 (N2180, N2168, N1162, N11);
and AND2 (N2181, N2149, N1136);
nor NOR2 (N2182, N2142, N1896);
nand NAND2 (N2183, N2167, N86);
not NOT1 (N2184, N2178);
buf BUF1 (N2185, N2182);
nand NAND3 (N2186, N2156, N593, N146);
not NOT1 (N2187, N2183);
nand NAND4 (N2188, N2179, N991, N2020, N1111);
buf BUF1 (N2189, N2185);
or OR2 (N2190, N2180, N939);
nor NOR2 (N2191, N2188, N1459);
not NOT1 (N2192, N2189);
nor NOR4 (N2193, N2184, N1179, N535, N31);
nor NOR4 (N2194, N2176, N319, N1838, N268);
and AND2 (N2195, N2191, N1423);
buf BUF1 (N2196, N2181);
not NOT1 (N2197, N2196);
xor XOR2 (N2198, N2195, N1764);
nor NOR3 (N2199, N2177, N1558, N1503);
nor NOR3 (N2200, N2193, N1016, N2019);
or OR4 (N2201, N2199, N1796, N74, N1892);
nor NOR2 (N2202, N2192, N1229);
nor NOR2 (N2203, N2198, N1384);
buf BUF1 (N2204, N2194);
buf BUF1 (N2205, N2204);
and AND3 (N2206, N2187, N846, N510);
and AND4 (N2207, N2186, N1534, N1013, N609);
nand NAND2 (N2208, N2190, N1152);
or OR3 (N2209, N2207, N942, N2153);
not NOT1 (N2210, N2209);
nor NOR4 (N2211, N2202, N2041, N170, N1605);
not NOT1 (N2212, N2211);
and AND2 (N2213, N2200, N1974);
or OR3 (N2214, N2206, N622, N553);
xor XOR2 (N2215, N2205, N1954);
nor NOR2 (N2216, N2201, N1625);
not NOT1 (N2217, N2197);
xor XOR2 (N2218, N2213, N1934);
and AND3 (N2219, N2215, N433, N1610);
xor XOR2 (N2220, N2208, N1556);
and AND3 (N2221, N2217, N90, N580);
and AND4 (N2222, N2220, N2080, N1310, N1472);
nand NAND3 (N2223, N2210, N1960, N1942);
buf BUF1 (N2224, N2203);
nor NOR4 (N2225, N2214, N280, N1816, N1963);
buf BUF1 (N2226, N2219);
xor XOR2 (N2227, N2216, N1577);
nor NOR4 (N2228, N2226, N1194, N339, N641);
nand NAND2 (N2229, N2227, N1207);
buf BUF1 (N2230, N2212);
buf BUF1 (N2231, N2225);
nor NOR4 (N2232, N2170, N1792, N2009, N927);
nor NOR4 (N2233, N2232, N1251, N107, N1822);
not NOT1 (N2234, N2231);
xor XOR2 (N2235, N2234, N2186);
nor NOR4 (N2236, N2218, N619, N1006, N1277);
not NOT1 (N2237, N2236);
xor XOR2 (N2238, N2229, N1697);
xor XOR2 (N2239, N2237, N1296);
not NOT1 (N2240, N2221);
xor XOR2 (N2241, N2240, N1108);
and AND4 (N2242, N2222, N166, N1733, N67);
buf BUF1 (N2243, N2233);
and AND3 (N2244, N2223, N2196, N1721);
xor XOR2 (N2245, N2230, N924);
and AND3 (N2246, N2238, N488, N1292);
not NOT1 (N2247, N2228);
xor XOR2 (N2248, N2246, N142);
xor XOR2 (N2249, N2244, N103);
buf BUF1 (N2250, N2249);
not NOT1 (N2251, N2239);
xor XOR2 (N2252, N2247, N1295);
and AND3 (N2253, N2241, N141, N361);
and AND3 (N2254, N2242, N1940, N1570);
and AND2 (N2255, N2235, N1572);
or OR2 (N2256, N2254, N943);
and AND3 (N2257, N2251, N823, N1975);
xor XOR2 (N2258, N2243, N30);
xor XOR2 (N2259, N2224, N1446);
xor XOR2 (N2260, N2252, N1199);
xor XOR2 (N2261, N2253, N239);
xor XOR2 (N2262, N2250, N86);
xor XOR2 (N2263, N2248, N1574);
and AND2 (N2264, N2260, N1122);
nand NAND2 (N2265, N2258, N855);
buf BUF1 (N2266, N2259);
not NOT1 (N2267, N2257);
not NOT1 (N2268, N2266);
not NOT1 (N2269, N2256);
buf BUF1 (N2270, N2262);
xor XOR2 (N2271, N2267, N1841);
buf BUF1 (N2272, N2269);
or OR4 (N2273, N2268, N487, N522, N446);
nor NOR2 (N2274, N2261, N129);
not NOT1 (N2275, N2270);
buf BUF1 (N2276, N2264);
buf BUF1 (N2277, N2275);
not NOT1 (N2278, N2255);
or OR3 (N2279, N2272, N1991, N284);
and AND4 (N2280, N2263, N128, N1836, N1666);
and AND4 (N2281, N2277, N402, N1713, N404);
buf BUF1 (N2282, N2271);
xor XOR2 (N2283, N2276, N1898);
nor NOR4 (N2284, N2278, N386, N1521, N821);
xor XOR2 (N2285, N2284, N285);
nand NAND4 (N2286, N2285, N2050, N259, N176);
xor XOR2 (N2287, N2282, N348);
nand NAND2 (N2288, N2265, N1994);
not NOT1 (N2289, N2280);
nand NAND4 (N2290, N2245, N2117, N2219, N253);
buf BUF1 (N2291, N2287);
buf BUF1 (N2292, N2279);
not NOT1 (N2293, N2288);
and AND3 (N2294, N2293, N1413, N626);
and AND2 (N2295, N2292, N1141);
xor XOR2 (N2296, N2274, N1582);
and AND3 (N2297, N2273, N1378, N1743);
and AND3 (N2298, N2281, N2223, N1040);
and AND2 (N2299, N2294, N898);
or OR2 (N2300, N2286, N423);
xor XOR2 (N2301, N2296, N1707);
xor XOR2 (N2302, N2301, N1920);
nor NOR3 (N2303, N2297, N895, N753);
not NOT1 (N2304, N2298);
and AND2 (N2305, N2304, N2183);
buf BUF1 (N2306, N2289);
nand NAND3 (N2307, N2283, N2119, N80);
not NOT1 (N2308, N2305);
buf BUF1 (N2309, N2308);
xor XOR2 (N2310, N2299, N116);
nand NAND4 (N2311, N2302, N1058, N1221, N1890);
and AND2 (N2312, N2307, N979);
nand NAND3 (N2313, N2290, N797, N1214);
buf BUF1 (N2314, N2306);
not NOT1 (N2315, N2314);
not NOT1 (N2316, N2309);
or OR4 (N2317, N2311, N440, N739, N1670);
buf BUF1 (N2318, N2295);
and AND4 (N2319, N2313, N2201, N1503, N490);
nor NOR4 (N2320, N2317, N1690, N2240, N1866);
or OR3 (N2321, N2318, N70, N2099);
not NOT1 (N2322, N2316);
or OR2 (N2323, N2300, N1516);
or OR3 (N2324, N2291, N1293, N1337);
or OR2 (N2325, N2310, N1072);
nand NAND3 (N2326, N2325, N881, N2284);
and AND2 (N2327, N2323, N320);
nand NAND2 (N2328, N2321, N1043);
nor NOR4 (N2329, N2320, N564, N1199, N962);
nor NOR2 (N2330, N2312, N439);
nand NAND2 (N2331, N2322, N2102);
or OR3 (N2332, N2330, N2065, N559);
nor NOR3 (N2333, N2331, N301, N1265);
nor NOR2 (N2334, N2333, N1234);
buf BUF1 (N2335, N2326);
and AND3 (N2336, N2327, N625, N1383);
nor NOR3 (N2337, N2328, N1858, N1071);
xor XOR2 (N2338, N2332, N1933);
nand NAND3 (N2339, N2324, N470, N513);
xor XOR2 (N2340, N2303, N994);
not NOT1 (N2341, N2334);
nand NAND4 (N2342, N2337, N1836, N1347, N358);
or OR3 (N2343, N2319, N80, N859);
nor NOR2 (N2344, N2342, N1683);
not NOT1 (N2345, N2343);
or OR2 (N2346, N2315, N832);
nor NOR3 (N2347, N2340, N1795, N1278);
not NOT1 (N2348, N2344);
nor NOR3 (N2349, N2345, N723, N1682);
xor XOR2 (N2350, N2335, N1447);
buf BUF1 (N2351, N2329);
or OR4 (N2352, N2349, N180, N1957, N840);
nand NAND4 (N2353, N2351, N1815, N638, N2267);
nor NOR4 (N2354, N2346, N1895, N1179, N1289);
buf BUF1 (N2355, N2347);
nand NAND4 (N2356, N2348, N362, N257, N403);
not NOT1 (N2357, N2341);
nor NOR3 (N2358, N2336, N1032, N1674);
or OR2 (N2359, N2354, N714);
xor XOR2 (N2360, N2352, N2340);
nand NAND2 (N2361, N2350, N2225);
not NOT1 (N2362, N2355);
or OR4 (N2363, N2358, N373, N307, N1374);
buf BUF1 (N2364, N2363);
not NOT1 (N2365, N2353);
not NOT1 (N2366, N2361);
or OR4 (N2367, N2365, N296, N708, N41);
xor XOR2 (N2368, N2360, N814);
xor XOR2 (N2369, N2368, N852);
xor XOR2 (N2370, N2364, N1109);
and AND4 (N2371, N2339, N1409, N1006, N1397);
nand NAND2 (N2372, N2371, N1538);
nand NAND2 (N2373, N2356, N1536);
not NOT1 (N2374, N2357);
buf BUF1 (N2375, N2338);
and AND3 (N2376, N2373, N1643, N1704);
nor NOR3 (N2377, N2359, N66, N2307);
or OR3 (N2378, N2375, N349, N235);
buf BUF1 (N2379, N2362);
not NOT1 (N2380, N2369);
nor NOR2 (N2381, N2366, N87);
and AND4 (N2382, N2378, N1092, N398, N1480);
not NOT1 (N2383, N2370);
nand NAND4 (N2384, N2374, N1907, N810, N892);
buf BUF1 (N2385, N2381);
or OR4 (N2386, N2372, N1637, N2143, N1515);
xor XOR2 (N2387, N2385, N1099);
or OR3 (N2388, N2386, N799, N1077);
xor XOR2 (N2389, N2387, N2047);
buf BUF1 (N2390, N2379);
xor XOR2 (N2391, N2377, N1945);
or OR3 (N2392, N2367, N2216, N2358);
nor NOR2 (N2393, N2392, N2361);
nand NAND3 (N2394, N2384, N591, N928);
nor NOR2 (N2395, N2393, N1627);
nand NAND2 (N2396, N2394, N978);
buf BUF1 (N2397, N2389);
xor XOR2 (N2398, N2397, N34);
nand NAND4 (N2399, N2398, N1274, N747, N1822);
nand NAND3 (N2400, N2391, N2227, N1134);
nor NOR3 (N2401, N2399, N2309, N1495);
and AND4 (N2402, N2400, N374, N1021, N331);
buf BUF1 (N2403, N2401);
buf BUF1 (N2404, N2376);
buf BUF1 (N2405, N2390);
nor NOR3 (N2406, N2395, N1094, N2260);
xor XOR2 (N2407, N2406, N618);
not NOT1 (N2408, N2382);
or OR4 (N2409, N2396, N2084, N786, N2395);
buf BUF1 (N2410, N2407);
or OR2 (N2411, N2380, N1052);
or OR3 (N2412, N2409, N422, N814);
buf BUF1 (N2413, N2404);
xor XOR2 (N2414, N2410, N1528);
buf BUF1 (N2415, N2388);
buf BUF1 (N2416, N2415);
buf BUF1 (N2417, N2416);
buf BUF1 (N2418, N2412);
nor NOR3 (N2419, N2411, N998, N2364);
nand NAND2 (N2420, N2408, N816);
and AND2 (N2421, N2419, N82);
not NOT1 (N2422, N2383);
or OR2 (N2423, N2405, N991);
xor XOR2 (N2424, N2403, N516);
buf BUF1 (N2425, N2420);
and AND3 (N2426, N2414, N245, N2266);
nor NOR3 (N2427, N2425, N433, N2302);
nor NOR3 (N2428, N2422, N1597, N2114);
xor XOR2 (N2429, N2426, N1082);
not NOT1 (N2430, N2402);
not NOT1 (N2431, N2417);
or OR3 (N2432, N2431, N860, N1165);
not NOT1 (N2433, N2418);
not NOT1 (N2434, N2429);
xor XOR2 (N2435, N2424, N1323);
not NOT1 (N2436, N2423);
not NOT1 (N2437, N2432);
and AND3 (N2438, N2436, N1482, N1511);
not NOT1 (N2439, N2427);
nor NOR4 (N2440, N2428, N1934, N685, N2224);
buf BUF1 (N2441, N2430);
nand NAND2 (N2442, N2437, N584);
buf BUF1 (N2443, N2439);
nor NOR3 (N2444, N2438, N2125, N420);
xor XOR2 (N2445, N2434, N313);
xor XOR2 (N2446, N2421, N1990);
or OR3 (N2447, N2440, N374, N2102);
buf BUF1 (N2448, N2443);
not NOT1 (N2449, N2445);
not NOT1 (N2450, N2442);
and AND4 (N2451, N2433, N2294, N871, N955);
nor NOR4 (N2452, N2447, N967, N82, N970);
and AND4 (N2453, N2441, N939, N737, N37);
or OR2 (N2454, N2446, N346);
xor XOR2 (N2455, N2453, N1722);
not NOT1 (N2456, N2455);
and AND4 (N2457, N2452, N1003, N908, N2434);
and AND3 (N2458, N2457, N1783, N1348);
xor XOR2 (N2459, N2458, N443);
nand NAND4 (N2460, N2456, N2209, N1181, N764);
xor XOR2 (N2461, N2449, N2108);
and AND3 (N2462, N2435, N159, N2452);
not NOT1 (N2463, N2459);
nor NOR4 (N2464, N2448, N883, N1983, N1742);
xor XOR2 (N2465, N2451, N609);
nor NOR2 (N2466, N2454, N1319);
xor XOR2 (N2467, N2460, N636);
buf BUF1 (N2468, N2464);
and AND3 (N2469, N2465, N2038, N988);
or OR4 (N2470, N2461, N1783, N1412, N69);
or OR4 (N2471, N2469, N758, N1628, N176);
or OR3 (N2472, N2470, N150, N1238);
xor XOR2 (N2473, N2467, N1983);
or OR2 (N2474, N2413, N1804);
and AND3 (N2475, N2450, N40, N2214);
not NOT1 (N2476, N2468);
and AND4 (N2477, N2476, N1710, N819, N553);
nand NAND3 (N2478, N2463, N498, N1820);
nand NAND4 (N2479, N2473, N2190, N1548, N1158);
xor XOR2 (N2480, N2478, N354);
nand NAND4 (N2481, N2475, N1027, N74, N885);
nand NAND2 (N2482, N2474, N1525);
and AND2 (N2483, N2471, N17);
nand NAND2 (N2484, N2482, N176);
buf BUF1 (N2485, N2480);
buf BUF1 (N2486, N2481);
buf BUF1 (N2487, N2479);
nor NOR4 (N2488, N2477, N1589, N964, N1745);
nor NOR4 (N2489, N2487, N1515, N1786, N578);
nor NOR4 (N2490, N2483, N649, N1015, N2225);
and AND4 (N2491, N2490, N2049, N26, N1425);
not NOT1 (N2492, N2488);
and AND2 (N2493, N2472, N1489);
buf BUF1 (N2494, N2486);
nor NOR4 (N2495, N2489, N2033, N927, N975);
or OR3 (N2496, N2462, N712, N1119);
not NOT1 (N2497, N2492);
and AND2 (N2498, N2484, N1845);
xor XOR2 (N2499, N2444, N2338);
buf BUF1 (N2500, N2494);
or OR2 (N2501, N2491, N951);
nor NOR2 (N2502, N2500, N1301);
buf BUF1 (N2503, N2466);
or OR2 (N2504, N2498, N1869);
nand NAND3 (N2505, N2485, N848, N2032);
xor XOR2 (N2506, N2497, N2281);
nor NOR4 (N2507, N2504, N1506, N146, N1251);
nor NOR2 (N2508, N2502, N1037);
nand NAND2 (N2509, N2493, N1384);
or OR3 (N2510, N2501, N1712, N1416);
or OR2 (N2511, N2503, N877);
nor NOR4 (N2512, N2505, N275, N1376, N152);
and AND3 (N2513, N2507, N1650, N151);
not NOT1 (N2514, N2509);
xor XOR2 (N2515, N2496, N328);
nand NAND2 (N2516, N2513, N2370);
nand NAND4 (N2517, N2516, N1273, N702, N1344);
nor NOR4 (N2518, N2511, N1636, N523, N2127);
nand NAND4 (N2519, N2510, N791, N921, N1211);
not NOT1 (N2520, N2515);
xor XOR2 (N2521, N2499, N295);
nor NOR3 (N2522, N2520, N275, N2305);
nor NOR3 (N2523, N2521, N1483, N1512);
nand NAND3 (N2524, N2518, N955, N1738);
xor XOR2 (N2525, N2524, N1666);
xor XOR2 (N2526, N2512, N1762);
nand NAND2 (N2527, N2517, N129);
xor XOR2 (N2528, N2514, N2365);
not NOT1 (N2529, N2495);
not NOT1 (N2530, N2506);
or OR3 (N2531, N2519, N818, N779);
nand NAND2 (N2532, N2530, N2319);
nor NOR2 (N2533, N2522, N555);
xor XOR2 (N2534, N2523, N1856);
xor XOR2 (N2535, N2533, N381);
xor XOR2 (N2536, N2535, N2069);
nand NAND2 (N2537, N2529, N885);
nor NOR2 (N2538, N2531, N1729);
xor XOR2 (N2539, N2538, N1011);
buf BUF1 (N2540, N2534);
nor NOR4 (N2541, N2525, N645, N835, N1724);
xor XOR2 (N2542, N2532, N2177);
nor NOR3 (N2543, N2540, N2289, N1675);
xor XOR2 (N2544, N2536, N1606);
nor NOR3 (N2545, N2508, N608, N986);
not NOT1 (N2546, N2539);
xor XOR2 (N2547, N2537, N659);
nand NAND3 (N2548, N2527, N683, N1132);
not NOT1 (N2549, N2545);
nor NOR3 (N2550, N2547, N214, N1587);
nand NAND2 (N2551, N2542, N1444);
xor XOR2 (N2552, N2526, N1178);
nor NOR4 (N2553, N2548, N2250, N1353, N1980);
xor XOR2 (N2554, N2549, N1886);
xor XOR2 (N2555, N2550, N1613);
and AND4 (N2556, N2554, N1325, N1174, N1112);
nand NAND2 (N2557, N2555, N512);
xor XOR2 (N2558, N2544, N1976);
and AND3 (N2559, N2528, N2148, N2076);
nand NAND3 (N2560, N2558, N617, N1073);
and AND4 (N2561, N2553, N33, N1484, N1368);
xor XOR2 (N2562, N2551, N1757);
nand NAND4 (N2563, N2559, N981, N2549, N1905);
or OR3 (N2564, N2541, N1872, N249);
or OR4 (N2565, N2546, N1178, N1516, N2198);
buf BUF1 (N2566, N2564);
xor XOR2 (N2567, N2543, N1770);
and AND4 (N2568, N2566, N177, N1975, N437);
nor NOR2 (N2569, N2561, N1785);
xor XOR2 (N2570, N2568, N1763);
and AND3 (N2571, N2560, N1222, N520);
not NOT1 (N2572, N2552);
and AND3 (N2573, N2569, N2507, N1428);
nand NAND4 (N2574, N2556, N2372, N885, N1846);
and AND3 (N2575, N2573, N1299, N1299);
xor XOR2 (N2576, N2571, N1254);
and AND4 (N2577, N2567, N408, N2372, N878);
nand NAND2 (N2578, N2565, N2268);
nand NAND2 (N2579, N2557, N73);
nor NOR3 (N2580, N2563, N2115, N1124);
nand NAND4 (N2581, N2579, N2230, N866, N641);
buf BUF1 (N2582, N2581);
xor XOR2 (N2583, N2575, N206);
nand NAND4 (N2584, N2577, N1568, N902, N238);
buf BUF1 (N2585, N2584);
or OR3 (N2586, N2580, N1462, N2271);
nor NOR2 (N2587, N2578, N1694);
and AND3 (N2588, N2574, N2528, N2328);
nor NOR2 (N2589, N2572, N2336);
or OR3 (N2590, N2576, N1285, N365);
nor NOR3 (N2591, N2588, N441, N221);
not NOT1 (N2592, N2570);
or OR3 (N2593, N2592, N614, N2427);
buf BUF1 (N2594, N2582);
or OR3 (N2595, N2593, N1311, N1765);
buf BUF1 (N2596, N2589);
nor NOR3 (N2597, N2583, N151, N766);
xor XOR2 (N2598, N2590, N165);
xor XOR2 (N2599, N2585, N303);
xor XOR2 (N2600, N2594, N1795);
or OR2 (N2601, N2586, N1732);
nor NOR3 (N2602, N2599, N1411, N1285);
and AND4 (N2603, N2595, N1389, N1604, N1008);
and AND4 (N2604, N2597, N1068, N591, N91);
and AND4 (N2605, N2587, N1668, N2442, N2214);
and AND3 (N2606, N2598, N346, N774);
xor XOR2 (N2607, N2602, N151);
nand NAND3 (N2608, N2605, N2264, N2524);
nand NAND4 (N2609, N2603, N928, N349, N2284);
not NOT1 (N2610, N2609);
buf BUF1 (N2611, N2606);
buf BUF1 (N2612, N2611);
not NOT1 (N2613, N2610);
nand NAND2 (N2614, N2608, N502);
and AND4 (N2615, N2604, N2147, N1016, N742);
buf BUF1 (N2616, N2562);
and AND2 (N2617, N2596, N2320);
nand NAND4 (N2618, N2614, N1789, N1861, N376);
and AND3 (N2619, N2607, N251, N866);
not NOT1 (N2620, N2591);
not NOT1 (N2621, N2620);
xor XOR2 (N2622, N2621, N2390);
not NOT1 (N2623, N2618);
xor XOR2 (N2624, N2619, N326);
not NOT1 (N2625, N2601);
not NOT1 (N2626, N2624);
nand NAND3 (N2627, N2613, N301, N1625);
xor XOR2 (N2628, N2612, N1232);
nand NAND2 (N2629, N2615, N573);
not NOT1 (N2630, N2623);
or OR2 (N2631, N2617, N2319);
not NOT1 (N2632, N2631);
nand NAND2 (N2633, N2600, N156);
and AND2 (N2634, N2629, N402);
and AND2 (N2635, N2630, N1929);
xor XOR2 (N2636, N2626, N2217);
and AND3 (N2637, N2625, N927, N556);
buf BUF1 (N2638, N2633);
not NOT1 (N2639, N2634);
xor XOR2 (N2640, N2637, N670);
and AND3 (N2641, N2627, N1025, N1237);
nor NOR3 (N2642, N2622, N1280, N46);
buf BUF1 (N2643, N2636);
or OR3 (N2644, N2628, N322, N1298);
nor NOR3 (N2645, N2639, N1815, N5);
or OR3 (N2646, N2632, N1605, N1651);
buf BUF1 (N2647, N2645);
buf BUF1 (N2648, N2646);
xor XOR2 (N2649, N2616, N1787);
and AND4 (N2650, N2638, N768, N1592, N229);
nor NOR3 (N2651, N2644, N2273, N1669);
nor NOR2 (N2652, N2650, N2210);
and AND2 (N2653, N2652, N683);
not NOT1 (N2654, N2647);
or OR4 (N2655, N2635, N346, N1818, N1989);
or OR3 (N2656, N2654, N749, N1501);
or OR2 (N2657, N2642, N1107);
buf BUF1 (N2658, N2641);
or OR4 (N2659, N2653, N554, N2540, N540);
nor NOR3 (N2660, N2655, N194, N957);
or OR2 (N2661, N2643, N568);
buf BUF1 (N2662, N2661);
xor XOR2 (N2663, N2662, N53);
xor XOR2 (N2664, N2660, N982);
and AND2 (N2665, N2663, N2213);
not NOT1 (N2666, N2657);
nand NAND4 (N2667, N2651, N660, N906, N2606);
nand NAND2 (N2668, N2666, N2429);
not NOT1 (N2669, N2665);
and AND3 (N2670, N2640, N526, N420);
nor NOR2 (N2671, N2670, N806);
or OR3 (N2672, N2658, N582, N2473);
nor NOR2 (N2673, N2672, N49);
and AND3 (N2674, N2664, N503, N609);
buf BUF1 (N2675, N2648);
and AND3 (N2676, N2674, N630, N1781);
xor XOR2 (N2677, N2667, N163);
nor NOR4 (N2678, N2656, N345, N2374, N394);
buf BUF1 (N2679, N2678);
nand NAND3 (N2680, N2673, N1635, N1898);
nor NOR4 (N2681, N2649, N1279, N2090, N367);
or OR3 (N2682, N2668, N1039, N1791);
buf BUF1 (N2683, N2669);
nand NAND2 (N2684, N2681, N1154);
and AND3 (N2685, N2677, N1816, N2358);
not NOT1 (N2686, N2671);
or OR4 (N2687, N2659, N105, N1370, N176);
not NOT1 (N2688, N2685);
or OR2 (N2689, N2679, N2525);
xor XOR2 (N2690, N2680, N610);
nor NOR4 (N2691, N2690, N309, N255, N1888);
nand NAND2 (N2692, N2691, N657);
nor NOR3 (N2693, N2687, N1646, N2307);
and AND2 (N2694, N2675, N593);
buf BUF1 (N2695, N2684);
buf BUF1 (N2696, N2682);
not NOT1 (N2697, N2689);
buf BUF1 (N2698, N2692);
or OR3 (N2699, N2688, N2088, N789);
nor NOR2 (N2700, N2694, N707);
nor NOR4 (N2701, N2697, N492, N937, N2072);
buf BUF1 (N2702, N2700);
buf BUF1 (N2703, N2698);
not NOT1 (N2704, N2686);
nand NAND4 (N2705, N2701, N1409, N1999, N1886);
buf BUF1 (N2706, N2705);
or OR4 (N2707, N2702, N1876, N1559, N2148);
nand NAND2 (N2708, N2704, N1419);
buf BUF1 (N2709, N2707);
nor NOR2 (N2710, N2703, N1249);
and AND4 (N2711, N2676, N2667, N2503, N2038);
buf BUF1 (N2712, N2711);
or OR3 (N2713, N2699, N897, N366);
or OR3 (N2714, N2693, N1843, N418);
or OR4 (N2715, N2712, N328, N1697, N1264);
buf BUF1 (N2716, N2715);
buf BUF1 (N2717, N2710);
buf BUF1 (N2718, N2714);
nor NOR3 (N2719, N2716, N2235, N2070);
buf BUF1 (N2720, N2683);
nand NAND3 (N2721, N2709, N1374, N1217);
or OR3 (N2722, N2719, N2334, N1900);
and AND3 (N2723, N2695, N1385, N1795);
xor XOR2 (N2724, N2720, N1386);
not NOT1 (N2725, N2713);
nand NAND3 (N2726, N2722, N2703, N275);
not NOT1 (N2727, N2726);
xor XOR2 (N2728, N2727, N701);
xor XOR2 (N2729, N2718, N1591);
or OR2 (N2730, N2696, N2277);
not NOT1 (N2731, N2723);
nor NOR2 (N2732, N2708, N1103);
or OR2 (N2733, N2721, N2466);
not NOT1 (N2734, N2732);
buf BUF1 (N2735, N2728);
nor NOR4 (N2736, N2735, N577, N91, N1262);
and AND4 (N2737, N2729, N2453, N1382, N85);
not NOT1 (N2738, N2706);
nand NAND2 (N2739, N2738, N1052);
nor NOR4 (N2740, N2737, N1384, N1133, N417);
nor NOR3 (N2741, N2736, N2520, N2443);
and AND4 (N2742, N2734, N1645, N971, N121);
nand NAND3 (N2743, N2733, N1322, N1887);
buf BUF1 (N2744, N2717);
buf BUF1 (N2745, N2744);
nor NOR3 (N2746, N2724, N1540, N904);
or OR4 (N2747, N2731, N2012, N1813, N801);
not NOT1 (N2748, N2747);
buf BUF1 (N2749, N2739);
nand NAND2 (N2750, N2749, N441);
or OR2 (N2751, N2743, N29);
nand NAND3 (N2752, N2740, N2292, N49);
or OR4 (N2753, N2730, N915, N827, N1196);
xor XOR2 (N2754, N2750, N1599);
not NOT1 (N2755, N2754);
xor XOR2 (N2756, N2725, N2610);
nand NAND3 (N2757, N2741, N1926, N670);
and AND2 (N2758, N2751, N2713);
or OR4 (N2759, N2756, N1321, N800, N158);
nor NOR4 (N2760, N2742, N2314, N1275, N842);
not NOT1 (N2761, N2745);
nor NOR3 (N2762, N2760, N1853, N1937);
xor XOR2 (N2763, N2746, N2328);
nor NOR3 (N2764, N2763, N520, N2291);
buf BUF1 (N2765, N2762);
not NOT1 (N2766, N2755);
not NOT1 (N2767, N2757);
nand NAND2 (N2768, N2759, N654);
or OR4 (N2769, N2766, N1782, N2575, N1958);
and AND3 (N2770, N2761, N49, N2408);
xor XOR2 (N2771, N2770, N279);
nor NOR4 (N2772, N2768, N717, N1635, N678);
nor NOR4 (N2773, N2753, N1986, N2031, N459);
nand NAND2 (N2774, N2758, N141);
nor NOR2 (N2775, N2767, N2362);
nor NOR2 (N2776, N2771, N2495);
xor XOR2 (N2777, N2769, N1726);
not NOT1 (N2778, N2772);
buf BUF1 (N2779, N2775);
not NOT1 (N2780, N2778);
and AND2 (N2781, N2752, N1761);
or OR4 (N2782, N2777, N1770, N404, N2163);
or OR2 (N2783, N2781, N1433);
and AND3 (N2784, N2779, N1715, N1516);
xor XOR2 (N2785, N2782, N262);
and AND2 (N2786, N2776, N2193);
not NOT1 (N2787, N2785);
and AND2 (N2788, N2787, N2428);
not NOT1 (N2789, N2783);
or OR4 (N2790, N2773, N2122, N102, N444);
xor XOR2 (N2791, N2774, N2099);
nor NOR3 (N2792, N2786, N2566, N2137);
buf BUF1 (N2793, N2748);
nand NAND3 (N2794, N2788, N311, N1463);
not NOT1 (N2795, N2765);
nor NOR3 (N2796, N2784, N1309, N134);
or OR2 (N2797, N2790, N1943);
not NOT1 (N2798, N2796);
buf BUF1 (N2799, N2793);
buf BUF1 (N2800, N2764);
xor XOR2 (N2801, N2780, N2112);
not NOT1 (N2802, N2794);
or OR2 (N2803, N2798, N660);
buf BUF1 (N2804, N2802);
nor NOR4 (N2805, N2801, N2561, N2046, N2089);
and AND3 (N2806, N2792, N1823, N976);
buf BUF1 (N2807, N2805);
xor XOR2 (N2808, N2795, N2251);
nand NAND3 (N2809, N2791, N2263, N1149);
nor NOR2 (N2810, N2808, N2608);
and AND2 (N2811, N2799, N2058);
and AND2 (N2812, N2803, N1773);
xor XOR2 (N2813, N2812, N640);
nand NAND3 (N2814, N2797, N339, N613);
nor NOR2 (N2815, N2813, N1732);
xor XOR2 (N2816, N2810, N2271);
and AND2 (N2817, N2815, N953);
nor NOR4 (N2818, N2809, N993, N354, N1758);
nand NAND3 (N2819, N2804, N1388, N1835);
nand NAND2 (N2820, N2806, N603);
nand NAND2 (N2821, N2817, N1709);
nor NOR3 (N2822, N2789, N2790, N2652);
xor XOR2 (N2823, N2821, N909);
nand NAND4 (N2824, N2814, N1389, N2689, N20);
and AND4 (N2825, N2823, N290, N1926, N2603);
nand NAND3 (N2826, N2822, N2369, N1314);
xor XOR2 (N2827, N2816, N148);
or OR4 (N2828, N2824, N1945, N1902, N344);
xor XOR2 (N2829, N2820, N589);
xor XOR2 (N2830, N2826, N970);
not NOT1 (N2831, N2828);
xor XOR2 (N2832, N2829, N2064);
or OR2 (N2833, N2832, N1740);
nor NOR2 (N2834, N2830, N1125);
and AND4 (N2835, N2825, N406, N391, N839);
xor XOR2 (N2836, N2833, N1900);
or OR3 (N2837, N2807, N1603, N1645);
nor NOR2 (N2838, N2800, N1956);
not NOT1 (N2839, N2811);
not NOT1 (N2840, N2838);
nand NAND2 (N2841, N2836, N546);
buf BUF1 (N2842, N2819);
nor NOR3 (N2843, N2835, N2184, N336);
and AND3 (N2844, N2831, N1261, N1146);
buf BUF1 (N2845, N2842);
buf BUF1 (N2846, N2827);
nand NAND4 (N2847, N2841, N147, N1948, N2027);
or OR4 (N2848, N2845, N1319, N1639, N2308);
xor XOR2 (N2849, N2834, N2009);
nor NOR4 (N2850, N2843, N947, N1322, N429);
nor NOR2 (N2851, N2848, N1571);
nor NOR3 (N2852, N2839, N2214, N2377);
or OR4 (N2853, N2850, N1084, N797, N539);
not NOT1 (N2854, N2844);
xor XOR2 (N2855, N2840, N540);
and AND2 (N2856, N2849, N31);
buf BUF1 (N2857, N2847);
not NOT1 (N2858, N2851);
nor NOR3 (N2859, N2858, N154, N979);
buf BUF1 (N2860, N2846);
buf BUF1 (N2861, N2854);
or OR4 (N2862, N2852, N430, N1038, N68);
and AND4 (N2863, N2837, N207, N1953, N928);
not NOT1 (N2864, N2818);
or OR3 (N2865, N2855, N1077, N666);
xor XOR2 (N2866, N2864, N1607);
buf BUF1 (N2867, N2863);
not NOT1 (N2868, N2867);
nor NOR4 (N2869, N2862, N756, N148, N547);
nand NAND4 (N2870, N2857, N1598, N1675, N469);
xor XOR2 (N2871, N2866, N2282);
buf BUF1 (N2872, N2865);
nand NAND4 (N2873, N2870, N1233, N248, N2237);
xor XOR2 (N2874, N2853, N437);
xor XOR2 (N2875, N2868, N2282);
not NOT1 (N2876, N2859);
nand NAND2 (N2877, N2860, N229);
xor XOR2 (N2878, N2871, N840);
not NOT1 (N2879, N2875);
nor NOR3 (N2880, N2856, N146, N423);
nand NAND3 (N2881, N2876, N507, N1959);
xor XOR2 (N2882, N2881, N1147);
nand NAND4 (N2883, N2861, N1079, N2750, N848);
nand NAND2 (N2884, N2878, N1896);
xor XOR2 (N2885, N2874, N501);
and AND3 (N2886, N2885, N1481, N2462);
buf BUF1 (N2887, N2880);
nand NAND4 (N2888, N2869, N1530, N1969, N1931);
buf BUF1 (N2889, N2886);
nand NAND4 (N2890, N2873, N2813, N720, N2165);
or OR3 (N2891, N2882, N2142, N2811);
buf BUF1 (N2892, N2890);
nand NAND3 (N2893, N2889, N1467, N31);
buf BUF1 (N2894, N2892);
xor XOR2 (N2895, N2891, N2170);
or OR3 (N2896, N2887, N1135, N825);
xor XOR2 (N2897, N2895, N1344);
xor XOR2 (N2898, N2893, N1901);
not NOT1 (N2899, N2884);
buf BUF1 (N2900, N2872);
or OR3 (N2901, N2879, N458, N430);
buf BUF1 (N2902, N2898);
or OR3 (N2903, N2877, N706, N1743);
not NOT1 (N2904, N2899);
and AND4 (N2905, N2897, N932, N39, N2837);
or OR2 (N2906, N2905, N1678);
buf BUF1 (N2907, N2901);
buf BUF1 (N2908, N2903);
xor XOR2 (N2909, N2908, N2167);
not NOT1 (N2910, N2909);
not NOT1 (N2911, N2904);
xor XOR2 (N2912, N2907, N286);
or OR2 (N2913, N2900, N198);
buf BUF1 (N2914, N2910);
nand NAND4 (N2915, N2902, N370, N1894, N346);
buf BUF1 (N2916, N2914);
nor NOR2 (N2917, N2888, N2);
or OR2 (N2918, N2913, N1657);
nor NOR2 (N2919, N2917, N1940);
nand NAND2 (N2920, N2916, N115);
not NOT1 (N2921, N2918);
and AND3 (N2922, N2906, N415, N1812);
nor NOR2 (N2923, N2915, N1698);
not NOT1 (N2924, N2894);
nor NOR3 (N2925, N2920, N2912, N2825);
nor NOR4 (N2926, N1892, N2359, N1263, N621);
xor XOR2 (N2927, N2896, N916);
nor NOR4 (N2928, N2911, N747, N368, N162);
nor NOR4 (N2929, N2919, N1769, N2676, N227);
nand NAND2 (N2930, N2925, N2552);
not NOT1 (N2931, N2926);
xor XOR2 (N2932, N2931, N825);
nor NOR2 (N2933, N2932, N2076);
and AND2 (N2934, N2933, N296);
buf BUF1 (N2935, N2934);
buf BUF1 (N2936, N2927);
nor NOR3 (N2937, N2936, N2698, N2210);
and AND4 (N2938, N2935, N1816, N2843, N779);
xor XOR2 (N2939, N2923, N2083);
xor XOR2 (N2940, N2924, N322);
nand NAND2 (N2941, N2938, N1275);
nand NAND4 (N2942, N2883, N1748, N2494, N591);
buf BUF1 (N2943, N2940);
or OR4 (N2944, N2941, N186, N2782, N847);
buf BUF1 (N2945, N2944);
or OR4 (N2946, N2929, N2933, N1075, N2134);
xor XOR2 (N2947, N2939, N804);
not NOT1 (N2948, N2942);
buf BUF1 (N2949, N2921);
nand NAND4 (N2950, N2949, N970, N2239, N221);
nand NAND2 (N2951, N2945, N2237);
buf BUF1 (N2952, N2930);
nor NOR3 (N2953, N2952, N2100, N710);
buf BUF1 (N2954, N2946);
xor XOR2 (N2955, N2954, N770);
and AND2 (N2956, N2948, N9);
buf BUF1 (N2957, N2950);
xor XOR2 (N2958, N2956, N624);
or OR2 (N2959, N2953, N2104);
xor XOR2 (N2960, N2928, N2018);
nor NOR4 (N2961, N2959, N802, N1854, N527);
nand NAND3 (N2962, N2958, N820, N2772);
xor XOR2 (N2963, N2955, N1111);
buf BUF1 (N2964, N2947);
nand NAND2 (N2965, N2957, N2584);
nor NOR4 (N2966, N2963, N2410, N1040, N301);
nor NOR3 (N2967, N2966, N1230, N1645);
or OR3 (N2968, N2965, N2237, N1192);
buf BUF1 (N2969, N2962);
nor NOR2 (N2970, N2969, N1996);
buf BUF1 (N2971, N2951);
nand NAND3 (N2972, N2960, N1047, N1810);
nand NAND4 (N2973, N2972, N1306, N190, N1029);
xor XOR2 (N2974, N2943, N2436);
nor NOR4 (N2975, N2968, N506, N2699, N2917);
nor NOR4 (N2976, N2973, N2864, N2460, N2043);
buf BUF1 (N2977, N2970);
xor XOR2 (N2978, N2961, N2007);
nand NAND2 (N2979, N2937, N286);
not NOT1 (N2980, N2967);
xor XOR2 (N2981, N2980, N2841);
nand NAND4 (N2982, N2964, N2973, N222, N91);
nor NOR4 (N2983, N2981, N2608, N2050, N368);
or OR2 (N2984, N2979, N2653);
nor NOR2 (N2985, N2971, N1828);
xor XOR2 (N2986, N2975, N587);
buf BUF1 (N2987, N2986);
and AND3 (N2988, N2978, N864, N928);
or OR3 (N2989, N2977, N957, N1086);
not NOT1 (N2990, N2984);
nor NOR3 (N2991, N2983, N1169, N142);
nand NAND4 (N2992, N2991, N530, N1086, N119);
or OR2 (N2993, N2989, N2476);
nand NAND4 (N2994, N2992, N2890, N1914, N1785);
not NOT1 (N2995, N2974);
nor NOR4 (N2996, N2993, N389, N2711, N2759);
not NOT1 (N2997, N2985);
buf BUF1 (N2998, N2994);
buf BUF1 (N2999, N2995);
buf BUF1 (N3000, N2976);
nand NAND3 (N3001, N2982, N1804, N2474);
nor NOR4 (N3002, N3000, N2632, N2820, N561);
nand NAND4 (N3003, N2996, N2102, N2357, N583);
and AND2 (N3004, N2987, N1704);
xor XOR2 (N3005, N2988, N1615);
nor NOR3 (N3006, N2922, N2782, N210);
and AND3 (N3007, N3004, N1819, N2515);
and AND3 (N3008, N3002, N1727, N1932);
or OR2 (N3009, N3008, N2432);
buf BUF1 (N3010, N3007);
nand NAND3 (N3011, N3006, N406, N2446);
not NOT1 (N3012, N3009);
or OR4 (N3013, N2997, N659, N274, N1831);
xor XOR2 (N3014, N3005, N2290);
nand NAND3 (N3015, N3014, N409, N1984);
not NOT1 (N3016, N2999);
or OR4 (N3017, N3001, N993, N222, N2559);
and AND2 (N3018, N3003, N1412);
or OR4 (N3019, N3015, N1397, N1885, N188);
or OR4 (N3020, N3019, N90, N3012, N597);
and AND4 (N3021, N94, N1025, N292, N1749);
buf BUF1 (N3022, N2990);
nand NAND4 (N3023, N3022, N680, N2248, N2155);
and AND3 (N3024, N3016, N2674, N2835);
or OR4 (N3025, N3018, N455, N1489, N1241);
nand NAND4 (N3026, N3025, N2199, N2440, N2662);
xor XOR2 (N3027, N3024, N4);
or OR3 (N3028, N3011, N680, N2129);
or OR2 (N3029, N3020, N632);
nand NAND2 (N3030, N3021, N43);
nand NAND4 (N3031, N3026, N2265, N102, N2774);
nor NOR4 (N3032, N3017, N424, N1638, N2015);
nor NOR4 (N3033, N3027, N1105, N1444, N38);
nand NAND3 (N3034, N3031, N2518, N1625);
nand NAND4 (N3035, N3032, N2726, N1305, N897);
xor XOR2 (N3036, N3028, N296);
xor XOR2 (N3037, N3035, N2745);
or OR3 (N3038, N3013, N2629, N821);
and AND2 (N3039, N3034, N2967);
not NOT1 (N3040, N3037);
xor XOR2 (N3041, N3030, N1305);
nand NAND2 (N3042, N3033, N2534);
nand NAND3 (N3043, N3040, N513, N2952);
nor NOR2 (N3044, N3039, N2067);
or OR3 (N3045, N3042, N2192, N2134);
nor NOR4 (N3046, N2998, N1566, N2467, N2847);
buf BUF1 (N3047, N3010);
and AND4 (N3048, N3045, N2004, N569, N1264);
and AND4 (N3049, N3041, N1644, N19, N2185);
xor XOR2 (N3050, N3046, N1740);
and AND4 (N3051, N3044, N1222, N358, N1935);
xor XOR2 (N3052, N3029, N975);
nor NOR4 (N3053, N3051, N739, N2684, N3022);
not NOT1 (N3054, N3023);
nand NAND4 (N3055, N3050, N40, N119, N231);
buf BUF1 (N3056, N3036);
buf BUF1 (N3057, N3056);
buf BUF1 (N3058, N3043);
nand NAND2 (N3059, N3058, N1272);
nor NOR2 (N3060, N3048, N2392);
nand NAND3 (N3061, N3060, N849, N2095);
and AND3 (N3062, N3054, N182, N786);
and AND3 (N3063, N3061, N2420, N2981);
not NOT1 (N3064, N3053);
nand NAND4 (N3065, N3064, N96, N167, N2926);
nand NAND3 (N3066, N3055, N470, N2466);
nor NOR3 (N3067, N3047, N445, N2568);
not NOT1 (N3068, N3049);
or OR2 (N3069, N3068, N1036);
and AND3 (N3070, N3057, N1703, N339);
buf BUF1 (N3071, N3059);
or OR4 (N3072, N3067, N2381, N605, N1882);
nor NOR4 (N3073, N3070, N2259, N2751, N611);
nand NAND4 (N3074, N3073, N277, N2748, N1653);
not NOT1 (N3075, N3072);
nand NAND4 (N3076, N3075, N405, N2817, N63);
xor XOR2 (N3077, N3052, N1519);
xor XOR2 (N3078, N3074, N297);
not NOT1 (N3079, N3078);
or OR3 (N3080, N3077, N2361, N1799);
xor XOR2 (N3081, N3071, N277);
xor XOR2 (N3082, N3069, N2882);
nand NAND3 (N3083, N3080, N2425, N1372);
buf BUF1 (N3084, N3079);
nor NOR3 (N3085, N3084, N735, N1239);
and AND2 (N3086, N3081, N2152);
not NOT1 (N3087, N3086);
xor XOR2 (N3088, N3062, N809);
nor NOR2 (N3089, N3065, N1056);
not NOT1 (N3090, N3063);
nor NOR2 (N3091, N3087, N1677);
nor NOR3 (N3092, N3083, N889, N1308);
nor NOR3 (N3093, N3066, N2561, N850);
xor XOR2 (N3094, N3076, N2673);
xor XOR2 (N3095, N3093, N1759);
not NOT1 (N3096, N3038);
or OR2 (N3097, N3091, N674);
and AND2 (N3098, N3085, N1952);
buf BUF1 (N3099, N3088);
and AND2 (N3100, N3097, N1853);
or OR3 (N3101, N3082, N633, N1382);
not NOT1 (N3102, N3094);
xor XOR2 (N3103, N3101, N82);
xor XOR2 (N3104, N3089, N563);
and AND4 (N3105, N3096, N2311, N1638, N1576);
xor XOR2 (N3106, N3092, N2643);
buf BUF1 (N3107, N3106);
nand NAND4 (N3108, N3104, N366, N2325, N621);
nand NAND2 (N3109, N3107, N1992);
xor XOR2 (N3110, N3095, N827);
xor XOR2 (N3111, N3102, N187);
buf BUF1 (N3112, N3090);
nand NAND2 (N3113, N3098, N1355);
not NOT1 (N3114, N3109);
buf BUF1 (N3115, N3103);
or OR2 (N3116, N3108, N2372);
buf BUF1 (N3117, N3105);
nor NOR4 (N3118, N3112, N61, N2638, N81);
or OR3 (N3119, N3099, N2823, N2812);
xor XOR2 (N3120, N3119, N1127);
and AND3 (N3121, N3114, N257, N2);
not NOT1 (N3122, N3110);
or OR2 (N3123, N3122, N2071);
not NOT1 (N3124, N3120);
nand NAND4 (N3125, N3123, N517, N2774, N236);
xor XOR2 (N3126, N3118, N12);
not NOT1 (N3127, N3117);
buf BUF1 (N3128, N3113);
not NOT1 (N3129, N3124);
buf BUF1 (N3130, N3126);
nor NOR3 (N3131, N3125, N1389, N1154);
and AND3 (N3132, N3128, N1829, N731);
or OR4 (N3133, N3115, N474, N514, N2938);
not NOT1 (N3134, N3131);
nor NOR4 (N3135, N3134, N2420, N2313, N2674);
xor XOR2 (N3136, N3100, N1864);
or OR4 (N3137, N3111, N393, N430, N1479);
nor NOR4 (N3138, N3136, N1658, N1024, N2563);
nor NOR3 (N3139, N3127, N1842, N2641);
not NOT1 (N3140, N3129);
or OR4 (N3141, N3135, N509, N1940, N1882);
not NOT1 (N3142, N3133);
and AND3 (N3143, N3132, N400, N2227);
nor NOR2 (N3144, N3141, N1511);
or OR4 (N3145, N3139, N70, N799, N2591);
xor XOR2 (N3146, N3143, N479);
or OR2 (N3147, N3121, N2654);
xor XOR2 (N3148, N3130, N695);
buf BUF1 (N3149, N3147);
or OR4 (N3150, N3148, N3004, N1736, N2388);
buf BUF1 (N3151, N3140);
or OR3 (N3152, N3145, N1113, N975);
not NOT1 (N3153, N3144);
not NOT1 (N3154, N3146);
not NOT1 (N3155, N3154);
and AND4 (N3156, N3116, N2886, N1646, N1795);
xor XOR2 (N3157, N3152, N1700);
buf BUF1 (N3158, N3138);
nand NAND2 (N3159, N3149, N770);
nor NOR3 (N3160, N3158, N1253, N82);
buf BUF1 (N3161, N3153);
or OR3 (N3162, N3159, N129, N1678);
not NOT1 (N3163, N3142);
buf BUF1 (N3164, N3162);
not NOT1 (N3165, N3137);
nor NOR4 (N3166, N3151, N534, N1611, N2354);
and AND3 (N3167, N3156, N493, N2091);
nand NAND3 (N3168, N3150, N1996, N2748);
not NOT1 (N3169, N3157);
nand NAND4 (N3170, N3167, N3105, N1480, N1079);
nor NOR4 (N3171, N3161, N1926, N754, N2570);
or OR4 (N3172, N3170, N1162, N146, N2501);
or OR4 (N3173, N3171, N3068, N1517, N989);
not NOT1 (N3174, N3163);
not NOT1 (N3175, N3166);
nand NAND2 (N3176, N3165, N1573);
nand NAND2 (N3177, N3169, N134);
and AND2 (N3178, N3164, N1670);
xor XOR2 (N3179, N3155, N618);
nor NOR2 (N3180, N3173, N1119);
and AND2 (N3181, N3160, N2305);
nand NAND4 (N3182, N3168, N1826, N2650, N2084);
nand NAND2 (N3183, N3174, N2048);
xor XOR2 (N3184, N3179, N198);
or OR3 (N3185, N3176, N573, N678);
or OR3 (N3186, N3172, N1099, N2778);
buf BUF1 (N3187, N3177);
not NOT1 (N3188, N3181);
and AND2 (N3189, N3187, N1814);
not NOT1 (N3190, N3175);
and AND3 (N3191, N3184, N285, N1131);
and AND4 (N3192, N3189, N963, N1191, N2255);
xor XOR2 (N3193, N3185, N2740);
buf BUF1 (N3194, N3188);
and AND4 (N3195, N3178, N2923, N2284, N1360);
or OR3 (N3196, N3193, N1023, N1624);
nor NOR3 (N3197, N3186, N501, N372);
buf BUF1 (N3198, N3197);
xor XOR2 (N3199, N3196, N2357);
nor NOR4 (N3200, N3192, N1469, N682, N1713);
nor NOR3 (N3201, N3191, N1691, N544);
nor NOR4 (N3202, N3183, N1134, N2455, N2117);
nand NAND4 (N3203, N3201, N1127, N2353, N3092);
and AND3 (N3204, N3198, N2643, N636);
xor XOR2 (N3205, N3182, N2715);
xor XOR2 (N3206, N3203, N2708);
nor NOR3 (N3207, N3202, N2301, N212);
and AND3 (N3208, N3200, N2159, N2838);
nand NAND2 (N3209, N3207, N439);
nand NAND3 (N3210, N3194, N1161, N1788);
not NOT1 (N3211, N3205);
not NOT1 (N3212, N3206);
nand NAND2 (N3213, N3211, N2350);
xor XOR2 (N3214, N3180, N1686);
or OR2 (N3215, N3195, N1571);
or OR2 (N3216, N3210, N51);
nand NAND3 (N3217, N3216, N2254, N645);
or OR2 (N3218, N3209, N699);
nand NAND2 (N3219, N3215, N292);
or OR2 (N3220, N3208, N742);
xor XOR2 (N3221, N3214, N2633);
nor NOR4 (N3222, N3190, N1656, N616, N2175);
not NOT1 (N3223, N3212);
xor XOR2 (N3224, N3222, N2724);
not NOT1 (N3225, N3219);
nand NAND3 (N3226, N3224, N2419, N1254);
not NOT1 (N3227, N3217);
not NOT1 (N3228, N3227);
buf BUF1 (N3229, N3213);
nand NAND3 (N3230, N3221, N2557, N1450);
nand NAND2 (N3231, N3223, N1767);
xor XOR2 (N3232, N3225, N2826);
buf BUF1 (N3233, N3204);
or OR4 (N3234, N3231, N720, N102, N124);
nor NOR4 (N3235, N3199, N1610, N1329, N2471);
not NOT1 (N3236, N3228);
and AND3 (N3237, N3232, N1112, N1507);
or OR4 (N3238, N3234, N1905, N1964, N985);
xor XOR2 (N3239, N3235, N1255);
xor XOR2 (N3240, N3238, N3038);
nor NOR2 (N3241, N3237, N1184);
nor NOR4 (N3242, N3241, N1944, N2243, N1297);
nand NAND4 (N3243, N3229, N2950, N966, N986);
nor NOR2 (N3244, N3218, N2482);
nor NOR4 (N3245, N3240, N99, N2537, N2154);
nand NAND2 (N3246, N3220, N3115);
nand NAND3 (N3247, N3246, N143, N456);
nand NAND4 (N3248, N3226, N883, N2848, N418);
nor NOR4 (N3249, N3230, N683, N1371, N2852);
or OR3 (N3250, N3236, N2980, N1060);
not NOT1 (N3251, N3250);
buf BUF1 (N3252, N3233);
xor XOR2 (N3253, N3249, N2601);
buf BUF1 (N3254, N3253);
nand NAND2 (N3255, N3252, N972);
nor NOR4 (N3256, N3239, N1827, N339, N2812);
not NOT1 (N3257, N3245);
buf BUF1 (N3258, N3242);
buf BUF1 (N3259, N3248);
or OR2 (N3260, N3256, N1869);
and AND4 (N3261, N3257, N758, N278, N1967);
not NOT1 (N3262, N3244);
or OR2 (N3263, N3262, N1623);
and AND3 (N3264, N3251, N1437, N2068);
xor XOR2 (N3265, N3247, N2762);
or OR2 (N3266, N3261, N2064);
or OR2 (N3267, N3243, N1278);
nand NAND2 (N3268, N3264, N1488);
not NOT1 (N3269, N3263);
nor NOR4 (N3270, N3259, N2538, N432, N3215);
nor NOR3 (N3271, N3265, N91, N15);
buf BUF1 (N3272, N3267);
not NOT1 (N3273, N3270);
xor XOR2 (N3274, N3269, N1062);
buf BUF1 (N3275, N3268);
and AND3 (N3276, N3271, N2590, N1326);
nor NOR2 (N3277, N3273, N528);
not NOT1 (N3278, N3276);
buf BUF1 (N3279, N3260);
or OR4 (N3280, N3275, N298, N19, N1267);
or OR3 (N3281, N3255, N2238, N392);
not NOT1 (N3282, N3279);
nor NOR2 (N3283, N3277, N3088);
or OR2 (N3284, N3266, N2054);
xor XOR2 (N3285, N3284, N1826);
nor NOR4 (N3286, N3272, N181, N3204, N1227);
not NOT1 (N3287, N3280);
not NOT1 (N3288, N3278);
or OR3 (N3289, N3283, N3234, N2646);
or OR3 (N3290, N3254, N2544, N220);
nand NAND2 (N3291, N3290, N2605);
buf BUF1 (N3292, N3287);
buf BUF1 (N3293, N3292);
or OR2 (N3294, N3282, N1994);
nand NAND2 (N3295, N3286, N2823);
xor XOR2 (N3296, N3281, N2937);
not NOT1 (N3297, N3288);
nand NAND3 (N3298, N3285, N465, N1824);
and AND2 (N3299, N3294, N2770);
nand NAND2 (N3300, N3289, N1037);
or OR2 (N3301, N3258, N699);
or OR2 (N3302, N3291, N3188);
buf BUF1 (N3303, N3298);
not NOT1 (N3304, N3303);
nor NOR3 (N3305, N3302, N136, N2974);
nor NOR4 (N3306, N3296, N433, N1716, N2893);
nor NOR2 (N3307, N3297, N227);
nand NAND3 (N3308, N3300, N2568, N2769);
nor NOR3 (N3309, N3305, N474, N448);
and AND2 (N3310, N3299, N3256);
xor XOR2 (N3311, N3308, N3275);
or OR2 (N3312, N3307, N590);
buf BUF1 (N3313, N3295);
nand NAND3 (N3314, N3301, N2329, N527);
nor NOR4 (N3315, N3274, N1895, N2237, N899);
nand NAND4 (N3316, N3304, N327, N2808, N1204);
or OR2 (N3317, N3313, N2115);
buf BUF1 (N3318, N3309);
xor XOR2 (N3319, N3317, N2602);
nand NAND4 (N3320, N3315, N2665, N433, N325);
nand NAND3 (N3321, N3316, N259, N1453);
nand NAND4 (N3322, N3306, N2404, N3102, N161);
or OR4 (N3323, N3321, N765, N2611, N2215);
nand NAND3 (N3324, N3310, N2489, N135);
buf BUF1 (N3325, N3293);
nand NAND4 (N3326, N3322, N191, N639, N240);
and AND4 (N3327, N3311, N2662, N2952, N585);
nand NAND4 (N3328, N3314, N588, N1790, N904);
or OR2 (N3329, N3318, N204);
nor NOR2 (N3330, N3326, N2534);
xor XOR2 (N3331, N3325, N2077);
or OR3 (N3332, N3331, N562, N3170);
not NOT1 (N3333, N3320);
and AND2 (N3334, N3332, N2360);
and AND3 (N3335, N3328, N442, N892);
nand NAND4 (N3336, N3333, N843, N2687, N2775);
and AND4 (N3337, N3324, N3015, N231, N2866);
xor XOR2 (N3338, N3323, N1429);
nor NOR2 (N3339, N3329, N2734);
not NOT1 (N3340, N3336);
or OR3 (N3341, N3330, N3265, N3012);
and AND3 (N3342, N3335, N1157, N525);
and AND2 (N3343, N3340, N1465);
not NOT1 (N3344, N3341);
nand NAND4 (N3345, N3312, N1254, N2185, N853);
buf BUF1 (N3346, N3344);
buf BUF1 (N3347, N3342);
xor XOR2 (N3348, N3319, N1504);
buf BUF1 (N3349, N3327);
not NOT1 (N3350, N3338);
or OR4 (N3351, N3334, N740, N3318, N2028);
or OR2 (N3352, N3345, N2511);
nand NAND4 (N3353, N3349, N1030, N687, N2052);
not NOT1 (N3354, N3351);
or OR4 (N3355, N3348, N3141, N2320, N3094);
xor XOR2 (N3356, N3353, N1215);
buf BUF1 (N3357, N3354);
not NOT1 (N3358, N3337);
buf BUF1 (N3359, N3352);
and AND3 (N3360, N3358, N3280, N2731);
or OR2 (N3361, N3343, N2044);
nor NOR4 (N3362, N3350, N2112, N1584, N361);
and AND3 (N3363, N3347, N620, N590);
or OR4 (N3364, N3356, N1207, N486, N437);
buf BUF1 (N3365, N3357);
nor NOR4 (N3366, N3361, N255, N1281, N2753);
nand NAND3 (N3367, N3365, N1960, N2508);
or OR4 (N3368, N3367, N1591, N1368, N610);
not NOT1 (N3369, N3366);
not NOT1 (N3370, N3369);
buf BUF1 (N3371, N3370);
not NOT1 (N3372, N3362);
not NOT1 (N3373, N3372);
or OR2 (N3374, N3346, N719);
and AND4 (N3375, N3360, N51, N1256, N1189);
nand NAND2 (N3376, N3339, N1518);
buf BUF1 (N3377, N3359);
or OR2 (N3378, N3373, N1071);
nand NAND4 (N3379, N3371, N20, N832, N2528);
or OR2 (N3380, N3355, N584);
or OR4 (N3381, N3375, N2794, N1341, N2913);
or OR4 (N3382, N3378, N1835, N1185, N1429);
nor NOR3 (N3383, N3381, N1305, N97);
and AND3 (N3384, N3368, N79, N2680);
not NOT1 (N3385, N3380);
or OR3 (N3386, N3377, N73, N2690);
or OR3 (N3387, N3364, N3257, N1984);
not NOT1 (N3388, N3376);
nor NOR3 (N3389, N3386, N2432, N2566);
or OR3 (N3390, N3388, N3250, N2246);
or OR2 (N3391, N3384, N1969);
and AND4 (N3392, N3379, N1484, N2342, N2926);
xor XOR2 (N3393, N3374, N1654);
buf BUF1 (N3394, N3382);
buf BUF1 (N3395, N3390);
nand NAND4 (N3396, N3394, N3145, N2220, N1633);
nand NAND4 (N3397, N3383, N3119, N1966, N2203);
and AND4 (N3398, N3397, N2116, N2344, N2405);
nand NAND4 (N3399, N3387, N542, N1040, N2761);
buf BUF1 (N3400, N3363);
not NOT1 (N3401, N3385);
nor NOR4 (N3402, N3395, N3068, N2214, N2150);
nand NAND4 (N3403, N3393, N321, N1281, N2062);
and AND3 (N3404, N3403, N1644, N3179);
not NOT1 (N3405, N3400);
not NOT1 (N3406, N3402);
not NOT1 (N3407, N3405);
xor XOR2 (N3408, N3389, N2769);
or OR4 (N3409, N3392, N3195, N3266, N3062);
nand NAND2 (N3410, N3404, N3252);
or OR4 (N3411, N3410, N1909, N1353, N1945);
nand NAND2 (N3412, N3391, N891);
xor XOR2 (N3413, N3399, N776);
nor NOR2 (N3414, N3407, N824);
nand NAND3 (N3415, N3401, N1954, N2152);
and AND2 (N3416, N3408, N2266);
not NOT1 (N3417, N3412);
xor XOR2 (N3418, N3416, N2381);
and AND4 (N3419, N3396, N3006, N2229, N2323);
or OR2 (N3420, N3419, N139);
nor NOR3 (N3421, N3409, N26, N2699);
xor XOR2 (N3422, N3411, N873);
not NOT1 (N3423, N3418);
buf BUF1 (N3424, N3414);
nand NAND3 (N3425, N3406, N1489, N818);
and AND3 (N3426, N3415, N1705, N2954);
xor XOR2 (N3427, N3426, N1900);
nand NAND4 (N3428, N3427, N1098, N1209, N102);
nor NOR3 (N3429, N3423, N1961, N3237);
nor NOR2 (N3430, N3413, N3070);
not NOT1 (N3431, N3425);
or OR2 (N3432, N3398, N2100);
buf BUF1 (N3433, N3428);
and AND4 (N3434, N3421, N2125, N422, N3334);
or OR3 (N3435, N3430, N2974, N680);
nand NAND3 (N3436, N3429, N1956, N1199);
and AND4 (N3437, N3424, N2845, N3223, N2336);
buf BUF1 (N3438, N3417);
not NOT1 (N3439, N3420);
not NOT1 (N3440, N3436);
buf BUF1 (N3441, N3440);
not NOT1 (N3442, N3431);
xor XOR2 (N3443, N3422, N2648);
not NOT1 (N3444, N3439);
or OR4 (N3445, N3438, N318, N819, N1650);
not NOT1 (N3446, N3441);
or OR2 (N3447, N3446, N2967);
or OR4 (N3448, N3444, N2676, N980, N1933);
not NOT1 (N3449, N3437);
nand NAND2 (N3450, N3449, N874);
nand NAND4 (N3451, N3432, N2038, N402, N54);
buf BUF1 (N3452, N3445);
nand NAND3 (N3453, N3433, N2234, N1083);
nand NAND4 (N3454, N3450, N2834, N1262, N787);
and AND4 (N3455, N3452, N512, N570, N3368);
or OR3 (N3456, N3447, N1322, N29);
nand NAND3 (N3457, N3454, N457, N2020);
and AND3 (N3458, N3435, N83, N617);
nor NOR2 (N3459, N3458, N2639);
nand NAND4 (N3460, N3455, N3391, N2582, N528);
not NOT1 (N3461, N3453);
nand NAND3 (N3462, N3443, N2776, N320);
nor NOR2 (N3463, N3460, N870);
nand NAND4 (N3464, N3448, N1851, N822, N226);
not NOT1 (N3465, N3462);
and AND2 (N3466, N3465, N2629);
or OR2 (N3467, N3459, N2085);
buf BUF1 (N3468, N3457);
nand NAND2 (N3469, N3461, N467);
xor XOR2 (N3470, N3434, N1291);
or OR4 (N3471, N3467, N332, N3276, N1549);
and AND2 (N3472, N3442, N166);
nand NAND2 (N3473, N3456, N1651);
buf BUF1 (N3474, N3471);
and AND4 (N3475, N3466, N2535, N1701, N3265);
nand NAND3 (N3476, N3473, N1152, N1514);
and AND3 (N3477, N3463, N2968, N3136);
nor NOR4 (N3478, N3451, N1071, N127, N1544);
nand NAND4 (N3479, N3468, N480, N851, N1894);
nand NAND2 (N3480, N3477, N273);
nor NOR3 (N3481, N3464, N2042, N3057);
nor NOR3 (N3482, N3475, N619, N2576);
buf BUF1 (N3483, N3474);
buf BUF1 (N3484, N3481);
nand NAND3 (N3485, N3476, N969, N2084);
or OR2 (N3486, N3478, N3037);
buf BUF1 (N3487, N3484);
nand NAND2 (N3488, N3480, N1932);
or OR2 (N3489, N3485, N515);
buf BUF1 (N3490, N3487);
and AND3 (N3491, N3488, N2541, N3031);
xor XOR2 (N3492, N3486, N2244);
not NOT1 (N3493, N3483);
nor NOR3 (N3494, N3479, N2704, N3368);
not NOT1 (N3495, N3472);
buf BUF1 (N3496, N3490);
buf BUF1 (N3497, N3496);
or OR2 (N3498, N3469, N1104);
xor XOR2 (N3499, N3493, N138);
nor NOR2 (N3500, N3482, N858);
or OR3 (N3501, N3497, N1484, N1605);
nand NAND4 (N3502, N3494, N2829, N1631, N1533);
not NOT1 (N3503, N3495);
nor NOR2 (N3504, N3499, N804);
nor NOR4 (N3505, N3492, N1416, N2699, N2117);
nand NAND3 (N3506, N3505, N870, N3224);
or OR3 (N3507, N3470, N3088, N507);
nor NOR2 (N3508, N3501, N175);
not NOT1 (N3509, N3489);
or OR2 (N3510, N3502, N312);
and AND2 (N3511, N3498, N1294);
nand NAND4 (N3512, N3511, N2025, N3183, N2889);
nand NAND3 (N3513, N3500, N3148, N2833);
nor NOR3 (N3514, N3509, N826, N2843);
and AND2 (N3515, N3504, N2027);
not NOT1 (N3516, N3510);
xor XOR2 (N3517, N3507, N284);
buf BUF1 (N3518, N3517);
nand NAND3 (N3519, N3506, N2589, N3362);
not NOT1 (N3520, N3508);
nor NOR3 (N3521, N3520, N1831, N2501);
nor NOR2 (N3522, N3516, N2179);
or OR2 (N3523, N3522, N2209);
nand NAND3 (N3524, N3512, N1104, N2792);
endmodule