// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N1502,N1495,N1510,N1499,N1513,N1506,N1494,N1512,N1509,N1515;

or OR2 (N16, N7, N2);
or OR2 (N17, N8, N8);
xor XOR2 (N18, N1, N8);
xor XOR2 (N19, N11, N10);
nor NOR3 (N20, N14, N10, N6);
not NOT1 (N21, N7);
and AND3 (N22, N8, N11, N21);
nand NAND3 (N23, N3, N15, N2);
not NOT1 (N24, N15);
not NOT1 (N25, N12);
and AND3 (N26, N11, N5, N18);
xor XOR2 (N27, N3, N22);
nor NOR2 (N28, N13, N27);
or OR4 (N29, N21, N5, N5, N19);
nor NOR4 (N30, N25, N21, N24, N24);
and AND3 (N31, N2, N14, N22);
nor NOR4 (N32, N8, N24, N22, N5);
or OR4 (N33, N17, N28, N8, N27);
or OR2 (N34, N6, N31);
and AND4 (N35, N5, N14, N17, N2);
buf BUF1 (N36, N32);
not NOT1 (N37, N34);
nand NAND4 (N38, N23, N2, N32, N32);
not NOT1 (N39, N16);
and AND4 (N40, N37, N17, N19, N28);
or OR4 (N41, N26, N26, N24, N30);
or OR2 (N42, N20, N23);
or OR2 (N43, N20, N9);
or OR3 (N44, N29, N23, N22);
nor NOR3 (N45, N36, N25, N11);
xor XOR2 (N46, N38, N14);
buf BUF1 (N47, N46);
not NOT1 (N48, N43);
nor NOR4 (N49, N44, N7, N43, N10);
xor XOR2 (N50, N47, N32);
or OR3 (N51, N39, N10, N8);
nand NAND2 (N52, N45, N14);
nand NAND4 (N53, N48, N40, N30, N13);
xor XOR2 (N54, N37, N22);
nor NOR2 (N55, N52, N42);
nand NAND2 (N56, N30, N33);
nand NAND3 (N57, N10, N45, N55);
or OR4 (N58, N56, N34, N5, N53);
and AND2 (N59, N17, N50);
or OR3 (N60, N44, N18, N44);
and AND3 (N61, N59, N45, N16);
xor XOR2 (N62, N6, N43);
and AND3 (N63, N54, N26, N16);
nand NAND2 (N64, N61, N37);
or OR2 (N65, N63, N29);
or OR2 (N66, N49, N8);
nand NAND4 (N67, N64, N47, N54, N35);
buf BUF1 (N68, N31);
not NOT1 (N69, N62);
nand NAND4 (N70, N68, N17, N39, N59);
nand NAND3 (N71, N66, N68, N65);
or OR2 (N72, N51, N44);
nand NAND4 (N73, N26, N13, N1, N23);
not NOT1 (N74, N67);
not NOT1 (N75, N74);
and AND2 (N76, N57, N18);
xor XOR2 (N77, N75, N49);
xor XOR2 (N78, N70, N55);
not NOT1 (N79, N69);
buf BUF1 (N80, N58);
and AND3 (N81, N41, N78, N13);
xor XOR2 (N82, N79, N46);
nor NOR2 (N83, N31, N75);
buf BUF1 (N84, N81);
buf BUF1 (N85, N84);
not NOT1 (N86, N76);
nor NOR4 (N87, N83, N61, N79, N15);
nor NOR3 (N88, N87, N61, N60);
not NOT1 (N89, N66);
not NOT1 (N90, N73);
xor XOR2 (N91, N71, N3);
xor XOR2 (N92, N90, N7);
nor NOR3 (N93, N86, N60, N14);
nor NOR4 (N94, N82, N53, N42, N47);
nor NOR4 (N95, N91, N28, N76, N10);
buf BUF1 (N96, N92);
nor NOR4 (N97, N95, N25, N54, N64);
buf BUF1 (N98, N89);
nor NOR3 (N99, N77, N29, N65);
xor XOR2 (N100, N88, N91);
buf BUF1 (N101, N85);
not NOT1 (N102, N97);
buf BUF1 (N103, N99);
buf BUF1 (N104, N98);
xor XOR2 (N105, N72, N16);
nor NOR2 (N106, N104, N79);
nor NOR3 (N107, N100, N60, N1);
buf BUF1 (N108, N106);
nor NOR2 (N109, N102, N59);
or OR4 (N110, N96, N102, N22, N103);
or OR4 (N111, N36, N93, N76, N52);
or OR4 (N112, N111, N77, N73, N40);
and AND2 (N113, N38, N99);
and AND4 (N114, N105, N76, N68, N48);
buf BUF1 (N115, N109);
or OR4 (N116, N94, N4, N104, N67);
or OR3 (N117, N114, N3, N74);
nand NAND4 (N118, N112, N108, N26, N58);
or OR3 (N119, N48, N75, N83);
nand NAND3 (N120, N117, N18, N34);
and AND3 (N121, N120, N62, N101);
or OR4 (N122, N75, N4, N1, N14);
or OR4 (N123, N115, N32, N28, N57);
xor XOR2 (N124, N80, N78);
buf BUF1 (N125, N107);
xor XOR2 (N126, N118, N124);
nand NAND3 (N127, N49, N45, N99);
xor XOR2 (N128, N122, N2);
or OR2 (N129, N110, N116);
nand NAND2 (N130, N10, N35);
and AND3 (N131, N113, N55, N3);
and AND3 (N132, N128, N29, N84);
or OR2 (N133, N129, N21);
and AND4 (N134, N126, N65, N72, N91);
buf BUF1 (N135, N127);
and AND3 (N136, N125, N75, N53);
nand NAND2 (N137, N132, N125);
xor XOR2 (N138, N123, N55);
nand NAND3 (N139, N135, N66, N62);
and AND3 (N140, N137, N34, N125);
xor XOR2 (N141, N139, N117);
or OR2 (N142, N141, N80);
nand NAND2 (N143, N131, N129);
xor XOR2 (N144, N134, N28);
buf BUF1 (N145, N143);
not NOT1 (N146, N138);
or OR4 (N147, N136, N116, N19, N120);
nor NOR4 (N148, N121, N86, N7, N123);
nand NAND2 (N149, N133, N115);
nand NAND2 (N150, N149, N51);
nand NAND3 (N151, N130, N33, N125);
or OR3 (N152, N144, N122, N8);
or OR3 (N153, N150, N27, N52);
xor XOR2 (N154, N145, N114);
buf BUF1 (N155, N140);
xor XOR2 (N156, N153, N5);
or OR3 (N157, N155, N20, N47);
xor XOR2 (N158, N157, N10);
not NOT1 (N159, N151);
or OR3 (N160, N147, N16, N78);
buf BUF1 (N161, N159);
and AND4 (N162, N156, N108, N85, N1);
xor XOR2 (N163, N161, N92);
buf BUF1 (N164, N148);
or OR4 (N165, N119, N106, N123, N127);
nor NOR2 (N166, N152, N133);
nand NAND4 (N167, N165, N65, N110, N4);
xor XOR2 (N168, N146, N27);
nand NAND3 (N169, N162, N70, N33);
or OR2 (N170, N154, N97);
xor XOR2 (N171, N170, N112);
xor XOR2 (N172, N160, N59);
and AND2 (N173, N167, N81);
nor NOR4 (N174, N164, N3, N23, N99);
or OR2 (N175, N158, N22);
and AND3 (N176, N174, N56, N93);
and AND2 (N177, N163, N139);
nor NOR4 (N178, N166, N48, N152, N96);
xor XOR2 (N179, N177, N159);
and AND3 (N180, N179, N95, N34);
nor NOR4 (N181, N169, N126, N46, N43);
and AND2 (N182, N168, N8);
buf BUF1 (N183, N181);
buf BUF1 (N184, N183);
or OR4 (N185, N184, N141, N98, N4);
buf BUF1 (N186, N175);
nand NAND3 (N187, N171, N76, N4);
xor XOR2 (N188, N178, N55);
or OR4 (N189, N187, N50, N132, N149);
xor XOR2 (N190, N185, N108);
not NOT1 (N191, N190);
nor NOR2 (N192, N182, N148);
not NOT1 (N193, N192);
not NOT1 (N194, N186);
xor XOR2 (N195, N176, N103);
nand NAND2 (N196, N189, N107);
not NOT1 (N197, N196);
and AND4 (N198, N188, N20, N38, N118);
not NOT1 (N199, N191);
buf BUF1 (N200, N195);
xor XOR2 (N201, N173, N100);
nor NOR4 (N202, N201, N150, N177, N46);
or OR3 (N203, N197, N123, N169);
nand NAND3 (N204, N142, N112, N42);
or OR2 (N205, N200, N74);
and AND4 (N206, N202, N195, N39, N106);
nand NAND3 (N207, N198, N135, N41);
not NOT1 (N208, N180);
xor XOR2 (N209, N194, N124);
nand NAND4 (N210, N206, N66, N70, N3);
buf BUF1 (N211, N208);
not NOT1 (N212, N205);
xor XOR2 (N213, N212, N84);
xor XOR2 (N214, N207, N90);
and AND3 (N215, N214, N210, N150);
not NOT1 (N216, N193);
xor XOR2 (N217, N209, N108);
nand NAND2 (N218, N199, N169);
not NOT1 (N219, N17);
nand NAND2 (N220, N216, N173);
buf BUF1 (N221, N213);
nand NAND4 (N222, N203, N220, N52, N70);
nor NOR2 (N223, N128, N209);
xor XOR2 (N224, N222, N124);
xor XOR2 (N225, N172, N46);
nand NAND2 (N226, N225, N48);
nand NAND3 (N227, N219, N218, N165);
or OR4 (N228, N5, N26, N200, N189);
nand NAND2 (N229, N226, N42);
not NOT1 (N230, N215);
and AND4 (N231, N229, N43, N45, N171);
or OR3 (N232, N227, N133, N15);
buf BUF1 (N233, N224);
or OR2 (N234, N228, N196);
nor NOR4 (N235, N233, N225, N197, N126);
nand NAND3 (N236, N234, N206, N99);
not NOT1 (N237, N217);
nor NOR4 (N238, N211, N170, N221, N165);
not NOT1 (N239, N97);
buf BUF1 (N240, N239);
or OR4 (N241, N240, N145, N40, N163);
and AND3 (N242, N238, N157, N207);
buf BUF1 (N243, N241);
nor NOR3 (N244, N242, N118, N15);
buf BUF1 (N245, N237);
not NOT1 (N246, N232);
nor NOR4 (N247, N235, N54, N239, N204);
nor NOR4 (N248, N165, N197, N89, N228);
not NOT1 (N249, N247);
xor XOR2 (N250, N223, N206);
buf BUF1 (N251, N244);
and AND4 (N252, N231, N206, N217, N47);
not NOT1 (N253, N243);
or OR4 (N254, N252, N22, N82, N247);
nand NAND3 (N255, N253, N32, N131);
or OR2 (N256, N248, N198);
buf BUF1 (N257, N249);
xor XOR2 (N258, N236, N220);
and AND4 (N259, N256, N51, N76, N172);
nand NAND3 (N260, N250, N144, N108);
and AND2 (N261, N255, N14);
buf BUF1 (N262, N251);
and AND2 (N263, N262, N74);
nor NOR3 (N264, N254, N85, N161);
nor NOR2 (N265, N258, N54);
buf BUF1 (N266, N246);
not NOT1 (N267, N257);
or OR3 (N268, N261, N67, N171);
and AND4 (N269, N267, N152, N16, N258);
not NOT1 (N270, N260);
not NOT1 (N271, N259);
not NOT1 (N272, N245);
and AND2 (N273, N265, N57);
or OR2 (N274, N271, N212);
nand NAND3 (N275, N273, N71, N96);
nand NAND3 (N276, N264, N171, N270);
nor NOR2 (N277, N78, N125);
nand NAND4 (N278, N276, N220, N120, N12);
nor NOR3 (N279, N274, N157, N16);
and AND2 (N280, N279, N129);
buf BUF1 (N281, N263);
nand NAND4 (N282, N266, N125, N104, N119);
not NOT1 (N283, N230);
buf BUF1 (N284, N272);
or OR4 (N285, N283, N91, N226, N236);
nor NOR2 (N286, N277, N157);
xor XOR2 (N287, N284, N224);
nand NAND3 (N288, N286, N13, N150);
not NOT1 (N289, N269);
xor XOR2 (N290, N288, N85);
buf BUF1 (N291, N290);
or OR4 (N292, N291, N257, N17, N258);
or OR3 (N293, N280, N28, N139);
and AND3 (N294, N281, N93, N290);
xor XOR2 (N295, N278, N278);
nand NAND2 (N296, N282, N12);
and AND3 (N297, N295, N62, N246);
or OR3 (N298, N275, N141, N162);
buf BUF1 (N299, N287);
nor NOR4 (N300, N298, N15, N208, N75);
or OR2 (N301, N296, N89);
nor NOR4 (N302, N294, N22, N196, N191);
buf BUF1 (N303, N292);
or OR3 (N304, N300, N31, N102);
xor XOR2 (N305, N268, N70);
nand NAND3 (N306, N302, N42, N47);
nor NOR3 (N307, N306, N200, N232);
nand NAND2 (N308, N293, N128);
not NOT1 (N309, N285);
or OR3 (N310, N297, N273, N302);
xor XOR2 (N311, N299, N87);
nand NAND4 (N312, N311, N150, N12, N194);
or OR3 (N313, N289, N45, N260);
nand NAND2 (N314, N301, N103);
buf BUF1 (N315, N313);
not NOT1 (N316, N310);
nand NAND3 (N317, N303, N103, N212);
buf BUF1 (N318, N312);
not NOT1 (N319, N308);
xor XOR2 (N320, N315, N10);
or OR2 (N321, N314, N186);
and AND3 (N322, N317, N117, N303);
or OR2 (N323, N318, N274);
nor NOR4 (N324, N309, N128, N210, N261);
buf BUF1 (N325, N307);
and AND4 (N326, N321, N322, N91, N162);
not NOT1 (N327, N97);
and AND4 (N328, N327, N266, N252, N190);
or OR2 (N329, N320, N73);
not NOT1 (N330, N319);
or OR2 (N331, N316, N201);
xor XOR2 (N332, N323, N217);
nand NAND3 (N333, N330, N43, N134);
nand NAND3 (N334, N328, N104, N42);
nand NAND2 (N335, N325, N190);
not NOT1 (N336, N304);
or OR2 (N337, N333, N106);
and AND3 (N338, N329, N85, N316);
not NOT1 (N339, N336);
or OR4 (N340, N326, N266, N190, N129);
nand NAND4 (N341, N339, N203, N93, N247);
and AND2 (N342, N341, N38);
buf BUF1 (N343, N338);
nor NOR4 (N344, N331, N242, N156, N212);
xor XOR2 (N345, N332, N61);
or OR3 (N346, N334, N213, N3);
not NOT1 (N347, N340);
nor NOR2 (N348, N335, N152);
buf BUF1 (N349, N344);
or OR4 (N350, N346, N267, N99, N190);
not NOT1 (N351, N345);
xor XOR2 (N352, N351, N108);
not NOT1 (N353, N324);
or OR3 (N354, N349, N29, N127);
buf BUF1 (N355, N354);
or OR4 (N356, N350, N160, N225, N105);
and AND3 (N357, N342, N195, N156);
or OR2 (N358, N356, N268);
buf BUF1 (N359, N353);
buf BUF1 (N360, N359);
nand NAND2 (N361, N348, N339);
and AND2 (N362, N357, N303);
or OR2 (N363, N358, N33);
not NOT1 (N364, N362);
nand NAND4 (N365, N363, N327, N129, N283);
nor NOR4 (N366, N355, N237, N285, N132);
not NOT1 (N367, N343);
or OR3 (N368, N367, N327, N84);
buf BUF1 (N369, N337);
and AND4 (N370, N366, N118, N230, N55);
and AND4 (N371, N364, N316, N167, N58);
or OR2 (N372, N347, N18);
or OR2 (N373, N368, N370);
xor XOR2 (N374, N331, N107);
nand NAND4 (N375, N352, N106, N316, N81);
nor NOR4 (N376, N369, N44, N172, N83);
not NOT1 (N377, N372);
buf BUF1 (N378, N373);
buf BUF1 (N379, N360);
or OR2 (N380, N305, N13);
nor NOR4 (N381, N365, N136, N366, N77);
nand NAND4 (N382, N361, N318, N361, N94);
not NOT1 (N383, N374);
or OR2 (N384, N371, N253);
not NOT1 (N385, N384);
and AND2 (N386, N383, N368);
buf BUF1 (N387, N381);
not NOT1 (N388, N375);
or OR2 (N389, N382, N261);
not NOT1 (N390, N389);
and AND2 (N391, N387, N191);
nand NAND3 (N392, N379, N253, N135);
or OR3 (N393, N386, N315, N64);
nand NAND3 (N394, N388, N324, N9);
xor XOR2 (N395, N380, N81);
xor XOR2 (N396, N376, N46);
or OR4 (N397, N390, N22, N226, N25);
nor NOR4 (N398, N391, N365, N327, N29);
nor NOR3 (N399, N392, N118, N291);
or OR3 (N400, N394, N99, N163);
and AND2 (N401, N396, N387);
nand NAND4 (N402, N393, N138, N372, N219);
or OR3 (N403, N400, N109, N47);
not NOT1 (N404, N385);
or OR2 (N405, N402, N398);
xor XOR2 (N406, N164, N63);
or OR2 (N407, N406, N208);
buf BUF1 (N408, N378);
nor NOR4 (N409, N407, N314, N76, N246);
or OR3 (N410, N403, N333, N12);
xor XOR2 (N411, N397, N274);
nand NAND4 (N412, N377, N162, N184, N318);
and AND4 (N413, N404, N308, N289, N224);
xor XOR2 (N414, N413, N217);
and AND3 (N415, N409, N174, N323);
buf BUF1 (N416, N412);
nand NAND2 (N417, N410, N283);
nor NOR4 (N418, N408, N13, N179, N345);
and AND3 (N419, N414, N316, N252);
buf BUF1 (N420, N405);
buf BUF1 (N421, N411);
buf BUF1 (N422, N421);
nor NOR4 (N423, N415, N244, N314, N196);
buf BUF1 (N424, N395);
nor NOR2 (N425, N420, N11);
and AND2 (N426, N399, N241);
nor NOR2 (N427, N416, N75);
nor NOR4 (N428, N401, N9, N352, N307);
buf BUF1 (N429, N422);
or OR3 (N430, N428, N21, N186);
xor XOR2 (N431, N419, N126);
not NOT1 (N432, N425);
nand NAND2 (N433, N429, N166);
and AND3 (N434, N430, N52, N286);
nor NOR2 (N435, N426, N368);
nand NAND3 (N436, N432, N282, N215);
not NOT1 (N437, N424);
or OR2 (N438, N435, N311);
nand NAND3 (N439, N418, N276, N261);
and AND2 (N440, N431, N359);
buf BUF1 (N441, N438);
xor XOR2 (N442, N439, N217);
and AND4 (N443, N417, N73, N264, N406);
buf BUF1 (N444, N433);
not NOT1 (N445, N444);
nand NAND4 (N446, N427, N86, N315, N314);
buf BUF1 (N447, N441);
nand NAND3 (N448, N442, N159, N137);
not NOT1 (N449, N437);
xor XOR2 (N450, N447, N56);
nor NOR4 (N451, N440, N13, N196, N219);
and AND4 (N452, N445, N278, N136, N382);
not NOT1 (N453, N434);
and AND4 (N454, N451, N314, N112, N221);
xor XOR2 (N455, N448, N307);
or OR4 (N456, N443, N99, N36, N439);
buf BUF1 (N457, N446);
buf BUF1 (N458, N423);
or OR3 (N459, N449, N285, N20);
nor NOR2 (N460, N453, N225);
nand NAND4 (N461, N450, N62, N304, N51);
or OR3 (N462, N460, N234, N329);
not NOT1 (N463, N452);
xor XOR2 (N464, N436, N416);
nand NAND4 (N465, N463, N152, N209, N408);
and AND2 (N466, N464, N377);
buf BUF1 (N467, N459);
or OR3 (N468, N462, N241, N185);
nand NAND3 (N469, N466, N92, N73);
not NOT1 (N470, N467);
nand NAND3 (N471, N470, N177, N85);
buf BUF1 (N472, N455);
or OR3 (N473, N471, N346, N390);
nor NOR2 (N474, N468, N473);
not NOT1 (N475, N306);
and AND3 (N476, N465, N190, N176);
xor XOR2 (N477, N474, N405);
buf BUF1 (N478, N472);
and AND3 (N479, N461, N249, N115);
not NOT1 (N480, N475);
nor NOR2 (N481, N477, N461);
or OR4 (N482, N479, N456, N402, N195);
buf BUF1 (N483, N322);
or OR2 (N484, N481, N43);
nand NAND3 (N485, N458, N393, N372);
or OR2 (N486, N484, N286);
not NOT1 (N487, N469);
buf BUF1 (N488, N485);
buf BUF1 (N489, N486);
or OR2 (N490, N482, N255);
buf BUF1 (N491, N488);
not NOT1 (N492, N490);
and AND4 (N493, N492, N482, N144, N73);
nand NAND2 (N494, N493, N249);
buf BUF1 (N495, N454);
nor NOR4 (N496, N494, N1, N334, N35);
and AND4 (N497, N491, N227, N265, N326);
buf BUF1 (N498, N476);
and AND2 (N499, N496, N109);
buf BUF1 (N500, N499);
nor NOR4 (N501, N480, N255, N401, N324);
not NOT1 (N502, N487);
or OR4 (N503, N457, N209, N393, N365);
nand NAND4 (N504, N500, N344, N44, N374);
nor NOR3 (N505, N504, N77, N134);
buf BUF1 (N506, N498);
nand NAND4 (N507, N503, N245, N220, N128);
xor XOR2 (N508, N489, N478);
not NOT1 (N509, N158);
and AND4 (N510, N505, N155, N402, N178);
or OR3 (N511, N483, N143, N125);
not NOT1 (N512, N511);
xor XOR2 (N513, N501, N260);
nand NAND2 (N514, N506, N239);
not NOT1 (N515, N502);
buf BUF1 (N516, N512);
xor XOR2 (N517, N508, N381);
nand NAND2 (N518, N495, N166);
and AND4 (N519, N514, N160, N75, N496);
xor XOR2 (N520, N509, N230);
xor XOR2 (N521, N518, N406);
nand NAND3 (N522, N515, N234, N477);
not NOT1 (N523, N521);
not NOT1 (N524, N517);
not NOT1 (N525, N497);
buf BUF1 (N526, N520);
nand NAND3 (N527, N526, N340, N49);
or OR3 (N528, N527, N188, N25);
buf BUF1 (N529, N523);
and AND2 (N530, N522, N477);
not NOT1 (N531, N510);
nand NAND3 (N532, N530, N183, N511);
and AND2 (N533, N528, N335);
nand NAND2 (N534, N531, N422);
nor NOR4 (N535, N516, N419, N24, N15);
buf BUF1 (N536, N535);
nand NAND4 (N537, N532, N321, N443, N151);
nand NAND3 (N538, N534, N196, N148);
nand NAND4 (N539, N538, N460, N436, N275);
and AND2 (N540, N507, N445);
xor XOR2 (N541, N533, N63);
xor XOR2 (N542, N539, N432);
or OR2 (N543, N519, N524);
or OR3 (N544, N445, N58, N406);
buf BUF1 (N545, N544);
or OR2 (N546, N525, N309);
nand NAND3 (N547, N536, N98, N175);
not NOT1 (N548, N545);
nand NAND4 (N549, N537, N232, N250, N142);
or OR4 (N550, N543, N270, N358, N324);
and AND4 (N551, N540, N303, N70, N115);
or OR4 (N552, N513, N225, N185, N200);
xor XOR2 (N553, N552, N45);
or OR4 (N554, N546, N207, N100, N218);
and AND2 (N555, N553, N131);
nor NOR2 (N556, N542, N156);
and AND2 (N557, N541, N36);
buf BUF1 (N558, N557);
nand NAND4 (N559, N529, N322, N138, N132);
and AND4 (N560, N550, N249, N431, N476);
nand NAND3 (N561, N548, N305, N418);
buf BUF1 (N562, N555);
xor XOR2 (N563, N554, N523);
nor NOR3 (N564, N551, N412, N316);
xor XOR2 (N565, N561, N82);
not NOT1 (N566, N547);
or OR4 (N567, N563, N211, N512, N379);
not NOT1 (N568, N567);
xor XOR2 (N569, N549, N126);
nor NOR2 (N570, N559, N195);
xor XOR2 (N571, N566, N248);
or OR2 (N572, N568, N195);
not NOT1 (N573, N556);
nor NOR2 (N574, N562, N68);
or OR4 (N575, N565, N266, N9, N133);
buf BUF1 (N576, N560);
buf BUF1 (N577, N576);
buf BUF1 (N578, N574);
and AND3 (N579, N571, N385, N297);
nor NOR2 (N580, N577, N148);
buf BUF1 (N581, N572);
buf BUF1 (N582, N581);
buf BUF1 (N583, N580);
or OR3 (N584, N578, N201, N458);
buf BUF1 (N585, N564);
buf BUF1 (N586, N583);
and AND4 (N587, N569, N424, N191, N462);
buf BUF1 (N588, N587);
buf BUF1 (N589, N586);
nor NOR3 (N590, N585, N379, N104);
not NOT1 (N591, N589);
buf BUF1 (N592, N591);
and AND3 (N593, N573, N533, N479);
not NOT1 (N594, N590);
and AND2 (N595, N582, N77);
not NOT1 (N596, N579);
or OR2 (N597, N584, N263);
nor NOR4 (N598, N558, N488, N498, N329);
nand NAND3 (N599, N595, N429, N434);
or OR4 (N600, N588, N237, N116, N122);
or OR2 (N601, N575, N163);
buf BUF1 (N602, N597);
nand NAND3 (N603, N570, N137, N447);
and AND2 (N604, N603, N224);
nand NAND4 (N605, N601, N342, N491, N248);
not NOT1 (N606, N599);
and AND2 (N607, N598, N77);
and AND4 (N608, N605, N445, N284, N548);
and AND3 (N609, N608, N394, N26);
xor XOR2 (N610, N600, N484);
not NOT1 (N611, N609);
buf BUF1 (N612, N611);
nor NOR3 (N613, N594, N133, N122);
not NOT1 (N614, N592);
and AND2 (N615, N607, N98);
nand NAND3 (N616, N612, N569, N234);
nor NOR3 (N617, N593, N297, N475);
xor XOR2 (N618, N615, N37);
or OR2 (N619, N613, N537);
nor NOR3 (N620, N614, N561, N577);
nand NAND4 (N621, N602, N144, N590, N164);
xor XOR2 (N622, N617, N304);
nor NOR4 (N623, N621, N588, N267, N384);
and AND3 (N624, N610, N568, N266);
xor XOR2 (N625, N606, N94);
nand NAND3 (N626, N622, N456, N17);
xor XOR2 (N627, N623, N38);
buf BUF1 (N628, N604);
nand NAND4 (N629, N627, N55, N608, N580);
nand NAND3 (N630, N629, N584, N141);
or OR4 (N631, N618, N613, N293, N460);
buf BUF1 (N632, N628);
nor NOR3 (N633, N631, N359, N120);
or OR4 (N634, N619, N491, N440, N290);
and AND4 (N635, N620, N483, N513, N474);
buf BUF1 (N636, N616);
xor XOR2 (N637, N636, N308);
or OR3 (N638, N624, N359, N503);
nor NOR3 (N639, N630, N473, N436);
buf BUF1 (N640, N637);
and AND2 (N641, N633, N332);
buf BUF1 (N642, N639);
nor NOR4 (N643, N596, N6, N315, N44);
xor XOR2 (N644, N635, N199);
and AND2 (N645, N642, N2);
nand NAND4 (N646, N645, N553, N290, N228);
nand NAND4 (N647, N646, N201, N90, N361);
or OR3 (N648, N644, N94, N533);
or OR2 (N649, N638, N100);
or OR3 (N650, N625, N533, N600);
nand NAND3 (N651, N641, N463, N488);
buf BUF1 (N652, N640);
nand NAND4 (N653, N652, N371, N92, N602);
nand NAND2 (N654, N647, N58);
buf BUF1 (N655, N649);
not NOT1 (N656, N654);
not NOT1 (N657, N655);
not NOT1 (N658, N656);
xor XOR2 (N659, N658, N650);
buf BUF1 (N660, N402);
not NOT1 (N661, N648);
nor NOR2 (N662, N657, N105);
buf BUF1 (N663, N651);
nand NAND2 (N664, N634, N452);
nand NAND3 (N665, N632, N642, N491);
not NOT1 (N666, N660);
or OR3 (N667, N664, N275, N432);
xor XOR2 (N668, N661, N426);
not NOT1 (N669, N665);
buf BUF1 (N670, N643);
not NOT1 (N671, N653);
nand NAND3 (N672, N671, N386, N46);
and AND4 (N673, N626, N469, N658, N185);
not NOT1 (N674, N672);
xor XOR2 (N675, N666, N68);
nor NOR4 (N676, N662, N571, N512, N485);
buf BUF1 (N677, N668);
not NOT1 (N678, N663);
buf BUF1 (N679, N674);
or OR3 (N680, N677, N470, N122);
nor NOR3 (N681, N676, N261, N573);
buf BUF1 (N682, N675);
and AND3 (N683, N682, N168, N380);
not NOT1 (N684, N659);
and AND4 (N685, N681, N3, N92, N629);
and AND3 (N686, N684, N295, N603);
and AND2 (N687, N673, N449);
not NOT1 (N688, N667);
and AND4 (N689, N680, N394, N227, N562);
buf BUF1 (N690, N685);
not NOT1 (N691, N670);
nor NOR3 (N692, N689, N499, N1);
nor NOR3 (N693, N683, N377, N57);
buf BUF1 (N694, N686);
xor XOR2 (N695, N691, N411);
or OR2 (N696, N695, N665);
xor XOR2 (N697, N679, N451);
nor NOR3 (N698, N692, N249, N78);
xor XOR2 (N699, N693, N499);
xor XOR2 (N700, N696, N269);
buf BUF1 (N701, N687);
nor NOR2 (N702, N697, N351);
not NOT1 (N703, N699);
nand NAND4 (N704, N688, N23, N393, N286);
not NOT1 (N705, N678);
nor NOR3 (N706, N704, N515, N118);
nand NAND3 (N707, N669, N420, N703);
or OR3 (N708, N268, N514, N692);
xor XOR2 (N709, N707, N652);
nand NAND4 (N710, N709, N335, N641, N547);
nand NAND3 (N711, N690, N281, N618);
or OR3 (N712, N705, N428, N534);
buf BUF1 (N713, N711);
buf BUF1 (N714, N700);
and AND4 (N715, N712, N150, N293, N203);
or OR3 (N716, N694, N458, N285);
nor NOR3 (N717, N715, N451, N287);
and AND2 (N718, N706, N447);
or OR3 (N719, N701, N352, N601);
or OR2 (N720, N719, N166);
xor XOR2 (N721, N718, N211);
nand NAND3 (N722, N717, N453, N281);
xor XOR2 (N723, N716, N46);
nor NOR2 (N724, N721, N302);
or OR2 (N725, N714, N123);
not NOT1 (N726, N723);
buf BUF1 (N727, N713);
and AND4 (N728, N720, N511, N200, N182);
nand NAND3 (N729, N725, N223, N141);
xor XOR2 (N730, N729, N279);
or OR4 (N731, N698, N594, N184, N94);
nor NOR4 (N732, N728, N714, N586, N149);
and AND3 (N733, N708, N409, N259);
nand NAND4 (N734, N726, N668, N707, N205);
nor NOR2 (N735, N727, N409);
nor NOR4 (N736, N724, N491, N464, N277);
nand NAND4 (N737, N731, N13, N251, N551);
not NOT1 (N738, N737);
or OR2 (N739, N702, N700);
not NOT1 (N740, N736);
nand NAND2 (N741, N722, N406);
nand NAND4 (N742, N730, N212, N417, N8);
nor NOR2 (N743, N732, N185);
xor XOR2 (N744, N738, N525);
and AND3 (N745, N743, N672, N274);
nor NOR3 (N746, N742, N397, N703);
and AND3 (N747, N734, N453, N50);
not NOT1 (N748, N735);
nand NAND2 (N749, N747, N429);
nor NOR4 (N750, N746, N458, N696, N218);
nor NOR4 (N751, N745, N155, N431, N129);
not NOT1 (N752, N751);
xor XOR2 (N753, N744, N478);
and AND2 (N754, N733, N566);
xor XOR2 (N755, N741, N158);
not NOT1 (N756, N740);
nand NAND4 (N757, N749, N654, N478, N649);
not NOT1 (N758, N756);
nand NAND2 (N759, N748, N715);
nand NAND3 (N760, N753, N720, N696);
xor XOR2 (N761, N755, N494);
buf BUF1 (N762, N757);
xor XOR2 (N763, N761, N752);
nand NAND3 (N764, N218, N662, N337);
buf BUF1 (N765, N754);
or OR3 (N766, N759, N41, N132);
nand NAND2 (N767, N764, N88);
not NOT1 (N768, N766);
or OR3 (N769, N750, N721, N716);
nand NAND4 (N770, N767, N702, N311, N203);
buf BUF1 (N771, N758);
nor NOR2 (N772, N710, N674);
not NOT1 (N773, N769);
xor XOR2 (N774, N772, N720);
or OR3 (N775, N763, N88, N308);
nand NAND4 (N776, N771, N436, N603, N416);
not NOT1 (N777, N770);
not NOT1 (N778, N762);
xor XOR2 (N779, N778, N465);
nand NAND4 (N780, N760, N777, N724, N61);
buf BUF1 (N781, N640);
not NOT1 (N782, N781);
not NOT1 (N783, N780);
or OR3 (N784, N765, N389, N599);
buf BUF1 (N785, N775);
or OR3 (N786, N785, N738, N520);
not NOT1 (N787, N768);
xor XOR2 (N788, N783, N95);
not NOT1 (N789, N774);
nand NAND2 (N790, N782, N605);
not NOT1 (N791, N789);
nand NAND4 (N792, N790, N540, N693, N10);
not NOT1 (N793, N788);
nor NOR2 (N794, N787, N463);
buf BUF1 (N795, N792);
buf BUF1 (N796, N795);
buf BUF1 (N797, N786);
buf BUF1 (N798, N776);
nor NOR2 (N799, N794, N288);
xor XOR2 (N800, N739, N749);
nor NOR2 (N801, N793, N790);
xor XOR2 (N802, N801, N377);
nand NAND4 (N803, N784, N361, N574, N218);
not NOT1 (N804, N797);
not NOT1 (N805, N799);
or OR4 (N806, N798, N298, N144, N499);
nor NOR2 (N807, N802, N112);
not NOT1 (N808, N779);
and AND4 (N809, N773, N673, N465, N302);
not NOT1 (N810, N806);
xor XOR2 (N811, N804, N732);
nor NOR3 (N812, N808, N518, N275);
nand NAND4 (N813, N800, N143, N170, N692);
or OR4 (N814, N812, N326, N284, N44);
or OR2 (N815, N805, N39);
and AND2 (N816, N815, N266);
nor NOR3 (N817, N791, N335, N365);
or OR2 (N818, N814, N98);
or OR2 (N819, N803, N657);
and AND4 (N820, N818, N192, N326, N1);
not NOT1 (N821, N813);
xor XOR2 (N822, N810, N811);
nand NAND3 (N823, N59, N564, N259);
nand NAND2 (N824, N819, N501);
or OR3 (N825, N809, N188, N486);
or OR2 (N826, N816, N746);
and AND4 (N827, N796, N238, N391, N732);
not NOT1 (N828, N820);
nand NAND2 (N829, N821, N503);
buf BUF1 (N830, N824);
and AND3 (N831, N825, N698, N445);
nor NOR2 (N832, N822, N41);
xor XOR2 (N833, N807, N254);
buf BUF1 (N834, N828);
or OR3 (N835, N834, N827, N296);
xor XOR2 (N836, N206, N277);
xor XOR2 (N837, N826, N719);
buf BUF1 (N838, N817);
nor NOR4 (N839, N829, N375, N196, N349);
or OR3 (N840, N833, N798, N530);
xor XOR2 (N841, N837, N358);
nand NAND4 (N842, N841, N253, N250, N202);
xor XOR2 (N843, N835, N520);
or OR2 (N844, N842, N814);
not NOT1 (N845, N839);
nor NOR3 (N846, N823, N396, N196);
xor XOR2 (N847, N838, N155);
and AND2 (N848, N840, N377);
nor NOR3 (N849, N845, N165, N604);
and AND2 (N850, N830, N574);
nand NAND3 (N851, N844, N566, N811);
or OR3 (N852, N847, N447, N726);
and AND2 (N853, N843, N768);
or OR4 (N854, N836, N117, N434, N514);
xor XOR2 (N855, N850, N270);
and AND3 (N856, N849, N801, N292);
xor XOR2 (N857, N832, N627);
xor XOR2 (N858, N857, N657);
nand NAND4 (N859, N852, N688, N441, N234);
nor NOR2 (N860, N858, N720);
xor XOR2 (N861, N859, N206);
buf BUF1 (N862, N851);
and AND3 (N863, N860, N411, N757);
nand NAND2 (N864, N861, N200);
or OR2 (N865, N863, N87);
xor XOR2 (N866, N862, N171);
xor XOR2 (N867, N865, N636);
not NOT1 (N868, N853);
nor NOR4 (N869, N831, N181, N858, N497);
nor NOR3 (N870, N846, N56, N25);
buf BUF1 (N871, N848);
nand NAND3 (N872, N855, N533, N431);
not NOT1 (N873, N872);
nand NAND4 (N874, N869, N239, N620, N329);
xor XOR2 (N875, N870, N609);
xor XOR2 (N876, N871, N248);
and AND4 (N877, N875, N611, N615, N68);
nor NOR2 (N878, N867, N295);
not NOT1 (N879, N874);
xor XOR2 (N880, N868, N810);
nor NOR4 (N881, N879, N801, N181, N290);
and AND4 (N882, N854, N217, N141, N471);
buf BUF1 (N883, N880);
or OR2 (N884, N883, N455);
or OR3 (N885, N864, N346, N623);
nand NAND4 (N886, N876, N845, N95, N106);
nand NAND2 (N887, N884, N776);
nand NAND2 (N888, N885, N663);
buf BUF1 (N889, N873);
xor XOR2 (N890, N877, N642);
and AND3 (N891, N856, N724, N289);
and AND2 (N892, N888, N518);
buf BUF1 (N893, N892);
nor NOR3 (N894, N887, N237, N647);
and AND2 (N895, N882, N713);
nor NOR4 (N896, N894, N86, N779, N288);
nor NOR3 (N897, N866, N36, N50);
xor XOR2 (N898, N878, N282);
and AND2 (N899, N895, N444);
nor NOR2 (N900, N897, N752);
and AND3 (N901, N891, N777, N755);
and AND3 (N902, N890, N579, N478);
or OR4 (N903, N889, N423, N545, N885);
nand NAND3 (N904, N881, N545, N89);
xor XOR2 (N905, N899, N739);
xor XOR2 (N906, N901, N270);
nand NAND2 (N907, N886, N707);
xor XOR2 (N908, N900, N656);
nor NOR4 (N909, N904, N399, N51, N121);
buf BUF1 (N910, N896);
or OR4 (N911, N905, N160, N703, N495);
nor NOR4 (N912, N907, N231, N440, N334);
not NOT1 (N913, N908);
buf BUF1 (N914, N902);
nand NAND2 (N915, N903, N457);
not NOT1 (N916, N893);
nor NOR4 (N917, N911, N410, N534, N862);
and AND2 (N918, N898, N64);
and AND4 (N919, N915, N429, N336, N673);
nand NAND4 (N920, N910, N740, N503, N463);
not NOT1 (N921, N913);
buf BUF1 (N922, N914);
buf BUF1 (N923, N922);
xor XOR2 (N924, N916, N804);
buf BUF1 (N925, N920);
and AND3 (N926, N925, N906, N834);
nand NAND3 (N927, N707, N348, N190);
nand NAND2 (N928, N921, N122);
and AND4 (N929, N928, N850, N555, N878);
nor NOR3 (N930, N927, N352, N380);
not NOT1 (N931, N917);
buf BUF1 (N932, N929);
not NOT1 (N933, N931);
or OR2 (N934, N918, N336);
not NOT1 (N935, N934);
not NOT1 (N936, N933);
nor NOR4 (N937, N930, N575, N700, N308);
and AND3 (N938, N936, N509, N749);
not NOT1 (N939, N919);
nand NAND4 (N940, N926, N855, N115, N679);
nand NAND3 (N941, N937, N879, N879);
buf BUF1 (N942, N941);
xor XOR2 (N943, N923, N43);
nor NOR2 (N944, N942, N398);
buf BUF1 (N945, N939);
nand NAND3 (N946, N924, N156, N199);
buf BUF1 (N947, N912);
not NOT1 (N948, N945);
not NOT1 (N949, N944);
or OR4 (N950, N946, N396, N114, N340);
nor NOR3 (N951, N948, N874, N905);
nand NAND2 (N952, N949, N284);
nand NAND2 (N953, N940, N353);
or OR2 (N954, N953, N380);
or OR3 (N955, N954, N753, N627);
or OR2 (N956, N943, N886);
and AND3 (N957, N955, N574, N89);
and AND4 (N958, N951, N894, N134, N158);
and AND3 (N959, N950, N803, N564);
nand NAND4 (N960, N952, N478, N171, N356);
buf BUF1 (N961, N960);
and AND2 (N962, N958, N735);
xor XOR2 (N963, N959, N447);
and AND2 (N964, N909, N191);
buf BUF1 (N965, N961);
buf BUF1 (N966, N938);
not NOT1 (N967, N957);
xor XOR2 (N968, N947, N686);
buf BUF1 (N969, N932);
nand NAND3 (N970, N935, N924, N749);
nor NOR4 (N971, N962, N95, N558, N262);
not NOT1 (N972, N966);
xor XOR2 (N973, N967, N675);
not NOT1 (N974, N969);
or OR3 (N975, N968, N142, N664);
nor NOR4 (N976, N965, N894, N336, N221);
buf BUF1 (N977, N963);
xor XOR2 (N978, N974, N9);
nand NAND2 (N979, N970, N822);
nand NAND3 (N980, N975, N652, N520);
and AND3 (N981, N964, N63, N799);
nor NOR2 (N982, N980, N941);
and AND3 (N983, N981, N809, N368);
nand NAND3 (N984, N978, N61, N816);
buf BUF1 (N985, N956);
buf BUF1 (N986, N971);
and AND2 (N987, N982, N660);
or OR4 (N988, N985, N577, N758, N174);
nor NOR3 (N989, N979, N136, N611);
not NOT1 (N990, N983);
buf BUF1 (N991, N987);
buf BUF1 (N992, N990);
nor NOR3 (N993, N988, N441, N193);
and AND2 (N994, N991, N349);
and AND2 (N995, N994, N173);
buf BUF1 (N996, N984);
not NOT1 (N997, N996);
and AND3 (N998, N997, N440, N270);
nand NAND3 (N999, N976, N380, N524);
xor XOR2 (N1000, N999, N408);
xor XOR2 (N1001, N986, N945);
not NOT1 (N1002, N989);
nor NOR4 (N1003, N993, N885, N712, N388);
xor XOR2 (N1004, N1002, N930);
nand NAND2 (N1005, N977, N528);
or OR3 (N1006, N992, N343, N909);
and AND3 (N1007, N1001, N724, N587);
nand NAND2 (N1008, N998, N352);
and AND3 (N1009, N1008, N481, N567);
nand NAND3 (N1010, N1005, N77, N565);
buf BUF1 (N1011, N995);
xor XOR2 (N1012, N1010, N764);
and AND2 (N1013, N973, N288);
or OR4 (N1014, N1004, N631, N778, N981);
nand NAND4 (N1015, N1000, N178, N288, N981);
nor NOR3 (N1016, N1015, N234, N689);
xor XOR2 (N1017, N1009, N374);
buf BUF1 (N1018, N1011);
nor NOR4 (N1019, N1018, N3, N684, N69);
buf BUF1 (N1020, N1017);
not NOT1 (N1021, N1006);
buf BUF1 (N1022, N1003);
xor XOR2 (N1023, N1014, N295);
xor XOR2 (N1024, N1023, N960);
buf BUF1 (N1025, N1007);
or OR2 (N1026, N1021, N282);
not NOT1 (N1027, N1012);
nor NOR2 (N1028, N1019, N440);
or OR3 (N1029, N972, N884, N664);
nor NOR3 (N1030, N1025, N946, N40);
xor XOR2 (N1031, N1022, N612);
buf BUF1 (N1032, N1024);
or OR2 (N1033, N1026, N593);
not NOT1 (N1034, N1029);
and AND3 (N1035, N1033, N974, N822);
and AND3 (N1036, N1034, N532, N681);
or OR3 (N1037, N1030, N355, N544);
nand NAND4 (N1038, N1028, N347, N404, N237);
or OR4 (N1039, N1037, N1021, N434, N270);
buf BUF1 (N1040, N1032);
and AND2 (N1041, N1038, N517);
buf BUF1 (N1042, N1035);
nand NAND3 (N1043, N1041, N637, N939);
nand NAND4 (N1044, N1020, N813, N437, N856);
buf BUF1 (N1045, N1039);
nor NOR2 (N1046, N1043, N681);
or OR4 (N1047, N1013, N455, N509, N351);
not NOT1 (N1048, N1042);
nand NAND3 (N1049, N1048, N573, N212);
xor XOR2 (N1050, N1016, N314);
nor NOR4 (N1051, N1045, N864, N905, N90);
xor XOR2 (N1052, N1031, N424);
or OR3 (N1053, N1049, N361, N652);
xor XOR2 (N1054, N1052, N1024);
not NOT1 (N1055, N1036);
nand NAND2 (N1056, N1027, N960);
buf BUF1 (N1057, N1056);
or OR3 (N1058, N1057, N11, N1037);
nand NAND4 (N1059, N1055, N580, N750, N895);
or OR2 (N1060, N1054, N220);
xor XOR2 (N1061, N1060, N700);
or OR2 (N1062, N1051, N336);
or OR2 (N1063, N1046, N292);
or OR2 (N1064, N1061, N167);
and AND3 (N1065, N1062, N252, N858);
nor NOR4 (N1066, N1040, N570, N664, N606);
or OR2 (N1067, N1058, N79);
nand NAND3 (N1068, N1053, N626, N789);
xor XOR2 (N1069, N1068, N812);
or OR2 (N1070, N1063, N998);
buf BUF1 (N1071, N1069);
or OR2 (N1072, N1067, N884);
or OR2 (N1073, N1044, N269);
or OR2 (N1074, N1071, N1031);
or OR2 (N1075, N1074, N60);
nand NAND3 (N1076, N1072, N840, N218);
buf BUF1 (N1077, N1073);
and AND3 (N1078, N1047, N522, N550);
xor XOR2 (N1079, N1075, N25);
nor NOR2 (N1080, N1059, N568);
nor NOR2 (N1081, N1080, N1078);
nor NOR4 (N1082, N606, N308, N804, N632);
not NOT1 (N1083, N1064);
buf BUF1 (N1084, N1081);
nor NOR4 (N1085, N1083, N348, N1062, N115);
nand NAND2 (N1086, N1085, N13);
xor XOR2 (N1087, N1086, N802);
or OR3 (N1088, N1084, N942, N224);
xor XOR2 (N1089, N1077, N713);
or OR3 (N1090, N1050, N798, N1011);
not NOT1 (N1091, N1088);
xor XOR2 (N1092, N1070, N247);
nand NAND4 (N1093, N1076, N78, N716, N85);
and AND2 (N1094, N1091, N382);
not NOT1 (N1095, N1094);
not NOT1 (N1096, N1082);
buf BUF1 (N1097, N1065);
nor NOR4 (N1098, N1093, N254, N197, N630);
xor XOR2 (N1099, N1089, N796);
not NOT1 (N1100, N1090);
nand NAND4 (N1101, N1087, N738, N471, N170);
xor XOR2 (N1102, N1099, N1017);
buf BUF1 (N1103, N1102);
buf BUF1 (N1104, N1100);
nor NOR2 (N1105, N1079, N9);
and AND2 (N1106, N1095, N531);
nor NOR4 (N1107, N1104, N1061, N673, N210);
xor XOR2 (N1108, N1107, N531);
buf BUF1 (N1109, N1103);
nand NAND3 (N1110, N1101, N327, N739);
buf BUF1 (N1111, N1108);
nor NOR4 (N1112, N1106, N821, N423, N1051);
not NOT1 (N1113, N1109);
nor NOR4 (N1114, N1097, N881, N288, N1096);
not NOT1 (N1115, N1038);
xor XOR2 (N1116, N1114, N938);
and AND4 (N1117, N1110, N721, N861, N120);
nand NAND2 (N1118, N1112, N432);
nand NAND4 (N1119, N1098, N418, N521, N512);
xor XOR2 (N1120, N1105, N187);
xor XOR2 (N1121, N1111, N840);
nand NAND2 (N1122, N1118, N1000);
and AND3 (N1123, N1122, N718, N687);
buf BUF1 (N1124, N1119);
xor XOR2 (N1125, N1124, N614);
xor XOR2 (N1126, N1120, N773);
nor NOR2 (N1127, N1113, N43);
nor NOR3 (N1128, N1127, N970, N519);
and AND4 (N1129, N1128, N1092, N663, N326);
buf BUF1 (N1130, N950);
or OR3 (N1131, N1066, N158, N785);
or OR4 (N1132, N1115, N754, N51, N721);
not NOT1 (N1133, N1125);
xor XOR2 (N1134, N1121, N715);
buf BUF1 (N1135, N1123);
and AND2 (N1136, N1132, N172);
or OR4 (N1137, N1126, N179, N954, N843);
nor NOR4 (N1138, N1116, N431, N482, N235);
and AND2 (N1139, N1135, N773);
not NOT1 (N1140, N1137);
not NOT1 (N1141, N1130);
buf BUF1 (N1142, N1129);
not NOT1 (N1143, N1142);
and AND4 (N1144, N1140, N1004, N667, N519);
nand NAND4 (N1145, N1144, N775, N138, N337);
or OR3 (N1146, N1138, N732, N1001);
nand NAND3 (N1147, N1136, N749, N507);
not NOT1 (N1148, N1146);
nand NAND4 (N1149, N1147, N796, N693, N344);
buf BUF1 (N1150, N1117);
not NOT1 (N1151, N1133);
nand NAND4 (N1152, N1139, N72, N1115, N707);
and AND2 (N1153, N1145, N569);
nor NOR2 (N1154, N1150, N660);
and AND3 (N1155, N1143, N790, N629);
nand NAND3 (N1156, N1151, N759, N961);
nor NOR4 (N1157, N1149, N1072, N854, N926);
not NOT1 (N1158, N1153);
buf BUF1 (N1159, N1141);
xor XOR2 (N1160, N1134, N682);
xor XOR2 (N1161, N1160, N620);
and AND3 (N1162, N1152, N471, N21);
and AND2 (N1163, N1162, N1119);
xor XOR2 (N1164, N1161, N591);
and AND3 (N1165, N1158, N99, N500);
or OR3 (N1166, N1164, N417, N483);
not NOT1 (N1167, N1148);
and AND4 (N1168, N1157, N639, N257, N467);
and AND4 (N1169, N1154, N1086, N850, N1058);
buf BUF1 (N1170, N1159);
nand NAND4 (N1171, N1167, N247, N195, N1049);
not NOT1 (N1172, N1155);
nand NAND2 (N1173, N1170, N737);
and AND2 (N1174, N1172, N994);
nand NAND4 (N1175, N1173, N39, N257, N102);
nor NOR2 (N1176, N1163, N24);
nor NOR3 (N1177, N1174, N150, N613);
and AND2 (N1178, N1171, N466);
or OR3 (N1179, N1166, N674, N231);
or OR4 (N1180, N1177, N776, N524, N942);
or OR3 (N1181, N1175, N318, N82);
nand NAND3 (N1182, N1169, N123, N1067);
xor XOR2 (N1183, N1179, N36);
buf BUF1 (N1184, N1176);
nand NAND2 (N1185, N1165, N33);
or OR4 (N1186, N1180, N455, N301, N365);
and AND4 (N1187, N1185, N402, N623, N192);
nor NOR4 (N1188, N1183, N1114, N442, N1148);
and AND3 (N1189, N1156, N937, N394);
nand NAND3 (N1190, N1181, N1071, N1182);
and AND4 (N1191, N324, N78, N1051, N541);
and AND3 (N1192, N1131, N15, N173);
and AND2 (N1193, N1184, N597);
buf BUF1 (N1194, N1187);
and AND3 (N1195, N1168, N1190, N400);
or OR4 (N1196, N1138, N164, N1188, N419);
and AND4 (N1197, N133, N519, N836, N60);
buf BUF1 (N1198, N1195);
and AND3 (N1199, N1192, N1027, N526);
xor XOR2 (N1200, N1178, N841);
buf BUF1 (N1201, N1191);
buf BUF1 (N1202, N1194);
buf BUF1 (N1203, N1196);
nor NOR3 (N1204, N1199, N1168, N529);
or OR3 (N1205, N1204, N1024, N748);
nand NAND2 (N1206, N1198, N137);
buf BUF1 (N1207, N1193);
not NOT1 (N1208, N1203);
nand NAND3 (N1209, N1207, N635, N836);
nand NAND2 (N1210, N1189, N1108);
not NOT1 (N1211, N1210);
nor NOR4 (N1212, N1186, N1207, N368, N83);
xor XOR2 (N1213, N1202, N869);
not NOT1 (N1214, N1213);
nor NOR2 (N1215, N1201, N14);
nand NAND2 (N1216, N1215, N239);
and AND3 (N1217, N1216, N901, N44);
xor XOR2 (N1218, N1197, N606);
not NOT1 (N1219, N1217);
and AND3 (N1220, N1200, N1022, N508);
nand NAND2 (N1221, N1218, N582);
or OR2 (N1222, N1220, N1055);
not NOT1 (N1223, N1211);
nor NOR4 (N1224, N1209, N761, N395, N6);
and AND3 (N1225, N1208, N271, N1087);
and AND2 (N1226, N1212, N532);
not NOT1 (N1227, N1224);
nand NAND2 (N1228, N1205, N732);
nand NAND4 (N1229, N1222, N754, N420, N584);
not NOT1 (N1230, N1229);
nand NAND4 (N1231, N1206, N108, N1131, N74);
or OR4 (N1232, N1228, N479, N46, N523);
and AND4 (N1233, N1221, N900, N651, N864);
buf BUF1 (N1234, N1232);
not NOT1 (N1235, N1219);
xor XOR2 (N1236, N1233, N1012);
or OR2 (N1237, N1235, N172);
or OR4 (N1238, N1214, N761, N199, N824);
not NOT1 (N1239, N1236);
nor NOR2 (N1240, N1237, N677);
nor NOR2 (N1241, N1227, N941);
and AND3 (N1242, N1239, N685, N77);
xor XOR2 (N1243, N1234, N661);
or OR2 (N1244, N1243, N61);
nor NOR2 (N1245, N1241, N952);
buf BUF1 (N1246, N1226);
or OR2 (N1247, N1245, N101);
not NOT1 (N1248, N1238);
buf BUF1 (N1249, N1247);
not NOT1 (N1250, N1248);
and AND2 (N1251, N1242, N829);
nand NAND2 (N1252, N1249, N557);
and AND2 (N1253, N1244, N242);
and AND2 (N1254, N1225, N433);
buf BUF1 (N1255, N1251);
nand NAND2 (N1256, N1254, N373);
nand NAND2 (N1257, N1240, N1237);
nor NOR4 (N1258, N1253, N757, N258, N559);
xor XOR2 (N1259, N1246, N1226);
xor XOR2 (N1260, N1257, N76);
nand NAND3 (N1261, N1223, N409, N862);
nor NOR2 (N1262, N1250, N131);
nor NOR4 (N1263, N1260, N564, N753, N302);
nand NAND4 (N1264, N1263, N737, N1060, N758);
xor XOR2 (N1265, N1256, N134);
not NOT1 (N1266, N1262);
nand NAND2 (N1267, N1259, N117);
not NOT1 (N1268, N1258);
or OR3 (N1269, N1267, N349, N367);
not NOT1 (N1270, N1261);
xor XOR2 (N1271, N1268, N974);
or OR3 (N1272, N1266, N167, N1001);
buf BUF1 (N1273, N1252);
buf BUF1 (N1274, N1270);
or OR4 (N1275, N1269, N508, N47, N744);
or OR3 (N1276, N1272, N752, N869);
and AND3 (N1277, N1255, N352, N158);
not NOT1 (N1278, N1230);
xor XOR2 (N1279, N1271, N10);
xor XOR2 (N1280, N1264, N693);
or OR3 (N1281, N1279, N220, N807);
or OR2 (N1282, N1276, N739);
or OR4 (N1283, N1278, N1227, N959, N905);
xor XOR2 (N1284, N1280, N718);
not NOT1 (N1285, N1284);
or OR2 (N1286, N1285, N1239);
buf BUF1 (N1287, N1281);
nor NOR3 (N1288, N1275, N578, N312);
not NOT1 (N1289, N1265);
nor NOR2 (N1290, N1274, N372);
and AND4 (N1291, N1288, N443, N1203, N596);
buf BUF1 (N1292, N1286);
not NOT1 (N1293, N1282);
buf BUF1 (N1294, N1283);
xor XOR2 (N1295, N1289, N15);
nor NOR2 (N1296, N1293, N1008);
and AND4 (N1297, N1231, N93, N517, N71);
or OR4 (N1298, N1297, N610, N790, N686);
nor NOR2 (N1299, N1277, N1156);
buf BUF1 (N1300, N1292);
not NOT1 (N1301, N1273);
nor NOR4 (N1302, N1295, N1273, N1151, N1178);
nor NOR2 (N1303, N1291, N832);
and AND3 (N1304, N1298, N1224, N1140);
xor XOR2 (N1305, N1304, N487);
xor XOR2 (N1306, N1303, N430);
or OR2 (N1307, N1290, N155);
not NOT1 (N1308, N1296);
buf BUF1 (N1309, N1302);
nand NAND4 (N1310, N1306, N158, N10, N807);
nor NOR2 (N1311, N1301, N794);
xor XOR2 (N1312, N1308, N1212);
buf BUF1 (N1313, N1294);
buf BUF1 (N1314, N1311);
not NOT1 (N1315, N1305);
not NOT1 (N1316, N1309);
buf BUF1 (N1317, N1300);
nor NOR4 (N1318, N1314, N803, N1215, N202);
or OR4 (N1319, N1318, N649, N153, N275);
nor NOR4 (N1320, N1287, N1128, N538, N80);
and AND4 (N1321, N1299, N607, N714, N769);
nand NAND4 (N1322, N1321, N1048, N630, N290);
xor XOR2 (N1323, N1317, N5);
buf BUF1 (N1324, N1310);
xor XOR2 (N1325, N1324, N1175);
buf BUF1 (N1326, N1307);
or OR2 (N1327, N1316, N895);
not NOT1 (N1328, N1327);
buf BUF1 (N1329, N1322);
nand NAND3 (N1330, N1326, N17, N1326);
buf BUF1 (N1331, N1312);
nand NAND3 (N1332, N1319, N508, N1112);
not NOT1 (N1333, N1323);
xor XOR2 (N1334, N1315, N1159);
nor NOR2 (N1335, N1333, N527);
nand NAND4 (N1336, N1328, N869, N415, N443);
xor XOR2 (N1337, N1335, N1095);
nand NAND2 (N1338, N1337, N110);
not NOT1 (N1339, N1338);
nand NAND3 (N1340, N1334, N556, N1200);
nand NAND2 (N1341, N1332, N1009);
xor XOR2 (N1342, N1340, N789);
nand NAND4 (N1343, N1336, N66, N638, N1058);
xor XOR2 (N1344, N1329, N834);
nor NOR2 (N1345, N1344, N396);
not NOT1 (N1346, N1320);
buf BUF1 (N1347, N1345);
or OR2 (N1348, N1343, N613);
nor NOR2 (N1349, N1313, N1152);
xor XOR2 (N1350, N1325, N703);
not NOT1 (N1351, N1350);
nand NAND4 (N1352, N1351, N1295, N853, N823);
nand NAND2 (N1353, N1352, N859);
nor NOR3 (N1354, N1341, N987, N519);
and AND3 (N1355, N1330, N717, N1052);
buf BUF1 (N1356, N1331);
nand NAND3 (N1357, N1346, N212, N646);
buf BUF1 (N1358, N1348);
or OR4 (N1359, N1347, N289, N769, N255);
xor XOR2 (N1360, N1354, N196);
nand NAND2 (N1361, N1355, N403);
not NOT1 (N1362, N1359);
not NOT1 (N1363, N1349);
xor XOR2 (N1364, N1363, N1292);
xor XOR2 (N1365, N1361, N432);
and AND2 (N1366, N1339, N642);
not NOT1 (N1367, N1360);
buf BUF1 (N1368, N1358);
xor XOR2 (N1369, N1365, N388);
buf BUF1 (N1370, N1362);
and AND3 (N1371, N1370, N450, N861);
nand NAND2 (N1372, N1364, N1203);
or OR4 (N1373, N1357, N25, N1118, N889);
xor XOR2 (N1374, N1373, N978);
not NOT1 (N1375, N1342);
nor NOR3 (N1376, N1366, N1130, N350);
buf BUF1 (N1377, N1353);
or OR2 (N1378, N1372, N477);
and AND2 (N1379, N1369, N786);
nor NOR3 (N1380, N1378, N1240, N786);
buf BUF1 (N1381, N1368);
not NOT1 (N1382, N1367);
buf BUF1 (N1383, N1382);
buf BUF1 (N1384, N1377);
nand NAND4 (N1385, N1376, N225, N36, N1320);
and AND2 (N1386, N1384, N1155);
and AND4 (N1387, N1356, N1182, N802, N960);
and AND3 (N1388, N1387, N1111, N150);
buf BUF1 (N1389, N1380);
nor NOR4 (N1390, N1374, N934, N1173, N1334);
xor XOR2 (N1391, N1381, N711);
buf BUF1 (N1392, N1371);
nor NOR2 (N1393, N1392, N1325);
nor NOR2 (N1394, N1391, N30);
not NOT1 (N1395, N1394);
and AND3 (N1396, N1395, N185, N604);
or OR2 (N1397, N1386, N234);
nand NAND2 (N1398, N1388, N1245);
not NOT1 (N1399, N1398);
not NOT1 (N1400, N1379);
buf BUF1 (N1401, N1393);
and AND2 (N1402, N1375, N389);
nor NOR3 (N1403, N1397, N1358, N1004);
and AND3 (N1404, N1401, N52, N344);
and AND3 (N1405, N1403, N911, N600);
xor XOR2 (N1406, N1396, N829);
not NOT1 (N1407, N1405);
or OR4 (N1408, N1407, N386, N654, N808);
nand NAND3 (N1409, N1402, N170, N1397);
xor XOR2 (N1410, N1406, N1330);
xor XOR2 (N1411, N1404, N714);
or OR3 (N1412, N1385, N217, N1086);
and AND2 (N1413, N1410, N72);
buf BUF1 (N1414, N1412);
and AND2 (N1415, N1414, N868);
or OR3 (N1416, N1411, N1036, N50);
not NOT1 (N1417, N1415);
or OR2 (N1418, N1400, N1350);
buf BUF1 (N1419, N1416);
and AND2 (N1420, N1413, N1346);
nand NAND3 (N1421, N1409, N273, N86);
not NOT1 (N1422, N1420);
nor NOR3 (N1423, N1422, N271, N919);
xor XOR2 (N1424, N1390, N913);
or OR4 (N1425, N1419, N274, N1222, N284);
xor XOR2 (N1426, N1424, N55);
not NOT1 (N1427, N1399);
nor NOR3 (N1428, N1418, N695, N1063);
or OR2 (N1429, N1426, N285);
not NOT1 (N1430, N1383);
nand NAND2 (N1431, N1417, N1404);
not NOT1 (N1432, N1421);
buf BUF1 (N1433, N1430);
not NOT1 (N1434, N1425);
buf BUF1 (N1435, N1428);
buf BUF1 (N1436, N1408);
nand NAND2 (N1437, N1389, N144);
not NOT1 (N1438, N1433);
not NOT1 (N1439, N1436);
buf BUF1 (N1440, N1429);
not NOT1 (N1441, N1435);
and AND4 (N1442, N1431, N648, N1176, N752);
nand NAND3 (N1443, N1439, N442, N501);
xor XOR2 (N1444, N1434, N211);
buf BUF1 (N1445, N1438);
nor NOR4 (N1446, N1442, N108, N118, N366);
nand NAND3 (N1447, N1427, N16, N413);
buf BUF1 (N1448, N1446);
nand NAND4 (N1449, N1447, N836, N750, N404);
nand NAND4 (N1450, N1449, N515, N323, N799);
nor NOR3 (N1451, N1437, N594, N1019);
buf BUF1 (N1452, N1440);
nor NOR3 (N1453, N1444, N1022, N509);
nor NOR3 (N1454, N1451, N14, N1276);
or OR4 (N1455, N1432, N240, N496, N1015);
or OR4 (N1456, N1452, N738, N1360, N1307);
buf BUF1 (N1457, N1453);
xor XOR2 (N1458, N1445, N1308);
or OR3 (N1459, N1457, N891, N1151);
nor NOR3 (N1460, N1458, N806, N532);
buf BUF1 (N1461, N1456);
xor XOR2 (N1462, N1459, N268);
buf BUF1 (N1463, N1443);
and AND2 (N1464, N1448, N378);
or OR4 (N1465, N1423, N207, N551, N1053);
or OR4 (N1466, N1465, N1152, N408, N253);
nand NAND4 (N1467, N1454, N1075, N169, N372);
not NOT1 (N1468, N1467);
nor NOR4 (N1469, N1463, N104, N605, N1305);
xor XOR2 (N1470, N1455, N854);
buf BUF1 (N1471, N1460);
or OR4 (N1472, N1462, N1437, N1390, N548);
and AND4 (N1473, N1450, N715, N1446, N1072);
nor NOR2 (N1474, N1441, N249);
nand NAND3 (N1475, N1474, N252, N389);
or OR2 (N1476, N1466, N964);
buf BUF1 (N1477, N1470);
buf BUF1 (N1478, N1464);
and AND2 (N1479, N1472, N1435);
not NOT1 (N1480, N1471);
and AND2 (N1481, N1461, N1266);
or OR4 (N1482, N1473, N1220, N985, N1298);
nor NOR4 (N1483, N1477, N911, N493, N1255);
buf BUF1 (N1484, N1480);
and AND4 (N1485, N1468, N1066, N587, N760);
or OR3 (N1486, N1478, N167, N1340);
not NOT1 (N1487, N1484);
nor NOR2 (N1488, N1476, N893);
nor NOR3 (N1489, N1487, N1141, N421);
buf BUF1 (N1490, N1469);
or OR4 (N1491, N1483, N57, N1211, N824);
or OR4 (N1492, N1479, N479, N192, N471);
or OR3 (N1493, N1481, N1075, N1002);
nor NOR3 (N1494, N1482, N1424, N1259);
nand NAND3 (N1495, N1491, N1293, N1106);
nand NAND2 (N1496, N1488, N360);
nor NOR2 (N1497, N1493, N443);
or OR4 (N1498, N1492, N1239, N525, N1482);
nand NAND3 (N1499, N1497, N691, N1334);
xor XOR2 (N1500, N1475, N628);
xor XOR2 (N1501, N1486, N468);
nand NAND4 (N1502, N1500, N592, N281, N541);
or OR2 (N1503, N1496, N979);
or OR4 (N1504, N1490, N1257, N375, N1234);
xor XOR2 (N1505, N1501, N255);
xor XOR2 (N1506, N1504, N268);
not NOT1 (N1507, N1503);
or OR3 (N1508, N1485, N934, N63);
and AND4 (N1509, N1508, N550, N162, N718);
xor XOR2 (N1510, N1505, N521);
nand NAND3 (N1511, N1489, N27, N1289);
and AND4 (N1512, N1511, N1407, N28, N229);
not NOT1 (N1513, N1498);
buf BUF1 (N1514, N1507);
not NOT1 (N1515, N1514);
endmodule