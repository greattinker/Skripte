// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N8008,N8018,N8020,N8005,N8009,N8016,N8011,N7993,N8019,N8021;

nor NOR4 (N22, N15, N19, N5, N3);
not NOT1 (N23, N9);
nor NOR4 (N24, N2, N7, N4, N2);
not NOT1 (N25, N11);
buf BUF1 (N26, N11);
nand NAND2 (N27, N8, N4);
nor NOR2 (N28, N7, N21);
not NOT1 (N29, N6);
nor NOR4 (N30, N8, N8, N1, N20);
or OR2 (N31, N6, N26);
or OR4 (N32, N5, N29, N18, N27);
nand NAND2 (N33, N20, N27);
buf BUF1 (N34, N26);
and AND2 (N35, N31, N21);
nand NAND3 (N36, N32, N10, N7);
nand NAND3 (N37, N33, N25, N23);
nand NAND3 (N38, N27, N8, N2);
nand NAND2 (N39, N6, N31);
xor XOR2 (N40, N39, N6);
xor XOR2 (N41, N38, N8);
not NOT1 (N42, N28);
buf BUF1 (N43, N34);
not NOT1 (N44, N41);
buf BUF1 (N45, N42);
or OR2 (N46, N22, N19);
xor XOR2 (N47, N40, N41);
nor NOR3 (N48, N44, N28, N34);
buf BUF1 (N49, N36);
nor NOR4 (N50, N49, N27, N38, N23);
and AND4 (N51, N37, N7, N47, N6);
nor NOR4 (N52, N25, N8, N36, N30);
and AND3 (N53, N12, N48, N20);
buf BUF1 (N54, N13);
and AND2 (N55, N43, N7);
not NOT1 (N56, N51);
nor NOR2 (N57, N52, N28);
and AND2 (N58, N55, N57);
and AND3 (N59, N48, N57, N43);
not NOT1 (N60, N46);
or OR4 (N61, N60, N18, N27, N37);
not NOT1 (N62, N54);
or OR2 (N63, N56, N21);
or OR2 (N64, N63, N38);
not NOT1 (N65, N53);
nor NOR2 (N66, N64, N11);
not NOT1 (N67, N58);
or OR2 (N68, N45, N42);
nand NAND4 (N69, N65, N10, N12, N45);
nor NOR3 (N70, N66, N24, N50);
nor NOR4 (N71, N41, N39, N57, N69);
nor NOR2 (N72, N15, N56);
buf BUF1 (N73, N71);
nor NOR3 (N74, N25, N39, N17);
nand NAND2 (N75, N62, N44);
nand NAND3 (N76, N67, N61, N39);
xor XOR2 (N77, N57, N71);
not NOT1 (N78, N75);
xor XOR2 (N79, N72, N19);
nor NOR4 (N80, N35, N79, N65, N44);
nand NAND3 (N81, N60, N39, N35);
buf BUF1 (N82, N74);
not NOT1 (N83, N73);
and AND3 (N84, N82, N17, N64);
nor NOR4 (N85, N81, N79, N22, N30);
or OR2 (N86, N77, N62);
not NOT1 (N87, N84);
and AND2 (N88, N68, N37);
buf BUF1 (N89, N87);
nand NAND3 (N90, N59, N25, N66);
buf BUF1 (N91, N89);
buf BUF1 (N92, N83);
buf BUF1 (N93, N92);
or OR4 (N94, N78, N69, N91, N29);
not NOT1 (N95, N27);
xor XOR2 (N96, N94, N66);
nand NAND3 (N97, N86, N39, N96);
nor NOR3 (N98, N57, N72, N8);
buf BUF1 (N99, N70);
nor NOR3 (N100, N98, N90, N53);
nand NAND4 (N101, N58, N10, N77, N32);
and AND4 (N102, N99, N32, N90, N80);
and AND3 (N103, N73, N14, N28);
nor NOR2 (N104, N88, N34);
nand NAND4 (N105, N103, N27, N39, N15);
buf BUF1 (N106, N85);
not NOT1 (N107, N97);
not NOT1 (N108, N102);
and AND3 (N109, N100, N88, N53);
or OR4 (N110, N101, N26, N58, N15);
buf BUF1 (N111, N110);
xor XOR2 (N112, N104, N2);
buf BUF1 (N113, N106);
not NOT1 (N114, N111);
or OR2 (N115, N93, N10);
nand NAND3 (N116, N105, N22, N37);
buf BUF1 (N117, N107);
nand NAND2 (N118, N113, N40);
buf BUF1 (N119, N117);
xor XOR2 (N120, N108, N8);
buf BUF1 (N121, N119);
nand NAND4 (N122, N121, N10, N25, N12);
nand NAND3 (N123, N116, N111, N2);
nand NAND4 (N124, N115, N78, N63, N94);
nand NAND4 (N125, N109, N116, N113, N34);
nand NAND4 (N126, N76, N57, N41, N12);
nor NOR4 (N127, N95, N45, N80, N45);
xor XOR2 (N128, N118, N89);
buf BUF1 (N129, N122);
nand NAND4 (N130, N127, N46, N29, N118);
or OR3 (N131, N123, N22, N122);
or OR3 (N132, N130, N1, N21);
nor NOR3 (N133, N125, N24, N128);
xor XOR2 (N134, N35, N5);
and AND4 (N135, N126, N97, N30, N132);
and AND2 (N136, N33, N3);
nor NOR4 (N137, N129, N110, N135, N81);
or OR4 (N138, N124, N120, N76, N27);
not NOT1 (N139, N13);
buf BUF1 (N140, N78);
nand NAND2 (N141, N140, N22);
and AND2 (N142, N131, N15);
and AND4 (N143, N137, N75, N75, N23);
or OR3 (N144, N112, N117, N85);
xor XOR2 (N145, N144, N110);
nand NAND3 (N146, N143, N139, N60);
buf BUF1 (N147, N13);
and AND3 (N148, N142, N87, N123);
or OR2 (N149, N148, N146);
nor NOR3 (N150, N140, N131, N32);
buf BUF1 (N151, N145);
and AND3 (N152, N136, N8, N120);
xor XOR2 (N153, N133, N136);
buf BUF1 (N154, N138);
nand NAND3 (N155, N141, N113, N59);
not NOT1 (N156, N154);
nor NOR2 (N157, N155, N23);
buf BUF1 (N158, N150);
xor XOR2 (N159, N157, N136);
xor XOR2 (N160, N147, N99);
or OR4 (N161, N153, N155, N81, N149);
buf BUF1 (N162, N83);
or OR2 (N163, N162, N142);
xor XOR2 (N164, N161, N158);
and AND4 (N165, N74, N53, N21, N73);
and AND3 (N166, N156, N104, N149);
not NOT1 (N167, N163);
and AND4 (N168, N167, N159, N69, N44);
buf BUF1 (N169, N79);
or OR4 (N170, N151, N159, N42, N107);
buf BUF1 (N171, N165);
nor NOR3 (N172, N160, N106, N58);
and AND2 (N173, N134, N167);
xor XOR2 (N174, N172, N134);
nand NAND3 (N175, N173, N162, N91);
buf BUF1 (N176, N170);
not NOT1 (N177, N166);
or OR2 (N178, N177, N110);
buf BUF1 (N179, N169);
buf BUF1 (N180, N168);
buf BUF1 (N181, N180);
and AND4 (N182, N164, N20, N106, N37);
not NOT1 (N183, N175);
xor XOR2 (N184, N183, N7);
xor XOR2 (N185, N179, N122);
buf BUF1 (N186, N171);
nor NOR3 (N187, N184, N28, N130);
xor XOR2 (N188, N178, N107);
nor NOR2 (N189, N181, N19);
or OR4 (N190, N188, N94, N88, N13);
nor NOR2 (N191, N187, N61);
not NOT1 (N192, N186);
xor XOR2 (N193, N152, N8);
not NOT1 (N194, N185);
nor NOR3 (N195, N191, N13, N113);
not NOT1 (N196, N182);
nand NAND3 (N197, N192, N26, N24);
or OR3 (N198, N174, N6, N23);
nand NAND2 (N199, N194, N193);
nor NOR4 (N200, N69, N183, N43, N54);
and AND2 (N201, N197, N151);
or OR3 (N202, N199, N200, N109);
nor NOR3 (N203, N40, N22, N157);
xor XOR2 (N204, N201, N159);
or OR3 (N205, N202, N113, N87);
nand NAND4 (N206, N195, N89, N45, N108);
nor NOR3 (N207, N196, N82, N185);
buf BUF1 (N208, N206);
nand NAND3 (N209, N207, N154, N187);
nand NAND4 (N210, N209, N204, N67, N207);
xor XOR2 (N211, N43, N112);
not NOT1 (N212, N205);
xor XOR2 (N213, N176, N138);
and AND3 (N214, N208, N52, N39);
and AND3 (N215, N213, N161, N71);
nand NAND4 (N216, N214, N24, N52, N82);
buf BUF1 (N217, N211);
and AND4 (N218, N190, N111, N63, N91);
or OR2 (N219, N198, N32);
and AND4 (N220, N219, N13, N73, N103);
nor NOR2 (N221, N114, N163);
and AND3 (N222, N215, N115, N159);
and AND4 (N223, N216, N97, N108, N162);
nor NOR4 (N224, N189, N92, N36, N87);
and AND3 (N225, N223, N125, N92);
nand NAND3 (N226, N221, N29, N185);
buf BUF1 (N227, N225);
and AND3 (N228, N222, N192, N188);
or OR2 (N229, N228, N108);
not NOT1 (N230, N227);
xor XOR2 (N231, N212, N125);
buf BUF1 (N232, N226);
buf BUF1 (N233, N203);
not NOT1 (N234, N232);
not NOT1 (N235, N231);
nand NAND3 (N236, N234, N150, N177);
and AND4 (N237, N218, N207, N162, N176);
or OR2 (N238, N217, N160);
not NOT1 (N239, N220);
nand NAND3 (N240, N233, N218, N157);
or OR2 (N241, N224, N221);
and AND4 (N242, N238, N214, N96, N13);
and AND4 (N243, N240, N22, N98, N102);
xor XOR2 (N244, N236, N134);
nand NAND4 (N245, N242, N69, N89, N232);
nor NOR2 (N246, N245, N125);
not NOT1 (N247, N237);
buf BUF1 (N248, N246);
and AND2 (N249, N235, N152);
nor NOR4 (N250, N210, N8, N87, N132);
nor NOR3 (N251, N230, N55, N243);
buf BUF1 (N252, N166);
xor XOR2 (N253, N247, N41);
nor NOR2 (N254, N251, N238);
not NOT1 (N255, N254);
xor XOR2 (N256, N248, N155);
xor XOR2 (N257, N250, N97);
or OR3 (N258, N229, N49, N46);
not NOT1 (N259, N256);
nand NAND4 (N260, N259, N26, N139, N225);
or OR3 (N261, N260, N149, N119);
nand NAND3 (N262, N249, N130, N122);
not NOT1 (N263, N261);
not NOT1 (N264, N263);
xor XOR2 (N265, N239, N214);
not NOT1 (N266, N253);
xor XOR2 (N267, N262, N165);
xor XOR2 (N268, N257, N145);
nand NAND4 (N269, N265, N187, N179, N82);
nand NAND3 (N270, N258, N188, N35);
nand NAND3 (N271, N269, N263, N80);
nand NAND4 (N272, N268, N157, N28, N76);
nand NAND4 (N273, N241, N29, N74, N168);
nand NAND4 (N274, N272, N247, N252, N236);
and AND3 (N275, N123, N222, N232);
and AND2 (N276, N270, N212);
and AND3 (N277, N274, N273, N203);
xor XOR2 (N278, N110, N110);
nor NOR3 (N279, N275, N238, N167);
xor XOR2 (N280, N276, N232);
nor NOR2 (N281, N278, N241);
not NOT1 (N282, N281);
xor XOR2 (N283, N255, N122);
not NOT1 (N284, N244);
not NOT1 (N285, N284);
not NOT1 (N286, N267);
or OR2 (N287, N271, N254);
and AND4 (N288, N285, N175, N48, N146);
or OR2 (N289, N266, N242);
not NOT1 (N290, N280);
xor XOR2 (N291, N287, N180);
or OR2 (N292, N283, N24);
not NOT1 (N293, N291);
not NOT1 (N294, N288);
nor NOR4 (N295, N290, N260, N187, N200);
buf BUF1 (N296, N286);
nor NOR4 (N297, N292, N294, N80, N128);
or OR3 (N298, N192, N278, N181);
nand NAND4 (N299, N296, N54, N9, N266);
not NOT1 (N300, N277);
buf BUF1 (N301, N300);
nand NAND2 (N302, N297, N269);
and AND3 (N303, N279, N296, N227);
or OR2 (N304, N298, N114);
buf BUF1 (N305, N282);
nor NOR2 (N306, N289, N6);
or OR2 (N307, N302, N286);
and AND3 (N308, N299, N301, N141);
buf BUF1 (N309, N192);
and AND4 (N310, N306, N288, N136, N127);
not NOT1 (N311, N310);
not NOT1 (N312, N304);
nor NOR3 (N313, N311, N34, N240);
xor XOR2 (N314, N293, N271);
buf BUF1 (N315, N295);
or OR4 (N316, N312, N105, N121, N33);
xor XOR2 (N317, N264, N276);
or OR2 (N318, N307, N272);
nor NOR2 (N319, N314, N122);
xor XOR2 (N320, N317, N19);
nand NAND4 (N321, N316, N191, N165, N190);
buf BUF1 (N322, N308);
buf BUF1 (N323, N322);
not NOT1 (N324, N320);
xor XOR2 (N325, N303, N48);
not NOT1 (N326, N325);
nor NOR4 (N327, N319, N153, N304, N75);
not NOT1 (N328, N309);
or OR3 (N329, N315, N56, N327);
xor XOR2 (N330, N160, N295);
or OR2 (N331, N326, N300);
not NOT1 (N332, N330);
and AND4 (N333, N323, N207, N298, N84);
buf BUF1 (N334, N329);
nand NAND2 (N335, N321, N18);
and AND2 (N336, N334, N331);
not NOT1 (N337, N155);
not NOT1 (N338, N333);
buf BUF1 (N339, N332);
or OR3 (N340, N324, N195, N249);
or OR3 (N341, N337, N238, N335);
buf BUF1 (N342, N110);
nand NAND4 (N343, N338, N229, N46, N154);
buf BUF1 (N344, N339);
nor NOR4 (N345, N343, N284, N321, N302);
nand NAND2 (N346, N345, N261);
not NOT1 (N347, N305);
buf BUF1 (N348, N336);
not NOT1 (N349, N341);
nand NAND2 (N350, N342, N39);
nor NOR4 (N351, N328, N141, N246, N205);
xor XOR2 (N352, N350, N19);
xor XOR2 (N353, N313, N245);
nand NAND4 (N354, N351, N182, N68, N42);
and AND2 (N355, N346, N237);
xor XOR2 (N356, N355, N14);
nand NAND2 (N357, N344, N309);
nand NAND2 (N358, N357, N281);
nand NAND4 (N359, N358, N39, N102, N147);
or OR2 (N360, N354, N184);
buf BUF1 (N361, N359);
and AND3 (N362, N353, N346, N6);
not NOT1 (N363, N347);
buf BUF1 (N364, N340);
xor XOR2 (N365, N348, N296);
buf BUF1 (N366, N356);
nor NOR4 (N367, N318, N90, N354, N230);
not NOT1 (N368, N366);
xor XOR2 (N369, N361, N90);
and AND2 (N370, N362, N283);
nor NOR4 (N371, N369, N256, N21, N322);
nand NAND3 (N372, N371, N359, N346);
nand NAND2 (N373, N370, N313);
buf BUF1 (N374, N352);
not NOT1 (N375, N364);
nor NOR2 (N376, N367, N181);
xor XOR2 (N377, N375, N162);
nor NOR4 (N378, N373, N121, N340, N275);
xor XOR2 (N379, N360, N2);
or OR4 (N380, N368, N47, N317, N281);
nand NAND3 (N381, N377, N267, N19);
nor NOR3 (N382, N365, N343, N292);
nand NAND3 (N383, N363, N82, N207);
buf BUF1 (N384, N383);
not NOT1 (N385, N376);
not NOT1 (N386, N380);
or OR4 (N387, N372, N172, N374, N103);
nor NOR2 (N388, N357, N281);
xor XOR2 (N389, N384, N235);
buf BUF1 (N390, N389);
and AND2 (N391, N382, N72);
xor XOR2 (N392, N386, N207);
and AND2 (N393, N387, N295);
not NOT1 (N394, N349);
and AND2 (N395, N378, N93);
nand NAND2 (N396, N385, N344);
and AND3 (N397, N393, N396, N49);
and AND4 (N398, N265, N337, N125, N75);
buf BUF1 (N399, N391);
buf BUF1 (N400, N398);
not NOT1 (N401, N392);
not NOT1 (N402, N395);
nand NAND4 (N403, N400, N251, N210, N10);
buf BUF1 (N404, N403);
or OR3 (N405, N394, N204, N258);
xor XOR2 (N406, N404, N21);
nor NOR3 (N407, N399, N51, N17);
and AND3 (N408, N388, N305, N31);
or OR4 (N409, N405, N159, N98, N233);
not NOT1 (N410, N407);
nand NAND4 (N411, N408, N222, N304, N150);
nand NAND4 (N412, N381, N15, N218, N74);
buf BUF1 (N413, N390);
nor NOR2 (N414, N402, N409);
not NOT1 (N415, N288);
nor NOR2 (N416, N415, N219);
or OR2 (N417, N411, N45);
buf BUF1 (N418, N413);
nand NAND2 (N419, N401, N159);
nand NAND2 (N420, N379, N163);
nand NAND2 (N421, N420, N99);
nand NAND4 (N422, N414, N67, N256, N56);
nor NOR3 (N423, N397, N285, N212);
nand NAND2 (N424, N416, N193);
not NOT1 (N425, N419);
not NOT1 (N426, N423);
buf BUF1 (N427, N422);
xor XOR2 (N428, N425, N139);
xor XOR2 (N429, N418, N263);
and AND4 (N430, N426, N313, N198, N215);
nand NAND3 (N431, N428, N113, N239);
nand NAND2 (N432, N412, N230);
or OR2 (N433, N430, N222);
not NOT1 (N434, N406);
not NOT1 (N435, N410);
nor NOR2 (N436, N417, N40);
or OR4 (N437, N434, N137, N188, N409);
nor NOR2 (N438, N435, N323);
or OR4 (N439, N433, N91, N57, N342);
nor NOR2 (N440, N439, N192);
xor XOR2 (N441, N440, N55);
not NOT1 (N442, N429);
and AND3 (N443, N427, N413, N303);
nor NOR2 (N444, N436, N125);
nand NAND4 (N445, N421, N366, N53, N245);
nor NOR2 (N446, N441, N383);
buf BUF1 (N447, N437);
nor NOR3 (N448, N444, N62, N432);
nor NOR2 (N449, N292, N48);
xor XOR2 (N450, N449, N335);
not NOT1 (N451, N424);
nand NAND2 (N452, N446, N264);
nor NOR2 (N453, N452, N223);
nor NOR3 (N454, N438, N317, N227);
nor NOR3 (N455, N431, N239, N391);
not NOT1 (N456, N450);
nand NAND2 (N457, N451, N168);
buf BUF1 (N458, N447);
buf BUF1 (N459, N456);
or OR4 (N460, N448, N133, N184, N294);
nor NOR2 (N461, N453, N23);
nor NOR3 (N462, N445, N182, N342);
not NOT1 (N463, N455);
nand NAND2 (N464, N461, N387);
xor XOR2 (N465, N443, N406);
xor XOR2 (N466, N462, N7);
or OR4 (N467, N463, N22, N98, N188);
and AND3 (N468, N464, N44, N397);
buf BUF1 (N469, N467);
nand NAND2 (N470, N465, N189);
not NOT1 (N471, N469);
xor XOR2 (N472, N457, N65);
buf BUF1 (N473, N454);
xor XOR2 (N474, N466, N164);
nor NOR3 (N475, N468, N193, N116);
nand NAND2 (N476, N475, N82);
nor NOR2 (N477, N459, N399);
and AND4 (N478, N442, N130, N283, N175);
nand NAND4 (N479, N458, N358, N149, N154);
buf BUF1 (N480, N471);
buf BUF1 (N481, N473);
not NOT1 (N482, N472);
xor XOR2 (N483, N477, N51);
xor XOR2 (N484, N483, N30);
xor XOR2 (N485, N481, N278);
not NOT1 (N486, N480);
not NOT1 (N487, N474);
and AND3 (N488, N482, N100, N144);
and AND3 (N489, N486, N130, N435);
or OR2 (N490, N476, N304);
xor XOR2 (N491, N488, N348);
xor XOR2 (N492, N460, N475);
or OR4 (N493, N489, N59, N313, N217);
buf BUF1 (N494, N485);
nand NAND3 (N495, N484, N492, N261);
nand NAND2 (N496, N431, N128);
not NOT1 (N497, N470);
not NOT1 (N498, N479);
and AND2 (N499, N496, N447);
and AND2 (N500, N491, N64);
nand NAND2 (N501, N493, N139);
xor XOR2 (N502, N490, N440);
nor NOR2 (N503, N499, N421);
not NOT1 (N504, N500);
buf BUF1 (N505, N487);
xor XOR2 (N506, N505, N123);
xor XOR2 (N507, N478, N172);
and AND2 (N508, N494, N221);
buf BUF1 (N509, N501);
not NOT1 (N510, N509);
and AND2 (N511, N504, N424);
nor NOR2 (N512, N498, N292);
and AND4 (N513, N497, N387, N478, N319);
xor XOR2 (N514, N513, N437);
nor NOR2 (N515, N502, N468);
not NOT1 (N516, N511);
or OR4 (N517, N506, N462, N461, N399);
buf BUF1 (N518, N503);
nor NOR2 (N519, N518, N25);
nand NAND2 (N520, N495, N350);
nand NAND3 (N521, N510, N264, N473);
not NOT1 (N522, N516);
or OR3 (N523, N515, N129, N259);
nand NAND3 (N524, N507, N364, N129);
buf BUF1 (N525, N519);
or OR3 (N526, N525, N373, N7);
buf BUF1 (N527, N524);
not NOT1 (N528, N514);
xor XOR2 (N529, N528, N102);
nor NOR3 (N530, N521, N331, N178);
or OR2 (N531, N508, N433);
buf BUF1 (N532, N527);
nand NAND3 (N533, N520, N24, N9);
buf BUF1 (N534, N517);
or OR2 (N535, N523, N129);
xor XOR2 (N536, N512, N258);
not NOT1 (N537, N536);
nor NOR2 (N538, N522, N144);
nand NAND4 (N539, N532, N160, N68, N428);
xor XOR2 (N540, N530, N39);
buf BUF1 (N541, N533);
and AND2 (N542, N541, N302);
nor NOR4 (N543, N542, N182, N405, N170);
not NOT1 (N544, N540);
nor NOR2 (N545, N529, N367);
and AND4 (N546, N545, N454, N529, N252);
nor NOR4 (N547, N544, N433, N289, N154);
and AND4 (N548, N534, N214, N312, N415);
xor XOR2 (N549, N535, N536);
buf BUF1 (N550, N548);
nor NOR3 (N551, N538, N487, N211);
xor XOR2 (N552, N546, N362);
and AND2 (N553, N550, N351);
nand NAND4 (N554, N553, N231, N368, N184);
not NOT1 (N555, N551);
not NOT1 (N556, N555);
buf BUF1 (N557, N537);
nand NAND4 (N558, N554, N21, N101, N191);
nor NOR2 (N559, N547, N233);
nor NOR2 (N560, N557, N139);
buf BUF1 (N561, N543);
buf BUF1 (N562, N559);
not NOT1 (N563, N539);
nor NOR4 (N564, N552, N409, N65, N154);
and AND2 (N565, N549, N345);
nand NAND2 (N566, N561, N207);
nor NOR3 (N567, N562, N90, N242);
xor XOR2 (N568, N567, N365);
not NOT1 (N569, N566);
nand NAND2 (N570, N563, N504);
and AND2 (N571, N558, N66);
xor XOR2 (N572, N560, N259);
buf BUF1 (N573, N531);
xor XOR2 (N574, N565, N309);
xor XOR2 (N575, N573, N141);
or OR4 (N576, N575, N232, N127, N97);
or OR3 (N577, N570, N476, N331);
nor NOR4 (N578, N576, N379, N65, N104);
or OR3 (N579, N571, N363, N163);
or OR4 (N580, N556, N496, N514, N1);
or OR2 (N581, N564, N81);
buf BUF1 (N582, N580);
xor XOR2 (N583, N572, N248);
nand NAND4 (N584, N574, N34, N256, N40);
buf BUF1 (N585, N583);
not NOT1 (N586, N579);
nor NOR2 (N587, N568, N559);
nand NAND3 (N588, N584, N177, N226);
nand NAND3 (N589, N581, N507, N40);
not NOT1 (N590, N588);
nand NAND2 (N591, N589, N4);
xor XOR2 (N592, N569, N62);
or OR3 (N593, N592, N193, N221);
buf BUF1 (N594, N582);
nor NOR2 (N595, N577, N269);
xor XOR2 (N596, N578, N432);
not NOT1 (N597, N594);
or OR2 (N598, N590, N212);
not NOT1 (N599, N587);
nor NOR2 (N600, N591, N400);
nor NOR3 (N601, N586, N70, N209);
or OR4 (N602, N595, N114, N331, N268);
buf BUF1 (N603, N585);
or OR2 (N604, N602, N289);
buf BUF1 (N605, N600);
buf BUF1 (N606, N605);
or OR2 (N607, N598, N173);
nor NOR2 (N608, N597, N468);
or OR3 (N609, N608, N271, N2);
nor NOR2 (N610, N599, N147);
buf BUF1 (N611, N610);
not NOT1 (N612, N603);
xor XOR2 (N613, N593, N343);
or OR4 (N614, N609, N336, N215, N551);
nand NAND4 (N615, N614, N261, N611, N291);
xor XOR2 (N616, N245, N14);
not NOT1 (N617, N526);
and AND3 (N618, N613, N40, N115);
xor XOR2 (N619, N612, N522);
and AND2 (N620, N607, N527);
not NOT1 (N621, N616);
nand NAND2 (N622, N620, N614);
buf BUF1 (N623, N621);
not NOT1 (N624, N604);
buf BUF1 (N625, N619);
nand NAND2 (N626, N624, N468);
buf BUF1 (N627, N622);
nand NAND4 (N628, N618, N383, N444, N413);
not NOT1 (N629, N615);
nor NOR2 (N630, N601, N356);
and AND2 (N631, N627, N614);
buf BUF1 (N632, N629);
and AND3 (N633, N623, N595, N180);
not NOT1 (N634, N632);
and AND3 (N635, N630, N72, N412);
or OR2 (N636, N628, N217);
or OR4 (N637, N633, N47, N416, N76);
nor NOR2 (N638, N634, N377);
not NOT1 (N639, N606);
buf BUF1 (N640, N626);
xor XOR2 (N641, N636, N360);
xor XOR2 (N642, N641, N190);
nand NAND4 (N643, N625, N524, N238, N14);
nand NAND4 (N644, N638, N251, N162, N52);
xor XOR2 (N645, N644, N159);
nand NAND4 (N646, N645, N378, N246, N64);
not NOT1 (N647, N646);
or OR4 (N648, N637, N97, N507, N316);
xor XOR2 (N649, N640, N5);
nand NAND2 (N650, N631, N578);
nor NOR3 (N651, N639, N319, N524);
and AND4 (N652, N649, N406, N480, N373);
buf BUF1 (N653, N642);
nor NOR2 (N654, N643, N239);
nor NOR2 (N655, N647, N116);
xor XOR2 (N656, N635, N11);
not NOT1 (N657, N652);
nor NOR4 (N658, N650, N390, N477, N625);
and AND4 (N659, N657, N156, N269, N398);
xor XOR2 (N660, N656, N159);
or OR2 (N661, N659, N70);
and AND4 (N662, N651, N136, N18, N434);
and AND2 (N663, N658, N51);
or OR4 (N664, N660, N317, N612, N279);
or OR3 (N665, N655, N542, N483);
buf BUF1 (N666, N596);
buf BUF1 (N667, N617);
buf BUF1 (N668, N654);
nand NAND2 (N669, N653, N326);
or OR3 (N670, N663, N505, N42);
not NOT1 (N671, N665);
and AND4 (N672, N661, N133, N391, N602);
and AND2 (N673, N666, N276);
buf BUF1 (N674, N667);
or OR2 (N675, N672, N443);
nor NOR3 (N676, N674, N629, N584);
nand NAND3 (N677, N670, N430, N271);
xor XOR2 (N678, N669, N274);
not NOT1 (N679, N675);
xor XOR2 (N680, N664, N571);
or OR2 (N681, N668, N449);
xor XOR2 (N682, N678, N368);
nand NAND2 (N683, N677, N159);
or OR2 (N684, N662, N127);
or OR2 (N685, N676, N35);
xor XOR2 (N686, N681, N675);
or OR4 (N687, N671, N604, N389, N559);
buf BUF1 (N688, N673);
or OR4 (N689, N680, N11, N639, N575);
nand NAND2 (N690, N684, N124);
buf BUF1 (N691, N679);
nor NOR4 (N692, N689, N262, N429, N97);
nand NAND2 (N693, N648, N517);
not NOT1 (N694, N690);
and AND4 (N695, N693, N290, N688, N402);
nor NOR4 (N696, N615, N493, N92, N63);
xor XOR2 (N697, N696, N132);
nand NAND2 (N698, N694, N460);
xor XOR2 (N699, N687, N144);
xor XOR2 (N700, N691, N40);
not NOT1 (N701, N699);
not NOT1 (N702, N700);
not NOT1 (N703, N698);
xor XOR2 (N704, N683, N457);
or OR3 (N705, N697, N178, N465);
xor XOR2 (N706, N703, N557);
nor NOR4 (N707, N705, N596, N522, N45);
buf BUF1 (N708, N692);
or OR3 (N709, N695, N497, N520);
nand NAND3 (N710, N708, N197, N204);
and AND2 (N711, N707, N486);
not NOT1 (N712, N701);
xor XOR2 (N713, N706, N550);
xor XOR2 (N714, N682, N491);
and AND4 (N715, N686, N468, N10, N98);
not NOT1 (N716, N711);
xor XOR2 (N717, N709, N1);
not NOT1 (N718, N685);
or OR3 (N719, N718, N345, N692);
nand NAND2 (N720, N719, N640);
and AND3 (N721, N716, N57, N670);
nor NOR3 (N722, N721, N79, N234);
and AND3 (N723, N715, N257, N70);
or OR3 (N724, N717, N139, N342);
buf BUF1 (N725, N713);
nor NOR2 (N726, N722, N545);
nor NOR4 (N727, N710, N77, N430, N448);
or OR2 (N728, N725, N430);
buf BUF1 (N729, N728);
not NOT1 (N730, N726);
nor NOR2 (N731, N714, N225);
xor XOR2 (N732, N730, N365);
buf BUF1 (N733, N727);
or OR3 (N734, N733, N442, N677);
xor XOR2 (N735, N702, N210);
nor NOR2 (N736, N732, N435);
and AND2 (N737, N734, N544);
or OR2 (N738, N735, N154);
nand NAND4 (N739, N712, N531, N405, N259);
nand NAND4 (N740, N739, N358, N551, N705);
and AND2 (N741, N724, N526);
and AND4 (N742, N704, N171, N385, N215);
xor XOR2 (N743, N738, N33);
and AND3 (N744, N720, N414, N389);
or OR4 (N745, N731, N225, N81, N632);
nand NAND2 (N746, N745, N229);
xor XOR2 (N747, N744, N664);
xor XOR2 (N748, N741, N31);
xor XOR2 (N749, N742, N344);
buf BUF1 (N750, N740);
buf BUF1 (N751, N736);
nor NOR3 (N752, N748, N517, N154);
buf BUF1 (N753, N743);
or OR2 (N754, N751, N343);
xor XOR2 (N755, N723, N464);
nand NAND2 (N756, N746, N219);
nand NAND2 (N757, N747, N129);
xor XOR2 (N758, N737, N136);
nor NOR4 (N759, N752, N108, N262, N643);
buf BUF1 (N760, N758);
and AND4 (N761, N760, N717, N342, N114);
not NOT1 (N762, N754);
not NOT1 (N763, N761);
buf BUF1 (N764, N750);
and AND4 (N765, N755, N234, N648, N124);
and AND2 (N766, N765, N560);
buf BUF1 (N767, N749);
nor NOR2 (N768, N764, N623);
and AND4 (N769, N757, N559, N539, N104);
or OR2 (N770, N759, N416);
not NOT1 (N771, N729);
xor XOR2 (N772, N763, N353);
xor XOR2 (N773, N756, N197);
nand NAND2 (N774, N768, N634);
and AND2 (N775, N767, N295);
buf BUF1 (N776, N762);
nor NOR2 (N777, N774, N319);
xor XOR2 (N778, N771, N625);
and AND3 (N779, N773, N549, N90);
nand NAND2 (N780, N778, N304);
nand NAND4 (N781, N776, N38, N674, N110);
nand NAND2 (N782, N769, N614);
xor XOR2 (N783, N753, N574);
buf BUF1 (N784, N781);
buf BUF1 (N785, N770);
nand NAND2 (N786, N766, N135);
not NOT1 (N787, N784);
nand NAND2 (N788, N780, N286);
and AND2 (N789, N775, N204);
nor NOR2 (N790, N789, N381);
not NOT1 (N791, N772);
buf BUF1 (N792, N790);
buf BUF1 (N793, N786);
nor NOR4 (N794, N788, N786, N571, N244);
not NOT1 (N795, N779);
buf BUF1 (N796, N777);
or OR2 (N797, N795, N704);
not NOT1 (N798, N796);
and AND4 (N799, N783, N185, N307, N792);
buf BUF1 (N800, N667);
not NOT1 (N801, N800);
not NOT1 (N802, N801);
and AND3 (N803, N802, N748, N422);
nand NAND3 (N804, N787, N17, N40);
nor NOR2 (N805, N803, N113);
buf BUF1 (N806, N799);
xor XOR2 (N807, N798, N362);
nor NOR3 (N808, N797, N516, N313);
not NOT1 (N809, N808);
nand NAND3 (N810, N794, N30, N727);
nor NOR4 (N811, N782, N557, N568, N752);
buf BUF1 (N812, N811);
or OR4 (N813, N809, N725, N17, N49);
nor NOR4 (N814, N806, N330, N554, N131);
buf BUF1 (N815, N814);
nand NAND3 (N816, N785, N20, N737);
buf BUF1 (N817, N793);
xor XOR2 (N818, N817, N738);
and AND4 (N819, N812, N398, N382, N507);
not NOT1 (N820, N810);
not NOT1 (N821, N816);
buf BUF1 (N822, N815);
nand NAND2 (N823, N820, N177);
and AND4 (N824, N807, N112, N415, N208);
and AND4 (N825, N822, N181, N477, N537);
or OR4 (N826, N819, N457, N23, N629);
buf BUF1 (N827, N825);
or OR4 (N828, N818, N560, N788, N756);
and AND4 (N829, N804, N254, N683, N176);
not NOT1 (N830, N824);
xor XOR2 (N831, N823, N828);
nand NAND2 (N832, N469, N38);
buf BUF1 (N833, N827);
and AND2 (N834, N813, N819);
not NOT1 (N835, N791);
buf BUF1 (N836, N834);
nand NAND4 (N837, N830, N178, N172, N648);
and AND2 (N838, N835, N398);
nor NOR4 (N839, N836, N358, N705, N672);
buf BUF1 (N840, N821);
nand NAND2 (N841, N831, N118);
xor XOR2 (N842, N805, N300);
nor NOR4 (N843, N841, N792, N643, N387);
nor NOR4 (N844, N833, N279, N265, N246);
and AND2 (N845, N843, N31);
nand NAND2 (N846, N837, N40);
xor XOR2 (N847, N840, N697);
nor NOR4 (N848, N829, N472, N521, N179);
xor XOR2 (N849, N847, N419);
xor XOR2 (N850, N846, N630);
nor NOR2 (N851, N844, N310);
nand NAND2 (N852, N832, N590);
xor XOR2 (N853, N848, N848);
xor XOR2 (N854, N851, N99);
nand NAND3 (N855, N850, N439, N755);
nand NAND4 (N856, N839, N829, N607, N851);
nand NAND4 (N857, N856, N501, N533, N18);
nor NOR4 (N858, N845, N237, N90, N463);
or OR3 (N859, N854, N599, N646);
and AND3 (N860, N852, N441, N400);
buf BUF1 (N861, N855);
nor NOR2 (N862, N861, N241);
or OR4 (N863, N842, N53, N75, N595);
and AND3 (N864, N858, N98, N472);
not NOT1 (N865, N863);
or OR2 (N866, N860, N354);
buf BUF1 (N867, N853);
xor XOR2 (N868, N849, N712);
or OR2 (N869, N867, N556);
not NOT1 (N870, N866);
and AND3 (N871, N870, N627, N800);
nand NAND4 (N872, N838, N566, N624, N625);
nand NAND3 (N873, N864, N834, N354);
nand NAND3 (N874, N873, N311, N174);
nand NAND2 (N875, N868, N611);
not NOT1 (N876, N826);
nand NAND2 (N877, N865, N568);
nand NAND2 (N878, N874, N827);
nor NOR4 (N879, N877, N177, N414, N196);
buf BUF1 (N880, N878);
or OR2 (N881, N876, N449);
or OR4 (N882, N879, N747, N244, N76);
or OR4 (N883, N880, N390, N156, N439);
xor XOR2 (N884, N875, N508);
nor NOR3 (N885, N857, N131, N591);
and AND3 (N886, N859, N281, N136);
buf BUF1 (N887, N871);
not NOT1 (N888, N883);
nand NAND3 (N889, N888, N594, N260);
nand NAND3 (N890, N881, N513, N854);
nand NAND3 (N891, N887, N787, N885);
xor XOR2 (N892, N345, N221);
or OR4 (N893, N882, N156, N661, N193);
nand NAND3 (N894, N872, N616, N664);
and AND4 (N895, N886, N185, N63, N204);
not NOT1 (N896, N890);
nor NOR2 (N897, N862, N17);
nand NAND3 (N898, N894, N489, N863);
nor NOR3 (N899, N897, N690, N85);
buf BUF1 (N900, N892);
buf BUF1 (N901, N898);
or OR4 (N902, N901, N180, N508, N546);
nand NAND4 (N903, N902, N518, N260, N824);
buf BUF1 (N904, N899);
or OR4 (N905, N893, N510, N673, N866);
and AND2 (N906, N889, N368);
xor XOR2 (N907, N903, N606);
and AND4 (N908, N891, N871, N337, N264);
or OR2 (N909, N908, N485);
not NOT1 (N910, N884);
xor XOR2 (N911, N909, N694);
nand NAND2 (N912, N900, N108);
not NOT1 (N913, N869);
or OR2 (N914, N906, N416);
nand NAND3 (N915, N914, N812, N357);
and AND3 (N916, N912, N784, N298);
xor XOR2 (N917, N916, N12);
or OR4 (N918, N904, N644, N761, N755);
nand NAND2 (N919, N913, N538);
not NOT1 (N920, N896);
nand NAND2 (N921, N917, N417);
nor NOR3 (N922, N920, N410, N223);
or OR4 (N923, N922, N755, N360, N647);
or OR3 (N924, N919, N622, N651);
buf BUF1 (N925, N910);
nand NAND3 (N926, N925, N276, N614);
not NOT1 (N927, N918);
nor NOR4 (N928, N895, N66, N597, N578);
nand NAND2 (N929, N907, N408);
and AND3 (N930, N928, N448, N846);
nand NAND2 (N931, N927, N553);
nand NAND3 (N932, N926, N422, N397);
nor NOR2 (N933, N905, N595);
not NOT1 (N934, N924);
not NOT1 (N935, N932);
xor XOR2 (N936, N934, N208);
nor NOR3 (N937, N931, N663, N47);
and AND4 (N938, N935, N776, N819, N761);
not NOT1 (N939, N921);
nand NAND3 (N940, N936, N192, N501);
not NOT1 (N941, N939);
and AND4 (N942, N911, N575, N775, N509);
xor XOR2 (N943, N938, N578);
xor XOR2 (N944, N940, N373);
nand NAND4 (N945, N944, N744, N48, N457);
and AND2 (N946, N915, N452);
and AND2 (N947, N937, N705);
buf BUF1 (N948, N933);
and AND4 (N949, N930, N724, N18, N831);
nor NOR4 (N950, N943, N936, N349, N164);
nand NAND2 (N951, N946, N100);
not NOT1 (N952, N942);
xor XOR2 (N953, N947, N256);
or OR2 (N954, N948, N565);
and AND4 (N955, N954, N271, N946, N714);
nor NOR4 (N956, N950, N400, N374, N47);
nand NAND3 (N957, N945, N149, N207);
buf BUF1 (N958, N941);
nand NAND3 (N959, N957, N931, N384);
xor XOR2 (N960, N923, N651);
xor XOR2 (N961, N949, N33);
not NOT1 (N962, N955);
or OR4 (N963, N959, N192, N728, N641);
nand NAND2 (N964, N953, N411);
buf BUF1 (N965, N951);
or OR4 (N966, N962, N433, N761, N24);
nor NOR3 (N967, N961, N102, N60);
nor NOR3 (N968, N965, N291, N382);
nand NAND2 (N969, N929, N9);
and AND2 (N970, N956, N11);
nand NAND4 (N971, N963, N93, N95, N948);
xor XOR2 (N972, N958, N476);
nand NAND2 (N973, N968, N570);
not NOT1 (N974, N971);
nor NOR2 (N975, N970, N89);
buf BUF1 (N976, N952);
and AND3 (N977, N976, N281, N441);
nand NAND4 (N978, N974, N458, N765, N860);
nand NAND3 (N979, N977, N474, N641);
buf BUF1 (N980, N966);
and AND3 (N981, N972, N471, N492);
not NOT1 (N982, N980);
buf BUF1 (N983, N975);
xor XOR2 (N984, N982, N880);
and AND3 (N985, N978, N212, N165);
and AND4 (N986, N967, N254, N67, N443);
buf BUF1 (N987, N960);
buf BUF1 (N988, N987);
and AND2 (N989, N979, N747);
and AND3 (N990, N981, N493, N808);
buf BUF1 (N991, N973);
not NOT1 (N992, N990);
xor XOR2 (N993, N984, N152);
or OR3 (N994, N985, N778, N992);
nand NAND2 (N995, N791, N944);
buf BUF1 (N996, N964);
nand NAND2 (N997, N969, N48);
nand NAND2 (N998, N996, N242);
and AND4 (N999, N998, N173, N249, N603);
nor NOR3 (N1000, N991, N998, N542);
nand NAND4 (N1001, N983, N516, N844, N354);
not NOT1 (N1002, N994);
nor NOR2 (N1003, N989, N91);
nand NAND3 (N1004, N997, N562, N179);
buf BUF1 (N1005, N988);
not NOT1 (N1006, N1005);
or OR4 (N1007, N995, N327, N362, N196);
or OR3 (N1008, N1003, N904, N503);
or OR2 (N1009, N993, N754);
xor XOR2 (N1010, N1000, N853);
and AND4 (N1011, N1008, N330, N437, N562);
not NOT1 (N1012, N1006);
xor XOR2 (N1013, N1001, N549);
xor XOR2 (N1014, N999, N791);
or OR2 (N1015, N1013, N480);
nor NOR2 (N1016, N1004, N264);
nand NAND3 (N1017, N1012, N298, N790);
or OR2 (N1018, N1007, N184);
and AND2 (N1019, N1002, N986);
nor NOR4 (N1020, N376, N253, N582, N238);
and AND3 (N1021, N1020, N25, N968);
not NOT1 (N1022, N1009);
xor XOR2 (N1023, N1019, N802);
buf BUF1 (N1024, N1010);
or OR4 (N1025, N1022, N921, N184, N270);
not NOT1 (N1026, N1021);
not NOT1 (N1027, N1016);
nor NOR2 (N1028, N1026, N31);
buf BUF1 (N1029, N1011);
or OR3 (N1030, N1017, N536, N779);
not NOT1 (N1031, N1014);
or OR3 (N1032, N1018, N159, N228);
nor NOR4 (N1033, N1027, N926, N258, N541);
xor XOR2 (N1034, N1024, N970);
nand NAND4 (N1035, N1034, N961, N546, N83);
nor NOR2 (N1036, N1032, N186);
or OR4 (N1037, N1031, N104, N204, N396);
and AND4 (N1038, N1028, N889, N712, N718);
and AND3 (N1039, N1023, N629, N1026);
not NOT1 (N1040, N1039);
not NOT1 (N1041, N1015);
nand NAND3 (N1042, N1037, N107, N168);
buf BUF1 (N1043, N1025);
nand NAND3 (N1044, N1042, N837, N1027);
buf BUF1 (N1045, N1035);
buf BUF1 (N1046, N1030);
and AND3 (N1047, N1044, N999, N359);
nor NOR2 (N1048, N1045, N164);
buf BUF1 (N1049, N1041);
xor XOR2 (N1050, N1048, N70);
nor NOR3 (N1051, N1038, N458, N925);
buf BUF1 (N1052, N1050);
xor XOR2 (N1053, N1051, N75);
and AND2 (N1054, N1053, N979);
not NOT1 (N1055, N1046);
and AND3 (N1056, N1055, N244, N444);
nor NOR3 (N1057, N1040, N1027, N10);
not NOT1 (N1058, N1029);
or OR3 (N1059, N1036, N35, N290);
nor NOR3 (N1060, N1049, N380, N802);
buf BUF1 (N1061, N1056);
and AND2 (N1062, N1043, N367);
buf BUF1 (N1063, N1033);
and AND4 (N1064, N1057, N18, N7, N933);
or OR2 (N1065, N1054, N281);
and AND3 (N1066, N1063, N286, N533);
or OR4 (N1067, N1065, N295, N616, N365);
not NOT1 (N1068, N1059);
or OR3 (N1069, N1062, N1067, N451);
and AND4 (N1070, N544, N746, N538, N53);
nor NOR4 (N1071, N1066, N770, N463, N640);
or OR3 (N1072, N1064, N582, N164);
xor XOR2 (N1073, N1052, N156);
not NOT1 (N1074, N1072);
and AND2 (N1075, N1068, N346);
buf BUF1 (N1076, N1047);
nor NOR2 (N1077, N1060, N520);
nor NOR3 (N1078, N1058, N40, N701);
buf BUF1 (N1079, N1076);
buf BUF1 (N1080, N1075);
or OR3 (N1081, N1080, N757, N98);
and AND4 (N1082, N1079, N776, N860, N168);
or OR3 (N1083, N1082, N467, N279);
or OR3 (N1084, N1083, N634, N709);
and AND2 (N1085, N1081, N994);
and AND3 (N1086, N1070, N118, N461);
or OR4 (N1087, N1061, N499, N881, N856);
nor NOR3 (N1088, N1087, N406, N408);
not NOT1 (N1089, N1088);
or OR4 (N1090, N1071, N833, N931, N1003);
nand NAND3 (N1091, N1073, N333, N495);
buf BUF1 (N1092, N1084);
and AND4 (N1093, N1085, N197, N306, N564);
or OR3 (N1094, N1069, N1089, N1027);
and AND3 (N1095, N934, N396, N770);
xor XOR2 (N1096, N1093, N817);
xor XOR2 (N1097, N1077, N350);
nand NAND2 (N1098, N1090, N33);
not NOT1 (N1099, N1086);
nor NOR2 (N1100, N1091, N91);
and AND4 (N1101, N1074, N16, N563, N153);
nand NAND3 (N1102, N1098, N485, N559);
xor XOR2 (N1103, N1096, N574);
not NOT1 (N1104, N1101);
or OR2 (N1105, N1103, N818);
nor NOR2 (N1106, N1092, N460);
nor NOR3 (N1107, N1095, N998, N202);
or OR2 (N1108, N1099, N269);
xor XOR2 (N1109, N1100, N303);
buf BUF1 (N1110, N1106);
not NOT1 (N1111, N1078);
not NOT1 (N1112, N1097);
nand NAND2 (N1113, N1109, N962);
not NOT1 (N1114, N1112);
not NOT1 (N1115, N1114);
not NOT1 (N1116, N1115);
or OR4 (N1117, N1116, N545, N413, N406);
nand NAND3 (N1118, N1108, N142, N300);
nor NOR4 (N1119, N1111, N82, N691, N615);
nand NAND3 (N1120, N1102, N458, N759);
nor NOR4 (N1121, N1113, N528, N13, N1024);
buf BUF1 (N1122, N1120);
not NOT1 (N1123, N1117);
not NOT1 (N1124, N1104);
and AND3 (N1125, N1118, N501, N655);
and AND2 (N1126, N1110, N212);
and AND2 (N1127, N1122, N1006);
not NOT1 (N1128, N1127);
and AND4 (N1129, N1125, N1008, N39, N641);
not NOT1 (N1130, N1094);
buf BUF1 (N1131, N1124);
nand NAND3 (N1132, N1123, N785, N938);
nor NOR4 (N1133, N1130, N831, N502, N543);
buf BUF1 (N1134, N1129);
and AND3 (N1135, N1119, N216, N663);
nor NOR4 (N1136, N1134, N814, N672, N583);
nor NOR2 (N1137, N1131, N209);
or OR3 (N1138, N1126, N693, N476);
or OR2 (N1139, N1107, N634);
and AND4 (N1140, N1133, N964, N1109, N69);
or OR3 (N1141, N1121, N316, N814);
and AND2 (N1142, N1140, N893);
nand NAND3 (N1143, N1138, N213, N758);
nor NOR3 (N1144, N1139, N929, N77);
nor NOR4 (N1145, N1128, N945, N74, N431);
or OR3 (N1146, N1143, N282, N494);
and AND2 (N1147, N1135, N1112);
nor NOR2 (N1148, N1142, N564);
and AND4 (N1149, N1146, N534, N1005, N850);
xor XOR2 (N1150, N1137, N600);
nor NOR2 (N1151, N1150, N306);
not NOT1 (N1152, N1136);
and AND4 (N1153, N1149, N214, N1070, N394);
nor NOR4 (N1154, N1105, N1126, N914, N794);
buf BUF1 (N1155, N1147);
not NOT1 (N1156, N1152);
and AND4 (N1157, N1145, N46, N918, N284);
or OR2 (N1158, N1154, N825);
nor NOR3 (N1159, N1141, N765, N37);
nand NAND4 (N1160, N1159, N691, N1039, N846);
xor XOR2 (N1161, N1132, N41);
nor NOR2 (N1162, N1151, N442);
and AND4 (N1163, N1162, N641, N673, N895);
or OR3 (N1164, N1158, N876, N429);
nand NAND2 (N1165, N1161, N374);
nor NOR3 (N1166, N1165, N146, N459);
nor NOR4 (N1167, N1155, N150, N691, N1012);
nand NAND2 (N1168, N1148, N513);
not NOT1 (N1169, N1166);
not NOT1 (N1170, N1164);
and AND2 (N1171, N1170, N621);
or OR2 (N1172, N1160, N830);
nor NOR2 (N1173, N1169, N914);
and AND2 (N1174, N1167, N476);
and AND3 (N1175, N1168, N1046, N704);
buf BUF1 (N1176, N1174);
not NOT1 (N1177, N1176);
nor NOR4 (N1178, N1172, N438, N1049, N1108);
nand NAND4 (N1179, N1163, N375, N498, N681);
xor XOR2 (N1180, N1153, N1075);
not NOT1 (N1181, N1178);
not NOT1 (N1182, N1179);
or OR3 (N1183, N1181, N707, N705);
or OR4 (N1184, N1173, N10, N243, N794);
xor XOR2 (N1185, N1156, N707);
xor XOR2 (N1186, N1185, N1183);
or OR2 (N1187, N1094, N960);
nand NAND2 (N1188, N1182, N622);
and AND2 (N1189, N1187, N11);
nor NOR4 (N1190, N1177, N305, N24, N240);
not NOT1 (N1191, N1144);
not NOT1 (N1192, N1171);
xor XOR2 (N1193, N1180, N471);
and AND2 (N1194, N1175, N933);
buf BUF1 (N1195, N1192);
buf BUF1 (N1196, N1189);
nor NOR3 (N1197, N1184, N1187, N174);
not NOT1 (N1198, N1196);
buf BUF1 (N1199, N1191);
buf BUF1 (N1200, N1197);
xor XOR2 (N1201, N1195, N454);
or OR4 (N1202, N1199, N513, N597, N1030);
and AND4 (N1203, N1201, N707, N346, N40);
nand NAND4 (N1204, N1202, N189, N415, N361);
not NOT1 (N1205, N1188);
and AND2 (N1206, N1200, N505);
nand NAND2 (N1207, N1198, N649);
nor NOR2 (N1208, N1157, N244);
nand NAND2 (N1209, N1193, N1006);
and AND2 (N1210, N1204, N859);
nor NOR3 (N1211, N1208, N1199, N1072);
nand NAND3 (N1212, N1194, N611, N220);
or OR2 (N1213, N1210, N982);
buf BUF1 (N1214, N1206);
nor NOR4 (N1215, N1190, N816, N741, N405);
and AND4 (N1216, N1211, N178, N1031, N41);
buf BUF1 (N1217, N1209);
or OR4 (N1218, N1216, N462, N131, N38);
or OR3 (N1219, N1213, N915, N431);
nand NAND4 (N1220, N1219, N52, N434, N667);
buf BUF1 (N1221, N1207);
not NOT1 (N1222, N1215);
xor XOR2 (N1223, N1221, N734);
and AND2 (N1224, N1205, N26);
not NOT1 (N1225, N1220);
xor XOR2 (N1226, N1186, N180);
not NOT1 (N1227, N1214);
buf BUF1 (N1228, N1227);
xor XOR2 (N1229, N1203, N272);
not NOT1 (N1230, N1223);
not NOT1 (N1231, N1228);
or OR2 (N1232, N1224, N399);
not NOT1 (N1233, N1222);
nor NOR4 (N1234, N1229, N80, N824, N1069);
or OR3 (N1235, N1225, N503, N212);
or OR3 (N1236, N1226, N546, N531);
or OR3 (N1237, N1217, N653, N151);
or OR4 (N1238, N1235, N645, N1060, N1116);
xor XOR2 (N1239, N1212, N915);
nor NOR2 (N1240, N1234, N1217);
not NOT1 (N1241, N1230);
or OR4 (N1242, N1233, N831, N1160, N1083);
nor NOR3 (N1243, N1237, N911, N930);
xor XOR2 (N1244, N1243, N1053);
not NOT1 (N1245, N1241);
xor XOR2 (N1246, N1239, N1147);
or OR2 (N1247, N1232, N905);
nor NOR2 (N1248, N1231, N81);
nor NOR4 (N1249, N1240, N296, N1152, N975);
and AND4 (N1250, N1244, N130, N1118, N151);
buf BUF1 (N1251, N1218);
xor XOR2 (N1252, N1236, N474);
nand NAND2 (N1253, N1245, N630);
nor NOR3 (N1254, N1238, N120, N528);
nand NAND3 (N1255, N1249, N731, N522);
xor XOR2 (N1256, N1255, N570);
nand NAND4 (N1257, N1242, N333, N696, N445);
and AND3 (N1258, N1256, N903, N136);
not NOT1 (N1259, N1257);
buf BUF1 (N1260, N1258);
buf BUF1 (N1261, N1259);
and AND4 (N1262, N1250, N364, N1144, N759);
nand NAND3 (N1263, N1252, N267, N707);
not NOT1 (N1264, N1260);
or OR3 (N1265, N1247, N68, N292);
xor XOR2 (N1266, N1265, N744);
buf BUF1 (N1267, N1246);
buf BUF1 (N1268, N1253);
or OR3 (N1269, N1261, N308, N449);
xor XOR2 (N1270, N1268, N1199);
buf BUF1 (N1271, N1248);
nor NOR4 (N1272, N1269, N3, N39, N922);
and AND4 (N1273, N1251, N809, N475, N712);
not NOT1 (N1274, N1266);
or OR2 (N1275, N1273, N520);
nor NOR4 (N1276, N1271, N105, N1123, N465);
and AND4 (N1277, N1267, N501, N577, N336);
xor XOR2 (N1278, N1254, N1163);
xor XOR2 (N1279, N1270, N1146);
and AND4 (N1280, N1275, N138, N240, N318);
nand NAND3 (N1281, N1279, N482, N836);
not NOT1 (N1282, N1278);
or OR2 (N1283, N1263, N406);
buf BUF1 (N1284, N1280);
or OR3 (N1285, N1282, N37, N90);
nand NAND4 (N1286, N1284, N404, N100, N469);
nor NOR2 (N1287, N1285, N340);
not NOT1 (N1288, N1287);
nor NOR4 (N1289, N1281, N358, N444, N365);
buf BUF1 (N1290, N1286);
nor NOR2 (N1291, N1272, N58);
and AND3 (N1292, N1289, N808, N842);
buf BUF1 (N1293, N1290);
buf BUF1 (N1294, N1293);
nor NOR3 (N1295, N1294, N447, N111);
xor XOR2 (N1296, N1262, N1046);
nand NAND3 (N1297, N1283, N1157, N1196);
and AND3 (N1298, N1264, N239, N1037);
buf BUF1 (N1299, N1277);
nor NOR4 (N1300, N1276, N1279, N414, N105);
nand NAND2 (N1301, N1298, N188);
not NOT1 (N1302, N1296);
and AND2 (N1303, N1297, N14);
and AND3 (N1304, N1295, N150, N1277);
not NOT1 (N1305, N1292);
nand NAND3 (N1306, N1291, N1254, N260);
nand NAND4 (N1307, N1302, N1143, N1141, N282);
not NOT1 (N1308, N1306);
buf BUF1 (N1309, N1274);
or OR3 (N1310, N1288, N267, N498);
nor NOR2 (N1311, N1299, N400);
buf BUF1 (N1312, N1305);
xor XOR2 (N1313, N1308, N60);
nand NAND3 (N1314, N1303, N381, N492);
not NOT1 (N1315, N1301);
buf BUF1 (N1316, N1304);
xor XOR2 (N1317, N1309, N127);
not NOT1 (N1318, N1310);
and AND4 (N1319, N1318, N1275, N354, N1112);
buf BUF1 (N1320, N1311);
nor NOR3 (N1321, N1315, N549, N1094);
xor XOR2 (N1322, N1320, N581);
xor XOR2 (N1323, N1316, N196);
nand NAND4 (N1324, N1319, N864, N427, N989);
and AND2 (N1325, N1300, N213);
or OR4 (N1326, N1321, N1229, N841, N739);
nand NAND3 (N1327, N1317, N748, N25);
not NOT1 (N1328, N1307);
xor XOR2 (N1329, N1328, N225);
nand NAND4 (N1330, N1326, N322, N121, N1021);
and AND3 (N1331, N1313, N795, N874);
or OR2 (N1332, N1323, N1008);
nand NAND2 (N1333, N1322, N657);
nand NAND3 (N1334, N1314, N785, N1221);
xor XOR2 (N1335, N1330, N30);
xor XOR2 (N1336, N1329, N863);
nor NOR3 (N1337, N1325, N1256, N663);
not NOT1 (N1338, N1335);
nor NOR4 (N1339, N1334, N1294, N195, N1042);
xor XOR2 (N1340, N1336, N1050);
nand NAND3 (N1341, N1324, N179, N1150);
buf BUF1 (N1342, N1340);
or OR3 (N1343, N1339, N1285, N957);
or OR3 (N1344, N1342, N345, N1274);
and AND4 (N1345, N1312, N1237, N879, N1143);
xor XOR2 (N1346, N1337, N713);
nand NAND4 (N1347, N1343, N449, N397, N819);
nand NAND3 (N1348, N1345, N622, N65);
buf BUF1 (N1349, N1331);
xor XOR2 (N1350, N1332, N301);
buf BUF1 (N1351, N1348);
or OR2 (N1352, N1349, N685);
xor XOR2 (N1353, N1341, N324);
nand NAND3 (N1354, N1347, N1135, N1318);
nand NAND2 (N1355, N1344, N347);
not NOT1 (N1356, N1327);
nand NAND2 (N1357, N1333, N1226);
or OR3 (N1358, N1338, N94, N256);
xor XOR2 (N1359, N1352, N47);
buf BUF1 (N1360, N1355);
or OR4 (N1361, N1350, N681, N1335, N862);
and AND4 (N1362, N1357, N712, N1289, N1241);
not NOT1 (N1363, N1356);
not NOT1 (N1364, N1359);
and AND4 (N1365, N1346, N472, N1085, N954);
buf BUF1 (N1366, N1362);
nand NAND2 (N1367, N1358, N18);
nand NAND3 (N1368, N1351, N731, N1214);
xor XOR2 (N1369, N1366, N829);
nand NAND4 (N1370, N1367, N1012, N565, N599);
nand NAND3 (N1371, N1365, N618, N646);
nor NOR3 (N1372, N1368, N984, N397);
nand NAND2 (N1373, N1360, N1219);
not NOT1 (N1374, N1369);
and AND4 (N1375, N1374, N87, N640, N890);
nand NAND2 (N1376, N1353, N330);
and AND2 (N1377, N1370, N708);
nor NOR2 (N1378, N1371, N1130);
or OR2 (N1379, N1361, N539);
not NOT1 (N1380, N1377);
and AND3 (N1381, N1378, N343, N736);
xor XOR2 (N1382, N1376, N778);
and AND3 (N1383, N1372, N84, N154);
and AND2 (N1384, N1381, N414);
or OR2 (N1385, N1354, N1208);
or OR2 (N1386, N1385, N952);
xor XOR2 (N1387, N1379, N1061);
nand NAND3 (N1388, N1382, N601, N951);
buf BUF1 (N1389, N1363);
not NOT1 (N1390, N1388);
or OR3 (N1391, N1380, N146, N600);
xor XOR2 (N1392, N1375, N734);
nand NAND2 (N1393, N1373, N110);
and AND4 (N1394, N1391, N1029, N226, N144);
and AND3 (N1395, N1386, N1143, N105);
or OR3 (N1396, N1389, N1056, N634);
not NOT1 (N1397, N1396);
not NOT1 (N1398, N1384);
not NOT1 (N1399, N1364);
and AND4 (N1400, N1398, N1069, N762, N724);
xor XOR2 (N1401, N1394, N1259);
and AND4 (N1402, N1395, N634, N513, N1332);
or OR2 (N1403, N1387, N1381);
and AND3 (N1404, N1399, N1193, N429);
or OR4 (N1405, N1393, N85, N1260, N144);
xor XOR2 (N1406, N1401, N803);
xor XOR2 (N1407, N1405, N689);
buf BUF1 (N1408, N1407);
nor NOR2 (N1409, N1397, N1293);
nand NAND4 (N1410, N1408, N548, N1315, N244);
nand NAND3 (N1411, N1392, N348, N685);
or OR4 (N1412, N1403, N1093, N501, N659);
xor XOR2 (N1413, N1402, N199);
not NOT1 (N1414, N1390);
or OR2 (N1415, N1411, N565);
xor XOR2 (N1416, N1400, N1137);
xor XOR2 (N1417, N1414, N175);
nor NOR4 (N1418, N1410, N463, N310, N23);
not NOT1 (N1419, N1383);
nor NOR4 (N1420, N1404, N306, N780, N808);
xor XOR2 (N1421, N1412, N117);
or OR4 (N1422, N1416, N1354, N644, N741);
or OR3 (N1423, N1419, N747, N928);
nand NAND4 (N1424, N1421, N833, N1020, N135);
xor XOR2 (N1425, N1413, N510);
and AND3 (N1426, N1409, N590, N713);
not NOT1 (N1427, N1418);
nor NOR2 (N1428, N1415, N1141);
xor XOR2 (N1429, N1427, N1347);
and AND3 (N1430, N1428, N936, N1057);
nand NAND3 (N1431, N1424, N2, N610);
and AND3 (N1432, N1423, N702, N37);
buf BUF1 (N1433, N1420);
not NOT1 (N1434, N1429);
xor XOR2 (N1435, N1422, N1203);
and AND4 (N1436, N1435, N544, N1160, N542);
not NOT1 (N1437, N1431);
buf BUF1 (N1438, N1437);
xor XOR2 (N1439, N1430, N532);
nor NOR2 (N1440, N1425, N283);
nand NAND3 (N1441, N1426, N1048, N645);
buf BUF1 (N1442, N1434);
nand NAND4 (N1443, N1417, N554, N1357, N728);
xor XOR2 (N1444, N1441, N109);
xor XOR2 (N1445, N1444, N176);
nand NAND3 (N1446, N1438, N523, N1261);
and AND3 (N1447, N1446, N830, N876);
nand NAND3 (N1448, N1432, N380, N1206);
and AND3 (N1449, N1440, N330, N898);
and AND2 (N1450, N1433, N1135);
not NOT1 (N1451, N1450);
xor XOR2 (N1452, N1448, N945);
and AND3 (N1453, N1445, N531, N1396);
not NOT1 (N1454, N1449);
nand NAND2 (N1455, N1443, N533);
xor XOR2 (N1456, N1453, N1378);
nor NOR2 (N1457, N1451, N1017);
or OR2 (N1458, N1439, N564);
buf BUF1 (N1459, N1454);
not NOT1 (N1460, N1459);
nor NOR3 (N1461, N1447, N1305, N594);
not NOT1 (N1462, N1457);
not NOT1 (N1463, N1458);
nor NOR3 (N1464, N1455, N1283, N217);
nor NOR3 (N1465, N1436, N1041, N859);
xor XOR2 (N1466, N1463, N1367);
and AND4 (N1467, N1406, N388, N77, N1172);
or OR3 (N1468, N1452, N1396, N1396);
nor NOR4 (N1469, N1461, N286, N1388, N775);
xor XOR2 (N1470, N1462, N1095);
not NOT1 (N1471, N1465);
nor NOR2 (N1472, N1466, N246);
buf BUF1 (N1473, N1456);
nor NOR3 (N1474, N1471, N77, N977);
and AND2 (N1475, N1470, N1343);
nor NOR2 (N1476, N1464, N1325);
nor NOR3 (N1477, N1473, N626, N200);
or OR2 (N1478, N1468, N271);
not NOT1 (N1479, N1460);
nand NAND2 (N1480, N1472, N149);
and AND2 (N1481, N1478, N842);
xor XOR2 (N1482, N1480, N676);
not NOT1 (N1483, N1482);
not NOT1 (N1484, N1474);
buf BUF1 (N1485, N1476);
nor NOR4 (N1486, N1467, N99, N112, N158);
nor NOR2 (N1487, N1469, N1460);
xor XOR2 (N1488, N1475, N23);
buf BUF1 (N1489, N1488);
xor XOR2 (N1490, N1479, N188);
and AND3 (N1491, N1483, N646, N596);
or OR3 (N1492, N1490, N1450, N334);
or OR4 (N1493, N1484, N126, N88, N1245);
xor XOR2 (N1494, N1491, N240);
or OR3 (N1495, N1485, N1353, N1417);
or OR4 (N1496, N1487, N1061, N1186, N67);
or OR3 (N1497, N1442, N946, N1406);
nor NOR2 (N1498, N1486, N156);
and AND2 (N1499, N1477, N314);
nor NOR3 (N1500, N1499, N346, N1107);
nand NAND4 (N1501, N1500, N1026, N687, N726);
and AND3 (N1502, N1498, N198, N1005);
and AND3 (N1503, N1489, N604, N388);
buf BUF1 (N1504, N1492);
not NOT1 (N1505, N1503);
xor XOR2 (N1506, N1495, N799);
buf BUF1 (N1507, N1504);
not NOT1 (N1508, N1502);
not NOT1 (N1509, N1494);
xor XOR2 (N1510, N1496, N396);
nand NAND2 (N1511, N1497, N795);
nand NAND3 (N1512, N1510, N659, N1113);
nor NOR2 (N1513, N1507, N452);
nor NOR2 (N1514, N1505, N1197);
and AND4 (N1515, N1481, N771, N863, N131);
buf BUF1 (N1516, N1508);
nand NAND4 (N1517, N1514, N315, N919, N1271);
not NOT1 (N1518, N1515);
or OR3 (N1519, N1509, N874, N1285);
nand NAND3 (N1520, N1506, N1164, N559);
nand NAND4 (N1521, N1519, N612, N897, N826);
nor NOR3 (N1522, N1521, N1418, N343);
nor NOR4 (N1523, N1522, N562, N1328, N778);
xor XOR2 (N1524, N1518, N1181);
buf BUF1 (N1525, N1524);
nor NOR2 (N1526, N1520, N727);
nand NAND2 (N1527, N1512, N1488);
and AND2 (N1528, N1525, N1095);
nand NAND3 (N1529, N1493, N92, N346);
nor NOR3 (N1530, N1523, N1245, N814);
not NOT1 (N1531, N1517);
buf BUF1 (N1532, N1531);
not NOT1 (N1533, N1513);
xor XOR2 (N1534, N1511, N575);
nor NOR2 (N1535, N1529, N274);
and AND4 (N1536, N1501, N706, N1521, N797);
nand NAND4 (N1537, N1516, N562, N1367, N746);
and AND2 (N1538, N1535, N326);
and AND4 (N1539, N1527, N212, N661, N819);
not NOT1 (N1540, N1530);
buf BUF1 (N1541, N1536);
buf BUF1 (N1542, N1541);
buf BUF1 (N1543, N1537);
nand NAND2 (N1544, N1542, N330);
buf BUF1 (N1545, N1540);
xor XOR2 (N1546, N1532, N1509);
and AND2 (N1547, N1538, N1225);
nor NOR2 (N1548, N1534, N384);
not NOT1 (N1549, N1547);
or OR2 (N1550, N1528, N160);
xor XOR2 (N1551, N1548, N114);
not NOT1 (N1552, N1544);
and AND3 (N1553, N1550, N1149, N666);
xor XOR2 (N1554, N1551, N1220);
or OR3 (N1555, N1549, N1258, N1511);
not NOT1 (N1556, N1539);
nand NAND3 (N1557, N1556, N492, N1145);
buf BUF1 (N1558, N1553);
or OR2 (N1559, N1533, N485);
and AND2 (N1560, N1554, N358);
and AND2 (N1561, N1552, N140);
and AND3 (N1562, N1545, N57, N369);
nor NOR2 (N1563, N1555, N761);
and AND2 (N1564, N1562, N864);
nand NAND4 (N1565, N1557, N355, N504, N1444);
xor XOR2 (N1566, N1543, N1163);
buf BUF1 (N1567, N1546);
buf BUF1 (N1568, N1566);
or OR4 (N1569, N1559, N953, N1117, N1160);
nor NOR4 (N1570, N1526, N324, N490, N2);
buf BUF1 (N1571, N1568);
not NOT1 (N1572, N1567);
or OR4 (N1573, N1561, N1288, N305, N374);
and AND4 (N1574, N1558, N1299, N1537, N620);
xor XOR2 (N1575, N1565, N602);
or OR3 (N1576, N1564, N1170, N1265);
nor NOR3 (N1577, N1576, N1054, N735);
nand NAND2 (N1578, N1560, N859);
nand NAND4 (N1579, N1574, N1204, N1139, N403);
xor XOR2 (N1580, N1570, N391);
nor NOR3 (N1581, N1571, N418, N1275);
and AND3 (N1582, N1579, N728, N1017);
and AND3 (N1583, N1581, N753, N647);
nand NAND4 (N1584, N1578, N1435, N524, N474);
xor XOR2 (N1585, N1572, N1005);
and AND3 (N1586, N1583, N356, N691);
nand NAND2 (N1587, N1584, N1583);
or OR3 (N1588, N1563, N1041, N1145);
not NOT1 (N1589, N1575);
not NOT1 (N1590, N1589);
xor XOR2 (N1591, N1577, N833);
not NOT1 (N1592, N1580);
xor XOR2 (N1593, N1592, N1422);
buf BUF1 (N1594, N1586);
and AND4 (N1595, N1594, N665, N1209, N725);
not NOT1 (N1596, N1585);
nand NAND3 (N1597, N1587, N1064, N689);
or OR4 (N1598, N1595, N289, N1260, N1436);
nor NOR3 (N1599, N1590, N811, N287);
or OR3 (N1600, N1596, N1555, N369);
nor NOR3 (N1601, N1600, N1055, N342);
buf BUF1 (N1602, N1591);
buf BUF1 (N1603, N1601);
not NOT1 (N1604, N1569);
nor NOR4 (N1605, N1573, N303, N812, N1185);
buf BUF1 (N1606, N1593);
buf BUF1 (N1607, N1605);
nor NOR2 (N1608, N1606, N220);
buf BUF1 (N1609, N1588);
not NOT1 (N1610, N1602);
nand NAND4 (N1611, N1604, N1266, N1519, N139);
nor NOR3 (N1612, N1608, N505, N192);
xor XOR2 (N1613, N1612, N743);
nand NAND4 (N1614, N1598, N1168, N47, N806);
xor XOR2 (N1615, N1599, N1090);
not NOT1 (N1616, N1582);
xor XOR2 (N1617, N1613, N524);
nand NAND2 (N1618, N1597, N939);
xor XOR2 (N1619, N1616, N79);
buf BUF1 (N1620, N1607);
buf BUF1 (N1621, N1614);
nand NAND3 (N1622, N1611, N883, N1451);
xor XOR2 (N1623, N1610, N978);
buf BUF1 (N1624, N1617);
nor NOR2 (N1625, N1621, N453);
nand NAND2 (N1626, N1625, N1319);
not NOT1 (N1627, N1609);
nand NAND4 (N1628, N1627, N535, N748, N1414);
buf BUF1 (N1629, N1623);
or OR4 (N1630, N1622, N1490, N865, N647);
or OR3 (N1631, N1619, N553, N8);
not NOT1 (N1632, N1624);
nor NOR4 (N1633, N1629, N1036, N1328, N1446);
xor XOR2 (N1634, N1620, N554);
xor XOR2 (N1635, N1603, N1527);
nand NAND2 (N1636, N1630, N1299);
nand NAND2 (N1637, N1633, N589);
nand NAND2 (N1638, N1631, N112);
buf BUF1 (N1639, N1636);
buf BUF1 (N1640, N1639);
and AND3 (N1641, N1638, N332, N1429);
and AND3 (N1642, N1632, N282, N1358);
buf BUF1 (N1643, N1615);
and AND3 (N1644, N1641, N1036, N1617);
buf BUF1 (N1645, N1640);
and AND4 (N1646, N1644, N184, N1207, N1612);
nor NOR3 (N1647, N1645, N1053, N624);
nand NAND2 (N1648, N1634, N560);
buf BUF1 (N1649, N1618);
nor NOR2 (N1650, N1642, N716);
and AND3 (N1651, N1649, N191, N134);
xor XOR2 (N1652, N1648, N648);
buf BUF1 (N1653, N1646);
not NOT1 (N1654, N1653);
nand NAND3 (N1655, N1650, N24, N178);
nor NOR4 (N1656, N1651, N707, N1594, N631);
nand NAND3 (N1657, N1655, N466, N737);
xor XOR2 (N1658, N1656, N809);
or OR3 (N1659, N1643, N1216, N1172);
xor XOR2 (N1660, N1628, N1190);
not NOT1 (N1661, N1659);
not NOT1 (N1662, N1660);
not NOT1 (N1663, N1657);
xor XOR2 (N1664, N1652, N1237);
nor NOR4 (N1665, N1663, N763, N573, N278);
xor XOR2 (N1666, N1664, N1552);
nand NAND4 (N1667, N1661, N1074, N356, N161);
buf BUF1 (N1668, N1654);
not NOT1 (N1669, N1635);
xor XOR2 (N1670, N1662, N580);
or OR3 (N1671, N1670, N347, N1319);
or OR3 (N1672, N1667, N366, N877);
not NOT1 (N1673, N1669);
nor NOR2 (N1674, N1658, N581);
buf BUF1 (N1675, N1665);
nor NOR2 (N1676, N1672, N991);
buf BUF1 (N1677, N1673);
xor XOR2 (N1678, N1671, N573);
not NOT1 (N1679, N1677);
buf BUF1 (N1680, N1668);
buf BUF1 (N1681, N1666);
and AND2 (N1682, N1674, N329);
buf BUF1 (N1683, N1675);
not NOT1 (N1684, N1683);
xor XOR2 (N1685, N1682, N244);
nand NAND3 (N1686, N1637, N849, N1224);
not NOT1 (N1687, N1647);
buf BUF1 (N1688, N1680);
or OR4 (N1689, N1687, N1365, N974, N569);
buf BUF1 (N1690, N1679);
xor XOR2 (N1691, N1689, N1126);
and AND4 (N1692, N1676, N73, N634, N1588);
and AND3 (N1693, N1685, N452, N124);
or OR3 (N1694, N1684, N620, N637);
buf BUF1 (N1695, N1690);
buf BUF1 (N1696, N1678);
not NOT1 (N1697, N1696);
nand NAND3 (N1698, N1681, N1354, N640);
or OR4 (N1699, N1693, N1488, N1186, N266);
nand NAND4 (N1700, N1686, N1282, N1309, N235);
not NOT1 (N1701, N1691);
xor XOR2 (N1702, N1700, N799);
not NOT1 (N1703, N1688);
buf BUF1 (N1704, N1697);
not NOT1 (N1705, N1692);
or OR2 (N1706, N1695, N428);
nand NAND4 (N1707, N1706, N1207, N1384, N470);
and AND4 (N1708, N1707, N1138, N149, N1357);
xor XOR2 (N1709, N1701, N736);
nor NOR4 (N1710, N1694, N108, N450, N645);
nand NAND3 (N1711, N1709, N1579, N215);
not NOT1 (N1712, N1710);
nor NOR2 (N1713, N1699, N1457);
nand NAND4 (N1714, N1705, N649, N883, N568);
nor NOR2 (N1715, N1708, N947);
or OR4 (N1716, N1626, N840, N133, N569);
and AND4 (N1717, N1714, N1052, N273, N1024);
or OR3 (N1718, N1704, N1107, N536);
xor XOR2 (N1719, N1711, N1559);
xor XOR2 (N1720, N1717, N980);
nor NOR3 (N1721, N1718, N590, N1272);
buf BUF1 (N1722, N1702);
and AND4 (N1723, N1698, N211, N178, N1167);
and AND3 (N1724, N1719, N1657, N637);
buf BUF1 (N1725, N1723);
nor NOR3 (N1726, N1716, N996, N1136);
nand NAND2 (N1727, N1725, N251);
buf BUF1 (N1728, N1720);
or OR3 (N1729, N1728, N448, N1682);
buf BUF1 (N1730, N1727);
nor NOR3 (N1731, N1724, N709, N1188);
or OR2 (N1732, N1721, N395);
xor XOR2 (N1733, N1712, N865);
nor NOR3 (N1734, N1715, N738, N1345);
nand NAND3 (N1735, N1726, N720, N388);
nor NOR3 (N1736, N1735, N1472, N1624);
buf BUF1 (N1737, N1703);
buf BUF1 (N1738, N1730);
nand NAND4 (N1739, N1722, N50, N1566, N1416);
nand NAND3 (N1740, N1734, N668, N226);
buf BUF1 (N1741, N1732);
xor XOR2 (N1742, N1731, N1260);
not NOT1 (N1743, N1736);
xor XOR2 (N1744, N1729, N946);
or OR4 (N1745, N1742, N351, N1551, N879);
buf BUF1 (N1746, N1738);
xor XOR2 (N1747, N1740, N876);
nand NAND4 (N1748, N1747, N1274, N1460, N530);
nor NOR4 (N1749, N1744, N1228, N364, N1076);
and AND4 (N1750, N1746, N1476, N1145, N353);
buf BUF1 (N1751, N1737);
nand NAND3 (N1752, N1739, N1079, N1385);
or OR2 (N1753, N1733, N1007);
or OR2 (N1754, N1750, N304);
and AND2 (N1755, N1752, N1439);
xor XOR2 (N1756, N1743, N337);
not NOT1 (N1757, N1713);
nor NOR3 (N1758, N1749, N734, N620);
not NOT1 (N1759, N1745);
nand NAND3 (N1760, N1753, N249, N1072);
and AND2 (N1761, N1759, N506);
not NOT1 (N1762, N1757);
not NOT1 (N1763, N1751);
or OR2 (N1764, N1748, N1019);
or OR3 (N1765, N1762, N288, N464);
or OR4 (N1766, N1764, N143, N1765, N1067);
and AND3 (N1767, N777, N1489, N186);
and AND2 (N1768, N1766, N800);
and AND2 (N1769, N1767, N480);
buf BUF1 (N1770, N1760);
buf BUF1 (N1771, N1770);
and AND4 (N1772, N1771, N1588, N1635, N1658);
nor NOR3 (N1773, N1763, N1635, N1266);
buf BUF1 (N1774, N1741);
xor XOR2 (N1775, N1755, N913);
xor XOR2 (N1776, N1775, N194);
or OR2 (N1777, N1772, N764);
nor NOR2 (N1778, N1754, N151);
nand NAND4 (N1779, N1774, N552, N1549, N251);
nor NOR3 (N1780, N1773, N304, N166);
and AND4 (N1781, N1779, N160, N1564, N1598);
and AND4 (N1782, N1776, N222, N1492, N202);
not NOT1 (N1783, N1756);
buf BUF1 (N1784, N1783);
buf BUF1 (N1785, N1777);
xor XOR2 (N1786, N1782, N1502);
or OR4 (N1787, N1781, N502, N823, N139);
nor NOR3 (N1788, N1780, N580, N870);
and AND3 (N1789, N1769, N656, N1631);
and AND3 (N1790, N1787, N818, N277);
nand NAND4 (N1791, N1786, N1187, N755, N280);
buf BUF1 (N1792, N1758);
xor XOR2 (N1793, N1785, N63);
not NOT1 (N1794, N1793);
not NOT1 (N1795, N1791);
not NOT1 (N1796, N1788);
nor NOR4 (N1797, N1784, N1537, N677, N462);
xor XOR2 (N1798, N1778, N985);
xor XOR2 (N1799, N1789, N828);
nand NAND4 (N1800, N1792, N1124, N724, N1517);
nand NAND3 (N1801, N1799, N1634, N1361);
nor NOR4 (N1802, N1798, N577, N185, N1476);
not NOT1 (N1803, N1800);
nor NOR2 (N1804, N1768, N819);
nand NAND2 (N1805, N1796, N840);
and AND4 (N1806, N1802, N1245, N367, N299);
xor XOR2 (N1807, N1804, N915);
nor NOR4 (N1808, N1797, N1054, N495, N1064);
not NOT1 (N1809, N1761);
xor XOR2 (N1810, N1790, N1317);
not NOT1 (N1811, N1794);
or OR4 (N1812, N1806, N1101, N1588, N1809);
and AND3 (N1813, N1716, N1503, N540);
not NOT1 (N1814, N1795);
and AND3 (N1815, N1811, N813, N1555);
buf BUF1 (N1816, N1813);
and AND3 (N1817, N1807, N1510, N1381);
buf BUF1 (N1818, N1816);
not NOT1 (N1819, N1814);
not NOT1 (N1820, N1810);
not NOT1 (N1821, N1805);
xor XOR2 (N1822, N1819, N1749);
xor XOR2 (N1823, N1812, N1160);
or OR4 (N1824, N1821, N1659, N485, N1070);
nand NAND2 (N1825, N1824, N922);
or OR3 (N1826, N1801, N1647, N1385);
nand NAND4 (N1827, N1803, N1396, N434, N712);
and AND3 (N1828, N1808, N670, N76);
or OR4 (N1829, N1817, N1221, N1219, N1675);
nand NAND4 (N1830, N1827, N502, N196, N1446);
nand NAND3 (N1831, N1818, N332, N1168);
xor XOR2 (N1832, N1822, N1428);
nand NAND2 (N1833, N1820, N654);
not NOT1 (N1834, N1831);
buf BUF1 (N1835, N1834);
not NOT1 (N1836, N1826);
or OR2 (N1837, N1828, N597);
or OR3 (N1838, N1835, N1318, N331);
and AND2 (N1839, N1825, N6);
or OR3 (N1840, N1815, N221, N127);
nor NOR4 (N1841, N1829, N186, N1039, N867);
nand NAND3 (N1842, N1832, N161, N832);
buf BUF1 (N1843, N1840);
buf BUF1 (N1844, N1838);
buf BUF1 (N1845, N1833);
buf BUF1 (N1846, N1841);
not NOT1 (N1847, N1830);
xor XOR2 (N1848, N1823, N1052);
and AND3 (N1849, N1843, N957, N933);
not NOT1 (N1850, N1839);
xor XOR2 (N1851, N1848, N152);
or OR4 (N1852, N1836, N1506, N1821, N126);
nor NOR3 (N1853, N1847, N1712, N791);
and AND3 (N1854, N1842, N1388, N321);
nand NAND2 (N1855, N1844, N1133);
nor NOR3 (N1856, N1855, N1260, N227);
nand NAND4 (N1857, N1845, N473, N838, N276);
not NOT1 (N1858, N1849);
or OR4 (N1859, N1837, N1062, N101, N464);
nand NAND3 (N1860, N1853, N498, N1140);
and AND2 (N1861, N1858, N1832);
and AND2 (N1862, N1861, N716);
nand NAND2 (N1863, N1859, N206);
and AND2 (N1864, N1852, N151);
not NOT1 (N1865, N1860);
and AND2 (N1866, N1854, N952);
xor XOR2 (N1867, N1856, N1167);
buf BUF1 (N1868, N1850);
buf BUF1 (N1869, N1857);
not NOT1 (N1870, N1865);
nand NAND3 (N1871, N1866, N1437, N456);
not NOT1 (N1872, N1862);
and AND4 (N1873, N1864, N1397, N1430, N1234);
nor NOR4 (N1874, N1867, N999, N1802, N101);
not NOT1 (N1875, N1871);
and AND4 (N1876, N1863, N1265, N1102, N962);
or OR2 (N1877, N1874, N12);
and AND4 (N1878, N1851, N1003, N1786, N1154);
buf BUF1 (N1879, N1877);
buf BUF1 (N1880, N1872);
xor XOR2 (N1881, N1868, N1467);
or OR4 (N1882, N1876, N1170, N1039, N118);
nor NOR3 (N1883, N1870, N1680, N1104);
not NOT1 (N1884, N1880);
nand NAND3 (N1885, N1883, N1014, N103);
buf BUF1 (N1886, N1882);
or OR4 (N1887, N1879, N1125, N147, N436);
and AND4 (N1888, N1873, N1457, N1470, N823);
xor XOR2 (N1889, N1875, N1477);
nand NAND4 (N1890, N1869, N643, N1255, N272);
xor XOR2 (N1891, N1884, N43);
nand NAND2 (N1892, N1890, N1523);
nor NOR4 (N1893, N1846, N889, N72, N1447);
not NOT1 (N1894, N1891);
nor NOR2 (N1895, N1878, N1425);
not NOT1 (N1896, N1893);
xor XOR2 (N1897, N1895, N261);
xor XOR2 (N1898, N1881, N464);
xor XOR2 (N1899, N1887, N1062);
not NOT1 (N1900, N1898);
not NOT1 (N1901, N1899);
nor NOR3 (N1902, N1889, N1314, N505);
nor NOR4 (N1903, N1897, N1290, N1115, N337);
or OR3 (N1904, N1901, N319, N1067);
xor XOR2 (N1905, N1903, N1318);
not NOT1 (N1906, N1904);
not NOT1 (N1907, N1905);
and AND2 (N1908, N1892, N1402);
nor NOR4 (N1909, N1900, N1120, N1006, N315);
nor NOR3 (N1910, N1906, N813, N514);
not NOT1 (N1911, N1886);
or OR3 (N1912, N1910, N1378, N1234);
not NOT1 (N1913, N1907);
not NOT1 (N1914, N1896);
and AND4 (N1915, N1913, N43, N525, N1446);
buf BUF1 (N1916, N1914);
not NOT1 (N1917, N1902);
not NOT1 (N1918, N1909);
or OR4 (N1919, N1915, N7, N1216, N344);
nand NAND4 (N1920, N1894, N520, N1791, N1364);
not NOT1 (N1921, N1908);
nor NOR3 (N1922, N1888, N195, N1181);
and AND2 (N1923, N1885, N1303);
nand NAND3 (N1924, N1919, N986, N1224);
buf BUF1 (N1925, N1917);
not NOT1 (N1926, N1921);
buf BUF1 (N1927, N1924);
or OR4 (N1928, N1918, N400, N836, N131);
xor XOR2 (N1929, N1912, N751);
or OR2 (N1930, N1925, N1300);
nor NOR3 (N1931, N1922, N110, N939);
xor XOR2 (N1932, N1929, N673);
nor NOR3 (N1933, N1926, N1521, N1532);
not NOT1 (N1934, N1931);
nor NOR2 (N1935, N1911, N1313);
nor NOR4 (N1936, N1934, N1053, N1032, N1356);
not NOT1 (N1937, N1935);
xor XOR2 (N1938, N1916, N459);
not NOT1 (N1939, N1920);
or OR3 (N1940, N1936, N1692, N564);
xor XOR2 (N1941, N1933, N1762);
nor NOR3 (N1942, N1932, N1154, N676);
nand NAND2 (N1943, N1923, N141);
nor NOR3 (N1944, N1938, N129, N951);
nor NOR2 (N1945, N1944, N278);
not NOT1 (N1946, N1927);
not NOT1 (N1947, N1930);
nand NAND4 (N1948, N1945, N1505, N236, N684);
not NOT1 (N1949, N1948);
not NOT1 (N1950, N1947);
buf BUF1 (N1951, N1940);
xor XOR2 (N1952, N1939, N1017);
not NOT1 (N1953, N1942);
not NOT1 (N1954, N1950);
and AND4 (N1955, N1951, N642, N1170, N9);
nand NAND3 (N1956, N1946, N1675, N1625);
nor NOR4 (N1957, N1955, N683, N1350, N882);
or OR2 (N1958, N1928, N1598);
nand NAND2 (N1959, N1949, N1926);
not NOT1 (N1960, N1959);
xor XOR2 (N1961, N1943, N1425);
buf BUF1 (N1962, N1960);
or OR3 (N1963, N1956, N1228, N424);
buf BUF1 (N1964, N1941);
nor NOR4 (N1965, N1964, N1165, N1206, N55);
nor NOR3 (N1966, N1963, N1895, N988);
nand NAND3 (N1967, N1962, N1201, N208);
not NOT1 (N1968, N1966);
or OR2 (N1969, N1965, N1273);
or OR4 (N1970, N1958, N1262, N1045, N1495);
not NOT1 (N1971, N1952);
or OR4 (N1972, N1967, N943, N717, N180);
and AND2 (N1973, N1971, N1628);
nand NAND3 (N1974, N1970, N1047, N1251);
xor XOR2 (N1975, N1961, N989);
or OR4 (N1976, N1974, N1503, N1455, N1351);
or OR2 (N1977, N1973, N363);
nand NAND4 (N1978, N1972, N1718, N870, N964);
and AND2 (N1979, N1957, N1289);
not NOT1 (N1980, N1976);
nand NAND4 (N1981, N1953, N1407, N596, N42);
xor XOR2 (N1982, N1954, N482);
not NOT1 (N1983, N1969);
xor XOR2 (N1984, N1981, N1963);
and AND2 (N1985, N1977, N1654);
xor XOR2 (N1986, N1985, N336);
buf BUF1 (N1987, N1978);
nor NOR3 (N1988, N1986, N493, N673);
xor XOR2 (N1989, N1983, N1424);
xor XOR2 (N1990, N1968, N1772);
nand NAND3 (N1991, N1989, N1648, N619);
nor NOR4 (N1992, N1987, N161, N1616, N1813);
and AND3 (N1993, N1982, N752, N602);
buf BUF1 (N1994, N1980);
not NOT1 (N1995, N1994);
nand NAND2 (N1996, N1993, N1296);
buf BUF1 (N1997, N1937);
or OR3 (N1998, N1990, N1642, N1764);
not NOT1 (N1999, N1984);
not NOT1 (N2000, N1995);
nor NOR3 (N2001, N1991, N1710, N129);
and AND4 (N2002, N1988, N1043, N1337, N1444);
xor XOR2 (N2003, N1998, N682);
xor XOR2 (N2004, N2000, N115);
xor XOR2 (N2005, N1992, N1720);
xor XOR2 (N2006, N2004, N1615);
buf BUF1 (N2007, N1996);
or OR3 (N2008, N1975, N911, N299);
buf BUF1 (N2009, N2002);
buf BUF1 (N2010, N1979);
buf BUF1 (N2011, N2009);
nor NOR2 (N2012, N2005, N867);
not NOT1 (N2013, N1999);
buf BUF1 (N2014, N2012);
nor NOR3 (N2015, N2003, N1816, N946);
xor XOR2 (N2016, N2001, N1507);
or OR3 (N2017, N2011, N1632, N879);
nand NAND4 (N2018, N1997, N1445, N606, N620);
and AND4 (N2019, N2017, N1098, N153, N32);
nor NOR2 (N2020, N2006, N622);
and AND3 (N2021, N2013, N1313, N1706);
xor XOR2 (N2022, N2016, N429);
nand NAND4 (N2023, N2019, N1853, N1790, N1060);
not NOT1 (N2024, N2007);
buf BUF1 (N2025, N2021);
xor XOR2 (N2026, N2018, N1172);
and AND3 (N2027, N2010, N1117, N312);
not NOT1 (N2028, N2008);
nor NOR2 (N2029, N2028, N1307);
not NOT1 (N2030, N2025);
buf BUF1 (N2031, N2027);
and AND2 (N2032, N2022, N1700);
not NOT1 (N2033, N2014);
buf BUF1 (N2034, N2031);
nor NOR2 (N2035, N2032, N1832);
nor NOR3 (N2036, N2030, N560, N817);
and AND2 (N2037, N2020, N948);
or OR2 (N2038, N2036, N835);
nor NOR3 (N2039, N2015, N1832, N682);
nor NOR2 (N2040, N2034, N1615);
or OR4 (N2041, N2033, N1734, N1573, N202);
nand NAND2 (N2042, N2039, N1054);
or OR4 (N2043, N2042, N1820, N1931, N1226);
nand NAND2 (N2044, N2037, N305);
xor XOR2 (N2045, N2038, N251);
and AND3 (N2046, N2045, N1614, N1495);
xor XOR2 (N2047, N2023, N105);
buf BUF1 (N2048, N2043);
nor NOR4 (N2049, N2044, N223, N453, N907);
and AND4 (N2050, N2029, N147, N1544, N517);
nand NAND2 (N2051, N2040, N1607);
and AND3 (N2052, N2046, N859, N1976);
nor NOR2 (N2053, N2052, N143);
not NOT1 (N2054, N2047);
not NOT1 (N2055, N2049);
not NOT1 (N2056, N2055);
nand NAND3 (N2057, N2051, N1504, N1915);
not NOT1 (N2058, N2048);
buf BUF1 (N2059, N2041);
and AND2 (N2060, N2024, N547);
and AND4 (N2061, N2060, N1181, N914, N88);
or OR2 (N2062, N2061, N1687);
buf BUF1 (N2063, N2026);
not NOT1 (N2064, N2054);
buf BUF1 (N2065, N2053);
xor XOR2 (N2066, N2050, N1672);
and AND2 (N2067, N2065, N390);
buf BUF1 (N2068, N2057);
buf BUF1 (N2069, N2062);
not NOT1 (N2070, N2063);
xor XOR2 (N2071, N2035, N294);
nor NOR2 (N2072, N2056, N129);
not NOT1 (N2073, N2069);
nor NOR2 (N2074, N2073, N985);
nand NAND3 (N2075, N2066, N1981, N444);
and AND3 (N2076, N2068, N377, N824);
or OR3 (N2077, N2058, N1604, N1497);
buf BUF1 (N2078, N2077);
nor NOR3 (N2079, N2074, N181, N812);
buf BUF1 (N2080, N2076);
nor NOR3 (N2081, N2079, N1790, N1557);
nand NAND2 (N2082, N2075, N649);
and AND2 (N2083, N2067, N1920);
buf BUF1 (N2084, N2071);
buf BUF1 (N2085, N2084);
nand NAND4 (N2086, N2080, N187, N2043, N725);
nor NOR2 (N2087, N2083, N1409);
or OR3 (N2088, N2081, N317, N1308);
and AND4 (N2089, N2086, N1749, N1102, N755);
and AND4 (N2090, N2088, N457, N53, N753);
xor XOR2 (N2091, N2064, N1321);
nand NAND2 (N2092, N2078, N788);
or OR2 (N2093, N2090, N1952);
nor NOR4 (N2094, N2093, N299, N51, N306);
not NOT1 (N2095, N2070);
or OR4 (N2096, N2091, N1075, N1075, N1110);
nor NOR4 (N2097, N2059, N1408, N1570, N120);
buf BUF1 (N2098, N2082);
and AND2 (N2099, N2094, N1166);
xor XOR2 (N2100, N2085, N2051);
not NOT1 (N2101, N2095);
nand NAND3 (N2102, N2099, N2038, N166);
and AND2 (N2103, N2087, N1045);
and AND3 (N2104, N2100, N57, N1911);
xor XOR2 (N2105, N2096, N918);
xor XOR2 (N2106, N2104, N462);
not NOT1 (N2107, N2102);
xor XOR2 (N2108, N2072, N1392);
xor XOR2 (N2109, N2103, N213);
or OR3 (N2110, N2097, N358, N1431);
nor NOR3 (N2111, N2105, N1419, N1356);
nand NAND3 (N2112, N2107, N265, N558);
or OR3 (N2113, N2111, N498, N1197);
not NOT1 (N2114, N2108);
nor NOR3 (N2115, N2092, N1393, N172);
nand NAND4 (N2116, N2089, N617, N643, N255);
nor NOR4 (N2117, N2109, N731, N1646, N1624);
or OR4 (N2118, N2114, N723, N1753, N37);
not NOT1 (N2119, N2113);
xor XOR2 (N2120, N2101, N1367);
and AND2 (N2121, N2112, N1795);
not NOT1 (N2122, N2115);
buf BUF1 (N2123, N2106);
nor NOR4 (N2124, N2110, N223, N1196, N308);
or OR4 (N2125, N2116, N457, N1019, N516);
or OR3 (N2126, N2124, N1508, N863);
nor NOR2 (N2127, N2118, N447);
not NOT1 (N2128, N2123);
nand NAND4 (N2129, N2119, N596, N38, N424);
not NOT1 (N2130, N2126);
nand NAND2 (N2131, N2098, N785);
nand NAND2 (N2132, N2125, N1483);
nor NOR3 (N2133, N2130, N821, N668);
not NOT1 (N2134, N2117);
nor NOR3 (N2135, N2122, N767, N1170);
or OR4 (N2136, N2129, N498, N1389, N1425);
or OR4 (N2137, N2131, N1958, N1486, N153);
not NOT1 (N2138, N2120);
nand NAND2 (N2139, N2135, N941);
nor NOR4 (N2140, N2127, N808, N1443, N1894);
nor NOR4 (N2141, N2133, N1207, N801, N888);
not NOT1 (N2142, N2139);
xor XOR2 (N2143, N2141, N480);
buf BUF1 (N2144, N2143);
not NOT1 (N2145, N2140);
not NOT1 (N2146, N2137);
buf BUF1 (N2147, N2132);
buf BUF1 (N2148, N2142);
nand NAND2 (N2149, N2134, N789);
not NOT1 (N2150, N2144);
or OR2 (N2151, N2148, N1003);
xor XOR2 (N2152, N2146, N1428);
or OR4 (N2153, N2151, N2084, N1386, N147);
not NOT1 (N2154, N2149);
nor NOR4 (N2155, N2153, N794, N1224, N1723);
and AND4 (N2156, N2128, N1921, N1953, N926);
or OR4 (N2157, N2152, N2014, N1235, N2064);
not NOT1 (N2158, N2147);
xor XOR2 (N2159, N2145, N1001);
nor NOR4 (N2160, N2159, N754, N117, N1180);
and AND3 (N2161, N2154, N1907, N148);
xor XOR2 (N2162, N2160, N207);
xor XOR2 (N2163, N2161, N1790);
not NOT1 (N2164, N2162);
not NOT1 (N2165, N2136);
nand NAND4 (N2166, N2138, N660, N1055, N468);
buf BUF1 (N2167, N2164);
buf BUF1 (N2168, N2167);
not NOT1 (N2169, N2155);
xor XOR2 (N2170, N2166, N442);
and AND4 (N2171, N2165, N929, N196, N291);
buf BUF1 (N2172, N2168);
not NOT1 (N2173, N2169);
not NOT1 (N2174, N2163);
not NOT1 (N2175, N2158);
and AND2 (N2176, N2150, N1050);
or OR4 (N2177, N2170, N761, N949, N594);
not NOT1 (N2178, N2172);
and AND3 (N2179, N2176, N1364, N1856);
nor NOR3 (N2180, N2178, N36, N1373);
and AND3 (N2181, N2180, N1851, N1664);
or OR2 (N2182, N2179, N1412);
not NOT1 (N2183, N2174);
nor NOR4 (N2184, N2173, N1617, N1475, N2070);
not NOT1 (N2185, N2182);
xor XOR2 (N2186, N2181, N948);
nor NOR3 (N2187, N2175, N373, N2103);
and AND2 (N2188, N2183, N670);
nand NAND2 (N2189, N2121, N137);
nand NAND2 (N2190, N2157, N1556);
not NOT1 (N2191, N2187);
not NOT1 (N2192, N2190);
xor XOR2 (N2193, N2184, N1309);
xor XOR2 (N2194, N2156, N1456);
buf BUF1 (N2195, N2185);
nor NOR3 (N2196, N2189, N2047, N271);
buf BUF1 (N2197, N2196);
buf BUF1 (N2198, N2195);
and AND2 (N2199, N2171, N1112);
xor XOR2 (N2200, N2177, N44);
xor XOR2 (N2201, N2186, N1941);
or OR3 (N2202, N2193, N441, N1297);
buf BUF1 (N2203, N2192);
or OR2 (N2204, N2202, N500);
buf BUF1 (N2205, N2197);
nor NOR2 (N2206, N2201, N1592);
and AND2 (N2207, N2206, N707);
nand NAND3 (N2208, N2200, N953, N1512);
not NOT1 (N2209, N2199);
or OR4 (N2210, N2205, N1011, N1371, N1922);
nor NOR4 (N2211, N2207, N811, N1085, N520);
xor XOR2 (N2212, N2210, N1105);
buf BUF1 (N2213, N2211);
and AND4 (N2214, N2212, N700, N1237, N231);
xor XOR2 (N2215, N2194, N1676);
xor XOR2 (N2216, N2203, N1589);
nand NAND2 (N2217, N2214, N978);
nor NOR4 (N2218, N2204, N985, N1720, N1954);
nand NAND2 (N2219, N2213, N1754);
or OR3 (N2220, N2188, N934, N2173);
and AND4 (N2221, N2217, N699, N2166, N56);
nor NOR3 (N2222, N2198, N907, N1806);
nor NOR3 (N2223, N2221, N345, N381);
xor XOR2 (N2224, N2208, N1738);
xor XOR2 (N2225, N2216, N1194);
and AND4 (N2226, N2219, N1776, N1079, N1017);
and AND2 (N2227, N2220, N585);
xor XOR2 (N2228, N2215, N469);
and AND3 (N2229, N2209, N1733, N186);
not NOT1 (N2230, N2191);
nand NAND4 (N2231, N2224, N1977, N2004, N92);
xor XOR2 (N2232, N2229, N1098);
nor NOR3 (N2233, N2222, N1260, N618);
nor NOR4 (N2234, N2233, N1207, N520, N1226);
or OR2 (N2235, N2225, N1310);
buf BUF1 (N2236, N2230);
or OR2 (N2237, N2227, N1099);
not NOT1 (N2238, N2226);
and AND2 (N2239, N2223, N626);
or OR4 (N2240, N2239, N1033, N2233, N432);
nor NOR4 (N2241, N2236, N1781, N309, N273);
or OR4 (N2242, N2241, N2040, N1132, N2010);
buf BUF1 (N2243, N2232);
buf BUF1 (N2244, N2234);
or OR4 (N2245, N2244, N1185, N356, N1138);
nor NOR2 (N2246, N2245, N422);
nand NAND2 (N2247, N2238, N778);
xor XOR2 (N2248, N2243, N1621);
and AND3 (N2249, N2231, N42, N1752);
nor NOR2 (N2250, N2240, N634);
xor XOR2 (N2251, N2237, N534);
and AND4 (N2252, N2251, N665, N1186, N2047);
xor XOR2 (N2253, N2246, N2205);
not NOT1 (N2254, N2242);
not NOT1 (N2255, N2235);
or OR3 (N2256, N2248, N1675, N2106);
not NOT1 (N2257, N2247);
and AND2 (N2258, N2253, N2036);
or OR2 (N2259, N2252, N305);
nand NAND3 (N2260, N2257, N1748, N1585);
nor NOR3 (N2261, N2249, N1244, N1103);
buf BUF1 (N2262, N2261);
xor XOR2 (N2263, N2262, N66);
buf BUF1 (N2264, N2255);
nor NOR3 (N2265, N2263, N544, N2000);
nor NOR3 (N2266, N2254, N43, N1281);
and AND3 (N2267, N2260, N1588, N1906);
buf BUF1 (N2268, N2266);
or OR3 (N2269, N2267, N1925, N31);
xor XOR2 (N2270, N2264, N897);
or OR2 (N2271, N2228, N45);
xor XOR2 (N2272, N2265, N2174);
nor NOR4 (N2273, N2270, N1914, N302, N585);
or OR4 (N2274, N2256, N146, N2216, N1039);
nand NAND2 (N2275, N2271, N146);
or OR2 (N2276, N2268, N2178);
or OR4 (N2277, N2218, N2204, N1557, N1336);
and AND2 (N2278, N2269, N2061);
buf BUF1 (N2279, N2272);
nor NOR2 (N2280, N2277, N2127);
buf BUF1 (N2281, N2280);
nand NAND2 (N2282, N2274, N325);
nor NOR2 (N2283, N2275, N677);
not NOT1 (N2284, N2258);
nand NAND3 (N2285, N2281, N1530, N867);
nor NOR2 (N2286, N2278, N33);
and AND3 (N2287, N2283, N491, N4);
xor XOR2 (N2288, N2273, N736);
buf BUF1 (N2289, N2276);
xor XOR2 (N2290, N2282, N476);
nor NOR3 (N2291, N2288, N1997, N1285);
or OR2 (N2292, N2289, N2203);
and AND3 (N2293, N2287, N1996, N2285);
nand NAND4 (N2294, N899, N371, N1452, N985);
xor XOR2 (N2295, N2291, N1099);
not NOT1 (N2296, N2293);
not NOT1 (N2297, N2292);
buf BUF1 (N2298, N2259);
buf BUF1 (N2299, N2290);
nor NOR4 (N2300, N2295, N592, N1096, N148);
not NOT1 (N2301, N2284);
nand NAND3 (N2302, N2286, N749, N378);
nor NOR2 (N2303, N2297, N2051);
xor XOR2 (N2304, N2302, N2071);
nand NAND4 (N2305, N2303, N978, N1, N1170);
not NOT1 (N2306, N2300);
not NOT1 (N2307, N2296);
nand NAND3 (N2308, N2250, N1434, N2291);
xor XOR2 (N2309, N2306, N688);
and AND2 (N2310, N2307, N938);
or OR2 (N2311, N2279, N497);
nand NAND2 (N2312, N2304, N885);
buf BUF1 (N2313, N2299);
nor NOR4 (N2314, N2313, N803, N1418, N2079);
nor NOR4 (N2315, N2298, N2083, N1012, N1300);
xor XOR2 (N2316, N2305, N1757);
and AND2 (N2317, N2315, N1382);
nor NOR2 (N2318, N2308, N1787);
buf BUF1 (N2319, N2311);
not NOT1 (N2320, N2310);
nor NOR4 (N2321, N2314, N2271, N1787, N154);
and AND4 (N2322, N2309, N1318, N967, N2042);
not NOT1 (N2323, N2318);
buf BUF1 (N2324, N2301);
and AND4 (N2325, N2321, N2194, N1154, N1410);
nor NOR2 (N2326, N2312, N1156);
nand NAND2 (N2327, N2317, N1188);
buf BUF1 (N2328, N2324);
nor NOR3 (N2329, N2328, N664, N939);
or OR2 (N2330, N2319, N1536);
or OR3 (N2331, N2327, N2184, N2031);
nand NAND4 (N2332, N2320, N467, N219, N2260);
buf BUF1 (N2333, N2330);
buf BUF1 (N2334, N2323);
nand NAND4 (N2335, N2332, N2148, N47, N726);
buf BUF1 (N2336, N2334);
nor NOR2 (N2337, N2333, N1703);
not NOT1 (N2338, N2294);
not NOT1 (N2339, N2331);
buf BUF1 (N2340, N2339);
or OR4 (N2341, N2322, N154, N2056, N608);
not NOT1 (N2342, N2338);
not NOT1 (N2343, N2340);
nand NAND2 (N2344, N2342, N956);
and AND4 (N2345, N2329, N61, N838, N2031);
not NOT1 (N2346, N2345);
not NOT1 (N2347, N2343);
xor XOR2 (N2348, N2337, N373);
xor XOR2 (N2349, N2341, N590);
or OR3 (N2350, N2326, N1765, N1726);
nand NAND3 (N2351, N2344, N548, N1805);
and AND2 (N2352, N2349, N2093);
nand NAND3 (N2353, N2335, N2330, N442);
not NOT1 (N2354, N2346);
not NOT1 (N2355, N2350);
buf BUF1 (N2356, N2355);
or OR4 (N2357, N2316, N1036, N1990, N1884);
nor NOR2 (N2358, N2348, N1581);
nand NAND4 (N2359, N2351, N708, N1320, N1906);
xor XOR2 (N2360, N2354, N1747);
and AND4 (N2361, N2357, N131, N990, N1669);
and AND4 (N2362, N2353, N1102, N487, N525);
not NOT1 (N2363, N2358);
or OR3 (N2364, N2347, N1180, N326);
buf BUF1 (N2365, N2360);
not NOT1 (N2366, N2362);
or OR4 (N2367, N2325, N304, N144, N1225);
buf BUF1 (N2368, N2363);
or OR3 (N2369, N2356, N383, N2283);
xor XOR2 (N2370, N2359, N729);
buf BUF1 (N2371, N2366);
and AND2 (N2372, N2371, N504);
nor NOR4 (N2373, N2365, N2049, N431, N1438);
nand NAND3 (N2374, N2367, N1654, N1363);
or OR3 (N2375, N2368, N2172, N1385);
not NOT1 (N2376, N2373);
nand NAND4 (N2377, N2370, N195, N1091, N71);
not NOT1 (N2378, N2364);
or OR3 (N2379, N2375, N1007, N1170);
nor NOR3 (N2380, N2374, N2034, N999);
or OR4 (N2381, N2378, N1259, N2366, N2184);
nor NOR2 (N2382, N2336, N2183);
nor NOR2 (N2383, N2372, N532);
nand NAND3 (N2384, N2379, N1101, N1934);
buf BUF1 (N2385, N2381);
xor XOR2 (N2386, N2361, N589);
and AND2 (N2387, N2382, N632);
xor XOR2 (N2388, N2384, N722);
not NOT1 (N2389, N2369);
nor NOR2 (N2390, N2385, N817);
and AND3 (N2391, N2383, N1319, N2098);
xor XOR2 (N2392, N2376, N1640);
nor NOR4 (N2393, N2387, N847, N815, N606);
xor XOR2 (N2394, N2377, N863);
not NOT1 (N2395, N2394);
nor NOR4 (N2396, N2389, N1978, N2138, N1257);
or OR2 (N2397, N2392, N15);
not NOT1 (N2398, N2380);
nand NAND2 (N2399, N2396, N1708);
or OR3 (N2400, N2395, N1926, N68);
nor NOR3 (N2401, N2399, N2148, N1202);
and AND2 (N2402, N2391, N1546);
nor NOR4 (N2403, N2388, N1355, N139, N455);
not NOT1 (N2404, N2402);
xor XOR2 (N2405, N2386, N193);
xor XOR2 (N2406, N2401, N2160);
buf BUF1 (N2407, N2398);
buf BUF1 (N2408, N2404);
or OR2 (N2409, N2352, N1138);
nand NAND3 (N2410, N2408, N1706, N1673);
xor XOR2 (N2411, N2390, N767);
not NOT1 (N2412, N2393);
buf BUF1 (N2413, N2406);
buf BUF1 (N2414, N2400);
nor NOR2 (N2415, N2409, N1877);
xor XOR2 (N2416, N2411, N2072);
xor XOR2 (N2417, N2415, N900);
and AND4 (N2418, N2397, N180, N392, N1746);
nand NAND3 (N2419, N2410, N1294, N1091);
and AND2 (N2420, N2414, N838);
nor NOR3 (N2421, N2417, N1462, N1917);
nor NOR3 (N2422, N2416, N1032, N1053);
and AND3 (N2423, N2405, N1621, N1122);
nor NOR4 (N2424, N2421, N1733, N1801, N454);
and AND4 (N2425, N2420, N2111, N1969, N1670);
or OR2 (N2426, N2407, N768);
or OR4 (N2427, N2426, N51, N2324, N2275);
nand NAND3 (N2428, N2423, N478, N2164);
or OR3 (N2429, N2413, N2291, N42);
not NOT1 (N2430, N2422);
buf BUF1 (N2431, N2403);
nand NAND3 (N2432, N2412, N2053, N1775);
xor XOR2 (N2433, N2427, N101);
xor XOR2 (N2434, N2432, N773);
buf BUF1 (N2435, N2430);
buf BUF1 (N2436, N2425);
not NOT1 (N2437, N2429);
or OR4 (N2438, N2419, N2247, N1448, N796);
buf BUF1 (N2439, N2434);
or OR2 (N2440, N2437, N221);
and AND3 (N2441, N2438, N2061, N1946);
and AND4 (N2442, N2418, N228, N222, N208);
nor NOR4 (N2443, N2436, N1901, N241, N2112);
and AND4 (N2444, N2433, N2220, N601, N622);
and AND2 (N2445, N2435, N2296);
nand NAND2 (N2446, N2424, N764);
buf BUF1 (N2447, N2440);
xor XOR2 (N2448, N2442, N150);
nor NOR3 (N2449, N2428, N586, N2442);
buf BUF1 (N2450, N2444);
and AND4 (N2451, N2449, N2227, N742, N516);
buf BUF1 (N2452, N2441);
nor NOR2 (N2453, N2448, N2026);
not NOT1 (N2454, N2443);
nor NOR4 (N2455, N2452, N1727, N596, N2264);
or OR4 (N2456, N2447, N601, N1687, N1174);
nand NAND3 (N2457, N2455, N431, N1459);
or OR2 (N2458, N2446, N1759);
or OR3 (N2459, N2453, N374, N1685);
or OR2 (N2460, N2450, N1423);
or OR4 (N2461, N2458, N730, N1139, N523);
xor XOR2 (N2462, N2457, N2224);
not NOT1 (N2463, N2431);
and AND4 (N2464, N2459, N837, N633, N2101);
and AND4 (N2465, N2461, N2027, N2425, N829);
xor XOR2 (N2466, N2460, N1437);
or OR2 (N2467, N2451, N383);
or OR2 (N2468, N2454, N1642);
nand NAND3 (N2469, N2467, N317, N1063);
xor XOR2 (N2470, N2462, N1002);
not NOT1 (N2471, N2464);
nor NOR2 (N2472, N2456, N2471);
or OR3 (N2473, N1959, N2395, N401);
buf BUF1 (N2474, N2465);
nor NOR2 (N2475, N2463, N2038);
and AND4 (N2476, N2474, N2386, N2191, N1233);
xor XOR2 (N2477, N2470, N1922);
xor XOR2 (N2478, N2466, N1988);
buf BUF1 (N2479, N2473);
nor NOR3 (N2480, N2469, N742, N2450);
not NOT1 (N2481, N2472);
nor NOR4 (N2482, N2468, N1082, N1705, N1737);
nand NAND4 (N2483, N2482, N2121, N2208, N1865);
not NOT1 (N2484, N2477);
not NOT1 (N2485, N2475);
not NOT1 (N2486, N2485);
or OR2 (N2487, N2483, N1108);
xor XOR2 (N2488, N2478, N1417);
buf BUF1 (N2489, N2480);
xor XOR2 (N2490, N2484, N940);
nand NAND3 (N2491, N2490, N749, N1147);
nand NAND4 (N2492, N2487, N1742, N1256, N2307);
not NOT1 (N2493, N2491);
or OR3 (N2494, N2481, N2316, N509);
buf BUF1 (N2495, N2445);
and AND3 (N2496, N2486, N1573, N2116);
and AND2 (N2497, N2494, N430);
buf BUF1 (N2498, N2489);
xor XOR2 (N2499, N2492, N2287);
not NOT1 (N2500, N2498);
nor NOR2 (N2501, N2497, N231);
or OR4 (N2502, N2500, N134, N1150, N578);
nand NAND4 (N2503, N2439, N1419, N2270, N2488);
not NOT1 (N2504, N2226);
and AND2 (N2505, N2499, N1552);
and AND3 (N2506, N2479, N1279, N1710);
nand NAND2 (N2507, N2496, N2303);
or OR4 (N2508, N2493, N2010, N413, N1008);
or OR4 (N2509, N2501, N1532, N1889, N1381);
not NOT1 (N2510, N2506);
or OR2 (N2511, N2476, N414);
nand NAND3 (N2512, N2503, N1951, N374);
nand NAND3 (N2513, N2511, N2147, N1356);
and AND4 (N2514, N2495, N565, N253, N1572);
nor NOR3 (N2515, N2509, N552, N1110);
and AND2 (N2516, N2507, N1425);
xor XOR2 (N2517, N2515, N2323);
nor NOR3 (N2518, N2516, N437, N357);
xor XOR2 (N2519, N2518, N980);
xor XOR2 (N2520, N2510, N1057);
buf BUF1 (N2521, N2513);
nor NOR3 (N2522, N2517, N599, N1375);
not NOT1 (N2523, N2512);
or OR4 (N2524, N2523, N1849, N2281, N136);
and AND3 (N2525, N2502, N1115, N2076);
buf BUF1 (N2526, N2504);
or OR4 (N2527, N2505, N1953, N1259, N2378);
buf BUF1 (N2528, N2522);
nor NOR2 (N2529, N2526, N2272);
or OR4 (N2530, N2521, N1402, N2420, N1673);
nand NAND2 (N2531, N2514, N1370);
xor XOR2 (N2532, N2528, N1727);
and AND2 (N2533, N2527, N151);
nand NAND3 (N2534, N2525, N2223, N1499);
and AND3 (N2535, N2508, N2402, N841);
xor XOR2 (N2536, N2529, N1678);
nor NOR4 (N2537, N2533, N2064, N990, N475);
buf BUF1 (N2538, N2524);
nand NAND4 (N2539, N2519, N853, N2275, N1660);
xor XOR2 (N2540, N2532, N680);
nor NOR4 (N2541, N2540, N1376, N778, N359);
not NOT1 (N2542, N2535);
nand NAND4 (N2543, N2534, N518, N396, N457);
nor NOR2 (N2544, N2542, N824);
xor XOR2 (N2545, N2539, N298);
xor XOR2 (N2546, N2520, N1463);
or OR4 (N2547, N2543, N2391, N2541, N1014);
xor XOR2 (N2548, N1605, N152);
nor NOR2 (N2549, N2538, N1253);
not NOT1 (N2550, N2549);
xor XOR2 (N2551, N2545, N759);
xor XOR2 (N2552, N2531, N2228);
nor NOR3 (N2553, N2551, N340, N913);
and AND3 (N2554, N2548, N100, N2020);
buf BUF1 (N2555, N2554);
and AND4 (N2556, N2550, N1200, N1261, N1272);
and AND3 (N2557, N2553, N2395, N203);
or OR3 (N2558, N2544, N1168, N522);
or OR4 (N2559, N2546, N297, N1689, N2246);
nand NAND3 (N2560, N2547, N1691, N1431);
and AND3 (N2561, N2537, N319, N149);
and AND2 (N2562, N2556, N1546);
not NOT1 (N2563, N2559);
xor XOR2 (N2564, N2561, N2524);
xor XOR2 (N2565, N2562, N1418);
and AND3 (N2566, N2564, N1336, N1603);
nor NOR4 (N2567, N2563, N1929, N813, N962);
and AND2 (N2568, N2565, N1965);
xor XOR2 (N2569, N2560, N412);
nand NAND2 (N2570, N2557, N1842);
nand NAND2 (N2571, N2558, N1490);
nand NAND4 (N2572, N2552, N1293, N2555, N1106);
buf BUF1 (N2573, N2103);
not NOT1 (N2574, N2570);
nand NAND3 (N2575, N2567, N681, N1159);
nand NAND3 (N2576, N2575, N1264, N682);
buf BUF1 (N2577, N2530);
not NOT1 (N2578, N2571);
or OR3 (N2579, N2569, N1079, N1300);
or OR4 (N2580, N2577, N1481, N1596, N1557);
xor XOR2 (N2581, N2566, N1775);
not NOT1 (N2582, N2536);
nor NOR2 (N2583, N2581, N2224);
xor XOR2 (N2584, N2578, N2400);
nor NOR2 (N2585, N2576, N1425);
nand NAND2 (N2586, N2583, N811);
nor NOR4 (N2587, N2573, N723, N825, N784);
nor NOR3 (N2588, N2580, N307, N706);
nand NAND3 (N2589, N2587, N1959, N946);
nand NAND2 (N2590, N2586, N201);
or OR3 (N2591, N2590, N453, N855);
xor XOR2 (N2592, N2582, N1252);
and AND4 (N2593, N2591, N420, N1786, N604);
buf BUF1 (N2594, N2574);
nand NAND2 (N2595, N2589, N1692);
or OR3 (N2596, N2568, N825, N726);
or OR4 (N2597, N2594, N1606, N1443, N1091);
nor NOR3 (N2598, N2585, N1005, N1143);
and AND2 (N2599, N2596, N1298);
and AND3 (N2600, N2572, N824, N2493);
buf BUF1 (N2601, N2597);
nand NAND3 (N2602, N2599, N1684, N1394);
or OR4 (N2603, N2592, N926, N1038, N33);
xor XOR2 (N2604, N2603, N656);
nand NAND4 (N2605, N2598, N2302, N1797, N1636);
not NOT1 (N2606, N2601);
and AND3 (N2607, N2606, N1128, N1343);
or OR4 (N2608, N2593, N458, N490, N648);
nand NAND2 (N2609, N2595, N869);
or OR2 (N2610, N2609, N636);
buf BUF1 (N2611, N2607);
and AND3 (N2612, N2602, N2445, N2031);
buf BUF1 (N2613, N2579);
nor NOR4 (N2614, N2588, N1224, N1425, N476);
xor XOR2 (N2615, N2608, N921);
not NOT1 (N2616, N2604);
or OR4 (N2617, N2614, N126, N23, N668);
buf BUF1 (N2618, N2613);
nor NOR4 (N2619, N2610, N255, N1869, N1246);
buf BUF1 (N2620, N2617);
or OR3 (N2621, N2605, N2138, N1774);
nand NAND4 (N2622, N2616, N1110, N580, N1184);
xor XOR2 (N2623, N2584, N1551);
not NOT1 (N2624, N2622);
nor NOR3 (N2625, N2600, N2442, N535);
nand NAND4 (N2626, N2620, N2078, N190, N213);
xor XOR2 (N2627, N2624, N520);
and AND4 (N2628, N2627, N673, N2038, N1150);
buf BUF1 (N2629, N2619);
nor NOR2 (N2630, N2621, N1529);
buf BUF1 (N2631, N2612);
not NOT1 (N2632, N2629);
and AND3 (N2633, N2611, N2028, N1167);
nor NOR4 (N2634, N2632, N1039, N2542, N451);
buf BUF1 (N2635, N2630);
nor NOR2 (N2636, N2626, N2572);
not NOT1 (N2637, N2615);
nand NAND3 (N2638, N2623, N430, N816);
xor XOR2 (N2639, N2618, N1734);
xor XOR2 (N2640, N2639, N1660);
nor NOR2 (N2641, N2634, N1878);
buf BUF1 (N2642, N2641);
xor XOR2 (N2643, N2636, N2030);
nand NAND4 (N2644, N2625, N1558, N1857, N2611);
nand NAND4 (N2645, N2633, N493, N1578, N1156);
nor NOR3 (N2646, N2631, N642, N11);
nand NAND2 (N2647, N2643, N1425);
nand NAND3 (N2648, N2635, N150, N80);
xor XOR2 (N2649, N2648, N1027);
not NOT1 (N2650, N2638);
xor XOR2 (N2651, N2645, N1751);
not NOT1 (N2652, N2646);
nor NOR2 (N2653, N2651, N407);
and AND3 (N2654, N2653, N2649, N1243);
and AND4 (N2655, N2307, N70, N2464, N61);
nor NOR2 (N2656, N2628, N1693);
nor NOR3 (N2657, N2650, N1342, N2348);
not NOT1 (N2658, N2647);
xor XOR2 (N2659, N2644, N1392);
xor XOR2 (N2660, N2658, N2390);
and AND3 (N2661, N2654, N1740, N2453);
buf BUF1 (N2662, N2661);
xor XOR2 (N2663, N2656, N2542);
or OR2 (N2664, N2652, N2064);
xor XOR2 (N2665, N2662, N981);
or OR4 (N2666, N2660, N1391, N2360, N2464);
nor NOR4 (N2667, N2659, N563, N1548, N426);
and AND4 (N2668, N2665, N2482, N1416, N2090);
nor NOR4 (N2669, N2640, N268, N1534, N1477);
not NOT1 (N2670, N2655);
not NOT1 (N2671, N2637);
buf BUF1 (N2672, N2669);
or OR3 (N2673, N2671, N2265, N940);
nor NOR4 (N2674, N2673, N2035, N1566, N2026);
or OR3 (N2675, N2672, N75, N1879);
or OR4 (N2676, N2674, N1777, N2512, N2143);
nor NOR2 (N2677, N2668, N1310);
and AND2 (N2678, N2663, N2055);
not NOT1 (N2679, N2666);
xor XOR2 (N2680, N2657, N1539);
buf BUF1 (N2681, N2679);
nor NOR4 (N2682, N2681, N873, N2115, N1306);
not NOT1 (N2683, N2667);
nor NOR3 (N2684, N2680, N1117, N1253);
buf BUF1 (N2685, N2683);
not NOT1 (N2686, N2676);
buf BUF1 (N2687, N2642);
and AND4 (N2688, N2664, N558, N761, N206);
or OR2 (N2689, N2678, N1637);
or OR3 (N2690, N2670, N1340, N527);
buf BUF1 (N2691, N2689);
and AND4 (N2692, N2690, N942, N164, N2428);
not NOT1 (N2693, N2692);
not NOT1 (N2694, N2687);
nand NAND4 (N2695, N2686, N1395, N1709, N1762);
xor XOR2 (N2696, N2675, N432);
not NOT1 (N2697, N2694);
not NOT1 (N2698, N2684);
and AND2 (N2699, N2698, N451);
nand NAND2 (N2700, N2693, N2520);
nor NOR3 (N2701, N2685, N2567, N2451);
xor XOR2 (N2702, N2688, N2607);
xor XOR2 (N2703, N2677, N733);
nand NAND2 (N2704, N2697, N254);
not NOT1 (N2705, N2700);
xor XOR2 (N2706, N2704, N1601);
nor NOR3 (N2707, N2699, N1819, N862);
not NOT1 (N2708, N2703);
xor XOR2 (N2709, N2696, N473);
buf BUF1 (N2710, N2708);
nand NAND4 (N2711, N2710, N432, N2373, N2619);
nand NAND3 (N2712, N2691, N2699, N1735);
or OR3 (N2713, N2682, N2110, N1935);
buf BUF1 (N2714, N2713);
not NOT1 (N2715, N2714);
xor XOR2 (N2716, N2707, N1117);
buf BUF1 (N2717, N2706);
and AND4 (N2718, N2702, N867, N1564, N324);
or OR3 (N2719, N2701, N1707, N2311);
xor XOR2 (N2720, N2718, N285);
not NOT1 (N2721, N2709);
not NOT1 (N2722, N2695);
nor NOR2 (N2723, N2722, N2639);
buf BUF1 (N2724, N2712);
xor XOR2 (N2725, N2716, N1952);
nor NOR4 (N2726, N2717, N175, N1951, N1540);
or OR2 (N2727, N2719, N1887);
nand NAND4 (N2728, N2715, N974, N265, N1222);
xor XOR2 (N2729, N2723, N375);
or OR4 (N2730, N2711, N1832, N2424, N2285);
not NOT1 (N2731, N2705);
not NOT1 (N2732, N2731);
nor NOR2 (N2733, N2728, N2363);
xor XOR2 (N2734, N2726, N2224);
not NOT1 (N2735, N2734);
or OR2 (N2736, N2730, N2483);
nand NAND2 (N2737, N2729, N1480);
and AND4 (N2738, N2735, N2032, N2505, N2179);
and AND3 (N2739, N2727, N1391, N2569);
not NOT1 (N2740, N2721);
nand NAND2 (N2741, N2720, N163);
nor NOR4 (N2742, N2738, N2648, N1012, N2470);
nor NOR3 (N2743, N2737, N1107, N621);
and AND3 (N2744, N2724, N515, N1039);
nand NAND3 (N2745, N2725, N391, N2619);
buf BUF1 (N2746, N2745);
nand NAND4 (N2747, N2743, N2517, N2048, N2683);
and AND4 (N2748, N2744, N2261, N368, N505);
not NOT1 (N2749, N2736);
xor XOR2 (N2750, N2741, N2291);
buf BUF1 (N2751, N2742);
or OR3 (N2752, N2747, N1385, N2446);
buf BUF1 (N2753, N2751);
nor NOR2 (N2754, N2750, N2577);
not NOT1 (N2755, N2748);
or OR4 (N2756, N2749, N2650, N2609, N2426);
nor NOR2 (N2757, N2733, N1175);
not NOT1 (N2758, N2732);
or OR2 (N2759, N2757, N940);
not NOT1 (N2760, N2753);
and AND4 (N2761, N2739, N2662, N2431, N203);
nor NOR4 (N2762, N2746, N2739, N1955, N1528);
nand NAND2 (N2763, N2752, N367);
buf BUF1 (N2764, N2759);
nor NOR4 (N2765, N2761, N2383, N2497, N2020);
not NOT1 (N2766, N2756);
nor NOR3 (N2767, N2766, N2190, N2138);
and AND4 (N2768, N2754, N480, N740, N2265);
not NOT1 (N2769, N2764);
not NOT1 (N2770, N2768);
or OR2 (N2771, N2760, N1529);
xor XOR2 (N2772, N2740, N1080);
xor XOR2 (N2773, N2765, N1485);
not NOT1 (N2774, N2771);
xor XOR2 (N2775, N2763, N858);
buf BUF1 (N2776, N2769);
nand NAND3 (N2777, N2755, N1271, N929);
nand NAND2 (N2778, N2770, N798);
or OR2 (N2779, N2775, N1301);
xor XOR2 (N2780, N2777, N2139);
nand NAND3 (N2781, N2772, N389, N2715);
and AND3 (N2782, N2767, N1141, N234);
nor NOR3 (N2783, N2778, N1290, N2583);
xor XOR2 (N2784, N2781, N2693);
and AND2 (N2785, N2779, N2030);
buf BUF1 (N2786, N2776);
nor NOR4 (N2787, N2785, N2550, N1566, N1114);
xor XOR2 (N2788, N2773, N811);
buf BUF1 (N2789, N2782);
nor NOR4 (N2790, N2786, N1873, N1854, N195);
nor NOR3 (N2791, N2762, N2753, N2505);
not NOT1 (N2792, N2788);
or OR4 (N2793, N2758, N977, N935, N2493);
nand NAND3 (N2794, N2787, N1773, N2584);
nand NAND4 (N2795, N2794, N2043, N2184, N355);
xor XOR2 (N2796, N2784, N2531);
or OR2 (N2797, N2780, N340);
xor XOR2 (N2798, N2793, N773);
xor XOR2 (N2799, N2798, N2236);
or OR2 (N2800, N2791, N1728);
nor NOR4 (N2801, N2783, N1091, N1218, N1878);
and AND4 (N2802, N2795, N1513, N1909, N2677);
nor NOR4 (N2803, N2789, N1263, N1994, N2654);
not NOT1 (N2804, N2800);
and AND2 (N2805, N2792, N217);
xor XOR2 (N2806, N2803, N220);
xor XOR2 (N2807, N2804, N1153);
or OR3 (N2808, N2802, N1371, N2411);
xor XOR2 (N2809, N2808, N37);
nor NOR4 (N2810, N2807, N2639, N1593, N2786);
and AND4 (N2811, N2806, N1240, N2005, N1471);
and AND4 (N2812, N2811, N377, N281, N1887);
xor XOR2 (N2813, N2812, N115);
xor XOR2 (N2814, N2790, N652);
buf BUF1 (N2815, N2797);
or OR3 (N2816, N2813, N280, N401);
buf BUF1 (N2817, N2799);
xor XOR2 (N2818, N2810, N2513);
buf BUF1 (N2819, N2774);
not NOT1 (N2820, N2796);
and AND2 (N2821, N2814, N2295);
and AND4 (N2822, N2819, N2677, N555, N520);
or OR3 (N2823, N2821, N1528, N2740);
xor XOR2 (N2824, N2823, N2474);
nor NOR4 (N2825, N2822, N1577, N279, N1673);
or OR2 (N2826, N2809, N324);
and AND4 (N2827, N2801, N142, N384, N41);
and AND2 (N2828, N2826, N26);
not NOT1 (N2829, N2825);
buf BUF1 (N2830, N2818);
and AND4 (N2831, N2820, N78, N1883, N2578);
xor XOR2 (N2832, N2805, N1277);
not NOT1 (N2833, N2828);
or OR4 (N2834, N2831, N1194, N1246, N2034);
nand NAND2 (N2835, N2824, N234);
buf BUF1 (N2836, N2833);
not NOT1 (N2837, N2827);
xor XOR2 (N2838, N2834, N1216);
and AND3 (N2839, N2832, N689, N2737);
nand NAND2 (N2840, N2815, N1557);
buf BUF1 (N2841, N2830);
buf BUF1 (N2842, N2817);
nand NAND3 (N2843, N2829, N832, N297);
buf BUF1 (N2844, N2816);
or OR3 (N2845, N2837, N1108, N924);
xor XOR2 (N2846, N2840, N1843);
buf BUF1 (N2847, N2845);
xor XOR2 (N2848, N2844, N2146);
nand NAND4 (N2849, N2838, N1223, N856, N2584);
buf BUF1 (N2850, N2849);
buf BUF1 (N2851, N2848);
nand NAND3 (N2852, N2836, N2304, N2319);
and AND4 (N2853, N2841, N2040, N1278, N1880);
or OR4 (N2854, N2850, N842, N2243, N764);
nor NOR2 (N2855, N2851, N2521);
and AND3 (N2856, N2853, N793, N1123);
nor NOR2 (N2857, N2855, N1541);
xor XOR2 (N2858, N2854, N205);
or OR2 (N2859, N2839, N1725);
xor XOR2 (N2860, N2857, N1263);
nor NOR2 (N2861, N2856, N2203);
nor NOR3 (N2862, N2847, N1700, N2025);
xor XOR2 (N2863, N2862, N798);
xor XOR2 (N2864, N2843, N1499);
xor XOR2 (N2865, N2858, N1520);
not NOT1 (N2866, N2846);
nand NAND3 (N2867, N2860, N1033, N1978);
buf BUF1 (N2868, N2842);
nand NAND3 (N2869, N2864, N2342, N1647);
nand NAND2 (N2870, N2869, N2625);
nand NAND2 (N2871, N2868, N2238);
and AND4 (N2872, N2867, N2788, N573, N1438);
or OR2 (N2873, N2835, N737);
not NOT1 (N2874, N2861);
xor XOR2 (N2875, N2872, N1532);
xor XOR2 (N2876, N2852, N537);
not NOT1 (N2877, N2875);
not NOT1 (N2878, N2863);
nand NAND2 (N2879, N2878, N835);
or OR2 (N2880, N2871, N2405);
nand NAND3 (N2881, N2877, N201, N2669);
nor NOR2 (N2882, N2873, N593);
not NOT1 (N2883, N2876);
or OR4 (N2884, N2865, N1220, N2406, N564);
nand NAND4 (N2885, N2884, N2594, N2280, N1093);
or OR4 (N2886, N2874, N340, N429, N1167);
nand NAND3 (N2887, N2879, N1407, N1543);
buf BUF1 (N2888, N2880);
nor NOR4 (N2889, N2888, N2160, N1449, N2332);
nor NOR4 (N2890, N2886, N82, N1660, N1565);
buf BUF1 (N2891, N2889);
and AND2 (N2892, N2887, N2654);
and AND3 (N2893, N2866, N581, N1763);
nor NOR3 (N2894, N2892, N2692, N2419);
xor XOR2 (N2895, N2870, N1628);
nor NOR4 (N2896, N2891, N2710, N1155, N1372);
or OR4 (N2897, N2883, N2025, N1159, N2229);
xor XOR2 (N2898, N2897, N2796);
not NOT1 (N2899, N2896);
and AND4 (N2900, N2890, N339, N2698, N2141);
and AND3 (N2901, N2894, N2201, N2382);
xor XOR2 (N2902, N2901, N332);
or OR2 (N2903, N2900, N495);
buf BUF1 (N2904, N2903);
or OR2 (N2905, N2902, N963);
and AND3 (N2906, N2893, N1435, N1671);
and AND4 (N2907, N2859, N2282, N2509, N2341);
and AND2 (N2908, N2905, N81);
nor NOR3 (N2909, N2907, N2768, N1917);
or OR4 (N2910, N2895, N1159, N2796, N1676);
not NOT1 (N2911, N2881);
or OR4 (N2912, N2911, N993, N1489, N1852);
buf BUF1 (N2913, N2882);
and AND2 (N2914, N2910, N2848);
or OR4 (N2915, N2908, N1844, N746, N2003);
and AND3 (N2916, N2909, N2693, N744);
buf BUF1 (N2917, N2912);
buf BUF1 (N2918, N2914);
nor NOR2 (N2919, N2898, N518);
nor NOR2 (N2920, N2885, N728);
buf BUF1 (N2921, N2916);
buf BUF1 (N2922, N2906);
nor NOR2 (N2923, N2919, N1216);
buf BUF1 (N2924, N2921);
and AND2 (N2925, N2917, N2355);
not NOT1 (N2926, N2924);
buf BUF1 (N2927, N2904);
and AND3 (N2928, N2915, N2687, N681);
nor NOR4 (N2929, N2928, N2356, N2536, N2694);
xor XOR2 (N2930, N2929, N798);
buf BUF1 (N2931, N2920);
or OR4 (N2932, N2931, N2893, N523, N745);
xor XOR2 (N2933, N2922, N326);
nand NAND3 (N2934, N2933, N90, N1054);
nor NOR3 (N2935, N2913, N2219, N835);
nand NAND2 (N2936, N2932, N269);
buf BUF1 (N2937, N2936);
xor XOR2 (N2938, N2937, N1985);
and AND3 (N2939, N2923, N1523, N1668);
buf BUF1 (N2940, N2918);
xor XOR2 (N2941, N2930, N1071);
xor XOR2 (N2942, N2927, N1786);
xor XOR2 (N2943, N2926, N2597);
and AND2 (N2944, N2935, N1521);
nand NAND2 (N2945, N2942, N947);
and AND2 (N2946, N2925, N663);
or OR3 (N2947, N2934, N1697, N2798);
and AND2 (N2948, N2943, N1562);
buf BUF1 (N2949, N2945);
nand NAND4 (N2950, N2938, N475, N2670, N2048);
and AND4 (N2951, N2949, N1522, N1436, N2264);
xor XOR2 (N2952, N2950, N2020);
nor NOR3 (N2953, N2941, N482, N1322);
buf BUF1 (N2954, N2948);
buf BUF1 (N2955, N2940);
nor NOR3 (N2956, N2947, N1334, N2011);
and AND4 (N2957, N2952, N2492, N28, N952);
not NOT1 (N2958, N2939);
xor XOR2 (N2959, N2957, N2897);
not NOT1 (N2960, N2956);
buf BUF1 (N2961, N2960);
nor NOR3 (N2962, N2955, N1715, N2840);
nand NAND3 (N2963, N2944, N2357, N1358);
and AND3 (N2964, N2963, N408, N167);
xor XOR2 (N2965, N2951, N960);
nor NOR4 (N2966, N2946, N2562, N560, N638);
nand NAND3 (N2967, N2966, N1776, N928);
nor NOR2 (N2968, N2967, N561);
buf BUF1 (N2969, N2961);
xor XOR2 (N2970, N2969, N168);
not NOT1 (N2971, N2954);
and AND2 (N2972, N2899, N1432);
buf BUF1 (N2973, N2971);
nor NOR3 (N2974, N2968, N2547, N268);
not NOT1 (N2975, N2974);
or OR2 (N2976, N2953, N980);
nand NAND3 (N2977, N2958, N570, N1594);
nor NOR4 (N2978, N2976, N2914, N2565, N1330);
buf BUF1 (N2979, N2965);
not NOT1 (N2980, N2975);
xor XOR2 (N2981, N2959, N1029);
buf BUF1 (N2982, N2962);
nor NOR4 (N2983, N2973, N2463, N559, N186);
xor XOR2 (N2984, N2982, N398);
not NOT1 (N2985, N2981);
nand NAND2 (N2986, N2978, N1959);
or OR3 (N2987, N2980, N2016, N281);
and AND3 (N2988, N2977, N1927, N1742);
not NOT1 (N2989, N2970);
and AND4 (N2990, N2988, N426, N439, N1978);
or OR3 (N2991, N2989, N1202, N1654);
or OR2 (N2992, N2990, N660);
buf BUF1 (N2993, N2986);
not NOT1 (N2994, N2985);
and AND4 (N2995, N2993, N2830, N431, N516);
xor XOR2 (N2996, N2987, N2278);
xor XOR2 (N2997, N2972, N618);
nand NAND3 (N2998, N2991, N2230, N2592);
or OR3 (N2999, N2983, N222, N880);
nor NOR2 (N3000, N2997, N2326);
xor XOR2 (N3001, N3000, N2753);
or OR4 (N3002, N2984, N2383, N2064, N1978);
nand NAND4 (N3003, N2979, N1275, N964, N2169);
buf BUF1 (N3004, N2964);
and AND3 (N3005, N2994, N2307, N2734);
nor NOR4 (N3006, N3001, N1742, N106, N931);
and AND2 (N3007, N2998, N284);
or OR3 (N3008, N2996, N264, N214);
xor XOR2 (N3009, N3007, N2693);
or OR2 (N3010, N3005, N2833);
xor XOR2 (N3011, N3004, N2402);
buf BUF1 (N3012, N3008);
nand NAND3 (N3013, N3003, N551, N1881);
xor XOR2 (N3014, N3006, N2996);
or OR3 (N3015, N3012, N2261, N505);
and AND4 (N3016, N2992, N1886, N2645, N2156);
not NOT1 (N3017, N2999);
buf BUF1 (N3018, N3011);
buf BUF1 (N3019, N3010);
and AND4 (N3020, N3009, N1408, N1855, N1290);
nor NOR4 (N3021, N3019, N290, N1318, N243);
not NOT1 (N3022, N3020);
xor XOR2 (N3023, N3015, N658);
or OR2 (N3024, N3018, N744);
not NOT1 (N3025, N2995);
or OR4 (N3026, N3013, N591, N1888, N2932);
or OR3 (N3027, N3017, N1176, N2013);
nor NOR2 (N3028, N3002, N695);
or OR4 (N3029, N3028, N1483, N1423, N1774);
xor XOR2 (N3030, N3023, N1426);
xor XOR2 (N3031, N3030, N2377);
or OR3 (N3032, N3014, N1621, N2604);
nor NOR4 (N3033, N3025, N1779, N772, N397);
or OR2 (N3034, N3021, N2669);
not NOT1 (N3035, N3022);
xor XOR2 (N3036, N3035, N2689);
not NOT1 (N3037, N3016);
nor NOR2 (N3038, N3034, N2256);
not NOT1 (N3039, N3031);
or OR2 (N3040, N3029, N2205);
nor NOR4 (N3041, N3032, N2415, N187, N2800);
not NOT1 (N3042, N3041);
nand NAND2 (N3043, N3024, N259);
nand NAND4 (N3044, N3027, N2633, N2242, N445);
xor XOR2 (N3045, N3026, N788);
xor XOR2 (N3046, N3037, N2157);
and AND3 (N3047, N3036, N898, N1084);
or OR2 (N3048, N3038, N329);
buf BUF1 (N3049, N3042);
and AND3 (N3050, N3043, N1586, N902);
buf BUF1 (N3051, N3049);
buf BUF1 (N3052, N3046);
xor XOR2 (N3053, N3045, N148);
or OR4 (N3054, N3047, N1467, N2132, N2255);
nor NOR4 (N3055, N3040, N533, N1817, N372);
or OR3 (N3056, N3053, N2333, N190);
nand NAND2 (N3057, N3052, N1245);
and AND2 (N3058, N3055, N1284);
nand NAND2 (N3059, N3039, N458);
xor XOR2 (N3060, N3033, N432);
not NOT1 (N3061, N3048);
xor XOR2 (N3062, N3056, N782);
nor NOR3 (N3063, N3059, N2351, N268);
nand NAND4 (N3064, N3050, N755, N2597, N2702);
nor NOR3 (N3065, N3061, N1520, N829);
not NOT1 (N3066, N3054);
nand NAND4 (N3067, N3066, N1073, N425, N1918);
xor XOR2 (N3068, N3060, N2289);
buf BUF1 (N3069, N3044);
nor NOR4 (N3070, N3069, N1505, N1870, N1852);
xor XOR2 (N3071, N3064, N1575);
xor XOR2 (N3072, N3067, N2581);
buf BUF1 (N3073, N3071);
xor XOR2 (N3074, N3070, N850);
nand NAND4 (N3075, N3058, N2539, N349, N293);
and AND3 (N3076, N3065, N2600, N1084);
nor NOR3 (N3077, N3051, N78, N703);
not NOT1 (N3078, N3075);
nor NOR4 (N3079, N3076, N2797, N1944, N1313);
buf BUF1 (N3080, N3068);
buf BUF1 (N3081, N3074);
not NOT1 (N3082, N3062);
or OR3 (N3083, N3077, N1949, N1719);
or OR4 (N3084, N3078, N57, N648, N2974);
not NOT1 (N3085, N3084);
nor NOR4 (N3086, N3085, N2327, N1186, N463);
nor NOR3 (N3087, N3080, N829, N1125);
or OR2 (N3088, N3063, N582);
nor NOR4 (N3089, N3081, N2757, N1752, N2389);
nor NOR3 (N3090, N3089, N349, N2605);
nor NOR4 (N3091, N3057, N3036, N1192, N133);
not NOT1 (N3092, N3079);
xor XOR2 (N3093, N3082, N1027);
buf BUF1 (N3094, N3072);
nand NAND2 (N3095, N3092, N2064);
nor NOR2 (N3096, N3073, N2572);
nor NOR4 (N3097, N3091, N720, N52, N1029);
and AND3 (N3098, N3090, N2584, N1033);
and AND2 (N3099, N3096, N529);
nand NAND2 (N3100, N3094, N280);
or OR4 (N3101, N3088, N2925, N2458, N1221);
and AND4 (N3102, N3095, N444, N917, N2489);
buf BUF1 (N3103, N3083);
nor NOR4 (N3104, N3087, N2164, N2827, N1411);
and AND4 (N3105, N3104, N244, N165, N1946);
nand NAND3 (N3106, N3097, N634, N253);
and AND2 (N3107, N3093, N1086);
buf BUF1 (N3108, N3105);
and AND2 (N3109, N3086, N1232);
nor NOR4 (N3110, N3101, N10, N1296, N2108);
or OR2 (N3111, N3107, N2829);
nand NAND3 (N3112, N3100, N2983, N2640);
nand NAND3 (N3113, N3103, N2284, N346);
buf BUF1 (N3114, N3108);
and AND3 (N3115, N3114, N1790, N1167);
nor NOR4 (N3116, N3098, N2166, N1914, N593);
xor XOR2 (N3117, N3112, N1775);
nor NOR4 (N3118, N3109, N1290, N1946, N899);
or OR2 (N3119, N3111, N352);
xor XOR2 (N3120, N3113, N1980);
nand NAND3 (N3121, N3102, N2687, N560);
nor NOR2 (N3122, N3121, N2056);
nor NOR2 (N3123, N3110, N1986);
nor NOR3 (N3124, N3119, N1167, N1527);
nor NOR4 (N3125, N3123, N1115, N1527, N1423);
nor NOR3 (N3126, N3106, N1058, N431);
buf BUF1 (N3127, N3122);
and AND3 (N3128, N3118, N623, N999);
and AND4 (N3129, N3124, N1233, N2817, N1144);
or OR3 (N3130, N3127, N2108, N386);
nor NOR4 (N3131, N3126, N2113, N1139, N2457);
or OR3 (N3132, N3129, N2700, N280);
and AND4 (N3133, N3099, N729, N1571, N1463);
and AND2 (N3134, N3116, N1689);
not NOT1 (N3135, N3117);
and AND4 (N3136, N3115, N161, N2711, N2416);
nand NAND2 (N3137, N3128, N1325);
nand NAND3 (N3138, N3120, N1901, N181);
or OR4 (N3139, N3133, N1449, N805, N685);
not NOT1 (N3140, N3131);
and AND3 (N3141, N3130, N1127, N2102);
or OR2 (N3142, N3137, N3067);
xor XOR2 (N3143, N3142, N2995);
buf BUF1 (N3144, N3125);
nand NAND3 (N3145, N3141, N582, N1972);
and AND3 (N3146, N3143, N1600, N2905);
buf BUF1 (N3147, N3146);
nor NOR2 (N3148, N3145, N2113);
or OR3 (N3149, N3144, N1162, N3038);
xor XOR2 (N3150, N3135, N2386);
and AND3 (N3151, N3149, N2292, N1616);
nor NOR2 (N3152, N3134, N1758);
nor NOR3 (N3153, N3140, N410, N763);
nand NAND4 (N3154, N3132, N1156, N586, N230);
buf BUF1 (N3155, N3136);
xor XOR2 (N3156, N3153, N869);
nand NAND4 (N3157, N3139, N967, N1577, N2711);
or OR2 (N3158, N3138, N2138);
nand NAND4 (N3159, N3148, N1472, N2333, N1436);
not NOT1 (N3160, N3151);
or OR4 (N3161, N3160, N2407, N1844, N726);
xor XOR2 (N3162, N3156, N3101);
nand NAND3 (N3163, N3147, N98, N1095);
nor NOR4 (N3164, N3163, N1611, N199, N2654);
nor NOR2 (N3165, N3157, N661);
not NOT1 (N3166, N3155);
nand NAND3 (N3167, N3162, N972, N1097);
nor NOR2 (N3168, N3167, N2205);
buf BUF1 (N3169, N3168);
and AND2 (N3170, N3159, N179);
or OR4 (N3171, N3152, N1300, N1665, N2976);
nor NOR2 (N3172, N3171, N228);
not NOT1 (N3173, N3164);
nand NAND4 (N3174, N3166, N1378, N1519, N125);
nand NAND4 (N3175, N3169, N1370, N2217, N2351);
or OR4 (N3176, N3154, N1687, N1337, N450);
not NOT1 (N3177, N3170);
nor NOR2 (N3178, N3175, N2218);
nor NOR4 (N3179, N3165, N213, N107, N2237);
and AND3 (N3180, N3176, N3118, N964);
or OR3 (N3181, N3158, N1971, N2873);
not NOT1 (N3182, N3177);
nand NAND3 (N3183, N3174, N1022, N649);
and AND4 (N3184, N3173, N3182, N2244, N2579);
or OR3 (N3185, N1102, N2752, N2896);
xor XOR2 (N3186, N3179, N260);
buf BUF1 (N3187, N3180);
not NOT1 (N3188, N3150);
xor XOR2 (N3189, N3187, N1084);
and AND2 (N3190, N3186, N2796);
xor XOR2 (N3191, N3161, N357);
nand NAND3 (N3192, N3184, N2060, N1590);
nand NAND2 (N3193, N3192, N2825);
buf BUF1 (N3194, N3189);
nor NOR3 (N3195, N3194, N2701, N781);
and AND4 (N3196, N3188, N1238, N2683, N1417);
or OR4 (N3197, N3195, N2136, N555, N440);
not NOT1 (N3198, N3197);
nand NAND2 (N3199, N3183, N1925);
and AND2 (N3200, N3172, N3097);
nor NOR3 (N3201, N3178, N2318, N437);
buf BUF1 (N3202, N3185);
and AND2 (N3203, N3181, N1725);
and AND4 (N3204, N3193, N2271, N2379, N2041);
xor XOR2 (N3205, N3200, N2317);
nor NOR2 (N3206, N3196, N656);
buf BUF1 (N3207, N3190);
xor XOR2 (N3208, N3201, N314);
xor XOR2 (N3209, N3203, N1649);
not NOT1 (N3210, N3198);
not NOT1 (N3211, N3207);
nor NOR2 (N3212, N3199, N2420);
xor XOR2 (N3213, N3211, N1798);
not NOT1 (N3214, N3206);
xor XOR2 (N3215, N3214, N2369);
or OR2 (N3216, N3209, N1987);
and AND3 (N3217, N3202, N3179, N2087);
not NOT1 (N3218, N3217);
not NOT1 (N3219, N3213);
buf BUF1 (N3220, N3215);
nand NAND2 (N3221, N3204, N383);
xor XOR2 (N3222, N3210, N3194);
or OR3 (N3223, N3205, N2587, N607);
buf BUF1 (N3224, N3221);
not NOT1 (N3225, N3218);
and AND3 (N3226, N3208, N1844, N2833);
xor XOR2 (N3227, N3222, N2942);
and AND2 (N3228, N3220, N2996);
buf BUF1 (N3229, N3219);
buf BUF1 (N3230, N3227);
xor XOR2 (N3231, N3226, N2623);
buf BUF1 (N3232, N3191);
nand NAND3 (N3233, N3232, N1743, N2168);
nand NAND4 (N3234, N3223, N2416, N605, N716);
xor XOR2 (N3235, N3234, N1972);
not NOT1 (N3236, N3228);
nand NAND2 (N3237, N3230, N877);
and AND3 (N3238, N3235, N1266, N879);
nand NAND4 (N3239, N3237, N1448, N805, N1339);
not NOT1 (N3240, N3233);
xor XOR2 (N3241, N3238, N1003);
not NOT1 (N3242, N3225);
xor XOR2 (N3243, N3231, N420);
buf BUF1 (N3244, N3239);
not NOT1 (N3245, N3236);
or OR2 (N3246, N3242, N1499);
buf BUF1 (N3247, N3241);
or OR4 (N3248, N3212, N1426, N561, N41);
nand NAND4 (N3249, N3229, N3159, N2734, N949);
nand NAND2 (N3250, N3216, N2828);
and AND3 (N3251, N3245, N2744, N1496);
xor XOR2 (N3252, N3240, N2146);
buf BUF1 (N3253, N3250);
and AND2 (N3254, N3246, N518);
or OR2 (N3255, N3247, N2320);
xor XOR2 (N3256, N3224, N2710);
xor XOR2 (N3257, N3244, N1973);
and AND2 (N3258, N3249, N836);
buf BUF1 (N3259, N3254);
not NOT1 (N3260, N3251);
or OR2 (N3261, N3243, N1227);
nor NOR3 (N3262, N3256, N2914, N1829);
nor NOR3 (N3263, N3255, N1787, N2292);
or OR3 (N3264, N3263, N1037, N280);
and AND2 (N3265, N3252, N478);
not NOT1 (N3266, N3258);
and AND3 (N3267, N3248, N3066, N2624);
or OR4 (N3268, N3259, N96, N870, N3118);
nor NOR4 (N3269, N3261, N1584, N1477, N754);
xor XOR2 (N3270, N3268, N1100);
nand NAND3 (N3271, N3253, N827, N173);
xor XOR2 (N3272, N3270, N1711);
and AND2 (N3273, N3265, N1566);
nand NAND4 (N3274, N3260, N2478, N1846, N2927);
buf BUF1 (N3275, N3267);
not NOT1 (N3276, N3257);
xor XOR2 (N3277, N3269, N1324);
xor XOR2 (N3278, N3277, N1801);
buf BUF1 (N3279, N3274);
not NOT1 (N3280, N3279);
nand NAND2 (N3281, N3278, N80);
or OR2 (N3282, N3275, N1661);
nand NAND2 (N3283, N3276, N2994);
nand NAND2 (N3284, N3272, N1349);
or OR4 (N3285, N3281, N2439, N1260, N1821);
and AND4 (N3286, N3262, N1413, N294, N597);
or OR2 (N3287, N3286, N1331);
not NOT1 (N3288, N3285);
and AND2 (N3289, N3282, N3212);
buf BUF1 (N3290, N3284);
or OR4 (N3291, N3288, N892, N1802, N494);
buf BUF1 (N3292, N3264);
and AND3 (N3293, N3271, N361, N3188);
buf BUF1 (N3294, N3280);
buf BUF1 (N3295, N3273);
and AND4 (N3296, N3292, N2868, N2513, N1491);
and AND2 (N3297, N3266, N1697);
nand NAND3 (N3298, N3287, N3232, N2659);
and AND4 (N3299, N3294, N328, N1996, N2973);
or OR2 (N3300, N3283, N419);
xor XOR2 (N3301, N3299, N483);
or OR3 (N3302, N3295, N804, N2879);
or OR4 (N3303, N3298, N1187, N2169, N1214);
xor XOR2 (N3304, N3293, N2232);
buf BUF1 (N3305, N3290);
nand NAND2 (N3306, N3303, N2191);
buf BUF1 (N3307, N3304);
nand NAND3 (N3308, N3296, N2932, N2815);
buf BUF1 (N3309, N3302);
or OR3 (N3310, N3300, N2023, N683);
nand NAND3 (N3311, N3301, N631, N2015);
not NOT1 (N3312, N3311);
nor NOR2 (N3313, N3308, N3276);
or OR3 (N3314, N3309, N1489, N1327);
nor NOR4 (N3315, N3312, N2369, N862, N198);
buf BUF1 (N3316, N3315);
buf BUF1 (N3317, N3306);
nand NAND4 (N3318, N3313, N1519, N1733, N3180);
xor XOR2 (N3319, N3305, N3144);
xor XOR2 (N3320, N3310, N969);
nor NOR2 (N3321, N3318, N3140);
nor NOR2 (N3322, N3321, N603);
and AND4 (N3323, N3319, N2992, N1539, N710);
buf BUF1 (N3324, N3322);
xor XOR2 (N3325, N3307, N2131);
buf BUF1 (N3326, N3317);
buf BUF1 (N3327, N3314);
xor XOR2 (N3328, N3297, N3184);
buf BUF1 (N3329, N3326);
or OR2 (N3330, N3325, N3290);
buf BUF1 (N3331, N3329);
xor XOR2 (N3332, N3323, N1547);
or OR4 (N3333, N3330, N2987, N3091, N605);
buf BUF1 (N3334, N3331);
or OR2 (N3335, N3332, N1161);
xor XOR2 (N3336, N3327, N1244);
xor XOR2 (N3337, N3328, N3222);
or OR2 (N3338, N3324, N2816);
nand NAND4 (N3339, N3338, N3238, N161, N3035);
nand NAND4 (N3340, N3336, N157, N643, N2809);
not NOT1 (N3341, N3339);
nand NAND3 (N3342, N3316, N1703, N3250);
and AND4 (N3343, N3335, N2651, N3065, N2673);
nor NOR3 (N3344, N3289, N424, N2558);
buf BUF1 (N3345, N3342);
nor NOR3 (N3346, N3333, N1783, N2493);
nor NOR2 (N3347, N3320, N2962);
nand NAND2 (N3348, N3334, N2376);
or OR4 (N3349, N3341, N2183, N3234, N2337);
nand NAND4 (N3350, N3345, N171, N1863, N639);
not NOT1 (N3351, N3337);
or OR4 (N3352, N3344, N1883, N2328, N1809);
or OR4 (N3353, N3348, N1456, N703, N947);
nand NAND2 (N3354, N3343, N2172);
and AND2 (N3355, N3340, N2758);
or OR2 (N3356, N3355, N983);
and AND2 (N3357, N3351, N515);
and AND2 (N3358, N3291, N1813);
xor XOR2 (N3359, N3347, N1428);
nor NOR2 (N3360, N3356, N631);
buf BUF1 (N3361, N3350);
and AND4 (N3362, N3349, N2950, N2135, N3249);
nor NOR3 (N3363, N3357, N2112, N1800);
and AND2 (N3364, N3360, N1988);
and AND3 (N3365, N3364, N340, N282);
or OR3 (N3366, N3346, N3349, N477);
xor XOR2 (N3367, N3352, N2107);
and AND2 (N3368, N3363, N547);
xor XOR2 (N3369, N3353, N625);
or OR4 (N3370, N3362, N2479, N2175, N319);
and AND3 (N3371, N3359, N2399, N1511);
and AND4 (N3372, N3370, N2254, N1679, N1777);
nand NAND3 (N3373, N3361, N2480, N345);
and AND3 (N3374, N3367, N1005, N3120);
xor XOR2 (N3375, N3354, N804);
xor XOR2 (N3376, N3358, N3046);
buf BUF1 (N3377, N3369);
not NOT1 (N3378, N3376);
nor NOR3 (N3379, N3371, N1407, N1393);
nand NAND2 (N3380, N3375, N148);
buf BUF1 (N3381, N3378);
not NOT1 (N3382, N3380);
buf BUF1 (N3383, N3365);
and AND2 (N3384, N3383, N210);
xor XOR2 (N3385, N3368, N1849);
nand NAND2 (N3386, N3379, N139);
nand NAND2 (N3387, N3382, N2714);
nand NAND4 (N3388, N3377, N873, N2816, N174);
buf BUF1 (N3389, N3384);
nand NAND2 (N3390, N3389, N1458);
not NOT1 (N3391, N3385);
or OR4 (N3392, N3373, N544, N828, N2387);
xor XOR2 (N3393, N3388, N2654);
and AND2 (N3394, N3390, N566);
and AND3 (N3395, N3366, N617, N1222);
nor NOR3 (N3396, N3374, N3271, N949);
nand NAND4 (N3397, N3372, N20, N3000, N2827);
or OR2 (N3398, N3395, N1480);
nor NOR4 (N3399, N3392, N288, N1830, N615);
nand NAND2 (N3400, N3396, N520);
not NOT1 (N3401, N3400);
and AND2 (N3402, N3391, N1811);
or OR4 (N3403, N3399, N2910, N1688, N3101);
nand NAND4 (N3404, N3402, N3115, N807, N2648);
xor XOR2 (N3405, N3394, N965);
buf BUF1 (N3406, N3405);
or OR2 (N3407, N3386, N2971);
or OR2 (N3408, N3406, N1544);
buf BUF1 (N3409, N3408);
xor XOR2 (N3410, N3398, N378);
nor NOR4 (N3411, N3409, N3257, N2384, N418);
nand NAND4 (N3412, N3393, N179, N50, N1919);
nor NOR4 (N3413, N3407, N1233, N877, N143);
and AND3 (N3414, N3411, N903, N3205);
nand NAND3 (N3415, N3414, N711, N409);
not NOT1 (N3416, N3401);
buf BUF1 (N3417, N3397);
or OR3 (N3418, N3417, N1148, N3409);
nor NOR4 (N3419, N3412, N1904, N3402, N949);
not NOT1 (N3420, N3387);
xor XOR2 (N3421, N3418, N3223);
nand NAND4 (N3422, N3420, N1614, N1267, N2280);
nand NAND3 (N3423, N3403, N3024, N1454);
xor XOR2 (N3424, N3381, N2991);
nand NAND3 (N3425, N3404, N368, N3376);
nand NAND2 (N3426, N3419, N1335);
xor XOR2 (N3427, N3415, N2375);
xor XOR2 (N3428, N3416, N1232);
not NOT1 (N3429, N3428);
not NOT1 (N3430, N3423);
buf BUF1 (N3431, N3427);
buf BUF1 (N3432, N3426);
or OR2 (N3433, N3431, N202);
not NOT1 (N3434, N3433);
nand NAND3 (N3435, N3429, N2115, N1832);
or OR2 (N3436, N3421, N658);
nand NAND2 (N3437, N3410, N1461);
buf BUF1 (N3438, N3437);
xor XOR2 (N3439, N3434, N3029);
or OR3 (N3440, N3422, N1125, N2591);
not NOT1 (N3441, N3413);
xor XOR2 (N3442, N3432, N3319);
xor XOR2 (N3443, N3425, N1792);
nor NOR2 (N3444, N3442, N1381);
not NOT1 (N3445, N3424);
nand NAND4 (N3446, N3440, N458, N1251, N2680);
xor XOR2 (N3447, N3438, N3232);
buf BUF1 (N3448, N3444);
and AND4 (N3449, N3446, N2593, N2042, N1272);
nand NAND2 (N3450, N3447, N2143);
and AND2 (N3451, N3436, N1546);
xor XOR2 (N3452, N3450, N219);
and AND2 (N3453, N3451, N1187);
nor NOR2 (N3454, N3439, N838);
or OR4 (N3455, N3448, N1029, N565, N2955);
nand NAND4 (N3456, N3454, N2152, N1194, N1963);
xor XOR2 (N3457, N3455, N3414);
nand NAND4 (N3458, N3441, N437, N621, N714);
nor NOR2 (N3459, N3458, N1817);
buf BUF1 (N3460, N3445);
and AND4 (N3461, N3430, N2724, N1785, N1591);
or OR4 (N3462, N3453, N1489, N1094, N2978);
buf BUF1 (N3463, N3459);
xor XOR2 (N3464, N3457, N771);
not NOT1 (N3465, N3463);
nand NAND4 (N3466, N3456, N1278, N1308, N3083);
nor NOR4 (N3467, N3466, N3313, N2272, N1319);
buf BUF1 (N3468, N3464);
buf BUF1 (N3469, N3449);
or OR2 (N3470, N3443, N2281);
or OR2 (N3471, N3467, N1907);
or OR4 (N3472, N3465, N2848, N1633, N2177);
nor NOR3 (N3473, N3435, N3193, N111);
nor NOR3 (N3474, N3471, N2511, N2732);
or OR2 (N3475, N3474, N2493);
xor XOR2 (N3476, N3462, N39);
and AND4 (N3477, N3460, N3330, N3112, N2356);
nand NAND3 (N3478, N3470, N811, N2860);
nand NAND2 (N3479, N3478, N1457);
buf BUF1 (N3480, N3468);
buf BUF1 (N3481, N3452);
nand NAND4 (N3482, N3469, N3143, N882, N1445);
buf BUF1 (N3483, N3480);
or OR3 (N3484, N3473, N2658, N115);
xor XOR2 (N3485, N3472, N3311);
nand NAND3 (N3486, N3461, N2624, N60);
not NOT1 (N3487, N3485);
buf BUF1 (N3488, N3482);
or OR2 (N3489, N3476, N2610);
or OR2 (N3490, N3488, N1998);
nor NOR4 (N3491, N3489, N2918, N2158, N527);
not NOT1 (N3492, N3490);
not NOT1 (N3493, N3479);
not NOT1 (N3494, N3491);
not NOT1 (N3495, N3494);
buf BUF1 (N3496, N3483);
nor NOR3 (N3497, N3487, N2816, N2800);
nor NOR3 (N3498, N3475, N2149, N2785);
buf BUF1 (N3499, N3481);
nand NAND3 (N3500, N3492, N1104, N3479);
buf BUF1 (N3501, N3495);
not NOT1 (N3502, N3484);
and AND4 (N3503, N3496, N1202, N2050, N1286);
buf BUF1 (N3504, N3502);
and AND3 (N3505, N3486, N2628, N2895);
nor NOR4 (N3506, N3505, N1547, N1304, N1005);
and AND4 (N3507, N3503, N1629, N962, N3073);
xor XOR2 (N3508, N3501, N1618);
or OR2 (N3509, N3498, N1800);
xor XOR2 (N3510, N3493, N1690);
buf BUF1 (N3511, N3477);
or OR2 (N3512, N3507, N3314);
and AND3 (N3513, N3506, N1215, N3271);
nor NOR2 (N3514, N3508, N62);
buf BUF1 (N3515, N3500);
and AND4 (N3516, N3511, N1939, N2739, N629);
or OR2 (N3517, N3512, N283);
nand NAND2 (N3518, N3516, N2914);
nand NAND4 (N3519, N3497, N3417, N125, N407);
not NOT1 (N3520, N3514);
nand NAND4 (N3521, N3513, N3159, N1155, N900);
xor XOR2 (N3522, N3504, N1593);
buf BUF1 (N3523, N3510);
or OR3 (N3524, N3518, N2900, N2663);
nand NAND3 (N3525, N3524, N22, N442);
or OR2 (N3526, N3525, N3131);
nor NOR4 (N3527, N3526, N3015, N3370, N2631);
not NOT1 (N3528, N3517);
buf BUF1 (N3529, N3528);
and AND4 (N3530, N3515, N514, N1057, N1730);
xor XOR2 (N3531, N3509, N2563);
or OR4 (N3532, N3531, N3523, N778, N320);
and AND2 (N3533, N1223, N1378);
not NOT1 (N3534, N3520);
nor NOR4 (N3535, N3522, N2696, N1167, N1990);
and AND4 (N3536, N3529, N3311, N2559, N2038);
or OR3 (N3537, N3527, N3216, N1756);
nor NOR3 (N3538, N3533, N1882, N1597);
nor NOR4 (N3539, N3534, N3515, N1593, N674);
nor NOR3 (N3540, N3519, N753, N2342);
or OR3 (N3541, N3537, N3165, N757);
nand NAND2 (N3542, N3536, N303);
or OR2 (N3543, N3540, N1070);
or OR4 (N3544, N3499, N1021, N705, N1021);
nand NAND2 (N3545, N3530, N1998);
and AND4 (N3546, N3545, N1572, N2693, N431);
not NOT1 (N3547, N3532);
xor XOR2 (N3548, N3539, N3102);
xor XOR2 (N3549, N3544, N1541);
and AND3 (N3550, N3548, N2693, N152);
and AND4 (N3551, N3535, N3034, N3243, N143);
nor NOR4 (N3552, N3551, N1446, N3219, N2163);
or OR2 (N3553, N3543, N2694);
nor NOR2 (N3554, N3542, N1282);
not NOT1 (N3555, N3546);
nand NAND4 (N3556, N3538, N828, N1587, N88);
and AND4 (N3557, N3554, N2041, N2769, N1182);
nor NOR2 (N3558, N3549, N2585);
or OR2 (N3559, N3552, N2465);
buf BUF1 (N3560, N3541);
xor XOR2 (N3561, N3555, N2283);
xor XOR2 (N3562, N3547, N2419);
not NOT1 (N3563, N3553);
nand NAND3 (N3564, N3561, N437, N1964);
and AND2 (N3565, N3559, N3107);
xor XOR2 (N3566, N3556, N1718);
xor XOR2 (N3567, N3563, N655);
nor NOR4 (N3568, N3567, N3042, N844, N2051);
and AND4 (N3569, N3562, N1989, N339, N482);
xor XOR2 (N3570, N3568, N3422);
not NOT1 (N3571, N3521);
nand NAND4 (N3572, N3564, N384, N2849, N3247);
and AND2 (N3573, N3572, N854);
xor XOR2 (N3574, N3573, N2454);
buf BUF1 (N3575, N3566);
nand NAND2 (N3576, N3575, N634);
nand NAND2 (N3577, N3550, N440);
or OR2 (N3578, N3577, N3413);
not NOT1 (N3579, N3576);
nand NAND2 (N3580, N3570, N2682);
buf BUF1 (N3581, N3558);
and AND4 (N3582, N3569, N2845, N1472, N3046);
buf BUF1 (N3583, N3557);
not NOT1 (N3584, N3560);
not NOT1 (N3585, N3581);
nand NAND4 (N3586, N3583, N2791, N333, N2722);
or OR4 (N3587, N3584, N2675, N2554, N1732);
nor NOR2 (N3588, N3578, N1565);
and AND4 (N3589, N3571, N593, N784, N3050);
xor XOR2 (N3590, N3582, N1667);
not NOT1 (N3591, N3588);
nand NAND4 (N3592, N3591, N1366, N1228, N2520);
or OR4 (N3593, N3586, N2087, N1196, N3310);
or OR2 (N3594, N3592, N604);
not NOT1 (N3595, N3565);
nand NAND3 (N3596, N3589, N2010, N1188);
or OR4 (N3597, N3574, N2157, N145, N431);
nor NOR2 (N3598, N3593, N663);
or OR2 (N3599, N3595, N2624);
and AND2 (N3600, N3587, N12);
nor NOR2 (N3601, N3599, N2188);
or OR2 (N3602, N3590, N218);
and AND3 (N3603, N3600, N550, N3535);
buf BUF1 (N3604, N3596);
and AND2 (N3605, N3585, N568);
nand NAND4 (N3606, N3579, N1342, N2836, N1547);
buf BUF1 (N3607, N3604);
and AND2 (N3608, N3605, N1497);
not NOT1 (N3609, N3603);
nor NOR3 (N3610, N3598, N3396, N2396);
nand NAND4 (N3611, N3609, N2593, N2974, N1205);
xor XOR2 (N3612, N3580, N1302);
buf BUF1 (N3613, N3610);
buf BUF1 (N3614, N3602);
nor NOR2 (N3615, N3612, N189);
buf BUF1 (N3616, N3594);
and AND3 (N3617, N3614, N1604, N482);
nor NOR4 (N3618, N3608, N1073, N3235, N1842);
or OR4 (N3619, N3618, N1633, N1932, N2601);
and AND3 (N3620, N3617, N428, N3113);
nand NAND4 (N3621, N3597, N3361, N2003, N3135);
or OR2 (N3622, N3607, N1398);
xor XOR2 (N3623, N3622, N772);
buf BUF1 (N3624, N3621);
or OR3 (N3625, N3615, N2173, N1904);
not NOT1 (N3626, N3613);
nand NAND2 (N3627, N3606, N1055);
nand NAND3 (N3628, N3624, N1787, N2975);
xor XOR2 (N3629, N3628, N2355);
and AND4 (N3630, N3619, N2286, N460, N914);
and AND2 (N3631, N3611, N536);
xor XOR2 (N3632, N3623, N1227);
or OR3 (N3633, N3631, N2432, N728);
nor NOR4 (N3634, N3632, N1022, N927, N1741);
nor NOR4 (N3635, N3629, N431, N929, N2006);
and AND3 (N3636, N3626, N1591, N1881);
not NOT1 (N3637, N3627);
buf BUF1 (N3638, N3633);
and AND4 (N3639, N3634, N3602, N436, N3134);
not NOT1 (N3640, N3638);
buf BUF1 (N3641, N3635);
nand NAND4 (N3642, N3639, N1214, N1618, N2313);
nor NOR2 (N3643, N3640, N181);
or OR2 (N3644, N3620, N2856);
or OR3 (N3645, N3641, N2367, N1776);
buf BUF1 (N3646, N3644);
or OR3 (N3647, N3630, N1971, N2046);
not NOT1 (N3648, N3637);
buf BUF1 (N3649, N3646);
xor XOR2 (N3650, N3648, N1127);
nand NAND4 (N3651, N3642, N1613, N2032, N3215);
not NOT1 (N3652, N3647);
nand NAND2 (N3653, N3651, N2115);
buf BUF1 (N3654, N3650);
nor NOR3 (N3655, N3654, N3364, N2113);
and AND4 (N3656, N3601, N458, N3531, N2550);
not NOT1 (N3657, N3649);
nor NOR2 (N3658, N3636, N2847);
or OR4 (N3659, N3657, N2246, N2712, N1237);
or OR3 (N3660, N3658, N124, N1875);
xor XOR2 (N3661, N3653, N1121);
xor XOR2 (N3662, N3659, N3650);
nor NOR3 (N3663, N3656, N2262, N806);
xor XOR2 (N3664, N3662, N1183);
nor NOR4 (N3665, N3661, N2276, N2696, N3002);
not NOT1 (N3666, N3645);
not NOT1 (N3667, N3625);
not NOT1 (N3668, N3663);
or OR4 (N3669, N3643, N3421, N3226, N662);
xor XOR2 (N3670, N3660, N2236);
buf BUF1 (N3671, N3665);
xor XOR2 (N3672, N3655, N2581);
not NOT1 (N3673, N3672);
not NOT1 (N3674, N3671);
not NOT1 (N3675, N3674);
or OR4 (N3676, N3667, N1825, N248, N3604);
nand NAND2 (N3677, N3664, N2581);
xor XOR2 (N3678, N3676, N2867);
or OR4 (N3679, N3670, N711, N1486, N3545);
or OR3 (N3680, N3652, N1823, N865);
and AND4 (N3681, N3679, N418, N2268, N1673);
or OR4 (N3682, N3666, N1448, N481, N1627);
and AND3 (N3683, N3673, N2792, N1374);
nand NAND2 (N3684, N3669, N1923);
not NOT1 (N3685, N3682);
xor XOR2 (N3686, N3668, N2656);
buf BUF1 (N3687, N3616);
and AND4 (N3688, N3685, N1560, N2772, N2913);
nand NAND4 (N3689, N3675, N1341, N1811, N2830);
nor NOR2 (N3690, N3686, N2801);
nand NAND3 (N3691, N3689, N292, N991);
nor NOR2 (N3692, N3677, N791);
buf BUF1 (N3693, N3681);
or OR3 (N3694, N3690, N273, N1475);
not NOT1 (N3695, N3693);
xor XOR2 (N3696, N3687, N2553);
xor XOR2 (N3697, N3695, N2874);
xor XOR2 (N3698, N3684, N1654);
or OR2 (N3699, N3688, N3430);
nor NOR3 (N3700, N3691, N3620, N295);
xor XOR2 (N3701, N3700, N203);
nor NOR4 (N3702, N3680, N1662, N3152, N883);
or OR3 (N3703, N3696, N3666, N1326);
nor NOR3 (N3704, N3694, N1487, N3101);
not NOT1 (N3705, N3701);
and AND3 (N3706, N3702, N2164, N3524);
nor NOR2 (N3707, N3692, N3039);
not NOT1 (N3708, N3699);
buf BUF1 (N3709, N3698);
buf BUF1 (N3710, N3705);
xor XOR2 (N3711, N3683, N1163);
buf BUF1 (N3712, N3706);
nand NAND4 (N3713, N3712, N2543, N22, N3023);
and AND2 (N3714, N3708, N453);
xor XOR2 (N3715, N3709, N2635);
buf BUF1 (N3716, N3703);
xor XOR2 (N3717, N3704, N1374);
xor XOR2 (N3718, N3714, N2213);
nand NAND3 (N3719, N3710, N915, N1521);
or OR2 (N3720, N3697, N894);
nor NOR3 (N3721, N3707, N1202, N1997);
nor NOR4 (N3722, N3713, N3030, N149, N1255);
buf BUF1 (N3723, N3722);
xor XOR2 (N3724, N3720, N2154);
buf BUF1 (N3725, N3721);
nor NOR3 (N3726, N3716, N2094, N2934);
not NOT1 (N3727, N3726);
and AND3 (N3728, N3717, N1430, N3485);
and AND2 (N3729, N3711, N381);
and AND3 (N3730, N3715, N1607, N664);
nand NAND2 (N3731, N3718, N2329);
nor NOR2 (N3732, N3678, N720);
or OR2 (N3733, N3731, N938);
xor XOR2 (N3734, N3728, N3362);
not NOT1 (N3735, N3733);
nor NOR4 (N3736, N3730, N3654, N255, N1968);
nor NOR4 (N3737, N3732, N2596, N469, N2952);
and AND4 (N3738, N3737, N2349, N1192, N1667);
and AND4 (N3739, N3734, N2568, N3698, N2585);
buf BUF1 (N3740, N3739);
buf BUF1 (N3741, N3738);
and AND3 (N3742, N3719, N2467, N556);
or OR2 (N3743, N3724, N2856);
and AND3 (N3744, N3729, N1708, N2312);
nor NOR4 (N3745, N3743, N2498, N2648, N779);
or OR3 (N3746, N3744, N2543, N2620);
not NOT1 (N3747, N3741);
xor XOR2 (N3748, N3723, N377);
and AND4 (N3749, N3736, N2686, N2466, N1441);
buf BUF1 (N3750, N3742);
xor XOR2 (N3751, N3747, N858);
buf BUF1 (N3752, N3725);
xor XOR2 (N3753, N3746, N525);
not NOT1 (N3754, N3745);
nand NAND2 (N3755, N3752, N2050);
nor NOR2 (N3756, N3727, N3479);
nor NOR4 (N3757, N3756, N2682, N3607, N1021);
xor XOR2 (N3758, N3751, N1797);
nand NAND2 (N3759, N3755, N867);
not NOT1 (N3760, N3757);
and AND3 (N3761, N3740, N3376, N2565);
buf BUF1 (N3762, N3758);
nand NAND2 (N3763, N3749, N163);
nor NOR3 (N3764, N3748, N684, N3529);
buf BUF1 (N3765, N3763);
nor NOR2 (N3766, N3759, N2491);
xor XOR2 (N3767, N3735, N2450);
xor XOR2 (N3768, N3760, N1017);
xor XOR2 (N3769, N3767, N2418);
nand NAND2 (N3770, N3766, N3036);
xor XOR2 (N3771, N3750, N3183);
not NOT1 (N3772, N3768);
or OR3 (N3773, N3769, N2056, N1384);
not NOT1 (N3774, N3764);
nor NOR3 (N3775, N3770, N1353, N3312);
nor NOR3 (N3776, N3762, N2738, N3104);
or OR2 (N3777, N3754, N2303);
and AND3 (N3778, N3777, N3141, N2137);
or OR2 (N3779, N3776, N310);
buf BUF1 (N3780, N3772);
or OR4 (N3781, N3778, N1167, N1044, N81);
nand NAND2 (N3782, N3780, N1605);
xor XOR2 (N3783, N3773, N2495);
buf BUF1 (N3784, N3765);
nor NOR3 (N3785, N3782, N2987, N1711);
not NOT1 (N3786, N3761);
xor XOR2 (N3787, N3785, N1826);
and AND4 (N3788, N3783, N3329, N678, N3532);
nand NAND3 (N3789, N3781, N1885, N2479);
buf BUF1 (N3790, N3771);
not NOT1 (N3791, N3788);
nor NOR2 (N3792, N3774, N2319);
not NOT1 (N3793, N3753);
nand NAND4 (N3794, N3784, N3522, N1745, N2814);
buf BUF1 (N3795, N3775);
buf BUF1 (N3796, N3791);
not NOT1 (N3797, N3796);
nand NAND2 (N3798, N3795, N722);
nor NOR4 (N3799, N3779, N17, N473, N3215);
or OR2 (N3800, N3794, N3227);
and AND4 (N3801, N3789, N3535, N3384, N1644);
nand NAND2 (N3802, N3786, N455);
nor NOR4 (N3803, N3792, N783, N465, N1758);
and AND3 (N3804, N3801, N557, N2030);
buf BUF1 (N3805, N3790);
and AND2 (N3806, N3798, N308);
nand NAND2 (N3807, N3806, N3279);
or OR3 (N3808, N3804, N1859, N630);
and AND2 (N3809, N3799, N3781);
not NOT1 (N3810, N3808);
xor XOR2 (N3811, N3787, N619);
buf BUF1 (N3812, N3809);
xor XOR2 (N3813, N3793, N349);
not NOT1 (N3814, N3802);
nor NOR3 (N3815, N3813, N20, N1605);
and AND3 (N3816, N3797, N1904, N2079);
nand NAND4 (N3817, N3807, N427, N1009, N1984);
nand NAND4 (N3818, N3817, N787, N711, N2867);
not NOT1 (N3819, N3810);
buf BUF1 (N3820, N3819);
not NOT1 (N3821, N3805);
nor NOR3 (N3822, N3803, N1757, N2794);
or OR3 (N3823, N3811, N2133, N2349);
nand NAND3 (N3824, N3822, N1810, N3596);
or OR4 (N3825, N3815, N1077, N1068, N3786);
xor XOR2 (N3826, N3816, N2528);
buf BUF1 (N3827, N3823);
nand NAND3 (N3828, N3818, N1492, N2065);
nor NOR2 (N3829, N3824, N1296);
or OR4 (N3830, N3800, N6, N502, N3114);
nand NAND2 (N3831, N3821, N2057);
nand NAND4 (N3832, N3812, N2534, N909, N2056);
nor NOR3 (N3833, N3832, N3020, N1629);
nand NAND4 (N3834, N3827, N2089, N2023, N1414);
not NOT1 (N3835, N3820);
xor XOR2 (N3836, N3835, N3255);
or OR2 (N3837, N3828, N2336);
not NOT1 (N3838, N3826);
buf BUF1 (N3839, N3825);
nor NOR3 (N3840, N3834, N1578, N3190);
buf BUF1 (N3841, N3838);
nor NOR4 (N3842, N3829, N482, N1138, N3703);
and AND2 (N3843, N3831, N1738);
buf BUF1 (N3844, N3842);
nor NOR3 (N3845, N3839, N2845, N2139);
not NOT1 (N3846, N3836);
xor XOR2 (N3847, N3837, N1226);
and AND3 (N3848, N3814, N3408, N865);
xor XOR2 (N3849, N3843, N3639);
xor XOR2 (N3850, N3849, N1134);
nor NOR4 (N3851, N3841, N2689, N1325, N2138);
not NOT1 (N3852, N3848);
nor NOR2 (N3853, N3833, N102);
buf BUF1 (N3854, N3830);
nor NOR3 (N3855, N3847, N1006, N3733);
nand NAND4 (N3856, N3840, N2789, N2952, N1133);
buf BUF1 (N3857, N3852);
xor XOR2 (N3858, N3846, N1676);
nor NOR2 (N3859, N3858, N2934);
buf BUF1 (N3860, N3845);
xor XOR2 (N3861, N3851, N1706);
xor XOR2 (N3862, N3859, N1988);
or OR4 (N3863, N3855, N3487, N510, N2772);
xor XOR2 (N3864, N3854, N521);
nor NOR2 (N3865, N3863, N3379);
xor XOR2 (N3866, N3856, N1822);
nor NOR2 (N3867, N3866, N2362);
xor XOR2 (N3868, N3850, N3329);
not NOT1 (N3869, N3860);
not NOT1 (N3870, N3864);
nand NAND4 (N3871, N3862, N87, N1624, N1573);
xor XOR2 (N3872, N3871, N955);
or OR2 (N3873, N3868, N2167);
nand NAND3 (N3874, N3861, N2278, N1473);
or OR2 (N3875, N3873, N3487);
nor NOR2 (N3876, N3865, N1259);
nand NAND3 (N3877, N3844, N187, N1125);
and AND3 (N3878, N3869, N2443, N1558);
or OR2 (N3879, N3878, N60);
or OR2 (N3880, N3872, N2903);
nor NOR3 (N3881, N3867, N693, N1113);
not NOT1 (N3882, N3870);
nand NAND2 (N3883, N3881, N622);
buf BUF1 (N3884, N3877);
nor NOR4 (N3885, N3876, N3539, N3719, N2698);
buf BUF1 (N3886, N3883);
buf BUF1 (N3887, N3853);
nor NOR2 (N3888, N3884, N861);
xor XOR2 (N3889, N3887, N656);
xor XOR2 (N3890, N3888, N3355);
not NOT1 (N3891, N3890);
nand NAND4 (N3892, N3875, N2501, N3356, N484);
buf BUF1 (N3893, N3889);
not NOT1 (N3894, N3880);
or OR2 (N3895, N3882, N246);
not NOT1 (N3896, N3874);
nand NAND3 (N3897, N3886, N2146, N567);
and AND3 (N3898, N3892, N716, N832);
nor NOR4 (N3899, N3891, N2192, N3572, N511);
buf BUF1 (N3900, N3898);
nor NOR4 (N3901, N3894, N1725, N1663, N3264);
and AND4 (N3902, N3896, N2508, N1903, N790);
buf BUF1 (N3903, N3893);
not NOT1 (N3904, N3897);
nor NOR2 (N3905, N3901, N981);
xor XOR2 (N3906, N3904, N2094);
nand NAND2 (N3907, N3903, N98);
and AND2 (N3908, N3907, N3491);
and AND4 (N3909, N3908, N1174, N18, N811);
and AND2 (N3910, N3895, N2455);
buf BUF1 (N3911, N3900);
not NOT1 (N3912, N3910);
xor XOR2 (N3913, N3911, N797);
and AND4 (N3914, N3885, N84, N2337, N296);
nor NOR3 (N3915, N3905, N3356, N1897);
nor NOR3 (N3916, N3914, N2061, N1598);
nand NAND4 (N3917, N3879, N3263, N1928, N1183);
nand NAND4 (N3918, N3906, N2254, N2665, N3012);
or OR4 (N3919, N3917, N1623, N620, N529);
nor NOR4 (N3920, N3913, N1976, N1689, N2346);
not NOT1 (N3921, N3919);
and AND4 (N3922, N3918, N2275, N336, N338);
buf BUF1 (N3923, N3921);
nand NAND4 (N3924, N3912, N2189, N2884, N378);
nand NAND4 (N3925, N3899, N232, N1749, N1578);
nand NAND3 (N3926, N3909, N1264, N1615);
buf BUF1 (N3927, N3922);
nor NOR4 (N3928, N3925, N751, N1261, N138);
and AND4 (N3929, N3857, N1199, N501, N30);
and AND4 (N3930, N3924, N932, N323, N2645);
not NOT1 (N3931, N3927);
or OR4 (N3932, N3915, N834, N551, N1402);
or OR3 (N3933, N3916, N2876, N3143);
and AND2 (N3934, N3920, N3653);
xor XOR2 (N3935, N3923, N3268);
nor NOR2 (N3936, N3926, N2975);
or OR4 (N3937, N3934, N947, N1153, N1715);
buf BUF1 (N3938, N3930);
buf BUF1 (N3939, N3929);
nand NAND3 (N3940, N3937, N2474, N1747);
nor NOR3 (N3941, N3902, N2789, N557);
xor XOR2 (N3942, N3932, N1290);
not NOT1 (N3943, N3935);
or OR3 (N3944, N3933, N3720, N597);
nor NOR4 (N3945, N3931, N385, N1541, N1015);
and AND2 (N3946, N3942, N2372);
and AND2 (N3947, N3928, N453);
nor NOR3 (N3948, N3938, N1775, N414);
xor XOR2 (N3949, N3948, N3727);
or OR4 (N3950, N3936, N543, N2955, N1132);
and AND3 (N3951, N3941, N330, N3067);
nor NOR3 (N3952, N3945, N1572, N1517);
not NOT1 (N3953, N3947);
nand NAND4 (N3954, N3953, N1545, N2088, N1033);
buf BUF1 (N3955, N3939);
or OR2 (N3956, N3949, N882);
or OR4 (N3957, N3954, N1465, N1024, N361);
xor XOR2 (N3958, N3943, N3514);
nor NOR3 (N3959, N3952, N3251, N2601);
and AND3 (N3960, N3955, N1091, N3951);
not NOT1 (N3961, N1616);
and AND4 (N3962, N3946, N78, N3937, N670);
nor NOR2 (N3963, N3960, N1585);
nand NAND3 (N3964, N3963, N1602, N816);
xor XOR2 (N3965, N3957, N2250);
not NOT1 (N3966, N3961);
xor XOR2 (N3967, N3966, N1398);
buf BUF1 (N3968, N3940);
or OR3 (N3969, N3958, N3724, N2480);
nand NAND2 (N3970, N3944, N3914);
and AND4 (N3971, N3964, N2901, N846, N3961);
not NOT1 (N3972, N3969);
nand NAND4 (N3973, N3959, N2124, N870, N1599);
or OR4 (N3974, N3973, N3807, N3158, N3889);
or OR3 (N3975, N3965, N903, N2819);
xor XOR2 (N3976, N3950, N3024);
buf BUF1 (N3977, N3968);
not NOT1 (N3978, N3972);
not NOT1 (N3979, N3970);
and AND4 (N3980, N3967, N1894, N2465, N167);
buf BUF1 (N3981, N3975);
xor XOR2 (N3982, N3974, N1523);
buf BUF1 (N3983, N3977);
nand NAND2 (N3984, N3980, N3114);
or OR4 (N3985, N3981, N3161, N2335, N812);
xor XOR2 (N3986, N3985, N2728);
not NOT1 (N3987, N3956);
or OR4 (N3988, N3984, N2176, N1921, N1953);
nand NAND4 (N3989, N3971, N3514, N3737, N371);
nor NOR4 (N3990, N3988, N901, N2413, N469);
and AND2 (N3991, N3983, N2740);
not NOT1 (N3992, N3962);
buf BUF1 (N3993, N3986);
and AND3 (N3994, N3990, N2635, N1517);
and AND4 (N3995, N3982, N2927, N3544, N3573);
and AND2 (N3996, N3994, N2358);
not NOT1 (N3997, N3978);
buf BUF1 (N3998, N3987);
not NOT1 (N3999, N3998);
nor NOR4 (N4000, N3997, N3832, N2630, N225);
xor XOR2 (N4001, N3999, N3966);
and AND2 (N4002, N3993, N634);
or OR3 (N4003, N4002, N1756, N2434);
nor NOR4 (N4004, N3996, N2610, N2053, N2069);
or OR2 (N4005, N3992, N524);
not NOT1 (N4006, N3991);
and AND3 (N4007, N4004, N2107, N3159);
xor XOR2 (N4008, N3995, N3225);
xor XOR2 (N4009, N4003, N1114);
buf BUF1 (N4010, N3989);
buf BUF1 (N4011, N4006);
buf BUF1 (N4012, N4001);
xor XOR2 (N4013, N4007, N3250);
not NOT1 (N4014, N3976);
and AND4 (N4015, N4010, N1977, N2664, N2170);
xor XOR2 (N4016, N4005, N2603);
xor XOR2 (N4017, N4011, N2074);
buf BUF1 (N4018, N4013);
nand NAND3 (N4019, N4008, N3090, N3112);
and AND2 (N4020, N4017, N3530);
buf BUF1 (N4021, N4018);
buf BUF1 (N4022, N4016);
buf BUF1 (N4023, N4012);
or OR3 (N4024, N4022, N2196, N2062);
not NOT1 (N4025, N4009);
xor XOR2 (N4026, N4014, N1010);
not NOT1 (N4027, N4026);
nand NAND2 (N4028, N4019, N1312);
not NOT1 (N4029, N4020);
not NOT1 (N4030, N4028);
not NOT1 (N4031, N3979);
buf BUF1 (N4032, N4031);
xor XOR2 (N4033, N4015, N896);
and AND2 (N4034, N4021, N2411);
or OR2 (N4035, N4032, N766);
or OR4 (N4036, N4023, N1488, N3893, N2753);
or OR2 (N4037, N4000, N2483);
nor NOR2 (N4038, N4036, N2230);
buf BUF1 (N4039, N4030);
nand NAND3 (N4040, N4038, N351, N2052);
xor XOR2 (N4041, N4035, N3893);
nor NOR2 (N4042, N4041, N1527);
not NOT1 (N4043, N4027);
or OR2 (N4044, N4039, N537);
or OR2 (N4045, N4043, N343);
nand NAND2 (N4046, N4024, N3179);
not NOT1 (N4047, N4040);
and AND4 (N4048, N4033, N1086, N1694, N1198);
xor XOR2 (N4049, N4047, N1767);
or OR4 (N4050, N4034, N1510, N2746, N4009);
or OR4 (N4051, N4050, N2138, N2191, N623);
buf BUF1 (N4052, N4046);
nor NOR2 (N4053, N4029, N661);
nor NOR2 (N4054, N4042, N1904);
not NOT1 (N4055, N4054);
or OR3 (N4056, N4048, N507, N3335);
and AND3 (N4057, N4053, N702, N562);
nand NAND3 (N4058, N4045, N3872, N109);
or OR3 (N4059, N4058, N1883, N991);
nor NOR4 (N4060, N4059, N409, N2620, N3703);
or OR2 (N4061, N4052, N1585);
and AND2 (N4062, N4049, N172);
nor NOR4 (N4063, N4057, N1786, N2532, N3227);
buf BUF1 (N4064, N4063);
not NOT1 (N4065, N4061);
nand NAND4 (N4066, N4051, N4041, N1562, N881);
buf BUF1 (N4067, N4062);
not NOT1 (N4068, N4056);
nand NAND2 (N4069, N4066, N163);
xor XOR2 (N4070, N4055, N752);
nor NOR2 (N4071, N4067, N30);
or OR4 (N4072, N4044, N3712, N3412, N3817);
nor NOR4 (N4073, N4037, N2734, N2784, N770);
xor XOR2 (N4074, N4060, N1223);
nand NAND2 (N4075, N4025, N1694);
xor XOR2 (N4076, N4072, N3992);
nor NOR4 (N4077, N4074, N1885, N1255, N2928);
xor XOR2 (N4078, N4077, N3094);
nand NAND2 (N4079, N4069, N687);
and AND3 (N4080, N4076, N1301, N2003);
or OR3 (N4081, N4068, N771, N2815);
not NOT1 (N4082, N4070);
buf BUF1 (N4083, N4079);
xor XOR2 (N4084, N4082, N1322);
xor XOR2 (N4085, N4065, N582);
buf BUF1 (N4086, N4085);
not NOT1 (N4087, N4083);
or OR3 (N4088, N4086, N3804, N3211);
nand NAND3 (N4089, N4073, N3947, N2186);
nand NAND2 (N4090, N4075, N2985);
nand NAND2 (N4091, N4081, N2148);
xor XOR2 (N4092, N4087, N2309);
nand NAND2 (N4093, N4064, N3905);
or OR3 (N4094, N4092, N2781, N3470);
or OR2 (N4095, N4089, N1308);
nand NAND4 (N4096, N4093, N385, N466, N1840);
or OR2 (N4097, N4091, N2054);
xor XOR2 (N4098, N4071, N538);
and AND2 (N4099, N4080, N2928);
nand NAND3 (N4100, N4097, N3296, N1892);
nand NAND2 (N4101, N4084, N3211);
nand NAND3 (N4102, N4088, N2903, N2458);
and AND3 (N4103, N4100, N3911, N444);
nand NAND2 (N4104, N4095, N1785);
nand NAND4 (N4105, N4098, N1215, N2042, N3793);
or OR4 (N4106, N4094, N2515, N1096, N48);
xor XOR2 (N4107, N4102, N1385);
buf BUF1 (N4108, N4106);
or OR2 (N4109, N4090, N747);
or OR4 (N4110, N4104, N3658, N3824, N1038);
nand NAND3 (N4111, N4099, N1638, N2911);
nor NOR2 (N4112, N4096, N3623);
nor NOR2 (N4113, N4112, N780);
xor XOR2 (N4114, N4078, N1638);
nand NAND3 (N4115, N4107, N1125, N1418);
and AND3 (N4116, N4111, N3263, N3003);
nand NAND2 (N4117, N4101, N1307);
nor NOR4 (N4118, N4105, N1660, N1288, N2225);
nand NAND2 (N4119, N4115, N2710);
xor XOR2 (N4120, N4110, N1342);
buf BUF1 (N4121, N4120);
not NOT1 (N4122, N4103);
nand NAND3 (N4123, N4108, N2547, N1508);
xor XOR2 (N4124, N4123, N1969);
buf BUF1 (N4125, N4114);
or OR4 (N4126, N4121, N1234, N87, N1333);
xor XOR2 (N4127, N4116, N3922);
not NOT1 (N4128, N4122);
buf BUF1 (N4129, N4119);
buf BUF1 (N4130, N4127);
nor NOR4 (N4131, N4126, N1420, N2195, N2711);
nand NAND3 (N4132, N4125, N1385, N2941);
xor XOR2 (N4133, N4132, N591);
nor NOR2 (N4134, N4131, N4003);
xor XOR2 (N4135, N4124, N1556);
nand NAND3 (N4136, N4134, N1661, N324);
buf BUF1 (N4137, N4113);
buf BUF1 (N4138, N4109);
and AND4 (N4139, N4118, N938, N2696, N2264);
buf BUF1 (N4140, N4136);
or OR2 (N4141, N4137, N420);
and AND4 (N4142, N4140, N3512, N2328, N1932);
and AND4 (N4143, N4128, N1597, N1475, N2679);
not NOT1 (N4144, N4142);
xor XOR2 (N4145, N4135, N3152);
xor XOR2 (N4146, N4130, N1847);
not NOT1 (N4147, N4146);
or OR4 (N4148, N4138, N3171, N1694, N1379);
and AND2 (N4149, N4117, N1059);
xor XOR2 (N4150, N4148, N4112);
nand NAND4 (N4151, N4139, N733, N1194, N112);
and AND3 (N4152, N4147, N2001, N3701);
not NOT1 (N4153, N4149);
nand NAND2 (N4154, N4133, N629);
or OR4 (N4155, N4153, N9, N1439, N2832);
nor NOR2 (N4156, N4150, N27);
not NOT1 (N4157, N4141);
xor XOR2 (N4158, N4145, N478);
and AND3 (N4159, N4154, N4030, N2683);
buf BUF1 (N4160, N4156);
buf BUF1 (N4161, N4155);
not NOT1 (N4162, N4159);
xor XOR2 (N4163, N4160, N2559);
nor NOR2 (N4164, N4152, N1953);
not NOT1 (N4165, N4129);
or OR4 (N4166, N4144, N3180, N2847, N2246);
buf BUF1 (N4167, N4161);
not NOT1 (N4168, N4158);
buf BUF1 (N4169, N4165);
and AND2 (N4170, N4162, N1943);
buf BUF1 (N4171, N4163);
nand NAND4 (N4172, N4167, N568, N2329, N1745);
not NOT1 (N4173, N4169);
nand NAND2 (N4174, N4170, N2365);
xor XOR2 (N4175, N4174, N2916);
buf BUF1 (N4176, N4171);
not NOT1 (N4177, N4166);
nand NAND3 (N4178, N4176, N3680, N2286);
buf BUF1 (N4179, N4175);
nor NOR2 (N4180, N4143, N934);
nor NOR3 (N4181, N4180, N3631, N634);
or OR3 (N4182, N4168, N4096, N310);
xor XOR2 (N4183, N4157, N4080);
or OR4 (N4184, N4164, N561, N3057, N2021);
xor XOR2 (N4185, N4178, N97);
nor NOR3 (N4186, N4184, N247, N3145);
not NOT1 (N4187, N4185);
xor XOR2 (N4188, N4151, N120);
and AND4 (N4189, N4179, N2554, N2273, N899);
and AND4 (N4190, N4186, N2566, N2526, N2942);
and AND3 (N4191, N4172, N578, N15);
buf BUF1 (N4192, N4181);
nor NOR4 (N4193, N4189, N3480, N232, N880);
xor XOR2 (N4194, N4173, N2019);
or OR3 (N4195, N4188, N726, N732);
xor XOR2 (N4196, N4194, N2658);
and AND3 (N4197, N4191, N1867, N179);
xor XOR2 (N4198, N4190, N1802);
or OR4 (N4199, N4187, N1819, N3712, N2735);
buf BUF1 (N4200, N4193);
buf BUF1 (N4201, N4182);
not NOT1 (N4202, N4198);
or OR2 (N4203, N4200, N751);
nand NAND4 (N4204, N4203, N3043, N3868, N3059);
not NOT1 (N4205, N4201);
nand NAND4 (N4206, N4199, N3014, N743, N3017);
xor XOR2 (N4207, N4183, N1058);
and AND3 (N4208, N4204, N1071, N3156);
nor NOR4 (N4209, N4206, N28, N4060, N2306);
xor XOR2 (N4210, N4208, N3791);
nor NOR3 (N4211, N4192, N2492, N3804);
not NOT1 (N4212, N4195);
nand NAND2 (N4213, N4212, N1079);
or OR4 (N4214, N4211, N2868, N3713, N780);
buf BUF1 (N4215, N4209);
xor XOR2 (N4216, N4197, N2916);
not NOT1 (N4217, N4215);
or OR4 (N4218, N4210, N1040, N4026, N1264);
nand NAND4 (N4219, N4196, N2256, N3007, N535);
or OR4 (N4220, N4213, N3939, N2283, N3354);
buf BUF1 (N4221, N4177);
and AND4 (N4222, N4217, N2302, N2878, N530);
not NOT1 (N4223, N4214);
nor NOR3 (N4224, N4220, N2212, N669);
nor NOR3 (N4225, N4216, N1495, N4208);
nor NOR3 (N4226, N4221, N264, N356);
xor XOR2 (N4227, N4218, N620);
nand NAND3 (N4228, N4222, N518, N2908);
buf BUF1 (N4229, N4205);
nor NOR2 (N4230, N4207, N3290);
buf BUF1 (N4231, N4224);
nand NAND3 (N4232, N4229, N1070, N1068);
or OR4 (N4233, N4231, N3185, N1652, N3892);
buf BUF1 (N4234, N4202);
and AND4 (N4235, N4225, N3755, N2583, N2353);
or OR3 (N4236, N4232, N67, N349);
not NOT1 (N4237, N4228);
not NOT1 (N4238, N4234);
or OR2 (N4239, N4236, N1047);
nand NAND2 (N4240, N4239, N3639);
not NOT1 (N4241, N4230);
not NOT1 (N4242, N4219);
nor NOR2 (N4243, N4238, N3618);
nand NAND3 (N4244, N4243, N1387, N1920);
xor XOR2 (N4245, N4244, N579);
and AND3 (N4246, N4241, N184, N1757);
or OR3 (N4247, N4226, N3116, N3026);
and AND3 (N4248, N4240, N2018, N445);
not NOT1 (N4249, N4223);
nor NOR4 (N4250, N4247, N3057, N1916, N237);
nor NOR2 (N4251, N4242, N3427);
nor NOR3 (N4252, N4233, N3607, N2667);
or OR4 (N4253, N4237, N3869, N1616, N1941);
buf BUF1 (N4254, N4253);
not NOT1 (N4255, N4249);
or OR3 (N4256, N4248, N2796, N4063);
nor NOR3 (N4257, N4235, N3075, N987);
not NOT1 (N4258, N4252);
nand NAND4 (N4259, N4258, N381, N2746, N2519);
xor XOR2 (N4260, N4250, N3162);
not NOT1 (N4261, N4227);
and AND4 (N4262, N4261, N490, N4257, N2939);
nand NAND4 (N4263, N138, N428, N2339, N2787);
xor XOR2 (N4264, N4255, N3188);
xor XOR2 (N4265, N4263, N4090);
nand NAND3 (N4266, N4246, N2020, N441);
xor XOR2 (N4267, N4251, N376);
and AND3 (N4268, N4245, N2494, N560);
nand NAND2 (N4269, N4265, N1536);
nor NOR2 (N4270, N4260, N1407);
not NOT1 (N4271, N4270);
and AND4 (N4272, N4259, N3913, N2969, N1045);
not NOT1 (N4273, N4268);
not NOT1 (N4274, N4273);
xor XOR2 (N4275, N4274, N2719);
and AND4 (N4276, N4264, N1164, N165, N2139);
or OR3 (N4277, N4272, N2378, N3503);
nand NAND4 (N4278, N4269, N2722, N420, N2249);
and AND4 (N4279, N4276, N2674, N3871, N4007);
nor NOR2 (N4280, N4254, N3814);
and AND3 (N4281, N4262, N1953, N4148);
not NOT1 (N4282, N4281);
nor NOR4 (N4283, N4266, N1808, N4048, N1546);
not NOT1 (N4284, N4256);
xor XOR2 (N4285, N4279, N601);
or OR2 (N4286, N4271, N1502);
xor XOR2 (N4287, N4277, N2277);
xor XOR2 (N4288, N4287, N3587);
nand NAND2 (N4289, N4288, N816);
nor NOR3 (N4290, N4289, N3261, N845);
not NOT1 (N4291, N4282);
nor NOR4 (N4292, N4291, N1497, N454, N903);
and AND3 (N4293, N4290, N4270, N1444);
buf BUF1 (N4294, N4286);
or OR4 (N4295, N4267, N1164, N1126, N1626);
xor XOR2 (N4296, N4275, N726);
nor NOR3 (N4297, N4280, N3172, N622);
buf BUF1 (N4298, N4284);
and AND4 (N4299, N4292, N663, N3441, N1275);
buf BUF1 (N4300, N4295);
or OR3 (N4301, N4300, N1178, N3193);
nor NOR3 (N4302, N4293, N2790, N1311);
not NOT1 (N4303, N4278);
nor NOR3 (N4304, N4294, N1770, N2576);
xor XOR2 (N4305, N4285, N2421);
and AND3 (N4306, N4298, N1827, N1766);
not NOT1 (N4307, N4301);
and AND2 (N4308, N4304, N675);
and AND4 (N4309, N4308, N2974, N1507, N871);
and AND4 (N4310, N4297, N6, N3401, N3062);
buf BUF1 (N4311, N4305);
not NOT1 (N4312, N4302);
not NOT1 (N4313, N4283);
buf BUF1 (N4314, N4312);
nand NAND4 (N4315, N4309, N45, N3614, N2812);
and AND4 (N4316, N4315, N922, N853, N1766);
or OR4 (N4317, N4313, N317, N2966, N2954);
xor XOR2 (N4318, N4310, N12);
buf BUF1 (N4319, N4296);
nor NOR2 (N4320, N4299, N816);
xor XOR2 (N4321, N4307, N2812);
or OR2 (N4322, N4314, N1152);
nor NOR2 (N4323, N4306, N4210);
or OR4 (N4324, N4316, N3212, N1280, N1138);
nand NAND2 (N4325, N4321, N1461);
nand NAND4 (N4326, N4322, N2346, N1339, N3324);
or OR2 (N4327, N4318, N3399);
buf BUF1 (N4328, N4320);
and AND2 (N4329, N4324, N3249);
xor XOR2 (N4330, N4325, N3189);
and AND3 (N4331, N4328, N603, N990);
and AND4 (N4332, N4329, N428, N2801, N3619);
not NOT1 (N4333, N4317);
xor XOR2 (N4334, N4330, N306);
nand NAND4 (N4335, N4323, N3448, N904, N2991);
and AND4 (N4336, N4311, N977, N3937, N4012);
buf BUF1 (N4337, N4327);
xor XOR2 (N4338, N4335, N3982);
xor XOR2 (N4339, N4331, N761);
and AND2 (N4340, N4333, N3796);
xor XOR2 (N4341, N4339, N2556);
and AND3 (N4342, N4326, N3802, N1971);
nor NOR3 (N4343, N4341, N1948, N2771);
nand NAND3 (N4344, N4336, N811, N3960);
and AND3 (N4345, N4344, N209, N1463);
xor XOR2 (N4346, N4338, N356);
nor NOR2 (N4347, N4319, N3556);
buf BUF1 (N4348, N4340);
nor NOR4 (N4349, N4343, N2711, N2517, N234);
nand NAND3 (N4350, N4346, N3078, N3135);
nand NAND4 (N4351, N4350, N3013, N4288, N2024);
buf BUF1 (N4352, N4342);
and AND3 (N4353, N4349, N779, N2604);
and AND3 (N4354, N4332, N4200, N3458);
buf BUF1 (N4355, N4351);
not NOT1 (N4356, N4353);
not NOT1 (N4357, N4334);
or OR3 (N4358, N4303, N3512, N1990);
not NOT1 (N4359, N4337);
or OR3 (N4360, N4356, N4305, N2453);
and AND4 (N4361, N4357, N4136, N178, N3636);
not NOT1 (N4362, N4358);
nor NOR3 (N4363, N4352, N3273, N769);
xor XOR2 (N4364, N4363, N788);
and AND3 (N4365, N4362, N1406, N2664);
nand NAND4 (N4366, N4345, N3565, N4017, N3475);
not NOT1 (N4367, N4365);
xor XOR2 (N4368, N4355, N2732);
and AND4 (N4369, N4361, N4295, N3429, N4001);
and AND2 (N4370, N4348, N1495);
not NOT1 (N4371, N4369);
nor NOR3 (N4372, N4347, N849, N3215);
and AND4 (N4373, N4354, N3999, N2688, N2640);
nand NAND2 (N4374, N4368, N4038);
or OR3 (N4375, N4372, N689, N656);
or OR4 (N4376, N4374, N2924, N513, N3923);
buf BUF1 (N4377, N4373);
nand NAND2 (N4378, N4364, N3702);
xor XOR2 (N4379, N4371, N2502);
nor NOR4 (N4380, N4377, N1279, N3071, N971);
buf BUF1 (N4381, N4360);
nand NAND3 (N4382, N4367, N1207, N1307);
xor XOR2 (N4383, N4375, N1764);
and AND2 (N4384, N4379, N29);
buf BUF1 (N4385, N4384);
not NOT1 (N4386, N4380);
and AND3 (N4387, N4366, N3146, N1385);
nor NOR3 (N4388, N4385, N2489, N3464);
not NOT1 (N4389, N4359);
not NOT1 (N4390, N4383);
or OR4 (N4391, N4378, N3667, N4319, N1626);
nand NAND3 (N4392, N4386, N1129, N164);
not NOT1 (N4393, N4388);
buf BUF1 (N4394, N4382);
buf BUF1 (N4395, N4381);
nand NAND2 (N4396, N4392, N310);
nand NAND4 (N4397, N4376, N1382, N4324, N997);
and AND3 (N4398, N4395, N2199, N1422);
not NOT1 (N4399, N4370);
not NOT1 (N4400, N4398);
or OR4 (N4401, N4399, N3315, N458, N3099);
or OR3 (N4402, N4397, N1980, N586);
nand NAND3 (N4403, N4387, N3403, N3494);
not NOT1 (N4404, N4390);
xor XOR2 (N4405, N4393, N3075);
not NOT1 (N4406, N4402);
nand NAND4 (N4407, N4404, N115, N1958, N459);
nand NAND3 (N4408, N4396, N3983, N3870);
or OR4 (N4409, N4406, N2324, N2557, N2563);
xor XOR2 (N4410, N4391, N3655);
and AND4 (N4411, N4394, N1188, N2727, N2321);
nand NAND4 (N4412, N4389, N2436, N2088, N1546);
not NOT1 (N4413, N4412);
or OR3 (N4414, N4411, N3241, N3424);
nand NAND4 (N4415, N4400, N394, N2749, N2014);
and AND3 (N4416, N4403, N2565, N2833);
or OR2 (N4417, N4410, N3704);
or OR3 (N4418, N4408, N1083, N2322);
or OR3 (N4419, N4409, N1745, N2597);
and AND2 (N4420, N4415, N640);
and AND3 (N4421, N4413, N720, N938);
buf BUF1 (N4422, N4414);
not NOT1 (N4423, N4405);
and AND3 (N4424, N4416, N1052, N1017);
xor XOR2 (N4425, N4420, N909);
and AND3 (N4426, N4419, N2450, N2035);
and AND2 (N4427, N4426, N248);
and AND3 (N4428, N4401, N2949, N292);
xor XOR2 (N4429, N4424, N3888);
not NOT1 (N4430, N4427);
buf BUF1 (N4431, N4418);
and AND2 (N4432, N4407, N1814);
and AND2 (N4433, N4417, N1220);
xor XOR2 (N4434, N4428, N924);
nor NOR3 (N4435, N4425, N2832, N2803);
nor NOR2 (N4436, N4421, N105);
nand NAND2 (N4437, N4431, N749);
nor NOR2 (N4438, N4435, N1270);
nand NAND2 (N4439, N4422, N3280);
nand NAND2 (N4440, N4434, N2403);
nor NOR4 (N4441, N4432, N1519, N2741, N1068);
xor XOR2 (N4442, N4436, N3979);
xor XOR2 (N4443, N4438, N2883);
not NOT1 (N4444, N4423);
not NOT1 (N4445, N4437);
buf BUF1 (N4446, N4445);
nor NOR4 (N4447, N4441, N1123, N2880, N2821);
or OR2 (N4448, N4440, N3382);
xor XOR2 (N4449, N4430, N4095);
not NOT1 (N4450, N4443);
nand NAND2 (N4451, N4448, N4286);
xor XOR2 (N4452, N4451, N2385);
xor XOR2 (N4453, N4449, N2654);
or OR3 (N4454, N4433, N1689, N2088);
xor XOR2 (N4455, N4453, N2260);
buf BUF1 (N4456, N4439);
nor NOR2 (N4457, N4450, N2583);
nor NOR4 (N4458, N4447, N1643, N1714, N628);
nand NAND4 (N4459, N4458, N1305, N920, N93);
nor NOR4 (N4460, N4459, N2871, N3616, N693);
and AND2 (N4461, N4452, N3663);
nand NAND4 (N4462, N4455, N1575, N562, N4329);
nor NOR3 (N4463, N4456, N3437, N3549);
buf BUF1 (N4464, N4444);
and AND3 (N4465, N4464, N3042, N4094);
and AND2 (N4466, N4460, N3761);
or OR2 (N4467, N4429, N3989);
buf BUF1 (N4468, N4466);
buf BUF1 (N4469, N4465);
nand NAND4 (N4470, N4468, N1454, N4070, N1641);
nor NOR3 (N4471, N4461, N1866, N3803);
and AND2 (N4472, N4470, N966);
buf BUF1 (N4473, N4454);
nand NAND3 (N4474, N4442, N4071, N1452);
buf BUF1 (N4475, N4474);
buf BUF1 (N4476, N4446);
nand NAND3 (N4477, N4476, N1868, N3242);
or OR4 (N4478, N4475, N1087, N1499, N4297);
and AND4 (N4479, N4471, N2071, N3479, N2201);
nor NOR3 (N4480, N4472, N1353, N1341);
and AND3 (N4481, N4469, N3424, N4013);
xor XOR2 (N4482, N4478, N1685);
and AND3 (N4483, N4467, N1203, N4047);
xor XOR2 (N4484, N4457, N1131);
or OR4 (N4485, N4477, N3223, N2701, N3453);
nor NOR2 (N4486, N4473, N1018);
nor NOR4 (N4487, N4485, N3465, N3799, N2250);
nor NOR3 (N4488, N4483, N1214, N2329);
nand NAND2 (N4489, N4462, N2328);
buf BUF1 (N4490, N4479);
nand NAND2 (N4491, N4482, N1291);
and AND2 (N4492, N4490, N4135);
xor XOR2 (N4493, N4491, N3092);
not NOT1 (N4494, N4488);
not NOT1 (N4495, N4492);
not NOT1 (N4496, N4480);
nor NOR3 (N4497, N4487, N221, N3398);
and AND4 (N4498, N4494, N3685, N1277, N646);
not NOT1 (N4499, N4493);
xor XOR2 (N4500, N4496, N3551);
nor NOR3 (N4501, N4499, N1607, N1164);
or OR3 (N4502, N4495, N3127, N3762);
or OR4 (N4503, N4501, N2858, N2167, N4162);
buf BUF1 (N4504, N4503);
nor NOR3 (N4505, N4489, N3208, N4141);
xor XOR2 (N4506, N4504, N2715);
xor XOR2 (N4507, N4498, N2602);
xor XOR2 (N4508, N4484, N3282);
or OR4 (N4509, N4508, N3929, N459, N4430);
and AND3 (N4510, N4509, N1020, N440);
xor XOR2 (N4511, N4497, N2644);
and AND2 (N4512, N4511, N754);
nand NAND2 (N4513, N4507, N2459);
or OR2 (N4514, N4510, N1103);
xor XOR2 (N4515, N4500, N548);
and AND2 (N4516, N4512, N810);
xor XOR2 (N4517, N4481, N843);
or OR4 (N4518, N4517, N3004, N1306, N3103);
nor NOR4 (N4519, N4506, N2241, N1754, N2560);
nand NAND3 (N4520, N4515, N2364, N2764);
and AND2 (N4521, N4518, N477);
nor NOR4 (N4522, N4519, N3385, N2249, N4235);
not NOT1 (N4523, N4514);
xor XOR2 (N4524, N4522, N2874);
or OR3 (N4525, N4502, N2845, N2267);
not NOT1 (N4526, N4525);
buf BUF1 (N4527, N4486);
not NOT1 (N4528, N4505);
or OR3 (N4529, N4520, N3877, N3112);
or OR2 (N4530, N4513, N1636);
nand NAND2 (N4531, N4524, N3439);
nand NAND4 (N4532, N4527, N1502, N1776, N504);
or OR4 (N4533, N4521, N4289, N2451, N2203);
buf BUF1 (N4534, N4530);
nor NOR2 (N4535, N4534, N3333);
not NOT1 (N4536, N4463);
nor NOR4 (N4537, N4528, N331, N114, N221);
buf BUF1 (N4538, N4536);
not NOT1 (N4539, N4531);
or OR4 (N4540, N4516, N747, N2582, N2935);
xor XOR2 (N4541, N4537, N3374);
and AND4 (N4542, N4523, N798, N3764, N1918);
not NOT1 (N4543, N4540);
nor NOR3 (N4544, N4539, N1701, N3154);
or OR2 (N4545, N4532, N401);
nor NOR3 (N4546, N4542, N470, N1071);
not NOT1 (N4547, N4535);
not NOT1 (N4548, N4538);
or OR2 (N4549, N4541, N2380);
not NOT1 (N4550, N4544);
xor XOR2 (N4551, N4543, N1064);
xor XOR2 (N4552, N4550, N2806);
xor XOR2 (N4553, N4545, N3782);
or OR4 (N4554, N4529, N987, N1837, N3176);
nand NAND2 (N4555, N4547, N3900);
xor XOR2 (N4556, N4554, N3276);
and AND3 (N4557, N4548, N1029, N274);
xor XOR2 (N4558, N4533, N2105);
or OR2 (N4559, N4557, N3814);
nor NOR3 (N4560, N4555, N1365, N3942);
or OR2 (N4561, N4526, N3142);
and AND2 (N4562, N4546, N398);
and AND2 (N4563, N4561, N3004);
or OR2 (N4564, N4553, N2728);
xor XOR2 (N4565, N4559, N1369);
or OR3 (N4566, N4563, N3998, N2958);
buf BUF1 (N4567, N4560);
or OR2 (N4568, N4566, N3731);
and AND4 (N4569, N4558, N3001, N4226, N691);
not NOT1 (N4570, N4556);
buf BUF1 (N4571, N4567);
and AND2 (N4572, N4551, N3785);
nand NAND2 (N4573, N4572, N4308);
nor NOR4 (N4574, N4564, N388, N1700, N2220);
nand NAND2 (N4575, N4570, N640);
not NOT1 (N4576, N4569);
xor XOR2 (N4577, N4552, N3694);
buf BUF1 (N4578, N4562);
nand NAND3 (N4579, N4568, N2002, N230);
nor NOR3 (N4580, N4574, N3757, N889);
xor XOR2 (N4581, N4577, N3727);
buf BUF1 (N4582, N4573);
nor NOR2 (N4583, N4580, N3699);
and AND2 (N4584, N4579, N2057);
and AND2 (N4585, N4581, N3739);
buf BUF1 (N4586, N4578);
buf BUF1 (N4587, N4549);
xor XOR2 (N4588, N4575, N3433);
xor XOR2 (N4589, N4582, N4579);
nor NOR4 (N4590, N4583, N4379, N213, N2955);
or OR4 (N4591, N4588, N1856, N1192, N1298);
xor XOR2 (N4592, N4591, N685);
and AND4 (N4593, N4571, N2411, N3412, N2759);
buf BUF1 (N4594, N4589);
nand NAND4 (N4595, N4584, N3551, N3558, N2990);
nor NOR3 (N4596, N4590, N428, N199);
nor NOR2 (N4597, N4596, N2527);
or OR2 (N4598, N4586, N44);
nor NOR4 (N4599, N4576, N32, N3088, N4177);
or OR3 (N4600, N4565, N2586, N1022);
and AND4 (N4601, N4593, N3675, N31, N2928);
buf BUF1 (N4602, N4592);
not NOT1 (N4603, N4585);
and AND2 (N4604, N4595, N2983);
buf BUF1 (N4605, N4594);
nor NOR2 (N4606, N4605, N55);
and AND4 (N4607, N4601, N4142, N987, N3094);
nand NAND4 (N4608, N4600, N8, N1433, N2676);
xor XOR2 (N4609, N4598, N2331);
nor NOR3 (N4610, N4602, N1761, N2072);
buf BUF1 (N4611, N4609);
nand NAND2 (N4612, N4604, N2765);
xor XOR2 (N4613, N4611, N1879);
or OR3 (N4614, N4613, N3966, N2412);
xor XOR2 (N4615, N4612, N334);
nor NOR2 (N4616, N4615, N1898);
xor XOR2 (N4617, N4603, N3838);
or OR2 (N4618, N4587, N1596);
or OR4 (N4619, N4607, N879, N1121, N2573);
nor NOR4 (N4620, N4619, N321, N3643, N410);
or OR2 (N4621, N4606, N2067);
nor NOR4 (N4622, N4610, N3527, N4278, N1061);
xor XOR2 (N4623, N4620, N3237);
buf BUF1 (N4624, N4597);
and AND3 (N4625, N4621, N3992, N2354);
nor NOR4 (N4626, N4616, N2071, N25, N4488);
not NOT1 (N4627, N4618);
buf BUF1 (N4628, N4627);
buf BUF1 (N4629, N4628);
buf BUF1 (N4630, N4599);
buf BUF1 (N4631, N4629);
not NOT1 (N4632, N4631);
nand NAND4 (N4633, N4626, N1993, N3876, N745);
and AND3 (N4634, N4624, N30, N81);
or OR3 (N4635, N4634, N273, N1720);
and AND2 (N4636, N4614, N1513);
nand NAND3 (N4637, N4623, N1845, N917);
nand NAND4 (N4638, N4633, N3261, N4084, N2705);
and AND4 (N4639, N4635, N3435, N2957, N1059);
or OR4 (N4640, N4625, N3785, N2783, N2089);
buf BUF1 (N4641, N4640);
nor NOR4 (N4642, N4630, N304, N164, N2371);
buf BUF1 (N4643, N4637);
buf BUF1 (N4644, N4639);
not NOT1 (N4645, N4632);
buf BUF1 (N4646, N4644);
nand NAND2 (N4647, N4617, N1768);
nand NAND2 (N4648, N4646, N2233);
nand NAND2 (N4649, N4647, N3946);
not NOT1 (N4650, N4636);
buf BUF1 (N4651, N4649);
xor XOR2 (N4652, N4651, N1200);
buf BUF1 (N4653, N4643);
not NOT1 (N4654, N4641);
xor XOR2 (N4655, N4648, N2297);
xor XOR2 (N4656, N4638, N939);
nand NAND3 (N4657, N4650, N805, N206);
xor XOR2 (N4658, N4655, N2496);
xor XOR2 (N4659, N4658, N2505);
nor NOR3 (N4660, N4656, N1239, N957);
xor XOR2 (N4661, N4660, N2599);
and AND3 (N4662, N4608, N2953, N773);
xor XOR2 (N4663, N4642, N2548);
xor XOR2 (N4664, N4663, N1214);
not NOT1 (N4665, N4654);
buf BUF1 (N4666, N4652);
buf BUF1 (N4667, N4622);
nand NAND2 (N4668, N4664, N3870);
not NOT1 (N4669, N4665);
or OR3 (N4670, N4668, N2990, N313);
nor NOR4 (N4671, N4653, N3566, N1476, N982);
nor NOR3 (N4672, N4662, N4488, N1782);
xor XOR2 (N4673, N4669, N3634);
buf BUF1 (N4674, N4670);
not NOT1 (N4675, N4659);
xor XOR2 (N4676, N4661, N906);
xor XOR2 (N4677, N4667, N3056);
or OR4 (N4678, N4676, N1710, N4070, N3765);
xor XOR2 (N4679, N4672, N2575);
or OR2 (N4680, N4657, N1425);
nor NOR4 (N4681, N4671, N3829, N1161, N641);
nor NOR4 (N4682, N4679, N133, N588, N3793);
xor XOR2 (N4683, N4680, N2125);
nand NAND4 (N4684, N4681, N4164, N1263, N857);
xor XOR2 (N4685, N4675, N2337);
xor XOR2 (N4686, N4685, N4066);
xor XOR2 (N4687, N4686, N3770);
and AND4 (N4688, N4684, N4287, N1366, N4574);
buf BUF1 (N4689, N4645);
and AND3 (N4690, N4678, N487, N3300);
not NOT1 (N4691, N4682);
not NOT1 (N4692, N4688);
not NOT1 (N4693, N4692);
and AND4 (N4694, N4689, N1092, N2188, N4399);
or OR3 (N4695, N4691, N1054, N1727);
or OR4 (N4696, N4693, N1869, N996, N1574);
nand NAND3 (N4697, N4673, N2497, N253);
or OR3 (N4698, N4666, N3428, N4483);
or OR2 (N4699, N4674, N604);
or OR2 (N4700, N4694, N1986);
nand NAND3 (N4701, N4687, N219, N692);
and AND2 (N4702, N4683, N103);
nor NOR2 (N4703, N4696, N1861);
not NOT1 (N4704, N4690);
nor NOR2 (N4705, N4702, N41);
and AND3 (N4706, N4695, N2577, N3463);
buf BUF1 (N4707, N4697);
nand NAND4 (N4708, N4699, N416, N1563, N3606);
buf BUF1 (N4709, N4701);
or OR3 (N4710, N4705, N2027, N2749);
buf BUF1 (N4711, N4677);
or OR3 (N4712, N4709, N218, N3328);
xor XOR2 (N4713, N4700, N1270);
buf BUF1 (N4714, N4713);
and AND3 (N4715, N4703, N1283, N1246);
xor XOR2 (N4716, N4711, N1122);
not NOT1 (N4717, N4710);
not NOT1 (N4718, N4706);
nor NOR3 (N4719, N4698, N2966, N1799);
buf BUF1 (N4720, N4707);
xor XOR2 (N4721, N4716, N2448);
and AND2 (N4722, N4718, N1624);
and AND4 (N4723, N4719, N485, N114, N880);
nor NOR4 (N4724, N4714, N2457, N686, N3861);
xor XOR2 (N4725, N4712, N2939);
nand NAND4 (N4726, N4723, N3735, N4335, N1192);
nand NAND4 (N4727, N4725, N3948, N4224, N3230);
xor XOR2 (N4728, N4724, N670);
xor XOR2 (N4729, N4715, N1233);
and AND3 (N4730, N4729, N844, N341);
nor NOR4 (N4731, N4708, N346, N389, N4687);
not NOT1 (N4732, N4726);
nor NOR2 (N4733, N4727, N2809);
buf BUF1 (N4734, N4720);
and AND2 (N4735, N4731, N1673);
and AND2 (N4736, N4735, N4324);
xor XOR2 (N4737, N4730, N4473);
nand NAND3 (N4738, N4734, N2608, N1277);
buf BUF1 (N4739, N4704);
not NOT1 (N4740, N4737);
not NOT1 (N4741, N4740);
not NOT1 (N4742, N4736);
nand NAND2 (N4743, N4739, N2436);
not NOT1 (N4744, N4742);
or OR2 (N4745, N4744, N4628);
nand NAND2 (N4746, N4741, N1707);
nand NAND4 (N4747, N4721, N2361, N2517, N818);
and AND3 (N4748, N4728, N2224, N1653);
and AND2 (N4749, N4738, N2160);
nor NOR2 (N4750, N4717, N2687);
not NOT1 (N4751, N4749);
not NOT1 (N4752, N4722);
nand NAND2 (N4753, N4748, N2443);
not NOT1 (N4754, N4752);
xor XOR2 (N4755, N4746, N3304);
nand NAND2 (N4756, N4745, N2286);
xor XOR2 (N4757, N4743, N109);
xor XOR2 (N4758, N4751, N2999);
not NOT1 (N4759, N4756);
nor NOR3 (N4760, N4759, N3972, N4387);
or OR3 (N4761, N4750, N2540, N1467);
not NOT1 (N4762, N4758);
xor XOR2 (N4763, N4755, N4407);
and AND3 (N4764, N4732, N2057, N3050);
xor XOR2 (N4765, N4763, N2991);
and AND4 (N4766, N4753, N2116, N4709, N3707);
xor XOR2 (N4767, N4733, N4308);
buf BUF1 (N4768, N4766);
xor XOR2 (N4769, N4764, N3923);
buf BUF1 (N4770, N4762);
not NOT1 (N4771, N4770);
nand NAND4 (N4772, N4757, N4071, N4251, N2345);
xor XOR2 (N4773, N4771, N2232);
nand NAND3 (N4774, N4754, N1439, N3489);
buf BUF1 (N4775, N4772);
nand NAND4 (N4776, N4768, N3429, N1209, N2440);
xor XOR2 (N4777, N4775, N1269);
and AND3 (N4778, N4760, N3419, N3610);
nor NOR2 (N4779, N4761, N423);
not NOT1 (N4780, N4773);
xor XOR2 (N4781, N4767, N1198);
buf BUF1 (N4782, N4776);
xor XOR2 (N4783, N4769, N1578);
buf BUF1 (N4784, N4778);
or OR4 (N4785, N4779, N4722, N3082, N2850);
not NOT1 (N4786, N4774);
or OR2 (N4787, N4777, N3887);
or OR2 (N4788, N4780, N277);
nor NOR4 (N4789, N4785, N2746, N969, N2423);
nand NAND2 (N4790, N4787, N553);
not NOT1 (N4791, N4786);
xor XOR2 (N4792, N4791, N3325);
buf BUF1 (N4793, N4788);
or OR4 (N4794, N4789, N3927, N2701, N1210);
nand NAND3 (N4795, N4792, N770, N2002);
nand NAND4 (N4796, N4783, N246, N1432, N645);
not NOT1 (N4797, N4747);
and AND4 (N4798, N4794, N1500, N861, N115);
buf BUF1 (N4799, N4790);
nand NAND4 (N4800, N4782, N3808, N3088, N4538);
or OR2 (N4801, N4784, N62);
not NOT1 (N4802, N4781);
or OR4 (N4803, N4798, N1914, N2943, N1624);
or OR2 (N4804, N4795, N3954);
and AND3 (N4805, N4800, N2158, N112);
nand NAND3 (N4806, N4801, N1611, N4769);
buf BUF1 (N4807, N4806);
nand NAND2 (N4808, N4799, N3717);
xor XOR2 (N4809, N4793, N1618);
or OR2 (N4810, N4809, N3459);
nand NAND4 (N4811, N4796, N3863, N172, N2240);
nand NAND4 (N4812, N4807, N2739, N3276, N3796);
nand NAND2 (N4813, N4810, N3326);
not NOT1 (N4814, N4803);
xor XOR2 (N4815, N4811, N2976);
or OR4 (N4816, N4813, N1545, N3981, N3537);
nor NOR2 (N4817, N4815, N3586);
xor XOR2 (N4818, N4802, N1042);
nand NAND2 (N4819, N4812, N2004);
buf BUF1 (N4820, N4817);
buf BUF1 (N4821, N4818);
buf BUF1 (N4822, N4819);
or OR2 (N4823, N4804, N1639);
not NOT1 (N4824, N4808);
nor NOR4 (N4825, N4822, N4619, N3183, N1181);
nand NAND3 (N4826, N4820, N4548, N440);
not NOT1 (N4827, N4824);
nand NAND4 (N4828, N4797, N539, N3650, N123);
not NOT1 (N4829, N4805);
xor XOR2 (N4830, N4828, N348);
nand NAND4 (N4831, N4821, N4301, N2871, N2981);
nor NOR4 (N4832, N4829, N937, N1452, N852);
xor XOR2 (N4833, N4831, N378);
and AND4 (N4834, N4814, N3589, N1354, N2416);
not NOT1 (N4835, N4826);
not NOT1 (N4836, N4765);
nor NOR2 (N4837, N4835, N1361);
not NOT1 (N4838, N4830);
nor NOR2 (N4839, N4838, N405);
nand NAND4 (N4840, N4816, N442, N2083, N4278);
nand NAND3 (N4841, N4833, N613, N2193);
not NOT1 (N4842, N4825);
xor XOR2 (N4843, N4839, N1130);
or OR4 (N4844, N4823, N3070, N2308, N1161);
nand NAND2 (N4845, N4840, N2739);
not NOT1 (N4846, N4832);
nand NAND4 (N4847, N4836, N4800, N4507, N867);
nand NAND2 (N4848, N4843, N2083);
or OR4 (N4849, N4841, N1232, N3243, N3736);
xor XOR2 (N4850, N4845, N534);
nor NOR2 (N4851, N4827, N1013);
nand NAND4 (N4852, N4837, N3378, N3409, N3941);
xor XOR2 (N4853, N4850, N4076);
not NOT1 (N4854, N4853);
nand NAND4 (N4855, N4844, N1927, N3898, N5);
not NOT1 (N4856, N4854);
nand NAND4 (N4857, N4856, N2935, N1285, N328);
not NOT1 (N4858, N4855);
not NOT1 (N4859, N4834);
and AND2 (N4860, N4849, N1609);
nand NAND3 (N4861, N4848, N1620, N652);
xor XOR2 (N4862, N4847, N3851);
nand NAND4 (N4863, N4851, N3873, N3861, N338);
nand NAND4 (N4864, N4863, N2877, N3470, N1497);
xor XOR2 (N4865, N4842, N3700);
nand NAND4 (N4866, N4865, N2920, N2190, N3005);
not NOT1 (N4867, N4861);
xor XOR2 (N4868, N4852, N3449);
not NOT1 (N4869, N4862);
nor NOR4 (N4870, N4859, N2903, N3025, N3957);
nand NAND4 (N4871, N4864, N1545, N3569, N3473);
nand NAND2 (N4872, N4869, N4156);
or OR2 (N4873, N4860, N4765);
not NOT1 (N4874, N4870);
nand NAND3 (N4875, N4872, N4139, N3708);
nor NOR3 (N4876, N4867, N254, N4830);
nor NOR4 (N4877, N4858, N2536, N3610, N4775);
xor XOR2 (N4878, N4846, N1863);
nor NOR2 (N4879, N4873, N1089);
nor NOR3 (N4880, N4875, N4263, N136);
buf BUF1 (N4881, N4868);
buf BUF1 (N4882, N4878);
buf BUF1 (N4883, N4871);
or OR4 (N4884, N4876, N1063, N340, N618);
not NOT1 (N4885, N4884);
or OR2 (N4886, N4879, N4748);
not NOT1 (N4887, N4880);
xor XOR2 (N4888, N4885, N277);
xor XOR2 (N4889, N4883, N3174);
xor XOR2 (N4890, N4886, N2105);
or OR2 (N4891, N4888, N1314);
or OR2 (N4892, N4891, N2645);
nand NAND2 (N4893, N4890, N3017);
buf BUF1 (N4894, N4881);
and AND4 (N4895, N4857, N4540, N3406, N1035);
and AND3 (N4896, N4882, N2857, N2619);
not NOT1 (N4897, N4866);
xor XOR2 (N4898, N4895, N1869);
buf BUF1 (N4899, N4887);
buf BUF1 (N4900, N4896);
nor NOR4 (N4901, N4900, N2924, N550, N3727);
buf BUF1 (N4902, N4892);
buf BUF1 (N4903, N4897);
and AND3 (N4904, N4874, N3072, N12);
nand NAND4 (N4905, N4898, N512, N4456, N1458);
nand NAND4 (N4906, N4902, N2369, N1356, N4799);
or OR3 (N4907, N4904, N2024, N4209);
and AND2 (N4908, N4903, N720);
not NOT1 (N4909, N4906);
nor NOR4 (N4910, N4899, N3629, N36, N86);
or OR2 (N4911, N4909, N2705);
not NOT1 (N4912, N4905);
nand NAND4 (N4913, N4911, N2476, N2343, N3238);
nand NAND3 (N4914, N4893, N3454, N4315);
nand NAND3 (N4915, N4908, N3631, N4326);
not NOT1 (N4916, N4889);
xor XOR2 (N4917, N4877, N3337);
nor NOR2 (N4918, N4915, N3014);
buf BUF1 (N4919, N4914);
not NOT1 (N4920, N4913);
or OR3 (N4921, N4910, N1117, N3765);
not NOT1 (N4922, N4920);
nor NOR4 (N4923, N4907, N468, N1904, N3974);
nor NOR2 (N4924, N4919, N4708);
xor XOR2 (N4925, N4916, N2306);
not NOT1 (N4926, N4918);
nor NOR3 (N4927, N4924, N1914, N1708);
or OR3 (N4928, N4926, N4927, N2638);
and AND4 (N4929, N2056, N870, N1703, N2416);
and AND2 (N4930, N4925, N4260);
nor NOR2 (N4931, N4922, N584);
buf BUF1 (N4932, N4917);
nand NAND4 (N4933, N4932, N1432, N4707, N3299);
nor NOR4 (N4934, N4931, N4471, N2747, N4604);
and AND3 (N4935, N4930, N4349, N403);
buf BUF1 (N4936, N4929);
xor XOR2 (N4937, N4928, N3531);
buf BUF1 (N4938, N4921);
or OR2 (N4939, N4936, N4097);
nor NOR4 (N4940, N4937, N2401, N4145, N915);
nor NOR2 (N4941, N4933, N3312);
and AND4 (N4942, N4941, N1519, N4131, N1850);
xor XOR2 (N4943, N4894, N4578);
buf BUF1 (N4944, N4912);
not NOT1 (N4945, N4943);
or OR4 (N4946, N4940, N3059, N1532, N3629);
buf BUF1 (N4947, N4935);
buf BUF1 (N4948, N4947);
xor XOR2 (N4949, N4942, N3382);
not NOT1 (N4950, N4938);
nor NOR4 (N4951, N4944, N261, N2178, N3059);
buf BUF1 (N4952, N4945);
and AND3 (N4953, N4946, N2211, N1575);
not NOT1 (N4954, N4901);
not NOT1 (N4955, N4934);
and AND3 (N4956, N4949, N2014, N534);
or OR2 (N4957, N4950, N3336);
buf BUF1 (N4958, N4952);
buf BUF1 (N4959, N4958);
nor NOR3 (N4960, N4957, N4218, N206);
not NOT1 (N4961, N4956);
buf BUF1 (N4962, N4959);
or OR2 (N4963, N4953, N4896);
and AND4 (N4964, N4960, N1801, N4254, N1822);
nand NAND2 (N4965, N4955, N349);
nand NAND2 (N4966, N4948, N2049);
and AND4 (N4967, N4963, N2693, N4608, N2938);
buf BUF1 (N4968, N4964);
nor NOR4 (N4969, N4923, N3485, N953, N2177);
nand NAND2 (N4970, N4966, N1699);
not NOT1 (N4971, N4954);
buf BUF1 (N4972, N4967);
xor XOR2 (N4973, N4968, N3186);
nand NAND3 (N4974, N4969, N2440, N600);
not NOT1 (N4975, N4971);
buf BUF1 (N4976, N4965);
xor XOR2 (N4977, N4939, N558);
nor NOR4 (N4978, N4973, N2175, N1248, N2088);
xor XOR2 (N4979, N4977, N3355);
nand NAND2 (N4980, N4951, N1206);
nand NAND3 (N4981, N4972, N2971, N2886);
not NOT1 (N4982, N4981);
nor NOR3 (N4983, N4974, N2429, N2605);
and AND3 (N4984, N4970, N3148, N1488);
and AND3 (N4985, N4979, N437, N3842);
and AND2 (N4986, N4962, N2307);
nand NAND4 (N4987, N4976, N1370, N1350, N3643);
xor XOR2 (N4988, N4986, N3079);
or OR3 (N4989, N4985, N3009, N2245);
buf BUF1 (N4990, N4988);
not NOT1 (N4991, N4961);
and AND4 (N4992, N4975, N4610, N2218, N3520);
nand NAND4 (N4993, N4989, N922, N450, N2522);
nand NAND2 (N4994, N4982, N4808);
nand NAND2 (N4995, N4992, N4976);
nand NAND4 (N4996, N4991, N3286, N3464, N713);
and AND4 (N4997, N4987, N1456, N3104, N831);
and AND2 (N4998, N4978, N369);
nand NAND2 (N4999, N4983, N1861);
or OR2 (N5000, N4997, N25);
or OR3 (N5001, N4984, N2871, N4274);
nor NOR2 (N5002, N4994, N4218);
xor XOR2 (N5003, N5001, N1973);
nand NAND3 (N5004, N4980, N663, N4618);
nand NAND4 (N5005, N5000, N3324, N3954, N2621);
and AND3 (N5006, N5003, N2978, N1590);
xor XOR2 (N5007, N4999, N3867);
buf BUF1 (N5008, N4998);
or OR3 (N5009, N4990, N4481, N4148);
not NOT1 (N5010, N5002);
nand NAND3 (N5011, N5007, N4376, N807);
nand NAND2 (N5012, N5005, N1775);
or OR4 (N5013, N5009, N4282, N3583, N2287);
nand NAND2 (N5014, N4995, N1522);
or OR4 (N5015, N5013, N4289, N3103, N3455);
nor NOR2 (N5016, N5010, N2621);
nor NOR2 (N5017, N5014, N3763);
buf BUF1 (N5018, N5015);
xor XOR2 (N5019, N4996, N2562);
and AND3 (N5020, N5019, N2949, N3883);
nand NAND3 (N5021, N5018, N990, N2222);
not NOT1 (N5022, N5004);
nor NOR3 (N5023, N5017, N4166, N2130);
and AND4 (N5024, N5006, N4135, N2010, N2331);
and AND2 (N5025, N5022, N2529);
or OR4 (N5026, N5020, N1589, N3633, N4596);
xor XOR2 (N5027, N5024, N997);
or OR2 (N5028, N5011, N1750);
nand NAND3 (N5029, N5023, N4369, N3539);
xor XOR2 (N5030, N5016, N4501);
nor NOR3 (N5031, N5025, N1597, N1666);
nand NAND4 (N5032, N5027, N3865, N2377, N2884);
nand NAND3 (N5033, N5021, N3007, N4223);
and AND4 (N5034, N4993, N4024, N815, N440);
or OR3 (N5035, N5029, N4092, N4719);
nand NAND3 (N5036, N5035, N3782, N362);
xor XOR2 (N5037, N5032, N2270);
not NOT1 (N5038, N5031);
buf BUF1 (N5039, N5028);
xor XOR2 (N5040, N5033, N2993);
buf BUF1 (N5041, N5034);
nor NOR2 (N5042, N5040, N995);
and AND2 (N5043, N5042, N2828);
nand NAND2 (N5044, N5043, N3927);
nand NAND2 (N5045, N5030, N4402);
xor XOR2 (N5046, N5039, N1287);
xor XOR2 (N5047, N5044, N3567);
nor NOR4 (N5048, N5008, N2378, N1215, N1302);
nor NOR4 (N5049, N5012, N5019, N748, N1911);
nand NAND4 (N5050, N5041, N1484, N2729, N276);
buf BUF1 (N5051, N5050);
not NOT1 (N5052, N5038);
nor NOR2 (N5053, N5047, N4079);
not NOT1 (N5054, N5052);
xor XOR2 (N5055, N5053, N2500);
not NOT1 (N5056, N5045);
not NOT1 (N5057, N5055);
nand NAND4 (N5058, N5048, N2279, N4264, N2221);
and AND3 (N5059, N5058, N3912, N399);
or OR2 (N5060, N5059, N4416);
nor NOR4 (N5061, N5057, N3295, N3065, N1119);
nand NAND2 (N5062, N5049, N660);
and AND4 (N5063, N5061, N1251, N5017, N3209);
not NOT1 (N5064, N5060);
buf BUF1 (N5065, N5063);
nand NAND3 (N5066, N5046, N3129, N1801);
and AND3 (N5067, N5066, N2411, N3750);
nor NOR4 (N5068, N5067, N1257, N2900, N3518);
xor XOR2 (N5069, N5037, N225);
or OR3 (N5070, N5054, N2850, N2962);
or OR2 (N5071, N5026, N3097);
not NOT1 (N5072, N5070);
not NOT1 (N5073, N5036);
or OR4 (N5074, N5068, N4723, N412, N4054);
not NOT1 (N5075, N5056);
nand NAND4 (N5076, N5069, N446, N3025, N3567);
xor XOR2 (N5077, N5062, N2722);
buf BUF1 (N5078, N5076);
xor XOR2 (N5079, N5071, N166);
or OR3 (N5080, N5065, N2498, N3846);
and AND2 (N5081, N5079, N2422);
or OR3 (N5082, N5081, N611, N3423);
xor XOR2 (N5083, N5073, N3548);
nor NOR3 (N5084, N5074, N4075, N942);
xor XOR2 (N5085, N5075, N1920);
or OR4 (N5086, N5084, N4089, N5041, N3899);
nand NAND2 (N5087, N5072, N3836);
buf BUF1 (N5088, N5078);
xor XOR2 (N5089, N5077, N1656);
nor NOR2 (N5090, N5051, N347);
nand NAND2 (N5091, N5080, N2164);
and AND3 (N5092, N5091, N4634, N2143);
or OR3 (N5093, N5089, N2989, N1067);
and AND3 (N5094, N5064, N3427, N2944);
not NOT1 (N5095, N5088);
not NOT1 (N5096, N5086);
buf BUF1 (N5097, N5087);
buf BUF1 (N5098, N5095);
nand NAND4 (N5099, N5096, N2456, N4065, N2379);
and AND4 (N5100, N5090, N496, N4807, N4580);
nor NOR3 (N5101, N5082, N751, N1671);
nand NAND3 (N5102, N5092, N1978, N174);
nand NAND3 (N5103, N5083, N224, N4245);
buf BUF1 (N5104, N5098);
or OR2 (N5105, N5102, N2267);
nor NOR4 (N5106, N5100, N4441, N118, N4746);
or OR3 (N5107, N5103, N2249, N672);
buf BUF1 (N5108, N5097);
nand NAND2 (N5109, N5104, N963);
and AND4 (N5110, N5093, N1261, N1086, N4637);
xor XOR2 (N5111, N5099, N3743);
and AND2 (N5112, N5094, N1144);
and AND2 (N5113, N5105, N3675);
xor XOR2 (N5114, N5109, N4813);
nor NOR3 (N5115, N5106, N4799, N2988);
nand NAND4 (N5116, N5108, N3382, N3339, N4751);
buf BUF1 (N5117, N5111);
nand NAND4 (N5118, N5110, N3183, N3734, N3667);
and AND3 (N5119, N5112, N3082, N3029);
and AND3 (N5120, N5101, N4543, N3850);
xor XOR2 (N5121, N5117, N2277);
not NOT1 (N5122, N5116);
nor NOR2 (N5123, N5085, N2811);
and AND2 (N5124, N5113, N4720);
or OR2 (N5125, N5114, N152);
not NOT1 (N5126, N5123);
nand NAND2 (N5127, N5126, N2838);
and AND4 (N5128, N5124, N2922, N191, N1231);
nor NOR4 (N5129, N5107, N904, N2966, N1487);
or OR3 (N5130, N5115, N2981, N2863);
nor NOR2 (N5131, N5128, N2023);
nor NOR3 (N5132, N5118, N854, N4109);
nor NOR2 (N5133, N5119, N4210);
xor XOR2 (N5134, N5131, N5080);
buf BUF1 (N5135, N5130);
and AND2 (N5136, N5125, N2457);
xor XOR2 (N5137, N5120, N2074);
nor NOR3 (N5138, N5122, N851, N3710);
xor XOR2 (N5139, N5127, N4970);
and AND3 (N5140, N5135, N3976, N4912);
nand NAND2 (N5141, N5133, N2104);
xor XOR2 (N5142, N5137, N3184);
or OR2 (N5143, N5132, N3796);
nand NAND4 (N5144, N5129, N4659, N2820, N2534);
and AND2 (N5145, N5141, N1016);
or OR3 (N5146, N5142, N681, N1275);
or OR4 (N5147, N5138, N3217, N236, N3217);
nand NAND3 (N5148, N5134, N4684, N4380);
and AND3 (N5149, N5144, N3909, N684);
or OR4 (N5150, N5139, N3734, N428, N4342);
and AND3 (N5151, N5121, N595, N2593);
not NOT1 (N5152, N5148);
buf BUF1 (N5153, N5140);
nand NAND3 (N5154, N5151, N1382, N4661);
not NOT1 (N5155, N5150);
or OR3 (N5156, N5153, N5007, N693);
or OR2 (N5157, N5154, N1513);
xor XOR2 (N5158, N5146, N134);
nand NAND4 (N5159, N5156, N318, N4250, N1788);
xor XOR2 (N5160, N5152, N1595);
xor XOR2 (N5161, N5149, N3969);
or OR2 (N5162, N5161, N1390);
not NOT1 (N5163, N5155);
buf BUF1 (N5164, N5136);
buf BUF1 (N5165, N5163);
and AND4 (N5166, N5162, N4916, N830, N3933);
nand NAND4 (N5167, N5157, N2696, N4381, N725);
nand NAND2 (N5168, N5166, N2209);
xor XOR2 (N5169, N5145, N4097);
nor NOR4 (N5170, N5164, N1442, N4129, N2422);
nor NOR4 (N5171, N5160, N3471, N2029, N4434);
xor XOR2 (N5172, N5169, N62);
nand NAND2 (N5173, N5172, N3946);
nand NAND3 (N5174, N5143, N3374, N251);
nor NOR4 (N5175, N5170, N3192, N3282, N4914);
buf BUF1 (N5176, N5171);
or OR2 (N5177, N5167, N904);
nand NAND3 (N5178, N5147, N1587, N2841);
and AND2 (N5179, N5177, N1715);
nor NOR2 (N5180, N5158, N2894);
and AND4 (N5181, N5179, N1847, N3311, N4821);
nor NOR4 (N5182, N5175, N4054, N3669, N1470);
or OR3 (N5183, N5178, N4593, N1537);
nor NOR2 (N5184, N5176, N5032);
and AND2 (N5185, N5174, N4407);
or OR3 (N5186, N5183, N2752, N3230);
buf BUF1 (N5187, N5180);
and AND4 (N5188, N5165, N1236, N5109, N2047);
or OR3 (N5189, N5188, N482, N4971);
nor NOR3 (N5190, N5181, N3625, N2526);
and AND4 (N5191, N5187, N3573, N2158, N142);
not NOT1 (N5192, N5184);
or OR4 (N5193, N5189, N216, N3245, N3037);
nand NAND4 (N5194, N5193, N3862, N1780, N5109);
and AND4 (N5195, N5191, N3102, N5016, N2252);
or OR4 (N5196, N5192, N4774, N5167, N5014);
nor NOR2 (N5197, N5190, N691);
xor XOR2 (N5198, N5186, N4661);
not NOT1 (N5199, N5196);
nand NAND3 (N5200, N5197, N4340, N4410);
nor NOR4 (N5201, N5198, N3095, N2011, N3181);
nand NAND4 (N5202, N5185, N1195, N3613, N1890);
and AND3 (N5203, N5194, N116, N2796);
buf BUF1 (N5204, N5200);
xor XOR2 (N5205, N5201, N4155);
xor XOR2 (N5206, N5203, N3954);
and AND4 (N5207, N5204, N3877, N3692, N1903);
not NOT1 (N5208, N5182);
nor NOR2 (N5209, N5208, N3486);
or OR2 (N5210, N5173, N3897);
and AND2 (N5211, N5207, N1426);
xor XOR2 (N5212, N5206, N907);
not NOT1 (N5213, N5168);
and AND2 (N5214, N5202, N3846);
not NOT1 (N5215, N5214);
xor XOR2 (N5216, N5205, N3574);
nand NAND4 (N5217, N5210, N3704, N3880, N82);
not NOT1 (N5218, N5217);
nand NAND4 (N5219, N5159, N3000, N1385, N2851);
nand NAND2 (N5220, N5209, N5098);
and AND2 (N5221, N5211, N4690);
nor NOR4 (N5222, N5216, N3412, N2065, N501);
not NOT1 (N5223, N5219);
buf BUF1 (N5224, N5221);
nor NOR2 (N5225, N5218, N3771);
and AND4 (N5226, N5195, N1974, N4137, N3657);
or OR4 (N5227, N5226, N3559, N1018, N4572);
or OR2 (N5228, N5215, N423);
and AND2 (N5229, N5223, N2011);
and AND2 (N5230, N5222, N1684);
or OR3 (N5231, N5212, N4734, N1574);
not NOT1 (N5232, N5224);
nor NOR3 (N5233, N5213, N3276, N4542);
and AND4 (N5234, N5227, N288, N5106, N4437);
not NOT1 (N5235, N5234);
not NOT1 (N5236, N5230);
xor XOR2 (N5237, N5199, N2128);
not NOT1 (N5238, N5231);
nor NOR4 (N5239, N5233, N1093, N915, N2559);
or OR3 (N5240, N5228, N3257, N5166);
nand NAND4 (N5241, N5232, N2841, N3917, N4702);
nand NAND2 (N5242, N5236, N223);
nand NAND4 (N5243, N5235, N619, N4971, N2736);
or OR4 (N5244, N5229, N1759, N4380, N4393);
buf BUF1 (N5245, N5241);
nand NAND4 (N5246, N5237, N2443, N323, N3935);
buf BUF1 (N5247, N5225);
nor NOR4 (N5248, N5239, N2295, N3155, N2156);
or OR4 (N5249, N5238, N4713, N1300, N4181);
nand NAND4 (N5250, N5248, N303, N4040, N1198);
xor XOR2 (N5251, N5243, N674);
or OR4 (N5252, N5220, N3935, N1701, N762);
buf BUF1 (N5253, N5240);
xor XOR2 (N5254, N5242, N4406);
nand NAND4 (N5255, N5250, N4062, N2127, N2723);
xor XOR2 (N5256, N5253, N2586);
and AND4 (N5257, N5245, N2911, N443, N3548);
not NOT1 (N5258, N5247);
nor NOR4 (N5259, N5249, N5144, N3957, N4630);
nand NAND2 (N5260, N5256, N4797);
nand NAND3 (N5261, N5259, N2542, N817);
not NOT1 (N5262, N5251);
xor XOR2 (N5263, N5261, N4420);
or OR3 (N5264, N5263, N1489, N4234);
not NOT1 (N5265, N5244);
xor XOR2 (N5266, N5254, N1944);
not NOT1 (N5267, N5246);
not NOT1 (N5268, N5258);
xor XOR2 (N5269, N5268, N3162);
nor NOR4 (N5270, N5252, N2121, N2363, N5118);
and AND2 (N5271, N5266, N291);
buf BUF1 (N5272, N5262);
nand NAND3 (N5273, N5265, N3982, N4554);
nor NOR2 (N5274, N5273, N468);
nor NOR4 (N5275, N5264, N2363, N952, N4830);
or OR4 (N5276, N5257, N3448, N2512, N1588);
not NOT1 (N5277, N5260);
buf BUF1 (N5278, N5255);
nor NOR3 (N5279, N5275, N519, N3646);
and AND4 (N5280, N5276, N3877, N2240, N1360);
nor NOR4 (N5281, N5280, N3834, N5062, N947);
not NOT1 (N5282, N5274);
nor NOR2 (N5283, N5270, N2007);
not NOT1 (N5284, N5281);
not NOT1 (N5285, N5278);
nand NAND3 (N5286, N5284, N125, N4135);
xor XOR2 (N5287, N5271, N906);
buf BUF1 (N5288, N5272);
xor XOR2 (N5289, N5286, N4736);
nand NAND4 (N5290, N5282, N145, N87, N3702);
xor XOR2 (N5291, N5289, N5193);
nand NAND2 (N5292, N5291, N3979);
buf BUF1 (N5293, N5269);
nor NOR3 (N5294, N5277, N2038, N5020);
xor XOR2 (N5295, N5290, N945);
and AND3 (N5296, N5283, N4701, N4488);
or OR4 (N5297, N5288, N1800, N963, N884);
and AND2 (N5298, N5297, N5047);
and AND3 (N5299, N5267, N462, N3554);
or OR2 (N5300, N5279, N1945);
nor NOR4 (N5301, N5298, N5177, N4450, N820);
and AND2 (N5302, N5285, N3734);
and AND4 (N5303, N5296, N1744, N438, N905);
and AND4 (N5304, N5295, N1396, N2569, N2322);
nor NOR2 (N5305, N5301, N3084);
nand NAND2 (N5306, N5302, N3785);
nand NAND4 (N5307, N5294, N2855, N1275, N4614);
nor NOR3 (N5308, N5292, N3702, N3326);
nand NAND3 (N5309, N5300, N42, N1298);
xor XOR2 (N5310, N5303, N2841);
xor XOR2 (N5311, N5307, N2806);
and AND4 (N5312, N5293, N4852, N4685, N2912);
or OR4 (N5313, N5308, N4733, N2567, N2361);
xor XOR2 (N5314, N5305, N3785);
or OR3 (N5315, N5309, N1326, N2125);
buf BUF1 (N5316, N5304);
nand NAND4 (N5317, N5314, N4457, N315, N3623);
nor NOR4 (N5318, N5317, N1005, N126, N110);
nor NOR4 (N5319, N5318, N1644, N5162, N4696);
nor NOR3 (N5320, N5315, N3898, N1480);
or OR2 (N5321, N5319, N2483);
not NOT1 (N5322, N5306);
nor NOR2 (N5323, N5287, N639);
xor XOR2 (N5324, N5323, N1187);
not NOT1 (N5325, N5322);
nor NOR3 (N5326, N5310, N1377, N1760);
not NOT1 (N5327, N5320);
buf BUF1 (N5328, N5311);
nand NAND2 (N5329, N5316, N38);
buf BUF1 (N5330, N5325);
buf BUF1 (N5331, N5327);
not NOT1 (N5332, N5330);
and AND3 (N5333, N5331, N5047, N3185);
not NOT1 (N5334, N5332);
or OR3 (N5335, N5326, N1887, N4721);
and AND2 (N5336, N5335, N3915);
not NOT1 (N5337, N5328);
or OR2 (N5338, N5324, N2403);
nor NOR4 (N5339, N5338, N1956, N5046, N2654);
or OR4 (N5340, N5299, N5034, N1509, N541);
xor XOR2 (N5341, N5336, N3839);
not NOT1 (N5342, N5333);
xor XOR2 (N5343, N5341, N159);
nand NAND2 (N5344, N5329, N1432);
xor XOR2 (N5345, N5321, N876);
xor XOR2 (N5346, N5340, N3872);
or OR3 (N5347, N5339, N1319, N4287);
buf BUF1 (N5348, N5344);
or OR2 (N5349, N5334, N524);
not NOT1 (N5350, N5313);
not NOT1 (N5351, N5347);
not NOT1 (N5352, N5345);
nand NAND2 (N5353, N5337, N2745);
nand NAND4 (N5354, N5343, N2132, N3538, N1562);
not NOT1 (N5355, N5349);
nand NAND4 (N5356, N5351, N1266, N2394, N1740);
or OR4 (N5357, N5354, N3546, N148, N1871);
nand NAND2 (N5358, N5355, N2811);
buf BUF1 (N5359, N5358);
nor NOR2 (N5360, N5357, N3854);
or OR2 (N5361, N5360, N2829);
xor XOR2 (N5362, N5352, N1946);
buf BUF1 (N5363, N5312);
nand NAND3 (N5364, N5346, N1319, N3731);
or OR4 (N5365, N5342, N1541, N122, N2121);
and AND2 (N5366, N5350, N2378);
not NOT1 (N5367, N5353);
nor NOR2 (N5368, N5362, N1014);
nand NAND4 (N5369, N5368, N2022, N2331, N4466);
not NOT1 (N5370, N5366);
nand NAND4 (N5371, N5356, N3191, N4096, N4142);
buf BUF1 (N5372, N5371);
or OR4 (N5373, N5372, N3407, N4196, N3974);
nand NAND4 (N5374, N5373, N2186, N42, N646);
nand NAND3 (N5375, N5369, N3136, N393);
nand NAND4 (N5376, N5361, N4730, N2419, N4027);
nand NAND4 (N5377, N5364, N5054, N1148, N2614);
or OR3 (N5378, N5348, N2709, N3525);
buf BUF1 (N5379, N5367);
and AND4 (N5380, N5377, N3967, N1919, N1157);
nor NOR4 (N5381, N5370, N1396, N1295, N3488);
nor NOR2 (N5382, N5375, N1962);
or OR4 (N5383, N5359, N1931, N3085, N2688);
or OR4 (N5384, N5363, N1976, N2180, N4659);
or OR3 (N5385, N5380, N1771, N2632);
buf BUF1 (N5386, N5374);
or OR4 (N5387, N5385, N1590, N4656, N205);
nor NOR4 (N5388, N5378, N3765, N1026, N3460);
xor XOR2 (N5389, N5365, N4188);
not NOT1 (N5390, N5387);
xor XOR2 (N5391, N5386, N4167);
xor XOR2 (N5392, N5389, N1732);
not NOT1 (N5393, N5390);
xor XOR2 (N5394, N5392, N2532);
nor NOR2 (N5395, N5394, N111);
nor NOR4 (N5396, N5381, N4000, N2294, N4981);
nand NAND3 (N5397, N5376, N4710, N4378);
buf BUF1 (N5398, N5379);
nand NAND4 (N5399, N5382, N113, N1020, N336);
buf BUF1 (N5400, N5393);
not NOT1 (N5401, N5391);
nor NOR3 (N5402, N5400, N4119, N4593);
and AND4 (N5403, N5398, N4495, N4924, N1431);
or OR4 (N5404, N5401, N288, N1357, N3775);
not NOT1 (N5405, N5404);
not NOT1 (N5406, N5399);
not NOT1 (N5407, N5388);
not NOT1 (N5408, N5396);
or OR4 (N5409, N5402, N3214, N959, N4414);
nand NAND2 (N5410, N5383, N41);
and AND4 (N5411, N5409, N4293, N1411, N1980);
and AND2 (N5412, N5384, N4435);
buf BUF1 (N5413, N5411);
xor XOR2 (N5414, N5412, N2897);
buf BUF1 (N5415, N5406);
not NOT1 (N5416, N5395);
nand NAND4 (N5417, N5403, N2402, N3764, N3164);
or OR4 (N5418, N5410, N4294, N4796, N3685);
nand NAND3 (N5419, N5414, N3294, N2555);
buf BUF1 (N5420, N5417);
nand NAND3 (N5421, N5408, N4698, N1752);
nor NOR2 (N5422, N5418, N3340);
nand NAND4 (N5423, N5407, N2167, N1500, N3282);
nor NOR4 (N5424, N5422, N1097, N506, N268);
xor XOR2 (N5425, N5416, N3177);
not NOT1 (N5426, N5425);
buf BUF1 (N5427, N5420);
xor XOR2 (N5428, N5413, N737);
and AND3 (N5429, N5415, N4533, N2922);
nand NAND4 (N5430, N5428, N3691, N4470, N4575);
not NOT1 (N5431, N5397);
not NOT1 (N5432, N5426);
xor XOR2 (N5433, N5431, N1995);
nand NAND2 (N5434, N5433, N1116);
nand NAND3 (N5435, N5429, N1423, N1504);
nor NOR3 (N5436, N5405, N4535, N4736);
or OR4 (N5437, N5432, N597, N4542, N4678);
not NOT1 (N5438, N5430);
xor XOR2 (N5439, N5421, N2077);
and AND3 (N5440, N5438, N877, N951);
buf BUF1 (N5441, N5435);
nor NOR4 (N5442, N5427, N4327, N262, N2366);
xor XOR2 (N5443, N5436, N870);
nor NOR3 (N5444, N5440, N4152, N5052);
buf BUF1 (N5445, N5443);
or OR3 (N5446, N5423, N79, N5346);
xor XOR2 (N5447, N5439, N2886);
nor NOR4 (N5448, N5419, N1666, N3060, N5002);
nor NOR2 (N5449, N5442, N1639);
and AND3 (N5450, N5444, N3533, N175);
buf BUF1 (N5451, N5424);
nor NOR2 (N5452, N5437, N5228);
buf BUF1 (N5453, N5448);
and AND3 (N5454, N5447, N1327, N1621);
and AND4 (N5455, N5434, N2080, N2335, N2231);
nor NOR3 (N5456, N5451, N3377, N1962);
buf BUF1 (N5457, N5452);
nor NOR4 (N5458, N5445, N5415, N423, N4929);
or OR4 (N5459, N5456, N2285, N3540, N254);
nand NAND4 (N5460, N5453, N4884, N5283, N4256);
not NOT1 (N5461, N5446);
buf BUF1 (N5462, N5455);
nand NAND2 (N5463, N5458, N3458);
buf BUF1 (N5464, N5449);
xor XOR2 (N5465, N5450, N2651);
or OR4 (N5466, N5463, N820, N542, N4853);
and AND4 (N5467, N5454, N4524, N3930, N2529);
nor NOR4 (N5468, N5464, N5441, N5094, N2291);
xor XOR2 (N5469, N3202, N4847);
buf BUF1 (N5470, N5466);
or OR2 (N5471, N5469, N517);
buf BUF1 (N5472, N5468);
nand NAND4 (N5473, N5471, N4923, N4932, N4709);
and AND3 (N5474, N5460, N3992, N3845);
or OR3 (N5475, N5470, N673, N202);
not NOT1 (N5476, N5465);
xor XOR2 (N5477, N5459, N2089);
nand NAND2 (N5478, N5462, N420);
xor XOR2 (N5479, N5472, N2624);
xor XOR2 (N5480, N5461, N1121);
and AND2 (N5481, N5480, N2790);
and AND2 (N5482, N5473, N897);
xor XOR2 (N5483, N5482, N1108);
and AND4 (N5484, N5457, N2340, N1320, N1996);
or OR4 (N5485, N5474, N1075, N2734, N5250);
or OR3 (N5486, N5478, N1786, N1442);
and AND2 (N5487, N5486, N5208);
xor XOR2 (N5488, N5467, N1945);
buf BUF1 (N5489, N5488);
buf BUF1 (N5490, N5481);
not NOT1 (N5491, N5485);
or OR2 (N5492, N5476, N243);
and AND2 (N5493, N5483, N143);
nand NAND2 (N5494, N5477, N3603);
xor XOR2 (N5495, N5489, N3054);
or OR2 (N5496, N5494, N1068);
xor XOR2 (N5497, N5484, N5306);
not NOT1 (N5498, N5497);
not NOT1 (N5499, N5498);
and AND2 (N5500, N5479, N5155);
xor XOR2 (N5501, N5490, N975);
nand NAND3 (N5502, N5495, N3045, N1837);
xor XOR2 (N5503, N5475, N4559);
and AND3 (N5504, N5503, N1409, N2475);
not NOT1 (N5505, N5493);
nor NOR2 (N5506, N5502, N4682);
and AND2 (N5507, N5491, N2059);
or OR2 (N5508, N5507, N4933);
or OR2 (N5509, N5496, N1691);
not NOT1 (N5510, N5508);
nand NAND3 (N5511, N5500, N1568, N951);
and AND3 (N5512, N5492, N1904, N4484);
buf BUF1 (N5513, N5511);
nand NAND2 (N5514, N5501, N1975);
nand NAND2 (N5515, N5513, N3848);
not NOT1 (N5516, N5504);
or OR2 (N5517, N5487, N1248);
nor NOR4 (N5518, N5499, N2218, N2806, N4424);
xor XOR2 (N5519, N5516, N2913);
and AND3 (N5520, N5514, N1078, N1566);
xor XOR2 (N5521, N5506, N1764);
xor XOR2 (N5522, N5521, N2425);
or OR3 (N5523, N5505, N4079, N2062);
nor NOR3 (N5524, N5518, N5016, N3489);
nor NOR2 (N5525, N5523, N1517);
and AND3 (N5526, N5512, N1569, N3926);
nor NOR3 (N5527, N5522, N3389, N4407);
nand NAND4 (N5528, N5510, N5015, N5015, N1063);
nor NOR2 (N5529, N5515, N4627);
not NOT1 (N5530, N5509);
and AND2 (N5531, N5529, N312);
and AND4 (N5532, N5517, N1347, N5508, N2857);
nor NOR3 (N5533, N5524, N3982, N865);
not NOT1 (N5534, N5527);
not NOT1 (N5535, N5525);
nand NAND4 (N5536, N5534, N241, N2524, N1197);
not NOT1 (N5537, N5520);
not NOT1 (N5538, N5528);
or OR4 (N5539, N5537, N3519, N3637, N1672);
not NOT1 (N5540, N5539);
nor NOR2 (N5541, N5530, N5011);
xor XOR2 (N5542, N5541, N2003);
nor NOR3 (N5543, N5535, N3858, N2086);
nand NAND3 (N5544, N5526, N377, N3059);
xor XOR2 (N5545, N5532, N1555);
or OR2 (N5546, N5545, N82);
xor XOR2 (N5547, N5543, N1205);
buf BUF1 (N5548, N5536);
and AND2 (N5549, N5547, N2476);
or OR4 (N5550, N5546, N389, N1968, N1134);
and AND3 (N5551, N5548, N3507, N2755);
not NOT1 (N5552, N5531);
nor NOR4 (N5553, N5533, N3633, N2384, N5109);
buf BUF1 (N5554, N5550);
xor XOR2 (N5555, N5519, N263);
nor NOR4 (N5556, N5552, N4237, N4362, N5191);
nor NOR3 (N5557, N5555, N4078, N4498);
not NOT1 (N5558, N5551);
nor NOR4 (N5559, N5540, N800, N2427, N4128);
or OR4 (N5560, N5558, N1288, N5395, N3934);
buf BUF1 (N5561, N5553);
nand NAND2 (N5562, N5560, N5124);
not NOT1 (N5563, N5544);
nand NAND2 (N5564, N5542, N1162);
and AND3 (N5565, N5556, N194, N69);
nor NOR3 (N5566, N5557, N4074, N4516);
and AND3 (N5567, N5559, N3286, N699);
nand NAND3 (N5568, N5566, N3753, N5372);
or OR3 (N5569, N5538, N1923, N4387);
buf BUF1 (N5570, N5563);
buf BUF1 (N5571, N5567);
xor XOR2 (N5572, N5562, N5327);
not NOT1 (N5573, N5561);
and AND3 (N5574, N5571, N3621, N1509);
buf BUF1 (N5575, N5564);
and AND3 (N5576, N5569, N3828, N4034);
nor NOR3 (N5577, N5570, N3673, N835);
nor NOR2 (N5578, N5572, N2453);
buf BUF1 (N5579, N5578);
nand NAND3 (N5580, N5576, N1440, N5061);
not NOT1 (N5581, N5574);
nor NOR2 (N5582, N5581, N2197);
not NOT1 (N5583, N5580);
buf BUF1 (N5584, N5565);
or OR3 (N5585, N5554, N233, N411);
nor NOR2 (N5586, N5585, N2264);
nor NOR4 (N5587, N5577, N2248, N711, N2657);
nor NOR4 (N5588, N5579, N3782, N2991, N948);
and AND4 (N5589, N5586, N3711, N3125, N3996);
buf BUF1 (N5590, N5583);
not NOT1 (N5591, N5589);
nor NOR2 (N5592, N5575, N1409);
not NOT1 (N5593, N5590);
and AND3 (N5594, N5592, N4678, N2185);
nor NOR4 (N5595, N5594, N3988, N3274, N4164);
buf BUF1 (N5596, N5582);
xor XOR2 (N5597, N5595, N3476);
or OR2 (N5598, N5549, N4810);
not NOT1 (N5599, N5588);
or OR4 (N5600, N5596, N2536, N2754, N3946);
buf BUF1 (N5601, N5593);
nor NOR3 (N5602, N5573, N223, N2313);
xor XOR2 (N5603, N5584, N2658);
not NOT1 (N5604, N5600);
buf BUF1 (N5605, N5604);
buf BUF1 (N5606, N5603);
nor NOR2 (N5607, N5606, N3453);
buf BUF1 (N5608, N5598);
nand NAND4 (N5609, N5568, N2598, N3043, N743);
xor XOR2 (N5610, N5607, N4);
and AND4 (N5611, N5605, N3458, N3050, N1590);
not NOT1 (N5612, N5587);
nor NOR3 (N5613, N5597, N5177, N3564);
nand NAND3 (N5614, N5602, N4349, N2263);
nor NOR3 (N5615, N5611, N5541, N1091);
not NOT1 (N5616, N5608);
and AND4 (N5617, N5610, N380, N4257, N1139);
nor NOR2 (N5618, N5591, N1718);
nand NAND2 (N5619, N5615, N5211);
nor NOR2 (N5620, N5609, N411);
buf BUF1 (N5621, N5613);
nand NAND2 (N5622, N5618, N4825);
nor NOR2 (N5623, N5616, N4222);
not NOT1 (N5624, N5612);
or OR3 (N5625, N5620, N2758, N1378);
nand NAND3 (N5626, N5624, N1057, N527);
buf BUF1 (N5627, N5626);
buf BUF1 (N5628, N5614);
xor XOR2 (N5629, N5617, N542);
nand NAND3 (N5630, N5619, N3404, N3595);
nor NOR3 (N5631, N5629, N2423, N3185);
nor NOR4 (N5632, N5631, N4943, N4591, N832);
or OR4 (N5633, N5622, N1203, N3014, N164);
buf BUF1 (N5634, N5632);
buf BUF1 (N5635, N5599);
and AND4 (N5636, N5630, N3519, N4747, N16);
xor XOR2 (N5637, N5633, N2669);
nand NAND4 (N5638, N5634, N2231, N1604, N879);
or OR2 (N5639, N5601, N5083);
nand NAND4 (N5640, N5627, N3316, N2545, N3750);
nand NAND2 (N5641, N5625, N5143);
xor XOR2 (N5642, N5636, N3466);
nand NAND4 (N5643, N5639, N1425, N4597, N4026);
or OR4 (N5644, N5621, N3543, N5063, N1605);
or OR3 (N5645, N5641, N5444, N3704);
nand NAND3 (N5646, N5638, N754, N4179);
and AND2 (N5647, N5640, N2189);
nand NAND3 (N5648, N5647, N4967, N2659);
and AND2 (N5649, N5643, N2167);
and AND4 (N5650, N5645, N2505, N2694, N2776);
nor NOR4 (N5651, N5649, N4668, N2279, N1511);
buf BUF1 (N5652, N5644);
nor NOR2 (N5653, N5650, N1791);
xor XOR2 (N5654, N5646, N4988);
or OR2 (N5655, N5653, N3454);
not NOT1 (N5656, N5623);
not NOT1 (N5657, N5654);
or OR3 (N5658, N5637, N5283, N1195);
not NOT1 (N5659, N5648);
xor XOR2 (N5660, N5659, N5461);
nor NOR2 (N5661, N5660, N1716);
xor XOR2 (N5662, N5642, N1196);
or OR4 (N5663, N5662, N4444, N4370, N1591);
or OR3 (N5664, N5651, N3793, N1269);
not NOT1 (N5665, N5663);
or OR4 (N5666, N5656, N211, N4805, N2133);
and AND3 (N5667, N5655, N5178, N5003);
nand NAND4 (N5668, N5665, N4127, N4096, N1720);
nand NAND4 (N5669, N5657, N2087, N2415, N6);
nand NAND2 (N5670, N5669, N3416);
and AND2 (N5671, N5628, N963);
and AND3 (N5672, N5671, N4203, N3145);
and AND4 (N5673, N5635, N4211, N4563, N2068);
and AND3 (N5674, N5672, N2708, N981);
or OR4 (N5675, N5674, N121, N4130, N2647);
or OR3 (N5676, N5673, N3692, N2299);
not NOT1 (N5677, N5664);
xor XOR2 (N5678, N5670, N1038);
nor NOR3 (N5679, N5658, N703, N4100);
or OR3 (N5680, N5652, N3067, N2219);
nor NOR2 (N5681, N5680, N1213);
buf BUF1 (N5682, N5679);
nand NAND4 (N5683, N5668, N2357, N4801, N1622);
xor XOR2 (N5684, N5682, N894);
buf BUF1 (N5685, N5676);
xor XOR2 (N5686, N5684, N176);
nand NAND2 (N5687, N5685, N5312);
xor XOR2 (N5688, N5681, N4948);
or OR4 (N5689, N5678, N2384, N5669, N2100);
or OR2 (N5690, N5687, N2210);
nand NAND3 (N5691, N5690, N3914, N3119);
buf BUF1 (N5692, N5686);
not NOT1 (N5693, N5689);
or OR2 (N5694, N5688, N2601);
nor NOR4 (N5695, N5675, N738, N451, N840);
not NOT1 (N5696, N5683);
or OR2 (N5697, N5694, N452);
and AND3 (N5698, N5696, N5041, N636);
not NOT1 (N5699, N5695);
and AND4 (N5700, N5677, N1683, N3921, N1312);
nand NAND3 (N5701, N5700, N5076, N3842);
or OR4 (N5702, N5666, N725, N1049, N3824);
or OR2 (N5703, N5698, N2047);
not NOT1 (N5704, N5667);
or OR2 (N5705, N5703, N3405);
nand NAND4 (N5706, N5704, N5557, N1686, N5117);
not NOT1 (N5707, N5702);
or OR3 (N5708, N5691, N2341, N3070);
xor XOR2 (N5709, N5708, N3414);
or OR3 (N5710, N5693, N5176, N2208);
nand NAND3 (N5711, N5661, N2320, N1788);
and AND3 (N5712, N5711, N2118, N199);
xor XOR2 (N5713, N5699, N3103);
nor NOR3 (N5714, N5707, N731, N800);
not NOT1 (N5715, N5706);
xor XOR2 (N5716, N5709, N2528);
and AND2 (N5717, N5701, N4540);
or OR3 (N5718, N5705, N251, N1226);
nor NOR2 (N5719, N5712, N3785);
or OR4 (N5720, N5715, N1063, N3139, N2460);
xor XOR2 (N5721, N5717, N2896);
or OR4 (N5722, N5720, N286, N4953, N4770);
not NOT1 (N5723, N5721);
xor XOR2 (N5724, N5722, N3057);
nor NOR4 (N5725, N5724, N3573, N3333, N4105);
nand NAND4 (N5726, N5713, N3502, N3151, N5114);
not NOT1 (N5727, N5719);
nand NAND2 (N5728, N5718, N2437);
buf BUF1 (N5729, N5723);
nor NOR3 (N5730, N5728, N4977, N2108);
buf BUF1 (N5731, N5716);
xor XOR2 (N5732, N5726, N3098);
not NOT1 (N5733, N5730);
not NOT1 (N5734, N5732);
and AND3 (N5735, N5725, N1496, N426);
nand NAND2 (N5736, N5733, N4754);
nand NAND2 (N5737, N5736, N4451);
xor XOR2 (N5738, N5692, N5580);
buf BUF1 (N5739, N5734);
nor NOR4 (N5740, N5727, N121, N5634, N5522);
nor NOR4 (N5741, N5737, N5198, N2053, N4248);
nand NAND2 (N5742, N5731, N1741);
or OR3 (N5743, N5729, N4835, N4029);
xor XOR2 (N5744, N5740, N2634);
buf BUF1 (N5745, N5714);
and AND4 (N5746, N5710, N2832, N1466, N2438);
buf BUF1 (N5747, N5746);
buf BUF1 (N5748, N5745);
not NOT1 (N5749, N5697);
and AND2 (N5750, N5735, N3562);
not NOT1 (N5751, N5739);
or OR2 (N5752, N5750, N2810);
not NOT1 (N5753, N5752);
or OR2 (N5754, N5741, N369);
nand NAND3 (N5755, N5743, N1014, N3595);
and AND4 (N5756, N5751, N646, N2455, N347);
or OR3 (N5757, N5742, N4010, N395);
nand NAND2 (N5758, N5738, N2292);
or OR4 (N5759, N5754, N3541, N2463, N2330);
nand NAND3 (N5760, N5748, N3926, N5715);
or OR3 (N5761, N5758, N5665, N3696);
buf BUF1 (N5762, N5753);
xor XOR2 (N5763, N5757, N4244);
not NOT1 (N5764, N5762);
buf BUF1 (N5765, N5747);
nand NAND2 (N5766, N5763, N4931);
buf BUF1 (N5767, N5764);
or OR3 (N5768, N5767, N1654, N5613);
not NOT1 (N5769, N5749);
xor XOR2 (N5770, N5761, N1298);
buf BUF1 (N5771, N5770);
nand NAND3 (N5772, N5766, N5688, N4837);
nand NAND3 (N5773, N5759, N2212, N855);
xor XOR2 (N5774, N5765, N2060);
nand NAND4 (N5775, N5744, N5710, N1588, N4430);
nand NAND2 (N5776, N5771, N3985);
not NOT1 (N5777, N5768);
buf BUF1 (N5778, N5773);
not NOT1 (N5779, N5777);
not NOT1 (N5780, N5774);
buf BUF1 (N5781, N5755);
buf BUF1 (N5782, N5775);
and AND2 (N5783, N5782, N152);
xor XOR2 (N5784, N5780, N5775);
nand NAND4 (N5785, N5776, N1173, N5406, N4026);
buf BUF1 (N5786, N5784);
and AND2 (N5787, N5760, N1080);
and AND4 (N5788, N5779, N1368, N5288, N5426);
nand NAND3 (N5789, N5785, N109, N1747);
buf BUF1 (N5790, N5781);
xor XOR2 (N5791, N5756, N3963);
or OR4 (N5792, N5783, N3827, N1788, N2492);
nand NAND4 (N5793, N5778, N2963, N133, N181);
not NOT1 (N5794, N5787);
or OR4 (N5795, N5789, N804, N5722, N2915);
and AND4 (N5796, N5794, N1407, N5027, N4696);
nor NOR4 (N5797, N5790, N2411, N1407, N4007);
not NOT1 (N5798, N5786);
nand NAND4 (N5799, N5769, N3624, N5745, N2762);
nor NOR2 (N5800, N5797, N410);
not NOT1 (N5801, N5798);
nor NOR3 (N5802, N5793, N1378, N2258);
xor XOR2 (N5803, N5795, N1267);
and AND3 (N5804, N5800, N933, N1964);
and AND2 (N5805, N5801, N3510);
nand NAND3 (N5806, N5805, N3508, N3695);
nand NAND3 (N5807, N5802, N552, N463);
buf BUF1 (N5808, N5791);
or OR4 (N5809, N5808, N4249, N1399, N953);
nand NAND4 (N5810, N5788, N2745, N5714, N4065);
or OR2 (N5811, N5809, N4464);
nor NOR3 (N5812, N5772, N3640, N4458);
and AND3 (N5813, N5796, N5016, N4287);
xor XOR2 (N5814, N5807, N869);
nor NOR3 (N5815, N5814, N5606, N330);
nor NOR2 (N5816, N5815, N3783);
nand NAND2 (N5817, N5811, N2055);
nor NOR4 (N5818, N5799, N4524, N497, N1836);
xor XOR2 (N5819, N5792, N5687);
and AND4 (N5820, N5818, N1273, N290, N4274);
buf BUF1 (N5821, N5803);
not NOT1 (N5822, N5813);
not NOT1 (N5823, N5819);
nand NAND3 (N5824, N5812, N4345, N5512);
nor NOR3 (N5825, N5806, N4356, N1753);
xor XOR2 (N5826, N5817, N4793);
nand NAND4 (N5827, N5816, N1674, N3032, N4276);
xor XOR2 (N5828, N5827, N3006);
not NOT1 (N5829, N5823);
nor NOR4 (N5830, N5829, N2597, N4888, N4309);
or OR4 (N5831, N5804, N3034, N2407, N1955);
nand NAND3 (N5832, N5810, N3065, N702);
not NOT1 (N5833, N5825);
and AND4 (N5834, N5824, N2592, N4103, N1863);
nand NAND4 (N5835, N5830, N3667, N4638, N1523);
or OR2 (N5836, N5831, N5701);
buf BUF1 (N5837, N5832);
or OR3 (N5838, N5822, N4245, N1272);
and AND4 (N5839, N5834, N5736, N3089, N1327);
buf BUF1 (N5840, N5837);
not NOT1 (N5841, N5838);
and AND4 (N5842, N5835, N5417, N5708, N4875);
or OR4 (N5843, N5840, N1014, N1585, N4128);
nand NAND4 (N5844, N5839, N3489, N1462, N2295);
not NOT1 (N5845, N5842);
not NOT1 (N5846, N5843);
and AND4 (N5847, N5845, N5604, N5065, N4801);
or OR4 (N5848, N5836, N664, N806, N5578);
xor XOR2 (N5849, N5841, N1815);
nand NAND2 (N5850, N5849, N4268);
nor NOR3 (N5851, N5848, N2126, N5301);
and AND3 (N5852, N5833, N340, N2295);
or OR3 (N5853, N5821, N3504, N2057);
or OR3 (N5854, N5826, N2872, N5815);
nor NOR4 (N5855, N5828, N869, N4168, N2857);
nand NAND2 (N5856, N5850, N3431);
buf BUF1 (N5857, N5847);
or OR2 (N5858, N5846, N584);
nor NOR2 (N5859, N5851, N3891);
not NOT1 (N5860, N5857);
xor XOR2 (N5861, N5852, N4334);
nor NOR4 (N5862, N5844, N2336, N3345, N4808);
and AND4 (N5863, N5855, N4872, N3517, N3507);
and AND3 (N5864, N5860, N1342, N1997);
buf BUF1 (N5865, N5853);
nand NAND3 (N5866, N5865, N1651, N5830);
not NOT1 (N5867, N5866);
and AND4 (N5868, N5858, N1713, N527, N1053);
not NOT1 (N5869, N5867);
not NOT1 (N5870, N5864);
not NOT1 (N5871, N5870);
not NOT1 (N5872, N5863);
not NOT1 (N5873, N5871);
xor XOR2 (N5874, N5820, N3116);
and AND2 (N5875, N5861, N5760);
or OR3 (N5876, N5875, N5323, N5324);
or OR2 (N5877, N5859, N5602);
nand NAND2 (N5878, N5872, N4487);
buf BUF1 (N5879, N5878);
xor XOR2 (N5880, N5873, N1656);
or OR4 (N5881, N5862, N1572, N4508, N2877);
not NOT1 (N5882, N5879);
or OR4 (N5883, N5880, N738, N5693, N5874);
not NOT1 (N5884, N2802);
and AND3 (N5885, N5856, N4934, N2018);
not NOT1 (N5886, N5881);
buf BUF1 (N5887, N5884);
not NOT1 (N5888, N5854);
not NOT1 (N5889, N5868);
nand NAND3 (N5890, N5883, N5747, N3190);
buf BUF1 (N5891, N5890);
or OR2 (N5892, N5876, N5389);
nand NAND2 (N5893, N5887, N5315);
or OR4 (N5894, N5893, N4415, N2910, N2685);
and AND3 (N5895, N5886, N603, N820);
not NOT1 (N5896, N5869);
nor NOR4 (N5897, N5882, N1726, N1900, N1950);
not NOT1 (N5898, N5897);
nor NOR3 (N5899, N5889, N4540, N2991);
nor NOR3 (N5900, N5888, N3569, N3332);
buf BUF1 (N5901, N5896);
not NOT1 (N5902, N5892);
and AND2 (N5903, N5895, N3277);
xor XOR2 (N5904, N5894, N5762);
or OR4 (N5905, N5903, N676, N5431, N214);
and AND2 (N5906, N5904, N3086);
xor XOR2 (N5907, N5898, N256);
buf BUF1 (N5908, N5905);
xor XOR2 (N5909, N5908, N3984);
not NOT1 (N5910, N5885);
xor XOR2 (N5911, N5909, N4174);
nor NOR3 (N5912, N5902, N3575, N5883);
xor XOR2 (N5913, N5910, N806);
or OR3 (N5914, N5877, N1505, N4065);
buf BUF1 (N5915, N5911);
not NOT1 (N5916, N5906);
nand NAND3 (N5917, N5915, N4651, N5624);
xor XOR2 (N5918, N5899, N1577);
buf BUF1 (N5919, N5918);
or OR3 (N5920, N5917, N2602, N1428);
not NOT1 (N5921, N5914);
and AND2 (N5922, N5913, N2888);
nand NAND2 (N5923, N5916, N2932);
nor NOR2 (N5924, N5907, N5515);
and AND2 (N5925, N5901, N3052);
nand NAND3 (N5926, N5920, N5283, N1829);
or OR2 (N5927, N5891, N1939);
nor NOR2 (N5928, N5927, N2432);
nor NOR3 (N5929, N5923, N5059, N2308);
not NOT1 (N5930, N5922);
buf BUF1 (N5931, N5928);
and AND3 (N5932, N5926, N5108, N131);
not NOT1 (N5933, N5900);
nand NAND2 (N5934, N5912, N5336);
xor XOR2 (N5935, N5930, N5577);
nor NOR2 (N5936, N5932, N5258);
nor NOR4 (N5937, N5935, N4329, N1773, N2498);
buf BUF1 (N5938, N5921);
or OR3 (N5939, N5933, N2481, N5098);
xor XOR2 (N5940, N5937, N4351);
or OR4 (N5941, N5919, N1208, N2915, N1407);
buf BUF1 (N5942, N5939);
nor NOR2 (N5943, N5929, N3346);
and AND3 (N5944, N5936, N5098, N332);
and AND3 (N5945, N5942, N2722, N4606);
nor NOR4 (N5946, N5924, N98, N777, N1377);
and AND2 (N5947, N5943, N2697);
or OR2 (N5948, N5945, N2819);
and AND3 (N5949, N5948, N253, N2850);
nor NOR4 (N5950, N5938, N3534, N1354, N1849);
or OR2 (N5951, N5931, N198);
nand NAND4 (N5952, N5946, N1723, N3528, N4756);
and AND3 (N5953, N5925, N5777, N2511);
or OR4 (N5954, N5934, N5161, N4985, N1333);
and AND3 (N5955, N5950, N5669, N2978);
xor XOR2 (N5956, N5954, N3436);
buf BUF1 (N5957, N5947);
buf BUF1 (N5958, N5951);
buf BUF1 (N5959, N5955);
buf BUF1 (N5960, N5956);
xor XOR2 (N5961, N5958, N3076);
buf BUF1 (N5962, N5953);
xor XOR2 (N5963, N5952, N1467);
not NOT1 (N5964, N5959);
or OR3 (N5965, N5960, N2708, N2231);
not NOT1 (N5966, N5941);
buf BUF1 (N5967, N5962);
buf BUF1 (N5968, N5967);
or OR3 (N5969, N5944, N440, N2374);
and AND3 (N5970, N5957, N3951, N2197);
and AND4 (N5971, N5965, N3477, N4406, N1500);
and AND4 (N5972, N5970, N4432, N1194, N3007);
nor NOR3 (N5973, N5972, N4910, N4179);
or OR3 (N5974, N5971, N5286, N5318);
and AND4 (N5975, N5966, N126, N769, N3616);
or OR2 (N5976, N5940, N2662);
or OR3 (N5977, N5974, N1109, N4131);
not NOT1 (N5978, N5961);
nand NAND3 (N5979, N5976, N1469, N4300);
nor NOR4 (N5980, N5968, N3017, N1964, N3472);
nor NOR4 (N5981, N5978, N3196, N3432, N2496);
buf BUF1 (N5982, N5975);
buf BUF1 (N5983, N5977);
or OR4 (N5984, N5979, N3163, N3896, N2231);
nor NOR4 (N5985, N5969, N4563, N4154, N677);
or OR2 (N5986, N5984, N1772);
buf BUF1 (N5987, N5963);
not NOT1 (N5988, N5949);
nor NOR4 (N5989, N5986, N1314, N244, N4549);
xor XOR2 (N5990, N5985, N1283);
nor NOR4 (N5991, N5981, N5744, N43, N5782);
buf BUF1 (N5992, N5987);
not NOT1 (N5993, N5990);
buf BUF1 (N5994, N5988);
nand NAND4 (N5995, N5989, N3502, N122, N5781);
or OR2 (N5996, N5991, N3082);
nor NOR4 (N5997, N5993, N3177, N5741, N3306);
nor NOR4 (N5998, N5983, N3904, N4429, N5123);
or OR3 (N5999, N5998, N3565, N4928);
and AND2 (N6000, N5999, N4016);
nor NOR3 (N6001, N5992, N260, N4591);
xor XOR2 (N6002, N5964, N3817);
and AND3 (N6003, N6001, N5181, N565);
not NOT1 (N6004, N6002);
and AND2 (N6005, N5995, N3947);
buf BUF1 (N6006, N5973);
nor NOR3 (N6007, N6005, N2470, N972);
nand NAND2 (N6008, N5982, N4767);
or OR3 (N6009, N5996, N5891, N4837);
buf BUF1 (N6010, N6008);
and AND2 (N6011, N6000, N1090);
and AND4 (N6012, N6007, N3423, N3190, N181);
xor XOR2 (N6013, N5994, N2210);
xor XOR2 (N6014, N6006, N3459);
or OR3 (N6015, N6010, N4183, N4555);
or OR4 (N6016, N6012, N3722, N5382, N5253);
nand NAND2 (N6017, N6013, N4956);
and AND2 (N6018, N5980, N3767);
buf BUF1 (N6019, N6017);
or OR2 (N6020, N6019, N67);
buf BUF1 (N6021, N6020);
xor XOR2 (N6022, N6004, N5726);
nor NOR4 (N6023, N6016, N4918, N4821, N361);
not NOT1 (N6024, N6009);
xor XOR2 (N6025, N6023, N5645);
nor NOR2 (N6026, N6011, N2626);
nand NAND2 (N6027, N6025, N5797);
or OR3 (N6028, N6027, N1454, N3464);
and AND3 (N6029, N6021, N2603, N688);
and AND3 (N6030, N5997, N2793, N3120);
xor XOR2 (N6031, N6029, N3938);
and AND3 (N6032, N6014, N3582, N5641);
nor NOR2 (N6033, N6003, N2950);
xor XOR2 (N6034, N6033, N2673);
and AND2 (N6035, N6030, N2425);
nand NAND2 (N6036, N6032, N5990);
and AND4 (N6037, N6035, N1058, N3051, N5134);
buf BUF1 (N6038, N6028);
nand NAND4 (N6039, N6037, N4153, N5269, N3248);
not NOT1 (N6040, N6024);
nor NOR4 (N6041, N6031, N3158, N701, N5972);
xor XOR2 (N6042, N6022, N637);
nand NAND3 (N6043, N6015, N870, N2538);
and AND4 (N6044, N6042, N2486, N1484, N4553);
nand NAND2 (N6045, N6040, N2229);
nand NAND2 (N6046, N6044, N1134);
buf BUF1 (N6047, N6018);
not NOT1 (N6048, N6046);
nand NAND4 (N6049, N6034, N5100, N2419, N401);
xor XOR2 (N6050, N6049, N352);
xor XOR2 (N6051, N6047, N1070);
xor XOR2 (N6052, N6051, N4237);
and AND4 (N6053, N6043, N2659, N660, N1142);
or OR3 (N6054, N6039, N5181, N915);
or OR2 (N6055, N6045, N3638);
nand NAND4 (N6056, N6026, N3643, N5869, N1826);
buf BUF1 (N6057, N6041);
nand NAND3 (N6058, N6056, N4905, N3640);
not NOT1 (N6059, N6038);
and AND4 (N6060, N6052, N2696, N1990, N4356);
not NOT1 (N6061, N6055);
and AND2 (N6062, N6061, N3408);
buf BUF1 (N6063, N6054);
or OR4 (N6064, N6057, N4284, N3267, N2170);
xor XOR2 (N6065, N6048, N4925);
or OR2 (N6066, N6050, N5739);
or OR4 (N6067, N6058, N1158, N1277, N6012);
buf BUF1 (N6068, N6065);
xor XOR2 (N6069, N6059, N546);
and AND4 (N6070, N6067, N2059, N2564, N3151);
and AND2 (N6071, N6036, N2386);
xor XOR2 (N6072, N6060, N5640);
or OR4 (N6073, N6066, N1375, N2389, N1632);
not NOT1 (N6074, N6053);
and AND3 (N6075, N6072, N3029, N3359);
nand NAND2 (N6076, N6069, N3020);
and AND2 (N6077, N6068, N82);
nor NOR3 (N6078, N6071, N3482, N360);
nand NAND4 (N6079, N6074, N1632, N5864, N2820);
nor NOR3 (N6080, N6070, N3176, N2856);
nand NAND3 (N6081, N6078, N3208, N3765);
xor XOR2 (N6082, N6063, N455);
buf BUF1 (N6083, N6064);
xor XOR2 (N6084, N6080, N2268);
not NOT1 (N6085, N6082);
not NOT1 (N6086, N6084);
buf BUF1 (N6087, N6062);
xor XOR2 (N6088, N6075, N3317);
buf BUF1 (N6089, N6079);
nor NOR2 (N6090, N6086, N3005);
not NOT1 (N6091, N6087);
nor NOR3 (N6092, N6090, N1232, N2051);
and AND2 (N6093, N6089, N5143);
nor NOR2 (N6094, N6081, N2761);
buf BUF1 (N6095, N6088);
nor NOR2 (N6096, N6073, N5184);
and AND4 (N6097, N6096, N2416, N845, N4769);
not NOT1 (N6098, N6097);
not NOT1 (N6099, N6076);
xor XOR2 (N6100, N6083, N4779);
xor XOR2 (N6101, N6091, N1421);
xor XOR2 (N6102, N6085, N1867);
buf BUF1 (N6103, N6099);
nor NOR4 (N6104, N6094, N196, N1392, N1681);
and AND2 (N6105, N6103, N1924);
nor NOR3 (N6106, N6077, N2544, N1630);
nand NAND3 (N6107, N6092, N5659, N612);
buf BUF1 (N6108, N6101);
not NOT1 (N6109, N6093);
xor XOR2 (N6110, N6100, N216);
or OR3 (N6111, N6108, N1557, N3552);
not NOT1 (N6112, N6098);
nor NOR3 (N6113, N6105, N2527, N3523);
nor NOR2 (N6114, N6095, N1323);
nand NAND3 (N6115, N6107, N4672, N3157);
xor XOR2 (N6116, N6109, N5148);
nor NOR2 (N6117, N6115, N1935);
nor NOR2 (N6118, N6110, N5951);
nand NAND2 (N6119, N6102, N1350);
nor NOR3 (N6120, N6114, N4121, N4037);
not NOT1 (N6121, N6106);
xor XOR2 (N6122, N6111, N1468);
xor XOR2 (N6123, N6116, N5220);
nand NAND4 (N6124, N6117, N2959, N2840, N5110);
xor XOR2 (N6125, N6123, N1543);
nor NOR2 (N6126, N6120, N5565);
not NOT1 (N6127, N6119);
and AND3 (N6128, N6121, N2496, N2927);
not NOT1 (N6129, N6112);
xor XOR2 (N6130, N6129, N2805);
nand NAND4 (N6131, N6130, N1220, N5530, N5717);
nand NAND4 (N6132, N6126, N661, N3607, N4612);
nor NOR4 (N6133, N6132, N4982, N5705, N710);
nand NAND4 (N6134, N6113, N5093, N1909, N3998);
nor NOR2 (N6135, N6128, N4497);
or OR4 (N6136, N6118, N3346, N4441, N1758);
and AND3 (N6137, N6133, N4784, N4649);
buf BUF1 (N6138, N6104);
nand NAND4 (N6139, N6135, N4770, N5135, N2663);
not NOT1 (N6140, N6137);
nand NAND4 (N6141, N6122, N4716, N273, N3636);
not NOT1 (N6142, N6125);
xor XOR2 (N6143, N6141, N5354);
buf BUF1 (N6144, N6139);
xor XOR2 (N6145, N6143, N4294);
buf BUF1 (N6146, N6144);
and AND2 (N6147, N6131, N5154);
buf BUF1 (N6148, N6142);
buf BUF1 (N6149, N6134);
nor NOR2 (N6150, N6138, N3636);
buf BUF1 (N6151, N6149);
xor XOR2 (N6152, N6140, N1285);
or OR4 (N6153, N6127, N1462, N1072, N2167);
not NOT1 (N6154, N6145);
or OR2 (N6155, N6152, N710);
nor NOR4 (N6156, N6154, N4377, N4117, N4477);
and AND2 (N6157, N6124, N5465);
and AND2 (N6158, N6150, N6047);
buf BUF1 (N6159, N6157);
and AND2 (N6160, N6159, N672);
xor XOR2 (N6161, N6153, N779);
and AND3 (N6162, N6156, N5637, N3734);
buf BUF1 (N6163, N6158);
not NOT1 (N6164, N6148);
nor NOR2 (N6165, N6155, N3996);
or OR3 (N6166, N6165, N1450, N2876);
nand NAND2 (N6167, N6166, N2399);
nand NAND3 (N6168, N6163, N3707, N3204);
not NOT1 (N6169, N6161);
not NOT1 (N6170, N6162);
not NOT1 (N6171, N6151);
and AND4 (N6172, N6167, N2126, N3347, N6013);
not NOT1 (N6173, N6168);
and AND3 (N6174, N6160, N1186, N5358);
and AND4 (N6175, N6169, N2800, N969, N1588);
nand NAND2 (N6176, N6147, N3834);
nor NOR3 (N6177, N6170, N624, N4322);
nor NOR2 (N6178, N6172, N5067);
xor XOR2 (N6179, N6171, N1490);
nand NAND3 (N6180, N6173, N4454, N5665);
xor XOR2 (N6181, N6175, N5526);
and AND2 (N6182, N6136, N4999);
or OR3 (N6183, N6179, N63, N4987);
or OR2 (N6184, N6178, N2141);
xor XOR2 (N6185, N6174, N1224);
and AND4 (N6186, N6183, N4393, N5742, N3597);
and AND2 (N6187, N6181, N3633);
or OR4 (N6188, N6184, N5602, N2250, N5394);
or OR3 (N6189, N6180, N1742, N6114);
and AND4 (N6190, N6188, N6184, N1628, N2746);
nand NAND2 (N6191, N6185, N1429);
not NOT1 (N6192, N6176);
not NOT1 (N6193, N6187);
xor XOR2 (N6194, N6190, N201);
buf BUF1 (N6195, N6191);
nor NOR2 (N6196, N6192, N1768);
nand NAND2 (N6197, N6186, N1434);
or OR4 (N6198, N6182, N5165, N3816, N3889);
nand NAND3 (N6199, N6164, N4126, N637);
nor NOR3 (N6200, N6194, N5373, N2901);
not NOT1 (N6201, N6193);
xor XOR2 (N6202, N6146, N1733);
nand NAND3 (N6203, N6198, N5957, N359);
or OR3 (N6204, N6203, N6045, N3787);
or OR3 (N6205, N6197, N1870, N5794);
xor XOR2 (N6206, N6177, N18);
nor NOR3 (N6207, N6196, N3816, N3583);
not NOT1 (N6208, N6202);
or OR3 (N6209, N6199, N4251, N3494);
nor NOR4 (N6210, N6195, N4591, N2024, N4902);
or OR4 (N6211, N6201, N2660, N3250, N5853);
or OR4 (N6212, N6200, N5436, N1691, N1593);
buf BUF1 (N6213, N6207);
not NOT1 (N6214, N6204);
or OR3 (N6215, N6213, N2472, N2794);
nand NAND4 (N6216, N6211, N5227, N581, N724);
nand NAND2 (N6217, N6212, N4197);
or OR4 (N6218, N6215, N380, N130, N962);
or OR3 (N6219, N6214, N1030, N3011);
nor NOR2 (N6220, N6219, N5602);
buf BUF1 (N6221, N6206);
and AND2 (N6222, N6216, N3965);
xor XOR2 (N6223, N6218, N50);
nand NAND4 (N6224, N6208, N327, N3537, N5757);
nor NOR3 (N6225, N6221, N6137, N2184);
buf BUF1 (N6226, N6189);
nor NOR3 (N6227, N6205, N1037, N3176);
nand NAND4 (N6228, N6222, N2541, N813, N2235);
nand NAND3 (N6229, N6210, N554, N3032);
not NOT1 (N6230, N6209);
nand NAND4 (N6231, N6225, N4372, N245, N6122);
buf BUF1 (N6232, N6227);
buf BUF1 (N6233, N6232);
buf BUF1 (N6234, N6220);
or OR4 (N6235, N6226, N3627, N6166, N4555);
nand NAND3 (N6236, N6234, N3179, N3840);
not NOT1 (N6237, N6217);
or OR2 (N6238, N6230, N2833);
not NOT1 (N6239, N6237);
xor XOR2 (N6240, N6239, N2150);
buf BUF1 (N6241, N6233);
xor XOR2 (N6242, N6241, N982);
or OR4 (N6243, N6238, N3869, N3491, N3668);
buf BUF1 (N6244, N6235);
xor XOR2 (N6245, N6229, N5922);
not NOT1 (N6246, N6240);
and AND4 (N6247, N6223, N183, N4102, N3237);
and AND2 (N6248, N6243, N5568);
not NOT1 (N6249, N6224);
and AND2 (N6250, N6228, N703);
and AND4 (N6251, N6246, N5667, N3234, N3219);
and AND2 (N6252, N6231, N4687);
nand NAND4 (N6253, N6248, N3329, N1268, N4454);
nand NAND4 (N6254, N6247, N3092, N43, N53);
not NOT1 (N6255, N6236);
nor NOR4 (N6256, N6252, N1122, N5914, N5118);
nor NOR3 (N6257, N6245, N2262, N5177);
or OR2 (N6258, N6242, N5785);
nor NOR2 (N6259, N6251, N790);
buf BUF1 (N6260, N6244);
and AND4 (N6261, N6249, N4856, N2863, N1575);
and AND3 (N6262, N6255, N1745, N3037);
buf BUF1 (N6263, N6253);
or OR3 (N6264, N6259, N4702, N5055);
not NOT1 (N6265, N6250);
or OR2 (N6266, N6258, N5209);
not NOT1 (N6267, N6264);
or OR2 (N6268, N6257, N5621);
and AND4 (N6269, N6261, N4726, N3332, N4823);
not NOT1 (N6270, N6256);
nor NOR4 (N6271, N6268, N3722, N3697, N4953);
not NOT1 (N6272, N6260);
xor XOR2 (N6273, N6272, N602);
or OR4 (N6274, N6273, N3806, N3851, N2296);
nor NOR4 (N6275, N6274, N3943, N1493, N363);
buf BUF1 (N6276, N6262);
buf BUF1 (N6277, N6267);
or OR2 (N6278, N6254, N3855);
buf BUF1 (N6279, N6269);
and AND2 (N6280, N6279, N1998);
xor XOR2 (N6281, N6278, N4556);
buf BUF1 (N6282, N6280);
buf BUF1 (N6283, N6281);
xor XOR2 (N6284, N6277, N1694);
nor NOR4 (N6285, N6270, N3915, N5547, N5715);
nand NAND3 (N6286, N6275, N6010, N2316);
and AND3 (N6287, N6266, N3146, N5593);
and AND4 (N6288, N6276, N4507, N5128, N3102);
and AND2 (N6289, N6286, N4332);
and AND4 (N6290, N6283, N1664, N2987, N633);
xor XOR2 (N6291, N6263, N5453);
and AND3 (N6292, N6288, N2762, N854);
xor XOR2 (N6293, N6282, N4781);
or OR2 (N6294, N6292, N3075);
and AND4 (N6295, N6284, N2634, N3594, N6166);
xor XOR2 (N6296, N6265, N3699);
xor XOR2 (N6297, N6296, N5019);
xor XOR2 (N6298, N6285, N4857);
xor XOR2 (N6299, N6294, N1816);
or OR4 (N6300, N6290, N1865, N2790, N2300);
buf BUF1 (N6301, N6299);
nor NOR4 (N6302, N6289, N5517, N4388, N241);
nor NOR2 (N6303, N6300, N3228);
xor XOR2 (N6304, N6298, N5221);
nor NOR4 (N6305, N6287, N5984, N4403, N5024);
or OR2 (N6306, N6303, N3544);
buf BUF1 (N6307, N6293);
nor NOR2 (N6308, N6306, N619);
and AND2 (N6309, N6304, N4149);
nor NOR3 (N6310, N6305, N4703, N964);
nand NAND4 (N6311, N6308, N5102, N563, N350);
buf BUF1 (N6312, N6302);
not NOT1 (N6313, N6301);
buf BUF1 (N6314, N6297);
buf BUF1 (N6315, N6271);
not NOT1 (N6316, N6315);
nor NOR2 (N6317, N6307, N567);
and AND3 (N6318, N6313, N3925, N2533);
not NOT1 (N6319, N6316);
xor XOR2 (N6320, N6318, N5236);
buf BUF1 (N6321, N6317);
not NOT1 (N6322, N6309);
xor XOR2 (N6323, N6312, N6318);
xor XOR2 (N6324, N6295, N6318);
buf BUF1 (N6325, N6324);
nand NAND4 (N6326, N6320, N3254, N823, N3223);
or OR2 (N6327, N6322, N1329);
nand NAND2 (N6328, N6326, N1604);
xor XOR2 (N6329, N6291, N26);
and AND2 (N6330, N6319, N4818);
buf BUF1 (N6331, N6314);
nand NAND3 (N6332, N6325, N4877, N5336);
nor NOR3 (N6333, N6330, N5927, N4178);
or OR3 (N6334, N6323, N189, N2989);
and AND3 (N6335, N6329, N5660, N5003);
and AND4 (N6336, N6332, N3552, N4707, N2258);
or OR2 (N6337, N6333, N3328);
nand NAND3 (N6338, N6321, N4131, N319);
nand NAND2 (N6339, N6336, N5935);
not NOT1 (N6340, N6328);
xor XOR2 (N6341, N6337, N2839);
xor XOR2 (N6342, N6341, N5361);
nand NAND3 (N6343, N6327, N1482, N173);
and AND4 (N6344, N6311, N2258, N4313, N1738);
nand NAND3 (N6345, N6334, N5070, N2790);
not NOT1 (N6346, N6340);
xor XOR2 (N6347, N6345, N483);
nand NAND2 (N6348, N6346, N4354);
and AND4 (N6349, N6348, N2312, N2675, N1143);
nand NAND4 (N6350, N6347, N3360, N3340, N5566);
xor XOR2 (N6351, N6349, N4385);
and AND2 (N6352, N6343, N3767);
or OR3 (N6353, N6339, N768, N879);
nand NAND2 (N6354, N6335, N2839);
buf BUF1 (N6355, N6350);
nor NOR4 (N6356, N6342, N5009, N5363, N855);
nand NAND4 (N6357, N6353, N5234, N3220, N953);
buf BUF1 (N6358, N6310);
and AND2 (N6359, N6355, N5618);
not NOT1 (N6360, N6351);
nor NOR4 (N6361, N6356, N1714, N4037, N619);
or OR2 (N6362, N6354, N4782);
or OR2 (N6363, N6357, N226);
or OR2 (N6364, N6360, N3351);
not NOT1 (N6365, N6362);
and AND4 (N6366, N6352, N3340, N727, N2065);
nor NOR4 (N6367, N6344, N876, N452, N6128);
and AND2 (N6368, N6364, N1445);
not NOT1 (N6369, N6365);
nor NOR2 (N6370, N6358, N2588);
nand NAND4 (N6371, N6359, N5516, N264, N246);
nand NAND4 (N6372, N6338, N5723, N767, N5787);
or OR2 (N6373, N6372, N1945);
or OR4 (N6374, N6368, N5914, N6331, N151);
buf BUF1 (N6375, N4581);
buf BUF1 (N6376, N6370);
buf BUF1 (N6377, N6371);
nand NAND3 (N6378, N6377, N982, N6265);
nand NAND2 (N6379, N6361, N2052);
and AND4 (N6380, N6374, N5658, N548, N610);
xor XOR2 (N6381, N6366, N4721);
xor XOR2 (N6382, N6378, N5881);
and AND4 (N6383, N6381, N2481, N925, N4360);
buf BUF1 (N6384, N6383);
nor NOR2 (N6385, N6369, N438);
nor NOR4 (N6386, N6373, N2517, N3889, N2094);
not NOT1 (N6387, N6375);
xor XOR2 (N6388, N6385, N3984);
xor XOR2 (N6389, N6363, N6379);
buf BUF1 (N6390, N5414);
nand NAND2 (N6391, N6376, N1851);
nand NAND4 (N6392, N6390, N4961, N1298, N1733);
nand NAND4 (N6393, N6392, N3324, N1278, N1833);
xor XOR2 (N6394, N6382, N3123);
xor XOR2 (N6395, N6387, N4479);
or OR2 (N6396, N6380, N5944);
not NOT1 (N6397, N6396);
and AND4 (N6398, N6388, N6032, N3562, N1293);
xor XOR2 (N6399, N6391, N1828);
xor XOR2 (N6400, N6389, N5141);
or OR3 (N6401, N6367, N1271, N1389);
buf BUF1 (N6402, N6401);
not NOT1 (N6403, N6399);
xor XOR2 (N6404, N6386, N1001);
not NOT1 (N6405, N6402);
buf BUF1 (N6406, N6405);
xor XOR2 (N6407, N6393, N4907);
and AND4 (N6408, N6384, N5632, N1486, N3359);
nand NAND4 (N6409, N6400, N1953, N1771, N5413);
or OR2 (N6410, N6409, N3582);
not NOT1 (N6411, N6395);
nor NOR3 (N6412, N6398, N5073, N761);
not NOT1 (N6413, N6403);
or OR4 (N6414, N6404, N3977, N4485, N3561);
not NOT1 (N6415, N6412);
or OR3 (N6416, N6410, N5974, N162);
or OR2 (N6417, N6408, N6242);
nand NAND3 (N6418, N6407, N5343, N6254);
or OR3 (N6419, N6413, N6418, N1909);
and AND3 (N6420, N6046, N3940, N4448);
buf BUF1 (N6421, N6394);
or OR3 (N6422, N6419, N3762, N4672);
buf BUF1 (N6423, N6411);
not NOT1 (N6424, N6414);
nor NOR4 (N6425, N6420, N1618, N1967, N5729);
buf BUF1 (N6426, N6406);
not NOT1 (N6427, N6426);
not NOT1 (N6428, N6397);
xor XOR2 (N6429, N6425, N2001);
or OR4 (N6430, N6424, N4251, N2195, N5454);
not NOT1 (N6431, N6421);
nor NOR2 (N6432, N6427, N4461);
buf BUF1 (N6433, N6428);
nor NOR3 (N6434, N6417, N1828, N3499);
and AND2 (N6435, N6430, N1841);
buf BUF1 (N6436, N6433);
not NOT1 (N6437, N6416);
xor XOR2 (N6438, N6437, N3233);
and AND3 (N6439, N6436, N3557, N1662);
nor NOR4 (N6440, N6435, N507, N4359, N444);
or OR3 (N6441, N6429, N3866, N5073);
nand NAND4 (N6442, N6440, N948, N6410, N1054);
nor NOR2 (N6443, N6438, N1188);
buf BUF1 (N6444, N6442);
or OR4 (N6445, N6415, N184, N3396, N3579);
and AND3 (N6446, N6423, N4722, N5778);
xor XOR2 (N6447, N6422, N3391);
and AND2 (N6448, N6445, N1859);
and AND4 (N6449, N6434, N5983, N5079, N4914);
and AND3 (N6450, N6447, N265, N4200);
nand NAND2 (N6451, N6443, N705);
not NOT1 (N6452, N6444);
or OR4 (N6453, N6452, N2585, N2289, N1340);
or OR2 (N6454, N6439, N5637);
nand NAND3 (N6455, N6432, N2909, N24);
or OR3 (N6456, N6446, N6151, N3140);
xor XOR2 (N6457, N6431, N918);
xor XOR2 (N6458, N6449, N948);
not NOT1 (N6459, N6456);
and AND2 (N6460, N6448, N5155);
nor NOR2 (N6461, N6450, N5199);
xor XOR2 (N6462, N6441, N4726);
nor NOR4 (N6463, N6455, N578, N2591, N2984);
nand NAND2 (N6464, N6454, N6073);
nor NOR3 (N6465, N6451, N2089, N957);
not NOT1 (N6466, N6461);
and AND2 (N6467, N6464, N4750);
nor NOR3 (N6468, N6462, N4700, N4100);
and AND4 (N6469, N6467, N5970, N5644, N4969);
or OR4 (N6470, N6463, N1587, N2022, N5407);
xor XOR2 (N6471, N6466, N54);
and AND2 (N6472, N6458, N5075);
and AND4 (N6473, N6472, N5283, N6054, N6027);
not NOT1 (N6474, N6469);
buf BUF1 (N6475, N6471);
or OR4 (N6476, N6475, N240, N1154, N597);
and AND3 (N6477, N6460, N3234, N5998);
xor XOR2 (N6478, N6453, N3438);
or OR2 (N6479, N6476, N2922);
buf BUF1 (N6480, N6478);
nand NAND3 (N6481, N6474, N5022, N6421);
not NOT1 (N6482, N6465);
nand NAND4 (N6483, N6473, N6460, N5589, N210);
nand NAND3 (N6484, N6479, N613, N3851);
nor NOR4 (N6485, N6483, N4985, N162, N6208);
or OR2 (N6486, N6457, N4223);
buf BUF1 (N6487, N6482);
not NOT1 (N6488, N6470);
buf BUF1 (N6489, N6481);
and AND2 (N6490, N6484, N1183);
not NOT1 (N6491, N6489);
or OR4 (N6492, N6486, N5429, N3183, N5389);
or OR3 (N6493, N6491, N2998, N3713);
or OR4 (N6494, N6459, N3262, N6015, N5861);
not NOT1 (N6495, N6477);
and AND4 (N6496, N6480, N4601, N2635, N1738);
nor NOR4 (N6497, N6495, N464, N6373, N219);
nor NOR3 (N6498, N6485, N2461, N2627);
not NOT1 (N6499, N6498);
and AND2 (N6500, N6496, N5259);
or OR4 (N6501, N6487, N4920, N1742, N1674);
or OR4 (N6502, N6494, N3328, N5500, N2604);
not NOT1 (N6503, N6490);
xor XOR2 (N6504, N6503, N4730);
or OR3 (N6505, N6488, N262, N3031);
and AND4 (N6506, N6492, N4096, N3197, N5072);
nor NOR4 (N6507, N6506, N5514, N1370, N104);
or OR2 (N6508, N6501, N4083);
nand NAND4 (N6509, N6468, N6039, N940, N2405);
nor NOR2 (N6510, N6500, N139);
xor XOR2 (N6511, N6505, N68);
nand NAND4 (N6512, N6499, N1323, N3338, N1497);
nand NAND4 (N6513, N6511, N3644, N2957, N6266);
xor XOR2 (N6514, N6508, N3720);
xor XOR2 (N6515, N6513, N2124);
nor NOR4 (N6516, N6509, N5894, N2583, N4372);
xor XOR2 (N6517, N6502, N125);
nand NAND4 (N6518, N6497, N2019, N218, N5256);
and AND2 (N6519, N6504, N421);
or OR3 (N6520, N6514, N447, N4158);
buf BUF1 (N6521, N6517);
xor XOR2 (N6522, N6507, N3040);
and AND2 (N6523, N6512, N3116);
buf BUF1 (N6524, N6518);
not NOT1 (N6525, N6510);
and AND4 (N6526, N6524, N29, N1512, N4792);
nor NOR4 (N6527, N6525, N2825, N3303, N1181);
not NOT1 (N6528, N6523);
xor XOR2 (N6529, N6521, N608);
or OR2 (N6530, N6527, N6159);
or OR4 (N6531, N6528, N4808, N432, N2612);
nand NAND3 (N6532, N6515, N842, N4103);
buf BUF1 (N6533, N6520);
or OR2 (N6534, N6531, N26);
or OR3 (N6535, N6533, N3215, N6035);
nor NOR2 (N6536, N6530, N4226);
xor XOR2 (N6537, N6526, N4815);
and AND4 (N6538, N6529, N4731, N4241, N4340);
or OR2 (N6539, N6536, N2141);
or OR4 (N6540, N6538, N3681, N3705, N4779);
not NOT1 (N6541, N6519);
xor XOR2 (N6542, N6532, N3926);
or OR3 (N6543, N6539, N4179, N755);
buf BUF1 (N6544, N6534);
nand NAND2 (N6545, N6544, N2596);
nor NOR2 (N6546, N6540, N3825);
xor XOR2 (N6547, N6535, N2326);
xor XOR2 (N6548, N6522, N18);
xor XOR2 (N6549, N6516, N3208);
and AND2 (N6550, N6543, N2553);
buf BUF1 (N6551, N6548);
nor NOR3 (N6552, N6542, N3277, N5651);
buf BUF1 (N6553, N6550);
nand NAND3 (N6554, N6549, N2255, N1115);
nand NAND3 (N6555, N6553, N552, N1064);
and AND3 (N6556, N6551, N2342, N3777);
xor XOR2 (N6557, N6545, N3698);
not NOT1 (N6558, N6555);
xor XOR2 (N6559, N6546, N1781);
xor XOR2 (N6560, N6557, N401);
or OR2 (N6561, N6537, N4092);
not NOT1 (N6562, N6558);
and AND4 (N6563, N6556, N1902, N3111, N1354);
xor XOR2 (N6564, N6559, N3316);
xor XOR2 (N6565, N6493, N5383);
or OR4 (N6566, N6554, N1331, N4101, N3336);
and AND3 (N6567, N6560, N4442, N5439);
or OR4 (N6568, N6552, N2651, N387, N2959);
nor NOR2 (N6569, N6568, N4808);
or OR3 (N6570, N6564, N3375, N479);
not NOT1 (N6571, N6567);
nand NAND3 (N6572, N6571, N5273, N1491);
buf BUF1 (N6573, N6566);
xor XOR2 (N6574, N6561, N6496);
nand NAND3 (N6575, N6569, N5557, N4039);
and AND4 (N6576, N6575, N3826, N5553, N459);
or OR2 (N6577, N6570, N3721);
nor NOR4 (N6578, N6563, N24, N5375, N1814);
and AND2 (N6579, N6576, N3348);
nor NOR4 (N6580, N6579, N3649, N3708, N4872);
buf BUF1 (N6581, N6580);
and AND4 (N6582, N6574, N4497, N87, N1545);
or OR2 (N6583, N6581, N3771);
not NOT1 (N6584, N6577);
nand NAND3 (N6585, N6582, N4772, N4613);
not NOT1 (N6586, N6585);
nor NOR2 (N6587, N6565, N374);
xor XOR2 (N6588, N6573, N1830);
nor NOR2 (N6589, N6547, N4712);
xor XOR2 (N6590, N6572, N5811);
buf BUF1 (N6591, N6588);
xor XOR2 (N6592, N6586, N899);
buf BUF1 (N6593, N6584);
xor XOR2 (N6594, N6583, N3457);
nor NOR3 (N6595, N6594, N3491, N631);
or OR2 (N6596, N6562, N6495);
and AND3 (N6597, N6596, N2530, N2665);
nand NAND3 (N6598, N6578, N3862, N4817);
or OR2 (N6599, N6591, N5279);
buf BUF1 (N6600, N6592);
not NOT1 (N6601, N6589);
and AND2 (N6602, N6598, N2146);
xor XOR2 (N6603, N6595, N1286);
nor NOR4 (N6604, N6541, N3247, N6479, N1855);
nand NAND3 (N6605, N6603, N3386, N548);
and AND3 (N6606, N6605, N1410, N1063);
nor NOR3 (N6607, N6587, N4826, N2370);
nor NOR3 (N6608, N6590, N5080, N1329);
buf BUF1 (N6609, N6599);
nor NOR2 (N6610, N6607, N3595);
nor NOR3 (N6611, N6597, N3404, N2556);
and AND4 (N6612, N6601, N3391, N2773, N3972);
and AND3 (N6613, N6609, N3078, N5949);
or OR3 (N6614, N6602, N741, N5355);
xor XOR2 (N6615, N6606, N3145);
and AND2 (N6616, N6610, N3886);
or OR3 (N6617, N6614, N4133, N2283);
buf BUF1 (N6618, N6616);
not NOT1 (N6619, N6613);
and AND2 (N6620, N6617, N774);
nand NAND4 (N6621, N6612, N2009, N4461, N4558);
buf BUF1 (N6622, N6615);
xor XOR2 (N6623, N6622, N6316);
or OR2 (N6624, N6619, N6158);
buf BUF1 (N6625, N6621);
not NOT1 (N6626, N6623);
buf BUF1 (N6627, N6611);
nand NAND3 (N6628, N6627, N5075, N4393);
or OR4 (N6629, N6625, N3557, N1743, N5693);
and AND2 (N6630, N6629, N6496);
or OR3 (N6631, N6626, N2257, N2021);
xor XOR2 (N6632, N6620, N746);
not NOT1 (N6633, N6618);
and AND4 (N6634, N6631, N4339, N6503, N4690);
nand NAND4 (N6635, N6632, N3595, N2168, N2546);
or OR4 (N6636, N6634, N5226, N6378, N3491);
or OR2 (N6637, N6628, N2505);
and AND2 (N6638, N6633, N1547);
or OR4 (N6639, N6593, N2457, N6397, N4648);
and AND3 (N6640, N6637, N1839, N3080);
nor NOR3 (N6641, N6639, N849, N6402);
and AND4 (N6642, N6638, N3502, N4923, N593);
or OR2 (N6643, N6635, N2318);
and AND2 (N6644, N6608, N6428);
and AND4 (N6645, N6643, N4518, N4650, N3594);
buf BUF1 (N6646, N6624);
nor NOR3 (N6647, N6600, N3700, N1147);
or OR2 (N6648, N6644, N6404);
or OR3 (N6649, N6630, N3613, N3940);
nor NOR2 (N6650, N6640, N5264);
or OR3 (N6651, N6650, N3120, N2641);
or OR3 (N6652, N6647, N538, N4343);
nor NOR2 (N6653, N6652, N5200);
and AND3 (N6654, N6641, N1470, N6112);
not NOT1 (N6655, N6645);
nand NAND4 (N6656, N6654, N2395, N3264, N5077);
or OR3 (N6657, N6646, N3062, N4270);
nand NAND3 (N6658, N6642, N5089, N439);
nand NAND2 (N6659, N6648, N3864);
and AND2 (N6660, N6656, N5679);
or OR2 (N6661, N6604, N565);
or OR3 (N6662, N6655, N1885, N3298);
not NOT1 (N6663, N6649);
or OR2 (N6664, N6653, N2920);
nor NOR4 (N6665, N6660, N395, N1665, N4182);
nor NOR3 (N6666, N6661, N5635, N1914);
nor NOR3 (N6667, N6664, N2251, N2615);
buf BUF1 (N6668, N6665);
buf BUF1 (N6669, N6662);
nand NAND2 (N6670, N6651, N4513);
or OR3 (N6671, N6668, N5297, N2118);
nand NAND2 (N6672, N6667, N97);
nor NOR4 (N6673, N6672, N796, N6416, N6275);
xor XOR2 (N6674, N6663, N628);
and AND4 (N6675, N6658, N577, N4541, N1398);
buf BUF1 (N6676, N6659);
xor XOR2 (N6677, N6670, N5252);
buf BUF1 (N6678, N6666);
xor XOR2 (N6679, N6669, N6074);
buf BUF1 (N6680, N6677);
and AND3 (N6681, N6674, N429, N5409);
xor XOR2 (N6682, N6679, N6219);
or OR3 (N6683, N6676, N688, N2281);
nand NAND2 (N6684, N6683, N1096);
and AND3 (N6685, N6680, N480, N1813);
xor XOR2 (N6686, N6682, N769);
xor XOR2 (N6687, N6636, N110);
buf BUF1 (N6688, N6678);
or OR4 (N6689, N6657, N3318, N606, N6274);
buf BUF1 (N6690, N6686);
not NOT1 (N6691, N6673);
xor XOR2 (N6692, N6684, N2858);
buf BUF1 (N6693, N6691);
nor NOR2 (N6694, N6687, N6097);
xor XOR2 (N6695, N6694, N5972);
nor NOR3 (N6696, N6689, N5382, N2848);
nor NOR2 (N6697, N6685, N2936);
buf BUF1 (N6698, N6688);
xor XOR2 (N6699, N6697, N5880);
xor XOR2 (N6700, N6695, N4861);
buf BUF1 (N6701, N6675);
nor NOR2 (N6702, N6692, N5511);
not NOT1 (N6703, N6693);
xor XOR2 (N6704, N6690, N509);
buf BUF1 (N6705, N6698);
buf BUF1 (N6706, N6699);
nor NOR2 (N6707, N6704, N6263);
nor NOR2 (N6708, N6701, N3351);
buf BUF1 (N6709, N6700);
buf BUF1 (N6710, N6696);
and AND2 (N6711, N6708, N31);
xor XOR2 (N6712, N6707, N1944);
xor XOR2 (N6713, N6711, N2874);
nand NAND4 (N6714, N6706, N383, N1358, N3748);
nor NOR2 (N6715, N6671, N5261);
or OR2 (N6716, N6709, N6228);
or OR2 (N6717, N6715, N1880);
nand NAND3 (N6718, N6712, N4841, N3200);
nor NOR2 (N6719, N6705, N1537);
nand NAND4 (N6720, N6702, N4178, N2108, N1973);
nor NOR2 (N6721, N6703, N57);
not NOT1 (N6722, N6714);
not NOT1 (N6723, N6721);
nor NOR2 (N6724, N6719, N1890);
buf BUF1 (N6725, N6724);
nand NAND2 (N6726, N6681, N6616);
nor NOR3 (N6727, N6718, N659, N3178);
and AND4 (N6728, N6710, N5668, N2929, N4315);
xor XOR2 (N6729, N6722, N312);
xor XOR2 (N6730, N6725, N6028);
nor NOR3 (N6731, N6720, N6653, N1555);
or OR2 (N6732, N6723, N1673);
not NOT1 (N6733, N6728);
not NOT1 (N6734, N6727);
nand NAND3 (N6735, N6731, N3708, N3286);
nand NAND2 (N6736, N6730, N4273);
nor NOR4 (N6737, N6733, N5804, N1692, N4091);
buf BUF1 (N6738, N6736);
nand NAND2 (N6739, N6713, N911);
not NOT1 (N6740, N6737);
and AND4 (N6741, N6740, N1330, N6591, N3445);
not NOT1 (N6742, N6734);
not NOT1 (N6743, N6742);
nor NOR4 (N6744, N6741, N787, N946, N787);
xor XOR2 (N6745, N6735, N2330);
nor NOR4 (N6746, N6716, N625, N5255, N1773);
or OR3 (N6747, N6729, N5390, N5654);
nand NAND2 (N6748, N6747, N4761);
nor NOR3 (N6749, N6732, N6689, N2010);
nand NAND3 (N6750, N6743, N111, N6340);
and AND4 (N6751, N6750, N4794, N2276, N2524);
or OR3 (N6752, N6748, N5548, N4382);
and AND3 (N6753, N6738, N2264, N2702);
and AND4 (N6754, N6749, N3506, N3863, N2464);
nand NAND2 (N6755, N6752, N5142);
nand NAND3 (N6756, N6745, N2347, N4255);
nor NOR2 (N6757, N6717, N1399);
buf BUF1 (N6758, N6751);
not NOT1 (N6759, N6758);
and AND2 (N6760, N6759, N2453);
xor XOR2 (N6761, N6760, N3501);
nand NAND3 (N6762, N6757, N501, N33);
xor XOR2 (N6763, N6755, N5723);
and AND4 (N6764, N6763, N5137, N3598, N1793);
xor XOR2 (N6765, N6739, N620);
and AND3 (N6766, N6756, N5882, N4985);
or OR2 (N6767, N6726, N2227);
buf BUF1 (N6768, N6762);
buf BUF1 (N6769, N6767);
nor NOR3 (N6770, N6765, N4923, N6243);
and AND3 (N6771, N6769, N3769, N2832);
nand NAND4 (N6772, N6746, N3556, N2204, N2556);
and AND3 (N6773, N6753, N5057, N3052);
xor XOR2 (N6774, N6772, N3609);
and AND2 (N6775, N6764, N504);
or OR2 (N6776, N6773, N1879);
buf BUF1 (N6777, N6754);
nand NAND4 (N6778, N6770, N5486, N1513, N595);
nor NOR2 (N6779, N6778, N1892);
and AND4 (N6780, N6777, N3327, N995, N5609);
buf BUF1 (N6781, N6779);
and AND3 (N6782, N6781, N1005, N1978);
nor NOR3 (N6783, N6766, N2501, N5702);
and AND4 (N6784, N6771, N5694, N296, N2278);
xor XOR2 (N6785, N6774, N5141);
or OR4 (N6786, N6783, N6662, N2258, N2936);
nand NAND2 (N6787, N6768, N6662);
and AND4 (N6788, N6776, N3457, N992, N1195);
not NOT1 (N6789, N6782);
or OR4 (N6790, N6789, N2510, N516, N4373);
not NOT1 (N6791, N6787);
or OR3 (N6792, N6744, N1083, N239);
and AND3 (N6793, N6786, N3640, N5043);
nand NAND4 (N6794, N6790, N6595, N4493, N2000);
nand NAND4 (N6795, N6784, N5053, N62, N6301);
buf BUF1 (N6796, N6791);
and AND4 (N6797, N6788, N2938, N5070, N1313);
not NOT1 (N6798, N6796);
and AND4 (N6799, N6794, N2655, N6294, N1158);
buf BUF1 (N6800, N6792);
buf BUF1 (N6801, N6780);
xor XOR2 (N6802, N6785, N5987);
xor XOR2 (N6803, N6802, N1762);
and AND2 (N6804, N6761, N5736);
not NOT1 (N6805, N6799);
not NOT1 (N6806, N6800);
nor NOR2 (N6807, N6803, N707);
buf BUF1 (N6808, N6807);
buf BUF1 (N6809, N6805);
nand NAND4 (N6810, N6797, N681, N144, N3655);
xor XOR2 (N6811, N6809, N6449);
and AND2 (N6812, N6810, N5784);
or OR2 (N6813, N6793, N1225);
buf BUF1 (N6814, N6808);
nand NAND4 (N6815, N6804, N6461, N1725, N2336);
nand NAND4 (N6816, N6812, N1676, N3796, N4302);
not NOT1 (N6817, N6795);
nand NAND2 (N6818, N6798, N919);
nand NAND4 (N6819, N6817, N1967, N6760, N6744);
nor NOR2 (N6820, N6815, N5953);
and AND2 (N6821, N6801, N4583);
xor XOR2 (N6822, N6821, N5923);
buf BUF1 (N6823, N6822);
or OR2 (N6824, N6823, N5082);
xor XOR2 (N6825, N6814, N2662);
nand NAND3 (N6826, N6816, N440, N582);
xor XOR2 (N6827, N6819, N5584);
and AND3 (N6828, N6824, N1624, N6629);
and AND4 (N6829, N6825, N401, N4549, N4987);
and AND3 (N6830, N6829, N4303, N6793);
buf BUF1 (N6831, N6828);
not NOT1 (N6832, N6775);
nor NOR2 (N6833, N6820, N5341);
nor NOR4 (N6834, N6811, N5425, N5, N1412);
buf BUF1 (N6835, N6831);
buf BUF1 (N6836, N6833);
and AND2 (N6837, N6813, N1805);
not NOT1 (N6838, N6818);
and AND2 (N6839, N6832, N6230);
or OR4 (N6840, N6806, N1128, N3609, N1607);
not NOT1 (N6841, N6834);
and AND4 (N6842, N6830, N3126, N4242, N1256);
not NOT1 (N6843, N6836);
nand NAND3 (N6844, N6835, N6670, N5918);
buf BUF1 (N6845, N6841);
buf BUF1 (N6846, N6837);
nand NAND3 (N6847, N6840, N6545, N6297);
and AND2 (N6848, N6842, N4419);
buf BUF1 (N6849, N6843);
not NOT1 (N6850, N6847);
buf BUF1 (N6851, N6848);
not NOT1 (N6852, N6826);
not NOT1 (N6853, N6852);
nor NOR2 (N6854, N6853, N1343);
nor NOR4 (N6855, N6838, N4603, N6056, N2778);
xor XOR2 (N6856, N6827, N3072);
nor NOR3 (N6857, N6856, N4629, N6525);
buf BUF1 (N6858, N6855);
nand NAND3 (N6859, N6844, N5673, N6836);
nand NAND4 (N6860, N6858, N3666, N1739, N1328);
xor XOR2 (N6861, N6850, N2738);
or OR3 (N6862, N6839, N3751, N6832);
nor NOR4 (N6863, N6860, N3329, N2896, N458);
xor XOR2 (N6864, N6862, N533);
nor NOR2 (N6865, N6864, N5365);
not NOT1 (N6866, N6849);
nand NAND4 (N6867, N6859, N1208, N6691, N5455);
xor XOR2 (N6868, N6865, N4507);
or OR2 (N6869, N6854, N3874);
or OR2 (N6870, N6857, N5608);
not NOT1 (N6871, N6863);
xor XOR2 (N6872, N6869, N4392);
xor XOR2 (N6873, N6867, N4395);
nor NOR3 (N6874, N6846, N4869, N4786);
not NOT1 (N6875, N6874);
xor XOR2 (N6876, N6870, N344);
xor XOR2 (N6877, N6845, N5337);
nand NAND3 (N6878, N6866, N2311, N1352);
not NOT1 (N6879, N6871);
buf BUF1 (N6880, N6861);
nand NAND4 (N6881, N6880, N5446, N2734, N6429);
nor NOR2 (N6882, N6873, N4143);
nor NOR4 (N6883, N6882, N3262, N6052, N5188);
or OR4 (N6884, N6879, N1084, N5995, N2250);
and AND4 (N6885, N6881, N4321, N6721, N4490);
not NOT1 (N6886, N6878);
nor NOR3 (N6887, N6868, N5602, N6874);
xor XOR2 (N6888, N6885, N4790);
xor XOR2 (N6889, N6876, N1352);
nor NOR3 (N6890, N6886, N5181, N703);
or OR2 (N6891, N6872, N3902);
xor XOR2 (N6892, N6887, N2862);
not NOT1 (N6893, N6892);
buf BUF1 (N6894, N6875);
or OR3 (N6895, N6893, N4751, N3668);
buf BUF1 (N6896, N6883);
or OR2 (N6897, N6851, N4850);
buf BUF1 (N6898, N6889);
xor XOR2 (N6899, N6898, N4815);
or OR2 (N6900, N6895, N4805);
buf BUF1 (N6901, N6891);
and AND2 (N6902, N6896, N6553);
xor XOR2 (N6903, N6894, N4887);
xor XOR2 (N6904, N6884, N1550);
xor XOR2 (N6905, N6897, N4279);
xor XOR2 (N6906, N6888, N223);
nand NAND3 (N6907, N6890, N5607, N3271);
and AND4 (N6908, N6900, N4062, N3939, N2795);
nand NAND4 (N6909, N6904, N558, N3309, N5283);
buf BUF1 (N6910, N6899);
buf BUF1 (N6911, N6903);
xor XOR2 (N6912, N6902, N729);
and AND3 (N6913, N6911, N6009, N1380);
or OR4 (N6914, N6908, N3362, N2478, N1156);
nor NOR2 (N6915, N6914, N1903);
buf BUF1 (N6916, N6907);
and AND4 (N6917, N6905, N239, N609, N4228);
or OR2 (N6918, N6915, N6741);
or OR4 (N6919, N6917, N4496, N1611, N1472);
or OR4 (N6920, N6910, N2214, N6778, N3407);
or OR2 (N6921, N6909, N1159);
and AND4 (N6922, N6877, N5579, N3371, N6121);
and AND3 (N6923, N6901, N39, N811);
or OR3 (N6924, N6921, N2001, N2914);
nor NOR4 (N6925, N6923, N1843, N3813, N4648);
and AND3 (N6926, N6906, N1656, N3984);
xor XOR2 (N6927, N6913, N1220);
nand NAND3 (N6928, N6924, N1714, N161);
not NOT1 (N6929, N6919);
nor NOR4 (N6930, N6926, N303, N5132, N3453);
xor XOR2 (N6931, N6927, N3577);
xor XOR2 (N6932, N6918, N5008);
nand NAND2 (N6933, N6930, N2202);
buf BUF1 (N6934, N6916);
buf BUF1 (N6935, N6912);
nor NOR4 (N6936, N6920, N3262, N5769, N1642);
not NOT1 (N6937, N6922);
nor NOR2 (N6938, N6931, N2174);
buf BUF1 (N6939, N6933);
xor XOR2 (N6940, N6928, N2948);
xor XOR2 (N6941, N6940, N5747);
buf BUF1 (N6942, N6925);
nor NOR3 (N6943, N6938, N4576, N5095);
not NOT1 (N6944, N6943);
xor XOR2 (N6945, N6944, N265);
nor NOR4 (N6946, N6932, N606, N2741, N3042);
buf BUF1 (N6947, N6942);
nand NAND3 (N6948, N6946, N4810, N1246);
xor XOR2 (N6949, N6945, N4217);
xor XOR2 (N6950, N6937, N720);
or OR4 (N6951, N6950, N802, N2375, N6860);
not NOT1 (N6952, N6936);
buf BUF1 (N6953, N6929);
nor NOR2 (N6954, N6949, N1205);
nor NOR2 (N6955, N6935, N5814);
nand NAND2 (N6956, N6947, N5461);
and AND3 (N6957, N6956, N205, N4176);
xor XOR2 (N6958, N6939, N6020);
or OR2 (N6959, N6951, N1029);
nand NAND4 (N6960, N6958, N4382, N5233, N998);
not NOT1 (N6961, N6954);
nor NOR4 (N6962, N6960, N5095, N4568, N5841);
xor XOR2 (N6963, N6941, N5676);
buf BUF1 (N6964, N6959);
nand NAND3 (N6965, N6934, N4663, N4249);
buf BUF1 (N6966, N6963);
nor NOR3 (N6967, N6948, N4589, N6821);
or OR2 (N6968, N6952, N5442);
nor NOR3 (N6969, N6957, N4590, N307);
nand NAND3 (N6970, N6955, N2016, N6016);
nand NAND4 (N6971, N6962, N3206, N6194, N4283);
not NOT1 (N6972, N6964);
xor XOR2 (N6973, N6966, N234);
nor NOR3 (N6974, N6953, N5830, N3607);
buf BUF1 (N6975, N6973);
buf BUF1 (N6976, N6968);
buf BUF1 (N6977, N6974);
and AND3 (N6978, N6967, N4477, N6958);
not NOT1 (N6979, N6978);
nor NOR4 (N6980, N6977, N1113, N4595, N6835);
nand NAND3 (N6981, N6969, N1972, N1282);
nor NOR4 (N6982, N6979, N6464, N4181, N2580);
xor XOR2 (N6983, N6982, N4106);
not NOT1 (N6984, N6976);
nand NAND3 (N6985, N6965, N2228, N5810);
and AND4 (N6986, N6970, N5555, N2354, N4169);
not NOT1 (N6987, N6985);
buf BUF1 (N6988, N6986);
xor XOR2 (N6989, N6987, N2812);
buf BUF1 (N6990, N6975);
and AND2 (N6991, N6984, N6010);
or OR4 (N6992, N6983, N3813, N2470, N1223);
buf BUF1 (N6993, N6981);
nand NAND2 (N6994, N6992, N3550);
or OR4 (N6995, N6988, N6054, N4999, N6121);
or OR4 (N6996, N6961, N4793, N5889, N923);
or OR4 (N6997, N6993, N3298, N5375, N6319);
xor XOR2 (N6998, N6996, N828);
not NOT1 (N6999, N6971);
or OR2 (N7000, N6995, N5124);
nor NOR3 (N7001, N6989, N2070, N2227);
or OR2 (N7002, N6994, N4911);
nor NOR4 (N7003, N6991, N495, N329, N1199);
nand NAND4 (N7004, N7000, N1800, N4302, N2506);
not NOT1 (N7005, N6997);
nand NAND4 (N7006, N7004, N3671, N3661, N3783);
xor XOR2 (N7007, N7002, N964);
nand NAND4 (N7008, N6980, N436, N6188, N70);
nand NAND3 (N7009, N6999, N5705, N3560);
nor NOR4 (N7010, N7003, N446, N5482, N5614);
not NOT1 (N7011, N7009);
nor NOR3 (N7012, N7010, N6739, N5869);
nand NAND2 (N7013, N6972, N2149);
not NOT1 (N7014, N7006);
and AND4 (N7015, N7005, N2711, N2166, N3576);
xor XOR2 (N7016, N7007, N1146);
or OR3 (N7017, N7001, N5835, N472);
buf BUF1 (N7018, N7016);
and AND4 (N7019, N7014, N1287, N5228, N5587);
nor NOR3 (N7020, N7012, N4986, N1605);
or OR4 (N7021, N7013, N1850, N3942, N6215);
buf BUF1 (N7022, N7018);
not NOT1 (N7023, N7015);
or OR4 (N7024, N7019, N4319, N112, N2483);
or OR3 (N7025, N7020, N6066, N5005);
buf BUF1 (N7026, N7022);
and AND2 (N7027, N6998, N3639);
and AND3 (N7028, N6990, N3798, N208);
xor XOR2 (N7029, N7027, N3578);
nand NAND2 (N7030, N7025, N4241);
and AND4 (N7031, N7028, N3511, N2297, N3724);
xor XOR2 (N7032, N7008, N4921);
or OR4 (N7033, N7024, N3252, N5279, N2951);
and AND3 (N7034, N7017, N6268, N4182);
and AND4 (N7035, N7021, N6889, N2198, N6869);
not NOT1 (N7036, N7035);
nor NOR2 (N7037, N7011, N2739);
not NOT1 (N7038, N7023);
nand NAND2 (N7039, N7033, N4970);
nand NAND2 (N7040, N7034, N75);
nand NAND2 (N7041, N7039, N3446);
nor NOR4 (N7042, N7032, N6317, N734, N6102);
xor XOR2 (N7043, N7038, N3120);
and AND2 (N7044, N7037, N1872);
nor NOR3 (N7045, N7029, N4391, N4023);
and AND4 (N7046, N7043, N5672, N904, N2352);
or OR4 (N7047, N7041, N3295, N4448, N3384);
or OR2 (N7048, N7046, N1358);
nor NOR4 (N7049, N7044, N1408, N6676, N435);
nand NAND2 (N7050, N7049, N2159);
nand NAND3 (N7051, N7047, N3115, N5320);
xor XOR2 (N7052, N7030, N2666);
not NOT1 (N7053, N7048);
and AND3 (N7054, N7045, N314, N893);
buf BUF1 (N7055, N7052);
nor NOR2 (N7056, N7053, N1401);
nor NOR3 (N7057, N7040, N1021, N660);
buf BUF1 (N7058, N7031);
and AND3 (N7059, N7036, N6911, N3698);
xor XOR2 (N7060, N7057, N3551);
not NOT1 (N7061, N7060);
nand NAND2 (N7062, N7050, N5175);
nand NAND2 (N7063, N7056, N3335);
buf BUF1 (N7064, N7055);
nand NAND4 (N7065, N7054, N604, N1781, N3340);
xor XOR2 (N7066, N7065, N1397);
nand NAND3 (N7067, N7062, N3130, N2022);
and AND3 (N7068, N7063, N1309, N1528);
nand NAND3 (N7069, N7064, N3088, N6219);
and AND4 (N7070, N7069, N4854, N2035, N6022);
xor XOR2 (N7071, N7066, N2947);
xor XOR2 (N7072, N7067, N6339);
buf BUF1 (N7073, N7071);
or OR2 (N7074, N7051, N5490);
and AND3 (N7075, N7059, N6500, N6770);
or OR3 (N7076, N7026, N2700, N6308);
nor NOR2 (N7077, N7070, N3247);
and AND4 (N7078, N7076, N2843, N7000, N2985);
nand NAND3 (N7079, N7061, N6850, N5592);
and AND2 (N7080, N7072, N1970);
buf BUF1 (N7081, N7042);
buf BUF1 (N7082, N7058);
nand NAND4 (N7083, N7075, N5456, N6263, N2971);
and AND4 (N7084, N7080, N1345, N3560, N4313);
nor NOR3 (N7085, N7081, N1434, N5900);
not NOT1 (N7086, N7083);
xor XOR2 (N7087, N7074, N464);
nand NAND3 (N7088, N7073, N4610, N4208);
and AND2 (N7089, N7082, N3092);
and AND2 (N7090, N7086, N143);
buf BUF1 (N7091, N7068);
buf BUF1 (N7092, N7077);
or OR4 (N7093, N7092, N5654, N6600, N2580);
or OR4 (N7094, N7089, N1408, N2048, N1498);
not NOT1 (N7095, N7094);
nor NOR4 (N7096, N7078, N6251, N3739, N5051);
buf BUF1 (N7097, N7093);
or OR4 (N7098, N7079, N516, N1254, N1260);
nor NOR4 (N7099, N7090, N6770, N2022, N6585);
not NOT1 (N7100, N7084);
nor NOR2 (N7101, N7087, N5901);
not NOT1 (N7102, N7088);
and AND3 (N7103, N7096, N5749, N1120);
nand NAND4 (N7104, N7102, N5977, N3636, N463);
not NOT1 (N7105, N7085);
and AND4 (N7106, N7100, N5092, N2810, N3174);
or OR3 (N7107, N7104, N706, N6106);
and AND2 (N7108, N7097, N1151);
nor NOR4 (N7109, N7107, N200, N2760, N3264);
xor XOR2 (N7110, N7101, N7023);
buf BUF1 (N7111, N7110);
nand NAND4 (N7112, N7099, N485, N5249, N2606);
and AND2 (N7113, N7098, N1650);
or OR2 (N7114, N7105, N6309);
buf BUF1 (N7115, N7106);
xor XOR2 (N7116, N7111, N5836);
buf BUF1 (N7117, N7091);
or OR4 (N7118, N7095, N1482, N3450, N2120);
buf BUF1 (N7119, N7113);
and AND2 (N7120, N7112, N5367);
not NOT1 (N7121, N7118);
buf BUF1 (N7122, N7109);
not NOT1 (N7123, N7119);
or OR4 (N7124, N7116, N2151, N2887, N5595);
nand NAND4 (N7125, N7114, N534, N1504, N921);
or OR4 (N7126, N7124, N616, N5332, N522);
and AND3 (N7127, N7125, N6570, N6077);
nand NAND3 (N7128, N7117, N697, N4555);
buf BUF1 (N7129, N7122);
xor XOR2 (N7130, N7129, N6434);
buf BUF1 (N7131, N7115);
buf BUF1 (N7132, N7123);
and AND4 (N7133, N7126, N6846, N5547, N6084);
or OR2 (N7134, N7132, N691);
nand NAND2 (N7135, N7108, N6907);
nor NOR2 (N7136, N7135, N2728);
nand NAND4 (N7137, N7128, N1661, N1488, N261);
buf BUF1 (N7138, N7121);
nor NOR3 (N7139, N7130, N2271, N369);
nor NOR3 (N7140, N7134, N6347, N1925);
and AND2 (N7141, N7133, N4025);
xor XOR2 (N7142, N7139, N5624);
not NOT1 (N7143, N7137);
buf BUF1 (N7144, N7136);
or OR4 (N7145, N7127, N1771, N5562, N3596);
nor NOR2 (N7146, N7141, N1404);
and AND3 (N7147, N7131, N1729, N6760);
nor NOR2 (N7148, N7120, N3745);
xor XOR2 (N7149, N7146, N4140);
or OR2 (N7150, N7140, N632);
xor XOR2 (N7151, N7150, N635);
nor NOR2 (N7152, N7144, N5472);
or OR2 (N7153, N7147, N4631);
xor XOR2 (N7154, N7143, N4408);
not NOT1 (N7155, N7148);
nand NAND4 (N7156, N7103, N4652, N2773, N4306);
xor XOR2 (N7157, N7152, N783);
not NOT1 (N7158, N7145);
nor NOR2 (N7159, N7142, N6876);
not NOT1 (N7160, N7138);
nand NAND2 (N7161, N7151, N7018);
nand NAND3 (N7162, N7153, N2607, N4751);
and AND2 (N7163, N7154, N5766);
buf BUF1 (N7164, N7155);
nor NOR2 (N7165, N7159, N6757);
not NOT1 (N7166, N7156);
not NOT1 (N7167, N7149);
nand NAND3 (N7168, N7164, N5688, N2434);
nand NAND3 (N7169, N7168, N2414, N2696);
nand NAND4 (N7170, N7162, N6751, N1495, N40);
xor XOR2 (N7171, N7166, N5800);
or OR3 (N7172, N7169, N2074, N670);
nand NAND3 (N7173, N7172, N3677, N674);
buf BUF1 (N7174, N7173);
nand NAND4 (N7175, N7167, N3150, N6337, N3156);
nand NAND2 (N7176, N7171, N4758);
nor NOR2 (N7177, N7165, N4446);
buf BUF1 (N7178, N7176);
not NOT1 (N7179, N7177);
and AND2 (N7180, N7157, N1748);
and AND4 (N7181, N7175, N2224, N5888, N426);
and AND4 (N7182, N7179, N2214, N7092, N5038);
not NOT1 (N7183, N7160);
nor NOR3 (N7184, N7163, N1823, N2200);
xor XOR2 (N7185, N7170, N2318);
xor XOR2 (N7186, N7178, N7073);
buf BUF1 (N7187, N7180);
buf BUF1 (N7188, N7187);
and AND4 (N7189, N7188, N3312, N1482, N1245);
xor XOR2 (N7190, N7185, N4346);
buf BUF1 (N7191, N7183);
nor NOR2 (N7192, N7191, N1790);
or OR2 (N7193, N7184, N1214);
xor XOR2 (N7194, N7189, N3237);
nor NOR4 (N7195, N7192, N745, N6063, N6904);
and AND3 (N7196, N7194, N2086, N3687);
xor XOR2 (N7197, N7174, N6062);
and AND4 (N7198, N7158, N2172, N4047, N2513);
or OR3 (N7199, N7186, N5590, N1532);
and AND2 (N7200, N7193, N4549);
buf BUF1 (N7201, N7200);
buf BUF1 (N7202, N7181);
nand NAND4 (N7203, N7201, N7008, N4247, N1388);
or OR2 (N7204, N7197, N4233);
nand NAND3 (N7205, N7195, N1747, N5904);
and AND3 (N7206, N7190, N3562, N5009);
and AND2 (N7207, N7203, N4450);
nand NAND3 (N7208, N7207, N3913, N2818);
nor NOR2 (N7209, N7182, N7184);
nor NOR2 (N7210, N7204, N7005);
xor XOR2 (N7211, N7210, N1746);
buf BUF1 (N7212, N7202);
buf BUF1 (N7213, N7209);
xor XOR2 (N7214, N7199, N209);
or OR4 (N7215, N7208, N7157, N2868, N4139);
nand NAND2 (N7216, N7212, N4293);
xor XOR2 (N7217, N7214, N6165);
xor XOR2 (N7218, N7205, N1539);
nand NAND2 (N7219, N7213, N4259);
xor XOR2 (N7220, N7217, N2383);
and AND2 (N7221, N7196, N4454);
not NOT1 (N7222, N7206);
not NOT1 (N7223, N7216);
nand NAND3 (N7224, N7222, N3626, N12);
not NOT1 (N7225, N7223);
nand NAND2 (N7226, N7224, N553);
or OR3 (N7227, N7219, N4175, N6438);
and AND2 (N7228, N7227, N6491);
nand NAND3 (N7229, N7221, N5750, N2099);
or OR3 (N7230, N7211, N6289, N6839);
or OR3 (N7231, N7220, N5547, N6572);
and AND2 (N7232, N7198, N2163);
not NOT1 (N7233, N7215);
and AND2 (N7234, N7228, N1099);
nor NOR4 (N7235, N7218, N4916, N224, N5669);
not NOT1 (N7236, N7235);
buf BUF1 (N7237, N7226);
not NOT1 (N7238, N7229);
and AND2 (N7239, N7237, N4879);
buf BUF1 (N7240, N7238);
nor NOR2 (N7241, N7232, N5693);
buf BUF1 (N7242, N7161);
nand NAND4 (N7243, N7233, N4506, N2191, N754);
nand NAND2 (N7244, N7240, N3739);
nand NAND3 (N7245, N7243, N6949, N5961);
nand NAND4 (N7246, N7225, N4605, N7, N3662);
or OR4 (N7247, N7245, N2280, N1942, N436);
nor NOR3 (N7248, N7230, N4102, N4076);
xor XOR2 (N7249, N7236, N3610);
nor NOR4 (N7250, N7249, N7106, N915, N3992);
nor NOR4 (N7251, N7234, N6727, N2558, N3338);
or OR3 (N7252, N7247, N2084, N6568);
or OR4 (N7253, N7239, N1641, N3506, N6065);
or OR2 (N7254, N7241, N3891);
buf BUF1 (N7255, N7252);
xor XOR2 (N7256, N7254, N1908);
buf BUF1 (N7257, N7242);
xor XOR2 (N7258, N7248, N4992);
or OR4 (N7259, N7256, N1138, N5157, N3575);
nor NOR2 (N7260, N7253, N6321);
buf BUF1 (N7261, N7246);
nand NAND3 (N7262, N7258, N2562, N4904);
not NOT1 (N7263, N7262);
not NOT1 (N7264, N7260);
nor NOR3 (N7265, N7255, N2877, N4814);
buf BUF1 (N7266, N7231);
nor NOR3 (N7267, N7265, N3763, N2639);
buf BUF1 (N7268, N7267);
and AND3 (N7269, N7263, N2892, N816);
or OR2 (N7270, N7268, N4473);
nand NAND4 (N7271, N7257, N2689, N3191, N6236);
and AND2 (N7272, N7269, N4992);
not NOT1 (N7273, N7266);
buf BUF1 (N7274, N7251);
nand NAND3 (N7275, N7259, N5237, N3134);
not NOT1 (N7276, N7264);
xor XOR2 (N7277, N7271, N6978);
nand NAND3 (N7278, N7244, N6924, N567);
buf BUF1 (N7279, N7273);
nand NAND2 (N7280, N7250, N5550);
or OR2 (N7281, N7280, N6813);
nor NOR2 (N7282, N7274, N4397);
xor XOR2 (N7283, N7272, N5394);
buf BUF1 (N7284, N7275);
nor NOR2 (N7285, N7281, N6298);
and AND4 (N7286, N7278, N6228, N5305, N2880);
nor NOR3 (N7287, N7282, N1278, N2601);
or OR3 (N7288, N7286, N6483, N3543);
or OR3 (N7289, N7283, N2280, N5236);
nand NAND3 (N7290, N7284, N7217, N2990);
and AND2 (N7291, N7279, N330);
nor NOR4 (N7292, N7287, N6965, N6528, N2728);
xor XOR2 (N7293, N7270, N3499);
not NOT1 (N7294, N7289);
buf BUF1 (N7295, N7276);
nor NOR3 (N7296, N7295, N4058, N7011);
nor NOR3 (N7297, N7294, N2853, N456);
buf BUF1 (N7298, N7291);
not NOT1 (N7299, N7290);
xor XOR2 (N7300, N7277, N1867);
xor XOR2 (N7301, N7293, N1441);
not NOT1 (N7302, N7300);
buf BUF1 (N7303, N7302);
buf BUF1 (N7304, N7296);
or OR4 (N7305, N7285, N7148, N6067, N3449);
and AND2 (N7306, N7298, N3706);
not NOT1 (N7307, N7288);
or OR3 (N7308, N7304, N6447, N189);
or OR3 (N7309, N7299, N3846, N2500);
and AND2 (N7310, N7292, N3992);
xor XOR2 (N7311, N7305, N4517);
xor XOR2 (N7312, N7261, N540);
buf BUF1 (N7313, N7310);
nand NAND2 (N7314, N7313, N2046);
nor NOR3 (N7315, N7308, N1092, N2806);
or OR3 (N7316, N7309, N2094, N420);
xor XOR2 (N7317, N7303, N3495);
buf BUF1 (N7318, N7301);
xor XOR2 (N7319, N7297, N799);
not NOT1 (N7320, N7314);
nor NOR3 (N7321, N7316, N3394, N5843);
and AND2 (N7322, N7321, N4780);
buf BUF1 (N7323, N7319);
not NOT1 (N7324, N7318);
buf BUF1 (N7325, N7320);
not NOT1 (N7326, N7306);
not NOT1 (N7327, N7307);
or OR2 (N7328, N7327, N4013);
not NOT1 (N7329, N7317);
xor XOR2 (N7330, N7324, N3229);
or OR2 (N7331, N7330, N7082);
xor XOR2 (N7332, N7315, N3513);
and AND4 (N7333, N7329, N6033, N3315, N320);
xor XOR2 (N7334, N7311, N3268);
and AND2 (N7335, N7325, N5419);
xor XOR2 (N7336, N7312, N2184);
xor XOR2 (N7337, N7328, N5517);
and AND3 (N7338, N7322, N3151, N4761);
buf BUF1 (N7339, N7336);
nand NAND4 (N7340, N7335, N1498, N1193, N6646);
or OR4 (N7341, N7331, N5618, N452, N2018);
nand NAND4 (N7342, N7338, N3418, N3682, N7110);
and AND3 (N7343, N7333, N1274, N736);
or OR4 (N7344, N7326, N533, N6111, N1708);
xor XOR2 (N7345, N7344, N2103);
and AND3 (N7346, N7342, N101, N5118);
and AND4 (N7347, N7323, N1630, N1067, N383);
or OR3 (N7348, N7343, N1555, N431);
buf BUF1 (N7349, N7347);
xor XOR2 (N7350, N7348, N4727);
xor XOR2 (N7351, N7339, N4937);
buf BUF1 (N7352, N7350);
xor XOR2 (N7353, N7352, N1945);
or OR4 (N7354, N7337, N3888, N5250, N945);
nand NAND4 (N7355, N7345, N3687, N5497, N6705);
and AND2 (N7356, N7332, N7260);
xor XOR2 (N7357, N7353, N3442);
xor XOR2 (N7358, N7346, N2262);
or OR3 (N7359, N7351, N1648, N1548);
nor NOR2 (N7360, N7357, N7015);
and AND4 (N7361, N7341, N7028, N2430, N1349);
nor NOR4 (N7362, N7360, N4509, N6343, N5302);
or OR3 (N7363, N7362, N7216, N6554);
not NOT1 (N7364, N7361);
buf BUF1 (N7365, N7354);
buf BUF1 (N7366, N7359);
nor NOR3 (N7367, N7334, N1313, N2471);
or OR3 (N7368, N7355, N4872, N1822);
not NOT1 (N7369, N7365);
nand NAND4 (N7370, N7358, N7360, N463, N4113);
or OR4 (N7371, N7367, N7223, N2450, N94);
and AND4 (N7372, N7363, N2013, N6481, N3874);
or OR2 (N7373, N7366, N4232);
nor NOR3 (N7374, N7364, N7302, N1788);
nor NOR4 (N7375, N7372, N2437, N2320, N2985);
and AND4 (N7376, N7369, N3549, N5797, N6457);
not NOT1 (N7377, N7376);
buf BUF1 (N7378, N7377);
xor XOR2 (N7379, N7371, N4959);
not NOT1 (N7380, N7370);
not NOT1 (N7381, N7349);
and AND3 (N7382, N7368, N4035, N3039);
not NOT1 (N7383, N7380);
nor NOR3 (N7384, N7378, N7373, N6859);
or OR2 (N7385, N148, N3949);
nand NAND4 (N7386, N7356, N6927, N1487, N5761);
or OR2 (N7387, N7379, N563);
or OR4 (N7388, N7375, N806, N3827, N3264);
nor NOR4 (N7389, N7388, N859, N4326, N1292);
xor XOR2 (N7390, N7374, N4459);
buf BUF1 (N7391, N7382);
and AND2 (N7392, N7384, N3788);
not NOT1 (N7393, N7386);
xor XOR2 (N7394, N7381, N3891);
nand NAND2 (N7395, N7387, N5544);
not NOT1 (N7396, N7393);
or OR4 (N7397, N7385, N1296, N1368, N5200);
and AND4 (N7398, N7389, N6180, N6757, N2557);
nor NOR2 (N7399, N7340, N48);
buf BUF1 (N7400, N7383);
nor NOR2 (N7401, N7397, N6740);
nor NOR4 (N7402, N7394, N5928, N4280, N4826);
and AND2 (N7403, N7395, N5005);
nor NOR4 (N7404, N7403, N7331, N6496, N4009);
not NOT1 (N7405, N7404);
not NOT1 (N7406, N7401);
and AND4 (N7407, N7405, N1772, N3619, N2323);
buf BUF1 (N7408, N7407);
or OR3 (N7409, N7390, N1290, N878);
xor XOR2 (N7410, N7398, N2000);
nor NOR2 (N7411, N7392, N3781);
nor NOR4 (N7412, N7408, N83, N2584, N3691);
and AND4 (N7413, N7400, N3677, N1700, N2763);
xor XOR2 (N7414, N7412, N851);
xor XOR2 (N7415, N7399, N3626);
nor NOR2 (N7416, N7402, N1159);
not NOT1 (N7417, N7406);
buf BUF1 (N7418, N7413);
buf BUF1 (N7419, N7411);
buf BUF1 (N7420, N7410);
not NOT1 (N7421, N7415);
xor XOR2 (N7422, N7421, N5949);
or OR4 (N7423, N7418, N1040, N6727, N7148);
and AND3 (N7424, N7423, N62, N5905);
not NOT1 (N7425, N7417);
not NOT1 (N7426, N7425);
or OR2 (N7427, N7420, N5041);
xor XOR2 (N7428, N7424, N7326);
not NOT1 (N7429, N7409);
and AND2 (N7430, N7429, N4274);
nand NAND2 (N7431, N7427, N1916);
xor XOR2 (N7432, N7422, N1751);
not NOT1 (N7433, N7391);
nor NOR2 (N7434, N7414, N4944);
nand NAND3 (N7435, N7431, N4560, N119);
not NOT1 (N7436, N7432);
xor XOR2 (N7437, N7416, N5130);
and AND4 (N7438, N7437, N5692, N4577, N6965);
nand NAND2 (N7439, N7434, N1523);
not NOT1 (N7440, N7426);
not NOT1 (N7441, N7428);
not NOT1 (N7442, N7419);
nor NOR2 (N7443, N7436, N6715);
nand NAND2 (N7444, N7433, N7397);
not NOT1 (N7445, N7443);
not NOT1 (N7446, N7444);
or OR4 (N7447, N7435, N4056, N1196, N7035);
xor XOR2 (N7448, N7446, N3714);
or OR4 (N7449, N7441, N2356, N258, N4657);
buf BUF1 (N7450, N7449);
and AND4 (N7451, N7448, N2018, N5596, N4681);
nor NOR2 (N7452, N7447, N5876);
nand NAND3 (N7453, N7442, N1976, N2497);
nand NAND3 (N7454, N7450, N4290, N350);
nand NAND2 (N7455, N7439, N4417);
xor XOR2 (N7456, N7455, N5885);
nand NAND3 (N7457, N7438, N2712, N2586);
xor XOR2 (N7458, N7396, N2852);
and AND3 (N7459, N7430, N6679, N270);
nand NAND4 (N7460, N7453, N3327, N849, N7177);
nand NAND2 (N7461, N7458, N1668);
nor NOR2 (N7462, N7461, N5934);
or OR2 (N7463, N7460, N4256);
nor NOR3 (N7464, N7457, N3529, N5150);
and AND3 (N7465, N7462, N2578, N7284);
xor XOR2 (N7466, N7456, N1483);
nor NOR3 (N7467, N7452, N4569, N5908);
xor XOR2 (N7468, N7464, N808);
and AND2 (N7469, N7465, N3340);
and AND3 (N7470, N7451, N7118, N6419);
buf BUF1 (N7471, N7469);
nor NOR3 (N7472, N7454, N7019, N4380);
nor NOR2 (N7473, N7470, N3020);
nand NAND2 (N7474, N7471, N2681);
nand NAND4 (N7475, N7468, N7192, N7182, N3147);
not NOT1 (N7476, N7474);
nor NOR2 (N7477, N7476, N2241);
or OR3 (N7478, N7475, N3075, N6857);
nand NAND3 (N7479, N7445, N2897, N2105);
xor XOR2 (N7480, N7477, N1548);
not NOT1 (N7481, N7467);
or OR3 (N7482, N7481, N4736, N1511);
xor XOR2 (N7483, N7482, N5921);
or OR4 (N7484, N7463, N1822, N2059, N5075);
or OR4 (N7485, N7459, N2601, N1935, N3167);
or OR2 (N7486, N7473, N6300);
buf BUF1 (N7487, N7466);
buf BUF1 (N7488, N7487);
nand NAND2 (N7489, N7488, N6223);
nand NAND2 (N7490, N7478, N54);
not NOT1 (N7491, N7485);
buf BUF1 (N7492, N7480);
nand NAND2 (N7493, N7486, N3884);
xor XOR2 (N7494, N7440, N4008);
buf BUF1 (N7495, N7489);
xor XOR2 (N7496, N7483, N5752);
and AND2 (N7497, N7492, N2219);
nand NAND3 (N7498, N7496, N1315, N2097);
nand NAND3 (N7499, N7479, N2223, N5671);
nor NOR4 (N7500, N7494, N5064, N5688, N5456);
and AND3 (N7501, N7491, N5685, N3688);
or OR4 (N7502, N7484, N3122, N5221, N6983);
nand NAND3 (N7503, N7490, N4401, N6);
nor NOR3 (N7504, N7500, N3122, N4068);
not NOT1 (N7505, N7472);
or OR4 (N7506, N7497, N2895, N5316, N1729);
not NOT1 (N7507, N7495);
nor NOR4 (N7508, N7505, N4402, N6013, N5844);
or OR2 (N7509, N7502, N7268);
xor XOR2 (N7510, N7499, N6384);
buf BUF1 (N7511, N7509);
not NOT1 (N7512, N7493);
buf BUF1 (N7513, N7498);
or OR2 (N7514, N7513, N5066);
not NOT1 (N7515, N7506);
xor XOR2 (N7516, N7508, N3769);
and AND4 (N7517, N7510, N87, N101, N3708);
nand NAND2 (N7518, N7512, N1531);
and AND2 (N7519, N7515, N7201);
or OR4 (N7520, N7511, N5171, N299, N6684);
xor XOR2 (N7521, N7507, N605);
nand NAND2 (N7522, N7503, N3116);
and AND4 (N7523, N7516, N554, N5270, N686);
or OR2 (N7524, N7520, N592);
nand NAND3 (N7525, N7501, N6837, N6163);
not NOT1 (N7526, N7514);
nand NAND4 (N7527, N7519, N4418, N5331, N3349);
not NOT1 (N7528, N7518);
nor NOR2 (N7529, N7525, N4331);
or OR2 (N7530, N7529, N1851);
buf BUF1 (N7531, N7517);
not NOT1 (N7532, N7522);
not NOT1 (N7533, N7521);
nand NAND3 (N7534, N7532, N1866, N105);
nand NAND4 (N7535, N7523, N5303, N648, N3400);
or OR2 (N7536, N7526, N7383);
nor NOR3 (N7537, N7524, N6153, N3160);
buf BUF1 (N7538, N7536);
not NOT1 (N7539, N7528);
or OR4 (N7540, N7534, N5771, N5047, N76);
not NOT1 (N7541, N7533);
xor XOR2 (N7542, N7531, N3511);
buf BUF1 (N7543, N7535);
buf BUF1 (N7544, N7537);
not NOT1 (N7545, N7544);
nor NOR2 (N7546, N7542, N3608);
nor NOR2 (N7547, N7530, N5880);
or OR2 (N7548, N7543, N4379);
xor XOR2 (N7549, N7547, N2193);
and AND2 (N7550, N7527, N3890);
not NOT1 (N7551, N7550);
nor NOR2 (N7552, N7551, N604);
nor NOR2 (N7553, N7541, N5192);
or OR3 (N7554, N7549, N3984, N2162);
and AND4 (N7555, N7554, N711, N6437, N682);
xor XOR2 (N7556, N7546, N4419);
nand NAND3 (N7557, N7556, N2369, N4677);
buf BUF1 (N7558, N7557);
or OR2 (N7559, N7538, N7159);
and AND2 (N7560, N7548, N7152);
buf BUF1 (N7561, N7555);
not NOT1 (N7562, N7560);
xor XOR2 (N7563, N7561, N4711);
and AND2 (N7564, N7545, N5473);
nor NOR4 (N7565, N7559, N5108, N4309, N6778);
and AND3 (N7566, N7558, N3555, N3488);
nor NOR2 (N7567, N7540, N1156);
nand NAND3 (N7568, N7565, N6335, N5900);
buf BUF1 (N7569, N7566);
or OR4 (N7570, N7569, N6479, N952, N2170);
buf BUF1 (N7571, N7504);
buf BUF1 (N7572, N7567);
and AND2 (N7573, N7553, N7139);
or OR4 (N7574, N7552, N667, N7530, N5077);
or OR3 (N7575, N7568, N1996, N2355);
buf BUF1 (N7576, N7539);
buf BUF1 (N7577, N7575);
nor NOR2 (N7578, N7576, N1967);
nand NAND2 (N7579, N7571, N7200);
xor XOR2 (N7580, N7579, N555);
nor NOR3 (N7581, N7570, N806, N2021);
not NOT1 (N7582, N7562);
xor XOR2 (N7583, N7577, N5889);
not NOT1 (N7584, N7572);
xor XOR2 (N7585, N7580, N410);
xor XOR2 (N7586, N7583, N6931);
xor XOR2 (N7587, N7586, N4064);
nor NOR2 (N7588, N7574, N5267);
xor XOR2 (N7589, N7581, N5092);
and AND4 (N7590, N7585, N1168, N3971, N1307);
and AND2 (N7591, N7582, N5104);
not NOT1 (N7592, N7563);
nand NAND2 (N7593, N7584, N6949);
or OR3 (N7594, N7589, N6937, N7547);
nor NOR4 (N7595, N7588, N2099, N5883, N4439);
nand NAND2 (N7596, N7590, N918);
buf BUF1 (N7597, N7587);
not NOT1 (N7598, N7578);
buf BUF1 (N7599, N7598);
and AND3 (N7600, N7594, N2642, N4018);
and AND2 (N7601, N7593, N5655);
and AND4 (N7602, N7573, N131, N2577, N2262);
nor NOR2 (N7603, N7564, N6924);
and AND3 (N7604, N7596, N693, N3270);
nor NOR2 (N7605, N7591, N5456);
nand NAND2 (N7606, N7602, N4375);
not NOT1 (N7607, N7595);
xor XOR2 (N7608, N7599, N4563);
nand NAND2 (N7609, N7601, N6632);
or OR4 (N7610, N7606, N1026, N2666, N7066);
or OR2 (N7611, N7609, N5861);
and AND4 (N7612, N7597, N6158, N1009, N5748);
buf BUF1 (N7613, N7600);
nand NAND2 (N7614, N7607, N6507);
nand NAND2 (N7615, N7614, N5464);
or OR2 (N7616, N7611, N60);
or OR3 (N7617, N7605, N7511, N3733);
buf BUF1 (N7618, N7615);
or OR2 (N7619, N7617, N814);
buf BUF1 (N7620, N7592);
not NOT1 (N7621, N7619);
and AND2 (N7622, N7603, N2931);
or OR2 (N7623, N7618, N5485);
buf BUF1 (N7624, N7622);
and AND3 (N7625, N7616, N148, N6512);
nand NAND4 (N7626, N7613, N5947, N3869, N485);
xor XOR2 (N7627, N7621, N750);
xor XOR2 (N7628, N7625, N6670);
xor XOR2 (N7629, N7604, N4992);
buf BUF1 (N7630, N7612);
or OR4 (N7631, N7620, N4333, N6579, N648);
not NOT1 (N7632, N7610);
not NOT1 (N7633, N7632);
and AND3 (N7634, N7630, N7440, N6441);
not NOT1 (N7635, N7627);
nor NOR3 (N7636, N7629, N7585, N2788);
nand NAND4 (N7637, N7624, N2970, N3358, N3309);
nor NOR3 (N7638, N7634, N2619, N1441);
nand NAND4 (N7639, N7633, N4052, N7166, N288);
not NOT1 (N7640, N7608);
nor NOR4 (N7641, N7638, N1256, N915, N2401);
and AND3 (N7642, N7640, N4724, N4184);
nand NAND4 (N7643, N7626, N5139, N6228, N3297);
not NOT1 (N7644, N7628);
nor NOR3 (N7645, N7637, N2331, N4972);
xor XOR2 (N7646, N7645, N3290);
buf BUF1 (N7647, N7631);
nor NOR2 (N7648, N7623, N4824);
nand NAND3 (N7649, N7642, N239, N2721);
nor NOR3 (N7650, N7648, N2790, N5514);
or OR3 (N7651, N7649, N521, N4100);
xor XOR2 (N7652, N7650, N6277);
buf BUF1 (N7653, N7636);
nand NAND4 (N7654, N7643, N1578, N1269, N143);
nand NAND2 (N7655, N7639, N4673);
nor NOR3 (N7656, N7646, N1783, N3775);
nand NAND2 (N7657, N7647, N1663);
buf BUF1 (N7658, N7656);
xor XOR2 (N7659, N7657, N3451);
buf BUF1 (N7660, N7655);
xor XOR2 (N7661, N7635, N5754);
or OR3 (N7662, N7653, N5599, N2843);
nand NAND2 (N7663, N7651, N2735);
or OR2 (N7664, N7663, N5288);
buf BUF1 (N7665, N7641);
and AND4 (N7666, N7660, N1885, N2881, N657);
and AND3 (N7667, N7665, N6545, N6083);
not NOT1 (N7668, N7652);
xor XOR2 (N7669, N7662, N655);
nand NAND2 (N7670, N7669, N7626);
not NOT1 (N7671, N7661);
nand NAND2 (N7672, N7654, N7108);
nor NOR3 (N7673, N7670, N2533, N6710);
not NOT1 (N7674, N7671);
xor XOR2 (N7675, N7659, N3183);
or OR2 (N7676, N7674, N7126);
buf BUF1 (N7677, N7673);
or OR4 (N7678, N7675, N2740, N1923, N3023);
nand NAND4 (N7679, N7677, N2650, N7362, N4671);
buf BUF1 (N7680, N7664);
xor XOR2 (N7681, N7644, N2666);
and AND3 (N7682, N7680, N6452, N5141);
and AND3 (N7683, N7666, N6595, N3638);
nand NAND2 (N7684, N7678, N5159);
or OR4 (N7685, N7681, N6979, N7623, N7681);
buf BUF1 (N7686, N7676);
not NOT1 (N7687, N7684);
not NOT1 (N7688, N7667);
nand NAND2 (N7689, N7685, N2118);
nand NAND3 (N7690, N7679, N5197, N2661);
xor XOR2 (N7691, N7683, N4339);
or OR4 (N7692, N7672, N7609, N7543, N3365);
or OR4 (N7693, N7682, N4539, N2531, N7681);
nand NAND4 (N7694, N7693, N5616, N3327, N1409);
and AND2 (N7695, N7688, N6847);
nor NOR3 (N7696, N7692, N3904, N2215);
nor NOR4 (N7697, N7694, N4208, N4045, N1024);
not NOT1 (N7698, N7687);
xor XOR2 (N7699, N7689, N1676);
and AND2 (N7700, N7658, N3007);
or OR3 (N7701, N7691, N3980, N759);
not NOT1 (N7702, N7697);
and AND4 (N7703, N7702, N4957, N2998, N7426);
and AND4 (N7704, N7696, N4269, N6684, N1374);
and AND3 (N7705, N7700, N1675, N5165);
nand NAND4 (N7706, N7704, N4025, N983, N5253);
buf BUF1 (N7707, N7698);
and AND4 (N7708, N7706, N1004, N6188, N7204);
xor XOR2 (N7709, N7708, N6680);
nor NOR3 (N7710, N7668, N4232, N6277);
nand NAND3 (N7711, N7699, N6010, N5857);
buf BUF1 (N7712, N7709);
xor XOR2 (N7713, N7690, N1539);
xor XOR2 (N7714, N7707, N4588);
and AND3 (N7715, N7686, N44, N3914);
and AND3 (N7716, N7712, N4478, N4267);
not NOT1 (N7717, N7705);
not NOT1 (N7718, N7714);
or OR2 (N7719, N7701, N3687);
or OR2 (N7720, N7695, N925);
or OR2 (N7721, N7711, N1694);
nor NOR3 (N7722, N7718, N1792, N5400);
nor NOR2 (N7723, N7721, N1533);
buf BUF1 (N7724, N7703);
nor NOR2 (N7725, N7723, N5529);
buf BUF1 (N7726, N7719);
and AND3 (N7727, N7717, N6208, N1578);
xor XOR2 (N7728, N7725, N6553);
xor XOR2 (N7729, N7728, N828);
and AND3 (N7730, N7722, N7128, N6465);
nand NAND2 (N7731, N7713, N4042);
buf BUF1 (N7732, N7730);
xor XOR2 (N7733, N7732, N2787);
xor XOR2 (N7734, N7727, N6566);
not NOT1 (N7735, N7729);
or OR3 (N7736, N7731, N5533, N1872);
buf BUF1 (N7737, N7720);
xor XOR2 (N7738, N7737, N1361);
nor NOR2 (N7739, N7734, N3887);
buf BUF1 (N7740, N7736);
nor NOR2 (N7741, N7738, N7708);
nand NAND4 (N7742, N7716, N2377, N769, N7068);
or OR3 (N7743, N7726, N654, N4066);
nand NAND4 (N7744, N7715, N4221, N471, N5948);
not NOT1 (N7745, N7744);
nor NOR4 (N7746, N7739, N6413, N4924, N1728);
and AND4 (N7747, N7746, N6920, N327, N2787);
buf BUF1 (N7748, N7742);
xor XOR2 (N7749, N7733, N2925);
nand NAND4 (N7750, N7724, N2132, N5791, N5254);
and AND3 (N7751, N7748, N1031, N3693);
not NOT1 (N7752, N7710);
xor XOR2 (N7753, N7741, N7390);
or OR4 (N7754, N7752, N5113, N7247, N587);
or OR2 (N7755, N7750, N811);
nor NOR4 (N7756, N7743, N5239, N5809, N2996);
not NOT1 (N7757, N7751);
buf BUF1 (N7758, N7753);
buf BUF1 (N7759, N7756);
nand NAND3 (N7760, N7754, N7522, N7398);
nand NAND2 (N7761, N7735, N1992);
not NOT1 (N7762, N7747);
or OR2 (N7763, N7758, N3770);
or OR2 (N7764, N7757, N192);
and AND3 (N7765, N7740, N99, N970);
nand NAND2 (N7766, N7749, N1328);
xor XOR2 (N7767, N7761, N501);
nand NAND2 (N7768, N7766, N5484);
xor XOR2 (N7769, N7765, N4961);
xor XOR2 (N7770, N7767, N4562);
buf BUF1 (N7771, N7763);
nand NAND4 (N7772, N7771, N4825, N6345, N4708);
or OR3 (N7773, N7764, N5541, N6627);
nor NOR3 (N7774, N7759, N6445, N2773);
or OR3 (N7775, N7772, N1589, N2037);
xor XOR2 (N7776, N7745, N823);
nand NAND4 (N7777, N7760, N5998, N4169, N3211);
or OR3 (N7778, N7773, N7486, N6660);
or OR2 (N7779, N7755, N6345);
or OR3 (N7780, N7779, N5889, N3647);
and AND2 (N7781, N7762, N829);
or OR2 (N7782, N7775, N2497);
or OR4 (N7783, N7781, N2425, N7232, N7332);
and AND3 (N7784, N7778, N6854, N3817);
buf BUF1 (N7785, N7777);
nand NAND3 (N7786, N7782, N6836, N204);
xor XOR2 (N7787, N7784, N7001);
nor NOR3 (N7788, N7787, N7283, N5392);
nand NAND4 (N7789, N7783, N3598, N1109, N542);
nor NOR3 (N7790, N7788, N731, N6758);
or OR2 (N7791, N7769, N3248);
and AND4 (N7792, N7790, N5678, N7422, N3758);
or OR4 (N7793, N7780, N1175, N6271, N1414);
not NOT1 (N7794, N7774);
nand NAND2 (N7795, N7794, N1280);
xor XOR2 (N7796, N7768, N2775);
not NOT1 (N7797, N7786);
buf BUF1 (N7798, N7797);
or OR2 (N7799, N7791, N1990);
buf BUF1 (N7800, N7796);
nor NOR4 (N7801, N7800, N5244, N2738, N6708);
nand NAND3 (N7802, N7795, N5074, N2938);
nor NOR2 (N7803, N7801, N5496);
buf BUF1 (N7804, N7799);
nor NOR2 (N7805, N7789, N464);
buf BUF1 (N7806, N7785);
nor NOR3 (N7807, N7793, N3788, N951);
xor XOR2 (N7808, N7804, N1942);
and AND2 (N7809, N7806, N323);
nand NAND4 (N7810, N7803, N6890, N1750, N93);
nor NOR4 (N7811, N7770, N5835, N4237, N3370);
and AND4 (N7812, N7809, N7218, N121, N3795);
and AND2 (N7813, N7811, N1251);
not NOT1 (N7814, N7812);
or OR2 (N7815, N7798, N868);
xor XOR2 (N7816, N7805, N3445);
not NOT1 (N7817, N7807);
or OR4 (N7818, N7813, N2772, N2750, N7611);
nand NAND2 (N7819, N7792, N5713);
nand NAND3 (N7820, N7819, N2948, N1221);
nor NOR4 (N7821, N7818, N6796, N2635, N2722);
and AND4 (N7822, N7816, N7254, N1251, N4144);
nand NAND3 (N7823, N7821, N1835, N1465);
not NOT1 (N7824, N7814);
or OR3 (N7825, N7815, N702, N999);
buf BUF1 (N7826, N7825);
nor NOR4 (N7827, N7823, N1292, N910, N6884);
or OR4 (N7828, N7776, N7510, N3474, N4707);
nand NAND3 (N7829, N7827, N7109, N6272);
and AND3 (N7830, N7810, N4458, N393);
xor XOR2 (N7831, N7820, N4903);
or OR2 (N7832, N7828, N3910);
and AND3 (N7833, N7831, N3116, N4457);
not NOT1 (N7834, N7832);
xor XOR2 (N7835, N7822, N3676);
and AND2 (N7836, N7830, N1735);
and AND4 (N7837, N7835, N7073, N7672, N7354);
not NOT1 (N7838, N7833);
xor XOR2 (N7839, N7837, N1411);
not NOT1 (N7840, N7802);
nor NOR2 (N7841, N7838, N4565);
nor NOR4 (N7842, N7817, N6607, N2208, N2486);
nand NAND3 (N7843, N7842, N7811, N6496);
buf BUF1 (N7844, N7839);
and AND2 (N7845, N7843, N1487);
nor NOR2 (N7846, N7841, N2721);
nand NAND4 (N7847, N7844, N825, N786, N4753);
or OR4 (N7848, N7846, N7813, N676, N7638);
and AND3 (N7849, N7824, N1253, N3857);
not NOT1 (N7850, N7829);
buf BUF1 (N7851, N7826);
xor XOR2 (N7852, N7808, N5093);
xor XOR2 (N7853, N7848, N2463);
not NOT1 (N7854, N7853);
xor XOR2 (N7855, N7845, N5887);
buf BUF1 (N7856, N7852);
xor XOR2 (N7857, N7851, N5561);
xor XOR2 (N7858, N7854, N3121);
and AND4 (N7859, N7836, N6769, N3266, N7314);
or OR2 (N7860, N7858, N5206);
or OR2 (N7861, N7860, N6222);
nand NAND2 (N7862, N7857, N1560);
buf BUF1 (N7863, N7862);
nand NAND2 (N7864, N7859, N4996);
or OR4 (N7865, N7847, N3170, N3507, N341);
nand NAND2 (N7866, N7856, N1116);
xor XOR2 (N7867, N7861, N1128);
nand NAND3 (N7868, N7867, N6541, N6466);
nand NAND4 (N7869, N7863, N6486, N6250, N3532);
not NOT1 (N7870, N7834);
nand NAND3 (N7871, N7849, N7061, N15);
and AND2 (N7872, N7869, N396);
nor NOR2 (N7873, N7872, N4771);
not NOT1 (N7874, N7871);
nand NAND4 (N7875, N7840, N6368, N3453, N291);
or OR4 (N7876, N7874, N6081, N63, N271);
and AND2 (N7877, N7868, N7562);
nand NAND3 (N7878, N7866, N6228, N5661);
nand NAND2 (N7879, N7876, N5421);
or OR3 (N7880, N7875, N7594, N3071);
and AND4 (N7881, N7878, N2946, N3564, N1416);
nand NAND4 (N7882, N7864, N602, N1977, N6278);
or OR2 (N7883, N7879, N5744);
xor XOR2 (N7884, N7883, N6861);
buf BUF1 (N7885, N7865);
xor XOR2 (N7886, N7882, N1015);
nand NAND4 (N7887, N7886, N6587, N3879, N4974);
not NOT1 (N7888, N7880);
nor NOR4 (N7889, N7870, N3027, N6535, N3079);
buf BUF1 (N7890, N7885);
not NOT1 (N7891, N7890);
buf BUF1 (N7892, N7891);
or OR3 (N7893, N7887, N7430, N6659);
xor XOR2 (N7894, N7873, N2050);
nand NAND3 (N7895, N7892, N467, N4865);
not NOT1 (N7896, N7895);
buf BUF1 (N7897, N7893);
or OR2 (N7898, N7894, N2331);
nand NAND3 (N7899, N7889, N4916, N7643);
buf BUF1 (N7900, N7884);
or OR4 (N7901, N7896, N6143, N3878, N6633);
buf BUF1 (N7902, N7899);
buf BUF1 (N7903, N7855);
or OR4 (N7904, N7903, N4809, N7848, N3270);
not NOT1 (N7905, N7898);
nor NOR2 (N7906, N7881, N5765);
nand NAND3 (N7907, N7877, N5248, N3769);
or OR3 (N7908, N7907, N4343, N2097);
buf BUF1 (N7909, N7902);
xor XOR2 (N7910, N7906, N5058);
or OR3 (N7911, N7909, N1070, N6409);
nand NAND4 (N7912, N7897, N6489, N6429, N5063);
nand NAND3 (N7913, N7912, N7381, N2970);
not NOT1 (N7914, N7910);
and AND3 (N7915, N7901, N5345, N2417);
and AND2 (N7916, N7913, N912);
and AND4 (N7917, N7888, N1703, N1794, N729);
and AND4 (N7918, N7916, N3239, N5611, N5005);
not NOT1 (N7919, N7900);
buf BUF1 (N7920, N7914);
not NOT1 (N7921, N7850);
buf BUF1 (N7922, N7915);
not NOT1 (N7923, N7919);
not NOT1 (N7924, N7917);
not NOT1 (N7925, N7918);
and AND3 (N7926, N7923, N5627, N5228);
or OR2 (N7927, N7904, N2921);
or OR3 (N7928, N7908, N1058, N491);
or OR3 (N7929, N7925, N6701, N4400);
or OR3 (N7930, N7905, N5776, N2911);
not NOT1 (N7931, N7911);
and AND2 (N7932, N7929, N5518);
or OR3 (N7933, N7922, N5849, N5165);
not NOT1 (N7934, N7928);
nor NOR3 (N7935, N7921, N6182, N1933);
nand NAND4 (N7936, N7920, N1103, N2773, N5114);
or OR2 (N7937, N7933, N701);
and AND4 (N7938, N7934, N1466, N4348, N2323);
xor XOR2 (N7939, N7937, N6724);
nand NAND4 (N7940, N7935, N1380, N7039, N6853);
not NOT1 (N7941, N7939);
and AND4 (N7942, N7927, N5370, N7202, N7125);
nor NOR2 (N7943, N7942, N3783);
nand NAND2 (N7944, N7926, N6007);
xor XOR2 (N7945, N7944, N7254);
and AND3 (N7946, N7932, N4097, N5150);
nand NAND4 (N7947, N7936, N6405, N5966, N1879);
xor XOR2 (N7948, N7943, N449);
nor NOR3 (N7949, N7940, N7868, N2639);
xor XOR2 (N7950, N7947, N2057);
nand NAND3 (N7951, N7931, N3658, N5535);
buf BUF1 (N7952, N7930);
xor XOR2 (N7953, N7941, N2623);
buf BUF1 (N7954, N7950);
nor NOR4 (N7955, N7948, N712, N5373, N1518);
not NOT1 (N7956, N7955);
and AND3 (N7957, N7949, N7701, N6071);
nor NOR3 (N7958, N7954, N7301, N837);
or OR4 (N7959, N7958, N3502, N6316, N1102);
and AND3 (N7960, N7952, N1465, N5105);
buf BUF1 (N7961, N7960);
buf BUF1 (N7962, N7938);
not NOT1 (N7963, N7951);
xor XOR2 (N7964, N7945, N4629);
nand NAND2 (N7965, N7946, N1402);
or OR2 (N7966, N7964, N695);
and AND2 (N7967, N7963, N1561);
buf BUF1 (N7968, N7965);
buf BUF1 (N7969, N7956);
nor NOR4 (N7970, N7924, N6487, N1112, N1385);
or OR2 (N7971, N7962, N1061);
xor XOR2 (N7972, N7969, N4477);
nor NOR3 (N7973, N7959, N2679, N6471);
nand NAND4 (N7974, N7953, N6952, N4668, N5341);
not NOT1 (N7975, N7974);
buf BUF1 (N7976, N7968);
buf BUF1 (N7977, N7971);
xor XOR2 (N7978, N7977, N6004);
xor XOR2 (N7979, N7978, N7794);
xor XOR2 (N7980, N7972, N2124);
xor XOR2 (N7981, N7979, N1098);
and AND3 (N7982, N7981, N5827, N4576);
or OR3 (N7983, N7966, N2906, N847);
nand NAND3 (N7984, N7982, N2341, N1253);
xor XOR2 (N7985, N7973, N3920);
buf BUF1 (N7986, N7975);
buf BUF1 (N7987, N7961);
buf BUF1 (N7988, N7983);
nor NOR4 (N7989, N7957, N4688, N7772, N3321);
xor XOR2 (N7990, N7984, N468);
nor NOR4 (N7991, N7990, N7404, N4733, N2767);
not NOT1 (N7992, N7976);
xor XOR2 (N7993, N7970, N7433);
buf BUF1 (N7994, N7991);
buf BUF1 (N7995, N7967);
not NOT1 (N7996, N7987);
xor XOR2 (N7997, N7995, N2952);
not NOT1 (N7998, N7989);
nor NOR2 (N7999, N7996, N7595);
xor XOR2 (N8000, N7985, N5826);
buf BUF1 (N8001, N8000);
and AND2 (N8002, N8001, N6456);
or OR2 (N8003, N7986, N3711);
or OR3 (N8004, N7992, N2100, N5373);
buf BUF1 (N8005, N7999);
xor XOR2 (N8006, N8002, N7922);
or OR4 (N8007, N8003, N188, N4362, N7563);
and AND3 (N8008, N8007, N5992, N1010);
or OR3 (N8009, N8004, N5087, N3523);
nand NAND3 (N8010, N7988, N1583, N6337);
nor NOR2 (N8011, N7997, N2192);
buf BUF1 (N8012, N7994);
or OR4 (N8013, N7980, N1313, N4415, N2722);
not NOT1 (N8014, N7998);
nor NOR3 (N8015, N8013, N1415, N861);
buf BUF1 (N8016, N8006);
and AND3 (N8017, N8010, N4976, N2921);
buf BUF1 (N8018, N8012);
buf BUF1 (N8019, N8014);
not NOT1 (N8020, N8015);
and AND4 (N8021, N8017, N7154, N273, N2529);
endmodule