// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N3216,N3212,N3200,N3210,N3190,N3214,N3213,N3206,N3207,N3217;

buf BUF1 (N18, N10);
xor XOR2 (N19, N1, N16);
not NOT1 (N20, N8);
not NOT1 (N21, N12);
nor NOR2 (N22, N8, N12);
buf BUF1 (N23, N11);
not NOT1 (N24, N4);
or OR2 (N25, N2, N18);
or OR4 (N26, N7, N25, N19, N14);
and AND2 (N27, N19, N15);
nor NOR3 (N28, N9, N9, N24);
xor XOR2 (N29, N27, N25);
nand NAND2 (N30, N27, N17);
not NOT1 (N31, N22);
not NOT1 (N32, N8);
or OR4 (N33, N28, N16, N14, N18);
and AND4 (N34, N23, N24, N29, N9);
or OR2 (N35, N27, N13);
or OR2 (N36, N27, N10);
xor XOR2 (N37, N21, N20);
not NOT1 (N38, N22);
not NOT1 (N39, N34);
not NOT1 (N40, N37);
nand NAND2 (N41, N32, N21);
and AND2 (N42, N39, N35);
buf BUF1 (N43, N31);
nor NOR3 (N44, N29, N30, N7);
and AND4 (N45, N37, N27, N28, N9);
not NOT1 (N46, N43);
nor NOR3 (N47, N26, N45, N37);
not NOT1 (N48, N35);
xor XOR2 (N49, N40, N2);
nor NOR3 (N50, N38, N32, N11);
nand NAND4 (N51, N41, N10, N15, N41);
and AND3 (N52, N48, N43, N46);
or OR4 (N53, N27, N43, N5, N33);
nand NAND4 (N54, N35, N26, N27, N50);
nand NAND3 (N55, N7, N30, N52);
nor NOR4 (N56, N15, N1, N18, N24);
and AND2 (N57, N47, N11);
nor NOR2 (N58, N57, N49);
nor NOR2 (N59, N32, N28);
or OR4 (N60, N51, N46, N49, N34);
nand NAND2 (N61, N36, N23);
and AND4 (N62, N53, N20, N3, N27);
and AND4 (N63, N62, N3, N14, N37);
xor XOR2 (N64, N59, N32);
not NOT1 (N65, N64);
xor XOR2 (N66, N54, N42);
xor XOR2 (N67, N36, N23);
xor XOR2 (N68, N66, N1);
or OR2 (N69, N60, N39);
and AND4 (N70, N58, N33, N66, N4);
or OR4 (N71, N68, N3, N3, N22);
not NOT1 (N72, N63);
nor NOR4 (N73, N44, N63, N1, N37);
and AND2 (N74, N56, N30);
or OR2 (N75, N61, N56);
not NOT1 (N76, N71);
or OR3 (N77, N75, N49, N31);
not NOT1 (N78, N72);
not NOT1 (N79, N55);
nor NOR3 (N80, N76, N78, N19);
buf BUF1 (N81, N39);
and AND2 (N82, N77, N40);
or OR2 (N83, N70, N57);
or OR3 (N84, N83, N60, N42);
not NOT1 (N85, N67);
xor XOR2 (N86, N65, N11);
and AND4 (N87, N79, N4, N49, N46);
not NOT1 (N88, N84);
and AND2 (N89, N88, N79);
buf BUF1 (N90, N80);
nand NAND2 (N91, N81, N57);
nor NOR2 (N92, N69, N27);
buf BUF1 (N93, N82);
or OR3 (N94, N85, N11, N60);
or OR2 (N95, N92, N55);
xor XOR2 (N96, N90, N21);
or OR4 (N97, N89, N23, N47, N63);
nor NOR4 (N98, N87, N48, N6, N62);
nand NAND3 (N99, N97, N48, N69);
nand NAND3 (N100, N73, N51, N28);
nor NOR2 (N101, N95, N69);
buf BUF1 (N102, N91);
buf BUF1 (N103, N98);
not NOT1 (N104, N96);
or OR4 (N105, N74, N79, N64, N12);
and AND4 (N106, N100, N58, N10, N13);
not NOT1 (N107, N103);
or OR4 (N108, N104, N96, N15, N94);
xor XOR2 (N109, N22, N33);
buf BUF1 (N110, N108);
nand NAND4 (N111, N110, N50, N94, N41);
buf BUF1 (N112, N107);
or OR3 (N113, N99, N60, N99);
xor XOR2 (N114, N86, N6);
not NOT1 (N115, N112);
and AND4 (N116, N101, N37, N78, N49);
and AND4 (N117, N113, N116, N4, N63);
nor NOR4 (N118, N114, N8, N82, N3);
buf BUF1 (N119, N66);
not NOT1 (N120, N93);
or OR3 (N121, N118, N43, N108);
xor XOR2 (N122, N109, N42);
nand NAND3 (N123, N106, N97, N83);
and AND2 (N124, N120, N81);
and AND2 (N125, N121, N90);
nor NOR2 (N126, N124, N37);
buf BUF1 (N127, N117);
not NOT1 (N128, N122);
or OR3 (N129, N123, N90, N123);
buf BUF1 (N130, N127);
buf BUF1 (N131, N105);
nor NOR4 (N132, N128, N46, N69, N85);
and AND4 (N133, N115, N88, N58, N31);
and AND2 (N134, N130, N1);
and AND3 (N135, N119, N42, N35);
or OR2 (N136, N125, N120);
buf BUF1 (N137, N132);
nand NAND4 (N138, N111, N73, N71, N124);
xor XOR2 (N139, N136, N103);
nand NAND4 (N140, N139, N65, N101, N24);
buf BUF1 (N141, N135);
nand NAND3 (N142, N102, N140, N32);
buf BUF1 (N143, N43);
buf BUF1 (N144, N134);
nor NOR3 (N145, N129, N125, N123);
not NOT1 (N146, N145);
xor XOR2 (N147, N131, N122);
nor NOR3 (N148, N147, N22, N96);
and AND4 (N149, N144, N145, N55, N23);
and AND3 (N150, N133, N108, N121);
nand NAND3 (N151, N149, N111, N60);
and AND2 (N152, N137, N50);
or OR2 (N153, N152, N32);
nor NOR4 (N154, N143, N62, N6, N137);
xor XOR2 (N155, N150, N85);
nor NOR2 (N156, N155, N139);
and AND3 (N157, N141, N20, N138);
nor NOR2 (N158, N116, N142);
buf BUF1 (N159, N55);
nand NAND4 (N160, N151, N49, N92, N66);
xor XOR2 (N161, N156, N155);
nor NOR3 (N162, N158, N71, N36);
not NOT1 (N163, N159);
nor NOR2 (N164, N126, N120);
and AND2 (N165, N162, N26);
buf BUF1 (N166, N154);
nor NOR3 (N167, N160, N128, N84);
xor XOR2 (N168, N167, N60);
nand NAND4 (N169, N146, N21, N107, N144);
buf BUF1 (N170, N168);
and AND4 (N171, N165, N117, N88, N22);
xor XOR2 (N172, N148, N166);
nor NOR4 (N173, N38, N35, N132, N31);
and AND4 (N174, N173, N23, N26, N99);
or OR3 (N175, N157, N94, N78);
xor XOR2 (N176, N164, N146);
buf BUF1 (N177, N174);
and AND4 (N178, N177, N73, N5, N74);
nor NOR3 (N179, N171, N156, N41);
not NOT1 (N180, N163);
nand NAND4 (N181, N161, N80, N100, N28);
and AND2 (N182, N179, N29);
or OR4 (N183, N180, N29, N178, N181);
xor XOR2 (N184, N82, N58);
and AND3 (N185, N8, N18, N44);
buf BUF1 (N186, N153);
buf BUF1 (N187, N182);
xor XOR2 (N188, N170, N187);
nand NAND2 (N189, N140, N178);
or OR2 (N190, N183, N104);
and AND2 (N191, N184, N64);
not NOT1 (N192, N185);
nor NOR3 (N193, N192, N29, N98);
or OR2 (N194, N191, N21);
nor NOR4 (N195, N169, N9, N145, N22);
xor XOR2 (N196, N193, N50);
or OR3 (N197, N189, N61, N162);
not NOT1 (N198, N194);
xor XOR2 (N199, N186, N48);
or OR2 (N200, N175, N172);
buf BUF1 (N201, N124);
xor XOR2 (N202, N198, N193);
nand NAND3 (N203, N176, N47, N163);
or OR3 (N204, N201, N21, N100);
nand NAND3 (N205, N195, N44, N30);
nor NOR3 (N206, N197, N141, N118);
buf BUF1 (N207, N200);
not NOT1 (N208, N205);
not NOT1 (N209, N199);
buf BUF1 (N210, N190);
nand NAND2 (N211, N196, N1);
and AND4 (N212, N206, N158, N103, N204);
nand NAND4 (N213, N161, N113, N41, N42);
nand NAND4 (N214, N208, N171, N23, N91);
not NOT1 (N215, N203);
buf BUF1 (N216, N214);
or OR4 (N217, N209, N28, N67, N128);
nand NAND2 (N218, N215, N71);
nand NAND3 (N219, N210, N25, N183);
xor XOR2 (N220, N202, N67);
or OR4 (N221, N217, N69, N2, N205);
nand NAND4 (N222, N218, N35, N66, N33);
nor NOR3 (N223, N220, N172, N106);
xor XOR2 (N224, N221, N1);
or OR2 (N225, N216, N168);
xor XOR2 (N226, N224, N38);
nor NOR4 (N227, N223, N143, N7, N199);
xor XOR2 (N228, N207, N205);
not NOT1 (N229, N228);
nand NAND3 (N230, N226, N99, N41);
and AND3 (N231, N213, N207, N184);
not NOT1 (N232, N212);
nand NAND2 (N233, N229, N94);
nand NAND4 (N234, N219, N171, N218, N169);
buf BUF1 (N235, N211);
or OR3 (N236, N225, N95, N206);
nand NAND3 (N237, N232, N9, N122);
and AND2 (N238, N235, N52);
nor NOR3 (N239, N230, N34, N138);
or OR3 (N240, N239, N107, N48);
and AND3 (N241, N236, N145, N123);
and AND3 (N242, N227, N212, N210);
and AND2 (N243, N231, N201);
and AND3 (N244, N240, N53, N25);
or OR4 (N245, N244, N101, N159, N19);
buf BUF1 (N246, N245);
nor NOR2 (N247, N243, N155);
not NOT1 (N248, N246);
buf BUF1 (N249, N233);
and AND2 (N250, N237, N227);
or OR2 (N251, N188, N187);
buf BUF1 (N252, N242);
and AND2 (N253, N248, N148);
nor NOR3 (N254, N249, N58, N142);
nand NAND4 (N255, N234, N30, N122, N254);
buf BUF1 (N256, N84);
or OR2 (N257, N247, N6);
or OR2 (N258, N251, N14);
nor NOR3 (N259, N258, N252, N68);
not NOT1 (N260, N126);
or OR2 (N261, N241, N9);
or OR2 (N262, N261, N157);
nand NAND4 (N263, N257, N123, N20, N84);
not NOT1 (N264, N222);
and AND4 (N265, N253, N129, N39, N208);
buf BUF1 (N266, N264);
buf BUF1 (N267, N265);
xor XOR2 (N268, N238, N178);
nor NOR2 (N269, N262, N11);
or OR4 (N270, N260, N127, N86, N44);
nand NAND3 (N271, N263, N235, N262);
nand NAND4 (N272, N271, N126, N39, N216);
nor NOR3 (N273, N255, N27, N27);
nand NAND2 (N274, N269, N60);
nand NAND4 (N275, N268, N151, N73, N91);
not NOT1 (N276, N250);
and AND2 (N277, N272, N84);
or OR2 (N278, N256, N137);
or OR3 (N279, N278, N269, N14);
xor XOR2 (N280, N275, N99);
or OR4 (N281, N266, N55, N248, N276);
nor NOR3 (N282, N40, N156, N268);
buf BUF1 (N283, N270);
nor NOR3 (N284, N282, N140, N90);
or OR4 (N285, N274, N239, N259, N197);
nor NOR2 (N286, N260, N184);
nand NAND4 (N287, N283, N265, N45, N11);
nor NOR3 (N288, N287, N173, N115);
nand NAND3 (N289, N288, N129, N202);
or OR4 (N290, N279, N207, N276, N40);
xor XOR2 (N291, N289, N70);
nor NOR4 (N292, N284, N240, N236, N42);
nor NOR2 (N293, N285, N77);
buf BUF1 (N294, N273);
buf BUF1 (N295, N281);
not NOT1 (N296, N277);
not NOT1 (N297, N296);
nor NOR3 (N298, N294, N235, N103);
nand NAND4 (N299, N293, N26, N114, N9);
and AND3 (N300, N286, N147, N244);
xor XOR2 (N301, N300, N39);
buf BUF1 (N302, N292);
not NOT1 (N303, N291);
xor XOR2 (N304, N303, N279);
xor XOR2 (N305, N302, N286);
not NOT1 (N306, N301);
xor XOR2 (N307, N306, N283);
and AND3 (N308, N307, N121, N294);
buf BUF1 (N309, N305);
or OR3 (N310, N298, N239, N166);
or OR2 (N311, N290, N210);
not NOT1 (N312, N309);
xor XOR2 (N313, N297, N301);
xor XOR2 (N314, N299, N100);
not NOT1 (N315, N312);
xor XOR2 (N316, N315, N95);
xor XOR2 (N317, N280, N180);
buf BUF1 (N318, N304);
or OR3 (N319, N310, N134, N129);
nor NOR3 (N320, N267, N139, N286);
buf BUF1 (N321, N318);
or OR4 (N322, N311, N307, N10, N55);
nor NOR4 (N323, N321, N105, N93, N13);
nor NOR3 (N324, N313, N189, N122);
buf BUF1 (N325, N322);
not NOT1 (N326, N314);
buf BUF1 (N327, N325);
or OR2 (N328, N295, N171);
not NOT1 (N329, N317);
xor XOR2 (N330, N329, N178);
or OR2 (N331, N320, N300);
nor NOR2 (N332, N327, N145);
not NOT1 (N333, N316);
nor NOR3 (N334, N333, N129, N306);
buf BUF1 (N335, N334);
nor NOR3 (N336, N308, N214, N53);
xor XOR2 (N337, N326, N58);
buf BUF1 (N338, N331);
xor XOR2 (N339, N328, N201);
not NOT1 (N340, N335);
or OR3 (N341, N324, N287, N5);
and AND4 (N342, N340, N74, N178, N45);
xor XOR2 (N343, N332, N163);
not NOT1 (N344, N342);
nand NAND4 (N345, N339, N330, N81, N140);
buf BUF1 (N346, N155);
buf BUF1 (N347, N336);
and AND2 (N348, N347, N332);
not NOT1 (N349, N344);
not NOT1 (N350, N348);
buf BUF1 (N351, N349);
nor NOR4 (N352, N337, N298, N350, N172);
xor XOR2 (N353, N323, N23);
nor NOR4 (N354, N126, N175, N334, N254);
not NOT1 (N355, N346);
xor XOR2 (N356, N352, N45);
xor XOR2 (N357, N341, N89);
or OR3 (N358, N345, N258, N295);
or OR4 (N359, N354, N350, N105, N70);
or OR3 (N360, N355, N38, N204);
nor NOR4 (N361, N353, N87, N312, N113);
buf BUF1 (N362, N361);
xor XOR2 (N363, N356, N270);
nor NOR4 (N364, N360, N39, N275, N138);
nor NOR2 (N365, N338, N193);
nand NAND2 (N366, N357, N111);
not NOT1 (N367, N351);
and AND2 (N368, N366, N24);
or OR3 (N369, N367, N326, N321);
buf BUF1 (N370, N369);
xor XOR2 (N371, N362, N260);
and AND3 (N372, N319, N146, N75);
xor XOR2 (N373, N370, N31);
or OR4 (N374, N372, N40, N207, N208);
xor XOR2 (N375, N365, N278);
or OR2 (N376, N364, N304);
not NOT1 (N377, N363);
buf BUF1 (N378, N359);
nand NAND2 (N379, N378, N319);
xor XOR2 (N380, N371, N271);
buf BUF1 (N381, N379);
buf BUF1 (N382, N375);
not NOT1 (N383, N377);
nor NOR4 (N384, N380, N109, N127, N168);
and AND3 (N385, N358, N301, N78);
and AND3 (N386, N376, N99, N352);
and AND4 (N387, N374, N100, N281, N241);
or OR3 (N388, N383, N245, N378);
or OR3 (N389, N387, N272, N95);
buf BUF1 (N390, N384);
or OR4 (N391, N388, N12, N136, N290);
nor NOR4 (N392, N381, N267, N262, N190);
buf BUF1 (N393, N392);
and AND3 (N394, N393, N87, N48);
nor NOR4 (N395, N394, N256, N108, N16);
xor XOR2 (N396, N391, N392);
xor XOR2 (N397, N373, N101);
buf BUF1 (N398, N389);
nand NAND3 (N399, N385, N59, N337);
buf BUF1 (N400, N395);
nor NOR3 (N401, N398, N388, N374);
nor NOR3 (N402, N386, N224, N281);
not NOT1 (N403, N400);
nor NOR2 (N404, N399, N221);
xor XOR2 (N405, N401, N121);
xor XOR2 (N406, N396, N2);
xor XOR2 (N407, N405, N85);
xor XOR2 (N408, N404, N315);
nor NOR4 (N409, N403, N212, N311, N274);
not NOT1 (N410, N390);
nor NOR3 (N411, N406, N76, N369);
not NOT1 (N412, N397);
nand NAND4 (N413, N409, N351, N73, N185);
not NOT1 (N414, N412);
or OR3 (N415, N413, N39, N168);
nor NOR2 (N416, N414, N47);
xor XOR2 (N417, N411, N59);
nand NAND3 (N418, N407, N317, N243);
and AND4 (N419, N416, N281, N103, N297);
and AND2 (N420, N415, N244);
and AND2 (N421, N420, N382);
not NOT1 (N422, N18);
or OR3 (N423, N421, N295, N90);
buf BUF1 (N424, N418);
or OR2 (N425, N343, N64);
not NOT1 (N426, N417);
buf BUF1 (N427, N419);
or OR2 (N428, N422, N332);
nor NOR2 (N429, N408, N414);
xor XOR2 (N430, N427, N344);
nor NOR4 (N431, N426, N408, N70, N361);
nor NOR4 (N432, N429, N424, N337, N95);
not NOT1 (N433, N98);
nand NAND3 (N434, N431, N246, N361);
and AND3 (N435, N430, N173, N123);
not NOT1 (N436, N435);
nor NOR4 (N437, N428, N421, N7, N284);
nor NOR2 (N438, N410, N115);
and AND2 (N439, N436, N284);
nand NAND4 (N440, N425, N189, N351, N227);
buf BUF1 (N441, N432);
nand NAND3 (N442, N434, N56, N30);
and AND3 (N443, N439, N194, N267);
and AND4 (N444, N433, N116, N428, N33);
and AND2 (N445, N444, N319);
and AND3 (N446, N402, N410, N228);
nand NAND4 (N447, N443, N241, N229, N78);
nor NOR4 (N448, N441, N139, N406, N109);
nand NAND4 (N449, N442, N235, N411, N66);
nor NOR4 (N450, N448, N102, N71, N444);
buf BUF1 (N451, N368);
and AND2 (N452, N450, N103);
nor NOR4 (N453, N451, N254, N358, N359);
not NOT1 (N454, N453);
not NOT1 (N455, N440);
nand NAND3 (N456, N423, N298, N280);
and AND4 (N457, N449, N265, N26, N192);
xor XOR2 (N458, N454, N293);
and AND2 (N459, N447, N298);
or OR3 (N460, N456, N137, N180);
nand NAND4 (N461, N455, N1, N339, N109);
not NOT1 (N462, N461);
or OR2 (N463, N452, N441);
nand NAND2 (N464, N446, N54);
nor NOR3 (N465, N457, N21, N255);
nor NOR3 (N466, N459, N349, N233);
and AND4 (N467, N438, N424, N307, N408);
buf BUF1 (N468, N465);
nor NOR4 (N469, N460, N23, N447, N248);
buf BUF1 (N470, N469);
nor NOR3 (N471, N470, N398, N72);
xor XOR2 (N472, N463, N247);
or OR4 (N473, N458, N236, N446, N113);
and AND4 (N474, N466, N206, N130, N71);
not NOT1 (N475, N462);
nand NAND3 (N476, N467, N62, N126);
not NOT1 (N477, N472);
and AND3 (N478, N468, N452, N123);
nand NAND4 (N479, N437, N207, N475, N207);
or OR4 (N480, N404, N99, N58, N31);
nor NOR4 (N481, N471, N29, N76, N172);
and AND4 (N482, N477, N152, N284, N245);
nand NAND2 (N483, N445, N334);
xor XOR2 (N484, N483, N457);
buf BUF1 (N485, N481);
buf BUF1 (N486, N482);
and AND4 (N487, N476, N12, N176, N77);
nor NOR3 (N488, N485, N391, N297);
not NOT1 (N489, N479);
buf BUF1 (N490, N486);
and AND2 (N491, N487, N117);
or OR2 (N492, N464, N160);
xor XOR2 (N493, N488, N96);
and AND3 (N494, N474, N342, N400);
nand NAND4 (N495, N473, N482, N154, N433);
buf BUF1 (N496, N484);
or OR2 (N497, N490, N3);
nor NOR3 (N498, N491, N287, N454);
not NOT1 (N499, N496);
nor NOR4 (N500, N493, N259, N334, N323);
nor NOR2 (N501, N489, N198);
or OR3 (N502, N478, N450, N159);
or OR4 (N503, N492, N238, N54, N83);
or OR4 (N504, N497, N46, N211, N398);
xor XOR2 (N505, N500, N396);
xor XOR2 (N506, N498, N249);
and AND3 (N507, N499, N253, N346);
and AND2 (N508, N505, N76);
xor XOR2 (N509, N501, N430);
buf BUF1 (N510, N509);
xor XOR2 (N511, N495, N52);
xor XOR2 (N512, N511, N211);
not NOT1 (N513, N504);
nand NAND2 (N514, N502, N486);
nand NAND3 (N515, N503, N483, N495);
nor NOR2 (N516, N506, N349);
buf BUF1 (N517, N514);
or OR3 (N518, N510, N236, N228);
and AND3 (N519, N508, N254, N422);
xor XOR2 (N520, N519, N156);
xor XOR2 (N521, N512, N196);
nor NOR2 (N522, N480, N516);
xor XOR2 (N523, N100, N277);
nand NAND4 (N524, N518, N520, N396, N265);
nand NAND2 (N525, N214, N132);
not NOT1 (N526, N523);
or OR4 (N527, N517, N472, N76, N63);
nand NAND3 (N528, N524, N24, N209);
or OR4 (N529, N507, N104, N365, N161);
xor XOR2 (N530, N525, N29);
buf BUF1 (N531, N494);
not NOT1 (N532, N515);
nor NOR4 (N533, N528, N217, N501, N346);
xor XOR2 (N534, N530, N8);
or OR4 (N535, N522, N76, N345, N412);
not NOT1 (N536, N532);
buf BUF1 (N537, N534);
nand NAND2 (N538, N513, N185);
buf BUF1 (N539, N521);
nand NAND2 (N540, N538, N277);
not NOT1 (N541, N531);
xor XOR2 (N542, N535, N284);
and AND4 (N543, N533, N356, N46, N399);
and AND4 (N544, N529, N295, N196, N508);
nand NAND4 (N545, N527, N36, N540, N502);
not NOT1 (N546, N324);
or OR4 (N547, N542, N287, N310, N477);
buf BUF1 (N548, N547);
xor XOR2 (N549, N539, N113);
nor NOR4 (N550, N541, N8, N549, N186);
or OR3 (N551, N309, N452, N46);
nor NOR3 (N552, N548, N65, N121);
nand NAND3 (N553, N526, N142, N391);
or OR3 (N554, N552, N64, N362);
nand NAND2 (N555, N537, N265);
nand NAND3 (N556, N554, N200, N294);
or OR4 (N557, N544, N235, N378, N370);
and AND2 (N558, N556, N61);
buf BUF1 (N559, N558);
nor NOR4 (N560, N553, N80, N501, N452);
buf BUF1 (N561, N559);
not NOT1 (N562, N546);
and AND2 (N563, N551, N501);
and AND2 (N564, N536, N298);
and AND2 (N565, N550, N563);
not NOT1 (N566, N92);
buf BUF1 (N567, N560);
and AND4 (N568, N564, N64, N509, N8);
xor XOR2 (N569, N545, N263);
nor NOR4 (N570, N568, N76, N290, N120);
and AND4 (N571, N557, N355, N113, N240);
or OR3 (N572, N555, N7, N527);
nor NOR3 (N573, N567, N131, N345);
buf BUF1 (N574, N543);
nor NOR4 (N575, N569, N98, N222, N220);
nand NAND2 (N576, N574, N553);
nor NOR2 (N577, N575, N248);
buf BUF1 (N578, N572);
buf BUF1 (N579, N576);
buf BUF1 (N580, N571);
nand NAND3 (N581, N580, N10, N380);
and AND4 (N582, N562, N403, N279, N98);
buf BUF1 (N583, N566);
or OR3 (N584, N583, N369, N173);
not NOT1 (N585, N577);
or OR3 (N586, N579, N584, N292);
buf BUF1 (N587, N523);
xor XOR2 (N588, N587, N165);
or OR2 (N589, N586, N52);
and AND4 (N590, N570, N44, N130, N411);
nand NAND3 (N591, N573, N9, N257);
or OR4 (N592, N591, N56, N234, N236);
nor NOR4 (N593, N578, N453, N25, N448);
nor NOR4 (N594, N592, N277, N278, N296);
buf BUF1 (N595, N581);
xor XOR2 (N596, N585, N364);
nor NOR4 (N597, N561, N357, N395, N228);
nor NOR3 (N598, N588, N232, N63);
nand NAND4 (N599, N589, N537, N112, N407);
not NOT1 (N600, N597);
buf BUF1 (N601, N599);
buf BUF1 (N602, N596);
nor NOR2 (N603, N594, N513);
not NOT1 (N604, N593);
buf BUF1 (N605, N595);
buf BUF1 (N606, N600);
nand NAND4 (N607, N606, N247, N534, N69);
nand NAND4 (N608, N602, N443, N243, N249);
and AND3 (N609, N605, N232, N354);
and AND4 (N610, N582, N534, N171, N551);
and AND4 (N611, N609, N317, N314, N129);
nor NOR3 (N612, N604, N456, N544);
nor NOR3 (N613, N608, N484, N111);
nand NAND4 (N614, N598, N495, N549, N299);
or OR2 (N615, N565, N270);
nand NAND4 (N616, N590, N448, N230, N187);
buf BUF1 (N617, N613);
xor XOR2 (N618, N615, N155);
xor XOR2 (N619, N617, N268);
nor NOR3 (N620, N601, N161, N326);
not NOT1 (N621, N618);
xor XOR2 (N622, N621, N498);
nor NOR3 (N623, N610, N610, N225);
buf BUF1 (N624, N616);
nor NOR2 (N625, N603, N18);
or OR2 (N626, N620, N155);
nand NAND3 (N627, N607, N476, N175);
xor XOR2 (N628, N614, N620);
not NOT1 (N629, N624);
nand NAND2 (N630, N627, N263);
and AND4 (N631, N619, N220, N85, N269);
buf BUF1 (N632, N611);
or OR2 (N633, N630, N469);
xor XOR2 (N634, N631, N417);
buf BUF1 (N635, N623);
or OR2 (N636, N633, N430);
not NOT1 (N637, N628);
xor XOR2 (N638, N629, N522);
xor XOR2 (N639, N637, N630);
not NOT1 (N640, N612);
buf BUF1 (N641, N638);
or OR4 (N642, N641, N133, N449, N186);
nand NAND3 (N643, N640, N610, N421);
and AND4 (N644, N636, N63, N195, N529);
nand NAND3 (N645, N639, N545, N557);
and AND3 (N646, N626, N318, N450);
buf BUF1 (N647, N632);
nor NOR4 (N648, N622, N209, N311, N112);
buf BUF1 (N649, N646);
or OR4 (N650, N635, N116, N144, N410);
xor XOR2 (N651, N625, N75);
buf BUF1 (N652, N648);
not NOT1 (N653, N651);
and AND2 (N654, N653, N81);
nor NOR2 (N655, N652, N49);
xor XOR2 (N656, N644, N121);
buf BUF1 (N657, N656);
nor NOR2 (N658, N643, N80);
xor XOR2 (N659, N657, N441);
not NOT1 (N660, N655);
and AND3 (N661, N660, N396, N15);
not NOT1 (N662, N649);
nor NOR4 (N663, N654, N179, N367, N188);
nand NAND4 (N664, N647, N489, N541, N146);
buf BUF1 (N665, N634);
not NOT1 (N666, N665);
and AND2 (N667, N645, N46);
and AND2 (N668, N667, N217);
nand NAND3 (N669, N658, N527, N77);
nor NOR2 (N670, N664, N412);
nor NOR3 (N671, N668, N3, N179);
xor XOR2 (N672, N669, N157);
not NOT1 (N673, N663);
not NOT1 (N674, N661);
not NOT1 (N675, N672);
or OR3 (N676, N670, N301, N480);
not NOT1 (N677, N666);
not NOT1 (N678, N673);
nor NOR3 (N679, N676, N347, N28);
xor XOR2 (N680, N677, N428);
or OR4 (N681, N680, N290, N218, N76);
or OR2 (N682, N659, N575);
buf BUF1 (N683, N650);
not NOT1 (N684, N683);
or OR2 (N685, N642, N248);
or OR3 (N686, N674, N468, N95);
xor XOR2 (N687, N678, N232);
nand NAND4 (N688, N662, N524, N178, N571);
or OR4 (N689, N682, N596, N574, N179);
xor XOR2 (N690, N671, N278);
and AND4 (N691, N686, N435, N226, N375);
not NOT1 (N692, N688);
nor NOR3 (N693, N685, N637, N622);
xor XOR2 (N694, N693, N502);
not NOT1 (N695, N681);
xor XOR2 (N696, N691, N444);
not NOT1 (N697, N679);
nand NAND2 (N698, N692, N117);
buf BUF1 (N699, N695);
not NOT1 (N700, N698);
nand NAND4 (N701, N699, N287, N439, N32);
nand NAND3 (N702, N684, N61, N566);
xor XOR2 (N703, N702, N655);
and AND3 (N704, N703, N96, N305);
not NOT1 (N705, N701);
and AND3 (N706, N690, N213, N576);
or OR3 (N707, N675, N685, N698);
or OR2 (N708, N707, N37);
and AND4 (N709, N687, N90, N686, N361);
or OR3 (N710, N706, N552, N649);
nand NAND3 (N711, N697, N518, N437);
nor NOR4 (N712, N694, N623, N551, N68);
and AND2 (N713, N696, N169);
not NOT1 (N714, N708);
nand NAND4 (N715, N705, N483, N256, N633);
or OR2 (N716, N704, N592);
nand NAND4 (N717, N700, N611, N625, N711);
not NOT1 (N718, N104);
buf BUF1 (N719, N709);
or OR3 (N720, N717, N699, N126);
nor NOR3 (N721, N715, N519, N304);
nor NOR4 (N722, N716, N599, N515, N30);
nor NOR2 (N723, N714, N150);
and AND2 (N724, N721, N470);
and AND2 (N725, N713, N302);
or OR2 (N726, N723, N437);
or OR3 (N727, N724, N74, N407);
nor NOR2 (N728, N725, N123);
and AND3 (N729, N719, N273, N372);
xor XOR2 (N730, N712, N527);
xor XOR2 (N731, N730, N532);
buf BUF1 (N732, N731);
nor NOR2 (N733, N710, N268);
and AND3 (N734, N727, N725, N439);
not NOT1 (N735, N733);
and AND3 (N736, N734, N28, N66);
nand NAND3 (N737, N736, N291, N479);
xor XOR2 (N738, N722, N148);
and AND3 (N739, N729, N13, N347);
or OR3 (N740, N735, N389, N666);
or OR3 (N741, N740, N521, N441);
and AND2 (N742, N718, N487);
not NOT1 (N743, N738);
xor XOR2 (N744, N720, N598);
not NOT1 (N745, N739);
nand NAND3 (N746, N745, N141, N4);
nand NAND4 (N747, N741, N219, N480, N742);
or OR4 (N748, N555, N435, N447, N114);
nand NAND4 (N749, N743, N410, N79, N463);
and AND3 (N750, N689, N733, N734);
nand NAND4 (N751, N726, N708, N59, N712);
or OR4 (N752, N750, N366, N72, N262);
buf BUF1 (N753, N744);
not NOT1 (N754, N737);
buf BUF1 (N755, N732);
not NOT1 (N756, N755);
xor XOR2 (N757, N748, N404);
and AND2 (N758, N753, N199);
nor NOR3 (N759, N752, N681, N624);
not NOT1 (N760, N746);
not NOT1 (N761, N754);
buf BUF1 (N762, N760);
nand NAND3 (N763, N728, N598, N642);
and AND4 (N764, N762, N5, N523, N282);
xor XOR2 (N765, N757, N524);
nor NOR3 (N766, N747, N573, N639);
xor XOR2 (N767, N764, N626);
xor XOR2 (N768, N763, N33);
xor XOR2 (N769, N751, N345);
xor XOR2 (N770, N758, N195);
or OR3 (N771, N765, N99, N268);
and AND4 (N772, N768, N471, N431, N28);
not NOT1 (N773, N761);
buf BUF1 (N774, N759);
or OR4 (N775, N767, N470, N416, N13);
buf BUF1 (N776, N773);
or OR4 (N777, N776, N214, N73, N481);
or OR4 (N778, N774, N409, N719, N113);
not NOT1 (N779, N749);
or OR2 (N780, N778, N492);
nand NAND4 (N781, N756, N747, N58, N574);
or OR2 (N782, N770, N706);
nor NOR3 (N783, N771, N441, N308);
or OR4 (N784, N769, N472, N653, N327);
or OR2 (N785, N782, N132);
nor NOR4 (N786, N779, N648, N361, N82);
nand NAND4 (N787, N777, N163, N504, N123);
nand NAND3 (N788, N781, N512, N690);
or OR4 (N789, N785, N651, N129, N756);
buf BUF1 (N790, N784);
or OR2 (N791, N789, N683);
buf BUF1 (N792, N786);
or OR2 (N793, N766, N316);
and AND4 (N794, N792, N583, N219, N521);
nand NAND4 (N795, N788, N114, N545, N744);
nand NAND2 (N796, N775, N575);
nand NAND4 (N797, N795, N742, N347, N348);
or OR3 (N798, N791, N300, N216);
not NOT1 (N799, N783);
nand NAND3 (N800, N798, N540, N527);
xor XOR2 (N801, N780, N257);
and AND4 (N802, N796, N181, N261, N667);
and AND3 (N803, N790, N272, N750);
not NOT1 (N804, N801);
or OR3 (N805, N800, N394, N320);
buf BUF1 (N806, N805);
and AND2 (N807, N797, N146);
nand NAND4 (N808, N772, N397, N307, N467);
not NOT1 (N809, N799);
xor XOR2 (N810, N807, N681);
and AND2 (N811, N806, N700);
xor XOR2 (N812, N810, N647);
xor XOR2 (N813, N811, N49);
or OR4 (N814, N808, N508, N383, N296);
nand NAND4 (N815, N804, N452, N116, N294);
not NOT1 (N816, N813);
buf BUF1 (N817, N815);
and AND4 (N818, N802, N60, N389, N380);
nand NAND3 (N819, N803, N753, N782);
not NOT1 (N820, N818);
nor NOR3 (N821, N814, N357, N24);
xor XOR2 (N822, N787, N17);
not NOT1 (N823, N819);
nor NOR4 (N824, N812, N506, N421, N14);
and AND4 (N825, N793, N117, N280, N142);
or OR3 (N826, N809, N160, N566);
buf BUF1 (N827, N825);
xor XOR2 (N828, N827, N639);
xor XOR2 (N829, N794, N628);
and AND4 (N830, N821, N618, N636, N512);
nand NAND3 (N831, N823, N547, N536);
nand NAND4 (N832, N829, N512, N413, N401);
and AND2 (N833, N822, N817);
nor NOR4 (N834, N787, N696, N6, N254);
nand NAND3 (N835, N831, N660, N595);
not NOT1 (N836, N824);
not NOT1 (N837, N828);
not NOT1 (N838, N816);
xor XOR2 (N839, N838, N751);
and AND3 (N840, N820, N93, N339);
buf BUF1 (N841, N834);
nor NOR2 (N842, N830, N646);
not NOT1 (N843, N840);
or OR4 (N844, N832, N155, N485, N709);
xor XOR2 (N845, N841, N40);
and AND3 (N846, N845, N709, N587);
xor XOR2 (N847, N837, N539);
xor XOR2 (N848, N826, N30);
or OR2 (N849, N848, N273);
or OR3 (N850, N842, N89, N710);
not NOT1 (N851, N835);
and AND2 (N852, N836, N844);
buf BUF1 (N853, N342);
buf BUF1 (N854, N846);
buf BUF1 (N855, N833);
and AND2 (N856, N847, N684);
buf BUF1 (N857, N850);
and AND4 (N858, N854, N338, N735, N178);
buf BUF1 (N859, N853);
nor NOR4 (N860, N852, N208, N533, N225);
and AND3 (N861, N843, N184, N108);
or OR4 (N862, N856, N384, N29, N818);
nand NAND2 (N863, N860, N230);
not NOT1 (N864, N859);
or OR3 (N865, N849, N377, N309);
and AND3 (N866, N865, N105, N241);
nand NAND4 (N867, N862, N588, N59, N820);
xor XOR2 (N868, N866, N728);
not NOT1 (N869, N867);
nand NAND4 (N870, N863, N587, N40, N634);
not NOT1 (N871, N858);
buf BUF1 (N872, N870);
nor NOR3 (N873, N851, N455, N822);
buf BUF1 (N874, N861);
not NOT1 (N875, N839);
or OR2 (N876, N873, N14);
buf BUF1 (N877, N871);
xor XOR2 (N878, N872, N354);
buf BUF1 (N879, N855);
xor XOR2 (N880, N869, N616);
nor NOR2 (N881, N876, N548);
nor NOR2 (N882, N868, N78);
buf BUF1 (N883, N880);
nor NOR2 (N884, N879, N259);
not NOT1 (N885, N864);
nand NAND2 (N886, N874, N880);
nand NAND3 (N887, N885, N382, N733);
nand NAND4 (N888, N887, N510, N869, N179);
not NOT1 (N889, N882);
xor XOR2 (N890, N888, N449);
xor XOR2 (N891, N886, N890);
nand NAND3 (N892, N762, N3, N451);
or OR3 (N893, N892, N274, N570);
xor XOR2 (N894, N878, N319);
and AND4 (N895, N877, N449, N215, N77);
or OR4 (N896, N875, N398, N650, N321);
buf BUF1 (N897, N893);
not NOT1 (N898, N857);
xor XOR2 (N899, N898, N143);
not NOT1 (N900, N899);
nand NAND3 (N901, N897, N626, N58);
nor NOR2 (N902, N881, N441);
or OR3 (N903, N883, N325, N145);
nor NOR4 (N904, N884, N793, N352, N659);
or OR2 (N905, N896, N521);
xor XOR2 (N906, N902, N269);
xor XOR2 (N907, N905, N717);
nand NAND3 (N908, N900, N14, N733);
buf BUF1 (N909, N904);
xor XOR2 (N910, N895, N454);
nand NAND4 (N911, N894, N9, N400, N718);
buf BUF1 (N912, N901);
xor XOR2 (N913, N891, N484);
xor XOR2 (N914, N909, N264);
not NOT1 (N915, N908);
not NOT1 (N916, N913);
not NOT1 (N917, N915);
buf BUF1 (N918, N906);
and AND3 (N919, N903, N238, N837);
nand NAND3 (N920, N889, N488, N714);
xor XOR2 (N921, N917, N494);
buf BUF1 (N922, N911);
not NOT1 (N923, N920);
xor XOR2 (N924, N921, N751);
nor NOR2 (N925, N910, N35);
not NOT1 (N926, N923);
and AND3 (N927, N907, N503, N317);
xor XOR2 (N928, N925, N210);
xor XOR2 (N929, N919, N215);
nor NOR4 (N930, N916, N789, N385, N747);
xor XOR2 (N931, N927, N362);
nor NOR3 (N932, N922, N622, N318);
or OR4 (N933, N912, N2, N383, N205);
not NOT1 (N934, N933);
and AND4 (N935, N928, N20, N604, N774);
xor XOR2 (N936, N935, N693);
not NOT1 (N937, N931);
buf BUF1 (N938, N926);
not NOT1 (N939, N934);
or OR4 (N940, N929, N229, N216, N241);
xor XOR2 (N941, N914, N671);
nand NAND3 (N942, N941, N530, N307);
not NOT1 (N943, N942);
nand NAND3 (N944, N937, N106, N431);
nor NOR4 (N945, N938, N491, N837, N76);
nand NAND3 (N946, N944, N451, N643);
not NOT1 (N947, N946);
or OR2 (N948, N918, N590);
buf BUF1 (N949, N939);
or OR3 (N950, N945, N501, N806);
nand NAND2 (N951, N947, N339);
or OR3 (N952, N930, N60, N430);
xor XOR2 (N953, N943, N682);
xor XOR2 (N954, N950, N391);
not NOT1 (N955, N949);
buf BUF1 (N956, N953);
xor XOR2 (N957, N948, N311);
nand NAND3 (N958, N954, N883, N406);
nor NOR2 (N959, N924, N674);
or OR4 (N960, N952, N611, N599, N28);
buf BUF1 (N961, N959);
xor XOR2 (N962, N955, N450);
nor NOR2 (N963, N936, N228);
xor XOR2 (N964, N961, N806);
not NOT1 (N965, N960);
nor NOR4 (N966, N965, N607, N346, N157);
and AND3 (N967, N932, N359, N854);
and AND4 (N968, N956, N192, N792, N157);
nand NAND4 (N969, N958, N16, N269, N704);
or OR4 (N970, N969, N18, N961, N278);
nand NAND4 (N971, N964, N569, N846, N799);
and AND4 (N972, N967, N506, N891, N842);
or OR3 (N973, N966, N415, N529);
not NOT1 (N974, N963);
buf BUF1 (N975, N968);
xor XOR2 (N976, N957, N766);
nor NOR2 (N977, N970, N345);
nor NOR4 (N978, N973, N501, N461, N566);
buf BUF1 (N979, N971);
nor NOR2 (N980, N962, N840);
or OR4 (N981, N977, N370, N839, N954);
xor XOR2 (N982, N940, N522);
nor NOR3 (N983, N976, N113, N667);
and AND3 (N984, N972, N185, N574);
or OR4 (N985, N975, N611, N152, N380);
nand NAND4 (N986, N974, N41, N911, N620);
xor XOR2 (N987, N982, N276);
or OR4 (N988, N951, N353, N837, N118);
nor NOR4 (N989, N983, N885, N309, N500);
nor NOR4 (N990, N978, N144, N43, N943);
not NOT1 (N991, N989);
nor NOR3 (N992, N987, N198, N48);
nand NAND2 (N993, N988, N266);
or OR3 (N994, N986, N898, N101);
not NOT1 (N995, N985);
xor XOR2 (N996, N995, N443);
or OR4 (N997, N990, N406, N68, N391);
buf BUF1 (N998, N979);
nor NOR2 (N999, N980, N49);
or OR4 (N1000, N996, N148, N910, N304);
not NOT1 (N1001, N991);
xor XOR2 (N1002, N1001, N928);
or OR3 (N1003, N999, N438, N894);
nand NAND3 (N1004, N994, N778, N869);
nor NOR3 (N1005, N1003, N999, N28);
nand NAND3 (N1006, N1005, N717, N689);
nand NAND2 (N1007, N1002, N674);
or OR4 (N1008, N1006, N937, N700, N346);
nand NAND4 (N1009, N984, N350, N229, N806);
or OR3 (N1010, N992, N426, N746);
nor NOR3 (N1011, N1009, N806, N76);
not NOT1 (N1012, N981);
buf BUF1 (N1013, N1004);
or OR3 (N1014, N1012, N363, N519);
nand NAND2 (N1015, N1010, N908);
nand NAND4 (N1016, N993, N766, N515, N659);
or OR2 (N1017, N1014, N205);
buf BUF1 (N1018, N997);
not NOT1 (N1019, N1000);
xor XOR2 (N1020, N1018, N972);
buf BUF1 (N1021, N1008);
buf BUF1 (N1022, N1019);
not NOT1 (N1023, N1021);
buf BUF1 (N1024, N998);
or OR2 (N1025, N1016, N293);
buf BUF1 (N1026, N1007);
or OR4 (N1027, N1024, N926, N173, N697);
nor NOR4 (N1028, N1017, N823, N867, N791);
or OR4 (N1029, N1011, N40, N314, N201);
buf BUF1 (N1030, N1015);
nor NOR3 (N1031, N1013, N923, N553);
or OR2 (N1032, N1020, N630);
nor NOR2 (N1033, N1023, N224);
nor NOR3 (N1034, N1022, N958, N818);
or OR2 (N1035, N1034, N80);
buf BUF1 (N1036, N1026);
nand NAND4 (N1037, N1036, N5, N573, N256);
or OR4 (N1038, N1028, N1013, N509, N82);
nand NAND3 (N1039, N1027, N830, N804);
nor NOR2 (N1040, N1033, N441);
not NOT1 (N1041, N1030);
nand NAND2 (N1042, N1029, N448);
or OR4 (N1043, N1035, N573, N910, N601);
not NOT1 (N1044, N1043);
not NOT1 (N1045, N1040);
xor XOR2 (N1046, N1038, N688);
and AND4 (N1047, N1025, N381, N9, N474);
xor XOR2 (N1048, N1037, N76);
buf BUF1 (N1049, N1047);
xor XOR2 (N1050, N1045, N151);
buf BUF1 (N1051, N1050);
nor NOR2 (N1052, N1049, N767);
nor NOR2 (N1053, N1042, N351);
not NOT1 (N1054, N1044);
and AND2 (N1055, N1051, N671);
nor NOR4 (N1056, N1039, N782, N608, N188);
not NOT1 (N1057, N1054);
xor XOR2 (N1058, N1052, N465);
not NOT1 (N1059, N1032);
not NOT1 (N1060, N1056);
nand NAND4 (N1061, N1048, N476, N1015, N244);
nor NOR4 (N1062, N1057, N443, N590, N46);
not NOT1 (N1063, N1062);
not NOT1 (N1064, N1055);
xor XOR2 (N1065, N1063, N744);
xor XOR2 (N1066, N1065, N77);
not NOT1 (N1067, N1041);
not NOT1 (N1068, N1067);
or OR3 (N1069, N1064, N484, N391);
nor NOR2 (N1070, N1061, N489);
xor XOR2 (N1071, N1046, N651);
nor NOR2 (N1072, N1031, N546);
or OR4 (N1073, N1060, N861, N1038, N279);
nand NAND3 (N1074, N1068, N204, N695);
and AND3 (N1075, N1073, N524, N497);
or OR4 (N1076, N1070, N997, N67, N962);
nor NOR2 (N1077, N1066, N890);
and AND4 (N1078, N1076, N191, N247, N267);
or OR3 (N1079, N1059, N9, N323);
nand NAND2 (N1080, N1053, N1074);
xor XOR2 (N1081, N369, N615);
xor XOR2 (N1082, N1072, N37);
xor XOR2 (N1083, N1081, N644);
and AND4 (N1084, N1071, N841, N656, N878);
buf BUF1 (N1085, N1058);
and AND3 (N1086, N1083, N753, N958);
buf BUF1 (N1087, N1069);
nor NOR2 (N1088, N1080, N389);
xor XOR2 (N1089, N1084, N462);
nand NAND4 (N1090, N1078, N651, N667, N439);
nor NOR3 (N1091, N1087, N286, N434);
buf BUF1 (N1092, N1089);
and AND3 (N1093, N1090, N650, N800);
xor XOR2 (N1094, N1085, N279);
buf BUF1 (N1095, N1093);
or OR2 (N1096, N1095, N217);
xor XOR2 (N1097, N1079, N363);
buf BUF1 (N1098, N1082);
and AND3 (N1099, N1098, N796, N126);
not NOT1 (N1100, N1077);
nand NAND2 (N1101, N1099, N284);
or OR4 (N1102, N1088, N523, N399, N926);
buf BUF1 (N1103, N1097);
xor XOR2 (N1104, N1096, N266);
buf BUF1 (N1105, N1086);
not NOT1 (N1106, N1105);
buf BUF1 (N1107, N1103);
nor NOR3 (N1108, N1092, N779, N501);
buf BUF1 (N1109, N1107);
and AND4 (N1110, N1094, N189, N460, N420);
xor XOR2 (N1111, N1104, N96);
nand NAND4 (N1112, N1102, N804, N695, N805);
not NOT1 (N1113, N1111);
nand NAND2 (N1114, N1110, N374);
or OR4 (N1115, N1108, N807, N940, N1050);
nand NAND2 (N1116, N1115, N784);
or OR4 (N1117, N1106, N476, N686, N908);
nor NOR3 (N1118, N1117, N368, N1097);
xor XOR2 (N1119, N1091, N899);
not NOT1 (N1120, N1101);
nand NAND4 (N1121, N1109, N232, N250, N459);
buf BUF1 (N1122, N1100);
buf BUF1 (N1123, N1119);
or OR2 (N1124, N1118, N697);
and AND4 (N1125, N1121, N340, N538, N468);
nor NOR2 (N1126, N1124, N297);
not NOT1 (N1127, N1123);
nor NOR4 (N1128, N1114, N538, N1091, N72);
not NOT1 (N1129, N1127);
and AND3 (N1130, N1116, N530, N365);
and AND2 (N1131, N1075, N788);
nand NAND2 (N1132, N1129, N108);
buf BUF1 (N1133, N1130);
nor NOR2 (N1134, N1133, N603);
buf BUF1 (N1135, N1122);
buf BUF1 (N1136, N1134);
nand NAND2 (N1137, N1135, N190);
or OR3 (N1138, N1132, N918, N1128);
and AND3 (N1139, N246, N789, N8);
or OR4 (N1140, N1136, N121, N379, N1021);
not NOT1 (N1141, N1113);
xor XOR2 (N1142, N1125, N134);
buf BUF1 (N1143, N1138);
not NOT1 (N1144, N1112);
nand NAND2 (N1145, N1140, N771);
xor XOR2 (N1146, N1142, N629);
and AND3 (N1147, N1126, N1060, N622);
xor XOR2 (N1148, N1143, N244);
buf BUF1 (N1149, N1139);
and AND2 (N1150, N1148, N1125);
not NOT1 (N1151, N1137);
not NOT1 (N1152, N1141);
nor NOR4 (N1153, N1131, N1139, N954, N680);
and AND4 (N1154, N1120, N614, N350, N393);
or OR3 (N1155, N1149, N544, N789);
nand NAND2 (N1156, N1145, N846);
not NOT1 (N1157, N1150);
xor XOR2 (N1158, N1157, N414);
nand NAND2 (N1159, N1152, N706);
or OR2 (N1160, N1158, N776);
or OR4 (N1161, N1160, N796, N1007, N132);
nor NOR3 (N1162, N1153, N1018, N588);
not NOT1 (N1163, N1151);
and AND4 (N1164, N1162, N613, N956, N501);
nor NOR4 (N1165, N1161, N781, N987, N482);
xor XOR2 (N1166, N1156, N745);
buf BUF1 (N1167, N1165);
nor NOR3 (N1168, N1146, N361, N60);
buf BUF1 (N1169, N1144);
buf BUF1 (N1170, N1154);
buf BUF1 (N1171, N1169);
buf BUF1 (N1172, N1163);
and AND3 (N1173, N1167, N724, N283);
and AND4 (N1174, N1173, N1025, N992, N100);
xor XOR2 (N1175, N1155, N1103);
xor XOR2 (N1176, N1171, N395);
or OR3 (N1177, N1172, N601, N71);
not NOT1 (N1178, N1159);
not NOT1 (N1179, N1170);
or OR4 (N1180, N1175, N858, N1100, N660);
nor NOR3 (N1181, N1178, N627, N506);
not NOT1 (N1182, N1180);
nor NOR2 (N1183, N1166, N786);
not NOT1 (N1184, N1177);
not NOT1 (N1185, N1183);
and AND3 (N1186, N1164, N309, N511);
nand NAND3 (N1187, N1174, N373, N864);
xor XOR2 (N1188, N1179, N221);
xor XOR2 (N1189, N1184, N509);
nand NAND4 (N1190, N1185, N189, N63, N890);
or OR4 (N1191, N1190, N108, N1093, N982);
not NOT1 (N1192, N1191);
nor NOR3 (N1193, N1192, N928, N389);
and AND4 (N1194, N1182, N908, N1105, N2);
or OR3 (N1195, N1181, N810, N626);
nand NAND2 (N1196, N1194, N466);
not NOT1 (N1197, N1147);
not NOT1 (N1198, N1196);
or OR2 (N1199, N1198, N650);
xor XOR2 (N1200, N1199, N342);
nand NAND4 (N1201, N1195, N217, N985, N1192);
xor XOR2 (N1202, N1187, N691);
nand NAND4 (N1203, N1201, N414, N676, N738);
not NOT1 (N1204, N1203);
and AND3 (N1205, N1176, N1154, N1032);
not NOT1 (N1206, N1205);
or OR2 (N1207, N1206, N63);
nand NAND2 (N1208, N1204, N872);
xor XOR2 (N1209, N1197, N541);
or OR2 (N1210, N1188, N1177);
and AND2 (N1211, N1210, N1190);
or OR2 (N1212, N1207, N105);
buf BUF1 (N1213, N1209);
and AND3 (N1214, N1186, N698, N534);
and AND4 (N1215, N1208, N332, N175, N522);
nand NAND3 (N1216, N1211, N899, N480);
not NOT1 (N1217, N1212);
not NOT1 (N1218, N1189);
nand NAND4 (N1219, N1217, N185, N242, N146);
xor XOR2 (N1220, N1216, N1034);
not NOT1 (N1221, N1214);
or OR3 (N1222, N1168, N924, N492);
and AND4 (N1223, N1215, N261, N1195, N1188);
not NOT1 (N1224, N1193);
not NOT1 (N1225, N1213);
or OR4 (N1226, N1219, N225, N360, N738);
and AND3 (N1227, N1223, N960, N174);
nand NAND3 (N1228, N1202, N504, N237);
nor NOR3 (N1229, N1221, N520, N218);
and AND2 (N1230, N1229, N144);
not NOT1 (N1231, N1200);
not NOT1 (N1232, N1231);
nor NOR2 (N1233, N1220, N521);
nand NAND3 (N1234, N1222, N575, N1098);
or OR3 (N1235, N1225, N1055, N908);
nor NOR3 (N1236, N1232, N923, N335);
and AND2 (N1237, N1226, N1012);
nand NAND2 (N1238, N1234, N831);
nand NAND3 (N1239, N1233, N787, N1085);
nor NOR2 (N1240, N1218, N634);
buf BUF1 (N1241, N1230);
buf BUF1 (N1242, N1235);
nor NOR3 (N1243, N1236, N836, N1022);
buf BUF1 (N1244, N1227);
nor NOR3 (N1245, N1243, N688, N331);
not NOT1 (N1246, N1245);
xor XOR2 (N1247, N1238, N156);
buf BUF1 (N1248, N1228);
and AND2 (N1249, N1244, N1019);
or OR2 (N1250, N1242, N548);
buf BUF1 (N1251, N1248);
nand NAND4 (N1252, N1224, N853, N925, N189);
or OR4 (N1253, N1240, N236, N419, N920);
and AND4 (N1254, N1241, N117, N644, N795);
buf BUF1 (N1255, N1251);
and AND3 (N1256, N1247, N763, N988);
or OR4 (N1257, N1239, N82, N1120, N345);
not NOT1 (N1258, N1237);
xor XOR2 (N1259, N1246, N136);
or OR3 (N1260, N1252, N665, N987);
and AND2 (N1261, N1257, N845);
not NOT1 (N1262, N1258);
buf BUF1 (N1263, N1255);
buf BUF1 (N1264, N1259);
buf BUF1 (N1265, N1261);
or OR4 (N1266, N1256, N73, N496, N958);
not NOT1 (N1267, N1264);
buf BUF1 (N1268, N1262);
xor XOR2 (N1269, N1253, N1027);
not NOT1 (N1270, N1263);
nand NAND2 (N1271, N1254, N421);
xor XOR2 (N1272, N1267, N1211);
nand NAND2 (N1273, N1249, N1010);
xor XOR2 (N1274, N1260, N913);
xor XOR2 (N1275, N1265, N793);
buf BUF1 (N1276, N1269);
xor XOR2 (N1277, N1268, N1056);
or OR3 (N1278, N1275, N1076, N492);
or OR4 (N1279, N1276, N448, N206, N338);
not NOT1 (N1280, N1279);
xor XOR2 (N1281, N1272, N147);
nor NOR2 (N1282, N1281, N351);
buf BUF1 (N1283, N1282);
xor XOR2 (N1284, N1266, N543);
or OR3 (N1285, N1250, N870, N943);
nand NAND4 (N1286, N1284, N142, N264, N1158);
xor XOR2 (N1287, N1283, N528);
not NOT1 (N1288, N1280);
or OR2 (N1289, N1277, N54);
nor NOR2 (N1290, N1274, N751);
and AND3 (N1291, N1273, N382, N280);
nand NAND3 (N1292, N1291, N379, N931);
or OR4 (N1293, N1290, N401, N248, N1030);
and AND2 (N1294, N1278, N1213);
not NOT1 (N1295, N1286);
nand NAND3 (N1296, N1289, N1209, N1258);
nand NAND3 (N1297, N1294, N258, N354);
xor XOR2 (N1298, N1295, N1260);
or OR3 (N1299, N1292, N684, N811);
and AND2 (N1300, N1293, N21);
or OR3 (N1301, N1288, N268, N1071);
buf BUF1 (N1302, N1297);
nor NOR2 (N1303, N1302, N484);
nor NOR4 (N1304, N1270, N855, N1168, N250);
xor XOR2 (N1305, N1298, N90);
or OR4 (N1306, N1285, N629, N1146, N1178);
buf BUF1 (N1307, N1306);
xor XOR2 (N1308, N1287, N589);
nand NAND4 (N1309, N1305, N241, N992, N725);
buf BUF1 (N1310, N1301);
nand NAND3 (N1311, N1307, N7, N1073);
and AND2 (N1312, N1311, N1176);
xor XOR2 (N1313, N1299, N759);
or OR4 (N1314, N1304, N823, N39, N563);
nor NOR2 (N1315, N1271, N1297);
not NOT1 (N1316, N1315);
buf BUF1 (N1317, N1313);
or OR3 (N1318, N1317, N1165, N362);
not NOT1 (N1319, N1314);
xor XOR2 (N1320, N1308, N952);
not NOT1 (N1321, N1300);
nor NOR2 (N1322, N1312, N691);
xor XOR2 (N1323, N1321, N720);
and AND3 (N1324, N1320, N690, N1103);
nand NAND3 (N1325, N1310, N612, N360);
not NOT1 (N1326, N1322);
not NOT1 (N1327, N1303);
xor XOR2 (N1328, N1326, N603);
and AND2 (N1329, N1323, N1222);
nand NAND3 (N1330, N1316, N1153, N641);
nor NOR4 (N1331, N1296, N945, N639, N357);
and AND3 (N1332, N1327, N166, N15);
and AND2 (N1333, N1331, N463);
buf BUF1 (N1334, N1309);
buf BUF1 (N1335, N1330);
buf BUF1 (N1336, N1325);
buf BUF1 (N1337, N1328);
not NOT1 (N1338, N1333);
nand NAND4 (N1339, N1318, N880, N843, N1304);
buf BUF1 (N1340, N1335);
not NOT1 (N1341, N1329);
not NOT1 (N1342, N1319);
xor XOR2 (N1343, N1341, N719);
and AND2 (N1344, N1334, N1291);
xor XOR2 (N1345, N1336, N1208);
not NOT1 (N1346, N1344);
not NOT1 (N1347, N1324);
xor XOR2 (N1348, N1342, N745);
not NOT1 (N1349, N1338);
not NOT1 (N1350, N1337);
or OR3 (N1351, N1339, N3, N659);
xor XOR2 (N1352, N1332, N179);
and AND2 (N1353, N1343, N198);
or OR4 (N1354, N1350, N1227, N317, N732);
or OR3 (N1355, N1348, N501, N752);
or OR2 (N1356, N1351, N900);
and AND2 (N1357, N1353, N112);
nor NOR2 (N1358, N1340, N536);
xor XOR2 (N1359, N1356, N1077);
buf BUF1 (N1360, N1354);
nor NOR3 (N1361, N1346, N1088, N171);
or OR2 (N1362, N1355, N865);
nand NAND3 (N1363, N1361, N647, N1045);
and AND3 (N1364, N1362, N955, N1318);
or OR4 (N1365, N1363, N861, N749, N255);
xor XOR2 (N1366, N1359, N822);
buf BUF1 (N1367, N1352);
nand NAND3 (N1368, N1367, N32, N173);
buf BUF1 (N1369, N1368);
nor NOR3 (N1370, N1369, N82, N329);
buf BUF1 (N1371, N1357);
nand NAND4 (N1372, N1358, N773, N350, N537);
xor XOR2 (N1373, N1365, N1319);
nor NOR3 (N1374, N1371, N438, N367);
xor XOR2 (N1375, N1374, N1099);
not NOT1 (N1376, N1372);
xor XOR2 (N1377, N1376, N1081);
xor XOR2 (N1378, N1375, N213);
nand NAND4 (N1379, N1349, N962, N80, N479);
buf BUF1 (N1380, N1347);
buf BUF1 (N1381, N1380);
nor NOR4 (N1382, N1366, N857, N2, N619);
nor NOR2 (N1383, N1360, N1);
xor XOR2 (N1384, N1377, N254);
not NOT1 (N1385, N1381);
or OR4 (N1386, N1383, N15, N339, N1184);
or OR3 (N1387, N1386, N1122, N1018);
xor XOR2 (N1388, N1345, N1110);
nor NOR4 (N1389, N1364, N863, N675, N1293);
nand NAND3 (N1390, N1379, N314, N1288);
nand NAND3 (N1391, N1370, N624, N1087);
nor NOR2 (N1392, N1387, N1068);
not NOT1 (N1393, N1384);
nor NOR4 (N1394, N1390, N153, N125, N1389);
nand NAND3 (N1395, N824, N493, N223);
buf BUF1 (N1396, N1394);
and AND4 (N1397, N1378, N750, N1005, N639);
buf BUF1 (N1398, N1395);
not NOT1 (N1399, N1382);
or OR3 (N1400, N1397, N103, N202);
not NOT1 (N1401, N1396);
buf BUF1 (N1402, N1401);
nor NOR3 (N1403, N1393, N1218, N224);
nor NOR2 (N1404, N1402, N615);
nor NOR3 (N1405, N1400, N285, N817);
not NOT1 (N1406, N1399);
nor NOR3 (N1407, N1388, N835, N305);
nor NOR3 (N1408, N1406, N1116, N1234);
or OR4 (N1409, N1392, N1020, N591, N191);
not NOT1 (N1410, N1409);
nor NOR3 (N1411, N1404, N324, N1290);
not NOT1 (N1412, N1410);
or OR2 (N1413, N1403, N1367);
nor NOR3 (N1414, N1385, N403, N210);
or OR2 (N1415, N1412, N268);
and AND3 (N1416, N1413, N486, N246);
not NOT1 (N1417, N1411);
nand NAND3 (N1418, N1373, N1272, N370);
and AND3 (N1419, N1407, N837, N922);
xor XOR2 (N1420, N1417, N952);
xor XOR2 (N1421, N1416, N357);
and AND3 (N1422, N1408, N808, N78);
nor NOR2 (N1423, N1414, N491);
or OR4 (N1424, N1420, N1231, N1002, N495);
buf BUF1 (N1425, N1391);
not NOT1 (N1426, N1405);
nand NAND4 (N1427, N1398, N998, N789, N52);
or OR2 (N1428, N1424, N1062);
nor NOR3 (N1429, N1418, N980, N745);
not NOT1 (N1430, N1427);
nor NOR4 (N1431, N1430, N1213, N706, N1252);
xor XOR2 (N1432, N1419, N560);
buf BUF1 (N1433, N1429);
nor NOR4 (N1434, N1432, N409, N1058, N1318);
buf BUF1 (N1435, N1425);
buf BUF1 (N1436, N1433);
buf BUF1 (N1437, N1428);
xor XOR2 (N1438, N1423, N803);
and AND3 (N1439, N1426, N522, N724);
xor XOR2 (N1440, N1438, N1029);
nand NAND2 (N1441, N1437, N1185);
xor XOR2 (N1442, N1421, N258);
nand NAND2 (N1443, N1439, N538);
nor NOR4 (N1444, N1440, N607, N122, N853);
not NOT1 (N1445, N1431);
buf BUF1 (N1446, N1435);
xor XOR2 (N1447, N1445, N947);
buf BUF1 (N1448, N1441);
nand NAND3 (N1449, N1444, N106, N850);
xor XOR2 (N1450, N1422, N872);
xor XOR2 (N1451, N1447, N448);
and AND3 (N1452, N1415, N404, N160);
xor XOR2 (N1453, N1450, N1186);
not NOT1 (N1454, N1448);
buf BUF1 (N1455, N1434);
not NOT1 (N1456, N1454);
nor NOR4 (N1457, N1453, N484, N234, N63);
not NOT1 (N1458, N1452);
nand NAND2 (N1459, N1436, N248);
buf BUF1 (N1460, N1443);
xor XOR2 (N1461, N1458, N634);
nand NAND4 (N1462, N1461, N436, N621, N1395);
nand NAND3 (N1463, N1462, N673, N153);
and AND2 (N1464, N1446, N1027);
or OR3 (N1465, N1463, N1346, N501);
and AND2 (N1466, N1465, N406);
nor NOR3 (N1467, N1464, N97, N506);
nand NAND4 (N1468, N1459, N1313, N182, N1063);
xor XOR2 (N1469, N1467, N1161);
not NOT1 (N1470, N1460);
not NOT1 (N1471, N1468);
or OR3 (N1472, N1466, N147, N402);
nand NAND4 (N1473, N1451, N234, N1312, N75);
xor XOR2 (N1474, N1471, N1321);
not NOT1 (N1475, N1457);
xor XOR2 (N1476, N1472, N28);
buf BUF1 (N1477, N1449);
and AND4 (N1478, N1477, N813, N342, N1373);
buf BUF1 (N1479, N1469);
xor XOR2 (N1480, N1475, N1204);
or OR4 (N1481, N1476, N920, N1173, N853);
nand NAND4 (N1482, N1473, N1273, N787, N135);
and AND2 (N1483, N1480, N1123);
nor NOR2 (N1484, N1481, N509);
and AND2 (N1485, N1482, N49);
and AND4 (N1486, N1479, N468, N479, N1358);
buf BUF1 (N1487, N1478);
nand NAND2 (N1488, N1484, N1400);
or OR3 (N1489, N1442, N288, N50);
nand NAND2 (N1490, N1456, N1177);
nor NOR4 (N1491, N1488, N701, N1093, N1069);
buf BUF1 (N1492, N1474);
xor XOR2 (N1493, N1489, N576);
or OR4 (N1494, N1486, N546, N228, N486);
or OR3 (N1495, N1491, N835, N845);
and AND4 (N1496, N1495, N657, N1223, N1165);
and AND3 (N1497, N1496, N605, N1308);
or OR4 (N1498, N1493, N1048, N1184, N503);
buf BUF1 (N1499, N1494);
buf BUF1 (N1500, N1487);
nor NOR4 (N1501, N1455, N1231, N1234, N1252);
nor NOR2 (N1502, N1490, N336);
nor NOR3 (N1503, N1483, N1031, N1080);
nor NOR4 (N1504, N1500, N534, N830, N54);
or OR2 (N1505, N1504, N1331);
nand NAND4 (N1506, N1503, N717, N397, N82);
xor XOR2 (N1507, N1470, N568);
nor NOR4 (N1508, N1499, N1435, N162, N1487);
nor NOR4 (N1509, N1498, N1062, N1470, N996);
nor NOR2 (N1510, N1508, N763);
xor XOR2 (N1511, N1507, N1504);
not NOT1 (N1512, N1497);
and AND2 (N1513, N1506, N692);
and AND4 (N1514, N1510, N90, N668, N733);
not NOT1 (N1515, N1492);
nand NAND3 (N1516, N1513, N59, N1094);
nor NOR3 (N1517, N1502, N1104, N734);
or OR2 (N1518, N1512, N1047);
buf BUF1 (N1519, N1501);
buf BUF1 (N1520, N1517);
buf BUF1 (N1521, N1516);
and AND4 (N1522, N1515, N1437, N1409, N1016);
nor NOR4 (N1523, N1511, N862, N176, N256);
not NOT1 (N1524, N1520);
nand NAND3 (N1525, N1521, N306, N755);
and AND4 (N1526, N1523, N959, N438, N1329);
buf BUF1 (N1527, N1514);
and AND4 (N1528, N1527, N82, N650, N1065);
or OR4 (N1529, N1509, N1040, N1140, N1235);
xor XOR2 (N1530, N1485, N330);
not NOT1 (N1531, N1530);
buf BUF1 (N1532, N1531);
nor NOR3 (N1533, N1522, N147, N344);
not NOT1 (N1534, N1519);
nand NAND4 (N1535, N1505, N1015, N301, N428);
nand NAND2 (N1536, N1529, N429);
nor NOR2 (N1537, N1526, N829);
xor XOR2 (N1538, N1536, N85);
not NOT1 (N1539, N1538);
nand NAND3 (N1540, N1524, N1283, N1308);
or OR4 (N1541, N1535, N1002, N621, N165);
not NOT1 (N1542, N1532);
not NOT1 (N1543, N1540);
and AND4 (N1544, N1542, N342, N1276, N712);
xor XOR2 (N1545, N1534, N928);
nand NAND4 (N1546, N1541, N140, N980, N661);
or OR4 (N1547, N1539, N585, N1374, N781);
buf BUF1 (N1548, N1528);
and AND4 (N1549, N1533, N1454, N1327, N247);
nand NAND3 (N1550, N1543, N1008, N621);
nand NAND4 (N1551, N1547, N858, N739, N321);
buf BUF1 (N1552, N1551);
not NOT1 (N1553, N1548);
nor NOR2 (N1554, N1545, N134);
not NOT1 (N1555, N1546);
and AND2 (N1556, N1544, N785);
or OR3 (N1557, N1549, N1223, N463);
and AND4 (N1558, N1553, N1238, N1318, N223);
and AND2 (N1559, N1554, N1276);
nand NAND3 (N1560, N1559, N99, N483);
buf BUF1 (N1561, N1518);
or OR2 (N1562, N1537, N1407);
nor NOR2 (N1563, N1558, N1530);
nand NAND3 (N1564, N1560, N1341, N80);
nand NAND3 (N1565, N1557, N866, N45);
nor NOR3 (N1566, N1550, N576, N904);
or OR4 (N1567, N1552, N860, N514, N160);
and AND2 (N1568, N1556, N1341);
buf BUF1 (N1569, N1563);
xor XOR2 (N1570, N1568, N943);
nor NOR2 (N1571, N1565, N469);
xor XOR2 (N1572, N1555, N1033);
buf BUF1 (N1573, N1525);
xor XOR2 (N1574, N1571, N508);
xor XOR2 (N1575, N1566, N1464);
and AND4 (N1576, N1562, N44, N640, N133);
buf BUF1 (N1577, N1564);
nor NOR2 (N1578, N1576, N1430);
buf BUF1 (N1579, N1570);
buf BUF1 (N1580, N1567);
nor NOR4 (N1581, N1574, N272, N1134, N987);
nand NAND4 (N1582, N1580, N715, N44, N385);
and AND4 (N1583, N1572, N281, N39, N923);
or OR4 (N1584, N1573, N1541, N276, N503);
nand NAND4 (N1585, N1581, N979, N384, N790);
xor XOR2 (N1586, N1583, N1282);
buf BUF1 (N1587, N1582);
and AND4 (N1588, N1579, N1500, N1542, N406);
and AND4 (N1589, N1584, N420, N187, N610);
or OR2 (N1590, N1588, N25);
nand NAND2 (N1591, N1590, N476);
nor NOR4 (N1592, N1578, N399, N284, N748);
or OR4 (N1593, N1575, N828, N1584, N293);
nand NAND4 (N1594, N1589, N523, N1301, N1267);
or OR2 (N1595, N1592, N519);
nor NOR4 (N1596, N1577, N185, N702, N370);
xor XOR2 (N1597, N1561, N534);
not NOT1 (N1598, N1595);
xor XOR2 (N1599, N1585, N185);
and AND4 (N1600, N1594, N755, N350, N1217);
buf BUF1 (N1601, N1591);
buf BUF1 (N1602, N1569);
and AND2 (N1603, N1600, N165);
xor XOR2 (N1604, N1603, N40);
nand NAND4 (N1605, N1587, N129, N306, N1379);
or OR4 (N1606, N1596, N416, N874, N816);
nand NAND2 (N1607, N1602, N171);
nor NOR2 (N1608, N1586, N846);
and AND4 (N1609, N1597, N276, N1044, N1471);
buf BUF1 (N1610, N1601);
nand NAND4 (N1611, N1604, N1602, N919, N792);
xor XOR2 (N1612, N1611, N543);
and AND2 (N1613, N1612, N20);
and AND3 (N1614, N1609, N684, N942);
or OR2 (N1615, N1605, N1193);
not NOT1 (N1616, N1607);
buf BUF1 (N1617, N1610);
nand NAND2 (N1618, N1613, N266);
and AND4 (N1619, N1606, N1163, N1252, N902);
nor NOR2 (N1620, N1599, N1426);
or OR2 (N1621, N1619, N667);
or OR3 (N1622, N1615, N196, N1500);
not NOT1 (N1623, N1593);
xor XOR2 (N1624, N1618, N457);
xor XOR2 (N1625, N1622, N1325);
nor NOR4 (N1626, N1617, N410, N737, N951);
and AND4 (N1627, N1624, N162, N28, N910);
nand NAND2 (N1628, N1608, N96);
nand NAND2 (N1629, N1616, N1045);
or OR4 (N1630, N1628, N409, N193, N34);
not NOT1 (N1631, N1614);
or OR2 (N1632, N1598, N337);
or OR3 (N1633, N1627, N1027, N1094);
buf BUF1 (N1634, N1629);
buf BUF1 (N1635, N1626);
and AND3 (N1636, N1631, N1051, N1334);
nand NAND2 (N1637, N1632, N1074);
or OR2 (N1638, N1625, N221);
and AND4 (N1639, N1621, N971, N1437, N1539);
or OR3 (N1640, N1639, N176, N1468);
nand NAND2 (N1641, N1634, N546);
nand NAND3 (N1642, N1640, N1598, N285);
buf BUF1 (N1643, N1638);
and AND2 (N1644, N1636, N884);
or OR2 (N1645, N1635, N578);
not NOT1 (N1646, N1642);
xor XOR2 (N1647, N1644, N87);
or OR4 (N1648, N1641, N879, N1292, N176);
nand NAND3 (N1649, N1646, N1399, N1486);
nor NOR4 (N1650, N1637, N734, N1107, N474);
or OR2 (N1651, N1647, N256);
buf BUF1 (N1652, N1645);
and AND3 (N1653, N1643, N1318, N472);
buf BUF1 (N1654, N1633);
or OR4 (N1655, N1652, N601, N148, N212);
xor XOR2 (N1656, N1620, N1255);
not NOT1 (N1657, N1630);
not NOT1 (N1658, N1648);
nor NOR3 (N1659, N1623, N119, N304);
nand NAND4 (N1660, N1650, N17, N612, N371);
nor NOR2 (N1661, N1651, N1350);
not NOT1 (N1662, N1649);
or OR3 (N1663, N1658, N1097, N1536);
not NOT1 (N1664, N1655);
nand NAND3 (N1665, N1663, N1341, N1614);
nand NAND3 (N1666, N1653, N1526, N287);
nand NAND2 (N1667, N1661, N49);
buf BUF1 (N1668, N1657);
and AND2 (N1669, N1656, N1409);
nor NOR4 (N1670, N1665, N1153, N1597, N1061);
xor XOR2 (N1671, N1660, N278);
and AND4 (N1672, N1668, N1509, N820, N507);
nand NAND3 (N1673, N1669, N690, N690);
not NOT1 (N1674, N1672);
not NOT1 (N1675, N1673);
not NOT1 (N1676, N1667);
xor XOR2 (N1677, N1664, N1007);
nor NOR2 (N1678, N1666, N669);
not NOT1 (N1679, N1659);
nor NOR4 (N1680, N1678, N1591, N1141, N1105);
nor NOR4 (N1681, N1677, N1246, N1123, N341);
buf BUF1 (N1682, N1671);
buf BUF1 (N1683, N1654);
xor XOR2 (N1684, N1683, N367);
not NOT1 (N1685, N1674);
and AND2 (N1686, N1670, N449);
nor NOR4 (N1687, N1686, N724, N1126, N626);
nand NAND3 (N1688, N1684, N1371, N680);
nand NAND3 (N1689, N1682, N1149, N878);
or OR4 (N1690, N1681, N1099, N1077, N451);
nand NAND4 (N1691, N1662, N63, N865, N151);
and AND3 (N1692, N1688, N768, N115);
and AND2 (N1693, N1691, N184);
nand NAND2 (N1694, N1687, N1580);
and AND4 (N1695, N1693, N971, N1592, N1692);
nor NOR3 (N1696, N484, N1185, N859);
xor XOR2 (N1697, N1679, N1536);
not NOT1 (N1698, N1690);
xor XOR2 (N1699, N1695, N1198);
and AND2 (N1700, N1676, N1428);
nor NOR2 (N1701, N1697, N1093);
xor XOR2 (N1702, N1698, N1093);
xor XOR2 (N1703, N1702, N1160);
and AND3 (N1704, N1700, N40, N1511);
buf BUF1 (N1705, N1680);
nand NAND2 (N1706, N1701, N396);
nor NOR3 (N1707, N1704, N386, N864);
xor XOR2 (N1708, N1696, N709);
buf BUF1 (N1709, N1699);
buf BUF1 (N1710, N1703);
xor XOR2 (N1711, N1708, N768);
xor XOR2 (N1712, N1706, N449);
not NOT1 (N1713, N1685);
xor XOR2 (N1714, N1713, N306);
nand NAND2 (N1715, N1694, N1223);
xor XOR2 (N1716, N1707, N717);
and AND2 (N1717, N1675, N1491);
nand NAND4 (N1718, N1705, N1545, N520, N754);
nor NOR2 (N1719, N1717, N1409);
buf BUF1 (N1720, N1715);
nor NOR2 (N1721, N1718, N1123);
not NOT1 (N1722, N1712);
or OR2 (N1723, N1710, N135);
or OR3 (N1724, N1721, N23, N491);
and AND4 (N1725, N1720, N1531, N79, N1119);
nand NAND4 (N1726, N1714, N579, N1122, N633);
xor XOR2 (N1727, N1722, N718);
nand NAND3 (N1728, N1716, N486, N1286);
or OR2 (N1729, N1711, N732);
nor NOR2 (N1730, N1728, N1663);
xor XOR2 (N1731, N1729, N112);
or OR2 (N1732, N1689, N83);
and AND2 (N1733, N1730, N975);
buf BUF1 (N1734, N1733);
not NOT1 (N1735, N1725);
nor NOR3 (N1736, N1727, N1343, N551);
or OR4 (N1737, N1719, N1374, N210, N1670);
not NOT1 (N1738, N1737);
nand NAND3 (N1739, N1738, N4, N374);
not NOT1 (N1740, N1739);
and AND3 (N1741, N1723, N653, N797);
nor NOR4 (N1742, N1735, N701, N583, N679);
nand NAND3 (N1743, N1731, N120, N1504);
or OR3 (N1744, N1743, N1676, N1710);
not NOT1 (N1745, N1742);
xor XOR2 (N1746, N1736, N223);
or OR4 (N1747, N1741, N894, N196, N963);
not NOT1 (N1748, N1746);
and AND4 (N1749, N1724, N514, N1145, N1203);
xor XOR2 (N1750, N1726, N831);
buf BUF1 (N1751, N1747);
and AND4 (N1752, N1709, N749, N1556, N118);
buf BUF1 (N1753, N1750);
or OR3 (N1754, N1732, N891, N1590);
nor NOR2 (N1755, N1753, N1468);
xor XOR2 (N1756, N1744, N1211);
nor NOR2 (N1757, N1756, N1737);
or OR2 (N1758, N1749, N825);
or OR2 (N1759, N1745, N779);
not NOT1 (N1760, N1759);
buf BUF1 (N1761, N1754);
and AND2 (N1762, N1755, N330);
not NOT1 (N1763, N1760);
or OR3 (N1764, N1757, N372, N655);
or OR3 (N1765, N1734, N1125, N171);
xor XOR2 (N1766, N1748, N544);
nor NOR2 (N1767, N1751, N726);
nand NAND3 (N1768, N1765, N1055, N1175);
xor XOR2 (N1769, N1758, N381);
and AND4 (N1770, N1766, N52, N163, N1069);
and AND2 (N1771, N1769, N774);
buf BUF1 (N1772, N1752);
nor NOR2 (N1773, N1770, N424);
and AND4 (N1774, N1761, N826, N206, N69);
and AND4 (N1775, N1763, N1406, N1170, N910);
or OR2 (N1776, N1774, N73);
nor NOR2 (N1777, N1740, N689);
nor NOR2 (N1778, N1764, N583);
or OR2 (N1779, N1768, N702);
nor NOR4 (N1780, N1778, N266, N260, N385);
buf BUF1 (N1781, N1780);
nor NOR2 (N1782, N1779, N783);
and AND2 (N1783, N1776, N1692);
nand NAND4 (N1784, N1773, N716, N149, N1395);
nand NAND3 (N1785, N1783, N502, N741);
not NOT1 (N1786, N1781);
xor XOR2 (N1787, N1775, N311);
nor NOR2 (N1788, N1777, N574);
buf BUF1 (N1789, N1772);
buf BUF1 (N1790, N1785);
nand NAND2 (N1791, N1789, N943);
nor NOR4 (N1792, N1762, N49, N1098, N1507);
not NOT1 (N1793, N1771);
and AND2 (N1794, N1792, N846);
not NOT1 (N1795, N1791);
or OR3 (N1796, N1794, N283, N735);
and AND4 (N1797, N1786, N249, N558, N460);
buf BUF1 (N1798, N1788);
xor XOR2 (N1799, N1767, N235);
nor NOR4 (N1800, N1799, N109, N1327, N147);
and AND3 (N1801, N1784, N1106, N476);
xor XOR2 (N1802, N1798, N1056);
nand NAND2 (N1803, N1801, N1024);
and AND4 (N1804, N1795, N1496, N1196, N1010);
xor XOR2 (N1805, N1797, N371);
buf BUF1 (N1806, N1800);
xor XOR2 (N1807, N1790, N810);
buf BUF1 (N1808, N1787);
and AND2 (N1809, N1805, N120);
nor NOR4 (N1810, N1782, N936, N974, N937);
or OR4 (N1811, N1802, N1046, N491, N1030);
or OR4 (N1812, N1809, N1294, N366, N144);
and AND2 (N1813, N1804, N492);
xor XOR2 (N1814, N1803, N808);
nor NOR2 (N1815, N1793, N405);
xor XOR2 (N1816, N1813, N1651);
buf BUF1 (N1817, N1815);
nor NOR4 (N1818, N1796, N347, N240, N155);
nor NOR3 (N1819, N1817, N1508, N112);
not NOT1 (N1820, N1818);
not NOT1 (N1821, N1812);
xor XOR2 (N1822, N1821, N1489);
or OR2 (N1823, N1806, N412);
nand NAND4 (N1824, N1823, N1220, N884, N1108);
nand NAND4 (N1825, N1814, N1184, N89, N1074);
not NOT1 (N1826, N1808);
not NOT1 (N1827, N1826);
buf BUF1 (N1828, N1807);
not NOT1 (N1829, N1820);
xor XOR2 (N1830, N1824, N1741);
not NOT1 (N1831, N1828);
not NOT1 (N1832, N1831);
nor NOR3 (N1833, N1830, N1306, N1181);
not NOT1 (N1834, N1819);
or OR4 (N1835, N1822, N1237, N1768, N907);
not NOT1 (N1836, N1811);
nand NAND4 (N1837, N1816, N558, N991, N467);
nor NOR3 (N1838, N1827, N1478, N1571);
buf BUF1 (N1839, N1810);
nor NOR2 (N1840, N1833, N842);
or OR4 (N1841, N1838, N1767, N1090, N773);
nor NOR3 (N1842, N1835, N1376, N1226);
or OR2 (N1843, N1836, N1205);
nand NAND3 (N1844, N1837, N680, N1555);
nand NAND3 (N1845, N1839, N1790, N1289);
nor NOR2 (N1846, N1834, N398);
and AND4 (N1847, N1844, N583, N381, N1185);
xor XOR2 (N1848, N1845, N717);
nor NOR4 (N1849, N1829, N1764, N596, N824);
nor NOR2 (N1850, N1841, N1561);
nor NOR4 (N1851, N1843, N1761, N1829, N1186);
nand NAND3 (N1852, N1848, N1455, N74);
xor XOR2 (N1853, N1842, N1453);
xor XOR2 (N1854, N1847, N756);
or OR2 (N1855, N1852, N1606);
nand NAND2 (N1856, N1854, N231);
or OR3 (N1857, N1849, N383, N819);
nor NOR2 (N1858, N1857, N631);
and AND2 (N1859, N1858, N23);
nor NOR2 (N1860, N1855, N1630);
nor NOR2 (N1861, N1825, N1532);
and AND4 (N1862, N1856, N66, N1430, N784);
and AND3 (N1863, N1859, N225, N397);
or OR3 (N1864, N1840, N315, N430);
and AND4 (N1865, N1846, N880, N1303, N1484);
not NOT1 (N1866, N1863);
nor NOR2 (N1867, N1860, N363);
xor XOR2 (N1868, N1861, N1097);
buf BUF1 (N1869, N1866);
not NOT1 (N1870, N1853);
nand NAND4 (N1871, N1851, N85, N1451, N1840);
nand NAND3 (N1872, N1871, N1283, N1579);
not NOT1 (N1873, N1864);
xor XOR2 (N1874, N1850, N187);
and AND4 (N1875, N1832, N1292, N381, N808);
nand NAND4 (N1876, N1868, N108, N373, N317);
and AND4 (N1877, N1862, N954, N846, N1622);
nor NOR3 (N1878, N1867, N244, N1711);
and AND3 (N1879, N1872, N423, N411);
or OR2 (N1880, N1873, N1639);
not NOT1 (N1881, N1879);
buf BUF1 (N1882, N1869);
and AND3 (N1883, N1878, N616, N1334);
xor XOR2 (N1884, N1880, N695);
nor NOR3 (N1885, N1865, N594, N156);
xor XOR2 (N1886, N1884, N603);
buf BUF1 (N1887, N1883);
not NOT1 (N1888, N1877);
and AND3 (N1889, N1870, N1322, N1081);
nor NOR2 (N1890, N1886, N1591);
buf BUF1 (N1891, N1881);
not NOT1 (N1892, N1882);
nor NOR3 (N1893, N1889, N957, N1494);
and AND4 (N1894, N1890, N614, N1810, N426);
or OR3 (N1895, N1874, N620, N505);
not NOT1 (N1896, N1875);
xor XOR2 (N1897, N1876, N179);
and AND2 (N1898, N1896, N925);
nand NAND2 (N1899, N1898, N58);
nand NAND2 (N1900, N1885, N1170);
not NOT1 (N1901, N1899);
xor XOR2 (N1902, N1893, N22);
xor XOR2 (N1903, N1897, N866);
buf BUF1 (N1904, N1903);
or OR2 (N1905, N1887, N1898);
nand NAND2 (N1906, N1905, N73);
xor XOR2 (N1907, N1894, N568);
not NOT1 (N1908, N1895);
buf BUF1 (N1909, N1888);
nand NAND2 (N1910, N1908, N1457);
nor NOR4 (N1911, N1906, N86, N1751, N613);
buf BUF1 (N1912, N1911);
nand NAND3 (N1913, N1901, N1051, N101);
or OR2 (N1914, N1907, N1016);
nand NAND2 (N1915, N1904, N192);
and AND4 (N1916, N1912, N1309, N1004, N789);
xor XOR2 (N1917, N1913, N1841);
and AND2 (N1918, N1914, N1708);
nand NAND3 (N1919, N1902, N1547, N961);
buf BUF1 (N1920, N1900);
and AND2 (N1921, N1917, N625);
or OR2 (N1922, N1920, N569);
buf BUF1 (N1923, N1915);
buf BUF1 (N1924, N1921);
nand NAND4 (N1925, N1891, N967, N1780, N1236);
not NOT1 (N1926, N1924);
and AND4 (N1927, N1926, N860, N1056, N1608);
and AND4 (N1928, N1892, N1314, N1329, N328);
or OR3 (N1929, N1909, N320, N1901);
nor NOR3 (N1930, N1919, N285, N1693);
xor XOR2 (N1931, N1922, N1530);
and AND3 (N1932, N1930, N1598, N163);
not NOT1 (N1933, N1910);
buf BUF1 (N1934, N1916);
xor XOR2 (N1935, N1934, N44);
and AND4 (N1936, N1918, N1294, N924, N694);
nand NAND4 (N1937, N1927, N1927, N897, N1441);
nor NOR4 (N1938, N1929, N1638, N1013, N597);
xor XOR2 (N1939, N1935, N1272);
xor XOR2 (N1940, N1932, N1696);
or OR3 (N1941, N1925, N1520, N941);
or OR3 (N1942, N1938, N1232, N822);
not NOT1 (N1943, N1931);
buf BUF1 (N1944, N1939);
xor XOR2 (N1945, N1940, N1941);
or OR3 (N1946, N367, N51, N995);
xor XOR2 (N1947, N1928, N319);
nor NOR3 (N1948, N1943, N1633, N392);
and AND2 (N1949, N1947, N325);
not NOT1 (N1950, N1923);
and AND4 (N1951, N1936, N1011, N1885, N296);
or OR4 (N1952, N1944, N1571, N653, N237);
and AND2 (N1953, N1942, N1601);
buf BUF1 (N1954, N1952);
nand NAND4 (N1955, N1950, N721, N581, N1651);
xor XOR2 (N1956, N1933, N1846);
xor XOR2 (N1957, N1937, N638);
nor NOR2 (N1958, N1955, N1173);
and AND3 (N1959, N1957, N767, N223);
not NOT1 (N1960, N1958);
nand NAND4 (N1961, N1951, N193, N1750, N1563);
or OR3 (N1962, N1960, N1350, N437);
xor XOR2 (N1963, N1949, N243);
xor XOR2 (N1964, N1953, N129);
xor XOR2 (N1965, N1945, N754);
and AND3 (N1966, N1948, N1224, N1566);
nand NAND2 (N1967, N1962, N386);
nand NAND3 (N1968, N1954, N1526, N145);
buf BUF1 (N1969, N1961);
nor NOR2 (N1970, N1946, N92);
xor XOR2 (N1971, N1964, N1153);
nand NAND4 (N1972, N1970, N1128, N1212, N1880);
buf BUF1 (N1973, N1966);
xor XOR2 (N1974, N1959, N775);
and AND2 (N1975, N1972, N1551);
and AND2 (N1976, N1974, N1396);
xor XOR2 (N1977, N1969, N1947);
nor NOR4 (N1978, N1975, N31, N513, N306);
nand NAND2 (N1979, N1965, N75);
nor NOR3 (N1980, N1977, N1337, N1864);
not NOT1 (N1981, N1976);
not NOT1 (N1982, N1963);
and AND3 (N1983, N1967, N1748, N617);
and AND3 (N1984, N1982, N1900, N1147);
nor NOR3 (N1985, N1978, N931, N1387);
nand NAND3 (N1986, N1968, N1363, N797);
and AND3 (N1987, N1980, N830, N1736);
xor XOR2 (N1988, N1981, N707);
not NOT1 (N1989, N1984);
buf BUF1 (N1990, N1971);
buf BUF1 (N1991, N1988);
xor XOR2 (N1992, N1973, N973);
and AND4 (N1993, N1983, N1684, N656, N489);
buf BUF1 (N1994, N1992);
or OR3 (N1995, N1979, N1860, N159);
or OR2 (N1996, N1986, N1717);
buf BUF1 (N1997, N1994);
and AND3 (N1998, N1993, N1665, N422);
nand NAND3 (N1999, N1995, N11, N1405);
buf BUF1 (N2000, N1991);
nor NOR4 (N2001, N1998, N266, N1641, N240);
xor XOR2 (N2002, N1987, N674);
or OR2 (N2003, N1990, N1532);
nand NAND2 (N2004, N2000, N457);
xor XOR2 (N2005, N1956, N1524);
nor NOR4 (N2006, N2004, N761, N1688, N219);
and AND3 (N2007, N2001, N114, N1074);
and AND4 (N2008, N2007, N1759, N46, N819);
not NOT1 (N2009, N1985);
or OR2 (N2010, N1999, N1756);
nand NAND2 (N2011, N1997, N1628);
nand NAND2 (N2012, N2003, N1387);
nor NOR2 (N2013, N1996, N1347);
or OR3 (N2014, N2013, N1503, N175);
nor NOR2 (N2015, N2011, N1155);
not NOT1 (N2016, N2015);
buf BUF1 (N2017, N2012);
and AND4 (N2018, N2005, N828, N1690, N1594);
or OR3 (N2019, N2009, N435, N1611);
and AND4 (N2020, N2010, N486, N1207, N1365);
or OR4 (N2021, N2008, N372, N1133, N1874);
buf BUF1 (N2022, N2018);
buf BUF1 (N2023, N2019);
xor XOR2 (N2024, N2016, N1201);
xor XOR2 (N2025, N2023, N1094);
or OR4 (N2026, N2002, N1474, N1048, N1002);
xor XOR2 (N2027, N2006, N1889);
xor XOR2 (N2028, N2020, N1208);
nor NOR4 (N2029, N2024, N1784, N529, N1019);
buf BUF1 (N2030, N1989);
xor XOR2 (N2031, N2014, N826);
buf BUF1 (N2032, N2025);
xor XOR2 (N2033, N2027, N120);
or OR3 (N2034, N2028, N340, N101);
nand NAND4 (N2035, N2029, N1426, N1738, N1801);
xor XOR2 (N2036, N2022, N44);
and AND3 (N2037, N2026, N1473, N44);
buf BUF1 (N2038, N2034);
or OR2 (N2039, N2030, N562);
nand NAND2 (N2040, N2032, N178);
buf BUF1 (N2041, N2031);
and AND3 (N2042, N2039, N1284, N1810);
xor XOR2 (N2043, N2021, N138);
xor XOR2 (N2044, N2038, N1745);
and AND4 (N2045, N2044, N2020, N168, N362);
and AND2 (N2046, N2045, N291);
and AND2 (N2047, N2033, N135);
not NOT1 (N2048, N2043);
xor XOR2 (N2049, N2036, N1337);
and AND3 (N2050, N2046, N551, N891);
nor NOR2 (N2051, N2048, N880);
buf BUF1 (N2052, N2042);
nor NOR2 (N2053, N2037, N1445);
nand NAND2 (N2054, N2049, N1309);
and AND3 (N2055, N2050, N1414, N1922);
and AND3 (N2056, N2035, N1126, N1504);
nand NAND2 (N2057, N2053, N1207);
nand NAND4 (N2058, N2051, N244, N733, N1624);
not NOT1 (N2059, N2052);
or OR4 (N2060, N2054, N248, N413, N196);
not NOT1 (N2061, N2017);
xor XOR2 (N2062, N2061, N698);
nand NAND4 (N2063, N2058, N1825, N1664, N1022);
or OR4 (N2064, N2057, N337, N150, N267);
and AND3 (N2065, N2059, N410, N1368);
buf BUF1 (N2066, N2041);
nor NOR4 (N2067, N2065, N475, N1450, N961);
and AND4 (N2068, N2056, N964, N90, N761);
nand NAND4 (N2069, N2066, N1359, N1679, N1322);
or OR3 (N2070, N2047, N1392, N874);
buf BUF1 (N2071, N2063);
xor XOR2 (N2072, N2071, N2010);
xor XOR2 (N2073, N2055, N620);
nand NAND3 (N2074, N2067, N938, N863);
buf BUF1 (N2075, N2062);
not NOT1 (N2076, N2075);
not NOT1 (N2077, N2074);
and AND3 (N2078, N2068, N1782, N1342);
xor XOR2 (N2079, N2040, N1269);
or OR3 (N2080, N2073, N142, N925);
nor NOR4 (N2081, N2078, N94, N1752, N673);
and AND2 (N2082, N2077, N767);
buf BUF1 (N2083, N2076);
and AND2 (N2084, N2069, N1877);
and AND2 (N2085, N2083, N2030);
not NOT1 (N2086, N2080);
nand NAND2 (N2087, N2081, N1775);
not NOT1 (N2088, N2079);
nand NAND2 (N2089, N2060, N1000);
nor NOR2 (N2090, N2085, N1220);
nor NOR4 (N2091, N2087, N1182, N1463, N500);
xor XOR2 (N2092, N2091, N1938);
nor NOR3 (N2093, N2082, N150, N1771);
buf BUF1 (N2094, N2072);
nor NOR2 (N2095, N2086, N157);
and AND2 (N2096, N2089, N811);
buf BUF1 (N2097, N2090);
and AND3 (N2098, N2094, N1796, N228);
not NOT1 (N2099, N2097);
nor NOR3 (N2100, N2088, N1202, N1336);
not NOT1 (N2101, N2092);
buf BUF1 (N2102, N2096);
xor XOR2 (N2103, N2095, N570);
nand NAND4 (N2104, N2093, N1446, N2080, N1478);
buf BUF1 (N2105, N2099);
buf BUF1 (N2106, N2105);
nand NAND2 (N2107, N2101, N529);
nor NOR4 (N2108, N2107, N1211, N97, N2043);
and AND4 (N2109, N2104, N437, N1599, N768);
nor NOR2 (N2110, N2109, N1603);
nor NOR4 (N2111, N2070, N1543, N1575, N1116);
nor NOR3 (N2112, N2106, N1797, N162);
nand NAND4 (N2113, N2108, N1269, N1953, N266);
not NOT1 (N2114, N2113);
and AND2 (N2115, N2064, N1582);
nor NOR3 (N2116, N2115, N806, N771);
xor XOR2 (N2117, N2084, N1876);
not NOT1 (N2118, N2100);
not NOT1 (N2119, N2114);
buf BUF1 (N2120, N2111);
nor NOR4 (N2121, N2116, N1004, N776, N788);
or OR3 (N2122, N2098, N1652, N1299);
or OR2 (N2123, N2103, N158);
nor NOR3 (N2124, N2112, N1235, N627);
or OR3 (N2125, N2110, N583, N1844);
buf BUF1 (N2126, N2102);
or OR3 (N2127, N2122, N1703, N1447);
nor NOR3 (N2128, N2119, N1692, N174);
nor NOR3 (N2129, N2127, N292, N202);
xor XOR2 (N2130, N2125, N608);
and AND4 (N2131, N2117, N848, N888, N3);
or OR2 (N2132, N2131, N197);
xor XOR2 (N2133, N2126, N2035);
buf BUF1 (N2134, N2130);
nand NAND4 (N2135, N2120, N458, N1358, N1120);
and AND3 (N2136, N2129, N71, N1142);
or OR2 (N2137, N2128, N501);
not NOT1 (N2138, N2134);
nand NAND2 (N2139, N2123, N1915);
buf BUF1 (N2140, N2121);
nor NOR4 (N2141, N2139, N62, N1714, N1567);
and AND3 (N2142, N2141, N894, N511);
nor NOR3 (N2143, N2136, N1067, N1676);
and AND2 (N2144, N2138, N1503);
nor NOR3 (N2145, N2142, N861, N878);
not NOT1 (N2146, N2145);
not NOT1 (N2147, N2146);
not NOT1 (N2148, N2147);
and AND4 (N2149, N2135, N1651, N1525, N1277);
nor NOR2 (N2150, N2143, N47);
or OR2 (N2151, N2140, N366);
nor NOR2 (N2152, N2144, N797);
xor XOR2 (N2153, N2132, N1968);
xor XOR2 (N2154, N2149, N2022);
nor NOR3 (N2155, N2124, N981, N605);
buf BUF1 (N2156, N2118);
and AND4 (N2157, N2156, N1376, N867, N1381);
and AND2 (N2158, N2152, N564);
or OR3 (N2159, N2154, N1228, N1771);
not NOT1 (N2160, N2157);
and AND4 (N2161, N2160, N2119, N1162, N1318);
buf BUF1 (N2162, N2153);
nor NOR2 (N2163, N2162, N1997);
xor XOR2 (N2164, N2159, N60);
or OR4 (N2165, N2148, N1971, N212, N162);
buf BUF1 (N2166, N2158);
buf BUF1 (N2167, N2155);
nor NOR2 (N2168, N2161, N1744);
or OR2 (N2169, N2137, N1818);
xor XOR2 (N2170, N2167, N1585);
not NOT1 (N2171, N2165);
nor NOR2 (N2172, N2169, N1197);
and AND4 (N2173, N2168, N371, N1046, N1998);
or OR3 (N2174, N2172, N504, N141);
buf BUF1 (N2175, N2164);
buf BUF1 (N2176, N2163);
and AND3 (N2177, N2166, N555, N1848);
nor NOR4 (N2178, N2174, N1399, N1196, N1962);
and AND3 (N2179, N2175, N1164, N898);
not NOT1 (N2180, N2150);
and AND3 (N2181, N2173, N1881, N1440);
nand NAND2 (N2182, N2177, N669);
buf BUF1 (N2183, N2170);
buf BUF1 (N2184, N2180);
or OR3 (N2185, N2171, N1044, N1169);
and AND4 (N2186, N2151, N379, N1390, N539);
buf BUF1 (N2187, N2183);
xor XOR2 (N2188, N2133, N1418);
not NOT1 (N2189, N2187);
and AND2 (N2190, N2188, N1055);
or OR2 (N2191, N2179, N1191);
xor XOR2 (N2192, N2190, N1306);
not NOT1 (N2193, N2181);
buf BUF1 (N2194, N2186);
nand NAND2 (N2195, N2184, N674);
xor XOR2 (N2196, N2195, N1438);
not NOT1 (N2197, N2196);
nand NAND3 (N2198, N2197, N2182, N1443);
buf BUF1 (N2199, N1305);
or OR3 (N2200, N2193, N363, N150);
and AND4 (N2201, N2194, N1543, N1870, N1666);
buf BUF1 (N2202, N2198);
not NOT1 (N2203, N2176);
xor XOR2 (N2204, N2185, N1288);
not NOT1 (N2205, N2200);
xor XOR2 (N2206, N2191, N2013);
nand NAND2 (N2207, N2203, N246);
nor NOR3 (N2208, N2204, N2183, N1194);
or OR3 (N2209, N2189, N1711, N1380);
xor XOR2 (N2210, N2201, N1296);
buf BUF1 (N2211, N2210);
nand NAND3 (N2212, N2206, N1187, N2187);
not NOT1 (N2213, N2202);
xor XOR2 (N2214, N2178, N1446);
or OR3 (N2215, N2192, N1137, N1084);
nand NAND4 (N2216, N2207, N1349, N1675, N977);
not NOT1 (N2217, N2216);
buf BUF1 (N2218, N2209);
nor NOR3 (N2219, N2218, N1452, N22);
nand NAND4 (N2220, N2211, N1199, N304, N1469);
and AND2 (N2221, N2217, N908);
buf BUF1 (N2222, N2199);
buf BUF1 (N2223, N2222);
not NOT1 (N2224, N2220);
nor NOR4 (N2225, N2214, N1291, N1953, N589);
buf BUF1 (N2226, N2225);
nand NAND2 (N2227, N2219, N1084);
buf BUF1 (N2228, N2226);
buf BUF1 (N2229, N2224);
not NOT1 (N2230, N2213);
not NOT1 (N2231, N2205);
nor NOR3 (N2232, N2208, N234, N2135);
nor NOR2 (N2233, N2228, N1408);
not NOT1 (N2234, N2215);
nor NOR4 (N2235, N2221, N1826, N815, N1534);
not NOT1 (N2236, N2233);
xor XOR2 (N2237, N2223, N994);
xor XOR2 (N2238, N2230, N1074);
nand NAND2 (N2239, N2232, N1663);
nand NAND4 (N2240, N2234, N1379, N2185, N719);
xor XOR2 (N2241, N2236, N2157);
or OR3 (N2242, N2241, N1929, N920);
buf BUF1 (N2243, N2242);
and AND4 (N2244, N2235, N2167, N897, N1960);
and AND2 (N2245, N2212, N1837);
xor XOR2 (N2246, N2240, N412);
nor NOR4 (N2247, N2227, N1810, N396, N1358);
not NOT1 (N2248, N2238);
nand NAND4 (N2249, N2245, N1955, N888, N678);
buf BUF1 (N2250, N2229);
or OR3 (N2251, N2243, N134, N543);
not NOT1 (N2252, N2250);
or OR3 (N2253, N2247, N526, N1824);
and AND2 (N2254, N2239, N575);
or OR4 (N2255, N2237, N378, N1347, N836);
nor NOR4 (N2256, N2231, N1765, N1206, N1059);
nand NAND2 (N2257, N2251, N100);
nand NAND2 (N2258, N2256, N5);
or OR4 (N2259, N2252, N1133, N2170, N746);
buf BUF1 (N2260, N2258);
nor NOR3 (N2261, N2253, N876, N578);
nand NAND3 (N2262, N2248, N623, N2075);
nand NAND2 (N2263, N2257, N1593);
nand NAND2 (N2264, N2244, N1481);
buf BUF1 (N2265, N2262);
nor NOR4 (N2266, N2265, N1337, N11, N65);
and AND2 (N2267, N2249, N2259);
or OR4 (N2268, N1967, N893, N1324, N1359);
xor XOR2 (N2269, N2267, N354);
or OR4 (N2270, N2260, N1316, N2069, N623);
xor XOR2 (N2271, N2270, N2066);
nand NAND2 (N2272, N2266, N1426);
and AND3 (N2273, N2264, N1647, N248);
nor NOR3 (N2274, N2271, N740, N230);
nor NOR2 (N2275, N2263, N1744);
or OR3 (N2276, N2254, N1113, N894);
and AND2 (N2277, N2261, N282);
not NOT1 (N2278, N2272);
nand NAND3 (N2279, N2255, N1276, N1965);
or OR4 (N2280, N2275, N1553, N811, N2005);
buf BUF1 (N2281, N2276);
nand NAND3 (N2282, N2279, N2156, N1754);
xor XOR2 (N2283, N2281, N1108);
nand NAND4 (N2284, N2277, N400, N976, N887);
xor XOR2 (N2285, N2280, N1528);
nand NAND2 (N2286, N2285, N1774);
and AND3 (N2287, N2278, N841, N1080);
or OR3 (N2288, N2282, N1514, N1996);
not NOT1 (N2289, N2246);
not NOT1 (N2290, N2273);
and AND2 (N2291, N2269, N50);
nor NOR4 (N2292, N2291, N372, N684, N262);
and AND4 (N2293, N2286, N867, N1554, N1005);
or OR4 (N2294, N2284, N1520, N1813, N1367);
not NOT1 (N2295, N2294);
nor NOR4 (N2296, N2289, N1297, N1359, N859);
nor NOR2 (N2297, N2287, N985);
or OR3 (N2298, N2268, N624, N1160);
and AND4 (N2299, N2293, N1294, N1116, N2221);
not NOT1 (N2300, N2292);
nor NOR3 (N2301, N2297, N1049, N987);
not NOT1 (N2302, N2296);
or OR4 (N2303, N2288, N1418, N91, N1043);
nor NOR4 (N2304, N2295, N88, N457, N251);
nand NAND4 (N2305, N2304, N76, N120, N174);
nor NOR3 (N2306, N2283, N2139, N897);
or OR2 (N2307, N2299, N2029);
and AND2 (N2308, N2301, N1317);
or OR3 (N2309, N2305, N1412, N2290);
nor NOR3 (N2310, N85, N988, N2092);
nor NOR4 (N2311, N2306, N228, N2095, N1496);
xor XOR2 (N2312, N2311, N732);
or OR2 (N2313, N2308, N1768);
and AND3 (N2314, N2274, N549, N710);
xor XOR2 (N2315, N2314, N1044);
and AND4 (N2316, N2309, N1089, N1210, N1663);
buf BUF1 (N2317, N2313);
or OR4 (N2318, N2302, N624, N148, N483);
and AND3 (N2319, N2307, N2175, N304);
buf BUF1 (N2320, N2316);
not NOT1 (N2321, N2315);
buf BUF1 (N2322, N2303);
or OR4 (N2323, N2312, N1967, N247, N319);
nand NAND3 (N2324, N2300, N354, N1696);
not NOT1 (N2325, N2322);
xor XOR2 (N2326, N2325, N59);
or OR2 (N2327, N2326, N1415);
nor NOR3 (N2328, N2310, N1860, N2307);
or OR2 (N2329, N2320, N1851);
not NOT1 (N2330, N2329);
nor NOR2 (N2331, N2298, N696);
and AND3 (N2332, N2323, N1151, N2000);
xor XOR2 (N2333, N2321, N1223);
or OR4 (N2334, N2332, N1766, N208, N281);
buf BUF1 (N2335, N2319);
xor XOR2 (N2336, N2330, N1703);
and AND4 (N2337, N2335, N798, N673, N2143);
xor XOR2 (N2338, N2317, N1846);
nand NAND4 (N2339, N2328, N299, N1082, N1549);
xor XOR2 (N2340, N2339, N2207);
and AND4 (N2341, N2318, N72, N623, N234);
not NOT1 (N2342, N2340);
xor XOR2 (N2343, N2324, N510);
and AND3 (N2344, N2334, N2080, N1318);
buf BUF1 (N2345, N2343);
xor XOR2 (N2346, N2333, N1602);
xor XOR2 (N2347, N2345, N1056);
not NOT1 (N2348, N2347);
and AND2 (N2349, N2342, N1533);
nand NAND3 (N2350, N2331, N894, N1262);
not NOT1 (N2351, N2348);
not NOT1 (N2352, N2349);
buf BUF1 (N2353, N2336);
not NOT1 (N2354, N2346);
buf BUF1 (N2355, N2354);
buf BUF1 (N2356, N2350);
and AND2 (N2357, N2337, N2321);
nand NAND4 (N2358, N2353, N274, N277, N1290);
and AND4 (N2359, N2341, N2173, N1, N1972);
nand NAND3 (N2360, N2356, N2137, N495);
or OR3 (N2361, N2355, N2360, N251);
and AND4 (N2362, N1624, N30, N2008, N2204);
and AND3 (N2363, N2352, N1995, N52);
and AND2 (N2364, N2351, N388);
and AND3 (N2365, N2338, N1371, N187);
nand NAND4 (N2366, N2363, N289, N484, N381);
not NOT1 (N2367, N2362);
and AND4 (N2368, N2359, N2191, N2249, N1611);
and AND4 (N2369, N2344, N539, N2084, N1317);
and AND4 (N2370, N2367, N1348, N2225, N1652);
nand NAND2 (N2371, N2369, N1409);
buf BUF1 (N2372, N2371);
buf BUF1 (N2373, N2357);
nand NAND2 (N2374, N2368, N1916);
xor XOR2 (N2375, N2366, N1209);
and AND3 (N2376, N2375, N1795, N1450);
xor XOR2 (N2377, N2364, N1020);
nor NOR4 (N2378, N2377, N476, N325, N1330);
not NOT1 (N2379, N2361);
or OR2 (N2380, N2379, N1037);
not NOT1 (N2381, N2376);
nand NAND4 (N2382, N2372, N645, N256, N303);
or OR4 (N2383, N2374, N681, N415, N993);
or OR2 (N2384, N2378, N2079);
xor XOR2 (N2385, N2382, N1476);
or OR4 (N2386, N2373, N1442, N722, N615);
or OR2 (N2387, N2383, N2231);
buf BUF1 (N2388, N2365);
and AND2 (N2389, N2388, N1850);
nor NOR3 (N2390, N2389, N599, N1511);
xor XOR2 (N2391, N2385, N1879);
nand NAND3 (N2392, N2370, N2178, N1571);
nand NAND3 (N2393, N2384, N273, N2123);
xor XOR2 (N2394, N2327, N1060);
xor XOR2 (N2395, N2394, N1298);
nand NAND2 (N2396, N2386, N1752);
not NOT1 (N2397, N2396);
or OR4 (N2398, N2380, N1377, N1395, N2303);
nor NOR2 (N2399, N2358, N538);
or OR4 (N2400, N2391, N815, N44, N2393);
not NOT1 (N2401, N1513);
buf BUF1 (N2402, N2387);
xor XOR2 (N2403, N2402, N550);
nor NOR3 (N2404, N2399, N1682, N147);
and AND3 (N2405, N2390, N1876, N1683);
and AND3 (N2406, N2398, N697, N251);
buf BUF1 (N2407, N2397);
buf BUF1 (N2408, N2407);
and AND3 (N2409, N2403, N1951, N2408);
buf BUF1 (N2410, N2321);
buf BUF1 (N2411, N2405);
and AND3 (N2412, N2395, N769, N2306);
nor NOR2 (N2413, N2381, N2391);
not NOT1 (N2414, N2400);
nor NOR3 (N2415, N2409, N613, N740);
not NOT1 (N2416, N2413);
nor NOR4 (N2417, N2415, N2384, N195, N1661);
buf BUF1 (N2418, N2412);
nor NOR3 (N2419, N2401, N2306, N1218);
xor XOR2 (N2420, N2392, N523);
buf BUF1 (N2421, N2419);
nor NOR4 (N2422, N2404, N1137, N532, N347);
buf BUF1 (N2423, N2422);
and AND2 (N2424, N2418, N230);
and AND3 (N2425, N2417, N1684, N787);
not NOT1 (N2426, N2410);
nand NAND2 (N2427, N2420, N1772);
nor NOR4 (N2428, N2421, N2329, N728, N812);
buf BUF1 (N2429, N2411);
nor NOR3 (N2430, N2428, N120, N128);
buf BUF1 (N2431, N2427);
or OR4 (N2432, N2431, N407, N553, N1357);
and AND2 (N2433, N2425, N1476);
xor XOR2 (N2434, N2432, N1130);
or OR4 (N2435, N2426, N1109, N1126, N1716);
nand NAND3 (N2436, N2416, N1080, N552);
nor NOR2 (N2437, N2406, N1698);
nor NOR4 (N2438, N2436, N1777, N1788, N752);
nor NOR2 (N2439, N2429, N2187);
and AND4 (N2440, N2439, N1382, N1927, N2280);
buf BUF1 (N2441, N2435);
buf BUF1 (N2442, N2434);
xor XOR2 (N2443, N2438, N20);
or OR3 (N2444, N2433, N107, N618);
or OR4 (N2445, N2424, N1512, N1237, N811);
xor XOR2 (N2446, N2440, N991);
xor XOR2 (N2447, N2443, N1094);
buf BUF1 (N2448, N2441);
and AND3 (N2449, N2446, N308, N998);
not NOT1 (N2450, N2444);
not NOT1 (N2451, N2448);
xor XOR2 (N2452, N2449, N2352);
and AND4 (N2453, N2445, N1937, N175, N1458);
and AND3 (N2454, N2452, N2361, N110);
buf BUF1 (N2455, N2450);
and AND3 (N2456, N2455, N1276, N2091);
not NOT1 (N2457, N2454);
xor XOR2 (N2458, N2423, N483);
buf BUF1 (N2459, N2451);
buf BUF1 (N2460, N2414);
or OR3 (N2461, N2437, N1314, N2156);
and AND3 (N2462, N2456, N2053, N1536);
nand NAND2 (N2463, N2447, N248);
nand NAND2 (N2464, N2459, N696);
nor NOR2 (N2465, N2464, N2436);
not NOT1 (N2466, N2460);
xor XOR2 (N2467, N2466, N1237);
nand NAND4 (N2468, N2463, N1326, N1157, N864);
and AND4 (N2469, N2458, N571, N10, N801);
not NOT1 (N2470, N2461);
or OR3 (N2471, N2467, N1835, N44);
nor NOR3 (N2472, N2442, N155, N2242);
nor NOR3 (N2473, N2453, N677, N1890);
or OR4 (N2474, N2473, N611, N2418, N2238);
xor XOR2 (N2475, N2470, N1947);
and AND2 (N2476, N2471, N1403);
or OR2 (N2477, N2457, N614);
and AND3 (N2478, N2472, N1421, N453);
not NOT1 (N2479, N2477);
or OR2 (N2480, N2430, N527);
and AND3 (N2481, N2475, N174, N656);
nand NAND2 (N2482, N2462, N760);
or OR3 (N2483, N2480, N2065, N812);
nor NOR2 (N2484, N2465, N1842);
nand NAND4 (N2485, N2474, N470, N1001, N837);
nor NOR4 (N2486, N2484, N2417, N1070, N710);
and AND2 (N2487, N2469, N991);
buf BUF1 (N2488, N2481);
and AND3 (N2489, N2486, N747, N1446);
nand NAND4 (N2490, N2476, N1457, N455, N2106);
not NOT1 (N2491, N2488);
buf BUF1 (N2492, N2489);
not NOT1 (N2493, N2485);
nand NAND4 (N2494, N2493, N1607, N2301, N1157);
nor NOR2 (N2495, N2487, N2408);
or OR4 (N2496, N2491, N2262, N1900, N860);
nor NOR3 (N2497, N2482, N1200, N1600);
nand NAND2 (N2498, N2479, N2009);
buf BUF1 (N2499, N2492);
nand NAND3 (N2500, N2496, N780, N414);
nor NOR3 (N2501, N2483, N1053, N1609);
xor XOR2 (N2502, N2499, N1956);
nor NOR4 (N2503, N2490, N9, N1518, N507);
and AND3 (N2504, N2503, N505, N254);
nand NAND4 (N2505, N2500, N380, N530, N736);
and AND2 (N2506, N2498, N1922);
nor NOR2 (N2507, N2494, N1868);
not NOT1 (N2508, N2504);
buf BUF1 (N2509, N2505);
and AND4 (N2510, N2468, N783, N1301, N358);
not NOT1 (N2511, N2502);
not NOT1 (N2512, N2478);
nor NOR4 (N2513, N2510, N1907, N2205, N1763);
nand NAND2 (N2514, N2511, N1136);
nand NAND4 (N2515, N2507, N822, N615, N2272);
nor NOR4 (N2516, N2514, N665, N1054, N1798);
xor XOR2 (N2517, N2495, N1594);
not NOT1 (N2518, N2515);
nand NAND4 (N2519, N2518, N1473, N1103, N2009);
or OR4 (N2520, N2516, N161, N2212, N889);
and AND2 (N2521, N2501, N898);
and AND3 (N2522, N2509, N515, N816);
xor XOR2 (N2523, N2521, N2181);
buf BUF1 (N2524, N2517);
xor XOR2 (N2525, N2524, N1825);
and AND3 (N2526, N2523, N601, N1490);
and AND2 (N2527, N2513, N107);
xor XOR2 (N2528, N2520, N2133);
not NOT1 (N2529, N2519);
buf BUF1 (N2530, N2528);
and AND3 (N2531, N2522, N2046, N841);
nor NOR4 (N2532, N2506, N1595, N1235, N2340);
not NOT1 (N2533, N2497);
or OR3 (N2534, N2512, N1447, N211);
and AND3 (N2535, N2533, N1560, N2139);
nand NAND3 (N2536, N2530, N1393, N1034);
and AND4 (N2537, N2535, N1173, N1668, N7);
and AND2 (N2538, N2508, N1891);
or OR3 (N2539, N2532, N1406, N847);
nor NOR3 (N2540, N2537, N1544, N2332);
or OR4 (N2541, N2527, N574, N376, N38);
buf BUF1 (N2542, N2536);
nand NAND2 (N2543, N2539, N477);
and AND2 (N2544, N2534, N151);
nand NAND2 (N2545, N2526, N911);
or OR2 (N2546, N2541, N2485);
or OR4 (N2547, N2529, N959, N2386, N1693);
nor NOR2 (N2548, N2544, N1617);
nand NAND4 (N2549, N2540, N982, N135, N1409);
nor NOR2 (N2550, N2543, N1814);
or OR4 (N2551, N2545, N2505, N2283, N2416);
or OR4 (N2552, N2550, N1316, N57, N1603);
not NOT1 (N2553, N2542);
buf BUF1 (N2554, N2547);
buf BUF1 (N2555, N2538);
or OR4 (N2556, N2548, N711, N1891, N306);
nand NAND2 (N2557, N2552, N2215);
xor XOR2 (N2558, N2531, N58);
buf BUF1 (N2559, N2546);
xor XOR2 (N2560, N2559, N2113);
buf BUF1 (N2561, N2557);
xor XOR2 (N2562, N2561, N2550);
nand NAND4 (N2563, N2555, N614, N1200, N1710);
not NOT1 (N2564, N2554);
nand NAND4 (N2565, N2525, N2279, N511, N1701);
nor NOR2 (N2566, N2565, N2103);
nand NAND3 (N2567, N2558, N1262, N1086);
nor NOR2 (N2568, N2549, N520);
or OR3 (N2569, N2562, N2180, N780);
and AND4 (N2570, N2553, N543, N2538, N805);
and AND2 (N2571, N2560, N407);
nor NOR3 (N2572, N2567, N1830, N2208);
nor NOR3 (N2573, N2568, N2484, N785);
or OR4 (N2574, N2569, N828, N1122, N196);
xor XOR2 (N2575, N2551, N828);
nand NAND3 (N2576, N2564, N1600, N2460);
buf BUF1 (N2577, N2571);
xor XOR2 (N2578, N2574, N1665);
nand NAND4 (N2579, N2573, N2373, N1909, N1034);
and AND3 (N2580, N2575, N2344, N1640);
nor NOR3 (N2581, N2580, N70, N957);
and AND3 (N2582, N2556, N57, N454);
buf BUF1 (N2583, N2566);
xor XOR2 (N2584, N2572, N765);
buf BUF1 (N2585, N2579);
nand NAND3 (N2586, N2570, N422, N2317);
xor XOR2 (N2587, N2578, N592);
xor XOR2 (N2588, N2576, N1509);
nor NOR4 (N2589, N2577, N1078, N1346, N1523);
xor XOR2 (N2590, N2581, N2581);
buf BUF1 (N2591, N2588);
nand NAND3 (N2592, N2582, N1439, N2165);
nand NAND3 (N2593, N2590, N1875, N2398);
buf BUF1 (N2594, N2583);
buf BUF1 (N2595, N2586);
buf BUF1 (N2596, N2591);
not NOT1 (N2597, N2585);
and AND3 (N2598, N2587, N1627, N966);
or OR2 (N2599, N2584, N300);
buf BUF1 (N2600, N2589);
xor XOR2 (N2601, N2563, N465);
nand NAND4 (N2602, N2596, N2464, N1111, N358);
nand NAND2 (N2603, N2598, N2435);
or OR4 (N2604, N2592, N2438, N1134, N1478);
nand NAND4 (N2605, N2594, N2060, N2201, N1924);
nor NOR4 (N2606, N2597, N1719, N436, N2372);
xor XOR2 (N2607, N2602, N954);
buf BUF1 (N2608, N2607);
xor XOR2 (N2609, N2599, N2020);
nor NOR2 (N2610, N2608, N998);
not NOT1 (N2611, N2609);
nand NAND3 (N2612, N2605, N1120, N1392);
xor XOR2 (N2613, N2593, N2586);
nand NAND2 (N2614, N2606, N2113);
and AND4 (N2615, N2595, N1165, N2552, N1447);
nor NOR2 (N2616, N2612, N479);
buf BUF1 (N2617, N2613);
buf BUF1 (N2618, N2615);
and AND3 (N2619, N2611, N1307, N48);
and AND3 (N2620, N2601, N1079, N2581);
or OR4 (N2621, N2618, N2305, N524, N2499);
and AND2 (N2622, N2617, N1761);
and AND4 (N2623, N2619, N124, N1298, N242);
xor XOR2 (N2624, N2603, N2387);
and AND3 (N2625, N2610, N2606, N414);
and AND3 (N2626, N2625, N1892, N1670);
not NOT1 (N2627, N2616);
not NOT1 (N2628, N2614);
buf BUF1 (N2629, N2624);
not NOT1 (N2630, N2621);
and AND4 (N2631, N2627, N1190, N164, N1377);
and AND4 (N2632, N2626, N590, N2227, N722);
nor NOR4 (N2633, N2631, N803, N2466, N629);
nand NAND4 (N2634, N2604, N1838, N789, N615);
xor XOR2 (N2635, N2633, N279);
not NOT1 (N2636, N2628);
xor XOR2 (N2637, N2634, N675);
and AND2 (N2638, N2622, N1126);
xor XOR2 (N2639, N2632, N1441);
buf BUF1 (N2640, N2630);
or OR2 (N2641, N2629, N2484);
nand NAND4 (N2642, N2641, N2545, N1607, N2160);
and AND2 (N2643, N2638, N2585);
not NOT1 (N2644, N2635);
buf BUF1 (N2645, N2620);
and AND3 (N2646, N2644, N2635, N2556);
nor NOR3 (N2647, N2642, N43, N678);
or OR3 (N2648, N2645, N2031, N135);
nor NOR3 (N2649, N2600, N2309, N418);
and AND4 (N2650, N2647, N1571, N267, N134);
xor XOR2 (N2651, N2643, N1365);
nor NOR4 (N2652, N2648, N892, N2231, N703);
or OR3 (N2653, N2637, N2463, N2268);
nor NOR2 (N2654, N2652, N2425);
nor NOR3 (N2655, N2636, N1393, N2268);
nor NOR4 (N2656, N2646, N1146, N1984, N1274);
or OR3 (N2657, N2623, N968, N1576);
and AND3 (N2658, N2639, N2451, N2242);
or OR3 (N2659, N2657, N1239, N777);
nor NOR2 (N2660, N2656, N256);
or OR4 (N2661, N2640, N1668, N804, N2017);
or OR3 (N2662, N2653, N477, N1017);
or OR4 (N2663, N2659, N2549, N1990, N1670);
nand NAND2 (N2664, N2654, N985);
not NOT1 (N2665, N2661);
buf BUF1 (N2666, N2649);
or OR2 (N2667, N2660, N2593);
nor NOR2 (N2668, N2664, N2207);
buf BUF1 (N2669, N2651);
and AND4 (N2670, N2655, N1276, N1660, N1173);
or OR4 (N2671, N2667, N1690, N2342, N2333);
and AND4 (N2672, N2658, N1536, N201, N2337);
xor XOR2 (N2673, N2662, N663);
xor XOR2 (N2674, N2665, N567);
or OR4 (N2675, N2674, N1683, N1603, N1709);
nor NOR4 (N2676, N2650, N897, N2007, N617);
or OR4 (N2677, N2671, N2082, N419, N1615);
or OR3 (N2678, N2670, N1934, N683);
xor XOR2 (N2679, N2668, N651);
nor NOR2 (N2680, N2666, N1079);
not NOT1 (N2681, N2663);
not NOT1 (N2682, N2679);
or OR2 (N2683, N2672, N357);
nand NAND4 (N2684, N2676, N2389, N678, N2371);
and AND4 (N2685, N2673, N207, N2673, N1972);
buf BUF1 (N2686, N2681);
xor XOR2 (N2687, N2680, N1385);
nand NAND3 (N2688, N2677, N2092, N718);
nor NOR4 (N2689, N2687, N1369, N1986, N1248);
and AND4 (N2690, N2682, N360, N67, N115);
nand NAND2 (N2691, N2688, N2103);
nor NOR3 (N2692, N2683, N857, N2654);
and AND4 (N2693, N2678, N949, N471, N1876);
nand NAND2 (N2694, N2689, N990);
not NOT1 (N2695, N2686);
xor XOR2 (N2696, N2690, N1401);
or OR4 (N2697, N2675, N1472, N2589, N2290);
nand NAND2 (N2698, N2669, N2318);
buf BUF1 (N2699, N2696);
and AND4 (N2700, N2684, N2600, N1961, N1430);
not NOT1 (N2701, N2691);
xor XOR2 (N2702, N2694, N916);
or OR3 (N2703, N2685, N1879, N696);
not NOT1 (N2704, N2697);
nor NOR4 (N2705, N2702, N921, N2456, N2317);
buf BUF1 (N2706, N2698);
nor NOR3 (N2707, N2692, N764, N840);
nand NAND2 (N2708, N2703, N2565);
xor XOR2 (N2709, N2707, N2676);
nor NOR4 (N2710, N2699, N505, N1762, N2699);
and AND4 (N2711, N2708, N916, N828, N999);
not NOT1 (N2712, N2706);
buf BUF1 (N2713, N2710);
nand NAND4 (N2714, N2693, N1150, N1820, N1781);
or OR2 (N2715, N2709, N1182);
buf BUF1 (N2716, N2712);
xor XOR2 (N2717, N2711, N279);
xor XOR2 (N2718, N2717, N2156);
not NOT1 (N2719, N2713);
buf BUF1 (N2720, N2716);
and AND4 (N2721, N2715, N84, N467, N634);
and AND3 (N2722, N2719, N1251, N410);
or OR3 (N2723, N2721, N1215, N2309);
not NOT1 (N2724, N2720);
or OR3 (N2725, N2724, N1926, N513);
and AND4 (N2726, N2722, N313, N2246, N1780);
not NOT1 (N2727, N2695);
buf BUF1 (N2728, N2725);
xor XOR2 (N2729, N2727, N1063);
nor NOR3 (N2730, N2718, N246, N206);
nand NAND2 (N2731, N2723, N2288);
or OR3 (N2732, N2729, N1505, N1736);
or OR3 (N2733, N2701, N1668, N1174);
nand NAND3 (N2734, N2704, N320, N217);
and AND4 (N2735, N2726, N1006, N1474, N2705);
or OR2 (N2736, N1489, N1513);
xor XOR2 (N2737, N2734, N628);
or OR3 (N2738, N2733, N1989, N1295);
and AND3 (N2739, N2730, N1160, N1748);
nor NOR4 (N2740, N2714, N1691, N1605, N1654);
or OR3 (N2741, N2731, N1913, N947);
buf BUF1 (N2742, N2737);
nand NAND4 (N2743, N2738, N1646, N1619, N1850);
and AND3 (N2744, N2735, N1383, N174);
nor NOR3 (N2745, N2742, N2303, N82);
nand NAND4 (N2746, N2728, N562, N1027, N1327);
not NOT1 (N2747, N2739);
not NOT1 (N2748, N2732);
nand NAND2 (N2749, N2745, N964);
xor XOR2 (N2750, N2741, N1104);
nand NAND2 (N2751, N2746, N52);
not NOT1 (N2752, N2700);
and AND2 (N2753, N2752, N677);
xor XOR2 (N2754, N2744, N2495);
or OR4 (N2755, N2754, N2102, N194, N1003);
and AND3 (N2756, N2755, N2333, N1655);
buf BUF1 (N2757, N2753);
or OR2 (N2758, N2751, N2349);
xor XOR2 (N2759, N2757, N2453);
or OR2 (N2760, N2758, N2252);
or OR4 (N2761, N2740, N1751, N2413, N1786);
xor XOR2 (N2762, N2748, N2592);
or OR2 (N2763, N2756, N2105);
nand NAND4 (N2764, N2762, N360, N552, N2321);
nand NAND4 (N2765, N2747, N358, N2646, N1933);
buf BUF1 (N2766, N2759);
nor NOR4 (N2767, N2743, N1736, N1899, N960);
not NOT1 (N2768, N2750);
xor XOR2 (N2769, N2764, N872);
xor XOR2 (N2770, N2763, N1535);
nor NOR3 (N2771, N2770, N2027, N54);
nor NOR3 (N2772, N2765, N1889, N1328);
nand NAND3 (N2773, N2768, N1403, N175);
nor NOR3 (N2774, N2736, N1528, N176);
buf BUF1 (N2775, N2769);
or OR2 (N2776, N2775, N1640);
xor XOR2 (N2777, N2767, N1561);
buf BUF1 (N2778, N2771);
nand NAND2 (N2779, N2766, N1038);
or OR2 (N2780, N2778, N2276);
nand NAND3 (N2781, N2760, N549, N1234);
or OR2 (N2782, N2777, N1370);
or OR3 (N2783, N2782, N1530, N2725);
nor NOR2 (N2784, N2776, N1022);
not NOT1 (N2785, N2784);
nor NOR3 (N2786, N2785, N2411, N1183);
nor NOR4 (N2787, N2786, N2300, N922, N2163);
xor XOR2 (N2788, N2779, N1354);
buf BUF1 (N2789, N2787);
or OR4 (N2790, N2789, N2684, N2180, N2299);
nor NOR2 (N2791, N2772, N2117);
xor XOR2 (N2792, N2780, N1772);
not NOT1 (N2793, N2773);
and AND4 (N2794, N2774, N1310, N1905, N1578);
not NOT1 (N2795, N2794);
or OR2 (N2796, N2788, N2446);
not NOT1 (N2797, N2761);
not NOT1 (N2798, N2796);
buf BUF1 (N2799, N2749);
and AND2 (N2800, N2791, N425);
buf BUF1 (N2801, N2799);
and AND2 (N2802, N2783, N2047);
nor NOR2 (N2803, N2792, N265);
or OR4 (N2804, N2800, N1960, N1410, N2077);
or OR2 (N2805, N2798, N2108);
nand NAND2 (N2806, N2781, N1598);
or OR2 (N2807, N2790, N307);
or OR4 (N2808, N2795, N148, N31, N966);
not NOT1 (N2809, N2803);
not NOT1 (N2810, N2806);
and AND3 (N2811, N2802, N1658, N358);
nor NOR3 (N2812, N2793, N1407, N885);
not NOT1 (N2813, N2809);
xor XOR2 (N2814, N2813, N2033);
nand NAND3 (N2815, N2805, N224, N1281);
nor NOR2 (N2816, N2812, N2663);
or OR2 (N2817, N2816, N2646);
and AND4 (N2818, N2808, N716, N130, N1085);
not NOT1 (N2819, N2797);
nand NAND4 (N2820, N2819, N1150, N1702, N570);
buf BUF1 (N2821, N2807);
and AND3 (N2822, N2818, N2497, N833);
not NOT1 (N2823, N2811);
not NOT1 (N2824, N2801);
xor XOR2 (N2825, N2804, N2621);
xor XOR2 (N2826, N2815, N601);
buf BUF1 (N2827, N2824);
not NOT1 (N2828, N2814);
nand NAND4 (N2829, N2821, N135, N2760, N1236);
and AND3 (N2830, N2823, N1295, N1273);
buf BUF1 (N2831, N2826);
xor XOR2 (N2832, N2829, N863);
buf BUF1 (N2833, N2832);
buf BUF1 (N2834, N2820);
not NOT1 (N2835, N2831);
not NOT1 (N2836, N2810);
not NOT1 (N2837, N2835);
nor NOR3 (N2838, N2830, N2409, N1539);
xor XOR2 (N2839, N2836, N896);
nand NAND2 (N2840, N2822, N2577);
nand NAND3 (N2841, N2834, N126, N1948);
buf BUF1 (N2842, N2838);
and AND2 (N2843, N2839, N694);
and AND3 (N2844, N2827, N180, N2462);
or OR3 (N2845, N2817, N318, N1197);
not NOT1 (N2846, N2841);
buf BUF1 (N2847, N2846);
and AND2 (N2848, N2833, N1957);
buf BUF1 (N2849, N2840);
buf BUF1 (N2850, N2843);
xor XOR2 (N2851, N2842, N167);
or OR3 (N2852, N2844, N2148, N454);
xor XOR2 (N2853, N2852, N519);
or OR2 (N2854, N2825, N1364);
and AND2 (N2855, N2848, N1336);
and AND2 (N2856, N2850, N2459);
not NOT1 (N2857, N2851);
nand NAND4 (N2858, N2847, N2723, N1746, N790);
not NOT1 (N2859, N2837);
xor XOR2 (N2860, N2859, N1662);
nor NOR2 (N2861, N2853, N679);
nor NOR3 (N2862, N2860, N1509, N2126);
nor NOR2 (N2863, N2854, N2830);
nor NOR3 (N2864, N2845, N1796, N1878);
buf BUF1 (N2865, N2863);
not NOT1 (N2866, N2861);
nand NAND3 (N2867, N2865, N940, N2817);
nor NOR4 (N2868, N2857, N2194, N2035, N1566);
not NOT1 (N2869, N2855);
not NOT1 (N2870, N2828);
and AND3 (N2871, N2862, N567, N474);
nand NAND4 (N2872, N2849, N1371, N1508, N1951);
or OR3 (N2873, N2856, N1737, N2090);
nor NOR3 (N2874, N2872, N1576, N2569);
buf BUF1 (N2875, N2864);
and AND2 (N2876, N2873, N2796);
nand NAND2 (N2877, N2867, N1267);
nor NOR4 (N2878, N2874, N1021, N1189, N2068);
buf BUF1 (N2879, N2878);
and AND2 (N2880, N2866, N40);
buf BUF1 (N2881, N2875);
buf BUF1 (N2882, N2869);
and AND3 (N2883, N2871, N1451, N2253);
buf BUF1 (N2884, N2877);
buf BUF1 (N2885, N2882);
and AND3 (N2886, N2885, N2723, N2239);
not NOT1 (N2887, N2880);
nand NAND4 (N2888, N2887, N1218, N17, N2641);
not NOT1 (N2889, N2886);
and AND3 (N2890, N2870, N81, N1464);
or OR4 (N2891, N2879, N2340, N180, N2618);
or OR4 (N2892, N2890, N1352, N1646, N2719);
nor NOR2 (N2893, N2858, N1273);
not NOT1 (N2894, N2893);
nand NAND3 (N2895, N2892, N1596, N1058);
and AND2 (N2896, N2889, N1012);
and AND4 (N2897, N2883, N1511, N1045, N201);
xor XOR2 (N2898, N2876, N2620);
buf BUF1 (N2899, N2884);
or OR4 (N2900, N2899, N1766, N2538, N725);
nor NOR4 (N2901, N2888, N701, N2892, N1102);
nand NAND3 (N2902, N2897, N2310, N2181);
xor XOR2 (N2903, N2891, N2624);
xor XOR2 (N2904, N2868, N2601);
not NOT1 (N2905, N2903);
nor NOR4 (N2906, N2895, N2497, N2687, N2299);
nor NOR4 (N2907, N2904, N1039, N1404, N27);
nor NOR4 (N2908, N2905, N59, N2716, N2178);
nor NOR2 (N2909, N2894, N904);
nand NAND4 (N2910, N2896, N541, N2072, N1770);
or OR3 (N2911, N2908, N811, N2088);
or OR4 (N2912, N2911, N2159, N2237, N1103);
buf BUF1 (N2913, N2900);
or OR3 (N2914, N2898, N985, N538);
xor XOR2 (N2915, N2910, N1081);
not NOT1 (N2916, N2912);
xor XOR2 (N2917, N2915, N2814);
nand NAND2 (N2918, N2901, N1099);
xor XOR2 (N2919, N2902, N402);
nand NAND3 (N2920, N2907, N1861, N1443);
nand NAND4 (N2921, N2881, N2629, N1156, N2111);
and AND2 (N2922, N2906, N392);
or OR3 (N2923, N2916, N1976, N2907);
nand NAND4 (N2924, N2919, N2374, N222, N1916);
or OR3 (N2925, N2924, N594, N1654);
and AND4 (N2926, N2917, N2568, N1142, N1844);
buf BUF1 (N2927, N2926);
nor NOR2 (N2928, N2923, N225);
not NOT1 (N2929, N2918);
xor XOR2 (N2930, N2929, N41);
not NOT1 (N2931, N2909);
and AND3 (N2932, N2927, N74, N981);
not NOT1 (N2933, N2932);
xor XOR2 (N2934, N2921, N2236);
not NOT1 (N2935, N2933);
not NOT1 (N2936, N2914);
or OR3 (N2937, N2930, N208, N21);
or OR4 (N2938, N2920, N1624, N2037, N2224);
xor XOR2 (N2939, N2935, N2499);
or OR4 (N2940, N2936, N1694, N761, N1005);
nand NAND2 (N2941, N2938, N2192);
nor NOR3 (N2942, N2937, N419, N1644);
not NOT1 (N2943, N2942);
nor NOR3 (N2944, N2943, N1251, N2254);
buf BUF1 (N2945, N2925);
nor NOR4 (N2946, N2940, N2096, N2672, N1476);
and AND3 (N2947, N2922, N12, N449);
nand NAND4 (N2948, N2934, N917, N1347, N1788);
or OR4 (N2949, N2946, N2753, N79, N1957);
xor XOR2 (N2950, N2944, N1727);
or OR4 (N2951, N2949, N2621, N1892, N993);
or OR2 (N2952, N2948, N416);
or OR4 (N2953, N2928, N2832, N597, N2447);
and AND3 (N2954, N2950, N81, N1773);
nand NAND4 (N2955, N2947, N619, N1805, N1069);
or OR2 (N2956, N2951, N2288);
and AND4 (N2957, N2939, N2494, N2389, N1924);
or OR2 (N2958, N2956, N141);
nor NOR3 (N2959, N2954, N1376, N323);
and AND2 (N2960, N2952, N1990);
xor XOR2 (N2961, N2960, N2436);
not NOT1 (N2962, N2955);
and AND4 (N2963, N2941, N1391, N1826, N1927);
or OR2 (N2964, N2957, N526);
xor XOR2 (N2965, N2962, N879);
not NOT1 (N2966, N2959);
buf BUF1 (N2967, N2958);
or OR4 (N2968, N2967, N825, N2256, N2684);
and AND2 (N2969, N2913, N2186);
or OR2 (N2970, N2964, N2422);
nand NAND4 (N2971, N2965, N1784, N2054, N2089);
nor NOR3 (N2972, N2968, N664, N1731);
buf BUF1 (N2973, N2953);
buf BUF1 (N2974, N2972);
and AND4 (N2975, N2974, N1474, N67, N2959);
not NOT1 (N2976, N2969);
or OR2 (N2977, N2961, N926);
nor NOR4 (N2978, N2975, N2488, N1363, N648);
and AND2 (N2979, N2971, N963);
buf BUF1 (N2980, N2977);
or OR3 (N2981, N2970, N2475, N849);
or OR2 (N2982, N2945, N142);
buf BUF1 (N2983, N2963);
nand NAND4 (N2984, N2982, N2555, N2755, N1266);
nand NAND4 (N2985, N2931, N2604, N976, N926);
xor XOR2 (N2986, N2966, N671);
nand NAND4 (N2987, N2979, N1950, N2243, N1007);
buf BUF1 (N2988, N2984);
xor XOR2 (N2989, N2973, N152);
or OR2 (N2990, N2978, N2961);
or OR4 (N2991, N2976, N2242, N1621, N1172);
nand NAND3 (N2992, N2980, N2207, N1554);
and AND3 (N2993, N2983, N2708, N1235);
nand NAND3 (N2994, N2991, N1183, N2397);
nor NOR2 (N2995, N2992, N159);
not NOT1 (N2996, N2989);
not NOT1 (N2997, N2993);
nor NOR3 (N2998, N2987, N1648, N2447);
nor NOR2 (N2999, N2988, N153);
nor NOR2 (N3000, N2995, N473);
xor XOR2 (N3001, N3000, N2919);
and AND4 (N3002, N2996, N58, N2447, N1771);
buf BUF1 (N3003, N3001);
buf BUF1 (N3004, N2997);
nand NAND4 (N3005, N2994, N1281, N2727, N544);
xor XOR2 (N3006, N2990, N474);
nand NAND3 (N3007, N3003, N659, N853);
xor XOR2 (N3008, N3004, N616);
or OR3 (N3009, N2998, N3008, N506);
buf BUF1 (N3010, N54);
and AND3 (N3011, N3006, N99, N381);
nor NOR3 (N3012, N2999, N1691, N628);
xor XOR2 (N3013, N3002, N312);
nand NAND2 (N3014, N3010, N2779);
not NOT1 (N3015, N3009);
xor XOR2 (N3016, N2986, N115);
buf BUF1 (N3017, N2985);
not NOT1 (N3018, N3017);
xor XOR2 (N3019, N2981, N1627);
xor XOR2 (N3020, N3018, N1694);
nor NOR3 (N3021, N3005, N1780, N2363);
buf BUF1 (N3022, N3014);
or OR3 (N3023, N3019, N1126, N590);
nor NOR3 (N3024, N3023, N1282, N2351);
and AND2 (N3025, N3007, N1791);
or OR4 (N3026, N3016, N787, N736, N2357);
nand NAND4 (N3027, N3021, N1822, N2953, N2584);
or OR2 (N3028, N3027, N2231);
nand NAND4 (N3029, N3024, N2918, N1717, N213);
not NOT1 (N3030, N3028);
not NOT1 (N3031, N3029);
and AND2 (N3032, N3030, N2603);
nor NOR2 (N3033, N3011, N46);
and AND4 (N3034, N3022, N2889, N193, N1485);
not NOT1 (N3035, N3013);
and AND3 (N3036, N3012, N1753, N2072);
buf BUF1 (N3037, N3033);
xor XOR2 (N3038, N3025, N2413);
xor XOR2 (N3039, N3034, N212);
or OR2 (N3040, N3036, N1748);
or OR4 (N3041, N3020, N1834, N1723, N3022);
nor NOR2 (N3042, N3031, N1127);
nor NOR2 (N3043, N3037, N2985);
nor NOR2 (N3044, N3026, N2247);
not NOT1 (N3045, N3041);
and AND4 (N3046, N3032, N995, N2572, N1354);
buf BUF1 (N3047, N3046);
or OR3 (N3048, N3044, N324, N913);
buf BUF1 (N3049, N3043);
nor NOR3 (N3050, N3048, N2808, N774);
buf BUF1 (N3051, N3040);
nand NAND4 (N3052, N3035, N292, N1778, N2904);
and AND3 (N3053, N3039, N1355, N1834);
not NOT1 (N3054, N3042);
xor XOR2 (N3055, N3054, N858);
buf BUF1 (N3056, N3045);
not NOT1 (N3057, N3015);
or OR3 (N3058, N3052, N2778, N1103);
nand NAND2 (N3059, N3055, N154);
buf BUF1 (N3060, N3050);
nor NOR3 (N3061, N3059, N1002, N742);
not NOT1 (N3062, N3057);
buf BUF1 (N3063, N3060);
nor NOR2 (N3064, N3053, N1083);
nand NAND3 (N3065, N3062, N2027, N2168);
and AND3 (N3066, N3056, N2613, N1451);
nor NOR4 (N3067, N3064, N1604, N2288, N1056);
not NOT1 (N3068, N3051);
nor NOR3 (N3069, N3065, N165, N3058);
xor XOR2 (N3070, N2667, N251);
nand NAND2 (N3071, N3049, N2294);
and AND3 (N3072, N3063, N1249, N2693);
not NOT1 (N3073, N3069);
not NOT1 (N3074, N3066);
nor NOR4 (N3075, N3072, N488, N1541, N698);
and AND3 (N3076, N3038, N1969, N127);
not NOT1 (N3077, N3068);
and AND4 (N3078, N3067, N451, N1131, N970);
not NOT1 (N3079, N3047);
buf BUF1 (N3080, N3071);
not NOT1 (N3081, N3080);
not NOT1 (N3082, N3075);
not NOT1 (N3083, N3078);
nor NOR2 (N3084, N3073, N2837);
nand NAND4 (N3085, N3070, N913, N1590, N190);
nand NAND4 (N3086, N3082, N1275, N1552, N2608);
and AND2 (N3087, N3085, N2280);
buf BUF1 (N3088, N3079);
not NOT1 (N3089, N3084);
not NOT1 (N3090, N3076);
or OR4 (N3091, N3077, N182, N1413, N828);
buf BUF1 (N3092, N3061);
xor XOR2 (N3093, N3081, N1599);
xor XOR2 (N3094, N3088, N534);
or OR4 (N3095, N3094, N1623, N884, N871);
and AND3 (N3096, N3090, N1933, N369);
or OR4 (N3097, N3095, N286, N1055, N1002);
nand NAND2 (N3098, N3096, N1847);
xor XOR2 (N3099, N3097, N651);
or OR2 (N3100, N3098, N948);
nor NOR3 (N3101, N3091, N132, N410);
or OR3 (N3102, N3087, N619, N1235);
or OR4 (N3103, N3093, N2716, N2589, N730);
nand NAND3 (N3104, N3074, N2841, N2137);
nor NOR2 (N3105, N3104, N2340);
or OR3 (N3106, N3086, N1418, N533);
buf BUF1 (N3107, N3103);
and AND3 (N3108, N3107, N1028, N2763);
nand NAND3 (N3109, N3101, N2997, N1351);
nand NAND2 (N3110, N3106, N2635);
xor XOR2 (N3111, N3092, N1054);
nand NAND4 (N3112, N3102, N1166, N1864, N1931);
buf BUF1 (N3113, N3112);
buf BUF1 (N3114, N3089);
or OR4 (N3115, N3113, N736, N2127, N891);
nor NOR4 (N3116, N3114, N1190, N377, N1527);
and AND4 (N3117, N3116, N1963, N1856, N2490);
buf BUF1 (N3118, N3115);
buf BUF1 (N3119, N3099);
nor NOR3 (N3120, N3119, N2363, N2530);
not NOT1 (N3121, N3083);
nor NOR2 (N3122, N3117, N1588);
not NOT1 (N3123, N3105);
xor XOR2 (N3124, N3108, N1749);
not NOT1 (N3125, N3111);
and AND4 (N3126, N3100, N615, N23, N2505);
buf BUF1 (N3127, N3126);
buf BUF1 (N3128, N3121);
nor NOR3 (N3129, N3125, N2821, N1948);
nand NAND4 (N3130, N3128, N3003, N1765, N233);
nor NOR4 (N3131, N3124, N1441, N1879, N2814);
xor XOR2 (N3132, N3131, N2900);
not NOT1 (N3133, N3120);
nor NOR2 (N3134, N3127, N271);
not NOT1 (N3135, N3110);
not NOT1 (N3136, N3109);
and AND3 (N3137, N3134, N241, N1804);
and AND3 (N3138, N3133, N2963, N1093);
buf BUF1 (N3139, N3122);
not NOT1 (N3140, N3132);
not NOT1 (N3141, N3118);
nand NAND4 (N3142, N3130, N1890, N3111, N1940);
not NOT1 (N3143, N3138);
nand NAND4 (N3144, N3139, N468, N1611, N2455);
buf BUF1 (N3145, N3143);
buf BUF1 (N3146, N3136);
buf BUF1 (N3147, N3123);
or OR2 (N3148, N3146, N843);
or OR2 (N3149, N3147, N1828);
buf BUF1 (N3150, N3144);
buf BUF1 (N3151, N3142);
not NOT1 (N3152, N3141);
nor NOR2 (N3153, N3140, N826);
or OR4 (N3154, N3150, N1354, N3118, N1599);
not NOT1 (N3155, N3149);
nand NAND2 (N3156, N3154, N129);
or OR2 (N3157, N3129, N2422);
and AND3 (N3158, N3157, N468, N615);
nand NAND2 (N3159, N3135, N1977);
buf BUF1 (N3160, N3151);
buf BUF1 (N3161, N3152);
nand NAND4 (N3162, N3145, N226, N1884, N2570);
or OR4 (N3163, N3159, N1767, N335, N493);
not NOT1 (N3164, N3162);
or OR4 (N3165, N3148, N1462, N2772, N871);
nor NOR4 (N3166, N3160, N1123, N856, N31);
not NOT1 (N3167, N3163);
buf BUF1 (N3168, N3161);
not NOT1 (N3169, N3164);
and AND4 (N3170, N3168, N2834, N2243, N204);
not NOT1 (N3171, N3155);
buf BUF1 (N3172, N3169);
nor NOR3 (N3173, N3165, N390, N854);
and AND2 (N3174, N3137, N2884);
not NOT1 (N3175, N3173);
xor XOR2 (N3176, N3170, N1080);
nor NOR4 (N3177, N3156, N198, N139, N1636);
nand NAND2 (N3178, N3167, N2621);
nor NOR3 (N3179, N3171, N677, N2016);
nand NAND3 (N3180, N3153, N3087, N1341);
or OR3 (N3181, N3176, N1660, N2677);
not NOT1 (N3182, N3174);
nor NOR3 (N3183, N3175, N535, N1976);
nor NOR3 (N3184, N3180, N2768, N1174);
and AND4 (N3185, N3178, N146, N1002, N1675);
nor NOR2 (N3186, N3183, N2193);
or OR3 (N3187, N3186, N1207, N495);
not NOT1 (N3188, N3182);
or OR3 (N3189, N3187, N2680, N419);
nand NAND2 (N3190, N3181, N2815);
nand NAND3 (N3191, N3184, N3078, N2915);
xor XOR2 (N3192, N3166, N412);
nor NOR4 (N3193, N3189, N2078, N1261, N514);
nand NAND2 (N3194, N3191, N3134);
buf BUF1 (N3195, N3188);
buf BUF1 (N3196, N3195);
xor XOR2 (N3197, N3172, N678);
nor NOR2 (N3198, N3177, N1642);
or OR2 (N3199, N3185, N2316);
or OR4 (N3200, N3179, N275, N1319, N1978);
nand NAND2 (N3201, N3158, N1910);
or OR3 (N3202, N3194, N1249, N196);
buf BUF1 (N3203, N3197);
buf BUF1 (N3204, N3203);
buf BUF1 (N3205, N3201);
xor XOR2 (N3206, N3193, N3056);
nand NAND4 (N3207, N3205, N1374, N810, N1364);
not NOT1 (N3208, N3202);
buf BUF1 (N3209, N3208);
xor XOR2 (N3210, N3198, N2064);
buf BUF1 (N3211, N3192);
xor XOR2 (N3212, N3209, N947);
nand NAND3 (N3213, N3199, N788, N2233);
buf BUF1 (N3214, N3204);
and AND3 (N3215, N3211, N685, N2739);
not NOT1 (N3216, N3215);
nand NAND2 (N3217, N3196, N1772);
endmodule