// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N617,N607,N620,N622,N611,N623,N602,N619,N614,N624;

nor NOR2 (N25, N20, N16);
and AND2 (N26, N18, N14);
or OR2 (N27, N8, N1);
nor NOR3 (N28, N7, N9, N27);
nor NOR2 (N29, N9, N4);
and AND2 (N30, N19, N17);
nor NOR4 (N31, N1, N4, N10, N4);
not NOT1 (N32, N4);
or OR4 (N33, N12, N6, N9, N22);
nor NOR4 (N34, N17, N19, N21, N12);
xor XOR2 (N35, N30, N15);
not NOT1 (N36, N13);
not NOT1 (N37, N33);
nand NAND4 (N38, N37, N22, N10, N12);
or OR4 (N39, N29, N12, N15, N22);
xor XOR2 (N40, N25, N30);
not NOT1 (N41, N31);
buf BUF1 (N42, N28);
buf BUF1 (N43, N32);
or OR3 (N44, N39, N1, N28);
nor NOR2 (N45, N40, N3);
buf BUF1 (N46, N36);
nand NAND2 (N47, N45, N37);
xor XOR2 (N48, N35, N22);
or OR2 (N49, N46, N6);
nor NOR4 (N50, N34, N31, N13, N41);
not NOT1 (N51, N19);
nor NOR3 (N52, N44, N44, N51);
nand NAND4 (N53, N40, N17, N20, N52);
and AND3 (N54, N33, N3, N7);
or OR3 (N55, N53, N12, N50);
buf BUF1 (N56, N32);
xor XOR2 (N57, N26, N47);
not NOT1 (N58, N41);
and AND3 (N59, N48, N5, N10);
nand NAND3 (N60, N57, N41, N44);
xor XOR2 (N61, N56, N43);
and AND2 (N62, N51, N34);
buf BUF1 (N63, N61);
not NOT1 (N64, N42);
nand NAND4 (N65, N63, N40, N17, N9);
and AND2 (N66, N49, N48);
nor NOR3 (N67, N65, N16, N42);
and AND3 (N68, N58, N3, N35);
not NOT1 (N69, N62);
buf BUF1 (N70, N67);
or OR2 (N71, N69, N57);
xor XOR2 (N72, N55, N11);
nand NAND3 (N73, N38, N3, N33);
xor XOR2 (N74, N68, N3);
nand NAND2 (N75, N54, N62);
or OR2 (N76, N59, N22);
and AND3 (N77, N76, N73, N32);
and AND2 (N78, N22, N75);
xor XOR2 (N79, N39, N72);
and AND2 (N80, N12, N61);
and AND3 (N81, N70, N19, N65);
buf BUF1 (N82, N66);
not NOT1 (N83, N80);
nand NAND3 (N84, N60, N30, N10);
xor XOR2 (N85, N71, N81);
nand NAND3 (N86, N50, N33, N78);
nor NOR2 (N87, N41, N41);
nand NAND2 (N88, N82, N23);
and AND4 (N89, N83, N53, N25, N10);
not NOT1 (N90, N86);
and AND2 (N91, N79, N61);
nor NOR2 (N92, N84, N42);
xor XOR2 (N93, N77, N74);
and AND2 (N94, N21, N40);
not NOT1 (N95, N92);
or OR3 (N96, N91, N26, N23);
nor NOR2 (N97, N90, N65);
nand NAND3 (N98, N87, N60, N84);
or OR3 (N99, N97, N61, N20);
xor XOR2 (N100, N95, N42);
nor NOR3 (N101, N85, N13, N10);
nand NAND2 (N102, N93, N59);
nor NOR3 (N103, N88, N99, N90);
xor XOR2 (N104, N65, N80);
and AND4 (N105, N64, N85, N68, N61);
nor NOR4 (N106, N101, N85, N6, N80);
nand NAND3 (N107, N106, N30, N47);
buf BUF1 (N108, N104);
or OR2 (N109, N94, N37);
or OR3 (N110, N109, N3, N75);
not NOT1 (N111, N105);
nand NAND2 (N112, N111, N5);
nor NOR2 (N113, N112, N45);
nor NOR4 (N114, N107, N57, N62, N29);
and AND3 (N115, N103, N112, N53);
and AND3 (N116, N114, N55, N4);
xor XOR2 (N117, N102, N77);
nor NOR2 (N118, N96, N94);
nor NOR2 (N119, N113, N34);
or OR4 (N120, N98, N23, N119, N111);
nor NOR4 (N121, N20, N111, N35, N34);
not NOT1 (N122, N89);
or OR3 (N123, N116, N104, N1);
and AND2 (N124, N122, N112);
buf BUF1 (N125, N118);
or OR3 (N126, N115, N88, N13);
buf BUF1 (N127, N120);
and AND2 (N128, N126, N99);
nor NOR3 (N129, N121, N19, N43);
and AND4 (N130, N124, N22, N80, N46);
and AND3 (N131, N110, N76, N108);
and AND2 (N132, N56, N78);
not NOT1 (N133, N123);
nor NOR3 (N134, N130, N35, N103);
nand NAND2 (N135, N128, N124);
buf BUF1 (N136, N127);
xor XOR2 (N137, N100, N72);
or OR3 (N138, N129, N18, N63);
nor NOR3 (N139, N135, N104, N105);
xor XOR2 (N140, N131, N33);
buf BUF1 (N141, N136);
not NOT1 (N142, N117);
nand NAND2 (N143, N125, N125);
xor XOR2 (N144, N137, N61);
and AND3 (N145, N144, N3, N21);
xor XOR2 (N146, N145, N33);
or OR2 (N147, N142, N65);
not NOT1 (N148, N138);
xor XOR2 (N149, N148, N116);
xor XOR2 (N150, N140, N27);
nor NOR3 (N151, N133, N20, N53);
buf BUF1 (N152, N147);
and AND3 (N153, N146, N97, N116);
or OR3 (N154, N152, N64, N137);
buf BUF1 (N155, N153);
not NOT1 (N156, N141);
or OR4 (N157, N143, N109, N92, N104);
xor XOR2 (N158, N149, N118);
or OR3 (N159, N134, N96, N71);
buf BUF1 (N160, N132);
and AND4 (N161, N154, N124, N114, N154);
or OR2 (N162, N151, N16);
not NOT1 (N163, N150);
xor XOR2 (N164, N156, N96);
nand NAND2 (N165, N161, N66);
nor NOR4 (N166, N139, N46, N26, N33);
not NOT1 (N167, N165);
nand NAND2 (N168, N159, N37);
or OR3 (N169, N166, N142, N119);
nor NOR3 (N170, N164, N164, N90);
not NOT1 (N171, N158);
or OR4 (N172, N170, N56, N164, N93);
buf BUF1 (N173, N157);
buf BUF1 (N174, N172);
nor NOR3 (N175, N174, N152, N145);
nand NAND2 (N176, N169, N76);
and AND2 (N177, N175, N45);
xor XOR2 (N178, N162, N53);
or OR3 (N179, N155, N41, N104);
and AND3 (N180, N171, N96, N38);
or OR2 (N181, N167, N21);
or OR2 (N182, N180, N81);
and AND3 (N183, N163, N25, N89);
or OR4 (N184, N177, N147, N132, N21);
buf BUF1 (N185, N176);
xor XOR2 (N186, N181, N84);
xor XOR2 (N187, N179, N10);
or OR3 (N188, N187, N100, N118);
or OR3 (N189, N160, N68, N182);
not NOT1 (N190, N48);
not NOT1 (N191, N190);
and AND3 (N192, N191, N40, N174);
xor XOR2 (N193, N178, N54);
and AND4 (N194, N168, N163, N16, N46);
buf BUF1 (N195, N185);
nor NOR3 (N196, N189, N141, N153);
and AND3 (N197, N188, N140, N148);
nor NOR2 (N198, N197, N105);
nand NAND3 (N199, N183, N121, N129);
nor NOR4 (N200, N198, N46, N174, N74);
not NOT1 (N201, N195);
buf BUF1 (N202, N194);
nor NOR4 (N203, N200, N78, N143, N31);
buf BUF1 (N204, N201);
nand NAND3 (N205, N184, N57, N181);
or OR2 (N206, N186, N73);
xor XOR2 (N207, N205, N164);
nand NAND2 (N208, N207, N59);
not NOT1 (N209, N202);
or OR2 (N210, N192, N68);
nor NOR2 (N211, N209, N52);
and AND2 (N212, N204, N86);
nor NOR2 (N213, N208, N2);
xor XOR2 (N214, N193, N211);
buf BUF1 (N215, N184);
xor XOR2 (N216, N212, N117);
or OR2 (N217, N173, N206);
nand NAND2 (N218, N207, N201);
or OR2 (N219, N217, N174);
nor NOR4 (N220, N196, N209, N7, N15);
and AND3 (N221, N199, N38, N81);
buf BUF1 (N222, N210);
not NOT1 (N223, N213);
nor NOR4 (N224, N214, N34, N41, N206);
or OR3 (N225, N221, N222, N210);
xor XOR2 (N226, N94, N169);
nor NOR4 (N227, N226, N56, N32, N142);
xor XOR2 (N228, N220, N112);
and AND2 (N229, N215, N225);
not NOT1 (N230, N78);
not NOT1 (N231, N218);
and AND4 (N232, N223, N67, N169, N49);
not NOT1 (N233, N228);
xor XOR2 (N234, N232, N49);
nand NAND4 (N235, N219, N188, N113, N168);
and AND2 (N236, N224, N86);
not NOT1 (N237, N234);
nor NOR2 (N238, N236, N215);
or OR4 (N239, N227, N48, N147, N189);
nor NOR3 (N240, N239, N232, N201);
and AND3 (N241, N235, N57, N113);
not NOT1 (N242, N231);
buf BUF1 (N243, N216);
nor NOR4 (N244, N233, N102, N4, N241);
and AND4 (N245, N91, N154, N227, N33);
nor NOR3 (N246, N242, N109, N60);
nor NOR4 (N247, N243, N234, N114, N115);
or OR3 (N248, N245, N102, N173);
xor XOR2 (N249, N248, N139);
and AND3 (N250, N247, N68, N179);
or OR4 (N251, N203, N193, N61, N191);
xor XOR2 (N252, N240, N73);
buf BUF1 (N253, N230);
nor NOR3 (N254, N244, N231, N75);
not NOT1 (N255, N250);
xor XOR2 (N256, N252, N42);
buf BUF1 (N257, N251);
buf BUF1 (N258, N249);
or OR3 (N259, N257, N91, N173);
nor NOR3 (N260, N238, N36, N183);
or OR3 (N261, N254, N161, N49);
buf BUF1 (N262, N255);
or OR3 (N263, N261, N164, N24);
and AND3 (N264, N259, N88, N55);
buf BUF1 (N265, N262);
nand NAND2 (N266, N258, N218);
nor NOR4 (N267, N263, N227, N220, N81);
or OR3 (N268, N253, N160, N187);
buf BUF1 (N269, N237);
buf BUF1 (N270, N268);
nand NAND2 (N271, N256, N104);
or OR2 (N272, N267, N178);
buf BUF1 (N273, N270);
or OR2 (N274, N269, N91);
and AND2 (N275, N271, N189);
xor XOR2 (N276, N264, N209);
buf BUF1 (N277, N266);
or OR2 (N278, N246, N214);
nand NAND2 (N279, N272, N178);
nor NOR3 (N280, N275, N195, N277);
buf BUF1 (N281, N109);
xor XOR2 (N282, N278, N128);
and AND2 (N283, N281, N158);
or OR2 (N284, N279, N212);
buf BUF1 (N285, N282);
nand NAND4 (N286, N265, N41, N277, N103);
nand NAND3 (N287, N280, N133, N187);
nand NAND4 (N288, N285, N177, N68, N11);
nor NOR2 (N289, N229, N68);
buf BUF1 (N290, N276);
buf BUF1 (N291, N289);
nor NOR2 (N292, N287, N150);
not NOT1 (N293, N284);
buf BUF1 (N294, N286);
and AND2 (N295, N283, N202);
xor XOR2 (N296, N273, N83);
or OR2 (N297, N292, N228);
xor XOR2 (N298, N295, N130);
nor NOR3 (N299, N298, N239, N61);
xor XOR2 (N300, N299, N160);
xor XOR2 (N301, N290, N273);
or OR2 (N302, N274, N275);
nand NAND3 (N303, N288, N237, N252);
or OR2 (N304, N260, N245);
and AND4 (N305, N302, N210, N138, N54);
nor NOR4 (N306, N301, N141, N25, N226);
nand NAND2 (N307, N300, N133);
and AND4 (N308, N303, N22, N205, N28);
buf BUF1 (N309, N305);
or OR3 (N310, N309, N272, N99);
and AND2 (N311, N308, N23);
not NOT1 (N312, N307);
nor NOR3 (N313, N310, N92, N84);
xor XOR2 (N314, N311, N14);
and AND2 (N315, N314, N56);
not NOT1 (N316, N291);
not NOT1 (N317, N293);
xor XOR2 (N318, N296, N33);
nand NAND2 (N319, N306, N98);
or OR4 (N320, N312, N22, N250, N2);
nor NOR3 (N321, N318, N143, N140);
xor XOR2 (N322, N315, N12);
and AND2 (N323, N322, N253);
or OR3 (N324, N319, N32, N269);
xor XOR2 (N325, N323, N13);
xor XOR2 (N326, N324, N138);
buf BUF1 (N327, N326);
nand NAND4 (N328, N294, N227, N139, N69);
xor XOR2 (N329, N297, N90);
or OR3 (N330, N329, N155, N29);
or OR4 (N331, N316, N33, N209, N18);
or OR2 (N332, N327, N271);
buf BUF1 (N333, N321);
nand NAND2 (N334, N332, N58);
buf BUF1 (N335, N317);
not NOT1 (N336, N333);
nor NOR2 (N337, N328, N123);
or OR4 (N338, N337, N75, N20, N297);
xor XOR2 (N339, N335, N152);
and AND4 (N340, N334, N172, N202, N307);
buf BUF1 (N341, N325);
nand NAND2 (N342, N339, N6);
nor NOR2 (N343, N304, N52);
xor XOR2 (N344, N320, N279);
or OR2 (N345, N344, N17);
buf BUF1 (N346, N313);
xor XOR2 (N347, N343, N242);
xor XOR2 (N348, N340, N161);
buf BUF1 (N349, N338);
buf BUF1 (N350, N349);
not NOT1 (N351, N347);
buf BUF1 (N352, N351);
and AND2 (N353, N341, N52);
not NOT1 (N354, N336);
buf BUF1 (N355, N348);
nand NAND4 (N356, N342, N75, N213, N47);
buf BUF1 (N357, N350);
or OR4 (N358, N357, N40, N274, N277);
buf BUF1 (N359, N358);
or OR4 (N360, N352, N357, N139, N295);
xor XOR2 (N361, N355, N64);
nor NOR4 (N362, N345, N357, N62, N103);
nand NAND2 (N363, N354, N211);
not NOT1 (N364, N356);
nor NOR3 (N365, N362, N36, N132);
buf BUF1 (N366, N361);
nand NAND4 (N367, N359, N291, N325, N238);
xor XOR2 (N368, N330, N85);
xor XOR2 (N369, N367, N135);
buf BUF1 (N370, N365);
xor XOR2 (N371, N346, N15);
buf BUF1 (N372, N369);
or OR2 (N373, N370, N77);
not NOT1 (N374, N366);
xor XOR2 (N375, N360, N351);
not NOT1 (N376, N372);
nand NAND3 (N377, N363, N75, N172);
xor XOR2 (N378, N377, N104);
or OR4 (N379, N373, N358, N105, N59);
not NOT1 (N380, N331);
not NOT1 (N381, N378);
xor XOR2 (N382, N381, N335);
not NOT1 (N383, N374);
and AND2 (N384, N382, N8);
not NOT1 (N385, N376);
nand NAND2 (N386, N385, N366);
not NOT1 (N387, N353);
nand NAND2 (N388, N384, N180);
xor XOR2 (N389, N380, N88);
or OR3 (N390, N368, N348, N359);
or OR3 (N391, N364, N92, N339);
nor NOR2 (N392, N389, N243);
not NOT1 (N393, N379);
not NOT1 (N394, N371);
and AND3 (N395, N386, N5, N225);
xor XOR2 (N396, N375, N332);
nor NOR4 (N397, N387, N253, N272, N321);
nor NOR3 (N398, N393, N193, N18);
not NOT1 (N399, N388);
xor XOR2 (N400, N398, N68);
xor XOR2 (N401, N394, N120);
nor NOR3 (N402, N391, N332, N350);
or OR2 (N403, N400, N326);
nand NAND3 (N404, N401, N117, N235);
nor NOR3 (N405, N404, N231, N181);
and AND2 (N406, N405, N188);
nor NOR3 (N407, N406, N386, N20);
nand NAND3 (N408, N383, N260, N209);
nor NOR4 (N409, N407, N347, N32, N366);
and AND2 (N410, N397, N97);
buf BUF1 (N411, N402);
nand NAND4 (N412, N399, N226, N208, N166);
nor NOR4 (N413, N396, N16, N382, N89);
nor NOR4 (N414, N409, N67, N271, N239);
xor XOR2 (N415, N395, N338);
or OR2 (N416, N390, N263);
or OR2 (N417, N411, N158);
nor NOR3 (N418, N392, N209, N416);
xor XOR2 (N419, N246, N239);
nand NAND2 (N420, N410, N121);
nor NOR4 (N421, N403, N225, N26, N137);
nand NAND2 (N422, N421, N22);
nand NAND2 (N423, N417, N194);
xor XOR2 (N424, N422, N216);
not NOT1 (N425, N424);
nand NAND2 (N426, N418, N278);
nor NOR3 (N427, N412, N320, N230);
buf BUF1 (N428, N427);
nor NOR3 (N429, N426, N353, N270);
nor NOR3 (N430, N429, N258, N125);
buf BUF1 (N431, N425);
and AND4 (N432, N419, N276, N50, N133);
not NOT1 (N433, N415);
nand NAND3 (N434, N408, N307, N9);
or OR3 (N435, N434, N329, N293);
or OR2 (N436, N433, N143);
or OR4 (N437, N423, N193, N209, N86);
and AND4 (N438, N420, N264, N199, N62);
or OR2 (N439, N430, N407);
and AND4 (N440, N435, N364, N295, N131);
or OR2 (N441, N440, N257);
or OR4 (N442, N438, N146, N355, N97);
and AND3 (N443, N442, N210, N219);
or OR3 (N444, N428, N143, N430);
not NOT1 (N445, N441);
buf BUF1 (N446, N437);
nor NOR3 (N447, N436, N236, N392);
buf BUF1 (N448, N444);
nor NOR4 (N449, N431, N360, N170, N166);
and AND3 (N450, N445, N416, N367);
nor NOR2 (N451, N450, N314);
nor NOR3 (N452, N443, N111, N345);
xor XOR2 (N453, N452, N301);
and AND2 (N454, N432, N415);
nor NOR2 (N455, N451, N425);
not NOT1 (N456, N454);
nor NOR2 (N457, N439, N20);
not NOT1 (N458, N457);
nand NAND4 (N459, N447, N425, N247, N229);
and AND2 (N460, N453, N135);
or OR2 (N461, N456, N130);
nor NOR4 (N462, N458, N1, N401, N311);
nor NOR4 (N463, N414, N376, N161, N320);
nor NOR3 (N464, N461, N91, N188);
nor NOR3 (N465, N463, N296, N383);
and AND4 (N466, N459, N204, N182, N448);
not NOT1 (N467, N380);
xor XOR2 (N468, N464, N55);
not NOT1 (N469, N466);
buf BUF1 (N470, N462);
nand NAND3 (N471, N469, N81, N32);
or OR3 (N472, N470, N109, N469);
nand NAND4 (N473, N449, N331, N382, N104);
nand NAND2 (N474, N471, N38);
and AND2 (N475, N413, N361);
not NOT1 (N476, N446);
not NOT1 (N477, N465);
buf BUF1 (N478, N460);
or OR4 (N479, N475, N371, N316, N379);
or OR4 (N480, N477, N269, N183, N327);
xor XOR2 (N481, N467, N209);
nor NOR3 (N482, N476, N435, N308);
not NOT1 (N483, N468);
and AND3 (N484, N481, N298, N176);
not NOT1 (N485, N482);
buf BUF1 (N486, N478);
or OR2 (N487, N455, N341);
xor XOR2 (N488, N483, N36);
xor XOR2 (N489, N472, N433);
buf BUF1 (N490, N479);
buf BUF1 (N491, N490);
nor NOR3 (N492, N486, N11, N7);
xor XOR2 (N493, N485, N426);
not NOT1 (N494, N489);
not NOT1 (N495, N474);
not NOT1 (N496, N487);
nand NAND3 (N497, N494, N352, N193);
xor XOR2 (N498, N497, N100);
buf BUF1 (N499, N480);
not NOT1 (N500, N492);
buf BUF1 (N501, N491);
not NOT1 (N502, N493);
not NOT1 (N503, N499);
not NOT1 (N504, N495);
or OR3 (N505, N473, N403, N144);
xor XOR2 (N506, N505, N102);
not NOT1 (N507, N498);
xor XOR2 (N508, N502, N186);
nand NAND4 (N509, N488, N226, N493, N211);
nor NOR2 (N510, N508, N326);
buf BUF1 (N511, N496);
nand NAND3 (N512, N503, N277, N424);
buf BUF1 (N513, N500);
nand NAND3 (N514, N484, N247, N50);
and AND3 (N515, N513, N416, N141);
xor XOR2 (N516, N515, N476);
not NOT1 (N517, N501);
nand NAND4 (N518, N516, N27, N158, N39);
and AND3 (N519, N518, N278, N331);
and AND2 (N520, N519, N4);
buf BUF1 (N521, N517);
not NOT1 (N522, N520);
xor XOR2 (N523, N510, N393);
nor NOR3 (N524, N511, N18, N134);
xor XOR2 (N525, N522, N499);
nand NAND2 (N526, N521, N330);
buf BUF1 (N527, N504);
nor NOR4 (N528, N509, N41, N487, N506);
nor NOR2 (N529, N384, N433);
nor NOR3 (N530, N529, N392, N312);
and AND2 (N531, N528, N226);
xor XOR2 (N532, N527, N272);
nand NAND3 (N533, N531, N439, N61);
xor XOR2 (N534, N526, N398);
nor NOR2 (N535, N523, N103);
buf BUF1 (N536, N512);
nand NAND4 (N537, N525, N494, N407, N451);
not NOT1 (N538, N530);
not NOT1 (N539, N534);
buf BUF1 (N540, N524);
nand NAND3 (N541, N532, N238, N536);
nor NOR3 (N542, N497, N504, N126);
nand NAND2 (N543, N542, N540);
buf BUF1 (N544, N418);
not NOT1 (N545, N537);
nor NOR2 (N546, N541, N365);
buf BUF1 (N547, N533);
nand NAND2 (N548, N545, N167);
nor NOR2 (N549, N543, N487);
not NOT1 (N550, N549);
and AND2 (N551, N514, N53);
and AND3 (N552, N550, N308, N112);
and AND3 (N553, N538, N66, N372);
xor XOR2 (N554, N507, N306);
nand NAND3 (N555, N551, N216, N387);
nand NAND4 (N556, N553, N211, N546, N17);
not NOT1 (N557, N60);
nor NOR3 (N558, N535, N402, N8);
xor XOR2 (N559, N548, N417);
or OR4 (N560, N552, N288, N30, N448);
nor NOR3 (N561, N555, N378, N16);
or OR4 (N562, N547, N84, N249, N91);
buf BUF1 (N563, N561);
or OR3 (N564, N544, N180, N438);
xor XOR2 (N565, N557, N71);
nand NAND3 (N566, N565, N288, N143);
nand NAND2 (N567, N560, N120);
xor XOR2 (N568, N562, N8);
xor XOR2 (N569, N567, N264);
not NOT1 (N570, N556);
xor XOR2 (N571, N563, N38);
and AND2 (N572, N571, N548);
and AND2 (N573, N569, N327);
buf BUF1 (N574, N568);
not NOT1 (N575, N574);
nor NOR4 (N576, N539, N356, N25, N135);
nand NAND4 (N577, N573, N417, N289, N90);
nand NAND4 (N578, N558, N207, N527, N193);
nor NOR2 (N579, N575, N240);
xor XOR2 (N580, N566, N444);
or OR4 (N581, N554, N62, N541, N366);
buf BUF1 (N582, N564);
buf BUF1 (N583, N581);
or OR4 (N584, N570, N427, N344, N313);
not NOT1 (N585, N584);
or OR4 (N586, N583, N341, N7, N223);
xor XOR2 (N587, N576, N57);
and AND4 (N588, N579, N487, N541, N462);
nor NOR4 (N589, N582, N206, N196, N247);
xor XOR2 (N590, N578, N204);
xor XOR2 (N591, N572, N287);
not NOT1 (N592, N580);
buf BUF1 (N593, N585);
nand NAND3 (N594, N593, N185, N427);
nor NOR3 (N595, N591, N292, N507);
and AND3 (N596, N587, N343, N375);
or OR4 (N597, N586, N180, N168, N533);
or OR2 (N598, N592, N227);
nand NAND4 (N599, N590, N119, N539, N139);
xor XOR2 (N600, N598, N115);
nand NAND4 (N601, N596, N121, N556, N411);
or OR2 (N602, N597, N163);
xor XOR2 (N603, N577, N130);
or OR3 (N604, N559, N472, N456);
nor NOR3 (N605, N595, N430, N469);
xor XOR2 (N606, N604, N105);
not NOT1 (N607, N606);
buf BUF1 (N608, N599);
nor NOR4 (N609, N594, N605, N570, N367);
nor NOR4 (N610, N24, N563, N294, N294);
xor XOR2 (N611, N600, N447);
buf BUF1 (N612, N610);
not NOT1 (N613, N609);
buf BUF1 (N614, N603);
or OR4 (N615, N608, N559, N192, N108);
nor NOR2 (N616, N589, N541);
and AND2 (N617, N613, N565);
nor NOR2 (N618, N612, N308);
and AND3 (N619, N615, N343, N227);
xor XOR2 (N620, N616, N269);
or OR4 (N621, N588, N160, N94, N598);
nor NOR2 (N622, N601, N122);
nor NOR3 (N623, N618, N106, N422);
not NOT1 (N624, N621);
endmodule