// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N1619,N1611,N1596,N1615,N1618,N1616,N1604,N1602,N1620,N1622;

not NOT1 (N23, N8);
buf BUF1 (N24, N21);
nand NAND2 (N25, N6, N17);
and AND3 (N26, N20, N21, N13);
buf BUF1 (N27, N14);
not NOT1 (N28, N23);
or OR3 (N29, N27, N15, N22);
nor NOR3 (N30, N13, N24, N25);
or OR2 (N31, N17, N30);
not NOT1 (N32, N16);
and AND3 (N33, N30, N24, N9);
and AND4 (N34, N28, N31, N24, N29);
not NOT1 (N35, N12);
or OR4 (N36, N21, N8, N26, N4);
and AND2 (N37, N8, N11);
not NOT1 (N38, N9);
nand NAND4 (N39, N29, N31, N35, N1);
or OR4 (N40, N15, N10, N31, N38);
and AND4 (N41, N30, N22, N30, N19);
not NOT1 (N42, N31);
nand NAND4 (N43, N38, N16, N39, N11);
and AND3 (N44, N16, N27, N40);
or OR4 (N45, N38, N25, N11, N6);
xor XOR2 (N46, N33, N36);
nand NAND3 (N47, N34, N46, N46);
or OR3 (N48, N34, N5, N15);
nor NOR2 (N49, N30, N35);
or OR2 (N50, N41, N42);
or OR3 (N51, N49, N8, N32);
and AND2 (N52, N19, N20);
and AND3 (N53, N10, N39, N8);
not NOT1 (N54, N53);
buf BUF1 (N55, N47);
buf BUF1 (N56, N55);
or OR3 (N57, N50, N25, N9);
not NOT1 (N58, N54);
xor XOR2 (N59, N48, N1);
nand NAND3 (N60, N45, N19, N9);
not NOT1 (N61, N57);
nand NAND4 (N62, N44, N26, N25, N40);
or OR4 (N63, N58, N57, N10, N33);
buf BUF1 (N64, N52);
or OR4 (N65, N64, N52, N49, N18);
buf BUF1 (N66, N62);
not NOT1 (N67, N51);
nand NAND3 (N68, N60, N35, N23);
not NOT1 (N69, N66);
nand NAND3 (N70, N37, N50, N37);
and AND3 (N71, N69, N35, N25);
xor XOR2 (N72, N61, N67);
nand NAND2 (N73, N69, N63);
buf BUF1 (N74, N63);
or OR3 (N75, N70, N68, N64);
buf BUF1 (N76, N8);
not NOT1 (N77, N72);
and AND4 (N78, N73, N71, N22, N64);
buf BUF1 (N79, N50);
and AND3 (N80, N59, N39, N37);
xor XOR2 (N81, N65, N37);
not NOT1 (N82, N56);
nor NOR4 (N83, N79, N40, N62, N60);
or OR4 (N84, N78, N25, N41, N75);
nand NAND3 (N85, N30, N24, N56);
and AND3 (N86, N85, N10, N63);
nor NOR3 (N87, N83, N13, N53);
not NOT1 (N88, N84);
or OR4 (N89, N43, N35, N15, N18);
nor NOR3 (N90, N87, N64, N16);
or OR3 (N91, N81, N45, N50);
and AND3 (N92, N91, N42, N24);
xor XOR2 (N93, N88, N52);
not NOT1 (N94, N80);
not NOT1 (N95, N94);
or OR2 (N96, N74, N89);
and AND2 (N97, N43, N91);
nor NOR2 (N98, N82, N75);
nand NAND3 (N99, N90, N81, N72);
not NOT1 (N100, N96);
buf BUF1 (N101, N92);
xor XOR2 (N102, N77, N53);
buf BUF1 (N103, N76);
buf BUF1 (N104, N102);
and AND3 (N105, N93, N13, N37);
or OR2 (N106, N86, N34);
nor NOR3 (N107, N101, N68, N44);
xor XOR2 (N108, N97, N63);
and AND3 (N109, N98, N108, N3);
or OR3 (N110, N17, N77, N18);
and AND2 (N111, N107, N48);
nor NOR3 (N112, N106, N103, N71);
xor XOR2 (N113, N87, N105);
and AND3 (N114, N26, N6, N103);
not NOT1 (N115, N113);
not NOT1 (N116, N112);
or OR2 (N117, N109, N104);
xor XOR2 (N118, N41, N1);
xor XOR2 (N119, N100, N106);
buf BUF1 (N120, N116);
nand NAND4 (N121, N117, N110, N116, N93);
or OR3 (N122, N8, N77, N118);
and AND3 (N123, N97, N118, N9);
nand NAND2 (N124, N111, N2);
buf BUF1 (N125, N122);
or OR2 (N126, N120, N89);
buf BUF1 (N127, N121);
not NOT1 (N128, N99);
not NOT1 (N129, N115);
nor NOR4 (N130, N128, N22, N99, N5);
or OR2 (N131, N130, N108);
and AND2 (N132, N131, N50);
nand NAND3 (N133, N114, N99, N85);
and AND2 (N134, N119, N51);
nor NOR3 (N135, N95, N38, N60);
and AND3 (N136, N127, N64, N52);
nor NOR2 (N137, N125, N88);
nand NAND4 (N138, N133, N30, N84, N11);
xor XOR2 (N139, N138, N8);
nand NAND4 (N140, N134, N107, N27, N84);
xor XOR2 (N141, N132, N93);
or OR4 (N142, N136, N113, N81, N96);
xor XOR2 (N143, N139, N125);
nand NAND3 (N144, N143, N133, N97);
not NOT1 (N145, N123);
xor XOR2 (N146, N141, N65);
not NOT1 (N147, N145);
not NOT1 (N148, N137);
not NOT1 (N149, N124);
xor XOR2 (N150, N126, N141);
xor XOR2 (N151, N150, N3);
and AND4 (N152, N129, N100, N28, N65);
buf BUF1 (N153, N146);
or OR2 (N154, N147, N55);
buf BUF1 (N155, N152);
buf BUF1 (N156, N140);
nand NAND2 (N157, N142, N37);
not NOT1 (N158, N154);
nand NAND4 (N159, N156, N44, N115, N118);
not NOT1 (N160, N148);
or OR3 (N161, N153, N135, N90);
or OR4 (N162, N137, N47, N110, N90);
nand NAND2 (N163, N151, N8);
nand NAND2 (N164, N163, N8);
xor XOR2 (N165, N161, N121);
buf BUF1 (N166, N165);
buf BUF1 (N167, N144);
or OR3 (N168, N157, N148, N86);
or OR3 (N169, N149, N94, N149);
buf BUF1 (N170, N159);
xor XOR2 (N171, N168, N34);
nor NOR2 (N172, N169, N35);
or OR3 (N173, N171, N132, N42);
nand NAND2 (N174, N173, N138);
nor NOR4 (N175, N164, N46, N85, N85);
nand NAND3 (N176, N172, N70, N89);
not NOT1 (N177, N160);
buf BUF1 (N178, N166);
xor XOR2 (N179, N176, N3);
or OR2 (N180, N162, N170);
xor XOR2 (N181, N32, N171);
or OR2 (N182, N167, N16);
not NOT1 (N183, N182);
not NOT1 (N184, N183);
and AND4 (N185, N180, N86, N55, N69);
nor NOR4 (N186, N155, N31, N106, N98);
or OR3 (N187, N174, N53, N146);
and AND4 (N188, N185, N187, N10, N63);
xor XOR2 (N189, N53, N92);
buf BUF1 (N190, N175);
nor NOR2 (N191, N186, N71);
and AND3 (N192, N181, N3, N40);
xor XOR2 (N193, N177, N97);
and AND3 (N194, N191, N175, N125);
and AND3 (N195, N190, N39, N32);
nor NOR3 (N196, N158, N187, N36);
nand NAND4 (N197, N192, N188, N149, N58);
buf BUF1 (N198, N121);
xor XOR2 (N199, N195, N145);
nand NAND3 (N200, N198, N72, N12);
nand NAND3 (N201, N194, N25, N39);
nor NOR4 (N202, N199, N2, N181, N119);
not NOT1 (N203, N197);
buf BUF1 (N204, N184);
xor XOR2 (N205, N189, N29);
buf BUF1 (N206, N179);
or OR3 (N207, N202, N15, N92);
nor NOR4 (N208, N193, N173, N3, N115);
buf BUF1 (N209, N205);
xor XOR2 (N210, N196, N120);
buf BUF1 (N211, N208);
nor NOR2 (N212, N210, N164);
buf BUF1 (N213, N211);
or OR3 (N214, N203, N137, N14);
or OR3 (N215, N178, N156, N160);
or OR3 (N216, N214, N162, N204);
buf BUF1 (N217, N24);
xor XOR2 (N218, N201, N205);
nor NOR4 (N219, N215, N180, N123, N34);
or OR2 (N220, N219, N189);
xor XOR2 (N221, N218, N165);
not NOT1 (N222, N220);
buf BUF1 (N223, N213);
buf BUF1 (N224, N209);
and AND2 (N225, N221, N161);
not NOT1 (N226, N207);
nand NAND3 (N227, N200, N179, N48);
not NOT1 (N228, N217);
nor NOR3 (N229, N206, N106, N24);
xor XOR2 (N230, N223, N32);
and AND2 (N231, N224, N136);
not NOT1 (N232, N222);
or OR4 (N233, N226, N214, N224, N66);
nor NOR2 (N234, N231, N205);
xor XOR2 (N235, N225, N140);
xor XOR2 (N236, N227, N3);
nor NOR4 (N237, N233, N167, N3, N167);
nor NOR3 (N238, N230, N117, N224);
not NOT1 (N239, N237);
not NOT1 (N240, N236);
nor NOR4 (N241, N228, N125, N16, N97);
nor NOR2 (N242, N235, N238);
and AND3 (N243, N204, N115, N122);
or OR2 (N244, N234, N125);
xor XOR2 (N245, N243, N129);
or OR3 (N246, N239, N185, N209);
and AND3 (N247, N245, N207, N170);
nor NOR2 (N248, N241, N119);
buf BUF1 (N249, N240);
nand NAND3 (N250, N248, N199, N220);
xor XOR2 (N251, N232, N147);
nand NAND4 (N252, N250, N133, N175, N238);
and AND3 (N253, N242, N139, N115);
buf BUF1 (N254, N246);
or OR2 (N255, N244, N232);
and AND4 (N256, N255, N131, N203, N78);
or OR4 (N257, N249, N153, N106, N158);
xor XOR2 (N258, N254, N4);
nand NAND2 (N259, N257, N122);
nor NOR3 (N260, N247, N47, N101);
xor XOR2 (N261, N251, N212);
or OR2 (N262, N134, N80);
or OR4 (N263, N259, N99, N203, N214);
nand NAND3 (N264, N216, N54, N169);
not NOT1 (N265, N253);
or OR4 (N266, N265, N244, N81, N264);
not NOT1 (N267, N58);
xor XOR2 (N268, N256, N19);
xor XOR2 (N269, N260, N172);
and AND3 (N270, N263, N100, N204);
nor NOR3 (N271, N266, N96, N58);
buf BUF1 (N272, N269);
nor NOR3 (N273, N258, N229, N252);
xor XOR2 (N274, N22, N174);
nand NAND2 (N275, N34, N129);
not NOT1 (N276, N270);
or OR4 (N277, N273, N87, N206, N231);
nor NOR3 (N278, N261, N4, N130);
nor NOR3 (N279, N267, N144, N213);
not NOT1 (N280, N271);
xor XOR2 (N281, N278, N267);
and AND4 (N282, N281, N76, N89, N45);
and AND2 (N283, N276, N45);
and AND3 (N284, N262, N60, N235);
buf BUF1 (N285, N279);
and AND2 (N286, N283, N284);
nand NAND2 (N287, N63, N113);
not NOT1 (N288, N268);
xor XOR2 (N289, N275, N211);
or OR4 (N290, N289, N266, N7, N69);
not NOT1 (N291, N285);
nor NOR4 (N292, N290, N274, N103, N1);
xor XOR2 (N293, N79, N141);
buf BUF1 (N294, N282);
buf BUF1 (N295, N292);
not NOT1 (N296, N288);
buf BUF1 (N297, N280);
not NOT1 (N298, N287);
nand NAND4 (N299, N294, N166, N13, N150);
not NOT1 (N300, N293);
or OR2 (N301, N300, N150);
and AND3 (N302, N291, N172, N161);
nor NOR3 (N303, N277, N254, N195);
nand NAND3 (N304, N286, N240, N292);
not NOT1 (N305, N295);
not NOT1 (N306, N301);
or OR3 (N307, N296, N206, N41);
nand NAND2 (N308, N307, N197);
not NOT1 (N309, N272);
and AND2 (N310, N299, N211);
xor XOR2 (N311, N304, N268);
nand NAND4 (N312, N311, N168, N75, N45);
or OR4 (N313, N312, N95, N295, N188);
and AND3 (N314, N313, N173, N285);
xor XOR2 (N315, N305, N55);
and AND3 (N316, N303, N64, N62);
nor NOR2 (N317, N302, N1);
nor NOR3 (N318, N306, N55, N253);
and AND4 (N319, N297, N41, N30, N184);
xor XOR2 (N320, N317, N293);
nor NOR4 (N321, N320, N11, N9, N232);
buf BUF1 (N322, N316);
buf BUF1 (N323, N298);
not NOT1 (N324, N323);
not NOT1 (N325, N310);
or OR3 (N326, N308, N121, N303);
xor XOR2 (N327, N315, N276);
xor XOR2 (N328, N322, N215);
and AND4 (N329, N314, N39, N21, N173);
and AND4 (N330, N329, N232, N270, N16);
nor NOR4 (N331, N319, N269, N167, N169);
and AND3 (N332, N324, N167, N17);
or OR2 (N333, N318, N76);
nor NOR3 (N334, N327, N194, N226);
or OR2 (N335, N331, N24);
nand NAND3 (N336, N335, N157, N176);
or OR2 (N337, N334, N201);
and AND4 (N338, N326, N277, N205, N59);
buf BUF1 (N339, N321);
nand NAND3 (N340, N333, N15, N256);
xor XOR2 (N341, N337, N238);
buf BUF1 (N342, N341);
and AND3 (N343, N342, N231, N53);
buf BUF1 (N344, N338);
xor XOR2 (N345, N325, N44);
not NOT1 (N346, N340);
not NOT1 (N347, N343);
or OR4 (N348, N346, N313, N258, N72);
nand NAND3 (N349, N332, N204, N14);
xor XOR2 (N350, N347, N303);
nor NOR2 (N351, N309, N206);
xor XOR2 (N352, N349, N314);
xor XOR2 (N353, N336, N64);
xor XOR2 (N354, N351, N334);
nand NAND2 (N355, N348, N130);
nand NAND4 (N356, N353, N198, N36, N175);
not NOT1 (N357, N352);
and AND2 (N358, N354, N321);
and AND2 (N359, N344, N107);
xor XOR2 (N360, N350, N236);
nand NAND4 (N361, N328, N59, N95, N323);
and AND2 (N362, N356, N155);
and AND2 (N363, N358, N113);
nor NOR4 (N364, N357, N298, N301, N342);
xor XOR2 (N365, N359, N354);
not NOT1 (N366, N363);
not NOT1 (N367, N360);
nor NOR3 (N368, N367, N157, N119);
nor NOR2 (N369, N362, N157);
nand NAND2 (N370, N368, N203);
not NOT1 (N371, N345);
xor XOR2 (N372, N330, N151);
or OR4 (N373, N365, N344, N154, N23);
not NOT1 (N374, N366);
or OR2 (N375, N364, N3);
or OR2 (N376, N369, N306);
nand NAND3 (N377, N374, N329, N241);
buf BUF1 (N378, N377);
nand NAND4 (N379, N376, N89, N205, N25);
nand NAND3 (N380, N371, N93, N337);
nor NOR4 (N381, N370, N305, N84, N307);
xor XOR2 (N382, N339, N246);
buf BUF1 (N383, N380);
buf BUF1 (N384, N373);
not NOT1 (N385, N384);
nand NAND2 (N386, N355, N353);
and AND2 (N387, N375, N311);
buf BUF1 (N388, N361);
buf BUF1 (N389, N381);
not NOT1 (N390, N387);
nand NAND3 (N391, N388, N24, N344);
and AND2 (N392, N383, N23);
and AND3 (N393, N391, N186, N97);
nor NOR4 (N394, N389, N156, N141, N349);
buf BUF1 (N395, N386);
nand NAND3 (N396, N395, N22, N348);
nor NOR2 (N397, N385, N86);
or OR3 (N398, N372, N304, N300);
xor XOR2 (N399, N394, N196);
nor NOR3 (N400, N392, N330, N349);
buf BUF1 (N401, N378);
xor XOR2 (N402, N398, N312);
buf BUF1 (N403, N401);
or OR3 (N404, N393, N142, N324);
nor NOR2 (N405, N379, N140);
and AND4 (N406, N403, N322, N93, N289);
or OR2 (N407, N390, N29);
not NOT1 (N408, N407);
xor XOR2 (N409, N399, N355);
buf BUF1 (N410, N404);
xor XOR2 (N411, N410, N31);
or OR3 (N412, N397, N406, N67);
and AND3 (N413, N293, N205, N271);
xor XOR2 (N414, N402, N104);
or OR2 (N415, N382, N142);
or OR4 (N416, N400, N2, N161, N328);
xor XOR2 (N417, N413, N261);
not NOT1 (N418, N405);
and AND3 (N419, N414, N386, N75);
not NOT1 (N420, N411);
not NOT1 (N421, N419);
nor NOR4 (N422, N408, N357, N136, N124);
nand NAND3 (N423, N416, N322, N222);
xor XOR2 (N424, N423, N402);
xor XOR2 (N425, N396, N192);
and AND4 (N426, N421, N272, N139, N16);
not NOT1 (N427, N420);
nor NOR2 (N428, N418, N62);
nand NAND3 (N429, N425, N340, N205);
or OR4 (N430, N412, N284, N188, N296);
nand NAND3 (N431, N429, N411, N198);
buf BUF1 (N432, N415);
nor NOR3 (N433, N417, N292, N9);
nor NOR3 (N434, N427, N186, N248);
nand NAND2 (N435, N432, N416);
not NOT1 (N436, N422);
buf BUF1 (N437, N431);
not NOT1 (N438, N428);
nand NAND2 (N439, N438, N435);
buf BUF1 (N440, N80);
nor NOR2 (N441, N437, N235);
nand NAND4 (N442, N436, N434, N129, N348);
and AND3 (N443, N221, N390, N328);
or OR4 (N444, N430, N22, N335, N139);
xor XOR2 (N445, N442, N230);
or OR2 (N446, N439, N410);
xor XOR2 (N447, N441, N2);
nand NAND2 (N448, N444, N215);
and AND3 (N449, N447, N176, N145);
nor NOR3 (N450, N448, N407, N317);
and AND4 (N451, N443, N64, N305, N409);
or OR4 (N452, N306, N186, N93, N412);
and AND3 (N453, N449, N129, N313);
nand NAND3 (N454, N433, N262, N342);
xor XOR2 (N455, N446, N28);
or OR3 (N456, N455, N61, N355);
or OR2 (N457, N426, N437);
nor NOR4 (N458, N454, N25, N237, N16);
buf BUF1 (N459, N450);
nor NOR4 (N460, N424, N102, N79, N13);
xor XOR2 (N461, N460, N137);
nor NOR3 (N462, N452, N205, N63);
nand NAND3 (N463, N440, N167, N68);
buf BUF1 (N464, N456);
and AND2 (N465, N459, N193);
xor XOR2 (N466, N461, N106);
or OR2 (N467, N451, N44);
or OR2 (N468, N457, N261);
xor XOR2 (N469, N463, N388);
not NOT1 (N470, N464);
buf BUF1 (N471, N467);
and AND4 (N472, N470, N435, N218, N429);
xor XOR2 (N473, N469, N10);
nor NOR4 (N474, N453, N234, N229, N263);
and AND3 (N475, N473, N65, N435);
xor XOR2 (N476, N471, N370);
nor NOR2 (N477, N462, N115);
not NOT1 (N478, N476);
xor XOR2 (N479, N478, N33);
or OR4 (N480, N475, N261, N39, N121);
nor NOR3 (N481, N458, N374, N388);
and AND3 (N482, N472, N172, N251);
and AND2 (N483, N466, N399);
and AND4 (N484, N481, N115, N157, N354);
or OR3 (N485, N468, N309, N458);
not NOT1 (N486, N445);
not NOT1 (N487, N480);
nor NOR4 (N488, N479, N251, N397, N180);
xor XOR2 (N489, N485, N216);
nand NAND3 (N490, N484, N62, N241);
nor NOR4 (N491, N482, N32, N454, N289);
or OR4 (N492, N487, N167, N447, N177);
nand NAND4 (N493, N488, N189, N389, N57);
not NOT1 (N494, N493);
and AND4 (N495, N465, N322, N54, N342);
or OR2 (N496, N483, N303);
nand NAND3 (N497, N491, N313, N376);
not NOT1 (N498, N496);
or OR2 (N499, N498, N495);
and AND3 (N500, N261, N23, N316);
xor XOR2 (N501, N492, N114);
nor NOR4 (N502, N500, N252, N362, N150);
nand NAND2 (N503, N501, N487);
buf BUF1 (N504, N503);
xor XOR2 (N505, N504, N180);
nand NAND2 (N506, N490, N476);
and AND4 (N507, N494, N373, N244, N240);
nand NAND4 (N508, N505, N81, N93, N315);
nor NOR3 (N509, N497, N502, N29);
or OR2 (N510, N18, N164);
nand NAND4 (N511, N510, N262, N456, N132);
nand NAND3 (N512, N511, N427, N235);
or OR2 (N513, N486, N369);
not NOT1 (N514, N509);
or OR3 (N515, N474, N111, N487);
nor NOR4 (N516, N489, N41, N275, N205);
buf BUF1 (N517, N513);
or OR2 (N518, N508, N302);
nor NOR2 (N519, N516, N246);
buf BUF1 (N520, N515);
nor NOR2 (N521, N512, N255);
buf BUF1 (N522, N518);
nand NAND3 (N523, N517, N22, N413);
buf BUF1 (N524, N506);
not NOT1 (N525, N524);
nand NAND2 (N526, N525, N446);
nor NOR3 (N527, N477, N471, N494);
buf BUF1 (N528, N523);
nand NAND4 (N529, N527, N280, N247, N70);
and AND4 (N530, N520, N273, N304, N128);
nand NAND4 (N531, N522, N57, N235, N501);
buf BUF1 (N532, N514);
nor NOR3 (N533, N528, N348, N523);
nor NOR2 (N534, N507, N98);
or OR4 (N535, N521, N76, N365, N471);
not NOT1 (N536, N533);
buf BUF1 (N537, N531);
not NOT1 (N538, N499);
and AND4 (N539, N536, N31, N133, N353);
nor NOR4 (N540, N535, N423, N462, N57);
xor XOR2 (N541, N530, N269);
xor XOR2 (N542, N537, N298);
not NOT1 (N543, N534);
xor XOR2 (N544, N519, N276);
and AND3 (N545, N538, N460, N241);
and AND3 (N546, N532, N289, N333);
nor NOR3 (N547, N543, N356, N386);
nor NOR4 (N548, N526, N174, N354, N530);
nand NAND2 (N549, N529, N131);
nor NOR3 (N550, N541, N2, N159);
nor NOR4 (N551, N539, N59, N365, N50);
not NOT1 (N552, N547);
or OR4 (N553, N545, N454, N476, N92);
nor NOR2 (N554, N552, N142);
xor XOR2 (N555, N548, N246);
and AND3 (N556, N540, N361, N453);
not NOT1 (N557, N554);
nor NOR2 (N558, N553, N103);
nand NAND3 (N559, N550, N531, N72);
and AND4 (N560, N544, N212, N211, N262);
nor NOR4 (N561, N542, N450, N14, N2);
buf BUF1 (N562, N560);
or OR3 (N563, N549, N409, N187);
buf BUF1 (N564, N557);
buf BUF1 (N565, N562);
or OR3 (N566, N564, N403, N72);
or OR2 (N567, N559, N176);
nand NAND4 (N568, N561, N179, N114, N365);
buf BUF1 (N569, N567);
not NOT1 (N570, N546);
or OR3 (N571, N565, N342, N11);
xor XOR2 (N572, N556, N239);
nand NAND2 (N573, N558, N496);
xor XOR2 (N574, N551, N243);
buf BUF1 (N575, N563);
buf BUF1 (N576, N568);
xor XOR2 (N577, N570, N468);
or OR3 (N578, N566, N263, N247);
nor NOR3 (N579, N578, N325, N229);
nor NOR3 (N580, N575, N254, N175);
xor XOR2 (N581, N576, N551);
or OR2 (N582, N572, N213);
nand NAND4 (N583, N577, N474, N389, N173);
xor XOR2 (N584, N571, N506);
not NOT1 (N585, N584);
and AND3 (N586, N574, N130, N344);
or OR4 (N587, N582, N259, N78, N348);
or OR2 (N588, N585, N167);
and AND4 (N589, N580, N67, N171, N178);
nand NAND2 (N590, N555, N16);
nand NAND2 (N591, N587, N354);
buf BUF1 (N592, N589);
or OR2 (N593, N579, N242);
and AND2 (N594, N593, N574);
nand NAND4 (N595, N573, N83, N504, N135);
nor NOR4 (N596, N595, N167, N12, N358);
buf BUF1 (N597, N569);
nand NAND4 (N598, N594, N257, N180, N518);
xor XOR2 (N599, N596, N267);
not NOT1 (N600, N592);
and AND3 (N601, N598, N212, N67);
not NOT1 (N602, N588);
xor XOR2 (N603, N586, N227);
or OR4 (N604, N583, N43, N535, N593);
and AND4 (N605, N590, N262, N346, N138);
nor NOR3 (N606, N597, N146, N168);
buf BUF1 (N607, N581);
nand NAND2 (N608, N602, N254);
and AND4 (N609, N605, N248, N97, N118);
not NOT1 (N610, N591);
nand NAND3 (N611, N600, N27, N117);
and AND3 (N612, N608, N183, N508);
xor XOR2 (N613, N601, N516);
xor XOR2 (N614, N599, N84);
xor XOR2 (N615, N614, N538);
or OR3 (N616, N609, N270, N91);
nor NOR3 (N617, N611, N405, N385);
nand NAND3 (N618, N615, N436, N605);
buf BUF1 (N619, N607);
buf BUF1 (N620, N616);
not NOT1 (N621, N620);
xor XOR2 (N622, N610, N75);
nand NAND4 (N623, N603, N226, N451, N545);
nor NOR3 (N624, N618, N134, N578);
not NOT1 (N625, N621);
not NOT1 (N626, N625);
nand NAND3 (N627, N606, N504, N119);
or OR4 (N628, N604, N370, N301, N504);
xor XOR2 (N629, N623, N65);
nand NAND2 (N630, N617, N132);
and AND2 (N631, N626, N62);
nand NAND3 (N632, N628, N108, N212);
xor XOR2 (N633, N629, N183);
buf BUF1 (N634, N627);
and AND4 (N635, N619, N619, N58, N284);
nand NAND3 (N636, N613, N101, N418);
and AND3 (N637, N624, N150, N91);
or OR2 (N638, N622, N471);
or OR2 (N639, N635, N118);
xor XOR2 (N640, N637, N239);
nand NAND3 (N641, N631, N389, N415);
nand NAND3 (N642, N632, N552, N531);
nor NOR2 (N643, N636, N564);
nand NAND4 (N644, N634, N589, N79, N153);
buf BUF1 (N645, N643);
buf BUF1 (N646, N642);
or OR2 (N647, N640, N391);
not NOT1 (N648, N612);
or OR3 (N649, N641, N280, N246);
and AND4 (N650, N647, N66, N68, N599);
not NOT1 (N651, N648);
nand NAND3 (N652, N630, N84, N359);
not NOT1 (N653, N633);
and AND2 (N654, N649, N155);
not NOT1 (N655, N653);
xor XOR2 (N656, N655, N598);
nand NAND3 (N657, N650, N421, N631);
xor XOR2 (N658, N651, N358);
nand NAND4 (N659, N646, N101, N310, N552);
not NOT1 (N660, N645);
nand NAND3 (N661, N654, N595, N592);
and AND2 (N662, N656, N212);
buf BUF1 (N663, N657);
or OR3 (N664, N660, N14, N440);
or OR4 (N665, N639, N452, N146, N500);
nor NOR2 (N666, N658, N365);
xor XOR2 (N667, N644, N437);
not NOT1 (N668, N659);
xor XOR2 (N669, N652, N197);
not NOT1 (N670, N665);
not NOT1 (N671, N664);
buf BUF1 (N672, N666);
not NOT1 (N673, N661);
and AND3 (N674, N638, N535, N257);
nor NOR2 (N675, N672, N99);
xor XOR2 (N676, N671, N458);
not NOT1 (N677, N676);
or OR4 (N678, N677, N48, N447, N434);
xor XOR2 (N679, N662, N322);
and AND2 (N680, N673, N528);
or OR2 (N681, N680, N320);
not NOT1 (N682, N681);
and AND2 (N683, N668, N170);
not NOT1 (N684, N669);
or OR4 (N685, N667, N462, N369, N570);
nand NAND4 (N686, N670, N503, N252, N327);
nand NAND2 (N687, N663, N221);
not NOT1 (N688, N675);
xor XOR2 (N689, N686, N230);
nand NAND2 (N690, N687, N521);
not NOT1 (N691, N674);
xor XOR2 (N692, N684, N448);
buf BUF1 (N693, N690);
buf BUF1 (N694, N693);
buf BUF1 (N695, N694);
not NOT1 (N696, N689);
xor XOR2 (N697, N679, N123);
buf BUF1 (N698, N688);
buf BUF1 (N699, N697);
not NOT1 (N700, N695);
or OR3 (N701, N691, N488, N493);
nand NAND3 (N702, N701, N273, N625);
or OR3 (N703, N700, N614, N93);
nor NOR2 (N704, N678, N75);
nand NAND3 (N705, N685, N69, N268);
nor NOR4 (N706, N683, N372, N160, N259);
and AND3 (N707, N682, N129, N118);
not NOT1 (N708, N702);
xor XOR2 (N709, N696, N126);
or OR4 (N710, N707, N57, N413, N371);
nor NOR3 (N711, N710, N573, N13);
and AND3 (N712, N711, N377, N108);
nor NOR3 (N713, N698, N248, N385);
not NOT1 (N714, N704);
buf BUF1 (N715, N709);
or OR3 (N716, N708, N278, N143);
and AND4 (N717, N715, N393, N153, N438);
not NOT1 (N718, N717);
nor NOR2 (N719, N718, N487);
not NOT1 (N720, N705);
not NOT1 (N721, N706);
and AND2 (N722, N692, N612);
nand NAND3 (N723, N720, N91, N266);
or OR3 (N724, N722, N136, N38);
nand NAND3 (N725, N703, N518, N277);
nand NAND3 (N726, N716, N279, N589);
nor NOR3 (N727, N714, N395, N202);
nand NAND2 (N728, N719, N10);
or OR4 (N729, N713, N221, N270, N56);
xor XOR2 (N730, N699, N575);
buf BUF1 (N731, N725);
and AND2 (N732, N712, N493);
buf BUF1 (N733, N727);
and AND2 (N734, N733, N372);
buf BUF1 (N735, N732);
xor XOR2 (N736, N721, N255);
nand NAND2 (N737, N726, N670);
and AND3 (N738, N730, N466, N460);
nor NOR3 (N739, N738, N463, N573);
and AND4 (N740, N736, N707, N545, N346);
and AND2 (N741, N740, N422);
not NOT1 (N742, N737);
nor NOR4 (N743, N723, N456, N338, N225);
xor XOR2 (N744, N731, N10);
or OR3 (N745, N729, N596, N232);
and AND2 (N746, N735, N236);
or OR3 (N747, N728, N713, N745);
xor XOR2 (N748, N20, N736);
nand NAND3 (N749, N743, N585, N139);
xor XOR2 (N750, N739, N255);
nor NOR3 (N751, N724, N533, N351);
xor XOR2 (N752, N750, N255);
nand NAND4 (N753, N742, N409, N230, N91);
not NOT1 (N754, N741);
nor NOR2 (N755, N746, N361);
or OR2 (N756, N744, N37);
and AND4 (N757, N753, N338, N366, N205);
nor NOR2 (N758, N754, N456);
nand NAND2 (N759, N748, N522);
nor NOR4 (N760, N759, N644, N558, N356);
nand NAND3 (N761, N760, N329, N43);
xor XOR2 (N762, N761, N12);
or OR2 (N763, N751, N196);
or OR2 (N764, N749, N682);
xor XOR2 (N765, N734, N481);
not NOT1 (N766, N755);
nor NOR4 (N767, N757, N204, N603, N240);
not NOT1 (N768, N766);
nor NOR4 (N769, N768, N213, N20, N511);
buf BUF1 (N770, N752);
xor XOR2 (N771, N765, N407);
not NOT1 (N772, N770);
buf BUF1 (N773, N771);
not NOT1 (N774, N763);
xor XOR2 (N775, N769, N684);
buf BUF1 (N776, N747);
nor NOR3 (N777, N758, N59, N389);
nor NOR4 (N778, N762, N120, N468, N585);
and AND2 (N779, N772, N457);
nor NOR2 (N780, N767, N27);
buf BUF1 (N781, N780);
xor XOR2 (N782, N775, N137);
not NOT1 (N783, N782);
or OR3 (N784, N774, N228, N337);
buf BUF1 (N785, N776);
nor NOR4 (N786, N778, N380, N584, N685);
xor XOR2 (N787, N779, N340);
not NOT1 (N788, N783);
buf BUF1 (N789, N781);
xor XOR2 (N790, N788, N309);
nor NOR4 (N791, N764, N677, N633, N506);
nor NOR2 (N792, N791, N76);
nand NAND2 (N793, N773, N505);
or OR4 (N794, N793, N110, N170, N551);
xor XOR2 (N795, N784, N469);
and AND2 (N796, N787, N35);
buf BUF1 (N797, N785);
and AND4 (N798, N777, N557, N96, N201);
xor XOR2 (N799, N790, N656);
not NOT1 (N800, N794);
or OR4 (N801, N789, N377, N549, N667);
nor NOR4 (N802, N798, N700, N729, N139);
and AND3 (N803, N796, N417, N346);
nor NOR2 (N804, N803, N548);
not NOT1 (N805, N795);
not NOT1 (N806, N800);
or OR2 (N807, N804, N273);
nand NAND2 (N808, N792, N349);
and AND2 (N809, N756, N278);
or OR2 (N810, N806, N428);
not NOT1 (N811, N799);
buf BUF1 (N812, N786);
xor XOR2 (N813, N805, N333);
and AND4 (N814, N808, N298, N92, N209);
xor XOR2 (N815, N812, N737);
xor XOR2 (N816, N807, N396);
and AND2 (N817, N809, N235);
xor XOR2 (N818, N810, N340);
nor NOR4 (N819, N811, N310, N694, N489);
xor XOR2 (N820, N816, N646);
buf BUF1 (N821, N820);
and AND4 (N822, N813, N174, N550, N393);
buf BUF1 (N823, N822);
and AND3 (N824, N823, N613, N285);
or OR4 (N825, N818, N330, N384, N352);
buf BUF1 (N826, N821);
xor XOR2 (N827, N817, N140);
nand NAND2 (N828, N819, N238);
or OR2 (N829, N826, N172);
and AND4 (N830, N814, N480, N764, N734);
buf BUF1 (N831, N802);
not NOT1 (N832, N830);
nand NAND3 (N833, N827, N388, N500);
nor NOR4 (N834, N832, N817, N442, N162);
nor NOR2 (N835, N828, N553);
not NOT1 (N836, N835);
xor XOR2 (N837, N797, N407);
buf BUF1 (N838, N833);
and AND3 (N839, N834, N698, N135);
buf BUF1 (N840, N815);
not NOT1 (N841, N838);
nor NOR4 (N842, N829, N416, N488, N648);
nor NOR3 (N843, N824, N746, N305);
not NOT1 (N844, N837);
nor NOR4 (N845, N831, N16, N811, N752);
nor NOR2 (N846, N843, N82);
buf BUF1 (N847, N840);
and AND3 (N848, N847, N505, N500);
buf BUF1 (N849, N848);
or OR2 (N850, N841, N266);
nor NOR4 (N851, N844, N107, N221, N798);
nor NOR3 (N852, N846, N805, N632);
and AND3 (N853, N842, N338, N135);
not NOT1 (N854, N801);
not NOT1 (N855, N851);
and AND3 (N856, N854, N475, N493);
or OR3 (N857, N845, N533, N565);
nor NOR4 (N858, N825, N423, N768, N418);
and AND2 (N859, N857, N375);
not NOT1 (N860, N856);
buf BUF1 (N861, N853);
nor NOR2 (N862, N836, N679);
or OR2 (N863, N839, N550);
nor NOR4 (N864, N863, N305, N282, N391);
nand NAND4 (N865, N864, N210, N618, N168);
xor XOR2 (N866, N858, N118);
nor NOR4 (N867, N849, N791, N746, N825);
buf BUF1 (N868, N860);
nand NAND4 (N869, N850, N833, N39, N102);
xor XOR2 (N870, N867, N411);
buf BUF1 (N871, N861);
not NOT1 (N872, N855);
not NOT1 (N873, N862);
buf BUF1 (N874, N872);
or OR4 (N875, N859, N136, N253, N352);
nand NAND3 (N876, N873, N708, N403);
not NOT1 (N877, N866);
not NOT1 (N878, N870);
nand NAND3 (N879, N877, N606, N125);
or OR3 (N880, N878, N537, N411);
not NOT1 (N881, N874);
xor XOR2 (N882, N881, N538);
and AND2 (N883, N879, N35);
xor XOR2 (N884, N883, N740);
buf BUF1 (N885, N884);
and AND2 (N886, N865, N443);
buf BUF1 (N887, N882);
and AND2 (N888, N875, N406);
nand NAND2 (N889, N880, N539);
not NOT1 (N890, N889);
and AND3 (N891, N869, N407, N827);
buf BUF1 (N892, N868);
and AND4 (N893, N887, N835, N440, N526);
and AND3 (N894, N892, N179, N590);
nor NOR2 (N895, N890, N763);
and AND4 (N896, N894, N345, N847, N422);
or OR4 (N897, N876, N496, N826, N92);
nor NOR4 (N898, N891, N235, N52, N67);
nor NOR3 (N899, N897, N720, N723);
or OR4 (N900, N886, N118, N231, N895);
xor XOR2 (N901, N665, N664);
nand NAND2 (N902, N896, N111);
nor NOR2 (N903, N871, N573);
nor NOR4 (N904, N898, N400, N354, N607);
nor NOR2 (N905, N904, N596);
nand NAND2 (N906, N903, N358);
and AND3 (N907, N900, N686, N636);
or OR3 (N908, N852, N786, N662);
not NOT1 (N909, N905);
nor NOR3 (N910, N893, N190, N260);
not NOT1 (N911, N910);
nor NOR2 (N912, N907, N1);
nand NAND3 (N913, N885, N244, N480);
and AND4 (N914, N888, N674, N17, N902);
not NOT1 (N915, N339);
or OR4 (N916, N909, N490, N433, N476);
buf BUF1 (N917, N914);
buf BUF1 (N918, N915);
nor NOR2 (N919, N918, N578);
nor NOR2 (N920, N908, N725);
xor XOR2 (N921, N913, N889);
not NOT1 (N922, N901);
and AND4 (N923, N922, N553, N286, N79);
nand NAND3 (N924, N916, N385, N475);
buf BUF1 (N925, N911);
and AND3 (N926, N919, N402, N212);
or OR4 (N927, N925, N431, N846, N318);
or OR3 (N928, N924, N677, N194);
nand NAND4 (N929, N912, N465, N542, N98);
xor XOR2 (N930, N929, N155);
buf BUF1 (N931, N917);
not NOT1 (N932, N906);
xor XOR2 (N933, N923, N433);
buf BUF1 (N934, N933);
and AND3 (N935, N920, N529, N528);
or OR4 (N936, N921, N237, N487, N669);
buf BUF1 (N937, N931);
nand NAND4 (N938, N927, N736, N681, N812);
nand NAND2 (N939, N938, N138);
nand NAND3 (N940, N936, N644, N335);
or OR3 (N941, N899, N496, N637);
nor NOR4 (N942, N928, N124, N189, N749);
nand NAND4 (N943, N932, N229, N442, N148);
buf BUF1 (N944, N942);
nand NAND3 (N945, N941, N646, N237);
not NOT1 (N946, N930);
nor NOR2 (N947, N944, N322);
xor XOR2 (N948, N937, N807);
xor XOR2 (N949, N940, N683);
and AND2 (N950, N939, N119);
buf BUF1 (N951, N943);
and AND2 (N952, N947, N310);
or OR3 (N953, N950, N527, N928);
nor NOR3 (N954, N935, N698, N499);
xor XOR2 (N955, N949, N49);
buf BUF1 (N956, N948);
nand NAND2 (N957, N955, N672);
and AND2 (N958, N926, N199);
and AND3 (N959, N951, N4, N244);
buf BUF1 (N960, N946);
nor NOR4 (N961, N956, N887, N572, N454);
or OR4 (N962, N954, N289, N381, N612);
and AND2 (N963, N959, N210);
nor NOR3 (N964, N957, N281, N377);
or OR2 (N965, N934, N169);
nor NOR2 (N966, N945, N885);
and AND3 (N967, N958, N295, N145);
xor XOR2 (N968, N962, N89);
and AND4 (N969, N963, N215, N696, N373);
not NOT1 (N970, N960);
buf BUF1 (N971, N953);
not NOT1 (N972, N971);
and AND2 (N973, N967, N339);
not NOT1 (N974, N966);
not NOT1 (N975, N961);
xor XOR2 (N976, N969, N166);
and AND2 (N977, N968, N110);
and AND2 (N978, N970, N813);
and AND2 (N979, N973, N580);
buf BUF1 (N980, N977);
xor XOR2 (N981, N975, N4);
or OR4 (N982, N979, N177, N247, N163);
xor XOR2 (N983, N976, N269);
not NOT1 (N984, N983);
nor NOR4 (N985, N965, N922, N830, N817);
not NOT1 (N986, N964);
nand NAND2 (N987, N984, N173);
buf BUF1 (N988, N978);
xor XOR2 (N989, N985, N552);
not NOT1 (N990, N972);
not NOT1 (N991, N990);
or OR4 (N992, N952, N355, N25, N768);
nand NAND4 (N993, N986, N861, N53, N758);
or OR4 (N994, N987, N308, N571, N635);
or OR3 (N995, N994, N272, N980);
not NOT1 (N996, N594);
nand NAND2 (N997, N974, N87);
xor XOR2 (N998, N993, N189);
nor NOR4 (N999, N992, N236, N764, N620);
and AND4 (N1000, N988, N660, N673, N649);
buf BUF1 (N1001, N998);
not NOT1 (N1002, N1001);
nand NAND3 (N1003, N996, N81, N342);
nand NAND4 (N1004, N991, N156, N546, N527);
or OR2 (N1005, N982, N882);
buf BUF1 (N1006, N995);
or OR3 (N1007, N1006, N767, N948);
not NOT1 (N1008, N1007);
xor XOR2 (N1009, N1005, N619);
nor NOR2 (N1010, N1009, N831);
not NOT1 (N1011, N1008);
and AND4 (N1012, N1010, N259, N164, N339);
xor XOR2 (N1013, N1012, N60);
xor XOR2 (N1014, N1004, N248);
or OR4 (N1015, N981, N833, N227, N140);
buf BUF1 (N1016, N997);
buf BUF1 (N1017, N1000);
nand NAND3 (N1018, N1003, N121, N446);
and AND3 (N1019, N999, N180, N490);
nand NAND4 (N1020, N1019, N44, N388, N483);
not NOT1 (N1021, N1014);
not NOT1 (N1022, N1017);
nand NAND3 (N1023, N1020, N357, N31);
not NOT1 (N1024, N1002);
not NOT1 (N1025, N1015);
xor XOR2 (N1026, N1016, N306);
nor NOR3 (N1027, N1013, N947, N857);
nor NOR4 (N1028, N1022, N13, N163, N656);
not NOT1 (N1029, N989);
not NOT1 (N1030, N1027);
not NOT1 (N1031, N1023);
nor NOR4 (N1032, N1011, N191, N877, N175);
not NOT1 (N1033, N1018);
not NOT1 (N1034, N1028);
nand NAND2 (N1035, N1026, N450);
or OR4 (N1036, N1030, N919, N704, N705);
buf BUF1 (N1037, N1035);
or OR2 (N1038, N1034, N216);
buf BUF1 (N1039, N1025);
and AND3 (N1040, N1038, N369, N727);
not NOT1 (N1041, N1036);
or OR4 (N1042, N1021, N46, N597, N744);
nand NAND4 (N1043, N1029, N432, N798, N855);
buf BUF1 (N1044, N1024);
nand NAND4 (N1045, N1031, N320, N102, N449);
and AND3 (N1046, N1041, N247, N66);
not NOT1 (N1047, N1045);
not NOT1 (N1048, N1033);
buf BUF1 (N1049, N1046);
nor NOR2 (N1050, N1037, N884);
xor XOR2 (N1051, N1039, N528);
nand NAND4 (N1052, N1048, N595, N681, N386);
nand NAND3 (N1053, N1052, N328, N1016);
not NOT1 (N1054, N1050);
not NOT1 (N1055, N1053);
xor XOR2 (N1056, N1047, N579);
not NOT1 (N1057, N1049);
xor XOR2 (N1058, N1043, N445);
and AND3 (N1059, N1032, N820, N49);
not NOT1 (N1060, N1057);
not NOT1 (N1061, N1054);
xor XOR2 (N1062, N1040, N886);
and AND3 (N1063, N1042, N988, N813);
buf BUF1 (N1064, N1044);
nor NOR2 (N1065, N1062, N715);
nand NAND4 (N1066, N1059, N670, N824, N437);
buf BUF1 (N1067, N1065);
nand NAND4 (N1068, N1060, N254, N797, N94);
buf BUF1 (N1069, N1061);
and AND3 (N1070, N1069, N811, N486);
nand NAND3 (N1071, N1070, N166, N14);
buf BUF1 (N1072, N1055);
or OR3 (N1073, N1051, N131, N949);
or OR3 (N1074, N1072, N528, N823);
buf BUF1 (N1075, N1058);
buf BUF1 (N1076, N1067);
nor NOR4 (N1077, N1073, N351, N266, N730);
nor NOR2 (N1078, N1076, N132);
not NOT1 (N1079, N1074);
xor XOR2 (N1080, N1063, N548);
buf BUF1 (N1081, N1071);
not NOT1 (N1082, N1079);
nor NOR3 (N1083, N1077, N868, N66);
and AND4 (N1084, N1082, N591, N391, N214);
nor NOR2 (N1085, N1084, N842);
not NOT1 (N1086, N1068);
and AND2 (N1087, N1083, N851);
and AND3 (N1088, N1078, N865, N418);
not NOT1 (N1089, N1086);
nor NOR2 (N1090, N1085, N824);
and AND3 (N1091, N1056, N685, N71);
xor XOR2 (N1092, N1064, N1084);
nand NAND3 (N1093, N1087, N546, N1058);
or OR2 (N1094, N1066, N146);
nor NOR4 (N1095, N1094, N1093, N381, N698);
nor NOR4 (N1096, N762, N143, N741, N155);
xor XOR2 (N1097, N1088, N838);
buf BUF1 (N1098, N1080);
nor NOR4 (N1099, N1096, N139, N770, N1087);
not NOT1 (N1100, N1097);
or OR3 (N1101, N1091, N192, N885);
and AND4 (N1102, N1098, N695, N782, N1070);
and AND3 (N1103, N1095, N802, N186);
nand NAND2 (N1104, N1100, N520);
xor XOR2 (N1105, N1075, N3);
or OR4 (N1106, N1092, N250, N889, N143);
buf BUF1 (N1107, N1105);
or OR3 (N1108, N1104, N431, N875);
not NOT1 (N1109, N1099);
nand NAND3 (N1110, N1106, N98, N871);
nand NAND2 (N1111, N1081, N280);
or OR3 (N1112, N1103, N737, N967);
nand NAND4 (N1113, N1110, N627, N26, N771);
or OR4 (N1114, N1113, N895, N171, N184);
or OR2 (N1115, N1109, N98);
nand NAND2 (N1116, N1111, N994);
nand NAND4 (N1117, N1089, N971, N485, N496);
nand NAND2 (N1118, N1112, N295);
buf BUF1 (N1119, N1118);
buf BUF1 (N1120, N1119);
buf BUF1 (N1121, N1116);
or OR2 (N1122, N1121, N393);
nor NOR4 (N1123, N1114, N142, N612, N875);
xor XOR2 (N1124, N1120, N1013);
or OR4 (N1125, N1122, N169, N592, N494);
not NOT1 (N1126, N1124);
or OR4 (N1127, N1117, N1020, N6, N942);
or OR4 (N1128, N1108, N1095, N857, N516);
or OR3 (N1129, N1123, N175, N1033);
or OR3 (N1130, N1102, N225, N737);
and AND4 (N1131, N1125, N660, N801, N557);
buf BUF1 (N1132, N1090);
not NOT1 (N1133, N1101);
or OR2 (N1134, N1126, N152);
nand NAND2 (N1135, N1130, N837);
not NOT1 (N1136, N1135);
not NOT1 (N1137, N1134);
or OR3 (N1138, N1129, N1046, N15);
buf BUF1 (N1139, N1133);
or OR4 (N1140, N1128, N580, N758, N857);
and AND3 (N1141, N1115, N598, N633);
xor XOR2 (N1142, N1131, N337);
xor XOR2 (N1143, N1138, N52);
and AND2 (N1144, N1143, N119);
not NOT1 (N1145, N1141);
xor XOR2 (N1146, N1107, N120);
nor NOR3 (N1147, N1139, N564, N447);
nand NAND4 (N1148, N1145, N580, N926, N1089);
buf BUF1 (N1149, N1147);
not NOT1 (N1150, N1144);
not NOT1 (N1151, N1148);
xor XOR2 (N1152, N1146, N841);
buf BUF1 (N1153, N1137);
or OR2 (N1154, N1150, N20);
not NOT1 (N1155, N1140);
and AND3 (N1156, N1127, N859, N96);
nand NAND3 (N1157, N1142, N170, N938);
not NOT1 (N1158, N1156);
not NOT1 (N1159, N1155);
nand NAND4 (N1160, N1132, N131, N415, N174);
nor NOR4 (N1161, N1160, N614, N846, N876);
buf BUF1 (N1162, N1152);
nor NOR3 (N1163, N1161, N510, N320);
and AND3 (N1164, N1154, N429, N529);
or OR2 (N1165, N1149, N523);
nand NAND2 (N1166, N1165, N48);
nand NAND3 (N1167, N1162, N243, N482);
not NOT1 (N1168, N1157);
and AND4 (N1169, N1166, N933, N173, N283);
nand NAND2 (N1170, N1169, N974);
buf BUF1 (N1171, N1151);
nor NOR3 (N1172, N1159, N46, N315);
nor NOR2 (N1173, N1170, N213);
or OR2 (N1174, N1171, N399);
and AND4 (N1175, N1172, N460, N131, N929);
nand NAND3 (N1176, N1136, N375, N282);
nand NAND4 (N1177, N1163, N137, N81, N427);
nand NAND4 (N1178, N1164, N383, N59, N202);
nor NOR2 (N1179, N1175, N881);
not NOT1 (N1180, N1174);
buf BUF1 (N1181, N1178);
not NOT1 (N1182, N1181);
xor XOR2 (N1183, N1179, N412);
or OR4 (N1184, N1153, N272, N469, N18);
and AND3 (N1185, N1168, N840, N39);
buf BUF1 (N1186, N1167);
nor NOR2 (N1187, N1185, N64);
xor XOR2 (N1188, N1183, N215);
xor XOR2 (N1189, N1158, N1008);
buf BUF1 (N1190, N1173);
buf BUF1 (N1191, N1188);
and AND2 (N1192, N1187, N1078);
nand NAND4 (N1193, N1180, N115, N762, N241);
nand NAND2 (N1194, N1182, N1007);
buf BUF1 (N1195, N1192);
nor NOR2 (N1196, N1193, N1017);
nand NAND3 (N1197, N1190, N1154, N732);
and AND3 (N1198, N1195, N294, N557);
not NOT1 (N1199, N1189);
xor XOR2 (N1200, N1194, N689);
xor XOR2 (N1201, N1200, N1163);
xor XOR2 (N1202, N1197, N469);
buf BUF1 (N1203, N1176);
not NOT1 (N1204, N1201);
nand NAND2 (N1205, N1196, N716);
buf BUF1 (N1206, N1199);
or OR3 (N1207, N1204, N16, N1188);
nor NOR3 (N1208, N1205, N847, N458);
nor NOR2 (N1209, N1208, N50);
and AND4 (N1210, N1177, N592, N296, N152);
not NOT1 (N1211, N1186);
or OR3 (N1212, N1184, N770, N87);
nor NOR3 (N1213, N1203, N710, N713);
not NOT1 (N1214, N1209);
nand NAND4 (N1215, N1206, N185, N673, N112);
and AND3 (N1216, N1198, N129, N650);
nor NOR4 (N1217, N1211, N453, N770, N1001);
or OR4 (N1218, N1215, N1004, N14, N1112);
not NOT1 (N1219, N1217);
xor XOR2 (N1220, N1213, N708);
or OR4 (N1221, N1202, N340, N144, N1071);
nand NAND2 (N1222, N1191, N70);
nor NOR4 (N1223, N1212, N457, N342, N137);
buf BUF1 (N1224, N1214);
and AND4 (N1225, N1222, N1190, N937, N542);
and AND3 (N1226, N1223, N754, N954);
nand NAND4 (N1227, N1224, N201, N826, N798);
not NOT1 (N1228, N1227);
xor XOR2 (N1229, N1219, N1158);
not NOT1 (N1230, N1220);
nand NAND4 (N1231, N1221, N631, N135, N278);
nor NOR3 (N1232, N1230, N768, N543);
nand NAND4 (N1233, N1210, N1081, N945, N540);
nand NAND3 (N1234, N1229, N975, N1210);
nand NAND3 (N1235, N1216, N765, N441);
nand NAND2 (N1236, N1234, N377);
and AND2 (N1237, N1226, N663);
or OR2 (N1238, N1231, N555);
not NOT1 (N1239, N1232);
or OR2 (N1240, N1236, N571);
nand NAND4 (N1241, N1233, N1011, N184, N32);
or OR3 (N1242, N1238, N222, N210);
and AND3 (N1243, N1207, N377, N394);
xor XOR2 (N1244, N1241, N689);
or OR4 (N1245, N1237, N251, N501, N650);
nor NOR3 (N1246, N1225, N636, N583);
nor NOR2 (N1247, N1242, N77);
and AND3 (N1248, N1246, N1079, N368);
nand NAND3 (N1249, N1240, N170, N865);
or OR4 (N1250, N1243, N378, N148, N535);
buf BUF1 (N1251, N1247);
or OR3 (N1252, N1245, N134, N137);
buf BUF1 (N1253, N1239);
nand NAND4 (N1254, N1244, N731, N434, N579);
and AND4 (N1255, N1228, N953, N1203, N938);
nand NAND4 (N1256, N1254, N7, N169, N65);
and AND3 (N1257, N1218, N351, N301);
or OR2 (N1258, N1235, N1216);
and AND3 (N1259, N1249, N171, N342);
not NOT1 (N1260, N1258);
and AND3 (N1261, N1257, N141, N1151);
nand NAND4 (N1262, N1260, N746, N77, N947);
buf BUF1 (N1263, N1248);
or OR4 (N1264, N1253, N983, N233, N1124);
not NOT1 (N1265, N1256);
not NOT1 (N1266, N1250);
nor NOR4 (N1267, N1263, N876, N759, N1024);
or OR2 (N1268, N1264, N973);
not NOT1 (N1269, N1255);
nand NAND3 (N1270, N1262, N41, N1110);
nor NOR3 (N1271, N1267, N584, N544);
nand NAND4 (N1272, N1251, N57, N586, N1062);
nand NAND4 (N1273, N1270, N596, N1236, N60);
nor NOR4 (N1274, N1259, N149, N1060, N502);
nand NAND3 (N1275, N1269, N591, N34);
buf BUF1 (N1276, N1274);
not NOT1 (N1277, N1273);
not NOT1 (N1278, N1266);
not NOT1 (N1279, N1265);
nand NAND4 (N1280, N1278, N251, N989, N544);
nor NOR4 (N1281, N1271, N1041, N782, N1115);
xor XOR2 (N1282, N1272, N297);
xor XOR2 (N1283, N1282, N392);
nor NOR4 (N1284, N1277, N218, N886, N48);
buf BUF1 (N1285, N1280);
buf BUF1 (N1286, N1275);
xor XOR2 (N1287, N1261, N257);
nor NOR4 (N1288, N1276, N497, N1220, N184);
not NOT1 (N1289, N1268);
buf BUF1 (N1290, N1286);
not NOT1 (N1291, N1289);
xor XOR2 (N1292, N1281, N836);
buf BUF1 (N1293, N1285);
or OR4 (N1294, N1291, N393, N542, N737);
nand NAND4 (N1295, N1284, N1041, N802, N568);
buf BUF1 (N1296, N1293);
buf BUF1 (N1297, N1295);
not NOT1 (N1298, N1287);
nor NOR4 (N1299, N1252, N1141, N610, N792);
and AND2 (N1300, N1290, N989);
nand NAND4 (N1301, N1299, N1227, N85, N1291);
not NOT1 (N1302, N1288);
nand NAND2 (N1303, N1297, N146);
nor NOR4 (N1304, N1279, N405, N124, N795);
nand NAND4 (N1305, N1301, N961, N542, N908);
and AND3 (N1306, N1303, N414, N1048);
nand NAND2 (N1307, N1305, N652);
buf BUF1 (N1308, N1302);
nor NOR4 (N1309, N1294, N161, N427, N232);
and AND2 (N1310, N1309, N555);
and AND2 (N1311, N1296, N100);
nand NAND3 (N1312, N1283, N1021, N856);
nor NOR2 (N1313, N1311, N1175);
or OR3 (N1314, N1304, N555, N3);
or OR2 (N1315, N1306, N788);
and AND4 (N1316, N1314, N101, N615, N456);
nand NAND3 (N1317, N1312, N539, N837);
nor NOR2 (N1318, N1307, N899);
nand NAND2 (N1319, N1292, N514);
or OR3 (N1320, N1319, N479, N982);
nand NAND2 (N1321, N1308, N983);
xor XOR2 (N1322, N1315, N396);
not NOT1 (N1323, N1298);
and AND2 (N1324, N1321, N1041);
and AND4 (N1325, N1300, N1146, N884, N1010);
and AND3 (N1326, N1316, N387, N314);
and AND2 (N1327, N1318, N316);
nand NAND2 (N1328, N1320, N304);
nand NAND4 (N1329, N1328, N1127, N181, N207);
nor NOR4 (N1330, N1324, N394, N850, N1250);
and AND2 (N1331, N1330, N76);
xor XOR2 (N1332, N1322, N65);
nand NAND2 (N1333, N1310, N789);
not NOT1 (N1334, N1313);
not NOT1 (N1335, N1326);
xor XOR2 (N1336, N1335, N860);
xor XOR2 (N1337, N1325, N978);
xor XOR2 (N1338, N1334, N1170);
or OR4 (N1339, N1337, N1234, N210, N1258);
nand NAND2 (N1340, N1339, N1121);
buf BUF1 (N1341, N1329);
not NOT1 (N1342, N1332);
or OR3 (N1343, N1317, N1190, N26);
and AND3 (N1344, N1333, N97, N466);
not NOT1 (N1345, N1327);
nand NAND2 (N1346, N1345, N237);
xor XOR2 (N1347, N1342, N286);
and AND3 (N1348, N1323, N622, N411);
nor NOR4 (N1349, N1346, N688, N635, N582);
nor NOR4 (N1350, N1340, N260, N1094, N1252);
buf BUF1 (N1351, N1350);
or OR2 (N1352, N1343, N204);
nor NOR3 (N1353, N1341, N206, N872);
or OR2 (N1354, N1331, N463);
xor XOR2 (N1355, N1353, N105);
or OR3 (N1356, N1344, N664, N1023);
and AND3 (N1357, N1336, N363, N1332);
buf BUF1 (N1358, N1354);
or OR3 (N1359, N1352, N16, N882);
buf BUF1 (N1360, N1349);
or OR3 (N1361, N1356, N1262, N272);
or OR2 (N1362, N1361, N1118);
nand NAND3 (N1363, N1362, N693, N1307);
xor XOR2 (N1364, N1351, N1092);
not NOT1 (N1365, N1355);
not NOT1 (N1366, N1348);
not NOT1 (N1367, N1358);
or OR4 (N1368, N1367, N1194, N100, N23);
xor XOR2 (N1369, N1357, N314);
and AND2 (N1370, N1359, N80);
buf BUF1 (N1371, N1365);
and AND2 (N1372, N1371, N1008);
xor XOR2 (N1373, N1347, N1029);
nand NAND4 (N1374, N1370, N1058, N223, N788);
buf BUF1 (N1375, N1360);
buf BUF1 (N1376, N1368);
nand NAND3 (N1377, N1369, N1074, N307);
or OR3 (N1378, N1364, N1280, N1232);
or OR2 (N1379, N1373, N560);
or OR3 (N1380, N1338, N1319, N913);
or OR2 (N1381, N1376, N1004);
not NOT1 (N1382, N1377);
nand NAND4 (N1383, N1378, N1240, N68, N987);
xor XOR2 (N1384, N1375, N1075);
or OR2 (N1385, N1381, N799);
xor XOR2 (N1386, N1382, N658);
nand NAND2 (N1387, N1363, N1269);
xor XOR2 (N1388, N1386, N1116);
and AND4 (N1389, N1380, N731, N104, N913);
buf BUF1 (N1390, N1383);
xor XOR2 (N1391, N1385, N492);
not NOT1 (N1392, N1366);
xor XOR2 (N1393, N1372, N1210);
nand NAND4 (N1394, N1390, N134, N990, N62);
nand NAND4 (N1395, N1384, N1246, N282, N619);
not NOT1 (N1396, N1374);
nand NAND4 (N1397, N1379, N1377, N626, N350);
xor XOR2 (N1398, N1393, N217);
not NOT1 (N1399, N1395);
or OR4 (N1400, N1391, N491, N1214, N1130);
nor NOR4 (N1401, N1397, N936, N1390, N1042);
buf BUF1 (N1402, N1396);
or OR2 (N1403, N1402, N407);
or OR3 (N1404, N1388, N669, N537);
or OR4 (N1405, N1400, N263, N561, N798);
or OR3 (N1406, N1403, N350, N458);
nor NOR2 (N1407, N1392, N541);
and AND4 (N1408, N1404, N995, N1302, N169);
buf BUF1 (N1409, N1398);
and AND2 (N1410, N1399, N117);
not NOT1 (N1411, N1409);
nor NOR3 (N1412, N1408, N885, N97);
and AND3 (N1413, N1411, N837, N662);
not NOT1 (N1414, N1406);
nand NAND4 (N1415, N1389, N968, N778, N303);
or OR2 (N1416, N1412, N49);
not NOT1 (N1417, N1414);
or OR3 (N1418, N1405, N136, N646);
buf BUF1 (N1419, N1417);
nand NAND3 (N1420, N1387, N273, N1410);
buf BUF1 (N1421, N220);
nor NOR3 (N1422, N1401, N229, N936);
not NOT1 (N1423, N1416);
xor XOR2 (N1424, N1418, N1363);
or OR2 (N1425, N1419, N291);
and AND4 (N1426, N1413, N980, N380, N665);
nor NOR2 (N1427, N1426, N965);
and AND4 (N1428, N1394, N333, N1126, N706);
or OR2 (N1429, N1425, N761);
or OR3 (N1430, N1424, N1048, N200);
xor XOR2 (N1431, N1415, N475);
nand NAND4 (N1432, N1422, N887, N832, N835);
nor NOR3 (N1433, N1428, N244, N338);
buf BUF1 (N1434, N1430);
and AND3 (N1435, N1433, N514, N262);
or OR2 (N1436, N1423, N112);
or OR4 (N1437, N1434, N864, N756, N877);
nand NAND2 (N1438, N1420, N141);
nor NOR3 (N1439, N1435, N66, N859);
nor NOR3 (N1440, N1438, N397, N691);
xor XOR2 (N1441, N1429, N831);
nor NOR2 (N1442, N1439, N1226);
and AND3 (N1443, N1407, N267, N190);
nand NAND2 (N1444, N1440, N220);
and AND4 (N1445, N1441, N773, N662, N1085);
and AND2 (N1446, N1437, N218);
nand NAND2 (N1447, N1446, N816);
nor NOR3 (N1448, N1436, N489, N157);
or OR3 (N1449, N1421, N1439, N219);
buf BUF1 (N1450, N1448);
nand NAND4 (N1451, N1427, N1323, N1439, N208);
nor NOR2 (N1452, N1449, N1450);
nand NAND2 (N1453, N1075, N705);
not NOT1 (N1454, N1451);
and AND3 (N1455, N1444, N215, N832);
not NOT1 (N1456, N1455);
nand NAND4 (N1457, N1443, N770, N1301, N1107);
or OR3 (N1458, N1453, N878, N1333);
nor NOR2 (N1459, N1432, N819);
and AND2 (N1460, N1458, N446);
xor XOR2 (N1461, N1454, N735);
xor XOR2 (N1462, N1459, N186);
not NOT1 (N1463, N1445);
buf BUF1 (N1464, N1457);
buf BUF1 (N1465, N1456);
xor XOR2 (N1466, N1431, N1462);
buf BUF1 (N1467, N160);
nand NAND3 (N1468, N1463, N1391, N1301);
xor XOR2 (N1469, N1464, N725);
or OR2 (N1470, N1466, N200);
nor NOR4 (N1471, N1447, N1265, N319, N325);
and AND3 (N1472, N1468, N678, N66);
buf BUF1 (N1473, N1470);
nor NOR4 (N1474, N1442, N418, N1451, N1420);
and AND2 (N1475, N1473, N1272);
nor NOR2 (N1476, N1461, N170);
or OR4 (N1477, N1452, N186, N439, N1045);
xor XOR2 (N1478, N1467, N894);
not NOT1 (N1479, N1475);
nor NOR4 (N1480, N1460, N869, N903, N1356);
nand NAND2 (N1481, N1479, N250);
buf BUF1 (N1482, N1465);
nor NOR4 (N1483, N1471, N1098, N34, N207);
nor NOR4 (N1484, N1482, N875, N694, N886);
nor NOR3 (N1485, N1480, N472, N306);
not NOT1 (N1486, N1484);
and AND3 (N1487, N1477, N167, N1468);
or OR2 (N1488, N1483, N653);
nand NAND4 (N1489, N1485, N80, N524, N841);
nor NOR3 (N1490, N1476, N937, N658);
or OR4 (N1491, N1489, N574, N1039, N1394);
nand NAND4 (N1492, N1469, N540, N895, N1486);
and AND2 (N1493, N233, N1346);
and AND3 (N1494, N1474, N1022, N377);
xor XOR2 (N1495, N1478, N106);
buf BUF1 (N1496, N1487);
buf BUF1 (N1497, N1488);
or OR2 (N1498, N1492, N162);
or OR2 (N1499, N1496, N998);
buf BUF1 (N1500, N1491);
not NOT1 (N1501, N1497);
and AND2 (N1502, N1498, N106);
nand NAND2 (N1503, N1495, N11);
and AND4 (N1504, N1493, N1377, N1384, N159);
nand NAND3 (N1505, N1472, N924, N2);
or OR2 (N1506, N1501, N82);
nor NOR4 (N1507, N1500, N1192, N1194, N256);
and AND4 (N1508, N1490, N880, N930, N1488);
or OR3 (N1509, N1504, N1215, N664);
not NOT1 (N1510, N1494);
nor NOR4 (N1511, N1503, N1331, N425, N413);
nor NOR3 (N1512, N1499, N672, N176);
xor XOR2 (N1513, N1507, N376);
not NOT1 (N1514, N1481);
and AND3 (N1515, N1511, N814, N346);
nand NAND3 (N1516, N1510, N651, N666);
xor XOR2 (N1517, N1516, N435);
nand NAND3 (N1518, N1505, N897, N419);
nand NAND3 (N1519, N1502, N665, N59);
or OR4 (N1520, N1519, N1261, N1190, N161);
or OR4 (N1521, N1508, N713, N69, N607);
not NOT1 (N1522, N1512);
or OR4 (N1523, N1518, N266, N1285, N12);
or OR4 (N1524, N1522, N458, N1094, N1264);
nand NAND3 (N1525, N1509, N605, N320);
not NOT1 (N1526, N1525);
nand NAND2 (N1527, N1513, N301);
or OR4 (N1528, N1520, N800, N91, N1304);
nand NAND2 (N1529, N1514, N1190);
xor XOR2 (N1530, N1506, N621);
or OR2 (N1531, N1528, N75);
not NOT1 (N1532, N1531);
nor NOR3 (N1533, N1521, N689, N689);
buf BUF1 (N1534, N1524);
and AND3 (N1535, N1517, N1390, N1195);
or OR3 (N1536, N1534, N688, N1291);
and AND2 (N1537, N1536, N1346);
and AND2 (N1538, N1530, N1277);
and AND3 (N1539, N1533, N1257, N265);
not NOT1 (N1540, N1532);
and AND2 (N1541, N1535, N85);
buf BUF1 (N1542, N1541);
nand NAND4 (N1543, N1539, N1507, N625, N29);
not NOT1 (N1544, N1543);
buf BUF1 (N1545, N1537);
nand NAND4 (N1546, N1515, N801, N130, N574);
nor NOR3 (N1547, N1540, N252, N1261);
not NOT1 (N1548, N1546);
nor NOR2 (N1549, N1545, N393);
xor XOR2 (N1550, N1526, N220);
not NOT1 (N1551, N1548);
and AND2 (N1552, N1527, N222);
xor XOR2 (N1553, N1538, N1235);
nor NOR3 (N1554, N1551, N967, N4);
buf BUF1 (N1555, N1542);
not NOT1 (N1556, N1549);
not NOT1 (N1557, N1556);
nand NAND2 (N1558, N1523, N1537);
nand NAND2 (N1559, N1555, N536);
not NOT1 (N1560, N1529);
or OR3 (N1561, N1553, N1539, N147);
nor NOR2 (N1562, N1550, N1090);
nand NAND2 (N1563, N1554, N120);
and AND4 (N1564, N1558, N1454, N904, N818);
and AND3 (N1565, N1562, N1539, N1344);
not NOT1 (N1566, N1547);
xor XOR2 (N1567, N1564, N1163);
buf BUF1 (N1568, N1557);
nand NAND2 (N1569, N1568, N61);
not NOT1 (N1570, N1569);
or OR3 (N1571, N1544, N188, N182);
and AND4 (N1572, N1560, N1480, N560, N798);
buf BUF1 (N1573, N1559);
buf BUF1 (N1574, N1561);
and AND3 (N1575, N1566, N708, N959);
and AND2 (N1576, N1575, N1468);
not NOT1 (N1577, N1576);
or OR4 (N1578, N1572, N1072, N166, N1117);
and AND3 (N1579, N1574, N1127, N1054);
xor XOR2 (N1580, N1573, N541);
and AND2 (N1581, N1578, N724);
nor NOR4 (N1582, N1565, N1101, N716, N1501);
or OR4 (N1583, N1552, N1235, N1320, N327);
nand NAND3 (N1584, N1571, N1198, N391);
and AND3 (N1585, N1567, N18, N1355);
nor NOR4 (N1586, N1563, N1255, N1003, N647);
not NOT1 (N1587, N1582);
xor XOR2 (N1588, N1586, N1445);
nand NAND4 (N1589, N1579, N905, N825, N1099);
xor XOR2 (N1590, N1581, N1000);
buf BUF1 (N1591, N1570);
xor XOR2 (N1592, N1587, N628);
xor XOR2 (N1593, N1580, N794);
nand NAND2 (N1594, N1590, N561);
or OR2 (N1595, N1583, N985);
buf BUF1 (N1596, N1584);
and AND2 (N1597, N1588, N601);
nor NOR4 (N1598, N1597, N612, N232, N1157);
and AND3 (N1599, N1592, N946, N731);
not NOT1 (N1600, N1595);
nor NOR3 (N1601, N1600, N1394, N898);
xor XOR2 (N1602, N1593, N1413);
or OR4 (N1603, N1601, N208, N946, N1108);
nand NAND2 (N1604, N1577, N1150);
buf BUF1 (N1605, N1591);
buf BUF1 (N1606, N1585);
nor NOR3 (N1607, N1589, N1149, N933);
or OR4 (N1608, N1594, N40, N1458, N597);
nand NAND4 (N1609, N1599, N147, N1217, N507);
nor NOR2 (N1610, N1606, N1548);
xor XOR2 (N1611, N1607, N1006);
nor NOR3 (N1612, N1598, N1073, N646);
or OR2 (N1613, N1609, N1128);
xor XOR2 (N1614, N1603, N855);
buf BUF1 (N1615, N1608);
and AND2 (N1616, N1610, N1469);
and AND2 (N1617, N1605, N1272);
buf BUF1 (N1618, N1612);
nand NAND2 (N1619, N1613, N169);
not NOT1 (N1620, N1614);
xor XOR2 (N1621, N1617, N566);
or OR4 (N1622, N1621, N1188, N87, N131);
endmodule