// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N408,N414,N421,N420,N415,N416,N418,N419,N422,N423;

nor NOR2 (N24, N9, N17);
buf BUF1 (N25, N20);
xor XOR2 (N26, N9, N2);
buf BUF1 (N27, N8);
nand NAND2 (N28, N13, N3);
nor NOR4 (N29, N6, N28, N26, N7);
and AND3 (N30, N27, N20, N6);
not NOT1 (N31, N6);
buf BUF1 (N32, N26);
or OR4 (N33, N28, N7, N4, N9);
or OR3 (N34, N31, N6, N21);
xor XOR2 (N35, N11, N23);
and AND3 (N36, N2, N29, N35);
nand NAND3 (N37, N31, N32, N12);
and AND2 (N38, N16, N25);
nor NOR2 (N39, N36, N7);
nor NOR2 (N40, N1, N31);
buf BUF1 (N41, N15);
nand NAND3 (N42, N27, N31, N33);
and AND2 (N43, N24, N24);
xor XOR2 (N44, N3, N13);
or OR2 (N45, N34, N11);
xor XOR2 (N46, N45, N38);
or OR4 (N47, N13, N32, N10, N31);
not NOT1 (N48, N47);
or OR3 (N49, N37, N30, N36);
or OR3 (N50, N16, N9, N18);
not NOT1 (N51, N49);
xor XOR2 (N52, N51, N45);
buf BUF1 (N53, N48);
buf BUF1 (N54, N52);
and AND4 (N55, N50, N36, N22, N43);
nand NAND4 (N56, N42, N25, N22, N4);
not NOT1 (N57, N39);
nand NAND3 (N58, N49, N1, N17);
buf BUF1 (N59, N46);
nor NOR3 (N60, N55, N49, N52);
or OR3 (N61, N41, N27, N55);
xor XOR2 (N62, N58, N22);
not NOT1 (N63, N61);
nor NOR4 (N64, N54, N7, N20, N30);
xor XOR2 (N65, N64, N50);
or OR4 (N66, N65, N3, N15, N61);
nor NOR2 (N67, N62, N33);
nand NAND4 (N68, N40, N5, N66, N58);
and AND2 (N69, N19, N23);
nor NOR4 (N70, N69, N50, N68, N10);
xor XOR2 (N71, N51, N5);
buf BUF1 (N72, N56);
xor XOR2 (N73, N53, N43);
nand NAND3 (N74, N71, N72, N40);
nor NOR2 (N75, N12, N60);
and AND3 (N76, N17, N68, N44);
not NOT1 (N77, N12);
nand NAND3 (N78, N57, N19, N51);
not NOT1 (N79, N77);
buf BUF1 (N80, N78);
nor NOR3 (N81, N79, N26, N1);
not NOT1 (N82, N59);
or OR4 (N83, N82, N18, N82, N53);
nor NOR3 (N84, N67, N78, N8);
nor NOR4 (N85, N70, N57, N83, N11);
nand NAND4 (N86, N68, N4, N73, N20);
xor XOR2 (N87, N11, N69);
not NOT1 (N88, N87);
xor XOR2 (N89, N80, N11);
and AND2 (N90, N86, N26);
xor XOR2 (N91, N63, N42);
and AND4 (N92, N84, N57, N18, N25);
nand NAND2 (N93, N88, N12);
or OR2 (N94, N89, N75);
not NOT1 (N95, N88);
buf BUF1 (N96, N93);
nand NAND2 (N97, N92, N22);
buf BUF1 (N98, N96);
not NOT1 (N99, N91);
nor NOR3 (N100, N85, N89, N83);
buf BUF1 (N101, N76);
xor XOR2 (N102, N98, N77);
nor NOR3 (N103, N90, N90, N75);
nor NOR2 (N104, N103, N55);
not NOT1 (N105, N74);
or OR4 (N106, N101, N104, N66, N15);
or OR2 (N107, N30, N97);
and AND4 (N108, N52, N89, N68, N12);
nor NOR4 (N109, N108, N9, N94, N32);
nand NAND3 (N110, N6, N62, N61);
buf BUF1 (N111, N102);
and AND4 (N112, N81, N79, N41, N47);
and AND3 (N113, N106, N73, N60);
nand NAND4 (N114, N95, N77, N30, N4);
and AND2 (N115, N111, N41);
xor XOR2 (N116, N109, N73);
nor NOR2 (N117, N107, N7);
buf BUF1 (N118, N99);
xor XOR2 (N119, N113, N5);
xor XOR2 (N120, N117, N67);
or OR2 (N121, N112, N32);
buf BUF1 (N122, N115);
buf BUF1 (N123, N100);
xor XOR2 (N124, N122, N72);
nand NAND2 (N125, N116, N110);
nor NOR3 (N126, N30, N69, N11);
and AND3 (N127, N105, N78, N13);
and AND2 (N128, N127, N78);
buf BUF1 (N129, N118);
and AND4 (N130, N119, N92, N16, N47);
xor XOR2 (N131, N124, N47);
not NOT1 (N132, N126);
not NOT1 (N133, N123);
nand NAND2 (N134, N131, N45);
or OR3 (N135, N121, N123, N17);
not NOT1 (N136, N133);
nand NAND4 (N137, N128, N53, N85, N63);
and AND3 (N138, N125, N81, N10);
nor NOR2 (N139, N129, N86);
xor XOR2 (N140, N130, N104);
nor NOR2 (N141, N114, N85);
buf BUF1 (N142, N139);
or OR3 (N143, N135, N61, N71);
xor XOR2 (N144, N138, N5);
or OR3 (N145, N143, N131, N100);
nor NOR3 (N146, N137, N56, N87);
nor NOR2 (N147, N141, N7);
nor NOR4 (N148, N132, N98, N58, N107);
nor NOR2 (N149, N136, N51);
buf BUF1 (N150, N149);
buf BUF1 (N151, N146);
nor NOR3 (N152, N145, N11, N25);
or OR3 (N153, N120, N20, N112);
not NOT1 (N154, N151);
not NOT1 (N155, N153);
and AND3 (N156, N134, N147, N144);
or OR4 (N157, N37, N14, N85, N34);
buf BUF1 (N158, N89);
or OR3 (N159, N148, N134, N9);
nand NAND4 (N160, N158, N30, N86, N94);
nor NOR3 (N161, N142, N52, N53);
or OR4 (N162, N155, N7, N142, N83);
and AND2 (N163, N156, N126);
nor NOR4 (N164, N160, N58, N130, N76);
not NOT1 (N165, N159);
not NOT1 (N166, N157);
nand NAND2 (N167, N150, N36);
nor NOR2 (N168, N152, N131);
and AND3 (N169, N167, N106, N37);
buf BUF1 (N170, N162);
nor NOR3 (N171, N164, N24, N141);
or OR3 (N172, N166, N81, N18);
and AND2 (N173, N171, N68);
or OR4 (N174, N169, N140, N172, N84);
xor XOR2 (N175, N18, N85);
and AND2 (N176, N34, N125);
nor NOR2 (N177, N170, N17);
or OR2 (N178, N161, N105);
xor XOR2 (N179, N174, N83);
nand NAND3 (N180, N175, N39, N165);
or OR3 (N181, N101, N144, N120);
or OR3 (N182, N176, N43, N37);
xor XOR2 (N183, N180, N166);
nor NOR4 (N184, N182, N91, N106, N97);
or OR3 (N185, N183, N122, N77);
buf BUF1 (N186, N154);
nor NOR3 (N187, N178, N93, N164);
nand NAND3 (N188, N186, N54, N80);
or OR4 (N189, N181, N20, N182, N77);
or OR2 (N190, N187, N44);
nand NAND2 (N191, N168, N102);
and AND2 (N192, N191, N63);
buf BUF1 (N193, N192);
nand NAND3 (N194, N185, N51, N36);
or OR4 (N195, N193, N86, N181, N185);
not NOT1 (N196, N163);
xor XOR2 (N197, N195, N151);
not NOT1 (N198, N188);
nand NAND4 (N199, N196, N151, N2, N127);
nor NOR2 (N200, N184, N138);
or OR4 (N201, N199, N34, N89, N47);
xor XOR2 (N202, N190, N36);
xor XOR2 (N203, N177, N115);
nor NOR2 (N204, N198, N88);
nor NOR3 (N205, N201, N167, N106);
nand NAND2 (N206, N179, N176);
nand NAND4 (N207, N197, N172, N149, N102);
nand NAND2 (N208, N173, N118);
nor NOR4 (N209, N208, N193, N192, N135);
buf BUF1 (N210, N204);
and AND4 (N211, N189, N64, N137, N5);
nand NAND3 (N212, N203, N162, N123);
and AND2 (N213, N205, N22);
or OR4 (N214, N206, N196, N139, N47);
buf BUF1 (N215, N209);
xor XOR2 (N216, N211, N137);
or OR3 (N217, N207, N7, N15);
nor NOR2 (N218, N212, N111);
nand NAND2 (N219, N194, N216);
xor XOR2 (N220, N102, N134);
and AND4 (N221, N213, N155, N78, N8);
xor XOR2 (N222, N215, N95);
or OR4 (N223, N219, N182, N162, N97);
nor NOR4 (N224, N223, N196, N170, N202);
not NOT1 (N225, N37);
buf BUF1 (N226, N225);
or OR4 (N227, N214, N18, N83, N16);
nand NAND4 (N228, N220, N209, N184, N222);
and AND4 (N229, N198, N172, N177, N138);
and AND3 (N230, N221, N219, N140);
and AND2 (N231, N210, N218);
nor NOR4 (N232, N201, N14, N120, N199);
nand NAND3 (N233, N224, N221, N8);
buf BUF1 (N234, N200);
nand NAND2 (N235, N230, N104);
buf BUF1 (N236, N226);
buf BUF1 (N237, N236);
buf BUF1 (N238, N237);
and AND4 (N239, N229, N97, N179, N148);
or OR4 (N240, N217, N217, N7, N43);
or OR2 (N241, N238, N215);
nand NAND4 (N242, N232, N142, N119, N117);
and AND2 (N243, N239, N43);
not NOT1 (N244, N240);
nand NAND2 (N245, N234, N26);
nand NAND4 (N246, N233, N208, N216, N200);
not NOT1 (N247, N245);
xor XOR2 (N248, N246, N75);
xor XOR2 (N249, N228, N221);
buf BUF1 (N250, N241);
nand NAND3 (N251, N244, N73, N170);
or OR3 (N252, N247, N86, N53);
and AND3 (N253, N235, N231, N249);
nor NOR3 (N254, N63, N178, N101);
and AND2 (N255, N125, N118);
nand NAND3 (N256, N253, N239, N165);
and AND2 (N257, N243, N114);
nor NOR2 (N258, N250, N56);
and AND4 (N259, N257, N204, N142, N32);
nor NOR3 (N260, N258, N179, N127);
nand NAND4 (N261, N254, N141, N99, N201);
and AND2 (N262, N255, N35);
or OR3 (N263, N260, N133, N111);
and AND2 (N264, N251, N175);
and AND4 (N265, N261, N163, N238, N257);
nor NOR2 (N266, N248, N51);
nand NAND4 (N267, N264, N247, N52, N130);
xor XOR2 (N268, N259, N221);
or OR4 (N269, N267, N52, N160, N131);
nand NAND4 (N270, N265, N147, N69, N49);
or OR4 (N271, N270, N40, N71, N114);
and AND2 (N272, N227, N55);
buf BUF1 (N273, N271);
not NOT1 (N274, N242);
buf BUF1 (N275, N252);
nand NAND2 (N276, N262, N3);
xor XOR2 (N277, N273, N35);
nand NAND3 (N278, N275, N168, N143);
xor XOR2 (N279, N278, N223);
xor XOR2 (N280, N263, N54);
nor NOR4 (N281, N274, N179, N60, N201);
nor NOR3 (N282, N268, N87, N47);
nor NOR2 (N283, N272, N55);
or OR3 (N284, N277, N280, N106);
nand NAND2 (N285, N140, N266);
nor NOR3 (N286, N229, N213, N153);
xor XOR2 (N287, N283, N212);
not NOT1 (N288, N286);
or OR2 (N289, N284, N266);
not NOT1 (N290, N285);
nand NAND3 (N291, N279, N248, N51);
buf BUF1 (N292, N276);
and AND3 (N293, N290, N123, N203);
nor NOR4 (N294, N287, N103, N25, N37);
buf BUF1 (N295, N291);
not NOT1 (N296, N269);
nor NOR2 (N297, N293, N194);
nor NOR4 (N298, N282, N176, N12, N86);
xor XOR2 (N299, N294, N116);
buf BUF1 (N300, N288);
xor XOR2 (N301, N256, N155);
nand NAND4 (N302, N289, N233, N239, N192);
or OR2 (N303, N301, N50);
xor XOR2 (N304, N300, N165);
or OR3 (N305, N299, N124, N229);
nand NAND2 (N306, N304, N173);
or OR2 (N307, N306, N20);
not NOT1 (N308, N305);
not NOT1 (N309, N281);
and AND3 (N310, N297, N300, N122);
nand NAND3 (N311, N296, N63, N22);
nand NAND3 (N312, N292, N175, N157);
and AND3 (N313, N308, N236, N94);
xor XOR2 (N314, N310, N159);
nand NAND3 (N315, N313, N234, N73);
xor XOR2 (N316, N314, N175);
or OR4 (N317, N303, N268, N227, N88);
or OR2 (N318, N302, N228);
not NOT1 (N319, N298);
or OR2 (N320, N307, N142);
xor XOR2 (N321, N317, N62);
nor NOR4 (N322, N320, N243, N176, N67);
nand NAND4 (N323, N319, N155, N172, N199);
buf BUF1 (N324, N295);
not NOT1 (N325, N323);
or OR3 (N326, N311, N291, N223);
nand NAND2 (N327, N322, N8);
buf BUF1 (N328, N309);
buf BUF1 (N329, N315);
nor NOR2 (N330, N318, N266);
and AND3 (N331, N325, N183, N167);
nor NOR4 (N332, N328, N236, N317, N261);
nor NOR4 (N333, N327, N230, N314, N279);
xor XOR2 (N334, N331, N325);
xor XOR2 (N335, N326, N109);
xor XOR2 (N336, N335, N130);
not NOT1 (N337, N330);
buf BUF1 (N338, N316);
or OR2 (N339, N324, N164);
and AND3 (N340, N329, N36, N32);
nand NAND3 (N341, N321, N308, N21);
buf BUF1 (N342, N312);
and AND2 (N343, N342, N213);
not NOT1 (N344, N337);
or OR2 (N345, N336, N39);
and AND2 (N346, N343, N289);
not NOT1 (N347, N332);
nand NAND2 (N348, N346, N67);
and AND3 (N349, N334, N88, N144);
nand NAND4 (N350, N348, N220, N218, N302);
buf BUF1 (N351, N344);
nor NOR4 (N352, N338, N243, N28, N120);
buf BUF1 (N353, N339);
nor NOR3 (N354, N349, N89, N41);
xor XOR2 (N355, N352, N180);
not NOT1 (N356, N354);
nor NOR3 (N357, N333, N102, N3);
nor NOR3 (N358, N341, N63, N352);
and AND3 (N359, N353, N103, N328);
or OR4 (N360, N355, N206, N125, N329);
and AND3 (N361, N351, N215, N351);
and AND2 (N362, N361, N54);
nor NOR3 (N363, N340, N15, N272);
and AND2 (N364, N357, N75);
xor XOR2 (N365, N356, N228);
buf BUF1 (N366, N350);
and AND2 (N367, N358, N330);
or OR2 (N368, N363, N39);
and AND2 (N369, N345, N139);
or OR4 (N370, N362, N117, N35, N4);
nor NOR2 (N371, N366, N104);
nand NAND4 (N372, N360, N331, N314, N194);
and AND2 (N373, N367, N142);
or OR4 (N374, N371, N52, N281, N147);
buf BUF1 (N375, N370);
xor XOR2 (N376, N373, N311);
xor XOR2 (N377, N374, N199);
not NOT1 (N378, N372);
buf BUF1 (N379, N369);
not NOT1 (N380, N376);
nor NOR4 (N381, N378, N76, N157, N319);
nand NAND4 (N382, N359, N213, N110, N65);
buf BUF1 (N383, N347);
not NOT1 (N384, N381);
not NOT1 (N385, N379);
or OR4 (N386, N380, N149, N367, N244);
or OR3 (N387, N377, N250, N102);
or OR4 (N388, N365, N98, N283, N94);
nand NAND3 (N389, N368, N144, N112);
or OR2 (N390, N384, N180);
not NOT1 (N391, N386);
nand NAND3 (N392, N383, N337, N133);
nand NAND4 (N393, N388, N347, N41, N116);
or OR4 (N394, N393, N220, N149, N223);
or OR4 (N395, N392, N5, N56, N47);
not NOT1 (N396, N391);
and AND3 (N397, N396, N364, N162);
buf BUF1 (N398, N5);
xor XOR2 (N399, N394, N393);
buf BUF1 (N400, N399);
buf BUF1 (N401, N385);
nand NAND3 (N402, N390, N306, N335);
xor XOR2 (N403, N401, N301);
not NOT1 (N404, N400);
xor XOR2 (N405, N403, N378);
xor XOR2 (N406, N398, N267);
nand NAND4 (N407, N406, N264, N57, N94);
not NOT1 (N408, N397);
nor NOR4 (N409, N382, N284, N78, N81);
nor NOR2 (N410, N405, N188);
buf BUF1 (N411, N402);
not NOT1 (N412, N395);
xor XOR2 (N413, N375, N115);
and AND2 (N414, N410, N112);
xor XOR2 (N415, N409, N162);
nor NOR4 (N416, N404, N46, N163, N88);
and AND2 (N417, N412, N377);
and AND4 (N418, N411, N280, N213, N338);
nand NAND3 (N419, N407, N221, N8);
not NOT1 (N420, N417);
nand NAND4 (N421, N389, N304, N294, N98);
nor NOR4 (N422, N387, N50, N413, N394);
buf BUF1 (N423, N151);
endmodule