// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N2011,N2005,N2020,N2022,N2018,N2023,N2021,N2016,N2009,N2024;

nor NOR3 (N25, N13, N14, N6);
xor XOR2 (N26, N17, N15);
nand NAND3 (N27, N24, N25, N15);
nor NOR3 (N28, N8, N19, N13);
or OR2 (N29, N24, N28);
and AND3 (N30, N3, N5, N15);
not NOT1 (N31, N22);
or OR3 (N32, N31, N26, N14);
xor XOR2 (N33, N5, N15);
nor NOR3 (N34, N28, N17, N8);
and AND2 (N35, N5, N31);
buf BUF1 (N36, N12);
buf BUF1 (N37, N18);
nor NOR2 (N38, N3, N10);
and AND3 (N39, N37, N30, N8);
nor NOR2 (N40, N23, N1);
not NOT1 (N41, N40);
xor XOR2 (N42, N34, N19);
xor XOR2 (N43, N33, N41);
xor XOR2 (N44, N33, N42);
or OR4 (N45, N12, N39, N20, N21);
not NOT1 (N46, N8);
buf BUF1 (N47, N27);
xor XOR2 (N48, N43, N42);
buf BUF1 (N49, N44);
buf BUF1 (N50, N29);
not NOT1 (N51, N45);
not NOT1 (N52, N32);
buf BUF1 (N53, N38);
or OR3 (N54, N47, N37, N7);
and AND3 (N55, N49, N53, N8);
and AND4 (N56, N33, N49, N17, N26);
nor NOR3 (N57, N48, N3, N27);
and AND4 (N58, N35, N41, N15, N56);
not NOT1 (N59, N53);
xor XOR2 (N60, N52, N38);
xor XOR2 (N61, N55, N39);
xor XOR2 (N62, N50, N15);
not NOT1 (N63, N62);
nor NOR3 (N64, N51, N57, N22);
buf BUF1 (N65, N62);
xor XOR2 (N66, N46, N19);
not NOT1 (N67, N66);
nor NOR3 (N68, N60, N48, N32);
or OR4 (N69, N61, N8, N48, N24);
not NOT1 (N70, N63);
nor NOR4 (N71, N70, N52, N68, N3);
nor NOR3 (N72, N32, N53, N57);
not NOT1 (N73, N71);
nor NOR4 (N74, N72, N50, N60, N69);
or OR2 (N75, N22, N73);
xor XOR2 (N76, N57, N3);
not NOT1 (N77, N64);
not NOT1 (N78, N59);
and AND2 (N79, N65, N71);
or OR3 (N80, N67, N53, N19);
nand NAND2 (N81, N79, N17);
buf BUF1 (N82, N54);
or OR2 (N83, N76, N63);
nor NOR4 (N84, N74, N12, N44, N15);
buf BUF1 (N85, N84);
nand NAND3 (N86, N80, N73, N55);
buf BUF1 (N87, N36);
buf BUF1 (N88, N81);
and AND4 (N89, N82, N10, N34, N48);
and AND3 (N90, N58, N74, N28);
or OR3 (N91, N78, N15, N6);
nor NOR3 (N92, N89, N32, N53);
nand NAND4 (N93, N75, N8, N56, N85);
buf BUF1 (N94, N46);
nand NAND2 (N95, N86, N74);
xor XOR2 (N96, N77, N30);
or OR3 (N97, N93, N54, N53);
nor NOR3 (N98, N96, N75, N33);
and AND3 (N99, N98, N4, N56);
and AND3 (N100, N91, N47, N97);
buf BUF1 (N101, N7);
xor XOR2 (N102, N87, N24);
buf BUF1 (N103, N102);
nor NOR3 (N104, N83, N27, N30);
not NOT1 (N105, N104);
nor NOR3 (N106, N101, N93, N54);
or OR4 (N107, N90, N65, N37, N87);
and AND3 (N108, N95, N93, N101);
xor XOR2 (N109, N106, N29);
or OR2 (N110, N88, N85);
and AND4 (N111, N105, N49, N47, N13);
and AND2 (N112, N111, N38);
not NOT1 (N113, N94);
nand NAND4 (N114, N99, N45, N88, N4);
buf BUF1 (N115, N92);
or OR4 (N116, N114, N80, N73, N88);
nor NOR2 (N117, N110, N112);
nor NOR2 (N118, N36, N46);
and AND4 (N119, N109, N102, N78, N6);
nand NAND4 (N120, N100, N8, N82, N67);
or OR2 (N121, N113, N2);
xor XOR2 (N122, N119, N12);
or OR4 (N123, N103, N5, N20, N74);
not NOT1 (N124, N121);
and AND4 (N125, N117, N43, N110, N99);
not NOT1 (N126, N107);
and AND3 (N127, N126, N18, N100);
nand NAND4 (N128, N120, N85, N68, N73);
buf BUF1 (N129, N124);
nor NOR4 (N130, N122, N69, N124, N54);
or OR3 (N131, N130, N41, N27);
xor XOR2 (N132, N118, N73);
buf BUF1 (N133, N115);
and AND4 (N134, N123, N4, N104, N49);
nor NOR2 (N135, N116, N35);
xor XOR2 (N136, N134, N23);
and AND4 (N137, N129, N113, N16, N24);
or OR3 (N138, N128, N22, N128);
xor XOR2 (N139, N133, N75);
not NOT1 (N140, N132);
buf BUF1 (N141, N136);
and AND4 (N142, N138, N127, N100, N101);
buf BUF1 (N143, N31);
nor NOR3 (N144, N108, N97, N98);
buf BUF1 (N145, N125);
not NOT1 (N146, N145);
xor XOR2 (N147, N140, N39);
nand NAND2 (N148, N147, N26);
or OR3 (N149, N139, N132, N98);
xor XOR2 (N150, N135, N146);
nor NOR4 (N151, N10, N102, N57, N109);
and AND2 (N152, N144, N146);
nand NAND2 (N153, N131, N81);
nand NAND4 (N154, N151, N82, N113, N42);
buf BUF1 (N155, N142);
and AND2 (N156, N150, N107);
and AND4 (N157, N149, N31, N75, N9);
not NOT1 (N158, N137);
not NOT1 (N159, N158);
buf BUF1 (N160, N153);
and AND2 (N161, N152, N63);
nor NOR3 (N162, N155, N106, N15);
nor NOR2 (N163, N156, N63);
and AND4 (N164, N141, N29, N109, N37);
nor NOR3 (N165, N143, N56, N74);
or OR3 (N166, N163, N85, N75);
nor NOR3 (N167, N148, N125, N131);
not NOT1 (N168, N157);
nand NAND3 (N169, N162, N87, N59);
not NOT1 (N170, N161);
xor XOR2 (N171, N160, N95);
and AND3 (N172, N170, N160, N101);
or OR3 (N173, N164, N24, N162);
buf BUF1 (N174, N159);
and AND4 (N175, N154, N141, N114, N172);
not NOT1 (N176, N151);
xor XOR2 (N177, N166, N10);
nor NOR4 (N178, N165, N5, N29, N44);
nor NOR3 (N179, N169, N108, N65);
nor NOR3 (N180, N179, N35, N138);
and AND4 (N181, N171, N58, N56, N40);
and AND2 (N182, N168, N156);
nor NOR2 (N183, N180, N20);
not NOT1 (N184, N175);
nor NOR2 (N185, N176, N114);
not NOT1 (N186, N167);
xor XOR2 (N187, N181, N134);
xor XOR2 (N188, N184, N77);
and AND3 (N189, N187, N61, N60);
not NOT1 (N190, N174);
xor XOR2 (N191, N183, N69);
nor NOR2 (N192, N173, N99);
not NOT1 (N193, N185);
or OR2 (N194, N182, N33);
or OR4 (N195, N178, N162, N74, N80);
or OR3 (N196, N188, N29, N144);
not NOT1 (N197, N193);
and AND4 (N198, N192, N147, N168, N145);
or OR2 (N199, N190, N184);
xor XOR2 (N200, N199, N7);
nor NOR3 (N201, N195, N8, N41);
and AND2 (N202, N189, N188);
nand NAND3 (N203, N198, N48, N42);
and AND2 (N204, N201, N158);
not NOT1 (N205, N202);
or OR2 (N206, N191, N66);
and AND4 (N207, N197, N9, N120, N131);
or OR4 (N208, N200, N61, N204, N99);
nor NOR4 (N209, N11, N11, N39, N191);
not NOT1 (N210, N208);
buf BUF1 (N211, N186);
nor NOR4 (N212, N206, N17, N193, N150);
and AND3 (N213, N211, N127, N158);
buf BUF1 (N214, N205);
nor NOR4 (N215, N209, N178, N139, N23);
or OR2 (N216, N212, N67);
or OR4 (N217, N213, N131, N4, N145);
nor NOR2 (N218, N196, N212);
xor XOR2 (N219, N217, N36);
nor NOR2 (N220, N210, N113);
nand NAND2 (N221, N218, N189);
not NOT1 (N222, N207);
buf BUF1 (N223, N177);
not NOT1 (N224, N215);
nand NAND2 (N225, N224, N91);
buf BUF1 (N226, N222);
buf BUF1 (N227, N221);
nand NAND4 (N228, N223, N72, N27, N120);
buf BUF1 (N229, N220);
buf BUF1 (N230, N216);
or OR4 (N231, N214, N81, N205, N220);
and AND3 (N232, N229, N5, N77);
buf BUF1 (N233, N194);
and AND4 (N234, N203, N99, N135, N46);
or OR4 (N235, N233, N61, N189, N181);
nand NAND4 (N236, N219, N63, N9, N111);
xor XOR2 (N237, N227, N64);
not NOT1 (N238, N232);
nor NOR3 (N239, N238, N115, N30);
nand NAND4 (N240, N234, N201, N144, N50);
or OR3 (N241, N228, N11, N55);
nor NOR4 (N242, N225, N12, N31, N187);
buf BUF1 (N243, N236);
nand NAND3 (N244, N231, N166, N50);
nand NAND3 (N245, N239, N82, N235);
buf BUF1 (N246, N178);
xor XOR2 (N247, N242, N206);
nor NOR2 (N248, N244, N240);
or OR2 (N249, N100, N37);
and AND2 (N250, N230, N104);
xor XOR2 (N251, N247, N48);
xor XOR2 (N252, N243, N77);
xor XOR2 (N253, N248, N57);
and AND3 (N254, N251, N175, N29);
nand NAND3 (N255, N249, N27, N249);
nand NAND3 (N256, N241, N92, N184);
nor NOR4 (N257, N245, N149, N134, N235);
nor NOR4 (N258, N252, N180, N130, N161);
xor XOR2 (N259, N257, N15);
buf BUF1 (N260, N246);
or OR2 (N261, N253, N164);
xor XOR2 (N262, N256, N44);
nor NOR2 (N263, N262, N262);
not NOT1 (N264, N237);
nor NOR3 (N265, N260, N160, N256);
xor XOR2 (N266, N255, N10);
buf BUF1 (N267, N266);
nor NOR3 (N268, N259, N232, N126);
xor XOR2 (N269, N250, N150);
xor XOR2 (N270, N264, N245);
buf BUF1 (N271, N268);
xor XOR2 (N272, N261, N150);
nor NOR3 (N273, N272, N193, N231);
and AND4 (N274, N254, N178, N147, N95);
nand NAND4 (N275, N270, N235, N209, N74);
nor NOR3 (N276, N258, N34, N89);
nor NOR3 (N277, N226, N32, N27);
or OR3 (N278, N269, N147, N184);
not NOT1 (N279, N278);
nor NOR2 (N280, N277, N30);
and AND3 (N281, N275, N20, N182);
not NOT1 (N282, N267);
and AND4 (N283, N265, N41, N194, N134);
nand NAND4 (N284, N271, N15, N267, N199);
nand NAND2 (N285, N274, N143);
nor NOR2 (N286, N284, N58);
and AND4 (N287, N285, N134, N74, N276);
or OR2 (N288, N56, N222);
xor XOR2 (N289, N263, N54);
and AND3 (N290, N282, N247, N164);
not NOT1 (N291, N289);
or OR4 (N292, N290, N166, N265, N155);
nor NOR4 (N293, N288, N190, N112, N146);
xor XOR2 (N294, N287, N8);
and AND2 (N295, N283, N19);
not NOT1 (N296, N294);
xor XOR2 (N297, N293, N169);
nand NAND4 (N298, N281, N97, N67, N65);
buf BUF1 (N299, N296);
nor NOR3 (N300, N279, N212, N255);
nand NAND2 (N301, N295, N105);
xor XOR2 (N302, N301, N39);
and AND2 (N303, N302, N164);
and AND3 (N304, N300, N68, N90);
buf BUF1 (N305, N273);
nand NAND2 (N306, N292, N246);
or OR3 (N307, N280, N136, N86);
buf BUF1 (N308, N298);
buf BUF1 (N309, N305);
or OR2 (N310, N299, N279);
xor XOR2 (N311, N307, N286);
buf BUF1 (N312, N145);
not NOT1 (N313, N309);
nand NAND2 (N314, N306, N77);
and AND3 (N315, N291, N165, N127);
nor NOR2 (N316, N315, N313);
not NOT1 (N317, N267);
or OR3 (N318, N303, N213, N310);
and AND2 (N319, N187, N222);
not NOT1 (N320, N311);
or OR3 (N321, N316, N186, N184);
xor XOR2 (N322, N308, N99);
xor XOR2 (N323, N314, N102);
buf BUF1 (N324, N321);
nor NOR4 (N325, N320, N55, N194, N218);
nand NAND4 (N326, N325, N19, N113, N185);
and AND2 (N327, N297, N59);
buf BUF1 (N328, N304);
nand NAND3 (N329, N323, N260, N119);
buf BUF1 (N330, N324);
nor NOR2 (N331, N326, N166);
not NOT1 (N332, N331);
not NOT1 (N333, N329);
xor XOR2 (N334, N317, N55);
nand NAND4 (N335, N330, N169, N248, N69);
nand NAND4 (N336, N333, N114, N325, N37);
nor NOR4 (N337, N334, N6, N75, N299);
xor XOR2 (N338, N327, N91);
nor NOR2 (N339, N318, N96);
buf BUF1 (N340, N339);
nand NAND2 (N341, N322, N26);
and AND3 (N342, N332, N178, N220);
or OR3 (N343, N337, N207, N248);
nor NOR2 (N344, N319, N285);
nand NAND2 (N345, N340, N131);
not NOT1 (N346, N328);
not NOT1 (N347, N342);
or OR4 (N348, N336, N45, N316, N250);
not NOT1 (N349, N312);
nand NAND2 (N350, N341, N52);
nor NOR4 (N351, N338, N266, N288, N261);
nand NAND4 (N352, N343, N31, N5, N83);
or OR2 (N353, N347, N208);
xor XOR2 (N354, N346, N144);
not NOT1 (N355, N348);
not NOT1 (N356, N354);
or OR2 (N357, N352, N191);
nand NAND4 (N358, N349, N60, N74, N188);
nand NAND3 (N359, N353, N228, N66);
nor NOR3 (N360, N358, N7, N23);
or OR2 (N361, N344, N356);
or OR3 (N362, N214, N157, N28);
and AND3 (N363, N345, N266, N98);
buf BUF1 (N364, N357);
not NOT1 (N365, N360);
buf BUF1 (N366, N363);
nor NOR4 (N367, N351, N207, N20, N28);
buf BUF1 (N368, N365);
nand NAND2 (N369, N364, N214);
xor XOR2 (N370, N350, N292);
and AND4 (N371, N359, N68, N87, N195);
nor NOR4 (N372, N368, N67, N328, N36);
and AND3 (N373, N372, N157, N106);
buf BUF1 (N374, N369);
nor NOR4 (N375, N373, N324, N198, N211);
not NOT1 (N376, N335);
nor NOR2 (N377, N376, N327);
and AND3 (N378, N375, N306, N309);
or OR3 (N379, N378, N178, N190);
buf BUF1 (N380, N361);
buf BUF1 (N381, N374);
and AND4 (N382, N370, N362, N232, N3);
and AND3 (N383, N232, N20, N151);
or OR4 (N384, N382, N131, N89, N342);
or OR3 (N385, N366, N168, N36);
not NOT1 (N386, N381);
buf BUF1 (N387, N355);
not NOT1 (N388, N385);
not NOT1 (N389, N387);
buf BUF1 (N390, N379);
buf BUF1 (N391, N371);
nor NOR4 (N392, N386, N377, N373, N239);
or OR2 (N393, N282, N87);
nand NAND3 (N394, N388, N214, N112);
nand NAND2 (N395, N393, N70);
not NOT1 (N396, N383);
nand NAND2 (N397, N396, N349);
buf BUF1 (N398, N390);
not NOT1 (N399, N395);
not NOT1 (N400, N384);
and AND2 (N401, N398, N10);
not NOT1 (N402, N380);
buf BUF1 (N403, N391);
nand NAND4 (N404, N403, N232, N36, N384);
or OR4 (N405, N397, N308, N209, N319);
not NOT1 (N406, N394);
buf BUF1 (N407, N389);
or OR4 (N408, N401, N209, N279, N166);
or OR4 (N409, N407, N264, N53, N208);
buf BUF1 (N410, N408);
buf BUF1 (N411, N404);
buf BUF1 (N412, N409);
or OR2 (N413, N402, N291);
xor XOR2 (N414, N392, N126);
buf BUF1 (N415, N410);
xor XOR2 (N416, N412, N220);
and AND2 (N417, N411, N172);
and AND4 (N418, N413, N279, N226, N21);
and AND2 (N419, N417, N389);
nor NOR3 (N420, N406, N399, N217);
or OR3 (N421, N254, N158, N147);
xor XOR2 (N422, N419, N94);
xor XOR2 (N423, N422, N3);
nor NOR4 (N424, N405, N336, N145, N237);
not NOT1 (N425, N424);
nand NAND4 (N426, N418, N22, N365, N150);
or OR3 (N427, N415, N176, N320);
xor XOR2 (N428, N416, N110);
or OR3 (N429, N428, N376, N55);
nand NAND4 (N430, N421, N429, N136, N411);
buf BUF1 (N431, N115);
buf BUF1 (N432, N427);
xor XOR2 (N433, N432, N18);
buf BUF1 (N434, N426);
or OR2 (N435, N433, N221);
or OR4 (N436, N367, N23, N394, N208);
or OR2 (N437, N431, N155);
buf BUF1 (N438, N425);
or OR4 (N439, N434, N233, N378, N431);
or OR3 (N440, N423, N112, N319);
buf BUF1 (N441, N430);
xor XOR2 (N442, N441, N272);
buf BUF1 (N443, N436);
and AND4 (N444, N443, N144, N60, N100);
not NOT1 (N445, N442);
and AND3 (N446, N400, N384, N174);
nor NOR2 (N447, N420, N275);
nor NOR3 (N448, N440, N339, N75);
not NOT1 (N449, N414);
not NOT1 (N450, N446);
xor XOR2 (N451, N439, N142);
or OR4 (N452, N445, N199, N359, N355);
buf BUF1 (N453, N452);
not NOT1 (N454, N444);
nor NOR4 (N455, N437, N294, N49, N62);
nand NAND4 (N456, N454, N419, N244, N407);
and AND4 (N457, N450, N76, N7, N428);
nor NOR3 (N458, N449, N168, N43);
xor XOR2 (N459, N438, N414);
buf BUF1 (N460, N456);
nor NOR2 (N461, N447, N312);
and AND2 (N462, N451, N40);
nand NAND3 (N463, N457, N281, N29);
buf BUF1 (N464, N458);
and AND4 (N465, N435, N45, N142, N59);
xor XOR2 (N466, N455, N290);
xor XOR2 (N467, N466, N322);
not NOT1 (N468, N467);
nor NOR4 (N469, N453, N147, N9, N253);
and AND2 (N470, N465, N198);
xor XOR2 (N471, N460, N399);
and AND4 (N472, N463, N433, N395, N377);
or OR2 (N473, N461, N111);
buf BUF1 (N474, N472);
not NOT1 (N475, N468);
or OR2 (N476, N448, N398);
or OR4 (N477, N469, N94, N138, N155);
buf BUF1 (N478, N474);
and AND3 (N479, N475, N196, N121);
or OR2 (N480, N476, N380);
and AND4 (N481, N462, N170, N183, N89);
nor NOR3 (N482, N480, N52, N431);
nor NOR4 (N483, N459, N14, N300, N76);
not NOT1 (N484, N481);
or OR2 (N485, N470, N53);
or OR3 (N486, N482, N415, N334);
nor NOR3 (N487, N486, N328, N327);
nand NAND4 (N488, N464, N453, N355, N302);
not NOT1 (N489, N471);
buf BUF1 (N490, N479);
nor NOR2 (N491, N489, N264);
and AND3 (N492, N490, N187, N172);
buf BUF1 (N493, N492);
nor NOR4 (N494, N493, N200, N21, N304);
nand NAND3 (N495, N478, N142, N98);
nor NOR4 (N496, N473, N307, N213, N415);
buf BUF1 (N497, N485);
buf BUF1 (N498, N497);
not NOT1 (N499, N484);
xor XOR2 (N500, N499, N149);
and AND3 (N501, N494, N23, N389);
buf BUF1 (N502, N483);
nor NOR4 (N503, N491, N156, N496, N450);
nand NAND3 (N504, N141, N5, N37);
and AND3 (N505, N488, N91, N381);
nand NAND3 (N506, N477, N446, N490);
nor NOR4 (N507, N504, N299, N149, N374);
and AND3 (N508, N498, N105, N297);
not NOT1 (N509, N487);
nand NAND4 (N510, N505, N432, N490, N70);
not NOT1 (N511, N507);
nor NOR4 (N512, N503, N319, N96, N156);
and AND3 (N513, N512, N358, N439);
nand NAND3 (N514, N513, N231, N308);
buf BUF1 (N515, N510);
nand NAND3 (N516, N506, N336, N119);
buf BUF1 (N517, N501);
nand NAND4 (N518, N502, N175, N159, N255);
not NOT1 (N519, N500);
and AND4 (N520, N514, N135, N210, N59);
nor NOR3 (N521, N519, N421, N168);
nor NOR2 (N522, N516, N468);
nand NAND4 (N523, N515, N142, N274, N215);
xor XOR2 (N524, N518, N100);
buf BUF1 (N525, N517);
or OR4 (N526, N495, N42, N157, N33);
and AND2 (N527, N511, N88);
not NOT1 (N528, N527);
xor XOR2 (N529, N508, N87);
and AND3 (N530, N522, N383, N85);
nand NAND4 (N531, N509, N225, N43, N404);
xor XOR2 (N532, N528, N5);
or OR2 (N533, N531, N365);
xor XOR2 (N534, N524, N408);
buf BUF1 (N535, N532);
and AND4 (N536, N521, N329, N35, N5);
nand NAND4 (N537, N523, N496, N159, N66);
not NOT1 (N538, N529);
xor XOR2 (N539, N537, N418);
and AND3 (N540, N526, N238, N462);
buf BUF1 (N541, N539);
xor XOR2 (N542, N538, N270);
or OR2 (N543, N530, N188);
xor XOR2 (N544, N525, N306);
nand NAND3 (N545, N520, N425, N144);
nand NAND4 (N546, N536, N126, N287, N312);
nand NAND3 (N547, N544, N474, N179);
nand NAND4 (N548, N533, N364, N236, N286);
nand NAND3 (N549, N546, N25, N294);
not NOT1 (N550, N534);
or OR2 (N551, N548, N51);
xor XOR2 (N552, N540, N152);
xor XOR2 (N553, N551, N103);
or OR2 (N554, N543, N248);
nand NAND2 (N555, N535, N22);
nand NAND4 (N556, N554, N514, N361, N246);
xor XOR2 (N557, N556, N470);
not NOT1 (N558, N542);
and AND2 (N559, N541, N205);
nor NOR4 (N560, N547, N71, N123, N285);
nor NOR2 (N561, N552, N328);
xor XOR2 (N562, N553, N132);
and AND4 (N563, N562, N550, N483, N320);
buf BUF1 (N564, N360);
not NOT1 (N565, N549);
not NOT1 (N566, N557);
and AND3 (N567, N559, N476, N372);
buf BUF1 (N568, N567);
not NOT1 (N569, N558);
buf BUF1 (N570, N565);
not NOT1 (N571, N564);
xor XOR2 (N572, N566, N118);
nand NAND2 (N573, N571, N247);
nor NOR3 (N574, N568, N4, N321);
buf BUF1 (N575, N573);
or OR4 (N576, N572, N86, N424, N299);
or OR2 (N577, N555, N248);
or OR4 (N578, N574, N292, N82, N215);
and AND3 (N579, N570, N286, N229);
nand NAND4 (N580, N578, N381, N494, N13);
buf BUF1 (N581, N580);
buf BUF1 (N582, N577);
or OR3 (N583, N579, N393, N58);
nor NOR2 (N584, N576, N2);
buf BUF1 (N585, N575);
xor XOR2 (N586, N561, N30);
buf BUF1 (N587, N585);
nand NAND4 (N588, N587, N577, N547, N155);
buf BUF1 (N589, N583);
not NOT1 (N590, N588);
or OR4 (N591, N582, N58, N560, N289);
nor NOR2 (N592, N529, N563);
nand NAND2 (N593, N407, N265);
or OR3 (N594, N591, N346, N367);
not NOT1 (N595, N584);
not NOT1 (N596, N586);
buf BUF1 (N597, N581);
or OR4 (N598, N592, N228, N125, N328);
not NOT1 (N599, N590);
nand NAND2 (N600, N589, N589);
buf BUF1 (N601, N599);
nor NOR3 (N602, N600, N157, N390);
buf BUF1 (N603, N594);
not NOT1 (N604, N602);
not NOT1 (N605, N597);
nand NAND4 (N606, N569, N193, N221, N516);
xor XOR2 (N607, N605, N319);
buf BUF1 (N608, N593);
nand NAND4 (N609, N607, N445, N46, N221);
nand NAND2 (N610, N609, N350);
and AND4 (N611, N595, N544, N195, N488);
xor XOR2 (N612, N545, N243);
and AND2 (N613, N608, N21);
and AND2 (N614, N598, N41);
or OR3 (N615, N606, N323, N546);
not NOT1 (N616, N613);
buf BUF1 (N617, N601);
not NOT1 (N618, N603);
nor NOR3 (N619, N618, N324, N194);
nor NOR4 (N620, N596, N328, N405, N48);
buf BUF1 (N621, N610);
nor NOR3 (N622, N614, N34, N564);
xor XOR2 (N623, N619, N250);
xor XOR2 (N624, N612, N330);
xor XOR2 (N625, N617, N328);
buf BUF1 (N626, N616);
nand NAND3 (N627, N620, N121, N138);
buf BUF1 (N628, N621);
nand NAND2 (N629, N625, N275);
and AND4 (N630, N604, N47, N372, N553);
buf BUF1 (N631, N628);
buf BUF1 (N632, N611);
not NOT1 (N633, N631);
buf BUF1 (N634, N622);
not NOT1 (N635, N632);
nor NOR4 (N636, N634, N130, N201, N87);
buf BUF1 (N637, N630);
or OR2 (N638, N624, N577);
nand NAND4 (N639, N636, N410, N425, N30);
not NOT1 (N640, N615);
xor XOR2 (N641, N623, N260);
buf BUF1 (N642, N637);
and AND4 (N643, N629, N329, N36, N63);
nor NOR4 (N644, N626, N168, N28, N615);
not NOT1 (N645, N639);
and AND4 (N646, N635, N378, N230, N153);
xor XOR2 (N647, N641, N275);
or OR2 (N648, N643, N173);
and AND2 (N649, N644, N249);
nand NAND4 (N650, N649, N606, N470, N544);
buf BUF1 (N651, N650);
and AND3 (N652, N645, N369, N268);
buf BUF1 (N653, N648);
buf BUF1 (N654, N640);
xor XOR2 (N655, N651, N133);
buf BUF1 (N656, N633);
or OR3 (N657, N652, N4, N503);
nand NAND3 (N658, N653, N35, N132);
and AND3 (N659, N656, N531, N458);
or OR3 (N660, N658, N212, N54);
and AND4 (N661, N655, N157, N455, N138);
xor XOR2 (N662, N647, N608);
buf BUF1 (N663, N654);
not NOT1 (N664, N662);
or OR2 (N665, N657, N442);
nand NAND2 (N666, N661, N519);
not NOT1 (N667, N660);
xor XOR2 (N668, N663, N267);
nand NAND2 (N669, N642, N572);
not NOT1 (N670, N646);
nand NAND4 (N671, N670, N444, N68, N3);
xor XOR2 (N672, N659, N237);
buf BUF1 (N673, N668);
and AND2 (N674, N664, N23);
or OR4 (N675, N671, N89, N633, N184);
buf BUF1 (N676, N627);
and AND2 (N677, N672, N224);
buf BUF1 (N678, N667);
nand NAND4 (N679, N669, N441, N606, N401);
not NOT1 (N680, N638);
nand NAND4 (N681, N680, N635, N229, N609);
nor NOR3 (N682, N665, N144, N473);
buf BUF1 (N683, N673);
xor XOR2 (N684, N679, N145);
nor NOR3 (N685, N677, N614, N68);
xor XOR2 (N686, N681, N510);
not NOT1 (N687, N666);
nand NAND3 (N688, N678, N204, N299);
not NOT1 (N689, N686);
or OR2 (N690, N674, N301);
nand NAND3 (N691, N690, N134, N491);
not NOT1 (N692, N685);
xor XOR2 (N693, N675, N622);
xor XOR2 (N694, N693, N310);
nand NAND3 (N695, N684, N232, N289);
buf BUF1 (N696, N689);
nor NOR2 (N697, N688, N120);
nand NAND4 (N698, N697, N439, N177, N370);
or OR3 (N699, N682, N449, N493);
nand NAND2 (N700, N699, N238);
nor NOR2 (N701, N694, N190);
and AND4 (N702, N692, N221, N200, N477);
nor NOR2 (N703, N702, N25);
not NOT1 (N704, N687);
nand NAND2 (N705, N695, N204);
xor XOR2 (N706, N705, N424);
buf BUF1 (N707, N691);
buf BUF1 (N708, N698);
nand NAND2 (N709, N704, N590);
xor XOR2 (N710, N701, N40);
or OR4 (N711, N709, N168, N422, N412);
nor NOR4 (N712, N696, N145, N559, N649);
and AND2 (N713, N707, N705);
nor NOR2 (N714, N683, N454);
not NOT1 (N715, N714);
nand NAND3 (N716, N706, N303, N423);
and AND2 (N717, N715, N307);
nand NAND3 (N718, N710, N710, N536);
or OR4 (N719, N713, N351, N406, N680);
xor XOR2 (N720, N712, N275);
or OR3 (N721, N711, N106, N544);
xor XOR2 (N722, N720, N214);
not NOT1 (N723, N703);
not NOT1 (N724, N723);
buf BUF1 (N725, N716);
not NOT1 (N726, N722);
and AND2 (N727, N726, N321);
or OR4 (N728, N724, N533, N487, N189);
nand NAND3 (N729, N717, N502, N591);
buf BUF1 (N730, N718);
buf BUF1 (N731, N719);
xor XOR2 (N732, N727, N18);
not NOT1 (N733, N725);
nor NOR4 (N734, N730, N673, N323, N541);
and AND4 (N735, N728, N604, N27, N307);
buf BUF1 (N736, N732);
nor NOR2 (N737, N731, N690);
not NOT1 (N738, N721);
not NOT1 (N739, N736);
not NOT1 (N740, N738);
not NOT1 (N741, N739);
and AND4 (N742, N676, N234, N692, N597);
nand NAND2 (N743, N741, N521);
xor XOR2 (N744, N708, N381);
nor NOR4 (N745, N729, N584, N601, N131);
nand NAND3 (N746, N744, N237, N394);
nor NOR2 (N747, N700, N251);
xor XOR2 (N748, N746, N300);
nand NAND4 (N749, N748, N309, N429, N49);
buf BUF1 (N750, N737);
not NOT1 (N751, N749);
not NOT1 (N752, N750);
buf BUF1 (N753, N735);
or OR4 (N754, N740, N310, N527, N568);
nand NAND4 (N755, N742, N682, N121, N252);
nor NOR2 (N756, N755, N622);
nand NAND2 (N757, N751, N282);
xor XOR2 (N758, N757, N510);
xor XOR2 (N759, N747, N9);
or OR3 (N760, N753, N724, N325);
buf BUF1 (N761, N754);
or OR3 (N762, N760, N645, N133);
and AND3 (N763, N745, N630, N535);
nor NOR4 (N764, N758, N477, N99, N620);
and AND4 (N765, N761, N310, N312, N361);
xor XOR2 (N766, N765, N478);
buf BUF1 (N767, N759);
buf BUF1 (N768, N763);
not NOT1 (N769, N733);
and AND4 (N770, N756, N285, N225, N539);
xor XOR2 (N771, N743, N688);
nor NOR3 (N772, N766, N504, N425);
not NOT1 (N773, N771);
nand NAND3 (N774, N767, N239, N73);
and AND3 (N775, N769, N193, N108);
nor NOR2 (N776, N770, N393);
nor NOR2 (N777, N773, N1);
nor NOR4 (N778, N775, N59, N93, N143);
buf BUF1 (N779, N762);
xor XOR2 (N780, N734, N532);
nand NAND4 (N781, N768, N398, N339, N693);
not NOT1 (N782, N774);
and AND4 (N783, N782, N232, N680, N525);
nor NOR2 (N784, N779, N507);
nand NAND2 (N785, N784, N416);
or OR2 (N786, N778, N109);
and AND4 (N787, N781, N756, N452, N387);
or OR2 (N788, N777, N126);
buf BUF1 (N789, N776);
and AND4 (N790, N783, N642, N316, N775);
not NOT1 (N791, N786);
nor NOR3 (N792, N764, N781, N524);
or OR4 (N793, N780, N37, N78, N236);
buf BUF1 (N794, N785);
xor XOR2 (N795, N772, N229);
and AND2 (N796, N787, N713);
not NOT1 (N797, N794);
xor XOR2 (N798, N788, N696);
buf BUF1 (N799, N793);
not NOT1 (N800, N791);
xor XOR2 (N801, N798, N138);
not NOT1 (N802, N797);
buf BUF1 (N803, N795);
and AND4 (N804, N800, N588, N550, N545);
nand NAND4 (N805, N790, N31, N138, N383);
and AND2 (N806, N803, N336);
nor NOR4 (N807, N792, N415, N17, N236);
nand NAND2 (N808, N799, N525);
buf BUF1 (N809, N806);
and AND2 (N810, N796, N249);
buf BUF1 (N811, N752);
xor XOR2 (N812, N789, N336);
nor NOR3 (N813, N810, N277, N477);
nor NOR3 (N814, N802, N93, N749);
nor NOR4 (N815, N813, N394, N412, N269);
nor NOR3 (N816, N811, N5, N353);
not NOT1 (N817, N809);
and AND3 (N818, N816, N694, N624);
or OR2 (N819, N815, N189);
nor NOR2 (N820, N804, N228);
or OR2 (N821, N812, N543);
not NOT1 (N822, N820);
buf BUF1 (N823, N808);
nor NOR4 (N824, N818, N553, N211, N779);
and AND2 (N825, N817, N150);
xor XOR2 (N826, N805, N584);
xor XOR2 (N827, N814, N507);
nand NAND3 (N828, N801, N460, N635);
nor NOR2 (N829, N827, N655);
not NOT1 (N830, N826);
or OR4 (N831, N829, N525, N668, N578);
nand NAND4 (N832, N822, N791, N783, N277);
xor XOR2 (N833, N828, N792);
buf BUF1 (N834, N821);
or OR2 (N835, N823, N598);
or OR2 (N836, N831, N505);
nand NAND2 (N837, N825, N379);
nor NOR2 (N838, N824, N91);
nand NAND4 (N839, N807, N138, N142, N389);
nand NAND2 (N840, N839, N262);
nand NAND3 (N841, N830, N240, N312);
not NOT1 (N842, N832);
or OR3 (N843, N840, N305, N334);
buf BUF1 (N844, N819);
nand NAND2 (N845, N841, N636);
or OR2 (N846, N834, N707);
or OR4 (N847, N837, N564, N123, N667);
xor XOR2 (N848, N844, N336);
or OR3 (N849, N836, N621, N234);
nand NAND3 (N850, N846, N384, N35);
buf BUF1 (N851, N848);
and AND4 (N852, N842, N165, N548, N467);
buf BUF1 (N853, N835);
nor NOR4 (N854, N845, N280, N499, N429);
and AND3 (N855, N853, N339, N663);
buf BUF1 (N856, N852);
nor NOR2 (N857, N855, N333);
not NOT1 (N858, N833);
nor NOR4 (N859, N858, N158, N811, N617);
or OR4 (N860, N854, N392, N24, N306);
xor XOR2 (N861, N838, N314);
nand NAND3 (N862, N860, N674, N284);
nor NOR3 (N863, N859, N36, N42);
or OR4 (N864, N857, N708, N6, N683);
nand NAND2 (N865, N862, N689);
xor XOR2 (N866, N851, N629);
and AND4 (N867, N861, N102, N332, N391);
xor XOR2 (N868, N847, N693);
buf BUF1 (N869, N863);
and AND3 (N870, N864, N574, N826);
nor NOR4 (N871, N867, N451, N35, N417);
nand NAND3 (N872, N865, N77, N634);
xor XOR2 (N873, N868, N333);
and AND4 (N874, N870, N635, N648, N29);
and AND4 (N875, N843, N820, N186, N391);
xor XOR2 (N876, N873, N198);
nand NAND3 (N877, N874, N647, N514);
and AND4 (N878, N876, N264, N207, N503);
buf BUF1 (N879, N856);
nand NAND3 (N880, N871, N299, N681);
xor XOR2 (N881, N877, N19);
nor NOR3 (N882, N875, N831, N622);
nor NOR3 (N883, N850, N284, N775);
nand NAND4 (N884, N866, N293, N105, N530);
nor NOR2 (N885, N878, N756);
nand NAND2 (N886, N885, N111);
xor XOR2 (N887, N880, N230);
buf BUF1 (N888, N879);
not NOT1 (N889, N882);
or OR3 (N890, N887, N132, N119);
buf BUF1 (N891, N888);
and AND3 (N892, N890, N401, N443);
not NOT1 (N893, N889);
or OR3 (N894, N891, N454, N697);
and AND2 (N895, N886, N332);
and AND3 (N896, N895, N694, N712);
nand NAND4 (N897, N896, N517, N589, N863);
buf BUF1 (N898, N883);
and AND3 (N899, N898, N849, N586);
and AND3 (N900, N94, N55, N140);
xor XOR2 (N901, N869, N197);
buf BUF1 (N902, N893);
buf BUF1 (N903, N900);
xor XOR2 (N904, N903, N67);
not NOT1 (N905, N884);
buf BUF1 (N906, N899);
nor NOR4 (N907, N897, N573, N450, N797);
xor XOR2 (N908, N904, N69);
or OR4 (N909, N892, N390, N578, N533);
not NOT1 (N910, N906);
buf BUF1 (N911, N872);
buf BUF1 (N912, N911);
xor XOR2 (N913, N901, N639);
or OR2 (N914, N909, N740);
nand NAND4 (N915, N910, N301, N645, N616);
buf BUF1 (N916, N913);
and AND2 (N917, N908, N530);
buf BUF1 (N918, N894);
xor XOR2 (N919, N902, N345);
buf BUF1 (N920, N912);
nor NOR2 (N921, N916, N526);
nor NOR2 (N922, N907, N217);
or OR3 (N923, N920, N290, N161);
and AND4 (N924, N917, N68, N912, N831);
or OR2 (N925, N923, N215);
and AND4 (N926, N921, N835, N743, N590);
not NOT1 (N927, N922);
buf BUF1 (N928, N915);
nand NAND4 (N929, N918, N700, N245, N803);
not NOT1 (N930, N927);
buf BUF1 (N931, N925);
nand NAND2 (N932, N926, N163);
xor XOR2 (N933, N919, N21);
nand NAND3 (N934, N929, N166, N33);
or OR3 (N935, N933, N467, N278);
buf BUF1 (N936, N881);
or OR3 (N937, N924, N537, N81);
not NOT1 (N938, N935);
and AND3 (N939, N934, N565, N85);
xor XOR2 (N940, N932, N788);
nor NOR4 (N941, N936, N304, N637, N880);
nand NAND3 (N942, N928, N194, N735);
nand NAND3 (N943, N940, N333, N294);
buf BUF1 (N944, N914);
not NOT1 (N945, N930);
and AND3 (N946, N942, N510, N893);
nand NAND2 (N947, N941, N517);
nand NAND2 (N948, N945, N302);
nor NOR2 (N949, N943, N209);
buf BUF1 (N950, N931);
nor NOR4 (N951, N937, N242, N397, N281);
or OR3 (N952, N948, N649, N442);
nand NAND2 (N953, N950, N28);
nor NOR4 (N954, N947, N425, N139, N815);
xor XOR2 (N955, N949, N48);
nor NOR4 (N956, N905, N408, N797, N568);
or OR4 (N957, N944, N229, N365, N169);
nand NAND4 (N958, N939, N671, N466, N468);
nand NAND4 (N959, N952, N866, N868, N364);
nand NAND2 (N960, N953, N156);
and AND2 (N961, N956, N518);
not NOT1 (N962, N958);
nand NAND3 (N963, N938, N892, N81);
xor XOR2 (N964, N951, N153);
xor XOR2 (N965, N959, N814);
nor NOR3 (N966, N964, N341, N835);
not NOT1 (N967, N965);
or OR4 (N968, N954, N104, N868, N618);
buf BUF1 (N969, N955);
nand NAND3 (N970, N957, N691, N845);
nor NOR4 (N971, N968, N691, N508, N456);
xor XOR2 (N972, N961, N352);
or OR2 (N973, N960, N582);
not NOT1 (N974, N962);
nand NAND3 (N975, N972, N193, N302);
not NOT1 (N976, N973);
and AND3 (N977, N975, N595, N242);
xor XOR2 (N978, N971, N539);
nor NOR3 (N979, N966, N933, N415);
nand NAND2 (N980, N967, N30);
not NOT1 (N981, N976);
or OR3 (N982, N978, N823, N809);
or OR3 (N983, N980, N516, N75);
xor XOR2 (N984, N969, N49);
not NOT1 (N985, N974);
nor NOR4 (N986, N985, N426, N112, N417);
not NOT1 (N987, N963);
xor XOR2 (N988, N987, N946);
and AND4 (N989, N61, N807, N577, N73);
xor XOR2 (N990, N977, N335);
not NOT1 (N991, N988);
or OR4 (N992, N989, N10, N767, N937);
nand NAND3 (N993, N986, N228, N291);
xor XOR2 (N994, N970, N654);
buf BUF1 (N995, N991);
not NOT1 (N996, N981);
or OR2 (N997, N993, N536);
nor NOR3 (N998, N992, N868, N584);
buf BUF1 (N999, N990);
xor XOR2 (N1000, N979, N991);
not NOT1 (N1001, N1000);
not NOT1 (N1002, N982);
nor NOR2 (N1003, N996, N215);
nor NOR2 (N1004, N1002, N462);
nand NAND3 (N1005, N1004, N383, N850);
buf BUF1 (N1006, N997);
nor NOR4 (N1007, N995, N327, N27, N40);
buf BUF1 (N1008, N1006);
buf BUF1 (N1009, N994);
or OR3 (N1010, N1007, N574, N613);
nand NAND2 (N1011, N1010, N648);
xor XOR2 (N1012, N1005, N277);
buf BUF1 (N1013, N1001);
nand NAND4 (N1014, N1008, N971, N746, N396);
and AND4 (N1015, N1014, N930, N749, N813);
or OR4 (N1016, N984, N304, N542, N873);
or OR4 (N1017, N1012, N177, N33, N840);
xor XOR2 (N1018, N999, N993);
or OR2 (N1019, N1015, N195);
buf BUF1 (N1020, N1019);
or OR2 (N1021, N1009, N215);
nand NAND4 (N1022, N1016, N727, N79, N424);
or OR3 (N1023, N1018, N59, N304);
xor XOR2 (N1024, N1022, N476);
buf BUF1 (N1025, N1023);
or OR4 (N1026, N1017, N139, N313, N116);
nor NOR4 (N1027, N1011, N933, N419, N568);
xor XOR2 (N1028, N1025, N957);
nand NAND4 (N1029, N1024, N796, N929, N911);
not NOT1 (N1030, N1020);
not NOT1 (N1031, N998);
buf BUF1 (N1032, N1031);
nor NOR2 (N1033, N1032, N550);
buf BUF1 (N1034, N983);
nor NOR3 (N1035, N1003, N292, N695);
buf BUF1 (N1036, N1021);
xor XOR2 (N1037, N1030, N1010);
buf BUF1 (N1038, N1026);
nor NOR3 (N1039, N1036, N10, N257);
xor XOR2 (N1040, N1035, N60);
not NOT1 (N1041, N1039);
not NOT1 (N1042, N1028);
xor XOR2 (N1043, N1040, N732);
nor NOR4 (N1044, N1042, N998, N200, N1038);
nor NOR2 (N1045, N593, N264);
nand NAND2 (N1046, N1043, N990);
buf BUF1 (N1047, N1044);
nor NOR2 (N1048, N1037, N432);
xor XOR2 (N1049, N1041, N533);
nor NOR2 (N1050, N1029, N33);
xor XOR2 (N1051, N1046, N208);
not NOT1 (N1052, N1047);
and AND4 (N1053, N1013, N558, N1001, N1008);
xor XOR2 (N1054, N1049, N748);
and AND2 (N1055, N1045, N358);
buf BUF1 (N1056, N1055);
buf BUF1 (N1057, N1056);
or OR2 (N1058, N1052, N592);
not NOT1 (N1059, N1057);
nor NOR2 (N1060, N1050, N544);
xor XOR2 (N1061, N1048, N917);
not NOT1 (N1062, N1027);
nand NAND3 (N1063, N1054, N593, N244);
xor XOR2 (N1064, N1053, N1003);
xor XOR2 (N1065, N1059, N764);
buf BUF1 (N1066, N1063);
xor XOR2 (N1067, N1064, N392);
not NOT1 (N1068, N1034);
buf BUF1 (N1069, N1067);
nor NOR2 (N1070, N1051, N126);
xor XOR2 (N1071, N1061, N371);
nand NAND4 (N1072, N1070, N404, N1009, N497);
not NOT1 (N1073, N1069);
xor XOR2 (N1074, N1060, N972);
nor NOR4 (N1075, N1074, N501, N585, N342);
xor XOR2 (N1076, N1058, N1034);
and AND3 (N1077, N1075, N305, N760);
buf BUF1 (N1078, N1077);
not NOT1 (N1079, N1073);
and AND2 (N1080, N1071, N430);
and AND4 (N1081, N1079, N281, N515, N993);
nand NAND3 (N1082, N1068, N122, N961);
buf BUF1 (N1083, N1072);
xor XOR2 (N1084, N1066, N170);
not NOT1 (N1085, N1078);
nand NAND4 (N1086, N1033, N278, N666, N549);
nor NOR4 (N1087, N1065, N615, N1074, N90);
nor NOR2 (N1088, N1087, N1009);
buf BUF1 (N1089, N1085);
xor XOR2 (N1090, N1076, N361);
nand NAND4 (N1091, N1088, N257, N406, N844);
not NOT1 (N1092, N1080);
and AND2 (N1093, N1062, N292);
xor XOR2 (N1094, N1084, N236);
xor XOR2 (N1095, N1090, N837);
buf BUF1 (N1096, N1089);
buf BUF1 (N1097, N1096);
not NOT1 (N1098, N1093);
nor NOR3 (N1099, N1092, N999, N413);
nor NOR2 (N1100, N1095, N58);
nor NOR4 (N1101, N1091, N562, N96, N980);
and AND2 (N1102, N1100, N411);
nand NAND4 (N1103, N1097, N1072, N542, N276);
buf BUF1 (N1104, N1082);
nand NAND4 (N1105, N1102, N543, N465, N416);
not NOT1 (N1106, N1105);
buf BUF1 (N1107, N1104);
buf BUF1 (N1108, N1098);
not NOT1 (N1109, N1083);
and AND2 (N1110, N1103, N189);
xor XOR2 (N1111, N1110, N149);
or OR4 (N1112, N1106, N637, N689, N764);
xor XOR2 (N1113, N1112, N569);
nand NAND3 (N1114, N1107, N156, N441);
xor XOR2 (N1115, N1111, N172);
or OR2 (N1116, N1081, N585);
not NOT1 (N1117, N1099);
nand NAND2 (N1118, N1109, N579);
nand NAND3 (N1119, N1117, N338, N488);
nor NOR2 (N1120, N1108, N696);
or OR3 (N1121, N1094, N421, N490);
xor XOR2 (N1122, N1101, N16);
or OR3 (N1123, N1119, N370, N463);
buf BUF1 (N1124, N1086);
buf BUF1 (N1125, N1124);
or OR3 (N1126, N1125, N834, N1004);
or OR3 (N1127, N1126, N244, N600);
or OR4 (N1128, N1123, N368, N919, N316);
nor NOR2 (N1129, N1128, N828);
and AND3 (N1130, N1127, N856, N994);
and AND3 (N1131, N1130, N461, N277);
and AND2 (N1132, N1116, N1077);
and AND3 (N1133, N1121, N576, N345);
buf BUF1 (N1134, N1122);
not NOT1 (N1135, N1133);
not NOT1 (N1136, N1115);
and AND2 (N1137, N1120, N956);
xor XOR2 (N1138, N1132, N887);
or OR3 (N1139, N1114, N146, N709);
or OR3 (N1140, N1137, N1075, N365);
nor NOR3 (N1141, N1134, N679, N988);
buf BUF1 (N1142, N1113);
and AND2 (N1143, N1136, N855);
buf BUF1 (N1144, N1143);
not NOT1 (N1145, N1142);
nand NAND3 (N1146, N1140, N831, N651);
xor XOR2 (N1147, N1145, N411);
buf BUF1 (N1148, N1138);
nand NAND4 (N1149, N1148, N410, N427, N1094);
nor NOR2 (N1150, N1149, N442);
not NOT1 (N1151, N1118);
nand NAND2 (N1152, N1129, N822);
and AND2 (N1153, N1147, N354);
nand NAND4 (N1154, N1135, N633, N26, N671);
and AND4 (N1155, N1151, N1056, N384, N849);
and AND3 (N1156, N1155, N311, N544);
and AND4 (N1157, N1144, N571, N958, N486);
nor NOR4 (N1158, N1139, N1013, N423, N790);
not NOT1 (N1159, N1131);
buf BUF1 (N1160, N1146);
xor XOR2 (N1161, N1157, N730);
not NOT1 (N1162, N1141);
nand NAND3 (N1163, N1158, N875, N162);
xor XOR2 (N1164, N1156, N565);
nor NOR2 (N1165, N1153, N697);
nand NAND3 (N1166, N1165, N141, N62);
nand NAND4 (N1167, N1160, N937, N161, N475);
nor NOR2 (N1168, N1163, N134);
and AND3 (N1169, N1162, N901, N299);
xor XOR2 (N1170, N1168, N719);
buf BUF1 (N1171, N1152);
buf BUF1 (N1172, N1169);
nand NAND4 (N1173, N1161, N1169, N873, N286);
xor XOR2 (N1174, N1154, N992);
not NOT1 (N1175, N1166);
or OR3 (N1176, N1175, N988, N676);
xor XOR2 (N1177, N1164, N115);
nand NAND2 (N1178, N1170, N396);
nor NOR3 (N1179, N1172, N678, N358);
buf BUF1 (N1180, N1173);
buf BUF1 (N1181, N1177);
nand NAND2 (N1182, N1176, N556);
nor NOR4 (N1183, N1179, N869, N633, N248);
or OR4 (N1184, N1174, N1060, N1137, N705);
nor NOR3 (N1185, N1167, N624, N865);
xor XOR2 (N1186, N1178, N334);
buf BUF1 (N1187, N1182);
and AND4 (N1188, N1171, N1070, N1069, N1158);
buf BUF1 (N1189, N1159);
xor XOR2 (N1190, N1181, N1168);
buf BUF1 (N1191, N1150);
nand NAND4 (N1192, N1180, N204, N343, N961);
nand NAND3 (N1193, N1185, N43, N1114);
nor NOR3 (N1194, N1191, N231, N804);
or OR3 (N1195, N1192, N1090, N971);
nand NAND4 (N1196, N1193, N320, N902, N319);
and AND4 (N1197, N1183, N97, N1099, N794);
or OR4 (N1198, N1187, N8, N421, N229);
nor NOR4 (N1199, N1198, N895, N420, N1102);
xor XOR2 (N1200, N1196, N76);
not NOT1 (N1201, N1190);
or OR4 (N1202, N1189, N534, N61, N62);
or OR3 (N1203, N1186, N839, N244);
buf BUF1 (N1204, N1194);
xor XOR2 (N1205, N1203, N980);
nor NOR2 (N1206, N1205, N13);
xor XOR2 (N1207, N1201, N944);
buf BUF1 (N1208, N1200);
or OR3 (N1209, N1204, N865, N369);
nand NAND2 (N1210, N1197, N140);
buf BUF1 (N1211, N1188);
or OR3 (N1212, N1211, N1120, N1179);
buf BUF1 (N1213, N1209);
nand NAND3 (N1214, N1184, N454, N353);
and AND3 (N1215, N1213, N181, N688);
or OR3 (N1216, N1208, N647, N767);
not NOT1 (N1217, N1210);
nand NAND2 (N1218, N1195, N843);
xor XOR2 (N1219, N1207, N361);
buf BUF1 (N1220, N1218);
or OR2 (N1221, N1220, N274);
nor NOR2 (N1222, N1212, N888);
and AND3 (N1223, N1219, N151, N325);
nand NAND3 (N1224, N1215, N712, N196);
nor NOR4 (N1225, N1214, N774, N1085, N740);
and AND2 (N1226, N1202, N78);
and AND2 (N1227, N1224, N1008);
buf BUF1 (N1228, N1199);
and AND4 (N1229, N1223, N556, N1003, N896);
nand NAND3 (N1230, N1216, N82, N951);
nor NOR3 (N1231, N1226, N304, N859);
buf BUF1 (N1232, N1206);
nor NOR2 (N1233, N1221, N34);
and AND3 (N1234, N1222, N951, N964);
not NOT1 (N1235, N1229);
buf BUF1 (N1236, N1230);
not NOT1 (N1237, N1236);
buf BUF1 (N1238, N1225);
and AND2 (N1239, N1233, N400);
xor XOR2 (N1240, N1234, N862);
nor NOR4 (N1241, N1228, N298, N821, N367);
nor NOR3 (N1242, N1235, N17, N29);
and AND3 (N1243, N1240, N752, N678);
xor XOR2 (N1244, N1231, N1077);
xor XOR2 (N1245, N1238, N320);
nand NAND4 (N1246, N1232, N186, N821, N505);
or OR3 (N1247, N1246, N392, N1175);
and AND2 (N1248, N1217, N203);
not NOT1 (N1249, N1242);
or OR3 (N1250, N1248, N196, N633);
xor XOR2 (N1251, N1250, N1078);
not NOT1 (N1252, N1227);
not NOT1 (N1253, N1241);
or OR2 (N1254, N1251, N387);
nor NOR3 (N1255, N1243, N1181, N236);
buf BUF1 (N1256, N1249);
nand NAND4 (N1257, N1253, N615, N999, N283);
or OR2 (N1258, N1257, N883);
and AND4 (N1259, N1237, N30, N921, N1090);
or OR4 (N1260, N1247, N1081, N1114, N851);
not NOT1 (N1261, N1239);
nand NAND2 (N1262, N1254, N1058);
buf BUF1 (N1263, N1255);
buf BUF1 (N1264, N1259);
nand NAND2 (N1265, N1245, N462);
xor XOR2 (N1266, N1260, N1118);
or OR2 (N1267, N1256, N904);
nand NAND2 (N1268, N1244, N430);
nand NAND4 (N1269, N1252, N1151, N1130, N613);
or OR3 (N1270, N1268, N1062, N563);
buf BUF1 (N1271, N1258);
nor NOR3 (N1272, N1264, N1188, N900);
or OR3 (N1273, N1263, N804, N1035);
nor NOR3 (N1274, N1272, N1114, N1087);
nand NAND4 (N1275, N1266, N325, N1250, N1165);
nand NAND4 (N1276, N1274, N1089, N140, N601);
and AND2 (N1277, N1276, N404);
xor XOR2 (N1278, N1270, N646);
nand NAND2 (N1279, N1271, N1055);
nor NOR4 (N1280, N1278, N736, N1123, N305);
buf BUF1 (N1281, N1261);
nand NAND3 (N1282, N1275, N710, N627);
and AND2 (N1283, N1281, N944);
nand NAND2 (N1284, N1279, N679);
not NOT1 (N1285, N1269);
nor NOR2 (N1286, N1273, N470);
buf BUF1 (N1287, N1277);
nand NAND3 (N1288, N1284, N1045, N213);
xor XOR2 (N1289, N1288, N833);
buf BUF1 (N1290, N1280);
xor XOR2 (N1291, N1283, N602);
and AND3 (N1292, N1282, N1258, N134);
and AND4 (N1293, N1265, N526, N736, N994);
nand NAND2 (N1294, N1292, N857);
and AND2 (N1295, N1291, N141);
nand NAND2 (N1296, N1294, N899);
or OR3 (N1297, N1262, N996, N183);
and AND3 (N1298, N1285, N446, N924);
and AND3 (N1299, N1286, N339, N751);
nand NAND3 (N1300, N1295, N1132, N158);
not NOT1 (N1301, N1293);
buf BUF1 (N1302, N1290);
and AND4 (N1303, N1299, N205, N580, N1033);
not NOT1 (N1304, N1300);
not NOT1 (N1305, N1297);
buf BUF1 (N1306, N1301);
nand NAND4 (N1307, N1306, N1145, N640, N695);
or OR4 (N1308, N1303, N1058, N336, N1001);
buf BUF1 (N1309, N1287);
nor NOR4 (N1310, N1305, N529, N1303, N597);
not NOT1 (N1311, N1308);
nand NAND4 (N1312, N1311, N285, N408, N1185);
and AND2 (N1313, N1312, N208);
or OR3 (N1314, N1310, N166, N525);
nand NAND4 (N1315, N1267, N629, N1275, N711);
buf BUF1 (N1316, N1309);
nand NAND2 (N1317, N1296, N395);
not NOT1 (N1318, N1289);
xor XOR2 (N1319, N1304, N891);
or OR2 (N1320, N1316, N1144);
nand NAND4 (N1321, N1320, N368, N1095, N326);
and AND2 (N1322, N1298, N528);
not NOT1 (N1323, N1313);
and AND3 (N1324, N1319, N216, N1179);
or OR2 (N1325, N1317, N455);
and AND2 (N1326, N1315, N570);
xor XOR2 (N1327, N1323, N1203);
and AND2 (N1328, N1322, N1099);
and AND2 (N1329, N1314, N1045);
and AND2 (N1330, N1324, N588);
and AND4 (N1331, N1307, N279, N338, N299);
buf BUF1 (N1332, N1331);
xor XOR2 (N1333, N1321, N944);
nor NOR4 (N1334, N1326, N1312, N73, N1000);
and AND4 (N1335, N1334, N1167, N243, N700);
nor NOR4 (N1336, N1329, N244, N883, N114);
nor NOR3 (N1337, N1335, N245, N983);
and AND3 (N1338, N1327, N942, N973);
not NOT1 (N1339, N1325);
xor XOR2 (N1340, N1336, N1279);
nor NOR3 (N1341, N1338, N354, N1216);
xor XOR2 (N1342, N1318, N435);
nand NAND2 (N1343, N1337, N931);
or OR4 (N1344, N1333, N192, N1201, N513);
or OR2 (N1345, N1343, N1046);
not NOT1 (N1346, N1342);
nor NOR2 (N1347, N1345, N7);
and AND4 (N1348, N1340, N209, N862, N20);
buf BUF1 (N1349, N1339);
not NOT1 (N1350, N1302);
or OR2 (N1351, N1341, N121);
and AND2 (N1352, N1330, N670);
xor XOR2 (N1353, N1347, N488);
buf BUF1 (N1354, N1332);
or OR4 (N1355, N1353, N526, N370, N1034);
buf BUF1 (N1356, N1346);
and AND2 (N1357, N1349, N791);
nor NOR2 (N1358, N1350, N336);
buf BUF1 (N1359, N1328);
buf BUF1 (N1360, N1355);
nor NOR2 (N1361, N1352, N551);
nor NOR4 (N1362, N1348, N1232, N961, N1185);
buf BUF1 (N1363, N1351);
and AND4 (N1364, N1357, N1033, N1065, N486);
nand NAND3 (N1365, N1361, N804, N148);
and AND3 (N1366, N1358, N1203, N26);
buf BUF1 (N1367, N1362);
xor XOR2 (N1368, N1364, N1011);
nand NAND3 (N1369, N1368, N522, N1317);
or OR2 (N1370, N1367, N432);
or OR4 (N1371, N1356, N1100, N813, N931);
or OR2 (N1372, N1359, N94);
or OR2 (N1373, N1366, N6);
and AND2 (N1374, N1365, N1283);
buf BUF1 (N1375, N1354);
and AND3 (N1376, N1344, N249, N362);
or OR3 (N1377, N1370, N444, N906);
not NOT1 (N1378, N1376);
nand NAND4 (N1379, N1369, N97, N541, N1110);
buf BUF1 (N1380, N1377);
and AND3 (N1381, N1374, N470, N411);
and AND4 (N1382, N1375, N465, N1134, N904);
xor XOR2 (N1383, N1372, N263);
nor NOR4 (N1384, N1378, N627, N1081, N173);
nand NAND2 (N1385, N1382, N112);
nor NOR3 (N1386, N1381, N371, N102);
buf BUF1 (N1387, N1380);
nor NOR4 (N1388, N1373, N655, N876, N212);
not NOT1 (N1389, N1385);
not NOT1 (N1390, N1360);
xor XOR2 (N1391, N1390, N218);
or OR3 (N1392, N1387, N852, N1141);
not NOT1 (N1393, N1389);
nor NOR2 (N1394, N1379, N1013);
xor XOR2 (N1395, N1393, N899);
and AND3 (N1396, N1392, N934, N831);
xor XOR2 (N1397, N1394, N105);
or OR2 (N1398, N1396, N1257);
xor XOR2 (N1399, N1388, N264);
xor XOR2 (N1400, N1363, N367);
buf BUF1 (N1401, N1400);
xor XOR2 (N1402, N1386, N336);
or OR4 (N1403, N1401, N1367, N1134, N1059);
xor XOR2 (N1404, N1395, N1368);
xor XOR2 (N1405, N1397, N938);
and AND4 (N1406, N1399, N1139, N692, N386);
xor XOR2 (N1407, N1371, N1058);
buf BUF1 (N1408, N1383);
or OR4 (N1409, N1384, N140, N1201, N1012);
nor NOR2 (N1410, N1405, N515);
nand NAND2 (N1411, N1410, N634);
not NOT1 (N1412, N1398);
or OR3 (N1413, N1403, N67, N879);
xor XOR2 (N1414, N1402, N332);
nand NAND4 (N1415, N1408, N1235, N266, N472);
buf BUF1 (N1416, N1391);
buf BUF1 (N1417, N1411);
xor XOR2 (N1418, N1412, N213);
or OR4 (N1419, N1407, N1119, N187, N528);
not NOT1 (N1420, N1414);
and AND2 (N1421, N1415, N350);
nand NAND4 (N1422, N1417, N306, N922, N353);
not NOT1 (N1423, N1419);
and AND4 (N1424, N1416, N1395, N224, N1030);
nor NOR3 (N1425, N1409, N826, N1123);
nand NAND2 (N1426, N1406, N1418);
not NOT1 (N1427, N1304);
and AND3 (N1428, N1424, N1364, N48);
buf BUF1 (N1429, N1413);
buf BUF1 (N1430, N1425);
or OR3 (N1431, N1429, N1225, N1229);
nor NOR3 (N1432, N1426, N721, N190);
nor NOR2 (N1433, N1404, N885);
or OR2 (N1434, N1427, N358);
or OR2 (N1435, N1428, N436);
nor NOR4 (N1436, N1420, N81, N301, N1117);
nor NOR2 (N1437, N1435, N1004);
and AND3 (N1438, N1433, N844, N425);
buf BUF1 (N1439, N1430);
and AND4 (N1440, N1423, N229, N47, N860);
not NOT1 (N1441, N1422);
and AND3 (N1442, N1437, N733, N1001);
not NOT1 (N1443, N1441);
buf BUF1 (N1444, N1434);
nor NOR2 (N1445, N1440, N407);
or OR3 (N1446, N1439, N1043, N1168);
and AND4 (N1447, N1432, N1006, N1244, N540);
xor XOR2 (N1448, N1438, N326);
xor XOR2 (N1449, N1431, N210);
nor NOR3 (N1450, N1447, N597, N1011);
buf BUF1 (N1451, N1443);
buf BUF1 (N1452, N1421);
and AND4 (N1453, N1448, N187, N90, N809);
buf BUF1 (N1454, N1442);
nand NAND4 (N1455, N1444, N515, N673, N648);
buf BUF1 (N1456, N1454);
nand NAND2 (N1457, N1456, N1046);
nand NAND2 (N1458, N1451, N963);
not NOT1 (N1459, N1449);
or OR4 (N1460, N1452, N153, N694, N223);
or OR4 (N1461, N1446, N1323, N1, N71);
nor NOR3 (N1462, N1450, N169, N731);
buf BUF1 (N1463, N1462);
nor NOR3 (N1464, N1455, N161, N966);
buf BUF1 (N1465, N1460);
and AND2 (N1466, N1436, N389);
and AND3 (N1467, N1463, N973, N608);
xor XOR2 (N1468, N1459, N1116);
or OR4 (N1469, N1466, N1321, N405, N234);
or OR3 (N1470, N1458, N850, N471);
not NOT1 (N1471, N1445);
and AND4 (N1472, N1453, N849, N1080, N701);
nand NAND3 (N1473, N1468, N485, N236);
or OR2 (N1474, N1469, N100);
not NOT1 (N1475, N1461);
and AND2 (N1476, N1467, N912);
not NOT1 (N1477, N1473);
nor NOR3 (N1478, N1474, N988, N385);
nand NAND2 (N1479, N1471, N1146);
buf BUF1 (N1480, N1470);
xor XOR2 (N1481, N1480, N1396);
nor NOR2 (N1482, N1472, N1096);
and AND4 (N1483, N1478, N399, N840, N192);
xor XOR2 (N1484, N1479, N616);
not NOT1 (N1485, N1484);
or OR4 (N1486, N1483, N732, N359, N618);
buf BUF1 (N1487, N1464);
or OR3 (N1488, N1457, N1291, N17);
xor XOR2 (N1489, N1488, N18);
xor XOR2 (N1490, N1481, N614);
buf BUF1 (N1491, N1486);
nand NAND3 (N1492, N1477, N728, N497);
nand NAND4 (N1493, N1482, N1016, N575, N119);
or OR2 (N1494, N1465, N1148);
or OR4 (N1495, N1494, N1247, N1206, N807);
and AND4 (N1496, N1492, N1441, N391, N1120);
nor NOR2 (N1497, N1493, N1315);
nand NAND4 (N1498, N1497, N492, N52, N996);
nor NOR2 (N1499, N1476, N123);
not NOT1 (N1500, N1487);
or OR3 (N1501, N1499, N1321, N1431);
nand NAND4 (N1502, N1489, N45, N1019, N441);
nand NAND3 (N1503, N1475, N1160, N31);
and AND3 (N1504, N1485, N495, N745);
and AND3 (N1505, N1500, N1222, N435);
or OR4 (N1506, N1502, N583, N971, N1419);
or OR2 (N1507, N1498, N414);
nor NOR4 (N1508, N1491, N366, N1034, N164);
nor NOR2 (N1509, N1506, N85);
not NOT1 (N1510, N1504);
nand NAND4 (N1511, N1496, N62, N1137, N1481);
and AND4 (N1512, N1505, N211, N285, N436);
xor XOR2 (N1513, N1510, N1097);
nor NOR4 (N1514, N1501, N193, N912, N386);
xor XOR2 (N1515, N1507, N552);
nor NOR2 (N1516, N1512, N1174);
nand NAND4 (N1517, N1508, N467, N1345, N354);
or OR2 (N1518, N1517, N494);
xor XOR2 (N1519, N1515, N271);
buf BUF1 (N1520, N1513);
xor XOR2 (N1521, N1518, N1344);
buf BUF1 (N1522, N1511);
and AND3 (N1523, N1495, N1391, N1496);
buf BUF1 (N1524, N1523);
or OR4 (N1525, N1524, N765, N24, N388);
and AND3 (N1526, N1525, N1429, N746);
nor NOR2 (N1527, N1514, N384);
nor NOR2 (N1528, N1527, N885);
xor XOR2 (N1529, N1509, N1207);
not NOT1 (N1530, N1521);
not NOT1 (N1531, N1490);
xor XOR2 (N1532, N1526, N72);
xor XOR2 (N1533, N1532, N105);
nor NOR4 (N1534, N1530, N174, N297, N221);
xor XOR2 (N1535, N1529, N662);
nand NAND3 (N1536, N1533, N1170, N232);
nand NAND3 (N1537, N1535, N554, N302);
xor XOR2 (N1538, N1536, N813);
not NOT1 (N1539, N1503);
nor NOR2 (N1540, N1531, N868);
nor NOR4 (N1541, N1539, N396, N348, N1102);
and AND4 (N1542, N1519, N1034, N806, N59);
xor XOR2 (N1543, N1522, N808);
nand NAND3 (N1544, N1540, N215, N376);
nor NOR2 (N1545, N1528, N508);
nand NAND2 (N1546, N1538, N1351);
or OR4 (N1547, N1520, N1311, N1525, N135);
nand NAND3 (N1548, N1545, N1020, N1501);
and AND2 (N1549, N1544, N1516);
not NOT1 (N1550, N539);
and AND2 (N1551, N1550, N1258);
and AND4 (N1552, N1534, N1196, N845, N777);
and AND4 (N1553, N1543, N1033, N988, N1551);
not NOT1 (N1554, N703);
buf BUF1 (N1555, N1541);
not NOT1 (N1556, N1553);
not NOT1 (N1557, N1555);
not NOT1 (N1558, N1542);
buf BUF1 (N1559, N1554);
and AND3 (N1560, N1548, N489, N1057);
nor NOR3 (N1561, N1558, N1470, N900);
nand NAND2 (N1562, N1559, N1344);
xor XOR2 (N1563, N1561, N722);
not NOT1 (N1564, N1556);
not NOT1 (N1565, N1564);
or OR2 (N1566, N1563, N1357);
or OR2 (N1567, N1547, N803);
buf BUF1 (N1568, N1560);
and AND3 (N1569, N1567, N534, N301);
nand NAND4 (N1570, N1537, N1200, N36, N1132);
xor XOR2 (N1571, N1565, N113);
nor NOR3 (N1572, N1549, N1531, N1512);
buf BUF1 (N1573, N1572);
nor NOR4 (N1574, N1562, N967, N482, N784);
or OR4 (N1575, N1573, N1153, N873, N149);
or OR2 (N1576, N1568, N97);
not NOT1 (N1577, N1574);
xor XOR2 (N1578, N1570, N1270);
buf BUF1 (N1579, N1571);
buf BUF1 (N1580, N1576);
not NOT1 (N1581, N1578);
xor XOR2 (N1582, N1566, N427);
not NOT1 (N1583, N1581);
xor XOR2 (N1584, N1575, N293);
not NOT1 (N1585, N1569);
nand NAND2 (N1586, N1583, N1465);
xor XOR2 (N1587, N1585, N55);
and AND4 (N1588, N1582, N874, N765, N641);
xor XOR2 (N1589, N1546, N1041);
nor NOR4 (N1590, N1580, N1460, N920, N1519);
buf BUF1 (N1591, N1584);
xor XOR2 (N1592, N1587, N1148);
nor NOR2 (N1593, N1557, N751);
or OR3 (N1594, N1591, N286, N889);
buf BUF1 (N1595, N1579);
not NOT1 (N1596, N1590);
not NOT1 (N1597, N1589);
nand NAND2 (N1598, N1596, N638);
not NOT1 (N1599, N1597);
or OR4 (N1600, N1594, N508, N1322, N312);
or OR2 (N1601, N1592, N1161);
or OR2 (N1602, N1552, N383);
nor NOR3 (N1603, N1599, N937, N983);
nand NAND3 (N1604, N1598, N1102, N963);
nand NAND3 (N1605, N1595, N1019, N40);
xor XOR2 (N1606, N1604, N345);
or OR2 (N1607, N1603, N296);
xor XOR2 (N1608, N1601, N612);
or OR4 (N1609, N1608, N834, N863, N932);
or OR4 (N1610, N1602, N284, N13, N323);
nor NOR2 (N1611, N1607, N3);
and AND2 (N1612, N1611, N1195);
or OR2 (N1613, N1588, N1084);
xor XOR2 (N1614, N1613, N1299);
xor XOR2 (N1615, N1606, N1332);
buf BUF1 (N1616, N1610);
buf BUF1 (N1617, N1614);
not NOT1 (N1618, N1577);
and AND2 (N1619, N1616, N1578);
nand NAND3 (N1620, N1615, N1397, N1263);
or OR3 (N1621, N1612, N988, N1369);
nand NAND2 (N1622, N1609, N921);
or OR4 (N1623, N1600, N1039, N272, N676);
buf BUF1 (N1624, N1620);
nor NOR4 (N1625, N1605, N607, N232, N726);
or OR3 (N1626, N1625, N1284, N305);
and AND3 (N1627, N1624, N1392, N1074);
nor NOR4 (N1628, N1617, N724, N1494, N919);
nor NOR4 (N1629, N1622, N742, N12, N1146);
and AND2 (N1630, N1627, N1560);
not NOT1 (N1631, N1626);
and AND4 (N1632, N1628, N616, N6, N1108);
xor XOR2 (N1633, N1630, N791);
nor NOR4 (N1634, N1629, N596, N1251, N565);
nor NOR2 (N1635, N1623, N568);
nand NAND2 (N1636, N1586, N634);
or OR3 (N1637, N1593, N793, N885);
nor NOR2 (N1638, N1632, N203);
xor XOR2 (N1639, N1618, N486);
not NOT1 (N1640, N1636);
xor XOR2 (N1641, N1633, N269);
and AND3 (N1642, N1619, N375, N1610);
xor XOR2 (N1643, N1642, N748);
not NOT1 (N1644, N1634);
xor XOR2 (N1645, N1644, N49);
nor NOR3 (N1646, N1640, N1188, N573);
and AND4 (N1647, N1631, N1526, N1227, N1375);
not NOT1 (N1648, N1647);
nand NAND3 (N1649, N1621, N486, N1425);
nand NAND4 (N1650, N1645, N1382, N24, N1044);
xor XOR2 (N1651, N1637, N512);
not NOT1 (N1652, N1638);
nand NAND3 (N1653, N1635, N628, N190);
nand NAND4 (N1654, N1648, N1061, N461, N376);
xor XOR2 (N1655, N1639, N1057);
and AND4 (N1656, N1646, N594, N1654, N1103);
nand NAND4 (N1657, N992, N593, N1370, N211);
buf BUF1 (N1658, N1643);
buf BUF1 (N1659, N1641);
xor XOR2 (N1660, N1659, N532);
and AND4 (N1661, N1655, N1080, N702, N31);
nor NOR3 (N1662, N1652, N987, N127);
nor NOR2 (N1663, N1649, N113);
xor XOR2 (N1664, N1651, N1293);
nand NAND2 (N1665, N1663, N975);
or OR4 (N1666, N1653, N1512, N1518, N252);
buf BUF1 (N1667, N1661);
buf BUF1 (N1668, N1658);
nand NAND2 (N1669, N1660, N1648);
and AND4 (N1670, N1669, N1499, N1473, N482);
xor XOR2 (N1671, N1662, N529);
buf BUF1 (N1672, N1665);
or OR4 (N1673, N1664, N880, N430, N1387);
nand NAND4 (N1674, N1666, N1267, N1282, N965);
nor NOR4 (N1675, N1674, N169, N805, N589);
nand NAND2 (N1676, N1671, N63);
nand NAND4 (N1677, N1675, N1163, N155, N740);
xor XOR2 (N1678, N1670, N729);
buf BUF1 (N1679, N1676);
nand NAND2 (N1680, N1656, N991);
buf BUF1 (N1681, N1673);
and AND2 (N1682, N1672, N738);
nand NAND2 (N1683, N1681, N1306);
and AND4 (N1684, N1679, N449, N1580, N378);
nand NAND2 (N1685, N1650, N924);
nor NOR2 (N1686, N1668, N1146);
or OR3 (N1687, N1667, N908, N1420);
or OR2 (N1688, N1682, N31);
not NOT1 (N1689, N1686);
nand NAND2 (N1690, N1685, N1532);
xor XOR2 (N1691, N1689, N1349);
xor XOR2 (N1692, N1677, N46);
nand NAND3 (N1693, N1684, N653, N323);
buf BUF1 (N1694, N1691);
xor XOR2 (N1695, N1692, N674);
buf BUF1 (N1696, N1680);
buf BUF1 (N1697, N1696);
or OR4 (N1698, N1695, N1371, N110, N1641);
and AND3 (N1699, N1697, N1497, N14);
not NOT1 (N1700, N1688);
buf BUF1 (N1701, N1694);
nor NOR2 (N1702, N1700, N1055);
or OR4 (N1703, N1678, N921, N1308, N1520);
nand NAND2 (N1704, N1703, N373);
buf BUF1 (N1705, N1702);
nor NOR3 (N1706, N1687, N1339, N427);
nand NAND4 (N1707, N1693, N740, N1038, N1059);
or OR4 (N1708, N1707, N1673, N263, N741);
xor XOR2 (N1709, N1706, N1259);
not NOT1 (N1710, N1708);
nand NAND4 (N1711, N1710, N1396, N1128, N340);
xor XOR2 (N1712, N1657, N1272);
and AND4 (N1713, N1698, N39, N1071, N139);
and AND3 (N1714, N1701, N1095, N636);
buf BUF1 (N1715, N1712);
and AND4 (N1716, N1705, N313, N389, N1169);
and AND2 (N1717, N1713, N1666);
and AND2 (N1718, N1714, N1516);
not NOT1 (N1719, N1699);
not NOT1 (N1720, N1716);
and AND4 (N1721, N1709, N8, N695, N1072);
xor XOR2 (N1722, N1718, N1225);
and AND3 (N1723, N1717, N1252, N1100);
nand NAND4 (N1724, N1711, N598, N161, N1380);
and AND2 (N1725, N1704, N187);
or OR2 (N1726, N1723, N1170);
xor XOR2 (N1727, N1722, N233);
nor NOR3 (N1728, N1720, N1205, N949);
nand NAND3 (N1729, N1724, N148, N1058);
or OR4 (N1730, N1725, N912, N1129, N113);
not NOT1 (N1731, N1728);
xor XOR2 (N1732, N1729, N398);
nor NOR3 (N1733, N1727, N1695, N397);
xor XOR2 (N1734, N1715, N1451);
nand NAND3 (N1735, N1732, N1513, N281);
and AND3 (N1736, N1734, N1245, N1268);
and AND3 (N1737, N1719, N373, N486);
nand NAND3 (N1738, N1726, N1713, N1599);
nor NOR4 (N1739, N1690, N1392, N113, N1390);
nor NOR2 (N1740, N1730, N488);
xor XOR2 (N1741, N1731, N170);
nand NAND3 (N1742, N1740, N1231, N1190);
xor XOR2 (N1743, N1735, N1430);
xor XOR2 (N1744, N1742, N1664);
nor NOR4 (N1745, N1733, N396, N1585, N1436);
xor XOR2 (N1746, N1745, N144);
nor NOR4 (N1747, N1738, N162, N1735, N321);
nand NAND4 (N1748, N1746, N588, N408, N374);
not NOT1 (N1749, N1739);
or OR2 (N1750, N1721, N66);
and AND2 (N1751, N1743, N1632);
not NOT1 (N1752, N1750);
nand NAND4 (N1753, N1749, N266, N1231, N1170);
xor XOR2 (N1754, N1683, N258);
nand NAND2 (N1755, N1748, N293);
and AND2 (N1756, N1744, N175);
or OR2 (N1757, N1756, N1589);
nand NAND2 (N1758, N1737, N1476);
not NOT1 (N1759, N1754);
not NOT1 (N1760, N1752);
xor XOR2 (N1761, N1760, N955);
and AND4 (N1762, N1747, N1708, N72, N483);
nor NOR2 (N1763, N1755, N1294);
not NOT1 (N1764, N1758);
xor XOR2 (N1765, N1762, N934);
and AND4 (N1766, N1753, N1409, N677, N1251);
or OR4 (N1767, N1766, N1551, N1523, N546);
nor NOR4 (N1768, N1761, N1316, N1336, N1361);
or OR4 (N1769, N1757, N1183, N1762, N363);
buf BUF1 (N1770, N1741);
nor NOR3 (N1771, N1736, N727, N1097);
and AND3 (N1772, N1770, N251, N777);
xor XOR2 (N1773, N1759, N277);
not NOT1 (N1774, N1773);
buf BUF1 (N1775, N1767);
not NOT1 (N1776, N1768);
and AND2 (N1777, N1751, N285);
xor XOR2 (N1778, N1771, N875);
buf BUF1 (N1779, N1776);
and AND4 (N1780, N1764, N812, N1547, N626);
xor XOR2 (N1781, N1779, N623);
buf BUF1 (N1782, N1774);
or OR4 (N1783, N1763, N1181, N770, N402);
xor XOR2 (N1784, N1769, N1494);
xor XOR2 (N1785, N1784, N1470);
and AND3 (N1786, N1765, N721, N643);
not NOT1 (N1787, N1786);
and AND2 (N1788, N1780, N633);
buf BUF1 (N1789, N1788);
buf BUF1 (N1790, N1782);
nand NAND3 (N1791, N1777, N1042, N75);
nand NAND3 (N1792, N1778, N743, N893);
nand NAND4 (N1793, N1775, N8, N671, N351);
not NOT1 (N1794, N1791);
and AND2 (N1795, N1772, N1352);
xor XOR2 (N1796, N1781, N998);
not NOT1 (N1797, N1783);
buf BUF1 (N1798, N1792);
and AND4 (N1799, N1794, N893, N553, N988);
nand NAND4 (N1800, N1789, N890, N1031, N1672);
not NOT1 (N1801, N1785);
buf BUF1 (N1802, N1787);
and AND3 (N1803, N1798, N55, N1679);
and AND3 (N1804, N1802, N407, N828);
nor NOR3 (N1805, N1800, N148, N1621);
and AND4 (N1806, N1793, N778, N1237, N869);
nand NAND3 (N1807, N1799, N27, N310);
and AND4 (N1808, N1806, N1195, N442, N180);
or OR2 (N1809, N1795, N1734);
and AND4 (N1810, N1809, N1807, N837, N514);
and AND3 (N1811, N1514, N804, N1202);
or OR4 (N1812, N1790, N1009, N374, N28);
xor XOR2 (N1813, N1796, N1504);
or OR4 (N1814, N1804, N163, N548, N1387);
and AND3 (N1815, N1805, N340, N555);
not NOT1 (N1816, N1814);
or OR3 (N1817, N1803, N385, N1074);
and AND3 (N1818, N1801, N352, N1332);
or OR4 (N1819, N1810, N939, N1305, N1545);
nand NAND2 (N1820, N1816, N1716);
nand NAND4 (N1821, N1815, N1350, N159, N1121);
buf BUF1 (N1822, N1812);
and AND3 (N1823, N1818, N604, N473);
nor NOR3 (N1824, N1817, N1511, N1797);
and AND2 (N1825, N1231, N1424);
and AND2 (N1826, N1819, N1305);
and AND4 (N1827, N1826, N1049, N1344, N133);
not NOT1 (N1828, N1820);
or OR3 (N1829, N1821, N1741, N87);
or OR2 (N1830, N1822, N328);
buf BUF1 (N1831, N1823);
and AND2 (N1832, N1827, N1034);
nor NOR3 (N1833, N1811, N691, N280);
or OR3 (N1834, N1824, N1237, N558);
or OR2 (N1835, N1833, N914);
nand NAND3 (N1836, N1828, N1805, N286);
not NOT1 (N1837, N1834);
and AND3 (N1838, N1808, N446, N844);
and AND2 (N1839, N1835, N1241);
xor XOR2 (N1840, N1839, N172);
xor XOR2 (N1841, N1831, N1820);
and AND4 (N1842, N1840, N1298, N80, N977);
not NOT1 (N1843, N1832);
not NOT1 (N1844, N1843);
xor XOR2 (N1845, N1830, N707);
xor XOR2 (N1846, N1837, N1030);
or OR4 (N1847, N1844, N921, N299, N818);
not NOT1 (N1848, N1841);
and AND3 (N1849, N1845, N1021, N62);
and AND3 (N1850, N1829, N1268, N1276);
buf BUF1 (N1851, N1813);
and AND2 (N1852, N1838, N223);
buf BUF1 (N1853, N1846);
nor NOR3 (N1854, N1852, N580, N1477);
nand NAND4 (N1855, N1853, N1383, N70, N1241);
xor XOR2 (N1856, N1855, N882);
or OR2 (N1857, N1825, N1785);
nand NAND3 (N1858, N1854, N447, N393);
not NOT1 (N1859, N1848);
buf BUF1 (N1860, N1859);
nand NAND4 (N1861, N1851, N1161, N1661, N41);
buf BUF1 (N1862, N1842);
xor XOR2 (N1863, N1847, N579);
xor XOR2 (N1864, N1850, N804);
buf BUF1 (N1865, N1858);
not NOT1 (N1866, N1864);
nand NAND4 (N1867, N1836, N994, N1254, N1467);
or OR4 (N1868, N1866, N1121, N891, N175);
and AND4 (N1869, N1860, N349, N1791, N770);
xor XOR2 (N1870, N1868, N1226);
or OR2 (N1871, N1870, N682);
nand NAND2 (N1872, N1871, N769);
xor XOR2 (N1873, N1856, N8);
and AND2 (N1874, N1865, N1384);
and AND2 (N1875, N1874, N197);
nor NOR3 (N1876, N1862, N606, N734);
or OR4 (N1877, N1873, N1356, N813, N1488);
and AND2 (N1878, N1877, N1304);
or OR2 (N1879, N1861, N102);
or OR4 (N1880, N1867, N563, N1615, N1432);
buf BUF1 (N1881, N1857);
nor NOR3 (N1882, N1863, N1045, N1260);
xor XOR2 (N1883, N1872, N316);
buf BUF1 (N1884, N1878);
or OR4 (N1885, N1881, N50, N294, N5);
not NOT1 (N1886, N1876);
nor NOR4 (N1887, N1885, N1485, N943, N945);
buf BUF1 (N1888, N1880);
xor XOR2 (N1889, N1884, N1675);
not NOT1 (N1890, N1879);
nand NAND2 (N1891, N1887, N84);
buf BUF1 (N1892, N1875);
nor NOR2 (N1893, N1889, N1086);
buf BUF1 (N1894, N1869);
or OR4 (N1895, N1888, N1186, N1703, N663);
xor XOR2 (N1896, N1894, N908);
xor XOR2 (N1897, N1893, N1771);
and AND4 (N1898, N1890, N197, N1746, N1895);
buf BUF1 (N1899, N1787);
buf BUF1 (N1900, N1891);
or OR4 (N1901, N1892, N206, N992, N310);
buf BUF1 (N1902, N1900);
nor NOR4 (N1903, N1882, N1275, N449, N169);
buf BUF1 (N1904, N1899);
buf BUF1 (N1905, N1897);
nor NOR2 (N1906, N1849, N1776);
or OR3 (N1907, N1886, N1266, N1455);
xor XOR2 (N1908, N1898, N1324);
nand NAND3 (N1909, N1906, N1120, N900);
nor NOR4 (N1910, N1907, N1357, N174, N1109);
nand NAND3 (N1911, N1902, N482, N1664);
not NOT1 (N1912, N1910);
and AND2 (N1913, N1901, N1498);
not NOT1 (N1914, N1903);
xor XOR2 (N1915, N1909, N696);
not NOT1 (N1916, N1896);
nor NOR3 (N1917, N1915, N1015, N1575);
buf BUF1 (N1918, N1883);
nor NOR4 (N1919, N1918, N283, N570, N1143);
or OR4 (N1920, N1919, N964, N1499, N1265);
xor XOR2 (N1921, N1914, N1270);
not NOT1 (N1922, N1911);
and AND4 (N1923, N1917, N1077, N1144, N328);
buf BUF1 (N1924, N1923);
buf BUF1 (N1925, N1916);
nand NAND4 (N1926, N1913, N1773, N1689, N1480);
and AND2 (N1927, N1926, N915);
not NOT1 (N1928, N1924);
not NOT1 (N1929, N1927);
and AND2 (N1930, N1921, N876);
and AND2 (N1931, N1905, N95);
buf BUF1 (N1932, N1920);
not NOT1 (N1933, N1928);
nor NOR2 (N1934, N1912, N461);
or OR3 (N1935, N1922, N1602, N1354);
xor XOR2 (N1936, N1935, N981);
nor NOR4 (N1937, N1929, N747, N1316, N1554);
xor XOR2 (N1938, N1936, N1718);
not NOT1 (N1939, N1932);
nand NAND4 (N1940, N1934, N29, N270, N922);
or OR2 (N1941, N1933, N411);
not NOT1 (N1942, N1931);
not NOT1 (N1943, N1930);
buf BUF1 (N1944, N1941);
not NOT1 (N1945, N1904);
buf BUF1 (N1946, N1938);
not NOT1 (N1947, N1946);
nand NAND4 (N1948, N1945, N1153, N1066, N1683);
or OR4 (N1949, N1937, N294, N64, N1117);
xor XOR2 (N1950, N1939, N820);
not NOT1 (N1951, N1949);
and AND4 (N1952, N1943, N1909, N822, N1287);
xor XOR2 (N1953, N1947, N245);
and AND2 (N1954, N1940, N409);
and AND4 (N1955, N1908, N1455, N455, N1275);
xor XOR2 (N1956, N1948, N964);
and AND4 (N1957, N1950, N1784, N1290, N821);
buf BUF1 (N1958, N1956);
not NOT1 (N1959, N1944);
xor XOR2 (N1960, N1925, N1036);
nand NAND4 (N1961, N1942, N1095, N1910, N974);
not NOT1 (N1962, N1952);
nand NAND3 (N1963, N1959, N1591, N606);
xor XOR2 (N1964, N1955, N1303);
or OR4 (N1965, N1960, N1825, N694, N1277);
nand NAND3 (N1966, N1963, N1545, N1469);
and AND4 (N1967, N1951, N1429, N405, N1356);
nand NAND3 (N1968, N1961, N402, N1343);
or OR4 (N1969, N1953, N1232, N656, N683);
and AND2 (N1970, N1957, N1483);
not NOT1 (N1971, N1958);
buf BUF1 (N1972, N1971);
nor NOR2 (N1973, N1965, N419);
nand NAND3 (N1974, N1970, N1932, N905);
nor NOR4 (N1975, N1974, N708, N1493, N447);
nand NAND2 (N1976, N1968, N411);
not NOT1 (N1977, N1976);
not NOT1 (N1978, N1975);
nor NOR4 (N1979, N1954, N46, N1700, N1397);
xor XOR2 (N1980, N1966, N900);
buf BUF1 (N1981, N1969);
and AND4 (N1982, N1977, N1477, N821, N1917);
not NOT1 (N1983, N1979);
and AND4 (N1984, N1983, N1595, N656, N745);
not NOT1 (N1985, N1980);
buf BUF1 (N1986, N1973);
xor XOR2 (N1987, N1985, N787);
xor XOR2 (N1988, N1981, N50);
or OR2 (N1989, N1962, N304);
and AND2 (N1990, N1984, N84);
buf BUF1 (N1991, N1964);
not NOT1 (N1992, N1991);
or OR2 (N1993, N1972, N48);
nand NAND2 (N1994, N1990, N206);
xor XOR2 (N1995, N1988, N1475);
nand NAND2 (N1996, N1989, N1125);
and AND4 (N1997, N1986, N1721, N1109, N1216);
nand NAND3 (N1998, N1982, N365, N1950);
or OR2 (N1999, N1993, N1906);
nor NOR2 (N2000, N1978, N214);
nor NOR4 (N2001, N1996, N777, N998, N23);
or OR2 (N2002, N1997, N49);
xor XOR2 (N2003, N2000, N143);
and AND4 (N2004, N1992, N1456, N921, N1422);
xor XOR2 (N2005, N2002, N570);
or OR2 (N2006, N1998, N156);
and AND3 (N2007, N1994, N1175, N1057);
buf BUF1 (N2008, N2006);
and AND3 (N2009, N1995, N695, N814);
nand NAND2 (N2010, N2003, N65);
nand NAND2 (N2011, N2007, N1684);
nand NAND4 (N2012, N2010, N685, N1798, N475);
not NOT1 (N2013, N2008);
xor XOR2 (N2014, N1987, N784);
not NOT1 (N2015, N2013);
nor NOR4 (N2016, N2015, N1455, N1222, N332);
nor NOR2 (N2017, N1967, N1689);
nand NAND4 (N2018, N2014, N407, N1731, N1748);
not NOT1 (N2019, N2004);
or OR2 (N2020, N2019, N1786);
nand NAND2 (N2021, N2017, N1466);
xor XOR2 (N2022, N2012, N684);
and AND4 (N2023, N2001, N483, N326, N959);
and AND4 (N2024, N1999, N71, N7, N1532);
endmodule