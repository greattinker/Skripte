// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N3994,N4008,N4002,N4001,N3987,N4012,N4006,N4011,N4005,N4013;

or OR4 (N14, N12, N1, N11, N6);
or OR2 (N15, N12, N8);
nand NAND3 (N16, N4, N14, N6);
or OR2 (N17, N12, N13);
nand NAND2 (N18, N1, N1);
nand NAND3 (N19, N10, N14, N18);
nand NAND3 (N20, N6, N4, N3);
and AND3 (N21, N16, N5, N12);
nand NAND4 (N22, N18, N2, N10, N8);
and AND2 (N23, N9, N10);
buf BUF1 (N24, N17);
xor XOR2 (N25, N17, N1);
nor NOR2 (N26, N4, N5);
and AND4 (N27, N17, N24, N19, N13);
or OR4 (N28, N20, N11, N9, N18);
nand NAND4 (N29, N1, N23, N18, N25);
or OR2 (N30, N8, N14);
xor XOR2 (N31, N4, N17);
nand NAND4 (N32, N21, N23, N20, N10);
not NOT1 (N33, N13);
not NOT1 (N34, N15);
or OR3 (N35, N30, N11, N9);
xor XOR2 (N36, N31, N18);
and AND4 (N37, N34, N14, N14, N12);
xor XOR2 (N38, N36, N17);
buf BUF1 (N39, N26);
xor XOR2 (N40, N33, N33);
not NOT1 (N41, N29);
xor XOR2 (N42, N22, N34);
not NOT1 (N43, N42);
not NOT1 (N44, N37);
buf BUF1 (N45, N43);
and AND3 (N46, N35, N5, N33);
not NOT1 (N47, N40);
buf BUF1 (N48, N27);
not NOT1 (N49, N32);
buf BUF1 (N50, N28);
not NOT1 (N51, N41);
and AND3 (N52, N51, N22, N49);
buf BUF1 (N53, N19);
nand NAND2 (N54, N52, N45);
nand NAND4 (N55, N52, N48, N3, N12);
nor NOR4 (N56, N7, N27, N24, N19);
not NOT1 (N57, N53);
xor XOR2 (N58, N56, N9);
not NOT1 (N59, N58);
nor NOR2 (N60, N57, N21);
and AND4 (N61, N39, N19, N29, N25);
or OR2 (N62, N60, N44);
or OR2 (N63, N19, N49);
xor XOR2 (N64, N47, N60);
buf BUF1 (N65, N59);
xor XOR2 (N66, N50, N27);
nor NOR2 (N67, N63, N43);
or OR2 (N68, N66, N13);
buf BUF1 (N69, N61);
and AND2 (N70, N62, N40);
or OR4 (N71, N38, N59, N9, N61);
nand NAND4 (N72, N65, N25, N19, N71);
xor XOR2 (N73, N57, N64);
xor XOR2 (N74, N39, N37);
and AND2 (N75, N46, N42);
not NOT1 (N76, N67);
nand NAND2 (N77, N70, N6);
not NOT1 (N78, N69);
nor NOR2 (N79, N76, N15);
or OR3 (N80, N68, N61, N59);
or OR4 (N81, N80, N30, N26, N13);
and AND3 (N82, N79, N2, N2);
xor XOR2 (N83, N55, N66);
and AND4 (N84, N72, N2, N9, N46);
xor XOR2 (N85, N54, N68);
or OR2 (N86, N82, N14);
buf BUF1 (N87, N86);
nand NAND3 (N88, N74, N47, N3);
buf BUF1 (N89, N83);
xor XOR2 (N90, N75, N22);
and AND3 (N91, N73, N71, N28);
nand NAND3 (N92, N84, N25, N57);
or OR4 (N93, N87, N7, N37, N43);
nor NOR2 (N94, N81, N5);
and AND2 (N95, N90, N72);
buf BUF1 (N96, N85);
nand NAND4 (N97, N88, N21, N21, N81);
and AND4 (N98, N94, N69, N95, N73);
and AND4 (N99, N5, N22, N83, N40);
nor NOR4 (N100, N91, N76, N24, N95);
and AND4 (N101, N96, N21, N17, N80);
or OR2 (N102, N77, N87);
or OR2 (N103, N99, N97);
not NOT1 (N104, N74);
nor NOR3 (N105, N103, N36, N67);
buf BUF1 (N106, N89);
not NOT1 (N107, N101);
nand NAND4 (N108, N98, N20, N10, N64);
not NOT1 (N109, N93);
not NOT1 (N110, N107);
nand NAND3 (N111, N78, N41, N100);
xor XOR2 (N112, N43, N87);
not NOT1 (N113, N111);
nand NAND3 (N114, N102, N2, N110);
nor NOR4 (N115, N83, N98, N98, N94);
nor NOR3 (N116, N109, N21, N60);
or OR4 (N117, N116, N66, N8, N36);
nor NOR2 (N118, N92, N55);
xor XOR2 (N119, N104, N79);
buf BUF1 (N120, N118);
nand NAND3 (N121, N105, N29, N66);
nor NOR4 (N122, N117, N106, N38, N37);
buf BUF1 (N123, N15);
nand NAND4 (N124, N122, N100, N87, N86);
or OR2 (N125, N124, N15);
or OR4 (N126, N120, N86, N80, N106);
or OR3 (N127, N108, N126, N53);
nor NOR4 (N128, N36, N107, N28, N119);
xor XOR2 (N129, N12, N123);
not NOT1 (N130, N62);
nand NAND3 (N131, N127, N74, N14);
not NOT1 (N132, N112);
nor NOR3 (N133, N114, N47, N99);
nor NOR3 (N134, N133, N11, N97);
not NOT1 (N135, N125);
or OR3 (N136, N115, N84, N102);
or OR4 (N137, N129, N30, N97, N96);
nor NOR2 (N138, N130, N108);
nand NAND3 (N139, N121, N65, N52);
buf BUF1 (N140, N132);
xor XOR2 (N141, N137, N99);
nor NOR3 (N142, N141, N108, N120);
nand NAND4 (N143, N142, N82, N2, N102);
buf BUF1 (N144, N143);
nor NOR3 (N145, N131, N142, N25);
or OR3 (N146, N128, N112, N34);
or OR2 (N147, N144, N65);
not NOT1 (N148, N140);
nand NAND3 (N149, N145, N32, N31);
nand NAND2 (N150, N135, N142);
or OR4 (N151, N113, N20, N24, N44);
nor NOR3 (N152, N149, N4, N122);
xor XOR2 (N153, N136, N112);
or OR4 (N154, N146, N6, N2, N78);
nor NOR4 (N155, N154, N51, N119, N151);
xor XOR2 (N156, N49, N11);
or OR2 (N157, N153, N84);
xor XOR2 (N158, N152, N150);
or OR3 (N159, N17, N16, N21);
xor XOR2 (N160, N159, N75);
xor XOR2 (N161, N139, N34);
or OR4 (N162, N147, N51, N34, N38);
buf BUF1 (N163, N161);
nor NOR3 (N164, N162, N5, N10);
nand NAND4 (N165, N156, N53, N98, N73);
not NOT1 (N166, N148);
buf BUF1 (N167, N163);
nand NAND2 (N168, N160, N40);
xor XOR2 (N169, N164, N136);
buf BUF1 (N170, N168);
nor NOR2 (N171, N166, N55);
buf BUF1 (N172, N171);
nand NAND4 (N173, N169, N161, N134, N122);
or OR3 (N174, N40, N136, N35);
or OR4 (N175, N165, N27, N138, N61);
xor XOR2 (N176, N158, N87);
xor XOR2 (N177, N95, N6);
nand NAND3 (N178, N167, N70, N34);
xor XOR2 (N179, N155, N1);
nor NOR2 (N180, N172, N25);
not NOT1 (N181, N177);
xor XOR2 (N182, N176, N121);
buf BUF1 (N183, N181);
not NOT1 (N184, N182);
not NOT1 (N185, N178);
nand NAND4 (N186, N183, N137, N80, N171);
xor XOR2 (N187, N186, N179);
not NOT1 (N188, N111);
and AND3 (N189, N173, N146, N20);
buf BUF1 (N190, N174);
not NOT1 (N191, N190);
not NOT1 (N192, N189);
buf BUF1 (N193, N180);
nand NAND2 (N194, N175, N33);
or OR2 (N195, N191, N89);
xor XOR2 (N196, N188, N187);
nand NAND3 (N197, N46, N110, N196);
not NOT1 (N198, N114);
and AND2 (N199, N170, N163);
nor NOR3 (N200, N199, N36, N107);
buf BUF1 (N201, N194);
nor NOR4 (N202, N200, N181, N87, N1);
nand NAND3 (N203, N184, N16, N110);
not NOT1 (N204, N195);
nand NAND4 (N205, N204, N39, N167, N13);
not NOT1 (N206, N192);
buf BUF1 (N207, N202);
xor XOR2 (N208, N201, N74);
nand NAND4 (N209, N157, N41, N97, N106);
and AND2 (N210, N193, N202);
buf BUF1 (N211, N198);
not NOT1 (N212, N185);
buf BUF1 (N213, N203);
or OR4 (N214, N208, N115, N63, N175);
and AND4 (N215, N211, N37, N136, N171);
xor XOR2 (N216, N215, N82);
buf BUF1 (N217, N205);
buf BUF1 (N218, N210);
and AND3 (N219, N212, N22, N132);
xor XOR2 (N220, N206, N74);
or OR2 (N221, N209, N198);
or OR2 (N222, N216, N39);
buf BUF1 (N223, N220);
nand NAND2 (N224, N214, N92);
or OR2 (N225, N219, N128);
or OR4 (N226, N207, N16, N134, N206);
and AND4 (N227, N226, N133, N136, N148);
and AND2 (N228, N218, N205);
not NOT1 (N229, N222);
xor XOR2 (N230, N224, N149);
and AND2 (N231, N217, N155);
xor XOR2 (N232, N229, N113);
and AND4 (N233, N223, N224, N180, N202);
and AND2 (N234, N231, N183);
buf BUF1 (N235, N233);
buf BUF1 (N236, N221);
not NOT1 (N237, N197);
and AND3 (N238, N227, N182, N96);
or OR3 (N239, N237, N102, N159);
nand NAND4 (N240, N232, N125, N7, N29);
xor XOR2 (N241, N213, N56);
buf BUF1 (N242, N228);
nor NOR3 (N243, N230, N75, N148);
not NOT1 (N244, N242);
and AND3 (N245, N241, N219, N82);
buf BUF1 (N246, N240);
and AND4 (N247, N236, N140, N152, N90);
or OR2 (N248, N239, N194);
nand NAND3 (N249, N244, N90, N189);
not NOT1 (N250, N243);
or OR2 (N251, N249, N192);
buf BUF1 (N252, N246);
xor XOR2 (N253, N247, N215);
not NOT1 (N254, N225);
nor NOR3 (N255, N254, N146, N112);
or OR2 (N256, N238, N9);
nand NAND4 (N257, N234, N65, N173, N92);
or OR4 (N258, N248, N162, N120, N51);
buf BUF1 (N259, N255);
not NOT1 (N260, N253);
xor XOR2 (N261, N251, N62);
and AND3 (N262, N261, N29, N219);
not NOT1 (N263, N252);
not NOT1 (N264, N257);
not NOT1 (N265, N264);
xor XOR2 (N266, N259, N167);
buf BUF1 (N267, N260);
nor NOR3 (N268, N263, N136, N255);
and AND3 (N269, N250, N222, N152);
xor XOR2 (N270, N235, N210);
buf BUF1 (N271, N267);
not NOT1 (N272, N266);
not NOT1 (N273, N265);
or OR2 (N274, N269, N8);
nor NOR2 (N275, N270, N212);
buf BUF1 (N276, N258);
nand NAND4 (N277, N256, N22, N2, N172);
nand NAND2 (N278, N274, N234);
nand NAND3 (N279, N262, N117, N5);
or OR4 (N280, N272, N74, N196, N6);
and AND3 (N281, N280, N73, N68);
xor XOR2 (N282, N275, N52);
nand NAND2 (N283, N278, N112);
nand NAND3 (N284, N276, N264, N268);
or OR4 (N285, N256, N159, N19, N65);
buf BUF1 (N286, N279);
not NOT1 (N287, N285);
nand NAND3 (N288, N284, N86, N134);
or OR2 (N289, N277, N122);
nor NOR3 (N290, N281, N118, N218);
not NOT1 (N291, N283);
nand NAND4 (N292, N290, N189, N180, N243);
or OR4 (N293, N286, N5, N104, N177);
not NOT1 (N294, N293);
buf BUF1 (N295, N291);
xor XOR2 (N296, N294, N100);
and AND3 (N297, N271, N21, N188);
or OR4 (N298, N245, N138, N223, N273);
xor XOR2 (N299, N80, N6);
xor XOR2 (N300, N287, N64);
buf BUF1 (N301, N297);
nand NAND3 (N302, N282, N36, N10);
buf BUF1 (N303, N298);
or OR4 (N304, N303, N65, N168, N79);
or OR3 (N305, N302, N133, N81);
buf BUF1 (N306, N288);
and AND4 (N307, N306, N286, N73, N20);
and AND4 (N308, N296, N90, N235, N47);
buf BUF1 (N309, N295);
not NOT1 (N310, N300);
nor NOR3 (N311, N304, N122, N267);
and AND4 (N312, N310, N84, N231, N8);
xor XOR2 (N313, N312, N77);
and AND3 (N314, N305, N139, N280);
buf BUF1 (N315, N313);
nor NOR3 (N316, N301, N210, N98);
and AND3 (N317, N315, N144, N306);
and AND3 (N318, N292, N160, N260);
nand NAND3 (N319, N317, N302, N133);
not NOT1 (N320, N318);
nor NOR4 (N321, N314, N16, N95, N237);
not NOT1 (N322, N319);
not NOT1 (N323, N316);
buf BUF1 (N324, N309);
and AND2 (N325, N307, N159);
and AND4 (N326, N320, N187, N257, N179);
or OR3 (N327, N321, N179, N217);
nor NOR4 (N328, N299, N166, N102, N181);
buf BUF1 (N329, N308);
nand NAND3 (N330, N324, N71, N245);
or OR3 (N331, N323, N72, N255);
buf BUF1 (N332, N322);
xor XOR2 (N333, N330, N103);
buf BUF1 (N334, N332);
xor XOR2 (N335, N329, N106);
nand NAND2 (N336, N333, N124);
nor NOR3 (N337, N336, N302, N218);
xor XOR2 (N338, N337, N82);
buf BUF1 (N339, N335);
nor NOR3 (N340, N334, N45, N289);
buf BUF1 (N341, N248);
or OR2 (N342, N327, N36);
not NOT1 (N343, N342);
nand NAND3 (N344, N311, N290, N91);
buf BUF1 (N345, N341);
buf BUF1 (N346, N338);
buf BUF1 (N347, N325);
or OR3 (N348, N346, N95, N186);
nand NAND2 (N349, N331, N96);
nand NAND2 (N350, N343, N73);
xor XOR2 (N351, N344, N85);
nor NOR3 (N352, N326, N230, N144);
buf BUF1 (N353, N339);
nand NAND3 (N354, N345, N50, N314);
not NOT1 (N355, N340);
buf BUF1 (N356, N347);
or OR4 (N357, N351, N37, N52, N135);
buf BUF1 (N358, N350);
or OR2 (N359, N353, N231);
nand NAND2 (N360, N328, N53);
nand NAND2 (N361, N352, N13);
nor NOR4 (N362, N355, N311, N348, N262);
nand NAND2 (N363, N76, N26);
nor NOR4 (N364, N361, N166, N236, N135);
or OR2 (N365, N357, N227);
nor NOR4 (N366, N360, N57, N182, N105);
nor NOR2 (N367, N363, N256);
xor XOR2 (N368, N349, N25);
or OR4 (N369, N364, N35, N215, N123);
and AND3 (N370, N365, N215, N365);
xor XOR2 (N371, N368, N75);
not NOT1 (N372, N362);
nor NOR3 (N373, N370, N61, N11);
buf BUF1 (N374, N371);
or OR4 (N375, N354, N20, N348, N325);
buf BUF1 (N376, N356);
nand NAND4 (N377, N358, N297, N88, N352);
and AND3 (N378, N375, N152, N260);
xor XOR2 (N379, N378, N71);
or OR2 (N380, N359, N228);
nor NOR3 (N381, N373, N93, N189);
nand NAND3 (N382, N379, N315, N89);
nand NAND2 (N383, N366, N207);
buf BUF1 (N384, N369);
and AND3 (N385, N383, N378, N358);
nor NOR2 (N386, N372, N48);
or OR2 (N387, N385, N217);
xor XOR2 (N388, N381, N154);
nor NOR4 (N389, N380, N85, N216, N80);
nor NOR3 (N390, N388, N148, N101);
nand NAND3 (N391, N390, N376, N65);
and AND4 (N392, N196, N255, N228, N183);
xor XOR2 (N393, N387, N375);
nor NOR3 (N394, N377, N304, N151);
not NOT1 (N395, N394);
nor NOR4 (N396, N389, N138, N347, N257);
xor XOR2 (N397, N392, N301);
and AND4 (N398, N386, N226, N37, N234);
not NOT1 (N399, N393);
not NOT1 (N400, N395);
or OR4 (N401, N396, N393, N151, N226);
nor NOR2 (N402, N401, N85);
and AND3 (N403, N391, N327, N160);
buf BUF1 (N404, N374);
nand NAND4 (N405, N384, N273, N330, N71);
or OR2 (N406, N399, N115);
buf BUF1 (N407, N398);
nor NOR2 (N408, N406, N302);
and AND2 (N409, N367, N397);
buf BUF1 (N410, N171);
or OR3 (N411, N408, N51, N353);
not NOT1 (N412, N400);
not NOT1 (N413, N403);
and AND2 (N414, N410, N14);
or OR2 (N415, N412, N278);
or OR3 (N416, N413, N137, N283);
not NOT1 (N417, N407);
nand NAND2 (N418, N409, N93);
not NOT1 (N419, N405);
xor XOR2 (N420, N414, N384);
nand NAND4 (N421, N402, N60, N304, N346);
not NOT1 (N422, N416);
nor NOR4 (N423, N417, N380, N56, N395);
nand NAND3 (N424, N404, N75, N234);
and AND4 (N425, N420, N16, N328, N38);
and AND4 (N426, N415, N83, N174, N364);
nand NAND2 (N427, N424, N33);
or OR4 (N428, N427, N78, N287, N13);
buf BUF1 (N429, N421);
nand NAND3 (N430, N418, N146, N310);
nand NAND4 (N431, N425, N417, N203, N49);
or OR2 (N432, N423, N352);
nand NAND2 (N433, N422, N19);
and AND2 (N434, N429, N328);
and AND4 (N435, N382, N319, N404, N83);
buf BUF1 (N436, N430);
xor XOR2 (N437, N434, N341);
xor XOR2 (N438, N432, N288);
nand NAND3 (N439, N428, N145, N244);
nor NOR3 (N440, N433, N405, N242);
nand NAND3 (N441, N438, N63, N264);
and AND2 (N442, N439, N72);
nor NOR2 (N443, N431, N415);
nor NOR3 (N444, N441, N8, N58);
xor XOR2 (N445, N437, N275);
buf BUF1 (N446, N442);
nor NOR3 (N447, N436, N293, N211);
or OR3 (N448, N419, N333, N296);
and AND2 (N449, N440, N171);
and AND2 (N450, N447, N99);
and AND2 (N451, N445, N63);
xor XOR2 (N452, N451, N302);
nand NAND3 (N453, N448, N162, N244);
xor XOR2 (N454, N435, N92);
nand NAND2 (N455, N450, N248);
not NOT1 (N456, N449);
buf BUF1 (N457, N452);
buf BUF1 (N458, N457);
nor NOR2 (N459, N411, N196);
not NOT1 (N460, N456);
nor NOR4 (N461, N426, N374, N38, N115);
nor NOR3 (N462, N458, N237, N205);
xor XOR2 (N463, N444, N391);
not NOT1 (N464, N459);
and AND2 (N465, N463, N421);
xor XOR2 (N466, N455, N316);
and AND2 (N467, N461, N430);
buf BUF1 (N468, N466);
buf BUF1 (N469, N460);
nor NOR4 (N470, N454, N193, N299, N157);
nand NAND2 (N471, N443, N231);
not NOT1 (N472, N462);
or OR2 (N473, N469, N370);
and AND4 (N474, N446, N45, N392, N56);
nand NAND4 (N475, N467, N407, N288, N241);
nor NOR2 (N476, N465, N273);
or OR2 (N477, N468, N94);
and AND3 (N478, N473, N368, N345);
buf BUF1 (N479, N474);
or OR4 (N480, N475, N112, N233, N415);
or OR3 (N481, N479, N28, N261);
or OR4 (N482, N464, N11, N159, N412);
and AND2 (N483, N481, N295);
xor XOR2 (N484, N472, N209);
xor XOR2 (N485, N478, N462);
and AND3 (N486, N482, N236, N328);
xor XOR2 (N487, N484, N22);
or OR4 (N488, N480, N107, N175, N274);
nor NOR3 (N489, N485, N402, N244);
nor NOR2 (N490, N487, N75);
nand NAND4 (N491, N453, N461, N222, N187);
not NOT1 (N492, N470);
xor XOR2 (N493, N471, N417);
xor XOR2 (N494, N491, N217);
or OR3 (N495, N488, N155, N355);
buf BUF1 (N496, N495);
not NOT1 (N497, N490);
xor XOR2 (N498, N493, N293);
or OR3 (N499, N498, N24, N122);
and AND3 (N500, N494, N141, N465);
buf BUF1 (N501, N489);
or OR2 (N502, N499, N329);
nand NAND3 (N503, N500, N62, N287);
or OR3 (N504, N492, N53, N302);
and AND2 (N505, N496, N283);
xor XOR2 (N506, N476, N217);
and AND4 (N507, N506, N117, N214, N361);
nand NAND3 (N508, N477, N290, N356);
nand NAND3 (N509, N505, N69, N503);
not NOT1 (N510, N184);
or OR4 (N511, N510, N464, N303, N197);
and AND2 (N512, N509, N239);
not NOT1 (N513, N504);
not NOT1 (N514, N512);
not NOT1 (N515, N514);
and AND3 (N516, N501, N110, N9);
nand NAND4 (N517, N508, N246, N450, N472);
not NOT1 (N518, N513);
xor XOR2 (N519, N517, N6);
buf BUF1 (N520, N507);
xor XOR2 (N521, N511, N97);
or OR4 (N522, N497, N28, N370, N57);
not NOT1 (N523, N521);
buf BUF1 (N524, N519);
nand NAND3 (N525, N524, N383, N381);
buf BUF1 (N526, N515);
xor XOR2 (N527, N520, N141);
xor XOR2 (N528, N502, N226);
nand NAND2 (N529, N516, N523);
nand NAND3 (N530, N270, N479, N171);
xor XOR2 (N531, N528, N103);
buf BUF1 (N532, N522);
or OR4 (N533, N483, N451, N8, N197);
and AND4 (N534, N525, N139, N137, N384);
and AND4 (N535, N531, N254, N176, N194);
xor XOR2 (N536, N532, N205);
buf BUF1 (N537, N486);
nor NOR4 (N538, N535, N409, N426, N287);
buf BUF1 (N539, N530);
or OR2 (N540, N518, N117);
not NOT1 (N541, N529);
not NOT1 (N542, N527);
nor NOR2 (N543, N533, N259);
nor NOR3 (N544, N526, N92, N30);
xor XOR2 (N545, N537, N541);
nand NAND4 (N546, N262, N303, N325, N520);
buf BUF1 (N547, N542);
xor XOR2 (N548, N544, N67);
not NOT1 (N549, N540);
xor XOR2 (N550, N543, N364);
nor NOR3 (N551, N534, N489, N257);
or OR4 (N552, N551, N7, N148, N297);
nor NOR3 (N553, N536, N366, N470);
or OR3 (N554, N553, N258, N255);
xor XOR2 (N555, N550, N535);
not NOT1 (N556, N552);
or OR2 (N557, N539, N428);
nand NAND3 (N558, N546, N160, N511);
or OR4 (N559, N548, N20, N432, N313);
or OR4 (N560, N559, N93, N514, N477);
and AND4 (N561, N554, N47, N545, N407);
or OR2 (N562, N108, N160);
or OR4 (N563, N555, N434, N83, N290);
nor NOR3 (N564, N549, N18, N37);
nor NOR4 (N565, N560, N319, N89, N439);
nor NOR2 (N566, N561, N383);
buf BUF1 (N567, N538);
and AND2 (N568, N558, N339);
xor XOR2 (N569, N547, N53);
xor XOR2 (N570, N567, N451);
xor XOR2 (N571, N562, N422);
not NOT1 (N572, N571);
nand NAND2 (N573, N556, N441);
nor NOR3 (N574, N572, N490, N160);
nor NOR4 (N575, N569, N180, N45, N465);
not NOT1 (N576, N575);
buf BUF1 (N577, N568);
nor NOR2 (N578, N566, N271);
or OR4 (N579, N570, N262, N396, N166);
nand NAND3 (N580, N574, N79, N561);
nand NAND2 (N581, N563, N128);
and AND4 (N582, N564, N452, N369, N423);
nand NAND4 (N583, N573, N562, N345, N494);
nor NOR2 (N584, N578, N264);
and AND2 (N585, N577, N261);
or OR3 (N586, N579, N322, N424);
or OR4 (N587, N583, N196, N248, N570);
buf BUF1 (N588, N585);
and AND4 (N589, N581, N304, N200, N526);
not NOT1 (N590, N586);
nand NAND4 (N591, N587, N390, N479, N257);
nor NOR2 (N592, N584, N481);
or OR2 (N593, N589, N117);
buf BUF1 (N594, N593);
not NOT1 (N595, N594);
and AND4 (N596, N595, N589, N368, N537);
not NOT1 (N597, N557);
nor NOR3 (N598, N597, N84, N534);
nand NAND3 (N599, N592, N24, N466);
and AND3 (N600, N565, N76, N82);
xor XOR2 (N601, N600, N340);
nor NOR3 (N602, N599, N347, N377);
buf BUF1 (N603, N590);
buf BUF1 (N604, N603);
nand NAND2 (N605, N580, N518);
and AND2 (N606, N598, N226);
nand NAND3 (N607, N591, N409, N55);
nand NAND2 (N608, N606, N340);
nand NAND3 (N609, N596, N24, N203);
not NOT1 (N610, N582);
buf BUF1 (N611, N576);
xor XOR2 (N612, N608, N141);
or OR3 (N613, N605, N348, N362);
buf BUF1 (N614, N610);
nand NAND4 (N615, N604, N362, N204, N604);
xor XOR2 (N616, N613, N97);
or OR2 (N617, N614, N537);
xor XOR2 (N618, N615, N381);
xor XOR2 (N619, N588, N336);
buf BUF1 (N620, N607);
nand NAND4 (N621, N609, N612, N399, N508);
nand NAND2 (N622, N273, N96);
and AND3 (N623, N622, N540, N53);
nor NOR2 (N624, N620, N105);
not NOT1 (N625, N601);
and AND2 (N626, N619, N344);
nor NOR3 (N627, N623, N13, N510);
not NOT1 (N628, N626);
and AND3 (N629, N625, N42, N418);
xor XOR2 (N630, N627, N60);
nor NOR2 (N631, N628, N538);
not NOT1 (N632, N602);
not NOT1 (N633, N629);
xor XOR2 (N634, N611, N414);
nand NAND4 (N635, N632, N364, N565, N580);
and AND3 (N636, N634, N204, N616);
not NOT1 (N637, N125);
nor NOR4 (N638, N624, N380, N95, N65);
buf BUF1 (N639, N631);
not NOT1 (N640, N635);
nand NAND3 (N641, N633, N30, N294);
not NOT1 (N642, N636);
and AND2 (N643, N641, N164);
nand NAND4 (N644, N640, N471, N182, N533);
or OR4 (N645, N617, N68, N359, N617);
or OR4 (N646, N621, N233, N250, N610);
nor NOR4 (N647, N646, N177, N16, N548);
or OR4 (N648, N642, N354, N176, N566);
buf BUF1 (N649, N643);
buf BUF1 (N650, N638);
or OR2 (N651, N649, N46);
xor XOR2 (N652, N651, N183);
xor XOR2 (N653, N618, N643);
or OR2 (N654, N652, N163);
nand NAND2 (N655, N639, N122);
xor XOR2 (N656, N647, N543);
buf BUF1 (N657, N630);
not NOT1 (N658, N657);
and AND3 (N659, N654, N592, N387);
nand NAND4 (N660, N637, N218, N221, N642);
nand NAND4 (N661, N660, N460, N300, N277);
and AND4 (N662, N655, N506, N513, N412);
or OR4 (N663, N653, N636, N125, N289);
or OR3 (N664, N656, N161, N208);
xor XOR2 (N665, N658, N615);
or OR2 (N666, N648, N650);
or OR4 (N667, N190, N7, N547, N420);
nor NOR4 (N668, N662, N155, N445, N429);
buf BUF1 (N669, N645);
xor XOR2 (N670, N644, N624);
or OR3 (N671, N667, N315, N359);
nand NAND2 (N672, N671, N332);
buf BUF1 (N673, N661);
xor XOR2 (N674, N668, N479);
xor XOR2 (N675, N666, N332);
nor NOR2 (N676, N669, N667);
and AND3 (N677, N665, N262, N519);
nor NOR4 (N678, N672, N415, N405, N5);
nor NOR3 (N679, N659, N85, N306);
and AND3 (N680, N678, N603, N570);
nor NOR3 (N681, N676, N469, N676);
or OR2 (N682, N674, N26);
buf BUF1 (N683, N663);
xor XOR2 (N684, N675, N452);
not NOT1 (N685, N679);
not NOT1 (N686, N685);
xor XOR2 (N687, N686, N291);
or OR4 (N688, N664, N490, N94, N405);
and AND3 (N689, N677, N273, N216);
xor XOR2 (N690, N670, N568);
nor NOR2 (N691, N687, N184);
not NOT1 (N692, N689);
not NOT1 (N693, N692);
or OR3 (N694, N682, N130, N449);
xor XOR2 (N695, N693, N413);
nand NAND4 (N696, N683, N446, N313, N254);
or OR4 (N697, N680, N353, N312, N528);
nor NOR3 (N698, N681, N492, N417);
not NOT1 (N699, N691);
nor NOR4 (N700, N688, N23, N361, N618);
or OR4 (N701, N697, N311, N49, N449);
xor XOR2 (N702, N694, N630);
nor NOR3 (N703, N684, N250, N132);
nor NOR4 (N704, N696, N34, N42, N300);
nand NAND3 (N705, N704, N519, N246);
xor XOR2 (N706, N701, N695);
not NOT1 (N707, N400);
or OR2 (N708, N705, N464);
xor XOR2 (N709, N702, N166);
buf BUF1 (N710, N708);
and AND3 (N711, N703, N551, N285);
nor NOR3 (N712, N698, N564, N292);
not NOT1 (N713, N707);
not NOT1 (N714, N711);
not NOT1 (N715, N690);
nor NOR2 (N716, N709, N358);
or OR2 (N717, N716, N700);
nor NOR3 (N718, N436, N43, N659);
buf BUF1 (N719, N706);
nor NOR4 (N720, N719, N131, N174, N458);
and AND3 (N721, N715, N449, N644);
nor NOR4 (N722, N712, N636, N397, N692);
not NOT1 (N723, N717);
and AND2 (N724, N721, N553);
xor XOR2 (N725, N723, N320);
nor NOR3 (N726, N720, N383, N331);
buf BUF1 (N727, N726);
and AND4 (N728, N727, N197, N29, N671);
and AND2 (N729, N714, N371);
and AND3 (N730, N728, N125, N182);
nand NAND4 (N731, N713, N717, N275, N188);
nand NAND4 (N732, N710, N46, N598, N244);
or OR4 (N733, N673, N487, N562, N423);
buf BUF1 (N734, N733);
not NOT1 (N735, N722);
not NOT1 (N736, N732);
not NOT1 (N737, N724);
buf BUF1 (N738, N734);
nor NOR3 (N739, N729, N236, N157);
xor XOR2 (N740, N735, N292);
or OR3 (N741, N730, N342, N226);
nor NOR2 (N742, N736, N362);
nand NAND4 (N743, N699, N645, N2, N663);
nand NAND4 (N744, N742, N456, N687, N647);
xor XOR2 (N745, N731, N556);
or OR3 (N746, N718, N226, N503);
nand NAND2 (N747, N745, N539);
buf BUF1 (N748, N738);
and AND4 (N749, N725, N400, N712, N421);
and AND4 (N750, N746, N521, N174, N446);
nor NOR4 (N751, N747, N320, N67, N543);
nor NOR4 (N752, N750, N260, N119, N599);
buf BUF1 (N753, N740);
buf BUF1 (N754, N749);
xor XOR2 (N755, N748, N601);
or OR3 (N756, N737, N469, N167);
and AND2 (N757, N751, N377);
nand NAND3 (N758, N739, N423, N636);
buf BUF1 (N759, N744);
nand NAND3 (N760, N757, N285, N436);
and AND3 (N761, N743, N682, N201);
nor NOR3 (N762, N759, N405, N226);
not NOT1 (N763, N762);
not NOT1 (N764, N763);
buf BUF1 (N765, N764);
and AND3 (N766, N756, N446, N223);
or OR2 (N767, N766, N97);
nand NAND3 (N768, N755, N492, N360);
buf BUF1 (N769, N767);
nand NAND3 (N770, N752, N463, N106);
xor XOR2 (N771, N761, N718);
nand NAND3 (N772, N768, N396, N629);
and AND3 (N773, N772, N110, N481);
and AND4 (N774, N765, N337, N157, N338);
nor NOR4 (N775, N758, N131, N324, N71);
nor NOR3 (N776, N741, N106, N285);
or OR4 (N777, N769, N630, N632, N683);
xor XOR2 (N778, N770, N114);
xor XOR2 (N779, N760, N551);
nor NOR2 (N780, N775, N503);
nor NOR2 (N781, N774, N767);
buf BUF1 (N782, N773);
buf BUF1 (N783, N781);
buf BUF1 (N784, N778);
or OR3 (N785, N779, N650, N217);
buf BUF1 (N786, N777);
buf BUF1 (N787, N780);
xor XOR2 (N788, N782, N155);
not NOT1 (N789, N754);
and AND4 (N790, N788, N321, N595, N655);
and AND4 (N791, N783, N115, N727, N421);
buf BUF1 (N792, N784);
and AND3 (N793, N787, N252, N348);
xor XOR2 (N794, N786, N780);
or OR2 (N795, N789, N12);
nor NOR3 (N796, N753, N459, N18);
and AND3 (N797, N793, N605, N357);
and AND2 (N798, N794, N177);
xor XOR2 (N799, N791, N647);
buf BUF1 (N800, N792);
or OR4 (N801, N776, N447, N609, N433);
buf BUF1 (N802, N795);
or OR2 (N803, N802, N606);
or OR2 (N804, N785, N372);
buf BUF1 (N805, N799);
nor NOR4 (N806, N797, N713, N370, N336);
and AND2 (N807, N790, N585);
not NOT1 (N808, N798);
buf BUF1 (N809, N771);
and AND2 (N810, N807, N217);
and AND2 (N811, N809, N267);
or OR3 (N812, N803, N29, N237);
buf BUF1 (N813, N801);
nand NAND3 (N814, N810, N357, N54);
nor NOR4 (N815, N806, N603, N419, N145);
nand NAND3 (N816, N812, N389, N196);
nor NOR2 (N817, N805, N692);
or OR2 (N818, N804, N160);
not NOT1 (N819, N815);
buf BUF1 (N820, N813);
not NOT1 (N821, N796);
nand NAND4 (N822, N814, N327, N304, N181);
nand NAND4 (N823, N822, N545, N547, N771);
nand NAND3 (N824, N816, N746, N174);
and AND4 (N825, N808, N587, N30, N482);
buf BUF1 (N826, N824);
xor XOR2 (N827, N820, N12);
buf BUF1 (N828, N818);
nor NOR4 (N829, N828, N19, N789, N689);
nand NAND4 (N830, N826, N354, N559, N419);
not NOT1 (N831, N811);
buf BUF1 (N832, N823);
xor XOR2 (N833, N819, N119);
buf BUF1 (N834, N829);
or OR3 (N835, N831, N249, N754);
xor XOR2 (N836, N835, N60);
nand NAND4 (N837, N833, N205, N527, N362);
and AND3 (N838, N800, N244, N637);
not NOT1 (N839, N838);
or OR4 (N840, N834, N541, N624, N623);
nor NOR2 (N841, N837, N660);
xor XOR2 (N842, N830, N822);
nor NOR2 (N843, N836, N826);
nor NOR4 (N844, N817, N391, N526, N521);
xor XOR2 (N845, N827, N433);
not NOT1 (N846, N825);
or OR4 (N847, N844, N638, N581, N468);
not NOT1 (N848, N839);
nor NOR4 (N849, N842, N2, N826, N819);
nand NAND4 (N850, N849, N61, N216, N790);
xor XOR2 (N851, N847, N354);
nor NOR3 (N852, N851, N523, N749);
xor XOR2 (N853, N848, N287);
nand NAND4 (N854, N852, N159, N478, N111);
not NOT1 (N855, N832);
and AND4 (N856, N850, N213, N725, N136);
nor NOR3 (N857, N845, N607, N234);
and AND2 (N858, N857, N657);
or OR3 (N859, N821, N620, N117);
or OR4 (N860, N856, N466, N834, N119);
not NOT1 (N861, N858);
or OR3 (N862, N853, N320, N205);
buf BUF1 (N863, N859);
not NOT1 (N864, N840);
and AND2 (N865, N846, N293);
not NOT1 (N866, N863);
buf BUF1 (N867, N862);
nand NAND3 (N868, N855, N501, N77);
nor NOR4 (N869, N865, N484, N79, N127);
xor XOR2 (N870, N841, N29);
and AND2 (N871, N867, N190);
and AND3 (N872, N868, N29, N316);
nor NOR3 (N873, N872, N814, N491);
xor XOR2 (N874, N869, N619);
nor NOR3 (N875, N854, N778, N868);
not NOT1 (N876, N874);
nand NAND3 (N877, N875, N539, N531);
nand NAND2 (N878, N871, N550);
buf BUF1 (N879, N864);
xor XOR2 (N880, N873, N295);
and AND4 (N881, N879, N479, N291, N262);
not NOT1 (N882, N870);
not NOT1 (N883, N861);
and AND4 (N884, N866, N213, N357, N321);
xor XOR2 (N885, N880, N237);
and AND2 (N886, N878, N877);
and AND2 (N887, N466, N380);
or OR3 (N888, N887, N700, N113);
buf BUF1 (N889, N882);
buf BUF1 (N890, N888);
not NOT1 (N891, N883);
and AND3 (N892, N889, N715, N489);
nand NAND2 (N893, N881, N414);
and AND4 (N894, N892, N183, N739, N499);
and AND4 (N895, N890, N383, N366, N639);
nand NAND3 (N896, N884, N251, N118);
nand NAND3 (N897, N896, N680, N99);
nand NAND2 (N898, N860, N196);
nor NOR2 (N899, N886, N598);
xor XOR2 (N900, N891, N791);
or OR4 (N901, N895, N385, N847, N843);
buf BUF1 (N902, N817);
nor NOR3 (N903, N885, N888, N872);
nand NAND4 (N904, N902, N333, N92, N585);
not NOT1 (N905, N903);
not NOT1 (N906, N899);
xor XOR2 (N907, N904, N231);
or OR2 (N908, N900, N561);
nor NOR3 (N909, N893, N222, N332);
xor XOR2 (N910, N901, N509);
and AND3 (N911, N897, N713, N286);
xor XOR2 (N912, N911, N647);
nand NAND3 (N913, N876, N201, N483);
nor NOR3 (N914, N910, N770, N721);
or OR4 (N915, N907, N418, N476, N496);
nand NAND2 (N916, N908, N248);
nand NAND4 (N917, N906, N840, N319, N892);
nand NAND4 (N918, N913, N379, N661, N796);
not NOT1 (N919, N898);
nand NAND3 (N920, N916, N776, N916);
and AND4 (N921, N919, N248, N715, N828);
nand NAND4 (N922, N921, N377, N509, N439);
not NOT1 (N923, N917);
or OR3 (N924, N918, N416, N255);
xor XOR2 (N925, N923, N522);
and AND3 (N926, N915, N527, N101);
xor XOR2 (N927, N925, N219);
nor NOR4 (N928, N894, N505, N187, N1);
buf BUF1 (N929, N909);
nand NAND2 (N930, N920, N614);
nor NOR2 (N931, N912, N246);
and AND2 (N932, N928, N607);
nand NAND4 (N933, N929, N219, N419, N211);
not NOT1 (N934, N905);
nand NAND2 (N935, N926, N156);
nand NAND3 (N936, N914, N899, N688);
xor XOR2 (N937, N934, N500);
nor NOR2 (N938, N933, N348);
and AND4 (N939, N930, N682, N160, N733);
buf BUF1 (N940, N935);
not NOT1 (N941, N939);
nor NOR3 (N942, N936, N808, N509);
nor NOR2 (N943, N927, N864);
nor NOR2 (N944, N931, N3);
not NOT1 (N945, N944);
buf BUF1 (N946, N938);
nand NAND3 (N947, N942, N775, N589);
not NOT1 (N948, N947);
and AND4 (N949, N946, N503, N589, N891);
or OR4 (N950, N940, N389, N656, N191);
xor XOR2 (N951, N932, N308);
or OR2 (N952, N943, N304);
xor XOR2 (N953, N949, N716);
xor XOR2 (N954, N950, N888);
or OR3 (N955, N922, N803, N701);
nand NAND4 (N956, N955, N233, N450, N787);
buf BUF1 (N957, N945);
nand NAND4 (N958, N954, N220, N386, N84);
and AND3 (N959, N952, N891, N886);
not NOT1 (N960, N956);
or OR2 (N961, N960, N905);
and AND2 (N962, N953, N140);
and AND4 (N963, N959, N814, N228, N648);
nand NAND3 (N964, N961, N605, N875);
nand NAND4 (N965, N957, N170, N955, N912);
not NOT1 (N966, N948);
or OR4 (N967, N965, N150, N963, N99);
nor NOR3 (N968, N19, N416, N724);
or OR3 (N969, N967, N545, N443);
not NOT1 (N970, N924);
nor NOR2 (N971, N966, N922);
or OR3 (N972, N964, N282, N618);
not NOT1 (N973, N941);
nand NAND3 (N974, N937, N593, N454);
and AND4 (N975, N972, N23, N135, N212);
xor XOR2 (N976, N968, N688);
xor XOR2 (N977, N958, N436);
or OR3 (N978, N973, N697, N358);
xor XOR2 (N979, N969, N378);
nand NAND3 (N980, N976, N574, N50);
xor XOR2 (N981, N971, N574);
and AND2 (N982, N979, N314);
nand NAND4 (N983, N980, N118, N234, N893);
xor XOR2 (N984, N978, N260);
nor NOR4 (N985, N977, N59, N978, N971);
not NOT1 (N986, N981);
buf BUF1 (N987, N984);
not NOT1 (N988, N975);
nand NAND4 (N989, N983, N227, N878, N49);
nand NAND4 (N990, N982, N736, N624, N409);
buf BUF1 (N991, N974);
not NOT1 (N992, N990);
not NOT1 (N993, N988);
nand NAND3 (N994, N987, N354, N547);
and AND4 (N995, N962, N199, N191, N289);
or OR2 (N996, N970, N302);
buf BUF1 (N997, N994);
nor NOR3 (N998, N951, N237, N621);
xor XOR2 (N999, N986, N300);
not NOT1 (N1000, N995);
not NOT1 (N1001, N993);
xor XOR2 (N1002, N1000, N774);
not NOT1 (N1003, N989);
and AND4 (N1004, N998, N302, N445, N1);
not NOT1 (N1005, N991);
and AND3 (N1006, N996, N976, N165);
and AND3 (N1007, N997, N331, N865);
not NOT1 (N1008, N1004);
not NOT1 (N1009, N1003);
and AND3 (N1010, N985, N603, N737);
and AND2 (N1011, N999, N43);
and AND2 (N1012, N1009, N781);
not NOT1 (N1013, N1001);
xor XOR2 (N1014, N1010, N559);
or OR2 (N1015, N1012, N755);
xor XOR2 (N1016, N1005, N150);
buf BUF1 (N1017, N1013);
xor XOR2 (N1018, N1008, N992);
not NOT1 (N1019, N76);
nand NAND3 (N1020, N1007, N787, N648);
not NOT1 (N1021, N1020);
buf BUF1 (N1022, N1014);
not NOT1 (N1023, N1018);
and AND3 (N1024, N1011, N205, N520);
buf BUF1 (N1025, N1023);
xor XOR2 (N1026, N1022, N962);
not NOT1 (N1027, N1024);
not NOT1 (N1028, N1026);
xor XOR2 (N1029, N1002, N635);
buf BUF1 (N1030, N1021);
not NOT1 (N1031, N1027);
and AND2 (N1032, N1019, N720);
nand NAND2 (N1033, N1028, N936);
or OR2 (N1034, N1015, N550);
nor NOR4 (N1035, N1030, N732, N875, N229);
not NOT1 (N1036, N1006);
nor NOR2 (N1037, N1034, N244);
nor NOR2 (N1038, N1031, N875);
nor NOR2 (N1039, N1038, N510);
and AND2 (N1040, N1037, N55);
buf BUF1 (N1041, N1017);
not NOT1 (N1042, N1040);
buf BUF1 (N1043, N1039);
xor XOR2 (N1044, N1016, N120);
or OR3 (N1045, N1035, N906, N971);
buf BUF1 (N1046, N1044);
not NOT1 (N1047, N1042);
or OR3 (N1048, N1033, N751, N850);
not NOT1 (N1049, N1041);
not NOT1 (N1050, N1029);
xor XOR2 (N1051, N1045, N532);
xor XOR2 (N1052, N1046, N660);
buf BUF1 (N1053, N1048);
xor XOR2 (N1054, N1049, N98);
not NOT1 (N1055, N1043);
nand NAND4 (N1056, N1051, N313, N567, N1025);
xor XOR2 (N1057, N923, N365);
xor XOR2 (N1058, N1054, N519);
or OR3 (N1059, N1052, N287, N505);
or OR3 (N1060, N1059, N403, N622);
not NOT1 (N1061, N1056);
nand NAND3 (N1062, N1055, N402, N420);
nor NOR3 (N1063, N1036, N201, N765);
xor XOR2 (N1064, N1053, N801);
and AND3 (N1065, N1047, N450, N914);
buf BUF1 (N1066, N1062);
and AND2 (N1067, N1057, N668);
not NOT1 (N1068, N1050);
nor NOR2 (N1069, N1063, N14);
buf BUF1 (N1070, N1066);
nor NOR2 (N1071, N1058, N1004);
not NOT1 (N1072, N1061);
buf BUF1 (N1073, N1071);
and AND4 (N1074, N1067, N543, N470, N105);
xor XOR2 (N1075, N1065, N468);
and AND3 (N1076, N1074, N1051, N179);
nand NAND2 (N1077, N1070, N70);
buf BUF1 (N1078, N1073);
nor NOR3 (N1079, N1069, N737, N98);
nand NAND3 (N1080, N1060, N234, N780);
nor NOR2 (N1081, N1072, N740);
not NOT1 (N1082, N1064);
xor XOR2 (N1083, N1079, N956);
nand NAND3 (N1084, N1083, N712, N937);
and AND3 (N1085, N1084, N536, N606);
nand NAND3 (N1086, N1082, N335, N1045);
nor NOR2 (N1087, N1085, N67);
nor NOR2 (N1088, N1087, N852);
xor XOR2 (N1089, N1076, N264);
or OR3 (N1090, N1075, N366, N926);
nor NOR2 (N1091, N1089, N942);
not NOT1 (N1092, N1080);
nor NOR3 (N1093, N1092, N327, N901);
and AND4 (N1094, N1090, N1057, N569, N431);
xor XOR2 (N1095, N1078, N461);
or OR4 (N1096, N1088, N1059, N331, N699);
nor NOR4 (N1097, N1068, N121, N473, N825);
not NOT1 (N1098, N1093);
nor NOR2 (N1099, N1086, N1025);
nand NAND3 (N1100, N1096, N632, N261);
not NOT1 (N1101, N1099);
nor NOR3 (N1102, N1032, N959, N842);
xor XOR2 (N1103, N1081, N344);
xor XOR2 (N1104, N1102, N403);
or OR2 (N1105, N1094, N313);
nor NOR3 (N1106, N1100, N266, N843);
buf BUF1 (N1107, N1095);
nand NAND2 (N1108, N1101, N294);
and AND3 (N1109, N1103, N387, N15);
and AND2 (N1110, N1105, N805);
buf BUF1 (N1111, N1108);
nor NOR3 (N1112, N1098, N834, N600);
nor NOR2 (N1113, N1106, N102);
nand NAND2 (N1114, N1091, N919);
nor NOR4 (N1115, N1110, N6, N992, N877);
buf BUF1 (N1116, N1112);
and AND2 (N1117, N1111, N701);
or OR3 (N1118, N1114, N325, N96);
xor XOR2 (N1119, N1107, N809);
not NOT1 (N1120, N1104);
xor XOR2 (N1121, N1113, N432);
nand NAND4 (N1122, N1097, N670, N285, N653);
not NOT1 (N1123, N1121);
xor XOR2 (N1124, N1120, N478);
nand NAND4 (N1125, N1115, N1008, N123, N870);
or OR2 (N1126, N1119, N291);
nor NOR3 (N1127, N1077, N236, N73);
or OR2 (N1128, N1123, N690);
or OR2 (N1129, N1126, N782);
or OR3 (N1130, N1129, N1037, N17);
xor XOR2 (N1131, N1116, N76);
nor NOR2 (N1132, N1122, N951);
and AND2 (N1133, N1125, N458);
or OR4 (N1134, N1118, N470, N331, N105);
xor XOR2 (N1135, N1117, N801);
and AND3 (N1136, N1131, N414, N311);
xor XOR2 (N1137, N1109, N688);
xor XOR2 (N1138, N1133, N920);
xor XOR2 (N1139, N1138, N216);
buf BUF1 (N1140, N1127);
and AND3 (N1141, N1136, N37, N192);
buf BUF1 (N1142, N1140);
not NOT1 (N1143, N1124);
nand NAND2 (N1144, N1137, N727);
not NOT1 (N1145, N1134);
not NOT1 (N1146, N1145);
buf BUF1 (N1147, N1141);
nor NOR2 (N1148, N1139, N188);
buf BUF1 (N1149, N1146);
or OR3 (N1150, N1144, N115, N367);
nand NAND2 (N1151, N1143, N545);
nand NAND4 (N1152, N1149, N374, N776, N228);
buf BUF1 (N1153, N1147);
nand NAND2 (N1154, N1151, N118);
and AND4 (N1155, N1154, N186, N836, N856);
not NOT1 (N1156, N1152);
not NOT1 (N1157, N1130);
buf BUF1 (N1158, N1148);
or OR3 (N1159, N1156, N605, N978);
not NOT1 (N1160, N1150);
not NOT1 (N1161, N1157);
and AND2 (N1162, N1128, N658);
and AND3 (N1163, N1158, N262, N386);
nor NOR2 (N1164, N1153, N83);
buf BUF1 (N1165, N1161);
nor NOR2 (N1166, N1159, N933);
xor XOR2 (N1167, N1132, N280);
or OR3 (N1168, N1167, N805, N349);
and AND2 (N1169, N1155, N148);
nor NOR2 (N1170, N1163, N414);
or OR3 (N1171, N1165, N862, N770);
and AND2 (N1172, N1171, N168);
xor XOR2 (N1173, N1169, N819);
xor XOR2 (N1174, N1135, N718);
buf BUF1 (N1175, N1142);
or OR3 (N1176, N1175, N932, N44);
nand NAND3 (N1177, N1162, N818, N499);
xor XOR2 (N1178, N1168, N166);
nor NOR4 (N1179, N1174, N159, N184, N510);
buf BUF1 (N1180, N1173);
nor NOR4 (N1181, N1166, N323, N282, N586);
nand NAND4 (N1182, N1180, N494, N945, N538);
or OR2 (N1183, N1181, N373);
or OR3 (N1184, N1183, N761, N455);
buf BUF1 (N1185, N1179);
or OR2 (N1186, N1170, N257);
nor NOR2 (N1187, N1184, N855);
not NOT1 (N1188, N1182);
xor XOR2 (N1189, N1178, N17);
buf BUF1 (N1190, N1189);
nor NOR3 (N1191, N1172, N909, N175);
or OR4 (N1192, N1160, N102, N1163, N1131);
xor XOR2 (N1193, N1186, N768);
buf BUF1 (N1194, N1177);
and AND3 (N1195, N1190, N596, N233);
and AND2 (N1196, N1194, N639);
not NOT1 (N1197, N1176);
nor NOR2 (N1198, N1195, N253);
and AND3 (N1199, N1193, N413, N1024);
not NOT1 (N1200, N1164);
xor XOR2 (N1201, N1191, N641);
or OR4 (N1202, N1185, N406, N154, N185);
or OR3 (N1203, N1196, N150, N475);
and AND3 (N1204, N1188, N200, N973);
buf BUF1 (N1205, N1187);
buf BUF1 (N1206, N1192);
nor NOR4 (N1207, N1203, N511, N823, N829);
nand NAND2 (N1208, N1204, N185);
and AND4 (N1209, N1200, N135, N817, N916);
nand NAND4 (N1210, N1201, N352, N900, N1072);
buf BUF1 (N1211, N1208);
buf BUF1 (N1212, N1205);
buf BUF1 (N1213, N1209);
and AND3 (N1214, N1212, N147, N349);
buf BUF1 (N1215, N1198);
or OR2 (N1216, N1202, N749);
and AND4 (N1217, N1211, N769, N1071, N1160);
xor XOR2 (N1218, N1213, N1138);
nand NAND4 (N1219, N1207, N1186, N675, N145);
xor XOR2 (N1220, N1199, N802);
xor XOR2 (N1221, N1216, N175);
nor NOR4 (N1222, N1210, N183, N310, N352);
nor NOR3 (N1223, N1197, N525, N931);
nor NOR2 (N1224, N1214, N575);
nand NAND2 (N1225, N1224, N459);
buf BUF1 (N1226, N1218);
buf BUF1 (N1227, N1215);
and AND2 (N1228, N1219, N791);
xor XOR2 (N1229, N1217, N548);
buf BUF1 (N1230, N1225);
buf BUF1 (N1231, N1228);
not NOT1 (N1232, N1206);
not NOT1 (N1233, N1223);
or OR3 (N1234, N1226, N614, N92);
xor XOR2 (N1235, N1233, N1068);
and AND3 (N1236, N1231, N14, N84);
xor XOR2 (N1237, N1222, N247);
or OR4 (N1238, N1234, N181, N814, N1125);
xor XOR2 (N1239, N1238, N421);
xor XOR2 (N1240, N1235, N511);
nor NOR4 (N1241, N1227, N528, N109, N557);
xor XOR2 (N1242, N1236, N1019);
buf BUF1 (N1243, N1221);
or OR4 (N1244, N1230, N1139, N1224, N733);
nand NAND2 (N1245, N1239, N126);
and AND4 (N1246, N1241, N307, N977, N1063);
buf BUF1 (N1247, N1244);
xor XOR2 (N1248, N1240, N1137);
xor XOR2 (N1249, N1245, N964);
and AND3 (N1250, N1232, N557, N908);
nor NOR4 (N1251, N1246, N464, N65, N67);
or OR2 (N1252, N1242, N134);
nand NAND2 (N1253, N1243, N171);
or OR4 (N1254, N1253, N1193, N355, N1223);
nor NOR3 (N1255, N1250, N69, N865);
not NOT1 (N1256, N1255);
and AND3 (N1257, N1254, N841, N159);
xor XOR2 (N1258, N1247, N213);
buf BUF1 (N1259, N1248);
not NOT1 (N1260, N1220);
or OR4 (N1261, N1251, N742, N998, N739);
or OR4 (N1262, N1261, N1230, N142, N448);
nand NAND4 (N1263, N1259, N460, N1067, N1125);
or OR2 (N1264, N1263, N900);
or OR3 (N1265, N1252, N155, N398);
buf BUF1 (N1266, N1249);
nand NAND4 (N1267, N1265, N440, N1102, N1080);
not NOT1 (N1268, N1260);
not NOT1 (N1269, N1257);
xor XOR2 (N1270, N1269, N164);
and AND2 (N1271, N1237, N864);
or OR2 (N1272, N1258, N1239);
not NOT1 (N1273, N1262);
buf BUF1 (N1274, N1270);
xor XOR2 (N1275, N1267, N780);
buf BUF1 (N1276, N1229);
buf BUF1 (N1277, N1256);
nor NOR4 (N1278, N1275, N512, N79, N431);
or OR2 (N1279, N1276, N1209);
or OR3 (N1280, N1264, N353, N112);
not NOT1 (N1281, N1278);
and AND2 (N1282, N1277, N56);
not NOT1 (N1283, N1274);
or OR4 (N1284, N1266, N1116, N323, N825);
xor XOR2 (N1285, N1279, N413);
nor NOR4 (N1286, N1282, N155, N593, N282);
or OR2 (N1287, N1283, N1141);
and AND4 (N1288, N1271, N841, N1235, N826);
or OR2 (N1289, N1287, N646);
buf BUF1 (N1290, N1289);
not NOT1 (N1291, N1290);
and AND2 (N1292, N1285, N551);
buf BUF1 (N1293, N1292);
nor NOR4 (N1294, N1284, N912, N199, N451);
or OR4 (N1295, N1268, N164, N412, N486);
buf BUF1 (N1296, N1281);
nor NOR2 (N1297, N1294, N312);
and AND2 (N1298, N1295, N1200);
buf BUF1 (N1299, N1298);
nand NAND4 (N1300, N1272, N894, N685, N1048);
and AND3 (N1301, N1293, N1142, N1143);
nor NOR2 (N1302, N1301, N398);
xor XOR2 (N1303, N1296, N1183);
buf BUF1 (N1304, N1302);
nand NAND4 (N1305, N1300, N898, N128, N1080);
and AND2 (N1306, N1299, N1153);
and AND2 (N1307, N1304, N382);
nand NAND4 (N1308, N1307, N163, N923, N484);
nor NOR2 (N1309, N1286, N136);
and AND3 (N1310, N1303, N92, N780);
nand NAND4 (N1311, N1308, N114, N481, N757);
and AND2 (N1312, N1309, N851);
and AND2 (N1313, N1311, N821);
nor NOR3 (N1314, N1305, N717, N481);
nand NAND2 (N1315, N1297, N654);
not NOT1 (N1316, N1280);
nand NAND3 (N1317, N1291, N459, N591);
xor XOR2 (N1318, N1314, N733);
and AND4 (N1319, N1288, N1291, N374, N1173);
or OR4 (N1320, N1315, N1107, N170, N396);
nor NOR3 (N1321, N1316, N664, N896);
and AND2 (N1322, N1317, N249);
or OR3 (N1323, N1321, N20, N123);
or OR4 (N1324, N1320, N730, N1263, N1162);
or OR3 (N1325, N1324, N833, N1287);
nand NAND4 (N1326, N1322, N236, N13, N820);
nand NAND2 (N1327, N1310, N1048);
xor XOR2 (N1328, N1318, N505);
and AND4 (N1329, N1312, N1303, N714, N713);
nor NOR3 (N1330, N1323, N1277, N489);
nor NOR4 (N1331, N1319, N1317, N132, N247);
or OR3 (N1332, N1329, N940, N869);
or OR4 (N1333, N1273, N1060, N223, N1227);
or OR2 (N1334, N1306, N1314);
or OR3 (N1335, N1327, N919, N1017);
buf BUF1 (N1336, N1335);
nand NAND3 (N1337, N1333, N1081, N1310);
buf BUF1 (N1338, N1325);
not NOT1 (N1339, N1313);
not NOT1 (N1340, N1328);
and AND2 (N1341, N1339, N19);
nand NAND3 (N1342, N1341, N474, N811);
or OR4 (N1343, N1331, N387, N1304, N659);
xor XOR2 (N1344, N1332, N1048);
nor NOR2 (N1345, N1344, N1121);
not NOT1 (N1346, N1338);
or OR4 (N1347, N1345, N137, N976, N809);
or OR4 (N1348, N1334, N1288, N782, N987);
buf BUF1 (N1349, N1326);
nor NOR4 (N1350, N1342, N1318, N803, N788);
buf BUF1 (N1351, N1347);
or OR2 (N1352, N1340, N887);
and AND3 (N1353, N1352, N651, N236);
or OR2 (N1354, N1346, N1243);
nor NOR2 (N1355, N1349, N178);
not NOT1 (N1356, N1354);
nand NAND4 (N1357, N1355, N801, N241, N116);
buf BUF1 (N1358, N1336);
and AND4 (N1359, N1353, N1182, N1356, N1159);
and AND4 (N1360, N432, N708, N1319, N1294);
nand NAND2 (N1361, N1360, N611);
buf BUF1 (N1362, N1358);
xor XOR2 (N1363, N1330, N515);
nor NOR2 (N1364, N1363, N243);
or OR3 (N1365, N1364, N495, N652);
xor XOR2 (N1366, N1357, N985);
nor NOR4 (N1367, N1343, N247, N568, N513);
buf BUF1 (N1368, N1362);
xor XOR2 (N1369, N1366, N879);
not NOT1 (N1370, N1361);
and AND3 (N1371, N1359, N902, N414);
not NOT1 (N1372, N1350);
not NOT1 (N1373, N1372);
not NOT1 (N1374, N1365);
nor NOR4 (N1375, N1348, N1157, N848, N376);
buf BUF1 (N1376, N1373);
xor XOR2 (N1377, N1374, N604);
not NOT1 (N1378, N1376);
nand NAND3 (N1379, N1375, N367, N1192);
not NOT1 (N1380, N1371);
not NOT1 (N1381, N1380);
xor XOR2 (N1382, N1367, N644);
and AND4 (N1383, N1370, N672, N1203, N86);
buf BUF1 (N1384, N1369);
nor NOR2 (N1385, N1381, N1130);
and AND3 (N1386, N1382, N151, N986);
xor XOR2 (N1387, N1368, N1037);
or OR2 (N1388, N1385, N1011);
xor XOR2 (N1389, N1351, N170);
xor XOR2 (N1390, N1379, N576);
or OR3 (N1391, N1378, N1036, N131);
or OR3 (N1392, N1383, N574, N715);
and AND4 (N1393, N1392, N1289, N739, N850);
nand NAND4 (N1394, N1389, N362, N820, N168);
nand NAND3 (N1395, N1377, N432, N309);
and AND3 (N1396, N1391, N105, N142);
and AND3 (N1397, N1337, N495, N942);
and AND3 (N1398, N1386, N725, N1326);
and AND3 (N1399, N1384, N483, N957);
nand NAND2 (N1400, N1390, N1180);
xor XOR2 (N1401, N1395, N1001);
not NOT1 (N1402, N1398);
nor NOR4 (N1403, N1402, N17, N593, N989);
nand NAND3 (N1404, N1403, N1322, N370);
buf BUF1 (N1405, N1393);
nand NAND2 (N1406, N1404, N1325);
nand NAND2 (N1407, N1387, N774);
nor NOR2 (N1408, N1388, N1301);
nand NAND3 (N1409, N1407, N1198, N1296);
not NOT1 (N1410, N1401);
or OR2 (N1411, N1409, N778);
nand NAND3 (N1412, N1405, N1198, N680);
nand NAND2 (N1413, N1400, N351);
nor NOR4 (N1414, N1406, N22, N933, N18);
nand NAND3 (N1415, N1399, N524, N1148);
nor NOR3 (N1416, N1412, N170, N5);
not NOT1 (N1417, N1410);
nor NOR2 (N1418, N1396, N26);
buf BUF1 (N1419, N1408);
xor XOR2 (N1420, N1415, N776);
buf BUF1 (N1421, N1397);
xor XOR2 (N1422, N1413, N1390);
not NOT1 (N1423, N1414);
nand NAND3 (N1424, N1421, N251, N1072);
not NOT1 (N1425, N1420);
nand NAND3 (N1426, N1417, N46, N1187);
xor XOR2 (N1427, N1394, N527);
buf BUF1 (N1428, N1416);
nand NAND3 (N1429, N1422, N1000, N255);
nor NOR3 (N1430, N1429, N1364, N968);
nand NAND4 (N1431, N1425, N622, N1134, N248);
and AND2 (N1432, N1418, N1276);
nor NOR3 (N1433, N1428, N460, N817);
nor NOR4 (N1434, N1430, N417, N839, N251);
buf BUF1 (N1435, N1423);
or OR3 (N1436, N1432, N235, N1120);
and AND3 (N1437, N1435, N945, N842);
nor NOR3 (N1438, N1437, N201, N52);
not NOT1 (N1439, N1434);
not NOT1 (N1440, N1419);
and AND4 (N1441, N1440, N998, N1167, N1357);
and AND3 (N1442, N1436, N392, N447);
or OR4 (N1443, N1427, N49, N451, N508);
nand NAND3 (N1444, N1411, N1396, N242);
not NOT1 (N1445, N1443);
or OR2 (N1446, N1431, N827);
buf BUF1 (N1447, N1433);
not NOT1 (N1448, N1439);
nand NAND4 (N1449, N1441, N1423, N1125, N928);
xor XOR2 (N1450, N1446, N1282);
nor NOR4 (N1451, N1445, N781, N482, N433);
nor NOR3 (N1452, N1448, N44, N1386);
and AND3 (N1453, N1449, N278, N370);
or OR2 (N1454, N1450, N1194);
not NOT1 (N1455, N1442);
xor XOR2 (N1456, N1424, N657);
nand NAND2 (N1457, N1452, N1041);
not NOT1 (N1458, N1444);
xor XOR2 (N1459, N1438, N1048);
buf BUF1 (N1460, N1458);
xor XOR2 (N1461, N1459, N114);
xor XOR2 (N1462, N1447, N355);
xor XOR2 (N1463, N1461, N823);
xor XOR2 (N1464, N1455, N1081);
xor XOR2 (N1465, N1456, N56);
buf BUF1 (N1466, N1426);
nor NOR2 (N1467, N1453, N868);
not NOT1 (N1468, N1467);
xor XOR2 (N1469, N1463, N1226);
buf BUF1 (N1470, N1466);
not NOT1 (N1471, N1451);
buf BUF1 (N1472, N1457);
not NOT1 (N1473, N1468);
or OR4 (N1474, N1469, N957, N996, N799);
buf BUF1 (N1475, N1462);
nor NOR3 (N1476, N1460, N272, N1410);
or OR2 (N1477, N1454, N579);
xor XOR2 (N1478, N1470, N137);
xor XOR2 (N1479, N1464, N882);
and AND2 (N1480, N1465, N1246);
xor XOR2 (N1481, N1474, N377);
or OR2 (N1482, N1472, N1167);
xor XOR2 (N1483, N1478, N598);
not NOT1 (N1484, N1482);
xor XOR2 (N1485, N1473, N394);
xor XOR2 (N1486, N1484, N244);
or OR2 (N1487, N1486, N70);
buf BUF1 (N1488, N1480);
nand NAND4 (N1489, N1487, N815, N1420, N1362);
not NOT1 (N1490, N1483);
nand NAND3 (N1491, N1489, N664, N234);
buf BUF1 (N1492, N1479);
buf BUF1 (N1493, N1475);
and AND4 (N1494, N1485, N920, N111, N72);
nand NAND2 (N1495, N1491, N49);
buf BUF1 (N1496, N1493);
and AND3 (N1497, N1492, N267, N14);
not NOT1 (N1498, N1495);
and AND2 (N1499, N1490, N106);
and AND4 (N1500, N1496, N984, N935, N1460);
not NOT1 (N1501, N1494);
buf BUF1 (N1502, N1471);
nand NAND3 (N1503, N1499, N121, N933);
or OR4 (N1504, N1497, N351, N123, N1340);
not NOT1 (N1505, N1476);
or OR4 (N1506, N1481, N1072, N869, N1379);
nand NAND2 (N1507, N1477, N460);
nor NOR2 (N1508, N1498, N293);
not NOT1 (N1509, N1508);
not NOT1 (N1510, N1507);
and AND2 (N1511, N1488, N126);
xor XOR2 (N1512, N1510, N957);
or OR3 (N1513, N1511, N219, N1407);
or OR3 (N1514, N1505, N142, N935);
and AND4 (N1515, N1504, N1378, N1025, N1091);
nor NOR4 (N1516, N1503, N1481, N832, N388);
nor NOR3 (N1517, N1512, N698, N1311);
nand NAND4 (N1518, N1500, N1501, N857, N1144);
not NOT1 (N1519, N1443);
nand NAND2 (N1520, N1519, N610);
or OR4 (N1521, N1518, N158, N835, N214);
nor NOR4 (N1522, N1514, N1416, N77, N902);
nand NAND2 (N1523, N1520, N607);
xor XOR2 (N1524, N1506, N1411);
nor NOR4 (N1525, N1523, N136, N729, N1191);
xor XOR2 (N1526, N1502, N551);
and AND3 (N1527, N1516, N195, N870);
xor XOR2 (N1528, N1521, N1306);
not NOT1 (N1529, N1527);
buf BUF1 (N1530, N1529);
buf BUF1 (N1531, N1525);
or OR2 (N1532, N1517, N821);
xor XOR2 (N1533, N1526, N649);
buf BUF1 (N1534, N1532);
nand NAND3 (N1535, N1509, N566, N1015);
nor NOR3 (N1536, N1530, N584, N1200);
or OR2 (N1537, N1533, N142);
or OR4 (N1538, N1536, N230, N889, N1334);
nand NAND3 (N1539, N1515, N422, N1051);
not NOT1 (N1540, N1538);
or OR3 (N1541, N1531, N437, N911);
and AND4 (N1542, N1534, N1170, N1003, N434);
nor NOR3 (N1543, N1524, N665, N1427);
not NOT1 (N1544, N1543);
buf BUF1 (N1545, N1544);
nor NOR4 (N1546, N1528, N272, N1500, N1013);
buf BUF1 (N1547, N1535);
nor NOR3 (N1548, N1537, N1066, N139);
and AND4 (N1549, N1547, N372, N822, N1175);
buf BUF1 (N1550, N1542);
or OR4 (N1551, N1539, N667, N1314, N1036);
nand NAND3 (N1552, N1513, N1143, N1163);
or OR3 (N1553, N1546, N1231, N1487);
and AND4 (N1554, N1551, N233, N439, N854);
and AND4 (N1555, N1552, N45, N1436, N7);
not NOT1 (N1556, N1522);
nor NOR4 (N1557, N1556, N1325, N1168, N34);
xor XOR2 (N1558, N1545, N1083);
and AND4 (N1559, N1550, N1325, N576, N343);
nor NOR3 (N1560, N1558, N290, N519);
or OR4 (N1561, N1548, N438, N567, N189);
nand NAND3 (N1562, N1554, N250, N859);
or OR3 (N1563, N1540, N541, N191);
xor XOR2 (N1564, N1555, N354);
xor XOR2 (N1565, N1563, N222);
or OR3 (N1566, N1549, N338, N355);
nor NOR3 (N1567, N1559, N1476, N146);
and AND4 (N1568, N1566, N329, N203, N432);
xor XOR2 (N1569, N1561, N60);
nor NOR2 (N1570, N1562, N1102);
and AND4 (N1571, N1553, N1020, N982, N1260);
buf BUF1 (N1572, N1568);
nand NAND2 (N1573, N1567, N888);
and AND2 (N1574, N1565, N200);
buf BUF1 (N1575, N1564);
nor NOR3 (N1576, N1560, N1437, N1240);
or OR4 (N1577, N1569, N661, N1353, N710);
and AND2 (N1578, N1570, N977);
nor NOR2 (N1579, N1571, N877);
not NOT1 (N1580, N1557);
nor NOR3 (N1581, N1576, N1031, N509);
nand NAND3 (N1582, N1580, N1031, N643);
nor NOR2 (N1583, N1581, N209);
not NOT1 (N1584, N1578);
not NOT1 (N1585, N1575);
nand NAND2 (N1586, N1583, N24);
nor NOR4 (N1587, N1541, N141, N1294, N1399);
or OR3 (N1588, N1587, N808, N305);
nand NAND3 (N1589, N1588, N1095, N222);
and AND2 (N1590, N1577, N717);
or OR3 (N1591, N1589, N893, N666);
nand NAND2 (N1592, N1590, N64);
nand NAND2 (N1593, N1586, N1314);
buf BUF1 (N1594, N1572);
nand NAND3 (N1595, N1585, N285, N51);
xor XOR2 (N1596, N1582, N25);
xor XOR2 (N1597, N1584, N1554);
nor NOR4 (N1598, N1591, N67, N264, N801);
nand NAND4 (N1599, N1573, N1035, N643, N587);
buf BUF1 (N1600, N1595);
buf BUF1 (N1601, N1600);
and AND2 (N1602, N1598, N1055);
not NOT1 (N1603, N1579);
nand NAND4 (N1604, N1596, N267, N1456, N197);
nor NOR4 (N1605, N1602, N177, N1159, N57);
xor XOR2 (N1606, N1593, N38);
xor XOR2 (N1607, N1597, N1354);
nor NOR3 (N1608, N1574, N1283, N1328);
and AND3 (N1609, N1607, N1509, N545);
buf BUF1 (N1610, N1606);
not NOT1 (N1611, N1594);
nand NAND3 (N1612, N1604, N1127, N183);
buf BUF1 (N1613, N1592);
not NOT1 (N1614, N1610);
not NOT1 (N1615, N1605);
not NOT1 (N1616, N1609);
nand NAND2 (N1617, N1611, N38);
nand NAND2 (N1618, N1613, N1071);
or OR2 (N1619, N1617, N1036);
nor NOR3 (N1620, N1615, N1514, N652);
nand NAND2 (N1621, N1608, N1525);
buf BUF1 (N1622, N1620);
and AND4 (N1623, N1622, N172, N1033, N1591);
xor XOR2 (N1624, N1603, N1031);
and AND4 (N1625, N1618, N1582, N136, N803);
nor NOR4 (N1626, N1601, N581, N214, N908);
or OR4 (N1627, N1616, N1338, N1118, N521);
nand NAND3 (N1628, N1627, N116, N125);
and AND4 (N1629, N1626, N1623, N312, N1265);
or OR2 (N1630, N842, N42);
not NOT1 (N1631, N1619);
buf BUF1 (N1632, N1621);
xor XOR2 (N1633, N1629, N1566);
nor NOR3 (N1634, N1630, N527, N1262);
nand NAND4 (N1635, N1625, N768, N717, N314);
not NOT1 (N1636, N1632);
xor XOR2 (N1637, N1631, N994);
nor NOR3 (N1638, N1633, N1357, N526);
not NOT1 (N1639, N1634);
buf BUF1 (N1640, N1637);
buf BUF1 (N1641, N1624);
nand NAND4 (N1642, N1641, N1475, N1131, N1596);
xor XOR2 (N1643, N1628, N306);
nor NOR3 (N1644, N1639, N580, N133);
nor NOR2 (N1645, N1599, N757);
xor XOR2 (N1646, N1644, N438);
or OR2 (N1647, N1640, N1322);
nor NOR4 (N1648, N1614, N520, N955, N532);
nand NAND3 (N1649, N1636, N1479, N458);
and AND4 (N1650, N1649, N1173, N759, N149);
not NOT1 (N1651, N1650);
or OR3 (N1652, N1643, N833, N1276);
nor NOR3 (N1653, N1648, N700, N1008);
buf BUF1 (N1654, N1646);
or OR4 (N1655, N1652, N1457, N380, N212);
or OR4 (N1656, N1647, N545, N581, N37);
and AND4 (N1657, N1638, N1086, N472, N475);
nand NAND3 (N1658, N1655, N300, N245);
and AND4 (N1659, N1642, N1357, N764, N923);
xor XOR2 (N1660, N1657, N1555);
or OR3 (N1661, N1654, N1335, N322);
and AND4 (N1662, N1612, N8, N92, N144);
buf BUF1 (N1663, N1660);
not NOT1 (N1664, N1635);
nand NAND2 (N1665, N1658, N192);
and AND4 (N1666, N1651, N491, N1606, N445);
nor NOR3 (N1667, N1665, N614, N513);
not NOT1 (N1668, N1653);
buf BUF1 (N1669, N1666);
or OR2 (N1670, N1645, N1456);
xor XOR2 (N1671, N1656, N279);
and AND4 (N1672, N1663, N1101, N1613, N1301);
buf BUF1 (N1673, N1669);
not NOT1 (N1674, N1671);
and AND2 (N1675, N1661, N1271);
xor XOR2 (N1676, N1674, N261);
nand NAND4 (N1677, N1675, N569, N113, N790);
nand NAND3 (N1678, N1672, N44, N693);
nand NAND4 (N1679, N1677, N1677, N335, N224);
xor XOR2 (N1680, N1668, N371);
nand NAND3 (N1681, N1678, N1203, N1248);
or OR2 (N1682, N1659, N767);
buf BUF1 (N1683, N1670);
nor NOR4 (N1684, N1680, N1237, N102, N112);
xor XOR2 (N1685, N1676, N1500);
or OR2 (N1686, N1684, N1046);
nand NAND4 (N1687, N1679, N1194, N140, N815);
nand NAND2 (N1688, N1682, N1357);
not NOT1 (N1689, N1662);
and AND4 (N1690, N1667, N293, N1379, N383);
nand NAND2 (N1691, N1690, N68);
nor NOR2 (N1692, N1689, N1682);
nor NOR3 (N1693, N1691, N218, N602);
nor NOR2 (N1694, N1693, N1666);
nand NAND3 (N1695, N1683, N736, N350);
nor NOR3 (N1696, N1692, N849, N1154);
not NOT1 (N1697, N1673);
and AND4 (N1698, N1686, N1520, N1143, N808);
nand NAND3 (N1699, N1694, N410, N227);
xor XOR2 (N1700, N1688, N1479);
not NOT1 (N1701, N1687);
not NOT1 (N1702, N1695);
xor XOR2 (N1703, N1698, N794);
not NOT1 (N1704, N1703);
nand NAND4 (N1705, N1704, N1245, N1270, N321);
buf BUF1 (N1706, N1702);
and AND3 (N1707, N1681, N140, N1457);
nor NOR4 (N1708, N1707, N788, N1035, N453);
xor XOR2 (N1709, N1701, N519);
and AND2 (N1710, N1705, N1672);
and AND4 (N1711, N1708, N620, N945, N354);
or OR3 (N1712, N1685, N58, N1054);
nor NOR2 (N1713, N1697, N857);
buf BUF1 (N1714, N1706);
not NOT1 (N1715, N1664);
nor NOR4 (N1716, N1709, N1315, N1068, N308);
or OR3 (N1717, N1716, N368, N102);
nor NOR3 (N1718, N1710, N741, N902);
xor XOR2 (N1719, N1713, N1463);
buf BUF1 (N1720, N1715);
xor XOR2 (N1721, N1696, N159);
or OR3 (N1722, N1719, N690, N456);
buf BUF1 (N1723, N1718);
buf BUF1 (N1724, N1711);
buf BUF1 (N1725, N1712);
nand NAND3 (N1726, N1721, N1072, N1196);
nor NOR4 (N1727, N1725, N500, N1224, N630);
and AND4 (N1728, N1727, N1433, N924, N1269);
or OR2 (N1729, N1700, N330);
not NOT1 (N1730, N1717);
not NOT1 (N1731, N1728);
xor XOR2 (N1732, N1730, N818);
nand NAND2 (N1733, N1729, N1350);
and AND2 (N1734, N1699, N432);
buf BUF1 (N1735, N1732);
not NOT1 (N1736, N1731);
not NOT1 (N1737, N1720);
and AND3 (N1738, N1736, N391, N772);
buf BUF1 (N1739, N1722);
nand NAND4 (N1740, N1726, N1033, N32, N1601);
and AND2 (N1741, N1734, N252);
nand NAND3 (N1742, N1738, N1454, N1610);
buf BUF1 (N1743, N1741);
and AND3 (N1744, N1735, N1708, N834);
buf BUF1 (N1745, N1740);
not NOT1 (N1746, N1737);
nor NOR3 (N1747, N1745, N874, N665);
xor XOR2 (N1748, N1744, N1534);
buf BUF1 (N1749, N1746);
xor XOR2 (N1750, N1724, N1090);
xor XOR2 (N1751, N1733, N1710);
not NOT1 (N1752, N1742);
not NOT1 (N1753, N1714);
buf BUF1 (N1754, N1723);
nor NOR2 (N1755, N1753, N1492);
nand NAND2 (N1756, N1751, N1681);
xor XOR2 (N1757, N1748, N119);
and AND3 (N1758, N1743, N76, N1381);
nor NOR2 (N1759, N1750, N37);
and AND2 (N1760, N1747, N797);
buf BUF1 (N1761, N1749);
and AND4 (N1762, N1757, N71, N428, N760);
not NOT1 (N1763, N1739);
xor XOR2 (N1764, N1756, N1450);
nand NAND4 (N1765, N1764, N159, N1152, N945);
xor XOR2 (N1766, N1762, N371);
or OR4 (N1767, N1755, N109, N989, N1017);
buf BUF1 (N1768, N1760);
not NOT1 (N1769, N1754);
xor XOR2 (N1770, N1758, N443);
buf BUF1 (N1771, N1765);
xor XOR2 (N1772, N1763, N44);
xor XOR2 (N1773, N1759, N125);
xor XOR2 (N1774, N1761, N379);
xor XOR2 (N1775, N1766, N584);
xor XOR2 (N1776, N1772, N330);
buf BUF1 (N1777, N1770);
or OR2 (N1778, N1777, N1559);
buf BUF1 (N1779, N1752);
buf BUF1 (N1780, N1775);
xor XOR2 (N1781, N1767, N1308);
and AND4 (N1782, N1776, N1440, N739, N982);
xor XOR2 (N1783, N1779, N1035);
or OR3 (N1784, N1774, N550, N845);
nor NOR4 (N1785, N1768, N867, N1776, N42);
nor NOR3 (N1786, N1785, N39, N1301);
xor XOR2 (N1787, N1778, N1328);
or OR2 (N1788, N1787, N1024);
and AND3 (N1789, N1784, N1293, N1560);
nor NOR2 (N1790, N1781, N1240);
buf BUF1 (N1791, N1769);
nand NAND3 (N1792, N1788, N1210, N1375);
nand NAND3 (N1793, N1791, N261, N157);
not NOT1 (N1794, N1792);
and AND4 (N1795, N1793, N979, N12, N588);
xor XOR2 (N1796, N1795, N161);
nor NOR2 (N1797, N1783, N487);
or OR3 (N1798, N1789, N231, N1539);
or OR4 (N1799, N1773, N353, N1181, N1409);
and AND4 (N1800, N1798, N914, N35, N115);
or OR2 (N1801, N1800, N821);
and AND4 (N1802, N1794, N1311, N1639, N51);
nand NAND4 (N1803, N1771, N1086, N151, N1801);
not NOT1 (N1804, N489);
nand NAND4 (N1805, N1796, N303, N707, N240);
or OR2 (N1806, N1802, N596);
xor XOR2 (N1807, N1797, N340);
xor XOR2 (N1808, N1799, N1633);
or OR4 (N1809, N1780, N134, N559, N777);
or OR2 (N1810, N1790, N1388);
xor XOR2 (N1811, N1786, N242);
or OR3 (N1812, N1807, N3, N196);
xor XOR2 (N1813, N1803, N709);
and AND4 (N1814, N1813, N936, N1049, N367);
not NOT1 (N1815, N1804);
xor XOR2 (N1816, N1808, N1434);
or OR4 (N1817, N1806, N1285, N1444, N928);
nor NOR3 (N1818, N1810, N621, N1171);
buf BUF1 (N1819, N1809);
xor XOR2 (N1820, N1782, N1362);
or OR3 (N1821, N1805, N1507, N1564);
or OR3 (N1822, N1816, N724, N1550);
buf BUF1 (N1823, N1821);
not NOT1 (N1824, N1822);
and AND2 (N1825, N1812, N1173);
buf BUF1 (N1826, N1820);
nor NOR4 (N1827, N1817, N460, N1033, N1717);
nand NAND2 (N1828, N1815, N1089);
or OR3 (N1829, N1828, N1233, N234);
and AND3 (N1830, N1824, N668, N1764);
xor XOR2 (N1831, N1823, N144);
or OR4 (N1832, N1830, N1543, N661, N364);
nor NOR2 (N1833, N1827, N1033);
nor NOR2 (N1834, N1811, N928);
nor NOR4 (N1835, N1832, N476, N404, N617);
nor NOR4 (N1836, N1814, N1691, N1563, N1432);
nor NOR2 (N1837, N1833, N1562);
and AND2 (N1838, N1837, N916);
xor XOR2 (N1839, N1818, N731);
not NOT1 (N1840, N1839);
buf BUF1 (N1841, N1826);
nor NOR4 (N1842, N1836, N689, N1537, N1078);
xor XOR2 (N1843, N1825, N1166);
nand NAND2 (N1844, N1840, N488);
buf BUF1 (N1845, N1843);
and AND4 (N1846, N1841, N21, N305, N436);
nand NAND2 (N1847, N1831, N721);
and AND3 (N1848, N1844, N836, N733);
or OR3 (N1849, N1847, N87, N1557);
xor XOR2 (N1850, N1835, N823);
xor XOR2 (N1851, N1846, N36);
not NOT1 (N1852, N1838);
and AND2 (N1853, N1834, N23);
nor NOR2 (N1854, N1852, N1780);
xor XOR2 (N1855, N1850, N894);
buf BUF1 (N1856, N1855);
nor NOR3 (N1857, N1845, N226, N710);
buf BUF1 (N1858, N1819);
or OR3 (N1859, N1842, N1831, N707);
or OR2 (N1860, N1829, N1545);
xor XOR2 (N1861, N1851, N1411);
buf BUF1 (N1862, N1858);
and AND4 (N1863, N1848, N1591, N1210, N424);
and AND4 (N1864, N1856, N668, N262, N471);
and AND2 (N1865, N1860, N130);
nor NOR4 (N1866, N1863, N1212, N901, N1820);
not NOT1 (N1867, N1859);
nand NAND2 (N1868, N1861, N154);
xor XOR2 (N1869, N1849, N407);
nand NAND3 (N1870, N1864, N580, N542);
buf BUF1 (N1871, N1857);
and AND2 (N1872, N1866, N1041);
and AND4 (N1873, N1871, N859, N782, N180);
and AND3 (N1874, N1862, N15, N1335);
nand NAND2 (N1875, N1865, N996);
not NOT1 (N1876, N1868);
and AND4 (N1877, N1867, N182, N48, N103);
or OR3 (N1878, N1854, N206, N1190);
not NOT1 (N1879, N1875);
or OR2 (N1880, N1872, N525);
or OR4 (N1881, N1874, N1140, N224, N850);
xor XOR2 (N1882, N1877, N512);
nor NOR3 (N1883, N1880, N654, N72);
buf BUF1 (N1884, N1869);
or OR4 (N1885, N1882, N1132, N267, N263);
and AND3 (N1886, N1878, N568, N1031);
nor NOR3 (N1887, N1853, N1134, N331);
xor XOR2 (N1888, N1884, N1241);
xor XOR2 (N1889, N1876, N875);
xor XOR2 (N1890, N1881, N1676);
and AND3 (N1891, N1885, N805, N952);
nor NOR3 (N1892, N1879, N382, N220);
or OR4 (N1893, N1890, N421, N808, N1042);
not NOT1 (N1894, N1888);
xor XOR2 (N1895, N1873, N592);
not NOT1 (N1896, N1889);
not NOT1 (N1897, N1893);
not NOT1 (N1898, N1887);
or OR2 (N1899, N1896, N590);
or OR3 (N1900, N1895, N1844, N430);
nor NOR3 (N1901, N1883, N1763, N1684);
and AND3 (N1902, N1870, N1427, N96);
xor XOR2 (N1903, N1897, N1377);
and AND3 (N1904, N1902, N372, N1820);
nor NOR4 (N1905, N1898, N667, N1071, N1677);
nor NOR3 (N1906, N1901, N1458, N1833);
buf BUF1 (N1907, N1906);
nand NAND2 (N1908, N1905, N812);
nand NAND4 (N1909, N1904, N454, N1576, N1846);
xor XOR2 (N1910, N1899, N102);
not NOT1 (N1911, N1891);
and AND4 (N1912, N1903, N867, N1522, N932);
not NOT1 (N1913, N1894);
nor NOR2 (N1914, N1910, N1546);
or OR3 (N1915, N1886, N368, N1891);
nand NAND4 (N1916, N1909, N1440, N885, N565);
xor XOR2 (N1917, N1913, N1795);
nor NOR3 (N1918, N1915, N1660, N1126);
nor NOR4 (N1919, N1907, N508, N61, N1634);
and AND2 (N1920, N1911, N875);
xor XOR2 (N1921, N1892, N1120);
buf BUF1 (N1922, N1908);
or OR2 (N1923, N1900, N1716);
nor NOR3 (N1924, N1919, N1405, N736);
buf BUF1 (N1925, N1918);
nor NOR3 (N1926, N1920, N1851, N1240);
not NOT1 (N1927, N1923);
not NOT1 (N1928, N1916);
xor XOR2 (N1929, N1914, N997);
buf BUF1 (N1930, N1924);
nor NOR2 (N1931, N1927, N133);
buf BUF1 (N1932, N1925);
nor NOR2 (N1933, N1922, N450);
xor XOR2 (N1934, N1930, N1257);
nor NOR2 (N1935, N1934, N1059);
buf BUF1 (N1936, N1933);
nand NAND4 (N1937, N1931, N1830, N470, N1139);
or OR4 (N1938, N1921, N1908, N671, N134);
and AND3 (N1939, N1932, N246, N575);
and AND4 (N1940, N1936, N605, N1890, N708);
and AND3 (N1941, N1929, N686, N1093);
nand NAND4 (N1942, N1939, N177, N1837, N1819);
not NOT1 (N1943, N1937);
and AND3 (N1944, N1917, N1640, N1800);
nor NOR2 (N1945, N1928, N678);
buf BUF1 (N1946, N1926);
and AND3 (N1947, N1945, N1477, N1252);
and AND3 (N1948, N1947, N159, N1342);
and AND3 (N1949, N1948, N1338, N1889);
and AND2 (N1950, N1949, N125);
nor NOR4 (N1951, N1941, N952, N1909, N1530);
nor NOR4 (N1952, N1942, N230, N1624, N760);
buf BUF1 (N1953, N1950);
xor XOR2 (N1954, N1938, N649);
nand NAND4 (N1955, N1935, N1099, N911, N563);
not NOT1 (N1956, N1940);
nand NAND4 (N1957, N1954, N707, N308, N105);
or OR3 (N1958, N1944, N1952, N96);
xor XOR2 (N1959, N509, N357);
buf BUF1 (N1960, N1946);
nand NAND3 (N1961, N1912, N119, N1773);
xor XOR2 (N1962, N1959, N841);
xor XOR2 (N1963, N1943, N400);
or OR2 (N1964, N1953, N268);
xor XOR2 (N1965, N1955, N1672);
nor NOR2 (N1966, N1961, N1015);
and AND2 (N1967, N1965, N228);
nand NAND3 (N1968, N1957, N1558, N1533);
or OR2 (N1969, N1964, N1537);
nand NAND4 (N1970, N1969, N668, N873, N1195);
nand NAND3 (N1971, N1960, N1486, N262);
not NOT1 (N1972, N1951);
not NOT1 (N1973, N1966);
nand NAND2 (N1974, N1968, N1514);
not NOT1 (N1975, N1972);
not NOT1 (N1976, N1971);
buf BUF1 (N1977, N1973);
nand NAND2 (N1978, N1963, N157);
and AND2 (N1979, N1962, N930);
xor XOR2 (N1980, N1974, N1315);
not NOT1 (N1981, N1980);
or OR2 (N1982, N1956, N1533);
not NOT1 (N1983, N1975);
nor NOR3 (N1984, N1979, N306, N1967);
not NOT1 (N1985, N1041);
and AND2 (N1986, N1985, N1746);
not NOT1 (N1987, N1981);
xor XOR2 (N1988, N1958, N440);
not NOT1 (N1989, N1978);
buf BUF1 (N1990, N1989);
xor XOR2 (N1991, N1988, N210);
and AND2 (N1992, N1987, N1239);
nand NAND3 (N1993, N1984, N993, N90);
xor XOR2 (N1994, N1991, N84);
nor NOR4 (N1995, N1976, N490, N1354, N299);
and AND3 (N1996, N1977, N581, N1123);
and AND4 (N1997, N1996, N923, N1707, N732);
buf BUF1 (N1998, N1997);
nand NAND4 (N1999, N1998, N214, N1794, N1996);
and AND4 (N2000, N1990, N164, N1557, N758);
xor XOR2 (N2001, N1986, N1015);
buf BUF1 (N2002, N1970);
xor XOR2 (N2003, N2002, N1969);
or OR3 (N2004, N1982, N1813, N623);
nor NOR3 (N2005, N2004, N1643, N219);
not NOT1 (N2006, N1993);
or OR3 (N2007, N1994, N1068, N92);
nor NOR2 (N2008, N1983, N758);
not NOT1 (N2009, N2006);
nand NAND3 (N2010, N2001, N1274, N1826);
xor XOR2 (N2011, N2005, N1617);
and AND2 (N2012, N2009, N415);
nor NOR2 (N2013, N1992, N1345);
buf BUF1 (N2014, N2012);
nor NOR3 (N2015, N2011, N177, N1184);
and AND3 (N2016, N2015, N1222, N85);
buf BUF1 (N2017, N2014);
nand NAND3 (N2018, N2013, N1007, N399);
buf BUF1 (N2019, N2010);
not NOT1 (N2020, N2007);
not NOT1 (N2021, N2018);
not NOT1 (N2022, N2019);
nor NOR2 (N2023, N2003, N879);
not NOT1 (N2024, N2016);
xor XOR2 (N2025, N2023, N1887);
nor NOR3 (N2026, N2020, N1656, N1801);
nand NAND2 (N2027, N1999, N32);
buf BUF1 (N2028, N2021);
not NOT1 (N2029, N2027);
and AND4 (N2030, N2008, N1560, N709, N1900);
xor XOR2 (N2031, N1995, N574);
nor NOR3 (N2032, N2029, N891, N1692);
nor NOR3 (N2033, N2017, N1507, N1603);
xor XOR2 (N2034, N2033, N1036);
or OR2 (N2035, N2028, N1766);
nor NOR2 (N2036, N2030, N1795);
xor XOR2 (N2037, N2022, N937);
or OR2 (N2038, N2031, N1814);
buf BUF1 (N2039, N2026);
buf BUF1 (N2040, N2039);
nor NOR3 (N2041, N2040, N1161, N1942);
not NOT1 (N2042, N2041);
or OR2 (N2043, N2036, N324);
nand NAND4 (N2044, N2038, N823, N1841, N1391);
not NOT1 (N2045, N2024);
buf BUF1 (N2046, N2000);
and AND3 (N2047, N2037, N8, N780);
xor XOR2 (N2048, N2043, N1759);
or OR2 (N2049, N2047, N322);
nand NAND3 (N2050, N2034, N695, N1513);
nand NAND3 (N2051, N2042, N921, N1549);
buf BUF1 (N2052, N2048);
nor NOR4 (N2053, N2044, N1113, N1733, N287);
or OR4 (N2054, N2035, N1214, N343, N1567);
not NOT1 (N2055, N2050);
nand NAND2 (N2056, N2046, N149);
and AND4 (N2057, N2032, N1120, N675, N890);
nor NOR2 (N2058, N2056, N1586);
nor NOR4 (N2059, N2049, N1662, N1581, N803);
nor NOR2 (N2060, N2058, N1924);
buf BUF1 (N2061, N2052);
nand NAND3 (N2062, N2051, N1029, N1892);
or OR2 (N2063, N2045, N112);
nor NOR3 (N2064, N2053, N588, N1733);
not NOT1 (N2065, N2057);
buf BUF1 (N2066, N2061);
or OR3 (N2067, N2054, N125, N40);
buf BUF1 (N2068, N2065);
nor NOR3 (N2069, N2059, N329, N235);
buf BUF1 (N2070, N2060);
buf BUF1 (N2071, N2068);
or OR2 (N2072, N2062, N1576);
nor NOR3 (N2073, N2064, N1466, N156);
not NOT1 (N2074, N2072);
nand NAND3 (N2075, N2073, N555, N586);
and AND4 (N2076, N2071, N122, N415, N1366);
buf BUF1 (N2077, N2067);
nand NAND3 (N2078, N2063, N1471, N300);
not NOT1 (N2079, N2025);
not NOT1 (N2080, N2076);
nand NAND3 (N2081, N2077, N133, N1371);
and AND3 (N2082, N2075, N1670, N1282);
xor XOR2 (N2083, N2069, N961);
nor NOR2 (N2084, N2066, N1280);
xor XOR2 (N2085, N2074, N1291);
buf BUF1 (N2086, N2080);
xor XOR2 (N2087, N2081, N85);
not NOT1 (N2088, N2055);
or OR3 (N2089, N2087, N386, N493);
not NOT1 (N2090, N2079);
not NOT1 (N2091, N2070);
nand NAND2 (N2092, N2090, N1116);
and AND4 (N2093, N2084, N1642, N1656, N2070);
nor NOR2 (N2094, N2089, N918);
and AND2 (N2095, N2093, N1887);
xor XOR2 (N2096, N2083, N1410);
buf BUF1 (N2097, N2095);
not NOT1 (N2098, N2097);
buf BUF1 (N2099, N2092);
buf BUF1 (N2100, N2094);
nand NAND2 (N2101, N2100, N909);
not NOT1 (N2102, N2085);
and AND3 (N2103, N2086, N1365, N352);
not NOT1 (N2104, N2101);
nand NAND3 (N2105, N2078, N746, N1080);
and AND2 (N2106, N2103, N1741);
buf BUF1 (N2107, N2106);
not NOT1 (N2108, N2105);
or OR4 (N2109, N2102, N1054, N474, N1851);
nand NAND4 (N2110, N2091, N178, N1636, N204);
or OR4 (N2111, N2108, N978, N392, N75);
or OR4 (N2112, N2088, N416, N1520, N88);
buf BUF1 (N2113, N2104);
not NOT1 (N2114, N2111);
or OR4 (N2115, N2099, N812, N1985, N1575);
xor XOR2 (N2116, N2112, N1557);
xor XOR2 (N2117, N2110, N1246);
buf BUF1 (N2118, N2096);
or OR4 (N2119, N2114, N1591, N227, N1512);
not NOT1 (N2120, N2109);
or OR3 (N2121, N2118, N1793, N2113);
or OR2 (N2122, N451, N1709);
xor XOR2 (N2123, N2122, N2102);
nor NOR2 (N2124, N2098, N201);
nand NAND3 (N2125, N2117, N435, N31);
not NOT1 (N2126, N2124);
nor NOR3 (N2127, N2125, N1214, N1164);
or OR2 (N2128, N2107, N796);
and AND4 (N2129, N2116, N122, N1759, N2059);
xor XOR2 (N2130, N2127, N2052);
buf BUF1 (N2131, N2130);
and AND2 (N2132, N2128, N503);
not NOT1 (N2133, N2120);
nand NAND2 (N2134, N2133, N1250);
nand NAND2 (N2135, N2082, N748);
nor NOR2 (N2136, N2123, N913);
xor XOR2 (N2137, N2115, N418);
not NOT1 (N2138, N2126);
nand NAND4 (N2139, N2121, N1635, N58, N455);
not NOT1 (N2140, N2138);
nand NAND4 (N2141, N2132, N185, N899, N1086);
and AND2 (N2142, N2139, N306);
buf BUF1 (N2143, N2129);
xor XOR2 (N2144, N2142, N555);
buf BUF1 (N2145, N2135);
or OR3 (N2146, N2134, N708, N1693);
xor XOR2 (N2147, N2136, N1010);
nand NAND4 (N2148, N2146, N861, N1680, N1091);
buf BUF1 (N2149, N2143);
xor XOR2 (N2150, N2137, N2014);
or OR2 (N2151, N2150, N113);
or OR2 (N2152, N2119, N36);
nand NAND3 (N2153, N2131, N1810, N1691);
nor NOR2 (N2154, N2144, N344);
or OR2 (N2155, N2149, N1101);
and AND2 (N2156, N2151, N1338);
nor NOR2 (N2157, N2153, N83);
nor NOR4 (N2158, N2140, N1341, N698, N843);
nor NOR3 (N2159, N2158, N1312, N1366);
xor XOR2 (N2160, N2154, N702);
or OR3 (N2161, N2145, N247, N314);
nor NOR3 (N2162, N2161, N1504, N1350);
not NOT1 (N2163, N2155);
xor XOR2 (N2164, N2152, N1104);
buf BUF1 (N2165, N2163);
not NOT1 (N2166, N2148);
not NOT1 (N2167, N2159);
or OR4 (N2168, N2147, N1582, N1592, N1817);
nand NAND2 (N2169, N2160, N2024);
nand NAND2 (N2170, N2165, N440);
not NOT1 (N2171, N2141);
or OR3 (N2172, N2168, N22, N1560);
buf BUF1 (N2173, N2162);
xor XOR2 (N2174, N2173, N16);
buf BUF1 (N2175, N2167);
and AND3 (N2176, N2164, N272, N1374);
and AND4 (N2177, N2174, N758, N1268, N1166);
and AND4 (N2178, N2176, N1272, N1340, N163);
or OR4 (N2179, N2172, N1036, N625, N861);
xor XOR2 (N2180, N2175, N73);
buf BUF1 (N2181, N2180);
and AND2 (N2182, N2177, N1790);
or OR3 (N2183, N2157, N2030, N210);
not NOT1 (N2184, N2178);
and AND3 (N2185, N2181, N1702, N2008);
and AND2 (N2186, N2169, N907);
or OR4 (N2187, N2184, N1813, N1266, N438);
buf BUF1 (N2188, N2171);
nand NAND4 (N2189, N2156, N1505, N1496, N329);
buf BUF1 (N2190, N2188);
and AND4 (N2191, N2190, N1783, N166, N2141);
or OR3 (N2192, N2185, N1329, N984);
and AND3 (N2193, N2186, N852, N174);
xor XOR2 (N2194, N2193, N1131);
or OR4 (N2195, N2179, N764, N2080, N1343);
and AND4 (N2196, N2183, N1487, N263, N1371);
or OR2 (N2197, N2196, N2063);
nor NOR4 (N2198, N2192, N718, N781, N1593);
and AND3 (N2199, N2191, N343, N1867);
and AND3 (N2200, N2197, N1840, N283);
nand NAND4 (N2201, N2198, N933, N2121, N962);
nor NOR3 (N2202, N2166, N57, N1557);
xor XOR2 (N2203, N2195, N870);
nand NAND2 (N2204, N2199, N987);
buf BUF1 (N2205, N2202);
not NOT1 (N2206, N2189);
nor NOR2 (N2207, N2204, N1645);
and AND2 (N2208, N2200, N887);
xor XOR2 (N2209, N2208, N336);
nor NOR2 (N2210, N2206, N1382);
buf BUF1 (N2211, N2170);
nand NAND2 (N2212, N2194, N1088);
or OR2 (N2213, N2205, N1608);
and AND3 (N2214, N2207, N173, N848);
or OR3 (N2215, N2209, N822, N756);
nor NOR2 (N2216, N2182, N1289);
not NOT1 (N2217, N2201);
buf BUF1 (N2218, N2211);
or OR3 (N2219, N2213, N456, N513);
or OR4 (N2220, N2210, N1124, N322, N2161);
nor NOR3 (N2221, N2219, N2218, N1995);
not NOT1 (N2222, N1331);
nand NAND4 (N2223, N2187, N1497, N1106, N517);
not NOT1 (N2224, N2212);
not NOT1 (N2225, N2217);
buf BUF1 (N2226, N2222);
nor NOR3 (N2227, N2215, N1961, N551);
or OR2 (N2228, N2224, N766);
nand NAND2 (N2229, N2226, N55);
buf BUF1 (N2230, N2228);
or OR3 (N2231, N2223, N131, N930);
and AND4 (N2232, N2221, N639, N933, N2027);
or OR3 (N2233, N2230, N589, N1502);
and AND4 (N2234, N2233, N1324, N713, N687);
buf BUF1 (N2235, N2220);
or OR3 (N2236, N2229, N1476, N2193);
and AND3 (N2237, N2231, N1906, N1131);
xor XOR2 (N2238, N2214, N885);
nand NAND3 (N2239, N2227, N854, N1688);
nor NOR3 (N2240, N2232, N687, N1106);
buf BUF1 (N2241, N2225);
buf BUF1 (N2242, N2241);
nand NAND3 (N2243, N2242, N461, N1504);
not NOT1 (N2244, N2238);
buf BUF1 (N2245, N2234);
xor XOR2 (N2246, N2244, N859);
xor XOR2 (N2247, N2235, N592);
xor XOR2 (N2248, N2245, N945);
nand NAND3 (N2249, N2216, N574, N2122);
not NOT1 (N2250, N2203);
not NOT1 (N2251, N2239);
nand NAND4 (N2252, N2247, N1002, N549, N2202);
and AND3 (N2253, N2243, N217, N2014);
not NOT1 (N2254, N2251);
nand NAND4 (N2255, N2253, N586, N31, N1711);
or OR4 (N2256, N2246, N1709, N349, N956);
and AND2 (N2257, N2252, N1260);
or OR4 (N2258, N2256, N1880, N661, N439);
xor XOR2 (N2259, N2257, N1026);
not NOT1 (N2260, N2240);
buf BUF1 (N2261, N2250);
not NOT1 (N2262, N2258);
buf BUF1 (N2263, N2259);
not NOT1 (N2264, N2262);
and AND2 (N2265, N2261, N1741);
buf BUF1 (N2266, N2264);
not NOT1 (N2267, N2260);
not NOT1 (N2268, N2249);
or OR3 (N2269, N2255, N898, N927);
and AND3 (N2270, N2263, N1281, N1346);
and AND3 (N2271, N2270, N530, N102);
not NOT1 (N2272, N2248);
buf BUF1 (N2273, N2267);
or OR4 (N2274, N2266, N894, N1211, N1103);
buf BUF1 (N2275, N2271);
xor XOR2 (N2276, N2268, N1678);
buf BUF1 (N2277, N2269);
or OR2 (N2278, N2277, N1290);
nor NOR4 (N2279, N2275, N1519, N34, N1855);
buf BUF1 (N2280, N2265);
or OR4 (N2281, N2278, N1725, N718, N677);
xor XOR2 (N2282, N2280, N578);
and AND2 (N2283, N2279, N1757);
not NOT1 (N2284, N2283);
nand NAND3 (N2285, N2282, N2249, N2119);
nand NAND3 (N2286, N2237, N1184, N2265);
nand NAND2 (N2287, N2281, N141);
nand NAND2 (N2288, N2254, N1400);
and AND2 (N2289, N2273, N661);
and AND3 (N2290, N2287, N237, N625);
nor NOR3 (N2291, N2276, N1339, N271);
not NOT1 (N2292, N2284);
or OR3 (N2293, N2274, N2023, N224);
not NOT1 (N2294, N2289);
not NOT1 (N2295, N2290);
xor XOR2 (N2296, N2236, N699);
not NOT1 (N2297, N2294);
or OR3 (N2298, N2288, N299, N231);
buf BUF1 (N2299, N2295);
and AND3 (N2300, N2286, N1538, N1688);
nand NAND2 (N2301, N2293, N1234);
not NOT1 (N2302, N2297);
nand NAND2 (N2303, N2300, N1095);
nand NAND2 (N2304, N2301, N2198);
nand NAND2 (N2305, N2304, N1875);
and AND4 (N2306, N2298, N1977, N2224, N258);
nor NOR4 (N2307, N2306, N180, N1292, N406);
and AND3 (N2308, N2303, N535, N2198);
buf BUF1 (N2309, N2292);
and AND4 (N2310, N2307, N1716, N53, N1398);
nand NAND4 (N2311, N2305, N1007, N721, N1297);
nand NAND2 (N2312, N2291, N959);
nor NOR2 (N2313, N2310, N760);
buf BUF1 (N2314, N2309);
xor XOR2 (N2315, N2272, N2091);
nand NAND2 (N2316, N2302, N1933);
and AND4 (N2317, N2299, N1142, N551, N611);
nor NOR3 (N2318, N2285, N962, N2199);
nand NAND4 (N2319, N2308, N54, N1502, N2087);
not NOT1 (N2320, N2312);
buf BUF1 (N2321, N2314);
nor NOR4 (N2322, N2319, N687, N1312, N1501);
or OR2 (N2323, N2315, N965);
nand NAND4 (N2324, N2320, N1691, N1951, N1523);
or OR2 (N2325, N2321, N788);
buf BUF1 (N2326, N2318);
not NOT1 (N2327, N2313);
nor NOR3 (N2328, N2296, N563, N1016);
nor NOR3 (N2329, N2328, N1939, N1851);
nor NOR3 (N2330, N2311, N147, N1416);
nor NOR2 (N2331, N2322, N561);
nand NAND2 (N2332, N2327, N2252);
xor XOR2 (N2333, N2324, N310);
xor XOR2 (N2334, N2332, N1461);
and AND3 (N2335, N2325, N2122, N1624);
xor XOR2 (N2336, N2317, N2030);
buf BUF1 (N2337, N2323);
and AND3 (N2338, N2326, N1646, N692);
and AND2 (N2339, N2334, N1650);
or OR4 (N2340, N2316, N1826, N1302, N506);
not NOT1 (N2341, N2335);
nand NAND2 (N2342, N2337, N1433);
or OR4 (N2343, N2341, N264, N566, N998);
and AND3 (N2344, N2331, N581, N133);
or OR4 (N2345, N2338, N867, N666, N1708);
nand NAND3 (N2346, N2345, N1805, N175);
or OR3 (N2347, N2329, N2316, N2195);
or OR3 (N2348, N2333, N2346, N1726);
xor XOR2 (N2349, N2225, N567);
buf BUF1 (N2350, N2340);
and AND3 (N2351, N2342, N1459, N1575);
nor NOR2 (N2352, N2351, N1891);
buf BUF1 (N2353, N2344);
xor XOR2 (N2354, N2353, N1486);
xor XOR2 (N2355, N2336, N348);
buf BUF1 (N2356, N2330);
nand NAND3 (N2357, N2355, N1260, N1176);
nor NOR2 (N2358, N2339, N770);
nor NOR2 (N2359, N2348, N1891);
or OR4 (N2360, N2343, N318, N1597, N1789);
nand NAND2 (N2361, N2356, N333);
and AND2 (N2362, N2359, N1667);
buf BUF1 (N2363, N2354);
nor NOR2 (N2364, N2360, N257);
nor NOR4 (N2365, N2349, N1376, N1195, N270);
not NOT1 (N2366, N2364);
and AND4 (N2367, N2357, N2046, N1377, N1749);
or OR4 (N2368, N2367, N2034, N1575, N1600);
and AND4 (N2369, N2361, N1503, N720, N2194);
and AND3 (N2370, N2365, N2363, N367);
nand NAND4 (N2371, N848, N1539, N856, N1091);
buf BUF1 (N2372, N2362);
and AND2 (N2373, N2370, N1330);
nand NAND2 (N2374, N2369, N666);
not NOT1 (N2375, N2350);
xor XOR2 (N2376, N2366, N2339);
nor NOR3 (N2377, N2375, N1547, N1924);
nor NOR2 (N2378, N2368, N1954);
and AND2 (N2379, N2358, N532);
buf BUF1 (N2380, N2352);
nand NAND4 (N2381, N2347, N1437, N1586, N393);
not NOT1 (N2382, N2374);
nand NAND2 (N2383, N2371, N58);
not NOT1 (N2384, N2380);
xor XOR2 (N2385, N2384, N584);
xor XOR2 (N2386, N2377, N841);
nand NAND3 (N2387, N2381, N2156, N618);
xor XOR2 (N2388, N2373, N829);
not NOT1 (N2389, N2385);
or OR3 (N2390, N2388, N1708, N977);
and AND2 (N2391, N2389, N2138);
or OR4 (N2392, N2378, N5, N1149, N1643);
nand NAND3 (N2393, N2390, N799, N349);
or OR3 (N2394, N2379, N1556, N1904);
nor NOR4 (N2395, N2372, N881, N1570, N1888);
nor NOR3 (N2396, N2376, N2143, N1876);
nand NAND4 (N2397, N2383, N188, N741, N327);
buf BUF1 (N2398, N2392);
or OR4 (N2399, N2396, N2186, N228, N1236);
buf BUF1 (N2400, N2397);
nor NOR2 (N2401, N2393, N1435);
buf BUF1 (N2402, N2401);
and AND4 (N2403, N2394, N562, N240, N6);
buf BUF1 (N2404, N2398);
or OR2 (N2405, N2387, N1027);
and AND2 (N2406, N2382, N732);
not NOT1 (N2407, N2391);
nor NOR4 (N2408, N2395, N1552, N1991, N901);
nand NAND4 (N2409, N2399, N893, N1195, N702);
not NOT1 (N2410, N2404);
nor NOR3 (N2411, N2409, N1301, N2231);
nor NOR2 (N2412, N2400, N1089);
buf BUF1 (N2413, N2403);
nor NOR4 (N2414, N2402, N1887, N2359, N1669);
or OR4 (N2415, N2407, N1892, N791, N222);
nor NOR2 (N2416, N2410, N1754);
nor NOR4 (N2417, N2408, N1180, N2269, N1272);
buf BUF1 (N2418, N2411);
nor NOR4 (N2419, N2413, N124, N1115, N470);
and AND4 (N2420, N2415, N717, N721, N493);
and AND2 (N2421, N2406, N1485);
nor NOR2 (N2422, N2405, N200);
and AND4 (N2423, N2419, N691, N1516, N526);
and AND2 (N2424, N2423, N1882);
buf BUF1 (N2425, N2417);
nand NAND3 (N2426, N2416, N2193, N2273);
xor XOR2 (N2427, N2426, N162);
nand NAND4 (N2428, N2424, N1541, N1832, N1876);
buf BUF1 (N2429, N2427);
and AND4 (N2430, N2428, N2170, N775, N194);
buf BUF1 (N2431, N2386);
buf BUF1 (N2432, N2414);
nor NOR4 (N2433, N2425, N618, N63, N1165);
nand NAND4 (N2434, N2429, N183, N790, N807);
and AND4 (N2435, N2433, N417, N1558, N876);
buf BUF1 (N2436, N2412);
xor XOR2 (N2437, N2432, N1858);
nor NOR4 (N2438, N2437, N413, N970, N1069);
and AND4 (N2439, N2431, N1181, N1864, N1455);
xor XOR2 (N2440, N2422, N196);
nor NOR3 (N2441, N2418, N456, N1737);
or OR2 (N2442, N2434, N935);
and AND2 (N2443, N2439, N835);
nor NOR3 (N2444, N2441, N1753, N1791);
nor NOR4 (N2445, N2443, N73, N302, N1884);
buf BUF1 (N2446, N2430);
nor NOR2 (N2447, N2420, N1938);
or OR3 (N2448, N2447, N500, N2391);
or OR3 (N2449, N2435, N808, N399);
not NOT1 (N2450, N2448);
xor XOR2 (N2451, N2436, N154);
xor XOR2 (N2452, N2450, N587);
nor NOR2 (N2453, N2451, N896);
nor NOR4 (N2454, N2421, N1379, N247, N1304);
buf BUF1 (N2455, N2452);
buf BUF1 (N2456, N2454);
not NOT1 (N2457, N2440);
xor XOR2 (N2458, N2444, N789);
or OR4 (N2459, N2456, N742, N1473, N1793);
xor XOR2 (N2460, N2455, N885);
or OR4 (N2461, N2460, N1705, N578, N1299);
nor NOR2 (N2462, N2459, N108);
or OR3 (N2463, N2453, N398, N333);
nand NAND3 (N2464, N2446, N252, N68);
not NOT1 (N2465, N2463);
and AND4 (N2466, N2457, N2358, N1069, N1492);
nor NOR2 (N2467, N2466, N486);
xor XOR2 (N2468, N2467, N623);
and AND4 (N2469, N2465, N470, N2196, N47);
xor XOR2 (N2470, N2458, N2237);
buf BUF1 (N2471, N2470);
or OR4 (N2472, N2445, N1793, N940, N1942);
nor NOR3 (N2473, N2464, N1201, N243);
not NOT1 (N2474, N2462);
and AND2 (N2475, N2438, N1151);
nand NAND3 (N2476, N2472, N928, N1889);
or OR2 (N2477, N2469, N2137);
nor NOR4 (N2478, N2473, N284, N1875, N374);
and AND4 (N2479, N2442, N1467, N2368, N1813);
not NOT1 (N2480, N2471);
xor XOR2 (N2481, N2474, N1084);
or OR4 (N2482, N2480, N1461, N967, N2108);
buf BUF1 (N2483, N2468);
buf BUF1 (N2484, N2477);
xor XOR2 (N2485, N2482, N1585);
or OR3 (N2486, N2461, N1879, N2134);
nor NOR4 (N2487, N2449, N1292, N1493, N1338);
xor XOR2 (N2488, N2475, N1924);
or OR4 (N2489, N2488, N844, N1879, N1448);
xor XOR2 (N2490, N2478, N2271);
xor XOR2 (N2491, N2476, N1624);
nor NOR2 (N2492, N2485, N1921);
not NOT1 (N2493, N2487);
xor XOR2 (N2494, N2491, N2079);
and AND2 (N2495, N2492, N1879);
not NOT1 (N2496, N2481);
buf BUF1 (N2497, N2490);
nor NOR4 (N2498, N2493, N1192, N109, N1442);
not NOT1 (N2499, N2495);
or OR2 (N2500, N2497, N2370);
nor NOR2 (N2501, N2486, N2445);
or OR4 (N2502, N2500, N1462, N1915, N1426);
xor XOR2 (N2503, N2483, N1358);
nand NAND2 (N2504, N2484, N1798);
nand NAND4 (N2505, N2498, N1439, N1335, N2478);
nand NAND3 (N2506, N2479, N1094, N850);
nand NAND2 (N2507, N2504, N73);
and AND4 (N2508, N2506, N167, N2369, N2306);
nand NAND4 (N2509, N2499, N333, N1130, N315);
buf BUF1 (N2510, N2489);
nand NAND4 (N2511, N2503, N423, N2379, N1763);
and AND4 (N2512, N2502, N828, N2265, N577);
xor XOR2 (N2513, N2501, N346);
buf BUF1 (N2514, N2505);
not NOT1 (N2515, N2510);
and AND3 (N2516, N2515, N149, N112);
not NOT1 (N2517, N2513);
or OR4 (N2518, N2512, N1172, N382, N2513);
nand NAND4 (N2519, N2518, N931, N606, N2107);
nor NOR4 (N2520, N2514, N1203, N1306, N1095);
nand NAND2 (N2521, N2508, N2148);
buf BUF1 (N2522, N2521);
xor XOR2 (N2523, N2494, N1616);
buf BUF1 (N2524, N2509);
and AND4 (N2525, N2519, N202, N1039, N332);
or OR4 (N2526, N2517, N132, N505, N125);
or OR4 (N2527, N2525, N380, N642, N571);
buf BUF1 (N2528, N2524);
or OR4 (N2529, N2520, N1700, N2116, N1850);
and AND3 (N2530, N2529, N611, N521);
xor XOR2 (N2531, N2523, N2079);
not NOT1 (N2532, N2511);
xor XOR2 (N2533, N2527, N1903);
not NOT1 (N2534, N2496);
and AND2 (N2535, N2526, N372);
buf BUF1 (N2536, N2528);
and AND3 (N2537, N2530, N2409, N2254);
xor XOR2 (N2538, N2522, N2147);
and AND2 (N2539, N2537, N2165);
and AND2 (N2540, N2536, N219);
buf BUF1 (N2541, N2538);
buf BUF1 (N2542, N2540);
not NOT1 (N2543, N2533);
or OR2 (N2544, N2532, N2356);
xor XOR2 (N2545, N2539, N755);
nand NAND4 (N2546, N2543, N2502, N552, N1780);
or OR4 (N2547, N2531, N2051, N970, N1690);
or OR4 (N2548, N2544, N1698, N2234, N1802);
or OR2 (N2549, N2542, N90);
xor XOR2 (N2550, N2535, N1036);
xor XOR2 (N2551, N2548, N1137);
nand NAND4 (N2552, N2547, N1479, N2089, N75);
nor NOR2 (N2553, N2516, N1892);
nor NOR2 (N2554, N2551, N1586);
not NOT1 (N2555, N2545);
not NOT1 (N2556, N2555);
xor XOR2 (N2557, N2549, N578);
not NOT1 (N2558, N2546);
xor XOR2 (N2559, N2558, N2440);
not NOT1 (N2560, N2553);
not NOT1 (N2561, N2556);
nor NOR3 (N2562, N2557, N961, N2329);
xor XOR2 (N2563, N2534, N960);
nand NAND2 (N2564, N2560, N2358);
buf BUF1 (N2565, N2564);
xor XOR2 (N2566, N2541, N1018);
nor NOR3 (N2567, N2562, N2548, N345);
or OR4 (N2568, N2561, N1474, N829, N1971);
and AND4 (N2569, N2552, N206, N1067, N2491);
and AND2 (N2570, N2559, N2499);
or OR4 (N2571, N2568, N1519, N663, N718);
and AND3 (N2572, N2569, N2530, N2274);
and AND4 (N2573, N2570, N1921, N221, N551);
xor XOR2 (N2574, N2566, N1264);
nor NOR3 (N2575, N2563, N1441, N2147);
not NOT1 (N2576, N2574);
or OR3 (N2577, N2567, N964, N2259);
xor XOR2 (N2578, N2571, N271);
or OR4 (N2579, N2507, N460, N1814, N745);
and AND2 (N2580, N2565, N1622);
xor XOR2 (N2581, N2577, N422);
not NOT1 (N2582, N2581);
buf BUF1 (N2583, N2576);
or OR2 (N2584, N2550, N610);
not NOT1 (N2585, N2572);
nor NOR2 (N2586, N2580, N544);
xor XOR2 (N2587, N2573, N942);
or OR4 (N2588, N2587, N2429, N1211, N2357);
nor NOR2 (N2589, N2588, N2211);
and AND2 (N2590, N2589, N773);
nand NAND3 (N2591, N2586, N751, N546);
xor XOR2 (N2592, N2584, N539);
nor NOR4 (N2593, N2585, N1136, N88, N416);
not NOT1 (N2594, N2591);
not NOT1 (N2595, N2583);
xor XOR2 (N2596, N2590, N867);
xor XOR2 (N2597, N2582, N2184);
xor XOR2 (N2598, N2596, N1683);
xor XOR2 (N2599, N2594, N878);
buf BUF1 (N2600, N2575);
not NOT1 (N2601, N2595);
xor XOR2 (N2602, N2554, N228);
or OR4 (N2603, N2599, N2321, N1268, N1888);
nor NOR3 (N2604, N2579, N1449, N1688);
buf BUF1 (N2605, N2592);
nand NAND2 (N2606, N2600, N1812);
or OR3 (N2607, N2598, N2557, N2194);
buf BUF1 (N2608, N2603);
xor XOR2 (N2609, N2578, N173);
or OR3 (N2610, N2597, N434, N1797);
or OR4 (N2611, N2610, N1203, N100, N947);
buf BUF1 (N2612, N2609);
nand NAND2 (N2613, N2612, N1363);
xor XOR2 (N2614, N2601, N798);
and AND2 (N2615, N2611, N585);
nand NAND3 (N2616, N2605, N1375, N1571);
buf BUF1 (N2617, N2608);
xor XOR2 (N2618, N2616, N1187);
or OR3 (N2619, N2607, N210, N1793);
buf BUF1 (N2620, N2604);
nand NAND4 (N2621, N2620, N1523, N799, N1401);
nand NAND3 (N2622, N2593, N783, N2447);
not NOT1 (N2623, N2615);
nor NOR4 (N2624, N2606, N1896, N605, N905);
and AND4 (N2625, N2624, N1994, N581, N1092);
nand NAND3 (N2626, N2602, N1457, N2283);
or OR4 (N2627, N2613, N2138, N2426, N541);
buf BUF1 (N2628, N2619);
buf BUF1 (N2629, N2627);
xor XOR2 (N2630, N2618, N2021);
and AND3 (N2631, N2626, N2253, N825);
and AND3 (N2632, N2617, N293, N891);
xor XOR2 (N2633, N2632, N1572);
buf BUF1 (N2634, N2614);
xor XOR2 (N2635, N2622, N790);
buf BUF1 (N2636, N2628);
not NOT1 (N2637, N2633);
and AND4 (N2638, N2634, N1760, N756, N206);
nor NOR3 (N2639, N2621, N1442, N963);
nand NAND3 (N2640, N2623, N1817, N1760);
and AND4 (N2641, N2635, N34, N12, N1940);
not NOT1 (N2642, N2629);
xor XOR2 (N2643, N2638, N581);
not NOT1 (N2644, N2639);
and AND3 (N2645, N2640, N1906, N1428);
and AND4 (N2646, N2636, N2120, N1421, N1131);
or OR3 (N2647, N2642, N574, N254);
buf BUF1 (N2648, N2641);
not NOT1 (N2649, N2644);
not NOT1 (N2650, N2643);
and AND3 (N2651, N2630, N1213, N793);
and AND4 (N2652, N2649, N330, N1509, N2328);
and AND4 (N2653, N2646, N247, N988, N845);
not NOT1 (N2654, N2650);
and AND4 (N2655, N2651, N1433, N382, N706);
not NOT1 (N2656, N2645);
not NOT1 (N2657, N2648);
xor XOR2 (N2658, N2654, N2081);
not NOT1 (N2659, N2625);
nor NOR3 (N2660, N2637, N823, N1948);
not NOT1 (N2661, N2659);
or OR4 (N2662, N2655, N1635, N554, N459);
buf BUF1 (N2663, N2658);
and AND2 (N2664, N2647, N1093);
nand NAND2 (N2665, N2663, N75);
xor XOR2 (N2666, N2652, N1067);
buf BUF1 (N2667, N2665);
and AND3 (N2668, N2661, N373, N2036);
nor NOR3 (N2669, N2656, N368, N2033);
nor NOR2 (N2670, N2631, N825);
not NOT1 (N2671, N2662);
or OR3 (N2672, N2664, N2390, N1889);
not NOT1 (N2673, N2667);
nor NOR2 (N2674, N2668, N14);
or OR4 (N2675, N2660, N1551, N88, N753);
nand NAND4 (N2676, N2666, N1972, N1071, N2203);
xor XOR2 (N2677, N2671, N1635);
nand NAND3 (N2678, N2657, N50, N331);
or OR3 (N2679, N2676, N306, N1525);
buf BUF1 (N2680, N2669);
not NOT1 (N2681, N2675);
and AND4 (N2682, N2672, N1385, N2055, N2051);
or OR4 (N2683, N2674, N1926, N123, N1316);
not NOT1 (N2684, N2653);
xor XOR2 (N2685, N2682, N2146);
or OR3 (N2686, N2678, N198, N2550);
and AND2 (N2687, N2684, N728);
xor XOR2 (N2688, N2670, N1278);
not NOT1 (N2689, N2683);
and AND2 (N2690, N2689, N2501);
not NOT1 (N2691, N2685);
or OR3 (N2692, N2681, N2585, N1399);
xor XOR2 (N2693, N2677, N755);
nand NAND2 (N2694, N2690, N1261);
nand NAND2 (N2695, N2694, N2561);
xor XOR2 (N2696, N2693, N2601);
not NOT1 (N2697, N2686);
nand NAND3 (N2698, N2688, N2300, N1795);
or OR2 (N2699, N2680, N2439);
buf BUF1 (N2700, N2699);
xor XOR2 (N2701, N2687, N1559);
and AND3 (N2702, N2696, N1113, N416);
buf BUF1 (N2703, N2700);
xor XOR2 (N2704, N2702, N2004);
xor XOR2 (N2705, N2703, N2378);
and AND3 (N2706, N2692, N1378, N2025);
nand NAND4 (N2707, N2695, N1636, N2178, N783);
or OR3 (N2708, N2697, N1234, N1975);
nor NOR4 (N2709, N2707, N1541, N2513, N341);
not NOT1 (N2710, N2701);
xor XOR2 (N2711, N2704, N1096);
buf BUF1 (N2712, N2691);
buf BUF1 (N2713, N2679);
nor NOR3 (N2714, N2673, N1942, N1686);
nand NAND3 (N2715, N2714, N7, N1159);
and AND2 (N2716, N2712, N684);
nor NOR4 (N2717, N2709, N803, N1490, N982);
and AND2 (N2718, N2717, N1122);
and AND3 (N2719, N2718, N2663, N2187);
or OR2 (N2720, N2713, N1614);
nor NOR4 (N2721, N2720, N1258, N2384, N234);
and AND2 (N2722, N2715, N1759);
not NOT1 (N2723, N2705);
nand NAND3 (N2724, N2698, N777, N2314);
not NOT1 (N2725, N2724);
or OR2 (N2726, N2708, N190);
and AND3 (N2727, N2716, N964, N516);
buf BUF1 (N2728, N2725);
nand NAND4 (N2729, N2710, N189, N1008, N2324);
and AND4 (N2730, N2711, N537, N1615, N1950);
not NOT1 (N2731, N2728);
nand NAND3 (N2732, N2730, N180, N1987);
xor XOR2 (N2733, N2721, N2308);
or OR4 (N2734, N2726, N650, N879, N2005);
xor XOR2 (N2735, N2723, N1135);
nor NOR3 (N2736, N2706, N247, N1621);
nand NAND4 (N2737, N2729, N2689, N93, N78);
or OR2 (N2738, N2732, N113);
nor NOR2 (N2739, N2719, N1869);
not NOT1 (N2740, N2734);
and AND2 (N2741, N2735, N1813);
buf BUF1 (N2742, N2722);
buf BUF1 (N2743, N2733);
nor NOR4 (N2744, N2743, N937, N2248, N780);
and AND4 (N2745, N2731, N1984, N2174, N2586);
and AND3 (N2746, N2736, N2473, N315);
buf BUF1 (N2747, N2737);
xor XOR2 (N2748, N2745, N294);
nand NAND2 (N2749, N2744, N488);
nand NAND3 (N2750, N2742, N2242, N1855);
nor NOR4 (N2751, N2740, N2683, N2167, N1564);
and AND3 (N2752, N2727, N1706, N1491);
nor NOR2 (N2753, N2746, N1488);
or OR4 (N2754, N2749, N2113, N369, N2301);
buf BUF1 (N2755, N2753);
nand NAND2 (N2756, N2739, N1407);
buf BUF1 (N2757, N2754);
and AND4 (N2758, N2752, N779, N1721, N1357);
nor NOR3 (N2759, N2757, N1340, N438);
xor XOR2 (N2760, N2758, N2413);
nor NOR3 (N2761, N2755, N217, N1360);
nor NOR3 (N2762, N2750, N611, N975);
nor NOR2 (N2763, N2760, N1222);
and AND3 (N2764, N2761, N1031, N2761);
and AND3 (N2765, N2764, N2502, N926);
nor NOR4 (N2766, N2748, N2139, N369, N2499);
xor XOR2 (N2767, N2765, N2318);
buf BUF1 (N2768, N2741);
nand NAND2 (N2769, N2762, N2727);
and AND3 (N2770, N2738, N542, N2078);
and AND3 (N2771, N2769, N577, N1510);
not NOT1 (N2772, N2766);
or OR4 (N2773, N2772, N1465, N1473, N669);
or OR4 (N2774, N2759, N36, N2380, N1357);
not NOT1 (N2775, N2768);
nand NAND3 (N2776, N2763, N232, N109);
xor XOR2 (N2777, N2770, N2110);
and AND3 (N2778, N2771, N593, N880);
or OR2 (N2779, N2756, N1407);
nand NAND2 (N2780, N2751, N299);
and AND3 (N2781, N2773, N865, N136);
nor NOR4 (N2782, N2775, N1352, N2587, N2762);
xor XOR2 (N2783, N2780, N2777);
buf BUF1 (N2784, N1140);
buf BUF1 (N2785, N2784);
nand NAND3 (N2786, N2785, N2210, N621);
not NOT1 (N2787, N2778);
nand NAND4 (N2788, N2781, N900, N1005, N74);
not NOT1 (N2789, N2776);
nand NAND4 (N2790, N2787, N594, N2206, N2155);
xor XOR2 (N2791, N2786, N232);
buf BUF1 (N2792, N2790);
nand NAND2 (N2793, N2782, N1621);
not NOT1 (N2794, N2774);
and AND3 (N2795, N2747, N2016, N1603);
or OR4 (N2796, N2795, N2471, N1823, N2175);
not NOT1 (N2797, N2783);
and AND2 (N2798, N2792, N2670);
not NOT1 (N2799, N2791);
xor XOR2 (N2800, N2767, N2726);
nand NAND2 (N2801, N2793, N438);
nand NAND4 (N2802, N2789, N1932, N1196, N1033);
not NOT1 (N2803, N2798);
not NOT1 (N2804, N2797);
and AND3 (N2805, N2788, N385, N1575);
buf BUF1 (N2806, N2802);
and AND2 (N2807, N2799, N2391);
or OR4 (N2808, N2779, N109, N2308, N2650);
nand NAND2 (N2809, N2804, N1577);
not NOT1 (N2810, N2800);
or OR4 (N2811, N2810, N1277, N495, N2086);
xor XOR2 (N2812, N2806, N1197);
nor NOR4 (N2813, N2811, N2528, N1746, N1227);
or OR2 (N2814, N2813, N1673);
or OR2 (N2815, N2801, N754);
nand NAND3 (N2816, N2807, N1408, N38);
or OR2 (N2817, N2805, N2211);
nor NOR4 (N2818, N2794, N546, N1990, N242);
xor XOR2 (N2819, N2809, N1855);
nor NOR4 (N2820, N2817, N843, N434, N296);
and AND2 (N2821, N2818, N2158);
buf BUF1 (N2822, N2819);
nand NAND3 (N2823, N2821, N2211, N916);
nor NOR4 (N2824, N2820, N245, N1730, N370);
or OR4 (N2825, N2815, N2404, N2037, N291);
or OR2 (N2826, N2796, N2226);
buf BUF1 (N2827, N2824);
nand NAND4 (N2828, N2825, N1025, N178, N1057);
and AND4 (N2829, N2803, N1637, N2423, N2745);
buf BUF1 (N2830, N2828);
buf BUF1 (N2831, N2829);
and AND4 (N2832, N2812, N1999, N932, N658);
buf BUF1 (N2833, N2832);
and AND4 (N2834, N2808, N756, N2272, N1615);
xor XOR2 (N2835, N2822, N2654);
nand NAND2 (N2836, N2833, N786);
and AND4 (N2837, N2834, N756, N1647, N191);
or OR4 (N2838, N2823, N1815, N197, N756);
and AND4 (N2839, N2830, N830, N2626, N285);
nand NAND4 (N2840, N2826, N1939, N2067, N1889);
or OR3 (N2841, N2814, N2628, N2561);
buf BUF1 (N2842, N2827);
xor XOR2 (N2843, N2837, N163);
not NOT1 (N2844, N2838);
nor NOR3 (N2845, N2842, N2814, N2488);
nand NAND2 (N2846, N2839, N455);
xor XOR2 (N2847, N2840, N1088);
not NOT1 (N2848, N2843);
buf BUF1 (N2849, N2846);
xor XOR2 (N2850, N2848, N593);
and AND4 (N2851, N2831, N2196, N2789, N2294);
nand NAND3 (N2852, N2841, N1522, N818);
nand NAND3 (N2853, N2844, N1190, N2777);
or OR3 (N2854, N2849, N149, N774);
buf BUF1 (N2855, N2853);
buf BUF1 (N2856, N2845);
xor XOR2 (N2857, N2835, N661);
xor XOR2 (N2858, N2847, N1963);
xor XOR2 (N2859, N2850, N1736);
not NOT1 (N2860, N2854);
and AND2 (N2861, N2856, N1028);
not NOT1 (N2862, N2855);
not NOT1 (N2863, N2858);
nor NOR2 (N2864, N2836, N2847);
xor XOR2 (N2865, N2864, N1524);
not NOT1 (N2866, N2865);
nor NOR3 (N2867, N2857, N1065, N2491);
not NOT1 (N2868, N2816);
or OR4 (N2869, N2859, N2513, N832, N469);
or OR3 (N2870, N2862, N2083, N456);
not NOT1 (N2871, N2863);
buf BUF1 (N2872, N2852);
and AND3 (N2873, N2851, N1031, N214);
and AND4 (N2874, N2866, N1663, N1615, N2753);
or OR3 (N2875, N2874, N1926, N550);
buf BUF1 (N2876, N2871);
buf BUF1 (N2877, N2870);
nand NAND2 (N2878, N2861, N1240);
not NOT1 (N2879, N2872);
buf BUF1 (N2880, N2876);
not NOT1 (N2881, N2878);
nand NAND2 (N2882, N2880, N308);
or OR4 (N2883, N2873, N707, N2302, N2708);
xor XOR2 (N2884, N2881, N1876);
or OR3 (N2885, N2883, N738, N1804);
or OR3 (N2886, N2885, N1771, N2272);
or OR2 (N2887, N2886, N1719);
not NOT1 (N2888, N2875);
and AND3 (N2889, N2860, N2423, N1284);
buf BUF1 (N2890, N2882);
not NOT1 (N2891, N2889);
nand NAND3 (N2892, N2867, N1302, N182);
buf BUF1 (N2893, N2877);
and AND4 (N2894, N2890, N1384, N979, N1293);
and AND3 (N2895, N2879, N2789, N2553);
and AND2 (N2896, N2887, N1058);
and AND4 (N2897, N2869, N2443, N2333, N1822);
and AND3 (N2898, N2895, N1559, N300);
xor XOR2 (N2899, N2892, N1924);
xor XOR2 (N2900, N2898, N1154);
nand NAND4 (N2901, N2899, N2257, N2549, N2315);
or OR4 (N2902, N2901, N1633, N1584, N680);
or OR4 (N2903, N2891, N543, N2628, N490);
nor NOR2 (N2904, N2897, N632);
or OR3 (N2905, N2888, N389, N585);
not NOT1 (N2906, N2904);
or OR3 (N2907, N2905, N1566, N433);
nand NAND4 (N2908, N2868, N1855, N2606, N971);
buf BUF1 (N2909, N2906);
or OR4 (N2910, N2894, N1356, N127, N2745);
buf BUF1 (N2911, N2903);
nand NAND4 (N2912, N2900, N1804, N145, N2733);
nor NOR3 (N2913, N2911, N1191, N2576);
or OR4 (N2914, N2896, N526, N2360, N566);
or OR3 (N2915, N2913, N380, N1525);
not NOT1 (N2916, N2912);
or OR3 (N2917, N2908, N2458, N706);
buf BUF1 (N2918, N2915);
and AND2 (N2919, N2917, N2222);
and AND4 (N2920, N2909, N2090, N1374, N2468);
and AND4 (N2921, N2919, N1694, N843, N70);
nor NOR3 (N2922, N2884, N740, N1073);
buf BUF1 (N2923, N2916);
buf BUF1 (N2924, N2920);
buf BUF1 (N2925, N2924);
xor XOR2 (N2926, N2918, N859);
nand NAND2 (N2927, N2923, N299);
and AND4 (N2928, N2914, N1993, N2293, N1307);
and AND2 (N2929, N2893, N178);
or OR3 (N2930, N2910, N1987, N1091);
xor XOR2 (N2931, N2921, N878);
buf BUF1 (N2932, N2931);
not NOT1 (N2933, N2929);
nor NOR3 (N2934, N2930, N2357, N2570);
or OR2 (N2935, N2934, N2776);
xor XOR2 (N2936, N2932, N1113);
buf BUF1 (N2937, N2927);
and AND4 (N2938, N2933, N2829, N900, N2061);
xor XOR2 (N2939, N2938, N2216);
buf BUF1 (N2940, N2935);
nand NAND3 (N2941, N2939, N2024, N1099);
not NOT1 (N2942, N2940);
nor NOR4 (N2943, N2937, N188, N1691, N179);
and AND4 (N2944, N2907, N2870, N18, N850);
nor NOR3 (N2945, N2941, N797, N2045);
nand NAND2 (N2946, N2902, N2198);
and AND2 (N2947, N2922, N1994);
nor NOR3 (N2948, N2947, N2082, N1053);
nand NAND3 (N2949, N2948, N2888, N823);
nor NOR2 (N2950, N2944, N284);
not NOT1 (N2951, N2928);
buf BUF1 (N2952, N2943);
xor XOR2 (N2953, N2936, N1654);
not NOT1 (N2954, N2949);
nor NOR4 (N2955, N2925, N2043, N291, N1230);
or OR2 (N2956, N2951, N2885);
nor NOR3 (N2957, N2942, N564, N870);
not NOT1 (N2958, N2926);
nor NOR3 (N2959, N2954, N843, N520);
and AND4 (N2960, N2946, N761, N1096, N963);
and AND2 (N2961, N2957, N2502);
nand NAND2 (N2962, N2956, N1417);
not NOT1 (N2963, N2959);
nor NOR3 (N2964, N2952, N2859, N2422);
nand NAND3 (N2965, N2958, N1901, N799);
and AND2 (N2966, N2964, N1030);
and AND3 (N2967, N2945, N2234, N2813);
nand NAND3 (N2968, N2961, N1544, N136);
and AND3 (N2969, N2966, N1776, N291);
nor NOR3 (N2970, N2968, N174, N69);
or OR3 (N2971, N2962, N2074, N407);
nand NAND4 (N2972, N2955, N196, N17, N410);
not NOT1 (N2973, N2963);
buf BUF1 (N2974, N2950);
xor XOR2 (N2975, N2971, N1439);
buf BUF1 (N2976, N2953);
or OR4 (N2977, N2967, N343, N943, N129);
or OR3 (N2978, N2969, N443, N1897);
not NOT1 (N2979, N2970);
or OR2 (N2980, N2975, N570);
or OR4 (N2981, N2973, N1249, N121, N2515);
not NOT1 (N2982, N2974);
buf BUF1 (N2983, N2978);
and AND4 (N2984, N2982, N2013, N741, N1147);
and AND4 (N2985, N2980, N2653, N428, N511);
xor XOR2 (N2986, N2983, N638);
nand NAND2 (N2987, N2986, N797);
and AND2 (N2988, N2984, N180);
xor XOR2 (N2989, N2965, N1966);
or OR2 (N2990, N2988, N639);
nor NOR2 (N2991, N2977, N1239);
nor NOR4 (N2992, N2981, N2028, N969, N328);
or OR3 (N2993, N2989, N1882, N204);
and AND3 (N2994, N2993, N31, N1695);
xor XOR2 (N2995, N2979, N2189);
nor NOR2 (N2996, N2992, N2032);
or OR3 (N2997, N2991, N2288, N2820);
buf BUF1 (N2998, N2976);
or OR2 (N2999, N2996, N1613);
xor XOR2 (N3000, N2990, N2685);
buf BUF1 (N3001, N2985);
xor XOR2 (N3002, N2999, N1960);
nor NOR4 (N3003, N3002, N467, N2936, N676);
or OR4 (N3004, N2987, N858, N1069, N1382);
or OR4 (N3005, N2960, N2240, N2082, N1085);
and AND4 (N3006, N2997, N2609, N2393, N1510);
buf BUF1 (N3007, N3006);
nor NOR3 (N3008, N2995, N2504, N853);
buf BUF1 (N3009, N3003);
nand NAND2 (N3010, N3001, N2303);
xor XOR2 (N3011, N2998, N2739);
nand NAND3 (N3012, N3004, N566, N861);
or OR3 (N3013, N3009, N205, N273);
not NOT1 (N3014, N3010);
xor XOR2 (N3015, N3012, N1630);
xor XOR2 (N3016, N3005, N82);
buf BUF1 (N3017, N3011);
xor XOR2 (N3018, N3008, N397);
not NOT1 (N3019, N3016);
xor XOR2 (N3020, N3017, N501);
and AND4 (N3021, N3019, N2522, N2261, N1887);
not NOT1 (N3022, N3015);
nor NOR4 (N3023, N3018, N2147, N2365, N929);
and AND2 (N3024, N3023, N1993);
or OR3 (N3025, N3021, N2231, N1649);
buf BUF1 (N3026, N3014);
and AND2 (N3027, N3026, N800);
nand NAND4 (N3028, N2972, N2273, N623, N1307);
nor NOR4 (N3029, N3022, N155, N670, N2855);
not NOT1 (N3030, N3013);
or OR3 (N3031, N3020, N1143, N2879);
or OR4 (N3032, N3030, N373, N1438, N478);
nor NOR3 (N3033, N3000, N1210, N2572);
nand NAND3 (N3034, N3033, N1265, N517);
or OR4 (N3035, N3032, N2255, N2663, N2966);
and AND2 (N3036, N3029, N935);
xor XOR2 (N3037, N2994, N190);
and AND3 (N3038, N3031, N2000, N1923);
buf BUF1 (N3039, N3036);
and AND2 (N3040, N3025, N2617);
nand NAND3 (N3041, N3037, N137, N494);
xor XOR2 (N3042, N3007, N2695);
xor XOR2 (N3043, N3035, N1890);
nand NAND2 (N3044, N3043, N1931);
xor XOR2 (N3045, N3040, N995);
buf BUF1 (N3046, N3041);
and AND3 (N3047, N3045, N2557, N638);
not NOT1 (N3048, N3028);
nand NAND4 (N3049, N3039, N212, N2695, N1692);
buf BUF1 (N3050, N3047);
and AND4 (N3051, N3046, N2521, N2539, N672);
and AND3 (N3052, N3051, N37, N35);
buf BUF1 (N3053, N3034);
or OR2 (N3054, N3027, N2273);
or OR3 (N3055, N3048, N2350, N2468);
or OR4 (N3056, N3054, N1053, N2066, N1077);
and AND3 (N3057, N3044, N1757, N2785);
not NOT1 (N3058, N3056);
nor NOR2 (N3059, N3042, N2477);
nand NAND4 (N3060, N3057, N592, N1119, N60);
xor XOR2 (N3061, N3050, N1529);
or OR4 (N3062, N3024, N1075, N1332, N1337);
not NOT1 (N3063, N3061);
not NOT1 (N3064, N3060);
or OR4 (N3065, N3049, N1177, N1863, N2089);
nand NAND4 (N3066, N3055, N2723, N1557, N829);
buf BUF1 (N3067, N3038);
xor XOR2 (N3068, N3064, N2144);
and AND3 (N3069, N3066, N2842, N1423);
buf BUF1 (N3070, N3065);
nor NOR3 (N3071, N3059, N1047, N273);
or OR4 (N3072, N3071, N1767, N2785, N1349);
or OR2 (N3073, N3070, N59);
and AND3 (N3074, N3073, N375, N2899);
buf BUF1 (N3075, N3063);
nand NAND4 (N3076, N3052, N756, N2635, N1953);
nor NOR4 (N3077, N3058, N2799, N1385, N2143);
or OR2 (N3078, N3076, N1420);
and AND2 (N3079, N3062, N3019);
and AND3 (N3080, N3072, N403, N1911);
or OR3 (N3081, N3078, N917, N13);
and AND2 (N3082, N3074, N2366);
xor XOR2 (N3083, N3067, N2721);
buf BUF1 (N3084, N3083);
xor XOR2 (N3085, N3082, N1538);
buf BUF1 (N3086, N3069);
and AND2 (N3087, N3077, N2415);
or OR4 (N3088, N3081, N2153, N537, N1190);
nand NAND3 (N3089, N3053, N1576, N2138);
buf BUF1 (N3090, N3089);
buf BUF1 (N3091, N3075);
buf BUF1 (N3092, N3084);
and AND3 (N3093, N3085, N289, N2556);
buf BUF1 (N3094, N3088);
xor XOR2 (N3095, N3068, N762);
not NOT1 (N3096, N3093);
nand NAND2 (N3097, N3079, N190);
not NOT1 (N3098, N3095);
nand NAND4 (N3099, N3087, N1846, N785, N350);
xor XOR2 (N3100, N3097, N2221);
or OR4 (N3101, N3092, N1005, N1624, N74);
nand NAND3 (N3102, N3094, N1366, N593);
or OR3 (N3103, N3080, N2403, N2472);
buf BUF1 (N3104, N3090);
or OR3 (N3105, N3086, N933, N2490);
buf BUF1 (N3106, N3104);
buf BUF1 (N3107, N3102);
buf BUF1 (N3108, N3106);
or OR4 (N3109, N3108, N2604, N828, N1081);
not NOT1 (N3110, N3098);
or OR2 (N3111, N3096, N1405);
buf BUF1 (N3112, N3111);
not NOT1 (N3113, N3110);
or OR4 (N3114, N3107, N2392, N2013, N313);
nand NAND3 (N3115, N3114, N2985, N2062);
nor NOR4 (N3116, N3112, N821, N453, N1716);
xor XOR2 (N3117, N3105, N430);
or OR2 (N3118, N3115, N1451);
nor NOR4 (N3119, N3117, N2774, N1930, N1445);
and AND4 (N3120, N3099, N2790, N1061, N152);
nand NAND2 (N3121, N3103, N3057);
not NOT1 (N3122, N3120);
not NOT1 (N3123, N3119);
nor NOR4 (N3124, N3100, N641, N835, N3072);
and AND2 (N3125, N3122, N857);
or OR4 (N3126, N3121, N1990, N675, N1000);
nor NOR2 (N3127, N3124, N1160);
buf BUF1 (N3128, N3101);
nand NAND4 (N3129, N3091, N1697, N591, N2478);
buf BUF1 (N3130, N3125);
and AND4 (N3131, N3123, N2212, N709, N983);
not NOT1 (N3132, N3127);
and AND3 (N3133, N3109, N2605, N60);
or OR4 (N3134, N3128, N404, N2504, N1680);
buf BUF1 (N3135, N3126);
or OR4 (N3136, N3118, N1293, N508, N2176);
not NOT1 (N3137, N3134);
nand NAND2 (N3138, N3135, N427);
and AND4 (N3139, N3138, N150, N2651, N921);
xor XOR2 (N3140, N3130, N2516);
or OR3 (N3141, N3136, N1936, N2871);
and AND3 (N3142, N3140, N793, N773);
xor XOR2 (N3143, N3133, N2797);
and AND2 (N3144, N3143, N2415);
or OR3 (N3145, N3139, N1590, N1152);
not NOT1 (N3146, N3113);
not NOT1 (N3147, N3129);
buf BUF1 (N3148, N3147);
not NOT1 (N3149, N3146);
nor NOR2 (N3150, N3149, N1176);
or OR3 (N3151, N3150, N1748, N314);
or OR2 (N3152, N3144, N1672);
nand NAND3 (N3153, N3132, N31, N2947);
and AND2 (N3154, N3152, N2654);
or OR4 (N3155, N3154, N133, N835, N1610);
nor NOR4 (N3156, N3137, N2136, N315, N1358);
nand NAND3 (N3157, N3142, N807, N2355);
and AND3 (N3158, N3157, N424, N2299);
buf BUF1 (N3159, N3153);
xor XOR2 (N3160, N3151, N1248);
and AND3 (N3161, N3156, N2666, N1859);
and AND4 (N3162, N3161, N408, N1782, N1513);
and AND4 (N3163, N3145, N2322, N2665, N608);
and AND2 (N3164, N3155, N2993);
nand NAND2 (N3165, N3131, N1780);
buf BUF1 (N3166, N3141);
nor NOR2 (N3167, N3166, N1410);
not NOT1 (N3168, N3162);
and AND3 (N3169, N3148, N1634, N1545);
xor XOR2 (N3170, N3160, N1049);
and AND2 (N3171, N3170, N1635);
buf BUF1 (N3172, N3169);
nor NOR2 (N3173, N3172, N2519);
and AND2 (N3174, N3116, N2438);
and AND4 (N3175, N3165, N370, N291, N2850);
or OR2 (N3176, N3168, N385);
nand NAND3 (N3177, N3175, N10, N1484);
buf BUF1 (N3178, N3159);
or OR3 (N3179, N3173, N373, N1758);
buf BUF1 (N3180, N3167);
and AND3 (N3181, N3158, N1001, N1218);
nand NAND2 (N3182, N3176, N2507);
and AND4 (N3183, N3178, N2213, N14, N3066);
or OR2 (N3184, N3181, N469);
not NOT1 (N3185, N3183);
nor NOR4 (N3186, N3177, N420, N1049, N886);
nor NOR4 (N3187, N3185, N2471, N125, N718);
not NOT1 (N3188, N3184);
xor XOR2 (N3189, N3187, N1987);
xor XOR2 (N3190, N3182, N537);
nand NAND4 (N3191, N3163, N3117, N2930, N978);
and AND3 (N3192, N3164, N1986, N2212);
nand NAND4 (N3193, N3189, N542, N1106, N1101);
nand NAND4 (N3194, N3186, N2660, N468, N1299);
nand NAND4 (N3195, N3180, N2953, N1553, N3182);
not NOT1 (N3196, N3188);
nor NOR4 (N3197, N3192, N1202, N2995, N512);
not NOT1 (N3198, N3195);
not NOT1 (N3199, N3197);
buf BUF1 (N3200, N3199);
or OR2 (N3201, N3194, N1061);
xor XOR2 (N3202, N3179, N1607);
nand NAND2 (N3203, N3202, N39);
xor XOR2 (N3204, N3190, N675);
nor NOR4 (N3205, N3191, N3040, N427, N2792);
nand NAND4 (N3206, N3201, N1474, N2686, N2063);
buf BUF1 (N3207, N3198);
buf BUF1 (N3208, N3204);
nor NOR2 (N3209, N3193, N20);
or OR4 (N3210, N3171, N1256, N676, N2863);
not NOT1 (N3211, N3174);
nor NOR3 (N3212, N3208, N1481, N2198);
xor XOR2 (N3213, N3200, N1073);
nand NAND4 (N3214, N3207, N1466, N1062, N1826);
not NOT1 (N3215, N3214);
buf BUF1 (N3216, N3203);
and AND3 (N3217, N3211, N2431, N1469);
xor XOR2 (N3218, N3216, N2958);
nand NAND3 (N3219, N3212, N2578, N802);
nand NAND3 (N3220, N3217, N550, N3212);
nor NOR2 (N3221, N3206, N152);
nor NOR4 (N3222, N3210, N3121, N445, N1952);
xor XOR2 (N3223, N3215, N2142);
not NOT1 (N3224, N3213);
nor NOR4 (N3225, N3209, N223, N1665, N3012);
not NOT1 (N3226, N3222);
and AND3 (N3227, N3221, N2014, N1120);
and AND3 (N3228, N3196, N844, N2748);
xor XOR2 (N3229, N3224, N1579);
not NOT1 (N3230, N3218);
and AND2 (N3231, N3220, N1354);
buf BUF1 (N3232, N3223);
xor XOR2 (N3233, N3225, N985);
or OR4 (N3234, N3233, N1043, N428, N46);
or OR4 (N3235, N3227, N2539, N859, N2943);
not NOT1 (N3236, N3234);
nor NOR4 (N3237, N3232, N1061, N1154, N2028);
or OR3 (N3238, N3235, N122, N2383);
xor XOR2 (N3239, N3238, N1258);
nand NAND3 (N3240, N3236, N1467, N1045);
not NOT1 (N3241, N3239);
or OR3 (N3242, N3226, N2685, N218);
nand NAND4 (N3243, N3205, N227, N1057, N519);
xor XOR2 (N3244, N3230, N1243);
xor XOR2 (N3245, N3231, N541);
xor XOR2 (N3246, N3229, N1118);
not NOT1 (N3247, N3237);
xor XOR2 (N3248, N3245, N383);
or OR3 (N3249, N3243, N2776, N2682);
nor NOR3 (N3250, N3228, N1899, N2651);
or OR2 (N3251, N3248, N3115);
nor NOR4 (N3252, N3240, N933, N191, N2716);
and AND3 (N3253, N3242, N1612, N789);
buf BUF1 (N3254, N3252);
nor NOR3 (N3255, N3249, N914, N1336);
buf BUF1 (N3256, N3244);
nand NAND3 (N3257, N3253, N1809, N404);
nor NOR2 (N3258, N3257, N2411);
or OR2 (N3259, N3256, N1542);
nand NAND2 (N3260, N3259, N428);
nand NAND2 (N3261, N3258, N1446);
and AND3 (N3262, N3255, N1892, N2467);
xor XOR2 (N3263, N3254, N1942);
xor XOR2 (N3264, N3246, N2268);
nand NAND4 (N3265, N3219, N1069, N1572, N1087);
xor XOR2 (N3266, N3251, N824);
or OR2 (N3267, N3262, N1552);
or OR4 (N3268, N3260, N2335, N2721, N1515);
buf BUF1 (N3269, N3266);
buf BUF1 (N3270, N3268);
xor XOR2 (N3271, N3263, N2330);
nand NAND2 (N3272, N3264, N2984);
or OR4 (N3273, N3250, N868, N2633, N1134);
nor NOR4 (N3274, N3261, N551, N854, N1144);
not NOT1 (N3275, N3273);
not NOT1 (N3276, N3265);
buf BUF1 (N3277, N3271);
and AND2 (N3278, N3277, N2032);
buf BUF1 (N3279, N3275);
nor NOR2 (N3280, N3269, N1948);
xor XOR2 (N3281, N3280, N1001);
nand NAND2 (N3282, N3267, N1455);
and AND3 (N3283, N3274, N2192, N1371);
not NOT1 (N3284, N3278);
and AND2 (N3285, N3247, N1423);
or OR3 (N3286, N3241, N2812, N2668);
xor XOR2 (N3287, N3270, N2288);
xor XOR2 (N3288, N3272, N2952);
and AND4 (N3289, N3287, N525, N1921, N3274);
nand NAND4 (N3290, N3282, N609, N595, N3247);
xor XOR2 (N3291, N3279, N3088);
or OR3 (N3292, N3281, N2297, N2602);
and AND2 (N3293, N3291, N2671);
nand NAND3 (N3294, N3283, N2277, N923);
xor XOR2 (N3295, N3289, N1644);
not NOT1 (N3296, N3290);
xor XOR2 (N3297, N3288, N2591);
nor NOR3 (N3298, N3286, N2826, N2673);
and AND4 (N3299, N3298, N2447, N1190, N916);
nand NAND3 (N3300, N3284, N2329, N1429);
buf BUF1 (N3301, N3295);
nor NOR2 (N3302, N3296, N2270);
or OR4 (N3303, N3276, N848, N1943, N1489);
and AND3 (N3304, N3301, N290, N2646);
and AND4 (N3305, N3293, N3099, N421, N986);
and AND4 (N3306, N3299, N2666, N1583, N1727);
buf BUF1 (N3307, N3304);
xor XOR2 (N3308, N3303, N2759);
or OR3 (N3309, N3300, N965, N1067);
nor NOR2 (N3310, N3292, N1153);
not NOT1 (N3311, N3310);
buf BUF1 (N3312, N3294);
not NOT1 (N3313, N3306);
or OR2 (N3314, N3305, N314);
nor NOR4 (N3315, N3309, N3006, N2219, N1735);
xor XOR2 (N3316, N3314, N1640);
or OR4 (N3317, N3316, N1386, N553, N1785);
not NOT1 (N3318, N3297);
nor NOR3 (N3319, N3313, N1537, N1337);
nor NOR3 (N3320, N3312, N2647, N2306);
xor XOR2 (N3321, N3308, N2731);
and AND3 (N3322, N3307, N59, N718);
or OR2 (N3323, N3317, N2893);
buf BUF1 (N3324, N3321);
nor NOR2 (N3325, N3320, N2749);
or OR4 (N3326, N3322, N1962, N2003, N3061);
nor NOR4 (N3327, N3326, N1199, N1396, N2997);
nor NOR3 (N3328, N3324, N3236, N2052);
xor XOR2 (N3329, N3302, N747);
not NOT1 (N3330, N3325);
and AND2 (N3331, N3311, N1598);
xor XOR2 (N3332, N3318, N2287);
and AND4 (N3333, N3327, N1501, N1019, N2122);
buf BUF1 (N3334, N3319);
nor NOR3 (N3335, N3330, N1461, N3151);
nor NOR3 (N3336, N3332, N2392, N1851);
and AND2 (N3337, N3336, N2389);
or OR4 (N3338, N3333, N373, N1480, N1970);
buf BUF1 (N3339, N3338);
buf BUF1 (N3340, N3315);
buf BUF1 (N3341, N3334);
or OR3 (N3342, N3285, N2873, N1196);
not NOT1 (N3343, N3328);
buf BUF1 (N3344, N3323);
not NOT1 (N3345, N3331);
nand NAND3 (N3346, N3335, N2384, N808);
nor NOR4 (N3347, N3342, N1572, N3082, N3273);
xor XOR2 (N3348, N3343, N144);
or OR2 (N3349, N3345, N646);
or OR4 (N3350, N3329, N2498, N49, N930);
buf BUF1 (N3351, N3341);
not NOT1 (N3352, N3346);
or OR3 (N3353, N3350, N734, N1983);
nand NAND3 (N3354, N3339, N2025, N1926);
nor NOR4 (N3355, N3351, N2720, N1843, N2453);
or OR2 (N3356, N3340, N3211);
buf BUF1 (N3357, N3348);
buf BUF1 (N3358, N3347);
buf BUF1 (N3359, N3353);
nor NOR4 (N3360, N3349, N3197, N537, N391);
not NOT1 (N3361, N3354);
or OR3 (N3362, N3356, N3191, N14);
nand NAND2 (N3363, N3337, N3358);
xor XOR2 (N3364, N1401, N3304);
or OR3 (N3365, N3363, N444, N1069);
or OR4 (N3366, N3359, N3203, N1018, N52);
nor NOR4 (N3367, N3344, N546, N3090, N144);
nand NAND3 (N3368, N3361, N1606, N3167);
buf BUF1 (N3369, N3352);
nor NOR2 (N3370, N3364, N2626);
and AND4 (N3371, N3366, N3343, N2927, N633);
buf BUF1 (N3372, N3357);
xor XOR2 (N3373, N3369, N618);
nand NAND3 (N3374, N3365, N2019, N1917);
or OR3 (N3375, N3355, N1220, N2323);
xor XOR2 (N3376, N3372, N2856);
or OR4 (N3377, N3376, N1807, N593, N559);
xor XOR2 (N3378, N3367, N1664);
nand NAND2 (N3379, N3360, N31);
xor XOR2 (N3380, N3368, N2678);
not NOT1 (N3381, N3375);
nand NAND4 (N3382, N3380, N1192, N1234, N2828);
or OR2 (N3383, N3379, N2925);
and AND2 (N3384, N3374, N2324);
not NOT1 (N3385, N3378);
buf BUF1 (N3386, N3385);
nand NAND4 (N3387, N3386, N821, N269, N1998);
nand NAND4 (N3388, N3371, N2960, N489, N2067);
and AND2 (N3389, N3388, N2976);
nand NAND3 (N3390, N3370, N2937, N896);
or OR2 (N3391, N3382, N2384);
and AND2 (N3392, N3383, N2471);
nand NAND3 (N3393, N3384, N2190, N1287);
and AND3 (N3394, N3381, N185, N195);
or OR3 (N3395, N3373, N128, N1024);
nand NAND3 (N3396, N3389, N1252, N3089);
buf BUF1 (N3397, N3377);
buf BUF1 (N3398, N3387);
buf BUF1 (N3399, N3392);
nand NAND4 (N3400, N3394, N743, N2855, N3241);
buf BUF1 (N3401, N3398);
nand NAND4 (N3402, N3395, N2737, N287, N2451);
xor XOR2 (N3403, N3391, N2814);
or OR4 (N3404, N3402, N817, N931, N1122);
buf BUF1 (N3405, N3362);
not NOT1 (N3406, N3393);
nand NAND4 (N3407, N3406, N3135, N465, N2382);
nor NOR4 (N3408, N3400, N192, N2983, N2843);
or OR3 (N3409, N3401, N3171, N1269);
not NOT1 (N3410, N3396);
or OR4 (N3411, N3397, N3024, N2478, N2773);
and AND2 (N3412, N3403, N1240);
nor NOR2 (N3413, N3399, N3113);
buf BUF1 (N3414, N3411);
not NOT1 (N3415, N3405);
not NOT1 (N3416, N3408);
buf BUF1 (N3417, N3390);
and AND2 (N3418, N3414, N130);
nand NAND4 (N3419, N3412, N3288, N2788, N1391);
and AND3 (N3420, N3415, N977, N673);
nand NAND3 (N3421, N3416, N1581, N3046);
buf BUF1 (N3422, N3419);
nand NAND2 (N3423, N3404, N42);
nand NAND4 (N3424, N3422, N1647, N2064, N2024);
nand NAND2 (N3425, N3417, N1358);
not NOT1 (N3426, N3409);
nand NAND2 (N3427, N3423, N2971);
not NOT1 (N3428, N3413);
and AND3 (N3429, N3418, N3331, N779);
nor NOR2 (N3430, N3410, N1992);
or OR3 (N3431, N3430, N2413, N3302);
and AND3 (N3432, N3428, N2777, N1921);
and AND4 (N3433, N3420, N1161, N901, N770);
buf BUF1 (N3434, N3425);
and AND2 (N3435, N3431, N2847);
xor XOR2 (N3436, N3421, N15);
not NOT1 (N3437, N3427);
nand NAND3 (N3438, N3424, N1461, N1340);
nand NAND4 (N3439, N3434, N338, N2972, N377);
nand NAND4 (N3440, N3426, N1484, N1382, N2839);
xor XOR2 (N3441, N3429, N915);
xor XOR2 (N3442, N3439, N450);
nor NOR4 (N3443, N3438, N2884, N3152, N1862);
xor XOR2 (N3444, N3437, N804);
buf BUF1 (N3445, N3443);
nand NAND2 (N3446, N3435, N1547);
and AND4 (N3447, N3441, N1032, N553, N1013);
buf BUF1 (N3448, N3445);
xor XOR2 (N3449, N3447, N2539);
nor NOR2 (N3450, N3442, N3210);
buf BUF1 (N3451, N3448);
not NOT1 (N3452, N3446);
nor NOR4 (N3453, N3433, N3099, N372, N31);
xor XOR2 (N3454, N3444, N1258);
and AND4 (N3455, N3451, N679, N2746, N1691);
nor NOR4 (N3456, N3436, N255, N94, N2264);
buf BUF1 (N3457, N3407);
xor XOR2 (N3458, N3454, N2284);
xor XOR2 (N3459, N3449, N929);
buf BUF1 (N3460, N3457);
nor NOR3 (N3461, N3453, N1047, N2466);
nand NAND2 (N3462, N3458, N3324);
buf BUF1 (N3463, N3460);
nor NOR4 (N3464, N3459, N2743, N294, N3127);
or OR3 (N3465, N3462, N2522, N1690);
buf BUF1 (N3466, N3452);
nand NAND2 (N3467, N3450, N2179);
nand NAND4 (N3468, N3432, N2839, N2606, N2244);
buf BUF1 (N3469, N3461);
nor NOR3 (N3470, N3464, N596, N747);
nand NAND3 (N3471, N3455, N291, N397);
nand NAND3 (N3472, N3465, N2868, N1726);
not NOT1 (N3473, N3463);
nand NAND3 (N3474, N3472, N684, N3291);
and AND2 (N3475, N3468, N1279);
xor XOR2 (N3476, N3471, N331);
and AND2 (N3477, N3476, N2503);
nand NAND3 (N3478, N3466, N835, N1474);
or OR3 (N3479, N3470, N2233, N3358);
xor XOR2 (N3480, N3478, N2529);
or OR4 (N3481, N3474, N1698, N3432, N999);
buf BUF1 (N3482, N3477);
or OR4 (N3483, N3481, N1509, N2326, N1205);
or OR4 (N3484, N3469, N362, N2744, N3303);
xor XOR2 (N3485, N3484, N1278);
or OR4 (N3486, N3467, N1255, N2390, N3423);
not NOT1 (N3487, N3486);
nor NOR2 (N3488, N3440, N2720);
buf BUF1 (N3489, N3482);
and AND3 (N3490, N3473, N2728, N134);
and AND3 (N3491, N3487, N2247, N1694);
nor NOR3 (N3492, N3485, N1420, N358);
or OR3 (N3493, N3492, N2198, N1510);
or OR4 (N3494, N3488, N2517, N1939, N2527);
nor NOR4 (N3495, N3489, N299, N3458, N3349);
or OR3 (N3496, N3494, N1036, N2457);
xor XOR2 (N3497, N3479, N3287);
or OR4 (N3498, N3496, N2882, N3343, N3094);
xor XOR2 (N3499, N3475, N869);
xor XOR2 (N3500, N3497, N1103);
buf BUF1 (N3501, N3498);
or OR2 (N3502, N3490, N2643);
nand NAND4 (N3503, N3502, N3171, N1475, N253);
nand NAND2 (N3504, N3501, N3150);
or OR3 (N3505, N3500, N270, N2626);
and AND4 (N3506, N3499, N699, N2176, N2913);
or OR3 (N3507, N3493, N1283, N2267);
or OR3 (N3508, N3456, N814, N3034);
and AND4 (N3509, N3507, N253, N384, N3084);
and AND3 (N3510, N3503, N1320, N3244);
nand NAND4 (N3511, N3505, N1193, N777, N3193);
nor NOR2 (N3512, N3509, N1427);
nand NAND2 (N3513, N3508, N975);
nand NAND4 (N3514, N3511, N1310, N694, N3421);
xor XOR2 (N3515, N3491, N1986);
nand NAND4 (N3516, N3506, N1189, N803, N2969);
nand NAND4 (N3517, N3513, N3100, N1037, N1724);
buf BUF1 (N3518, N3480);
nor NOR3 (N3519, N3483, N1650, N1339);
not NOT1 (N3520, N3517);
xor XOR2 (N3521, N3518, N1500);
or OR2 (N3522, N3520, N2498);
buf BUF1 (N3523, N3519);
not NOT1 (N3524, N3514);
nor NOR2 (N3525, N3524, N2782);
xor XOR2 (N3526, N3522, N2675);
or OR2 (N3527, N3526, N3334);
not NOT1 (N3528, N3512);
or OR2 (N3529, N3527, N138);
and AND3 (N3530, N3516, N1463, N2189);
not NOT1 (N3531, N3530);
not NOT1 (N3532, N3504);
nor NOR4 (N3533, N3523, N553, N186, N1794);
and AND4 (N3534, N3525, N3482, N3411, N2013);
buf BUF1 (N3535, N3510);
or OR3 (N3536, N3521, N1543, N3486);
and AND2 (N3537, N3535, N3370);
buf BUF1 (N3538, N3528);
xor XOR2 (N3539, N3538, N3113);
nand NAND2 (N3540, N3529, N233);
not NOT1 (N3541, N3539);
not NOT1 (N3542, N3533);
or OR2 (N3543, N3515, N3528);
or OR3 (N3544, N3543, N229, N1587);
or OR4 (N3545, N3532, N673, N2207, N1584);
not NOT1 (N3546, N3545);
buf BUF1 (N3547, N3537);
nor NOR4 (N3548, N3531, N1902, N878, N3229);
nor NOR4 (N3549, N3546, N1294, N1050, N336);
or OR2 (N3550, N3536, N1047);
not NOT1 (N3551, N3547);
xor XOR2 (N3552, N3495, N361);
not NOT1 (N3553, N3541);
not NOT1 (N3554, N3550);
and AND3 (N3555, N3540, N957, N2973);
not NOT1 (N3556, N3542);
nor NOR4 (N3557, N3556, N2169, N3151, N3182);
buf BUF1 (N3558, N3555);
not NOT1 (N3559, N3544);
nor NOR2 (N3560, N3553, N1529);
not NOT1 (N3561, N3549);
xor XOR2 (N3562, N3561, N905);
nor NOR3 (N3563, N3552, N1560, N1538);
or OR4 (N3564, N3560, N2607, N1, N235);
or OR2 (N3565, N3559, N128);
not NOT1 (N3566, N3548);
or OR4 (N3567, N3565, N877, N2775, N3520);
or OR4 (N3568, N3557, N941, N725, N2719);
and AND2 (N3569, N3551, N1962);
not NOT1 (N3570, N3568);
and AND3 (N3571, N3558, N3393, N238);
buf BUF1 (N3572, N3554);
nor NOR3 (N3573, N3567, N1679, N284);
buf BUF1 (N3574, N3563);
and AND3 (N3575, N3569, N649, N1939);
and AND3 (N3576, N3573, N3485, N1748);
xor XOR2 (N3577, N3564, N249);
buf BUF1 (N3578, N3575);
or OR4 (N3579, N3574, N3148, N2457, N75);
xor XOR2 (N3580, N3566, N527);
xor XOR2 (N3581, N3570, N3486);
nor NOR2 (N3582, N3571, N3129);
buf BUF1 (N3583, N3572);
xor XOR2 (N3584, N3579, N2053);
nand NAND3 (N3585, N3583, N1086, N973);
nand NAND4 (N3586, N3584, N304, N1518, N2733);
xor XOR2 (N3587, N3578, N3196);
nand NAND3 (N3588, N3587, N2828, N2762);
not NOT1 (N3589, N3580);
not NOT1 (N3590, N3585);
xor XOR2 (N3591, N3588, N2628);
or OR4 (N3592, N3590, N3108, N2430, N2425);
xor XOR2 (N3593, N3576, N1454);
buf BUF1 (N3594, N3589);
xor XOR2 (N3595, N3593, N2195);
nand NAND2 (N3596, N3577, N918);
not NOT1 (N3597, N3594);
and AND3 (N3598, N3591, N2603, N3216);
or OR4 (N3599, N3598, N1899, N3316, N1298);
not NOT1 (N3600, N3596);
xor XOR2 (N3601, N3586, N436);
xor XOR2 (N3602, N3599, N3495);
not NOT1 (N3603, N3600);
xor XOR2 (N3604, N3534, N2448);
nor NOR2 (N3605, N3592, N1685);
and AND4 (N3606, N3602, N1916, N897, N2651);
not NOT1 (N3607, N3603);
buf BUF1 (N3608, N3601);
nand NAND3 (N3609, N3581, N2690, N1140);
xor XOR2 (N3610, N3606, N2946);
or OR3 (N3611, N3597, N2177, N2480);
or OR2 (N3612, N3608, N901);
nor NOR4 (N3613, N3612, N687, N521, N172);
and AND2 (N3614, N3610, N2070);
nor NOR3 (N3615, N3611, N1713, N933);
and AND4 (N3616, N3607, N1275, N808, N3161);
or OR3 (N3617, N3604, N302, N3491);
buf BUF1 (N3618, N3582);
nand NAND2 (N3619, N3614, N2019);
nand NAND2 (N3620, N3616, N1847);
or OR3 (N3621, N3618, N2749, N1665);
nor NOR3 (N3622, N3605, N3273, N699);
or OR2 (N3623, N3617, N2752);
nor NOR2 (N3624, N3615, N704);
or OR3 (N3625, N3609, N1442, N758);
or OR3 (N3626, N3595, N706, N396);
and AND4 (N3627, N3622, N3406, N2481, N1788);
or OR2 (N3628, N3626, N3094);
or OR3 (N3629, N3620, N3131, N1276);
not NOT1 (N3630, N3625);
and AND4 (N3631, N3630, N511, N337, N1458);
nand NAND2 (N3632, N3613, N771);
buf BUF1 (N3633, N3629);
not NOT1 (N3634, N3623);
and AND4 (N3635, N3621, N2539, N1987, N1386);
or OR2 (N3636, N3631, N1906);
nand NAND2 (N3637, N3635, N856);
buf BUF1 (N3638, N3562);
or OR4 (N3639, N3627, N2657, N1118, N2868);
or OR4 (N3640, N3637, N3358, N470, N3010);
xor XOR2 (N3641, N3639, N3269);
not NOT1 (N3642, N3636);
nand NAND2 (N3643, N3642, N2748);
or OR2 (N3644, N3640, N1837);
nand NAND3 (N3645, N3633, N822, N3471);
or OR4 (N3646, N3645, N725, N962, N339);
nor NOR4 (N3647, N3619, N550, N2809, N2992);
or OR3 (N3648, N3624, N3486, N972);
or OR3 (N3649, N3632, N3328, N1035);
buf BUF1 (N3650, N3638);
buf BUF1 (N3651, N3628);
nor NOR4 (N3652, N3650, N121, N2213, N371);
buf BUF1 (N3653, N3643);
nor NOR2 (N3654, N3651, N452);
not NOT1 (N3655, N3646);
not NOT1 (N3656, N3653);
not NOT1 (N3657, N3652);
not NOT1 (N3658, N3648);
not NOT1 (N3659, N3649);
buf BUF1 (N3660, N3634);
and AND4 (N3661, N3654, N2687, N2127, N1321);
nand NAND3 (N3662, N3644, N2409, N3147);
not NOT1 (N3663, N3662);
xor XOR2 (N3664, N3660, N2793);
buf BUF1 (N3665, N3659);
not NOT1 (N3666, N3657);
xor XOR2 (N3667, N3664, N2967);
nand NAND4 (N3668, N3658, N1957, N420, N3606);
buf BUF1 (N3669, N3641);
or OR4 (N3670, N3666, N229, N1553, N1384);
buf BUF1 (N3671, N3669);
not NOT1 (N3672, N3668);
buf BUF1 (N3673, N3656);
nor NOR3 (N3674, N3673, N812, N3376);
nand NAND2 (N3675, N3674, N2079);
and AND4 (N3676, N3663, N3317, N1927, N3055);
nor NOR4 (N3677, N3655, N557, N1873, N3294);
not NOT1 (N3678, N3670);
buf BUF1 (N3679, N3676);
and AND2 (N3680, N3678, N1352);
nand NAND3 (N3681, N3661, N2019, N1048);
or OR4 (N3682, N3679, N774, N3305, N781);
nor NOR4 (N3683, N3682, N2846, N1534, N206);
or OR2 (N3684, N3665, N213);
buf BUF1 (N3685, N3683);
nand NAND4 (N3686, N3675, N492, N16, N2745);
buf BUF1 (N3687, N3647);
or OR2 (N3688, N3684, N1918);
xor XOR2 (N3689, N3672, N1788);
buf BUF1 (N3690, N3677);
xor XOR2 (N3691, N3680, N2014);
xor XOR2 (N3692, N3689, N2087);
not NOT1 (N3693, N3688);
and AND3 (N3694, N3685, N3513, N640);
buf BUF1 (N3695, N3671);
nand NAND2 (N3696, N3693, N2852);
buf BUF1 (N3697, N3691);
xor XOR2 (N3698, N3692, N3093);
or OR3 (N3699, N3681, N2618, N2150);
or OR2 (N3700, N3687, N1420);
or OR3 (N3701, N3698, N1330, N52);
buf BUF1 (N3702, N3667);
and AND2 (N3703, N3699, N251);
and AND2 (N3704, N3702, N1490);
and AND4 (N3705, N3695, N2747, N844, N351);
or OR4 (N3706, N3697, N1997, N2455, N1603);
buf BUF1 (N3707, N3704);
nand NAND4 (N3708, N3703, N400, N2875, N328);
nor NOR3 (N3709, N3707, N3707, N1307);
xor XOR2 (N3710, N3696, N623);
and AND3 (N3711, N3700, N2876, N1304);
and AND2 (N3712, N3708, N125);
nor NOR3 (N3713, N3686, N1991, N878);
nor NOR3 (N3714, N3706, N2407, N100);
buf BUF1 (N3715, N3709);
or OR4 (N3716, N3694, N2035, N3688, N1476);
not NOT1 (N3717, N3716);
buf BUF1 (N3718, N3714);
buf BUF1 (N3719, N3711);
nor NOR4 (N3720, N3719, N847, N3018, N224);
xor XOR2 (N3721, N3710, N2270);
xor XOR2 (N3722, N3713, N3595);
nor NOR4 (N3723, N3721, N907, N631, N168);
and AND2 (N3724, N3712, N2040);
and AND3 (N3725, N3718, N2996, N3715);
nor NOR4 (N3726, N249, N728, N829, N130);
or OR3 (N3727, N3723, N3021, N1198);
and AND2 (N3728, N3690, N1555);
and AND2 (N3729, N3720, N1640);
buf BUF1 (N3730, N3722);
or OR2 (N3731, N3730, N904);
not NOT1 (N3732, N3728);
or OR2 (N3733, N3725, N944);
nor NOR4 (N3734, N3717, N2245, N2311, N3396);
nor NOR4 (N3735, N3726, N3406, N2756, N613);
or OR4 (N3736, N3732, N447, N2071, N662);
nand NAND3 (N3737, N3705, N2983, N1414);
nand NAND4 (N3738, N3729, N1986, N3657, N108);
or OR3 (N3739, N3738, N294, N30);
nand NAND4 (N3740, N3727, N1937, N3365, N405);
xor XOR2 (N3741, N3734, N1795);
not NOT1 (N3742, N3737);
or OR3 (N3743, N3735, N3217, N920);
not NOT1 (N3744, N3731);
not NOT1 (N3745, N3724);
buf BUF1 (N3746, N3745);
or OR2 (N3747, N3740, N2786);
nor NOR4 (N3748, N3736, N3609, N1962, N381);
nor NOR2 (N3749, N3748, N2888);
xor XOR2 (N3750, N3739, N590);
not NOT1 (N3751, N3701);
or OR4 (N3752, N3742, N3524, N280, N2350);
not NOT1 (N3753, N3752);
buf BUF1 (N3754, N3750);
and AND2 (N3755, N3753, N2220);
xor XOR2 (N3756, N3744, N1712);
nor NOR3 (N3757, N3746, N132, N3354);
or OR4 (N3758, N3751, N3313, N2691, N137);
nand NAND3 (N3759, N3741, N2420, N2164);
or OR2 (N3760, N3758, N2359);
xor XOR2 (N3761, N3756, N1957);
buf BUF1 (N3762, N3761);
and AND4 (N3763, N3762, N2576, N3452, N575);
nand NAND3 (N3764, N3754, N188, N281);
buf BUF1 (N3765, N3759);
xor XOR2 (N3766, N3743, N971);
nand NAND3 (N3767, N3749, N1682, N234);
or OR3 (N3768, N3767, N1326, N574);
buf BUF1 (N3769, N3757);
nor NOR3 (N3770, N3766, N2320, N1494);
and AND3 (N3771, N3769, N104, N2202);
not NOT1 (N3772, N3770);
or OR2 (N3773, N3768, N2772);
buf BUF1 (N3774, N3772);
buf BUF1 (N3775, N3771);
and AND2 (N3776, N3763, N3094);
nor NOR2 (N3777, N3775, N2865);
not NOT1 (N3778, N3755);
nand NAND4 (N3779, N3774, N3039, N1431, N275);
nand NAND2 (N3780, N3764, N2950);
nor NOR3 (N3781, N3773, N353, N666);
xor XOR2 (N3782, N3779, N1661);
nor NOR3 (N3783, N3776, N195, N189);
buf BUF1 (N3784, N3778);
or OR4 (N3785, N3782, N1365, N1203, N2907);
and AND3 (N3786, N3785, N1302, N1794);
nand NAND2 (N3787, N3783, N1103);
nand NAND4 (N3788, N3786, N263, N2261, N2723);
not NOT1 (N3789, N3777);
buf BUF1 (N3790, N3788);
nand NAND2 (N3791, N3760, N341);
not NOT1 (N3792, N3790);
xor XOR2 (N3793, N3791, N2382);
nand NAND4 (N3794, N3733, N1272, N903, N2237);
nand NAND3 (N3795, N3765, N938, N2122);
xor XOR2 (N3796, N3781, N1437);
nand NAND3 (N3797, N3794, N3046, N3070);
nor NOR3 (N3798, N3796, N2801, N1634);
nor NOR3 (N3799, N3787, N3337, N2783);
nand NAND2 (N3800, N3780, N2941);
and AND2 (N3801, N3798, N1536);
or OR3 (N3802, N3784, N3068, N2716);
xor XOR2 (N3803, N3792, N3013);
or OR2 (N3804, N3799, N2281);
not NOT1 (N3805, N3800);
xor XOR2 (N3806, N3801, N45);
nand NAND2 (N3807, N3806, N2518);
or OR3 (N3808, N3805, N2391, N3494);
buf BUF1 (N3809, N3793);
and AND2 (N3810, N3803, N665);
nand NAND4 (N3811, N3789, N3141, N1206, N1634);
and AND2 (N3812, N3747, N3076);
not NOT1 (N3813, N3807);
buf BUF1 (N3814, N3811);
xor XOR2 (N3815, N3813, N639);
or OR3 (N3816, N3814, N2398, N384);
nor NOR2 (N3817, N3797, N1798);
xor XOR2 (N3818, N3809, N337);
xor XOR2 (N3819, N3804, N247);
buf BUF1 (N3820, N3819);
nand NAND2 (N3821, N3818, N3443);
or OR4 (N3822, N3812, N2290, N3720, N1000);
or OR2 (N3823, N3795, N2617);
not NOT1 (N3824, N3810);
nor NOR2 (N3825, N3816, N1670);
buf BUF1 (N3826, N3815);
or OR3 (N3827, N3821, N1634, N965);
nand NAND4 (N3828, N3808, N1665, N3365, N1805);
nor NOR2 (N3829, N3820, N2111);
not NOT1 (N3830, N3825);
buf BUF1 (N3831, N3823);
nand NAND2 (N3832, N3802, N3792);
xor XOR2 (N3833, N3822, N1748);
or OR3 (N3834, N3817, N478, N2790);
nor NOR2 (N3835, N3828, N623);
nor NOR2 (N3836, N3832, N3609);
or OR2 (N3837, N3824, N37);
buf BUF1 (N3838, N3837);
and AND2 (N3839, N3838, N2027);
nor NOR2 (N3840, N3834, N1923);
not NOT1 (N3841, N3831);
nor NOR3 (N3842, N3841, N2637, N2873);
xor XOR2 (N3843, N3836, N1710);
and AND3 (N3844, N3826, N2964, N2916);
xor XOR2 (N3845, N3827, N375);
nor NOR4 (N3846, N3839, N2560, N2370, N3061);
buf BUF1 (N3847, N3840);
xor XOR2 (N3848, N3829, N1620);
or OR2 (N3849, N3835, N3820);
nor NOR4 (N3850, N3833, N1683, N1481, N769);
nor NOR2 (N3851, N3849, N2550);
or OR4 (N3852, N3844, N3169, N3070, N1993);
xor XOR2 (N3853, N3830, N1896);
not NOT1 (N3854, N3843);
not NOT1 (N3855, N3845);
and AND4 (N3856, N3847, N3005, N1536, N1095);
nand NAND3 (N3857, N3854, N2974, N949);
nor NOR3 (N3858, N3848, N1751, N349);
nor NOR2 (N3859, N3852, N3536);
or OR2 (N3860, N3853, N2060);
nor NOR3 (N3861, N3846, N896, N756);
xor XOR2 (N3862, N3858, N3714);
xor XOR2 (N3863, N3857, N1271);
nor NOR4 (N3864, N3861, N3456, N2803, N3156);
xor XOR2 (N3865, N3851, N3589);
xor XOR2 (N3866, N3856, N3013);
not NOT1 (N3867, N3860);
or OR2 (N3868, N3842, N2063);
xor XOR2 (N3869, N3855, N2255);
nand NAND2 (N3870, N3862, N1010);
nor NOR2 (N3871, N3866, N1105);
buf BUF1 (N3872, N3864);
nand NAND4 (N3873, N3872, N2471, N1802, N2268);
xor XOR2 (N3874, N3867, N1851);
nor NOR3 (N3875, N3873, N1135, N2971);
or OR4 (N3876, N3869, N1343, N35, N3391);
xor XOR2 (N3877, N3874, N1597);
and AND2 (N3878, N3863, N2586);
not NOT1 (N3879, N3878);
xor XOR2 (N3880, N3865, N1617);
nand NAND4 (N3881, N3879, N1731, N1659, N3470);
and AND3 (N3882, N3868, N345, N930);
or OR2 (N3883, N3882, N3865);
xor XOR2 (N3884, N3850, N3194);
nor NOR2 (N3885, N3884, N708);
or OR2 (N3886, N3871, N986);
buf BUF1 (N3887, N3870);
and AND2 (N3888, N3885, N2132);
not NOT1 (N3889, N3880);
or OR2 (N3890, N3883, N3254);
buf BUF1 (N3891, N3887);
and AND4 (N3892, N3888, N1348, N3500, N2015);
buf BUF1 (N3893, N3892);
and AND2 (N3894, N3889, N3488);
not NOT1 (N3895, N3890);
nand NAND2 (N3896, N3894, N1678);
nand NAND4 (N3897, N3859, N310, N1875, N3074);
nor NOR2 (N3898, N3881, N2468);
or OR4 (N3899, N3898, N2720, N2672, N2496);
and AND3 (N3900, N3876, N1668, N2900);
nor NOR2 (N3901, N3877, N3772);
not NOT1 (N3902, N3899);
nor NOR4 (N3903, N3896, N3698, N1875, N1500);
xor XOR2 (N3904, N3875, N1680);
xor XOR2 (N3905, N3902, N2936);
not NOT1 (N3906, N3900);
and AND3 (N3907, N3901, N1965, N63);
not NOT1 (N3908, N3903);
buf BUF1 (N3909, N3886);
xor XOR2 (N3910, N3891, N3753);
xor XOR2 (N3911, N3909, N2891);
xor XOR2 (N3912, N3897, N436);
not NOT1 (N3913, N3908);
buf BUF1 (N3914, N3905);
not NOT1 (N3915, N3912);
or OR4 (N3916, N3907, N2168, N1161, N2338);
nor NOR4 (N3917, N3895, N1062, N482, N811);
buf BUF1 (N3918, N3917);
or OR4 (N3919, N3910, N2537, N56, N1544);
buf BUF1 (N3920, N3893);
nor NOR2 (N3921, N3920, N2070);
nand NAND3 (N3922, N3919, N21, N3003);
and AND2 (N3923, N3914, N2686);
or OR4 (N3924, N3904, N1637, N990, N2994);
xor XOR2 (N3925, N3918, N3881);
and AND3 (N3926, N3906, N698, N1760);
and AND2 (N3927, N3925, N266);
or OR4 (N3928, N3911, N444, N3086, N1242);
buf BUF1 (N3929, N3923);
nor NOR4 (N3930, N3921, N3352, N695, N3518);
buf BUF1 (N3931, N3922);
and AND2 (N3932, N3926, N3091);
not NOT1 (N3933, N3932);
nor NOR2 (N3934, N3931, N691);
not NOT1 (N3935, N3928);
nand NAND2 (N3936, N3916, N3450);
and AND3 (N3937, N3933, N355, N235);
nand NAND3 (N3938, N3913, N1369, N2962);
xor XOR2 (N3939, N3930, N3068);
not NOT1 (N3940, N3935);
nand NAND3 (N3941, N3937, N300, N1869);
or OR2 (N3942, N3936, N1651);
and AND3 (N3943, N3940, N2195, N1315);
nor NOR2 (N3944, N3941, N1106);
or OR2 (N3945, N3939, N3007);
or OR4 (N3946, N3927, N3605, N2054, N3245);
not NOT1 (N3947, N3938);
or OR2 (N3948, N3942, N415);
xor XOR2 (N3949, N3915, N373);
xor XOR2 (N3950, N3948, N2717);
nand NAND4 (N3951, N3946, N1847, N1573, N479);
not NOT1 (N3952, N3944);
or OR4 (N3953, N3949, N1620, N3341, N441);
nor NOR3 (N3954, N3952, N304, N2547);
or OR2 (N3955, N3951, N13);
nand NAND2 (N3956, N3947, N1072);
nor NOR2 (N3957, N3945, N3322);
not NOT1 (N3958, N3924);
nor NOR3 (N3959, N3953, N1455, N341);
nand NAND3 (N3960, N3959, N3805, N2890);
xor XOR2 (N3961, N3954, N3162);
nor NOR3 (N3962, N3960, N3592, N1769);
and AND2 (N3963, N3958, N699);
and AND2 (N3964, N3950, N1049);
buf BUF1 (N3965, N3934);
xor XOR2 (N3966, N3955, N1863);
buf BUF1 (N3967, N3965);
nand NAND2 (N3968, N3956, N2921);
or OR4 (N3969, N3943, N3007, N2703, N2925);
buf BUF1 (N3970, N3929);
and AND4 (N3971, N3964, N3423, N3737, N3538);
or OR4 (N3972, N3971, N2490, N2393, N128);
nor NOR4 (N3973, N3957, N3168, N408, N3116);
or OR2 (N3974, N3973, N1666);
nand NAND2 (N3975, N3970, N294);
buf BUF1 (N3976, N3975);
or OR3 (N3977, N3966, N193, N3488);
buf BUF1 (N3978, N3968);
nor NOR3 (N3979, N3977, N2468, N3504);
nand NAND4 (N3980, N3972, N322, N345, N1135);
not NOT1 (N3981, N3963);
nor NOR4 (N3982, N3969, N2731, N795, N564);
xor XOR2 (N3983, N3981, N135);
buf BUF1 (N3984, N3978);
not NOT1 (N3985, N3961);
and AND3 (N3986, N3982, N1077, N612);
buf BUF1 (N3987, N3980);
and AND2 (N3988, N3974, N1271);
and AND2 (N3989, N3976, N3577);
not NOT1 (N3990, N3984);
nor NOR2 (N3991, N3962, N417);
xor XOR2 (N3992, N3989, N2360);
not NOT1 (N3993, N3990);
nor NOR4 (N3994, N3985, N1095, N55, N3805);
nor NOR3 (N3995, N3988, N2536, N1063);
xor XOR2 (N3996, N3986, N1051);
or OR3 (N3997, N3992, N942, N2522);
xor XOR2 (N3998, N3979, N2125);
buf BUF1 (N3999, N3967);
nand NAND4 (N4000, N3999, N348, N3863, N599);
not NOT1 (N4001, N3996);
or OR4 (N4002, N3998, N1912, N126, N2144);
not NOT1 (N4003, N3993);
nor NOR2 (N4004, N3997, N3237);
nor NOR4 (N4005, N3995, N3900, N453, N1199);
nor NOR3 (N4006, N4004, N924, N158);
buf BUF1 (N4007, N4000);
not NOT1 (N4008, N3983);
nor NOR3 (N4009, N3991, N294, N2955);
xor XOR2 (N4010, N4009, N345);
nand NAND2 (N4011, N4007, N3130);
nand NAND3 (N4012, N4010, N2048, N296);
nand NAND2 (N4013, N4003, N3262);
endmodule