// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N706,N704,N707,N702,N699,N692,N697,N693,N703,N710;

not NOT1 (N11, N10);
not NOT1 (N12, N6);
or OR3 (N13, N7, N7, N4);
xor XOR2 (N14, N10, N8);
nor NOR2 (N15, N13, N10);
buf BUF1 (N16, N15);
nor NOR3 (N17, N12, N14, N5);
and AND3 (N18, N15, N16, N9);
nand NAND3 (N19, N18, N14, N13);
xor XOR2 (N20, N9, N9);
nand NAND2 (N21, N19, N14);
and AND2 (N22, N4, N11);
nand NAND2 (N23, N6, N14);
or OR4 (N24, N17, N2, N6, N5);
nand NAND2 (N25, N14, N10);
not NOT1 (N26, N15);
and AND2 (N27, N2, N10);
nand NAND4 (N28, N15, N14, N1, N8);
nand NAND4 (N29, N5, N11, N13, N8);
nand NAND4 (N30, N29, N19, N6, N20);
xor XOR2 (N31, N16, N16);
xor XOR2 (N32, N27, N18);
or OR2 (N33, N30, N21);
and AND2 (N34, N32, N8);
nand NAND3 (N35, N5, N26, N8);
and AND2 (N36, N29, N21);
and AND2 (N37, N23, N10);
or OR3 (N38, N36, N23, N5);
nor NOR3 (N39, N28, N10, N17);
buf BUF1 (N40, N31);
nand NAND2 (N41, N24, N31);
or OR3 (N42, N37, N20, N36);
and AND2 (N43, N42, N10);
xor XOR2 (N44, N43, N12);
buf BUF1 (N45, N35);
nor NOR2 (N46, N41, N8);
and AND4 (N47, N38, N17, N30, N26);
and AND2 (N48, N39, N14);
buf BUF1 (N49, N47);
and AND4 (N50, N45, N47, N10, N29);
xor XOR2 (N51, N48, N39);
and AND4 (N52, N44, N40, N44, N48);
nand NAND3 (N53, N33, N37, N38);
nor NOR4 (N54, N47, N18, N36, N29);
or OR4 (N55, N25, N50, N20, N49);
nand NAND4 (N56, N49, N29, N12, N22);
nand NAND3 (N57, N6, N25, N38);
xor XOR2 (N58, N50, N35);
nand NAND2 (N59, N55, N37);
nor NOR3 (N60, N59, N10, N44);
not NOT1 (N61, N52);
buf BUF1 (N62, N60);
nor NOR4 (N63, N58, N14, N60, N29);
buf BUF1 (N64, N62);
or OR3 (N65, N57, N56, N41);
not NOT1 (N66, N37);
xor XOR2 (N67, N34, N27);
buf BUF1 (N68, N65);
xor XOR2 (N69, N63, N57);
nor NOR3 (N70, N64, N3, N50);
xor XOR2 (N71, N66, N17);
nor NOR3 (N72, N54, N54, N63);
not NOT1 (N73, N67);
nor NOR2 (N74, N69, N51);
buf BUF1 (N75, N26);
not NOT1 (N76, N53);
xor XOR2 (N77, N76, N14);
nand NAND3 (N78, N46, N38, N9);
not NOT1 (N79, N71);
nor NOR2 (N80, N75, N53);
buf BUF1 (N81, N80);
nand NAND2 (N82, N73, N6);
xor XOR2 (N83, N70, N19);
or OR3 (N84, N78, N20, N55);
xor XOR2 (N85, N79, N74);
xor XOR2 (N86, N42, N17);
xor XOR2 (N87, N77, N80);
nor NOR2 (N88, N85, N55);
buf BUF1 (N89, N86);
or OR2 (N90, N83, N79);
xor XOR2 (N91, N90, N21);
buf BUF1 (N92, N89);
xor XOR2 (N93, N61, N17);
and AND2 (N94, N87, N53);
or OR2 (N95, N82, N40);
buf BUF1 (N96, N95);
and AND4 (N97, N93, N51, N82, N76);
nand NAND3 (N98, N84, N6, N53);
buf BUF1 (N99, N96);
nand NAND4 (N100, N88, N19, N94, N84);
or OR4 (N101, N44, N18, N81, N90);
nor NOR4 (N102, N62, N6, N27, N22);
or OR2 (N103, N92, N43);
nand NAND3 (N104, N100, N55, N25);
buf BUF1 (N105, N99);
nand NAND4 (N106, N101, N26, N99, N41);
or OR4 (N107, N91, N5, N93, N87);
not NOT1 (N108, N103);
and AND4 (N109, N68, N97, N9, N14);
not NOT1 (N110, N85);
not NOT1 (N111, N102);
not NOT1 (N112, N107);
nor NOR4 (N113, N108, N75, N70, N26);
and AND2 (N114, N111, N39);
nor NOR2 (N115, N109, N105);
buf BUF1 (N116, N1);
xor XOR2 (N117, N104, N45);
or OR3 (N118, N98, N30, N68);
and AND3 (N119, N118, N62, N75);
not NOT1 (N120, N119);
nor NOR4 (N121, N112, N119, N29, N48);
nor NOR2 (N122, N117, N48);
buf BUF1 (N123, N72);
nand NAND2 (N124, N121, N71);
nor NOR4 (N125, N115, N43, N31, N88);
buf BUF1 (N126, N106);
nor NOR3 (N127, N114, N13, N91);
xor XOR2 (N128, N123, N43);
nand NAND2 (N129, N110, N9);
xor XOR2 (N130, N116, N102);
and AND4 (N131, N125, N67, N99, N92);
not NOT1 (N132, N113);
buf BUF1 (N133, N120);
not NOT1 (N134, N127);
nand NAND2 (N135, N122, N101);
nor NOR3 (N136, N132, N35, N67);
nor NOR2 (N137, N130, N126);
xor XOR2 (N138, N75, N78);
not NOT1 (N139, N137);
not NOT1 (N140, N133);
or OR4 (N141, N128, N121, N78, N110);
nand NAND2 (N142, N138, N63);
nand NAND4 (N143, N142, N12, N89, N130);
not NOT1 (N144, N139);
or OR3 (N145, N136, N61, N124);
and AND3 (N146, N63, N117, N23);
buf BUF1 (N147, N145);
buf BUF1 (N148, N134);
nand NAND3 (N149, N129, N86, N49);
buf BUF1 (N150, N148);
and AND2 (N151, N150, N36);
buf BUF1 (N152, N131);
or OR3 (N153, N143, N107, N31);
nor NOR4 (N154, N141, N73, N107, N100);
and AND2 (N155, N152, N144);
buf BUF1 (N156, N99);
not NOT1 (N157, N153);
and AND2 (N158, N146, N119);
nor NOR4 (N159, N157, N132, N146, N86);
or OR2 (N160, N149, N132);
nand NAND4 (N161, N159, N91, N22, N54);
not NOT1 (N162, N156);
or OR4 (N163, N135, N131, N117, N144);
nor NOR4 (N164, N161, N85, N159, N33);
not NOT1 (N165, N155);
nor NOR4 (N166, N160, N8, N135, N91);
not NOT1 (N167, N140);
nor NOR3 (N168, N147, N14, N136);
or OR2 (N169, N167, N115);
not NOT1 (N170, N168);
nand NAND3 (N171, N164, N111, N170);
nand NAND3 (N172, N22, N128, N62);
nand NAND2 (N173, N151, N43);
not NOT1 (N174, N173);
nand NAND4 (N175, N163, N86, N21, N116);
xor XOR2 (N176, N162, N122);
or OR2 (N177, N171, N19);
nor NOR4 (N178, N166, N22, N134, N9);
or OR4 (N179, N165, N62, N19, N138);
nand NAND3 (N180, N158, N116, N127);
xor XOR2 (N181, N175, N71);
not NOT1 (N182, N172);
nand NAND2 (N183, N181, N128);
not NOT1 (N184, N169);
buf BUF1 (N185, N182);
nand NAND4 (N186, N174, N136, N164, N45);
and AND2 (N187, N179, N122);
or OR3 (N188, N185, N102, N33);
nand NAND3 (N189, N183, N169, N5);
or OR3 (N190, N176, N108, N44);
and AND2 (N191, N189, N19);
and AND3 (N192, N178, N147, N132);
buf BUF1 (N193, N180);
not NOT1 (N194, N193);
xor XOR2 (N195, N188, N95);
and AND4 (N196, N195, N174, N20, N183);
or OR3 (N197, N187, N17, N125);
not NOT1 (N198, N194);
not NOT1 (N199, N177);
nand NAND3 (N200, N186, N64, N103);
not NOT1 (N201, N184);
buf BUF1 (N202, N197);
nor NOR2 (N203, N202, N77);
not NOT1 (N204, N198);
nand NAND2 (N205, N199, N197);
xor XOR2 (N206, N205, N121);
or OR3 (N207, N192, N141, N76);
nand NAND4 (N208, N206, N165, N46, N84);
nand NAND2 (N209, N208, N70);
nand NAND4 (N210, N196, N161, N135, N72);
not NOT1 (N211, N210);
nand NAND2 (N212, N154, N138);
not NOT1 (N213, N209);
xor XOR2 (N214, N191, N125);
not NOT1 (N215, N203);
buf BUF1 (N216, N204);
nand NAND4 (N217, N215, N33, N125, N3);
nor NOR2 (N218, N211, N213);
not NOT1 (N219, N35);
buf BUF1 (N220, N190);
nand NAND4 (N221, N201, N187, N79, N192);
not NOT1 (N222, N216);
buf BUF1 (N223, N217);
nor NOR3 (N224, N207, N165, N65);
xor XOR2 (N225, N222, N142);
buf BUF1 (N226, N219);
nand NAND4 (N227, N221, N123, N3, N165);
nand NAND2 (N228, N218, N10);
nand NAND2 (N229, N226, N178);
and AND4 (N230, N229, N174, N53, N177);
nor NOR2 (N231, N224, N71);
nor NOR3 (N232, N230, N77, N152);
or OR4 (N233, N220, N40, N106, N190);
and AND3 (N234, N227, N195, N146);
not NOT1 (N235, N223);
and AND4 (N236, N200, N6, N141, N38);
xor XOR2 (N237, N228, N160);
not NOT1 (N238, N232);
nand NAND2 (N239, N236, N191);
nand NAND3 (N240, N238, N63, N160);
nor NOR3 (N241, N239, N195, N55);
and AND2 (N242, N233, N158);
or OR4 (N243, N234, N60, N182, N142);
or OR4 (N244, N241, N172, N164, N227);
xor XOR2 (N245, N237, N11);
or OR4 (N246, N243, N11, N106, N147);
xor XOR2 (N247, N245, N1);
nand NAND3 (N248, N214, N61, N7);
not NOT1 (N249, N225);
or OR4 (N250, N212, N222, N82, N143);
nand NAND3 (N251, N240, N170, N12);
nand NAND4 (N252, N251, N62, N125, N229);
and AND2 (N253, N250, N245);
and AND3 (N254, N249, N212, N80);
nand NAND2 (N255, N248, N120);
or OR4 (N256, N247, N248, N11, N222);
nand NAND4 (N257, N244, N207, N196, N181);
nor NOR4 (N258, N254, N250, N175, N161);
nor NOR2 (N259, N258, N137);
nand NAND2 (N260, N253, N220);
not NOT1 (N261, N231);
nor NOR3 (N262, N261, N141, N218);
nand NAND3 (N263, N262, N235, N65);
not NOT1 (N264, N232);
xor XOR2 (N265, N259, N223);
nor NOR4 (N266, N256, N99, N171, N180);
or OR4 (N267, N264, N5, N127, N144);
nand NAND4 (N268, N265, N253, N194, N32);
or OR3 (N269, N246, N164, N122);
nor NOR2 (N270, N252, N22);
nand NAND3 (N271, N270, N196, N250);
nor NOR3 (N272, N263, N75, N211);
nor NOR4 (N273, N271, N169, N29, N58);
nor NOR3 (N274, N268, N227, N187);
buf BUF1 (N275, N272);
buf BUF1 (N276, N273);
and AND3 (N277, N267, N49, N101);
buf BUF1 (N278, N276);
and AND2 (N279, N269, N134);
nand NAND4 (N280, N279, N279, N274, N220);
not NOT1 (N281, N100);
nand NAND3 (N282, N281, N30, N240);
and AND2 (N283, N266, N192);
not NOT1 (N284, N277);
or OR2 (N285, N260, N21);
nand NAND4 (N286, N255, N17, N250, N279);
nand NAND4 (N287, N280, N195, N225, N38);
nand NAND3 (N288, N285, N228, N58);
buf BUF1 (N289, N287);
or OR4 (N290, N288, N191, N30, N32);
and AND3 (N291, N275, N143, N95);
xor XOR2 (N292, N283, N35);
nor NOR4 (N293, N291, N123, N103, N235);
nand NAND3 (N294, N257, N236, N274);
and AND2 (N295, N284, N64);
xor XOR2 (N296, N295, N8);
or OR4 (N297, N286, N138, N27, N56);
not NOT1 (N298, N282);
or OR2 (N299, N297, N115);
nand NAND3 (N300, N293, N215, N145);
and AND3 (N301, N292, N159, N111);
buf BUF1 (N302, N296);
xor XOR2 (N303, N298, N155);
and AND3 (N304, N299, N220, N26);
and AND4 (N305, N301, N175, N235, N244);
nand NAND3 (N306, N305, N207, N120);
not NOT1 (N307, N300);
not NOT1 (N308, N306);
or OR3 (N309, N290, N34, N11);
and AND2 (N310, N308, N184);
not NOT1 (N311, N242);
buf BUF1 (N312, N303);
or OR4 (N313, N309, N22, N33, N179);
nand NAND2 (N314, N312, N8);
nand NAND4 (N315, N307, N141, N312, N56);
and AND4 (N316, N311, N173, N256, N295);
not NOT1 (N317, N278);
buf BUF1 (N318, N304);
nand NAND3 (N319, N294, N175, N154);
buf BUF1 (N320, N318);
buf BUF1 (N321, N320);
not NOT1 (N322, N302);
nand NAND2 (N323, N313, N16);
and AND2 (N324, N319, N6);
nand NAND2 (N325, N322, N163);
or OR2 (N326, N315, N96);
nand NAND2 (N327, N314, N286);
and AND3 (N328, N327, N306, N198);
buf BUF1 (N329, N323);
nand NAND2 (N330, N328, N222);
and AND4 (N331, N317, N323, N60, N233);
buf BUF1 (N332, N330);
buf BUF1 (N333, N332);
nand NAND4 (N334, N316, N227, N197, N225);
and AND3 (N335, N326, N137, N31);
and AND3 (N336, N310, N180, N256);
nor NOR2 (N337, N334, N297);
nand NAND4 (N338, N333, N182, N211, N136);
not NOT1 (N339, N289);
or OR3 (N340, N325, N272, N92);
nand NAND2 (N341, N329, N65);
buf BUF1 (N342, N341);
buf BUF1 (N343, N342);
xor XOR2 (N344, N340, N225);
xor XOR2 (N345, N338, N14);
buf BUF1 (N346, N321);
xor XOR2 (N347, N331, N321);
nor NOR4 (N348, N337, N269, N283, N53);
xor XOR2 (N349, N324, N105);
nor NOR3 (N350, N344, N202, N131);
nand NAND4 (N351, N348, N160, N122, N3);
nor NOR4 (N352, N351, N40, N198, N86);
or OR3 (N353, N335, N16, N178);
and AND4 (N354, N343, N151, N207, N350);
nor NOR2 (N355, N6, N312);
nor NOR4 (N356, N339, N213, N66, N136);
not NOT1 (N357, N347);
buf BUF1 (N358, N353);
nor NOR2 (N359, N346, N215);
buf BUF1 (N360, N345);
nor NOR3 (N361, N355, N285, N170);
not NOT1 (N362, N357);
and AND2 (N363, N360, N213);
xor XOR2 (N364, N336, N325);
and AND3 (N365, N363, N60, N233);
or OR4 (N366, N359, N302, N149, N197);
nand NAND3 (N367, N354, N98, N241);
buf BUF1 (N368, N362);
and AND2 (N369, N368, N107);
and AND4 (N370, N369, N312, N18, N190);
nor NOR2 (N371, N349, N21);
nand NAND3 (N372, N366, N364, N237);
and AND3 (N373, N53, N137, N162);
nor NOR4 (N374, N372, N162, N277, N295);
and AND3 (N375, N352, N334, N14);
buf BUF1 (N376, N373);
nor NOR3 (N377, N375, N345, N279);
not NOT1 (N378, N361);
and AND4 (N379, N367, N85, N259, N34);
buf BUF1 (N380, N371);
not NOT1 (N381, N370);
and AND4 (N382, N356, N296, N119, N39);
nand NAND2 (N383, N379, N321);
buf BUF1 (N384, N380);
nand NAND4 (N385, N383, N36, N201, N373);
and AND4 (N386, N376, N154, N184, N136);
and AND3 (N387, N358, N57, N86);
not NOT1 (N388, N377);
buf BUF1 (N389, N378);
and AND4 (N390, N374, N366, N99, N63);
and AND3 (N391, N384, N322, N375);
nor NOR3 (N392, N381, N10, N188);
and AND2 (N393, N392, N352);
and AND3 (N394, N388, N100, N80);
and AND4 (N395, N391, N46, N158, N252);
not NOT1 (N396, N390);
xor XOR2 (N397, N387, N113);
nor NOR2 (N398, N394, N22);
nor NOR2 (N399, N389, N85);
and AND4 (N400, N397, N74, N230, N268);
or OR3 (N401, N393, N118, N380);
and AND4 (N402, N401, N111, N11, N276);
and AND4 (N403, N385, N180, N181, N107);
not NOT1 (N404, N403);
buf BUF1 (N405, N402);
or OR4 (N406, N365, N70, N393, N149);
buf BUF1 (N407, N386);
xor XOR2 (N408, N398, N261);
xor XOR2 (N409, N405, N262);
nand NAND3 (N410, N409, N249, N328);
nor NOR3 (N411, N408, N45, N236);
not NOT1 (N412, N382);
and AND4 (N413, N407, N282, N174, N227);
buf BUF1 (N414, N400);
or OR3 (N415, N410, N5, N149);
or OR4 (N416, N399, N181, N91, N3);
or OR4 (N417, N413, N97, N412, N88);
nand NAND2 (N418, N219, N102);
nand NAND2 (N419, N416, N340);
buf BUF1 (N420, N396);
or OR4 (N421, N420, N266, N74, N195);
not NOT1 (N422, N417);
nand NAND4 (N423, N419, N186, N420, N290);
or OR3 (N424, N421, N310, N281);
xor XOR2 (N425, N395, N203);
nand NAND4 (N426, N414, N329, N176, N274);
and AND4 (N427, N422, N248, N316, N135);
not NOT1 (N428, N411);
not NOT1 (N429, N427);
nand NAND4 (N430, N424, N41, N134, N322);
nand NAND4 (N431, N418, N162, N126, N322);
buf BUF1 (N432, N404);
and AND3 (N433, N431, N375, N165);
nor NOR2 (N434, N428, N287);
not NOT1 (N435, N425);
not NOT1 (N436, N432);
nand NAND2 (N437, N433, N223);
and AND2 (N438, N437, N360);
buf BUF1 (N439, N406);
nor NOR2 (N440, N423, N116);
not NOT1 (N441, N426);
xor XOR2 (N442, N439, N187);
xor XOR2 (N443, N440, N359);
nand NAND4 (N444, N438, N296, N108, N113);
and AND4 (N445, N442, N119, N218, N338);
and AND2 (N446, N429, N273);
xor XOR2 (N447, N436, N230);
xor XOR2 (N448, N430, N296);
buf BUF1 (N449, N446);
xor XOR2 (N450, N445, N362);
or OR3 (N451, N447, N135, N313);
nand NAND4 (N452, N435, N97, N368, N407);
not NOT1 (N453, N448);
nand NAND3 (N454, N441, N430, N417);
nor NOR4 (N455, N443, N405, N216, N263);
or OR3 (N456, N455, N125, N442);
nand NAND3 (N457, N444, N150, N426);
or OR3 (N458, N454, N342, N438);
nor NOR2 (N459, N449, N452);
nor NOR4 (N460, N82, N372, N179, N161);
not NOT1 (N461, N456);
nor NOR3 (N462, N457, N167, N339);
not NOT1 (N463, N462);
or OR3 (N464, N453, N85, N295);
xor XOR2 (N465, N459, N157);
xor XOR2 (N466, N463, N300);
buf BUF1 (N467, N466);
xor XOR2 (N468, N460, N215);
or OR2 (N469, N415, N457);
xor XOR2 (N470, N450, N438);
nand NAND4 (N471, N467, N153, N182, N342);
and AND3 (N472, N461, N155, N464);
or OR4 (N473, N118, N14, N23, N203);
or OR2 (N474, N469, N56);
nor NOR4 (N475, N470, N297, N389, N270);
not NOT1 (N476, N434);
and AND4 (N477, N475, N56, N232, N107);
nor NOR4 (N478, N472, N80, N84, N247);
nor NOR3 (N479, N478, N432, N24);
xor XOR2 (N480, N468, N463);
buf BUF1 (N481, N474);
not NOT1 (N482, N481);
nor NOR3 (N483, N479, N149, N61);
not NOT1 (N484, N471);
and AND3 (N485, N473, N235, N224);
nor NOR2 (N486, N458, N344);
xor XOR2 (N487, N480, N462);
or OR3 (N488, N477, N201, N472);
buf BUF1 (N489, N485);
and AND4 (N490, N451, N158, N452, N194);
buf BUF1 (N491, N488);
xor XOR2 (N492, N489, N140);
or OR3 (N493, N483, N338, N298);
and AND2 (N494, N486, N272);
nand NAND2 (N495, N482, N102);
and AND3 (N496, N465, N182, N482);
and AND2 (N497, N493, N471);
buf BUF1 (N498, N476);
nand NAND2 (N499, N497, N453);
xor XOR2 (N500, N492, N9);
and AND4 (N501, N484, N213, N47, N400);
not NOT1 (N502, N487);
nor NOR4 (N503, N496, N428, N136, N32);
and AND3 (N504, N503, N54, N54);
or OR2 (N505, N502, N125);
nor NOR2 (N506, N498, N28);
not NOT1 (N507, N505);
nand NAND4 (N508, N494, N4, N234, N270);
nor NOR3 (N509, N499, N233, N197);
or OR2 (N510, N500, N206);
nor NOR4 (N511, N495, N359, N116, N173);
nand NAND2 (N512, N508, N245);
or OR2 (N513, N507, N103);
xor XOR2 (N514, N509, N235);
nand NAND2 (N515, N512, N2);
not NOT1 (N516, N510);
or OR2 (N517, N516, N395);
not NOT1 (N518, N515);
buf BUF1 (N519, N514);
and AND3 (N520, N517, N95, N10);
buf BUF1 (N521, N490);
or OR4 (N522, N513, N6, N13, N45);
or OR3 (N523, N521, N326, N289);
buf BUF1 (N524, N491);
not NOT1 (N525, N518);
and AND3 (N526, N511, N263, N510);
and AND2 (N527, N506, N92);
nand NAND2 (N528, N524, N434);
nor NOR3 (N529, N504, N165, N394);
nand NAND2 (N530, N529, N120);
not NOT1 (N531, N522);
xor XOR2 (N532, N525, N334);
xor XOR2 (N533, N519, N148);
and AND2 (N534, N531, N382);
nand NAND3 (N535, N532, N5, N455);
xor XOR2 (N536, N501, N254);
not NOT1 (N537, N535);
nand NAND2 (N538, N536, N116);
or OR3 (N539, N530, N68, N269);
buf BUF1 (N540, N539);
buf BUF1 (N541, N527);
or OR3 (N542, N540, N283, N144);
not NOT1 (N543, N526);
buf BUF1 (N544, N542);
and AND3 (N545, N537, N355, N300);
not NOT1 (N546, N533);
buf BUF1 (N547, N520);
nand NAND3 (N548, N545, N5, N402);
and AND3 (N549, N543, N307, N425);
not NOT1 (N550, N538);
nor NOR3 (N551, N541, N10, N424);
nand NAND3 (N552, N534, N437, N23);
buf BUF1 (N553, N547);
and AND4 (N554, N523, N508, N255, N523);
xor XOR2 (N555, N551, N97);
buf BUF1 (N556, N554);
nor NOR2 (N557, N548, N112);
and AND4 (N558, N557, N279, N407, N319);
nand NAND4 (N559, N544, N273, N518, N536);
and AND3 (N560, N555, N26, N176);
nand NAND4 (N561, N559, N184, N437, N16);
and AND2 (N562, N549, N68);
and AND4 (N563, N556, N478, N99, N450);
or OR4 (N564, N562, N52, N292, N270);
and AND3 (N565, N560, N467, N305);
nand NAND4 (N566, N565, N165, N211, N536);
xor XOR2 (N567, N528, N122);
xor XOR2 (N568, N550, N367);
buf BUF1 (N569, N564);
buf BUF1 (N570, N569);
xor XOR2 (N571, N546, N347);
nor NOR2 (N572, N571, N389);
not NOT1 (N573, N563);
nor NOR2 (N574, N572, N90);
or OR2 (N575, N558, N409);
and AND2 (N576, N566, N420);
or OR3 (N577, N568, N353, N323);
and AND4 (N578, N574, N235, N59, N421);
and AND2 (N579, N577, N565);
buf BUF1 (N580, N576);
or OR3 (N581, N579, N55, N434);
xor XOR2 (N582, N580, N61);
not NOT1 (N583, N578);
not NOT1 (N584, N552);
nor NOR4 (N585, N581, N459, N425, N454);
or OR4 (N586, N561, N75, N239, N110);
nor NOR2 (N587, N584, N183);
not NOT1 (N588, N586);
or OR2 (N589, N573, N12);
nor NOR4 (N590, N583, N176, N468, N354);
or OR3 (N591, N570, N355, N550);
and AND3 (N592, N591, N102, N412);
xor XOR2 (N593, N582, N551);
xor XOR2 (N594, N567, N577);
not NOT1 (N595, N588);
buf BUF1 (N596, N589);
nor NOR4 (N597, N590, N454, N270, N230);
xor XOR2 (N598, N575, N550);
or OR4 (N599, N593, N516, N531, N210);
or OR4 (N600, N598, N189, N168, N515);
xor XOR2 (N601, N597, N313);
buf BUF1 (N602, N600);
or OR4 (N603, N596, N467, N113, N438);
and AND2 (N604, N587, N249);
nand NAND2 (N605, N603, N127);
nor NOR2 (N606, N592, N139);
nor NOR3 (N607, N601, N544, N167);
xor XOR2 (N608, N605, N266);
buf BUF1 (N609, N594);
nor NOR3 (N610, N607, N388, N255);
buf BUF1 (N611, N608);
nor NOR4 (N612, N609, N144, N604, N490);
or OR2 (N613, N48, N290);
or OR2 (N614, N585, N122);
not NOT1 (N615, N612);
and AND4 (N616, N615, N1, N463, N230);
buf BUF1 (N617, N616);
buf BUF1 (N618, N606);
xor XOR2 (N619, N553, N74);
nand NAND4 (N620, N617, N451, N340, N67);
buf BUF1 (N621, N595);
buf BUF1 (N622, N611);
not NOT1 (N623, N599);
or OR4 (N624, N618, N365, N361, N524);
and AND4 (N625, N620, N594, N199, N7);
nand NAND4 (N626, N625, N16, N305, N266);
nand NAND2 (N627, N602, N216);
not NOT1 (N628, N614);
nand NAND2 (N629, N624, N55);
and AND2 (N630, N613, N257);
or OR3 (N631, N627, N330, N426);
buf BUF1 (N632, N621);
buf BUF1 (N633, N629);
not NOT1 (N634, N632);
buf BUF1 (N635, N626);
nand NAND2 (N636, N631, N308);
nand NAND3 (N637, N622, N430, N624);
xor XOR2 (N638, N633, N92);
xor XOR2 (N639, N610, N285);
and AND2 (N640, N637, N194);
or OR3 (N641, N634, N161, N3);
and AND2 (N642, N635, N73);
not NOT1 (N643, N640);
nand NAND2 (N644, N623, N293);
and AND4 (N645, N628, N123, N252, N356);
nand NAND2 (N646, N619, N118);
xor XOR2 (N647, N638, N54);
buf BUF1 (N648, N646);
not NOT1 (N649, N642);
and AND4 (N650, N643, N634, N321, N131);
and AND3 (N651, N639, N114, N156);
nand NAND2 (N652, N649, N477);
not NOT1 (N653, N648);
buf BUF1 (N654, N653);
and AND3 (N655, N630, N582, N226);
nor NOR4 (N656, N645, N328, N429, N539);
and AND2 (N657, N636, N602);
and AND3 (N658, N654, N478, N511);
xor XOR2 (N659, N651, N175);
and AND4 (N660, N659, N113, N280, N142);
xor XOR2 (N661, N656, N158);
and AND2 (N662, N661, N197);
not NOT1 (N663, N650);
and AND3 (N664, N662, N99, N410);
buf BUF1 (N665, N660);
buf BUF1 (N666, N655);
and AND4 (N667, N644, N411, N352, N398);
xor XOR2 (N668, N664, N255);
or OR3 (N669, N667, N445, N541);
xor XOR2 (N670, N663, N101);
xor XOR2 (N671, N657, N506);
xor XOR2 (N672, N665, N588);
xor XOR2 (N673, N652, N415);
not NOT1 (N674, N647);
nor NOR4 (N675, N658, N308, N73, N534);
and AND3 (N676, N641, N641, N50);
nor NOR3 (N677, N669, N92, N92);
and AND4 (N678, N675, N656, N469, N37);
buf BUF1 (N679, N670);
not NOT1 (N680, N674);
and AND4 (N681, N677, N489, N549, N215);
nand NAND2 (N682, N679, N126);
nor NOR4 (N683, N666, N163, N635, N400);
and AND3 (N684, N678, N544, N232);
buf BUF1 (N685, N680);
or OR4 (N686, N672, N451, N303, N578);
nor NOR2 (N687, N676, N525);
xor XOR2 (N688, N683, N300);
xor XOR2 (N689, N673, N82);
nand NAND3 (N690, N687, N302, N348);
nand NAND4 (N691, N671, N571, N5, N531);
nand NAND4 (N692, N684, N684, N9, N123);
nand NAND3 (N693, N682, N341, N291);
buf BUF1 (N694, N668);
or OR2 (N695, N691, N339);
not NOT1 (N696, N686);
nor NOR3 (N697, N688, N257, N422);
buf BUF1 (N698, N694);
nand NAND3 (N699, N695, N142, N55);
buf BUF1 (N700, N681);
or OR2 (N701, N690, N468);
nand NAND3 (N702, N689, N500, N295);
nor NOR4 (N703, N698, N171, N541, N360);
xor XOR2 (N704, N701, N533);
nand NAND4 (N705, N685, N613, N465, N535);
buf BUF1 (N706, N700);
xor XOR2 (N707, N705, N460);
or OR2 (N708, N696, N50);
xor XOR2 (N709, N708, N695);
not NOT1 (N710, N709);
endmodule