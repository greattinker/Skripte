// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N12810,N12812,N12797,N12819,N12816,N12817,N12803,N12809,N12811,N12820;

nor NOR2 (N21, N5, N9);
buf BUF1 (N22, N9);
nand NAND4 (N23, N16, N16, N1, N17);
buf BUF1 (N24, N21);
and AND3 (N25, N1, N3, N11);
buf BUF1 (N26, N9);
nand NAND3 (N27, N1, N12, N12);
nand NAND4 (N28, N4, N15, N22, N16);
and AND4 (N29, N24, N19, N14, N15);
or OR4 (N30, N29, N14, N19, N10);
or OR4 (N31, N5, N14, N18, N28);
not NOT1 (N32, N1);
xor XOR2 (N33, N2, N5);
nor NOR2 (N34, N31, N17);
and AND3 (N35, N33, N21, N15);
buf BUF1 (N36, N15);
not NOT1 (N37, N35);
and AND2 (N38, N26, N13);
xor XOR2 (N39, N3, N34);
buf BUF1 (N40, N29);
nand NAND4 (N41, N27, N33, N21, N10);
or OR3 (N42, N32, N32, N35);
nor NOR2 (N43, N25, N2);
buf BUF1 (N44, N41);
or OR3 (N45, N40, N31, N33);
nor NOR2 (N46, N45, N30);
xor XOR2 (N47, N3, N16);
nor NOR3 (N48, N46, N39, N6);
or OR3 (N49, N9, N15, N48);
nor NOR2 (N50, N48, N37);
nor NOR2 (N51, N3, N37);
and AND4 (N52, N36, N11, N12, N41);
xor XOR2 (N53, N49, N18);
not NOT1 (N54, N51);
xor XOR2 (N55, N47, N26);
or OR4 (N56, N38, N41, N44, N14);
buf BUF1 (N57, N32);
xor XOR2 (N58, N55, N51);
and AND3 (N59, N54, N39, N45);
buf BUF1 (N60, N58);
or OR2 (N61, N53, N45);
not NOT1 (N62, N60);
and AND2 (N63, N42, N6);
buf BUF1 (N64, N23);
and AND2 (N65, N59, N43);
nor NOR4 (N66, N63, N64, N3, N3);
nor NOR4 (N67, N60, N43, N16, N24);
buf BUF1 (N68, N59);
or OR2 (N69, N56, N4);
or OR2 (N70, N62, N44);
xor XOR2 (N71, N68, N5);
nor NOR2 (N72, N50, N59);
and AND2 (N73, N70, N60);
nand NAND3 (N74, N66, N57, N4);
nor NOR4 (N75, N28, N52, N53, N65);
buf BUF1 (N76, N3);
xor XOR2 (N77, N41, N59);
not NOT1 (N78, N67);
not NOT1 (N79, N77);
nor NOR2 (N80, N75, N44);
and AND2 (N81, N76, N61);
nor NOR2 (N82, N3, N25);
or OR3 (N83, N71, N7, N29);
nand NAND3 (N84, N79, N73, N14);
and AND4 (N85, N3, N59, N48, N31);
buf BUF1 (N86, N81);
nor NOR4 (N87, N83, N29, N60, N29);
nor NOR3 (N88, N85, N35, N56);
nand NAND4 (N89, N86, N19, N65, N7);
or OR3 (N90, N80, N39, N11);
buf BUF1 (N91, N90);
nor NOR2 (N92, N69, N12);
xor XOR2 (N93, N84, N56);
nand NAND3 (N94, N78, N14, N90);
not NOT1 (N95, N89);
not NOT1 (N96, N94);
not NOT1 (N97, N82);
xor XOR2 (N98, N87, N54);
and AND2 (N99, N97, N78);
buf BUF1 (N100, N91);
not NOT1 (N101, N74);
buf BUF1 (N102, N95);
nor NOR2 (N103, N100, N20);
nand NAND2 (N104, N96, N8);
xor XOR2 (N105, N104, N59);
and AND4 (N106, N88, N6, N15, N84);
or OR3 (N107, N72, N62, N90);
nand NAND3 (N108, N105, N10, N96);
not NOT1 (N109, N108);
or OR2 (N110, N109, N53);
not NOT1 (N111, N110);
xor XOR2 (N112, N99, N103);
buf BUF1 (N113, N63);
and AND2 (N114, N93, N10);
nand NAND3 (N115, N107, N16, N65);
not NOT1 (N116, N111);
buf BUF1 (N117, N92);
buf BUF1 (N118, N98);
not NOT1 (N119, N116);
or OR2 (N120, N117, N23);
xor XOR2 (N121, N112, N10);
nor NOR2 (N122, N121, N67);
nand NAND4 (N123, N106, N69, N29, N102);
or OR2 (N124, N38, N68);
and AND2 (N125, N119, N21);
buf BUF1 (N126, N118);
xor XOR2 (N127, N101, N115);
or OR3 (N128, N69, N8, N100);
nor NOR3 (N129, N122, N125, N91);
not NOT1 (N130, N103);
buf BUF1 (N131, N113);
nand NAND4 (N132, N124, N49, N117, N43);
nand NAND4 (N133, N132, N129, N81, N60);
nand NAND2 (N134, N130, N107);
nor NOR3 (N135, N27, N110, N133);
and AND4 (N136, N50, N107, N90, N78);
xor XOR2 (N137, N136, N88);
or OR4 (N138, N126, N96, N112, N136);
and AND3 (N139, N131, N22, N94);
and AND3 (N140, N134, N27, N113);
nor NOR4 (N141, N138, N96, N56, N5);
and AND4 (N142, N114, N10, N39, N124);
buf BUF1 (N143, N120);
xor XOR2 (N144, N140, N21);
nand NAND4 (N145, N137, N103, N2, N119);
xor XOR2 (N146, N144, N69);
buf BUF1 (N147, N135);
or OR4 (N148, N147, N100, N107, N67);
buf BUF1 (N149, N146);
nor NOR2 (N150, N123, N146);
not NOT1 (N151, N139);
or OR4 (N152, N149, N83, N40, N38);
xor XOR2 (N153, N141, N11);
xor XOR2 (N154, N143, N47);
xor XOR2 (N155, N127, N82);
nand NAND4 (N156, N153, N72, N123, N118);
xor XOR2 (N157, N155, N45);
or OR3 (N158, N151, N155, N114);
and AND2 (N159, N157, N37);
buf BUF1 (N160, N156);
buf BUF1 (N161, N128);
or OR2 (N162, N160, N152);
xor XOR2 (N163, N5, N134);
nand NAND4 (N164, N142, N26, N130, N124);
buf BUF1 (N165, N148);
buf BUF1 (N166, N158);
nand NAND4 (N167, N161, N32, N43, N15);
not NOT1 (N168, N165);
or OR2 (N169, N145, N143);
buf BUF1 (N170, N163);
xor XOR2 (N171, N167, N94);
and AND4 (N172, N171, N26, N90, N62);
or OR3 (N173, N150, N50, N87);
not NOT1 (N174, N172);
or OR4 (N175, N170, N140, N55, N24);
or OR3 (N176, N174, N17, N6);
not NOT1 (N177, N162);
nand NAND2 (N178, N173, N153);
or OR2 (N179, N175, N103);
or OR2 (N180, N169, N161);
buf BUF1 (N181, N159);
not NOT1 (N182, N164);
nand NAND2 (N183, N179, N21);
and AND4 (N184, N168, N83, N115, N134);
and AND3 (N185, N183, N73, N86);
and AND2 (N186, N184, N158);
buf BUF1 (N187, N185);
not NOT1 (N188, N177);
buf BUF1 (N189, N187);
or OR4 (N190, N176, N15, N86, N59);
or OR4 (N191, N166, N59, N36, N186);
and AND3 (N192, N27, N190, N69);
nor NOR2 (N193, N27, N186);
and AND4 (N194, N178, N171, N176, N100);
nor NOR2 (N195, N189, N94);
not NOT1 (N196, N193);
not NOT1 (N197, N188);
or OR3 (N198, N195, N83, N71);
xor XOR2 (N199, N198, N20);
or OR2 (N200, N199, N134);
not NOT1 (N201, N194);
buf BUF1 (N202, N181);
nor NOR4 (N203, N180, N140, N158, N85);
nand NAND4 (N204, N192, N170, N18, N134);
nand NAND4 (N205, N201, N125, N145, N103);
or OR4 (N206, N205, N58, N103, N137);
xor XOR2 (N207, N203, N180);
nor NOR2 (N208, N202, N188);
xor XOR2 (N209, N200, N2);
and AND2 (N210, N204, N12);
nor NOR3 (N211, N206, N142, N140);
not NOT1 (N212, N211);
or OR2 (N213, N191, N81);
nand NAND2 (N214, N210, N124);
and AND3 (N215, N208, N16, N154);
not NOT1 (N216, N151);
or OR2 (N217, N215, N186);
not NOT1 (N218, N209);
or OR4 (N219, N182, N49, N13, N165);
or OR4 (N220, N217, N75, N126, N171);
or OR3 (N221, N219, N209, N121);
and AND4 (N222, N214, N165, N79, N161);
or OR4 (N223, N197, N94, N95, N79);
not NOT1 (N224, N216);
or OR2 (N225, N218, N143);
and AND2 (N226, N223, N215);
or OR2 (N227, N212, N96);
buf BUF1 (N228, N222);
nor NOR3 (N229, N196, N180, N178);
not NOT1 (N230, N213);
and AND4 (N231, N226, N156, N43, N165);
nor NOR4 (N232, N230, N132, N146, N222);
not NOT1 (N233, N228);
not NOT1 (N234, N207);
not NOT1 (N235, N229);
buf BUF1 (N236, N231);
nor NOR3 (N237, N220, N207, N81);
nor NOR3 (N238, N221, N132, N36);
nor NOR4 (N239, N232, N75, N163, N75);
nand NAND2 (N240, N237, N163);
buf BUF1 (N241, N224);
not NOT1 (N242, N235);
nor NOR3 (N243, N240, N189, N56);
nor NOR2 (N244, N238, N195);
nand NAND2 (N245, N227, N92);
not NOT1 (N246, N239);
buf BUF1 (N247, N242);
not NOT1 (N248, N236);
xor XOR2 (N249, N241, N165);
nor NOR2 (N250, N245, N9);
xor XOR2 (N251, N250, N236);
and AND3 (N252, N246, N206, N170);
xor XOR2 (N253, N234, N200);
not NOT1 (N254, N225);
or OR3 (N255, N253, N4, N45);
buf BUF1 (N256, N252);
nor NOR3 (N257, N244, N178, N27);
not NOT1 (N258, N249);
not NOT1 (N259, N233);
and AND3 (N260, N258, N55, N227);
xor XOR2 (N261, N254, N187);
nand NAND2 (N262, N248, N166);
xor XOR2 (N263, N247, N46);
or OR2 (N264, N263, N118);
nand NAND4 (N265, N262, N71, N163, N246);
nand NAND4 (N266, N265, N181, N37, N198);
or OR2 (N267, N259, N242);
not NOT1 (N268, N243);
nand NAND3 (N269, N261, N251, N148);
and AND4 (N270, N175, N165, N212, N47);
or OR3 (N271, N269, N112, N181);
not NOT1 (N272, N260);
nor NOR4 (N273, N255, N97, N247, N63);
nand NAND3 (N274, N271, N88, N97);
buf BUF1 (N275, N256);
nand NAND2 (N276, N257, N67);
nand NAND4 (N277, N270, N76, N49, N229);
xor XOR2 (N278, N268, N109);
or OR3 (N279, N275, N80, N36);
nand NAND3 (N280, N279, N229, N52);
nand NAND4 (N281, N278, N64, N39, N279);
nand NAND4 (N282, N276, N209, N136, N274);
xor XOR2 (N283, N204, N67);
or OR2 (N284, N280, N235);
xor XOR2 (N285, N283, N276);
nand NAND3 (N286, N281, N256, N204);
nand NAND2 (N287, N282, N27);
not NOT1 (N288, N287);
not NOT1 (N289, N277);
or OR2 (N290, N267, N94);
or OR3 (N291, N290, N56, N176);
buf BUF1 (N292, N291);
not NOT1 (N293, N292);
nand NAND3 (N294, N272, N284, N20);
xor XOR2 (N295, N32, N63);
buf BUF1 (N296, N294);
and AND3 (N297, N295, N171, N135);
buf BUF1 (N298, N288);
xor XOR2 (N299, N285, N280);
or OR4 (N300, N264, N294, N160, N286);
not NOT1 (N301, N6);
xor XOR2 (N302, N266, N61);
and AND2 (N303, N289, N167);
or OR2 (N304, N298, N93);
xor XOR2 (N305, N304, N234);
and AND2 (N306, N293, N70);
nor NOR2 (N307, N306, N54);
nand NAND3 (N308, N273, N222, N148);
not NOT1 (N309, N305);
or OR4 (N310, N301, N212, N190, N65);
nor NOR3 (N311, N299, N35, N280);
or OR4 (N312, N310, N25, N120, N256);
nand NAND3 (N313, N303, N146, N78);
not NOT1 (N314, N308);
and AND4 (N315, N313, N304, N211, N44);
or OR4 (N316, N311, N141, N159, N45);
and AND2 (N317, N312, N175);
and AND2 (N318, N297, N182);
xor XOR2 (N319, N307, N62);
or OR3 (N320, N319, N291, N40);
nor NOR2 (N321, N300, N185);
buf BUF1 (N322, N318);
buf BUF1 (N323, N296);
or OR3 (N324, N322, N245, N60);
nor NOR4 (N325, N323, N179, N68, N16);
nand NAND2 (N326, N315, N302);
xor XOR2 (N327, N300, N72);
or OR4 (N328, N320, N243, N305, N90);
buf BUF1 (N329, N324);
nor NOR3 (N330, N316, N44, N50);
nand NAND2 (N331, N330, N26);
buf BUF1 (N332, N326);
xor XOR2 (N333, N332, N270);
nor NOR4 (N334, N327, N154, N126, N199);
and AND4 (N335, N317, N300, N68, N11);
buf BUF1 (N336, N325);
and AND3 (N337, N334, N153, N295);
buf BUF1 (N338, N333);
and AND3 (N339, N336, N158, N71);
nor NOR3 (N340, N335, N261, N135);
not NOT1 (N341, N314);
and AND2 (N342, N331, N4);
nor NOR4 (N343, N340, N338, N54, N6);
xor XOR2 (N344, N226, N336);
buf BUF1 (N345, N342);
nor NOR3 (N346, N321, N290, N194);
buf BUF1 (N347, N337);
and AND2 (N348, N339, N308);
buf BUF1 (N349, N309);
xor XOR2 (N350, N346, N186);
nor NOR4 (N351, N349, N127, N151, N18);
nor NOR4 (N352, N350, N63, N18, N266);
xor XOR2 (N353, N348, N42);
xor XOR2 (N354, N353, N207);
or OR4 (N355, N352, N141, N2, N316);
buf BUF1 (N356, N328);
xor XOR2 (N357, N343, N276);
buf BUF1 (N358, N351);
nand NAND4 (N359, N354, N112, N123, N134);
or OR4 (N360, N329, N260, N127, N180);
or OR3 (N361, N359, N253, N155);
and AND2 (N362, N360, N19);
and AND2 (N363, N358, N290);
xor XOR2 (N364, N362, N232);
and AND3 (N365, N347, N254, N334);
not NOT1 (N366, N361);
not NOT1 (N367, N365);
nor NOR4 (N368, N363, N364, N38, N229);
and AND2 (N369, N269, N250);
xor XOR2 (N370, N356, N330);
buf BUF1 (N371, N355);
nor NOR3 (N372, N357, N324, N155);
nand NAND2 (N373, N372, N295);
buf BUF1 (N374, N371);
buf BUF1 (N375, N368);
nand NAND2 (N376, N369, N242);
or OR3 (N377, N366, N301, N104);
and AND4 (N378, N376, N57, N248, N18);
nand NAND2 (N379, N373, N222);
nand NAND2 (N380, N345, N348);
or OR3 (N381, N377, N284, N251);
or OR2 (N382, N370, N193);
or OR2 (N383, N381, N116);
buf BUF1 (N384, N382);
buf BUF1 (N385, N383);
xor XOR2 (N386, N380, N130);
xor XOR2 (N387, N344, N7);
not NOT1 (N388, N385);
and AND2 (N389, N387, N305);
buf BUF1 (N390, N375);
nand NAND3 (N391, N390, N283, N57);
xor XOR2 (N392, N386, N208);
xor XOR2 (N393, N379, N366);
nor NOR4 (N394, N391, N369, N302, N299);
or OR4 (N395, N388, N115, N161, N94);
or OR2 (N396, N392, N17);
and AND3 (N397, N341, N270, N140);
not NOT1 (N398, N389);
buf BUF1 (N399, N398);
and AND3 (N400, N395, N232, N276);
not NOT1 (N401, N394);
and AND2 (N402, N400, N106);
buf BUF1 (N403, N401);
nand NAND2 (N404, N399, N28);
xor XOR2 (N405, N404, N189);
nor NOR4 (N406, N396, N263, N19, N404);
not NOT1 (N407, N403);
and AND2 (N408, N384, N340);
or OR2 (N409, N374, N378);
xor XOR2 (N410, N327, N258);
nand NAND2 (N411, N408, N333);
nor NOR4 (N412, N397, N46, N168, N312);
or OR3 (N413, N412, N123, N291);
buf BUF1 (N414, N413);
buf BUF1 (N415, N414);
or OR2 (N416, N415, N136);
nand NAND4 (N417, N416, N181, N78, N344);
or OR4 (N418, N402, N358, N313, N239);
nor NOR4 (N419, N367, N77, N137, N318);
nand NAND2 (N420, N410, N352);
nor NOR2 (N421, N419, N129);
nor NOR4 (N422, N409, N24, N278, N160);
and AND3 (N423, N411, N66, N29);
xor XOR2 (N424, N405, N184);
or OR4 (N425, N420, N287, N342, N287);
buf BUF1 (N426, N393);
not NOT1 (N427, N426);
xor XOR2 (N428, N417, N110);
nand NAND3 (N429, N421, N200, N157);
xor XOR2 (N430, N423, N322);
nor NOR2 (N431, N424, N208);
nand NAND2 (N432, N425, N240);
xor XOR2 (N433, N422, N181);
buf BUF1 (N434, N418);
nor NOR4 (N435, N429, N73, N273, N148);
buf BUF1 (N436, N434);
not NOT1 (N437, N430);
nor NOR4 (N438, N428, N382, N135, N123);
xor XOR2 (N439, N427, N415);
nand NAND3 (N440, N437, N368, N304);
nor NOR3 (N441, N436, N266, N59);
buf BUF1 (N442, N441);
nor NOR4 (N443, N439, N25, N345, N168);
not NOT1 (N444, N432);
and AND4 (N445, N407, N390, N52, N197);
nand NAND3 (N446, N433, N169, N229);
xor XOR2 (N447, N435, N183);
or OR3 (N448, N446, N234, N198);
and AND2 (N449, N442, N291);
buf BUF1 (N450, N406);
not NOT1 (N451, N450);
xor XOR2 (N452, N451, N357);
nor NOR4 (N453, N448, N394, N431, N219);
nand NAND3 (N454, N279, N425, N145);
xor XOR2 (N455, N443, N401);
nor NOR3 (N456, N447, N291, N416);
nand NAND3 (N457, N456, N247, N32);
not NOT1 (N458, N449);
nor NOR3 (N459, N438, N26, N100);
xor XOR2 (N460, N453, N237);
not NOT1 (N461, N440);
or OR3 (N462, N460, N370, N13);
and AND4 (N463, N459, N263, N412, N143);
xor XOR2 (N464, N455, N170);
not NOT1 (N465, N452);
xor XOR2 (N466, N465, N176);
or OR4 (N467, N444, N159, N164, N433);
nor NOR2 (N468, N457, N415);
nor NOR2 (N469, N462, N184);
or OR4 (N470, N467, N311, N35, N362);
xor XOR2 (N471, N468, N4);
nor NOR2 (N472, N469, N354);
nor NOR2 (N473, N471, N415);
buf BUF1 (N474, N464);
xor XOR2 (N475, N466, N53);
nand NAND4 (N476, N473, N191, N34, N315);
nand NAND4 (N477, N445, N362, N331, N309);
nand NAND4 (N478, N461, N153, N83, N219);
or OR3 (N479, N463, N436, N122);
buf BUF1 (N480, N454);
buf BUF1 (N481, N470);
xor XOR2 (N482, N472, N135);
nand NAND4 (N483, N477, N385, N446, N463);
nor NOR3 (N484, N483, N42, N424);
not NOT1 (N485, N476);
buf BUF1 (N486, N484);
nor NOR3 (N487, N482, N59, N61);
buf BUF1 (N488, N479);
buf BUF1 (N489, N480);
and AND2 (N490, N475, N484);
nor NOR2 (N491, N485, N288);
or OR4 (N492, N489, N31, N206, N345);
nor NOR2 (N493, N491, N315);
not NOT1 (N494, N478);
nand NAND2 (N495, N490, N58);
or OR4 (N496, N492, N64, N97, N44);
and AND2 (N497, N486, N344);
not NOT1 (N498, N496);
or OR3 (N499, N488, N469, N423);
nor NOR2 (N500, N474, N104);
not NOT1 (N501, N458);
nand NAND2 (N502, N499, N302);
buf BUF1 (N503, N493);
nor NOR3 (N504, N500, N133, N146);
and AND2 (N505, N498, N151);
not NOT1 (N506, N503);
or OR4 (N507, N495, N65, N21, N339);
buf BUF1 (N508, N507);
nor NOR2 (N509, N504, N87);
and AND2 (N510, N505, N324);
and AND3 (N511, N481, N155, N242);
nand NAND2 (N512, N502, N352);
nor NOR2 (N513, N494, N23);
buf BUF1 (N514, N497);
nand NAND2 (N515, N511, N325);
or OR4 (N516, N514, N467, N115, N499);
xor XOR2 (N517, N512, N516);
nor NOR2 (N518, N266, N176);
not NOT1 (N519, N487);
not NOT1 (N520, N518);
not NOT1 (N521, N510);
xor XOR2 (N522, N517, N341);
and AND4 (N523, N501, N254, N490, N290);
nand NAND3 (N524, N519, N190, N487);
or OR3 (N525, N513, N471, N203);
xor XOR2 (N526, N522, N358);
and AND2 (N527, N506, N157);
buf BUF1 (N528, N508);
and AND2 (N529, N515, N268);
nand NAND2 (N530, N523, N452);
nor NOR2 (N531, N530, N475);
not NOT1 (N532, N525);
not NOT1 (N533, N526);
nand NAND2 (N534, N531, N165);
buf BUF1 (N535, N532);
and AND4 (N536, N534, N269, N509, N503);
not NOT1 (N537, N46);
nor NOR3 (N538, N536, N254, N400);
and AND4 (N539, N528, N394, N286, N231);
not NOT1 (N540, N535);
nor NOR4 (N541, N538, N365, N382, N219);
nand NAND3 (N542, N529, N437, N459);
not NOT1 (N543, N533);
and AND4 (N544, N542, N40, N279, N182);
not NOT1 (N545, N541);
buf BUF1 (N546, N520);
xor XOR2 (N547, N524, N17);
or OR4 (N548, N543, N443, N170, N383);
nor NOR2 (N549, N537, N237);
or OR3 (N550, N545, N371, N225);
buf BUF1 (N551, N546);
or OR4 (N552, N527, N411, N71, N35);
not NOT1 (N553, N549);
not NOT1 (N554, N540);
nor NOR3 (N555, N551, N376, N362);
xor XOR2 (N556, N555, N521);
or OR3 (N557, N280, N16, N80);
buf BUF1 (N558, N550);
and AND2 (N559, N548, N519);
nor NOR2 (N560, N557, N349);
not NOT1 (N561, N559);
not NOT1 (N562, N547);
or OR3 (N563, N558, N382, N403);
nand NAND3 (N564, N563, N311, N407);
nor NOR4 (N565, N544, N307, N498, N72);
not NOT1 (N566, N564);
nand NAND3 (N567, N566, N494, N245);
or OR3 (N568, N539, N164, N182);
and AND4 (N569, N565, N318, N548, N411);
nand NAND2 (N570, N562, N523);
nand NAND4 (N571, N568, N348, N172, N559);
nand NAND2 (N572, N556, N46);
and AND2 (N573, N570, N433);
and AND2 (N574, N560, N101);
or OR4 (N575, N561, N176, N393, N330);
or OR3 (N576, N575, N571, N481);
and AND2 (N577, N537, N307);
not NOT1 (N578, N569);
nor NOR3 (N579, N576, N544, N266);
nand NAND3 (N580, N578, N76, N524);
not NOT1 (N581, N579);
buf BUF1 (N582, N580);
buf BUF1 (N583, N567);
not NOT1 (N584, N554);
nand NAND4 (N585, N577, N438, N298, N246);
xor XOR2 (N586, N552, N466);
xor XOR2 (N587, N553, N239);
buf BUF1 (N588, N572);
nor NOR3 (N589, N584, N422, N513);
and AND2 (N590, N588, N398);
nand NAND3 (N591, N586, N30, N367);
or OR4 (N592, N589, N295, N91, N362);
xor XOR2 (N593, N591, N481);
nor NOR2 (N594, N592, N45);
xor XOR2 (N595, N594, N241);
buf BUF1 (N596, N573);
xor XOR2 (N597, N574, N515);
xor XOR2 (N598, N593, N527);
or OR2 (N599, N597, N180);
nand NAND2 (N600, N599, N49);
and AND4 (N601, N582, N96, N205, N531);
not NOT1 (N602, N583);
nand NAND4 (N603, N587, N82, N352, N133);
nand NAND3 (N604, N581, N328, N227);
nor NOR3 (N605, N598, N359, N328);
and AND3 (N606, N590, N488, N451);
xor XOR2 (N607, N603, N136);
nand NAND4 (N608, N604, N235, N332, N88);
buf BUF1 (N609, N600);
nor NOR3 (N610, N601, N17, N301);
nand NAND4 (N611, N607, N467, N258, N174);
xor XOR2 (N612, N596, N442);
nand NAND2 (N613, N585, N189);
not NOT1 (N614, N610);
nor NOR3 (N615, N614, N333, N578);
xor XOR2 (N616, N611, N522);
nor NOR2 (N617, N613, N531);
buf BUF1 (N618, N615);
nor NOR4 (N619, N616, N275, N110, N296);
or OR4 (N620, N617, N114, N456, N254);
nand NAND3 (N621, N605, N78, N437);
nand NAND2 (N622, N606, N393);
and AND2 (N623, N622, N603);
nand NAND3 (N624, N620, N67, N565);
or OR4 (N625, N608, N570, N286, N202);
xor XOR2 (N626, N625, N145);
and AND4 (N627, N612, N88, N476, N491);
nor NOR4 (N628, N621, N358, N506, N563);
not NOT1 (N629, N623);
xor XOR2 (N630, N628, N221);
not NOT1 (N631, N618);
buf BUF1 (N632, N631);
nor NOR2 (N633, N629, N1);
and AND3 (N634, N632, N267, N104);
and AND3 (N635, N633, N204, N208);
and AND3 (N636, N635, N382, N166);
or OR4 (N637, N634, N211, N453, N375);
not NOT1 (N638, N609);
nand NAND2 (N639, N626, N469);
not NOT1 (N640, N638);
or OR4 (N641, N595, N204, N70, N142);
buf BUF1 (N642, N630);
nor NOR2 (N643, N641, N74);
or OR4 (N644, N624, N625, N319, N469);
and AND2 (N645, N644, N401);
and AND4 (N646, N636, N508, N329, N184);
nor NOR2 (N647, N637, N13);
and AND3 (N648, N643, N412, N456);
or OR2 (N649, N639, N556);
not NOT1 (N650, N647);
and AND2 (N651, N642, N558);
nand NAND4 (N652, N602, N3, N644, N181);
buf BUF1 (N653, N649);
and AND3 (N654, N646, N64, N315);
or OR4 (N655, N653, N174, N286, N338);
not NOT1 (N656, N640);
nand NAND2 (N657, N656, N304);
buf BUF1 (N658, N652);
nor NOR4 (N659, N658, N151, N242, N196);
buf BUF1 (N660, N659);
buf BUF1 (N661, N650);
and AND2 (N662, N657, N274);
or OR2 (N663, N627, N325);
xor XOR2 (N664, N654, N634);
nand NAND2 (N665, N661, N300);
nand NAND3 (N666, N665, N607, N627);
or OR4 (N667, N663, N653, N382, N407);
and AND2 (N668, N662, N16);
nor NOR2 (N669, N648, N647);
not NOT1 (N670, N645);
nand NAND3 (N671, N666, N415, N46);
buf BUF1 (N672, N671);
not NOT1 (N673, N655);
nor NOR2 (N674, N673, N158);
nand NAND3 (N675, N668, N237, N372);
nor NOR2 (N676, N619, N96);
nor NOR2 (N677, N672, N230);
and AND4 (N678, N675, N254, N143, N657);
nand NAND3 (N679, N667, N151, N498);
buf BUF1 (N680, N669);
nand NAND2 (N681, N660, N527);
nor NOR3 (N682, N679, N325, N168);
buf BUF1 (N683, N674);
buf BUF1 (N684, N670);
nand NAND2 (N685, N677, N604);
and AND3 (N686, N681, N359, N299);
nand NAND3 (N687, N676, N550, N145);
xor XOR2 (N688, N680, N383);
nand NAND4 (N689, N685, N2, N591, N29);
or OR4 (N690, N682, N430, N102, N437);
not NOT1 (N691, N651);
not NOT1 (N692, N664);
nor NOR3 (N693, N687, N648, N673);
nand NAND3 (N694, N689, N613, N464);
and AND2 (N695, N684, N151);
nand NAND2 (N696, N683, N685);
buf BUF1 (N697, N688);
buf BUF1 (N698, N690);
or OR3 (N699, N697, N627, N170);
buf BUF1 (N700, N696);
and AND4 (N701, N698, N82, N82, N396);
not NOT1 (N702, N686);
and AND4 (N703, N700, N28, N510, N108);
or OR4 (N704, N703, N159, N646, N357);
xor XOR2 (N705, N699, N555);
nor NOR2 (N706, N705, N328);
nor NOR2 (N707, N704, N265);
buf BUF1 (N708, N692);
xor XOR2 (N709, N707, N96);
buf BUF1 (N710, N691);
or OR4 (N711, N695, N655, N38, N678);
buf BUF1 (N712, N112);
nand NAND2 (N713, N706, N478);
xor XOR2 (N714, N709, N78);
xor XOR2 (N715, N708, N100);
or OR2 (N716, N701, N220);
xor XOR2 (N717, N712, N210);
nor NOR3 (N718, N713, N419, N290);
not NOT1 (N719, N710);
and AND3 (N720, N693, N192, N621);
not NOT1 (N721, N694);
nor NOR3 (N722, N711, N213, N308);
and AND2 (N723, N716, N122);
xor XOR2 (N724, N718, N17);
buf BUF1 (N725, N724);
xor XOR2 (N726, N714, N544);
not NOT1 (N727, N721);
or OR4 (N728, N727, N131, N538, N586);
buf BUF1 (N729, N720);
nor NOR3 (N730, N702, N218, N158);
nor NOR4 (N731, N725, N552, N680, N620);
not NOT1 (N732, N730);
nor NOR2 (N733, N722, N303);
not NOT1 (N734, N715);
xor XOR2 (N735, N731, N16);
and AND3 (N736, N732, N318, N140);
and AND2 (N737, N719, N284);
nor NOR2 (N738, N729, N97);
or OR2 (N739, N717, N122);
xor XOR2 (N740, N738, N434);
and AND2 (N741, N728, N712);
and AND4 (N742, N723, N14, N686, N163);
buf BUF1 (N743, N737);
buf BUF1 (N744, N734);
and AND4 (N745, N741, N703, N723, N446);
or OR4 (N746, N745, N50, N704, N605);
nor NOR3 (N747, N744, N666, N621);
xor XOR2 (N748, N733, N290);
not NOT1 (N749, N739);
or OR2 (N750, N740, N49);
or OR4 (N751, N726, N85, N487, N597);
not NOT1 (N752, N736);
not NOT1 (N753, N751);
buf BUF1 (N754, N746);
nand NAND4 (N755, N747, N629, N8, N484);
nor NOR3 (N756, N752, N596, N677);
nand NAND3 (N757, N750, N614, N375);
not NOT1 (N758, N753);
xor XOR2 (N759, N748, N475);
xor XOR2 (N760, N758, N693);
not NOT1 (N761, N756);
nand NAND2 (N762, N742, N597);
and AND4 (N763, N755, N14, N488, N380);
nor NOR2 (N764, N760, N190);
or OR4 (N765, N759, N339, N449, N177);
xor XOR2 (N766, N764, N135);
or OR4 (N767, N762, N485, N737, N139);
and AND2 (N768, N767, N491);
xor XOR2 (N769, N735, N376);
nand NAND4 (N770, N766, N389, N68, N251);
nor NOR2 (N771, N754, N322);
nand NAND4 (N772, N770, N38, N40, N496);
and AND3 (N773, N768, N111, N397);
or OR2 (N774, N749, N411);
buf BUF1 (N775, N761);
and AND2 (N776, N743, N563);
or OR2 (N777, N776, N627);
not NOT1 (N778, N773);
not NOT1 (N779, N775);
nand NAND2 (N780, N765, N201);
or OR3 (N781, N757, N14, N18);
buf BUF1 (N782, N780);
not NOT1 (N783, N779);
nor NOR3 (N784, N781, N164, N714);
xor XOR2 (N785, N782, N760);
not NOT1 (N786, N769);
xor XOR2 (N787, N786, N682);
buf BUF1 (N788, N784);
buf BUF1 (N789, N788);
nand NAND2 (N790, N783, N745);
nand NAND4 (N791, N778, N39, N756, N91);
and AND4 (N792, N790, N168, N420, N666);
and AND2 (N793, N789, N709);
nand NAND4 (N794, N774, N506, N489, N574);
and AND3 (N795, N791, N7, N760);
not NOT1 (N796, N772);
xor XOR2 (N797, N771, N428);
and AND3 (N798, N796, N556, N389);
buf BUF1 (N799, N787);
not NOT1 (N800, N799);
and AND2 (N801, N797, N232);
buf BUF1 (N802, N777);
not NOT1 (N803, N795);
buf BUF1 (N804, N800);
nand NAND4 (N805, N785, N290, N105, N324);
xor XOR2 (N806, N794, N467);
or OR3 (N807, N806, N467, N377);
nand NAND4 (N808, N792, N599, N234, N442);
nor NOR2 (N809, N798, N312);
xor XOR2 (N810, N763, N108);
nor NOR4 (N811, N793, N455, N63, N405);
or OR4 (N812, N805, N196, N679, N602);
and AND4 (N813, N808, N281, N155, N234);
and AND4 (N814, N812, N344, N7, N389);
not NOT1 (N815, N810);
nor NOR2 (N816, N814, N653);
buf BUF1 (N817, N803);
xor XOR2 (N818, N807, N94);
nor NOR4 (N819, N816, N431, N255, N112);
and AND4 (N820, N818, N738, N317, N168);
and AND3 (N821, N801, N76, N315);
nor NOR3 (N822, N811, N511, N178);
nand NAND4 (N823, N820, N298, N90, N8);
xor XOR2 (N824, N823, N579);
and AND2 (N825, N819, N707);
nor NOR3 (N826, N813, N556, N261);
or OR3 (N827, N825, N231, N572);
nand NAND2 (N828, N821, N760);
xor XOR2 (N829, N802, N393);
xor XOR2 (N830, N804, N463);
nand NAND2 (N831, N829, N269);
not NOT1 (N832, N817);
nor NOR2 (N833, N822, N125);
xor XOR2 (N834, N809, N764);
buf BUF1 (N835, N828);
nand NAND3 (N836, N826, N9, N345);
not NOT1 (N837, N835);
nor NOR3 (N838, N824, N438, N507);
nor NOR4 (N839, N836, N744, N774, N511);
and AND4 (N840, N831, N166, N369, N97);
xor XOR2 (N841, N840, N126);
not NOT1 (N842, N841);
buf BUF1 (N843, N834);
xor XOR2 (N844, N833, N44);
nand NAND3 (N845, N844, N680, N519);
not NOT1 (N846, N843);
nand NAND3 (N847, N827, N247, N534);
nand NAND4 (N848, N842, N370, N406, N679);
buf BUF1 (N849, N832);
not NOT1 (N850, N830);
xor XOR2 (N851, N837, N355);
not NOT1 (N852, N815);
not NOT1 (N853, N850);
nand NAND2 (N854, N845, N93);
nor NOR3 (N855, N854, N806, N177);
or OR4 (N856, N847, N458, N514, N179);
and AND3 (N857, N855, N378, N337);
not NOT1 (N858, N848);
xor XOR2 (N859, N852, N584);
nand NAND2 (N860, N851, N796);
not NOT1 (N861, N838);
buf BUF1 (N862, N856);
nand NAND2 (N863, N858, N196);
buf BUF1 (N864, N849);
xor XOR2 (N865, N846, N218);
and AND2 (N866, N862, N367);
not NOT1 (N867, N863);
not NOT1 (N868, N866);
xor XOR2 (N869, N857, N577);
nor NOR2 (N870, N868, N394);
not NOT1 (N871, N869);
or OR2 (N872, N839, N174);
buf BUF1 (N873, N865);
nand NAND4 (N874, N859, N738, N195, N14);
nor NOR3 (N875, N853, N773, N719);
nand NAND4 (N876, N860, N432, N376, N104);
xor XOR2 (N877, N872, N659);
xor XOR2 (N878, N876, N320);
or OR3 (N879, N870, N585, N485);
buf BUF1 (N880, N861);
nand NAND2 (N881, N871, N254);
buf BUF1 (N882, N873);
nand NAND4 (N883, N867, N376, N139, N457);
xor XOR2 (N884, N883, N667);
buf BUF1 (N885, N875);
not NOT1 (N886, N885);
not NOT1 (N887, N874);
buf BUF1 (N888, N880);
not NOT1 (N889, N881);
buf BUF1 (N890, N879);
not NOT1 (N891, N889);
nand NAND3 (N892, N886, N256, N261);
nor NOR4 (N893, N864, N854, N644, N488);
or OR2 (N894, N890, N836);
nor NOR3 (N895, N888, N821, N869);
or OR3 (N896, N877, N726, N371);
not NOT1 (N897, N891);
or OR2 (N898, N897, N143);
xor XOR2 (N899, N887, N705);
or OR4 (N900, N898, N327, N890, N709);
nand NAND3 (N901, N896, N304, N110);
not NOT1 (N902, N878);
nor NOR3 (N903, N892, N239, N640);
xor XOR2 (N904, N903, N91);
nand NAND4 (N905, N895, N242, N102, N82);
and AND2 (N906, N884, N494);
not NOT1 (N907, N882);
nor NOR2 (N908, N904, N79);
and AND4 (N909, N893, N872, N900, N157);
buf BUF1 (N910, N113);
nor NOR4 (N911, N905, N841, N379, N234);
xor XOR2 (N912, N901, N598);
not NOT1 (N913, N899);
nand NAND3 (N914, N909, N841, N88);
and AND3 (N915, N912, N359, N625);
nand NAND4 (N916, N913, N881, N73, N573);
or OR2 (N917, N915, N402);
buf BUF1 (N918, N894);
nand NAND2 (N919, N902, N13);
nor NOR3 (N920, N910, N712, N99);
nor NOR3 (N921, N916, N764, N359);
or OR4 (N922, N911, N257, N430, N127);
xor XOR2 (N923, N917, N701);
and AND4 (N924, N922, N277, N180, N466);
nor NOR4 (N925, N908, N698, N74, N500);
xor XOR2 (N926, N914, N626);
and AND4 (N927, N920, N98, N776, N134);
buf BUF1 (N928, N926);
not NOT1 (N929, N928);
xor XOR2 (N930, N923, N398);
not NOT1 (N931, N919);
nor NOR2 (N932, N929, N111);
or OR2 (N933, N932, N641);
and AND4 (N934, N927, N862, N580, N435);
nand NAND2 (N935, N934, N233);
nand NAND3 (N936, N918, N791, N916);
or OR4 (N937, N906, N75, N520, N705);
nand NAND2 (N938, N921, N293);
nand NAND2 (N939, N925, N723);
or OR4 (N940, N936, N476, N387, N290);
and AND4 (N941, N937, N934, N257, N568);
nor NOR2 (N942, N935, N303);
nand NAND2 (N943, N907, N52);
and AND4 (N944, N931, N270, N759, N75);
and AND3 (N945, N938, N374, N846);
and AND4 (N946, N924, N175, N82, N215);
nor NOR4 (N947, N941, N332, N883, N894);
buf BUF1 (N948, N945);
not NOT1 (N949, N944);
nor NOR2 (N950, N940, N694);
xor XOR2 (N951, N949, N455);
buf BUF1 (N952, N942);
not NOT1 (N953, N948);
xor XOR2 (N954, N930, N910);
and AND3 (N955, N953, N861, N945);
nor NOR2 (N956, N947, N524);
and AND4 (N957, N952, N115, N727, N620);
buf BUF1 (N958, N950);
or OR2 (N959, N939, N444);
nand NAND3 (N960, N954, N711, N21);
or OR3 (N961, N955, N113, N596);
xor XOR2 (N962, N958, N133);
xor XOR2 (N963, N946, N3);
nand NAND4 (N964, N959, N821, N251, N12);
or OR3 (N965, N957, N928, N40);
and AND2 (N966, N962, N950);
not NOT1 (N967, N943);
nor NOR2 (N968, N963, N581);
not NOT1 (N969, N951);
or OR2 (N970, N966, N610);
or OR2 (N971, N961, N85);
xor XOR2 (N972, N968, N836);
buf BUF1 (N973, N972);
xor XOR2 (N974, N971, N602);
nor NOR3 (N975, N967, N639, N919);
nor NOR3 (N976, N974, N221, N569);
not NOT1 (N977, N960);
or OR2 (N978, N970, N588);
nand NAND2 (N979, N965, N743);
xor XOR2 (N980, N933, N590);
buf BUF1 (N981, N956);
nor NOR3 (N982, N969, N460, N262);
buf BUF1 (N983, N980);
or OR3 (N984, N975, N711, N136);
and AND4 (N985, N978, N689, N662, N38);
nand NAND2 (N986, N973, N653);
not NOT1 (N987, N985);
nor NOR2 (N988, N976, N939);
nand NAND4 (N989, N977, N784, N689, N247);
xor XOR2 (N990, N988, N782);
or OR4 (N991, N987, N278, N142, N797);
not NOT1 (N992, N982);
buf BUF1 (N993, N990);
and AND3 (N994, N984, N689, N598);
nand NAND3 (N995, N983, N916, N212);
or OR4 (N996, N994, N432, N178, N236);
not NOT1 (N997, N986);
nor NOR4 (N998, N997, N67, N817, N587);
buf BUF1 (N999, N979);
not NOT1 (N1000, N989);
and AND4 (N1001, N993, N490, N279, N17);
xor XOR2 (N1002, N992, N805);
nand NAND3 (N1003, N1001, N232, N978);
nor NOR4 (N1004, N964, N788, N996, N825);
nand NAND4 (N1005, N105, N703, N204, N32);
or OR4 (N1006, N1004, N818, N709, N806);
not NOT1 (N1007, N995);
nor NOR3 (N1008, N1000, N674, N244);
or OR4 (N1009, N991, N941, N187, N617);
nand NAND4 (N1010, N1002, N800, N683, N249);
xor XOR2 (N1011, N981, N835);
nor NOR4 (N1012, N1011, N991, N378, N501);
not NOT1 (N1013, N1009);
xor XOR2 (N1014, N1010, N419);
not NOT1 (N1015, N1008);
nor NOR3 (N1016, N1005, N155, N630);
and AND2 (N1017, N1014, N277);
not NOT1 (N1018, N1007);
or OR2 (N1019, N1012, N544);
nand NAND2 (N1020, N1016, N553);
xor XOR2 (N1021, N1006, N914);
and AND2 (N1022, N1013, N174);
not NOT1 (N1023, N1019);
or OR4 (N1024, N999, N534, N207, N745);
nor NOR4 (N1025, N1017, N17, N176, N609);
buf BUF1 (N1026, N1024);
xor XOR2 (N1027, N1022, N387);
nand NAND3 (N1028, N1021, N372, N24);
and AND2 (N1029, N1003, N963);
and AND4 (N1030, N1026, N44, N799, N1014);
not NOT1 (N1031, N1015);
buf BUF1 (N1032, N1031);
not NOT1 (N1033, N1032);
or OR3 (N1034, N1028, N334, N591);
buf BUF1 (N1035, N1034);
not NOT1 (N1036, N1033);
or OR2 (N1037, N1027, N359);
and AND2 (N1038, N1018, N440);
nor NOR3 (N1039, N1038, N169, N433);
buf BUF1 (N1040, N1036);
or OR4 (N1041, N1025, N643, N831, N460);
nand NAND4 (N1042, N1023, N483, N740, N616);
nor NOR2 (N1043, N1039, N583);
nand NAND4 (N1044, N1029, N611, N344, N875);
or OR3 (N1045, N1035, N911, N753);
buf BUF1 (N1046, N1037);
or OR2 (N1047, N1040, N260);
not NOT1 (N1048, N1045);
or OR3 (N1049, N1020, N451, N859);
or OR4 (N1050, N1048, N370, N924, N667);
nand NAND2 (N1051, N1041, N18);
nand NAND4 (N1052, N1046, N684, N462, N180);
nand NAND3 (N1053, N1052, N180, N204);
nand NAND2 (N1054, N998, N873);
not NOT1 (N1055, N1053);
not NOT1 (N1056, N1047);
and AND3 (N1057, N1049, N442, N325);
xor XOR2 (N1058, N1043, N143);
and AND4 (N1059, N1057, N135, N549, N937);
buf BUF1 (N1060, N1054);
buf BUF1 (N1061, N1044);
and AND2 (N1062, N1030, N426);
and AND2 (N1063, N1056, N538);
xor XOR2 (N1064, N1042, N298);
nor NOR2 (N1065, N1063, N507);
or OR3 (N1066, N1061, N976, N920);
and AND2 (N1067, N1051, N766);
or OR4 (N1068, N1067, N66, N786, N526);
or OR4 (N1069, N1064, N1054, N846, N347);
nor NOR3 (N1070, N1058, N1049, N656);
or OR3 (N1071, N1065, N428, N507);
nor NOR4 (N1072, N1050, N817, N785, N925);
or OR2 (N1073, N1069, N393);
not NOT1 (N1074, N1068);
or OR2 (N1075, N1066, N404);
or OR3 (N1076, N1055, N679, N708);
nor NOR2 (N1077, N1059, N672);
nand NAND2 (N1078, N1071, N545);
nand NAND4 (N1079, N1070, N877, N971, N326);
buf BUF1 (N1080, N1079);
or OR4 (N1081, N1078, N1035, N211, N105);
xor XOR2 (N1082, N1062, N254);
buf BUF1 (N1083, N1082);
xor XOR2 (N1084, N1080, N849);
buf BUF1 (N1085, N1081);
xor XOR2 (N1086, N1077, N27);
nand NAND4 (N1087, N1072, N562, N697, N947);
not NOT1 (N1088, N1074);
nand NAND2 (N1089, N1083, N964);
and AND4 (N1090, N1089, N71, N637, N607);
buf BUF1 (N1091, N1090);
nand NAND2 (N1092, N1060, N595);
nand NAND4 (N1093, N1076, N778, N127, N813);
and AND3 (N1094, N1091, N631, N11);
or OR2 (N1095, N1092, N846);
xor XOR2 (N1096, N1088, N1022);
not NOT1 (N1097, N1087);
nor NOR3 (N1098, N1097, N268, N138);
buf BUF1 (N1099, N1086);
xor XOR2 (N1100, N1094, N47);
nor NOR2 (N1101, N1098, N888);
and AND2 (N1102, N1075, N804);
and AND4 (N1103, N1095, N993, N116, N326);
and AND3 (N1104, N1102, N856, N686);
nor NOR3 (N1105, N1093, N93, N166);
not NOT1 (N1106, N1103);
xor XOR2 (N1107, N1073, N927);
not NOT1 (N1108, N1085);
not NOT1 (N1109, N1099);
xor XOR2 (N1110, N1084, N689);
xor XOR2 (N1111, N1105, N954);
not NOT1 (N1112, N1111);
and AND4 (N1113, N1101, N762, N231, N1047);
nand NAND2 (N1114, N1108, N755);
buf BUF1 (N1115, N1114);
xor XOR2 (N1116, N1115, N983);
nand NAND4 (N1117, N1104, N897, N203, N816);
or OR2 (N1118, N1106, N217);
nand NAND4 (N1119, N1109, N414, N181, N553);
not NOT1 (N1120, N1118);
or OR2 (N1121, N1107, N636);
buf BUF1 (N1122, N1096);
and AND2 (N1123, N1110, N1003);
nand NAND3 (N1124, N1112, N1112, N1078);
not NOT1 (N1125, N1122);
or OR3 (N1126, N1124, N477, N1123);
nor NOR3 (N1127, N689, N134, N681);
and AND3 (N1128, N1100, N114, N1057);
or OR2 (N1129, N1127, N589);
buf BUF1 (N1130, N1119);
and AND3 (N1131, N1126, N548, N325);
or OR4 (N1132, N1130, N430, N773, N892);
buf BUF1 (N1133, N1121);
not NOT1 (N1134, N1113);
nor NOR3 (N1135, N1131, N348, N350);
and AND2 (N1136, N1129, N931);
nor NOR2 (N1137, N1134, N1017);
and AND3 (N1138, N1120, N686, N772);
buf BUF1 (N1139, N1137);
or OR4 (N1140, N1125, N852, N52, N643);
nand NAND3 (N1141, N1139, N226, N70);
nor NOR3 (N1142, N1128, N664, N676);
xor XOR2 (N1143, N1140, N528);
buf BUF1 (N1144, N1141);
or OR3 (N1145, N1116, N990, N165);
nand NAND4 (N1146, N1138, N1130, N465, N1015);
or OR3 (N1147, N1143, N776, N413);
nor NOR4 (N1148, N1135, N64, N297, N63);
nor NOR3 (N1149, N1145, N218, N864);
or OR2 (N1150, N1146, N456);
and AND3 (N1151, N1149, N945, N1087);
xor XOR2 (N1152, N1142, N1069);
not NOT1 (N1153, N1144);
not NOT1 (N1154, N1148);
not NOT1 (N1155, N1117);
buf BUF1 (N1156, N1150);
buf BUF1 (N1157, N1152);
not NOT1 (N1158, N1156);
buf BUF1 (N1159, N1151);
nor NOR4 (N1160, N1133, N330, N1025, N984);
xor XOR2 (N1161, N1132, N6);
or OR3 (N1162, N1161, N20, N637);
not NOT1 (N1163, N1157);
xor XOR2 (N1164, N1155, N659);
and AND3 (N1165, N1136, N778, N45);
nor NOR3 (N1166, N1164, N287, N167);
nor NOR4 (N1167, N1165, N301, N673, N1090);
xor XOR2 (N1168, N1158, N381);
buf BUF1 (N1169, N1154);
nor NOR3 (N1170, N1153, N212, N704);
nand NAND4 (N1171, N1169, N710, N950, N118);
and AND4 (N1172, N1166, N339, N578, N11);
buf BUF1 (N1173, N1167);
or OR2 (N1174, N1163, N234);
nand NAND3 (N1175, N1159, N1082, N868);
or OR3 (N1176, N1171, N1079, N459);
xor XOR2 (N1177, N1175, N204);
nor NOR4 (N1178, N1172, N679, N970, N954);
nor NOR3 (N1179, N1178, N662, N692);
or OR3 (N1180, N1168, N762, N1081);
not NOT1 (N1181, N1147);
or OR3 (N1182, N1160, N984, N130);
nand NAND2 (N1183, N1174, N796);
nor NOR2 (N1184, N1182, N426);
and AND4 (N1185, N1183, N176, N883, N22);
nor NOR4 (N1186, N1180, N376, N960, N1025);
buf BUF1 (N1187, N1173);
nand NAND4 (N1188, N1162, N671, N291, N335);
nand NAND2 (N1189, N1179, N90);
nand NAND3 (N1190, N1185, N281, N696);
nand NAND2 (N1191, N1189, N247);
and AND3 (N1192, N1177, N603, N60);
or OR2 (N1193, N1191, N86);
buf BUF1 (N1194, N1170);
and AND4 (N1195, N1186, N1054, N1039, N803);
nand NAND2 (N1196, N1190, N522);
nand NAND4 (N1197, N1181, N1171, N103, N108);
or OR4 (N1198, N1187, N49, N887, N456);
or OR3 (N1199, N1192, N785, N123);
nand NAND3 (N1200, N1188, N1186, N521);
not NOT1 (N1201, N1193);
nor NOR4 (N1202, N1199, N1187, N441, N508);
or OR3 (N1203, N1201, N883, N815);
and AND2 (N1204, N1198, N494);
not NOT1 (N1205, N1204);
nand NAND3 (N1206, N1197, N966, N1078);
buf BUF1 (N1207, N1184);
buf BUF1 (N1208, N1203);
buf BUF1 (N1209, N1205);
or OR3 (N1210, N1206, N500, N812);
or OR2 (N1211, N1200, N816);
nor NOR3 (N1212, N1176, N268, N392);
buf BUF1 (N1213, N1209);
or OR2 (N1214, N1211, N1156);
nor NOR4 (N1215, N1202, N572, N869, N312);
xor XOR2 (N1216, N1195, N400);
not NOT1 (N1217, N1212);
and AND2 (N1218, N1208, N358);
nor NOR4 (N1219, N1194, N343, N912, N631);
not NOT1 (N1220, N1217);
nand NAND2 (N1221, N1210, N235);
not NOT1 (N1222, N1214);
and AND3 (N1223, N1220, N342, N1033);
nand NAND2 (N1224, N1216, N673);
or OR2 (N1225, N1207, N1174);
and AND4 (N1226, N1224, N689, N24, N1157);
or OR2 (N1227, N1215, N850);
nand NAND4 (N1228, N1225, N411, N1000, N1060);
nand NAND3 (N1229, N1219, N12, N572);
or OR2 (N1230, N1229, N631);
buf BUF1 (N1231, N1230);
xor XOR2 (N1232, N1222, N725);
nor NOR2 (N1233, N1223, N369);
nand NAND3 (N1234, N1213, N132, N1146);
not NOT1 (N1235, N1228);
or OR3 (N1236, N1226, N153, N514);
buf BUF1 (N1237, N1196);
or OR3 (N1238, N1236, N672, N100);
and AND3 (N1239, N1227, N70, N350);
xor XOR2 (N1240, N1234, N379);
buf BUF1 (N1241, N1221);
nor NOR4 (N1242, N1231, N1175, N515, N687);
not NOT1 (N1243, N1242);
xor XOR2 (N1244, N1243, N1064);
xor XOR2 (N1245, N1218, N382);
not NOT1 (N1246, N1241);
or OR2 (N1247, N1246, N749);
nand NAND3 (N1248, N1232, N955, N400);
not NOT1 (N1249, N1244);
or OR4 (N1250, N1240, N614, N423, N591);
and AND2 (N1251, N1249, N736);
nand NAND3 (N1252, N1251, N835, N310);
not NOT1 (N1253, N1237);
nor NOR4 (N1254, N1250, N603, N730, N735);
or OR2 (N1255, N1253, N19);
and AND4 (N1256, N1233, N475, N519, N602);
and AND2 (N1257, N1252, N251);
not NOT1 (N1258, N1238);
nor NOR4 (N1259, N1248, N366, N978, N713);
buf BUF1 (N1260, N1247);
not NOT1 (N1261, N1256);
not NOT1 (N1262, N1235);
buf BUF1 (N1263, N1262);
and AND2 (N1264, N1245, N304);
not NOT1 (N1265, N1255);
or OR3 (N1266, N1259, N127, N847);
buf BUF1 (N1267, N1265);
and AND4 (N1268, N1267, N235, N989, N587);
and AND4 (N1269, N1254, N88, N1175, N1025);
buf BUF1 (N1270, N1268);
and AND2 (N1271, N1258, N155);
xor XOR2 (N1272, N1260, N304);
xor XOR2 (N1273, N1263, N300);
not NOT1 (N1274, N1273);
nand NAND2 (N1275, N1271, N247);
xor XOR2 (N1276, N1264, N704);
buf BUF1 (N1277, N1269);
or OR4 (N1278, N1274, N13, N353, N693);
buf BUF1 (N1279, N1266);
or OR3 (N1280, N1272, N466, N656);
buf BUF1 (N1281, N1279);
buf BUF1 (N1282, N1276);
and AND2 (N1283, N1282, N377);
xor XOR2 (N1284, N1277, N163);
buf BUF1 (N1285, N1281);
buf BUF1 (N1286, N1261);
buf BUF1 (N1287, N1286);
and AND3 (N1288, N1285, N857, N1140);
xor XOR2 (N1289, N1278, N803);
buf BUF1 (N1290, N1257);
not NOT1 (N1291, N1283);
not NOT1 (N1292, N1270);
xor XOR2 (N1293, N1289, N847);
or OR4 (N1294, N1291, N891, N102, N1211);
xor XOR2 (N1295, N1239, N360);
nor NOR4 (N1296, N1295, N737, N1226, N440);
and AND3 (N1297, N1287, N408, N660);
not NOT1 (N1298, N1284);
nand NAND2 (N1299, N1290, N332);
buf BUF1 (N1300, N1275);
not NOT1 (N1301, N1300);
xor XOR2 (N1302, N1296, N345);
and AND3 (N1303, N1298, N724, N197);
nand NAND3 (N1304, N1293, N1001, N444);
or OR2 (N1305, N1299, N299);
nand NAND4 (N1306, N1305, N190, N1146, N70);
or OR2 (N1307, N1292, N989);
nor NOR4 (N1308, N1297, N554, N827, N180);
and AND4 (N1309, N1304, N550, N534, N7);
or OR3 (N1310, N1306, N1220, N283);
nand NAND3 (N1311, N1288, N691, N674);
or OR3 (N1312, N1311, N727, N999);
nor NOR2 (N1313, N1309, N406);
buf BUF1 (N1314, N1308);
or OR3 (N1315, N1313, N1131, N379);
buf BUF1 (N1316, N1315);
buf BUF1 (N1317, N1310);
nor NOR2 (N1318, N1302, N975);
or OR2 (N1319, N1280, N317);
nand NAND4 (N1320, N1314, N623, N123, N1273);
or OR4 (N1321, N1312, N1291, N200, N868);
buf BUF1 (N1322, N1294);
xor XOR2 (N1323, N1317, N95);
buf BUF1 (N1324, N1303);
not NOT1 (N1325, N1307);
or OR2 (N1326, N1325, N328);
xor XOR2 (N1327, N1319, N4);
nor NOR3 (N1328, N1326, N560, N1056);
nand NAND3 (N1329, N1323, N1102, N871);
nand NAND4 (N1330, N1328, N848, N1099, N773);
not NOT1 (N1331, N1316);
nand NAND2 (N1332, N1318, N443);
and AND4 (N1333, N1301, N14, N1312, N1065);
not NOT1 (N1334, N1329);
or OR2 (N1335, N1324, N1231);
buf BUF1 (N1336, N1331);
nand NAND4 (N1337, N1330, N682, N1217, N272);
not NOT1 (N1338, N1327);
buf BUF1 (N1339, N1322);
xor XOR2 (N1340, N1320, N1178);
or OR2 (N1341, N1339, N1252);
and AND4 (N1342, N1340, N385, N753, N1295);
buf BUF1 (N1343, N1334);
nand NAND4 (N1344, N1321, N812, N1085, N689);
or OR4 (N1345, N1336, N1165, N959, N353);
nand NAND2 (N1346, N1344, N27);
xor XOR2 (N1347, N1333, N897);
nand NAND4 (N1348, N1347, N1111, N36, N821);
nor NOR3 (N1349, N1342, N1198, N403);
or OR4 (N1350, N1346, N1155, N97, N10);
buf BUF1 (N1351, N1343);
nor NOR4 (N1352, N1351, N1226, N1236, N1178);
nor NOR4 (N1353, N1345, N1149, N630, N343);
nand NAND3 (N1354, N1335, N861, N1288);
nand NAND4 (N1355, N1354, N1047, N445, N1217);
nor NOR3 (N1356, N1352, N949, N935);
nand NAND3 (N1357, N1332, N290, N1306);
and AND4 (N1358, N1350, N610, N25, N1015);
nand NAND2 (N1359, N1353, N660);
xor XOR2 (N1360, N1338, N902);
and AND4 (N1361, N1355, N682, N102, N1091);
not NOT1 (N1362, N1349);
nand NAND3 (N1363, N1357, N807, N613);
and AND2 (N1364, N1341, N792);
buf BUF1 (N1365, N1356);
nand NAND4 (N1366, N1348, N639, N594, N690);
nor NOR3 (N1367, N1359, N737, N56);
or OR4 (N1368, N1365, N690, N35, N578);
buf BUF1 (N1369, N1363);
nor NOR3 (N1370, N1362, N1141, N826);
and AND4 (N1371, N1367, N936, N685, N648);
not NOT1 (N1372, N1366);
and AND4 (N1373, N1361, N792, N164, N178);
buf BUF1 (N1374, N1337);
and AND3 (N1375, N1358, N1196, N483);
or OR4 (N1376, N1360, N1019, N1194, N1180);
buf BUF1 (N1377, N1376);
not NOT1 (N1378, N1371);
or OR3 (N1379, N1373, N306, N277);
xor XOR2 (N1380, N1375, N1332);
nand NAND3 (N1381, N1372, N358, N1);
not NOT1 (N1382, N1369);
nand NAND4 (N1383, N1364, N1104, N283, N646);
not NOT1 (N1384, N1381);
buf BUF1 (N1385, N1379);
or OR3 (N1386, N1382, N7, N40);
not NOT1 (N1387, N1386);
nor NOR3 (N1388, N1380, N873, N738);
or OR4 (N1389, N1374, N1314, N2, N1261);
xor XOR2 (N1390, N1377, N952);
and AND2 (N1391, N1387, N1130);
or OR4 (N1392, N1368, N1332, N317, N995);
buf BUF1 (N1393, N1388);
nor NOR4 (N1394, N1389, N547, N310, N606);
nand NAND4 (N1395, N1393, N1379, N1183, N979);
xor XOR2 (N1396, N1391, N83);
buf BUF1 (N1397, N1396);
or OR3 (N1398, N1383, N777, N1270);
buf BUF1 (N1399, N1392);
nor NOR2 (N1400, N1395, N497);
not NOT1 (N1401, N1385);
nand NAND3 (N1402, N1401, N1049, N290);
and AND2 (N1403, N1384, N410);
buf BUF1 (N1404, N1398);
and AND4 (N1405, N1404, N1005, N996, N531);
xor XOR2 (N1406, N1397, N952);
xor XOR2 (N1407, N1405, N74);
nor NOR3 (N1408, N1407, N1336, N458);
nand NAND4 (N1409, N1378, N1313, N677, N860);
nor NOR3 (N1410, N1406, N899, N257);
nor NOR2 (N1411, N1394, N1217);
or OR2 (N1412, N1411, N773);
not NOT1 (N1413, N1399);
nor NOR4 (N1414, N1410, N1330, N895, N491);
xor XOR2 (N1415, N1370, N670);
buf BUF1 (N1416, N1402);
buf BUF1 (N1417, N1413);
and AND3 (N1418, N1417, N428, N907);
buf BUF1 (N1419, N1415);
nand NAND2 (N1420, N1414, N32);
buf BUF1 (N1421, N1418);
and AND4 (N1422, N1420, N1329, N537, N128);
buf BUF1 (N1423, N1390);
nand NAND4 (N1424, N1421, N931, N17, N461);
not NOT1 (N1425, N1409);
not NOT1 (N1426, N1412);
nand NAND2 (N1427, N1424, N421);
not NOT1 (N1428, N1426);
xor XOR2 (N1429, N1422, N729);
xor XOR2 (N1430, N1419, N59);
not NOT1 (N1431, N1428);
xor XOR2 (N1432, N1427, N641);
xor XOR2 (N1433, N1400, N272);
nor NOR2 (N1434, N1433, N420);
nor NOR2 (N1435, N1432, N1427);
xor XOR2 (N1436, N1435, N860);
nand NAND3 (N1437, N1429, N1116, N1004);
nor NOR3 (N1438, N1431, N926, N615);
buf BUF1 (N1439, N1430);
not NOT1 (N1440, N1434);
buf BUF1 (N1441, N1436);
nand NAND3 (N1442, N1425, N700, N1145);
buf BUF1 (N1443, N1442);
nand NAND4 (N1444, N1416, N1274, N747, N666);
or OR2 (N1445, N1408, N1315);
nor NOR4 (N1446, N1440, N428, N1109, N40);
nand NAND3 (N1447, N1446, N112, N1164);
buf BUF1 (N1448, N1439);
buf BUF1 (N1449, N1444);
or OR3 (N1450, N1403, N787, N878);
or OR3 (N1451, N1423, N796, N1322);
or OR4 (N1452, N1441, N701, N1398, N326);
xor XOR2 (N1453, N1450, N1071);
buf BUF1 (N1454, N1445);
nand NAND3 (N1455, N1449, N324, N1290);
or OR4 (N1456, N1454, N150, N157, N227);
or OR4 (N1457, N1448, N1069, N851, N1099);
not NOT1 (N1458, N1438);
and AND3 (N1459, N1443, N1026, N1264);
buf BUF1 (N1460, N1437);
and AND3 (N1461, N1455, N1322, N866);
and AND3 (N1462, N1457, N690, N1308);
nand NAND2 (N1463, N1452, N156);
nor NOR4 (N1464, N1461, N919, N1208, N576);
nand NAND4 (N1465, N1459, N1160, N828, N881);
or OR2 (N1466, N1458, N1422);
not NOT1 (N1467, N1456);
xor XOR2 (N1468, N1462, N458);
buf BUF1 (N1469, N1447);
xor XOR2 (N1470, N1467, N45);
xor XOR2 (N1471, N1468, N814);
and AND4 (N1472, N1469, N601, N472, N306);
and AND2 (N1473, N1470, N756);
not NOT1 (N1474, N1471);
nand NAND4 (N1475, N1465, N333, N1327, N1429);
not NOT1 (N1476, N1475);
nand NAND3 (N1477, N1453, N74, N1377);
buf BUF1 (N1478, N1474);
buf BUF1 (N1479, N1476);
nand NAND3 (N1480, N1477, N1301, N1454);
buf BUF1 (N1481, N1472);
and AND4 (N1482, N1473, N717, N167, N741);
xor XOR2 (N1483, N1463, N216);
not NOT1 (N1484, N1466);
xor XOR2 (N1485, N1479, N1343);
xor XOR2 (N1486, N1482, N776);
nor NOR3 (N1487, N1483, N1357, N573);
xor XOR2 (N1488, N1485, N155);
buf BUF1 (N1489, N1460);
nand NAND2 (N1490, N1486, N27);
nor NOR4 (N1491, N1488, N2, N432, N1218);
nor NOR2 (N1492, N1489, N113);
buf BUF1 (N1493, N1464);
nor NOR4 (N1494, N1487, N561, N253, N765);
nand NAND4 (N1495, N1490, N313, N359, N680);
not NOT1 (N1496, N1495);
nand NAND3 (N1497, N1451, N939, N913);
and AND3 (N1498, N1492, N919, N1135);
buf BUF1 (N1499, N1481);
not NOT1 (N1500, N1484);
buf BUF1 (N1501, N1497);
and AND3 (N1502, N1491, N1118, N396);
or OR4 (N1503, N1500, N368, N167, N881);
nor NOR2 (N1504, N1502, N1314);
and AND2 (N1505, N1480, N1342);
buf BUF1 (N1506, N1498);
not NOT1 (N1507, N1506);
nand NAND3 (N1508, N1503, N1177, N150);
or OR2 (N1509, N1499, N968);
or OR2 (N1510, N1478, N1053);
buf BUF1 (N1511, N1507);
nand NAND4 (N1512, N1496, N1263, N797, N201);
buf BUF1 (N1513, N1504);
nand NAND2 (N1514, N1512, N579);
or OR4 (N1515, N1510, N117, N249, N101);
not NOT1 (N1516, N1509);
not NOT1 (N1517, N1493);
not NOT1 (N1518, N1508);
xor XOR2 (N1519, N1501, N603);
xor XOR2 (N1520, N1517, N627);
not NOT1 (N1521, N1505);
nor NOR3 (N1522, N1520, N838, N1482);
or OR2 (N1523, N1511, N978);
nor NOR2 (N1524, N1521, N653);
and AND2 (N1525, N1514, N1073);
xor XOR2 (N1526, N1523, N900);
nand NAND2 (N1527, N1525, N935);
nor NOR4 (N1528, N1526, N127, N1291, N751);
buf BUF1 (N1529, N1524);
or OR2 (N1530, N1527, N760);
nand NAND2 (N1531, N1513, N902);
or OR2 (N1532, N1518, N1046);
nor NOR3 (N1533, N1529, N1094, N916);
buf BUF1 (N1534, N1532);
xor XOR2 (N1535, N1494, N1138);
xor XOR2 (N1536, N1534, N1327);
xor XOR2 (N1537, N1531, N259);
and AND3 (N1538, N1533, N1132, N1233);
buf BUF1 (N1539, N1516);
nand NAND2 (N1540, N1536, N455);
or OR4 (N1541, N1540, N1370, N1103, N117);
buf BUF1 (N1542, N1519);
and AND3 (N1543, N1542, N564, N1288);
and AND4 (N1544, N1541, N584, N358, N320);
nor NOR2 (N1545, N1528, N743);
nor NOR2 (N1546, N1543, N262);
and AND2 (N1547, N1538, N1119);
xor XOR2 (N1548, N1545, N185);
and AND4 (N1549, N1544, N491, N571, N147);
nand NAND3 (N1550, N1548, N367, N57);
xor XOR2 (N1551, N1550, N552);
xor XOR2 (N1552, N1515, N506);
and AND4 (N1553, N1547, N1472, N642, N1464);
nor NOR4 (N1554, N1535, N718, N398, N326);
not NOT1 (N1555, N1537);
xor XOR2 (N1556, N1546, N811);
nand NAND3 (N1557, N1552, N321, N29);
nor NOR3 (N1558, N1556, N935, N341);
or OR3 (N1559, N1553, N1034, N1550);
or OR4 (N1560, N1551, N727, N1041, N952);
and AND3 (N1561, N1549, N453, N326);
not NOT1 (N1562, N1554);
or OR2 (N1563, N1558, N380);
nand NAND3 (N1564, N1539, N265, N35);
or OR4 (N1565, N1557, N1462, N472, N27);
or OR4 (N1566, N1564, N127, N1503, N1456);
not NOT1 (N1567, N1559);
nor NOR4 (N1568, N1563, N670, N1431, N1326);
buf BUF1 (N1569, N1530);
not NOT1 (N1570, N1568);
buf BUF1 (N1571, N1555);
nand NAND3 (N1572, N1560, N263, N871);
and AND4 (N1573, N1569, N997, N5, N340);
not NOT1 (N1574, N1562);
not NOT1 (N1575, N1565);
not NOT1 (N1576, N1574);
not NOT1 (N1577, N1573);
and AND3 (N1578, N1575, N223, N749);
nor NOR3 (N1579, N1522, N152, N1255);
nand NAND4 (N1580, N1571, N155, N133, N75);
buf BUF1 (N1581, N1579);
not NOT1 (N1582, N1566);
and AND4 (N1583, N1572, N1309, N650, N1096);
xor XOR2 (N1584, N1582, N700);
buf BUF1 (N1585, N1583);
xor XOR2 (N1586, N1581, N649);
nor NOR3 (N1587, N1578, N457, N1078);
not NOT1 (N1588, N1561);
and AND3 (N1589, N1584, N41, N199);
nor NOR4 (N1590, N1588, N410, N246, N1141);
and AND3 (N1591, N1590, N812, N305);
and AND3 (N1592, N1587, N284, N666);
and AND3 (N1593, N1577, N1546, N13);
or OR4 (N1594, N1593, N546, N1050, N766);
nand NAND2 (N1595, N1591, N1284);
nor NOR3 (N1596, N1570, N1562, N775);
nor NOR2 (N1597, N1576, N857);
and AND3 (N1598, N1580, N420, N365);
or OR2 (N1599, N1598, N188);
nor NOR2 (N1600, N1567, N289);
nand NAND4 (N1601, N1599, N1125, N61, N1431);
nor NOR3 (N1602, N1595, N999, N1059);
and AND4 (N1603, N1601, N38, N937, N878);
nand NAND3 (N1604, N1592, N623, N78);
nor NOR2 (N1605, N1600, N1480);
xor XOR2 (N1606, N1597, N628);
buf BUF1 (N1607, N1586);
or OR2 (N1608, N1603, N132);
buf BUF1 (N1609, N1596);
xor XOR2 (N1610, N1609, N1114);
or OR3 (N1611, N1604, N702, N1448);
nor NOR3 (N1612, N1585, N781, N346);
or OR3 (N1613, N1606, N662, N585);
nand NAND4 (N1614, N1605, N284, N531, N1407);
and AND4 (N1615, N1612, N259, N568, N474);
xor XOR2 (N1616, N1610, N1162);
not NOT1 (N1617, N1594);
not NOT1 (N1618, N1617);
buf BUF1 (N1619, N1615);
and AND2 (N1620, N1619, N1554);
not NOT1 (N1621, N1608);
not NOT1 (N1622, N1602);
not NOT1 (N1623, N1618);
buf BUF1 (N1624, N1589);
buf BUF1 (N1625, N1620);
xor XOR2 (N1626, N1623, N62);
or OR4 (N1627, N1614, N600, N111, N516);
and AND2 (N1628, N1625, N1110);
nor NOR4 (N1629, N1622, N1553, N928, N1021);
not NOT1 (N1630, N1628);
nand NAND4 (N1631, N1629, N1174, N623, N1311);
and AND2 (N1632, N1621, N1098);
nor NOR2 (N1633, N1616, N1281);
and AND2 (N1634, N1633, N820);
nor NOR2 (N1635, N1624, N1382);
not NOT1 (N1636, N1607);
not NOT1 (N1637, N1634);
not NOT1 (N1638, N1626);
or OR3 (N1639, N1611, N918, N519);
xor XOR2 (N1640, N1639, N1155);
buf BUF1 (N1641, N1631);
nor NOR2 (N1642, N1641, N632);
or OR4 (N1643, N1630, N1123, N556, N41);
xor XOR2 (N1644, N1635, N1001);
buf BUF1 (N1645, N1627);
nor NOR2 (N1646, N1637, N546);
or OR3 (N1647, N1646, N48, N901);
nor NOR3 (N1648, N1643, N578, N58);
nand NAND2 (N1649, N1648, N839);
xor XOR2 (N1650, N1649, N281);
xor XOR2 (N1651, N1638, N1221);
and AND4 (N1652, N1644, N1042, N742, N27);
buf BUF1 (N1653, N1640);
nor NOR3 (N1654, N1650, N1141, N1320);
not NOT1 (N1655, N1645);
xor XOR2 (N1656, N1647, N1596);
buf BUF1 (N1657, N1655);
nand NAND2 (N1658, N1653, N511);
or OR4 (N1659, N1651, N113, N1329, N77);
nand NAND4 (N1660, N1652, N435, N87, N964);
xor XOR2 (N1661, N1654, N892);
xor XOR2 (N1662, N1659, N1218);
buf BUF1 (N1663, N1660);
xor XOR2 (N1664, N1661, N1565);
nand NAND4 (N1665, N1657, N940, N507, N1129);
not NOT1 (N1666, N1664);
not NOT1 (N1667, N1656);
nor NOR2 (N1668, N1667, N548);
xor XOR2 (N1669, N1666, N294);
nand NAND3 (N1670, N1663, N818, N5);
nor NOR2 (N1671, N1669, N354);
not NOT1 (N1672, N1671);
nand NAND3 (N1673, N1636, N1169, N569);
not NOT1 (N1674, N1632);
and AND4 (N1675, N1672, N1249, N702, N1030);
and AND4 (N1676, N1665, N865, N946, N362);
nand NAND2 (N1677, N1642, N365);
buf BUF1 (N1678, N1674);
nor NOR4 (N1679, N1662, N158, N823, N1622);
nor NOR4 (N1680, N1679, N9, N1009, N27);
xor XOR2 (N1681, N1677, N26);
not NOT1 (N1682, N1675);
not NOT1 (N1683, N1668);
and AND2 (N1684, N1673, N802);
and AND3 (N1685, N1682, N657, N1490);
xor XOR2 (N1686, N1680, N1320);
not NOT1 (N1687, N1681);
buf BUF1 (N1688, N1676);
not NOT1 (N1689, N1687);
nor NOR2 (N1690, N1683, N997);
and AND2 (N1691, N1670, N482);
buf BUF1 (N1692, N1686);
and AND2 (N1693, N1689, N108);
buf BUF1 (N1694, N1690);
nor NOR2 (N1695, N1694, N1521);
nor NOR2 (N1696, N1613, N1612);
buf BUF1 (N1697, N1691);
buf BUF1 (N1698, N1685);
not NOT1 (N1699, N1658);
nand NAND3 (N1700, N1678, N1268, N47);
not NOT1 (N1701, N1688);
not NOT1 (N1702, N1696);
nand NAND4 (N1703, N1700, N459, N1666, N1376);
buf BUF1 (N1704, N1697);
nor NOR2 (N1705, N1701, N1282);
nor NOR3 (N1706, N1705, N170, N1344);
or OR3 (N1707, N1706, N843, N1166);
buf BUF1 (N1708, N1693);
xor XOR2 (N1709, N1699, N1366);
buf BUF1 (N1710, N1702);
not NOT1 (N1711, N1695);
or OR2 (N1712, N1704, N270);
and AND2 (N1713, N1708, N246);
xor XOR2 (N1714, N1711, N164);
not NOT1 (N1715, N1710);
buf BUF1 (N1716, N1714);
and AND3 (N1717, N1703, N1587, N650);
not NOT1 (N1718, N1684);
or OR4 (N1719, N1715, N1046, N643, N557);
nand NAND3 (N1720, N1718, N903, N394);
buf BUF1 (N1721, N1717);
buf BUF1 (N1722, N1719);
not NOT1 (N1723, N1707);
nand NAND4 (N1724, N1723, N717, N1313, N900);
buf BUF1 (N1725, N1724);
or OR3 (N1726, N1716, N963, N487);
xor XOR2 (N1727, N1698, N1037);
nor NOR3 (N1728, N1725, N1194, N1628);
buf BUF1 (N1729, N1692);
nor NOR3 (N1730, N1712, N936, N1050);
not NOT1 (N1731, N1728);
nand NAND4 (N1732, N1709, N1654, N1138, N685);
buf BUF1 (N1733, N1726);
and AND3 (N1734, N1727, N1286, N1600);
xor XOR2 (N1735, N1733, N712);
nand NAND4 (N1736, N1722, N990, N270, N1631);
not NOT1 (N1737, N1729);
xor XOR2 (N1738, N1720, N1317);
xor XOR2 (N1739, N1737, N46);
buf BUF1 (N1740, N1730);
nor NOR2 (N1741, N1735, N889);
not NOT1 (N1742, N1741);
and AND3 (N1743, N1739, N1640, N538);
nand NAND3 (N1744, N1736, N1328, N748);
and AND4 (N1745, N1731, N1076, N866, N907);
xor XOR2 (N1746, N1740, N1006);
and AND4 (N1747, N1746, N1152, N517, N1042);
or OR3 (N1748, N1721, N1156, N1646);
nor NOR3 (N1749, N1734, N1056, N1561);
or OR3 (N1750, N1713, N968, N292);
buf BUF1 (N1751, N1747);
not NOT1 (N1752, N1743);
buf BUF1 (N1753, N1751);
or OR3 (N1754, N1753, N159, N338);
buf BUF1 (N1755, N1732);
nand NAND3 (N1756, N1744, N893, N1473);
buf BUF1 (N1757, N1738);
nand NAND2 (N1758, N1745, N392);
buf BUF1 (N1759, N1754);
not NOT1 (N1760, N1752);
nand NAND4 (N1761, N1755, N318, N1608, N1315);
not NOT1 (N1762, N1749);
not NOT1 (N1763, N1748);
and AND3 (N1764, N1742, N463, N132);
buf BUF1 (N1765, N1763);
or OR3 (N1766, N1758, N1713, N1438);
nand NAND3 (N1767, N1765, N1448, N150);
buf BUF1 (N1768, N1750);
nand NAND4 (N1769, N1760, N1004, N1383, N917);
nand NAND3 (N1770, N1759, N1447, N448);
buf BUF1 (N1771, N1762);
buf BUF1 (N1772, N1757);
or OR2 (N1773, N1767, N1314);
xor XOR2 (N1774, N1756, N48);
nor NOR4 (N1775, N1761, N1604, N550, N134);
nand NAND2 (N1776, N1764, N838);
and AND2 (N1777, N1769, N48);
buf BUF1 (N1778, N1768);
not NOT1 (N1779, N1774);
not NOT1 (N1780, N1777);
nor NOR4 (N1781, N1779, N1197, N1564, N543);
xor XOR2 (N1782, N1766, N1186);
buf BUF1 (N1783, N1781);
nand NAND2 (N1784, N1773, N854);
xor XOR2 (N1785, N1776, N497);
or OR2 (N1786, N1785, N70);
not NOT1 (N1787, N1778);
not NOT1 (N1788, N1775);
or OR2 (N1789, N1770, N691);
nand NAND2 (N1790, N1771, N925);
nor NOR3 (N1791, N1789, N1506, N1157);
nand NAND3 (N1792, N1790, N974, N740);
or OR4 (N1793, N1786, N295, N1483, N715);
and AND4 (N1794, N1780, N698, N758, N19);
not NOT1 (N1795, N1791);
and AND4 (N1796, N1783, N999, N438, N1552);
not NOT1 (N1797, N1784);
or OR4 (N1798, N1796, N1132, N579, N98);
or OR4 (N1799, N1798, N305, N241, N901);
xor XOR2 (N1800, N1797, N1613);
and AND2 (N1801, N1799, N357);
buf BUF1 (N1802, N1793);
nor NOR2 (N1803, N1801, N45);
nand NAND4 (N1804, N1802, N795, N687, N1300);
and AND2 (N1805, N1772, N958);
or OR4 (N1806, N1788, N1196, N1596, N827);
xor XOR2 (N1807, N1804, N1036);
nand NAND2 (N1808, N1782, N1239);
not NOT1 (N1809, N1800);
xor XOR2 (N1810, N1792, N161);
or OR4 (N1811, N1807, N1655, N68, N1667);
nor NOR2 (N1812, N1809, N360);
buf BUF1 (N1813, N1795);
nand NAND3 (N1814, N1787, N1198, N387);
nor NOR4 (N1815, N1808, N910, N713, N453);
or OR3 (N1816, N1805, N1149, N1108);
and AND3 (N1817, N1816, N381, N483);
buf BUF1 (N1818, N1817);
or OR2 (N1819, N1810, N254);
or OR2 (N1820, N1813, N433);
nand NAND2 (N1821, N1803, N1438);
and AND2 (N1822, N1812, N398);
nor NOR2 (N1823, N1814, N46);
buf BUF1 (N1824, N1819);
nand NAND3 (N1825, N1823, N1764, N740);
or OR3 (N1826, N1794, N656, N897);
buf BUF1 (N1827, N1822);
nor NOR4 (N1828, N1825, N434, N1608, N1550);
nor NOR2 (N1829, N1827, N106);
and AND3 (N1830, N1829, N722, N185);
not NOT1 (N1831, N1828);
and AND4 (N1832, N1811, N1227, N322, N557);
xor XOR2 (N1833, N1824, N983);
buf BUF1 (N1834, N1833);
xor XOR2 (N1835, N1821, N295);
xor XOR2 (N1836, N1834, N1091);
or OR4 (N1837, N1818, N1464, N969, N1804);
buf BUF1 (N1838, N1835);
xor XOR2 (N1839, N1820, N1789);
nor NOR2 (N1840, N1836, N189);
nor NOR4 (N1841, N1839, N864, N610, N1352);
buf BUF1 (N1842, N1840);
not NOT1 (N1843, N1842);
buf BUF1 (N1844, N1806);
nor NOR3 (N1845, N1844, N713, N1142);
or OR2 (N1846, N1831, N173);
nor NOR3 (N1847, N1837, N687, N776);
xor XOR2 (N1848, N1847, N1580);
xor XOR2 (N1849, N1843, N1153);
nor NOR3 (N1850, N1849, N1558, N1339);
not NOT1 (N1851, N1841);
nand NAND2 (N1852, N1845, N1847);
or OR4 (N1853, N1846, N70, N307, N1233);
nand NAND2 (N1854, N1832, N102);
nand NAND2 (N1855, N1848, N1041);
or OR3 (N1856, N1854, N576, N505);
xor XOR2 (N1857, N1855, N1198);
not NOT1 (N1858, N1838);
and AND3 (N1859, N1830, N1772, N125);
or OR3 (N1860, N1858, N1729, N509);
nor NOR3 (N1861, N1850, N15, N1644);
nand NAND4 (N1862, N1859, N529, N1144, N1360);
xor XOR2 (N1863, N1860, N454);
nor NOR2 (N1864, N1856, N1107);
or OR3 (N1865, N1851, N1447, N1752);
buf BUF1 (N1866, N1865);
xor XOR2 (N1867, N1863, N798);
and AND3 (N1868, N1862, N793, N1499);
nor NOR2 (N1869, N1815, N181);
nand NAND3 (N1870, N1866, N1015, N1769);
buf BUF1 (N1871, N1826);
or OR4 (N1872, N1864, N1160, N326, N1395);
buf BUF1 (N1873, N1871);
or OR4 (N1874, N1870, N415, N178, N1370);
and AND3 (N1875, N1861, N173, N410);
not NOT1 (N1876, N1868);
nand NAND3 (N1877, N1874, N1039, N1065);
buf BUF1 (N1878, N1852);
and AND4 (N1879, N1876, N1360, N90, N1737);
or OR4 (N1880, N1877, N1495, N408, N1192);
nand NAND3 (N1881, N1879, N709, N442);
not NOT1 (N1882, N1873);
and AND2 (N1883, N1857, N407);
or OR2 (N1884, N1883, N404);
and AND2 (N1885, N1880, N1318);
xor XOR2 (N1886, N1884, N1689);
xor XOR2 (N1887, N1867, N412);
nor NOR3 (N1888, N1853, N428, N153);
not NOT1 (N1889, N1878);
not NOT1 (N1890, N1875);
not NOT1 (N1891, N1888);
nand NAND2 (N1892, N1872, N817);
xor XOR2 (N1893, N1890, N210);
xor XOR2 (N1894, N1885, N948);
or OR3 (N1895, N1891, N1149, N1712);
nand NAND3 (N1896, N1882, N1375, N1190);
nor NOR3 (N1897, N1895, N226, N997);
and AND2 (N1898, N1881, N579);
xor XOR2 (N1899, N1898, N1177);
or OR3 (N1900, N1887, N1838, N1174);
buf BUF1 (N1901, N1886);
buf BUF1 (N1902, N1889);
and AND2 (N1903, N1893, N1733);
buf BUF1 (N1904, N1897);
not NOT1 (N1905, N1899);
not NOT1 (N1906, N1903);
not NOT1 (N1907, N1869);
and AND3 (N1908, N1896, N1873, N202);
xor XOR2 (N1909, N1908, N987);
or OR4 (N1910, N1907, N235, N1411, N1488);
or OR3 (N1911, N1902, N1422, N1481);
nand NAND4 (N1912, N1900, N350, N241, N1198);
buf BUF1 (N1913, N1906);
or OR4 (N1914, N1905, N1450, N777, N1186);
nand NAND3 (N1915, N1904, N679, N594);
or OR3 (N1916, N1901, N1457, N514);
or OR2 (N1917, N1913, N402);
or OR4 (N1918, N1909, N49, N498, N458);
nand NAND2 (N1919, N1915, N117);
and AND4 (N1920, N1917, N159, N585, N1128);
or OR2 (N1921, N1911, N1785);
nand NAND2 (N1922, N1910, N447);
xor XOR2 (N1923, N1892, N1766);
or OR4 (N1924, N1914, N538, N1412, N1851);
nand NAND2 (N1925, N1916, N580);
buf BUF1 (N1926, N1923);
not NOT1 (N1927, N1894);
buf BUF1 (N1928, N1926);
xor XOR2 (N1929, N1924, N85);
and AND3 (N1930, N1920, N1155, N447);
xor XOR2 (N1931, N1918, N1713);
xor XOR2 (N1932, N1929, N1048);
not NOT1 (N1933, N1931);
nor NOR2 (N1934, N1922, N193);
or OR3 (N1935, N1925, N95, N1790);
nand NAND3 (N1936, N1919, N1313, N472);
nor NOR2 (N1937, N1933, N1689);
xor XOR2 (N1938, N1930, N1133);
and AND4 (N1939, N1921, N1308, N1584, N900);
buf BUF1 (N1940, N1939);
not NOT1 (N1941, N1912);
nor NOR2 (N1942, N1927, N1593);
or OR3 (N1943, N1928, N1385, N1174);
or OR2 (N1944, N1940, N25);
not NOT1 (N1945, N1938);
nor NOR4 (N1946, N1941, N1944, N1295, N1309);
or OR3 (N1947, N152, N1011, N865);
xor XOR2 (N1948, N1946, N1864);
or OR2 (N1949, N1945, N1460);
buf BUF1 (N1950, N1937);
nand NAND4 (N1951, N1934, N127, N152, N859);
nand NAND2 (N1952, N1935, N1155);
xor XOR2 (N1953, N1952, N1178);
or OR2 (N1954, N1936, N743);
xor XOR2 (N1955, N1950, N611);
and AND4 (N1956, N1942, N45, N835, N839);
nor NOR4 (N1957, N1932, N138, N1058, N550);
nand NAND4 (N1958, N1949, N286, N1601, N985);
or OR2 (N1959, N1956, N821);
and AND2 (N1960, N1948, N484);
or OR2 (N1961, N1943, N1910);
buf BUF1 (N1962, N1959);
and AND2 (N1963, N1958, N854);
nand NAND2 (N1964, N1963, N1804);
nand NAND3 (N1965, N1951, N421, N750);
or OR2 (N1966, N1961, N1043);
xor XOR2 (N1967, N1962, N337);
not NOT1 (N1968, N1947);
not NOT1 (N1969, N1964);
and AND2 (N1970, N1967, N1228);
not NOT1 (N1971, N1960);
buf BUF1 (N1972, N1969);
buf BUF1 (N1973, N1965);
nor NOR3 (N1974, N1972, N47, N549);
xor XOR2 (N1975, N1970, N1027);
and AND2 (N1976, N1973, N499);
xor XOR2 (N1977, N1976, N484);
buf BUF1 (N1978, N1966);
not NOT1 (N1979, N1977);
and AND3 (N1980, N1968, N923, N967);
nor NOR4 (N1981, N1975, N1915, N1954, N564);
buf BUF1 (N1982, N729);
and AND3 (N1983, N1980, N245, N1522);
not NOT1 (N1984, N1957);
nand NAND2 (N1985, N1981, N394);
buf BUF1 (N1986, N1955);
nor NOR4 (N1987, N1985, N1714, N1872, N1117);
or OR4 (N1988, N1983, N397, N1865, N454);
not NOT1 (N1989, N1978);
buf BUF1 (N1990, N1988);
buf BUF1 (N1991, N1986);
or OR3 (N1992, N1991, N1006, N1813);
and AND3 (N1993, N1953, N74, N1005);
nor NOR4 (N1994, N1979, N42, N996, N1613);
nand NAND3 (N1995, N1974, N1501, N1326);
and AND3 (N1996, N1982, N218, N673);
or OR2 (N1997, N1987, N1923);
or OR3 (N1998, N1990, N148, N525);
buf BUF1 (N1999, N1998);
or OR2 (N2000, N1999, N242);
buf BUF1 (N2001, N1992);
xor XOR2 (N2002, N1994, N1913);
nand NAND2 (N2003, N2002, N889);
buf BUF1 (N2004, N1984);
not NOT1 (N2005, N1995);
buf BUF1 (N2006, N2004);
xor XOR2 (N2007, N1989, N438);
nor NOR4 (N2008, N2006, N6, N76, N1411);
not NOT1 (N2009, N2000);
nor NOR4 (N2010, N2008, N1042, N1088, N1484);
and AND2 (N2011, N2009, N1423);
xor XOR2 (N2012, N2011, N2008);
not NOT1 (N2013, N2003);
nor NOR4 (N2014, N2013, N701, N1547, N1595);
xor XOR2 (N2015, N1971, N537);
or OR3 (N2016, N2001, N68, N207);
and AND2 (N2017, N2005, N315);
not NOT1 (N2018, N1996);
buf BUF1 (N2019, N2015);
not NOT1 (N2020, N2018);
not NOT1 (N2021, N2007);
nand NAND3 (N2022, N2017, N1104, N978);
nand NAND2 (N2023, N2010, N1351);
or OR3 (N2024, N2020, N1343, N1830);
buf BUF1 (N2025, N2016);
not NOT1 (N2026, N2021);
and AND3 (N2027, N1993, N461, N599);
nand NAND3 (N2028, N2024, N499, N141);
and AND2 (N2029, N2022, N589);
nand NAND4 (N2030, N2029, N496, N1359, N597);
or OR2 (N2031, N2030, N145);
buf BUF1 (N2032, N2014);
xor XOR2 (N2033, N2028, N306);
nor NOR3 (N2034, N1997, N427, N51);
not NOT1 (N2035, N2033);
xor XOR2 (N2036, N2035, N1555);
xor XOR2 (N2037, N2012, N546);
nor NOR4 (N2038, N2037, N1278, N740, N931);
nand NAND4 (N2039, N2034, N82, N669, N275);
not NOT1 (N2040, N2027);
not NOT1 (N2041, N2031);
xor XOR2 (N2042, N2038, N192);
nor NOR3 (N2043, N2042, N1636, N85);
buf BUF1 (N2044, N2039);
and AND4 (N2045, N2026, N309, N1764, N1870);
nor NOR4 (N2046, N2041, N556, N1857, N655);
nand NAND3 (N2047, N2044, N421, N681);
xor XOR2 (N2048, N2032, N1633);
nand NAND4 (N2049, N2048, N417, N532, N1221);
xor XOR2 (N2050, N2049, N990);
or OR4 (N2051, N2040, N30, N4, N640);
or OR3 (N2052, N2023, N421, N861);
or OR4 (N2053, N2043, N1778, N1257, N1005);
and AND3 (N2054, N2047, N1159, N120);
or OR3 (N2055, N2053, N1362, N424);
and AND3 (N2056, N2045, N932, N10);
nor NOR4 (N2057, N2050, N289, N73, N1455);
xor XOR2 (N2058, N2055, N157);
or OR4 (N2059, N2056, N496, N1191, N438);
nand NAND3 (N2060, N2025, N1401, N1754);
and AND3 (N2061, N2054, N1867, N2048);
or OR2 (N2062, N2061, N1298);
or OR3 (N2063, N2062, N608, N422);
buf BUF1 (N2064, N2046);
or OR4 (N2065, N2019, N1787, N1195, N1104);
xor XOR2 (N2066, N2052, N435);
nand NAND2 (N2067, N2063, N1344);
not NOT1 (N2068, N2065);
or OR4 (N2069, N2067, N142, N859, N1672);
and AND3 (N2070, N2036, N235, N959);
buf BUF1 (N2071, N2051);
or OR3 (N2072, N2069, N1086, N573);
and AND3 (N2073, N2060, N1738, N1411);
buf BUF1 (N2074, N2059);
not NOT1 (N2075, N2071);
nor NOR3 (N2076, N2066, N183, N1524);
xor XOR2 (N2077, N2073, N700);
or OR4 (N2078, N2077, N631, N805, N977);
or OR4 (N2079, N2068, N1608, N2070, N364);
or OR3 (N2080, N299, N1611, N1586);
not NOT1 (N2081, N2076);
nor NOR3 (N2082, N2058, N252, N24);
xor XOR2 (N2083, N2075, N1348);
or OR2 (N2084, N2072, N364);
nand NAND4 (N2085, N2083, N122, N846, N864);
nand NAND2 (N2086, N2085, N1600);
nand NAND4 (N2087, N2079, N231, N717, N728);
xor XOR2 (N2088, N2064, N1735);
buf BUF1 (N2089, N2082);
or OR3 (N2090, N2086, N370, N606);
nand NAND4 (N2091, N2088, N83, N2027, N1147);
not NOT1 (N2092, N2057);
and AND4 (N2093, N2087, N961, N1194, N1061);
not NOT1 (N2094, N2084);
buf BUF1 (N2095, N2094);
nand NAND2 (N2096, N2080, N1496);
or OR2 (N2097, N2093, N625);
buf BUF1 (N2098, N2097);
nor NOR4 (N2099, N2098, N1041, N1912, N2095);
nand NAND2 (N2100, N2037, N1529);
and AND2 (N2101, N2090, N120);
not NOT1 (N2102, N2074);
or OR2 (N2103, N2099, N917);
xor XOR2 (N2104, N2081, N1714);
or OR3 (N2105, N2102, N1699, N2002);
xor XOR2 (N2106, N2096, N1840);
not NOT1 (N2107, N2091);
xor XOR2 (N2108, N2089, N296);
nand NAND2 (N2109, N2107, N285);
buf BUF1 (N2110, N2078);
not NOT1 (N2111, N2100);
xor XOR2 (N2112, N2108, N175);
or OR3 (N2113, N2105, N1857, N1828);
buf BUF1 (N2114, N2110);
nor NOR4 (N2115, N2106, N1155, N768, N884);
xor XOR2 (N2116, N2103, N1460);
xor XOR2 (N2117, N2111, N991);
not NOT1 (N2118, N2101);
xor XOR2 (N2119, N2104, N1531);
and AND2 (N2120, N2109, N965);
xor XOR2 (N2121, N2118, N888);
not NOT1 (N2122, N2092);
not NOT1 (N2123, N2113);
nand NAND4 (N2124, N2121, N755, N436, N1480);
and AND3 (N2125, N2114, N2097, N2064);
and AND3 (N2126, N2116, N1455, N1008);
xor XOR2 (N2127, N2120, N1135);
not NOT1 (N2128, N2123);
nor NOR3 (N2129, N2112, N55, N1867);
xor XOR2 (N2130, N2115, N421);
xor XOR2 (N2131, N2117, N2015);
buf BUF1 (N2132, N2124);
nand NAND3 (N2133, N2130, N132, N1594);
nand NAND4 (N2134, N2128, N1358, N1166, N546);
nand NAND4 (N2135, N2119, N389, N1270, N1588);
not NOT1 (N2136, N2133);
and AND4 (N2137, N2131, N171, N757, N644);
not NOT1 (N2138, N2127);
nor NOR4 (N2139, N2125, N1079, N612, N1553);
xor XOR2 (N2140, N2134, N98);
buf BUF1 (N2141, N2126);
buf BUF1 (N2142, N2136);
not NOT1 (N2143, N2135);
nand NAND2 (N2144, N2140, N1367);
nand NAND3 (N2145, N2129, N768, N752);
not NOT1 (N2146, N2137);
nand NAND4 (N2147, N2122, N373, N1415, N817);
nor NOR2 (N2148, N2132, N1505);
buf BUF1 (N2149, N2145);
buf BUF1 (N2150, N2144);
or OR4 (N2151, N2146, N1102, N217, N833);
or OR2 (N2152, N2149, N134);
xor XOR2 (N2153, N2139, N1255);
nor NOR2 (N2154, N2138, N196);
or OR4 (N2155, N2151, N2132, N1518, N2135);
xor XOR2 (N2156, N2148, N1494);
xor XOR2 (N2157, N2150, N116);
nand NAND4 (N2158, N2142, N532, N568, N412);
nand NAND4 (N2159, N2154, N1460, N1637, N608);
not NOT1 (N2160, N2155);
buf BUF1 (N2161, N2153);
nand NAND3 (N2162, N2159, N282, N674);
xor XOR2 (N2163, N2156, N1211);
nor NOR2 (N2164, N2143, N1688);
nand NAND2 (N2165, N2147, N358);
or OR4 (N2166, N2160, N1566, N45, N890);
nor NOR3 (N2167, N2141, N1333, N838);
nand NAND2 (N2168, N2164, N1036);
not NOT1 (N2169, N2152);
xor XOR2 (N2170, N2168, N693);
xor XOR2 (N2171, N2167, N506);
nor NOR4 (N2172, N2171, N1196, N1986, N1056);
or OR3 (N2173, N2161, N1291, N275);
xor XOR2 (N2174, N2165, N251);
and AND3 (N2175, N2157, N820, N1590);
and AND3 (N2176, N2175, N65, N911);
nand NAND2 (N2177, N2174, N31);
nand NAND3 (N2178, N2176, N525, N248);
nand NAND3 (N2179, N2177, N666, N2018);
xor XOR2 (N2180, N2163, N1477);
buf BUF1 (N2181, N2179);
buf BUF1 (N2182, N2181);
not NOT1 (N2183, N2158);
not NOT1 (N2184, N2183);
buf BUF1 (N2185, N2162);
nand NAND4 (N2186, N2180, N1423, N1347, N656);
xor XOR2 (N2187, N2185, N140);
xor XOR2 (N2188, N2184, N1225);
not NOT1 (N2189, N2182);
or OR4 (N2190, N2166, N1403, N166, N1085);
xor XOR2 (N2191, N2190, N168);
nand NAND2 (N2192, N2178, N840);
buf BUF1 (N2193, N2186);
nand NAND4 (N2194, N2173, N853, N2184, N883);
buf BUF1 (N2195, N2170);
or OR2 (N2196, N2187, N995);
and AND3 (N2197, N2195, N1716, N1540);
nor NOR4 (N2198, N2172, N1484, N1388, N1378);
buf BUF1 (N2199, N2188);
xor XOR2 (N2200, N2189, N1031);
xor XOR2 (N2201, N2197, N514);
not NOT1 (N2202, N2194);
not NOT1 (N2203, N2192);
and AND2 (N2204, N2199, N466);
and AND2 (N2205, N2198, N1090);
or OR2 (N2206, N2200, N814);
xor XOR2 (N2207, N2201, N392);
not NOT1 (N2208, N2205);
and AND3 (N2209, N2202, N2200, N1845);
nand NAND4 (N2210, N2204, N269, N177, N735);
not NOT1 (N2211, N2191);
not NOT1 (N2212, N2169);
not NOT1 (N2213, N2206);
nand NAND3 (N2214, N2210, N405, N502);
buf BUF1 (N2215, N2207);
xor XOR2 (N2216, N2209, N724);
nor NOR3 (N2217, N2215, N848, N1576);
nor NOR4 (N2218, N2196, N1401, N1342, N279);
not NOT1 (N2219, N2211);
and AND4 (N2220, N2208, N583, N343, N1504);
and AND2 (N2221, N2220, N947);
xor XOR2 (N2222, N2213, N1419);
or OR3 (N2223, N2212, N1276, N2056);
buf BUF1 (N2224, N2222);
xor XOR2 (N2225, N2203, N1535);
buf BUF1 (N2226, N2217);
nand NAND3 (N2227, N2223, N1501, N1285);
and AND3 (N2228, N2221, N1205, N1013);
not NOT1 (N2229, N2228);
not NOT1 (N2230, N2193);
xor XOR2 (N2231, N2227, N16);
or OR2 (N2232, N2218, N1367);
buf BUF1 (N2233, N2230);
nand NAND3 (N2234, N2219, N439, N280);
and AND4 (N2235, N2214, N2204, N1988, N738);
and AND4 (N2236, N2234, N1503, N1435, N1160);
nor NOR2 (N2237, N2236, N195);
buf BUF1 (N2238, N2233);
and AND3 (N2239, N2238, N2086, N651);
and AND4 (N2240, N2231, N290, N31, N1439);
nor NOR2 (N2241, N2237, N1079);
and AND2 (N2242, N2240, N719);
xor XOR2 (N2243, N2239, N1341);
buf BUF1 (N2244, N2226);
xor XOR2 (N2245, N2242, N569);
xor XOR2 (N2246, N2235, N12);
buf BUF1 (N2247, N2225);
or OR3 (N2248, N2224, N100, N1396);
buf BUF1 (N2249, N2246);
nand NAND4 (N2250, N2229, N870, N1490, N190);
or OR4 (N2251, N2250, N1077, N679, N1356);
or OR3 (N2252, N2243, N29, N391);
buf BUF1 (N2253, N2216);
xor XOR2 (N2254, N2245, N2120);
xor XOR2 (N2255, N2247, N737);
nand NAND3 (N2256, N2254, N2151, N2077);
and AND2 (N2257, N2244, N304);
nor NOR4 (N2258, N2252, N439, N1279, N31);
not NOT1 (N2259, N2253);
buf BUF1 (N2260, N2241);
buf BUF1 (N2261, N2255);
not NOT1 (N2262, N2259);
nand NAND4 (N2263, N2249, N1736, N986, N789);
or OR4 (N2264, N2256, N864, N1576, N1364);
not NOT1 (N2265, N2260);
nand NAND3 (N2266, N2258, N625, N1158);
nand NAND2 (N2267, N2262, N702);
and AND4 (N2268, N2232, N1211, N1793, N632);
buf BUF1 (N2269, N2264);
nor NOR3 (N2270, N2268, N240, N1548);
buf BUF1 (N2271, N2263);
buf BUF1 (N2272, N2261);
nand NAND3 (N2273, N2272, N1885, N2067);
or OR3 (N2274, N2269, N1462, N1566);
or OR4 (N2275, N2248, N1284, N598, N871);
xor XOR2 (N2276, N2257, N7);
and AND3 (N2277, N2265, N429, N2189);
or OR4 (N2278, N2274, N410, N1064, N168);
not NOT1 (N2279, N2276);
nor NOR2 (N2280, N2251, N1008);
not NOT1 (N2281, N2279);
nor NOR2 (N2282, N2266, N1402);
and AND2 (N2283, N2270, N275);
xor XOR2 (N2284, N2275, N1146);
or OR4 (N2285, N2271, N2280, N1818, N1326);
and AND3 (N2286, N121, N731, N79);
not NOT1 (N2287, N2267);
and AND3 (N2288, N2286, N1853, N1846);
buf BUF1 (N2289, N2287);
nand NAND2 (N2290, N2278, N1422);
xor XOR2 (N2291, N2284, N1176);
not NOT1 (N2292, N2277);
buf BUF1 (N2293, N2283);
and AND3 (N2294, N2273, N2163, N809);
xor XOR2 (N2295, N2293, N1898);
nor NOR2 (N2296, N2288, N1759);
not NOT1 (N2297, N2282);
xor XOR2 (N2298, N2294, N637);
nand NAND2 (N2299, N2285, N1791);
nor NOR3 (N2300, N2292, N1696, N1098);
buf BUF1 (N2301, N2299);
or OR3 (N2302, N2290, N331, N2295);
xor XOR2 (N2303, N1857, N2189);
xor XOR2 (N2304, N2301, N1241);
not NOT1 (N2305, N2297);
not NOT1 (N2306, N2302);
nand NAND2 (N2307, N2300, N530);
not NOT1 (N2308, N2303);
buf BUF1 (N2309, N2296);
not NOT1 (N2310, N2289);
and AND3 (N2311, N2309, N74, N48);
buf BUF1 (N2312, N2306);
or OR3 (N2313, N2298, N1166, N364);
nand NAND4 (N2314, N2291, N1032, N1647, N1319);
buf BUF1 (N2315, N2313);
and AND3 (N2316, N2314, N1702, N801);
and AND3 (N2317, N2315, N2122, N1634);
buf BUF1 (N2318, N2311);
buf BUF1 (N2319, N2307);
nor NOR4 (N2320, N2310, N324, N1096, N1951);
or OR3 (N2321, N2316, N1216, N980);
nor NOR2 (N2322, N2304, N71);
and AND2 (N2323, N2312, N1354);
or OR4 (N2324, N2323, N2180, N813, N1621);
buf BUF1 (N2325, N2305);
nand NAND4 (N2326, N2321, N1944, N2207, N659);
and AND3 (N2327, N2322, N2213, N572);
xor XOR2 (N2328, N2325, N93);
buf BUF1 (N2329, N2326);
xor XOR2 (N2330, N2324, N675);
nor NOR3 (N2331, N2320, N509, N1273);
not NOT1 (N2332, N2308);
and AND4 (N2333, N2332, N2250, N662, N406);
not NOT1 (N2334, N2327);
or OR2 (N2335, N2331, N694);
nor NOR4 (N2336, N2328, N810, N1214, N1096);
xor XOR2 (N2337, N2318, N257);
xor XOR2 (N2338, N2333, N97);
and AND3 (N2339, N2319, N2255, N964);
or OR4 (N2340, N2281, N81, N1784, N198);
buf BUF1 (N2341, N2317);
nor NOR3 (N2342, N2338, N1250, N448);
and AND3 (N2343, N2329, N1441, N257);
xor XOR2 (N2344, N2339, N1962);
buf BUF1 (N2345, N2344);
xor XOR2 (N2346, N2341, N247);
nand NAND4 (N2347, N2337, N1647, N426, N600);
nand NAND2 (N2348, N2345, N36);
not NOT1 (N2349, N2348);
and AND2 (N2350, N2347, N1581);
or OR2 (N2351, N2336, N239);
buf BUF1 (N2352, N2349);
xor XOR2 (N2353, N2351, N1135);
buf BUF1 (N2354, N2352);
not NOT1 (N2355, N2335);
xor XOR2 (N2356, N2340, N1027);
buf BUF1 (N2357, N2355);
xor XOR2 (N2358, N2357, N695);
buf BUF1 (N2359, N2350);
nand NAND4 (N2360, N2353, N1893, N940, N388);
not NOT1 (N2361, N2330);
not NOT1 (N2362, N2343);
not NOT1 (N2363, N2361);
nor NOR2 (N2364, N2342, N1776);
nor NOR4 (N2365, N2354, N1506, N1844, N76);
xor XOR2 (N2366, N2360, N1);
and AND4 (N2367, N2362, N1171, N1865, N2311);
xor XOR2 (N2368, N2346, N1583);
buf BUF1 (N2369, N2366);
xor XOR2 (N2370, N2369, N1294);
nand NAND4 (N2371, N2358, N202, N582, N961);
buf BUF1 (N2372, N2356);
nor NOR4 (N2373, N2359, N2354, N1686, N2102);
xor XOR2 (N2374, N2370, N1724);
nor NOR4 (N2375, N2363, N884, N266, N2346);
nor NOR2 (N2376, N2367, N949);
nor NOR2 (N2377, N2374, N1349);
and AND3 (N2378, N2334, N797, N2198);
and AND4 (N2379, N2368, N2306, N744, N316);
not NOT1 (N2380, N2373);
or OR4 (N2381, N2365, N2188, N2078, N2004);
xor XOR2 (N2382, N2380, N107);
nand NAND3 (N2383, N2372, N1905, N1498);
buf BUF1 (N2384, N2382);
and AND3 (N2385, N2383, N2211, N1362);
not NOT1 (N2386, N2381);
not NOT1 (N2387, N2386);
nor NOR3 (N2388, N2385, N1622, N1835);
nand NAND3 (N2389, N2375, N674, N1650);
nor NOR4 (N2390, N2371, N2199, N1105, N1788);
and AND3 (N2391, N2387, N1652, N2138);
buf BUF1 (N2392, N2389);
nor NOR3 (N2393, N2391, N1910, N605);
buf BUF1 (N2394, N2393);
buf BUF1 (N2395, N2388);
nand NAND4 (N2396, N2377, N2299, N2269, N1874);
not NOT1 (N2397, N2392);
nor NOR3 (N2398, N2390, N1700, N2199);
nor NOR3 (N2399, N2394, N216, N1627);
xor XOR2 (N2400, N2376, N2082);
and AND3 (N2401, N2397, N1445, N1743);
xor XOR2 (N2402, N2401, N330);
buf BUF1 (N2403, N2400);
buf BUF1 (N2404, N2396);
and AND2 (N2405, N2399, N1306);
not NOT1 (N2406, N2384);
nor NOR3 (N2407, N2378, N223, N1575);
buf BUF1 (N2408, N2398);
not NOT1 (N2409, N2395);
and AND4 (N2410, N2405, N1789, N2268, N614);
buf BUF1 (N2411, N2404);
xor XOR2 (N2412, N2403, N1245);
nor NOR2 (N2413, N2364, N427);
not NOT1 (N2414, N2379);
or OR2 (N2415, N2407, N1180);
nand NAND3 (N2416, N2402, N844, N68);
or OR3 (N2417, N2406, N2328, N1635);
buf BUF1 (N2418, N2414);
buf BUF1 (N2419, N2410);
nand NAND2 (N2420, N2419, N408);
nand NAND2 (N2421, N2409, N48);
nand NAND3 (N2422, N2417, N2319, N193);
and AND2 (N2423, N2421, N215);
not NOT1 (N2424, N2416);
nor NOR2 (N2425, N2422, N1487);
nor NOR4 (N2426, N2425, N805, N722, N851);
xor XOR2 (N2427, N2418, N727);
and AND2 (N2428, N2411, N1072);
or OR2 (N2429, N2408, N959);
xor XOR2 (N2430, N2420, N52);
xor XOR2 (N2431, N2426, N1780);
and AND2 (N2432, N2430, N668);
nor NOR3 (N2433, N2428, N1684, N1243);
buf BUF1 (N2434, N2423);
xor XOR2 (N2435, N2434, N1771);
buf BUF1 (N2436, N2415);
nand NAND2 (N2437, N2433, N1424);
and AND3 (N2438, N2436, N2065, N371);
xor XOR2 (N2439, N2437, N720);
buf BUF1 (N2440, N2439);
buf BUF1 (N2441, N2413);
and AND4 (N2442, N2412, N2395, N23, N309);
buf BUF1 (N2443, N2435);
not NOT1 (N2444, N2427);
or OR2 (N2445, N2444, N1501);
nor NOR4 (N2446, N2432, N1241, N559, N170);
nand NAND2 (N2447, N2438, N2178);
buf BUF1 (N2448, N2424);
nand NAND3 (N2449, N2431, N1427, N1062);
or OR2 (N2450, N2448, N836);
or OR4 (N2451, N2440, N319, N1437, N778);
xor XOR2 (N2452, N2441, N1952);
nand NAND4 (N2453, N2452, N1052, N1663, N1608);
buf BUF1 (N2454, N2449);
nor NOR4 (N2455, N2446, N2306, N2210, N841);
nand NAND4 (N2456, N2429, N2200, N1576, N364);
and AND2 (N2457, N2453, N689);
not NOT1 (N2458, N2442);
and AND2 (N2459, N2454, N1724);
nand NAND2 (N2460, N2458, N2049);
or OR2 (N2461, N2450, N1022);
not NOT1 (N2462, N2459);
and AND2 (N2463, N2457, N2347);
xor XOR2 (N2464, N2445, N2078);
nor NOR3 (N2465, N2443, N1029, N1825);
nand NAND3 (N2466, N2463, N1421, N698);
buf BUF1 (N2467, N2461);
nor NOR2 (N2468, N2456, N1197);
nand NAND4 (N2469, N2462, N837, N1578, N616);
not NOT1 (N2470, N2467);
nor NOR2 (N2471, N2470, N1988);
not NOT1 (N2472, N2460);
nor NOR4 (N2473, N2466, N98, N717, N1514);
xor XOR2 (N2474, N2468, N85);
or OR4 (N2475, N2469, N2043, N1764, N1999);
nand NAND4 (N2476, N2471, N719, N59, N737);
nand NAND4 (N2477, N2465, N138, N2051, N1646);
or OR2 (N2478, N2476, N25);
xor XOR2 (N2479, N2475, N2037);
or OR4 (N2480, N2478, N754, N457, N876);
buf BUF1 (N2481, N2464);
or OR2 (N2482, N2481, N1653);
or OR4 (N2483, N2479, N2017, N614, N69);
nand NAND3 (N2484, N2483, N2458, N1660);
nor NOR4 (N2485, N2482, N1102, N283, N1515);
or OR4 (N2486, N2451, N1776, N862, N103);
and AND2 (N2487, N2447, N1752);
xor XOR2 (N2488, N2474, N363);
buf BUF1 (N2489, N2487);
xor XOR2 (N2490, N2486, N196);
nand NAND3 (N2491, N2480, N1671, N2473);
not NOT1 (N2492, N2133);
buf BUF1 (N2493, N2472);
or OR4 (N2494, N2484, N1268, N1100, N2393);
not NOT1 (N2495, N2488);
buf BUF1 (N2496, N2455);
nand NAND2 (N2497, N2491, N1613);
nand NAND2 (N2498, N2477, N1467);
buf BUF1 (N2499, N2485);
buf BUF1 (N2500, N2496);
nor NOR4 (N2501, N2499, N1327, N457, N308);
buf BUF1 (N2502, N2494);
nor NOR4 (N2503, N2498, N1881, N2152, N1025);
not NOT1 (N2504, N2495);
buf BUF1 (N2505, N2503);
or OR4 (N2506, N2493, N327, N207, N1855);
and AND4 (N2507, N2502, N2077, N2175, N2396);
and AND4 (N2508, N2490, N1014, N1768, N1683);
xor XOR2 (N2509, N2489, N1995);
nor NOR4 (N2510, N2505, N1672, N853, N2300);
buf BUF1 (N2511, N2507);
nand NAND4 (N2512, N2511, N2378, N604, N2286);
nor NOR2 (N2513, N2500, N1220);
or OR3 (N2514, N2508, N1703, N1653);
xor XOR2 (N2515, N2514, N2329);
buf BUF1 (N2516, N2506);
buf BUF1 (N2517, N2509);
nor NOR2 (N2518, N2504, N1110);
and AND4 (N2519, N2515, N301, N411, N608);
nor NOR2 (N2520, N2497, N126);
and AND3 (N2521, N2513, N100, N1592);
and AND3 (N2522, N2517, N290, N1950);
or OR3 (N2523, N2516, N1583, N1627);
xor XOR2 (N2524, N2519, N565);
nand NAND4 (N2525, N2523, N2268, N2342, N1851);
xor XOR2 (N2526, N2521, N1121);
and AND2 (N2527, N2510, N1533);
nor NOR2 (N2528, N2518, N2412);
xor XOR2 (N2529, N2524, N1251);
or OR4 (N2530, N2525, N1946, N923, N662);
and AND2 (N2531, N2522, N192);
nor NOR3 (N2532, N2526, N834, N233);
nor NOR4 (N2533, N2520, N1282, N101, N1861);
and AND3 (N2534, N2492, N1230, N1592);
buf BUF1 (N2535, N2501);
buf BUF1 (N2536, N2535);
nand NAND2 (N2537, N2530, N993);
and AND2 (N2538, N2536, N941);
not NOT1 (N2539, N2528);
nand NAND4 (N2540, N2533, N2070, N1974, N299);
not NOT1 (N2541, N2512);
or OR2 (N2542, N2527, N384);
xor XOR2 (N2543, N2534, N2163);
xor XOR2 (N2544, N2532, N720);
nor NOR4 (N2545, N2544, N843, N828, N1739);
nor NOR4 (N2546, N2531, N417, N112, N1211);
or OR3 (N2547, N2542, N1037, N1947);
and AND3 (N2548, N2529, N1173, N1707);
buf BUF1 (N2549, N2546);
nor NOR4 (N2550, N2549, N1397, N1263, N1754);
nor NOR3 (N2551, N2547, N1562, N1415);
and AND4 (N2552, N2538, N328, N2240, N1490);
not NOT1 (N2553, N2541);
not NOT1 (N2554, N2545);
not NOT1 (N2555, N2550);
buf BUF1 (N2556, N2548);
or OR4 (N2557, N2552, N1862, N727, N171);
buf BUF1 (N2558, N2543);
or OR3 (N2559, N2551, N2346, N1607);
nand NAND3 (N2560, N2540, N425, N351);
xor XOR2 (N2561, N2554, N488);
buf BUF1 (N2562, N2561);
or OR3 (N2563, N2537, N6, N2411);
and AND3 (N2564, N2558, N2391, N2441);
and AND4 (N2565, N2553, N649, N1329, N409);
xor XOR2 (N2566, N2556, N2110);
nor NOR2 (N2567, N2563, N1301);
nand NAND3 (N2568, N2539, N1902, N556);
nor NOR2 (N2569, N2560, N355);
or OR2 (N2570, N2566, N2378);
or OR3 (N2571, N2557, N21, N1111);
xor XOR2 (N2572, N2565, N376);
and AND2 (N2573, N2559, N1181);
not NOT1 (N2574, N2572);
nand NAND3 (N2575, N2570, N1435, N1285);
xor XOR2 (N2576, N2564, N732);
xor XOR2 (N2577, N2573, N1780);
not NOT1 (N2578, N2571);
or OR4 (N2579, N2576, N1691, N1820, N2135);
not NOT1 (N2580, N2575);
xor XOR2 (N2581, N2568, N62);
not NOT1 (N2582, N2577);
nor NOR3 (N2583, N2555, N1548, N2143);
buf BUF1 (N2584, N2580);
or OR2 (N2585, N2582, N1583);
not NOT1 (N2586, N2574);
not NOT1 (N2587, N2585);
nor NOR4 (N2588, N2578, N1273, N957, N828);
or OR2 (N2589, N2581, N283);
not NOT1 (N2590, N2579);
nand NAND4 (N2591, N2589, N2319, N1595, N2046);
buf BUF1 (N2592, N2583);
nor NOR3 (N2593, N2592, N2191, N348);
nor NOR4 (N2594, N2567, N1925, N2404, N48);
buf BUF1 (N2595, N2562);
buf BUF1 (N2596, N2588);
xor XOR2 (N2597, N2596, N1451);
buf BUF1 (N2598, N2584);
not NOT1 (N2599, N2595);
not NOT1 (N2600, N2593);
not NOT1 (N2601, N2590);
nand NAND2 (N2602, N2598, N2299);
or OR3 (N2603, N2586, N1926, N894);
or OR3 (N2604, N2587, N1226, N83);
and AND2 (N2605, N2603, N357);
and AND3 (N2606, N2599, N34, N782);
buf BUF1 (N2607, N2605);
or OR2 (N2608, N2606, N420);
nor NOR3 (N2609, N2604, N1349, N707);
or OR2 (N2610, N2601, N2005);
nor NOR3 (N2611, N2602, N580, N2106);
buf BUF1 (N2612, N2610);
xor XOR2 (N2613, N2612, N2468);
and AND2 (N2614, N2600, N859);
buf BUF1 (N2615, N2594);
nor NOR4 (N2616, N2614, N1164, N2267, N839);
nand NAND3 (N2617, N2609, N1159, N260);
nand NAND2 (N2618, N2613, N1947);
buf BUF1 (N2619, N2611);
not NOT1 (N2620, N2615);
buf BUF1 (N2621, N2619);
xor XOR2 (N2622, N2618, N2571);
nor NOR3 (N2623, N2607, N2208, N2395);
or OR3 (N2624, N2608, N1670, N1763);
or OR2 (N2625, N2591, N138);
and AND2 (N2626, N2620, N1646);
nor NOR4 (N2627, N2626, N2153, N2399, N2321);
and AND4 (N2628, N2624, N1799, N1141, N617);
nand NAND4 (N2629, N2617, N1504, N396, N1839);
or OR3 (N2630, N2597, N659, N1264);
and AND4 (N2631, N2621, N2126, N2265, N402);
nand NAND2 (N2632, N2627, N1733);
buf BUF1 (N2633, N2629);
and AND4 (N2634, N2623, N431, N975, N119);
nand NAND4 (N2635, N2625, N104, N648, N1992);
xor XOR2 (N2636, N2569, N1783);
nand NAND4 (N2637, N2633, N290, N1862, N860);
nor NOR3 (N2638, N2631, N2147, N785);
not NOT1 (N2639, N2632);
buf BUF1 (N2640, N2637);
nor NOR2 (N2641, N2638, N669);
nand NAND3 (N2642, N2636, N1190, N682);
or OR3 (N2643, N2616, N728, N1648);
not NOT1 (N2644, N2628);
nand NAND2 (N2645, N2641, N1776);
not NOT1 (N2646, N2642);
not NOT1 (N2647, N2630);
or OR2 (N2648, N2645, N1830);
nor NOR3 (N2649, N2644, N1321, N2038);
nor NOR3 (N2650, N2640, N1527, N1897);
nor NOR4 (N2651, N2639, N966, N1430, N1427);
or OR2 (N2652, N2651, N1011);
and AND3 (N2653, N2643, N1730, N951);
xor XOR2 (N2654, N2650, N339);
buf BUF1 (N2655, N2622);
not NOT1 (N2656, N2635);
or OR4 (N2657, N2634, N1418, N2371, N24);
buf BUF1 (N2658, N2649);
or OR2 (N2659, N2653, N828);
nor NOR2 (N2660, N2648, N1658);
xor XOR2 (N2661, N2652, N1428);
and AND2 (N2662, N2655, N1340);
buf BUF1 (N2663, N2646);
or OR3 (N2664, N2661, N1100, N1930);
and AND2 (N2665, N2663, N540);
buf BUF1 (N2666, N2660);
xor XOR2 (N2667, N2658, N703);
or OR3 (N2668, N2667, N1173, N1278);
nand NAND2 (N2669, N2665, N736);
nand NAND3 (N2670, N2656, N1990, N612);
or OR4 (N2671, N2647, N2165, N1462, N20);
and AND2 (N2672, N2669, N2254);
not NOT1 (N2673, N2664);
buf BUF1 (N2674, N2671);
nor NOR4 (N2675, N2674, N1502, N382, N451);
nor NOR4 (N2676, N2670, N495, N1335, N259);
or OR2 (N2677, N2668, N1894);
nor NOR4 (N2678, N2673, N2145, N1735, N1652);
xor XOR2 (N2679, N2657, N1180);
xor XOR2 (N2680, N2678, N1113);
buf BUF1 (N2681, N2679);
or OR4 (N2682, N2654, N139, N1258, N2642);
not NOT1 (N2683, N2677);
or OR3 (N2684, N2680, N1776, N1435);
not NOT1 (N2685, N2675);
and AND2 (N2686, N2682, N1431);
buf BUF1 (N2687, N2662);
nand NAND3 (N2688, N2666, N1261, N1535);
not NOT1 (N2689, N2684);
or OR3 (N2690, N2681, N1509, N2027);
not NOT1 (N2691, N2687);
xor XOR2 (N2692, N2686, N2536);
nand NAND2 (N2693, N2688, N1967);
nand NAND4 (N2694, N2672, N2603, N2664, N2255);
buf BUF1 (N2695, N2676);
buf BUF1 (N2696, N2690);
buf BUF1 (N2697, N2694);
xor XOR2 (N2698, N2685, N494);
nor NOR4 (N2699, N2691, N2125, N1958, N492);
and AND4 (N2700, N2692, N378, N1452, N2130);
buf BUF1 (N2701, N2698);
not NOT1 (N2702, N2683);
or OR2 (N2703, N2702, N1855);
and AND4 (N2704, N2689, N259, N1451, N857);
xor XOR2 (N2705, N2659, N850);
buf BUF1 (N2706, N2703);
and AND2 (N2707, N2700, N2473);
buf BUF1 (N2708, N2704);
and AND2 (N2709, N2705, N130);
or OR2 (N2710, N2695, N1534);
or OR4 (N2711, N2693, N7, N2077, N626);
nor NOR2 (N2712, N2699, N2611);
buf BUF1 (N2713, N2710);
or OR4 (N2714, N2697, N858, N2520, N2301);
xor XOR2 (N2715, N2709, N2444);
nand NAND3 (N2716, N2711, N441, N1205);
and AND2 (N2717, N2712, N939);
nand NAND2 (N2718, N2713, N1280);
and AND3 (N2719, N2717, N1659, N358);
and AND3 (N2720, N2718, N1550, N1459);
nor NOR3 (N2721, N2701, N158, N2059);
buf BUF1 (N2722, N2720);
nor NOR2 (N2723, N2707, N620);
nor NOR2 (N2724, N2696, N2473);
and AND4 (N2725, N2724, N2081, N2542, N1980);
or OR4 (N2726, N2706, N2579, N2067, N1704);
xor XOR2 (N2727, N2719, N2351);
xor XOR2 (N2728, N2722, N716);
nand NAND2 (N2729, N2715, N475);
buf BUF1 (N2730, N2727);
xor XOR2 (N2731, N2708, N2467);
xor XOR2 (N2732, N2716, N2723);
not NOT1 (N2733, N283);
or OR2 (N2734, N2726, N174);
nand NAND3 (N2735, N2728, N185, N13);
nand NAND4 (N2736, N2733, N909, N1355, N2043);
and AND2 (N2737, N2736, N1526);
xor XOR2 (N2738, N2731, N1751);
or OR3 (N2739, N2725, N639, N1940);
and AND4 (N2740, N2730, N1223, N1165, N869);
buf BUF1 (N2741, N2714);
buf BUF1 (N2742, N2734);
or OR4 (N2743, N2729, N2316, N2584, N2236);
not NOT1 (N2744, N2738);
not NOT1 (N2745, N2740);
not NOT1 (N2746, N2737);
not NOT1 (N2747, N2745);
xor XOR2 (N2748, N2732, N1356);
buf BUF1 (N2749, N2742);
nor NOR3 (N2750, N2735, N824, N676);
and AND2 (N2751, N2743, N2068);
nor NOR4 (N2752, N2744, N2365, N2111, N174);
xor XOR2 (N2753, N2739, N315);
and AND2 (N2754, N2741, N609);
and AND4 (N2755, N2746, N1204, N756, N2721);
not NOT1 (N2756, N670);
not NOT1 (N2757, N2748);
nand NAND2 (N2758, N2752, N2505);
buf BUF1 (N2759, N2758);
not NOT1 (N2760, N2759);
buf BUF1 (N2761, N2750);
or OR3 (N2762, N2747, N192, N971);
or OR4 (N2763, N2753, N224, N771, N1092);
buf BUF1 (N2764, N2760);
or OR2 (N2765, N2764, N366);
and AND3 (N2766, N2762, N844, N628);
and AND4 (N2767, N2757, N2267, N38, N1310);
and AND2 (N2768, N2761, N1070);
or OR3 (N2769, N2749, N1484, N1214);
or OR2 (N2770, N2768, N841);
nor NOR2 (N2771, N2755, N1627);
not NOT1 (N2772, N2765);
not NOT1 (N2773, N2763);
nand NAND2 (N2774, N2756, N544);
not NOT1 (N2775, N2772);
and AND4 (N2776, N2754, N37, N1105, N968);
nand NAND4 (N2777, N2776, N2157, N107, N2693);
nor NOR2 (N2778, N2777, N1621);
buf BUF1 (N2779, N2775);
nand NAND2 (N2780, N2769, N2483);
buf BUF1 (N2781, N2774);
buf BUF1 (N2782, N2779);
or OR3 (N2783, N2770, N1745, N994);
nand NAND4 (N2784, N2766, N2489, N2268, N885);
nand NAND2 (N2785, N2784, N2219);
xor XOR2 (N2786, N2782, N1820);
buf BUF1 (N2787, N2751);
nor NOR4 (N2788, N2787, N225, N1782, N2406);
xor XOR2 (N2789, N2771, N1937);
or OR2 (N2790, N2780, N2605);
and AND4 (N2791, N2786, N330, N731, N933);
xor XOR2 (N2792, N2785, N1921);
buf BUF1 (N2793, N2792);
or OR3 (N2794, N2791, N147, N1448);
buf BUF1 (N2795, N2794);
xor XOR2 (N2796, N2788, N2214);
buf BUF1 (N2797, N2773);
xor XOR2 (N2798, N2789, N2581);
buf BUF1 (N2799, N2781);
and AND2 (N2800, N2797, N2580);
nand NAND3 (N2801, N2790, N2494, N2671);
xor XOR2 (N2802, N2793, N2126);
xor XOR2 (N2803, N2783, N992);
or OR3 (N2804, N2801, N1734, N2007);
or OR3 (N2805, N2803, N1998, N2457);
nor NOR4 (N2806, N2798, N47, N1230, N26);
nor NOR2 (N2807, N2767, N65);
xor XOR2 (N2808, N2807, N1143);
xor XOR2 (N2809, N2808, N1116);
buf BUF1 (N2810, N2795);
buf BUF1 (N2811, N2809);
xor XOR2 (N2812, N2796, N605);
xor XOR2 (N2813, N2805, N580);
nand NAND3 (N2814, N2810, N1263, N2237);
nand NAND3 (N2815, N2812, N2785, N2573);
nand NAND4 (N2816, N2811, N2198, N42, N1300);
not NOT1 (N2817, N2799);
and AND3 (N2818, N2800, N578, N2589);
not NOT1 (N2819, N2817);
and AND4 (N2820, N2818, N439, N1523, N769);
buf BUF1 (N2821, N2814);
or OR4 (N2822, N2806, N889, N1568, N2341);
or OR4 (N2823, N2778, N2438, N497, N1788);
and AND2 (N2824, N2816, N1714);
or OR4 (N2825, N2823, N2350, N2262, N1523);
nor NOR2 (N2826, N2819, N293);
not NOT1 (N2827, N2824);
buf BUF1 (N2828, N2802);
nor NOR2 (N2829, N2828, N1166);
not NOT1 (N2830, N2822);
buf BUF1 (N2831, N2804);
buf BUF1 (N2832, N2813);
and AND3 (N2833, N2815, N757, N1636);
nor NOR3 (N2834, N2827, N1779, N2182);
or OR3 (N2835, N2829, N2334, N1493);
nor NOR3 (N2836, N2830, N1685, N1099);
nor NOR2 (N2837, N2831, N516);
buf BUF1 (N2838, N2836);
and AND2 (N2839, N2825, N92);
nand NAND4 (N2840, N2833, N1050, N2026, N2307);
not NOT1 (N2841, N2821);
and AND4 (N2842, N2835, N687, N1249, N804);
and AND3 (N2843, N2826, N2562, N366);
xor XOR2 (N2844, N2839, N2627);
buf BUF1 (N2845, N2837);
not NOT1 (N2846, N2845);
nand NAND4 (N2847, N2834, N1683, N6, N1985);
nor NOR4 (N2848, N2843, N390, N1820, N2587);
buf BUF1 (N2849, N2838);
xor XOR2 (N2850, N2844, N9);
not NOT1 (N2851, N2849);
xor XOR2 (N2852, N2850, N621);
nand NAND4 (N2853, N2842, N412, N1733, N172);
or OR4 (N2854, N2847, N576, N652, N1697);
and AND3 (N2855, N2846, N2084, N2691);
nand NAND4 (N2856, N2832, N986, N1940, N2560);
nor NOR3 (N2857, N2840, N187, N1937);
buf BUF1 (N2858, N2853);
not NOT1 (N2859, N2852);
buf BUF1 (N2860, N2854);
nor NOR3 (N2861, N2859, N2498, N2665);
or OR2 (N2862, N2860, N509);
buf BUF1 (N2863, N2862);
and AND2 (N2864, N2856, N2809);
nand NAND3 (N2865, N2857, N989, N104);
not NOT1 (N2866, N2865);
nand NAND3 (N2867, N2848, N1425, N1847);
and AND2 (N2868, N2861, N2407);
xor XOR2 (N2869, N2867, N527);
nand NAND2 (N2870, N2858, N1321);
and AND4 (N2871, N2855, N1599, N1531, N2097);
not NOT1 (N2872, N2870);
buf BUF1 (N2873, N2820);
nand NAND2 (N2874, N2851, N1988);
not NOT1 (N2875, N2863);
and AND3 (N2876, N2874, N975, N259);
nor NOR2 (N2877, N2875, N1031);
nor NOR4 (N2878, N2872, N206, N1728, N1506);
not NOT1 (N2879, N2878);
xor XOR2 (N2880, N2841, N2310);
nand NAND4 (N2881, N2871, N1983, N300, N1113);
xor XOR2 (N2882, N2879, N2676);
and AND3 (N2883, N2877, N257, N1377);
nand NAND2 (N2884, N2876, N669);
nand NAND2 (N2885, N2883, N2133);
and AND2 (N2886, N2864, N1746);
and AND4 (N2887, N2868, N412, N1466, N1778);
or OR4 (N2888, N2887, N695, N1297, N1742);
xor XOR2 (N2889, N2884, N1883);
xor XOR2 (N2890, N2880, N2439);
nand NAND4 (N2891, N2866, N374, N851, N1849);
buf BUF1 (N2892, N2885);
and AND3 (N2893, N2891, N249, N2746);
or OR4 (N2894, N2889, N1800, N2278, N108);
nand NAND3 (N2895, N2869, N2096, N51);
and AND2 (N2896, N2873, N335);
and AND3 (N2897, N2895, N2100, N125);
and AND2 (N2898, N2894, N2275);
nor NOR4 (N2899, N2886, N626, N2357, N2536);
nor NOR3 (N2900, N2882, N1210, N2059);
nand NAND3 (N2901, N2899, N2715, N805);
or OR3 (N2902, N2898, N955, N1620);
nor NOR4 (N2903, N2881, N2555, N1854, N1438);
nand NAND3 (N2904, N2903, N1168, N2299);
not NOT1 (N2905, N2893);
or OR3 (N2906, N2902, N2057, N590);
nor NOR2 (N2907, N2905, N2527);
not NOT1 (N2908, N2907);
nand NAND3 (N2909, N2888, N1857, N2271);
nor NOR4 (N2910, N2890, N1015, N1104, N2716);
buf BUF1 (N2911, N2892);
buf BUF1 (N2912, N2908);
not NOT1 (N2913, N2901);
xor XOR2 (N2914, N2900, N2514);
buf BUF1 (N2915, N2904);
nand NAND4 (N2916, N2911, N155, N2905, N2226);
and AND3 (N2917, N2897, N504, N2294);
and AND4 (N2918, N2912, N2373, N2492, N1568);
nand NAND2 (N2919, N2916, N603);
and AND2 (N2920, N2909, N2327);
buf BUF1 (N2921, N2917);
buf BUF1 (N2922, N2920);
not NOT1 (N2923, N2896);
and AND2 (N2924, N2910, N1654);
and AND3 (N2925, N2919, N2897, N2307);
buf BUF1 (N2926, N2921);
nand NAND4 (N2927, N2906, N736, N498, N2141);
not NOT1 (N2928, N2925);
xor XOR2 (N2929, N2927, N961);
not NOT1 (N2930, N2922);
nand NAND2 (N2931, N2929, N2307);
buf BUF1 (N2932, N2913);
nand NAND4 (N2933, N2924, N2167, N2583, N2108);
or OR4 (N2934, N2928, N2689, N1728, N1917);
buf BUF1 (N2935, N2933);
and AND2 (N2936, N2932, N2549);
not NOT1 (N2937, N2935);
and AND2 (N2938, N2915, N398);
and AND2 (N2939, N2926, N517);
nand NAND4 (N2940, N2930, N2561, N2374, N1874);
not NOT1 (N2941, N2931);
not NOT1 (N2942, N2914);
nor NOR2 (N2943, N2936, N2183);
or OR3 (N2944, N2918, N594, N44);
or OR3 (N2945, N2934, N1437, N1467);
not NOT1 (N2946, N2942);
xor XOR2 (N2947, N2939, N513);
nand NAND3 (N2948, N2947, N399, N2875);
not NOT1 (N2949, N2944);
not NOT1 (N2950, N2941);
buf BUF1 (N2951, N2948);
nor NOR3 (N2952, N2946, N2865, N2900);
not NOT1 (N2953, N2938);
or OR3 (N2954, N2945, N179, N1447);
or OR3 (N2955, N2950, N2717, N51);
buf BUF1 (N2956, N2937);
nor NOR2 (N2957, N2955, N129);
nand NAND3 (N2958, N2952, N395, N1349);
xor XOR2 (N2959, N2954, N288);
nand NAND4 (N2960, N2956, N2748, N1548, N832);
nor NOR2 (N2961, N2943, N708);
xor XOR2 (N2962, N2960, N14);
xor XOR2 (N2963, N2957, N2195);
nor NOR4 (N2964, N2953, N788, N110, N1050);
or OR3 (N2965, N2923, N313, N2803);
or OR3 (N2966, N2963, N1472, N18);
nor NOR4 (N2967, N2958, N2180, N1929, N1160);
or OR3 (N2968, N2965, N1843, N918);
xor XOR2 (N2969, N2961, N517);
nand NAND2 (N2970, N2940, N425);
xor XOR2 (N2971, N2966, N252);
or OR4 (N2972, N2949, N1667, N1213, N2188);
nor NOR3 (N2973, N2968, N1918, N2089);
nor NOR3 (N2974, N2970, N848, N1389);
buf BUF1 (N2975, N2969);
xor XOR2 (N2976, N2951, N116);
xor XOR2 (N2977, N2962, N2347);
buf BUF1 (N2978, N2976);
xor XOR2 (N2979, N2973, N2721);
xor XOR2 (N2980, N2975, N189);
or OR4 (N2981, N2971, N32, N1234, N2377);
and AND2 (N2982, N2964, N2125);
nor NOR4 (N2983, N2981, N164, N2349, N1411);
buf BUF1 (N2984, N2979);
and AND4 (N2985, N2984, N692, N2569, N2440);
and AND3 (N2986, N2972, N1192, N2268);
not NOT1 (N2987, N2967);
xor XOR2 (N2988, N2978, N26);
nor NOR2 (N2989, N2982, N2665);
not NOT1 (N2990, N2959);
or OR4 (N2991, N2985, N2326, N2783, N848);
and AND2 (N2992, N2983, N882);
or OR4 (N2993, N2989, N2171, N2617, N458);
xor XOR2 (N2994, N2990, N583);
or OR2 (N2995, N2987, N1238);
nand NAND2 (N2996, N2980, N2943);
buf BUF1 (N2997, N2974);
nand NAND2 (N2998, N2995, N56);
not NOT1 (N2999, N2993);
and AND3 (N3000, N2977, N2029, N2464);
and AND3 (N3001, N2998, N1685, N230);
not NOT1 (N3002, N2988);
or OR4 (N3003, N3001, N2451, N4, N973);
not NOT1 (N3004, N2991);
nor NOR3 (N3005, N2992, N304, N1611);
or OR3 (N3006, N2994, N300, N579);
xor XOR2 (N3007, N2997, N801);
xor XOR2 (N3008, N3004, N859);
nor NOR3 (N3009, N3002, N2147, N2821);
xor XOR2 (N3010, N2996, N817);
xor XOR2 (N3011, N2999, N1197);
not NOT1 (N3012, N3009);
not NOT1 (N3013, N3007);
or OR4 (N3014, N3005, N2546, N2450, N1386);
xor XOR2 (N3015, N3008, N2235);
nor NOR3 (N3016, N3011, N2596, N2205);
buf BUF1 (N3017, N3006);
or OR4 (N3018, N2986, N734, N2293, N2582);
not NOT1 (N3019, N3013);
nand NAND3 (N3020, N3015, N616, N494);
nand NAND4 (N3021, N3018, N1851, N607, N1118);
nor NOR2 (N3022, N3020, N837);
nor NOR2 (N3023, N3016, N506);
buf BUF1 (N3024, N3000);
buf BUF1 (N3025, N3022);
nor NOR2 (N3026, N3010, N368);
and AND3 (N3027, N3025, N2180, N1213);
nand NAND4 (N3028, N3019, N2972, N1225, N1971);
and AND4 (N3029, N3027, N2354, N1829, N419);
buf BUF1 (N3030, N3023);
nand NAND3 (N3031, N3029, N2577, N2716);
buf BUF1 (N3032, N3014);
nand NAND2 (N3033, N3028, N2903);
not NOT1 (N3034, N3032);
not NOT1 (N3035, N3021);
or OR4 (N3036, N3012, N436, N2677, N720);
nand NAND2 (N3037, N3026, N1976);
nand NAND3 (N3038, N3017, N422, N513);
and AND3 (N3039, N3003, N94, N1122);
and AND3 (N3040, N3033, N1932, N2381);
and AND4 (N3041, N3038, N2459, N1029, N2195);
buf BUF1 (N3042, N3039);
and AND4 (N3043, N3036, N2015, N2950, N880);
and AND2 (N3044, N3043, N2218);
not NOT1 (N3045, N3031);
and AND2 (N3046, N3037, N1387);
or OR4 (N3047, N3035, N752, N1233, N860);
not NOT1 (N3048, N3041);
xor XOR2 (N3049, N3042, N1646);
and AND4 (N3050, N3034, N2443, N1764, N334);
nor NOR3 (N3051, N3030, N2297, N2363);
xor XOR2 (N3052, N3040, N1985);
and AND3 (N3053, N3046, N1771, N2122);
xor XOR2 (N3054, N3050, N607);
and AND4 (N3055, N3052, N572, N1731, N3023);
or OR4 (N3056, N3049, N2346, N2655, N1886);
nand NAND4 (N3057, N3048, N2446, N1168, N972);
and AND2 (N3058, N3057, N694);
nand NAND2 (N3059, N3053, N2033);
or OR2 (N3060, N3051, N1330);
xor XOR2 (N3061, N3044, N1069);
xor XOR2 (N3062, N3056, N1885);
buf BUF1 (N3063, N3061);
or OR4 (N3064, N3059, N536, N184, N1527);
nand NAND3 (N3065, N3045, N157, N1811);
and AND2 (N3066, N3062, N433);
and AND4 (N3067, N3024, N2344, N2113, N2500);
and AND2 (N3068, N3067, N2454);
buf BUF1 (N3069, N3054);
not NOT1 (N3070, N3064);
and AND2 (N3071, N3065, N1717);
nand NAND2 (N3072, N3069, N2608);
xor XOR2 (N3073, N3055, N1462);
nor NOR4 (N3074, N3071, N2414, N1353, N447);
buf BUF1 (N3075, N3066);
xor XOR2 (N3076, N3074, N998);
and AND2 (N3077, N3070, N19);
not NOT1 (N3078, N3058);
nor NOR4 (N3079, N3047, N294, N2723, N2352);
nand NAND3 (N3080, N3063, N1430, N183);
and AND3 (N3081, N3080, N2118, N1364);
not NOT1 (N3082, N3076);
nand NAND4 (N3083, N3081, N3057, N676, N1432);
or OR4 (N3084, N3079, N2143, N2836, N303);
or OR4 (N3085, N3083, N413, N2597, N1464);
and AND3 (N3086, N3085, N2928, N727);
xor XOR2 (N3087, N3078, N2178);
or OR2 (N3088, N3086, N797);
and AND2 (N3089, N3088, N1977);
and AND3 (N3090, N3089, N2191, N3077);
xor XOR2 (N3091, N1842, N1012);
nand NAND4 (N3092, N3068, N827, N449, N2710);
not NOT1 (N3093, N3075);
nand NAND2 (N3094, N3087, N2257);
and AND3 (N3095, N3084, N846, N2529);
xor XOR2 (N3096, N3094, N1484);
nand NAND3 (N3097, N3073, N1107, N1398);
nor NOR3 (N3098, N3095, N1492, N363);
nor NOR3 (N3099, N3090, N3058, N3073);
or OR3 (N3100, N3097, N515, N2822);
or OR2 (N3101, N3091, N1793);
buf BUF1 (N3102, N3099);
buf BUF1 (N3103, N3101);
and AND2 (N3104, N3093, N2714);
nor NOR3 (N3105, N3096, N720, N64);
nor NOR2 (N3106, N3103, N2921);
xor XOR2 (N3107, N3092, N881);
nor NOR2 (N3108, N3104, N1169);
not NOT1 (N3109, N3106);
nor NOR3 (N3110, N3108, N2956, N727);
buf BUF1 (N3111, N3105);
xor XOR2 (N3112, N3072, N2433);
nand NAND4 (N3113, N3110, N2639, N1230, N254);
or OR3 (N3114, N3082, N3102, N50);
not NOT1 (N3115, N828);
xor XOR2 (N3116, N3112, N2830);
nor NOR2 (N3117, N3100, N228);
nor NOR4 (N3118, N3115, N95, N837, N1530);
nand NAND3 (N3119, N3109, N2301, N2721);
or OR2 (N3120, N3116, N3005);
and AND4 (N3121, N3111, N916, N426, N2500);
nor NOR2 (N3122, N3098, N1884);
nand NAND4 (N3123, N3113, N1629, N788, N976);
xor XOR2 (N3124, N3117, N2149);
nand NAND4 (N3125, N3123, N2329, N741, N2992);
or OR3 (N3126, N3119, N451, N746);
nor NOR3 (N3127, N3122, N1850, N2528);
nor NOR4 (N3128, N3060, N1165, N2472, N978);
xor XOR2 (N3129, N3125, N738);
nor NOR3 (N3130, N3120, N1821, N330);
nor NOR2 (N3131, N3130, N734);
nand NAND2 (N3132, N3114, N1098);
xor XOR2 (N3133, N3131, N1129);
nand NAND3 (N3134, N3132, N2641, N250);
buf BUF1 (N3135, N3127);
nor NOR2 (N3136, N3134, N96);
xor XOR2 (N3137, N3118, N1942);
nand NAND4 (N3138, N3126, N2891, N1565, N2229);
and AND2 (N3139, N3121, N1892);
nor NOR3 (N3140, N3136, N151, N420);
not NOT1 (N3141, N3107);
buf BUF1 (N3142, N3133);
xor XOR2 (N3143, N3124, N1884);
xor XOR2 (N3144, N3141, N2434);
or OR3 (N3145, N3139, N3049, N1965);
buf BUF1 (N3146, N3140);
xor XOR2 (N3147, N3142, N2165);
nor NOR3 (N3148, N3145, N2030, N2100);
xor XOR2 (N3149, N3128, N307);
not NOT1 (N3150, N3138);
and AND4 (N3151, N3150, N563, N114, N2760);
buf BUF1 (N3152, N3144);
buf BUF1 (N3153, N3137);
nor NOR4 (N3154, N3135, N2549, N2429, N1553);
nor NOR2 (N3155, N3149, N2028);
not NOT1 (N3156, N3151);
or OR2 (N3157, N3148, N1630);
nor NOR3 (N3158, N3152, N2921, N604);
not NOT1 (N3159, N3155);
or OR4 (N3160, N3147, N1000, N735, N283);
nand NAND2 (N3161, N3143, N2793);
buf BUF1 (N3162, N3146);
and AND3 (N3163, N3160, N2660, N480);
buf BUF1 (N3164, N3158);
nand NAND2 (N3165, N3129, N324);
not NOT1 (N3166, N3165);
nand NAND2 (N3167, N3161, N647);
xor XOR2 (N3168, N3166, N1178);
not NOT1 (N3169, N3168);
buf BUF1 (N3170, N3157);
buf BUF1 (N3171, N3170);
nor NOR2 (N3172, N3164, N2196);
nor NOR2 (N3173, N3156, N2064);
or OR4 (N3174, N3162, N2273, N344, N1921);
buf BUF1 (N3175, N3171);
buf BUF1 (N3176, N3167);
and AND3 (N3177, N3169, N1959, N2586);
and AND4 (N3178, N3173, N2015, N858, N478);
and AND3 (N3179, N3175, N2714, N666);
and AND4 (N3180, N3174, N2953, N503, N954);
or OR3 (N3181, N3179, N2271, N2632);
nor NOR2 (N3182, N3178, N1454);
nand NAND4 (N3183, N3181, N1462, N1739, N2611);
nor NOR3 (N3184, N3177, N2078, N2647);
and AND3 (N3185, N3180, N2163, N494);
nor NOR3 (N3186, N3159, N1944, N1379);
and AND4 (N3187, N3153, N2830, N1825, N265);
not NOT1 (N3188, N3187);
nand NAND2 (N3189, N3182, N3135);
or OR3 (N3190, N3154, N1972, N1661);
nor NOR3 (N3191, N3185, N1151, N3176);
or OR2 (N3192, N1079, N194);
xor XOR2 (N3193, N3163, N2035);
nand NAND4 (N3194, N3184, N194, N567, N1191);
buf BUF1 (N3195, N3191);
xor XOR2 (N3196, N3183, N2696);
or OR2 (N3197, N3194, N2183);
xor XOR2 (N3198, N3188, N1221);
buf BUF1 (N3199, N3172);
nand NAND4 (N3200, N3198, N1461, N2512, N2733);
nand NAND2 (N3201, N3190, N2588);
nor NOR2 (N3202, N3196, N630);
or OR2 (N3203, N3202, N2017);
buf BUF1 (N3204, N3203);
or OR4 (N3205, N3195, N1047, N1108, N44);
nor NOR4 (N3206, N3205, N2607, N622, N2195);
xor XOR2 (N3207, N3200, N2994);
nor NOR3 (N3208, N3189, N1203, N835);
nor NOR4 (N3209, N3197, N222, N2410, N159);
not NOT1 (N3210, N3192);
not NOT1 (N3211, N3201);
and AND3 (N3212, N3209, N2957, N1385);
not NOT1 (N3213, N3212);
and AND2 (N3214, N3208, N2195);
nor NOR2 (N3215, N3204, N694);
and AND2 (N3216, N3210, N55);
xor XOR2 (N3217, N3214, N865);
buf BUF1 (N3218, N3213);
not NOT1 (N3219, N3215);
nand NAND3 (N3220, N3199, N300, N984);
not NOT1 (N3221, N3206);
and AND2 (N3222, N3218, N1573);
or OR4 (N3223, N3221, N2760, N2869, N508);
xor XOR2 (N3224, N3193, N2537);
buf BUF1 (N3225, N3211);
not NOT1 (N3226, N3220);
nand NAND4 (N3227, N3186, N1125, N2841, N352);
nor NOR3 (N3228, N3207, N2698, N3216);
not NOT1 (N3229, N1353);
nor NOR2 (N3230, N3227, N1145);
buf BUF1 (N3231, N3217);
xor XOR2 (N3232, N3224, N64);
not NOT1 (N3233, N3229);
nor NOR3 (N3234, N3223, N3042, N2883);
buf BUF1 (N3235, N3222);
xor XOR2 (N3236, N3230, N1619);
not NOT1 (N3237, N3236);
not NOT1 (N3238, N3219);
buf BUF1 (N3239, N3238);
not NOT1 (N3240, N3226);
and AND4 (N3241, N3235, N3195, N3179, N672);
and AND2 (N3242, N3233, N554);
nor NOR2 (N3243, N3232, N2079);
xor XOR2 (N3244, N3243, N496);
or OR4 (N3245, N3242, N3226, N1665, N3088);
or OR2 (N3246, N3245, N498);
nand NAND2 (N3247, N3231, N809);
nand NAND4 (N3248, N3240, N2974, N848, N1254);
buf BUF1 (N3249, N3239);
nand NAND4 (N3250, N3241, N4, N890, N2866);
and AND3 (N3251, N3249, N1822, N2971);
and AND2 (N3252, N3237, N1566);
xor XOR2 (N3253, N3244, N2235);
nand NAND3 (N3254, N3246, N582, N219);
and AND4 (N3255, N3228, N2322, N2001, N3247);
nand NAND4 (N3256, N2283, N2371, N678, N3092);
not NOT1 (N3257, N3252);
xor XOR2 (N3258, N3250, N2263);
buf BUF1 (N3259, N3254);
and AND2 (N3260, N3256, N805);
and AND3 (N3261, N3234, N822, N2119);
nand NAND2 (N3262, N3259, N2658);
nor NOR3 (N3263, N3261, N221, N275);
or OR2 (N3264, N3255, N2894);
nand NAND4 (N3265, N3251, N2302, N916, N1448);
buf BUF1 (N3266, N3262);
nand NAND3 (N3267, N3260, N2098, N2597);
nor NOR2 (N3268, N3258, N3092);
not NOT1 (N3269, N3266);
nor NOR4 (N3270, N3248, N518, N442, N166);
and AND2 (N3271, N3265, N93);
nand NAND4 (N3272, N3268, N1963, N2704, N2812);
or OR4 (N3273, N3270, N2788, N2435, N2263);
or OR3 (N3274, N3263, N917, N2911);
not NOT1 (N3275, N3225);
nor NOR3 (N3276, N3275, N1169, N1467);
nand NAND4 (N3277, N3272, N463, N336, N1268);
buf BUF1 (N3278, N3276);
xor XOR2 (N3279, N3269, N1626);
nor NOR4 (N3280, N3264, N2318, N307, N678);
not NOT1 (N3281, N3274);
nand NAND4 (N3282, N3273, N3042, N1959, N2886);
and AND4 (N3283, N3253, N1737, N1506, N2479);
buf BUF1 (N3284, N3281);
or OR2 (N3285, N3284, N2457);
or OR2 (N3286, N3283, N729);
xor XOR2 (N3287, N3278, N3076);
or OR2 (N3288, N3285, N1111);
nor NOR2 (N3289, N3282, N2667);
nor NOR2 (N3290, N3257, N1920);
xor XOR2 (N3291, N3279, N2593);
buf BUF1 (N3292, N3287);
nor NOR4 (N3293, N3292, N1143, N1524, N2122);
xor XOR2 (N3294, N3293, N2509);
or OR2 (N3295, N3289, N109);
nand NAND4 (N3296, N3286, N1791, N3085, N2556);
nand NAND2 (N3297, N3280, N153);
xor XOR2 (N3298, N3267, N1317);
and AND4 (N3299, N3277, N1372, N2013, N2096);
nand NAND3 (N3300, N3295, N183, N111);
xor XOR2 (N3301, N3296, N1124);
xor XOR2 (N3302, N3294, N707);
buf BUF1 (N3303, N3288);
not NOT1 (N3304, N3303);
not NOT1 (N3305, N3299);
not NOT1 (N3306, N3298);
nand NAND2 (N3307, N3305, N482);
nor NOR3 (N3308, N3306, N2873, N1488);
buf BUF1 (N3309, N3271);
or OR4 (N3310, N3304, N1139, N545, N1182);
not NOT1 (N3311, N3307);
nand NAND3 (N3312, N3309, N1909, N1322);
not NOT1 (N3313, N3310);
nor NOR2 (N3314, N3290, N1997);
or OR3 (N3315, N3312, N2798, N838);
buf BUF1 (N3316, N3301);
buf BUF1 (N3317, N3297);
nor NOR2 (N3318, N3317, N2858);
nand NAND2 (N3319, N3313, N1018);
nand NAND4 (N3320, N3315, N846, N1271, N275);
or OR4 (N3321, N3311, N1478, N2486, N2374);
nand NAND4 (N3322, N3314, N3254, N1515, N1950);
nand NAND2 (N3323, N3302, N1077);
nor NOR2 (N3324, N3321, N1437);
or OR4 (N3325, N3324, N1058, N1470, N2431);
xor XOR2 (N3326, N3323, N2078);
nor NOR3 (N3327, N3318, N1445, N2807);
or OR4 (N3328, N3325, N1244, N337, N2524);
buf BUF1 (N3329, N3327);
nand NAND4 (N3330, N3328, N2900, N2338, N1892);
buf BUF1 (N3331, N3330);
and AND4 (N3332, N3308, N434, N2100, N726);
not NOT1 (N3333, N3322);
nand NAND4 (N3334, N3320, N211, N171, N2153);
and AND4 (N3335, N3316, N2455, N2270, N1918);
or OR2 (N3336, N3332, N1698);
buf BUF1 (N3337, N3291);
and AND3 (N3338, N3300, N1541, N1727);
nor NOR4 (N3339, N3329, N2350, N1596, N2246);
nor NOR3 (N3340, N3337, N492, N919);
nand NAND2 (N3341, N3339, N690);
nand NAND2 (N3342, N3331, N486);
nand NAND2 (N3343, N3333, N238);
and AND4 (N3344, N3334, N520, N1459, N1110);
nor NOR4 (N3345, N3342, N1678, N44, N249);
buf BUF1 (N3346, N3344);
nor NOR4 (N3347, N3340, N2069, N406, N2751);
xor XOR2 (N3348, N3336, N2745);
buf BUF1 (N3349, N3345);
or OR2 (N3350, N3343, N926);
or OR2 (N3351, N3319, N212);
and AND2 (N3352, N3326, N2807);
nand NAND2 (N3353, N3348, N2503);
and AND2 (N3354, N3335, N2585);
nand NAND4 (N3355, N3338, N2218, N3215, N705);
xor XOR2 (N3356, N3346, N1962);
buf BUF1 (N3357, N3354);
or OR2 (N3358, N3349, N1114);
buf BUF1 (N3359, N3356);
or OR2 (N3360, N3357, N522);
nor NOR3 (N3361, N3355, N2730, N3350);
nand NAND4 (N3362, N2595, N73, N1610, N2288);
nor NOR2 (N3363, N3352, N461);
and AND3 (N3364, N3359, N2157, N1480);
nand NAND4 (N3365, N3361, N2404, N283, N3063);
not NOT1 (N3366, N3365);
xor XOR2 (N3367, N3353, N1384);
not NOT1 (N3368, N3347);
xor XOR2 (N3369, N3362, N1850);
nand NAND2 (N3370, N3351, N1229);
xor XOR2 (N3371, N3366, N2720);
xor XOR2 (N3372, N3368, N3194);
xor XOR2 (N3373, N3370, N3354);
and AND4 (N3374, N3373, N1013, N3151, N1621);
nand NAND2 (N3375, N3372, N1265);
not NOT1 (N3376, N3363);
xor XOR2 (N3377, N3341, N1018);
xor XOR2 (N3378, N3377, N3190);
not NOT1 (N3379, N3374);
nor NOR4 (N3380, N3375, N1993, N908, N2206);
xor XOR2 (N3381, N3360, N1873);
or OR2 (N3382, N3378, N1717);
xor XOR2 (N3383, N3367, N2511);
buf BUF1 (N3384, N3376);
xor XOR2 (N3385, N3369, N1356);
xor XOR2 (N3386, N3379, N2353);
nand NAND2 (N3387, N3381, N1166);
not NOT1 (N3388, N3382);
buf BUF1 (N3389, N3383);
not NOT1 (N3390, N3386);
and AND2 (N3391, N3387, N1926);
and AND4 (N3392, N3380, N2432, N2431, N262);
nand NAND3 (N3393, N3390, N637, N140);
buf BUF1 (N3394, N3392);
and AND4 (N3395, N3371, N1175, N2090, N2782);
buf BUF1 (N3396, N3385);
and AND3 (N3397, N3391, N636, N2510);
and AND2 (N3398, N3393, N1163);
or OR3 (N3399, N3358, N1487, N2361);
or OR4 (N3400, N3394, N613, N2235, N2304);
xor XOR2 (N3401, N3364, N2431);
nand NAND2 (N3402, N3400, N1633);
buf BUF1 (N3403, N3389);
nor NOR4 (N3404, N3402, N965, N3102, N2617);
buf BUF1 (N3405, N3403);
and AND3 (N3406, N3384, N2298, N624);
nand NAND4 (N3407, N3398, N2093, N3222, N1624);
not NOT1 (N3408, N3395);
and AND2 (N3409, N3401, N931);
or OR4 (N3410, N3388, N3079, N762, N85);
nor NOR4 (N3411, N3399, N3002, N932, N3019);
not NOT1 (N3412, N3405);
xor XOR2 (N3413, N3410, N2403);
xor XOR2 (N3414, N3406, N2468);
nand NAND2 (N3415, N3407, N1051);
not NOT1 (N3416, N3414);
and AND4 (N3417, N3411, N136, N3370, N142);
and AND2 (N3418, N3409, N840);
or OR2 (N3419, N3416, N3345);
xor XOR2 (N3420, N3415, N3224);
and AND4 (N3421, N3408, N1674, N2509, N151);
nand NAND4 (N3422, N3412, N2151, N1682, N120);
buf BUF1 (N3423, N3397);
not NOT1 (N3424, N3404);
or OR2 (N3425, N3396, N1791);
not NOT1 (N3426, N3421);
nand NAND2 (N3427, N3423, N1751);
nor NOR4 (N3428, N3425, N794, N659, N1343);
not NOT1 (N3429, N3427);
or OR2 (N3430, N3428, N37);
nand NAND4 (N3431, N3420, N607, N2089, N463);
xor XOR2 (N3432, N3422, N2173);
or OR2 (N3433, N3431, N2093);
or OR3 (N3434, N3432, N2360, N215);
and AND3 (N3435, N3426, N2491, N1306);
buf BUF1 (N3436, N3430);
xor XOR2 (N3437, N3418, N794);
or OR2 (N3438, N3437, N77);
buf BUF1 (N3439, N3434);
and AND4 (N3440, N3435, N3315, N1746, N1590);
or OR3 (N3441, N3429, N356, N1207);
buf BUF1 (N3442, N3440);
not NOT1 (N3443, N3433);
buf BUF1 (N3444, N3417);
xor XOR2 (N3445, N3443, N96);
nand NAND4 (N3446, N3424, N3373, N762, N215);
nand NAND2 (N3447, N3444, N2887);
buf BUF1 (N3448, N3413);
buf BUF1 (N3449, N3441);
buf BUF1 (N3450, N3442);
not NOT1 (N3451, N3436);
nor NOR3 (N3452, N3438, N915, N2671);
or OR3 (N3453, N3451, N950, N517);
not NOT1 (N3454, N3447);
nor NOR4 (N3455, N3454, N2424, N3389, N662);
not NOT1 (N3456, N3452);
not NOT1 (N3457, N3450);
nor NOR2 (N3458, N3446, N1667);
xor XOR2 (N3459, N3456, N1224);
buf BUF1 (N3460, N3459);
or OR3 (N3461, N3460, N2802, N1400);
nand NAND2 (N3462, N3457, N2839);
or OR3 (N3463, N3462, N2530, N1193);
not NOT1 (N3464, N3449);
nor NOR4 (N3465, N3419, N2620, N1790, N1609);
buf BUF1 (N3466, N3448);
and AND4 (N3467, N3453, N99, N1437, N22);
not NOT1 (N3468, N3439);
and AND2 (N3469, N3445, N2712);
buf BUF1 (N3470, N3467);
xor XOR2 (N3471, N3466, N463);
buf BUF1 (N3472, N3469);
or OR2 (N3473, N3470, N1616);
xor XOR2 (N3474, N3455, N2108);
xor XOR2 (N3475, N3471, N1992);
xor XOR2 (N3476, N3458, N2737);
nor NOR4 (N3477, N3465, N1220, N1466, N84);
and AND3 (N3478, N3475, N1129, N826);
and AND2 (N3479, N3472, N3455);
buf BUF1 (N3480, N3464);
or OR4 (N3481, N3461, N1263, N292, N3225);
nand NAND3 (N3482, N3468, N1147, N27);
not NOT1 (N3483, N3482);
xor XOR2 (N3484, N3474, N2711);
or OR4 (N3485, N3478, N451, N1311, N3204);
or OR4 (N3486, N3483, N1271, N2162, N2313);
and AND4 (N3487, N3477, N1941, N3121, N3081);
not NOT1 (N3488, N3486);
buf BUF1 (N3489, N3487);
nor NOR3 (N3490, N3479, N1477, N1702);
buf BUF1 (N3491, N3476);
not NOT1 (N3492, N3484);
buf BUF1 (N3493, N3488);
nor NOR3 (N3494, N3480, N3049, N323);
and AND2 (N3495, N3493, N3333);
nor NOR3 (N3496, N3492, N3341, N3038);
not NOT1 (N3497, N3473);
or OR3 (N3498, N3497, N817, N1652);
xor XOR2 (N3499, N3495, N2704);
nor NOR2 (N3500, N3481, N499);
nor NOR2 (N3501, N3496, N1550);
and AND2 (N3502, N3489, N1949);
xor XOR2 (N3503, N3499, N11);
nand NAND4 (N3504, N3500, N217, N175, N3053);
buf BUF1 (N3505, N3491);
xor XOR2 (N3506, N3504, N1875);
buf BUF1 (N3507, N3485);
and AND4 (N3508, N3463, N3482, N2699, N323);
and AND3 (N3509, N3506, N2276, N824);
not NOT1 (N3510, N3505);
xor XOR2 (N3511, N3508, N834);
not NOT1 (N3512, N3511);
and AND2 (N3513, N3501, N3347);
or OR2 (N3514, N3503, N2509);
nor NOR2 (N3515, N3494, N1157);
not NOT1 (N3516, N3515);
xor XOR2 (N3517, N3509, N2865);
buf BUF1 (N3518, N3514);
nor NOR3 (N3519, N3490, N235, N591);
buf BUF1 (N3520, N3513);
and AND4 (N3521, N3502, N201, N2014, N1566);
not NOT1 (N3522, N3516);
nor NOR4 (N3523, N3521, N979, N1347, N1274);
nor NOR4 (N3524, N3510, N921, N1300, N2056);
nor NOR2 (N3525, N3523, N1618);
and AND4 (N3526, N3522, N2292, N3400, N3494);
nand NAND2 (N3527, N3518, N201);
not NOT1 (N3528, N3519);
and AND3 (N3529, N3525, N2383, N2121);
or OR4 (N3530, N3524, N3225, N409, N3132);
buf BUF1 (N3531, N3526);
nor NOR4 (N3532, N3528, N1983, N2969, N1345);
not NOT1 (N3533, N3517);
buf BUF1 (N3534, N3512);
xor XOR2 (N3535, N3507, N1484);
or OR3 (N3536, N3533, N154, N2014);
not NOT1 (N3537, N3531);
buf BUF1 (N3538, N3532);
not NOT1 (N3539, N3520);
buf BUF1 (N3540, N3537);
nand NAND3 (N3541, N3539, N1925, N770);
nor NOR3 (N3542, N3498, N270, N1928);
or OR4 (N3543, N3536, N678, N2164, N2516);
and AND4 (N3544, N3535, N2103, N250, N1518);
nor NOR2 (N3545, N3542, N1553);
not NOT1 (N3546, N3534);
and AND4 (N3547, N3545, N3138, N1225, N2345);
buf BUF1 (N3548, N3541);
and AND4 (N3549, N3538, N2418, N1806, N1426);
nor NOR3 (N3550, N3543, N3358, N2489);
and AND4 (N3551, N3544, N1183, N2841, N1520);
xor XOR2 (N3552, N3547, N1515);
xor XOR2 (N3553, N3551, N2107);
nand NAND4 (N3554, N3548, N1195, N80, N3126);
nand NAND3 (N3555, N3529, N1161, N3279);
xor XOR2 (N3556, N3550, N455);
buf BUF1 (N3557, N3527);
xor XOR2 (N3558, N3549, N663);
not NOT1 (N3559, N3554);
not NOT1 (N3560, N3530);
buf BUF1 (N3561, N3552);
nor NOR2 (N3562, N3555, N3225);
nor NOR2 (N3563, N3546, N2447);
nand NAND3 (N3564, N3561, N1037, N567);
buf BUF1 (N3565, N3563);
and AND3 (N3566, N3559, N1765, N3064);
not NOT1 (N3567, N3560);
and AND2 (N3568, N3562, N3291);
nor NOR4 (N3569, N3553, N2245, N1528, N3484);
buf BUF1 (N3570, N3566);
nand NAND4 (N3571, N3556, N831, N779, N3158);
xor XOR2 (N3572, N3569, N911);
xor XOR2 (N3573, N3572, N2005);
or OR2 (N3574, N3540, N51);
buf BUF1 (N3575, N3568);
buf BUF1 (N3576, N3564);
or OR2 (N3577, N3575, N1242);
not NOT1 (N3578, N3576);
xor XOR2 (N3579, N3565, N1437);
and AND3 (N3580, N3579, N1527, N102);
buf BUF1 (N3581, N3557);
buf BUF1 (N3582, N3573);
and AND2 (N3583, N3571, N2499);
nand NAND4 (N3584, N3582, N1086, N170, N3139);
nor NOR3 (N3585, N3574, N842, N2516);
not NOT1 (N3586, N3584);
and AND3 (N3587, N3567, N2088, N2981);
not NOT1 (N3588, N3583);
nand NAND2 (N3589, N3586, N2360);
nand NAND3 (N3590, N3587, N3191, N1743);
buf BUF1 (N3591, N3585);
not NOT1 (N3592, N3588);
nor NOR3 (N3593, N3581, N504, N2531);
xor XOR2 (N3594, N3590, N3563);
buf BUF1 (N3595, N3577);
buf BUF1 (N3596, N3591);
nor NOR4 (N3597, N3589, N2799, N235, N3088);
nor NOR2 (N3598, N3578, N2411);
buf BUF1 (N3599, N3558);
or OR2 (N3600, N3580, N3066);
nand NAND2 (N3601, N3600, N3270);
nor NOR2 (N3602, N3570, N1811);
or OR4 (N3603, N3598, N56, N1112, N2566);
or OR4 (N3604, N3602, N2002, N2200, N2258);
and AND4 (N3605, N3593, N3038, N1104, N1344);
nand NAND4 (N3606, N3592, N3562, N2027, N705);
nand NAND2 (N3607, N3596, N896);
nor NOR4 (N3608, N3599, N802, N3206, N3416);
xor XOR2 (N3609, N3597, N3260);
or OR4 (N3610, N3606, N1549, N2665, N3018);
nor NOR2 (N3611, N3601, N2887);
nor NOR3 (N3612, N3604, N1703, N2222);
not NOT1 (N3613, N3605);
or OR3 (N3614, N3612, N711, N1939);
xor XOR2 (N3615, N3607, N2918);
buf BUF1 (N3616, N3608);
xor XOR2 (N3617, N3603, N3136);
and AND3 (N3618, N3611, N2869, N2596);
xor XOR2 (N3619, N3618, N985);
nand NAND2 (N3620, N3613, N1036);
buf BUF1 (N3621, N3615);
nor NOR2 (N3622, N3614, N1257);
and AND4 (N3623, N3609, N535, N3183, N747);
nand NAND2 (N3624, N3620, N1547);
xor XOR2 (N3625, N3621, N2931);
buf BUF1 (N3626, N3595);
xor XOR2 (N3627, N3623, N2060);
and AND2 (N3628, N3626, N1770);
or OR4 (N3629, N3624, N2328, N2407, N3476);
and AND4 (N3630, N3616, N1294, N3414, N456);
not NOT1 (N3631, N3594);
and AND4 (N3632, N3627, N3160, N2293, N1976);
or OR2 (N3633, N3622, N252);
not NOT1 (N3634, N3619);
and AND3 (N3635, N3625, N1962, N682);
not NOT1 (N3636, N3629);
xor XOR2 (N3637, N3610, N604);
nand NAND2 (N3638, N3630, N1737);
and AND4 (N3639, N3632, N2978, N3136, N618);
not NOT1 (N3640, N3638);
buf BUF1 (N3641, N3628);
or OR2 (N3642, N3633, N2247);
or OR3 (N3643, N3617, N2222, N142);
not NOT1 (N3644, N3637);
buf BUF1 (N3645, N3634);
not NOT1 (N3646, N3631);
and AND2 (N3647, N3640, N3198);
xor XOR2 (N3648, N3647, N1467);
nand NAND3 (N3649, N3639, N476, N2311);
or OR4 (N3650, N3642, N1101, N218, N3502);
xor XOR2 (N3651, N3649, N3509);
not NOT1 (N3652, N3644);
nor NOR2 (N3653, N3651, N2624);
nor NOR2 (N3654, N3650, N3142);
not NOT1 (N3655, N3652);
and AND3 (N3656, N3654, N2459, N2906);
nand NAND3 (N3657, N3635, N851, N3305);
or OR2 (N3658, N3641, N3358);
nand NAND3 (N3659, N3646, N508, N1021);
nor NOR4 (N3660, N3648, N1005, N1602, N1619);
buf BUF1 (N3661, N3659);
or OR4 (N3662, N3643, N1163, N636, N1021);
nor NOR2 (N3663, N3658, N2075);
or OR3 (N3664, N3653, N3515, N3456);
nand NAND3 (N3665, N3664, N3024, N2495);
buf BUF1 (N3666, N3665);
nand NAND4 (N3667, N3657, N1588, N463, N105);
nor NOR3 (N3668, N3666, N2662, N268);
xor XOR2 (N3669, N3660, N3176);
buf BUF1 (N3670, N3655);
xor XOR2 (N3671, N3662, N582);
nand NAND2 (N3672, N3671, N2219);
not NOT1 (N3673, N3667);
nand NAND3 (N3674, N3673, N8, N1610);
buf BUF1 (N3675, N3670);
buf BUF1 (N3676, N3674);
and AND2 (N3677, N3668, N1577);
buf BUF1 (N3678, N3676);
nand NAND2 (N3679, N3678, N1348);
nand NAND2 (N3680, N3663, N2024);
or OR2 (N3681, N3675, N1082);
not NOT1 (N3682, N3677);
xor XOR2 (N3683, N3681, N2264);
nand NAND4 (N3684, N3679, N2094, N1039, N1387);
buf BUF1 (N3685, N3672);
and AND2 (N3686, N3656, N762);
not NOT1 (N3687, N3686);
or OR2 (N3688, N3682, N3318);
xor XOR2 (N3689, N3687, N2332);
xor XOR2 (N3690, N3689, N688);
and AND2 (N3691, N3661, N790);
and AND2 (N3692, N3684, N2095);
buf BUF1 (N3693, N3669);
xor XOR2 (N3694, N3692, N220);
xor XOR2 (N3695, N3693, N1240);
buf BUF1 (N3696, N3680);
and AND3 (N3697, N3636, N278, N1706);
xor XOR2 (N3698, N3695, N1910);
nand NAND3 (N3699, N3690, N3377, N2763);
and AND4 (N3700, N3698, N3214, N2074, N2880);
buf BUF1 (N3701, N3685);
buf BUF1 (N3702, N3697);
buf BUF1 (N3703, N3645);
nor NOR3 (N3704, N3701, N3020, N2589);
nand NAND2 (N3705, N3691, N2239);
not NOT1 (N3706, N3700);
or OR2 (N3707, N3688, N2536);
not NOT1 (N3708, N3705);
buf BUF1 (N3709, N3696);
not NOT1 (N3710, N3704);
and AND4 (N3711, N3699, N1697, N2944, N1259);
and AND2 (N3712, N3683, N132);
nor NOR2 (N3713, N3706, N810);
and AND3 (N3714, N3703, N3396, N325);
nor NOR2 (N3715, N3711, N245);
or OR3 (N3716, N3709, N3098, N2143);
not NOT1 (N3717, N3715);
or OR3 (N3718, N3694, N966, N3489);
and AND2 (N3719, N3712, N470);
xor XOR2 (N3720, N3717, N3624);
nor NOR4 (N3721, N3720, N2702, N1324, N951);
buf BUF1 (N3722, N3713);
nand NAND3 (N3723, N3710, N2973, N3573);
not NOT1 (N3724, N3716);
not NOT1 (N3725, N3707);
or OR4 (N3726, N3714, N2490, N2956, N1461);
nand NAND4 (N3727, N3721, N3702, N2338, N1697);
not NOT1 (N3728, N2270);
xor XOR2 (N3729, N3719, N674);
xor XOR2 (N3730, N3722, N3044);
and AND3 (N3731, N3730, N45, N855);
nand NAND4 (N3732, N3728, N3393, N538, N2710);
nor NOR3 (N3733, N3723, N3099, N3168);
nor NOR4 (N3734, N3718, N1312, N247, N3559);
buf BUF1 (N3735, N3726);
or OR3 (N3736, N3734, N1574, N1911);
not NOT1 (N3737, N3736);
xor XOR2 (N3738, N3735, N3538);
buf BUF1 (N3739, N3738);
and AND3 (N3740, N3724, N2157, N3712);
xor XOR2 (N3741, N3727, N2067);
not NOT1 (N3742, N3741);
not NOT1 (N3743, N3708);
nor NOR3 (N3744, N3731, N3450, N2332);
nor NOR2 (N3745, N3742, N865);
xor XOR2 (N3746, N3740, N526);
buf BUF1 (N3747, N3746);
xor XOR2 (N3748, N3733, N1902);
not NOT1 (N3749, N3725);
nand NAND4 (N3750, N3737, N3640, N3705, N1182);
xor XOR2 (N3751, N3729, N1184);
nand NAND3 (N3752, N3749, N2096, N2181);
not NOT1 (N3753, N3732);
or OR4 (N3754, N3753, N2656, N283, N1858);
nand NAND2 (N3755, N3752, N3272);
nand NAND4 (N3756, N3739, N2805, N3026, N168);
not NOT1 (N3757, N3750);
and AND4 (N3758, N3756, N86, N12, N3278);
nor NOR4 (N3759, N3744, N3473, N25, N2040);
or OR4 (N3760, N3757, N2886, N2067, N2762);
not NOT1 (N3761, N3754);
nor NOR4 (N3762, N3758, N3097, N377, N2777);
not NOT1 (N3763, N3761);
and AND4 (N3764, N3743, N385, N773, N1711);
buf BUF1 (N3765, N3763);
or OR2 (N3766, N3751, N2529);
or OR3 (N3767, N3748, N1486, N2371);
xor XOR2 (N3768, N3766, N145);
nand NAND2 (N3769, N3759, N1522);
not NOT1 (N3770, N3768);
and AND2 (N3771, N3755, N2317);
buf BUF1 (N3772, N3764);
nand NAND2 (N3773, N3771, N3363);
or OR3 (N3774, N3767, N336, N3477);
buf BUF1 (N3775, N3769);
xor XOR2 (N3776, N3760, N660);
or OR4 (N3777, N3773, N980, N357, N1536);
buf BUF1 (N3778, N3776);
not NOT1 (N3779, N3774);
xor XOR2 (N3780, N3765, N3319);
xor XOR2 (N3781, N3778, N62);
not NOT1 (N3782, N3779);
or OR4 (N3783, N3747, N2973, N874, N1824);
and AND4 (N3784, N3780, N2182, N2015, N2995);
and AND3 (N3785, N3777, N101, N2883);
nor NOR4 (N3786, N3783, N1295, N1304, N3171);
buf BUF1 (N3787, N3772);
buf BUF1 (N3788, N3745);
buf BUF1 (N3789, N3762);
nor NOR2 (N3790, N3787, N3439);
not NOT1 (N3791, N3789);
nand NAND3 (N3792, N3791, N1439, N1253);
nor NOR4 (N3793, N3781, N2634, N1125, N45);
and AND2 (N3794, N3790, N1330);
xor XOR2 (N3795, N3786, N3525);
nand NAND4 (N3796, N3775, N2883, N541, N1345);
not NOT1 (N3797, N3788);
buf BUF1 (N3798, N3782);
nor NOR3 (N3799, N3794, N413, N767);
nand NAND2 (N3800, N3784, N721);
not NOT1 (N3801, N3785);
nand NAND2 (N3802, N3800, N3362);
and AND4 (N3803, N3770, N127, N3149, N197);
nor NOR4 (N3804, N3798, N1863, N2977, N30);
nand NAND4 (N3805, N3797, N56, N1939, N2469);
and AND2 (N3806, N3805, N383);
buf BUF1 (N3807, N3795);
xor XOR2 (N3808, N3796, N811);
not NOT1 (N3809, N3806);
or OR2 (N3810, N3804, N1914);
or OR3 (N3811, N3807, N3233, N3251);
xor XOR2 (N3812, N3792, N784);
nor NOR4 (N3813, N3799, N2404, N3043, N1858);
nand NAND4 (N3814, N3801, N2776, N2288, N3139);
xor XOR2 (N3815, N3811, N1746);
and AND3 (N3816, N3802, N3178, N3411);
nor NOR3 (N3817, N3803, N852, N153);
nand NAND2 (N3818, N3813, N305);
nor NOR2 (N3819, N3815, N1618);
nor NOR2 (N3820, N3810, N2256);
buf BUF1 (N3821, N3820);
nor NOR2 (N3822, N3808, N2915);
buf BUF1 (N3823, N3816);
buf BUF1 (N3824, N3809);
or OR4 (N3825, N3819, N2428, N1453, N794);
buf BUF1 (N3826, N3814);
or OR2 (N3827, N3821, N3294);
buf BUF1 (N3828, N3793);
and AND4 (N3829, N3822, N1025, N1002, N2323);
buf BUF1 (N3830, N3828);
buf BUF1 (N3831, N3826);
xor XOR2 (N3832, N3827, N2641);
xor XOR2 (N3833, N3823, N3392);
xor XOR2 (N3834, N3825, N1970);
or OR4 (N3835, N3833, N1478, N498, N463);
and AND3 (N3836, N3829, N3544, N1065);
not NOT1 (N3837, N3824);
xor XOR2 (N3838, N3817, N2832);
nor NOR4 (N3839, N3832, N2395, N2142, N2954);
buf BUF1 (N3840, N3812);
not NOT1 (N3841, N3835);
nand NAND4 (N3842, N3838, N3327, N1579, N3429);
nor NOR2 (N3843, N3837, N43);
and AND4 (N3844, N3830, N1975, N2906, N385);
nor NOR3 (N3845, N3844, N3749, N3214);
xor XOR2 (N3846, N3842, N889);
and AND2 (N3847, N3843, N2685);
nor NOR3 (N3848, N3846, N2608, N2725);
and AND3 (N3849, N3848, N754, N2251);
xor XOR2 (N3850, N3834, N3734);
not NOT1 (N3851, N3841);
or OR2 (N3852, N3836, N123);
not NOT1 (N3853, N3852);
xor XOR2 (N3854, N3845, N3762);
nor NOR4 (N3855, N3850, N452, N2754, N792);
and AND2 (N3856, N3840, N2893);
buf BUF1 (N3857, N3839);
buf BUF1 (N3858, N3818);
xor XOR2 (N3859, N3857, N2320);
nand NAND2 (N3860, N3849, N48);
nand NAND3 (N3861, N3853, N1066, N3675);
xor XOR2 (N3862, N3860, N843);
or OR2 (N3863, N3831, N1636);
nand NAND4 (N3864, N3855, N2164, N845, N1001);
xor XOR2 (N3865, N3861, N3148);
or OR3 (N3866, N3854, N1308, N2378);
nor NOR2 (N3867, N3858, N3580);
or OR2 (N3868, N3847, N3330);
nand NAND3 (N3869, N3868, N2817, N58);
or OR3 (N3870, N3851, N2722, N1169);
nor NOR4 (N3871, N3864, N3414, N389, N1223);
and AND3 (N3872, N3865, N2835, N3835);
not NOT1 (N3873, N3866);
nor NOR4 (N3874, N3862, N2398, N2610, N1998);
nand NAND3 (N3875, N3869, N3793, N594);
buf BUF1 (N3876, N3871);
not NOT1 (N3877, N3867);
buf BUF1 (N3878, N3863);
xor XOR2 (N3879, N3856, N3728);
buf BUF1 (N3880, N3877);
buf BUF1 (N3881, N3879);
not NOT1 (N3882, N3875);
xor XOR2 (N3883, N3874, N1560);
not NOT1 (N3884, N3882);
buf BUF1 (N3885, N3881);
not NOT1 (N3886, N3878);
or OR2 (N3887, N3880, N3753);
or OR3 (N3888, N3870, N3488, N1677);
xor XOR2 (N3889, N3859, N397);
nand NAND3 (N3890, N3876, N418, N2749);
nand NAND4 (N3891, N3887, N3642, N2032, N1702);
nand NAND3 (N3892, N3884, N2202, N801);
and AND3 (N3893, N3888, N100, N942);
nand NAND4 (N3894, N3885, N1836, N3013, N1164);
and AND4 (N3895, N3872, N374, N3323, N777);
nand NAND4 (N3896, N3895, N3881, N2133, N672);
or OR4 (N3897, N3889, N1171, N3821, N583);
or OR2 (N3898, N3894, N257);
and AND3 (N3899, N3892, N361, N3776);
nor NOR2 (N3900, N3883, N166);
buf BUF1 (N3901, N3890);
and AND2 (N3902, N3873, N344);
or OR4 (N3903, N3893, N2199, N2720, N3095);
not NOT1 (N3904, N3898);
and AND4 (N3905, N3896, N2020, N1032, N1912);
xor XOR2 (N3906, N3900, N3869);
buf BUF1 (N3907, N3899);
nor NOR2 (N3908, N3886, N2854);
nand NAND4 (N3909, N3908, N168, N845, N1446);
and AND2 (N3910, N3907, N2978);
nand NAND2 (N3911, N3904, N1458);
buf BUF1 (N3912, N3897);
not NOT1 (N3913, N3902);
xor XOR2 (N3914, N3905, N1686);
or OR3 (N3915, N3901, N2646, N1306);
or OR3 (N3916, N3910, N1488, N1232);
and AND2 (N3917, N3916, N3582);
nand NAND4 (N3918, N3891, N2558, N2343, N2354);
not NOT1 (N3919, N3913);
xor XOR2 (N3920, N3915, N1938);
buf BUF1 (N3921, N3917);
not NOT1 (N3922, N3911);
not NOT1 (N3923, N3920);
and AND2 (N3924, N3919, N2668);
or OR2 (N3925, N3924, N3295);
nand NAND3 (N3926, N3922, N2144, N2518);
or OR3 (N3927, N3903, N2877, N594);
and AND2 (N3928, N3923, N1606);
or OR3 (N3929, N3909, N2455, N2466);
nand NAND2 (N3930, N3925, N2706);
and AND2 (N3931, N3930, N3072);
xor XOR2 (N3932, N3914, N1912);
and AND4 (N3933, N3929, N3183, N1206, N829);
or OR3 (N3934, N3912, N3813, N3281);
not NOT1 (N3935, N3928);
or OR4 (N3936, N3927, N1667, N295, N2595);
and AND3 (N3937, N3934, N3568, N1180);
not NOT1 (N3938, N3906);
nand NAND3 (N3939, N3918, N906, N225);
nor NOR3 (N3940, N3933, N1672, N3345);
buf BUF1 (N3941, N3940);
nor NOR4 (N3942, N3932, N1143, N2725, N1434);
nand NAND2 (N3943, N3937, N1404);
or OR4 (N3944, N3921, N2975, N3396, N1242);
and AND4 (N3945, N3935, N203, N3914, N3502);
and AND4 (N3946, N3938, N1486, N2760, N2939);
nor NOR2 (N3947, N3926, N3114);
or OR4 (N3948, N3945, N3461, N3179, N3543);
or OR4 (N3949, N3946, N600, N359, N1790);
not NOT1 (N3950, N3948);
and AND2 (N3951, N3936, N797);
not NOT1 (N3952, N3931);
nand NAND4 (N3953, N3951, N2497, N3867, N3709);
not NOT1 (N3954, N3953);
not NOT1 (N3955, N3944);
nor NOR3 (N3956, N3955, N425, N2911);
xor XOR2 (N3957, N3943, N2891);
xor XOR2 (N3958, N3949, N886);
or OR3 (N3959, N3956, N1714, N846);
buf BUF1 (N3960, N3957);
buf BUF1 (N3961, N3939);
buf BUF1 (N3962, N3961);
and AND2 (N3963, N3960, N2487);
nor NOR2 (N3964, N3950, N3095);
or OR2 (N3965, N3959, N3114);
buf BUF1 (N3966, N3962);
and AND4 (N3967, N3947, N2463, N2711, N2275);
not NOT1 (N3968, N3964);
xor XOR2 (N3969, N3942, N3333);
nor NOR3 (N3970, N3963, N1419, N3774);
and AND4 (N3971, N3941, N1787, N2660, N1058);
nand NAND3 (N3972, N3952, N3581, N2400);
buf BUF1 (N3973, N3958);
or OR4 (N3974, N3967, N1566, N2024, N859);
nand NAND4 (N3975, N3966, N2061, N319, N985);
buf BUF1 (N3976, N3968);
or OR3 (N3977, N3970, N1870, N1113);
buf BUF1 (N3978, N3973);
nand NAND3 (N3979, N3976, N54, N2648);
and AND3 (N3980, N3969, N2637, N732);
xor XOR2 (N3981, N3974, N2647);
and AND4 (N3982, N3978, N617, N3194, N734);
xor XOR2 (N3983, N3954, N2231);
or OR4 (N3984, N3983, N2466, N3806, N852);
not NOT1 (N3985, N3979);
or OR2 (N3986, N3971, N1346);
and AND3 (N3987, N3985, N960, N866);
xor XOR2 (N3988, N3977, N839);
xor XOR2 (N3989, N3965, N1445);
xor XOR2 (N3990, N3980, N3851);
not NOT1 (N3991, N3988);
and AND4 (N3992, N3972, N3084, N2769, N389);
nand NAND2 (N3993, N3989, N2356);
buf BUF1 (N3994, N3981);
nor NOR3 (N3995, N3991, N3954, N2330);
nand NAND3 (N3996, N3990, N1131, N2043);
xor XOR2 (N3997, N3994, N135);
xor XOR2 (N3998, N3997, N2250);
not NOT1 (N3999, N3998);
and AND2 (N4000, N3987, N288);
or OR4 (N4001, N3984, N2351, N3584, N778);
nor NOR2 (N4002, N4001, N144);
xor XOR2 (N4003, N3999, N3209);
nand NAND3 (N4004, N3992, N835, N1149);
buf BUF1 (N4005, N4002);
nor NOR2 (N4006, N3995, N2143);
and AND2 (N4007, N4003, N2386);
not NOT1 (N4008, N3996);
and AND2 (N4009, N4007, N2831);
buf BUF1 (N4010, N4009);
and AND4 (N4011, N4000, N1154, N1727, N2967);
xor XOR2 (N4012, N4011, N2961);
and AND3 (N4013, N3975, N779, N268);
nor NOR2 (N4014, N4012, N3855);
nor NOR2 (N4015, N3982, N1046);
nand NAND2 (N4016, N4004, N3064);
not NOT1 (N4017, N3993);
or OR2 (N4018, N4005, N3019);
nand NAND3 (N4019, N4016, N3035, N560);
buf BUF1 (N4020, N4015);
and AND4 (N4021, N4020, N2479, N3958, N1921);
buf BUF1 (N4022, N4006);
buf BUF1 (N4023, N4008);
nor NOR3 (N4024, N3986, N3981, N4011);
nor NOR4 (N4025, N4024, N3338, N3357, N866);
nor NOR4 (N4026, N4013, N3884, N2898, N606);
not NOT1 (N4027, N4026);
or OR3 (N4028, N4018, N3595, N1527);
or OR4 (N4029, N4019, N1135, N1549, N2550);
or OR3 (N4030, N4014, N1473, N3703);
or OR3 (N4031, N4017, N1702, N493);
or OR3 (N4032, N4023, N2337, N140);
and AND3 (N4033, N4021, N46, N3086);
buf BUF1 (N4034, N4022);
nor NOR2 (N4035, N4027, N948);
xor XOR2 (N4036, N4030, N965);
or OR2 (N4037, N4032, N2617);
nand NAND3 (N4038, N4033, N1826, N732);
or OR4 (N4039, N4036, N40, N1186, N1378);
or OR4 (N4040, N4034, N3797, N1103, N2626);
nor NOR4 (N4041, N4035, N659, N594, N687);
not NOT1 (N4042, N4041);
not NOT1 (N4043, N4028);
and AND3 (N4044, N4039, N1179, N2586);
or OR4 (N4045, N4029, N3422, N1271, N2168);
or OR3 (N4046, N4038, N3904, N2839);
xor XOR2 (N4047, N4044, N2438);
not NOT1 (N4048, N4025);
not NOT1 (N4049, N4045);
nand NAND3 (N4050, N4047, N258, N2055);
nand NAND4 (N4051, N4050, N2466, N2576, N2105);
nor NOR2 (N4052, N4051, N2148);
and AND2 (N4053, N4037, N2910);
xor XOR2 (N4054, N4053, N900);
or OR2 (N4055, N4049, N3813);
not NOT1 (N4056, N4054);
buf BUF1 (N4057, N4046);
or OR4 (N4058, N4048, N2694, N1062, N928);
nand NAND4 (N4059, N4042, N183, N2118, N3382);
or OR3 (N4060, N4031, N260, N3055);
not NOT1 (N4061, N4052);
not NOT1 (N4062, N4056);
or OR3 (N4063, N4061, N746, N2942);
nor NOR2 (N4064, N4040, N2415);
nor NOR4 (N4065, N4010, N253, N3457, N2189);
not NOT1 (N4066, N4055);
xor XOR2 (N4067, N4057, N1158);
and AND2 (N4068, N4066, N3850);
buf BUF1 (N4069, N4059);
nand NAND3 (N4070, N4064, N2979, N2424);
not NOT1 (N4071, N4069);
nand NAND2 (N4072, N4067, N3408);
xor XOR2 (N4073, N4062, N3021);
nand NAND4 (N4074, N4072, N2154, N2871, N2569);
and AND3 (N4075, N4060, N203, N1307);
and AND2 (N4076, N4074, N1455);
xor XOR2 (N4077, N4070, N1904);
xor XOR2 (N4078, N4075, N3562);
nand NAND3 (N4079, N4078, N2440, N482);
nand NAND2 (N4080, N4077, N553);
nand NAND4 (N4081, N4073, N450, N4058, N1226);
buf BUF1 (N4082, N3101);
not NOT1 (N4083, N4071);
or OR2 (N4084, N4081, N1706);
nand NAND2 (N4085, N4084, N1589);
not NOT1 (N4086, N4079);
xor XOR2 (N4087, N4043, N3430);
nor NOR2 (N4088, N4080, N3585);
buf BUF1 (N4089, N4085);
or OR3 (N4090, N4086, N1948, N214);
or OR3 (N4091, N4087, N3601, N1810);
and AND2 (N4092, N4082, N1896);
and AND3 (N4093, N4091, N2700, N1338);
not NOT1 (N4094, N4076);
or OR4 (N4095, N4093, N853, N2410, N2884);
not NOT1 (N4096, N4095);
not NOT1 (N4097, N4083);
buf BUF1 (N4098, N4068);
buf BUF1 (N4099, N4094);
and AND2 (N4100, N4088, N2596);
not NOT1 (N4101, N4090);
xor XOR2 (N4102, N4097, N3226);
or OR4 (N4103, N4099, N1248, N2186, N3749);
not NOT1 (N4104, N4089);
nand NAND2 (N4105, N4104, N3218);
not NOT1 (N4106, N4105);
nor NOR4 (N4107, N4103, N2390, N1674, N3787);
or OR4 (N4108, N4065, N3425, N2214, N1780);
buf BUF1 (N4109, N4108);
buf BUF1 (N4110, N4063);
nand NAND4 (N4111, N4092, N3478, N3112, N1763);
not NOT1 (N4112, N4098);
or OR3 (N4113, N4100, N2154, N576);
xor XOR2 (N4114, N4102, N3599);
buf BUF1 (N4115, N4096);
not NOT1 (N4116, N4111);
or OR4 (N4117, N4109, N2075, N1386, N2556);
and AND3 (N4118, N4114, N581, N3558);
or OR4 (N4119, N4115, N3444, N1127, N236);
not NOT1 (N4120, N4113);
or OR3 (N4121, N4106, N1766, N3698);
xor XOR2 (N4122, N4116, N1015);
buf BUF1 (N4123, N4122);
and AND4 (N4124, N4117, N664, N3251, N2598);
buf BUF1 (N4125, N4118);
or OR4 (N4126, N4110, N296, N1756, N655);
or OR4 (N4127, N4123, N2859, N564, N840);
nor NOR3 (N4128, N4120, N1952, N667);
nor NOR3 (N4129, N4125, N3324, N544);
or OR2 (N4130, N4128, N582);
or OR4 (N4131, N4129, N110, N2930, N3443);
and AND4 (N4132, N4112, N950, N2809, N1856);
xor XOR2 (N4133, N4119, N1751);
buf BUF1 (N4134, N4124);
buf BUF1 (N4135, N4121);
and AND4 (N4136, N4133, N1620, N2532, N2002);
xor XOR2 (N4137, N4107, N3964);
not NOT1 (N4138, N4132);
buf BUF1 (N4139, N4130);
xor XOR2 (N4140, N4134, N441);
nand NAND2 (N4141, N4140, N1066);
and AND4 (N4142, N4131, N1425, N2584, N3057);
buf BUF1 (N4143, N4101);
buf BUF1 (N4144, N4136);
not NOT1 (N4145, N4127);
and AND4 (N4146, N4135, N148, N668, N3745);
nand NAND2 (N4147, N4144, N1632);
and AND4 (N4148, N4139, N308, N2147, N2674);
buf BUF1 (N4149, N4147);
and AND2 (N4150, N4149, N875);
buf BUF1 (N4151, N4145);
xor XOR2 (N4152, N4151, N3274);
not NOT1 (N4153, N4138);
xor XOR2 (N4154, N4148, N2327);
and AND2 (N4155, N4143, N156);
nor NOR4 (N4156, N4141, N736, N2494, N1799);
not NOT1 (N4157, N4152);
nand NAND4 (N4158, N4157, N178, N1390, N1977);
nor NOR3 (N4159, N4137, N2335, N3240);
or OR2 (N4160, N4126, N1110);
nand NAND2 (N4161, N4153, N3822);
buf BUF1 (N4162, N4146);
nor NOR2 (N4163, N4154, N1841);
xor XOR2 (N4164, N4161, N3056);
nor NOR4 (N4165, N4142, N3068, N2675, N3376);
nor NOR3 (N4166, N4159, N1886, N1482);
or OR2 (N4167, N4155, N4106);
buf BUF1 (N4168, N4156);
xor XOR2 (N4169, N4166, N7);
or OR2 (N4170, N4165, N288);
nand NAND4 (N4171, N4164, N2888, N2325, N3202);
nand NAND4 (N4172, N4160, N3776, N405, N131);
nand NAND3 (N4173, N4170, N2726, N1458);
buf BUF1 (N4174, N4158);
buf BUF1 (N4175, N4150);
or OR3 (N4176, N4173, N434, N2912);
nor NOR4 (N4177, N4171, N2027, N3802, N3401);
buf BUF1 (N4178, N4167);
buf BUF1 (N4179, N4168);
not NOT1 (N4180, N4162);
not NOT1 (N4181, N4176);
and AND4 (N4182, N4177, N431, N2242, N654);
buf BUF1 (N4183, N4174);
nor NOR4 (N4184, N4169, N299, N91, N3813);
xor XOR2 (N4185, N4178, N874);
and AND4 (N4186, N4185, N1105, N1067, N80);
nor NOR3 (N4187, N4184, N2173, N1720);
xor XOR2 (N4188, N4186, N1426);
nand NAND2 (N4189, N4183, N1541);
not NOT1 (N4190, N4188);
and AND4 (N4191, N4180, N295, N1299, N1704);
or OR3 (N4192, N4181, N399, N1497);
or OR3 (N4193, N4172, N1780, N1453);
and AND4 (N4194, N4187, N1342, N2679, N1959);
nand NAND2 (N4195, N4175, N1116);
buf BUF1 (N4196, N4179);
and AND3 (N4197, N4195, N2279, N3801);
xor XOR2 (N4198, N4189, N3253);
xor XOR2 (N4199, N4198, N3076);
or OR4 (N4200, N4194, N1130, N3166, N3097);
xor XOR2 (N4201, N4196, N3826);
and AND3 (N4202, N4193, N1509, N2448);
nand NAND2 (N4203, N4201, N2671);
and AND2 (N4204, N4197, N2244);
nand NAND2 (N4205, N4203, N522);
nand NAND2 (N4206, N4202, N1490);
xor XOR2 (N4207, N4192, N751);
nand NAND2 (N4208, N4204, N3334);
or OR2 (N4209, N4199, N3156);
buf BUF1 (N4210, N4163);
xor XOR2 (N4211, N4190, N2918);
and AND2 (N4212, N4209, N3033);
nand NAND2 (N4213, N4205, N351);
or OR3 (N4214, N4208, N1168, N201);
or OR2 (N4215, N4212, N1685);
not NOT1 (N4216, N4200);
and AND4 (N4217, N4216, N1660, N780, N2651);
nand NAND4 (N4218, N4211, N1556, N2884, N1960);
or OR2 (N4219, N4210, N948);
and AND3 (N4220, N4206, N2317, N1546);
and AND4 (N4221, N4218, N3387, N3033, N1451);
or OR3 (N4222, N4213, N1262, N2390);
and AND3 (N4223, N4214, N2445, N3297);
or OR3 (N4224, N4207, N29, N2022);
nand NAND2 (N4225, N4182, N404);
nand NAND4 (N4226, N4219, N208, N3075, N814);
xor XOR2 (N4227, N4222, N3509);
or OR3 (N4228, N4226, N3918, N2457);
or OR3 (N4229, N4227, N3163, N1361);
buf BUF1 (N4230, N4217);
nor NOR2 (N4231, N4228, N209);
buf BUF1 (N4232, N4231);
not NOT1 (N4233, N4223);
and AND3 (N4234, N4220, N1019, N2164);
nand NAND4 (N4235, N4225, N3476, N3409, N1493);
nor NOR3 (N4236, N4224, N3888, N635);
buf BUF1 (N4237, N4191);
xor XOR2 (N4238, N4236, N3217);
nor NOR2 (N4239, N4233, N963);
and AND2 (N4240, N4235, N2748);
nor NOR4 (N4241, N4234, N3182, N3287, N323);
xor XOR2 (N4242, N4237, N1155);
buf BUF1 (N4243, N4230);
nand NAND2 (N4244, N4229, N2143);
nor NOR2 (N4245, N4241, N487);
buf BUF1 (N4246, N4239);
nor NOR4 (N4247, N4232, N1748, N1514, N4058);
xor XOR2 (N4248, N4245, N2630);
nand NAND2 (N4249, N4248, N3140);
and AND2 (N4250, N4238, N928);
not NOT1 (N4251, N4249);
buf BUF1 (N4252, N4215);
xor XOR2 (N4253, N4246, N1377);
not NOT1 (N4254, N4240);
xor XOR2 (N4255, N4253, N3355);
not NOT1 (N4256, N4255);
nand NAND4 (N4257, N4242, N2734, N703, N2506);
and AND4 (N4258, N4256, N3849, N1782, N2632);
xor XOR2 (N4259, N4247, N2629);
xor XOR2 (N4260, N4250, N1683);
nor NOR4 (N4261, N4244, N1502, N658, N2951);
not NOT1 (N4262, N4258);
xor XOR2 (N4263, N4261, N1238);
not NOT1 (N4264, N4259);
nor NOR4 (N4265, N4221, N715, N111, N858);
nor NOR4 (N4266, N4260, N4091, N2734, N2885);
xor XOR2 (N4267, N4265, N375);
nand NAND3 (N4268, N4266, N2872, N1799);
nor NOR3 (N4269, N4251, N3104, N3406);
nand NAND2 (N4270, N4269, N3394);
not NOT1 (N4271, N4263);
not NOT1 (N4272, N4264);
xor XOR2 (N4273, N4272, N754);
not NOT1 (N4274, N4271);
or OR3 (N4275, N4243, N2950, N2758);
or OR2 (N4276, N4268, N1284);
buf BUF1 (N4277, N4257);
xor XOR2 (N4278, N4273, N4070);
nor NOR2 (N4279, N4275, N3003);
xor XOR2 (N4280, N4278, N4027);
not NOT1 (N4281, N4280);
and AND3 (N4282, N4267, N2941, N1542);
xor XOR2 (N4283, N4282, N2911);
not NOT1 (N4284, N4276);
or OR3 (N4285, N4254, N1673, N1722);
not NOT1 (N4286, N4277);
nor NOR4 (N4287, N4285, N3832, N528, N809);
buf BUF1 (N4288, N4281);
nor NOR3 (N4289, N4288, N4256, N3824);
buf BUF1 (N4290, N4286);
and AND4 (N4291, N4283, N3166, N985, N939);
nor NOR4 (N4292, N4284, N3330, N3886, N2416);
xor XOR2 (N4293, N4279, N427);
or OR2 (N4294, N4293, N3276);
and AND3 (N4295, N4274, N3077, N1111);
xor XOR2 (N4296, N4289, N63);
not NOT1 (N4297, N4296);
xor XOR2 (N4298, N4294, N1918);
and AND3 (N4299, N4252, N2931, N1167);
not NOT1 (N4300, N4299);
nor NOR2 (N4301, N4300, N3248);
buf BUF1 (N4302, N4291);
xor XOR2 (N4303, N4302, N3105);
not NOT1 (N4304, N4290);
or OR3 (N4305, N4295, N1244, N2702);
and AND3 (N4306, N4298, N1634, N2692);
xor XOR2 (N4307, N4306, N3837);
or OR3 (N4308, N4303, N1970, N1825);
or OR3 (N4309, N4270, N878, N581);
or OR4 (N4310, N4305, N2725, N575, N2904);
xor XOR2 (N4311, N4262, N1439);
not NOT1 (N4312, N4301);
buf BUF1 (N4313, N4312);
nand NAND4 (N4314, N4313, N2972, N2850, N2051);
and AND3 (N4315, N4304, N2630, N1191);
nand NAND4 (N4316, N4287, N706, N2328, N559);
and AND4 (N4317, N4311, N4301, N3969, N2256);
and AND4 (N4318, N4292, N1169, N3434, N1041);
buf BUF1 (N4319, N4318);
or OR4 (N4320, N4319, N3033, N3028, N1977);
xor XOR2 (N4321, N4309, N3652);
not NOT1 (N4322, N4317);
xor XOR2 (N4323, N4307, N3965);
nand NAND2 (N4324, N4297, N4026);
or OR4 (N4325, N4321, N3647, N1008, N3865);
not NOT1 (N4326, N4320);
nand NAND4 (N4327, N4310, N3358, N1560, N853);
xor XOR2 (N4328, N4324, N1302);
xor XOR2 (N4329, N4326, N2958);
nor NOR4 (N4330, N4316, N2915, N720, N2136);
xor XOR2 (N4331, N4325, N4256);
nand NAND2 (N4332, N4330, N1516);
buf BUF1 (N4333, N4332);
buf BUF1 (N4334, N4333);
not NOT1 (N4335, N4315);
nor NOR2 (N4336, N4334, N2158);
or OR3 (N4337, N4314, N1177, N3607);
not NOT1 (N4338, N4331);
and AND3 (N4339, N4308, N3125, N4235);
not NOT1 (N4340, N4338);
and AND2 (N4341, N4322, N2516);
nand NAND2 (N4342, N4336, N163);
nand NAND2 (N4343, N4340, N2370);
not NOT1 (N4344, N4337);
or OR2 (N4345, N4344, N2676);
not NOT1 (N4346, N4323);
and AND4 (N4347, N4342, N2378, N140, N177);
or OR3 (N4348, N4328, N2919, N3534);
buf BUF1 (N4349, N4339);
or OR4 (N4350, N4329, N3953, N2463, N3405);
and AND4 (N4351, N4350, N2167, N3915, N3328);
and AND4 (N4352, N4343, N1565, N3318, N2981);
or OR4 (N4353, N4327, N1480, N1879, N2872);
xor XOR2 (N4354, N4346, N3828);
and AND4 (N4355, N4348, N642, N1668, N975);
and AND3 (N4356, N4352, N3766, N2970);
nand NAND3 (N4357, N4347, N1340, N1706);
nor NOR4 (N4358, N4357, N3628, N527, N601);
and AND2 (N4359, N4356, N922);
buf BUF1 (N4360, N4341);
not NOT1 (N4361, N4359);
or OR4 (N4362, N4351, N112, N1936, N1010);
not NOT1 (N4363, N4360);
buf BUF1 (N4364, N4363);
buf BUF1 (N4365, N4358);
not NOT1 (N4366, N4353);
buf BUF1 (N4367, N4355);
xor XOR2 (N4368, N4365, N1152);
nor NOR3 (N4369, N4349, N1947, N1735);
nor NOR2 (N4370, N4368, N2456);
buf BUF1 (N4371, N4361);
nand NAND2 (N4372, N4370, N1041);
or OR4 (N4373, N4345, N2593, N1549, N3436);
nor NOR3 (N4374, N4371, N808, N3033);
and AND2 (N4375, N4354, N2089);
and AND4 (N4376, N4372, N1824, N3546, N4186);
xor XOR2 (N4377, N4373, N1923);
nor NOR4 (N4378, N4369, N1496, N733, N3603);
buf BUF1 (N4379, N4362);
nand NAND2 (N4380, N4367, N3020);
xor XOR2 (N4381, N4374, N1921);
nor NOR2 (N4382, N4377, N3207);
not NOT1 (N4383, N4381);
and AND3 (N4384, N4378, N676, N340);
xor XOR2 (N4385, N4375, N3491);
xor XOR2 (N4386, N4384, N4027);
xor XOR2 (N4387, N4380, N4087);
nand NAND2 (N4388, N4387, N9);
or OR3 (N4389, N4388, N2892, N2038);
nor NOR2 (N4390, N4386, N3906);
buf BUF1 (N4391, N4364);
xor XOR2 (N4392, N4385, N1023);
and AND4 (N4393, N4382, N716, N3629, N1396);
and AND3 (N4394, N4393, N1740, N4076);
and AND2 (N4395, N4394, N1410);
or OR3 (N4396, N4392, N897, N849);
and AND3 (N4397, N4335, N2680, N1521);
and AND4 (N4398, N4366, N4070, N1353, N2870);
nand NAND3 (N4399, N4376, N3402, N1095);
and AND2 (N4400, N4391, N1643);
or OR4 (N4401, N4390, N3158, N1672, N1184);
buf BUF1 (N4402, N4401);
nand NAND4 (N4403, N4396, N3483, N2944, N2295);
not NOT1 (N4404, N4398);
buf BUF1 (N4405, N4400);
buf BUF1 (N4406, N4383);
xor XOR2 (N4407, N4389, N2485);
nand NAND2 (N4408, N4402, N3434);
xor XOR2 (N4409, N4379, N578);
nor NOR4 (N4410, N4403, N3693, N665, N623);
nand NAND4 (N4411, N4397, N936, N1993, N4150);
not NOT1 (N4412, N4404);
nor NOR4 (N4413, N4410, N2835, N4029, N1394);
and AND3 (N4414, N4406, N1008, N2852);
nor NOR3 (N4415, N4407, N1489, N2428);
nand NAND4 (N4416, N4411, N1718, N295, N4370);
nand NAND4 (N4417, N4399, N3010, N2845, N2152);
or OR3 (N4418, N4415, N3676, N3976);
buf BUF1 (N4419, N4408);
and AND4 (N4420, N4413, N3221, N361, N2538);
xor XOR2 (N4421, N4417, N2422);
nor NOR3 (N4422, N4418, N1011, N980);
nor NOR3 (N4423, N4419, N1020, N3991);
buf BUF1 (N4424, N4412);
nor NOR3 (N4425, N4395, N4357, N18);
xor XOR2 (N4426, N4405, N719);
xor XOR2 (N4427, N4414, N2646);
not NOT1 (N4428, N4424);
xor XOR2 (N4429, N4409, N4171);
nand NAND4 (N4430, N4428, N837, N3021, N2949);
nand NAND3 (N4431, N4421, N4275, N1037);
or OR3 (N4432, N4420, N1953, N3576);
and AND2 (N4433, N4427, N2318);
nand NAND4 (N4434, N4433, N3286, N593, N3953);
buf BUF1 (N4435, N4430);
xor XOR2 (N4436, N4431, N3049);
xor XOR2 (N4437, N4426, N1961);
xor XOR2 (N4438, N4437, N2434);
not NOT1 (N4439, N4438);
not NOT1 (N4440, N4434);
nand NAND4 (N4441, N4432, N2790, N3477, N1876);
nor NOR4 (N4442, N4435, N3720, N1472, N944);
nand NAND4 (N4443, N4425, N4350, N1384, N1294);
buf BUF1 (N4444, N4442);
and AND2 (N4445, N4416, N4141);
and AND3 (N4446, N4444, N2904, N1148);
or OR3 (N4447, N4441, N2445, N3919);
buf BUF1 (N4448, N4446);
nand NAND4 (N4449, N4445, N982, N1545, N2467);
or OR3 (N4450, N4422, N2058, N572);
nor NOR2 (N4451, N4436, N1882);
and AND2 (N4452, N4450, N4445);
buf BUF1 (N4453, N4449);
nor NOR3 (N4454, N4443, N3918, N3012);
or OR3 (N4455, N4429, N384, N792);
nor NOR3 (N4456, N4454, N3242, N2865);
nor NOR2 (N4457, N4452, N207);
and AND3 (N4458, N4451, N4412, N3551);
not NOT1 (N4459, N4440);
and AND3 (N4460, N4423, N3562, N3238);
not NOT1 (N4461, N4455);
nor NOR4 (N4462, N4453, N757, N378, N639);
xor XOR2 (N4463, N4460, N591);
nor NOR4 (N4464, N4459, N4272, N663, N497);
buf BUF1 (N4465, N4463);
nor NOR4 (N4466, N4461, N489, N4069, N3043);
nor NOR3 (N4467, N4447, N2793, N1458);
or OR2 (N4468, N4448, N3418);
nand NAND4 (N4469, N4466, N3988, N591, N1757);
nand NAND2 (N4470, N4458, N203);
buf BUF1 (N4471, N4467);
buf BUF1 (N4472, N4465);
and AND2 (N4473, N4469, N488);
or OR2 (N4474, N4471, N2654);
or OR3 (N4475, N4456, N268, N3183);
and AND3 (N4476, N4462, N1652, N3548);
and AND2 (N4477, N4464, N63);
nand NAND3 (N4478, N4439, N2877, N3462);
buf BUF1 (N4479, N4478);
nand NAND3 (N4480, N4472, N584, N1646);
and AND2 (N4481, N4479, N1525);
and AND3 (N4482, N4470, N1964, N2048);
nand NAND2 (N4483, N4482, N38);
and AND3 (N4484, N4481, N2623, N3092);
nand NAND2 (N4485, N4484, N1747);
xor XOR2 (N4486, N4480, N2683);
and AND3 (N4487, N4486, N912, N4270);
nand NAND3 (N4488, N4487, N2074, N1634);
or OR4 (N4489, N4488, N845, N656, N2413);
nand NAND3 (N4490, N4489, N1286, N963);
and AND4 (N4491, N4485, N985, N1577, N1275);
nand NAND3 (N4492, N4476, N2932, N2815);
and AND3 (N4493, N4492, N192, N4271);
not NOT1 (N4494, N4493);
nor NOR4 (N4495, N4473, N3745, N1930, N2320);
and AND3 (N4496, N4490, N3607, N2447);
or OR4 (N4497, N4494, N3968, N1875, N849);
or OR4 (N4498, N4474, N3415, N2450, N3653);
not NOT1 (N4499, N4468);
nand NAND2 (N4500, N4496, N788);
and AND4 (N4501, N4498, N4193, N4101, N1523);
nand NAND2 (N4502, N4499, N1722);
not NOT1 (N4503, N4500);
and AND2 (N4504, N4497, N287);
nand NAND4 (N4505, N4457, N2797, N295, N3363);
or OR3 (N4506, N4483, N3029, N2296);
or OR2 (N4507, N4504, N1502);
or OR4 (N4508, N4507, N4029, N352, N1491);
nand NAND3 (N4509, N4505, N4313, N3280);
xor XOR2 (N4510, N4501, N3740);
buf BUF1 (N4511, N4495);
not NOT1 (N4512, N4477);
nand NAND4 (N4513, N4502, N2946, N3007, N3341);
and AND4 (N4514, N4506, N2248, N2930, N2162);
not NOT1 (N4515, N4508);
or OR4 (N4516, N4491, N832, N1373, N1147);
not NOT1 (N4517, N4513);
or OR2 (N4518, N4516, N3826);
and AND4 (N4519, N4503, N3550, N2978, N1590);
nand NAND2 (N4520, N4518, N528);
buf BUF1 (N4521, N4520);
nand NAND3 (N4522, N4512, N2833, N3121);
buf BUF1 (N4523, N4510);
nand NAND4 (N4524, N4519, N2422, N583, N4250);
and AND4 (N4525, N4524, N2279, N4354, N2230);
nor NOR4 (N4526, N4525, N2057, N3755, N1206);
buf BUF1 (N4527, N4526);
not NOT1 (N4528, N4521);
xor XOR2 (N4529, N4514, N3509);
not NOT1 (N4530, N4529);
xor XOR2 (N4531, N4522, N2589);
and AND3 (N4532, N4511, N2040, N3830);
nand NAND2 (N4533, N4517, N3631);
nand NAND2 (N4534, N4527, N2271);
buf BUF1 (N4535, N4534);
buf BUF1 (N4536, N4515);
nand NAND2 (N4537, N4536, N1588);
xor XOR2 (N4538, N4530, N2573);
xor XOR2 (N4539, N4532, N816);
nor NOR2 (N4540, N4475, N1005);
nand NAND2 (N4541, N4538, N4170);
xor XOR2 (N4542, N4533, N3908);
and AND3 (N4543, N4531, N1195, N558);
buf BUF1 (N4544, N4540);
nand NAND4 (N4545, N4509, N551, N2807, N4295);
nor NOR2 (N4546, N4543, N4419);
nor NOR3 (N4547, N4544, N1581, N3795);
and AND3 (N4548, N4535, N1336, N3988);
nand NAND4 (N4549, N4539, N4069, N1199, N3175);
nor NOR4 (N4550, N4541, N1953, N2564, N3896);
not NOT1 (N4551, N4546);
or OR2 (N4552, N4542, N1997);
nand NAND3 (N4553, N4551, N1797, N1671);
xor XOR2 (N4554, N4548, N3576);
and AND2 (N4555, N4537, N713);
and AND2 (N4556, N4552, N3324);
or OR4 (N4557, N4528, N2578, N1324, N342);
xor XOR2 (N4558, N4523, N1137);
and AND2 (N4559, N4558, N1180);
or OR4 (N4560, N4547, N1134, N2230, N1774);
nor NOR3 (N4561, N4559, N2354, N890);
buf BUF1 (N4562, N4555);
and AND2 (N4563, N4553, N1482);
nor NOR4 (N4564, N4556, N1582, N3010, N4403);
buf BUF1 (N4565, N4550);
buf BUF1 (N4566, N4560);
xor XOR2 (N4567, N4564, N1050);
or OR4 (N4568, N4549, N1050, N2667, N2998);
and AND2 (N4569, N4561, N2492);
xor XOR2 (N4570, N4566, N3502);
and AND2 (N4571, N4567, N4396);
nor NOR2 (N4572, N4565, N4017);
xor XOR2 (N4573, N4557, N3702);
xor XOR2 (N4574, N4545, N4418);
and AND4 (N4575, N4568, N4287, N3488, N406);
nand NAND4 (N4576, N4573, N1573, N4466, N1852);
not NOT1 (N4577, N4562);
xor XOR2 (N4578, N4576, N4133);
or OR3 (N4579, N4571, N4387, N1865);
buf BUF1 (N4580, N4572);
buf BUF1 (N4581, N4578);
not NOT1 (N4582, N4563);
buf BUF1 (N4583, N4574);
not NOT1 (N4584, N4577);
xor XOR2 (N4585, N4579, N475);
or OR3 (N4586, N4570, N2948, N1802);
xor XOR2 (N4587, N4583, N1390);
xor XOR2 (N4588, N4584, N243);
xor XOR2 (N4589, N4575, N3124);
nor NOR4 (N4590, N4585, N1387, N2062, N545);
and AND2 (N4591, N4586, N2149);
not NOT1 (N4592, N4591);
or OR3 (N4593, N4554, N3920, N2050);
not NOT1 (N4594, N4581);
or OR4 (N4595, N4588, N3062, N3017, N3131);
nand NAND4 (N4596, N4582, N266, N1675, N3086);
and AND2 (N4597, N4580, N4304);
or OR4 (N4598, N4569, N1939, N3302, N2807);
buf BUF1 (N4599, N4587);
xor XOR2 (N4600, N4598, N3368);
buf BUF1 (N4601, N4599);
nand NAND4 (N4602, N4596, N2986, N3749, N947);
and AND4 (N4603, N4594, N3483, N2078, N3045);
nand NAND3 (N4604, N4595, N3179, N577);
nor NOR3 (N4605, N4590, N1332, N1920);
and AND4 (N4606, N4601, N1841, N2416, N2741);
nand NAND3 (N4607, N4597, N808, N4455);
buf BUF1 (N4608, N4592);
and AND3 (N4609, N4589, N4154, N2462);
and AND2 (N4610, N4606, N2150);
buf BUF1 (N4611, N4593);
and AND4 (N4612, N4600, N2715, N2983, N1426);
buf BUF1 (N4613, N4602);
nand NAND2 (N4614, N4604, N2748);
nand NAND4 (N4615, N4610, N3252, N2217, N3075);
nand NAND4 (N4616, N4605, N342, N3067, N1380);
nand NAND4 (N4617, N4616, N1801, N4305, N4571);
buf BUF1 (N4618, N4612);
not NOT1 (N4619, N4607);
nand NAND4 (N4620, N4613, N3505, N3798, N1518);
buf BUF1 (N4621, N4609);
xor XOR2 (N4622, N4615, N998);
xor XOR2 (N4623, N4618, N433);
and AND4 (N4624, N4614, N3180, N380, N2034);
and AND4 (N4625, N4624, N2415, N849, N934);
xor XOR2 (N4626, N4623, N777);
xor XOR2 (N4627, N4621, N3225);
and AND4 (N4628, N4622, N1771, N977, N854);
nor NOR4 (N4629, N4603, N1337, N853, N4598);
nor NOR2 (N4630, N4620, N2824);
or OR4 (N4631, N4628, N3660, N1748, N1582);
nand NAND2 (N4632, N4625, N1452);
not NOT1 (N4633, N4617);
xor XOR2 (N4634, N4633, N2464);
nand NAND2 (N4635, N4627, N129);
or OR2 (N4636, N4619, N676);
xor XOR2 (N4637, N4630, N1186);
or OR4 (N4638, N4629, N269, N292, N4348);
or OR3 (N4639, N4632, N2069, N4611);
nand NAND2 (N4640, N2705, N4628);
not NOT1 (N4641, N4639);
nand NAND3 (N4642, N4641, N4570, N3197);
or OR2 (N4643, N4626, N2371);
nand NAND3 (N4644, N4638, N3533, N1820);
xor XOR2 (N4645, N4640, N4253);
xor XOR2 (N4646, N4642, N4541);
nor NOR2 (N4647, N4608, N2066);
and AND4 (N4648, N4637, N333, N3031, N324);
buf BUF1 (N4649, N4644);
or OR3 (N4650, N4631, N4449, N1016);
nand NAND3 (N4651, N4634, N1043, N4426);
and AND4 (N4652, N4635, N2226, N3957, N1689);
buf BUF1 (N4653, N4648);
nor NOR2 (N4654, N4643, N1346);
or OR3 (N4655, N4654, N3401, N811);
or OR2 (N4656, N4650, N3285);
not NOT1 (N4657, N4636);
or OR2 (N4658, N4655, N2559);
xor XOR2 (N4659, N4657, N2978);
nor NOR3 (N4660, N4646, N3071, N2034);
nor NOR4 (N4661, N4651, N3408, N92, N2919);
buf BUF1 (N4662, N4656);
or OR2 (N4663, N4659, N2628);
or OR2 (N4664, N4645, N3345);
nor NOR2 (N4665, N4663, N1990);
xor XOR2 (N4666, N4662, N2137);
or OR3 (N4667, N4649, N937, N1764);
buf BUF1 (N4668, N4667);
buf BUF1 (N4669, N4661);
not NOT1 (N4670, N4666);
xor XOR2 (N4671, N4665, N209);
and AND3 (N4672, N4652, N1069, N1848);
or OR2 (N4673, N4670, N1294);
nand NAND2 (N4674, N4664, N2380);
and AND2 (N4675, N4660, N3001);
nand NAND2 (N4676, N4674, N134);
and AND3 (N4677, N4647, N1825, N3517);
not NOT1 (N4678, N4668);
or OR2 (N4679, N4677, N4369);
buf BUF1 (N4680, N4679);
nor NOR4 (N4681, N4673, N12, N4190, N1565);
buf BUF1 (N4682, N4681);
and AND4 (N4683, N4682, N3551, N74, N1222);
nor NOR2 (N4684, N4658, N1372);
nor NOR2 (N4685, N4684, N4074);
nor NOR4 (N4686, N4676, N1825, N224, N1460);
nand NAND2 (N4687, N4686, N3743);
not NOT1 (N4688, N4687);
nor NOR3 (N4689, N4672, N4437, N4568);
and AND3 (N4690, N4669, N2620, N3213);
nand NAND3 (N4691, N4683, N900, N271);
nor NOR3 (N4692, N4678, N1957, N2706);
xor XOR2 (N4693, N4653, N1231);
not NOT1 (N4694, N4688);
nor NOR2 (N4695, N4693, N4061);
xor XOR2 (N4696, N4680, N3353);
not NOT1 (N4697, N4691);
and AND4 (N4698, N4697, N872, N4244, N1661);
nand NAND2 (N4699, N4675, N2704);
xor XOR2 (N4700, N4689, N3946);
buf BUF1 (N4701, N4694);
xor XOR2 (N4702, N4696, N3162);
buf BUF1 (N4703, N4685);
nand NAND3 (N4704, N4698, N255, N2171);
nand NAND4 (N4705, N4692, N1956, N2221, N692);
nand NAND4 (N4706, N4700, N2471, N4565, N2880);
buf BUF1 (N4707, N4671);
xor XOR2 (N4708, N4690, N3053);
xor XOR2 (N4709, N4695, N3867);
or OR4 (N4710, N4704, N4592, N3326, N3850);
buf BUF1 (N4711, N4701);
or OR2 (N4712, N4703, N860);
nor NOR4 (N4713, N4707, N1902, N1089, N1510);
buf BUF1 (N4714, N4708);
xor XOR2 (N4715, N4702, N10);
nand NAND2 (N4716, N4710, N427);
buf BUF1 (N4717, N4714);
buf BUF1 (N4718, N4705);
xor XOR2 (N4719, N4706, N4662);
nor NOR2 (N4720, N4719, N2752);
nor NOR4 (N4721, N4713, N1035, N4376, N599);
or OR3 (N4722, N4709, N1299, N952);
not NOT1 (N4723, N4711);
nand NAND4 (N4724, N4712, N2521, N67, N1837);
nand NAND3 (N4725, N4722, N1501, N2903);
buf BUF1 (N4726, N4720);
or OR3 (N4727, N4699, N1528, N2460);
nor NOR2 (N4728, N4724, N3106);
and AND4 (N4729, N4728, N3716, N3963, N456);
nor NOR4 (N4730, N4715, N4211, N365, N2197);
buf BUF1 (N4731, N4730);
buf BUF1 (N4732, N4727);
not NOT1 (N4733, N4717);
buf BUF1 (N4734, N4733);
nand NAND2 (N4735, N4716, N4058);
xor XOR2 (N4736, N4735, N1726);
xor XOR2 (N4737, N4736, N2000);
xor XOR2 (N4738, N4731, N4549);
buf BUF1 (N4739, N4721);
not NOT1 (N4740, N4737);
xor XOR2 (N4741, N4725, N3979);
xor XOR2 (N4742, N4718, N1843);
nand NAND3 (N4743, N4739, N1603, N4474);
and AND3 (N4744, N4726, N1015, N4633);
not NOT1 (N4745, N4729);
or OR4 (N4746, N4741, N960, N2436, N2340);
xor XOR2 (N4747, N4746, N4387);
and AND4 (N4748, N4738, N117, N1604, N1916);
nor NOR3 (N4749, N4743, N1258, N4737);
buf BUF1 (N4750, N4740);
buf BUF1 (N4751, N4749);
nor NOR2 (N4752, N4734, N2071);
nand NAND2 (N4753, N4752, N1865);
not NOT1 (N4754, N4753);
and AND2 (N4755, N4754, N2636);
xor XOR2 (N4756, N4755, N1283);
xor XOR2 (N4757, N4723, N2081);
or OR4 (N4758, N4751, N265, N377, N1351);
buf BUF1 (N4759, N4732);
xor XOR2 (N4760, N4757, N2022);
or OR4 (N4761, N4742, N3221, N2487, N1986);
buf BUF1 (N4762, N4747);
nor NOR3 (N4763, N4758, N537, N478);
nand NAND3 (N4764, N4761, N1527, N2392);
and AND3 (N4765, N4763, N3397, N3610);
xor XOR2 (N4766, N4760, N247);
not NOT1 (N4767, N4765);
or OR3 (N4768, N4767, N996, N3187);
or OR2 (N4769, N4764, N4176);
buf BUF1 (N4770, N4756);
buf BUF1 (N4771, N4762);
or OR3 (N4772, N4745, N383, N3391);
nor NOR3 (N4773, N4766, N2138, N3873);
nand NAND4 (N4774, N4750, N2517, N3947, N3704);
nand NAND3 (N4775, N4768, N1430, N2081);
not NOT1 (N4776, N4748);
xor XOR2 (N4777, N4769, N4218);
nor NOR4 (N4778, N4772, N447, N1591, N1433);
nor NOR2 (N4779, N4744, N3833);
or OR4 (N4780, N4774, N729, N3058, N1683);
and AND2 (N4781, N4780, N1565);
and AND3 (N4782, N4773, N3721, N2515);
nor NOR3 (N4783, N4771, N3193, N3426);
nand NAND3 (N4784, N4778, N3137, N4147);
and AND3 (N4785, N4782, N4264, N4094);
not NOT1 (N4786, N4776);
xor XOR2 (N4787, N4784, N2997);
nor NOR2 (N4788, N4781, N2927);
not NOT1 (N4789, N4770);
xor XOR2 (N4790, N4777, N443);
not NOT1 (N4791, N4783);
nand NAND2 (N4792, N4785, N109);
not NOT1 (N4793, N4787);
xor XOR2 (N4794, N4793, N2923);
nand NAND4 (N4795, N4759, N4098, N4057, N1360);
xor XOR2 (N4796, N4788, N3287);
buf BUF1 (N4797, N4775);
nor NOR4 (N4798, N4794, N4113, N384, N1548);
not NOT1 (N4799, N4796);
not NOT1 (N4800, N4795);
or OR2 (N4801, N4792, N726);
buf BUF1 (N4802, N4799);
not NOT1 (N4803, N4779);
not NOT1 (N4804, N4791);
or OR2 (N4805, N4798, N116);
buf BUF1 (N4806, N4797);
not NOT1 (N4807, N4800);
or OR2 (N4808, N4802, N1827);
buf BUF1 (N4809, N4805);
xor XOR2 (N4810, N4808, N2727);
nand NAND3 (N4811, N4801, N1566, N1536);
and AND2 (N4812, N4809, N2333);
and AND2 (N4813, N4806, N4587);
buf BUF1 (N4814, N4803);
nand NAND3 (N4815, N4804, N3747, N2878);
nand NAND3 (N4816, N4790, N801, N4375);
not NOT1 (N4817, N4811);
buf BUF1 (N4818, N4817);
or OR3 (N4819, N4813, N446, N798);
not NOT1 (N4820, N4789);
buf BUF1 (N4821, N4819);
buf BUF1 (N4822, N4812);
xor XOR2 (N4823, N4807, N2796);
nor NOR4 (N4824, N4786, N2658, N733, N514);
nor NOR2 (N4825, N4816, N2371);
xor XOR2 (N4826, N4824, N3404);
nor NOR3 (N4827, N4822, N809, N138);
xor XOR2 (N4828, N4821, N1171);
xor XOR2 (N4829, N4823, N3552);
nand NAND4 (N4830, N4818, N1648, N2489, N741);
xor XOR2 (N4831, N4826, N859);
nor NOR3 (N4832, N4831, N255, N1282);
or OR4 (N4833, N4828, N1653, N522, N2646);
not NOT1 (N4834, N4827);
nand NAND4 (N4835, N4815, N2985, N4267, N269);
nor NOR2 (N4836, N4820, N2313);
or OR3 (N4837, N4825, N160, N3530);
nand NAND3 (N4838, N4833, N4698, N2125);
and AND2 (N4839, N4836, N4211);
not NOT1 (N4840, N4829);
nor NOR2 (N4841, N4838, N4468);
not NOT1 (N4842, N4840);
xor XOR2 (N4843, N4814, N4417);
not NOT1 (N4844, N4832);
or OR2 (N4845, N4810, N2709);
buf BUF1 (N4846, N4842);
not NOT1 (N4847, N4846);
nor NOR3 (N4848, N4830, N492, N3964);
xor XOR2 (N4849, N4847, N1966);
buf BUF1 (N4850, N4835);
or OR4 (N4851, N4848, N4446, N4644, N745);
not NOT1 (N4852, N4843);
buf BUF1 (N4853, N4849);
nand NAND2 (N4854, N4851, N1493);
and AND4 (N4855, N4845, N4464, N2975, N3793);
nor NOR3 (N4856, N4841, N3204, N2955);
nor NOR3 (N4857, N4852, N3706, N369);
not NOT1 (N4858, N4853);
not NOT1 (N4859, N4850);
and AND4 (N4860, N4854, N364, N888, N4332);
not NOT1 (N4861, N4857);
nor NOR3 (N4862, N4861, N2871, N1381);
nand NAND3 (N4863, N4862, N121, N1264);
or OR3 (N4864, N4844, N2500, N1771);
buf BUF1 (N4865, N4834);
buf BUF1 (N4866, N4839);
and AND4 (N4867, N4856, N3606, N1978, N2917);
or OR4 (N4868, N4860, N815, N4268, N1326);
nor NOR4 (N4869, N4866, N382, N1880, N534);
not NOT1 (N4870, N4865);
or OR2 (N4871, N4869, N2031);
not NOT1 (N4872, N4859);
xor XOR2 (N4873, N4870, N3484);
not NOT1 (N4874, N4868);
or OR2 (N4875, N4855, N1610);
not NOT1 (N4876, N4863);
xor XOR2 (N4877, N4864, N2334);
or OR4 (N4878, N4874, N1318, N4757, N2606);
nand NAND2 (N4879, N4878, N4495);
nand NAND4 (N4880, N4879, N1368, N1941, N4582);
nor NOR3 (N4881, N4872, N939, N4482);
xor XOR2 (N4882, N4873, N1701);
nor NOR3 (N4883, N4882, N2354, N2604);
or OR4 (N4884, N4837, N4393, N2775, N3537);
or OR4 (N4885, N4876, N3955, N3002, N2321);
nand NAND4 (N4886, N4877, N2551, N42, N290);
and AND3 (N4887, N4885, N4761, N299);
buf BUF1 (N4888, N4881);
nor NOR3 (N4889, N4858, N3351, N4389);
nor NOR2 (N4890, N4867, N1824);
or OR2 (N4891, N4883, N2296);
xor XOR2 (N4892, N4875, N414);
xor XOR2 (N4893, N4892, N4190);
xor XOR2 (N4894, N4880, N4304);
buf BUF1 (N4895, N4890);
or OR3 (N4896, N4871, N1842, N2029);
nand NAND4 (N4897, N4891, N3294, N1483, N3330);
nor NOR4 (N4898, N4887, N568, N4172, N58);
nand NAND4 (N4899, N4897, N2286, N3835, N2606);
and AND3 (N4900, N4886, N2613, N4248);
or OR2 (N4901, N4895, N3450);
nor NOR2 (N4902, N4899, N446);
nand NAND2 (N4903, N4889, N3417);
buf BUF1 (N4904, N4888);
nor NOR2 (N4905, N4902, N4448);
nor NOR4 (N4906, N4884, N692, N3346, N3417);
buf BUF1 (N4907, N4893);
or OR2 (N4908, N4907, N2266);
nand NAND2 (N4909, N4894, N1652);
or OR2 (N4910, N4901, N1399);
nor NOR2 (N4911, N4900, N2129);
xor XOR2 (N4912, N4909, N618);
not NOT1 (N4913, N4910);
buf BUF1 (N4914, N4912);
not NOT1 (N4915, N4913);
xor XOR2 (N4916, N4898, N2150);
buf BUF1 (N4917, N4905);
buf BUF1 (N4918, N4911);
or OR3 (N4919, N4915, N1495, N1357);
and AND2 (N4920, N4904, N1737);
or OR3 (N4921, N4903, N3480, N2170);
xor XOR2 (N4922, N4917, N3247);
not NOT1 (N4923, N4908);
or OR3 (N4924, N4914, N297, N3475);
nor NOR2 (N4925, N4923, N2462);
not NOT1 (N4926, N4919);
nor NOR2 (N4927, N4926, N1211);
nand NAND2 (N4928, N4916, N4071);
not NOT1 (N4929, N4925);
buf BUF1 (N4930, N4928);
not NOT1 (N4931, N4930);
not NOT1 (N4932, N4929);
buf BUF1 (N4933, N4921);
and AND2 (N4934, N4906, N216);
and AND3 (N4935, N4933, N4431, N2184);
nand NAND2 (N4936, N4935, N70);
not NOT1 (N4937, N4927);
buf BUF1 (N4938, N4922);
not NOT1 (N4939, N4896);
not NOT1 (N4940, N4920);
nor NOR2 (N4941, N4939, N56);
nor NOR2 (N4942, N4931, N803);
and AND2 (N4943, N4940, N2265);
nor NOR3 (N4944, N4918, N1584, N743);
nor NOR3 (N4945, N4937, N3964, N1974);
buf BUF1 (N4946, N4936);
or OR2 (N4947, N4924, N4524);
xor XOR2 (N4948, N4943, N4324);
nand NAND4 (N4949, N4948, N4493, N3586, N3187);
buf BUF1 (N4950, N4932);
nor NOR3 (N4951, N4945, N4137, N4013);
not NOT1 (N4952, N4946);
nor NOR2 (N4953, N4952, N4928);
not NOT1 (N4954, N4938);
nor NOR2 (N4955, N4944, N1665);
nand NAND2 (N4956, N4953, N3275);
and AND2 (N4957, N4950, N3293);
and AND3 (N4958, N4942, N1889, N1833);
not NOT1 (N4959, N4949);
nand NAND4 (N4960, N4958, N522, N4302, N3866);
xor XOR2 (N4961, N4955, N683);
nand NAND4 (N4962, N4957, N4627, N7, N2164);
xor XOR2 (N4963, N4962, N47);
or OR2 (N4964, N4960, N1252);
not NOT1 (N4965, N4954);
nand NAND2 (N4966, N4956, N4660);
or OR4 (N4967, N4959, N4860, N40, N3285);
or OR2 (N4968, N4963, N1569);
buf BUF1 (N4969, N4941);
nand NAND2 (N4970, N4965, N2021);
and AND2 (N4971, N4961, N4170);
xor XOR2 (N4972, N4970, N806);
or OR2 (N4973, N4966, N2604);
not NOT1 (N4974, N4972);
not NOT1 (N4975, N4968);
nand NAND4 (N4976, N4973, N3993, N2124, N4162);
or OR4 (N4977, N4975, N4028, N249, N970);
nor NOR2 (N4978, N4951, N2881);
not NOT1 (N4979, N4964);
nor NOR2 (N4980, N4976, N1257);
nand NAND4 (N4981, N4967, N1148, N3792, N3390);
buf BUF1 (N4982, N4947);
not NOT1 (N4983, N4978);
not NOT1 (N4984, N4974);
buf BUF1 (N4985, N4934);
nor NOR4 (N4986, N4984, N1293, N3979, N463);
buf BUF1 (N4987, N4985);
nor NOR4 (N4988, N4983, N4111, N2931, N344);
xor XOR2 (N4989, N4980, N1240);
not NOT1 (N4990, N4982);
xor XOR2 (N4991, N4969, N4319);
buf BUF1 (N4992, N4977);
not NOT1 (N4993, N4989);
or OR3 (N4994, N4979, N493, N3877);
nand NAND4 (N4995, N4993, N3536, N4858, N1993);
not NOT1 (N4996, N4994);
or OR3 (N4997, N4981, N4912, N1575);
nand NAND2 (N4998, N4986, N435);
nor NOR4 (N4999, N4997, N685, N4988, N3900);
nand NAND2 (N5000, N3612, N3684);
xor XOR2 (N5001, N4998, N342);
not NOT1 (N5002, N4996);
nor NOR3 (N5003, N4990, N3681, N2351);
buf BUF1 (N5004, N5001);
nand NAND2 (N5005, N4971, N3581);
not NOT1 (N5006, N5005);
or OR2 (N5007, N4999, N1640);
xor XOR2 (N5008, N4987, N4872);
buf BUF1 (N5009, N5006);
xor XOR2 (N5010, N4991, N3385);
not NOT1 (N5011, N5007);
nor NOR3 (N5012, N5004, N4198, N2355);
xor XOR2 (N5013, N5012, N4793);
buf BUF1 (N5014, N5013);
not NOT1 (N5015, N5009);
nand NAND3 (N5016, N4995, N576, N323);
buf BUF1 (N5017, N5014);
and AND2 (N5018, N5016, N4883);
xor XOR2 (N5019, N5008, N3028);
not NOT1 (N5020, N5017);
not NOT1 (N5021, N5020);
buf BUF1 (N5022, N5000);
buf BUF1 (N5023, N5003);
not NOT1 (N5024, N5015);
buf BUF1 (N5025, N5023);
nand NAND3 (N5026, N5022, N848, N1656);
xor XOR2 (N5027, N5021, N1680);
or OR3 (N5028, N5024, N1677, N1781);
or OR2 (N5029, N5011, N1889);
xor XOR2 (N5030, N5010, N1006);
nor NOR4 (N5031, N5018, N4430, N1561, N3679);
nor NOR2 (N5032, N5030, N4203);
nor NOR3 (N5033, N5027, N325, N4989);
buf BUF1 (N5034, N5029);
or OR3 (N5035, N5026, N4784, N1120);
or OR2 (N5036, N5019, N13);
or OR4 (N5037, N5025, N87, N4518, N430);
not NOT1 (N5038, N5035);
nor NOR3 (N5039, N5034, N2283, N1908);
not NOT1 (N5040, N5031);
xor XOR2 (N5041, N5039, N2404);
or OR3 (N5042, N5041, N1321, N657);
nor NOR2 (N5043, N5042, N2341);
nand NAND3 (N5044, N5038, N4184, N3025);
xor XOR2 (N5045, N5040, N3240);
nand NAND4 (N5046, N5028, N1645, N1005, N3104);
nand NAND2 (N5047, N5002, N4258);
xor XOR2 (N5048, N5047, N1238);
xor XOR2 (N5049, N5043, N1255);
and AND3 (N5050, N5044, N3282, N1470);
and AND4 (N5051, N5037, N1907, N695, N154);
nor NOR3 (N5052, N5046, N2995, N3234);
or OR2 (N5053, N4992, N1114);
nor NOR2 (N5054, N5033, N3338);
and AND2 (N5055, N5048, N4373);
or OR3 (N5056, N5053, N3416, N924);
or OR2 (N5057, N5055, N1555);
and AND4 (N5058, N5050, N733, N4166, N4397);
nand NAND3 (N5059, N5056, N4708, N3476);
buf BUF1 (N5060, N5052);
not NOT1 (N5061, N5045);
buf BUF1 (N5062, N5059);
nor NOR3 (N5063, N5051, N2723, N4047);
not NOT1 (N5064, N5032);
xor XOR2 (N5065, N5064, N1917);
and AND3 (N5066, N5063, N2579, N3383);
or OR4 (N5067, N5049, N1727, N3887, N3365);
buf BUF1 (N5068, N5062);
not NOT1 (N5069, N5060);
nand NAND3 (N5070, N5058, N3736, N2826);
xor XOR2 (N5071, N5068, N5054);
or OR4 (N5072, N2047, N4160, N846, N4484);
xor XOR2 (N5073, N5066, N2183);
nor NOR2 (N5074, N5071, N1541);
or OR4 (N5075, N5070, N433, N497, N49);
or OR2 (N5076, N5074, N746);
nor NOR3 (N5077, N5073, N1767, N2424);
not NOT1 (N5078, N5075);
xor XOR2 (N5079, N5067, N4518);
and AND2 (N5080, N5061, N4828);
not NOT1 (N5081, N5079);
and AND4 (N5082, N5072, N1779, N2289, N4530);
and AND3 (N5083, N5069, N4888, N953);
not NOT1 (N5084, N5065);
not NOT1 (N5085, N5084);
and AND2 (N5086, N5082, N2086);
or OR2 (N5087, N5080, N3387);
and AND4 (N5088, N5076, N347, N2224, N3587);
and AND4 (N5089, N5088, N2720, N3653, N2595);
nor NOR3 (N5090, N5077, N958, N3123);
xor XOR2 (N5091, N5085, N3331);
not NOT1 (N5092, N5089);
or OR3 (N5093, N5086, N1197, N3517);
or OR2 (N5094, N5091, N2756);
xor XOR2 (N5095, N5094, N4946);
buf BUF1 (N5096, N5083);
xor XOR2 (N5097, N5090, N212);
or OR2 (N5098, N5097, N122);
buf BUF1 (N5099, N5095);
not NOT1 (N5100, N5092);
and AND4 (N5101, N5100, N2682, N3724, N1087);
nand NAND4 (N5102, N5098, N1698, N5046, N3807);
not NOT1 (N5103, N5101);
buf BUF1 (N5104, N5087);
nand NAND2 (N5105, N5078, N1095);
xor XOR2 (N5106, N5103, N1047);
buf BUF1 (N5107, N5036);
buf BUF1 (N5108, N5099);
xor XOR2 (N5109, N5104, N4349);
nor NOR2 (N5110, N5102, N4162);
xor XOR2 (N5111, N5107, N2530);
xor XOR2 (N5112, N5096, N2648);
nor NOR4 (N5113, N5108, N3380, N3726, N4863);
and AND4 (N5114, N5112, N2006, N2016, N1879);
nor NOR3 (N5115, N5113, N4436, N2723);
nand NAND3 (N5116, N5115, N4786, N3190);
buf BUF1 (N5117, N5057);
and AND3 (N5118, N5111, N2463, N4098);
or OR3 (N5119, N5106, N1769, N438);
nor NOR2 (N5120, N5116, N3202);
buf BUF1 (N5121, N5118);
nor NOR3 (N5122, N5117, N733, N202);
buf BUF1 (N5123, N5093);
or OR3 (N5124, N5122, N1717, N1001);
or OR2 (N5125, N5109, N2471);
nor NOR3 (N5126, N5120, N4237, N5008);
or OR3 (N5127, N5105, N3875, N1711);
and AND2 (N5128, N5114, N581);
nand NAND4 (N5129, N5125, N508, N3177, N3410);
xor XOR2 (N5130, N5126, N2160);
not NOT1 (N5131, N5081);
buf BUF1 (N5132, N5127);
not NOT1 (N5133, N5119);
buf BUF1 (N5134, N5128);
not NOT1 (N5135, N5133);
not NOT1 (N5136, N5130);
nor NOR3 (N5137, N5124, N4758, N1650);
or OR3 (N5138, N5137, N1649, N2350);
buf BUF1 (N5139, N5110);
nand NAND3 (N5140, N5138, N162, N1405);
buf BUF1 (N5141, N5139);
nand NAND3 (N5142, N5141, N1616, N4609);
nor NOR3 (N5143, N5121, N1557, N2376);
nand NAND3 (N5144, N5131, N4105, N844);
nor NOR2 (N5145, N5129, N1383);
nor NOR2 (N5146, N5144, N849);
not NOT1 (N5147, N5123);
not NOT1 (N5148, N5142);
nand NAND4 (N5149, N5140, N4582, N4040, N2651);
or OR2 (N5150, N5134, N4461);
nand NAND3 (N5151, N5148, N4270, N4068);
not NOT1 (N5152, N5145);
not NOT1 (N5153, N5135);
nand NAND3 (N5154, N5152, N983, N142);
not NOT1 (N5155, N5132);
buf BUF1 (N5156, N5146);
buf BUF1 (N5157, N5156);
buf BUF1 (N5158, N5155);
nand NAND4 (N5159, N5158, N2873, N4192, N4072);
nand NAND4 (N5160, N5136, N1155, N2928, N4972);
nor NOR3 (N5161, N5160, N3823, N2453);
or OR2 (N5162, N5150, N1196);
or OR3 (N5163, N5149, N3, N2283);
nor NOR3 (N5164, N5159, N927, N4881);
or OR4 (N5165, N5162, N5134, N3046, N1316);
not NOT1 (N5166, N5154);
or OR2 (N5167, N5161, N3004);
nand NAND4 (N5168, N5157, N1512, N4047, N432);
or OR2 (N5169, N5153, N3595);
nor NOR2 (N5170, N5143, N3051);
and AND3 (N5171, N5168, N2063, N2330);
buf BUF1 (N5172, N5164);
and AND2 (N5173, N5151, N1793);
nor NOR3 (N5174, N5173, N2927, N4692);
nand NAND3 (N5175, N5170, N1854, N2771);
xor XOR2 (N5176, N5174, N2532);
nand NAND2 (N5177, N5166, N539);
not NOT1 (N5178, N5175);
not NOT1 (N5179, N5176);
nor NOR2 (N5180, N5163, N4876);
or OR2 (N5181, N5172, N575);
xor XOR2 (N5182, N5178, N4397);
nor NOR2 (N5183, N5167, N1278);
and AND2 (N5184, N5147, N1708);
buf BUF1 (N5185, N5181);
nand NAND4 (N5186, N5184, N1012, N4896, N3834);
xor XOR2 (N5187, N5185, N3830);
not NOT1 (N5188, N5183);
not NOT1 (N5189, N5182);
nand NAND3 (N5190, N5171, N4895, N2106);
xor XOR2 (N5191, N5177, N405);
or OR3 (N5192, N5180, N4256, N3196);
buf BUF1 (N5193, N5179);
and AND4 (N5194, N5189, N3624, N4649, N2990);
not NOT1 (N5195, N5169);
nand NAND4 (N5196, N5192, N2774, N3055, N3890);
buf BUF1 (N5197, N5194);
xor XOR2 (N5198, N5187, N1927);
nand NAND3 (N5199, N5196, N2774, N807);
nor NOR4 (N5200, N5195, N4919, N1301, N3791);
xor XOR2 (N5201, N5188, N1120);
buf BUF1 (N5202, N5193);
or OR3 (N5203, N5186, N578, N3701);
nand NAND3 (N5204, N5191, N1190, N1303);
xor XOR2 (N5205, N5204, N2956);
and AND3 (N5206, N5190, N4194, N1887);
xor XOR2 (N5207, N5165, N979);
xor XOR2 (N5208, N5203, N3007);
and AND4 (N5209, N5201, N3545, N2409, N1026);
xor XOR2 (N5210, N5206, N5015);
and AND3 (N5211, N5209, N1596, N3103);
nand NAND4 (N5212, N5211, N2308, N1947, N3224);
nand NAND3 (N5213, N5205, N2904, N4035);
not NOT1 (N5214, N5210);
xor XOR2 (N5215, N5212, N1729);
nor NOR4 (N5216, N5215, N2886, N553, N3954);
not NOT1 (N5217, N5216);
nand NAND4 (N5218, N5200, N4787, N282, N2145);
and AND4 (N5219, N5218, N1026, N4820, N2251);
not NOT1 (N5220, N5217);
or OR3 (N5221, N5219, N548, N1596);
buf BUF1 (N5222, N5197);
buf BUF1 (N5223, N5220);
and AND2 (N5224, N5207, N3649);
nor NOR2 (N5225, N5223, N519);
buf BUF1 (N5226, N5225);
not NOT1 (N5227, N5202);
nor NOR3 (N5228, N5214, N1062, N43);
and AND3 (N5229, N5213, N3128, N548);
and AND2 (N5230, N5228, N2610);
nor NOR2 (N5231, N5222, N681);
and AND4 (N5232, N5231, N3642, N3761, N1806);
not NOT1 (N5233, N5224);
nor NOR2 (N5234, N5233, N871);
nand NAND2 (N5235, N5198, N4555);
xor XOR2 (N5236, N5199, N5234);
or OR2 (N5237, N2447, N3831);
or OR4 (N5238, N5230, N4066, N1421, N1536);
xor XOR2 (N5239, N5236, N2613);
not NOT1 (N5240, N5239);
xor XOR2 (N5241, N5232, N8);
or OR3 (N5242, N5237, N133, N1068);
nand NAND2 (N5243, N5221, N3167);
nor NOR2 (N5244, N5227, N1960);
nor NOR2 (N5245, N5235, N1501);
nor NOR3 (N5246, N5238, N1368, N4181);
buf BUF1 (N5247, N5208);
not NOT1 (N5248, N5240);
xor XOR2 (N5249, N5242, N1127);
and AND3 (N5250, N5226, N1764, N2080);
nor NOR3 (N5251, N5249, N1545, N4690);
xor XOR2 (N5252, N5251, N4134);
and AND2 (N5253, N5250, N2136);
or OR2 (N5254, N5229, N716);
nand NAND4 (N5255, N5246, N1674, N4530, N1407);
not NOT1 (N5256, N5244);
xor XOR2 (N5257, N5243, N2726);
nand NAND4 (N5258, N5257, N3771, N3929, N772);
nand NAND4 (N5259, N5248, N3905, N4792, N4126);
xor XOR2 (N5260, N5247, N4694);
nand NAND3 (N5261, N5259, N2160, N4160);
nand NAND4 (N5262, N5256, N2715, N5092, N4911);
buf BUF1 (N5263, N5254);
nor NOR4 (N5264, N5262, N4044, N2398, N3052);
buf BUF1 (N5265, N5263);
and AND2 (N5266, N5252, N4703);
not NOT1 (N5267, N5264);
not NOT1 (N5268, N5265);
nor NOR4 (N5269, N5258, N4667, N1186, N1178);
buf BUF1 (N5270, N5268);
and AND4 (N5271, N5260, N739, N3240, N1165);
nand NAND2 (N5272, N5269, N2473);
nor NOR3 (N5273, N5245, N5260, N557);
or OR3 (N5274, N5270, N4303, N1466);
or OR4 (N5275, N5271, N1696, N2871, N4862);
buf BUF1 (N5276, N5272);
or OR2 (N5277, N5273, N2371);
not NOT1 (N5278, N5253);
buf BUF1 (N5279, N5278);
or OR4 (N5280, N5261, N1892, N5267, N4967);
xor XOR2 (N5281, N1130, N2203);
not NOT1 (N5282, N5279);
and AND3 (N5283, N5281, N1038, N1686);
nor NOR2 (N5284, N5266, N2537);
nor NOR4 (N5285, N5283, N3444, N4359, N2283);
and AND4 (N5286, N5275, N52, N791, N841);
nand NAND4 (N5287, N5277, N3041, N179, N1439);
xor XOR2 (N5288, N5274, N3011);
and AND2 (N5289, N5241, N5170);
buf BUF1 (N5290, N5276);
and AND2 (N5291, N5255, N1363);
and AND2 (N5292, N5289, N2611);
or OR3 (N5293, N5292, N1298, N1313);
buf BUF1 (N5294, N5290);
nor NOR2 (N5295, N5284, N2615);
not NOT1 (N5296, N5280);
or OR3 (N5297, N5285, N4210, N3553);
not NOT1 (N5298, N5295);
and AND3 (N5299, N5288, N2978, N725);
nand NAND4 (N5300, N5298, N351, N1505, N949);
buf BUF1 (N5301, N5291);
buf BUF1 (N5302, N5297);
nor NOR4 (N5303, N5287, N4963, N3105, N3318);
nand NAND2 (N5304, N5286, N4642);
and AND4 (N5305, N5299, N2286, N3198, N4184);
xor XOR2 (N5306, N5296, N3021);
buf BUF1 (N5307, N5294);
nor NOR3 (N5308, N5303, N1301, N1900);
and AND2 (N5309, N5304, N3255);
xor XOR2 (N5310, N5308, N2650);
nand NAND2 (N5311, N5305, N3995);
or OR2 (N5312, N5310, N268);
xor XOR2 (N5313, N5309, N1423);
xor XOR2 (N5314, N5301, N4471);
nand NAND2 (N5315, N5307, N2585);
nor NOR2 (N5316, N5312, N5146);
not NOT1 (N5317, N5313);
nor NOR4 (N5318, N5302, N972, N2533, N1413);
buf BUF1 (N5319, N5316);
nand NAND4 (N5320, N5282, N371, N1826, N1742);
nand NAND3 (N5321, N5319, N3500, N1600);
buf BUF1 (N5322, N5293);
nor NOR4 (N5323, N5315, N3417, N2511, N2112);
xor XOR2 (N5324, N5323, N2400);
and AND3 (N5325, N5320, N883, N1652);
nand NAND2 (N5326, N5324, N4273);
or OR4 (N5327, N5322, N957, N376, N4569);
and AND3 (N5328, N5318, N3959, N2704);
and AND2 (N5329, N5328, N2062);
nor NOR4 (N5330, N5300, N637, N4, N2817);
xor XOR2 (N5331, N5330, N4129);
nand NAND3 (N5332, N5327, N746, N4177);
buf BUF1 (N5333, N5325);
buf BUF1 (N5334, N5314);
not NOT1 (N5335, N5306);
buf BUF1 (N5336, N5332);
xor XOR2 (N5337, N5336, N4154);
nand NAND3 (N5338, N5311, N1212, N3015);
xor XOR2 (N5339, N5337, N4213);
or OR4 (N5340, N5329, N3543, N974, N1870);
or OR3 (N5341, N5340, N3661, N1687);
and AND3 (N5342, N5326, N76, N3512);
not NOT1 (N5343, N5333);
and AND2 (N5344, N5335, N5199);
nand NAND2 (N5345, N5344, N3330);
xor XOR2 (N5346, N5331, N2306);
xor XOR2 (N5347, N5345, N3977);
not NOT1 (N5348, N5343);
buf BUF1 (N5349, N5334);
xor XOR2 (N5350, N5348, N4993);
nand NAND2 (N5351, N5339, N311);
not NOT1 (N5352, N5341);
nor NOR2 (N5353, N5338, N4182);
or OR4 (N5354, N5353, N113, N4317, N3413);
buf BUF1 (N5355, N5347);
nand NAND3 (N5356, N5352, N2606, N115);
xor XOR2 (N5357, N5355, N4694);
nand NAND4 (N5358, N5354, N85, N2793, N1427);
nor NOR4 (N5359, N5358, N4030, N2724, N1105);
nor NOR3 (N5360, N5342, N5302, N3312);
xor XOR2 (N5361, N5321, N3051);
or OR2 (N5362, N5361, N2235);
xor XOR2 (N5363, N5346, N3937);
buf BUF1 (N5364, N5349);
nand NAND2 (N5365, N5359, N194);
buf BUF1 (N5366, N5363);
xor XOR2 (N5367, N5357, N3203);
xor XOR2 (N5368, N5351, N3523);
not NOT1 (N5369, N5350);
or OR2 (N5370, N5367, N3943);
buf BUF1 (N5371, N5356);
and AND3 (N5372, N5370, N1952, N5231);
not NOT1 (N5373, N5372);
nor NOR2 (N5374, N5365, N5106);
xor XOR2 (N5375, N5366, N5350);
not NOT1 (N5376, N5375);
xor XOR2 (N5377, N5373, N1387);
not NOT1 (N5378, N5377);
and AND3 (N5379, N5374, N2005, N1711);
nand NAND3 (N5380, N5362, N3589, N5304);
not NOT1 (N5381, N5364);
nand NAND2 (N5382, N5317, N4243);
and AND3 (N5383, N5379, N2608, N4706);
nor NOR3 (N5384, N5378, N5158, N1917);
nand NAND4 (N5385, N5368, N701, N3549, N5339);
nor NOR3 (N5386, N5360, N868, N2888);
or OR2 (N5387, N5376, N3305);
nand NAND2 (N5388, N5380, N682);
not NOT1 (N5389, N5381);
and AND4 (N5390, N5371, N3451, N3154, N4698);
nor NOR4 (N5391, N5382, N797, N3824, N1142);
buf BUF1 (N5392, N5383);
not NOT1 (N5393, N5369);
or OR3 (N5394, N5386, N2623, N2154);
not NOT1 (N5395, N5394);
and AND3 (N5396, N5390, N3213, N655);
nor NOR2 (N5397, N5391, N2507);
and AND3 (N5398, N5393, N690, N716);
nor NOR3 (N5399, N5388, N464, N3910);
not NOT1 (N5400, N5384);
not NOT1 (N5401, N5389);
and AND2 (N5402, N5387, N1618);
buf BUF1 (N5403, N5397);
not NOT1 (N5404, N5398);
xor XOR2 (N5405, N5395, N2023);
nor NOR2 (N5406, N5401, N3077);
buf BUF1 (N5407, N5406);
not NOT1 (N5408, N5404);
buf BUF1 (N5409, N5385);
or OR3 (N5410, N5396, N2301, N300);
nand NAND3 (N5411, N5392, N4011, N3354);
not NOT1 (N5412, N5409);
not NOT1 (N5413, N5405);
or OR4 (N5414, N5399, N2258, N2040, N2710);
and AND4 (N5415, N5410, N4873, N1756, N283);
and AND2 (N5416, N5407, N440);
not NOT1 (N5417, N5415);
not NOT1 (N5418, N5413);
nor NOR3 (N5419, N5417, N840, N4789);
nor NOR3 (N5420, N5400, N1338, N4498);
nand NAND2 (N5421, N5416, N1308);
not NOT1 (N5422, N5420);
and AND2 (N5423, N5412, N2089);
nor NOR3 (N5424, N5411, N2058, N1123);
nor NOR4 (N5425, N5403, N3831, N2128, N1744);
not NOT1 (N5426, N5424);
or OR3 (N5427, N5425, N4728, N1423);
nand NAND2 (N5428, N5426, N2952);
nor NOR2 (N5429, N5408, N4479);
xor XOR2 (N5430, N5414, N3371);
nor NOR2 (N5431, N5422, N3630);
nor NOR2 (N5432, N5429, N204);
buf BUF1 (N5433, N5423);
xor XOR2 (N5434, N5428, N881);
or OR2 (N5435, N5434, N1158);
or OR2 (N5436, N5435, N1911);
and AND3 (N5437, N5421, N1049, N4921);
xor XOR2 (N5438, N5436, N2803);
buf BUF1 (N5439, N5402);
and AND4 (N5440, N5433, N3111, N5085, N5405);
and AND3 (N5441, N5432, N1313, N673);
or OR2 (N5442, N5438, N3313);
nor NOR4 (N5443, N5440, N3894, N1036, N4452);
buf BUF1 (N5444, N5441);
xor XOR2 (N5445, N5442, N4087);
buf BUF1 (N5446, N5444);
and AND2 (N5447, N5427, N5385);
or OR2 (N5448, N5419, N1548);
and AND4 (N5449, N5443, N1639, N2928, N3898);
or OR3 (N5450, N5430, N98, N1467);
not NOT1 (N5451, N5445);
nand NAND3 (N5452, N5449, N2298, N2307);
not NOT1 (N5453, N5431);
and AND4 (N5454, N5451, N4490, N3748, N1462);
or OR2 (N5455, N5450, N5448);
not NOT1 (N5456, N3149);
and AND3 (N5457, N5439, N930, N988);
and AND3 (N5458, N5454, N5326, N1618);
xor XOR2 (N5459, N5458, N896);
or OR2 (N5460, N5457, N5258);
nand NAND3 (N5461, N5460, N3598, N831);
xor XOR2 (N5462, N5446, N3079);
and AND2 (N5463, N5418, N477);
or OR4 (N5464, N5452, N1731, N4782, N5251);
xor XOR2 (N5465, N5463, N1300);
xor XOR2 (N5466, N5447, N4057);
and AND2 (N5467, N5437, N4092);
and AND3 (N5468, N5466, N1573, N417);
xor XOR2 (N5469, N5453, N170);
xor XOR2 (N5470, N5468, N3071);
xor XOR2 (N5471, N5469, N2913);
or OR4 (N5472, N5461, N2188, N1326, N199);
and AND2 (N5473, N5470, N4843);
not NOT1 (N5474, N5472);
xor XOR2 (N5475, N5464, N2178);
or OR4 (N5476, N5474, N4124, N2699, N4340);
buf BUF1 (N5477, N5476);
buf BUF1 (N5478, N5473);
buf BUF1 (N5479, N5456);
not NOT1 (N5480, N5475);
buf BUF1 (N5481, N5462);
not NOT1 (N5482, N5455);
nand NAND2 (N5483, N5467, N3155);
not NOT1 (N5484, N5459);
not NOT1 (N5485, N5481);
not NOT1 (N5486, N5482);
or OR2 (N5487, N5478, N5329);
xor XOR2 (N5488, N5484, N1337);
or OR3 (N5489, N5465, N755, N3016);
not NOT1 (N5490, N5477);
nor NOR3 (N5491, N5480, N2438, N3437);
nor NOR4 (N5492, N5479, N1834, N4756, N5409);
and AND2 (N5493, N5487, N5198);
or OR4 (N5494, N5491, N1775, N3924, N1481);
and AND2 (N5495, N5488, N5021);
and AND3 (N5496, N5490, N5036, N4945);
xor XOR2 (N5497, N5496, N4558);
not NOT1 (N5498, N5483);
xor XOR2 (N5499, N5497, N1993);
xor XOR2 (N5500, N5499, N3183);
nor NOR2 (N5501, N5500, N2243);
xor XOR2 (N5502, N5471, N5072);
not NOT1 (N5503, N5495);
xor XOR2 (N5504, N5486, N3553);
not NOT1 (N5505, N5503);
buf BUF1 (N5506, N5498);
xor XOR2 (N5507, N5505, N5053);
nor NOR3 (N5508, N5501, N5217, N2975);
xor XOR2 (N5509, N5502, N3533);
xor XOR2 (N5510, N5485, N3428);
and AND3 (N5511, N5494, N2054, N2179);
nor NOR2 (N5512, N5506, N374);
buf BUF1 (N5513, N5508);
xor XOR2 (N5514, N5493, N1487);
or OR3 (N5515, N5511, N1772, N4681);
buf BUF1 (N5516, N5509);
buf BUF1 (N5517, N5513);
nand NAND4 (N5518, N5512, N135, N594, N5506);
or OR4 (N5519, N5510, N159, N3691, N2311);
buf BUF1 (N5520, N5518);
xor XOR2 (N5521, N5517, N3871);
xor XOR2 (N5522, N5504, N5275);
and AND2 (N5523, N5521, N2995);
nor NOR2 (N5524, N5515, N3290);
and AND2 (N5525, N5523, N4981);
xor XOR2 (N5526, N5492, N5203);
nor NOR2 (N5527, N5526, N456);
not NOT1 (N5528, N5519);
nand NAND2 (N5529, N5525, N2937);
xor XOR2 (N5530, N5489, N2940);
xor XOR2 (N5531, N5524, N5148);
not NOT1 (N5532, N5516);
nor NOR4 (N5533, N5531, N4750, N5309, N5406);
not NOT1 (N5534, N5514);
buf BUF1 (N5535, N5520);
or OR3 (N5536, N5533, N1039, N4955);
not NOT1 (N5537, N5522);
not NOT1 (N5538, N5537);
not NOT1 (N5539, N5532);
or OR2 (N5540, N5528, N3332);
xor XOR2 (N5541, N5535, N2117);
or OR2 (N5542, N5538, N4109);
or OR2 (N5543, N5542, N3421);
nor NOR2 (N5544, N5541, N4536);
buf BUF1 (N5545, N5529);
nor NOR2 (N5546, N5507, N2672);
xor XOR2 (N5547, N5544, N326);
buf BUF1 (N5548, N5534);
buf BUF1 (N5549, N5536);
nand NAND2 (N5550, N5549, N1539);
xor XOR2 (N5551, N5540, N5468);
or OR3 (N5552, N5527, N955, N1179);
xor XOR2 (N5553, N5550, N5060);
xor XOR2 (N5554, N5551, N3904);
not NOT1 (N5555, N5552);
buf BUF1 (N5556, N5530);
nor NOR4 (N5557, N5553, N4785, N1551, N5515);
buf BUF1 (N5558, N5548);
or OR3 (N5559, N5558, N3221, N5279);
or OR4 (N5560, N5539, N2550, N3194, N1129);
nor NOR4 (N5561, N5557, N862, N2212, N173);
nor NOR2 (N5562, N5543, N4506);
buf BUF1 (N5563, N5547);
buf BUF1 (N5564, N5546);
or OR3 (N5565, N5555, N2982, N4643);
and AND2 (N5566, N5554, N4199);
nor NOR4 (N5567, N5566, N1132, N1024, N2710);
and AND2 (N5568, N5545, N4110);
or OR3 (N5569, N5562, N1580, N3596);
or OR3 (N5570, N5563, N4714, N5532);
or OR4 (N5571, N5559, N3053, N5563, N2811);
and AND2 (N5572, N5565, N3573);
or OR3 (N5573, N5567, N4240, N4582);
not NOT1 (N5574, N5561);
or OR3 (N5575, N5574, N2710, N1947);
xor XOR2 (N5576, N5575, N2451);
buf BUF1 (N5577, N5570);
xor XOR2 (N5578, N5556, N187);
not NOT1 (N5579, N5568);
buf BUF1 (N5580, N5564);
or OR2 (N5581, N5573, N4799);
buf BUF1 (N5582, N5580);
or OR4 (N5583, N5579, N3509, N243, N4611);
buf BUF1 (N5584, N5582);
nand NAND2 (N5585, N5569, N1880);
nor NOR4 (N5586, N5571, N1630, N139, N1365);
nor NOR4 (N5587, N5578, N2262, N1349, N201);
not NOT1 (N5588, N5560);
or OR2 (N5589, N5587, N2252);
or OR4 (N5590, N5588, N4348, N1689, N533);
xor XOR2 (N5591, N5586, N3981);
nor NOR2 (N5592, N5583, N4839);
xor XOR2 (N5593, N5592, N4613);
not NOT1 (N5594, N5590);
or OR4 (N5595, N5594, N3737, N1648, N1839);
or OR2 (N5596, N5581, N3627);
nand NAND3 (N5597, N5585, N2204, N1763);
not NOT1 (N5598, N5576);
buf BUF1 (N5599, N5593);
nor NOR3 (N5600, N5596, N839, N2551);
and AND4 (N5601, N5595, N2634, N4733, N434);
buf BUF1 (N5602, N5601);
or OR2 (N5603, N5598, N3229);
and AND3 (N5604, N5591, N2419, N3399);
or OR4 (N5605, N5600, N1460, N1701, N2381);
nand NAND4 (N5606, N5605, N3991, N780, N1952);
nand NAND2 (N5607, N5603, N1034);
or OR2 (N5608, N5572, N3468);
or OR4 (N5609, N5599, N1644, N4922, N88);
buf BUF1 (N5610, N5607);
xor XOR2 (N5611, N5604, N1047);
buf BUF1 (N5612, N5597);
xor XOR2 (N5613, N5602, N1820);
not NOT1 (N5614, N5613);
not NOT1 (N5615, N5584);
xor XOR2 (N5616, N5606, N4316);
or OR4 (N5617, N5609, N5578, N210, N1893);
not NOT1 (N5618, N5615);
and AND4 (N5619, N5611, N4490, N4509, N562);
or OR3 (N5620, N5619, N1265, N5065);
nor NOR3 (N5621, N5589, N448, N2351);
not NOT1 (N5622, N5577);
nand NAND2 (N5623, N5617, N4018);
and AND3 (N5624, N5620, N1696, N4259);
not NOT1 (N5625, N5614);
nand NAND3 (N5626, N5616, N4767, N3939);
xor XOR2 (N5627, N5624, N4147);
nand NAND3 (N5628, N5621, N4566, N3349);
not NOT1 (N5629, N5612);
xor XOR2 (N5630, N5625, N118);
nand NAND4 (N5631, N5626, N707, N399, N627);
not NOT1 (N5632, N5630);
not NOT1 (N5633, N5622);
not NOT1 (N5634, N5628);
nand NAND4 (N5635, N5631, N1893, N1657, N2407);
xor XOR2 (N5636, N5633, N5371);
xor XOR2 (N5637, N5627, N3976);
and AND3 (N5638, N5610, N4521, N2236);
xor XOR2 (N5639, N5634, N737);
nor NOR3 (N5640, N5608, N4225, N1558);
and AND4 (N5641, N5623, N2186, N2862, N2958);
nor NOR2 (N5642, N5641, N783);
nand NAND4 (N5643, N5618, N3850, N2032, N4500);
or OR4 (N5644, N5639, N2620, N1448, N1236);
nand NAND2 (N5645, N5637, N2484);
nand NAND2 (N5646, N5629, N3183);
or OR4 (N5647, N5636, N55, N366, N967);
or OR3 (N5648, N5642, N250, N2201);
and AND2 (N5649, N5632, N4060);
not NOT1 (N5650, N5648);
nor NOR2 (N5651, N5650, N185);
or OR4 (N5652, N5645, N244, N5056, N1807);
xor XOR2 (N5653, N5646, N4037);
buf BUF1 (N5654, N5643);
buf BUF1 (N5655, N5640);
xor XOR2 (N5656, N5635, N5132);
not NOT1 (N5657, N5655);
and AND3 (N5658, N5657, N863, N270);
not NOT1 (N5659, N5651);
nand NAND2 (N5660, N5638, N4751);
and AND3 (N5661, N5649, N2765, N2254);
not NOT1 (N5662, N5653);
nor NOR3 (N5663, N5654, N4397, N4408);
not NOT1 (N5664, N5656);
nor NOR2 (N5665, N5644, N5326);
not NOT1 (N5666, N5659);
not NOT1 (N5667, N5663);
not NOT1 (N5668, N5666);
and AND3 (N5669, N5647, N1317, N1013);
or OR3 (N5670, N5664, N2967, N2744);
xor XOR2 (N5671, N5665, N5626);
and AND4 (N5672, N5658, N1260, N5183, N3359);
xor XOR2 (N5673, N5661, N475);
nand NAND4 (N5674, N5670, N4666, N4823, N3166);
nand NAND3 (N5675, N5674, N3047, N2670);
or OR2 (N5676, N5652, N3972);
or OR2 (N5677, N5669, N4392);
buf BUF1 (N5678, N5671);
nor NOR3 (N5679, N5677, N3750, N1315);
not NOT1 (N5680, N5667);
nor NOR3 (N5681, N5673, N4459, N2016);
xor XOR2 (N5682, N5679, N1252);
nand NAND3 (N5683, N5682, N4239, N4334);
not NOT1 (N5684, N5683);
or OR2 (N5685, N5680, N3013);
not NOT1 (N5686, N5672);
xor XOR2 (N5687, N5676, N2261);
nor NOR4 (N5688, N5686, N318, N4233, N1581);
not NOT1 (N5689, N5688);
nand NAND2 (N5690, N5678, N3622);
nor NOR2 (N5691, N5681, N1268);
xor XOR2 (N5692, N5691, N5432);
xor XOR2 (N5693, N5660, N2207);
buf BUF1 (N5694, N5689);
buf BUF1 (N5695, N5668);
or OR3 (N5696, N5662, N1888, N3588);
xor XOR2 (N5697, N5695, N3088);
not NOT1 (N5698, N5690);
buf BUF1 (N5699, N5694);
buf BUF1 (N5700, N5687);
xor XOR2 (N5701, N5696, N3928);
not NOT1 (N5702, N5698);
nand NAND3 (N5703, N5685, N1477, N5268);
xor XOR2 (N5704, N5692, N4350);
nand NAND4 (N5705, N5675, N4698, N1380, N3191);
xor XOR2 (N5706, N5697, N4904);
and AND2 (N5707, N5693, N3884);
or OR3 (N5708, N5684, N2009, N4937);
not NOT1 (N5709, N5703);
nor NOR3 (N5710, N5702, N361, N3909);
nand NAND3 (N5711, N5705, N1167, N2562);
xor XOR2 (N5712, N5704, N4358);
or OR3 (N5713, N5707, N2242, N659);
nand NAND4 (N5714, N5709, N2975, N4409, N3609);
and AND4 (N5715, N5712, N930, N4571, N5639);
nor NOR2 (N5716, N5700, N3350);
not NOT1 (N5717, N5701);
not NOT1 (N5718, N5706);
xor XOR2 (N5719, N5715, N4174);
nor NOR2 (N5720, N5717, N5485);
nor NOR2 (N5721, N5708, N4429);
or OR4 (N5722, N5714, N2144, N4165, N5520);
nand NAND3 (N5723, N5721, N1242, N2769);
buf BUF1 (N5724, N5710);
xor XOR2 (N5725, N5713, N4594);
or OR3 (N5726, N5722, N5172, N1310);
buf BUF1 (N5727, N5726);
nand NAND2 (N5728, N5718, N5593);
nand NAND4 (N5729, N5727, N3565, N227, N2568);
or OR3 (N5730, N5729, N3513, N2529);
and AND2 (N5731, N5725, N804);
buf BUF1 (N5732, N5711);
and AND3 (N5733, N5720, N3528, N4397);
nor NOR3 (N5734, N5732, N5230, N1896);
nand NAND3 (N5735, N5734, N126, N1997);
nand NAND3 (N5736, N5716, N2332, N3730);
or OR4 (N5737, N5731, N96, N2717, N4986);
and AND4 (N5738, N5724, N3337, N4381, N5102);
buf BUF1 (N5739, N5723);
xor XOR2 (N5740, N5738, N2909);
xor XOR2 (N5741, N5719, N352);
xor XOR2 (N5742, N5728, N3206);
nor NOR4 (N5743, N5733, N468, N3971, N4094);
nor NOR3 (N5744, N5741, N2782, N696);
nor NOR3 (N5745, N5730, N4400, N3388);
or OR4 (N5746, N5744, N1013, N182, N3109);
buf BUF1 (N5747, N5740);
xor XOR2 (N5748, N5746, N5133);
buf BUF1 (N5749, N5736);
nor NOR2 (N5750, N5735, N2292);
buf BUF1 (N5751, N5699);
or OR2 (N5752, N5751, N722);
xor XOR2 (N5753, N5747, N3596);
nor NOR2 (N5754, N5737, N4677);
nor NOR4 (N5755, N5750, N4701, N3239, N2768);
nor NOR2 (N5756, N5742, N333);
or OR3 (N5757, N5743, N236, N3758);
xor XOR2 (N5758, N5754, N737);
buf BUF1 (N5759, N5758);
xor XOR2 (N5760, N5739, N1185);
and AND2 (N5761, N5749, N2299);
and AND3 (N5762, N5760, N3866, N773);
nor NOR4 (N5763, N5762, N3880, N3809, N2479);
buf BUF1 (N5764, N5757);
nor NOR3 (N5765, N5748, N2068, N2568);
xor XOR2 (N5766, N5764, N4429);
xor XOR2 (N5767, N5753, N409);
nor NOR2 (N5768, N5759, N613);
buf BUF1 (N5769, N5763);
and AND3 (N5770, N5752, N2109, N3671);
or OR2 (N5771, N5770, N4191);
not NOT1 (N5772, N5745);
nor NOR4 (N5773, N5772, N2909, N721, N4392);
xor XOR2 (N5774, N5756, N3316);
and AND4 (N5775, N5767, N4728, N3467, N2540);
buf BUF1 (N5776, N5771);
not NOT1 (N5777, N5761);
nand NAND4 (N5778, N5765, N3129, N4779, N4760);
nand NAND3 (N5779, N5766, N4678, N1658);
buf BUF1 (N5780, N5779);
xor XOR2 (N5781, N5777, N4243);
buf BUF1 (N5782, N5768);
xor XOR2 (N5783, N5774, N655);
xor XOR2 (N5784, N5783, N921);
and AND2 (N5785, N5755, N731);
nand NAND3 (N5786, N5781, N392, N4088);
xor XOR2 (N5787, N5775, N5609);
xor XOR2 (N5788, N5769, N4720);
and AND2 (N5789, N5788, N4141);
xor XOR2 (N5790, N5776, N4586);
buf BUF1 (N5791, N5786);
xor XOR2 (N5792, N5773, N4642);
or OR2 (N5793, N5787, N4489);
nor NOR2 (N5794, N5789, N2622);
xor XOR2 (N5795, N5791, N4320);
and AND2 (N5796, N5793, N4862);
buf BUF1 (N5797, N5780);
not NOT1 (N5798, N5778);
nand NAND4 (N5799, N5785, N24, N3528, N4514);
and AND3 (N5800, N5792, N3067, N4769);
buf BUF1 (N5801, N5795);
not NOT1 (N5802, N5800);
nand NAND4 (N5803, N5798, N5646, N5029, N4070);
and AND4 (N5804, N5790, N475, N3322, N4021);
nor NOR2 (N5805, N5794, N1841);
nand NAND4 (N5806, N5803, N81, N3813, N2115);
or OR2 (N5807, N5799, N181);
xor XOR2 (N5808, N5796, N1803);
nor NOR2 (N5809, N5807, N4204);
xor XOR2 (N5810, N5784, N4107);
buf BUF1 (N5811, N5805);
nand NAND4 (N5812, N5811, N696, N5646, N4481);
nor NOR4 (N5813, N5810, N4708, N701, N254);
not NOT1 (N5814, N5782);
nand NAND4 (N5815, N5813, N4738, N577, N5717);
and AND4 (N5816, N5809, N861, N5048, N2772);
or OR4 (N5817, N5797, N2657, N4702, N1074);
nor NOR2 (N5818, N5812, N3770);
not NOT1 (N5819, N5818);
and AND2 (N5820, N5819, N1051);
or OR2 (N5821, N5820, N3490);
and AND3 (N5822, N5816, N1257, N3851);
nand NAND4 (N5823, N5802, N4451, N3025, N1200);
buf BUF1 (N5824, N5814);
nand NAND3 (N5825, N5824, N1921, N2762);
nor NOR4 (N5826, N5806, N4617, N3302, N314);
not NOT1 (N5827, N5801);
buf BUF1 (N5828, N5817);
nand NAND4 (N5829, N5827, N910, N3191, N1748);
nor NOR2 (N5830, N5821, N358);
xor XOR2 (N5831, N5822, N1865);
buf BUF1 (N5832, N5808);
xor XOR2 (N5833, N5815, N1598);
and AND4 (N5834, N5831, N3633, N1727, N2399);
and AND4 (N5835, N5826, N1819, N4721, N3316);
not NOT1 (N5836, N5825);
xor XOR2 (N5837, N5832, N4464);
buf BUF1 (N5838, N5823);
xor XOR2 (N5839, N5830, N2497);
or OR4 (N5840, N5829, N4444, N2141, N783);
buf BUF1 (N5841, N5839);
and AND2 (N5842, N5834, N2304);
xor XOR2 (N5843, N5841, N2796);
nor NOR3 (N5844, N5835, N2141, N3508);
nand NAND2 (N5845, N5844, N421);
nor NOR2 (N5846, N5845, N3274);
nand NAND2 (N5847, N5846, N1556);
not NOT1 (N5848, N5840);
and AND4 (N5849, N5838, N3615, N1354, N4156);
or OR3 (N5850, N5849, N2110, N2496);
and AND4 (N5851, N5828, N2944, N4163, N809);
xor XOR2 (N5852, N5850, N4825);
buf BUF1 (N5853, N5837);
xor XOR2 (N5854, N5851, N47);
buf BUF1 (N5855, N5842);
buf BUF1 (N5856, N5853);
or OR3 (N5857, N5855, N2527, N2139);
buf BUF1 (N5858, N5847);
buf BUF1 (N5859, N5854);
buf BUF1 (N5860, N5804);
nor NOR2 (N5861, N5860, N1767);
nor NOR2 (N5862, N5852, N384);
and AND4 (N5863, N5843, N5302, N407, N4010);
or OR3 (N5864, N5857, N4848, N307);
nor NOR4 (N5865, N5864, N5437, N759, N3437);
and AND3 (N5866, N5863, N1939, N4455);
buf BUF1 (N5867, N5862);
and AND4 (N5868, N5865, N2492, N2407, N2607);
xor XOR2 (N5869, N5848, N1624);
nand NAND4 (N5870, N5858, N1414, N2379, N2442);
xor XOR2 (N5871, N5866, N378);
and AND2 (N5872, N5870, N1585);
not NOT1 (N5873, N5859);
not NOT1 (N5874, N5872);
not NOT1 (N5875, N5868);
xor XOR2 (N5876, N5856, N5845);
nand NAND4 (N5877, N5869, N2735, N2562, N2955);
nor NOR3 (N5878, N5836, N763, N1714);
buf BUF1 (N5879, N5874);
or OR2 (N5880, N5879, N365);
or OR4 (N5881, N5876, N5719, N478, N2146);
buf BUF1 (N5882, N5880);
and AND3 (N5883, N5871, N894, N2191);
buf BUF1 (N5884, N5833);
buf BUF1 (N5885, N5877);
or OR4 (N5886, N5861, N4212, N4238, N1139);
and AND3 (N5887, N5881, N3656, N166);
or OR2 (N5888, N5884, N860);
or OR3 (N5889, N5882, N4810, N3976);
xor XOR2 (N5890, N5886, N1430);
nor NOR2 (N5891, N5873, N4779);
and AND2 (N5892, N5875, N4340);
buf BUF1 (N5893, N5878);
buf BUF1 (N5894, N5888);
nand NAND2 (N5895, N5867, N1894);
xor XOR2 (N5896, N5894, N4715);
buf BUF1 (N5897, N5890);
not NOT1 (N5898, N5889);
not NOT1 (N5899, N5885);
nand NAND4 (N5900, N5897, N2830, N3086, N2888);
buf BUF1 (N5901, N5893);
and AND2 (N5902, N5895, N5375);
xor XOR2 (N5903, N5900, N1315);
nand NAND4 (N5904, N5892, N1886, N3955, N1155);
nand NAND4 (N5905, N5902, N2105, N5408, N1443);
not NOT1 (N5906, N5903);
xor XOR2 (N5907, N5891, N4842);
xor XOR2 (N5908, N5906, N1440);
or OR2 (N5909, N5901, N1425);
xor XOR2 (N5910, N5883, N5552);
nand NAND4 (N5911, N5899, N3676, N457, N4432);
buf BUF1 (N5912, N5904);
nor NOR4 (N5913, N5905, N4800, N2559, N2379);
xor XOR2 (N5914, N5896, N4265);
nor NOR3 (N5915, N5898, N5775, N3994);
xor XOR2 (N5916, N5909, N1582);
buf BUF1 (N5917, N5915);
nand NAND2 (N5918, N5908, N740);
and AND4 (N5919, N5914, N2820, N4108, N3464);
and AND3 (N5920, N5907, N1906, N2695);
and AND3 (N5921, N5916, N1735, N587);
not NOT1 (N5922, N5912);
nand NAND3 (N5923, N5919, N725, N4215);
and AND4 (N5924, N5887, N2, N4120, N5142);
and AND3 (N5925, N5910, N4044, N561);
or OR4 (N5926, N5922, N954, N2601, N4690);
xor XOR2 (N5927, N5920, N3194);
nand NAND2 (N5928, N5927, N5139);
not NOT1 (N5929, N5926);
or OR4 (N5930, N5917, N4946, N1130, N958);
buf BUF1 (N5931, N5918);
or OR2 (N5932, N5921, N2011);
not NOT1 (N5933, N5930);
or OR4 (N5934, N5925, N2979, N1927, N1247);
buf BUF1 (N5935, N5934);
buf BUF1 (N5936, N5935);
nor NOR2 (N5937, N5933, N83);
not NOT1 (N5938, N5929);
not NOT1 (N5939, N5924);
not NOT1 (N5940, N5923);
buf BUF1 (N5941, N5939);
nand NAND4 (N5942, N5938, N2944, N3375, N2145);
xor XOR2 (N5943, N5941, N5171);
nor NOR4 (N5944, N5911, N4626, N4560, N4614);
or OR4 (N5945, N5931, N5792, N72, N1151);
xor XOR2 (N5946, N5932, N3969);
nor NOR3 (N5947, N5943, N4209, N4463);
nand NAND3 (N5948, N5928, N1764, N5919);
xor XOR2 (N5949, N5944, N2966);
and AND4 (N5950, N5937, N3901, N2350, N2592);
buf BUF1 (N5951, N5949);
nand NAND2 (N5952, N5951, N1942);
and AND4 (N5953, N5945, N942, N2219, N1587);
xor XOR2 (N5954, N5948, N3342);
or OR4 (N5955, N5947, N2788, N3157, N2693);
or OR2 (N5956, N5955, N4622);
and AND3 (N5957, N5950, N2437, N5478);
and AND2 (N5958, N5954, N2795);
nand NAND3 (N5959, N5956, N721, N2993);
nor NOR3 (N5960, N5953, N1925, N1707);
and AND3 (N5961, N5957, N3147, N3532);
nor NOR2 (N5962, N5952, N1102);
and AND4 (N5963, N5960, N4320, N3132, N5348);
or OR4 (N5964, N5959, N1156, N456, N2617);
xor XOR2 (N5965, N5958, N3879);
xor XOR2 (N5966, N5940, N2889);
or OR4 (N5967, N5965, N5529, N1360, N2305);
or OR4 (N5968, N5962, N3309, N670, N5183);
buf BUF1 (N5969, N5963);
nand NAND3 (N5970, N5969, N5400, N4871);
and AND4 (N5971, N5970, N1174, N2363, N2347);
buf BUF1 (N5972, N5913);
not NOT1 (N5973, N5968);
and AND2 (N5974, N5942, N4170);
and AND4 (N5975, N5967, N4991, N2228, N3719);
and AND2 (N5976, N5973, N1098);
buf BUF1 (N5977, N5946);
buf BUF1 (N5978, N5972);
nor NOR4 (N5979, N5971, N2964, N3466, N3521);
nand NAND4 (N5980, N5966, N2014, N3280, N3423);
not NOT1 (N5981, N5961);
xor XOR2 (N5982, N5981, N2966);
nand NAND2 (N5983, N5980, N69);
buf BUF1 (N5984, N5976);
or OR4 (N5985, N5979, N5791, N1369, N4557);
nand NAND3 (N5986, N5977, N3316, N5177);
buf BUF1 (N5987, N5936);
and AND4 (N5988, N5985, N1406, N3806, N5422);
nor NOR2 (N5989, N5983, N3496);
and AND2 (N5990, N5987, N1596);
and AND2 (N5991, N5974, N3267);
not NOT1 (N5992, N5988);
nand NAND2 (N5993, N5978, N35);
nor NOR4 (N5994, N5982, N5762, N3381, N949);
or OR2 (N5995, N5994, N2904);
xor XOR2 (N5996, N5964, N1502);
xor XOR2 (N5997, N5996, N2998);
xor XOR2 (N5998, N5984, N829);
and AND2 (N5999, N5995, N1474);
nor NOR4 (N6000, N5998, N3516, N2572, N871);
xor XOR2 (N6001, N5999, N2532);
not NOT1 (N6002, N6000);
or OR3 (N6003, N5993, N2491, N5286);
not NOT1 (N6004, N5990);
nor NOR4 (N6005, N5997, N1902, N4898, N1467);
and AND4 (N6006, N6005, N5178, N4599, N2501);
not NOT1 (N6007, N5991);
xor XOR2 (N6008, N5975, N2922);
not NOT1 (N6009, N5986);
not NOT1 (N6010, N6009);
not NOT1 (N6011, N6003);
or OR4 (N6012, N6001, N644, N3474, N2937);
nor NOR2 (N6013, N6008, N4797);
buf BUF1 (N6014, N6002);
and AND3 (N6015, N6013, N2615, N1320);
nand NAND4 (N6016, N6012, N3333, N1513, N4129);
buf BUF1 (N6017, N6004);
not NOT1 (N6018, N6016);
xor XOR2 (N6019, N5989, N1657);
nand NAND2 (N6020, N6015, N1465);
or OR3 (N6021, N6011, N5829, N646);
nor NOR2 (N6022, N6006, N1788);
and AND2 (N6023, N5992, N1116);
or OR3 (N6024, N6020, N95, N2579);
nand NAND3 (N6025, N6010, N4154, N4189);
and AND2 (N6026, N6014, N998);
not NOT1 (N6027, N6026);
not NOT1 (N6028, N6018);
and AND4 (N6029, N6019, N3544, N2883, N5560);
nor NOR3 (N6030, N6007, N1748, N1401);
buf BUF1 (N6031, N6025);
xor XOR2 (N6032, N6031, N874);
xor XOR2 (N6033, N6023, N2650);
nor NOR3 (N6034, N6024, N1428, N2091);
and AND3 (N6035, N6032, N69, N1067);
xor XOR2 (N6036, N6028, N2560);
or OR2 (N6037, N6017, N3513);
not NOT1 (N6038, N6022);
and AND2 (N6039, N6027, N1412);
not NOT1 (N6040, N6038);
nor NOR3 (N6041, N6021, N149, N1814);
nor NOR2 (N6042, N6039, N834);
or OR2 (N6043, N6041, N5699);
or OR4 (N6044, N6040, N452, N1203, N991);
nand NAND3 (N6045, N6030, N3551, N3046);
nand NAND2 (N6046, N6042, N2775);
or OR2 (N6047, N6037, N4182);
and AND3 (N6048, N6045, N1306, N803);
nor NOR2 (N6049, N6048, N4968);
nor NOR3 (N6050, N6036, N3369, N743);
or OR2 (N6051, N6050, N1806);
buf BUF1 (N6052, N6029);
buf BUF1 (N6053, N6044);
or OR3 (N6054, N6053, N518, N2614);
and AND4 (N6055, N6035, N4813, N5624, N3388);
nand NAND3 (N6056, N6043, N556, N5443);
and AND2 (N6057, N6047, N6003);
buf BUF1 (N6058, N6056);
nand NAND4 (N6059, N6033, N56, N3308, N2139);
not NOT1 (N6060, N6059);
xor XOR2 (N6061, N6057, N5149);
xor XOR2 (N6062, N6055, N1783);
nor NOR4 (N6063, N6061, N1481, N825, N634);
or OR2 (N6064, N6051, N5815);
not NOT1 (N6065, N6049);
buf BUF1 (N6066, N6058);
nand NAND3 (N6067, N6060, N607, N1348);
nand NAND3 (N6068, N6063, N5025, N263);
buf BUF1 (N6069, N6066);
and AND2 (N6070, N6064, N3288);
nor NOR4 (N6071, N6067, N3409, N5692, N843);
and AND3 (N6072, N6054, N4067, N4111);
not NOT1 (N6073, N6034);
or OR4 (N6074, N6052, N2728, N2116, N4030);
buf BUF1 (N6075, N6073);
xor XOR2 (N6076, N6071, N1811);
nand NAND2 (N6077, N6070, N2122);
nand NAND4 (N6078, N6068, N1241, N4984, N5650);
xor XOR2 (N6079, N6075, N4852);
nand NAND4 (N6080, N6077, N3605, N2624, N3660);
or OR3 (N6081, N6078, N2774, N6010);
nand NAND2 (N6082, N6069, N3826);
buf BUF1 (N6083, N6080);
not NOT1 (N6084, N6072);
nor NOR2 (N6085, N6062, N4181);
and AND4 (N6086, N6074, N2676, N1080, N4737);
and AND4 (N6087, N6081, N1808, N2709, N3956);
xor XOR2 (N6088, N6087, N3556);
or OR4 (N6089, N6046, N1047, N4834, N2219);
xor XOR2 (N6090, N6084, N2234);
xor XOR2 (N6091, N6076, N3528);
nor NOR4 (N6092, N6091, N2489, N5111, N867);
nand NAND3 (N6093, N6065, N1832, N2986);
nand NAND3 (N6094, N6086, N3210, N4550);
and AND4 (N6095, N6092, N855, N2942, N1952);
nor NOR2 (N6096, N6083, N2382);
and AND2 (N6097, N6088, N4589);
not NOT1 (N6098, N6094);
and AND2 (N6099, N6093, N2402);
nor NOR4 (N6100, N6090, N1047, N1849, N2018);
or OR4 (N6101, N6095, N3664, N5625, N4280);
nand NAND2 (N6102, N6089, N63);
and AND3 (N6103, N6079, N3482, N4553);
nand NAND4 (N6104, N6098, N3298, N221, N5789);
xor XOR2 (N6105, N6099, N4647);
nor NOR2 (N6106, N6096, N1052);
and AND4 (N6107, N6085, N487, N2131, N4137);
nand NAND2 (N6108, N6101, N4471);
nor NOR3 (N6109, N6107, N3024, N2503);
and AND3 (N6110, N6104, N4661, N3998);
nor NOR3 (N6111, N6109, N1161, N4283);
nand NAND4 (N6112, N6102, N2199, N5754, N4253);
buf BUF1 (N6113, N6103);
and AND2 (N6114, N6108, N4226);
not NOT1 (N6115, N6112);
buf BUF1 (N6116, N6110);
buf BUF1 (N6117, N6115);
buf BUF1 (N6118, N6116);
xor XOR2 (N6119, N6100, N2917);
or OR2 (N6120, N6082, N5937);
or OR4 (N6121, N6106, N1552, N4088, N1253);
nand NAND2 (N6122, N6120, N4785);
nor NOR3 (N6123, N6119, N2100, N2716);
or OR3 (N6124, N6111, N4348, N2579);
xor XOR2 (N6125, N6118, N3718);
xor XOR2 (N6126, N6114, N4752);
and AND4 (N6127, N6124, N5273, N480, N3779);
buf BUF1 (N6128, N6117);
and AND2 (N6129, N6097, N4293);
and AND3 (N6130, N6113, N1806, N5527);
or OR2 (N6131, N6128, N4352);
buf BUF1 (N6132, N6125);
buf BUF1 (N6133, N6130);
nor NOR3 (N6134, N6121, N157, N1319);
and AND4 (N6135, N6126, N5153, N907, N2779);
xor XOR2 (N6136, N6129, N5212);
buf BUF1 (N6137, N6122);
not NOT1 (N6138, N6132);
nor NOR4 (N6139, N6138, N3638, N5446, N2964);
not NOT1 (N6140, N6123);
not NOT1 (N6141, N6140);
nor NOR2 (N6142, N6105, N2939);
or OR3 (N6143, N6142, N154, N1136);
nand NAND4 (N6144, N6143, N1803, N188, N1267);
buf BUF1 (N6145, N6135);
nor NOR3 (N6146, N6145, N996, N3059);
and AND2 (N6147, N6146, N2274);
nor NOR2 (N6148, N6144, N4102);
nor NOR2 (N6149, N6133, N5167);
nor NOR3 (N6150, N6136, N911, N4201);
buf BUF1 (N6151, N6131);
nor NOR4 (N6152, N6148, N2244, N1669, N4374);
buf BUF1 (N6153, N6141);
nand NAND2 (N6154, N6127, N4442);
or OR2 (N6155, N6150, N5342);
and AND4 (N6156, N6151, N4909, N1983, N1902);
nor NOR3 (N6157, N6139, N544, N3718);
buf BUF1 (N6158, N6149);
and AND3 (N6159, N6154, N2372, N5457);
not NOT1 (N6160, N6157);
or OR2 (N6161, N6153, N2681);
and AND3 (N6162, N6155, N5943, N6144);
nand NAND3 (N6163, N6152, N5769, N3206);
or OR3 (N6164, N6156, N594, N2045);
and AND2 (N6165, N6147, N1399);
nor NOR3 (N6166, N6158, N4039, N2085);
nor NOR3 (N6167, N6165, N645, N4888);
nor NOR2 (N6168, N6162, N620);
nor NOR4 (N6169, N6163, N5362, N5667, N925);
not NOT1 (N6170, N6160);
xor XOR2 (N6171, N6134, N4134);
xor XOR2 (N6172, N6168, N2073);
or OR3 (N6173, N6170, N2218, N4510);
and AND4 (N6174, N6159, N2655, N4378, N3027);
buf BUF1 (N6175, N6161);
or OR2 (N6176, N6174, N353);
nand NAND2 (N6177, N6173, N1057);
or OR4 (N6178, N6137, N2741, N2258, N883);
or OR4 (N6179, N6166, N4462, N6105, N3401);
and AND4 (N6180, N6179, N4178, N5390, N3416);
not NOT1 (N6181, N6178);
not NOT1 (N6182, N6176);
nand NAND3 (N6183, N6177, N1094, N1822);
nand NAND3 (N6184, N6175, N2718, N4929);
not NOT1 (N6185, N6172);
or OR2 (N6186, N6181, N3381);
nand NAND4 (N6187, N6164, N4838, N2411, N1486);
and AND4 (N6188, N6182, N5187, N5805, N5158);
or OR2 (N6189, N6188, N3377);
nor NOR3 (N6190, N6169, N1251, N2865);
buf BUF1 (N6191, N6167);
and AND2 (N6192, N6171, N1535);
or OR2 (N6193, N6186, N1076);
xor XOR2 (N6194, N6190, N4806);
or OR3 (N6195, N6183, N841, N2140);
nand NAND4 (N6196, N6189, N4946, N1709, N2344);
xor XOR2 (N6197, N6184, N3692);
nand NAND4 (N6198, N6191, N5000, N2692, N5952);
not NOT1 (N6199, N6193);
nand NAND4 (N6200, N6192, N2545, N1836, N2966);
nand NAND3 (N6201, N6185, N6179, N1311);
xor XOR2 (N6202, N6194, N5528);
nor NOR2 (N6203, N6187, N3297);
nand NAND4 (N6204, N6196, N1018, N4383, N3378);
and AND3 (N6205, N6203, N795, N2434);
not NOT1 (N6206, N6199);
not NOT1 (N6207, N6204);
not NOT1 (N6208, N6197);
and AND4 (N6209, N6200, N476, N5400, N702);
or OR3 (N6210, N6202, N182, N154);
buf BUF1 (N6211, N6207);
buf BUF1 (N6212, N6201);
nor NOR2 (N6213, N6211, N965);
or OR4 (N6214, N6180, N177, N5822, N1992);
buf BUF1 (N6215, N6213);
nor NOR3 (N6216, N6210, N4195, N334);
and AND4 (N6217, N6205, N1859, N2682, N3175);
nand NAND4 (N6218, N6214, N2681, N4501, N4495);
or OR3 (N6219, N6206, N1003, N1276);
or OR2 (N6220, N6209, N265);
or OR4 (N6221, N6216, N6202, N2152, N5956);
or OR2 (N6222, N6217, N4168);
nand NAND3 (N6223, N6215, N1034, N1643);
and AND3 (N6224, N6220, N1508, N4894);
not NOT1 (N6225, N6195);
nand NAND2 (N6226, N6219, N163);
or OR4 (N6227, N6225, N1670, N3846, N5125);
or OR4 (N6228, N6223, N268, N5446, N5833);
or OR4 (N6229, N6224, N3560, N2414, N4132);
or OR3 (N6230, N6221, N3496, N31);
buf BUF1 (N6231, N6226);
not NOT1 (N6232, N6230);
buf BUF1 (N6233, N6218);
xor XOR2 (N6234, N6227, N352);
buf BUF1 (N6235, N6229);
and AND2 (N6236, N6208, N1833);
and AND4 (N6237, N6228, N306, N5822, N839);
nand NAND3 (N6238, N6233, N3500, N4443);
buf BUF1 (N6239, N6238);
and AND3 (N6240, N6235, N82, N3959);
nand NAND2 (N6241, N6212, N3664);
nor NOR3 (N6242, N6240, N2406, N1970);
xor XOR2 (N6243, N6222, N2153);
not NOT1 (N6244, N6242);
not NOT1 (N6245, N6237);
not NOT1 (N6246, N6234);
not NOT1 (N6247, N6241);
not NOT1 (N6248, N6246);
or OR2 (N6249, N6236, N2080);
nor NOR4 (N6250, N6198, N5972, N405, N957);
xor XOR2 (N6251, N6250, N3261);
or OR4 (N6252, N6249, N3414, N6037, N2722);
not NOT1 (N6253, N6244);
or OR3 (N6254, N6239, N3754, N377);
xor XOR2 (N6255, N6253, N1877);
nor NOR4 (N6256, N6232, N1933, N6216, N4125);
nand NAND2 (N6257, N6251, N4979);
and AND3 (N6258, N6248, N4222, N3192);
not NOT1 (N6259, N6247);
xor XOR2 (N6260, N6256, N5236);
buf BUF1 (N6261, N6258);
nor NOR3 (N6262, N6231, N3401, N1940);
and AND2 (N6263, N6254, N27);
nand NAND2 (N6264, N6255, N1232);
buf BUF1 (N6265, N6262);
and AND4 (N6266, N6259, N1993, N1540, N6133);
buf BUF1 (N6267, N6261);
nor NOR4 (N6268, N6265, N2689, N1699, N2289);
or OR3 (N6269, N6245, N3864, N2139);
or OR2 (N6270, N6269, N3418);
or OR2 (N6271, N6264, N1989);
nand NAND3 (N6272, N6260, N6067, N4986);
buf BUF1 (N6273, N6266);
xor XOR2 (N6274, N6267, N1020);
or OR2 (N6275, N6271, N4204);
or OR4 (N6276, N6263, N1609, N6039, N1796);
not NOT1 (N6277, N6272);
or OR2 (N6278, N6270, N1146);
not NOT1 (N6279, N6273);
nand NAND3 (N6280, N6243, N1387, N5720);
and AND2 (N6281, N6274, N2531);
not NOT1 (N6282, N6257);
xor XOR2 (N6283, N6276, N2808);
not NOT1 (N6284, N6280);
or OR2 (N6285, N6275, N2928);
nor NOR3 (N6286, N6281, N2780, N3586);
and AND2 (N6287, N6284, N5629);
or OR3 (N6288, N6278, N5238, N3089);
buf BUF1 (N6289, N6283);
xor XOR2 (N6290, N6268, N4839);
not NOT1 (N6291, N6285);
nor NOR2 (N6292, N6289, N502);
nor NOR4 (N6293, N6252, N263, N1915, N4221);
xor XOR2 (N6294, N6292, N3798);
or OR2 (N6295, N6290, N3595);
nand NAND2 (N6296, N6288, N1958);
xor XOR2 (N6297, N6277, N3417);
or OR2 (N6298, N6291, N2557);
nand NAND3 (N6299, N6298, N1649, N3705);
or OR4 (N6300, N6282, N3693, N2097, N675);
nand NAND3 (N6301, N6287, N6021, N663);
not NOT1 (N6302, N6300);
nand NAND2 (N6303, N6293, N190);
nand NAND3 (N6304, N6301, N2945, N6178);
not NOT1 (N6305, N6279);
nor NOR3 (N6306, N6294, N6015, N2120);
nand NAND2 (N6307, N6303, N2479);
nor NOR2 (N6308, N6305, N5040);
and AND4 (N6309, N6306, N701, N1211, N1984);
nor NOR3 (N6310, N6286, N4583, N2245);
nor NOR2 (N6311, N6308, N1579);
nand NAND2 (N6312, N6295, N1753);
xor XOR2 (N6313, N6296, N782);
buf BUF1 (N6314, N6299);
nand NAND3 (N6315, N6312, N5385, N2807);
buf BUF1 (N6316, N6310);
xor XOR2 (N6317, N6311, N1874);
and AND3 (N6318, N6304, N4838, N2661);
nand NAND2 (N6319, N6315, N2516);
buf BUF1 (N6320, N6297);
and AND4 (N6321, N6307, N2023, N1062, N4287);
nand NAND4 (N6322, N6319, N4270, N2337, N259);
nor NOR4 (N6323, N6322, N480, N5969, N6261);
or OR4 (N6324, N6314, N3254, N5728, N1980);
not NOT1 (N6325, N6317);
nand NAND4 (N6326, N6320, N5100, N5008, N5120);
not NOT1 (N6327, N6316);
buf BUF1 (N6328, N6325);
nand NAND4 (N6329, N6302, N1781, N1255, N4614);
or OR3 (N6330, N6328, N6006, N824);
nand NAND2 (N6331, N6323, N3941);
nand NAND4 (N6332, N6330, N5558, N586, N4962);
nand NAND3 (N6333, N6326, N1295, N2862);
nor NOR2 (N6334, N6321, N6230);
not NOT1 (N6335, N6318);
nor NOR3 (N6336, N6327, N2894, N4333);
not NOT1 (N6337, N6313);
not NOT1 (N6338, N6324);
not NOT1 (N6339, N6335);
nand NAND2 (N6340, N6337, N2023);
and AND4 (N6341, N6336, N4852, N2016, N2669);
nand NAND4 (N6342, N6329, N1781, N3757, N368);
and AND4 (N6343, N6342, N6064, N2706, N4729);
or OR4 (N6344, N6333, N4261, N1261, N3837);
not NOT1 (N6345, N6332);
nand NAND3 (N6346, N6344, N534, N4659);
or OR2 (N6347, N6339, N512);
not NOT1 (N6348, N6331);
and AND4 (N6349, N6348, N1920, N5050, N4314);
nand NAND2 (N6350, N6349, N1537);
buf BUF1 (N6351, N6347);
and AND2 (N6352, N6309, N5656);
xor XOR2 (N6353, N6346, N2757);
and AND4 (N6354, N6351, N3909, N5605, N3958);
or OR4 (N6355, N6341, N704, N3494, N6305);
buf BUF1 (N6356, N6340);
or OR4 (N6357, N6352, N6006, N1317, N139);
nand NAND2 (N6358, N6353, N1132);
nor NOR3 (N6359, N6357, N1300, N3315);
xor XOR2 (N6360, N6356, N2194);
and AND4 (N6361, N6354, N2726, N1821, N2626);
or OR4 (N6362, N6350, N1779, N983, N4105);
xor XOR2 (N6363, N6362, N5366);
nand NAND4 (N6364, N6360, N3375, N3515, N3983);
buf BUF1 (N6365, N6343);
not NOT1 (N6366, N6358);
nand NAND2 (N6367, N6359, N3049);
nor NOR4 (N6368, N6334, N5487, N1745, N2403);
or OR4 (N6369, N6367, N1719, N3030, N3656);
buf BUF1 (N6370, N6363);
or OR3 (N6371, N6338, N3834, N4839);
xor XOR2 (N6372, N6355, N245);
nand NAND3 (N6373, N6371, N4075, N4169);
nand NAND4 (N6374, N6368, N6153, N5405, N4550);
xor XOR2 (N6375, N6366, N2877);
or OR3 (N6376, N6370, N271, N5777);
buf BUF1 (N6377, N6376);
nand NAND3 (N6378, N6364, N4408, N2217);
and AND2 (N6379, N6365, N1546);
or OR4 (N6380, N6361, N1211, N2874, N6198);
or OR2 (N6381, N6378, N3397);
not NOT1 (N6382, N6372);
xor XOR2 (N6383, N6375, N7);
nor NOR3 (N6384, N6380, N301, N3943);
not NOT1 (N6385, N6382);
nor NOR4 (N6386, N6381, N4494, N5603, N4223);
xor XOR2 (N6387, N6369, N3500);
xor XOR2 (N6388, N6385, N2264);
or OR3 (N6389, N6384, N6102, N2039);
buf BUF1 (N6390, N6379);
nor NOR3 (N6391, N6389, N229, N814);
nor NOR4 (N6392, N6390, N6037, N1881, N4169);
nand NAND2 (N6393, N6383, N3907);
nand NAND3 (N6394, N6391, N3696, N4929);
and AND3 (N6395, N6393, N595, N4602);
nor NOR2 (N6396, N6387, N3105);
and AND4 (N6397, N6395, N2376, N1227, N5568);
not NOT1 (N6398, N6373);
xor XOR2 (N6399, N6377, N4195);
buf BUF1 (N6400, N6345);
nand NAND2 (N6401, N6374, N2055);
or OR2 (N6402, N6388, N5310);
not NOT1 (N6403, N6401);
xor XOR2 (N6404, N6392, N1923);
xor XOR2 (N6405, N6386, N919);
nor NOR2 (N6406, N6403, N2123);
not NOT1 (N6407, N6400);
and AND3 (N6408, N6397, N1799, N6359);
or OR4 (N6409, N6407, N1718, N2305, N3386);
and AND4 (N6410, N6406, N5592, N2614, N4115);
nand NAND3 (N6411, N6410, N3619, N1822);
nor NOR2 (N6412, N6398, N2471);
nand NAND2 (N6413, N6411, N3344);
and AND4 (N6414, N6399, N3556, N134, N2421);
nor NOR4 (N6415, N6408, N258, N4538, N5045);
nand NAND2 (N6416, N6409, N3781);
not NOT1 (N6417, N6394);
nand NAND3 (N6418, N6402, N3241, N4591);
buf BUF1 (N6419, N6412);
nor NOR3 (N6420, N6405, N4169, N6170);
buf BUF1 (N6421, N6404);
not NOT1 (N6422, N6416);
nor NOR4 (N6423, N6414, N4467, N2887, N1709);
buf BUF1 (N6424, N6396);
or OR4 (N6425, N6419, N200, N482, N4329);
and AND3 (N6426, N6417, N5702, N3836);
xor XOR2 (N6427, N6423, N1441);
xor XOR2 (N6428, N6418, N1333);
or OR3 (N6429, N6428, N2020, N1865);
nand NAND4 (N6430, N6421, N4209, N3980, N450);
buf BUF1 (N6431, N6429);
nand NAND4 (N6432, N6424, N5444, N426, N4535);
or OR3 (N6433, N6432, N1667, N1878);
buf BUF1 (N6434, N6427);
nor NOR4 (N6435, N6420, N4866, N1623, N2841);
xor XOR2 (N6436, N6425, N941);
xor XOR2 (N6437, N6435, N3529);
buf BUF1 (N6438, N6431);
buf BUF1 (N6439, N6422);
nand NAND4 (N6440, N6438, N2639, N3176, N2454);
xor XOR2 (N6441, N6436, N1771);
xor XOR2 (N6442, N6433, N1974);
nand NAND4 (N6443, N6426, N5020, N1848, N6031);
nor NOR4 (N6444, N6415, N2388, N1950, N3728);
not NOT1 (N6445, N6413);
xor XOR2 (N6446, N6440, N4698);
or OR2 (N6447, N6434, N6298);
or OR2 (N6448, N6446, N5030);
not NOT1 (N6449, N6448);
buf BUF1 (N6450, N6445);
not NOT1 (N6451, N6444);
xor XOR2 (N6452, N6450, N96);
nor NOR3 (N6453, N6442, N4794, N1881);
or OR4 (N6454, N6439, N4195, N1549, N4066);
not NOT1 (N6455, N6430);
or OR3 (N6456, N6443, N4073, N3560);
buf BUF1 (N6457, N6453);
nor NOR3 (N6458, N6452, N5939, N5266);
not NOT1 (N6459, N6449);
buf BUF1 (N6460, N6458);
buf BUF1 (N6461, N6460);
xor XOR2 (N6462, N6455, N1086);
xor XOR2 (N6463, N6461, N3292);
not NOT1 (N6464, N6447);
not NOT1 (N6465, N6441);
nand NAND2 (N6466, N6454, N5992);
or OR4 (N6467, N6466, N3658, N3381, N1833);
xor XOR2 (N6468, N6437, N2527);
and AND3 (N6469, N6464, N3233, N2296);
nor NOR4 (N6470, N6457, N3367, N5095, N4233);
nor NOR4 (N6471, N6469, N4300, N2785, N5474);
buf BUF1 (N6472, N6467);
nor NOR2 (N6473, N6451, N5206);
buf BUF1 (N6474, N6468);
not NOT1 (N6475, N6462);
or OR4 (N6476, N6470, N5312, N3452, N6119);
not NOT1 (N6477, N6472);
buf BUF1 (N6478, N6476);
or OR4 (N6479, N6465, N2696, N1309, N1752);
not NOT1 (N6480, N6459);
nand NAND3 (N6481, N6463, N2206, N6034);
or OR2 (N6482, N6478, N889);
and AND2 (N6483, N6480, N3714);
nor NOR3 (N6484, N6456, N580, N1546);
not NOT1 (N6485, N6479);
nor NOR2 (N6486, N6475, N3715);
xor XOR2 (N6487, N6474, N620);
xor XOR2 (N6488, N6477, N1374);
nor NOR2 (N6489, N6473, N547);
or OR3 (N6490, N6484, N2318, N2359);
not NOT1 (N6491, N6471);
buf BUF1 (N6492, N6489);
nand NAND2 (N6493, N6486, N2569);
buf BUF1 (N6494, N6490);
or OR3 (N6495, N6481, N1326, N501);
xor XOR2 (N6496, N6491, N1104);
buf BUF1 (N6497, N6487);
and AND4 (N6498, N6494, N730, N6228, N413);
nand NAND4 (N6499, N6492, N679, N3469, N4803);
and AND2 (N6500, N6493, N5967);
nor NOR2 (N6501, N6485, N4894);
nand NAND2 (N6502, N6495, N398);
nand NAND4 (N6503, N6482, N6218, N1010, N545);
xor XOR2 (N6504, N6499, N1033);
and AND2 (N6505, N6500, N1783);
nor NOR4 (N6506, N6498, N2156, N1467, N657);
and AND4 (N6507, N6501, N3802, N5373, N5779);
nand NAND2 (N6508, N6483, N4149);
not NOT1 (N6509, N6507);
xor XOR2 (N6510, N6488, N500);
and AND4 (N6511, N6506, N2075, N102, N6135);
and AND3 (N6512, N6503, N6157, N1441);
not NOT1 (N6513, N6504);
and AND4 (N6514, N6502, N4772, N3904, N1777);
nand NAND4 (N6515, N6497, N4831, N1177, N2965);
or OR2 (N6516, N6509, N2593);
or OR4 (N6517, N6510, N5199, N1273, N5102);
or OR3 (N6518, N6513, N6465, N1972);
nand NAND3 (N6519, N6512, N6188, N4612);
not NOT1 (N6520, N6519);
not NOT1 (N6521, N6520);
not NOT1 (N6522, N6511);
xor XOR2 (N6523, N6518, N1209);
not NOT1 (N6524, N6514);
xor XOR2 (N6525, N6521, N3295);
nor NOR2 (N6526, N6516, N5375);
nor NOR4 (N6527, N6525, N6393, N5072, N3190);
nor NOR4 (N6528, N6523, N2922, N3487, N4929);
and AND3 (N6529, N6508, N1469, N5984);
buf BUF1 (N6530, N6496);
and AND3 (N6531, N6526, N1831, N466);
and AND4 (N6532, N6529, N3227, N339, N2321);
xor XOR2 (N6533, N6532, N4915);
xor XOR2 (N6534, N6505, N3374);
and AND4 (N6535, N6527, N4512, N6367, N1448);
and AND2 (N6536, N6522, N3889);
xor XOR2 (N6537, N6536, N3662);
nand NAND4 (N6538, N6535, N4183, N3584, N2885);
or OR3 (N6539, N6524, N3680, N397);
nor NOR4 (N6540, N6530, N5408, N841, N3984);
and AND4 (N6541, N6533, N6137, N4490, N6013);
nand NAND4 (N6542, N6531, N3642, N5968, N3876);
and AND3 (N6543, N6541, N5101, N3567);
buf BUF1 (N6544, N6538);
not NOT1 (N6545, N6534);
buf BUF1 (N6546, N6543);
and AND2 (N6547, N6515, N5010);
or OR3 (N6548, N6539, N2058, N3245);
nor NOR4 (N6549, N6548, N1864, N234, N5284);
buf BUF1 (N6550, N6528);
and AND2 (N6551, N6542, N3797);
buf BUF1 (N6552, N6537);
nand NAND4 (N6553, N6551, N6442, N5076, N1069);
xor XOR2 (N6554, N6546, N2951);
not NOT1 (N6555, N6547);
and AND2 (N6556, N6517, N3930);
or OR2 (N6557, N6540, N2467);
or OR2 (N6558, N6552, N6204);
nand NAND4 (N6559, N6556, N628, N2070, N4745);
or OR4 (N6560, N6544, N4298, N590, N2069);
nor NOR2 (N6561, N6553, N3399);
not NOT1 (N6562, N6559);
not NOT1 (N6563, N6555);
or OR3 (N6564, N6558, N5747, N5776);
or OR4 (N6565, N6560, N1731, N970, N4740);
buf BUF1 (N6566, N6545);
nor NOR2 (N6567, N6562, N1782);
buf BUF1 (N6568, N6549);
not NOT1 (N6569, N6566);
and AND3 (N6570, N6567, N1980, N6113);
nand NAND4 (N6571, N6568, N2458, N6013, N3254);
nor NOR3 (N6572, N6570, N2410, N3717);
buf BUF1 (N6573, N6564);
nor NOR4 (N6574, N6569, N2509, N5160, N416);
xor XOR2 (N6575, N6572, N2659);
xor XOR2 (N6576, N6561, N4568);
or OR4 (N6577, N6563, N5923, N3050, N1646);
buf BUF1 (N6578, N6557);
xor XOR2 (N6579, N6554, N1666);
nand NAND4 (N6580, N6550, N840, N3661, N4537);
nor NOR3 (N6581, N6574, N6063, N1072);
not NOT1 (N6582, N6576);
buf BUF1 (N6583, N6580);
or OR2 (N6584, N6582, N1627);
nor NOR2 (N6585, N6583, N919);
buf BUF1 (N6586, N6565);
buf BUF1 (N6587, N6579);
or OR3 (N6588, N6585, N681, N248);
buf BUF1 (N6589, N6575);
or OR3 (N6590, N6587, N2743, N1158);
or OR2 (N6591, N6584, N2878);
nor NOR3 (N6592, N6589, N3704, N4787);
nor NOR2 (N6593, N6578, N161);
not NOT1 (N6594, N6577);
xor XOR2 (N6595, N6586, N944);
nor NOR2 (N6596, N6594, N2047);
buf BUF1 (N6597, N6573);
or OR2 (N6598, N6592, N3395);
buf BUF1 (N6599, N6581);
not NOT1 (N6600, N6588);
nand NAND4 (N6601, N6590, N4114, N415, N3090);
and AND2 (N6602, N6596, N5883);
nor NOR2 (N6603, N6591, N5029);
or OR2 (N6604, N6571, N4684);
or OR2 (N6605, N6600, N2146);
nor NOR2 (N6606, N6598, N6351);
nand NAND2 (N6607, N6593, N1743);
or OR4 (N6608, N6605, N3926, N3125, N5088);
or OR4 (N6609, N6601, N6218, N402, N6016);
xor XOR2 (N6610, N6597, N1586);
nor NOR4 (N6611, N6599, N5637, N3333, N2151);
xor XOR2 (N6612, N6609, N1887);
and AND2 (N6613, N6607, N2582);
nor NOR2 (N6614, N6610, N1702);
or OR2 (N6615, N6603, N4441);
nor NOR3 (N6616, N6614, N5063, N3435);
xor XOR2 (N6617, N6612, N5088);
nand NAND4 (N6618, N6602, N3164, N2323, N3565);
xor XOR2 (N6619, N6615, N2710);
nand NAND2 (N6620, N6618, N3736);
buf BUF1 (N6621, N6604);
and AND2 (N6622, N6620, N1295);
nor NOR2 (N6623, N6595, N4531);
xor XOR2 (N6624, N6621, N5402);
buf BUF1 (N6625, N6619);
or OR2 (N6626, N6608, N1902);
or OR4 (N6627, N6625, N6527, N2430, N2424);
nor NOR2 (N6628, N6622, N2889);
nand NAND2 (N6629, N6613, N5622);
and AND3 (N6630, N6626, N1922, N945);
xor XOR2 (N6631, N6623, N4240);
buf BUF1 (N6632, N6631);
nand NAND3 (N6633, N6630, N1481, N6583);
not NOT1 (N6634, N6616);
and AND3 (N6635, N6633, N4741, N5033);
nand NAND2 (N6636, N6624, N400);
and AND2 (N6637, N6611, N2696);
or OR3 (N6638, N6635, N2090, N6220);
or OR2 (N6639, N6628, N6608);
xor XOR2 (N6640, N6617, N4349);
nor NOR3 (N6641, N6632, N2374, N485);
and AND4 (N6642, N6606, N2251, N1266, N240);
xor XOR2 (N6643, N6642, N152);
and AND2 (N6644, N6627, N184);
not NOT1 (N6645, N6641);
and AND2 (N6646, N6644, N1065);
and AND3 (N6647, N6634, N1415, N2719);
and AND3 (N6648, N6647, N2633, N5014);
xor XOR2 (N6649, N6646, N1011);
and AND3 (N6650, N6637, N3202, N6550);
and AND4 (N6651, N6640, N1191, N5686, N3799);
buf BUF1 (N6652, N6639);
and AND4 (N6653, N6650, N2026, N522, N6413);
buf BUF1 (N6654, N6651);
or OR2 (N6655, N6636, N1591);
nand NAND3 (N6656, N6629, N6023, N5531);
buf BUF1 (N6657, N6643);
and AND4 (N6658, N6657, N979, N6016, N4162);
not NOT1 (N6659, N6649);
xor XOR2 (N6660, N6654, N2798);
or OR2 (N6661, N6655, N6109);
nor NOR4 (N6662, N6653, N1187, N6376, N4353);
not NOT1 (N6663, N6661);
buf BUF1 (N6664, N6658);
buf BUF1 (N6665, N6659);
or OR2 (N6666, N6663, N262);
or OR3 (N6667, N6648, N3142, N2269);
nor NOR2 (N6668, N6656, N5504);
or OR3 (N6669, N6665, N132, N6520);
not NOT1 (N6670, N6645);
not NOT1 (N6671, N6668);
nand NAND2 (N6672, N6664, N3743);
nor NOR3 (N6673, N6669, N1884, N3615);
or OR3 (N6674, N6662, N4410, N2522);
nand NAND3 (N6675, N6660, N1872, N4866);
xor XOR2 (N6676, N6638, N6286);
buf BUF1 (N6677, N6666);
nor NOR2 (N6678, N6652, N529);
nor NOR3 (N6679, N6674, N5295, N39);
and AND4 (N6680, N6676, N3948, N2627, N988);
xor XOR2 (N6681, N6667, N1853);
nand NAND4 (N6682, N6675, N5795, N1111, N3240);
buf BUF1 (N6683, N6678);
nand NAND4 (N6684, N6670, N1357, N1766, N3682);
nand NAND4 (N6685, N6673, N1409, N1992, N3407);
not NOT1 (N6686, N6671);
or OR4 (N6687, N6682, N2722, N2001, N192);
nand NAND3 (N6688, N6686, N3217, N5863);
not NOT1 (N6689, N6688);
buf BUF1 (N6690, N6685);
and AND3 (N6691, N6672, N5038, N4732);
or OR4 (N6692, N6690, N3289, N4304, N2684);
nor NOR4 (N6693, N6677, N5557, N6114, N5107);
xor XOR2 (N6694, N6680, N3187);
nor NOR4 (N6695, N6693, N5562, N1320, N91);
or OR2 (N6696, N6689, N5113);
nand NAND3 (N6697, N6684, N5572, N2185);
and AND2 (N6698, N6691, N4751);
buf BUF1 (N6699, N6687);
not NOT1 (N6700, N6683);
or OR2 (N6701, N6692, N3983);
not NOT1 (N6702, N6700);
nor NOR2 (N6703, N6701, N6647);
or OR2 (N6704, N6694, N5685);
nor NOR4 (N6705, N6695, N4122, N5704, N6303);
nor NOR2 (N6706, N6679, N3907);
or OR2 (N6707, N6702, N3258);
xor XOR2 (N6708, N6696, N776);
xor XOR2 (N6709, N6697, N3286);
nand NAND2 (N6710, N6706, N1129);
and AND4 (N6711, N6681, N3060, N2710, N1157);
nor NOR3 (N6712, N6698, N4354, N6101);
xor XOR2 (N6713, N6710, N5746);
nand NAND3 (N6714, N6704, N3158, N89);
nor NOR2 (N6715, N6714, N6684);
not NOT1 (N6716, N6699);
nor NOR4 (N6717, N6711, N3084, N2373, N4825);
or OR2 (N6718, N6703, N3740);
not NOT1 (N6719, N6705);
xor XOR2 (N6720, N6719, N918);
and AND2 (N6721, N6709, N5257);
nor NOR2 (N6722, N6717, N4049);
buf BUF1 (N6723, N6713);
or OR4 (N6724, N6718, N2122, N4710, N125);
nor NOR2 (N6725, N6723, N551);
xor XOR2 (N6726, N6720, N595);
nor NOR3 (N6727, N6722, N2970, N4857);
and AND2 (N6728, N6708, N4335);
or OR2 (N6729, N6707, N2129);
xor XOR2 (N6730, N6712, N2313);
and AND3 (N6731, N6715, N5469, N5338);
or OR4 (N6732, N6728, N6546, N6450, N1821);
not NOT1 (N6733, N6726);
nand NAND2 (N6734, N6716, N2925);
or OR4 (N6735, N6729, N5501, N4218, N6600);
xor XOR2 (N6736, N6735, N2726);
buf BUF1 (N6737, N6732);
and AND2 (N6738, N6730, N1725);
xor XOR2 (N6739, N6721, N3433);
buf BUF1 (N6740, N6731);
or OR4 (N6741, N6737, N2766, N5910, N42);
xor XOR2 (N6742, N6740, N727);
or OR2 (N6743, N6727, N6591);
not NOT1 (N6744, N6743);
or OR2 (N6745, N6725, N3282);
nor NOR3 (N6746, N6741, N5607, N894);
and AND2 (N6747, N6724, N5372);
buf BUF1 (N6748, N6738);
buf BUF1 (N6749, N6739);
or OR3 (N6750, N6742, N5876, N3090);
or OR3 (N6751, N6744, N5080, N1664);
buf BUF1 (N6752, N6733);
xor XOR2 (N6753, N6734, N4031);
and AND2 (N6754, N6752, N6409);
buf BUF1 (N6755, N6749);
xor XOR2 (N6756, N6748, N426);
nor NOR3 (N6757, N6747, N5643, N5983);
nor NOR3 (N6758, N6745, N6176, N1224);
nor NOR2 (N6759, N6756, N6424);
nor NOR2 (N6760, N6759, N3841);
buf BUF1 (N6761, N6750);
nand NAND3 (N6762, N6758, N4131, N3681);
not NOT1 (N6763, N6761);
and AND2 (N6764, N6746, N3693);
xor XOR2 (N6765, N6762, N2348);
not NOT1 (N6766, N6764);
nand NAND2 (N6767, N6755, N5547);
xor XOR2 (N6768, N6736, N5790);
nand NAND3 (N6769, N6763, N32, N5538);
xor XOR2 (N6770, N6754, N2171);
nor NOR3 (N6771, N6753, N146, N5029);
nor NOR4 (N6772, N6757, N547, N871, N4232);
or OR4 (N6773, N6772, N1572, N4962, N1937);
nand NAND3 (N6774, N6771, N6121, N2907);
not NOT1 (N6775, N6766);
xor XOR2 (N6776, N6760, N5504);
not NOT1 (N6777, N6765);
not NOT1 (N6778, N6774);
nand NAND3 (N6779, N6768, N1269, N875);
buf BUF1 (N6780, N6769);
or OR3 (N6781, N6776, N3820, N5594);
or OR3 (N6782, N6778, N45, N210);
and AND3 (N6783, N6773, N760, N4272);
nor NOR3 (N6784, N6783, N2227, N2182);
and AND2 (N6785, N6782, N5697);
nor NOR3 (N6786, N6767, N2437, N5131);
or OR4 (N6787, N6777, N5292, N626, N2650);
nor NOR3 (N6788, N6779, N6232, N1160);
nand NAND2 (N6789, N6787, N1984);
nand NAND3 (N6790, N6788, N3531, N3612);
nand NAND4 (N6791, N6790, N5319, N5030, N1352);
nor NOR3 (N6792, N6789, N2049, N2764);
nor NOR3 (N6793, N6775, N5785, N760);
not NOT1 (N6794, N6751);
and AND4 (N6795, N6785, N4412, N5051, N4298);
xor XOR2 (N6796, N6791, N5767);
nor NOR3 (N6797, N6780, N6134, N5967);
nand NAND2 (N6798, N6792, N3032);
nor NOR2 (N6799, N6784, N1218);
nor NOR2 (N6800, N6793, N2975);
nor NOR2 (N6801, N6795, N6043);
nor NOR2 (N6802, N6797, N2499);
and AND3 (N6803, N6796, N6370, N4313);
nor NOR2 (N6804, N6770, N868);
nor NOR3 (N6805, N6803, N5781, N6420);
or OR3 (N6806, N6804, N4611, N3818);
not NOT1 (N6807, N6801);
and AND3 (N6808, N6794, N6539, N6001);
xor XOR2 (N6809, N6799, N1909);
and AND2 (N6810, N6806, N2760);
and AND2 (N6811, N6798, N2736);
xor XOR2 (N6812, N6800, N6535);
buf BUF1 (N6813, N6812);
or OR3 (N6814, N6808, N162, N612);
xor XOR2 (N6815, N6781, N1851);
not NOT1 (N6816, N6815);
nor NOR4 (N6817, N6810, N4444, N4347, N5868);
not NOT1 (N6818, N6814);
and AND3 (N6819, N6802, N5581, N1647);
and AND4 (N6820, N6807, N2073, N2511, N6812);
buf BUF1 (N6821, N6820);
or OR2 (N6822, N6821, N2392);
or OR3 (N6823, N6813, N4514, N4351);
not NOT1 (N6824, N6822);
nand NAND4 (N6825, N6816, N6479, N2015, N5513);
buf BUF1 (N6826, N6786);
and AND2 (N6827, N6811, N2427);
not NOT1 (N6828, N6818);
nand NAND2 (N6829, N6823, N176);
not NOT1 (N6830, N6825);
buf BUF1 (N6831, N6819);
or OR2 (N6832, N6831, N1570);
nor NOR4 (N6833, N6829, N2716, N3902, N3208);
buf BUF1 (N6834, N6828);
not NOT1 (N6835, N6805);
buf BUF1 (N6836, N6834);
buf BUF1 (N6837, N6817);
nand NAND3 (N6838, N6826, N365, N1260);
nand NAND2 (N6839, N6832, N5823);
nor NOR2 (N6840, N6824, N3698);
nor NOR2 (N6841, N6833, N4338);
and AND3 (N6842, N6840, N332, N626);
xor XOR2 (N6843, N6836, N511);
and AND2 (N6844, N6837, N5432);
not NOT1 (N6845, N6809);
not NOT1 (N6846, N6838);
not NOT1 (N6847, N6846);
nand NAND4 (N6848, N6839, N4844, N5477, N6627);
or OR3 (N6849, N6830, N4897, N6125);
not NOT1 (N6850, N6848);
nand NAND2 (N6851, N6849, N3423);
nor NOR2 (N6852, N6842, N5040);
nor NOR3 (N6853, N6841, N2013, N3367);
not NOT1 (N6854, N6851);
xor XOR2 (N6855, N6827, N28);
nand NAND3 (N6856, N6855, N1013, N747);
buf BUF1 (N6857, N6856);
nor NOR2 (N6858, N6854, N5318);
or OR3 (N6859, N6845, N2421, N3496);
and AND3 (N6860, N6847, N2666, N1827);
nor NOR3 (N6861, N6843, N3683, N822);
or OR4 (N6862, N6844, N5762, N3285, N3325);
or OR2 (N6863, N6862, N3170);
nand NAND2 (N6864, N6863, N595);
nand NAND4 (N6865, N6859, N2531, N71, N1654);
nor NOR2 (N6866, N6860, N582);
and AND2 (N6867, N6865, N1380);
nor NOR2 (N6868, N6852, N4184);
xor XOR2 (N6869, N6850, N1209);
nand NAND2 (N6870, N6868, N411);
or OR2 (N6871, N6864, N5188);
nand NAND4 (N6872, N6858, N4026, N1811, N3384);
or OR4 (N6873, N6872, N5402, N4845, N6828);
or OR3 (N6874, N6873, N1851, N4451);
not NOT1 (N6875, N6861);
xor XOR2 (N6876, N6870, N2947);
buf BUF1 (N6877, N6835);
nand NAND2 (N6878, N6871, N5993);
not NOT1 (N6879, N6878);
xor XOR2 (N6880, N6866, N2536);
xor XOR2 (N6881, N6869, N2637);
not NOT1 (N6882, N6867);
nor NOR3 (N6883, N6875, N374, N2342);
xor XOR2 (N6884, N6879, N3871);
and AND3 (N6885, N6883, N1913, N5884);
buf BUF1 (N6886, N6884);
or OR3 (N6887, N6877, N5559, N809);
or OR2 (N6888, N6876, N4364);
nand NAND2 (N6889, N6888, N3456);
xor XOR2 (N6890, N6881, N1504);
or OR2 (N6891, N6874, N374);
and AND2 (N6892, N6885, N5298);
and AND3 (N6893, N6891, N5757, N5199);
xor XOR2 (N6894, N6886, N1088);
and AND2 (N6895, N6894, N1473);
or OR3 (N6896, N6892, N1130, N152);
nand NAND4 (N6897, N6890, N6820, N4092, N1357);
nor NOR3 (N6898, N6893, N4573, N6025);
buf BUF1 (N6899, N6898);
nor NOR3 (N6900, N6880, N1710, N1421);
or OR2 (N6901, N6899, N1636);
nand NAND3 (N6902, N6895, N414, N4421);
nand NAND4 (N6903, N6887, N5258, N4107, N2647);
and AND3 (N6904, N6901, N5287, N4065);
xor XOR2 (N6905, N6896, N2470);
xor XOR2 (N6906, N6900, N2093);
nor NOR2 (N6907, N6905, N983);
nor NOR3 (N6908, N6904, N333, N2037);
and AND2 (N6909, N6889, N596);
or OR2 (N6910, N6908, N6229);
buf BUF1 (N6911, N6906);
nand NAND3 (N6912, N6882, N4307, N6710);
xor XOR2 (N6913, N6910, N1369);
nor NOR2 (N6914, N6903, N606);
and AND2 (N6915, N6911, N4902);
xor XOR2 (N6916, N6914, N1285);
or OR2 (N6917, N6915, N719);
xor XOR2 (N6918, N6857, N998);
not NOT1 (N6919, N6912);
xor XOR2 (N6920, N6909, N1990);
nand NAND3 (N6921, N6853, N1907, N5652);
buf BUF1 (N6922, N6902);
not NOT1 (N6923, N6917);
xor XOR2 (N6924, N6913, N4808);
not NOT1 (N6925, N6907);
not NOT1 (N6926, N6922);
nand NAND2 (N6927, N6925, N5576);
nand NAND3 (N6928, N6916, N1049, N673);
not NOT1 (N6929, N6921);
nand NAND2 (N6930, N6927, N6873);
not NOT1 (N6931, N6897);
buf BUF1 (N6932, N6918);
nand NAND2 (N6933, N6923, N2046);
or OR2 (N6934, N6932, N6012);
and AND3 (N6935, N6934, N6145, N4503);
and AND4 (N6936, N6933, N887, N2181, N651);
xor XOR2 (N6937, N6935, N3340);
nand NAND4 (N6938, N6929, N6204, N6284, N533);
nor NOR2 (N6939, N6919, N4400);
nor NOR4 (N6940, N6926, N4268, N983, N5532);
and AND2 (N6941, N6930, N6590);
xor XOR2 (N6942, N6939, N3888);
nand NAND4 (N6943, N6940, N668, N1682, N1353);
buf BUF1 (N6944, N6931);
buf BUF1 (N6945, N6937);
nor NOR3 (N6946, N6920, N5315, N6495);
nor NOR4 (N6947, N6943, N5572, N1166, N4877);
or OR2 (N6948, N6942, N4663);
or OR2 (N6949, N6928, N3582);
and AND2 (N6950, N6924, N2763);
xor XOR2 (N6951, N6948, N2787);
nor NOR3 (N6952, N6947, N1502, N2556);
buf BUF1 (N6953, N6945);
nand NAND3 (N6954, N6951, N6313, N867);
xor XOR2 (N6955, N6946, N8);
nand NAND2 (N6956, N6949, N5736);
xor XOR2 (N6957, N6941, N4953);
not NOT1 (N6958, N6952);
buf BUF1 (N6959, N6944);
or OR3 (N6960, N6957, N616, N677);
buf BUF1 (N6961, N6959);
buf BUF1 (N6962, N6956);
xor XOR2 (N6963, N6936, N5128);
nor NOR3 (N6964, N6963, N3978, N6298);
nor NOR2 (N6965, N6954, N5838);
xor XOR2 (N6966, N6962, N3572);
or OR2 (N6967, N6955, N849);
and AND2 (N6968, N6961, N50);
or OR2 (N6969, N6953, N2461);
nor NOR2 (N6970, N6969, N4678);
nor NOR2 (N6971, N6938, N2224);
nand NAND4 (N6972, N6964, N1255, N2515, N4493);
xor XOR2 (N6973, N6971, N3816);
nor NOR3 (N6974, N6967, N3496, N2602);
nor NOR4 (N6975, N6958, N1882, N3200, N3452);
nand NAND4 (N6976, N6972, N400, N4031, N16);
and AND3 (N6977, N6950, N5580, N1525);
buf BUF1 (N6978, N6974);
nand NAND2 (N6979, N6970, N6085);
nand NAND4 (N6980, N6965, N2770, N2820, N3862);
and AND3 (N6981, N6979, N5316, N5451);
nor NOR3 (N6982, N6978, N5124, N4881);
nand NAND2 (N6983, N6968, N3906);
xor XOR2 (N6984, N6983, N2452);
or OR2 (N6985, N6980, N6021);
or OR3 (N6986, N6960, N5463, N861);
or OR4 (N6987, N6985, N3878, N1512, N6718);
nand NAND4 (N6988, N6975, N1447, N6230, N5112);
and AND4 (N6989, N6988, N1680, N6591, N4766);
and AND2 (N6990, N6982, N1267);
or OR2 (N6991, N6981, N1008);
buf BUF1 (N6992, N6991);
not NOT1 (N6993, N6984);
nand NAND2 (N6994, N6993, N1751);
nand NAND3 (N6995, N6977, N3718, N3845);
nor NOR2 (N6996, N6987, N5126);
nor NOR2 (N6997, N6990, N6989);
nor NOR3 (N6998, N5136, N2166, N1710);
nand NAND3 (N6999, N6996, N6699, N2138);
nor NOR3 (N7000, N6999, N5990, N5632);
nand NAND4 (N7001, N7000, N4830, N5783, N1066);
or OR2 (N7002, N6986, N1658);
nor NOR2 (N7003, N6998, N2549);
buf BUF1 (N7004, N6995);
nand NAND2 (N7005, N7001, N6042);
xor XOR2 (N7006, N7003, N6352);
xor XOR2 (N7007, N6992, N5341);
xor XOR2 (N7008, N6997, N6278);
or OR2 (N7009, N6976, N3705);
buf BUF1 (N7010, N7009);
or OR2 (N7011, N7007, N3265);
xor XOR2 (N7012, N6994, N474);
nand NAND4 (N7013, N7008, N4243, N4281, N6671);
and AND4 (N7014, N6973, N1696, N752, N636);
and AND2 (N7015, N7004, N2590);
not NOT1 (N7016, N7005);
xor XOR2 (N7017, N7012, N821);
nand NAND2 (N7018, N7014, N4644);
nor NOR4 (N7019, N7010, N2110, N5867, N2829);
and AND2 (N7020, N7006, N205);
and AND2 (N7021, N7020, N446);
or OR3 (N7022, N7018, N6599, N3937);
or OR4 (N7023, N7011, N6232, N384, N7);
nor NOR4 (N7024, N7021, N5243, N2432, N526);
not NOT1 (N7025, N6966);
nor NOR3 (N7026, N7019, N4110, N706);
not NOT1 (N7027, N7022);
nand NAND3 (N7028, N7026, N4758, N2350);
nand NAND2 (N7029, N7024, N4222);
or OR2 (N7030, N7023, N3043);
and AND2 (N7031, N7013, N1281);
nor NOR2 (N7032, N7002, N590);
not NOT1 (N7033, N7016);
nand NAND2 (N7034, N7033, N6892);
or OR3 (N7035, N7028, N1161, N2795);
and AND3 (N7036, N7030, N3323, N1279);
nor NOR3 (N7037, N7017, N1108, N1140);
buf BUF1 (N7038, N7032);
buf BUF1 (N7039, N7029);
xor XOR2 (N7040, N7039, N5644);
nor NOR2 (N7041, N7037, N2162);
buf BUF1 (N7042, N7031);
buf BUF1 (N7043, N7035);
xor XOR2 (N7044, N7040, N5464);
not NOT1 (N7045, N7044);
or OR4 (N7046, N7038, N2645, N227, N5004);
or OR2 (N7047, N7036, N634);
buf BUF1 (N7048, N7034);
not NOT1 (N7049, N7046);
not NOT1 (N7050, N7025);
and AND2 (N7051, N7049, N2777);
nor NOR2 (N7052, N7047, N5769);
xor XOR2 (N7053, N7015, N5455);
nand NAND4 (N7054, N7043, N466, N2117, N5113);
xor XOR2 (N7055, N7051, N2312);
and AND3 (N7056, N7055, N2374, N1377);
nand NAND3 (N7057, N7052, N5093, N4280);
and AND3 (N7058, N7048, N4406, N2400);
nand NAND3 (N7059, N7045, N7045, N4775);
not NOT1 (N7060, N7027);
nor NOR2 (N7061, N7057, N315);
not NOT1 (N7062, N7042);
nand NAND2 (N7063, N7060, N3463);
xor XOR2 (N7064, N7053, N3839);
or OR2 (N7065, N7061, N2074);
buf BUF1 (N7066, N7062);
not NOT1 (N7067, N7041);
nor NOR4 (N7068, N7058, N6476, N1173, N3485);
xor XOR2 (N7069, N7066, N2071);
not NOT1 (N7070, N7067);
nor NOR3 (N7071, N7063, N279, N2630);
nor NOR4 (N7072, N7056, N1589, N5537, N380);
buf BUF1 (N7073, N7054);
buf BUF1 (N7074, N7050);
or OR4 (N7075, N7074, N7050, N6434, N6699);
buf BUF1 (N7076, N7075);
nor NOR4 (N7077, N7064, N389, N1963, N2311);
xor XOR2 (N7078, N7069, N1056);
or OR2 (N7079, N7059, N2827);
or OR2 (N7080, N7078, N4832);
buf BUF1 (N7081, N7070);
nand NAND2 (N7082, N7080, N5028);
nor NOR2 (N7083, N7072, N6781);
or OR3 (N7084, N7065, N5788, N6294);
nor NOR2 (N7085, N7082, N955);
nand NAND4 (N7086, N7083, N6144, N6211, N6493);
nor NOR2 (N7087, N7085, N2928);
not NOT1 (N7088, N7087);
not NOT1 (N7089, N7068);
and AND4 (N7090, N7073, N2749, N2772, N6354);
nor NOR2 (N7091, N7089, N4483);
or OR2 (N7092, N7071, N4508);
not NOT1 (N7093, N7092);
not NOT1 (N7094, N7093);
not NOT1 (N7095, N7079);
not NOT1 (N7096, N7076);
and AND2 (N7097, N7096, N4602);
buf BUF1 (N7098, N7086);
or OR3 (N7099, N7084, N5097, N4578);
and AND4 (N7100, N7094, N4773, N5253, N1938);
nor NOR2 (N7101, N7081, N2881);
nand NAND2 (N7102, N7100, N3412);
or OR3 (N7103, N7090, N5626, N5826);
buf BUF1 (N7104, N7101);
not NOT1 (N7105, N7097);
and AND3 (N7106, N7105, N2941, N6616);
buf BUF1 (N7107, N7077);
and AND2 (N7108, N7098, N4556);
nand NAND4 (N7109, N7088, N6761, N5312, N2003);
nand NAND4 (N7110, N7103, N3155, N902, N5168);
buf BUF1 (N7111, N7095);
xor XOR2 (N7112, N7104, N4332);
nand NAND3 (N7113, N7099, N1353, N5380);
and AND4 (N7114, N7113, N4570, N3271, N3355);
buf BUF1 (N7115, N7112);
nor NOR3 (N7116, N7115, N2145, N1438);
buf BUF1 (N7117, N7102);
buf BUF1 (N7118, N7117);
or OR4 (N7119, N7108, N4844, N1653, N1879);
and AND3 (N7120, N7116, N5352, N2136);
and AND2 (N7121, N7109, N6597);
nand NAND2 (N7122, N7118, N3049);
buf BUF1 (N7123, N7121);
buf BUF1 (N7124, N7091);
nor NOR3 (N7125, N7119, N1169, N5848);
buf BUF1 (N7126, N7124);
nand NAND2 (N7127, N7106, N5935);
buf BUF1 (N7128, N7120);
and AND4 (N7129, N7111, N918, N825, N5150);
xor XOR2 (N7130, N7122, N1406);
buf BUF1 (N7131, N7114);
and AND3 (N7132, N7127, N4934, N4304);
nor NOR4 (N7133, N7107, N6594, N7109, N6560);
buf BUF1 (N7134, N7133);
and AND3 (N7135, N7128, N679, N3588);
and AND4 (N7136, N7110, N6017, N5703, N6306);
or OR4 (N7137, N7130, N4143, N6227, N2781);
buf BUF1 (N7138, N7137);
buf BUF1 (N7139, N7131);
nor NOR3 (N7140, N7129, N803, N2930);
nand NAND4 (N7141, N7139, N5662, N6094, N3990);
not NOT1 (N7142, N7140);
not NOT1 (N7143, N7136);
and AND4 (N7144, N7132, N6, N2611, N2527);
nor NOR4 (N7145, N7126, N5430, N3009, N503);
or OR3 (N7146, N7135, N896, N3147);
not NOT1 (N7147, N7125);
nand NAND3 (N7148, N7138, N499, N592);
and AND2 (N7149, N7142, N1837);
and AND3 (N7150, N7148, N5480, N278);
buf BUF1 (N7151, N7145);
nand NAND2 (N7152, N7150, N1940);
nor NOR4 (N7153, N7152, N7089, N5902, N2688);
xor XOR2 (N7154, N7153, N5568);
and AND4 (N7155, N7154, N2530, N5776, N416);
nor NOR2 (N7156, N7155, N1096);
and AND4 (N7157, N7134, N4400, N386, N6425);
and AND4 (N7158, N7123, N5127, N4728, N1015);
not NOT1 (N7159, N7143);
nand NAND4 (N7160, N7156, N3101, N1403, N5179);
or OR3 (N7161, N7159, N6438, N3012);
xor XOR2 (N7162, N7157, N3568);
not NOT1 (N7163, N7141);
nor NOR3 (N7164, N7151, N4933, N3177);
xor XOR2 (N7165, N7144, N1110);
xor XOR2 (N7166, N7162, N4634);
and AND3 (N7167, N7146, N298, N6907);
nand NAND3 (N7168, N7147, N1472, N5898);
xor XOR2 (N7169, N7166, N1440);
nor NOR3 (N7170, N7160, N1999, N1845);
or OR4 (N7171, N7169, N5445, N2416, N5028);
nor NOR2 (N7172, N7158, N3443);
or OR3 (N7173, N7167, N232, N3190);
and AND2 (N7174, N7172, N4037);
nor NOR4 (N7175, N7165, N5349, N5453, N3821);
nor NOR4 (N7176, N7164, N6612, N4198, N1773);
nand NAND4 (N7177, N7161, N5994, N5760, N5321);
buf BUF1 (N7178, N7149);
and AND2 (N7179, N7178, N7169);
or OR4 (N7180, N7177, N5204, N6070, N6682);
and AND3 (N7181, N7163, N2061, N5014);
nor NOR4 (N7182, N7179, N427, N1254, N710);
and AND3 (N7183, N7173, N1236, N3549);
or OR4 (N7184, N7180, N5300, N5839, N3979);
buf BUF1 (N7185, N7184);
and AND3 (N7186, N7185, N4652, N5788);
nor NOR2 (N7187, N7170, N482);
or OR2 (N7188, N7187, N3745);
buf BUF1 (N7189, N7186);
nor NOR2 (N7190, N7168, N3862);
xor XOR2 (N7191, N7190, N524);
buf BUF1 (N7192, N7176);
buf BUF1 (N7193, N7183);
nand NAND4 (N7194, N7181, N2304, N3740, N4836);
not NOT1 (N7195, N7194);
not NOT1 (N7196, N7171);
nor NOR3 (N7197, N7174, N4063, N1808);
nor NOR3 (N7198, N7195, N5980, N6250);
buf BUF1 (N7199, N7197);
and AND2 (N7200, N7192, N5469);
nor NOR2 (N7201, N7188, N6635);
nand NAND2 (N7202, N7196, N2673);
not NOT1 (N7203, N7182);
and AND3 (N7204, N7191, N5419, N180);
or OR3 (N7205, N7203, N1420, N2091);
nand NAND2 (N7206, N7189, N2402);
xor XOR2 (N7207, N7202, N3631);
nor NOR3 (N7208, N7175, N6685, N439);
not NOT1 (N7209, N7206);
and AND4 (N7210, N7209, N6283, N4084, N2174);
not NOT1 (N7211, N7199);
and AND3 (N7212, N7200, N2338, N3251);
nor NOR2 (N7213, N7208, N4230);
or OR3 (N7214, N7213, N1398, N4814);
nor NOR4 (N7215, N7211, N7104, N6690, N1059);
nand NAND4 (N7216, N7215, N2411, N3397, N2089);
not NOT1 (N7217, N7205);
not NOT1 (N7218, N7204);
not NOT1 (N7219, N7207);
not NOT1 (N7220, N7214);
not NOT1 (N7221, N7219);
buf BUF1 (N7222, N7221);
or OR4 (N7223, N7193, N2298, N5425, N1644);
nor NOR3 (N7224, N7216, N5359, N5269);
and AND2 (N7225, N7210, N6283);
or OR3 (N7226, N7220, N3659, N73);
buf BUF1 (N7227, N7224);
nor NOR4 (N7228, N7223, N4424, N6918, N5950);
not NOT1 (N7229, N7225);
xor XOR2 (N7230, N7217, N3405);
and AND3 (N7231, N7227, N4152, N3641);
and AND3 (N7232, N7201, N2717, N6030);
nor NOR3 (N7233, N7226, N4849, N5617);
nand NAND2 (N7234, N7232, N1394);
xor XOR2 (N7235, N7231, N1666);
nand NAND2 (N7236, N7218, N4932);
and AND4 (N7237, N7234, N5457, N6556, N1127);
buf BUF1 (N7238, N7228);
or OR2 (N7239, N7212, N6615);
nor NOR2 (N7240, N7239, N907);
nand NAND4 (N7241, N7229, N5395, N2664, N3363);
xor XOR2 (N7242, N7241, N1651);
xor XOR2 (N7243, N7198, N6695);
nor NOR3 (N7244, N7222, N78, N1392);
or OR3 (N7245, N7237, N7104, N6779);
not NOT1 (N7246, N7245);
and AND2 (N7247, N7233, N4858);
nand NAND3 (N7248, N7243, N2734, N1777);
and AND2 (N7249, N7236, N2099);
not NOT1 (N7250, N7248);
nand NAND2 (N7251, N7235, N1278);
and AND2 (N7252, N7251, N4340);
nor NOR4 (N7253, N7247, N2903, N2465, N4173);
buf BUF1 (N7254, N7249);
buf BUF1 (N7255, N7250);
and AND2 (N7256, N7253, N2665);
nand NAND4 (N7257, N7254, N1347, N2105, N2220);
xor XOR2 (N7258, N7244, N6417);
nand NAND2 (N7259, N7252, N6235);
xor XOR2 (N7260, N7238, N3002);
nand NAND2 (N7261, N7257, N3104);
xor XOR2 (N7262, N7230, N1146);
nor NOR4 (N7263, N7255, N4447, N1674, N4429);
not NOT1 (N7264, N7240);
nor NOR4 (N7265, N7261, N3580, N3906, N7091);
nor NOR2 (N7266, N7246, N676);
or OR4 (N7267, N7266, N5406, N3022, N226);
and AND4 (N7268, N7267, N4760, N7193, N1080);
buf BUF1 (N7269, N7268);
nand NAND3 (N7270, N7262, N4867, N6720);
xor XOR2 (N7271, N7270, N2710);
buf BUF1 (N7272, N7259);
or OR4 (N7273, N7263, N5585, N1480, N6719);
and AND4 (N7274, N7264, N878, N1964, N351);
xor XOR2 (N7275, N7265, N545);
and AND2 (N7276, N7260, N1373);
xor XOR2 (N7277, N7256, N5040);
buf BUF1 (N7278, N7242);
or OR2 (N7279, N7258, N5160);
buf BUF1 (N7280, N7274);
buf BUF1 (N7281, N7280);
not NOT1 (N7282, N7272);
nand NAND3 (N7283, N7277, N3208, N5852);
not NOT1 (N7284, N7281);
nand NAND4 (N7285, N7271, N4760, N5307, N3846);
nor NOR3 (N7286, N7276, N6718, N706);
and AND2 (N7287, N7286, N5737);
buf BUF1 (N7288, N7282);
buf BUF1 (N7289, N7287);
nor NOR2 (N7290, N7269, N4935);
buf BUF1 (N7291, N7275);
or OR2 (N7292, N7278, N989);
xor XOR2 (N7293, N7290, N458);
buf BUF1 (N7294, N7285);
nand NAND4 (N7295, N7283, N4386, N904, N2247);
and AND2 (N7296, N7294, N110);
nand NAND2 (N7297, N7284, N1138);
buf BUF1 (N7298, N7292);
buf BUF1 (N7299, N7296);
buf BUF1 (N7300, N7297);
not NOT1 (N7301, N7293);
xor XOR2 (N7302, N7298, N4774);
and AND4 (N7303, N7301, N6455, N4657, N6181);
nor NOR2 (N7304, N7273, N3281);
buf BUF1 (N7305, N7289);
and AND2 (N7306, N7291, N1190);
or OR2 (N7307, N7299, N3287);
and AND2 (N7308, N7305, N458);
and AND2 (N7309, N7279, N3227);
nor NOR2 (N7310, N7304, N5333);
xor XOR2 (N7311, N7308, N4341);
and AND2 (N7312, N7302, N3916);
buf BUF1 (N7313, N7288);
xor XOR2 (N7314, N7307, N2593);
and AND2 (N7315, N7310, N4874);
and AND3 (N7316, N7314, N1189, N7168);
or OR4 (N7317, N7313, N5629, N2610, N6829);
buf BUF1 (N7318, N7309);
and AND4 (N7319, N7318, N4367, N4767, N7076);
nand NAND2 (N7320, N7319, N2965);
nor NOR4 (N7321, N7315, N355, N4543, N1384);
xor XOR2 (N7322, N7303, N5797);
and AND3 (N7323, N7311, N4211, N5184);
nor NOR2 (N7324, N7306, N6602);
buf BUF1 (N7325, N7322);
buf BUF1 (N7326, N7320);
buf BUF1 (N7327, N7295);
nor NOR2 (N7328, N7316, N4558);
or OR2 (N7329, N7328, N2740);
nor NOR3 (N7330, N7323, N307, N5086);
buf BUF1 (N7331, N7317);
and AND4 (N7332, N7321, N5489, N5826, N1882);
not NOT1 (N7333, N7331);
nor NOR3 (N7334, N7332, N3214, N6991);
or OR4 (N7335, N7330, N3281, N2502, N1671);
or OR4 (N7336, N7333, N5474, N5989, N7125);
not NOT1 (N7337, N7312);
not NOT1 (N7338, N7334);
nand NAND2 (N7339, N7335, N4106);
buf BUF1 (N7340, N7337);
nand NAND4 (N7341, N7339, N5808, N5715, N6570);
or OR3 (N7342, N7341, N1613, N6659);
buf BUF1 (N7343, N7326);
and AND4 (N7344, N7325, N2985, N2349, N112);
xor XOR2 (N7345, N7324, N5028);
and AND3 (N7346, N7340, N4811, N6203);
not NOT1 (N7347, N7345);
nand NAND3 (N7348, N7300, N6852, N7332);
xor XOR2 (N7349, N7347, N1068);
and AND2 (N7350, N7348, N3182);
buf BUF1 (N7351, N7327);
not NOT1 (N7352, N7342);
not NOT1 (N7353, N7351);
xor XOR2 (N7354, N7349, N3634);
nor NOR4 (N7355, N7350, N6239, N1415, N2843);
not NOT1 (N7356, N7352);
xor XOR2 (N7357, N7355, N5250);
or OR4 (N7358, N7354, N6236, N2150, N3909);
xor XOR2 (N7359, N7357, N4012);
and AND4 (N7360, N7358, N2884, N2811, N5810);
or OR3 (N7361, N7336, N3857, N425);
or OR3 (N7362, N7338, N3024, N4422);
not NOT1 (N7363, N7361);
xor XOR2 (N7364, N7344, N56);
and AND4 (N7365, N7356, N6920, N6639, N4946);
and AND3 (N7366, N7365, N4985, N1084);
not NOT1 (N7367, N7329);
nand NAND4 (N7368, N7364, N2881, N127, N1882);
xor XOR2 (N7369, N7362, N12);
nor NOR4 (N7370, N7346, N7012, N5457, N3810);
xor XOR2 (N7371, N7360, N3724);
buf BUF1 (N7372, N7363);
and AND4 (N7373, N7359, N1331, N5181, N1237);
buf BUF1 (N7374, N7372);
not NOT1 (N7375, N7353);
nand NAND4 (N7376, N7343, N3294, N2309, N2563);
and AND4 (N7377, N7374, N47, N1890, N6290);
xor XOR2 (N7378, N7368, N1564);
nor NOR4 (N7379, N7370, N5096, N223, N5998);
nor NOR2 (N7380, N7376, N6717);
nand NAND2 (N7381, N7371, N5394);
nand NAND4 (N7382, N7380, N5129, N68, N4510);
xor XOR2 (N7383, N7381, N3257);
and AND2 (N7384, N7366, N4418);
and AND3 (N7385, N7382, N6221, N1591);
xor XOR2 (N7386, N7383, N5579);
buf BUF1 (N7387, N7385);
xor XOR2 (N7388, N7369, N6346);
or OR4 (N7389, N7373, N3987, N5996, N7056);
xor XOR2 (N7390, N7379, N3519);
or OR4 (N7391, N7378, N6933, N7056, N7083);
not NOT1 (N7392, N7389);
nor NOR3 (N7393, N7388, N444, N17);
xor XOR2 (N7394, N7391, N7227);
buf BUF1 (N7395, N7392);
buf BUF1 (N7396, N7384);
and AND4 (N7397, N7396, N7123, N2344, N6631);
nor NOR4 (N7398, N7394, N7028, N6315, N348);
and AND4 (N7399, N7387, N4679, N7235, N4469);
nor NOR2 (N7400, N7398, N1094);
not NOT1 (N7401, N7395);
xor XOR2 (N7402, N7386, N3778);
xor XOR2 (N7403, N7393, N2679);
nand NAND2 (N7404, N7399, N3977);
buf BUF1 (N7405, N7367);
nor NOR3 (N7406, N7390, N5075, N1056);
not NOT1 (N7407, N7397);
and AND2 (N7408, N7407, N4082);
or OR4 (N7409, N7402, N3286, N5671, N4200);
buf BUF1 (N7410, N7400);
and AND2 (N7411, N7401, N6826);
and AND4 (N7412, N7406, N4660, N4421, N1983);
xor XOR2 (N7413, N7404, N4103);
nor NOR2 (N7414, N7403, N2630);
nor NOR2 (N7415, N7377, N4956);
nand NAND3 (N7416, N7408, N1692, N2296);
nor NOR4 (N7417, N7412, N6580, N6054, N1946);
xor XOR2 (N7418, N7416, N3296);
or OR2 (N7419, N7417, N689);
xor XOR2 (N7420, N7375, N5599);
xor XOR2 (N7421, N7405, N5989);
and AND2 (N7422, N7411, N1530);
nand NAND4 (N7423, N7413, N1927, N2581, N3692);
or OR3 (N7424, N7422, N6254, N3946);
nor NOR4 (N7425, N7415, N5915, N669, N1570);
xor XOR2 (N7426, N7414, N4880);
xor XOR2 (N7427, N7424, N2668);
not NOT1 (N7428, N7418);
and AND3 (N7429, N7423, N2170, N4868);
and AND2 (N7430, N7410, N478);
or OR2 (N7431, N7430, N5552);
xor XOR2 (N7432, N7429, N4499);
not NOT1 (N7433, N7432);
not NOT1 (N7434, N7420);
not NOT1 (N7435, N7434);
xor XOR2 (N7436, N7426, N6375);
nor NOR3 (N7437, N7427, N6300, N429);
nand NAND2 (N7438, N7433, N4615);
not NOT1 (N7439, N7431);
nand NAND2 (N7440, N7419, N3989);
nor NOR2 (N7441, N7428, N5195);
nor NOR3 (N7442, N7425, N952, N3306);
or OR3 (N7443, N7437, N5808, N1015);
xor XOR2 (N7444, N7443, N358);
xor XOR2 (N7445, N7421, N5698);
or OR2 (N7446, N7441, N4881);
nor NOR3 (N7447, N7445, N1964, N7242);
and AND3 (N7448, N7440, N2135, N2987);
buf BUF1 (N7449, N7435);
and AND3 (N7450, N7436, N5507, N331);
nor NOR3 (N7451, N7438, N3091, N3940);
buf BUF1 (N7452, N7449);
and AND3 (N7453, N7448, N1844, N5094);
buf BUF1 (N7454, N7446);
nand NAND3 (N7455, N7409, N5166, N5128);
or OR2 (N7456, N7451, N2717);
xor XOR2 (N7457, N7444, N5347);
nor NOR2 (N7458, N7457, N4977);
or OR4 (N7459, N7454, N5197, N4928, N1666);
nor NOR2 (N7460, N7456, N4675);
not NOT1 (N7461, N7453);
buf BUF1 (N7462, N7459);
or OR2 (N7463, N7452, N1093);
nor NOR4 (N7464, N7447, N4983, N3001, N6061);
nand NAND2 (N7465, N7461, N1114);
nand NAND2 (N7466, N7458, N3662);
and AND4 (N7467, N7466, N3929, N794, N6759);
buf BUF1 (N7468, N7442);
or OR3 (N7469, N7455, N6594, N2119);
xor XOR2 (N7470, N7462, N3254);
buf BUF1 (N7471, N7467);
nor NOR4 (N7472, N7439, N4563, N6315, N4862);
or OR4 (N7473, N7460, N5598, N4385, N1435);
xor XOR2 (N7474, N7468, N5592);
not NOT1 (N7475, N7463);
not NOT1 (N7476, N7465);
nand NAND3 (N7477, N7475, N5134, N6314);
buf BUF1 (N7478, N7472);
xor XOR2 (N7479, N7469, N7135);
buf BUF1 (N7480, N7478);
and AND2 (N7481, N7477, N3499);
buf BUF1 (N7482, N7470);
and AND2 (N7483, N7479, N2753);
and AND3 (N7484, N7480, N714, N4023);
or OR3 (N7485, N7474, N3257, N2770);
or OR3 (N7486, N7481, N1826, N3073);
buf BUF1 (N7487, N7476);
or OR2 (N7488, N7450, N551);
nand NAND4 (N7489, N7484, N4971, N2396, N5042);
nor NOR3 (N7490, N7485, N3404, N6410);
or OR4 (N7491, N7488, N1897, N5128, N1982);
buf BUF1 (N7492, N7489);
buf BUF1 (N7493, N7482);
xor XOR2 (N7494, N7490, N1822);
nand NAND3 (N7495, N7494, N7363, N5826);
nand NAND3 (N7496, N7483, N4318, N5183);
not NOT1 (N7497, N7491);
not NOT1 (N7498, N7493);
or OR2 (N7499, N7497, N3618);
and AND2 (N7500, N7496, N647);
nor NOR3 (N7501, N7499, N5252, N6683);
not NOT1 (N7502, N7495);
buf BUF1 (N7503, N7502);
and AND4 (N7504, N7487, N4951, N2447, N6968);
and AND4 (N7505, N7501, N2058, N1928, N4650);
or OR3 (N7506, N7464, N288, N2377);
buf BUF1 (N7507, N7498);
and AND2 (N7508, N7500, N2104);
and AND4 (N7509, N7503, N1903, N530, N3417);
buf BUF1 (N7510, N7486);
nand NAND3 (N7511, N7510, N3943, N2332);
buf BUF1 (N7512, N7508);
nand NAND3 (N7513, N7506, N4652, N6858);
not NOT1 (N7514, N7512);
and AND4 (N7515, N7504, N1668, N7479, N6856);
buf BUF1 (N7516, N7513);
buf BUF1 (N7517, N7514);
nand NAND3 (N7518, N7515, N3155, N1696);
nor NOR3 (N7519, N7507, N6288, N3159);
and AND2 (N7520, N7473, N3748);
nor NOR2 (N7521, N7509, N2133);
or OR2 (N7522, N7511, N1090);
or OR3 (N7523, N7516, N5469, N3488);
nor NOR2 (N7524, N7519, N1597);
buf BUF1 (N7525, N7518);
nor NOR2 (N7526, N7520, N3726);
or OR4 (N7527, N7505, N7443, N3207, N1374);
or OR3 (N7528, N7492, N3053, N4906);
not NOT1 (N7529, N7524);
nor NOR2 (N7530, N7526, N1017);
and AND4 (N7531, N7522, N2119, N5628, N7181);
buf BUF1 (N7532, N7471);
or OR3 (N7533, N7530, N4165, N668);
xor XOR2 (N7534, N7531, N3366);
nand NAND3 (N7535, N7533, N2045, N4480);
nand NAND2 (N7536, N7521, N1907);
nand NAND4 (N7537, N7517, N6704, N7440, N4655);
nor NOR3 (N7538, N7536, N6593, N7251);
and AND3 (N7539, N7525, N2996, N2448);
nand NAND2 (N7540, N7535, N2840);
xor XOR2 (N7541, N7529, N2374);
buf BUF1 (N7542, N7540);
nand NAND4 (N7543, N7541, N7426, N524, N7505);
nand NAND2 (N7544, N7528, N4127);
or OR4 (N7545, N7534, N2770, N4363, N3412);
and AND4 (N7546, N7542, N5801, N2168, N1740);
and AND3 (N7547, N7538, N308, N4630);
nand NAND3 (N7548, N7545, N3968, N1253);
and AND4 (N7549, N7544, N596, N30, N5623);
not NOT1 (N7550, N7539);
nor NOR2 (N7551, N7548, N3299);
not NOT1 (N7552, N7527);
and AND4 (N7553, N7551, N5291, N2921, N6652);
buf BUF1 (N7554, N7546);
buf BUF1 (N7555, N7532);
nand NAND4 (N7556, N7553, N6654, N6274, N767);
buf BUF1 (N7557, N7555);
not NOT1 (N7558, N7557);
nor NOR2 (N7559, N7549, N1602);
buf BUF1 (N7560, N7559);
or OR3 (N7561, N7543, N128, N5690);
nand NAND2 (N7562, N7554, N4544);
xor XOR2 (N7563, N7552, N2694);
or OR2 (N7564, N7563, N6864);
not NOT1 (N7565, N7537);
and AND3 (N7566, N7550, N3642, N7359);
and AND3 (N7567, N7561, N1777, N6184);
nand NAND4 (N7568, N7556, N4921, N512, N5190);
buf BUF1 (N7569, N7566);
or OR4 (N7570, N7523, N176, N6565, N2399);
and AND3 (N7571, N7565, N6923, N3912);
or OR2 (N7572, N7571, N7171);
not NOT1 (N7573, N7558);
nand NAND3 (N7574, N7562, N3703, N6008);
not NOT1 (N7575, N7560);
buf BUF1 (N7576, N7547);
buf BUF1 (N7577, N7575);
or OR3 (N7578, N7567, N4332, N2422);
not NOT1 (N7579, N7568);
nand NAND4 (N7580, N7579, N6849, N5382, N2890);
xor XOR2 (N7581, N7574, N1353);
buf BUF1 (N7582, N7572);
nand NAND4 (N7583, N7578, N1022, N4537, N2873);
nor NOR3 (N7584, N7564, N7061, N5728);
xor XOR2 (N7585, N7576, N526);
and AND2 (N7586, N7585, N5715);
buf BUF1 (N7587, N7582);
xor XOR2 (N7588, N7577, N1383);
nor NOR2 (N7589, N7583, N3200);
or OR4 (N7590, N7569, N7352, N4896, N5942);
nor NOR2 (N7591, N7589, N405);
or OR4 (N7592, N7580, N5391, N380, N1026);
buf BUF1 (N7593, N7581);
buf BUF1 (N7594, N7590);
nor NOR4 (N7595, N7573, N2294, N714, N4296);
nand NAND2 (N7596, N7584, N3482);
xor XOR2 (N7597, N7595, N6937);
not NOT1 (N7598, N7586);
xor XOR2 (N7599, N7594, N631);
and AND3 (N7600, N7587, N3497, N3497);
nor NOR2 (N7601, N7591, N5801);
and AND4 (N7602, N7600, N6868, N174, N4421);
or OR3 (N7603, N7601, N4025, N2252);
nor NOR3 (N7604, N7570, N3391, N3335);
buf BUF1 (N7605, N7597);
not NOT1 (N7606, N7588);
and AND3 (N7607, N7599, N1682, N4560);
nand NAND3 (N7608, N7592, N2681, N2086);
and AND2 (N7609, N7607, N5690);
not NOT1 (N7610, N7593);
nand NAND3 (N7611, N7603, N463, N4815);
not NOT1 (N7612, N7596);
nand NAND3 (N7613, N7609, N1405, N5538);
nor NOR3 (N7614, N7608, N6781, N640);
buf BUF1 (N7615, N7604);
nand NAND4 (N7616, N7602, N4784, N3370, N1597);
and AND4 (N7617, N7611, N6783, N4312, N3733);
not NOT1 (N7618, N7612);
nand NAND4 (N7619, N7605, N6870, N4918, N3246);
nand NAND4 (N7620, N7598, N5639, N3182, N2403);
xor XOR2 (N7621, N7618, N2275);
buf BUF1 (N7622, N7610);
nand NAND4 (N7623, N7613, N1428, N6860, N1379);
xor XOR2 (N7624, N7616, N6805);
and AND3 (N7625, N7621, N546, N4109);
not NOT1 (N7626, N7622);
not NOT1 (N7627, N7623);
or OR3 (N7628, N7620, N1697, N3017);
xor XOR2 (N7629, N7624, N3922);
nor NOR2 (N7630, N7617, N3077);
or OR2 (N7631, N7628, N2098);
nor NOR2 (N7632, N7626, N2684);
nand NAND4 (N7633, N7632, N3727, N6645, N2890);
or OR2 (N7634, N7619, N7048);
xor XOR2 (N7635, N7631, N7570);
buf BUF1 (N7636, N7634);
xor XOR2 (N7637, N7633, N5014);
nand NAND2 (N7638, N7614, N6558);
or OR2 (N7639, N7635, N3716);
and AND2 (N7640, N7637, N6906);
or OR3 (N7641, N7627, N1114, N6919);
nand NAND4 (N7642, N7629, N1028, N2039, N903);
nor NOR2 (N7643, N7630, N4571);
nand NAND3 (N7644, N7642, N5837, N268);
nand NAND3 (N7645, N7625, N4356, N1603);
nand NAND2 (N7646, N7606, N6667);
or OR3 (N7647, N7639, N6793, N4437);
buf BUF1 (N7648, N7646);
and AND2 (N7649, N7643, N6543);
nor NOR3 (N7650, N7640, N5469, N7637);
nor NOR4 (N7651, N7647, N154, N1500, N2489);
nor NOR4 (N7652, N7651, N7526, N5250, N1063);
and AND4 (N7653, N7638, N6647, N1468, N3912);
xor XOR2 (N7654, N7648, N3552);
not NOT1 (N7655, N7645);
not NOT1 (N7656, N7652);
or OR4 (N7657, N7615, N349, N7546, N6205);
nand NAND4 (N7658, N7644, N5389, N1109, N2283);
and AND2 (N7659, N7653, N192);
or OR3 (N7660, N7636, N3428, N6663);
nor NOR3 (N7661, N7656, N5409, N355);
nand NAND3 (N7662, N7649, N6699, N4951);
or OR4 (N7663, N7662, N1224, N69, N3292);
and AND2 (N7664, N7660, N4995);
buf BUF1 (N7665, N7641);
and AND4 (N7666, N7663, N4432, N5809, N2302);
nor NOR2 (N7667, N7654, N6544);
and AND2 (N7668, N7667, N4759);
buf BUF1 (N7669, N7650);
not NOT1 (N7670, N7661);
or OR3 (N7671, N7658, N5935, N1812);
buf BUF1 (N7672, N7657);
nand NAND3 (N7673, N7670, N3533, N3278);
buf BUF1 (N7674, N7673);
not NOT1 (N7675, N7672);
buf BUF1 (N7676, N7674);
or OR2 (N7677, N7675, N1066);
not NOT1 (N7678, N7665);
nor NOR3 (N7679, N7659, N7516, N6130);
not NOT1 (N7680, N7664);
xor XOR2 (N7681, N7668, N3226);
and AND2 (N7682, N7680, N6943);
and AND2 (N7683, N7677, N6945);
nor NOR2 (N7684, N7671, N395);
buf BUF1 (N7685, N7676);
xor XOR2 (N7686, N7682, N3206);
xor XOR2 (N7687, N7686, N4660);
xor XOR2 (N7688, N7684, N629);
nand NAND2 (N7689, N7681, N6387);
nor NOR4 (N7690, N7688, N6547, N1844, N7677);
nor NOR4 (N7691, N7666, N6086, N3295, N4948);
and AND4 (N7692, N7685, N1957, N3989, N4285);
or OR2 (N7693, N7687, N3266);
nand NAND3 (N7694, N7679, N4141, N5624);
or OR4 (N7695, N7691, N5548, N4667, N885);
not NOT1 (N7696, N7693);
and AND4 (N7697, N7695, N3551, N366, N5911);
or OR2 (N7698, N7692, N130);
nor NOR4 (N7699, N7697, N2248, N1303, N3318);
buf BUF1 (N7700, N7689);
not NOT1 (N7701, N7698);
xor XOR2 (N7702, N7701, N6637);
nand NAND3 (N7703, N7699, N5338, N5066);
or OR2 (N7704, N7655, N6011);
and AND4 (N7705, N7703, N6346, N1811, N7220);
buf BUF1 (N7706, N7678);
not NOT1 (N7707, N7700);
or OR4 (N7708, N7704, N5826, N532, N377);
and AND4 (N7709, N7694, N2084, N297, N2812);
buf BUF1 (N7710, N7708);
not NOT1 (N7711, N7683);
or OR2 (N7712, N7707, N7079);
nand NAND4 (N7713, N7711, N3928, N5749, N3626);
nor NOR4 (N7714, N7696, N1461, N6490, N757);
nor NOR3 (N7715, N7702, N4214, N2850);
buf BUF1 (N7716, N7715);
nand NAND2 (N7717, N7705, N4994);
nand NAND4 (N7718, N7712, N1720, N1774, N1761);
xor XOR2 (N7719, N7706, N6761);
not NOT1 (N7720, N7718);
nor NOR4 (N7721, N7716, N1789, N407, N3355);
nand NAND3 (N7722, N7717, N73, N5313);
xor XOR2 (N7723, N7690, N2876);
not NOT1 (N7724, N7709);
nand NAND3 (N7725, N7724, N4728, N252);
or OR2 (N7726, N7713, N4700);
nor NOR2 (N7727, N7669, N6549);
nand NAND3 (N7728, N7722, N3704, N2853);
and AND3 (N7729, N7719, N1231, N7526);
nor NOR2 (N7730, N7710, N4725);
xor XOR2 (N7731, N7725, N94);
xor XOR2 (N7732, N7721, N1948);
not NOT1 (N7733, N7720);
nor NOR3 (N7734, N7727, N1563, N1346);
xor XOR2 (N7735, N7714, N5642);
nand NAND2 (N7736, N7726, N7603);
xor XOR2 (N7737, N7728, N6988);
xor XOR2 (N7738, N7730, N761);
nor NOR4 (N7739, N7734, N3017, N4607, N1328);
nand NAND2 (N7740, N7733, N5483);
and AND2 (N7741, N7740, N3108);
buf BUF1 (N7742, N7729);
xor XOR2 (N7743, N7735, N3864);
nand NAND2 (N7744, N7741, N4578);
or OR4 (N7745, N7723, N1086, N6858, N253);
xor XOR2 (N7746, N7744, N714);
and AND3 (N7747, N7736, N5416, N3556);
or OR4 (N7748, N7743, N5774, N1455, N7557);
buf BUF1 (N7749, N7742);
nor NOR3 (N7750, N7738, N437, N5284);
xor XOR2 (N7751, N7745, N2545);
xor XOR2 (N7752, N7751, N2674);
not NOT1 (N7753, N7732);
and AND4 (N7754, N7737, N1388, N4652, N6890);
not NOT1 (N7755, N7748);
buf BUF1 (N7756, N7747);
not NOT1 (N7757, N7756);
or OR3 (N7758, N7752, N4309, N768);
nand NAND3 (N7759, N7739, N6564, N518);
nand NAND2 (N7760, N7757, N7637);
nand NAND3 (N7761, N7746, N826, N4077);
not NOT1 (N7762, N7755);
nand NAND2 (N7763, N7762, N252);
not NOT1 (N7764, N7759);
buf BUF1 (N7765, N7754);
nand NAND3 (N7766, N7758, N1438, N3037);
nand NAND2 (N7767, N7760, N6360);
xor XOR2 (N7768, N7764, N2334);
buf BUF1 (N7769, N7731);
and AND3 (N7770, N7753, N3470, N840);
nor NOR3 (N7771, N7765, N2511, N995);
xor XOR2 (N7772, N7767, N5594);
xor XOR2 (N7773, N7770, N603);
or OR4 (N7774, N7773, N239, N7385, N7151);
nor NOR2 (N7775, N7766, N7390);
nand NAND2 (N7776, N7772, N6556);
not NOT1 (N7777, N7768);
nor NOR3 (N7778, N7749, N5233, N166);
buf BUF1 (N7779, N7775);
and AND2 (N7780, N7776, N6289);
nor NOR4 (N7781, N7778, N3471, N7457, N1090);
buf BUF1 (N7782, N7750);
nor NOR3 (N7783, N7771, N4356, N830);
nand NAND4 (N7784, N7780, N5319, N275, N1199);
and AND2 (N7785, N7763, N570);
xor XOR2 (N7786, N7782, N5839);
xor XOR2 (N7787, N7774, N2880);
xor XOR2 (N7788, N7777, N5880);
nor NOR2 (N7789, N7761, N1178);
or OR3 (N7790, N7789, N1139, N3122);
not NOT1 (N7791, N7781);
nand NAND4 (N7792, N7769, N13, N299, N7231);
buf BUF1 (N7793, N7786);
xor XOR2 (N7794, N7783, N2987);
nand NAND4 (N7795, N7790, N4145, N3864, N4663);
and AND4 (N7796, N7794, N569, N1669, N3681);
or OR2 (N7797, N7785, N4877);
not NOT1 (N7798, N7791);
buf BUF1 (N7799, N7797);
xor XOR2 (N7800, N7787, N7183);
buf BUF1 (N7801, N7793);
nor NOR4 (N7802, N7798, N1798, N4064, N6354);
not NOT1 (N7803, N7802);
and AND3 (N7804, N7779, N281, N3590);
not NOT1 (N7805, N7803);
or OR3 (N7806, N7805, N7320, N968);
nand NAND2 (N7807, N7796, N3891);
xor XOR2 (N7808, N7804, N4673);
nor NOR4 (N7809, N7799, N7746, N1744, N7061);
not NOT1 (N7810, N7801);
not NOT1 (N7811, N7795);
buf BUF1 (N7812, N7808);
and AND4 (N7813, N7806, N5681, N5595, N170);
and AND4 (N7814, N7810, N4352, N1906, N2099);
buf BUF1 (N7815, N7792);
and AND3 (N7816, N7809, N4054, N7633);
nor NOR2 (N7817, N7788, N2422);
nand NAND4 (N7818, N7784, N4963, N7160, N404);
nand NAND3 (N7819, N7811, N1241, N6767);
nor NOR2 (N7820, N7815, N4769);
or OR4 (N7821, N7816, N6168, N4949, N6159);
not NOT1 (N7822, N7817);
nand NAND3 (N7823, N7813, N526, N1126);
nor NOR2 (N7824, N7821, N2226);
not NOT1 (N7825, N7800);
xor XOR2 (N7826, N7825, N4760);
not NOT1 (N7827, N7826);
or OR3 (N7828, N7807, N2168, N4618);
or OR4 (N7829, N7820, N4614, N1442, N3639);
xor XOR2 (N7830, N7812, N3541);
nand NAND3 (N7831, N7827, N7537, N1989);
and AND2 (N7832, N7830, N7043);
buf BUF1 (N7833, N7822);
and AND4 (N7834, N7829, N2748, N5726, N7133);
or OR4 (N7835, N7833, N6272, N6691, N869);
nor NOR4 (N7836, N7814, N3922, N3789, N53);
or OR4 (N7837, N7819, N5274, N2799, N2174);
and AND2 (N7838, N7836, N1502);
nor NOR2 (N7839, N7828, N5819);
xor XOR2 (N7840, N7823, N5362);
or OR2 (N7841, N7835, N835);
buf BUF1 (N7842, N7834);
or OR2 (N7843, N7842, N3588);
not NOT1 (N7844, N7838);
or OR2 (N7845, N7839, N39);
xor XOR2 (N7846, N7845, N2455);
nor NOR4 (N7847, N7843, N1202, N944, N3595);
nor NOR2 (N7848, N7831, N4998);
nand NAND4 (N7849, N7818, N5499, N7077, N6883);
nand NAND4 (N7850, N7832, N1866, N3004, N1192);
nand NAND4 (N7851, N7849, N5380, N6166, N2175);
xor XOR2 (N7852, N7847, N6477);
xor XOR2 (N7853, N7848, N1238);
or OR4 (N7854, N7846, N7350, N4322, N1280);
xor XOR2 (N7855, N7851, N5579);
not NOT1 (N7856, N7853);
nor NOR2 (N7857, N7841, N6022);
nor NOR2 (N7858, N7857, N1180);
or OR2 (N7859, N7840, N5626);
and AND4 (N7860, N7844, N2546, N780, N426);
or OR2 (N7861, N7850, N1741);
and AND3 (N7862, N7837, N2382, N5792);
nand NAND2 (N7863, N7824, N5044);
buf BUF1 (N7864, N7852);
nor NOR3 (N7865, N7862, N6225, N5606);
xor XOR2 (N7866, N7864, N5106);
and AND3 (N7867, N7858, N5172, N876);
or OR4 (N7868, N7859, N4051, N1411, N1390);
xor XOR2 (N7869, N7860, N874);
nor NOR3 (N7870, N7855, N2869, N5364);
not NOT1 (N7871, N7869);
xor XOR2 (N7872, N7866, N6686);
nand NAND3 (N7873, N7868, N4384, N187);
nor NOR2 (N7874, N7854, N6532);
nand NAND2 (N7875, N7874, N4328);
buf BUF1 (N7876, N7865);
or OR4 (N7877, N7875, N2884, N6326, N4768);
nand NAND4 (N7878, N7863, N4909, N2380, N7761);
and AND2 (N7879, N7861, N4594);
and AND4 (N7880, N7873, N5358, N7535, N4468);
not NOT1 (N7881, N7878);
buf BUF1 (N7882, N7871);
and AND3 (N7883, N7882, N5294, N1666);
or OR4 (N7884, N7883, N2117, N5066, N1954);
nor NOR4 (N7885, N7880, N2781, N1510, N2864);
not NOT1 (N7886, N7879);
or OR4 (N7887, N7885, N5309, N6823, N776);
and AND4 (N7888, N7884, N4406, N2181, N3579);
not NOT1 (N7889, N7867);
buf BUF1 (N7890, N7888);
or OR4 (N7891, N7890, N7257, N255, N3936);
nor NOR2 (N7892, N7881, N5151);
buf BUF1 (N7893, N7870);
and AND4 (N7894, N7876, N522, N4740, N3933);
buf BUF1 (N7895, N7889);
not NOT1 (N7896, N7892);
or OR2 (N7897, N7896, N6292);
and AND3 (N7898, N7894, N1652, N1587);
buf BUF1 (N7899, N7893);
and AND4 (N7900, N7872, N4705, N2260, N2199);
or OR3 (N7901, N7877, N2800, N4729);
buf BUF1 (N7902, N7899);
buf BUF1 (N7903, N7895);
or OR2 (N7904, N7902, N530);
or OR3 (N7905, N7897, N5356, N1410);
or OR2 (N7906, N7905, N7403);
xor XOR2 (N7907, N7904, N1195);
buf BUF1 (N7908, N7903);
or OR2 (N7909, N7887, N2210);
buf BUF1 (N7910, N7909);
or OR3 (N7911, N7908, N1455, N1314);
xor XOR2 (N7912, N7907, N4058);
or OR4 (N7913, N7891, N1915, N3576, N4817);
nand NAND4 (N7914, N7901, N5991, N5301, N2753);
buf BUF1 (N7915, N7906);
xor XOR2 (N7916, N7900, N6104);
nand NAND2 (N7917, N7910, N3470);
buf BUF1 (N7918, N7898);
buf BUF1 (N7919, N7918);
nor NOR2 (N7920, N7917, N1143);
or OR4 (N7921, N7914, N7681, N3177, N2643);
nand NAND3 (N7922, N7911, N2901, N6137);
buf BUF1 (N7923, N7915);
and AND2 (N7924, N7922, N1107);
nor NOR3 (N7925, N7919, N3860, N1468);
nor NOR2 (N7926, N7925, N5552);
nor NOR3 (N7927, N7916, N7088, N4741);
nor NOR2 (N7928, N7856, N6800);
not NOT1 (N7929, N7921);
xor XOR2 (N7930, N7924, N7411);
nand NAND4 (N7931, N7923, N7248, N5243, N4153);
and AND3 (N7932, N7927, N5811, N5865);
nand NAND3 (N7933, N7920, N1690, N6033);
or OR2 (N7934, N7913, N7421);
nand NAND4 (N7935, N7912, N7929, N4705, N3888);
nor NOR3 (N7936, N5643, N6823, N6857);
buf BUF1 (N7937, N7886);
not NOT1 (N7938, N7933);
nor NOR4 (N7939, N7928, N5414, N4065, N1313);
xor XOR2 (N7940, N7938, N5530);
nand NAND2 (N7941, N7932, N1101);
not NOT1 (N7942, N7939);
buf BUF1 (N7943, N7936);
not NOT1 (N7944, N7941);
buf BUF1 (N7945, N7937);
or OR2 (N7946, N7930, N4567);
or OR4 (N7947, N7945, N5850, N4657, N6564);
or OR2 (N7948, N7944, N5129);
or OR2 (N7949, N7934, N6951);
nor NOR3 (N7950, N7926, N2521, N4534);
and AND4 (N7951, N7931, N7300, N1980, N5719);
xor XOR2 (N7952, N7947, N4195);
and AND2 (N7953, N7952, N5792);
buf BUF1 (N7954, N7935);
nor NOR3 (N7955, N7954, N1671, N919);
not NOT1 (N7956, N7951);
and AND2 (N7957, N7956, N6731);
nand NAND2 (N7958, N7948, N663);
buf BUF1 (N7959, N7942);
or OR4 (N7960, N7958, N485, N813, N7193);
nand NAND2 (N7961, N7943, N6073);
buf BUF1 (N7962, N7953);
nor NOR3 (N7963, N7946, N3540, N5993);
nor NOR2 (N7964, N7961, N3538);
or OR2 (N7965, N7955, N6276);
xor XOR2 (N7966, N7962, N3984);
and AND3 (N7967, N7964, N1168, N3114);
or OR4 (N7968, N7963, N7443, N5708, N4014);
nor NOR3 (N7969, N7965, N6483, N3159);
and AND3 (N7970, N7966, N2166, N5865);
or OR2 (N7971, N7970, N3025);
and AND2 (N7972, N7971, N3720);
and AND4 (N7973, N7940, N4829, N2743, N2262);
nand NAND2 (N7974, N7968, N7721);
or OR2 (N7975, N7973, N7397);
xor XOR2 (N7976, N7957, N4261);
or OR2 (N7977, N7969, N561);
nor NOR3 (N7978, N7967, N894, N2897);
and AND4 (N7979, N7949, N5769, N205, N5256);
and AND2 (N7980, N7977, N4662);
nor NOR4 (N7981, N7975, N4688, N2057, N4856);
or OR4 (N7982, N7974, N1642, N1993, N2517);
nor NOR2 (N7983, N7959, N3746);
not NOT1 (N7984, N7976);
buf BUF1 (N7985, N7960);
nand NAND2 (N7986, N7950, N2839);
not NOT1 (N7987, N7984);
not NOT1 (N7988, N7986);
nor NOR3 (N7989, N7979, N3043, N1872);
not NOT1 (N7990, N7985);
or OR4 (N7991, N7982, N7618, N2638, N1533);
not NOT1 (N7992, N7990);
and AND4 (N7993, N7991, N7988, N3386, N4616);
buf BUF1 (N7994, N7084);
buf BUF1 (N7995, N7989);
or OR2 (N7996, N7980, N6968);
and AND2 (N7997, N7978, N7495);
and AND4 (N7998, N7972, N7622, N3312, N6728);
nand NAND4 (N7999, N7983, N4564, N1313, N5648);
nor NOR4 (N8000, N7993, N1412, N5965, N5942);
buf BUF1 (N8001, N8000);
buf BUF1 (N8002, N7997);
nor NOR4 (N8003, N7994, N6258, N2667, N1993);
nand NAND2 (N8004, N7981, N3457);
nor NOR4 (N8005, N8003, N7216, N2176, N5055);
nand NAND2 (N8006, N8001, N5732);
nor NOR4 (N8007, N8005, N2300, N3614, N7791);
nand NAND2 (N8008, N7998, N264);
nand NAND4 (N8009, N8006, N3035, N1573, N5677);
not NOT1 (N8010, N7999);
xor XOR2 (N8011, N8008, N7089);
and AND4 (N8012, N8009, N52, N1143, N6993);
and AND2 (N8013, N7992, N6439);
and AND4 (N8014, N8002, N5735, N7313, N6238);
nor NOR3 (N8015, N7987, N1737, N3302);
and AND3 (N8016, N8010, N5903, N6613);
nor NOR2 (N8017, N8016, N784);
buf BUF1 (N8018, N8007);
not NOT1 (N8019, N8015);
buf BUF1 (N8020, N8014);
and AND4 (N8021, N8018, N3877, N6619, N4544);
nor NOR2 (N8022, N8020, N2864);
not NOT1 (N8023, N7995);
not NOT1 (N8024, N8011);
xor XOR2 (N8025, N8021, N2004);
or OR4 (N8026, N8022, N3000, N634, N2105);
xor XOR2 (N8027, N8025, N6463);
nand NAND4 (N8028, N7996, N66, N6440, N6996);
and AND2 (N8029, N8027, N1526);
and AND4 (N8030, N8029, N5852, N2678, N1046);
or OR2 (N8031, N8019, N1391);
nand NAND3 (N8032, N8013, N1882, N7801);
nand NAND2 (N8033, N8030, N7405);
xor XOR2 (N8034, N8023, N5028);
nand NAND4 (N8035, N8031, N7375, N6015, N113);
not NOT1 (N8036, N8035);
buf BUF1 (N8037, N8033);
or OR3 (N8038, N8037, N5890, N6585);
buf BUF1 (N8039, N8028);
or OR3 (N8040, N8012, N3337, N6281);
or OR2 (N8041, N8038, N7530);
nor NOR4 (N8042, N8041, N3082, N1731, N221);
nor NOR2 (N8043, N8004, N2247);
nor NOR2 (N8044, N8039, N843);
xor XOR2 (N8045, N8044, N5951);
or OR2 (N8046, N8032, N691);
or OR4 (N8047, N8040, N5867, N7316, N2160);
not NOT1 (N8048, N8046);
nand NAND4 (N8049, N8042, N2071, N5913, N3873);
nor NOR3 (N8050, N8048, N6892, N1445);
or OR4 (N8051, N8050, N1520, N7215, N472);
buf BUF1 (N8052, N8049);
nand NAND3 (N8053, N8017, N7878, N5055);
and AND2 (N8054, N8047, N7314);
not NOT1 (N8055, N8034);
not NOT1 (N8056, N8045);
buf BUF1 (N8057, N8056);
not NOT1 (N8058, N8026);
nor NOR3 (N8059, N8055, N6583, N5238);
or OR3 (N8060, N8059, N802, N3469);
xor XOR2 (N8061, N8052, N354);
nor NOR2 (N8062, N8024, N593);
or OR4 (N8063, N8060, N2275, N1886, N7699);
buf BUF1 (N8064, N8054);
or OR2 (N8065, N8043, N6359);
and AND2 (N8066, N8063, N1466);
nand NAND3 (N8067, N8053, N7644, N2746);
and AND2 (N8068, N8036, N2547);
buf BUF1 (N8069, N8057);
and AND2 (N8070, N8058, N4865);
nor NOR4 (N8071, N8062, N2548, N2595, N2141);
nor NOR3 (N8072, N8066, N2287, N2611);
buf BUF1 (N8073, N8069);
or OR2 (N8074, N8070, N4237);
xor XOR2 (N8075, N8065, N8042);
and AND2 (N8076, N8068, N4232);
nor NOR4 (N8077, N8073, N4960, N4838, N5951);
or OR3 (N8078, N8067, N4031, N7984);
and AND4 (N8079, N8074, N1862, N545, N6115);
or OR4 (N8080, N8071, N1738, N6497, N8055);
nand NAND3 (N8081, N8051, N2915, N3045);
xor XOR2 (N8082, N8072, N5758);
buf BUF1 (N8083, N8079);
buf BUF1 (N8084, N8083);
xor XOR2 (N8085, N8061, N9);
nor NOR4 (N8086, N8064, N7948, N5201, N4568);
nand NAND2 (N8087, N8086, N5457);
buf BUF1 (N8088, N8084);
nand NAND2 (N8089, N8082, N2831);
xor XOR2 (N8090, N8089, N2949);
nand NAND3 (N8091, N8078, N4127, N1462);
nor NOR4 (N8092, N8080, N7857, N3097, N2654);
or OR4 (N8093, N8088, N197, N790, N2941);
and AND2 (N8094, N8090, N3266);
buf BUF1 (N8095, N8091);
xor XOR2 (N8096, N8077, N1557);
buf BUF1 (N8097, N8085);
or OR4 (N8098, N8095, N1837, N3724, N6981);
xor XOR2 (N8099, N8094, N7449);
nand NAND2 (N8100, N8097, N581);
or OR2 (N8101, N8087, N4304);
not NOT1 (N8102, N8092);
not NOT1 (N8103, N8075);
or OR2 (N8104, N8098, N1992);
and AND3 (N8105, N8100, N7612, N6221);
nand NAND4 (N8106, N8104, N7387, N2679, N5249);
nor NOR4 (N8107, N8099, N4404, N4330, N5060);
nand NAND2 (N8108, N8076, N5015);
nor NOR2 (N8109, N8093, N1163);
not NOT1 (N8110, N8109);
xor XOR2 (N8111, N8110, N409);
and AND4 (N8112, N8106, N6989, N2866, N7093);
nor NOR2 (N8113, N8081, N2328);
not NOT1 (N8114, N8096);
buf BUF1 (N8115, N8114);
xor XOR2 (N8116, N8107, N1832);
buf BUF1 (N8117, N8116);
or OR4 (N8118, N8102, N5898, N5169, N551);
not NOT1 (N8119, N8112);
nor NOR3 (N8120, N8118, N2759, N2646);
xor XOR2 (N8121, N8113, N6451);
buf BUF1 (N8122, N8121);
or OR3 (N8123, N8115, N5723, N1143);
nand NAND2 (N8124, N8111, N4968);
or OR4 (N8125, N8117, N5796, N2, N7363);
buf BUF1 (N8126, N8120);
buf BUF1 (N8127, N8101);
nand NAND3 (N8128, N8119, N1872, N7575);
or OR4 (N8129, N8103, N3622, N3754, N6135);
nand NAND3 (N8130, N8126, N5238, N1914);
xor XOR2 (N8131, N8122, N6918);
or OR3 (N8132, N8130, N5924, N6474);
nor NOR3 (N8133, N8131, N373, N1746);
not NOT1 (N8134, N8128);
xor XOR2 (N8135, N8133, N2849);
or OR3 (N8136, N8127, N3048, N5400);
xor XOR2 (N8137, N8136, N776);
nand NAND4 (N8138, N8132, N6592, N3965, N826);
xor XOR2 (N8139, N8137, N4969);
buf BUF1 (N8140, N8135);
buf BUF1 (N8141, N8138);
or OR2 (N8142, N8140, N7732);
and AND2 (N8143, N8129, N7891);
or OR4 (N8144, N8124, N3671, N7, N7587);
or OR3 (N8145, N8144, N6118, N6297);
not NOT1 (N8146, N8139);
buf BUF1 (N8147, N8146);
buf BUF1 (N8148, N8108);
and AND4 (N8149, N8105, N7870, N4890, N5220);
xor XOR2 (N8150, N8141, N3952);
xor XOR2 (N8151, N8125, N1371);
buf BUF1 (N8152, N8147);
xor XOR2 (N8153, N8148, N5909);
and AND3 (N8154, N8123, N6776, N7720);
nor NOR2 (N8155, N8152, N4863);
or OR3 (N8156, N8142, N1993, N385);
nand NAND4 (N8157, N8151, N3284, N5462, N6468);
or OR2 (N8158, N8154, N890);
or OR4 (N8159, N8155, N5726, N2349, N6176);
buf BUF1 (N8160, N8157);
or OR4 (N8161, N8134, N8095, N2861, N929);
or OR4 (N8162, N8149, N2651, N3459, N7934);
xor XOR2 (N8163, N8159, N2430);
nor NOR2 (N8164, N8143, N5413);
and AND3 (N8165, N8145, N6943, N6681);
or OR3 (N8166, N8161, N7225, N4373);
nor NOR2 (N8167, N8150, N1403);
nand NAND4 (N8168, N8156, N6063, N1609, N143);
or OR2 (N8169, N8166, N2443);
not NOT1 (N8170, N8160);
xor XOR2 (N8171, N8167, N403);
or OR3 (N8172, N8170, N3634, N2581);
or OR2 (N8173, N8169, N4784);
buf BUF1 (N8174, N8173);
and AND4 (N8175, N8174, N7889, N2299, N7173);
or OR3 (N8176, N8153, N6788, N3546);
nand NAND3 (N8177, N8172, N230, N4257);
nor NOR3 (N8178, N8164, N2455, N3142);
and AND3 (N8179, N8163, N3463, N6030);
nor NOR2 (N8180, N8165, N5983);
buf BUF1 (N8181, N8177);
and AND4 (N8182, N8171, N3815, N4118, N3592);
buf BUF1 (N8183, N8178);
xor XOR2 (N8184, N8158, N6634);
buf BUF1 (N8185, N8182);
and AND3 (N8186, N8176, N5955, N6221);
or OR3 (N8187, N8184, N5538, N7660);
nor NOR3 (N8188, N8180, N2430, N5622);
xor XOR2 (N8189, N8187, N4891);
and AND3 (N8190, N8168, N6279, N7389);
nor NOR2 (N8191, N8190, N6925);
not NOT1 (N8192, N8189);
nor NOR2 (N8193, N8192, N5259);
not NOT1 (N8194, N8183);
and AND2 (N8195, N8175, N4846);
nand NAND2 (N8196, N8195, N153);
xor XOR2 (N8197, N8186, N812);
or OR4 (N8198, N8179, N3495, N4650, N1318);
nand NAND2 (N8199, N8191, N6475);
and AND3 (N8200, N8197, N7143, N1318);
nor NOR4 (N8201, N8162, N7215, N718, N1591);
or OR4 (N8202, N8181, N4005, N3557, N5356);
xor XOR2 (N8203, N8199, N6817);
buf BUF1 (N8204, N8193);
buf BUF1 (N8205, N8185);
buf BUF1 (N8206, N8200);
nand NAND3 (N8207, N8203, N7836, N6408);
or OR2 (N8208, N8198, N6105);
nor NOR4 (N8209, N8207, N5749, N7533, N5513);
xor XOR2 (N8210, N8196, N1970);
not NOT1 (N8211, N8205);
buf BUF1 (N8212, N8204);
nand NAND4 (N8213, N8202, N4173, N7164, N7913);
not NOT1 (N8214, N8188);
nand NAND3 (N8215, N8210, N7827, N5878);
xor XOR2 (N8216, N8209, N2037);
nor NOR3 (N8217, N8206, N7866, N2891);
buf BUF1 (N8218, N8212);
buf BUF1 (N8219, N8211);
buf BUF1 (N8220, N8213);
nand NAND2 (N8221, N8216, N1392);
nand NAND4 (N8222, N8194, N7292, N7085, N2226);
xor XOR2 (N8223, N8222, N2109);
nor NOR3 (N8224, N8214, N1648, N4648);
buf BUF1 (N8225, N8219);
not NOT1 (N8226, N8201);
buf BUF1 (N8227, N8217);
or OR2 (N8228, N8223, N4258);
or OR3 (N8229, N8208, N4377, N4513);
buf BUF1 (N8230, N8228);
not NOT1 (N8231, N8227);
nor NOR2 (N8232, N8231, N5434);
not NOT1 (N8233, N8230);
or OR4 (N8234, N8224, N3712, N3658, N3623);
buf BUF1 (N8235, N8233);
nand NAND3 (N8236, N8226, N6362, N3286);
nand NAND2 (N8237, N8232, N1454);
not NOT1 (N8238, N8225);
buf BUF1 (N8239, N8215);
nor NOR3 (N8240, N8220, N6344, N6206);
not NOT1 (N8241, N8238);
xor XOR2 (N8242, N8237, N7966);
nor NOR4 (N8243, N8241, N3382, N3247, N6355);
xor XOR2 (N8244, N8229, N3248);
nor NOR2 (N8245, N8234, N7577);
nand NAND3 (N8246, N8243, N677, N1854);
nand NAND4 (N8247, N8236, N7936, N937, N66);
nand NAND2 (N8248, N8221, N7491);
buf BUF1 (N8249, N8248);
nor NOR4 (N8250, N8239, N169, N4797, N2124);
buf BUF1 (N8251, N8235);
or OR4 (N8252, N8247, N2528, N8155, N5658);
buf BUF1 (N8253, N8246);
nor NOR2 (N8254, N8240, N3613);
or OR4 (N8255, N8218, N3138, N6407, N8187);
not NOT1 (N8256, N8254);
xor XOR2 (N8257, N8251, N440);
buf BUF1 (N8258, N8252);
nor NOR4 (N8259, N8255, N2963, N6990, N915);
nor NOR4 (N8260, N8253, N6266, N5499, N6033);
xor XOR2 (N8261, N8256, N257);
nor NOR3 (N8262, N8245, N430, N2845);
nor NOR3 (N8263, N8242, N4976, N1220);
xor XOR2 (N8264, N8244, N5609);
nand NAND2 (N8265, N8264, N1982);
xor XOR2 (N8266, N8249, N5708);
xor XOR2 (N8267, N8261, N7195);
not NOT1 (N8268, N8260);
buf BUF1 (N8269, N8265);
xor XOR2 (N8270, N8258, N6205);
or OR2 (N8271, N8269, N897);
nor NOR3 (N8272, N8270, N2647, N1290);
buf BUF1 (N8273, N8259);
not NOT1 (N8274, N8267);
not NOT1 (N8275, N8263);
buf BUF1 (N8276, N8262);
buf BUF1 (N8277, N8272);
buf BUF1 (N8278, N8268);
not NOT1 (N8279, N8276);
not NOT1 (N8280, N8278);
nand NAND4 (N8281, N8274, N7399, N4578, N2774);
not NOT1 (N8282, N8277);
not NOT1 (N8283, N8280);
or OR2 (N8284, N8271, N2955);
buf BUF1 (N8285, N8250);
or OR3 (N8286, N8279, N6957, N4120);
or OR2 (N8287, N8282, N2433);
or OR3 (N8288, N8287, N6399, N3192);
or OR3 (N8289, N8285, N5082, N332);
not NOT1 (N8290, N8284);
xor XOR2 (N8291, N8290, N3897);
nand NAND3 (N8292, N8266, N3523, N6733);
nand NAND3 (N8293, N8257, N6195, N796);
buf BUF1 (N8294, N8289);
or OR4 (N8295, N8293, N5944, N7681, N4625);
not NOT1 (N8296, N8288);
not NOT1 (N8297, N8275);
nor NOR2 (N8298, N8283, N745);
xor XOR2 (N8299, N8286, N7819);
xor XOR2 (N8300, N8298, N1020);
xor XOR2 (N8301, N8291, N6864);
or OR4 (N8302, N8273, N5438, N2834, N2794);
buf BUF1 (N8303, N8281);
nor NOR4 (N8304, N8296, N5680, N5644, N4978);
or OR2 (N8305, N8299, N7788);
and AND4 (N8306, N8292, N7877, N6878, N412);
not NOT1 (N8307, N8295);
xor XOR2 (N8308, N8306, N1629);
buf BUF1 (N8309, N8294);
nor NOR2 (N8310, N8300, N7188);
xor XOR2 (N8311, N8305, N2710);
or OR2 (N8312, N8304, N4085);
not NOT1 (N8313, N8307);
buf BUF1 (N8314, N8309);
buf BUF1 (N8315, N8301);
and AND4 (N8316, N8297, N4193, N4552, N3698);
not NOT1 (N8317, N8308);
not NOT1 (N8318, N8317);
or OR2 (N8319, N8314, N7258);
or OR4 (N8320, N8313, N7118, N3645, N2658);
buf BUF1 (N8321, N8310);
and AND2 (N8322, N8315, N3864);
xor XOR2 (N8323, N8302, N5876);
and AND3 (N8324, N8322, N3257, N4651);
nor NOR3 (N8325, N8324, N7415, N6848);
and AND4 (N8326, N8321, N2955, N1022, N7197);
buf BUF1 (N8327, N8316);
xor XOR2 (N8328, N8311, N5183);
buf BUF1 (N8329, N8323);
nor NOR3 (N8330, N8320, N6157, N8165);
or OR3 (N8331, N8330, N5302, N925);
or OR2 (N8332, N8328, N571);
nand NAND2 (N8333, N8303, N1524);
or OR3 (N8334, N8325, N1003, N4134);
nand NAND2 (N8335, N8318, N7151);
or OR2 (N8336, N8329, N1744);
not NOT1 (N8337, N8334);
nand NAND4 (N8338, N8333, N6901, N5990, N2118);
buf BUF1 (N8339, N8336);
nor NOR3 (N8340, N8327, N5438, N6826);
xor XOR2 (N8341, N8338, N132);
not NOT1 (N8342, N8340);
and AND3 (N8343, N8331, N7770, N503);
not NOT1 (N8344, N8326);
nor NOR3 (N8345, N8343, N2515, N1370);
or OR2 (N8346, N8319, N4850);
not NOT1 (N8347, N8335);
nor NOR3 (N8348, N8312, N6196, N5600);
or OR3 (N8349, N8332, N11, N7408);
xor XOR2 (N8350, N8347, N562);
nor NOR3 (N8351, N8341, N395, N2243);
xor XOR2 (N8352, N8339, N2495);
buf BUF1 (N8353, N8337);
nor NOR3 (N8354, N8351, N3305, N2598);
and AND3 (N8355, N8353, N2596, N6090);
xor XOR2 (N8356, N8342, N4052);
nand NAND4 (N8357, N8345, N8044, N7975, N7612);
nand NAND4 (N8358, N8354, N2474, N6749, N2172);
and AND2 (N8359, N8352, N4939);
and AND4 (N8360, N8346, N7185, N5508, N7486);
and AND4 (N8361, N8358, N6784, N6071, N202);
not NOT1 (N8362, N8349);
or OR4 (N8363, N8356, N1216, N3143, N4057);
xor XOR2 (N8364, N8363, N841);
buf BUF1 (N8365, N8362);
nand NAND3 (N8366, N8365, N5100, N3026);
and AND4 (N8367, N8359, N7533, N5655, N4566);
xor XOR2 (N8368, N8344, N7078);
not NOT1 (N8369, N8350);
and AND3 (N8370, N8355, N23, N7335);
nor NOR4 (N8371, N8366, N6737, N4285, N2289);
buf BUF1 (N8372, N8348);
nand NAND3 (N8373, N8367, N6826, N4015);
nand NAND3 (N8374, N8360, N884, N3506);
buf BUF1 (N8375, N8368);
xor XOR2 (N8376, N8369, N6675);
or OR2 (N8377, N8357, N7112);
nand NAND2 (N8378, N8371, N6188);
and AND3 (N8379, N8370, N5358, N4697);
buf BUF1 (N8380, N8372);
buf BUF1 (N8381, N8373);
nor NOR2 (N8382, N8380, N7207);
or OR3 (N8383, N8374, N7578, N7987);
nand NAND4 (N8384, N8379, N2311, N1351, N7410);
buf BUF1 (N8385, N8376);
xor XOR2 (N8386, N8377, N7089);
nor NOR3 (N8387, N8361, N5711, N8248);
nor NOR3 (N8388, N8386, N5386, N5825);
nor NOR2 (N8389, N8364, N5209);
nand NAND3 (N8390, N8381, N7514, N6566);
and AND2 (N8391, N8388, N1665);
and AND4 (N8392, N8391, N7277, N6612, N3384);
xor XOR2 (N8393, N8384, N5294);
buf BUF1 (N8394, N8389);
or OR2 (N8395, N8375, N6917);
not NOT1 (N8396, N8390);
nand NAND4 (N8397, N8382, N3465, N175, N6303);
or OR4 (N8398, N8383, N5427, N656, N7582);
or OR3 (N8399, N8393, N3252, N1087);
and AND3 (N8400, N8385, N1104, N4389);
and AND4 (N8401, N8392, N7600, N4637, N7989);
xor XOR2 (N8402, N8378, N4599);
and AND3 (N8403, N8399, N2675, N5009);
not NOT1 (N8404, N8398);
or OR3 (N8405, N8403, N4640, N4136);
and AND4 (N8406, N8397, N3279, N2593, N1430);
and AND2 (N8407, N8405, N8279);
or OR3 (N8408, N8402, N6341, N2186);
or OR4 (N8409, N8407, N26, N1372, N4263);
buf BUF1 (N8410, N8396);
not NOT1 (N8411, N8406);
xor XOR2 (N8412, N8401, N4888);
and AND2 (N8413, N8411, N1290);
and AND3 (N8414, N8404, N1249, N5144);
nor NOR3 (N8415, N8413, N6080, N5759);
nor NOR2 (N8416, N8395, N8035);
or OR3 (N8417, N8400, N6718, N3108);
buf BUF1 (N8418, N8394);
or OR3 (N8419, N8412, N6149, N5231);
nand NAND4 (N8420, N8410, N5061, N4131, N3410);
and AND3 (N8421, N8419, N1268, N3803);
buf BUF1 (N8422, N8416);
nor NOR3 (N8423, N8414, N853, N2756);
or OR3 (N8424, N8387, N3672, N7149);
xor XOR2 (N8425, N8421, N1885);
or OR3 (N8426, N8418, N6537, N7989);
xor XOR2 (N8427, N8422, N4525);
nor NOR2 (N8428, N8427, N7369);
not NOT1 (N8429, N8415);
xor XOR2 (N8430, N8417, N3516);
not NOT1 (N8431, N8425);
buf BUF1 (N8432, N8430);
nor NOR3 (N8433, N8431, N2710, N6167);
and AND3 (N8434, N8409, N1206, N6835);
nand NAND3 (N8435, N8428, N6024, N4239);
nand NAND2 (N8436, N8434, N1971);
nor NOR3 (N8437, N8424, N8420, N378);
nor NOR2 (N8438, N3972, N1447);
not NOT1 (N8439, N8437);
xor XOR2 (N8440, N8423, N6014);
nand NAND2 (N8441, N8432, N1559);
not NOT1 (N8442, N8439);
xor XOR2 (N8443, N8442, N6706);
nor NOR3 (N8444, N8433, N1495, N5254);
or OR2 (N8445, N8426, N2811);
and AND4 (N8446, N8429, N6038, N4947, N2406);
or OR3 (N8447, N8446, N1394, N8043);
buf BUF1 (N8448, N8441);
nor NOR4 (N8449, N8440, N4978, N4641, N7518);
nor NOR2 (N8450, N8443, N2352);
not NOT1 (N8451, N8445);
nor NOR2 (N8452, N8450, N3759);
xor XOR2 (N8453, N8435, N2915);
and AND2 (N8454, N8452, N6631);
or OR2 (N8455, N8408, N4865);
nor NOR3 (N8456, N8454, N7376, N3990);
xor XOR2 (N8457, N8447, N3604);
nand NAND3 (N8458, N8451, N5207, N2568);
or OR4 (N8459, N8436, N1927, N3040, N7120);
nor NOR2 (N8460, N8457, N249);
nor NOR4 (N8461, N8453, N89, N2262, N2358);
or OR4 (N8462, N8460, N3748, N4655, N6136);
and AND4 (N8463, N8461, N7981, N3572, N2627);
xor XOR2 (N8464, N8462, N435);
nor NOR2 (N8465, N8455, N5769);
buf BUF1 (N8466, N8448);
nor NOR4 (N8467, N8466, N2433, N8433, N918);
nand NAND2 (N8468, N8459, N4587);
and AND2 (N8469, N8438, N2465);
nor NOR2 (N8470, N8465, N7274);
nor NOR4 (N8471, N8464, N2663, N4000, N1946);
nand NAND2 (N8472, N8471, N3019);
buf BUF1 (N8473, N8456);
nand NAND2 (N8474, N8468, N8357);
not NOT1 (N8475, N8449);
not NOT1 (N8476, N8470);
nor NOR3 (N8477, N8472, N7651, N3668);
not NOT1 (N8478, N8458);
xor XOR2 (N8479, N8469, N1676);
not NOT1 (N8480, N8444);
not NOT1 (N8481, N8477);
xor XOR2 (N8482, N8475, N7335);
buf BUF1 (N8483, N8478);
and AND3 (N8484, N8483, N7338, N4677);
buf BUF1 (N8485, N8481);
nand NAND2 (N8486, N8463, N4746);
xor XOR2 (N8487, N8480, N2853);
and AND2 (N8488, N8482, N3353);
xor XOR2 (N8489, N8484, N8394);
nand NAND2 (N8490, N8485, N8076);
xor XOR2 (N8491, N8486, N3446);
nor NOR2 (N8492, N8489, N7109);
xor XOR2 (N8493, N8479, N1972);
and AND4 (N8494, N8487, N323, N3281, N5970);
or OR4 (N8495, N8474, N6491, N3386, N6422);
not NOT1 (N8496, N8492);
xor XOR2 (N8497, N8495, N7818);
not NOT1 (N8498, N8476);
nand NAND2 (N8499, N8493, N4145);
buf BUF1 (N8500, N8494);
xor XOR2 (N8501, N8497, N2933);
or OR3 (N8502, N8501, N3518, N4512);
buf BUF1 (N8503, N8496);
xor XOR2 (N8504, N8473, N8376);
and AND4 (N8505, N8499, N4368, N759, N5234);
nand NAND2 (N8506, N8504, N6396);
xor XOR2 (N8507, N8503, N2682);
nand NAND3 (N8508, N8488, N3765, N3981);
buf BUF1 (N8509, N8502);
nand NAND2 (N8510, N8490, N4733);
nand NAND4 (N8511, N8508, N6676, N5364, N6991);
and AND4 (N8512, N8491, N140, N2351, N5968);
buf BUF1 (N8513, N8500);
not NOT1 (N8514, N8513);
and AND3 (N8515, N8509, N8259, N790);
and AND4 (N8516, N8510, N516, N415, N2367);
nand NAND4 (N8517, N8511, N547, N2622, N1162);
nor NOR4 (N8518, N8506, N4810, N4215, N1470);
nor NOR3 (N8519, N8512, N6970, N6719);
and AND3 (N8520, N8516, N4632, N5278);
nor NOR4 (N8521, N8505, N4901, N6018, N1185);
buf BUF1 (N8522, N8498);
and AND3 (N8523, N8515, N8002, N7533);
not NOT1 (N8524, N8518);
nand NAND4 (N8525, N8517, N5132, N4653, N4925);
or OR3 (N8526, N8514, N741, N5170);
nand NAND2 (N8527, N8523, N6379);
buf BUF1 (N8528, N8526);
not NOT1 (N8529, N8525);
and AND4 (N8530, N8467, N1984, N2805, N1590);
not NOT1 (N8531, N8519);
nand NAND4 (N8532, N8527, N3449, N5225, N6751);
not NOT1 (N8533, N8524);
not NOT1 (N8534, N8529);
nor NOR2 (N8535, N8534, N2173);
buf BUF1 (N8536, N8533);
and AND3 (N8537, N8522, N4089, N49);
nor NOR4 (N8538, N8521, N7670, N3464, N4161);
not NOT1 (N8539, N8532);
or OR3 (N8540, N8507, N3950, N1913);
buf BUF1 (N8541, N8539);
nor NOR4 (N8542, N8541, N5273, N5417, N6180);
not NOT1 (N8543, N8520);
and AND2 (N8544, N8543, N1741);
xor XOR2 (N8545, N8531, N3953);
not NOT1 (N8546, N8535);
and AND4 (N8547, N8546, N7031, N1914, N5189);
or OR2 (N8548, N8536, N7721);
nand NAND2 (N8549, N8547, N3904);
and AND3 (N8550, N8538, N1913, N3721);
xor XOR2 (N8551, N8530, N7299);
and AND2 (N8552, N8548, N7641);
xor XOR2 (N8553, N8551, N17);
nand NAND4 (N8554, N8549, N791, N2938, N2303);
not NOT1 (N8555, N8542);
nor NOR3 (N8556, N8528, N729, N730);
xor XOR2 (N8557, N8544, N248);
not NOT1 (N8558, N8554);
xor XOR2 (N8559, N8555, N1847);
and AND2 (N8560, N8537, N3997);
not NOT1 (N8561, N8552);
nor NOR4 (N8562, N8553, N5049, N5976, N7417);
xor XOR2 (N8563, N8560, N528);
nand NAND3 (N8564, N8561, N2676, N6382);
nand NAND2 (N8565, N8564, N3796);
nor NOR3 (N8566, N8559, N6877, N6651);
nor NOR4 (N8567, N8550, N2307, N8303, N3960);
and AND3 (N8568, N8556, N760, N1377);
and AND4 (N8569, N8566, N4207, N1225, N7499);
not NOT1 (N8570, N8567);
buf BUF1 (N8571, N8558);
not NOT1 (N8572, N8571);
nor NOR3 (N8573, N8568, N4161, N6417);
buf BUF1 (N8574, N8545);
or OR4 (N8575, N8557, N801, N4377, N1319);
or OR3 (N8576, N8562, N5276, N3812);
buf BUF1 (N8577, N8570);
buf BUF1 (N8578, N8540);
and AND2 (N8579, N8573, N3028);
not NOT1 (N8580, N8578);
nor NOR4 (N8581, N8565, N428, N3771, N5228);
nor NOR2 (N8582, N8580, N232);
not NOT1 (N8583, N8581);
xor XOR2 (N8584, N8572, N5122);
or OR3 (N8585, N8569, N3143, N474);
xor XOR2 (N8586, N8583, N6851);
xor XOR2 (N8587, N8584, N7887);
not NOT1 (N8588, N8574);
buf BUF1 (N8589, N8575);
or OR2 (N8590, N8589, N319);
buf BUF1 (N8591, N8588);
xor XOR2 (N8592, N8576, N1837);
or OR3 (N8593, N8579, N7628, N6688);
buf BUF1 (N8594, N8587);
and AND3 (N8595, N8577, N3295, N256);
not NOT1 (N8596, N8594);
xor XOR2 (N8597, N8593, N3347);
or OR3 (N8598, N8590, N6608, N3521);
not NOT1 (N8599, N8595);
and AND3 (N8600, N8591, N5083, N4516);
buf BUF1 (N8601, N8598);
xor XOR2 (N8602, N8596, N4561);
nand NAND2 (N8603, N8601, N5552);
xor XOR2 (N8604, N8600, N6564);
and AND4 (N8605, N8604, N3384, N4216, N6255);
and AND3 (N8606, N8592, N6892, N5845);
and AND3 (N8607, N8582, N4825, N2193);
xor XOR2 (N8608, N8605, N7244);
nand NAND2 (N8609, N8586, N3027);
not NOT1 (N8610, N8599);
xor XOR2 (N8611, N8606, N4489);
and AND3 (N8612, N8611, N2149, N8283);
nand NAND4 (N8613, N8612, N6759, N3905, N4332);
not NOT1 (N8614, N8602);
xor XOR2 (N8615, N8607, N3247);
nor NOR3 (N8616, N8603, N2825, N4318);
and AND4 (N8617, N8608, N7969, N7664, N2998);
nor NOR2 (N8618, N8616, N4530);
or OR3 (N8619, N8609, N2536, N4522);
or OR2 (N8620, N8615, N6720);
nand NAND2 (N8621, N8613, N1964);
and AND2 (N8622, N8614, N6144);
and AND3 (N8623, N8621, N5208, N4360);
nand NAND2 (N8624, N8622, N1783);
xor XOR2 (N8625, N8585, N1394);
not NOT1 (N8626, N8617);
not NOT1 (N8627, N8619);
not NOT1 (N8628, N8627);
and AND4 (N8629, N8618, N6749, N4900, N2439);
or OR2 (N8630, N8597, N1624);
or OR3 (N8631, N8628, N1680, N8489);
not NOT1 (N8632, N8630);
xor XOR2 (N8633, N8620, N6368);
nor NOR4 (N8634, N8610, N5908, N5565, N2535);
nor NOR2 (N8635, N8625, N8223);
xor XOR2 (N8636, N8634, N2396);
and AND2 (N8637, N8563, N2928);
and AND3 (N8638, N8632, N4812, N3462);
xor XOR2 (N8639, N8629, N5297);
or OR2 (N8640, N8638, N3644);
or OR4 (N8641, N8626, N855, N2955, N3035);
xor XOR2 (N8642, N8636, N1643);
xor XOR2 (N8643, N8639, N4647);
nor NOR3 (N8644, N8633, N3006, N3454);
buf BUF1 (N8645, N8637);
nor NOR2 (N8646, N8623, N1099);
nor NOR3 (N8647, N8640, N8056, N3793);
not NOT1 (N8648, N8644);
buf BUF1 (N8649, N8641);
and AND2 (N8650, N8631, N2997);
and AND2 (N8651, N8650, N2761);
xor XOR2 (N8652, N8645, N5108);
and AND2 (N8653, N8624, N6973);
buf BUF1 (N8654, N8647);
nor NOR4 (N8655, N8654, N5090, N3804, N6751);
buf BUF1 (N8656, N8655);
xor XOR2 (N8657, N8635, N3427);
not NOT1 (N8658, N8642);
buf BUF1 (N8659, N8658);
buf BUF1 (N8660, N8659);
or OR2 (N8661, N8652, N7494);
or OR3 (N8662, N8649, N7767, N8138);
and AND2 (N8663, N8661, N8531);
and AND3 (N8664, N8657, N1012, N6105);
or OR4 (N8665, N8648, N4408, N6575, N7230);
buf BUF1 (N8666, N8643);
nand NAND4 (N8667, N8664, N1750, N7617, N3701);
nand NAND4 (N8668, N8667, N5506, N6040, N4888);
nor NOR2 (N8669, N8662, N5433);
and AND3 (N8670, N8651, N2847, N5725);
and AND4 (N8671, N8660, N133, N7519, N6498);
nand NAND2 (N8672, N8663, N5799);
buf BUF1 (N8673, N8646);
nor NOR4 (N8674, N8672, N8526, N3824, N4121);
buf BUF1 (N8675, N8653);
nor NOR3 (N8676, N8666, N5954, N3429);
buf BUF1 (N8677, N8665);
or OR4 (N8678, N8675, N223, N2715, N8104);
nand NAND4 (N8679, N8670, N4806, N2695, N4864);
nand NAND2 (N8680, N8678, N7713);
not NOT1 (N8681, N8680);
nor NOR4 (N8682, N8674, N5565, N738, N4539);
nor NOR4 (N8683, N8668, N4554, N2841, N2930);
nand NAND4 (N8684, N8673, N3282, N3494, N2951);
xor XOR2 (N8685, N8677, N2287);
buf BUF1 (N8686, N8683);
buf BUF1 (N8687, N8682);
xor XOR2 (N8688, N8679, N60);
or OR2 (N8689, N8687, N3647);
and AND3 (N8690, N8671, N7546, N4540);
or OR3 (N8691, N8676, N2541, N3163);
xor XOR2 (N8692, N8684, N6136);
xor XOR2 (N8693, N8688, N4901);
and AND3 (N8694, N8691, N2868, N99);
and AND2 (N8695, N8686, N5819);
nor NOR4 (N8696, N8689, N962, N333, N2047);
or OR2 (N8697, N8656, N7058);
and AND3 (N8698, N8685, N3626, N6880);
nand NAND4 (N8699, N8697, N4688, N6526, N591);
nor NOR2 (N8700, N8695, N6406);
nand NAND3 (N8701, N8669, N7292, N7838);
buf BUF1 (N8702, N8681);
and AND4 (N8703, N8699, N1472, N5443, N1916);
xor XOR2 (N8704, N8700, N7420);
and AND3 (N8705, N8704, N3313, N2113);
not NOT1 (N8706, N8702);
not NOT1 (N8707, N8694);
nand NAND3 (N8708, N8705, N3561, N882);
xor XOR2 (N8709, N8692, N2920);
and AND4 (N8710, N8709, N3004, N4632, N590);
nor NOR2 (N8711, N8693, N8014);
nand NAND3 (N8712, N8710, N1310, N224);
or OR2 (N8713, N8698, N2298);
nand NAND3 (N8714, N8701, N1629, N8426);
xor XOR2 (N8715, N8712, N4439);
and AND4 (N8716, N8707, N844, N5021, N5032);
nor NOR4 (N8717, N8708, N1934, N1159, N6582);
and AND3 (N8718, N8711, N1986, N1234);
or OR3 (N8719, N8718, N4015, N7574);
nand NAND2 (N8720, N8696, N3857);
nor NOR4 (N8721, N8690, N1779, N2483, N3300);
not NOT1 (N8722, N8721);
or OR3 (N8723, N8714, N3745, N3612);
xor XOR2 (N8724, N8723, N4165);
nand NAND3 (N8725, N8715, N2486, N326);
nand NAND2 (N8726, N8722, N5221);
buf BUF1 (N8727, N8716);
xor XOR2 (N8728, N8724, N2124);
not NOT1 (N8729, N8713);
xor XOR2 (N8730, N8728, N5714);
nand NAND4 (N8731, N8725, N1245, N1900, N787);
and AND2 (N8732, N8729, N5960);
not NOT1 (N8733, N8706);
or OR2 (N8734, N8720, N1350);
nor NOR4 (N8735, N8732, N8223, N5505, N3664);
or OR2 (N8736, N8727, N3047);
buf BUF1 (N8737, N8703);
xor XOR2 (N8738, N8726, N4202);
nand NAND4 (N8739, N8737, N1945, N649, N4263);
not NOT1 (N8740, N8719);
or OR4 (N8741, N8738, N852, N5878, N2530);
nor NOR2 (N8742, N8740, N4338);
and AND2 (N8743, N8733, N8069);
not NOT1 (N8744, N8741);
or OR4 (N8745, N8744, N408, N7753, N4750);
nor NOR3 (N8746, N8739, N1273, N4179);
nand NAND3 (N8747, N8742, N5921, N8722);
and AND2 (N8748, N8734, N35);
and AND4 (N8749, N8748, N2343, N2679, N6469);
or OR2 (N8750, N8743, N1803);
xor XOR2 (N8751, N8731, N1873);
and AND4 (N8752, N8749, N8281, N4562, N4587);
nand NAND2 (N8753, N8736, N6504);
or OR3 (N8754, N8752, N8543, N3649);
and AND4 (N8755, N8754, N3152, N5267, N2633);
nor NOR2 (N8756, N8746, N666);
nand NAND4 (N8757, N8753, N3032, N3829, N6846);
nand NAND4 (N8758, N8730, N2581, N8493, N7651);
nand NAND3 (N8759, N8735, N3278, N1672);
xor XOR2 (N8760, N8759, N149);
and AND3 (N8761, N8751, N6719, N2756);
and AND2 (N8762, N8755, N2764);
nand NAND3 (N8763, N8747, N3342, N6709);
nor NOR2 (N8764, N8762, N3470);
not NOT1 (N8765, N8760);
and AND3 (N8766, N8750, N743, N3447);
and AND3 (N8767, N8766, N6532, N994);
buf BUF1 (N8768, N8745);
nor NOR4 (N8769, N8758, N2977, N6143, N2876);
nand NAND2 (N8770, N8756, N5472);
xor XOR2 (N8771, N8765, N3794);
not NOT1 (N8772, N8764);
nor NOR2 (N8773, N8771, N5907);
nor NOR2 (N8774, N8763, N7679);
buf BUF1 (N8775, N8772);
not NOT1 (N8776, N8775);
nor NOR3 (N8777, N8717, N6642, N54);
and AND2 (N8778, N8769, N5084);
and AND2 (N8779, N8761, N3759);
not NOT1 (N8780, N8774);
nand NAND3 (N8781, N8779, N6559, N5223);
nor NOR4 (N8782, N8773, N1929, N7571, N7080);
nor NOR2 (N8783, N8777, N5103);
not NOT1 (N8784, N8768);
buf BUF1 (N8785, N8757);
nor NOR2 (N8786, N8785, N1921);
nand NAND4 (N8787, N8784, N3612, N8195, N5935);
nor NOR2 (N8788, N8783, N6086);
nor NOR2 (N8789, N8770, N1357);
xor XOR2 (N8790, N8788, N5467);
nor NOR4 (N8791, N8787, N2256, N696, N3421);
nor NOR2 (N8792, N8767, N647);
nand NAND2 (N8793, N8778, N3761);
not NOT1 (N8794, N8776);
nor NOR3 (N8795, N8786, N1212, N1414);
not NOT1 (N8796, N8793);
buf BUF1 (N8797, N8794);
buf BUF1 (N8798, N8792);
and AND2 (N8799, N8791, N3680);
not NOT1 (N8800, N8797);
xor XOR2 (N8801, N8795, N1860);
or OR3 (N8802, N8782, N1987, N8169);
nand NAND3 (N8803, N8789, N5603, N6927);
nor NOR2 (N8804, N8799, N2048);
or OR4 (N8805, N8800, N4066, N249, N4871);
nand NAND2 (N8806, N8796, N7414);
and AND4 (N8807, N8803, N1043, N1709, N6994);
xor XOR2 (N8808, N8798, N4123);
and AND2 (N8809, N8802, N3857);
and AND3 (N8810, N8806, N5732, N7162);
and AND2 (N8811, N8805, N4461);
nand NAND3 (N8812, N8807, N6093, N6586);
xor XOR2 (N8813, N8812, N2408);
not NOT1 (N8814, N8808);
nand NAND4 (N8815, N8809, N7429, N7136, N4850);
not NOT1 (N8816, N8814);
and AND4 (N8817, N8813, N6668, N4774, N195);
buf BUF1 (N8818, N8815);
xor XOR2 (N8819, N8811, N7069);
nor NOR4 (N8820, N8780, N8713, N8103, N5861);
not NOT1 (N8821, N8810);
nor NOR3 (N8822, N8820, N6751, N2510);
and AND3 (N8823, N8804, N1711, N4421);
nor NOR3 (N8824, N8823, N2862, N5395);
not NOT1 (N8825, N8822);
nand NAND3 (N8826, N8816, N2087, N3163);
not NOT1 (N8827, N8818);
or OR2 (N8828, N8819, N8778);
not NOT1 (N8829, N8790);
buf BUF1 (N8830, N8827);
nor NOR2 (N8831, N8781, N1383);
xor XOR2 (N8832, N8817, N6652);
xor XOR2 (N8833, N8824, N8539);
xor XOR2 (N8834, N8831, N1129);
or OR2 (N8835, N8830, N2549);
not NOT1 (N8836, N8834);
and AND3 (N8837, N8832, N836, N5518);
and AND4 (N8838, N8829, N5975, N2169, N8220);
nand NAND2 (N8839, N8825, N7095);
nand NAND2 (N8840, N8837, N2571);
or OR4 (N8841, N8828, N5397, N2096, N4430);
or OR4 (N8842, N8840, N2576, N6853, N1265);
not NOT1 (N8843, N8842);
nand NAND4 (N8844, N8826, N1766, N7060, N8723);
or OR2 (N8845, N8821, N7608);
xor XOR2 (N8846, N8838, N1385);
buf BUF1 (N8847, N8835);
xor XOR2 (N8848, N8847, N4495);
and AND4 (N8849, N8801, N4654, N1622, N7353);
buf BUF1 (N8850, N8844);
nand NAND2 (N8851, N8839, N4145);
and AND4 (N8852, N8845, N2173, N330, N1038);
or OR4 (N8853, N8843, N4793, N1599, N993);
buf BUF1 (N8854, N8846);
and AND2 (N8855, N8854, N1519);
nor NOR3 (N8856, N8849, N723, N8618);
nor NOR4 (N8857, N8852, N2850, N2330, N2863);
not NOT1 (N8858, N8833);
buf BUF1 (N8859, N8855);
not NOT1 (N8860, N8851);
xor XOR2 (N8861, N8841, N5096);
not NOT1 (N8862, N8836);
and AND2 (N8863, N8862, N8792);
or OR3 (N8864, N8858, N8695, N7154);
or OR2 (N8865, N8859, N7209);
xor XOR2 (N8866, N8861, N3124);
xor XOR2 (N8867, N8863, N4938);
or OR3 (N8868, N8856, N3258, N5912);
nand NAND3 (N8869, N8857, N8812, N6517);
buf BUF1 (N8870, N8850);
and AND2 (N8871, N8864, N8651);
or OR4 (N8872, N8867, N8470, N8352, N198);
or OR3 (N8873, N8848, N1169, N167);
nand NAND4 (N8874, N8873, N3765, N3167, N2119);
nand NAND2 (N8875, N8868, N3625);
not NOT1 (N8876, N8865);
xor XOR2 (N8877, N8875, N3977);
nand NAND3 (N8878, N8870, N678, N8382);
or OR3 (N8879, N8878, N7480, N291);
not NOT1 (N8880, N8874);
nor NOR4 (N8881, N8879, N8386, N2375, N8554);
buf BUF1 (N8882, N8876);
nor NOR3 (N8883, N8871, N7122, N2408);
and AND2 (N8884, N8860, N2088);
nand NAND3 (N8885, N8877, N4709, N8572);
and AND2 (N8886, N8866, N3228);
nand NAND4 (N8887, N8853, N3707, N6620, N2845);
buf BUF1 (N8888, N8887);
not NOT1 (N8889, N8884);
nand NAND3 (N8890, N8889, N8848, N6569);
nand NAND2 (N8891, N8880, N7801);
xor XOR2 (N8892, N8883, N1225);
and AND3 (N8893, N8869, N156, N3471);
not NOT1 (N8894, N8882);
buf BUF1 (N8895, N8888);
not NOT1 (N8896, N8892);
xor XOR2 (N8897, N8894, N1706);
not NOT1 (N8898, N8881);
buf BUF1 (N8899, N8886);
xor XOR2 (N8900, N8899, N6522);
and AND4 (N8901, N8895, N951, N4334, N1844);
not NOT1 (N8902, N8893);
buf BUF1 (N8903, N8898);
buf BUF1 (N8904, N8890);
not NOT1 (N8905, N8897);
nor NOR4 (N8906, N8900, N5757, N3998, N2459);
or OR2 (N8907, N8904, N4125);
or OR4 (N8908, N8901, N5121, N3471, N5429);
nand NAND4 (N8909, N8905, N366, N3982, N4713);
or OR3 (N8910, N8909, N7748, N2324);
and AND2 (N8911, N8896, N7972);
buf BUF1 (N8912, N8891);
nand NAND3 (N8913, N8902, N7857, N4359);
not NOT1 (N8914, N8872);
buf BUF1 (N8915, N8913);
xor XOR2 (N8916, N8903, N6734);
nor NOR3 (N8917, N8906, N4877, N2912);
nor NOR4 (N8918, N8911, N8406, N6859, N5166);
and AND3 (N8919, N8915, N3476, N2633);
xor XOR2 (N8920, N8917, N351);
nor NOR4 (N8921, N8914, N1887, N3183, N8365);
and AND3 (N8922, N8912, N1412, N6217);
buf BUF1 (N8923, N8919);
and AND4 (N8924, N8907, N6566, N5854, N1034);
or OR2 (N8925, N8923, N950);
not NOT1 (N8926, N8916);
or OR3 (N8927, N8926, N4980, N7749);
xor XOR2 (N8928, N8910, N8880);
not NOT1 (N8929, N8918);
and AND3 (N8930, N8925, N7075, N7353);
or OR3 (N8931, N8924, N8493, N5222);
not NOT1 (N8932, N8929);
and AND2 (N8933, N8922, N6119);
nor NOR4 (N8934, N8908, N7420, N7783, N6398);
or OR3 (N8935, N8920, N4190, N7776);
xor XOR2 (N8936, N8932, N4628);
buf BUF1 (N8937, N8927);
and AND4 (N8938, N8885, N4374, N433, N3216);
nand NAND2 (N8939, N8931, N1382);
nor NOR4 (N8940, N8936, N2199, N865, N1449);
buf BUF1 (N8941, N8934);
or OR3 (N8942, N8930, N7169, N5237);
nand NAND2 (N8943, N8942, N5054);
nand NAND2 (N8944, N8943, N3745);
xor XOR2 (N8945, N8939, N5886);
not NOT1 (N8946, N8938);
not NOT1 (N8947, N8928);
or OR3 (N8948, N8940, N6819, N3533);
or OR4 (N8949, N8948, N31, N2685, N4684);
nand NAND2 (N8950, N8921, N7067);
not NOT1 (N8951, N8933);
buf BUF1 (N8952, N8947);
not NOT1 (N8953, N8951);
nand NAND3 (N8954, N8953, N7619, N4443);
nand NAND3 (N8955, N8935, N7263, N5568);
xor XOR2 (N8956, N8937, N3343);
buf BUF1 (N8957, N8949);
not NOT1 (N8958, N8945);
not NOT1 (N8959, N8958);
and AND4 (N8960, N8952, N6860, N1744, N6245);
xor XOR2 (N8961, N8960, N7303);
not NOT1 (N8962, N8957);
or OR3 (N8963, N8955, N6667, N5255);
nor NOR2 (N8964, N8941, N1414);
or OR2 (N8965, N8956, N1710);
and AND3 (N8966, N8944, N4946, N8955);
nor NOR3 (N8967, N8959, N795, N7794);
xor XOR2 (N8968, N8946, N2614);
nand NAND4 (N8969, N8965, N2695, N3714, N3262);
buf BUF1 (N8970, N8969);
and AND3 (N8971, N8967, N2146, N5908);
or OR3 (N8972, N8954, N5617, N6319);
xor XOR2 (N8973, N8971, N6089);
nor NOR3 (N8974, N8950, N3485, N6436);
and AND3 (N8975, N8964, N2617, N5577);
not NOT1 (N8976, N8961);
nand NAND2 (N8977, N8968, N6926);
xor XOR2 (N8978, N8975, N347);
nor NOR3 (N8979, N8978, N1890, N8454);
nor NOR4 (N8980, N8966, N6381, N4436, N7695);
and AND2 (N8981, N8970, N6982);
or OR4 (N8982, N8981, N541, N3913, N7983);
buf BUF1 (N8983, N8980);
and AND4 (N8984, N8973, N3172, N8413, N7121);
nor NOR4 (N8985, N8976, N246, N3749, N3299);
nand NAND2 (N8986, N8979, N6988);
not NOT1 (N8987, N8986);
xor XOR2 (N8988, N8972, N188);
and AND2 (N8989, N8974, N5813);
nor NOR3 (N8990, N8988, N5101, N1208);
nand NAND3 (N8991, N8990, N6207, N2967);
buf BUF1 (N8992, N8987);
nand NAND4 (N8993, N8962, N6147, N2530, N8065);
xor XOR2 (N8994, N8989, N1974);
not NOT1 (N8995, N8983);
not NOT1 (N8996, N8963);
or OR2 (N8997, N8985, N8639);
or OR4 (N8998, N8993, N6615, N6831, N1481);
nand NAND3 (N8999, N8991, N4826, N7074);
nor NOR2 (N9000, N8996, N898);
and AND3 (N9001, N8999, N1078, N3722);
or OR3 (N9002, N9000, N6668, N5723);
nand NAND3 (N9003, N9001, N3264, N6315);
xor XOR2 (N9004, N8982, N3282);
and AND2 (N9005, N8992, N8945);
not NOT1 (N9006, N9004);
or OR2 (N9007, N9003, N2082);
xor XOR2 (N9008, N8998, N700);
or OR3 (N9009, N8997, N1387, N901);
not NOT1 (N9010, N9006);
and AND3 (N9011, N9005, N3166, N4515);
and AND4 (N9012, N8977, N217, N8164, N1984);
buf BUF1 (N9013, N9008);
xor XOR2 (N9014, N9007, N5447);
and AND4 (N9015, N9010, N6401, N3744, N5358);
xor XOR2 (N9016, N9012, N6798);
buf BUF1 (N9017, N9014);
xor XOR2 (N9018, N9015, N7128);
xor XOR2 (N9019, N9013, N1583);
buf BUF1 (N9020, N8994);
or OR3 (N9021, N9017, N5727, N3245);
and AND4 (N9022, N9002, N3442, N3043, N319);
and AND4 (N9023, N9018, N6789, N5684, N2620);
nor NOR3 (N9024, N9019, N6092, N7101);
or OR4 (N9025, N9023, N5125, N7509, N6376);
nand NAND2 (N9026, N9021, N6139);
buf BUF1 (N9027, N9020);
buf BUF1 (N9028, N8995);
xor XOR2 (N9029, N9011, N1829);
nand NAND3 (N9030, N9024, N3585, N5029);
or OR4 (N9031, N9016, N2709, N6651, N2750);
or OR4 (N9032, N9022, N7726, N8174, N6682);
and AND3 (N9033, N9029, N4483, N114);
buf BUF1 (N9034, N9028);
not NOT1 (N9035, N9026);
buf BUF1 (N9036, N9031);
and AND4 (N9037, N9027, N2151, N2190, N3587);
or OR4 (N9038, N9034, N995, N572, N5288);
xor XOR2 (N9039, N9038, N3368);
buf BUF1 (N9040, N8984);
xor XOR2 (N9041, N9009, N6889);
not NOT1 (N9042, N9037);
nand NAND4 (N9043, N9040, N2313, N5949, N7691);
nand NAND2 (N9044, N9039, N441);
and AND2 (N9045, N9036, N2107);
not NOT1 (N9046, N9044);
xor XOR2 (N9047, N9045, N8734);
buf BUF1 (N9048, N9043);
xor XOR2 (N9049, N9041, N3876);
or OR4 (N9050, N9030, N761, N860, N540);
buf BUF1 (N9051, N9035);
and AND4 (N9052, N9032, N3525, N5806, N4850);
or OR4 (N9053, N9050, N6724, N3539, N13);
nand NAND2 (N9054, N9052, N2776);
nor NOR3 (N9055, N9053, N5683, N4380);
xor XOR2 (N9056, N9046, N3120);
or OR2 (N9057, N9033, N4493);
and AND4 (N9058, N9055, N538, N6767, N6485);
nand NAND4 (N9059, N9051, N5753, N5114, N6755);
nor NOR2 (N9060, N9059, N3879);
or OR2 (N9061, N9047, N8879);
buf BUF1 (N9062, N9061);
not NOT1 (N9063, N9060);
nand NAND2 (N9064, N9025, N3423);
xor XOR2 (N9065, N9054, N6405);
buf BUF1 (N9066, N9064);
not NOT1 (N9067, N9057);
xor XOR2 (N9068, N9063, N4892);
nand NAND4 (N9069, N9056, N8499, N8599, N8815);
or OR2 (N9070, N9066, N993);
buf BUF1 (N9071, N9067);
xor XOR2 (N9072, N9062, N8620);
and AND2 (N9073, N9048, N8757);
and AND3 (N9074, N9068, N8752, N1287);
and AND2 (N9075, N9065, N2108);
not NOT1 (N9076, N9058);
and AND4 (N9077, N9071, N6799, N3775, N1449);
not NOT1 (N9078, N9072);
or OR3 (N9079, N9042, N7672, N7867);
and AND3 (N9080, N9077, N8168, N4495);
xor XOR2 (N9081, N9076, N3259);
buf BUF1 (N9082, N9081);
xor XOR2 (N9083, N9074, N5904);
nor NOR2 (N9084, N9080, N5695);
buf BUF1 (N9085, N9069);
or OR3 (N9086, N9070, N2652, N396);
not NOT1 (N9087, N9073);
buf BUF1 (N9088, N9087);
buf BUF1 (N9089, N9082);
nand NAND4 (N9090, N9085, N640, N6990, N1923);
buf BUF1 (N9091, N9088);
and AND4 (N9092, N9091, N5678, N4173, N2588);
buf BUF1 (N9093, N9075);
xor XOR2 (N9094, N9089, N5254);
nor NOR2 (N9095, N9079, N9008);
not NOT1 (N9096, N9093);
buf BUF1 (N9097, N9094);
nor NOR3 (N9098, N9097, N5434, N6736);
nor NOR3 (N9099, N9086, N1539, N5247);
xor XOR2 (N9100, N9049, N135);
not NOT1 (N9101, N9100);
buf BUF1 (N9102, N9095);
nor NOR3 (N9103, N9098, N4711, N1235);
nor NOR2 (N9104, N9090, N7227);
buf BUF1 (N9105, N9099);
and AND4 (N9106, N9103, N1270, N2649, N3611);
or OR3 (N9107, N9092, N9100, N3871);
nor NOR2 (N9108, N9096, N7739);
buf BUF1 (N9109, N9101);
not NOT1 (N9110, N9104);
xor XOR2 (N9111, N9105, N2544);
nor NOR3 (N9112, N9106, N3504, N5161);
not NOT1 (N9113, N9083);
nand NAND2 (N9114, N9078, N3730);
buf BUF1 (N9115, N9114);
not NOT1 (N9116, N9109);
nor NOR3 (N9117, N9111, N1238, N6536);
nand NAND2 (N9118, N9107, N689);
nor NOR3 (N9119, N9108, N1816, N6777);
and AND4 (N9120, N9113, N6393, N8982, N5007);
and AND3 (N9121, N9115, N7140, N5143);
and AND4 (N9122, N9116, N1271, N2013, N3979);
nand NAND4 (N9123, N9121, N2588, N4979, N419);
and AND4 (N9124, N9118, N7125, N3508, N3729);
nand NAND3 (N9125, N9123, N4582, N8131);
xor XOR2 (N9126, N9084, N8634);
nand NAND3 (N9127, N9102, N1133, N2936);
buf BUF1 (N9128, N9110);
and AND2 (N9129, N9127, N2055);
and AND4 (N9130, N9126, N5993, N8528, N7499);
or OR2 (N9131, N9122, N9095);
and AND2 (N9132, N9125, N6963);
and AND2 (N9133, N9128, N102);
and AND4 (N9134, N9131, N2662, N7425, N6332);
and AND4 (N9135, N9117, N8855, N3839, N12);
nand NAND3 (N9136, N9129, N7090, N6619);
nand NAND3 (N9137, N9133, N842, N2225);
or OR3 (N9138, N9120, N1687, N4384);
buf BUF1 (N9139, N9134);
nor NOR4 (N9140, N9135, N8752, N2110, N6754);
not NOT1 (N9141, N9136);
or OR3 (N9142, N9138, N7369, N1454);
nand NAND3 (N9143, N9141, N7259, N5617);
and AND4 (N9144, N9119, N1506, N7365, N4788);
buf BUF1 (N9145, N9130);
nand NAND3 (N9146, N9144, N302, N8467);
buf BUF1 (N9147, N9143);
not NOT1 (N9148, N9139);
xor XOR2 (N9149, N9137, N8893);
buf BUF1 (N9150, N9142);
or OR2 (N9151, N9147, N6198);
xor XOR2 (N9152, N9149, N8569);
xor XOR2 (N9153, N9140, N7621);
not NOT1 (N9154, N9124);
or OR2 (N9155, N9152, N4259);
nand NAND3 (N9156, N9148, N4091, N7199);
not NOT1 (N9157, N9155);
buf BUF1 (N9158, N9146);
xor XOR2 (N9159, N9150, N9056);
or OR4 (N9160, N9151, N570, N7087, N6847);
or OR4 (N9161, N9112, N5563, N3998, N6126);
xor XOR2 (N9162, N9158, N3);
or OR2 (N9163, N9145, N1007);
xor XOR2 (N9164, N9154, N5888);
xor XOR2 (N9165, N9161, N5095);
nand NAND2 (N9166, N9164, N8404);
not NOT1 (N9167, N9160);
nand NAND3 (N9168, N9153, N582, N7572);
and AND3 (N9169, N9157, N6875, N5710);
buf BUF1 (N9170, N9163);
or OR3 (N9171, N9170, N7889, N6000);
xor XOR2 (N9172, N9162, N8711);
nand NAND2 (N9173, N9159, N4357);
and AND3 (N9174, N9169, N1186, N8777);
or OR4 (N9175, N9172, N2463, N9124, N7095);
xor XOR2 (N9176, N9167, N8110);
nor NOR4 (N9177, N9176, N305, N2296, N1112);
xor XOR2 (N9178, N9168, N6552);
or OR3 (N9179, N9174, N6544, N5723);
or OR3 (N9180, N9175, N8976, N4430);
buf BUF1 (N9181, N9173);
and AND4 (N9182, N9132, N4056, N3882, N1899);
not NOT1 (N9183, N9182);
and AND3 (N9184, N9178, N8729, N6619);
or OR4 (N9185, N9166, N1119, N5589, N8845);
not NOT1 (N9186, N9179);
not NOT1 (N9187, N9177);
and AND3 (N9188, N9184, N5340, N2197);
buf BUF1 (N9189, N9183);
not NOT1 (N9190, N9156);
or OR2 (N9191, N9188, N6555);
xor XOR2 (N9192, N9165, N260);
buf BUF1 (N9193, N9187);
nor NOR3 (N9194, N9185, N4232, N750);
and AND4 (N9195, N9194, N7295, N2180, N6660);
xor XOR2 (N9196, N9190, N7605);
nand NAND3 (N9197, N9191, N8924, N1850);
nand NAND3 (N9198, N9192, N4310, N5852);
not NOT1 (N9199, N9195);
buf BUF1 (N9200, N9198);
or OR4 (N9201, N9193, N3138, N126, N4153);
buf BUF1 (N9202, N9196);
buf BUF1 (N9203, N9197);
nand NAND2 (N9204, N9202, N5352);
xor XOR2 (N9205, N9171, N8723);
nand NAND4 (N9206, N9180, N6974, N1427, N7390);
buf BUF1 (N9207, N9205);
xor XOR2 (N9208, N9204, N6839);
and AND4 (N9209, N9203, N4523, N1253, N3872);
nand NAND3 (N9210, N9208, N5578, N7363);
xor XOR2 (N9211, N9201, N3828);
nor NOR3 (N9212, N9209, N1935, N7903);
xor XOR2 (N9213, N9189, N1462);
not NOT1 (N9214, N9211);
buf BUF1 (N9215, N9200);
buf BUF1 (N9216, N9199);
buf BUF1 (N9217, N9212);
nand NAND3 (N9218, N9217, N1005, N7274);
nor NOR3 (N9219, N9214, N2418, N1198);
nor NOR3 (N9220, N9207, N2454, N595);
or OR2 (N9221, N9218, N3729);
buf BUF1 (N9222, N9210);
and AND3 (N9223, N9222, N1346, N7880);
or OR3 (N9224, N9219, N5504, N7667);
not NOT1 (N9225, N9186);
nand NAND3 (N9226, N9206, N7056, N7056);
nor NOR2 (N9227, N9181, N4057);
nor NOR3 (N9228, N9215, N3727, N7128);
and AND3 (N9229, N9225, N1166, N2974);
and AND3 (N9230, N9228, N9104, N242);
buf BUF1 (N9231, N9216);
and AND3 (N9232, N9227, N6963, N1735);
or OR2 (N9233, N9213, N1425);
and AND4 (N9234, N9230, N5503, N2529, N6071);
buf BUF1 (N9235, N9223);
nor NOR2 (N9236, N9229, N1808);
or OR4 (N9237, N9224, N826, N8622, N1479);
buf BUF1 (N9238, N9236);
and AND2 (N9239, N9235, N4629);
and AND2 (N9240, N9221, N7369);
xor XOR2 (N9241, N9238, N2840);
nor NOR4 (N9242, N9241, N7337, N4910, N8311);
buf BUF1 (N9243, N9220);
nor NOR3 (N9244, N9231, N4028, N456);
or OR2 (N9245, N9242, N8222);
and AND4 (N9246, N9239, N5084, N4989, N7161);
buf BUF1 (N9247, N9234);
or OR3 (N9248, N9237, N1223, N5118);
not NOT1 (N9249, N9233);
or OR3 (N9250, N9240, N6454, N814);
and AND3 (N9251, N9248, N7085, N4652);
or OR2 (N9252, N9250, N8220);
buf BUF1 (N9253, N9232);
not NOT1 (N9254, N9243);
buf BUF1 (N9255, N9245);
nand NAND4 (N9256, N9226, N8802, N4014, N3541);
nand NAND4 (N9257, N9252, N4187, N9088, N7693);
nand NAND3 (N9258, N9253, N2272, N651);
xor XOR2 (N9259, N9251, N3074);
and AND4 (N9260, N9258, N492, N6373, N979);
and AND3 (N9261, N9257, N8837, N5785);
xor XOR2 (N9262, N9259, N5264);
xor XOR2 (N9263, N9249, N4429);
and AND4 (N9264, N9244, N1327, N7668, N1297);
nor NOR4 (N9265, N9264, N1466, N7770, N4692);
not NOT1 (N9266, N9261);
xor XOR2 (N9267, N9262, N1066);
nand NAND4 (N9268, N9255, N4745, N6319, N1162);
nor NOR4 (N9269, N9246, N8184, N124, N7341);
nand NAND2 (N9270, N9256, N4766);
or OR2 (N9271, N9270, N9009);
buf BUF1 (N9272, N9254);
or OR3 (N9273, N9266, N4008, N5285);
and AND2 (N9274, N9271, N2839);
and AND2 (N9275, N9265, N2981);
or OR4 (N9276, N9274, N4211, N8226, N5003);
xor XOR2 (N9277, N9275, N381);
nand NAND2 (N9278, N9273, N1091);
nand NAND3 (N9279, N9276, N2411, N3519);
buf BUF1 (N9280, N9278);
xor XOR2 (N9281, N9267, N3037);
nand NAND3 (N9282, N9260, N2606, N2782);
or OR2 (N9283, N9268, N7141);
xor XOR2 (N9284, N9263, N6672);
xor XOR2 (N9285, N9280, N3491);
nand NAND4 (N9286, N9285, N141, N7963, N8358);
xor XOR2 (N9287, N9282, N1142);
or OR3 (N9288, N9272, N820, N6939);
or OR2 (N9289, N9288, N2591);
xor XOR2 (N9290, N9269, N4395);
and AND2 (N9291, N9290, N6953);
xor XOR2 (N9292, N9286, N4817);
nand NAND2 (N9293, N9277, N884);
nand NAND3 (N9294, N9287, N7727, N4191);
buf BUF1 (N9295, N9281);
nand NAND4 (N9296, N9279, N1524, N5326, N4726);
or OR3 (N9297, N9292, N8986, N8933);
or OR3 (N9298, N9293, N1684, N6189);
and AND4 (N9299, N9296, N4535, N5113, N751);
not NOT1 (N9300, N9295);
or OR4 (N9301, N9299, N2426, N4419, N1866);
not NOT1 (N9302, N9301);
buf BUF1 (N9303, N9297);
nor NOR4 (N9304, N9284, N5145, N852, N8879);
not NOT1 (N9305, N9294);
xor XOR2 (N9306, N9289, N7847);
buf BUF1 (N9307, N9283);
nor NOR2 (N9308, N9298, N9261);
not NOT1 (N9309, N9303);
and AND4 (N9310, N9306, N9256, N611, N6098);
nand NAND4 (N9311, N9300, N1254, N4973, N8734);
and AND3 (N9312, N9308, N459, N5420);
and AND2 (N9313, N9302, N4914);
xor XOR2 (N9314, N9304, N5325);
not NOT1 (N9315, N9309);
or OR3 (N9316, N9315, N2933, N5694);
nand NAND3 (N9317, N9311, N6571, N2264);
or OR4 (N9318, N9307, N3459, N3262, N6115);
buf BUF1 (N9319, N9247);
and AND4 (N9320, N9317, N6195, N5352, N3291);
or OR3 (N9321, N9313, N8781, N4155);
xor XOR2 (N9322, N9305, N2771);
or OR2 (N9323, N9322, N1902);
buf BUF1 (N9324, N9320);
not NOT1 (N9325, N9310);
nor NOR3 (N9326, N9319, N2812, N1311);
or OR2 (N9327, N9318, N1167);
xor XOR2 (N9328, N9323, N6499);
nand NAND3 (N9329, N9328, N1698, N3426);
nand NAND3 (N9330, N9312, N9253, N2056);
nor NOR3 (N9331, N9330, N2975, N1664);
nand NAND3 (N9332, N9329, N6389, N1131);
buf BUF1 (N9333, N9332);
nor NOR3 (N9334, N9324, N6168, N1553);
nor NOR4 (N9335, N9331, N3922, N5594, N3948);
nand NAND3 (N9336, N9314, N9271, N8057);
buf BUF1 (N9337, N9336);
and AND2 (N9338, N9326, N7588);
and AND2 (N9339, N9335, N6079);
xor XOR2 (N9340, N9339, N3667);
or OR3 (N9341, N9340, N8860, N3809);
nor NOR2 (N9342, N9337, N9081);
not NOT1 (N9343, N9327);
xor XOR2 (N9344, N9343, N7518);
nand NAND3 (N9345, N9316, N6496, N4389);
or OR3 (N9346, N9291, N4177, N664);
or OR3 (N9347, N9344, N3166, N9192);
buf BUF1 (N9348, N9342);
or OR4 (N9349, N9348, N406, N8205, N6084);
nor NOR4 (N9350, N9321, N5503, N5476, N6448);
and AND4 (N9351, N9333, N5149, N2250, N2097);
not NOT1 (N9352, N9325);
xor XOR2 (N9353, N9341, N2579);
and AND3 (N9354, N9334, N4180, N2216);
nand NAND4 (N9355, N9346, N3786, N3525, N2902);
buf BUF1 (N9356, N9345);
nor NOR4 (N9357, N9352, N7011, N4414, N8186);
buf BUF1 (N9358, N9349);
or OR3 (N9359, N9353, N1463, N5791);
or OR2 (N9360, N9347, N6682);
and AND4 (N9361, N9351, N2546, N6575, N1932);
nor NOR2 (N9362, N9360, N2455);
or OR3 (N9363, N9362, N4060, N3954);
xor XOR2 (N9364, N9358, N6795);
nand NAND3 (N9365, N9350, N8404, N7057);
nand NAND4 (N9366, N9363, N4825, N4951, N8161);
nor NOR2 (N9367, N9364, N1497);
not NOT1 (N9368, N9359);
nand NAND3 (N9369, N9365, N6976, N9276);
not NOT1 (N9370, N9369);
nor NOR2 (N9371, N9356, N7350);
buf BUF1 (N9372, N9368);
or OR4 (N9373, N9361, N8307, N2285, N6402);
nand NAND2 (N9374, N9367, N7879);
nand NAND4 (N9375, N9373, N839, N1750, N7259);
or OR4 (N9376, N9370, N7622, N5390, N130);
and AND4 (N9377, N9338, N2842, N6132, N8605);
buf BUF1 (N9378, N9377);
buf BUF1 (N9379, N9355);
buf BUF1 (N9380, N9371);
and AND2 (N9381, N9374, N7406);
xor XOR2 (N9382, N9380, N7443);
nand NAND3 (N9383, N9354, N1129, N8635);
and AND3 (N9384, N9378, N6267, N5232);
not NOT1 (N9385, N9379);
nor NOR2 (N9386, N9372, N9005);
and AND4 (N9387, N9381, N7447, N5910, N2688);
nor NOR3 (N9388, N9376, N260, N565);
and AND2 (N9389, N9384, N718);
xor XOR2 (N9390, N9388, N8913);
not NOT1 (N9391, N9383);
and AND2 (N9392, N9375, N388);
nor NOR4 (N9393, N9392, N7130, N780, N1381);
not NOT1 (N9394, N9389);
buf BUF1 (N9395, N9394);
nand NAND4 (N9396, N9385, N1305, N970, N6227);
xor XOR2 (N9397, N9386, N2010);
or OR3 (N9398, N9391, N6316, N4127);
and AND4 (N9399, N9357, N5466, N4463, N2603);
buf BUF1 (N9400, N9390);
buf BUF1 (N9401, N9398);
or OR2 (N9402, N9401, N324);
or OR2 (N9403, N9399, N8659);
buf BUF1 (N9404, N9403);
not NOT1 (N9405, N9402);
xor XOR2 (N9406, N9387, N2699);
not NOT1 (N9407, N9366);
nand NAND3 (N9408, N9396, N4179, N3192);
buf BUF1 (N9409, N9400);
nor NOR3 (N9410, N9405, N1585, N628);
or OR2 (N9411, N9407, N5203);
nor NOR3 (N9412, N9406, N4181, N6756);
or OR3 (N9413, N9393, N1070, N3277);
nor NOR2 (N9414, N9404, N4018);
nor NOR4 (N9415, N9413, N6961, N8986, N4792);
nor NOR2 (N9416, N9397, N8507);
not NOT1 (N9417, N9409);
or OR2 (N9418, N9411, N4108);
and AND4 (N9419, N9418, N8043, N4945, N4168);
not NOT1 (N9420, N9410);
and AND3 (N9421, N9412, N8183, N8469);
not NOT1 (N9422, N9421);
and AND2 (N9423, N9416, N794);
not NOT1 (N9424, N9417);
nor NOR4 (N9425, N9382, N1403, N2405, N7985);
not NOT1 (N9426, N9425);
and AND2 (N9427, N9422, N5447);
nand NAND2 (N9428, N9408, N7510);
not NOT1 (N9429, N9426);
nand NAND2 (N9430, N9427, N9137);
nor NOR2 (N9431, N9395, N8076);
xor XOR2 (N9432, N9424, N7054);
buf BUF1 (N9433, N9420);
buf BUF1 (N9434, N9423);
xor XOR2 (N9435, N9433, N2091);
and AND3 (N9436, N9434, N8094, N2562);
buf BUF1 (N9437, N9428);
buf BUF1 (N9438, N9429);
nor NOR4 (N9439, N9438, N5024, N8387, N4539);
xor XOR2 (N9440, N9437, N5748);
not NOT1 (N9441, N9431);
nand NAND3 (N9442, N9436, N2875, N5495);
nand NAND2 (N9443, N9432, N7474);
nor NOR4 (N9444, N9415, N6120, N7391, N7169);
not NOT1 (N9445, N9444);
xor XOR2 (N9446, N9445, N9372);
or OR3 (N9447, N9439, N9119, N7482);
xor XOR2 (N9448, N9446, N1136);
xor XOR2 (N9449, N9419, N4501);
xor XOR2 (N9450, N9447, N2115);
and AND3 (N9451, N9442, N4631, N4235);
not NOT1 (N9452, N9449);
and AND4 (N9453, N9414, N8387, N6141, N5949);
nor NOR3 (N9454, N9452, N3272, N55);
or OR4 (N9455, N9450, N4417, N4817, N1534);
or OR3 (N9456, N9443, N8046, N4677);
not NOT1 (N9457, N9430);
and AND4 (N9458, N9435, N4374, N1383, N6688);
and AND2 (N9459, N9456, N4404);
or OR3 (N9460, N9440, N67, N3908);
nor NOR3 (N9461, N9457, N3590, N1170);
or OR4 (N9462, N9455, N5203, N3736, N1778);
buf BUF1 (N9463, N9448);
nand NAND3 (N9464, N9441, N5001, N7366);
xor XOR2 (N9465, N9454, N2608);
buf BUF1 (N9466, N9458);
buf BUF1 (N9467, N9460);
xor XOR2 (N9468, N9453, N960);
not NOT1 (N9469, N9466);
buf BUF1 (N9470, N9463);
buf BUF1 (N9471, N9451);
not NOT1 (N9472, N9469);
nor NOR4 (N9473, N9470, N300, N1390, N3497);
not NOT1 (N9474, N9464);
xor XOR2 (N9475, N9465, N4911);
nand NAND2 (N9476, N9467, N8519);
or OR3 (N9477, N9459, N7926, N2297);
buf BUF1 (N9478, N9475);
xor XOR2 (N9479, N9471, N5344);
or OR3 (N9480, N9473, N5749, N8197);
not NOT1 (N9481, N9479);
xor XOR2 (N9482, N9462, N2277);
or OR2 (N9483, N9477, N6291);
or OR3 (N9484, N9480, N6647, N8441);
or OR3 (N9485, N9472, N4272, N6015);
nor NOR4 (N9486, N9482, N5946, N7179, N3849);
xor XOR2 (N9487, N9485, N9451);
buf BUF1 (N9488, N9481);
xor XOR2 (N9489, N9474, N4751);
not NOT1 (N9490, N9484);
not NOT1 (N9491, N9488);
xor XOR2 (N9492, N9486, N9345);
or OR3 (N9493, N9468, N2159, N1743);
buf BUF1 (N9494, N9492);
nand NAND4 (N9495, N9489, N7050, N8667, N4951);
and AND2 (N9496, N9487, N7823);
nor NOR3 (N9497, N9491, N422, N5842);
buf BUF1 (N9498, N9495);
and AND3 (N9499, N9461, N628, N226);
not NOT1 (N9500, N9499);
buf BUF1 (N9501, N9476);
or OR2 (N9502, N9496, N7017);
nor NOR3 (N9503, N9490, N1226, N2731);
or OR4 (N9504, N9483, N2875, N8997, N6086);
nand NAND3 (N9505, N9498, N1138, N7808);
not NOT1 (N9506, N9505);
or OR3 (N9507, N9501, N9200, N3364);
buf BUF1 (N9508, N9504);
nand NAND3 (N9509, N9503, N8923, N705);
and AND4 (N9510, N9497, N1884, N64, N7428);
buf BUF1 (N9511, N9502);
buf BUF1 (N9512, N9509);
nor NOR4 (N9513, N9507, N17, N5092, N1585);
nand NAND3 (N9514, N9500, N7834, N2082);
xor XOR2 (N9515, N9478, N8168);
nor NOR2 (N9516, N9506, N5383);
nor NOR4 (N9517, N9511, N2183, N3631, N3522);
nor NOR3 (N9518, N9493, N7936, N1532);
and AND3 (N9519, N9514, N4094, N8235);
or OR3 (N9520, N9515, N4959, N5751);
nand NAND4 (N9521, N9516, N3299, N9347, N9195);
nor NOR3 (N9522, N9519, N2199, N2421);
and AND3 (N9523, N9512, N560, N8114);
not NOT1 (N9524, N9508);
nand NAND3 (N9525, N9523, N4617, N2474);
and AND2 (N9526, N9494, N6692);
or OR2 (N9527, N9520, N1075);
nand NAND3 (N9528, N9522, N6862, N8779);
xor XOR2 (N9529, N9513, N5105);
nand NAND2 (N9530, N9528, N2121);
and AND3 (N9531, N9527, N7101, N2934);
or OR2 (N9532, N9518, N2031);
nand NAND4 (N9533, N9532, N4571, N444, N8237);
nand NAND2 (N9534, N9529, N5992);
and AND3 (N9535, N9525, N5584, N5749);
and AND3 (N9536, N9521, N992, N8860);
or OR2 (N9537, N9510, N425);
nor NOR3 (N9538, N9531, N8850, N1032);
and AND4 (N9539, N9526, N238, N4010, N3382);
and AND4 (N9540, N9517, N1797, N1872, N1846);
xor XOR2 (N9541, N9524, N6837);
not NOT1 (N9542, N9537);
not NOT1 (N9543, N9534);
xor XOR2 (N9544, N9536, N5081);
nor NOR4 (N9545, N9540, N6640, N2767, N8129);
not NOT1 (N9546, N9538);
xor XOR2 (N9547, N9533, N8871);
xor XOR2 (N9548, N9530, N5203);
xor XOR2 (N9549, N9539, N7838);
not NOT1 (N9550, N9549);
buf BUF1 (N9551, N9548);
xor XOR2 (N9552, N9547, N163);
not NOT1 (N9553, N9543);
not NOT1 (N9554, N9553);
nand NAND2 (N9555, N9544, N923);
nand NAND2 (N9556, N9551, N175);
nor NOR3 (N9557, N9555, N7302, N8918);
nand NAND4 (N9558, N9545, N737, N3415, N514);
not NOT1 (N9559, N9550);
nor NOR4 (N9560, N9552, N1836, N4108, N4425);
nor NOR2 (N9561, N9554, N6327);
xor XOR2 (N9562, N9560, N2736);
or OR2 (N9563, N9559, N360);
nand NAND2 (N9564, N9535, N4880);
not NOT1 (N9565, N9557);
or OR2 (N9566, N9564, N7677);
not NOT1 (N9567, N9561);
nand NAND2 (N9568, N9565, N3117);
not NOT1 (N9569, N9556);
or OR4 (N9570, N9562, N6705, N2351, N7833);
nand NAND4 (N9571, N9567, N334, N8564, N2242);
xor XOR2 (N9572, N9546, N4248);
buf BUF1 (N9573, N9566);
and AND4 (N9574, N9571, N4260, N5228, N6362);
xor XOR2 (N9575, N9541, N676);
not NOT1 (N9576, N9563);
not NOT1 (N9577, N9569);
and AND3 (N9578, N9574, N1544, N473);
buf BUF1 (N9579, N9578);
nor NOR3 (N9580, N9575, N3402, N7500);
buf BUF1 (N9581, N9572);
nor NOR2 (N9582, N9576, N1665);
buf BUF1 (N9583, N9568);
xor XOR2 (N9584, N9573, N2959);
or OR2 (N9585, N9577, N4126);
or OR3 (N9586, N9570, N5367, N6007);
nor NOR4 (N9587, N9579, N2227, N1288, N5247);
not NOT1 (N9588, N9582);
and AND3 (N9589, N9580, N7597, N2987);
buf BUF1 (N9590, N9558);
nor NOR2 (N9591, N9586, N2330);
buf BUF1 (N9592, N9581);
or OR4 (N9593, N9587, N5743, N8288, N9513);
and AND2 (N9594, N9590, N5400);
nand NAND4 (N9595, N9584, N8166, N8412, N4308);
nor NOR2 (N9596, N9583, N8891);
buf BUF1 (N9597, N9595);
nor NOR3 (N9598, N9542, N933, N6490);
or OR2 (N9599, N9592, N7356);
nand NAND2 (N9600, N9585, N8492);
nand NAND2 (N9601, N9597, N8199);
and AND4 (N9602, N9599, N2813, N8446, N1189);
xor XOR2 (N9603, N9596, N1175);
not NOT1 (N9604, N9591);
not NOT1 (N9605, N9598);
and AND4 (N9606, N9601, N3508, N59, N6051);
or OR4 (N9607, N9606, N4473, N6335, N2376);
nand NAND2 (N9608, N9603, N6192);
nor NOR2 (N9609, N9588, N7211);
buf BUF1 (N9610, N9600);
nor NOR4 (N9611, N9589, N1153, N2276, N1009);
or OR4 (N9612, N9610, N5499, N7517, N390);
buf BUF1 (N9613, N9612);
and AND3 (N9614, N9608, N4258, N5142);
nand NAND2 (N9615, N9609, N1599);
not NOT1 (N9616, N9593);
not NOT1 (N9617, N9594);
xor XOR2 (N9618, N9616, N5608);
and AND4 (N9619, N9605, N7484, N6680, N316);
not NOT1 (N9620, N9618);
xor XOR2 (N9621, N9607, N8621);
nand NAND4 (N9622, N9617, N8284, N8269, N5882);
buf BUF1 (N9623, N9615);
nand NAND2 (N9624, N9614, N8622);
and AND4 (N9625, N9602, N1814, N312, N6718);
or OR4 (N9626, N9621, N1018, N3096, N1110);
nand NAND3 (N9627, N9626, N2332, N2507);
or OR2 (N9628, N9604, N2883);
xor XOR2 (N9629, N9625, N627);
nand NAND3 (N9630, N9624, N4507, N7952);
xor XOR2 (N9631, N9630, N5881);
nor NOR3 (N9632, N9619, N1966, N7296);
xor XOR2 (N9633, N9613, N7852);
not NOT1 (N9634, N9620);
or OR3 (N9635, N9628, N4273, N2351);
buf BUF1 (N9636, N9622);
not NOT1 (N9637, N9627);
and AND4 (N9638, N9611, N7773, N6918, N2407);
buf BUF1 (N9639, N9638);
and AND3 (N9640, N9635, N2587, N3959);
nor NOR3 (N9641, N9637, N3409, N3550);
not NOT1 (N9642, N9632);
or OR4 (N9643, N9640, N3604, N8439, N8035);
buf BUF1 (N9644, N9636);
or OR4 (N9645, N9639, N6454, N429, N3076);
nand NAND2 (N9646, N9631, N5905);
not NOT1 (N9647, N9641);
not NOT1 (N9648, N9647);
and AND4 (N9649, N9643, N5587, N9513, N8608);
not NOT1 (N9650, N9633);
nand NAND3 (N9651, N9629, N9340, N809);
nor NOR3 (N9652, N9648, N7444, N6937);
nand NAND3 (N9653, N9651, N4053, N7901);
nor NOR3 (N9654, N9634, N8072, N8628);
xor XOR2 (N9655, N9646, N5775);
nor NOR4 (N9656, N9649, N6535, N2051, N2150);
nor NOR4 (N9657, N9650, N7265, N5627, N5882);
or OR2 (N9658, N9656, N1924);
and AND4 (N9659, N9654, N444, N4497, N1325);
nor NOR4 (N9660, N9642, N9192, N6182, N1145);
xor XOR2 (N9661, N9659, N466);
xor XOR2 (N9662, N9645, N4036);
xor XOR2 (N9663, N9661, N1793);
buf BUF1 (N9664, N9657);
nand NAND4 (N9665, N9658, N7760, N6747, N8208);
not NOT1 (N9666, N9664);
or OR2 (N9667, N9660, N6500);
nor NOR3 (N9668, N9652, N124, N4072);
nor NOR4 (N9669, N9623, N7335, N8627, N4652);
xor XOR2 (N9670, N9666, N7510);
nand NAND4 (N9671, N9644, N7386, N9420, N8589);
nand NAND2 (N9672, N9667, N2772);
and AND3 (N9673, N9671, N4025, N7856);
xor XOR2 (N9674, N9672, N8921);
buf BUF1 (N9675, N9655);
nand NAND4 (N9676, N9668, N4975, N8785, N8867);
or OR3 (N9677, N9663, N7292, N1164);
not NOT1 (N9678, N9669);
or OR3 (N9679, N9675, N2287, N3870);
or OR3 (N9680, N9674, N6324, N1459);
nor NOR4 (N9681, N9678, N6707, N7356, N6017);
xor XOR2 (N9682, N9662, N7944);
nor NOR2 (N9683, N9676, N2277);
not NOT1 (N9684, N9665);
or OR3 (N9685, N9681, N2180, N2813);
and AND4 (N9686, N9682, N4935, N6314, N5545);
nand NAND3 (N9687, N9685, N8321, N3839);
and AND3 (N9688, N9683, N8274, N8632);
and AND2 (N9689, N9687, N2082);
nor NOR2 (N9690, N9677, N8239);
not NOT1 (N9691, N9690);
buf BUF1 (N9692, N9670);
nand NAND3 (N9693, N9686, N8958, N8394);
buf BUF1 (N9694, N9688);
nand NAND2 (N9695, N9684, N510);
and AND2 (N9696, N9692, N1501);
nand NAND4 (N9697, N9695, N445, N7268, N597);
and AND2 (N9698, N9694, N3687);
not NOT1 (N9699, N9691);
buf BUF1 (N9700, N9696);
buf BUF1 (N9701, N9693);
buf BUF1 (N9702, N9699);
nand NAND4 (N9703, N9700, N3327, N6410, N2042);
nor NOR2 (N9704, N9702, N5722);
xor XOR2 (N9705, N9653, N3468);
or OR3 (N9706, N9703, N6601, N1723);
xor XOR2 (N9707, N9701, N7056);
or OR4 (N9708, N9698, N4285, N3331, N5387);
buf BUF1 (N9709, N9679);
xor XOR2 (N9710, N9709, N8461);
or OR4 (N9711, N9710, N3158, N4946, N4745);
buf BUF1 (N9712, N9705);
nand NAND4 (N9713, N9697, N5219, N2331, N8512);
nand NAND2 (N9714, N9711, N2110);
buf BUF1 (N9715, N9713);
not NOT1 (N9716, N9706);
or OR2 (N9717, N9716, N8346);
nand NAND3 (N9718, N9707, N8839, N8112);
buf BUF1 (N9719, N9689);
nor NOR3 (N9720, N9712, N1979, N2959);
or OR3 (N9721, N9718, N2602, N1558);
or OR4 (N9722, N9680, N718, N584, N4112);
buf BUF1 (N9723, N9717);
nor NOR2 (N9724, N9721, N5337);
not NOT1 (N9725, N9714);
nand NAND3 (N9726, N9673, N6435, N8758);
nand NAND4 (N9727, N9719, N1284, N523, N7681);
and AND2 (N9728, N9725, N4528);
and AND2 (N9729, N9727, N9457);
nor NOR2 (N9730, N9708, N6652);
nand NAND2 (N9731, N9726, N6068);
nor NOR3 (N9732, N9720, N2597, N599);
xor XOR2 (N9733, N9731, N8701);
or OR4 (N9734, N9732, N2853, N6776, N4572);
xor XOR2 (N9735, N9728, N485);
nor NOR4 (N9736, N9724, N867, N867, N1288);
not NOT1 (N9737, N9735);
nor NOR3 (N9738, N9730, N1701, N3383);
or OR2 (N9739, N9723, N3078);
nand NAND2 (N9740, N9738, N6661);
buf BUF1 (N9741, N9737);
not NOT1 (N9742, N9739);
xor XOR2 (N9743, N9736, N4255);
nand NAND2 (N9744, N9722, N6301);
not NOT1 (N9745, N9743);
buf BUF1 (N9746, N9715);
xor XOR2 (N9747, N9741, N1962);
nor NOR4 (N9748, N9733, N1084, N7469, N1423);
nand NAND3 (N9749, N9744, N8074, N512);
xor XOR2 (N9750, N9742, N441);
not NOT1 (N9751, N9734);
xor XOR2 (N9752, N9750, N5481);
and AND3 (N9753, N9748, N4824, N5894);
nor NOR3 (N9754, N9752, N5905, N5978);
nand NAND4 (N9755, N9749, N6484, N2043, N1470);
or OR2 (N9756, N9745, N1616);
and AND3 (N9757, N9746, N2974, N9181);
not NOT1 (N9758, N9753);
xor XOR2 (N9759, N9729, N222);
buf BUF1 (N9760, N9759);
xor XOR2 (N9761, N9758, N8803);
xor XOR2 (N9762, N9756, N472);
and AND3 (N9763, N9761, N3202, N5080);
nand NAND4 (N9764, N9757, N8185, N833, N4312);
or OR2 (N9765, N9762, N3666);
and AND3 (N9766, N9704, N4202, N1002);
or OR3 (N9767, N9764, N3530, N1862);
buf BUF1 (N9768, N9767);
nand NAND4 (N9769, N9740, N8157, N3586, N5698);
nand NAND2 (N9770, N9755, N9004);
xor XOR2 (N9771, N9747, N409);
xor XOR2 (N9772, N9768, N141);
nand NAND3 (N9773, N9770, N6453, N4820);
nand NAND2 (N9774, N9765, N6968);
nor NOR2 (N9775, N9766, N9647);
buf BUF1 (N9776, N9751);
not NOT1 (N9777, N9763);
buf BUF1 (N9778, N9760);
xor XOR2 (N9779, N9772, N3006);
or OR2 (N9780, N9773, N2552);
buf BUF1 (N9781, N9778);
nand NAND4 (N9782, N9777, N4496, N3565, N674);
nand NAND4 (N9783, N9775, N5289, N4366, N4527);
and AND3 (N9784, N9780, N3198, N5365);
or OR3 (N9785, N9779, N3119, N3624);
not NOT1 (N9786, N9783);
buf BUF1 (N9787, N9769);
nand NAND4 (N9788, N9784, N2072, N5892, N7399);
not NOT1 (N9789, N9782);
buf BUF1 (N9790, N9788);
nand NAND3 (N9791, N9790, N9369, N543);
not NOT1 (N9792, N9791);
not NOT1 (N9793, N9785);
buf BUF1 (N9794, N9754);
nor NOR2 (N9795, N9789, N340);
nand NAND3 (N9796, N9776, N5427, N1081);
nor NOR3 (N9797, N9786, N3365, N9571);
not NOT1 (N9798, N9796);
xor XOR2 (N9799, N9794, N9446);
buf BUF1 (N9800, N9792);
buf BUF1 (N9801, N9781);
nand NAND4 (N9802, N9795, N8418, N4910, N3434);
not NOT1 (N9803, N9793);
nor NOR3 (N9804, N9797, N475, N9420);
buf BUF1 (N9805, N9799);
xor XOR2 (N9806, N9771, N669);
or OR3 (N9807, N9774, N4183, N7842);
nor NOR3 (N9808, N9807, N6102, N7101);
nand NAND2 (N9809, N9801, N8512);
nand NAND4 (N9810, N9798, N8501, N5945, N6218);
nand NAND3 (N9811, N9803, N4657, N3939);
xor XOR2 (N9812, N9787, N9420);
and AND2 (N9813, N9811, N7141);
and AND4 (N9814, N9813, N1138, N9063, N7555);
nand NAND3 (N9815, N9800, N2804, N1469);
xor XOR2 (N9816, N9804, N6720);
not NOT1 (N9817, N9808);
and AND3 (N9818, N9816, N4491, N4327);
xor XOR2 (N9819, N9812, N2311);
buf BUF1 (N9820, N9810);
or OR4 (N9821, N9809, N3480, N6384, N6921);
nand NAND4 (N9822, N9818, N6144, N4899, N5007);
xor XOR2 (N9823, N9817, N9434);
nand NAND3 (N9824, N9806, N6680, N6273);
nor NOR4 (N9825, N9814, N3121, N921, N9428);
xor XOR2 (N9826, N9822, N561);
not NOT1 (N9827, N9823);
nor NOR4 (N9828, N9802, N1054, N3719, N698);
nand NAND3 (N9829, N9825, N7394, N3805);
xor XOR2 (N9830, N9828, N5537);
not NOT1 (N9831, N9826);
nand NAND2 (N9832, N9805, N4871);
not NOT1 (N9833, N9830);
and AND3 (N9834, N9815, N4841, N236);
not NOT1 (N9835, N9831);
or OR2 (N9836, N9819, N3852);
nor NOR4 (N9837, N9836, N4137, N5914, N65);
not NOT1 (N9838, N9821);
buf BUF1 (N9839, N9838);
nand NAND2 (N9840, N9837, N762);
nand NAND3 (N9841, N9829, N256, N5972);
nor NOR4 (N9842, N9834, N1186, N1471, N8641);
not NOT1 (N9843, N9841);
not NOT1 (N9844, N9835);
or OR3 (N9845, N9832, N259, N893);
buf BUF1 (N9846, N9842);
nor NOR2 (N9847, N9845, N118);
xor XOR2 (N9848, N9833, N8336);
buf BUF1 (N9849, N9844);
or OR4 (N9850, N9847, N2316, N8762, N5500);
not NOT1 (N9851, N9846);
nand NAND2 (N9852, N9827, N6825);
nand NAND2 (N9853, N9851, N1852);
and AND3 (N9854, N9840, N1230, N1960);
nand NAND2 (N9855, N9850, N4463);
nand NAND4 (N9856, N9824, N8207, N5338, N853);
nand NAND3 (N9857, N9843, N5750, N5011);
xor XOR2 (N9858, N9854, N6127);
and AND3 (N9859, N9858, N853, N4591);
and AND2 (N9860, N9856, N6278);
buf BUF1 (N9861, N9849);
xor XOR2 (N9862, N9857, N3869);
nand NAND2 (N9863, N9852, N8062);
and AND4 (N9864, N9863, N2581, N4379, N479);
nor NOR2 (N9865, N9859, N7136);
nor NOR2 (N9866, N9861, N2987);
xor XOR2 (N9867, N9866, N1503);
not NOT1 (N9868, N9865);
xor XOR2 (N9869, N9855, N8268);
nor NOR2 (N9870, N9860, N7916);
not NOT1 (N9871, N9867);
nor NOR4 (N9872, N9848, N8265, N2549, N8223);
nor NOR2 (N9873, N9869, N3252);
buf BUF1 (N9874, N9871);
buf BUF1 (N9875, N9862);
not NOT1 (N9876, N9874);
not NOT1 (N9877, N9868);
and AND3 (N9878, N9870, N4570, N1654);
or OR2 (N9879, N9877, N2861);
or OR2 (N9880, N9875, N130);
xor XOR2 (N9881, N9876, N1321);
or OR3 (N9882, N9820, N2534, N1258);
buf BUF1 (N9883, N9882);
xor XOR2 (N9884, N9879, N6397);
not NOT1 (N9885, N9883);
nor NOR3 (N9886, N9873, N1834, N451);
not NOT1 (N9887, N9878);
and AND4 (N9888, N9864, N3847, N5997, N4661);
buf BUF1 (N9889, N9853);
or OR4 (N9890, N9887, N1528, N7126, N8054);
nor NOR3 (N9891, N9884, N756, N2566);
buf BUF1 (N9892, N9891);
buf BUF1 (N9893, N9885);
nand NAND3 (N9894, N9872, N4770, N9502);
or OR3 (N9895, N9890, N3526, N7802);
buf BUF1 (N9896, N9894);
or OR3 (N9897, N9881, N3191, N4774);
buf BUF1 (N9898, N9886);
not NOT1 (N9899, N9895);
or OR4 (N9900, N9896, N9400, N5504, N8666);
nor NOR3 (N9901, N9893, N303, N5443);
nor NOR2 (N9902, N9880, N5334);
nor NOR2 (N9903, N9902, N6748);
xor XOR2 (N9904, N9892, N722);
xor XOR2 (N9905, N9839, N6438);
nor NOR3 (N9906, N9904, N749, N5464);
nand NAND4 (N9907, N9889, N9740, N6708, N2168);
or OR3 (N9908, N9888, N6866, N8293);
not NOT1 (N9909, N9898);
nand NAND2 (N9910, N9900, N7353);
nand NAND3 (N9911, N9910, N3472, N9813);
not NOT1 (N9912, N9903);
or OR3 (N9913, N9912, N4579, N8550);
xor XOR2 (N9914, N9901, N8048);
and AND4 (N9915, N9899, N2237, N219, N5152);
buf BUF1 (N9916, N9911);
or OR3 (N9917, N9916, N7938, N9047);
or OR4 (N9918, N9905, N4071, N8793, N7226);
not NOT1 (N9919, N9897);
and AND2 (N9920, N9913, N2742);
nor NOR2 (N9921, N9915, N6033);
or OR2 (N9922, N9921, N7046);
buf BUF1 (N9923, N9906);
nand NAND4 (N9924, N9918, N3686, N4128, N557);
or OR4 (N9925, N9907, N6278, N9672, N6084);
not NOT1 (N9926, N9924);
or OR4 (N9927, N9917, N3677, N3361, N8336);
or OR2 (N9928, N9923, N9541);
not NOT1 (N9929, N9925);
or OR3 (N9930, N9927, N7422, N2774);
xor XOR2 (N9931, N9929, N9276);
or OR4 (N9932, N9930, N5568, N6525, N1200);
not NOT1 (N9933, N9932);
and AND3 (N9934, N9922, N1758, N8451);
buf BUF1 (N9935, N9920);
not NOT1 (N9936, N9919);
buf BUF1 (N9937, N9935);
nor NOR4 (N9938, N9931, N614, N248, N9324);
nor NOR3 (N9939, N9934, N9085, N9750);
nand NAND3 (N9940, N9914, N5753, N6659);
nand NAND2 (N9941, N9937, N594);
nand NAND4 (N9942, N9939, N4741, N1820, N2012);
or OR2 (N9943, N9933, N3591);
nor NOR4 (N9944, N9909, N1979, N7502, N6288);
xor XOR2 (N9945, N9908, N1336);
and AND2 (N9946, N9936, N7293);
and AND2 (N9947, N9943, N2022);
nor NOR3 (N9948, N9945, N1471, N7060);
not NOT1 (N9949, N9940);
and AND2 (N9950, N9938, N2688);
buf BUF1 (N9951, N9944);
nor NOR3 (N9952, N9948, N3151, N3233);
and AND2 (N9953, N9947, N1039);
or OR2 (N9954, N9950, N5354);
xor XOR2 (N9955, N9949, N3968);
and AND3 (N9956, N9952, N3978, N3327);
buf BUF1 (N9957, N9941);
nor NOR2 (N9958, N9942, N1543);
and AND2 (N9959, N9946, N5147);
buf BUF1 (N9960, N9954);
nand NAND4 (N9961, N9958, N9630, N8564, N3221);
xor XOR2 (N9962, N9928, N8555);
or OR4 (N9963, N9955, N2352, N8625, N532);
xor XOR2 (N9964, N9953, N3179);
or OR4 (N9965, N9959, N6816, N1082, N5607);
buf BUF1 (N9966, N9961);
buf BUF1 (N9967, N9963);
buf BUF1 (N9968, N9957);
buf BUF1 (N9969, N9967);
not NOT1 (N9970, N9965);
buf BUF1 (N9971, N9956);
xor XOR2 (N9972, N9962, N5903);
buf BUF1 (N9973, N9972);
buf BUF1 (N9974, N9951);
nand NAND3 (N9975, N9970, N9919, N8191);
nor NOR2 (N9976, N9926, N103);
nand NAND2 (N9977, N9966, N2382);
and AND4 (N9978, N9960, N9849, N4176, N4069);
nand NAND3 (N9979, N9977, N564, N2433);
xor XOR2 (N9980, N9969, N9627);
and AND3 (N9981, N9968, N6481, N3204);
nand NAND4 (N9982, N9981, N3515, N8606, N2828);
nor NOR3 (N9983, N9982, N7373, N6467);
not NOT1 (N9984, N9983);
buf BUF1 (N9985, N9971);
nor NOR3 (N9986, N9975, N9218, N6445);
nand NAND2 (N9987, N9976, N954);
xor XOR2 (N9988, N9985, N9307);
nor NOR4 (N9989, N9987, N7205, N6854, N2897);
not NOT1 (N9990, N9973);
not NOT1 (N9991, N9984);
buf BUF1 (N9992, N9991);
xor XOR2 (N9993, N9979, N4841);
nor NOR3 (N9994, N9964, N1350, N5168);
or OR3 (N9995, N9994, N6382, N4514);
or OR4 (N9996, N9989, N7806, N4101, N7757);
and AND2 (N9997, N9986, N2165);
nor NOR3 (N9998, N9974, N8695, N2971);
or OR2 (N9999, N9990, N8179);
xor XOR2 (N10000, N9996, N5288);
buf BUF1 (N10001, N9998);
nand NAND3 (N10002, N10001, N6582, N3318);
nor NOR3 (N10003, N9992, N3749, N7477);
nor NOR4 (N10004, N9997, N3534, N6943, N7883);
buf BUF1 (N10005, N9999);
not NOT1 (N10006, N10004);
or OR3 (N10007, N9995, N1747, N6209);
and AND2 (N10008, N9980, N9399);
xor XOR2 (N10009, N10006, N2001);
and AND2 (N10010, N9993, N8810);
nand NAND2 (N10011, N10002, N5451);
or OR2 (N10012, N10011, N9921);
and AND4 (N10013, N10007, N4922, N2634, N8468);
or OR4 (N10014, N10008, N7385, N7457, N530);
not NOT1 (N10015, N9978);
nor NOR4 (N10016, N10005, N645, N717, N9633);
xor XOR2 (N10017, N10009, N8748);
xor XOR2 (N10018, N10013, N1045);
not NOT1 (N10019, N10014);
not NOT1 (N10020, N10000);
or OR4 (N10021, N10019, N2265, N7963, N2579);
xor XOR2 (N10022, N10018, N3885);
or OR2 (N10023, N10017, N4607);
nand NAND2 (N10024, N10003, N7447);
and AND2 (N10025, N10015, N3266);
buf BUF1 (N10026, N10024);
not NOT1 (N10027, N9988);
or OR2 (N10028, N10027, N5249);
nor NOR4 (N10029, N10025, N3711, N6212, N1481);
or OR4 (N10030, N10022, N3005, N9853, N8692);
nor NOR2 (N10031, N10030, N9116);
buf BUF1 (N10032, N10029);
nor NOR3 (N10033, N10010, N9382, N9163);
xor XOR2 (N10034, N10031, N3437);
not NOT1 (N10035, N10028);
nand NAND2 (N10036, N10023, N3229);
or OR2 (N10037, N10036, N3396);
nand NAND2 (N10038, N10026, N908);
xor XOR2 (N10039, N10020, N5367);
buf BUF1 (N10040, N10033);
not NOT1 (N10041, N10035);
or OR2 (N10042, N10034, N2225);
xor XOR2 (N10043, N10038, N6526);
or OR4 (N10044, N10032, N2787, N3103, N8381);
buf BUF1 (N10045, N10040);
xor XOR2 (N10046, N10021, N6265);
xor XOR2 (N10047, N10045, N4989);
or OR4 (N10048, N10042, N4884, N2708, N9484);
xor XOR2 (N10049, N10037, N2640);
xor XOR2 (N10050, N10041, N2367);
and AND4 (N10051, N10046, N4903, N7569, N1682);
or OR2 (N10052, N10016, N5263);
buf BUF1 (N10053, N10012);
or OR4 (N10054, N10050, N5232, N3081, N7811);
and AND2 (N10055, N10052, N7428);
and AND2 (N10056, N10051, N8051);
not NOT1 (N10057, N10048);
nand NAND2 (N10058, N10057, N2482);
and AND2 (N10059, N10055, N5310);
not NOT1 (N10060, N10059);
not NOT1 (N10061, N10044);
not NOT1 (N10062, N10056);
xor XOR2 (N10063, N10049, N7824);
not NOT1 (N10064, N10054);
or OR3 (N10065, N10043, N6871, N8125);
nor NOR2 (N10066, N10047, N2261);
nand NAND4 (N10067, N10062, N1775, N2604, N5490);
or OR2 (N10068, N10063, N4599);
or OR2 (N10069, N10058, N7789);
or OR3 (N10070, N10065, N5228, N7361);
xor XOR2 (N10071, N10068, N1308);
not NOT1 (N10072, N10066);
buf BUF1 (N10073, N10039);
buf BUF1 (N10074, N10070);
and AND3 (N10075, N10072, N2684, N8194);
and AND4 (N10076, N10067, N9837, N312, N2771);
buf BUF1 (N10077, N10071);
not NOT1 (N10078, N10060);
xor XOR2 (N10079, N10076, N5443);
and AND4 (N10080, N10073, N5023, N2209, N7276);
and AND4 (N10081, N10080, N3194, N1833, N7166);
nor NOR2 (N10082, N10077, N9241);
nand NAND4 (N10083, N10064, N7881, N4579, N1286);
not NOT1 (N10084, N10074);
xor XOR2 (N10085, N10084, N5519);
xor XOR2 (N10086, N10061, N3458);
nand NAND3 (N10087, N10083, N7509, N1446);
xor XOR2 (N10088, N10085, N7725);
nand NAND3 (N10089, N10082, N9221, N5309);
nor NOR3 (N10090, N10078, N3083, N3586);
not NOT1 (N10091, N10088);
xor XOR2 (N10092, N10087, N1887);
xor XOR2 (N10093, N10079, N3531);
or OR3 (N10094, N10053, N1839, N7271);
or OR4 (N10095, N10092, N2576, N3860, N1910);
xor XOR2 (N10096, N10090, N9132);
or OR4 (N10097, N10086, N9821, N9268, N4494);
nand NAND4 (N10098, N10089, N7221, N3026, N6552);
nor NOR3 (N10099, N10094, N8602, N3062);
not NOT1 (N10100, N10095);
xor XOR2 (N10101, N10081, N166);
or OR4 (N10102, N10091, N7010, N1603, N833);
not NOT1 (N10103, N10093);
or OR2 (N10104, N10069, N5341);
buf BUF1 (N10105, N10075);
nor NOR2 (N10106, N10096, N4184);
and AND2 (N10107, N10098, N3090);
not NOT1 (N10108, N10103);
nor NOR3 (N10109, N10107, N9346, N3772);
nor NOR2 (N10110, N10097, N5047);
buf BUF1 (N10111, N10104);
or OR2 (N10112, N10100, N4433);
nor NOR4 (N10113, N10112, N8455, N1577, N3333);
xor XOR2 (N10114, N10106, N3557);
nand NAND3 (N10115, N10105, N1567, N9240);
nand NAND3 (N10116, N10108, N6313, N3693);
buf BUF1 (N10117, N10111);
not NOT1 (N10118, N10117);
nor NOR3 (N10119, N10114, N4603, N5832);
nor NOR4 (N10120, N10119, N1976, N7516, N3733);
nand NAND2 (N10121, N10116, N572);
buf BUF1 (N10122, N10110);
xor XOR2 (N10123, N10122, N1575);
or OR3 (N10124, N10109, N5477, N441);
buf BUF1 (N10125, N10115);
nand NAND2 (N10126, N10125, N5372);
and AND2 (N10127, N10101, N2441);
not NOT1 (N10128, N10124);
xor XOR2 (N10129, N10113, N3810);
or OR2 (N10130, N10128, N2511);
or OR3 (N10131, N10121, N3872, N6388);
nand NAND2 (N10132, N10102, N4247);
nor NOR2 (N10133, N10123, N767);
not NOT1 (N10134, N10129);
xor XOR2 (N10135, N10126, N126);
and AND3 (N10136, N10135, N4269, N4904);
and AND4 (N10137, N10127, N740, N9675, N1411);
buf BUF1 (N10138, N10130);
or OR3 (N10139, N10136, N670, N1050);
or OR4 (N10140, N10118, N2288, N961, N7841);
not NOT1 (N10141, N10133);
buf BUF1 (N10142, N10139);
or OR3 (N10143, N10137, N4001, N437);
or OR2 (N10144, N10143, N4456);
xor XOR2 (N10145, N10131, N8087);
xor XOR2 (N10146, N10141, N4289);
not NOT1 (N10147, N10134);
not NOT1 (N10148, N10146);
not NOT1 (N10149, N10132);
nor NOR2 (N10150, N10148, N2226);
nor NOR4 (N10151, N10144, N2794, N149, N5649);
and AND3 (N10152, N10142, N4212, N3304);
nand NAND4 (N10153, N10152, N4577, N7950, N8259);
buf BUF1 (N10154, N10151);
and AND2 (N10155, N10154, N4303);
or OR3 (N10156, N10145, N8075, N4686);
xor XOR2 (N10157, N10149, N3498);
and AND3 (N10158, N10157, N4586, N7491);
buf BUF1 (N10159, N10150);
buf BUF1 (N10160, N10158);
buf BUF1 (N10161, N10140);
or OR2 (N10162, N10138, N5123);
nand NAND3 (N10163, N10162, N7968, N5696);
and AND2 (N10164, N10153, N9463);
not NOT1 (N10165, N10161);
nand NAND4 (N10166, N10155, N1231, N4253, N5621);
not NOT1 (N10167, N10159);
or OR3 (N10168, N10147, N1899, N8779);
xor XOR2 (N10169, N10167, N5097);
not NOT1 (N10170, N10160);
or OR4 (N10171, N10166, N9529, N4454, N934);
nand NAND2 (N10172, N10163, N4913);
and AND4 (N10173, N10165, N8295, N1966, N1640);
or OR3 (N10174, N10120, N1412, N3332);
nand NAND4 (N10175, N10164, N4169, N4000, N6162);
not NOT1 (N10176, N10172);
buf BUF1 (N10177, N10156);
and AND2 (N10178, N10169, N3832);
nand NAND3 (N10179, N10177, N9166, N8108);
not NOT1 (N10180, N10173);
and AND4 (N10181, N10174, N6858, N1284, N9260);
not NOT1 (N10182, N10099);
nand NAND4 (N10183, N10179, N7277, N8528, N1698);
or OR4 (N10184, N10168, N3030, N9375, N10008);
buf BUF1 (N10185, N10182);
not NOT1 (N10186, N10184);
nand NAND4 (N10187, N10171, N3592, N3100, N8994);
buf BUF1 (N10188, N10185);
xor XOR2 (N10189, N10176, N4310);
and AND3 (N10190, N10188, N7393, N9219);
buf BUF1 (N10191, N10190);
xor XOR2 (N10192, N10189, N3570);
and AND4 (N10193, N10180, N456, N803, N9170);
not NOT1 (N10194, N10187);
nand NAND3 (N10195, N10175, N5429, N8400);
nand NAND2 (N10196, N10195, N4219);
not NOT1 (N10197, N10191);
not NOT1 (N10198, N10196);
or OR4 (N10199, N10198, N5797, N659, N2285);
buf BUF1 (N10200, N10183);
or OR4 (N10201, N10193, N3785, N10089, N7459);
not NOT1 (N10202, N10197);
or OR3 (N10203, N10202, N6095, N5829);
xor XOR2 (N10204, N10201, N7761);
not NOT1 (N10205, N10194);
not NOT1 (N10206, N10200);
nand NAND3 (N10207, N10203, N1416, N3949);
xor XOR2 (N10208, N10192, N1967);
and AND2 (N10209, N10181, N9440);
nor NOR2 (N10210, N10178, N7198);
and AND2 (N10211, N10210, N6193);
xor XOR2 (N10212, N10186, N9878);
nand NAND3 (N10213, N10211, N935, N9703);
buf BUF1 (N10214, N10212);
nand NAND4 (N10215, N10204, N9071, N8509, N6189);
xor XOR2 (N10216, N10205, N3453);
nand NAND2 (N10217, N10209, N4567);
buf BUF1 (N10218, N10214);
buf BUF1 (N10219, N10207);
nand NAND4 (N10220, N10219, N2029, N3199, N9573);
or OR4 (N10221, N10170, N8919, N1565, N1692);
xor XOR2 (N10222, N10199, N1271);
nor NOR4 (N10223, N10216, N4740, N551, N3354);
nor NOR3 (N10224, N10221, N7479, N5316);
nor NOR3 (N10225, N10220, N2497, N9239);
not NOT1 (N10226, N10208);
and AND2 (N10227, N10225, N6176);
buf BUF1 (N10228, N10226);
nor NOR2 (N10229, N10222, N3739);
or OR2 (N10230, N10224, N1358);
or OR2 (N10231, N10217, N10058);
or OR2 (N10232, N10231, N345);
or OR3 (N10233, N10213, N5991, N9605);
and AND3 (N10234, N10229, N1152, N5407);
xor XOR2 (N10235, N10227, N5295);
not NOT1 (N10236, N10230);
or OR4 (N10237, N10232, N7861, N10067, N8242);
xor XOR2 (N10238, N10236, N8195);
and AND2 (N10239, N10228, N7191);
xor XOR2 (N10240, N10223, N5620);
nand NAND4 (N10241, N10239, N5981, N7565, N10029);
nand NAND2 (N10242, N10240, N2200);
or OR4 (N10243, N10206, N7560, N2382, N2732);
nand NAND2 (N10244, N10243, N10238);
and AND2 (N10245, N7802, N8089);
buf BUF1 (N10246, N10237);
xor XOR2 (N10247, N10242, N1049);
not NOT1 (N10248, N10241);
buf BUF1 (N10249, N10234);
or OR4 (N10250, N10246, N5275, N2120, N180);
and AND4 (N10251, N10245, N2438, N7004, N5886);
not NOT1 (N10252, N10248);
and AND3 (N10253, N10247, N434, N795);
or OR2 (N10254, N10218, N1064);
not NOT1 (N10255, N10253);
nor NOR3 (N10256, N10254, N7481, N780);
nor NOR2 (N10257, N10251, N3028);
or OR2 (N10258, N10244, N569);
nand NAND3 (N10259, N10257, N676, N8711);
nand NAND3 (N10260, N10256, N5173, N4462);
not NOT1 (N10261, N10233);
or OR3 (N10262, N10259, N5681, N7359);
not NOT1 (N10263, N10262);
nor NOR3 (N10264, N10235, N3472, N550);
buf BUF1 (N10265, N10255);
xor XOR2 (N10266, N10250, N718);
xor XOR2 (N10267, N10264, N6693);
not NOT1 (N10268, N10263);
not NOT1 (N10269, N10265);
or OR2 (N10270, N10215, N5078);
and AND3 (N10271, N10268, N8515, N9750);
xor XOR2 (N10272, N10261, N2312);
and AND2 (N10273, N10266, N4733);
nor NOR2 (N10274, N10252, N7322);
xor XOR2 (N10275, N10249, N9727);
nand NAND3 (N10276, N10271, N5745, N1184);
not NOT1 (N10277, N10274);
not NOT1 (N10278, N10267);
not NOT1 (N10279, N10270);
xor XOR2 (N10280, N10272, N6831);
and AND4 (N10281, N10258, N1350, N5513, N122);
nor NOR2 (N10282, N10278, N4074);
buf BUF1 (N10283, N10269);
nand NAND2 (N10284, N10277, N3707);
or OR2 (N10285, N10283, N149);
and AND4 (N10286, N10282, N2745, N1398, N7057);
xor XOR2 (N10287, N10280, N1530);
nor NOR3 (N10288, N10275, N944, N8230);
nor NOR2 (N10289, N10284, N3993);
buf BUF1 (N10290, N10287);
nor NOR2 (N10291, N10279, N2986);
buf BUF1 (N10292, N10291);
xor XOR2 (N10293, N10289, N8827);
nand NAND4 (N10294, N10288, N7456, N6382, N3485);
buf BUF1 (N10295, N10285);
not NOT1 (N10296, N10276);
not NOT1 (N10297, N10273);
and AND2 (N10298, N10294, N5188);
or OR3 (N10299, N10297, N8985, N7788);
or OR2 (N10300, N10260, N3641);
nor NOR2 (N10301, N10299, N10042);
nor NOR4 (N10302, N10298, N6573, N4837, N3524);
buf BUF1 (N10303, N10300);
nor NOR2 (N10304, N10292, N7871);
not NOT1 (N10305, N10281);
xor XOR2 (N10306, N10304, N8452);
and AND3 (N10307, N10305, N8892, N395);
xor XOR2 (N10308, N10293, N2958);
nor NOR3 (N10309, N10303, N8425, N4514);
not NOT1 (N10310, N10301);
and AND2 (N10311, N10308, N8511);
xor XOR2 (N10312, N10286, N23);
nand NAND4 (N10313, N10312, N5820, N8848, N5999);
xor XOR2 (N10314, N10306, N4142);
not NOT1 (N10315, N10314);
nor NOR4 (N10316, N10295, N6263, N8651, N6927);
or OR3 (N10317, N10315, N940, N1540);
and AND4 (N10318, N10316, N10155, N4407, N5936);
and AND2 (N10319, N10310, N9361);
not NOT1 (N10320, N10302);
or OR3 (N10321, N10311, N2554, N10047);
nor NOR2 (N10322, N10318, N2344);
nand NAND2 (N10323, N10290, N9812);
nand NAND3 (N10324, N10323, N4342, N7496);
buf BUF1 (N10325, N10324);
nand NAND2 (N10326, N10307, N9000);
nor NOR3 (N10327, N10313, N10104, N10131);
xor XOR2 (N10328, N10296, N3231);
xor XOR2 (N10329, N10319, N2256);
xor XOR2 (N10330, N10321, N9853);
not NOT1 (N10331, N10325);
or OR4 (N10332, N10328, N3854, N5740, N4284);
or OR3 (N10333, N10317, N8694, N6502);
and AND3 (N10334, N10322, N5378, N5370);
not NOT1 (N10335, N10331);
nor NOR4 (N10336, N10335, N5405, N1522, N2193);
not NOT1 (N10337, N10327);
buf BUF1 (N10338, N10336);
and AND2 (N10339, N10334, N4471);
buf BUF1 (N10340, N10339);
nand NAND4 (N10341, N10340, N180, N6650, N657);
and AND4 (N10342, N10326, N2966, N9838, N764);
not NOT1 (N10343, N10309);
buf BUF1 (N10344, N10342);
or OR2 (N10345, N10337, N1303);
xor XOR2 (N10346, N10330, N8425);
nand NAND4 (N10347, N10345, N2516, N8947, N6956);
nand NAND4 (N10348, N10343, N5060, N1725, N5070);
nand NAND2 (N10349, N10347, N9019);
nand NAND3 (N10350, N10332, N2295, N9664);
or OR4 (N10351, N10329, N604, N5850, N5063);
xor XOR2 (N10352, N10351, N1070);
and AND4 (N10353, N10346, N571, N4069, N10005);
and AND4 (N10354, N10352, N2872, N7624, N8390);
or OR3 (N10355, N10354, N7648, N7784);
and AND4 (N10356, N10338, N4709, N4436, N7733);
buf BUF1 (N10357, N10356);
not NOT1 (N10358, N10349);
nand NAND4 (N10359, N10348, N8537, N1118, N6208);
or OR4 (N10360, N10350, N6742, N2693, N10035);
nor NOR3 (N10361, N10355, N10209, N4158);
xor XOR2 (N10362, N10358, N2527);
buf BUF1 (N10363, N10357);
and AND3 (N10364, N10362, N6635, N1794);
or OR3 (N10365, N10353, N10314, N7767);
not NOT1 (N10366, N10344);
and AND4 (N10367, N10366, N3836, N5044, N6894);
nor NOR3 (N10368, N10364, N543, N3356);
buf BUF1 (N10369, N10365);
not NOT1 (N10370, N10368);
nand NAND2 (N10371, N10320, N294);
buf BUF1 (N10372, N10370);
and AND2 (N10373, N10360, N2855);
xor XOR2 (N10374, N10341, N1783);
xor XOR2 (N10375, N10333, N1262);
nor NOR2 (N10376, N10372, N8139);
nor NOR4 (N10377, N10363, N7601, N7325, N1510);
nor NOR3 (N10378, N10369, N1331, N7362);
xor XOR2 (N10379, N10371, N7631);
xor XOR2 (N10380, N10378, N1585);
xor XOR2 (N10381, N10379, N4943);
and AND2 (N10382, N10381, N7356);
or OR2 (N10383, N10374, N7627);
nor NOR4 (N10384, N10380, N3014, N1852, N7112);
and AND2 (N10385, N10375, N520);
not NOT1 (N10386, N10377);
and AND3 (N10387, N10367, N4081, N927);
or OR4 (N10388, N10361, N1675, N5981, N548);
nor NOR4 (N10389, N10384, N3224, N5911, N6761);
and AND3 (N10390, N10376, N2717, N480);
buf BUF1 (N10391, N10386);
nand NAND3 (N10392, N10383, N2825, N9488);
or OR3 (N10393, N10385, N3463, N9132);
or OR4 (N10394, N10382, N10377, N3859, N5151);
nand NAND4 (N10395, N10388, N7444, N7021, N5693);
nor NOR4 (N10396, N10390, N1858, N1544, N5133);
nor NOR3 (N10397, N10359, N1807, N9339);
not NOT1 (N10398, N10397);
buf BUF1 (N10399, N10394);
and AND3 (N10400, N10373, N6650, N3528);
xor XOR2 (N10401, N10395, N7324);
not NOT1 (N10402, N10389);
nand NAND4 (N10403, N10391, N9536, N346, N2048);
and AND2 (N10404, N10403, N6743);
nor NOR2 (N10405, N10387, N5905);
not NOT1 (N10406, N10392);
nor NOR2 (N10407, N10401, N9109);
buf BUF1 (N10408, N10396);
not NOT1 (N10409, N10408);
or OR2 (N10410, N10404, N5442);
or OR4 (N10411, N10393, N510, N1234, N4809);
and AND2 (N10412, N10400, N4303);
and AND3 (N10413, N10405, N6885, N5360);
nor NOR4 (N10414, N10409, N69, N1402, N358);
not NOT1 (N10415, N10411);
buf BUF1 (N10416, N10407);
nand NAND2 (N10417, N10402, N4863);
and AND2 (N10418, N10414, N1426);
or OR4 (N10419, N10410, N8782, N2233, N10352);
nor NOR3 (N10420, N10417, N4076, N296);
buf BUF1 (N10421, N10416);
nor NOR4 (N10422, N10418, N363, N3023, N5434);
or OR3 (N10423, N10399, N1664, N3761);
xor XOR2 (N10424, N10413, N2051);
xor XOR2 (N10425, N10423, N4590);
buf BUF1 (N10426, N10420);
not NOT1 (N10427, N10422);
not NOT1 (N10428, N10424);
nor NOR4 (N10429, N10427, N3780, N2746, N5343);
buf BUF1 (N10430, N10428);
nor NOR3 (N10431, N10430, N3274, N1666);
or OR4 (N10432, N10415, N7881, N6511, N127);
or OR4 (N10433, N10429, N122, N5, N5791);
nand NAND2 (N10434, N10425, N10376);
nor NOR2 (N10435, N10434, N4602);
and AND3 (N10436, N10431, N411, N6966);
buf BUF1 (N10437, N10419);
nand NAND2 (N10438, N10406, N9595);
or OR3 (N10439, N10412, N4195, N5675);
xor XOR2 (N10440, N10438, N3748);
xor XOR2 (N10441, N10440, N3701);
or OR2 (N10442, N10437, N1398);
nor NOR4 (N10443, N10439, N5112, N8806, N9854);
xor XOR2 (N10444, N10436, N1918);
xor XOR2 (N10445, N10443, N6968);
not NOT1 (N10446, N10398);
buf BUF1 (N10447, N10432);
or OR3 (N10448, N10426, N9033, N6360);
nand NAND2 (N10449, N10445, N3750);
nor NOR2 (N10450, N10421, N5671);
or OR4 (N10451, N10433, N918, N4995, N5618);
and AND4 (N10452, N10441, N4936, N7204, N9208);
xor XOR2 (N10453, N10442, N4676);
and AND2 (N10454, N10453, N2641);
or OR2 (N10455, N10452, N10357);
buf BUF1 (N10456, N10450);
xor XOR2 (N10457, N10447, N9994);
xor XOR2 (N10458, N10454, N5952);
and AND3 (N10459, N10451, N48, N969);
buf BUF1 (N10460, N10446);
or OR4 (N10461, N10448, N587, N2194, N5747);
not NOT1 (N10462, N10435);
xor XOR2 (N10463, N10461, N2832);
and AND4 (N10464, N10463, N5889, N3971, N9937);
xor XOR2 (N10465, N10458, N4468);
buf BUF1 (N10466, N10459);
xor XOR2 (N10467, N10444, N8857);
or OR2 (N10468, N10460, N9277);
nor NOR3 (N10469, N10466, N9402, N4178);
nand NAND2 (N10470, N10467, N797);
nor NOR3 (N10471, N10465, N109, N2275);
xor XOR2 (N10472, N10464, N5288);
xor XOR2 (N10473, N10471, N1162);
not NOT1 (N10474, N10449);
xor XOR2 (N10475, N10472, N6952);
nor NOR4 (N10476, N10468, N6170, N8678, N7128);
or OR3 (N10477, N10470, N6549, N4683);
or OR2 (N10478, N10455, N7116);
buf BUF1 (N10479, N10478);
xor XOR2 (N10480, N10477, N9358);
and AND3 (N10481, N10462, N2016, N900);
not NOT1 (N10482, N10456);
nor NOR2 (N10483, N10480, N8545);
or OR3 (N10484, N10476, N5334, N5617);
nand NAND3 (N10485, N10469, N5693, N6039);
nor NOR2 (N10486, N10475, N7162);
xor XOR2 (N10487, N10481, N2142);
xor XOR2 (N10488, N10479, N1239);
or OR4 (N10489, N10486, N6919, N9837, N5985);
xor XOR2 (N10490, N10483, N4582);
and AND2 (N10491, N10489, N8829);
or OR3 (N10492, N10484, N9128, N5585);
buf BUF1 (N10493, N10487);
not NOT1 (N10494, N10457);
buf BUF1 (N10495, N10485);
not NOT1 (N10496, N10474);
xor XOR2 (N10497, N10495, N1953);
buf BUF1 (N10498, N10492);
not NOT1 (N10499, N10498);
nor NOR2 (N10500, N10494, N6480);
buf BUF1 (N10501, N10473);
xor XOR2 (N10502, N10488, N1604);
not NOT1 (N10503, N10490);
buf BUF1 (N10504, N10496);
and AND2 (N10505, N10493, N353);
buf BUF1 (N10506, N10491);
or OR4 (N10507, N10504, N1719, N3056, N4023);
nor NOR3 (N10508, N10503, N6851, N2525);
not NOT1 (N10509, N10508);
nand NAND4 (N10510, N10482, N3488, N261, N6395);
nand NAND3 (N10511, N10501, N6998, N2632);
xor XOR2 (N10512, N10510, N2115);
nand NAND3 (N10513, N10497, N10076, N5796);
or OR3 (N10514, N10505, N10463, N3575);
buf BUF1 (N10515, N10513);
and AND2 (N10516, N10511, N911);
and AND4 (N10517, N10516, N4587, N385, N9402);
and AND4 (N10518, N10507, N10307, N3303, N8600);
xor XOR2 (N10519, N10512, N5424);
and AND2 (N10520, N10499, N9139);
or OR2 (N10521, N10520, N3914);
or OR3 (N10522, N10509, N4018, N2072);
buf BUF1 (N10523, N10522);
buf BUF1 (N10524, N10515);
nand NAND2 (N10525, N10502, N25);
nor NOR4 (N10526, N10500, N5504, N1813, N3180);
not NOT1 (N10527, N10523);
xor XOR2 (N10528, N10526, N4400);
xor XOR2 (N10529, N10517, N4499);
xor XOR2 (N10530, N10519, N4177);
nand NAND2 (N10531, N10514, N2688);
or OR2 (N10532, N10524, N2602);
xor XOR2 (N10533, N10527, N5128);
not NOT1 (N10534, N10506);
nor NOR4 (N10535, N10533, N8133, N7300, N2299);
not NOT1 (N10536, N10521);
xor XOR2 (N10537, N10536, N4009);
and AND3 (N10538, N10525, N4492, N179);
nand NAND4 (N10539, N10537, N2777, N1350, N6161);
buf BUF1 (N10540, N10538);
xor XOR2 (N10541, N10540, N59);
nor NOR3 (N10542, N10534, N2298, N10237);
or OR4 (N10543, N10518, N9743, N1775, N2673);
or OR2 (N10544, N10529, N7182);
buf BUF1 (N10545, N10543);
buf BUF1 (N10546, N10528);
xor XOR2 (N10547, N10541, N9317);
or OR2 (N10548, N10547, N6449);
nor NOR3 (N10549, N10539, N6841, N9500);
and AND3 (N10550, N10548, N4971, N6758);
xor XOR2 (N10551, N10549, N9745);
not NOT1 (N10552, N10546);
not NOT1 (N10553, N10544);
or OR3 (N10554, N10545, N1880, N5193);
buf BUF1 (N10555, N10553);
buf BUF1 (N10556, N10531);
buf BUF1 (N10557, N10542);
buf BUF1 (N10558, N10551);
buf BUF1 (N10559, N10558);
and AND2 (N10560, N10557, N6751);
or OR4 (N10561, N10559, N4749, N3393, N6553);
and AND3 (N10562, N10554, N2685, N3674);
not NOT1 (N10563, N10555);
xor XOR2 (N10564, N10560, N3947);
nand NAND3 (N10565, N10532, N9060, N9947);
nor NOR2 (N10566, N10561, N5566);
xor XOR2 (N10567, N10564, N4841);
xor XOR2 (N10568, N10567, N6908);
xor XOR2 (N10569, N10565, N9919);
not NOT1 (N10570, N10568);
and AND2 (N10571, N10570, N5495);
nand NAND3 (N10572, N10535, N8862, N7534);
not NOT1 (N10573, N10550);
nor NOR4 (N10574, N10552, N3497, N5069, N5100);
or OR2 (N10575, N10530, N834);
and AND2 (N10576, N10572, N810);
buf BUF1 (N10577, N10573);
xor XOR2 (N10578, N10577, N1332);
and AND4 (N10579, N10556, N929, N8470, N5401);
nor NOR2 (N10580, N10562, N5232);
xor XOR2 (N10581, N10580, N3398);
and AND3 (N10582, N10571, N4817, N5021);
xor XOR2 (N10583, N10563, N4710);
or OR2 (N10584, N10576, N9907);
or OR4 (N10585, N10575, N4581, N2350, N5241);
not NOT1 (N10586, N10581);
and AND3 (N10587, N10582, N5534, N3890);
not NOT1 (N10588, N10574);
and AND4 (N10589, N10578, N8195, N2248, N6033);
not NOT1 (N10590, N10585);
xor XOR2 (N10591, N10584, N3932);
nor NOR3 (N10592, N10587, N7377, N97);
buf BUF1 (N10593, N10579);
not NOT1 (N10594, N10593);
xor XOR2 (N10595, N10583, N1276);
nor NOR2 (N10596, N10594, N3296);
and AND4 (N10597, N10589, N8494, N1418, N1885);
nor NOR2 (N10598, N10590, N5770);
nand NAND4 (N10599, N10595, N7380, N10149, N1897);
not NOT1 (N10600, N10599);
and AND2 (N10601, N10566, N5206);
nand NAND3 (N10602, N10592, N9939, N6908);
nand NAND4 (N10603, N10586, N9617, N7444, N1912);
or OR2 (N10604, N10591, N992);
not NOT1 (N10605, N10602);
buf BUF1 (N10606, N10604);
or OR3 (N10607, N10600, N6609, N5683);
xor XOR2 (N10608, N10588, N5673);
and AND3 (N10609, N10597, N3101, N8790);
nor NOR4 (N10610, N10609, N2843, N7077, N215);
buf BUF1 (N10611, N10605);
xor XOR2 (N10612, N10611, N9376);
or OR4 (N10613, N10607, N1002, N213, N4737);
nor NOR4 (N10614, N10612, N7320, N917, N2919);
nor NOR2 (N10615, N10596, N2989);
or OR4 (N10616, N10569, N10077, N8884, N9951);
nor NOR3 (N10617, N10606, N7338, N6100);
xor XOR2 (N10618, N10617, N7674);
nor NOR3 (N10619, N10614, N6391, N6072);
and AND3 (N10620, N10618, N2713, N1878);
nand NAND2 (N10621, N10601, N8474);
not NOT1 (N10622, N10610);
and AND4 (N10623, N10615, N1318, N259, N1457);
and AND3 (N10624, N10621, N6486, N2941);
nor NOR2 (N10625, N10598, N2470);
xor XOR2 (N10626, N10624, N8206);
nor NOR4 (N10627, N10619, N5979, N6707, N2411);
nand NAND4 (N10628, N10626, N4100, N4020, N304);
or OR2 (N10629, N10628, N2580);
and AND2 (N10630, N10608, N2120);
xor XOR2 (N10631, N10616, N2797);
and AND2 (N10632, N10613, N3414);
or OR3 (N10633, N10603, N3354, N7319);
nand NAND4 (N10634, N10629, N7012, N855, N9191);
or OR3 (N10635, N10632, N4692, N1889);
nand NAND2 (N10636, N10631, N4547);
nand NAND4 (N10637, N10623, N2764, N5943, N8631);
or OR2 (N10638, N10636, N2062);
nor NOR3 (N10639, N10630, N9266, N9273);
nor NOR4 (N10640, N10627, N6643, N6834, N1568);
nor NOR4 (N10641, N10640, N3044, N10349, N9196);
not NOT1 (N10642, N10633);
not NOT1 (N10643, N10638);
and AND2 (N10644, N10641, N3550);
xor XOR2 (N10645, N10634, N4350);
xor XOR2 (N10646, N10644, N7035);
not NOT1 (N10647, N10622);
buf BUF1 (N10648, N10642);
not NOT1 (N10649, N10635);
and AND2 (N10650, N10647, N5641);
and AND4 (N10651, N10639, N8956, N246, N8121);
not NOT1 (N10652, N10645);
and AND4 (N10653, N10637, N9201, N1490, N6886);
not NOT1 (N10654, N10650);
nand NAND2 (N10655, N10625, N409);
xor XOR2 (N10656, N10654, N704);
not NOT1 (N10657, N10656);
nor NOR3 (N10658, N10655, N10463, N6399);
and AND4 (N10659, N10643, N8104, N3895, N6765);
or OR3 (N10660, N10652, N5487, N9759);
and AND2 (N10661, N10657, N663);
or OR3 (N10662, N10661, N3788, N8406);
not NOT1 (N10663, N10651);
and AND3 (N10664, N10653, N5857, N10054);
or OR3 (N10665, N10620, N10419, N6550);
nor NOR4 (N10666, N10662, N5297, N840, N7575);
xor XOR2 (N10667, N10648, N3908);
or OR3 (N10668, N10665, N5615, N3736);
buf BUF1 (N10669, N10659);
or OR3 (N10670, N10668, N2821, N1056);
or OR4 (N10671, N10658, N97, N6001, N9428);
not NOT1 (N10672, N10646);
nand NAND4 (N10673, N10670, N5370, N10325, N4451);
not NOT1 (N10674, N10669);
xor XOR2 (N10675, N10672, N10147);
nand NAND3 (N10676, N10667, N2247, N3483);
nor NOR3 (N10677, N10674, N4604, N9044);
buf BUF1 (N10678, N10677);
and AND4 (N10679, N10671, N2973, N1807, N2215);
nor NOR2 (N10680, N10666, N163);
not NOT1 (N10681, N10676);
nand NAND4 (N10682, N10673, N8625, N1193, N996);
and AND3 (N10683, N10679, N7698, N2950);
not NOT1 (N10684, N10681);
xor XOR2 (N10685, N10664, N9433);
buf BUF1 (N10686, N10663);
nor NOR4 (N10687, N10682, N2168, N7578, N10012);
or OR2 (N10688, N10686, N2943);
nand NAND2 (N10689, N10688, N3232);
buf BUF1 (N10690, N10683);
or OR3 (N10691, N10684, N4576, N1258);
nand NAND2 (N10692, N10649, N5850);
or OR3 (N10693, N10675, N7478, N3160);
nor NOR4 (N10694, N10689, N9623, N3875, N7220);
nor NOR2 (N10695, N10693, N5133);
buf BUF1 (N10696, N10678);
not NOT1 (N10697, N10685);
xor XOR2 (N10698, N10694, N9134);
or OR4 (N10699, N10687, N6964, N8822, N4995);
not NOT1 (N10700, N10697);
nand NAND2 (N10701, N10690, N1275);
nand NAND2 (N10702, N10660, N337);
buf BUF1 (N10703, N10701);
nand NAND2 (N10704, N10680, N10064);
xor XOR2 (N10705, N10699, N8053);
nand NAND3 (N10706, N10695, N1696, N5063);
or OR2 (N10707, N10691, N463);
nor NOR2 (N10708, N10698, N7398);
not NOT1 (N10709, N10704);
or OR2 (N10710, N10709, N7730);
and AND4 (N10711, N10708, N10546, N6935, N91);
nor NOR2 (N10712, N10692, N4055);
xor XOR2 (N10713, N10702, N1050);
buf BUF1 (N10714, N10706);
or OR2 (N10715, N10710, N9292);
buf BUF1 (N10716, N10711);
xor XOR2 (N10717, N10713, N6591);
or OR4 (N10718, N10716, N3536, N1638, N6556);
or OR4 (N10719, N10715, N9945, N9820, N8976);
and AND4 (N10720, N10707, N9810, N1839, N4733);
nand NAND3 (N10721, N10719, N6286, N2288);
nor NOR2 (N10722, N10705, N3466);
nand NAND4 (N10723, N10720, N7072, N7263, N106);
buf BUF1 (N10724, N10700);
not NOT1 (N10725, N10718);
buf BUF1 (N10726, N10703);
nor NOR2 (N10727, N10696, N6494);
or OR4 (N10728, N10724, N9653, N159, N2382);
xor XOR2 (N10729, N10725, N8813);
nor NOR3 (N10730, N10723, N2240, N5692);
nor NOR3 (N10731, N10721, N7511, N9111);
or OR4 (N10732, N10712, N4484, N8581, N639);
not NOT1 (N10733, N10731);
xor XOR2 (N10734, N10733, N5196);
buf BUF1 (N10735, N10726);
and AND2 (N10736, N10728, N9049);
xor XOR2 (N10737, N10722, N6072);
xor XOR2 (N10738, N10732, N1932);
xor XOR2 (N10739, N10737, N3869);
not NOT1 (N10740, N10717);
xor XOR2 (N10741, N10736, N2209);
nor NOR4 (N10742, N10738, N2446, N3621, N4573);
nor NOR4 (N10743, N10734, N3755, N5026, N8921);
not NOT1 (N10744, N10742);
nand NAND4 (N10745, N10735, N6369, N3931, N8935);
nand NAND3 (N10746, N10739, N2156, N172);
and AND2 (N10747, N10729, N9348);
buf BUF1 (N10748, N10744);
or OR3 (N10749, N10747, N6263, N7963);
nand NAND2 (N10750, N10749, N3851);
xor XOR2 (N10751, N10741, N5272);
nor NOR4 (N10752, N10745, N1194, N6465, N4964);
and AND3 (N10753, N10743, N7890, N2600);
and AND4 (N10754, N10748, N707, N1239, N9920);
or OR4 (N10755, N10727, N9458, N2543, N2371);
xor XOR2 (N10756, N10714, N5187);
buf BUF1 (N10757, N10756);
buf BUF1 (N10758, N10730);
and AND4 (N10759, N10758, N8298, N5282, N4575);
nand NAND2 (N10760, N10754, N5593);
nor NOR4 (N10761, N10752, N1088, N1820, N4009);
and AND4 (N10762, N10740, N6620, N4459, N6113);
and AND4 (N10763, N10751, N9519, N2196, N7038);
or OR3 (N10764, N10757, N2268, N661);
nand NAND4 (N10765, N10753, N8379, N8991, N6659);
or OR3 (N10766, N10760, N7566, N10535);
not NOT1 (N10767, N10759);
buf BUF1 (N10768, N10755);
and AND4 (N10769, N10750, N3492, N3905, N435);
buf BUF1 (N10770, N10767);
xor XOR2 (N10771, N10770, N8733);
xor XOR2 (N10772, N10763, N128);
xor XOR2 (N10773, N10764, N3987);
not NOT1 (N10774, N10766);
or OR3 (N10775, N10773, N8748, N8953);
nand NAND2 (N10776, N10774, N9854);
or OR2 (N10777, N10768, N8709);
not NOT1 (N10778, N10775);
xor XOR2 (N10779, N10771, N4556);
nand NAND3 (N10780, N10777, N6718, N10083);
and AND2 (N10781, N10776, N4649);
buf BUF1 (N10782, N10779);
or OR4 (N10783, N10761, N6786, N3788, N1890);
buf BUF1 (N10784, N10780);
buf BUF1 (N10785, N10783);
buf BUF1 (N10786, N10785);
nand NAND3 (N10787, N10772, N2784, N9988);
nor NOR4 (N10788, N10769, N10605, N5795, N10668);
nand NAND2 (N10789, N10784, N4505);
and AND4 (N10790, N10778, N2766, N5864, N3736);
not NOT1 (N10791, N10788);
not NOT1 (N10792, N10762);
or OR2 (N10793, N10787, N879);
buf BUF1 (N10794, N10789);
xor XOR2 (N10795, N10782, N238);
buf BUF1 (N10796, N10765);
not NOT1 (N10797, N10794);
xor XOR2 (N10798, N10786, N1795);
and AND3 (N10799, N10792, N8124, N2690);
and AND3 (N10800, N10790, N399, N5290);
or OR4 (N10801, N10793, N4033, N10412, N8255);
xor XOR2 (N10802, N10791, N3670);
or OR4 (N10803, N10798, N5259, N4032, N57);
not NOT1 (N10804, N10803);
or OR4 (N10805, N10746, N4058, N4891, N7112);
buf BUF1 (N10806, N10800);
xor XOR2 (N10807, N10804, N7299);
nor NOR3 (N10808, N10799, N4715, N1804);
nor NOR2 (N10809, N10807, N5099);
or OR4 (N10810, N10806, N5981, N6300, N4795);
buf BUF1 (N10811, N10797);
not NOT1 (N10812, N10801);
buf BUF1 (N10813, N10812);
or OR4 (N10814, N10795, N1205, N8537, N3923);
nor NOR4 (N10815, N10810, N2550, N10772, N6804);
or OR3 (N10816, N10813, N5652, N7655);
nor NOR3 (N10817, N10796, N794, N4228);
buf BUF1 (N10818, N10809);
or OR4 (N10819, N10816, N7910, N8711, N4602);
buf BUF1 (N10820, N10818);
not NOT1 (N10821, N10814);
not NOT1 (N10822, N10815);
or OR4 (N10823, N10817, N3771, N9209, N5085);
buf BUF1 (N10824, N10802);
or OR4 (N10825, N10822, N6341, N10732, N2172);
not NOT1 (N10826, N10824);
nor NOR3 (N10827, N10821, N1619, N7837);
nor NOR3 (N10828, N10819, N850, N10337);
or OR4 (N10829, N10823, N9034, N1327, N6097);
not NOT1 (N10830, N10828);
and AND3 (N10831, N10805, N5274, N3698);
and AND2 (N10832, N10826, N10632);
not NOT1 (N10833, N10829);
nor NOR3 (N10834, N10811, N564, N8351);
not NOT1 (N10835, N10781);
xor XOR2 (N10836, N10825, N2886);
not NOT1 (N10837, N10827);
buf BUF1 (N10838, N10834);
not NOT1 (N10839, N10838);
and AND3 (N10840, N10830, N143, N3749);
or OR3 (N10841, N10840, N2810, N4622);
nand NAND4 (N10842, N10837, N9775, N2409, N6471);
or OR4 (N10843, N10833, N472, N1245, N9394);
nand NAND3 (N10844, N10835, N6499, N3573);
not NOT1 (N10845, N10841);
buf BUF1 (N10846, N10843);
nor NOR3 (N10847, N10844, N2813, N2311);
nor NOR2 (N10848, N10808, N5585);
nand NAND4 (N10849, N10847, N8062, N1904, N10838);
or OR3 (N10850, N10842, N676, N8892);
and AND2 (N10851, N10836, N8282);
not NOT1 (N10852, N10839);
nand NAND2 (N10853, N10851, N559);
nand NAND3 (N10854, N10853, N7840, N6740);
not NOT1 (N10855, N10854);
nand NAND2 (N10856, N10846, N6825);
buf BUF1 (N10857, N10831);
and AND2 (N10858, N10852, N2409);
or OR2 (N10859, N10856, N3654);
nand NAND3 (N10860, N10850, N7612, N4225);
nand NAND2 (N10861, N10855, N1854);
nor NOR2 (N10862, N10857, N443);
nor NOR4 (N10863, N10845, N2316, N7707, N2123);
nand NAND3 (N10864, N10858, N2679, N10578);
or OR2 (N10865, N10863, N1397);
buf BUF1 (N10866, N10849);
nand NAND3 (N10867, N10860, N7579, N3171);
nand NAND3 (N10868, N10866, N6475, N6175);
xor XOR2 (N10869, N10820, N5543);
buf BUF1 (N10870, N10865);
and AND3 (N10871, N10870, N6186, N2346);
not NOT1 (N10872, N10871);
or OR2 (N10873, N10861, N6756);
xor XOR2 (N10874, N10832, N5531);
not NOT1 (N10875, N10873);
or OR4 (N10876, N10848, N10272, N2609, N4876);
xor XOR2 (N10877, N10874, N6979);
and AND3 (N10878, N10868, N4938, N3591);
not NOT1 (N10879, N10867);
nor NOR4 (N10880, N10879, N753, N7507, N4992);
xor XOR2 (N10881, N10869, N8623);
buf BUF1 (N10882, N10876);
buf BUF1 (N10883, N10875);
xor XOR2 (N10884, N10878, N2701);
xor XOR2 (N10885, N10862, N6750);
nand NAND3 (N10886, N10882, N2135, N2710);
nand NAND4 (N10887, N10883, N5182, N7440, N734);
nand NAND2 (N10888, N10884, N6814);
nor NOR2 (N10889, N10872, N3164);
and AND2 (N10890, N10886, N6108);
nor NOR2 (N10891, N10864, N5293);
xor XOR2 (N10892, N10880, N1406);
nand NAND3 (N10893, N10877, N6319, N10770);
and AND3 (N10894, N10891, N2442, N7942);
not NOT1 (N10895, N10888);
or OR2 (N10896, N10885, N9248);
and AND4 (N10897, N10892, N10077, N9654, N7144);
nand NAND4 (N10898, N10859, N7164, N5618, N2757);
not NOT1 (N10899, N10887);
nor NOR2 (N10900, N10896, N4317);
xor XOR2 (N10901, N10899, N3653);
nor NOR4 (N10902, N10898, N8201, N9030, N1085);
not NOT1 (N10903, N10894);
xor XOR2 (N10904, N10895, N4838);
not NOT1 (N10905, N10889);
and AND3 (N10906, N10901, N4443, N4578);
or OR4 (N10907, N10890, N8783, N4243, N3551);
and AND3 (N10908, N10902, N2889, N6058);
nor NOR2 (N10909, N10905, N3314);
and AND4 (N10910, N10893, N8791, N10369, N9284);
nor NOR3 (N10911, N10900, N6866, N7049);
buf BUF1 (N10912, N10906);
not NOT1 (N10913, N10912);
nand NAND2 (N10914, N10903, N8039);
xor XOR2 (N10915, N10897, N9966);
xor XOR2 (N10916, N10914, N3623);
nor NOR3 (N10917, N10881, N5984, N2020);
xor XOR2 (N10918, N10909, N10124);
xor XOR2 (N10919, N10913, N2386);
nand NAND4 (N10920, N10911, N689, N5074, N3537);
not NOT1 (N10921, N10908);
buf BUF1 (N10922, N10920);
nand NAND2 (N10923, N10921, N10239);
xor XOR2 (N10924, N10910, N935);
buf BUF1 (N10925, N10924);
nor NOR3 (N10926, N10907, N5284, N2382);
xor XOR2 (N10927, N10923, N3551);
buf BUF1 (N10928, N10919);
nand NAND2 (N10929, N10904, N9263);
not NOT1 (N10930, N10917);
and AND4 (N10931, N10922, N1787, N3218, N7747);
and AND2 (N10932, N10925, N1704);
nor NOR4 (N10933, N10927, N1246, N1597, N9350);
and AND2 (N10934, N10932, N3540);
buf BUF1 (N10935, N10931);
buf BUF1 (N10936, N10930);
nand NAND2 (N10937, N10916, N2679);
buf BUF1 (N10938, N10926);
xor XOR2 (N10939, N10937, N5537);
and AND2 (N10940, N10935, N7262);
buf BUF1 (N10941, N10915);
nor NOR3 (N10942, N10928, N1704, N2759);
nor NOR2 (N10943, N10929, N3077);
nand NAND3 (N10944, N10918, N2615, N1156);
and AND2 (N10945, N10940, N3748);
or OR3 (N10946, N10943, N2605, N7484);
or OR2 (N10947, N10944, N2298);
not NOT1 (N10948, N10941);
xor XOR2 (N10949, N10933, N3830);
xor XOR2 (N10950, N10939, N540);
buf BUF1 (N10951, N10949);
not NOT1 (N10952, N10936);
nor NOR2 (N10953, N10942, N9956);
xor XOR2 (N10954, N10951, N9583);
xor XOR2 (N10955, N10948, N6035);
nand NAND4 (N10956, N10945, N6491, N27, N876);
nand NAND2 (N10957, N10938, N2030);
nor NOR4 (N10958, N10955, N10840, N962, N8087);
or OR2 (N10959, N10954, N7622);
not NOT1 (N10960, N10952);
xor XOR2 (N10961, N10956, N2102);
nor NOR2 (N10962, N10947, N2136);
buf BUF1 (N10963, N10934);
nand NAND4 (N10964, N10958, N7348, N2800, N4829);
not NOT1 (N10965, N10960);
xor XOR2 (N10966, N10963, N3172);
and AND2 (N10967, N10957, N7347);
and AND2 (N10968, N10950, N1825);
not NOT1 (N10969, N10961);
or OR2 (N10970, N10969, N10952);
nand NAND4 (N10971, N10962, N6754, N6615, N6890);
xor XOR2 (N10972, N10971, N6558);
and AND3 (N10973, N10964, N1454, N9805);
and AND4 (N10974, N10973, N1171, N1753, N1812);
not NOT1 (N10975, N10970);
or OR4 (N10976, N10974, N6269, N7374, N2893);
nand NAND4 (N10977, N10959, N1494, N1491, N2388);
or OR2 (N10978, N10968, N2059);
and AND4 (N10979, N10977, N2960, N10086, N2284);
not NOT1 (N10980, N10946);
nor NOR4 (N10981, N10980, N2161, N4197, N8481);
buf BUF1 (N10982, N10978);
not NOT1 (N10983, N10979);
and AND3 (N10984, N10972, N10287, N9178);
nor NOR2 (N10985, N10976, N3550);
nor NOR4 (N10986, N10953, N290, N2291, N4580);
xor XOR2 (N10987, N10985, N2421);
xor XOR2 (N10988, N10982, N9295);
nand NAND3 (N10989, N10983, N4850, N8112);
nand NAND3 (N10990, N10986, N2170, N585);
not NOT1 (N10991, N10987);
xor XOR2 (N10992, N10966, N8560);
nor NOR2 (N10993, N10989, N5293);
not NOT1 (N10994, N10988);
xor XOR2 (N10995, N10992, N681);
xor XOR2 (N10996, N10967, N4559);
and AND4 (N10997, N10994, N9722, N4458, N10408);
and AND3 (N10998, N10984, N10325, N8113);
nand NAND4 (N10999, N10996, N10036, N6573, N3745);
buf BUF1 (N11000, N10981);
not NOT1 (N11001, N10995);
and AND4 (N11002, N10999, N2900, N4230, N4662);
nand NAND4 (N11003, N10990, N2585, N6550, N424);
buf BUF1 (N11004, N10993);
or OR2 (N11005, N10997, N4955);
buf BUF1 (N11006, N10991);
and AND4 (N11007, N10975, N7367, N2588, N7328);
not NOT1 (N11008, N11001);
nor NOR3 (N11009, N11005, N244, N9941);
or OR2 (N11010, N11007, N6353);
not NOT1 (N11011, N11000);
not NOT1 (N11012, N11010);
not NOT1 (N11013, N10965);
nand NAND4 (N11014, N11013, N7772, N5310, N9771);
and AND2 (N11015, N11006, N233);
and AND2 (N11016, N11008, N8102);
buf BUF1 (N11017, N11011);
and AND3 (N11018, N10998, N10504, N3292);
and AND4 (N11019, N11009, N320, N1001, N10768);
and AND3 (N11020, N11018, N3195, N4085);
buf BUF1 (N11021, N11019);
not NOT1 (N11022, N11004);
xor XOR2 (N11023, N11014, N1659);
nor NOR4 (N11024, N11021, N4151, N3424, N967);
or OR2 (N11025, N11015, N901);
or OR2 (N11026, N11020, N10677);
nand NAND3 (N11027, N11022, N6613, N10179);
nor NOR3 (N11028, N11024, N1574, N3746);
xor XOR2 (N11029, N11027, N4766);
nor NOR4 (N11030, N11016, N1780, N3141, N3487);
buf BUF1 (N11031, N11002);
nand NAND3 (N11032, N11030, N7344, N4327);
or OR3 (N11033, N11026, N7677, N1133);
not NOT1 (N11034, N11031);
buf BUF1 (N11035, N11023);
nand NAND4 (N11036, N11012, N4380, N10421, N5418);
buf BUF1 (N11037, N11035);
nor NOR2 (N11038, N11034, N4717);
nor NOR4 (N11039, N11028, N3503, N8001, N4320);
not NOT1 (N11040, N11003);
nor NOR2 (N11041, N11025, N9672);
not NOT1 (N11042, N11029);
buf BUF1 (N11043, N11017);
and AND3 (N11044, N11041, N807, N5742);
or OR3 (N11045, N11033, N9981, N6552);
and AND2 (N11046, N11038, N8099);
and AND2 (N11047, N11045, N6278);
nand NAND3 (N11048, N11040, N2527, N3608);
nor NOR4 (N11049, N11043, N4637, N4617, N2396);
nand NAND4 (N11050, N11032, N8731, N6368, N2588);
buf BUF1 (N11051, N11042);
not NOT1 (N11052, N11049);
not NOT1 (N11053, N11037);
or OR4 (N11054, N11036, N424, N6371, N4375);
not NOT1 (N11055, N11039);
nor NOR4 (N11056, N11054, N7052, N5712, N1404);
or OR4 (N11057, N11056, N3533, N1685, N7263);
and AND2 (N11058, N11055, N4056);
buf BUF1 (N11059, N11058);
nand NAND4 (N11060, N11048, N1447, N8157, N9516);
and AND2 (N11061, N11059, N10240);
and AND4 (N11062, N11052, N4089, N7009, N214);
not NOT1 (N11063, N11053);
and AND3 (N11064, N11044, N7657, N1871);
nand NAND4 (N11065, N11050, N4548, N8724, N3790);
nand NAND4 (N11066, N11047, N574, N4959, N4685);
nand NAND3 (N11067, N11057, N6382, N3310);
nand NAND2 (N11068, N11060, N10787);
nor NOR3 (N11069, N11063, N3481, N1821);
not NOT1 (N11070, N11062);
or OR2 (N11071, N11061, N9832);
xor XOR2 (N11072, N11046, N8680);
and AND2 (N11073, N11071, N4530);
buf BUF1 (N11074, N11064);
xor XOR2 (N11075, N11065, N1132);
buf BUF1 (N11076, N11066);
and AND2 (N11077, N11068, N10366);
or OR4 (N11078, N11074, N6571, N4807, N292);
nand NAND2 (N11079, N11067, N10566);
nor NOR3 (N11080, N11076, N5151, N1863);
buf BUF1 (N11081, N11080);
buf BUF1 (N11082, N11073);
or OR2 (N11083, N11075, N8632);
or OR2 (N11084, N11072, N9755);
and AND3 (N11085, N11084, N4053, N3096);
nand NAND4 (N11086, N11083, N4230, N7218, N3787);
and AND3 (N11087, N11051, N6043, N2519);
not NOT1 (N11088, N11078);
xor XOR2 (N11089, N11070, N5074);
not NOT1 (N11090, N11081);
nor NOR3 (N11091, N11090, N5994, N10334);
nor NOR3 (N11092, N11069, N4447, N8559);
not NOT1 (N11093, N11087);
nor NOR3 (N11094, N11091, N1002, N1904);
buf BUF1 (N11095, N11086);
nor NOR2 (N11096, N11095, N5975);
or OR2 (N11097, N11094, N5862);
or OR4 (N11098, N11089, N10492, N8995, N3000);
buf BUF1 (N11099, N11077);
nor NOR3 (N11100, N11079, N5996, N7181);
nand NAND4 (N11101, N11085, N7636, N7942, N4683);
buf BUF1 (N11102, N11100);
buf BUF1 (N11103, N11101);
not NOT1 (N11104, N11082);
buf BUF1 (N11105, N11093);
nand NAND4 (N11106, N11098, N8812, N2833, N9243);
not NOT1 (N11107, N11103);
nor NOR3 (N11108, N11107, N4882, N10117);
nand NAND4 (N11109, N11108, N1518, N1961, N9923);
buf BUF1 (N11110, N11097);
xor XOR2 (N11111, N11099, N1518);
nand NAND4 (N11112, N11105, N8462, N5947, N843);
nand NAND3 (N11113, N11096, N9877, N6739);
buf BUF1 (N11114, N11106);
buf BUF1 (N11115, N11110);
nand NAND3 (N11116, N11104, N3047, N8741);
buf BUF1 (N11117, N11092);
or OR4 (N11118, N11117, N3238, N8149, N1286);
nor NOR2 (N11119, N11102, N604);
and AND2 (N11120, N11115, N8852);
nor NOR4 (N11121, N11114, N1369, N9406, N2522);
buf BUF1 (N11122, N11088);
buf BUF1 (N11123, N11121);
nand NAND2 (N11124, N11122, N5240);
nor NOR2 (N11125, N11120, N8350);
xor XOR2 (N11126, N11125, N6699);
buf BUF1 (N11127, N11118);
not NOT1 (N11128, N11127);
nor NOR2 (N11129, N11116, N3659);
xor XOR2 (N11130, N11109, N3108);
buf BUF1 (N11131, N11113);
nand NAND2 (N11132, N11123, N9230);
and AND3 (N11133, N11130, N4348, N7946);
buf BUF1 (N11134, N11129);
xor XOR2 (N11135, N11112, N10249);
buf BUF1 (N11136, N11131);
not NOT1 (N11137, N11136);
nand NAND3 (N11138, N11119, N8180, N1357);
xor XOR2 (N11139, N11111, N6883);
nor NOR3 (N11140, N11124, N9884, N7886);
buf BUF1 (N11141, N11128);
xor XOR2 (N11142, N11139, N2469);
or OR2 (N11143, N11134, N8688);
xor XOR2 (N11144, N11135, N2830);
xor XOR2 (N11145, N11138, N9237);
buf BUF1 (N11146, N11126);
buf BUF1 (N11147, N11145);
or OR4 (N11148, N11133, N5691, N7478, N1892);
not NOT1 (N11149, N11148);
buf BUF1 (N11150, N11144);
and AND3 (N11151, N11140, N1028, N9991);
nand NAND4 (N11152, N11143, N329, N4150, N6756);
xor XOR2 (N11153, N11132, N11018);
xor XOR2 (N11154, N11150, N3833);
xor XOR2 (N11155, N11153, N6707);
nand NAND4 (N11156, N11151, N6052, N7369, N7525);
nor NOR4 (N11157, N11156, N6821, N4325, N3117);
buf BUF1 (N11158, N11137);
and AND4 (N11159, N11152, N1797, N621, N11151);
nand NAND2 (N11160, N11149, N2210);
or OR2 (N11161, N11155, N9518);
xor XOR2 (N11162, N11161, N1029);
nor NOR4 (N11163, N11146, N3871, N3976, N5663);
nand NAND2 (N11164, N11163, N9226);
nand NAND2 (N11165, N11154, N9898);
nor NOR2 (N11166, N11142, N1623);
or OR4 (N11167, N11164, N962, N2781, N3966);
buf BUF1 (N11168, N11147);
xor XOR2 (N11169, N11159, N9945);
nand NAND4 (N11170, N11160, N3035, N10145, N2357);
or OR2 (N11171, N11165, N9004);
xor XOR2 (N11172, N11168, N7252);
nand NAND4 (N11173, N11171, N1663, N166, N6344);
nand NAND2 (N11174, N11162, N980);
and AND2 (N11175, N11172, N687);
not NOT1 (N11176, N11157);
not NOT1 (N11177, N11166);
xor XOR2 (N11178, N11174, N8867);
nand NAND3 (N11179, N11170, N1050, N1479);
and AND4 (N11180, N11173, N9721, N9826, N1634);
and AND3 (N11181, N11179, N11020, N3138);
not NOT1 (N11182, N11141);
xor XOR2 (N11183, N11167, N2406);
and AND2 (N11184, N11177, N2784);
nor NOR2 (N11185, N11184, N3138);
xor XOR2 (N11186, N11158, N8774);
nor NOR3 (N11187, N11176, N9964, N1826);
nand NAND2 (N11188, N11185, N10169);
xor XOR2 (N11189, N11188, N7147);
buf BUF1 (N11190, N11187);
nand NAND2 (N11191, N11181, N8778);
or OR2 (N11192, N11190, N8478);
nor NOR2 (N11193, N11183, N10792);
or OR2 (N11194, N11182, N6069);
or OR4 (N11195, N11186, N8864, N5891, N2832);
not NOT1 (N11196, N11180);
xor XOR2 (N11197, N11195, N7079);
nand NAND3 (N11198, N11196, N3341, N6670);
and AND2 (N11199, N11178, N9397);
nor NOR2 (N11200, N11199, N7841);
nand NAND4 (N11201, N11191, N4466, N3431, N531);
buf BUF1 (N11202, N11200);
nor NOR3 (N11203, N11201, N2137, N5834);
nand NAND4 (N11204, N11189, N10657, N2258, N3706);
nand NAND3 (N11205, N11204, N6287, N1873);
nand NAND3 (N11206, N11175, N1159, N6782);
buf BUF1 (N11207, N11205);
or OR2 (N11208, N11202, N5449);
nor NOR2 (N11209, N11206, N4116);
buf BUF1 (N11210, N11208);
and AND4 (N11211, N11193, N6930, N4224, N1831);
or OR3 (N11212, N11210, N5622, N7718);
nand NAND2 (N11213, N11198, N4842);
nor NOR3 (N11214, N11213, N4773, N565);
nor NOR2 (N11215, N11214, N8086);
nor NOR2 (N11216, N11194, N2584);
or OR2 (N11217, N11209, N7682);
and AND3 (N11218, N11207, N1390, N4268);
nand NAND4 (N11219, N11217, N2324, N1151, N10261);
or OR2 (N11220, N11219, N5158);
and AND2 (N11221, N11169, N9029);
xor XOR2 (N11222, N11197, N5683);
not NOT1 (N11223, N11220);
nor NOR3 (N11224, N11221, N1435, N4071);
and AND4 (N11225, N11211, N6385, N549, N9146);
not NOT1 (N11226, N11218);
nand NAND3 (N11227, N11224, N2735, N447);
buf BUF1 (N11228, N11203);
not NOT1 (N11229, N11216);
buf BUF1 (N11230, N11192);
nor NOR4 (N11231, N11222, N11162, N4783, N8431);
not NOT1 (N11232, N11231);
buf BUF1 (N11233, N11227);
and AND2 (N11234, N11232, N6435);
nand NAND4 (N11235, N11215, N6912, N3328, N3498);
or OR3 (N11236, N11229, N7404, N6169);
or OR3 (N11237, N11230, N9521, N10712);
or OR4 (N11238, N11225, N9544, N1310, N5156);
not NOT1 (N11239, N11233);
xor XOR2 (N11240, N11223, N473);
nand NAND4 (N11241, N11235, N4863, N5470, N5260);
not NOT1 (N11242, N11212);
not NOT1 (N11243, N11236);
and AND2 (N11244, N11240, N9475);
xor XOR2 (N11245, N11243, N10460);
or OR4 (N11246, N11228, N1532, N2562, N5105);
nand NAND2 (N11247, N11245, N7771);
xor XOR2 (N11248, N11226, N10455);
not NOT1 (N11249, N11239);
buf BUF1 (N11250, N11242);
nor NOR4 (N11251, N11244, N1513, N4953, N7009);
buf BUF1 (N11252, N11234);
xor XOR2 (N11253, N11246, N825);
or OR4 (N11254, N11248, N6107, N1723, N3567);
and AND2 (N11255, N11253, N920);
xor XOR2 (N11256, N11252, N4957);
or OR4 (N11257, N11250, N688, N5477, N10533);
buf BUF1 (N11258, N11251);
nor NOR3 (N11259, N11247, N6847, N26);
buf BUF1 (N11260, N11256);
and AND3 (N11261, N11255, N6081, N6739);
or OR2 (N11262, N11238, N2228);
nand NAND2 (N11263, N11261, N9391);
or OR3 (N11264, N11262, N617, N9651);
buf BUF1 (N11265, N11258);
nand NAND3 (N11266, N11264, N5919, N28);
and AND4 (N11267, N11257, N6174, N943, N3318);
nor NOR3 (N11268, N11266, N8017, N2711);
and AND4 (N11269, N11265, N11120, N730, N10427);
and AND2 (N11270, N11269, N2012);
nor NOR3 (N11271, N11241, N1961, N2048);
xor XOR2 (N11272, N11260, N3153);
nand NAND3 (N11273, N11259, N5692, N3099);
buf BUF1 (N11274, N11271);
xor XOR2 (N11275, N11268, N9270);
not NOT1 (N11276, N11237);
and AND2 (N11277, N11272, N3260);
or OR3 (N11278, N11270, N4085, N623);
not NOT1 (N11279, N11267);
nand NAND3 (N11280, N11279, N8358, N1316);
nand NAND2 (N11281, N11254, N3609);
or OR3 (N11282, N11273, N3371, N5697);
and AND2 (N11283, N11282, N108);
not NOT1 (N11284, N11278);
nor NOR4 (N11285, N11274, N592, N9628, N9820);
xor XOR2 (N11286, N11263, N4867);
nand NAND2 (N11287, N11275, N715);
not NOT1 (N11288, N11286);
nor NOR4 (N11289, N11276, N2978, N8065, N9516);
xor XOR2 (N11290, N11285, N2828);
buf BUF1 (N11291, N11249);
nand NAND2 (N11292, N11291, N8256);
nor NOR2 (N11293, N11277, N4053);
and AND4 (N11294, N11283, N3426, N9774, N3316);
nor NOR2 (N11295, N11281, N8168);
nand NAND3 (N11296, N11290, N9017, N639);
xor XOR2 (N11297, N11292, N2485);
nand NAND2 (N11298, N11294, N9306);
xor XOR2 (N11299, N11296, N5212);
nor NOR2 (N11300, N11284, N2123);
nand NAND3 (N11301, N11293, N6997, N10193);
nand NAND3 (N11302, N11301, N4479, N4202);
buf BUF1 (N11303, N11300);
or OR4 (N11304, N11289, N4475, N5870, N3982);
xor XOR2 (N11305, N11304, N2504);
not NOT1 (N11306, N11297);
nor NOR3 (N11307, N11302, N257, N8339);
and AND3 (N11308, N11299, N4411, N173);
or OR2 (N11309, N11308, N1323);
or OR3 (N11310, N11298, N8744, N6177);
or OR4 (N11311, N11307, N956, N5809, N1816);
xor XOR2 (N11312, N11305, N1317);
buf BUF1 (N11313, N11287);
not NOT1 (N11314, N11288);
or OR3 (N11315, N11313, N7892, N10806);
or OR2 (N11316, N11311, N6558);
nor NOR4 (N11317, N11310, N2889, N6869, N9669);
or OR2 (N11318, N11314, N10181);
xor XOR2 (N11319, N11312, N75);
xor XOR2 (N11320, N11280, N1914);
nand NAND3 (N11321, N11318, N8716, N10392);
buf BUF1 (N11322, N11319);
not NOT1 (N11323, N11320);
and AND2 (N11324, N11295, N1285);
buf BUF1 (N11325, N11309);
not NOT1 (N11326, N11324);
and AND2 (N11327, N11306, N11069);
or OR3 (N11328, N11323, N6549, N2554);
nor NOR3 (N11329, N11327, N7927, N10455);
nor NOR3 (N11330, N11325, N10976, N5596);
nor NOR2 (N11331, N11317, N7769);
not NOT1 (N11332, N11303);
not NOT1 (N11333, N11315);
and AND2 (N11334, N11316, N10066);
or OR2 (N11335, N11332, N1378);
nand NAND3 (N11336, N11329, N7974, N2358);
nor NOR2 (N11337, N11335, N9020);
not NOT1 (N11338, N11328);
xor XOR2 (N11339, N11337, N6891);
and AND3 (N11340, N11326, N8436, N7327);
buf BUF1 (N11341, N11322);
nand NAND2 (N11342, N11330, N7422);
not NOT1 (N11343, N11321);
xor XOR2 (N11344, N11341, N3626);
buf BUF1 (N11345, N11343);
xor XOR2 (N11346, N11338, N6856);
nand NAND3 (N11347, N11331, N502, N1630);
and AND4 (N11348, N11345, N4676, N5447, N10109);
nand NAND4 (N11349, N11347, N4797, N862, N675);
xor XOR2 (N11350, N11344, N1506);
nand NAND4 (N11351, N11339, N7945, N1748, N7637);
or OR2 (N11352, N11351, N9063);
xor XOR2 (N11353, N11342, N2233);
xor XOR2 (N11354, N11340, N2854);
or OR2 (N11355, N11350, N10520);
xor XOR2 (N11356, N11355, N954);
not NOT1 (N11357, N11334);
nor NOR4 (N11358, N11352, N11065, N4305, N7046);
not NOT1 (N11359, N11353);
buf BUF1 (N11360, N11357);
not NOT1 (N11361, N11346);
or OR2 (N11362, N11359, N10650);
or OR4 (N11363, N11358, N935, N7715, N7077);
xor XOR2 (N11364, N11348, N11016);
nor NOR4 (N11365, N11364, N6426, N8283, N8609);
nand NAND2 (N11366, N11365, N7689);
xor XOR2 (N11367, N11349, N10186);
xor XOR2 (N11368, N11362, N247);
not NOT1 (N11369, N11360);
not NOT1 (N11370, N11367);
nor NOR4 (N11371, N11370, N6433, N2596, N440);
xor XOR2 (N11372, N11361, N6345);
nor NOR4 (N11373, N11371, N4698, N4606, N109);
not NOT1 (N11374, N11369);
nor NOR3 (N11375, N11368, N6989, N8302);
nor NOR4 (N11376, N11374, N6257, N7953, N4517);
not NOT1 (N11377, N11333);
nand NAND2 (N11378, N11373, N9525);
nor NOR4 (N11379, N11372, N4382, N2032, N3615);
nor NOR4 (N11380, N11375, N8061, N1792, N635);
nor NOR4 (N11381, N11336, N8786, N10757, N2053);
and AND2 (N11382, N11378, N2122);
nor NOR4 (N11383, N11380, N6548, N1237, N10087);
or OR4 (N11384, N11363, N3860, N9224, N8152);
nor NOR4 (N11385, N11384, N928, N4763, N1127);
nor NOR4 (N11386, N11377, N6300, N1948, N5778);
not NOT1 (N11387, N11354);
nand NAND3 (N11388, N11356, N7548, N3734);
and AND2 (N11389, N11388, N9973);
or OR2 (N11390, N11383, N9883);
and AND3 (N11391, N11385, N7717, N9231);
buf BUF1 (N11392, N11386);
not NOT1 (N11393, N11381);
nand NAND3 (N11394, N11392, N9097, N652);
nand NAND4 (N11395, N11394, N5085, N806, N1780);
nor NOR4 (N11396, N11366, N3290, N1335, N1796);
nand NAND3 (N11397, N11393, N3805, N9280);
nand NAND2 (N11398, N11395, N9438);
buf BUF1 (N11399, N11389);
xor XOR2 (N11400, N11390, N1996);
nand NAND3 (N11401, N11379, N9069, N7572);
not NOT1 (N11402, N11398);
not NOT1 (N11403, N11391);
or OR2 (N11404, N11396, N8128);
buf BUF1 (N11405, N11401);
or OR2 (N11406, N11403, N5848);
and AND4 (N11407, N11402, N6401, N295, N3798);
nand NAND3 (N11408, N11405, N5927, N8106);
or OR4 (N11409, N11400, N11098, N7808, N6026);
xor XOR2 (N11410, N11387, N5595);
not NOT1 (N11411, N11407);
and AND3 (N11412, N11399, N3224, N7440);
buf BUF1 (N11413, N11409);
not NOT1 (N11414, N11408);
nand NAND4 (N11415, N11411, N5199, N6161, N5457);
nor NOR2 (N11416, N11406, N2460);
buf BUF1 (N11417, N11412);
not NOT1 (N11418, N11417);
nor NOR4 (N11419, N11397, N577, N2306, N2134);
and AND3 (N11420, N11404, N258, N8113);
and AND2 (N11421, N11418, N7680);
nand NAND4 (N11422, N11413, N8465, N9229, N3827);
or OR2 (N11423, N11415, N10841);
nor NOR2 (N11424, N11422, N4151);
nor NOR2 (N11425, N11423, N5617);
not NOT1 (N11426, N11424);
and AND3 (N11427, N11414, N3600, N1196);
and AND2 (N11428, N11425, N387);
not NOT1 (N11429, N11421);
or OR2 (N11430, N11427, N2815);
nand NAND4 (N11431, N11420, N650, N1855, N3154);
and AND3 (N11432, N11426, N7418, N6214);
buf BUF1 (N11433, N11429);
or OR2 (N11434, N11416, N7119);
nand NAND2 (N11435, N11434, N1961);
and AND3 (N11436, N11433, N5256, N10789);
nand NAND4 (N11437, N11430, N5835, N6987, N8805);
nand NAND4 (N11438, N11376, N5323, N215, N8839);
nor NOR4 (N11439, N11419, N7752, N2687, N9943);
nand NAND2 (N11440, N11437, N3458);
nor NOR2 (N11441, N11410, N6997);
xor XOR2 (N11442, N11428, N7365);
xor XOR2 (N11443, N11439, N3918);
nor NOR2 (N11444, N11441, N11403);
nor NOR2 (N11445, N11436, N7678);
nor NOR4 (N11446, N11382, N7244, N7889, N2160);
and AND3 (N11447, N11442, N3601, N3538);
buf BUF1 (N11448, N11444);
buf BUF1 (N11449, N11440);
or OR3 (N11450, N11431, N180, N2059);
nor NOR2 (N11451, N11445, N8012);
xor XOR2 (N11452, N11435, N11155);
xor XOR2 (N11453, N11447, N2999);
or OR4 (N11454, N11432, N3444, N3523, N753);
nor NOR3 (N11455, N11451, N7264, N8983);
nand NAND4 (N11456, N11452, N10033, N4218, N2066);
or OR2 (N11457, N11448, N10236);
nor NOR4 (N11458, N11449, N7199, N9299, N226);
nand NAND3 (N11459, N11455, N9410, N7683);
and AND2 (N11460, N11446, N4419);
buf BUF1 (N11461, N11459);
and AND2 (N11462, N11461, N11423);
buf BUF1 (N11463, N11438);
buf BUF1 (N11464, N11458);
nor NOR4 (N11465, N11464, N3949, N10008, N8986);
xor XOR2 (N11466, N11463, N2993);
not NOT1 (N11467, N11456);
xor XOR2 (N11468, N11466, N10275);
or OR2 (N11469, N11467, N2158);
xor XOR2 (N11470, N11469, N10882);
buf BUF1 (N11471, N11450);
or OR4 (N11472, N11470, N5644, N8251, N8447);
nor NOR2 (N11473, N11457, N10521);
or OR4 (N11474, N11454, N4135, N4929, N3294);
nor NOR3 (N11475, N11460, N4116, N9258);
not NOT1 (N11476, N11453);
nor NOR4 (N11477, N11465, N6722, N6292, N5260);
or OR4 (N11478, N11475, N3446, N10086, N118);
xor XOR2 (N11479, N11476, N9457);
buf BUF1 (N11480, N11472);
not NOT1 (N11481, N11477);
nand NAND4 (N11482, N11480, N149, N3184, N9360);
buf BUF1 (N11483, N11471);
nand NAND2 (N11484, N11474, N2024);
buf BUF1 (N11485, N11483);
nor NOR4 (N11486, N11479, N159, N11091, N1528);
xor XOR2 (N11487, N11486, N5587);
nor NOR3 (N11488, N11473, N9009, N9599);
nor NOR4 (N11489, N11487, N4301, N9722, N10940);
or OR4 (N11490, N11488, N1926, N3905, N9767);
nor NOR2 (N11491, N11485, N137);
and AND2 (N11492, N11491, N4231);
nor NOR2 (N11493, N11482, N2850);
and AND3 (N11494, N11493, N4400, N8972);
buf BUF1 (N11495, N11492);
and AND3 (N11496, N11462, N2378, N2791);
xor XOR2 (N11497, N11468, N5274);
or OR2 (N11498, N11495, N4536);
not NOT1 (N11499, N11478);
nand NAND2 (N11500, N11496, N8106);
nand NAND3 (N11501, N11484, N3240, N7165);
nor NOR2 (N11502, N11498, N7798);
buf BUF1 (N11503, N11501);
not NOT1 (N11504, N11500);
or OR3 (N11505, N11443, N430, N2773);
xor XOR2 (N11506, N11481, N6103);
nand NAND2 (N11507, N11503, N6382);
or OR4 (N11508, N11502, N285, N1610, N8097);
buf BUF1 (N11509, N11508);
and AND4 (N11510, N11504, N4617, N8432, N3064);
nand NAND3 (N11511, N11489, N7411, N756);
xor XOR2 (N11512, N11490, N8469);
nor NOR2 (N11513, N11506, N814);
xor XOR2 (N11514, N11505, N6652);
xor XOR2 (N11515, N11511, N6691);
and AND3 (N11516, N11512, N9008, N9488);
xor XOR2 (N11517, N11516, N7533);
nor NOR3 (N11518, N11513, N5888, N7506);
buf BUF1 (N11519, N11494);
buf BUF1 (N11520, N11518);
buf BUF1 (N11521, N11519);
buf BUF1 (N11522, N11515);
nand NAND3 (N11523, N11522, N10197, N9094);
xor XOR2 (N11524, N11499, N9789);
and AND4 (N11525, N11517, N9964, N1653, N3290);
and AND2 (N11526, N11521, N6602);
not NOT1 (N11527, N11507);
xor XOR2 (N11528, N11524, N8591);
or OR2 (N11529, N11497, N9072);
not NOT1 (N11530, N11523);
and AND3 (N11531, N11527, N4239, N5893);
not NOT1 (N11532, N11514);
not NOT1 (N11533, N11509);
buf BUF1 (N11534, N11525);
nand NAND2 (N11535, N11530, N7428);
nand NAND2 (N11536, N11529, N4461);
xor XOR2 (N11537, N11528, N9902);
not NOT1 (N11538, N11526);
nor NOR2 (N11539, N11538, N2757);
nor NOR4 (N11540, N11531, N9546, N10668, N10306);
not NOT1 (N11541, N11534);
not NOT1 (N11542, N11541);
xor XOR2 (N11543, N11532, N623);
nor NOR2 (N11544, N11510, N7362);
buf BUF1 (N11545, N11535);
buf BUF1 (N11546, N11545);
and AND4 (N11547, N11533, N3797, N2653, N9127);
nand NAND3 (N11548, N11537, N2869, N11193);
or OR4 (N11549, N11543, N4004, N9192, N2228);
buf BUF1 (N11550, N11536);
and AND4 (N11551, N11542, N2926, N5556, N4141);
nor NOR3 (N11552, N11540, N9796, N4086);
or OR3 (N11553, N11547, N10109, N9894);
nand NAND4 (N11554, N11553, N11268, N10413, N1743);
nand NAND3 (N11555, N11552, N9338, N3782);
xor XOR2 (N11556, N11549, N4482);
and AND4 (N11557, N11544, N3085, N6665, N5417);
xor XOR2 (N11558, N11551, N8334);
and AND2 (N11559, N11520, N10692);
nand NAND2 (N11560, N11546, N2463);
nor NOR4 (N11561, N11556, N5023, N2533, N9158);
or OR3 (N11562, N11554, N4923, N3794);
buf BUF1 (N11563, N11557);
not NOT1 (N11564, N11550);
nor NOR2 (N11565, N11539, N1844);
or OR2 (N11566, N11564, N9348);
and AND2 (N11567, N11561, N5031);
buf BUF1 (N11568, N11559);
nor NOR4 (N11569, N11558, N10461, N5779, N7859);
nor NOR3 (N11570, N11567, N5696, N4525);
not NOT1 (N11571, N11566);
and AND2 (N11572, N11570, N7309);
nand NAND3 (N11573, N11571, N7918, N3946);
not NOT1 (N11574, N11548);
xor XOR2 (N11575, N11560, N242);
or OR2 (N11576, N11574, N7487);
nand NAND4 (N11577, N11576, N7145, N11170, N10977);
nor NOR3 (N11578, N11568, N7172, N4171);
xor XOR2 (N11579, N11573, N7225);
or OR2 (N11580, N11563, N11061);
or OR4 (N11581, N11565, N11318, N10541, N4433);
and AND4 (N11582, N11580, N1548, N3013, N2700);
not NOT1 (N11583, N11577);
nor NOR4 (N11584, N11583, N2478, N4353, N2105);
xor XOR2 (N11585, N11569, N7454);
buf BUF1 (N11586, N11585);
buf BUF1 (N11587, N11584);
buf BUF1 (N11588, N11575);
not NOT1 (N11589, N11562);
nor NOR4 (N11590, N11572, N7493, N5525, N3540);
nor NOR3 (N11591, N11586, N11053, N8979);
nor NOR3 (N11592, N11555, N11238, N6412);
xor XOR2 (N11593, N11588, N3142);
buf BUF1 (N11594, N11579);
or OR2 (N11595, N11581, N3455);
nand NAND4 (N11596, N11582, N380, N10311, N1378);
nand NAND3 (N11597, N11592, N5854, N11388);
xor XOR2 (N11598, N11597, N5579);
nand NAND2 (N11599, N11589, N10201);
and AND2 (N11600, N11587, N3158);
and AND4 (N11601, N11578, N4167, N7648, N9901);
or OR2 (N11602, N11591, N11050);
not NOT1 (N11603, N11600);
nand NAND4 (N11604, N11599, N4409, N3176, N4120);
nor NOR4 (N11605, N11596, N4393, N8095, N7385);
and AND4 (N11606, N11603, N11407, N5244, N4051);
or OR2 (N11607, N11601, N11538);
nor NOR4 (N11608, N11604, N7490, N1495, N367);
and AND2 (N11609, N11605, N3477);
and AND2 (N11610, N11602, N9558);
nand NAND3 (N11611, N11608, N6678, N11170);
nor NOR4 (N11612, N11606, N10161, N2915, N9929);
xor XOR2 (N11613, N11612, N3699);
nor NOR2 (N11614, N11595, N2976);
and AND2 (N11615, N11593, N11497);
not NOT1 (N11616, N11609);
buf BUF1 (N11617, N11607);
nand NAND2 (N11618, N11616, N2300);
or OR4 (N11619, N11614, N11392, N7981, N2562);
or OR2 (N11620, N11610, N3753);
nand NAND2 (N11621, N11611, N2145);
buf BUF1 (N11622, N11598);
or OR4 (N11623, N11618, N1206, N8624, N8341);
and AND2 (N11624, N11613, N4478);
or OR3 (N11625, N11623, N10783, N4963);
buf BUF1 (N11626, N11615);
or OR3 (N11627, N11617, N8290, N11108);
nor NOR3 (N11628, N11627, N2248, N4779);
nand NAND4 (N11629, N11624, N10139, N11049, N9448);
not NOT1 (N11630, N11629);
or OR2 (N11631, N11621, N5527);
not NOT1 (N11632, N11625);
and AND4 (N11633, N11590, N11172, N11241, N5732);
nand NAND2 (N11634, N11594, N6648);
nor NOR3 (N11635, N11634, N6112, N4963);
buf BUF1 (N11636, N11630);
nor NOR4 (N11637, N11626, N954, N5903, N5567);
or OR3 (N11638, N11637, N6652, N4490);
and AND3 (N11639, N11631, N6864, N8353);
xor XOR2 (N11640, N11636, N6312);
and AND2 (N11641, N11633, N7355);
buf BUF1 (N11642, N11639);
nor NOR2 (N11643, N11641, N5524);
not NOT1 (N11644, N11638);
not NOT1 (N11645, N11644);
nor NOR3 (N11646, N11642, N11013, N7275);
nor NOR3 (N11647, N11622, N2595, N10271);
and AND2 (N11648, N11632, N1286);
xor XOR2 (N11649, N11647, N3398);
xor XOR2 (N11650, N11619, N5018);
and AND3 (N11651, N11648, N6997, N7259);
buf BUF1 (N11652, N11640);
nand NAND4 (N11653, N11620, N495, N6558, N4900);
buf BUF1 (N11654, N11646);
xor XOR2 (N11655, N11645, N8642);
xor XOR2 (N11656, N11650, N4261);
buf BUF1 (N11657, N11655);
nor NOR4 (N11658, N11654, N4437, N11567, N4090);
xor XOR2 (N11659, N11651, N4940);
xor XOR2 (N11660, N11628, N851);
buf BUF1 (N11661, N11658);
not NOT1 (N11662, N11656);
buf BUF1 (N11663, N11661);
buf BUF1 (N11664, N11652);
buf BUF1 (N11665, N11664);
not NOT1 (N11666, N11662);
not NOT1 (N11667, N11660);
buf BUF1 (N11668, N11663);
nand NAND4 (N11669, N11667, N5987, N4153, N8725);
nand NAND4 (N11670, N11643, N6836, N6958, N6100);
buf BUF1 (N11671, N11649);
and AND2 (N11672, N11653, N11315);
nor NOR3 (N11673, N11670, N9121, N5877);
xor XOR2 (N11674, N11657, N7927);
nor NOR3 (N11675, N11674, N5246, N3391);
buf BUF1 (N11676, N11668);
xor XOR2 (N11677, N11671, N277);
not NOT1 (N11678, N11635);
nor NOR4 (N11679, N11665, N11379, N4667, N7275);
or OR2 (N11680, N11677, N5846);
xor XOR2 (N11681, N11675, N8684);
buf BUF1 (N11682, N11669);
nand NAND2 (N11683, N11681, N4623);
nor NOR3 (N11684, N11679, N4304, N609);
and AND4 (N11685, N11676, N2630, N9259, N11289);
and AND4 (N11686, N11684, N5626, N3294, N4254);
buf BUF1 (N11687, N11672);
not NOT1 (N11688, N11666);
or OR2 (N11689, N11680, N8639);
buf BUF1 (N11690, N11659);
nor NOR4 (N11691, N11689, N6253, N3706, N10498);
nor NOR4 (N11692, N11685, N10835, N6430, N11523);
nor NOR2 (N11693, N11673, N9509);
nand NAND3 (N11694, N11692, N1843, N8585);
buf BUF1 (N11695, N11693);
or OR2 (N11696, N11686, N283);
and AND3 (N11697, N11696, N2940, N5865);
nand NAND2 (N11698, N11697, N4242);
not NOT1 (N11699, N11691);
nand NAND4 (N11700, N11695, N10104, N8532, N864);
and AND3 (N11701, N11687, N2713, N3597);
not NOT1 (N11702, N11682);
and AND2 (N11703, N11688, N6179);
not NOT1 (N11704, N11703);
nand NAND2 (N11705, N11701, N6569);
and AND4 (N11706, N11698, N477, N6357, N1030);
nor NOR3 (N11707, N11702, N2737, N810);
buf BUF1 (N11708, N11700);
not NOT1 (N11709, N11704);
not NOT1 (N11710, N11707);
nor NOR3 (N11711, N11706, N3408, N2262);
or OR4 (N11712, N11683, N6240, N3858, N11087);
nor NOR2 (N11713, N11711, N2323);
nor NOR3 (N11714, N11709, N1700, N10258);
or OR4 (N11715, N11712, N11571, N981, N9327);
xor XOR2 (N11716, N11710, N5414);
nor NOR3 (N11717, N11708, N7211, N3718);
nor NOR3 (N11718, N11699, N1317, N504);
and AND4 (N11719, N11678, N9371, N6755, N421);
and AND2 (N11720, N11714, N1982);
buf BUF1 (N11721, N11694);
and AND2 (N11722, N11717, N2398);
or OR2 (N11723, N11722, N9088);
or OR3 (N11724, N11690, N2110, N2529);
buf BUF1 (N11725, N11719);
and AND2 (N11726, N11716, N5609);
nand NAND4 (N11727, N11720, N4354, N129, N951);
nand NAND2 (N11728, N11705, N8381);
xor XOR2 (N11729, N11726, N2604);
nor NOR2 (N11730, N11724, N2541);
xor XOR2 (N11731, N11729, N10366);
nand NAND4 (N11732, N11728, N1075, N5739, N2191);
nor NOR2 (N11733, N11731, N7315);
or OR2 (N11734, N11713, N9963);
and AND3 (N11735, N11733, N4186, N9266);
buf BUF1 (N11736, N11725);
or OR3 (N11737, N11721, N5073, N8208);
buf BUF1 (N11738, N11732);
or OR3 (N11739, N11715, N11500, N7661);
nor NOR3 (N11740, N11723, N324, N6091);
nand NAND2 (N11741, N11736, N10000);
xor XOR2 (N11742, N11730, N2767);
xor XOR2 (N11743, N11735, N2081);
nand NAND2 (N11744, N11740, N695);
xor XOR2 (N11745, N11737, N2967);
or OR4 (N11746, N11741, N5947, N6576, N2474);
or OR3 (N11747, N11746, N5152, N11054);
nand NAND4 (N11748, N11743, N981, N3096, N4843);
nor NOR4 (N11749, N11744, N3635, N4189, N3839);
and AND2 (N11750, N11742, N660);
nor NOR4 (N11751, N11727, N2050, N2386, N6703);
xor XOR2 (N11752, N11738, N10435);
or OR3 (N11753, N11751, N3953, N6024);
and AND4 (N11754, N11718, N5183, N1173, N9902);
xor XOR2 (N11755, N11753, N9071);
and AND4 (N11756, N11752, N77, N9420, N3735);
and AND3 (N11757, N11734, N5676, N5270);
or OR4 (N11758, N11748, N10772, N6378, N3321);
buf BUF1 (N11759, N11755);
buf BUF1 (N11760, N11749);
or OR2 (N11761, N11758, N4942);
nor NOR4 (N11762, N11754, N2783, N3640, N10639);
nand NAND2 (N11763, N11757, N1025);
not NOT1 (N11764, N11761);
nor NOR3 (N11765, N11747, N10201, N2332);
not NOT1 (N11766, N11750);
not NOT1 (N11767, N11766);
nand NAND4 (N11768, N11764, N731, N3567, N10990);
nand NAND3 (N11769, N11765, N7144, N938);
nor NOR2 (N11770, N11769, N5688);
or OR3 (N11771, N11739, N4507, N4597);
or OR3 (N11772, N11745, N1501, N11078);
xor XOR2 (N11773, N11759, N2134);
not NOT1 (N11774, N11763);
xor XOR2 (N11775, N11771, N3643);
nand NAND4 (N11776, N11775, N11679, N9681, N7897);
not NOT1 (N11777, N11762);
buf BUF1 (N11778, N11770);
buf BUF1 (N11779, N11756);
xor XOR2 (N11780, N11776, N615);
and AND2 (N11781, N11760, N6875);
not NOT1 (N11782, N11767);
xor XOR2 (N11783, N11777, N4204);
buf BUF1 (N11784, N11779);
not NOT1 (N11785, N11780);
nand NAND2 (N11786, N11772, N249);
not NOT1 (N11787, N11778);
buf BUF1 (N11788, N11784);
not NOT1 (N11789, N11783);
xor XOR2 (N11790, N11782, N8467);
not NOT1 (N11791, N11774);
nand NAND3 (N11792, N11785, N8103, N11024);
xor XOR2 (N11793, N11781, N6371);
and AND2 (N11794, N11787, N181);
nor NOR2 (N11795, N11794, N158);
xor XOR2 (N11796, N11789, N7106);
xor XOR2 (N11797, N11790, N7201);
or OR4 (N11798, N11773, N7811, N7199, N3368);
not NOT1 (N11799, N11796);
not NOT1 (N11800, N11795);
not NOT1 (N11801, N11768);
or OR4 (N11802, N11797, N3837, N10513, N5369);
or OR4 (N11803, N11801, N9236, N10511, N2885);
nand NAND4 (N11804, N11802, N8694, N171, N8069);
and AND4 (N11805, N11799, N8966, N4376, N3616);
nor NOR3 (N11806, N11792, N2184, N7838);
not NOT1 (N11807, N11788);
xor XOR2 (N11808, N11786, N5722);
and AND3 (N11809, N11808, N11168, N4279);
and AND4 (N11810, N11807, N3914, N3021, N3066);
buf BUF1 (N11811, N11791);
nor NOR2 (N11812, N11804, N11125);
and AND2 (N11813, N11800, N6911);
not NOT1 (N11814, N11806);
and AND2 (N11815, N11812, N6940);
and AND4 (N11816, N11803, N6840, N9251, N7372);
not NOT1 (N11817, N11814);
or OR4 (N11818, N11811, N9414, N8428, N1311);
nand NAND3 (N11819, N11793, N3561, N4612);
not NOT1 (N11820, N11805);
not NOT1 (N11821, N11817);
nor NOR2 (N11822, N11810, N5444);
buf BUF1 (N11823, N11813);
nand NAND4 (N11824, N11823, N2762, N8778, N8558);
nor NOR4 (N11825, N11798, N4349, N960, N1765);
nand NAND4 (N11826, N11809, N7995, N4498, N7809);
and AND4 (N11827, N11821, N2065, N6150, N11739);
nor NOR3 (N11828, N11827, N4339, N3233);
or OR3 (N11829, N11816, N8892, N4310);
and AND3 (N11830, N11820, N11576, N10441);
nand NAND4 (N11831, N11829, N2649, N3504, N4661);
or OR3 (N11832, N11818, N426, N3945);
nor NOR2 (N11833, N11815, N1796);
nand NAND4 (N11834, N11828, N8726, N2667, N878);
or OR4 (N11835, N11822, N111, N8657, N3230);
xor XOR2 (N11836, N11833, N4040);
nand NAND4 (N11837, N11830, N6441, N933, N3520);
and AND3 (N11838, N11826, N2809, N2070);
not NOT1 (N11839, N11825);
and AND4 (N11840, N11838, N2047, N8033, N9835);
nand NAND3 (N11841, N11832, N106, N6198);
and AND3 (N11842, N11831, N643, N5318);
not NOT1 (N11843, N11834);
nand NAND2 (N11844, N11839, N2767);
and AND3 (N11845, N11819, N11441, N7577);
nand NAND2 (N11846, N11841, N6400);
not NOT1 (N11847, N11837);
xor XOR2 (N11848, N11843, N7839);
not NOT1 (N11849, N11836);
nand NAND4 (N11850, N11835, N10232, N11084, N6329);
not NOT1 (N11851, N11842);
not NOT1 (N11852, N11850);
not NOT1 (N11853, N11824);
xor XOR2 (N11854, N11847, N2965);
buf BUF1 (N11855, N11846);
nor NOR2 (N11856, N11851, N8457);
not NOT1 (N11857, N11856);
or OR3 (N11858, N11857, N855, N10478);
and AND2 (N11859, N11854, N8362);
xor XOR2 (N11860, N11849, N789);
and AND2 (N11861, N11860, N10969);
buf BUF1 (N11862, N11845);
buf BUF1 (N11863, N11853);
and AND4 (N11864, N11859, N11317, N1138, N5229);
or OR2 (N11865, N11848, N3530);
xor XOR2 (N11866, N11863, N345);
nor NOR3 (N11867, N11840, N10389, N8328);
or OR4 (N11868, N11861, N7982, N9136, N6073);
and AND4 (N11869, N11858, N1066, N6943, N5175);
and AND2 (N11870, N11868, N4771);
nand NAND2 (N11871, N11855, N10301);
buf BUF1 (N11872, N11870);
not NOT1 (N11873, N11844);
not NOT1 (N11874, N11852);
nor NOR4 (N11875, N11864, N8408, N7189, N11642);
nor NOR4 (N11876, N11869, N5967, N8941, N6527);
xor XOR2 (N11877, N11867, N7997);
or OR3 (N11878, N11871, N11498, N2783);
nand NAND2 (N11879, N11873, N6650);
or OR2 (N11880, N11874, N4510);
nand NAND3 (N11881, N11862, N10481, N806);
or OR4 (N11882, N11865, N2779, N7101, N7236);
buf BUF1 (N11883, N11877);
buf BUF1 (N11884, N11883);
buf BUF1 (N11885, N11880);
nand NAND3 (N11886, N11872, N3311, N6272);
buf BUF1 (N11887, N11885);
nand NAND4 (N11888, N11878, N9431, N11826, N9717);
or OR4 (N11889, N11866, N3400, N6133, N757);
nor NOR4 (N11890, N11875, N8843, N7274, N9657);
nand NAND4 (N11891, N11888, N6648, N7726, N9103);
nand NAND3 (N11892, N11890, N5136, N7206);
buf BUF1 (N11893, N11882);
nor NOR3 (N11894, N11879, N11300, N7823);
or OR3 (N11895, N11891, N6304, N5935);
xor XOR2 (N11896, N11881, N10978);
and AND4 (N11897, N11894, N2655, N6323, N4346);
buf BUF1 (N11898, N11895);
buf BUF1 (N11899, N11884);
buf BUF1 (N11900, N11876);
and AND4 (N11901, N11897, N7649, N11797, N4676);
nand NAND3 (N11902, N11899, N6722, N6407);
and AND4 (N11903, N11893, N7717, N10132, N9927);
xor XOR2 (N11904, N11903, N4434);
xor XOR2 (N11905, N11900, N10415);
and AND4 (N11906, N11892, N3046, N10828, N4732);
nand NAND2 (N11907, N11889, N7156);
or OR3 (N11908, N11886, N5745, N11571);
and AND2 (N11909, N11896, N7054);
buf BUF1 (N11910, N11898);
or OR4 (N11911, N11909, N1531, N9038, N11772);
buf BUF1 (N11912, N11906);
xor XOR2 (N11913, N11902, N10084);
nor NOR4 (N11914, N11907, N5989, N9062, N11616);
xor XOR2 (N11915, N11913, N3775);
nand NAND3 (N11916, N11915, N1044, N9467);
buf BUF1 (N11917, N11914);
xor XOR2 (N11918, N11910, N2002);
or OR4 (N11919, N11905, N7282, N3327, N8040);
nand NAND2 (N11920, N11904, N1094);
and AND3 (N11921, N11916, N6129, N11665);
and AND3 (N11922, N11911, N9534, N3905);
nor NOR3 (N11923, N11922, N9113, N7057);
and AND3 (N11924, N11908, N10798, N9716);
buf BUF1 (N11925, N11912);
nor NOR3 (N11926, N11921, N7, N10085);
not NOT1 (N11927, N11918);
and AND3 (N11928, N11925, N6982, N3541);
nand NAND3 (N11929, N11920, N6820, N5835);
buf BUF1 (N11930, N11887);
and AND4 (N11931, N11917, N7102, N3451, N10974);
nand NAND3 (N11932, N11919, N11552, N5017);
not NOT1 (N11933, N11932);
nor NOR2 (N11934, N11901, N9331);
xor XOR2 (N11935, N11928, N4241);
not NOT1 (N11936, N11934);
or OR3 (N11937, N11924, N8799, N10543);
xor XOR2 (N11938, N11930, N9389);
buf BUF1 (N11939, N11929);
or OR3 (N11940, N11927, N6446, N7206);
buf BUF1 (N11941, N11937);
not NOT1 (N11942, N11936);
or OR2 (N11943, N11933, N11040);
nand NAND2 (N11944, N11931, N5593);
nand NAND3 (N11945, N11944, N3284, N10898);
buf BUF1 (N11946, N11943);
buf BUF1 (N11947, N11946);
nand NAND4 (N11948, N11935, N1019, N2342, N7333);
xor XOR2 (N11949, N11938, N2824);
or OR4 (N11950, N11941, N2374, N10034, N7071);
nor NOR3 (N11951, N11949, N1615, N8293);
or OR4 (N11952, N11923, N2427, N7782, N650);
and AND2 (N11953, N11942, N2625);
or OR4 (N11954, N11948, N10879, N6093, N11831);
or OR2 (N11955, N11952, N5777);
xor XOR2 (N11956, N11951, N1093);
buf BUF1 (N11957, N11953);
nor NOR2 (N11958, N11939, N7505);
xor XOR2 (N11959, N11926, N5568);
not NOT1 (N11960, N11945);
or OR2 (N11961, N11959, N4235);
xor XOR2 (N11962, N11947, N9827);
or OR3 (N11963, N11955, N8376, N3110);
xor XOR2 (N11964, N11957, N8524);
or OR4 (N11965, N11960, N288, N10372, N451);
buf BUF1 (N11966, N11964);
buf BUF1 (N11967, N11958);
buf BUF1 (N11968, N11940);
and AND4 (N11969, N11962, N11852, N4465, N2745);
or OR3 (N11970, N11950, N3405, N9401);
nor NOR4 (N11971, N11966, N3449, N4655, N4560);
xor XOR2 (N11972, N11969, N9122);
or OR3 (N11973, N11963, N9542, N29);
or OR2 (N11974, N11961, N4901);
nand NAND4 (N11975, N11971, N6250, N1014, N2424);
or OR2 (N11976, N11975, N4484);
and AND3 (N11977, N11974, N7688, N5779);
and AND3 (N11978, N11968, N1676, N1652);
xor XOR2 (N11979, N11978, N7552);
nand NAND2 (N11980, N11973, N8539);
xor XOR2 (N11981, N11970, N10175);
or OR3 (N11982, N11954, N2915, N10764);
xor XOR2 (N11983, N11972, N8731);
nor NOR2 (N11984, N11981, N9244);
and AND3 (N11985, N11965, N11656, N2726);
nand NAND4 (N11986, N11977, N797, N6333, N10084);
or OR4 (N11987, N11985, N4178, N3042, N1027);
and AND3 (N11988, N11982, N4972, N1408);
or OR2 (N11989, N11988, N3808);
and AND3 (N11990, N11987, N4752, N9496);
not NOT1 (N11991, N11986);
or OR3 (N11992, N11984, N1418, N4385);
buf BUF1 (N11993, N11967);
or OR4 (N11994, N11993, N6722, N351, N2031);
nor NOR3 (N11995, N11994, N9186, N5583);
xor XOR2 (N11996, N11995, N1404);
and AND2 (N11997, N11990, N10259);
or OR3 (N11998, N11991, N3895, N5024);
buf BUF1 (N11999, N11956);
buf BUF1 (N12000, N11979);
and AND3 (N12001, N12000, N11344, N8023);
nor NOR4 (N12002, N12001, N8001, N6704, N5697);
nand NAND4 (N12003, N11999, N874, N1223, N9565);
nand NAND4 (N12004, N12002, N5418, N3812, N9342);
or OR4 (N12005, N11996, N570, N6662, N10182);
xor XOR2 (N12006, N12005, N7118);
nand NAND2 (N12007, N12006, N3849);
not NOT1 (N12008, N11980);
nor NOR4 (N12009, N11989, N6766, N226, N4397);
xor XOR2 (N12010, N11992, N4044);
buf BUF1 (N12011, N11998);
or OR3 (N12012, N12008, N9844, N10663);
nor NOR3 (N12013, N12003, N4210, N2670);
xor XOR2 (N12014, N12009, N7923);
or OR3 (N12015, N12014, N2524, N10956);
nor NOR4 (N12016, N12011, N11712, N9456, N6649);
buf BUF1 (N12017, N12010);
or OR2 (N12018, N12013, N1247);
nand NAND2 (N12019, N12004, N1852);
nor NOR2 (N12020, N11983, N3057);
buf BUF1 (N12021, N11976);
buf BUF1 (N12022, N12019);
not NOT1 (N12023, N12015);
xor XOR2 (N12024, N12021, N3065);
and AND3 (N12025, N12018, N11786, N3225);
nor NOR4 (N12026, N11997, N3683, N2854, N1601);
buf BUF1 (N12027, N12026);
xor XOR2 (N12028, N12016, N11298);
or OR2 (N12029, N12020, N10244);
not NOT1 (N12030, N12024);
or OR2 (N12031, N12023, N3619);
nand NAND4 (N12032, N12012, N7525, N1104, N5239);
buf BUF1 (N12033, N12030);
not NOT1 (N12034, N12007);
not NOT1 (N12035, N12027);
nand NAND4 (N12036, N12035, N11123, N4183, N8352);
nor NOR2 (N12037, N12017, N50);
not NOT1 (N12038, N12034);
xor XOR2 (N12039, N12033, N437);
or OR2 (N12040, N12028, N11314);
not NOT1 (N12041, N12039);
xor XOR2 (N12042, N12031, N8148);
nand NAND3 (N12043, N12032, N349, N218);
buf BUF1 (N12044, N12036);
xor XOR2 (N12045, N12043, N10355);
and AND3 (N12046, N12037, N989, N11077);
buf BUF1 (N12047, N12046);
not NOT1 (N12048, N12022);
not NOT1 (N12049, N12040);
not NOT1 (N12050, N12041);
nand NAND3 (N12051, N12050, N9091, N8922);
nand NAND4 (N12052, N12025, N7987, N4778, N8341);
nor NOR3 (N12053, N12029, N6635, N919);
nand NAND2 (N12054, N12053, N10181);
buf BUF1 (N12055, N12049);
nor NOR3 (N12056, N12052, N8875, N6049);
or OR3 (N12057, N12047, N10749, N3179);
nor NOR4 (N12058, N12056, N3041, N2008, N1354);
xor XOR2 (N12059, N12038, N2070);
or OR2 (N12060, N12058, N719);
and AND4 (N12061, N12054, N6021, N5689, N4492);
not NOT1 (N12062, N12055);
not NOT1 (N12063, N12061);
nor NOR3 (N12064, N12062, N11199, N1631);
buf BUF1 (N12065, N12064);
nand NAND4 (N12066, N12051, N7019, N3896, N4414);
nand NAND4 (N12067, N12057, N11757, N4576, N4636);
xor XOR2 (N12068, N12048, N11156);
or OR4 (N12069, N12059, N442, N2089, N6634);
buf BUF1 (N12070, N12045);
buf BUF1 (N12071, N12070);
xor XOR2 (N12072, N12065, N7863);
not NOT1 (N12073, N12044);
nand NAND2 (N12074, N12060, N10844);
or OR3 (N12075, N12063, N538, N4416);
not NOT1 (N12076, N12072);
nor NOR2 (N12077, N12042, N3108);
buf BUF1 (N12078, N12075);
nor NOR2 (N12079, N12067, N6040);
nand NAND2 (N12080, N12074, N1436);
or OR3 (N12081, N12066, N1788, N3307);
and AND2 (N12082, N12079, N6554);
not NOT1 (N12083, N12082);
nand NAND3 (N12084, N12083, N4821, N2847);
or OR2 (N12085, N12073, N1781);
nand NAND2 (N12086, N12085, N1962);
nand NAND3 (N12087, N12080, N5191, N5333);
and AND2 (N12088, N12071, N8548);
buf BUF1 (N12089, N12076);
nand NAND2 (N12090, N12078, N4469);
buf BUF1 (N12091, N12087);
nor NOR4 (N12092, N12068, N7245, N1095, N4893);
not NOT1 (N12093, N12092);
nor NOR2 (N12094, N12093, N8798);
nor NOR2 (N12095, N12077, N9996);
and AND3 (N12096, N12090, N11687, N1870);
nand NAND3 (N12097, N12086, N3933, N9672);
or OR4 (N12098, N12097, N6942, N1450, N8245);
nor NOR4 (N12099, N12098, N5768, N1302, N900);
buf BUF1 (N12100, N12099);
and AND4 (N12101, N12069, N3407, N9504, N142);
xor XOR2 (N12102, N12089, N2871);
buf BUF1 (N12103, N12101);
buf BUF1 (N12104, N12102);
buf BUF1 (N12105, N12100);
buf BUF1 (N12106, N12095);
not NOT1 (N12107, N12094);
or OR4 (N12108, N12091, N330, N11228, N4734);
not NOT1 (N12109, N12096);
xor XOR2 (N12110, N12084, N7270);
nor NOR2 (N12111, N12109, N9860);
and AND4 (N12112, N12088, N9592, N2841, N6527);
not NOT1 (N12113, N12105);
buf BUF1 (N12114, N12113);
xor XOR2 (N12115, N12103, N8678);
and AND2 (N12116, N12115, N1692);
xor XOR2 (N12117, N12116, N3764);
not NOT1 (N12118, N12111);
nor NOR2 (N12119, N12104, N6577);
and AND3 (N12120, N12117, N12078, N2797);
and AND3 (N12121, N12120, N9137, N2485);
nor NOR2 (N12122, N12107, N8780);
xor XOR2 (N12123, N12119, N9046);
nand NAND2 (N12124, N12108, N6464);
xor XOR2 (N12125, N12110, N7544);
nand NAND4 (N12126, N12122, N1599, N11487, N3727);
or OR3 (N12127, N12126, N95, N6051);
not NOT1 (N12128, N12123);
not NOT1 (N12129, N12121);
not NOT1 (N12130, N12081);
buf BUF1 (N12131, N12127);
nand NAND2 (N12132, N12114, N2760);
xor XOR2 (N12133, N12124, N3602);
not NOT1 (N12134, N12129);
nand NAND3 (N12135, N12131, N8251, N1169);
buf BUF1 (N12136, N12132);
and AND4 (N12137, N12133, N3123, N5045, N9796);
xor XOR2 (N12138, N12130, N7591);
and AND2 (N12139, N12137, N4962);
xor XOR2 (N12140, N12128, N3711);
buf BUF1 (N12141, N12125);
or OR4 (N12142, N12136, N8093, N1194, N1329);
and AND2 (N12143, N12140, N11493);
or OR2 (N12144, N12142, N8208);
nand NAND2 (N12145, N12138, N11700);
or OR3 (N12146, N12135, N2297, N7855);
buf BUF1 (N12147, N12139);
nor NOR2 (N12148, N12143, N8552);
xor XOR2 (N12149, N12147, N1861);
xor XOR2 (N12150, N12145, N5386);
nand NAND2 (N12151, N12144, N397);
and AND3 (N12152, N12151, N3107, N405);
buf BUF1 (N12153, N12152);
nor NOR4 (N12154, N12112, N664, N2662, N4147);
and AND3 (N12155, N12118, N3642, N3253);
buf BUF1 (N12156, N12148);
and AND2 (N12157, N12146, N12052);
nand NAND2 (N12158, N12156, N9838);
not NOT1 (N12159, N12157);
not NOT1 (N12160, N12153);
or OR3 (N12161, N12158, N548, N2238);
nand NAND2 (N12162, N12106, N1281);
not NOT1 (N12163, N12159);
and AND3 (N12164, N12161, N810, N6008);
and AND2 (N12165, N12155, N10066);
or OR2 (N12166, N12149, N5910);
not NOT1 (N12167, N12166);
nand NAND4 (N12168, N12165, N8093, N1613, N9904);
nand NAND3 (N12169, N12164, N10198, N6148);
and AND3 (N12170, N12160, N1077, N1909);
nand NAND4 (N12171, N12163, N1479, N2229, N10206);
not NOT1 (N12172, N12168);
xor XOR2 (N12173, N12162, N7414);
not NOT1 (N12174, N12167);
or OR2 (N12175, N12172, N6616);
nand NAND4 (N12176, N12170, N8368, N4858, N3276);
not NOT1 (N12177, N12174);
or OR3 (N12178, N12171, N10568, N6750);
nor NOR3 (N12179, N12154, N1200, N9455);
or OR4 (N12180, N12178, N9501, N2482, N1585);
and AND2 (N12181, N12141, N11797);
buf BUF1 (N12182, N12169);
nand NAND3 (N12183, N12182, N7088, N4987);
or OR3 (N12184, N12177, N838, N11069);
or OR2 (N12185, N12173, N731);
or OR3 (N12186, N12185, N6555, N2396);
and AND4 (N12187, N12179, N3139, N6614, N9095);
nor NOR4 (N12188, N12150, N8008, N9658, N9287);
xor XOR2 (N12189, N12188, N4142);
xor XOR2 (N12190, N12189, N11789);
and AND3 (N12191, N12175, N1806, N2251);
xor XOR2 (N12192, N12190, N8310);
buf BUF1 (N12193, N12187);
buf BUF1 (N12194, N12181);
nor NOR4 (N12195, N12186, N3446, N7436, N7789);
nor NOR2 (N12196, N12192, N7511);
nand NAND3 (N12197, N12193, N4916, N97);
buf BUF1 (N12198, N12196);
and AND4 (N12199, N12183, N519, N727, N4918);
xor XOR2 (N12200, N12198, N7878);
nor NOR2 (N12201, N12180, N8895);
buf BUF1 (N12202, N12184);
buf BUF1 (N12203, N12134);
or OR2 (N12204, N12176, N6214);
or OR3 (N12205, N12200, N4798, N7917);
or OR2 (N12206, N12202, N395);
and AND2 (N12207, N12204, N6401);
nor NOR2 (N12208, N12201, N10845);
and AND4 (N12209, N12205, N7917, N5267, N6212);
nand NAND4 (N12210, N12195, N9061, N1993, N4233);
nand NAND3 (N12211, N12209, N11401, N5374);
nand NAND2 (N12212, N12194, N6593);
nand NAND2 (N12213, N12191, N4524);
and AND4 (N12214, N12208, N3606, N10084, N5894);
buf BUF1 (N12215, N12212);
nor NOR3 (N12216, N12207, N380, N7367);
or OR2 (N12217, N12211, N11559);
xor XOR2 (N12218, N12216, N5931);
nor NOR2 (N12219, N12197, N463);
and AND3 (N12220, N12199, N1129, N4601);
and AND4 (N12221, N12213, N2790, N5956, N2336);
and AND3 (N12222, N12203, N6998, N684);
and AND3 (N12223, N12219, N4048, N3768);
nor NOR3 (N12224, N12223, N2523, N1052);
or OR4 (N12225, N12220, N9591, N6234, N6353);
or OR3 (N12226, N12215, N888, N3572);
buf BUF1 (N12227, N12224);
buf BUF1 (N12228, N12210);
buf BUF1 (N12229, N12217);
not NOT1 (N12230, N12225);
not NOT1 (N12231, N12221);
xor XOR2 (N12232, N12231, N3458);
or OR4 (N12233, N12229, N8416, N6024, N11214);
or OR2 (N12234, N12228, N5990);
nand NAND4 (N12235, N12230, N2066, N4266, N1515);
or OR4 (N12236, N12226, N11188, N1817, N6937);
or OR4 (N12237, N12236, N3035, N6985, N10603);
xor XOR2 (N12238, N12214, N535);
or OR2 (N12239, N12234, N11781);
or OR2 (N12240, N12233, N1875);
xor XOR2 (N12241, N12227, N6672);
nor NOR3 (N12242, N12222, N8152, N8156);
buf BUF1 (N12243, N12206);
nand NAND2 (N12244, N12243, N6968);
not NOT1 (N12245, N12240);
nand NAND3 (N12246, N12241, N6955, N5447);
or OR3 (N12247, N12218, N9766, N6448);
and AND4 (N12248, N12244, N1516, N4370, N2943);
and AND2 (N12249, N12237, N11943);
xor XOR2 (N12250, N12232, N2089);
nand NAND2 (N12251, N12248, N10392);
not NOT1 (N12252, N12242);
nand NAND4 (N12253, N12251, N6836, N9874, N2837);
or OR3 (N12254, N12253, N6230, N6132);
and AND2 (N12255, N12246, N5374);
xor XOR2 (N12256, N12254, N3635);
not NOT1 (N12257, N12249);
not NOT1 (N12258, N12235);
and AND3 (N12259, N12250, N8411, N11724);
not NOT1 (N12260, N12255);
nand NAND3 (N12261, N12260, N5601, N1344);
and AND3 (N12262, N12247, N1976, N4795);
or OR3 (N12263, N12238, N11467, N350);
and AND4 (N12264, N12239, N5690, N3227, N6744);
buf BUF1 (N12265, N12261);
and AND2 (N12266, N12259, N9272);
or OR4 (N12267, N12258, N1061, N10996, N8638);
not NOT1 (N12268, N12257);
or OR2 (N12269, N12264, N5351);
not NOT1 (N12270, N12268);
not NOT1 (N12271, N12265);
or OR4 (N12272, N12263, N793, N10148, N4767);
nand NAND2 (N12273, N12272, N4789);
buf BUF1 (N12274, N12273);
or OR2 (N12275, N12267, N12261);
and AND3 (N12276, N12269, N10814, N5143);
nand NAND3 (N12277, N12274, N11659, N8152);
buf BUF1 (N12278, N12266);
nor NOR2 (N12279, N12278, N6969);
not NOT1 (N12280, N12270);
or OR4 (N12281, N12271, N8013, N12250, N1945);
buf BUF1 (N12282, N12252);
or OR4 (N12283, N12262, N10251, N2715, N2976);
or OR3 (N12284, N12283, N3870, N4409);
or OR3 (N12285, N12256, N4926, N8253);
and AND4 (N12286, N12279, N981, N10083, N11533);
and AND3 (N12287, N12275, N6413, N3959);
buf BUF1 (N12288, N12282);
buf BUF1 (N12289, N12286);
nor NOR3 (N12290, N12280, N3782, N3891);
xor XOR2 (N12291, N12285, N4521);
or OR2 (N12292, N12276, N11725);
nand NAND4 (N12293, N12284, N3222, N7985, N8785);
nor NOR3 (N12294, N12245, N6262, N9662);
nor NOR3 (N12295, N12292, N3517, N4188);
and AND4 (N12296, N12294, N6488, N927, N10214);
nor NOR4 (N12297, N12293, N8155, N11829, N3427);
or OR3 (N12298, N12289, N1020, N9695);
nor NOR2 (N12299, N12277, N11502);
not NOT1 (N12300, N12281);
xor XOR2 (N12301, N12297, N7488);
nand NAND4 (N12302, N12290, N9318, N7280, N11903);
nand NAND4 (N12303, N12299, N2955, N10720, N7521);
buf BUF1 (N12304, N12300);
not NOT1 (N12305, N12304);
nor NOR2 (N12306, N12305, N8580);
nor NOR2 (N12307, N12295, N7695);
not NOT1 (N12308, N12288);
or OR4 (N12309, N12296, N7722, N11648, N6401);
not NOT1 (N12310, N12309);
nor NOR3 (N12311, N12302, N1509, N10468);
buf BUF1 (N12312, N12311);
and AND4 (N12313, N12291, N4593, N3646, N1571);
and AND3 (N12314, N12308, N4487, N12158);
nor NOR4 (N12315, N12301, N2962, N7586, N10926);
nand NAND2 (N12316, N12313, N2338);
not NOT1 (N12317, N12306);
nor NOR3 (N12318, N12314, N946, N7845);
buf BUF1 (N12319, N12315);
and AND2 (N12320, N12312, N10538);
nand NAND4 (N12321, N12310, N10774, N2326, N6497);
xor XOR2 (N12322, N12318, N6210);
buf BUF1 (N12323, N12298);
xor XOR2 (N12324, N12319, N9451);
buf BUF1 (N12325, N12322);
nor NOR2 (N12326, N12316, N9842);
or OR2 (N12327, N12324, N12198);
and AND3 (N12328, N12327, N541, N8703);
nand NAND2 (N12329, N12325, N2664);
not NOT1 (N12330, N12320);
or OR3 (N12331, N12317, N7370, N9092);
buf BUF1 (N12332, N12287);
buf BUF1 (N12333, N12330);
not NOT1 (N12334, N12331);
buf BUF1 (N12335, N12332);
nand NAND4 (N12336, N12326, N2371, N3369, N9842);
nand NAND4 (N12337, N12323, N9937, N12101, N1222);
nor NOR3 (N12338, N12334, N3043, N8022);
or OR2 (N12339, N12321, N10125);
nand NAND3 (N12340, N12333, N7672, N2325);
or OR2 (N12341, N12338, N1234);
and AND2 (N12342, N12340, N7315);
and AND2 (N12343, N12336, N6677);
nand NAND3 (N12344, N12341, N9160, N4123);
nand NAND4 (N12345, N12329, N3460, N11730, N7142);
xor XOR2 (N12346, N12342, N5099);
buf BUF1 (N12347, N12337);
and AND4 (N12348, N12346, N9305, N11662, N10182);
or OR4 (N12349, N12328, N8162, N4016, N6469);
nand NAND4 (N12350, N12344, N11334, N10603, N2797);
xor XOR2 (N12351, N12339, N2968);
not NOT1 (N12352, N12349);
nand NAND2 (N12353, N12350, N6868);
nand NAND2 (N12354, N12351, N12302);
nor NOR2 (N12355, N12303, N4236);
or OR3 (N12356, N12355, N3617, N3089);
or OR3 (N12357, N12348, N5648, N4439);
buf BUF1 (N12358, N12354);
nand NAND4 (N12359, N12343, N12311, N4018, N11184);
and AND4 (N12360, N12353, N4402, N8797, N978);
not NOT1 (N12361, N12335);
xor XOR2 (N12362, N12361, N10406);
not NOT1 (N12363, N12347);
nand NAND3 (N12364, N12352, N65, N3751);
buf BUF1 (N12365, N12307);
buf BUF1 (N12366, N12362);
xor XOR2 (N12367, N12357, N1028);
xor XOR2 (N12368, N12359, N5826);
buf BUF1 (N12369, N12360);
nand NAND3 (N12370, N12345, N1229, N6545);
or OR3 (N12371, N12356, N119, N6124);
nor NOR3 (N12372, N12364, N2762, N3532);
nor NOR3 (N12373, N12358, N4665, N10867);
buf BUF1 (N12374, N12373);
not NOT1 (N12375, N12365);
nand NAND2 (N12376, N12370, N7447);
nand NAND2 (N12377, N12363, N3586);
nor NOR2 (N12378, N12369, N5689);
or OR3 (N12379, N12378, N11851, N2231);
not NOT1 (N12380, N12376);
xor XOR2 (N12381, N12379, N3547);
xor XOR2 (N12382, N12372, N8703);
nor NOR2 (N12383, N12381, N97);
nand NAND2 (N12384, N12366, N5094);
nor NOR4 (N12385, N12368, N3873, N12033, N5872);
nand NAND4 (N12386, N12367, N3432, N6841, N6429);
nand NAND3 (N12387, N12375, N507, N5465);
and AND4 (N12388, N12377, N952, N7463, N1789);
buf BUF1 (N12389, N12385);
nand NAND2 (N12390, N12383, N8647);
xor XOR2 (N12391, N12382, N7944);
and AND2 (N12392, N12391, N9379);
xor XOR2 (N12393, N12384, N11160);
buf BUF1 (N12394, N12388);
nand NAND2 (N12395, N12389, N9784);
xor XOR2 (N12396, N12374, N8072);
or OR4 (N12397, N12395, N4897, N1779, N5897);
not NOT1 (N12398, N12392);
not NOT1 (N12399, N12380);
nand NAND3 (N12400, N12397, N3060, N3127);
xor XOR2 (N12401, N12394, N11847);
and AND2 (N12402, N12400, N8672);
nand NAND2 (N12403, N12393, N6873);
buf BUF1 (N12404, N12401);
or OR3 (N12405, N12403, N1281, N4243);
or OR4 (N12406, N12404, N7720, N1683, N6791);
not NOT1 (N12407, N12402);
xor XOR2 (N12408, N12386, N9649);
not NOT1 (N12409, N12407);
and AND2 (N12410, N12387, N11236);
not NOT1 (N12411, N12371);
nand NAND2 (N12412, N12398, N6518);
nand NAND4 (N12413, N12396, N1014, N5587, N999);
not NOT1 (N12414, N12409);
or OR3 (N12415, N12411, N614, N3369);
or OR4 (N12416, N12408, N2369, N7239, N10783);
nor NOR4 (N12417, N12410, N175, N3672, N4444);
and AND3 (N12418, N12412, N2769, N4283);
nor NOR3 (N12419, N12418, N10754, N4657);
nor NOR3 (N12420, N12414, N10244, N7306);
nand NAND3 (N12421, N12406, N7476, N6782);
nor NOR2 (N12422, N12416, N1177);
not NOT1 (N12423, N12413);
or OR2 (N12424, N12419, N10160);
not NOT1 (N12425, N12421);
not NOT1 (N12426, N12390);
buf BUF1 (N12427, N12405);
or OR2 (N12428, N12415, N1410);
nand NAND2 (N12429, N12428, N4645);
buf BUF1 (N12430, N12420);
nand NAND2 (N12431, N12423, N6300);
buf BUF1 (N12432, N12426);
nor NOR3 (N12433, N12429, N4855, N8346);
nor NOR4 (N12434, N12427, N11436, N6729, N10529);
or OR2 (N12435, N12422, N328);
or OR2 (N12436, N12435, N10397);
or OR4 (N12437, N12430, N8184, N12063, N8987);
and AND4 (N12438, N12424, N2328, N12274, N21);
or OR4 (N12439, N12399, N724, N6068, N65);
not NOT1 (N12440, N12437);
nand NAND3 (N12441, N12417, N10834, N8474);
nor NOR4 (N12442, N12432, N3223, N1581, N7443);
or OR4 (N12443, N12441, N4725, N5050, N11852);
and AND3 (N12444, N12443, N617, N9143);
or OR2 (N12445, N12431, N9122);
not NOT1 (N12446, N12425);
nor NOR3 (N12447, N12444, N5309, N8062);
buf BUF1 (N12448, N12442);
nand NAND4 (N12449, N12446, N1399, N9557, N9527);
xor XOR2 (N12450, N12439, N11153);
xor XOR2 (N12451, N12449, N1994);
nor NOR3 (N12452, N12447, N6327, N10622);
buf BUF1 (N12453, N12452);
and AND2 (N12454, N12453, N6527);
not NOT1 (N12455, N12438);
xor XOR2 (N12456, N12433, N5223);
buf BUF1 (N12457, N12455);
nor NOR3 (N12458, N12440, N2786, N490);
nor NOR3 (N12459, N12458, N3188, N142);
nand NAND2 (N12460, N12459, N6277);
xor XOR2 (N12461, N12436, N4436);
and AND4 (N12462, N12461, N10441, N8269, N4525);
not NOT1 (N12463, N12454);
nor NOR3 (N12464, N12434, N8501, N1522);
and AND2 (N12465, N12462, N1052);
buf BUF1 (N12466, N12451);
not NOT1 (N12467, N12448);
buf BUF1 (N12468, N12466);
xor XOR2 (N12469, N12468, N2864);
nor NOR2 (N12470, N12445, N1769);
and AND3 (N12471, N12467, N10113, N12336);
nor NOR3 (N12472, N12463, N3856, N2667);
buf BUF1 (N12473, N12465);
xor XOR2 (N12474, N12471, N11492);
buf BUF1 (N12475, N12456);
nand NAND3 (N12476, N12464, N5229, N10412);
xor XOR2 (N12477, N12450, N576);
xor XOR2 (N12478, N12473, N1019);
and AND3 (N12479, N12460, N1191, N1708);
nor NOR2 (N12480, N12474, N471);
nor NOR3 (N12481, N12477, N6316, N8366);
xor XOR2 (N12482, N12478, N10879);
xor XOR2 (N12483, N12481, N2979);
not NOT1 (N12484, N12469);
nand NAND4 (N12485, N12470, N2906, N3502, N12455);
xor XOR2 (N12486, N12472, N8181);
not NOT1 (N12487, N12480);
not NOT1 (N12488, N12475);
buf BUF1 (N12489, N12457);
xor XOR2 (N12490, N12476, N10054);
or OR3 (N12491, N12484, N4485, N7566);
buf BUF1 (N12492, N12491);
not NOT1 (N12493, N12488);
and AND3 (N12494, N12482, N12391, N8810);
or OR2 (N12495, N12492, N10953);
or OR4 (N12496, N12479, N12407, N9808, N1866);
and AND2 (N12497, N12486, N11429);
nand NAND4 (N12498, N12483, N10132, N3373, N2362);
or OR4 (N12499, N12497, N651, N5012, N10280);
not NOT1 (N12500, N12489);
xor XOR2 (N12501, N12495, N11456);
buf BUF1 (N12502, N12498);
not NOT1 (N12503, N12496);
nand NAND2 (N12504, N12499, N5177);
xor XOR2 (N12505, N12487, N9270);
xor XOR2 (N12506, N12502, N2548);
or OR3 (N12507, N12505, N6730, N9026);
nor NOR2 (N12508, N12506, N698);
buf BUF1 (N12509, N12493);
not NOT1 (N12510, N12507);
xor XOR2 (N12511, N12510, N9650);
nand NAND4 (N12512, N12504, N7941, N10165, N83);
xor XOR2 (N12513, N12511, N7348);
not NOT1 (N12514, N12490);
xor XOR2 (N12515, N12485, N10909);
or OR2 (N12516, N12501, N8059);
not NOT1 (N12517, N12503);
or OR4 (N12518, N12494, N11366, N8112, N10166);
or OR3 (N12519, N12508, N4576, N12146);
xor XOR2 (N12520, N12515, N429);
xor XOR2 (N12521, N12517, N8133);
nand NAND4 (N12522, N12520, N4200, N5789, N11994);
buf BUF1 (N12523, N12509);
and AND3 (N12524, N12523, N3834, N11899);
xor XOR2 (N12525, N12516, N11510);
or OR4 (N12526, N12518, N9061, N3354, N6763);
nor NOR3 (N12527, N12525, N6802, N8465);
buf BUF1 (N12528, N12522);
or OR2 (N12529, N12527, N5085);
or OR4 (N12530, N12524, N5629, N2658, N11175);
or OR2 (N12531, N12521, N5371);
xor XOR2 (N12532, N12528, N648);
or OR2 (N12533, N12529, N8980);
or OR3 (N12534, N12532, N3211, N9902);
xor XOR2 (N12535, N12519, N2859);
nor NOR4 (N12536, N12533, N8880, N2266, N6299);
or OR4 (N12537, N12514, N10915, N459, N7990);
xor XOR2 (N12538, N12534, N4453);
xor XOR2 (N12539, N12538, N807);
and AND4 (N12540, N12500, N12380, N8038, N910);
nor NOR2 (N12541, N12535, N3528);
and AND3 (N12542, N12539, N9754, N3811);
or OR4 (N12543, N12513, N11564, N8347, N7122);
nand NAND2 (N12544, N12530, N3956);
or OR2 (N12545, N12540, N9556);
buf BUF1 (N12546, N12537);
or OR4 (N12547, N12536, N10392, N5318, N2589);
or OR4 (N12548, N12543, N9151, N6474, N2226);
or OR3 (N12549, N12541, N2419, N1449);
buf BUF1 (N12550, N12547);
nor NOR4 (N12551, N12546, N3767, N6337, N10193);
not NOT1 (N12552, N12526);
buf BUF1 (N12553, N12551);
nor NOR4 (N12554, N12512, N2632, N12146, N1597);
xor XOR2 (N12555, N12552, N12363);
nand NAND2 (N12556, N12545, N12256);
not NOT1 (N12557, N12531);
or OR4 (N12558, N12557, N10905, N1512, N6256);
buf BUF1 (N12559, N12556);
nand NAND2 (N12560, N12559, N109);
nand NAND3 (N12561, N12550, N4902, N4901);
nor NOR3 (N12562, N12542, N11953, N5389);
xor XOR2 (N12563, N12555, N4184);
nand NAND4 (N12564, N12558, N11350, N2223, N8580);
or OR2 (N12565, N12561, N4304);
and AND2 (N12566, N12565, N2805);
not NOT1 (N12567, N12544);
xor XOR2 (N12568, N12564, N770);
or OR4 (N12569, N12554, N6966, N10216, N1709);
nand NAND3 (N12570, N12567, N8878, N1687);
nor NOR3 (N12571, N12562, N2446, N6428);
nor NOR4 (N12572, N12553, N5260, N6298, N11351);
xor XOR2 (N12573, N12569, N9501);
nor NOR3 (N12574, N12560, N2818, N7085);
xor XOR2 (N12575, N12548, N658);
and AND3 (N12576, N12570, N10502, N8837);
buf BUF1 (N12577, N12571);
buf BUF1 (N12578, N12577);
nor NOR3 (N12579, N12574, N1958, N8595);
or OR3 (N12580, N12579, N10478, N6979);
buf BUF1 (N12581, N12572);
xor XOR2 (N12582, N12575, N5963);
not NOT1 (N12583, N12576);
buf BUF1 (N12584, N12581);
and AND2 (N12585, N12578, N1218);
nor NOR3 (N12586, N12573, N1748, N1926);
not NOT1 (N12587, N12549);
buf BUF1 (N12588, N12587);
nor NOR4 (N12589, N12563, N8026, N11308, N3077);
nor NOR4 (N12590, N12568, N1259, N11797, N7102);
and AND4 (N12591, N12590, N124, N5192, N11224);
nor NOR2 (N12592, N12583, N10865);
or OR2 (N12593, N12591, N9762);
nand NAND4 (N12594, N12586, N5967, N5013, N7570);
not NOT1 (N12595, N12593);
and AND3 (N12596, N12589, N9301, N4188);
nor NOR2 (N12597, N12582, N11082);
nand NAND3 (N12598, N12584, N1184, N7273);
buf BUF1 (N12599, N12595);
and AND3 (N12600, N12596, N4813, N10818);
and AND3 (N12601, N12580, N9781, N10119);
and AND3 (N12602, N12592, N2532, N11671);
not NOT1 (N12603, N12601);
nand NAND4 (N12604, N12594, N791, N2705, N10240);
nor NOR2 (N12605, N12603, N11401);
xor XOR2 (N12606, N12600, N2476);
xor XOR2 (N12607, N12598, N7254);
nor NOR4 (N12608, N12604, N6804, N6876, N8013);
nor NOR2 (N12609, N12585, N1610);
nor NOR2 (N12610, N12607, N984);
and AND2 (N12611, N12608, N12057);
xor XOR2 (N12612, N12611, N5658);
nor NOR2 (N12613, N12609, N3137);
nor NOR4 (N12614, N12588, N2647, N10, N10384);
nor NOR4 (N12615, N12610, N1160, N3071, N5554);
and AND2 (N12616, N12614, N3728);
not NOT1 (N12617, N12615);
not NOT1 (N12618, N12606);
not NOT1 (N12619, N12602);
nor NOR4 (N12620, N12613, N11320, N7014, N10870);
nor NOR4 (N12621, N12605, N4728, N7917, N7459);
buf BUF1 (N12622, N12617);
or OR3 (N12623, N12620, N6722, N11167);
nor NOR3 (N12624, N12622, N6700, N739);
not NOT1 (N12625, N12599);
buf BUF1 (N12626, N12597);
not NOT1 (N12627, N12626);
xor XOR2 (N12628, N12566, N4746);
xor XOR2 (N12629, N12612, N6283);
buf BUF1 (N12630, N12623);
not NOT1 (N12631, N12618);
not NOT1 (N12632, N12619);
or OR2 (N12633, N12621, N10237);
nand NAND3 (N12634, N12628, N3021, N12397);
nand NAND4 (N12635, N12627, N7374, N7023, N3431);
xor XOR2 (N12636, N12631, N11226);
not NOT1 (N12637, N12634);
not NOT1 (N12638, N12629);
nand NAND4 (N12639, N12633, N10054, N10707, N979);
or OR3 (N12640, N12636, N6127, N7392);
or OR2 (N12641, N12625, N10020);
xor XOR2 (N12642, N12635, N4694);
buf BUF1 (N12643, N12641);
or OR3 (N12644, N12632, N3509, N383);
xor XOR2 (N12645, N12642, N10552);
nor NOR3 (N12646, N12637, N6149, N6218);
buf BUF1 (N12647, N12624);
or OR4 (N12648, N12644, N976, N2601, N4629);
not NOT1 (N12649, N12646);
and AND4 (N12650, N12639, N1332, N2473, N1391);
xor XOR2 (N12651, N12647, N4449);
nand NAND2 (N12652, N12645, N2004);
xor XOR2 (N12653, N12638, N5029);
not NOT1 (N12654, N12650);
or OR2 (N12655, N12630, N12521);
not NOT1 (N12656, N12654);
xor XOR2 (N12657, N12656, N1598);
nor NOR4 (N12658, N12652, N7149, N11524, N5486);
xor XOR2 (N12659, N12640, N7075);
and AND4 (N12660, N12648, N2700, N7266, N6824);
nor NOR4 (N12661, N12658, N8316, N690, N6490);
and AND4 (N12662, N12657, N8310, N6555, N5271);
nor NOR4 (N12663, N12616, N492, N10629, N12081);
xor XOR2 (N12664, N12653, N6294);
buf BUF1 (N12665, N12655);
nand NAND3 (N12666, N12661, N8941, N1198);
or OR3 (N12667, N12662, N6283, N9322);
buf BUF1 (N12668, N12664);
or OR4 (N12669, N12666, N9759, N9423, N2392);
and AND3 (N12670, N12668, N2569, N1310);
nand NAND3 (N12671, N12659, N4667, N11345);
not NOT1 (N12672, N12660);
xor XOR2 (N12673, N12671, N12100);
not NOT1 (N12674, N12670);
nor NOR2 (N12675, N12663, N5854);
xor XOR2 (N12676, N12665, N8494);
nand NAND4 (N12677, N12667, N8717, N4950, N965);
or OR2 (N12678, N12675, N7792);
not NOT1 (N12679, N12649);
and AND3 (N12680, N12679, N1599, N9005);
nand NAND2 (N12681, N12651, N9095);
not NOT1 (N12682, N12669);
or OR3 (N12683, N12674, N11836, N8710);
nand NAND2 (N12684, N12680, N11828);
nor NOR3 (N12685, N12673, N1388, N8466);
and AND3 (N12686, N12676, N1991, N8650);
nor NOR3 (N12687, N12643, N3127, N471);
xor XOR2 (N12688, N12677, N790);
and AND3 (N12689, N12683, N6346, N11852);
nor NOR3 (N12690, N12689, N3069, N12354);
not NOT1 (N12691, N12678);
nand NAND4 (N12692, N12685, N4591, N3337, N5672);
nor NOR2 (N12693, N12682, N4052);
xor XOR2 (N12694, N12681, N123);
or OR4 (N12695, N12686, N4204, N5164, N10545);
nor NOR2 (N12696, N12693, N5815);
and AND3 (N12697, N12692, N3374, N9054);
or OR2 (N12698, N12695, N2111);
or OR3 (N12699, N12688, N4324, N10500);
or OR3 (N12700, N12672, N4416, N1507);
buf BUF1 (N12701, N12690);
not NOT1 (N12702, N12698);
nor NOR3 (N12703, N12684, N7682, N4534);
or OR3 (N12704, N12697, N6270, N7309);
nand NAND2 (N12705, N12703, N8692);
not NOT1 (N12706, N12687);
or OR4 (N12707, N12700, N691, N6303, N2727);
or OR3 (N12708, N12704, N3413, N2446);
and AND2 (N12709, N12691, N4992);
buf BUF1 (N12710, N12709);
nand NAND2 (N12711, N12701, N4931);
or OR2 (N12712, N12705, N7656);
nor NOR4 (N12713, N12706, N1026, N10768, N10298);
nor NOR3 (N12714, N12694, N4028, N9299);
or OR2 (N12715, N12712, N8412);
nand NAND4 (N12716, N12696, N2033, N7639, N10924);
nand NAND4 (N12717, N12699, N10510, N7008, N2988);
xor XOR2 (N12718, N12713, N3914);
nor NOR2 (N12719, N12710, N355);
nand NAND2 (N12720, N12715, N9888);
or OR2 (N12721, N12711, N945);
xor XOR2 (N12722, N12720, N6357);
or OR3 (N12723, N12718, N12265, N10451);
or OR3 (N12724, N12719, N5449, N4061);
not NOT1 (N12725, N12717);
xor XOR2 (N12726, N12707, N2066);
or OR4 (N12727, N12722, N4333, N5116, N6401);
not NOT1 (N12728, N12725);
and AND4 (N12729, N12724, N3416, N1783, N11707);
nor NOR2 (N12730, N12728, N7961);
or OR2 (N12731, N12702, N6725);
or OR3 (N12732, N12727, N9276, N1603);
buf BUF1 (N12733, N12723);
buf BUF1 (N12734, N12716);
nand NAND3 (N12735, N12721, N2596, N8178);
and AND3 (N12736, N12733, N11888, N1015);
xor XOR2 (N12737, N12731, N823);
and AND4 (N12738, N12729, N5127, N7358, N7330);
buf BUF1 (N12739, N12732);
nand NAND2 (N12740, N12726, N5565);
nor NOR2 (N12741, N12735, N7948);
nand NAND2 (N12742, N12736, N3509);
or OR2 (N12743, N12730, N5535);
or OR4 (N12744, N12741, N10762, N664, N1349);
nand NAND4 (N12745, N12708, N4468, N7727, N2561);
nor NOR4 (N12746, N12742, N7829, N3905, N6507);
not NOT1 (N12747, N12737);
not NOT1 (N12748, N12744);
not NOT1 (N12749, N12746);
not NOT1 (N12750, N12743);
not NOT1 (N12751, N12750);
buf BUF1 (N12752, N12745);
nor NOR3 (N12753, N12749, N7489, N4164);
buf BUF1 (N12754, N12748);
or OR4 (N12755, N12739, N6113, N7699, N12428);
buf BUF1 (N12756, N12738);
and AND2 (N12757, N12747, N12036);
not NOT1 (N12758, N12714);
and AND3 (N12759, N12755, N4795, N3170);
xor XOR2 (N12760, N12756, N3015);
nor NOR2 (N12761, N12754, N10462);
nand NAND4 (N12762, N12740, N6051, N428, N806);
not NOT1 (N12763, N12760);
xor XOR2 (N12764, N12757, N4877);
nor NOR2 (N12765, N12762, N4802);
xor XOR2 (N12766, N12734, N7886);
or OR3 (N12767, N12766, N7118, N11012);
nor NOR3 (N12768, N12764, N10417, N12214);
and AND4 (N12769, N12753, N124, N11949, N1209);
xor XOR2 (N12770, N12758, N10485);
not NOT1 (N12771, N12770);
and AND3 (N12772, N12751, N12216, N12642);
xor XOR2 (N12773, N12759, N11477);
buf BUF1 (N12774, N12767);
not NOT1 (N12775, N12771);
or OR4 (N12776, N12752, N6698, N1549, N3594);
nor NOR4 (N12777, N12774, N4168, N10794, N4666);
or OR2 (N12778, N12776, N3025);
nand NAND3 (N12779, N12773, N12577, N8191);
nand NAND2 (N12780, N12775, N5630);
nor NOR3 (N12781, N12761, N11929, N9438);
nand NAND3 (N12782, N12780, N5535, N1804);
and AND3 (N12783, N12781, N2961, N11690);
nand NAND3 (N12784, N12778, N4839, N2846);
buf BUF1 (N12785, N12763);
and AND2 (N12786, N12782, N516);
and AND4 (N12787, N12772, N9717, N12566, N4574);
buf BUF1 (N12788, N12783);
or OR4 (N12789, N12769, N675, N6430, N5595);
nand NAND3 (N12790, N12787, N7236, N12668);
or OR2 (N12791, N12790, N8851);
or OR2 (N12792, N12786, N4235);
nand NAND4 (N12793, N12765, N9625, N2592, N4699);
or OR4 (N12794, N12792, N1155, N657, N5382);
xor XOR2 (N12795, N12793, N3265);
not NOT1 (N12796, N12779);
nand NAND4 (N12797, N12795, N8611, N10711, N12407);
and AND2 (N12798, N12785, N9495);
nand NAND2 (N12799, N12794, N9360);
nand NAND4 (N12800, N12788, N1829, N11964, N11070);
xor XOR2 (N12801, N12796, N8627);
xor XOR2 (N12802, N12777, N10866);
and AND3 (N12803, N12768, N1583, N82);
and AND4 (N12804, N12789, N10259, N1127, N10450);
not NOT1 (N12805, N12801);
xor XOR2 (N12806, N12798, N11812);
xor XOR2 (N12807, N12799, N8551);
and AND3 (N12808, N12806, N100, N3186);
not NOT1 (N12809, N12791);
and AND2 (N12810, N12802, N12302);
xor XOR2 (N12811, N12800, N12228);
nor NOR4 (N12812, N12808, N11371, N8273, N1815);
not NOT1 (N12813, N12805);
buf BUF1 (N12814, N12784);
buf BUF1 (N12815, N12807);
xor XOR2 (N12816, N12813, N9411);
buf BUF1 (N12817, N12804);
nor NOR4 (N12818, N12815, N1655, N6831, N3300);
buf BUF1 (N12819, N12818);
nand NAND4 (N12820, N12814, N5670, N2277, N4456);
endmodule