// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N3205,N3189,N3210,N3199,N3208,N3192,N3212,N3213,N3214,N3215;

not NOT1 (N16, N3);
not NOT1 (N17, N13);
xor XOR2 (N18, N2, N10);
nor NOR2 (N19, N11, N10);
and AND2 (N20, N2, N2);
buf BUF1 (N21, N6);
nor NOR4 (N22, N8, N16, N6, N7);
or OR2 (N23, N22, N7);
buf BUF1 (N24, N4);
nor NOR2 (N25, N22, N21);
nand NAND2 (N26, N23, N15);
nor NOR4 (N27, N10, N13, N1, N1);
buf BUF1 (N28, N1);
and AND4 (N29, N17, N1, N5, N16);
not NOT1 (N30, N17);
buf BUF1 (N31, N30);
nand NAND2 (N32, N25, N20);
and AND2 (N33, N25, N29);
nand NAND2 (N34, N14, N9);
or OR2 (N35, N26, N20);
not NOT1 (N36, N33);
nand NAND3 (N37, N18, N31, N22);
nor NOR2 (N38, N16, N9);
buf BUF1 (N39, N35);
or OR3 (N40, N34, N33, N8);
not NOT1 (N41, N27);
xor XOR2 (N42, N38, N13);
xor XOR2 (N43, N19, N21);
xor XOR2 (N44, N28, N20);
and AND3 (N45, N37, N10, N27);
not NOT1 (N46, N39);
or OR3 (N47, N44, N41, N4);
nor NOR4 (N48, N28, N30, N12, N43);
not NOT1 (N49, N43);
nor NOR4 (N50, N42, N17, N13, N26);
xor XOR2 (N51, N45, N28);
nand NAND4 (N52, N51, N47, N27, N34);
and AND3 (N53, N14, N19, N3);
not NOT1 (N54, N24);
not NOT1 (N55, N46);
nor NOR4 (N56, N36, N51, N6, N19);
xor XOR2 (N57, N55, N25);
nand NAND2 (N58, N50, N49);
nor NOR2 (N59, N37, N20);
xor XOR2 (N60, N53, N46);
and AND3 (N61, N57, N19, N57);
nand NAND3 (N62, N32, N40, N22);
nor NOR2 (N63, N61, N34);
or OR4 (N64, N13, N48, N33, N43);
nand NAND2 (N65, N32, N59);
and AND3 (N66, N37, N17, N13);
xor XOR2 (N67, N52, N33);
nand NAND3 (N68, N58, N22, N46);
buf BUF1 (N69, N66);
xor XOR2 (N70, N54, N51);
not NOT1 (N71, N60);
buf BUF1 (N72, N69);
or OR4 (N73, N72, N7, N65, N61);
xor XOR2 (N74, N7, N25);
nor NOR4 (N75, N63, N69, N61, N50);
nand NAND4 (N76, N74, N31, N34, N55);
or OR3 (N77, N67, N49, N57);
buf BUF1 (N78, N70);
or OR3 (N79, N75, N10, N29);
nor NOR2 (N80, N68, N9);
not NOT1 (N81, N76);
not NOT1 (N82, N71);
not NOT1 (N83, N56);
and AND3 (N84, N82, N3, N39);
not NOT1 (N85, N78);
nand NAND3 (N86, N80, N37, N55);
xor XOR2 (N87, N81, N82);
or OR3 (N88, N85, N22, N36);
nand NAND3 (N89, N77, N70, N16);
and AND4 (N90, N79, N8, N30, N64);
xor XOR2 (N91, N85, N51);
xor XOR2 (N92, N86, N8);
nor NOR4 (N93, N83, N35, N38, N64);
xor XOR2 (N94, N84, N31);
or OR2 (N95, N90, N14);
nor NOR3 (N96, N94, N70, N87);
or OR3 (N97, N90, N49, N13);
or OR2 (N98, N97, N28);
and AND4 (N99, N62, N77, N10, N19);
buf BUF1 (N100, N73);
and AND3 (N101, N99, N97, N36);
buf BUF1 (N102, N95);
or OR3 (N103, N101, N11, N19);
buf BUF1 (N104, N92);
and AND3 (N105, N88, N87, N83);
not NOT1 (N106, N93);
not NOT1 (N107, N100);
and AND3 (N108, N102, N23, N66);
and AND3 (N109, N98, N63, N82);
not NOT1 (N110, N105);
xor XOR2 (N111, N104, N60);
not NOT1 (N112, N109);
nand NAND2 (N113, N106, N29);
not NOT1 (N114, N103);
buf BUF1 (N115, N113);
buf BUF1 (N116, N112);
or OR3 (N117, N89, N106, N60);
not NOT1 (N118, N111);
xor XOR2 (N119, N115, N61);
not NOT1 (N120, N96);
xor XOR2 (N121, N108, N13);
or OR3 (N122, N116, N117, N48);
not NOT1 (N123, N87);
xor XOR2 (N124, N110, N18);
xor XOR2 (N125, N114, N1);
nor NOR3 (N126, N118, N14, N64);
and AND2 (N127, N107, N69);
nand NAND2 (N128, N120, N15);
nand NAND3 (N129, N124, N66, N84);
xor XOR2 (N130, N119, N44);
and AND2 (N131, N129, N123);
xor XOR2 (N132, N31, N81);
or OR3 (N133, N127, N92, N28);
and AND4 (N134, N91, N44, N92, N22);
xor XOR2 (N135, N134, N124);
buf BUF1 (N136, N128);
nand NAND3 (N137, N131, N101, N28);
and AND4 (N138, N133, N114, N6, N55);
xor XOR2 (N139, N130, N113);
buf BUF1 (N140, N121);
not NOT1 (N141, N138);
xor XOR2 (N142, N122, N63);
or OR3 (N143, N142, N18, N116);
buf BUF1 (N144, N140);
nand NAND4 (N145, N143, N28, N106, N137);
xor XOR2 (N146, N4, N111);
or OR3 (N147, N139, N98, N91);
not NOT1 (N148, N132);
not NOT1 (N149, N147);
buf BUF1 (N150, N126);
nor NOR4 (N151, N148, N6, N33, N6);
nor NOR2 (N152, N141, N62);
buf BUF1 (N153, N149);
not NOT1 (N154, N136);
not NOT1 (N155, N144);
not NOT1 (N156, N154);
nor NOR3 (N157, N145, N87, N24);
buf BUF1 (N158, N125);
xor XOR2 (N159, N156, N7);
and AND3 (N160, N151, N22, N101);
or OR3 (N161, N146, N141, N8);
and AND4 (N162, N158, N107, N117, N98);
nor NOR3 (N163, N150, N77, N1);
nor NOR2 (N164, N152, N156);
xor XOR2 (N165, N157, N88);
nor NOR3 (N166, N162, N95, N61);
or OR4 (N167, N155, N140, N79, N75);
or OR4 (N168, N167, N7, N85, N93);
not NOT1 (N169, N160);
and AND3 (N170, N166, N145, N161);
and AND3 (N171, N51, N71, N61);
xor XOR2 (N172, N159, N137);
and AND3 (N173, N170, N109, N41);
nand NAND3 (N174, N168, N85, N60);
nand NAND3 (N175, N173, N154, N102);
and AND4 (N176, N165, N157, N67, N117);
or OR4 (N177, N175, N126, N30, N132);
not NOT1 (N178, N174);
xor XOR2 (N179, N176, N156);
not NOT1 (N180, N164);
nand NAND2 (N181, N163, N36);
nor NOR4 (N182, N180, N74, N163, N154);
nor NOR2 (N183, N177, N177);
xor XOR2 (N184, N135, N131);
xor XOR2 (N185, N172, N26);
xor XOR2 (N186, N153, N154);
and AND4 (N187, N185, N71, N72, N161);
and AND3 (N188, N178, N28, N30);
nor NOR3 (N189, N183, N172, N70);
and AND3 (N190, N186, N165, N188);
not NOT1 (N191, N136);
xor XOR2 (N192, N187, N46);
not NOT1 (N193, N184);
buf BUF1 (N194, N179);
xor XOR2 (N195, N169, N58);
xor XOR2 (N196, N189, N191);
nand NAND4 (N197, N153, N156, N109, N110);
xor XOR2 (N198, N193, N135);
nor NOR3 (N199, N194, N10, N56);
or OR2 (N200, N190, N171);
or OR2 (N201, N5, N164);
and AND3 (N202, N195, N81, N143);
or OR3 (N203, N200, N102, N50);
and AND4 (N204, N197, N144, N198, N174);
and AND3 (N205, N160, N111, N2);
not NOT1 (N206, N196);
xor XOR2 (N207, N192, N151);
and AND3 (N208, N207, N118, N181);
nand NAND3 (N209, N29, N18, N53);
buf BUF1 (N210, N201);
not NOT1 (N211, N202);
and AND4 (N212, N209, N80, N21, N99);
or OR4 (N213, N199, N110, N76, N11);
or OR3 (N214, N204, N189, N144);
not NOT1 (N215, N206);
not NOT1 (N216, N215);
or OR4 (N217, N211, N121, N119, N176);
nand NAND3 (N218, N216, N52, N141);
buf BUF1 (N219, N203);
buf BUF1 (N220, N182);
not NOT1 (N221, N212);
or OR2 (N222, N218, N104);
and AND4 (N223, N222, N93, N125, N188);
nand NAND4 (N224, N219, N185, N161, N59);
nor NOR3 (N225, N217, N106, N133);
or OR3 (N226, N205, N118, N42);
or OR3 (N227, N214, N118, N29);
and AND3 (N228, N213, N11, N208);
and AND3 (N229, N225, N141, N142);
and AND3 (N230, N136, N147, N147);
or OR4 (N231, N223, N127, N22, N175);
and AND2 (N232, N231, N49);
nand NAND3 (N233, N226, N135, N40);
nand NAND3 (N234, N230, N198, N20);
not NOT1 (N235, N221);
nand NAND2 (N236, N224, N136);
nand NAND4 (N237, N233, N219, N106, N32);
or OR2 (N238, N210, N129);
nor NOR3 (N239, N227, N144, N78);
and AND2 (N240, N237, N21);
not NOT1 (N241, N220);
xor XOR2 (N242, N239, N188);
or OR4 (N243, N229, N229, N179, N228);
nor NOR2 (N244, N73, N18);
or OR3 (N245, N236, N180, N142);
not NOT1 (N246, N238);
or OR3 (N247, N240, N193, N52);
not NOT1 (N248, N242);
and AND3 (N249, N235, N215, N10);
not NOT1 (N250, N247);
nor NOR4 (N251, N243, N202, N17, N39);
nor NOR4 (N252, N234, N97, N41, N74);
buf BUF1 (N253, N248);
nor NOR4 (N254, N244, N246, N142, N116);
nand NAND4 (N255, N95, N189, N101, N60);
nor NOR2 (N256, N249, N223);
xor XOR2 (N257, N251, N8);
buf BUF1 (N258, N255);
nand NAND4 (N259, N254, N248, N19, N95);
buf BUF1 (N260, N252);
xor XOR2 (N261, N241, N14);
xor XOR2 (N262, N253, N193);
buf BUF1 (N263, N260);
xor XOR2 (N264, N232, N42);
not NOT1 (N265, N250);
and AND2 (N266, N261, N156);
nor NOR4 (N267, N266, N262, N182, N10);
nor NOR4 (N268, N247, N145, N181, N146);
nand NAND3 (N269, N263, N198, N29);
or OR2 (N270, N245, N23);
nor NOR4 (N271, N269, N230, N105, N243);
or OR3 (N272, N264, N149, N105);
or OR2 (N273, N258, N266);
nor NOR3 (N274, N265, N174, N102);
not NOT1 (N275, N273);
xor XOR2 (N276, N257, N103);
or OR4 (N277, N274, N137, N151, N170);
and AND3 (N278, N275, N159, N170);
buf BUF1 (N279, N270);
and AND2 (N280, N256, N12);
xor XOR2 (N281, N268, N44);
xor XOR2 (N282, N279, N148);
xor XOR2 (N283, N281, N55);
or OR3 (N284, N278, N268, N145);
nor NOR2 (N285, N271, N143);
xor XOR2 (N286, N283, N267);
buf BUF1 (N287, N192);
nand NAND3 (N288, N282, N146, N230);
and AND2 (N289, N276, N112);
buf BUF1 (N290, N288);
xor XOR2 (N291, N286, N170);
not NOT1 (N292, N289);
buf BUF1 (N293, N272);
and AND4 (N294, N280, N122, N154, N89);
xor XOR2 (N295, N294, N150);
nor NOR4 (N296, N287, N232, N287, N255);
buf BUF1 (N297, N259);
and AND2 (N298, N295, N158);
nor NOR3 (N299, N293, N292, N73);
buf BUF1 (N300, N291);
nand NAND2 (N301, N282, N26);
xor XOR2 (N302, N284, N14);
not NOT1 (N303, N302);
xor XOR2 (N304, N285, N217);
or OR3 (N305, N303, N227, N168);
xor XOR2 (N306, N299, N254);
nand NAND3 (N307, N305, N81, N96);
buf BUF1 (N308, N304);
buf BUF1 (N309, N298);
or OR4 (N310, N306, N114, N218, N225);
xor XOR2 (N311, N277, N207);
nand NAND2 (N312, N297, N101);
buf BUF1 (N313, N310);
not NOT1 (N314, N309);
not NOT1 (N315, N312);
not NOT1 (N316, N315);
not NOT1 (N317, N308);
xor XOR2 (N318, N296, N188);
not NOT1 (N319, N318);
or OR2 (N320, N301, N213);
and AND4 (N321, N311, N145, N190, N140);
and AND3 (N322, N307, N76, N167);
or OR3 (N323, N317, N215, N5);
not NOT1 (N324, N322);
xor XOR2 (N325, N320, N209);
xor XOR2 (N326, N314, N86);
or OR2 (N327, N316, N322);
nand NAND2 (N328, N290, N200);
buf BUF1 (N329, N326);
not NOT1 (N330, N319);
xor XOR2 (N331, N321, N60);
buf BUF1 (N332, N323);
xor XOR2 (N333, N332, N244);
or OR3 (N334, N328, N239, N289);
nor NOR2 (N335, N329, N169);
xor XOR2 (N336, N300, N99);
xor XOR2 (N337, N313, N5);
or OR2 (N338, N334, N123);
nor NOR2 (N339, N336, N54);
and AND2 (N340, N331, N109);
nand NAND4 (N341, N324, N261, N94, N174);
and AND2 (N342, N330, N300);
xor XOR2 (N343, N335, N39);
and AND3 (N344, N339, N288, N157);
nor NOR3 (N345, N341, N45, N184);
and AND2 (N346, N327, N319);
nand NAND3 (N347, N337, N200, N287);
not NOT1 (N348, N338);
or OR2 (N349, N347, N177);
buf BUF1 (N350, N333);
or OR4 (N351, N350, N18, N80, N332);
nand NAND2 (N352, N346, N219);
nor NOR3 (N353, N352, N226, N146);
buf BUF1 (N354, N343);
nand NAND4 (N355, N348, N182, N56, N18);
nand NAND4 (N356, N325, N135, N288, N224);
xor XOR2 (N357, N342, N297);
nor NOR3 (N358, N353, N157, N274);
xor XOR2 (N359, N340, N348);
or OR4 (N360, N351, N195, N111, N189);
or OR3 (N361, N344, N272, N209);
or OR3 (N362, N358, N241, N50);
buf BUF1 (N363, N360);
and AND4 (N364, N361, N177, N227, N307);
or OR2 (N365, N364, N182);
xor XOR2 (N366, N357, N143);
buf BUF1 (N367, N363);
or OR3 (N368, N354, N258, N317);
buf BUF1 (N369, N355);
and AND4 (N370, N362, N362, N132, N252);
and AND3 (N371, N356, N330, N16);
not NOT1 (N372, N365);
and AND4 (N373, N366, N147, N90, N233);
and AND4 (N374, N349, N135, N269, N17);
nor NOR3 (N375, N373, N244, N221);
not NOT1 (N376, N372);
nor NOR2 (N377, N370, N190);
not NOT1 (N378, N375);
nor NOR3 (N379, N376, N359, N28);
nor NOR4 (N380, N325, N307, N51, N37);
nor NOR4 (N381, N378, N164, N215, N39);
and AND4 (N382, N374, N190, N153, N93);
xor XOR2 (N383, N345, N318);
and AND4 (N384, N381, N293, N193, N4);
xor XOR2 (N385, N380, N76);
xor XOR2 (N386, N384, N230);
and AND2 (N387, N367, N154);
not NOT1 (N388, N369);
buf BUF1 (N389, N368);
and AND2 (N390, N377, N27);
and AND3 (N391, N386, N162, N206);
xor XOR2 (N392, N390, N292);
xor XOR2 (N393, N389, N325);
or OR3 (N394, N392, N314, N165);
nand NAND4 (N395, N379, N355, N14, N73);
and AND3 (N396, N383, N326, N364);
and AND2 (N397, N396, N167);
and AND4 (N398, N388, N41, N184, N364);
nor NOR4 (N399, N391, N266, N199, N258);
and AND3 (N400, N382, N314, N224);
or OR2 (N401, N394, N202);
or OR2 (N402, N395, N130);
or OR3 (N403, N401, N293, N183);
nor NOR3 (N404, N402, N293, N402);
nand NAND3 (N405, N399, N403, N351);
nand NAND3 (N406, N137, N234, N72);
nand NAND2 (N407, N385, N113);
nand NAND3 (N408, N371, N93, N283);
not NOT1 (N409, N408);
nor NOR3 (N410, N397, N260, N372);
and AND2 (N411, N406, N152);
not NOT1 (N412, N409);
nand NAND4 (N413, N405, N128, N321, N185);
buf BUF1 (N414, N404);
and AND4 (N415, N411, N334, N29, N414);
xor XOR2 (N416, N246, N104);
buf BUF1 (N417, N415);
buf BUF1 (N418, N393);
or OR2 (N419, N416, N248);
not NOT1 (N420, N418);
buf BUF1 (N421, N412);
nor NOR2 (N422, N410, N339);
nand NAND3 (N423, N421, N287, N226);
or OR2 (N424, N423, N255);
xor XOR2 (N425, N419, N113);
not NOT1 (N426, N417);
buf BUF1 (N427, N407);
xor XOR2 (N428, N400, N164);
and AND4 (N429, N387, N270, N321, N106);
and AND4 (N430, N429, N212, N114, N107);
nand NAND3 (N431, N425, N20, N333);
not NOT1 (N432, N424);
nor NOR3 (N433, N428, N293, N194);
xor XOR2 (N434, N426, N231);
nor NOR4 (N435, N427, N383, N411, N389);
and AND3 (N436, N434, N55, N34);
buf BUF1 (N437, N420);
or OR2 (N438, N430, N301);
xor XOR2 (N439, N431, N258);
xor XOR2 (N440, N398, N189);
not NOT1 (N441, N432);
xor XOR2 (N442, N435, N89);
or OR4 (N443, N436, N381, N176, N215);
or OR2 (N444, N433, N72);
not NOT1 (N445, N413);
xor XOR2 (N446, N440, N112);
or OR3 (N447, N445, N158, N360);
and AND4 (N448, N437, N239, N349, N305);
not NOT1 (N449, N443);
or OR4 (N450, N442, N303, N220, N399);
xor XOR2 (N451, N448, N15);
buf BUF1 (N452, N441);
and AND2 (N453, N446, N272);
xor XOR2 (N454, N449, N261);
xor XOR2 (N455, N438, N253);
buf BUF1 (N456, N450);
and AND3 (N457, N454, N413, N79);
and AND4 (N458, N451, N416, N309, N99);
and AND4 (N459, N457, N196, N71, N282);
nand NAND2 (N460, N459, N352);
and AND2 (N461, N458, N331);
nand NAND3 (N462, N456, N310, N211);
buf BUF1 (N463, N444);
nand NAND4 (N464, N462, N95, N401, N316);
and AND3 (N465, N455, N55, N449);
and AND4 (N466, N439, N148, N391, N52);
nor NOR3 (N467, N463, N366, N63);
buf BUF1 (N468, N447);
nor NOR2 (N469, N467, N76);
buf BUF1 (N470, N466);
and AND3 (N471, N465, N27, N372);
xor XOR2 (N472, N461, N467);
buf BUF1 (N473, N452);
buf BUF1 (N474, N422);
buf BUF1 (N475, N471);
or OR3 (N476, N474, N24, N88);
and AND3 (N477, N476, N295, N132);
not NOT1 (N478, N464);
or OR4 (N479, N460, N250, N312, N13);
and AND2 (N480, N478, N371);
buf BUF1 (N481, N475);
and AND3 (N482, N481, N337, N310);
nor NOR4 (N483, N472, N431, N86, N365);
not NOT1 (N484, N482);
and AND4 (N485, N469, N64, N217, N428);
or OR2 (N486, N468, N412);
buf BUF1 (N487, N473);
and AND3 (N488, N485, N91, N459);
not NOT1 (N489, N483);
and AND4 (N490, N488, N226, N270, N471);
not NOT1 (N491, N490);
xor XOR2 (N492, N489, N88);
and AND4 (N493, N479, N323, N448, N104);
or OR3 (N494, N487, N470, N34);
not NOT1 (N495, N168);
nor NOR4 (N496, N493, N141, N424, N254);
buf BUF1 (N497, N453);
xor XOR2 (N498, N486, N99);
not NOT1 (N499, N477);
buf BUF1 (N500, N499);
or OR3 (N501, N480, N69, N21);
not NOT1 (N502, N501);
or OR2 (N503, N495, N282);
not NOT1 (N504, N496);
nor NOR4 (N505, N498, N334, N113, N356);
xor XOR2 (N506, N505, N315);
or OR4 (N507, N491, N297, N304, N308);
and AND4 (N508, N494, N133, N107, N437);
nor NOR4 (N509, N507, N346, N393, N225);
not NOT1 (N510, N502);
buf BUF1 (N511, N492);
or OR3 (N512, N504, N72, N320);
nand NAND3 (N513, N503, N476, N149);
or OR3 (N514, N506, N342, N160);
or OR4 (N515, N512, N397, N484, N164);
buf BUF1 (N516, N318);
not NOT1 (N517, N510);
xor XOR2 (N518, N515, N302);
not NOT1 (N519, N508);
not NOT1 (N520, N514);
nand NAND2 (N521, N497, N228);
nand NAND2 (N522, N500, N366);
buf BUF1 (N523, N513);
or OR2 (N524, N522, N107);
and AND3 (N525, N516, N391, N451);
not NOT1 (N526, N518);
and AND4 (N527, N521, N96, N377, N16);
nor NOR2 (N528, N523, N294);
not NOT1 (N529, N511);
xor XOR2 (N530, N519, N398);
or OR4 (N531, N517, N204, N253, N434);
not NOT1 (N532, N527);
buf BUF1 (N533, N526);
not NOT1 (N534, N509);
nor NOR4 (N535, N533, N231, N370, N222);
not NOT1 (N536, N529);
not NOT1 (N537, N525);
and AND2 (N538, N534, N168);
not NOT1 (N539, N520);
or OR4 (N540, N528, N261, N286, N264);
buf BUF1 (N541, N535);
buf BUF1 (N542, N537);
not NOT1 (N543, N531);
nor NOR4 (N544, N530, N199, N355, N389);
or OR2 (N545, N539, N382);
or OR2 (N546, N538, N14);
xor XOR2 (N547, N545, N394);
nor NOR2 (N548, N543, N61);
nor NOR4 (N549, N541, N165, N165, N348);
or OR3 (N550, N549, N304, N545);
nand NAND2 (N551, N548, N137);
buf BUF1 (N552, N536);
nor NOR3 (N553, N546, N109, N427);
nor NOR4 (N554, N550, N285, N343, N467);
nand NAND2 (N555, N547, N52);
or OR3 (N556, N542, N502, N320);
nor NOR3 (N557, N554, N343, N361);
nand NAND2 (N558, N557, N85);
not NOT1 (N559, N524);
and AND3 (N560, N551, N542, N405);
buf BUF1 (N561, N559);
nand NAND3 (N562, N552, N33, N322);
or OR2 (N563, N556, N314);
or OR4 (N564, N553, N303, N23, N241);
not NOT1 (N565, N560);
xor XOR2 (N566, N555, N158);
buf BUF1 (N567, N532);
xor XOR2 (N568, N562, N251);
not NOT1 (N569, N544);
nor NOR4 (N570, N558, N308, N64, N482);
nor NOR2 (N571, N566, N505);
not NOT1 (N572, N569);
not NOT1 (N573, N564);
not NOT1 (N574, N565);
not NOT1 (N575, N573);
nand NAND2 (N576, N567, N10);
not NOT1 (N577, N574);
and AND3 (N578, N570, N149, N275);
nand NAND4 (N579, N577, N173, N30, N444);
not NOT1 (N580, N563);
nor NOR3 (N581, N579, N63, N487);
buf BUF1 (N582, N540);
not NOT1 (N583, N581);
xor XOR2 (N584, N571, N478);
xor XOR2 (N585, N583, N563);
xor XOR2 (N586, N580, N434);
not NOT1 (N587, N585);
nand NAND4 (N588, N586, N276, N6, N129);
or OR2 (N589, N588, N299);
or OR3 (N590, N576, N231, N1);
nor NOR4 (N591, N590, N268, N467, N7);
and AND4 (N592, N578, N39, N58, N138);
and AND3 (N593, N572, N358, N517);
xor XOR2 (N594, N584, N459);
or OR2 (N595, N568, N82);
or OR2 (N596, N582, N517);
or OR3 (N597, N561, N327, N253);
xor XOR2 (N598, N592, N287);
and AND2 (N599, N593, N98);
buf BUF1 (N600, N594);
and AND4 (N601, N591, N372, N588, N540);
nor NOR2 (N602, N596, N44);
nand NAND4 (N603, N587, N80, N409, N231);
xor XOR2 (N604, N598, N464);
and AND3 (N605, N599, N355, N538);
nand NAND2 (N606, N600, N38);
and AND2 (N607, N605, N85);
nor NOR2 (N608, N603, N270);
xor XOR2 (N609, N595, N56);
or OR3 (N610, N609, N338, N455);
not NOT1 (N611, N607);
nor NOR4 (N612, N610, N139, N216, N274);
and AND4 (N613, N608, N512, N368, N496);
not NOT1 (N614, N601);
nand NAND3 (N615, N604, N162, N514);
nor NOR2 (N616, N597, N562);
xor XOR2 (N617, N575, N398);
nand NAND3 (N618, N615, N419, N416);
or OR3 (N619, N606, N578, N222);
nor NOR4 (N620, N616, N92, N74, N99);
nor NOR4 (N621, N618, N57, N269, N611);
and AND2 (N622, N533, N510);
buf BUF1 (N623, N612);
and AND2 (N624, N621, N516);
buf BUF1 (N625, N613);
nand NAND2 (N626, N619, N619);
not NOT1 (N627, N617);
nor NOR2 (N628, N620, N312);
nor NOR2 (N629, N623, N174);
nor NOR4 (N630, N614, N335, N513, N378);
or OR4 (N631, N589, N573, N510, N583);
and AND4 (N632, N629, N316, N81, N496);
buf BUF1 (N633, N624);
nor NOR3 (N634, N602, N380, N177);
not NOT1 (N635, N626);
and AND3 (N636, N635, N494, N271);
nand NAND3 (N637, N622, N328, N82);
and AND4 (N638, N627, N179, N484, N198);
or OR3 (N639, N638, N445, N6);
or OR4 (N640, N637, N208, N363, N466);
or OR4 (N641, N631, N167, N504, N197);
or OR3 (N642, N640, N600, N34);
nor NOR2 (N643, N642, N187);
and AND2 (N644, N639, N394);
and AND4 (N645, N643, N400, N561, N539);
nand NAND2 (N646, N628, N600);
buf BUF1 (N647, N630);
not NOT1 (N648, N634);
nor NOR4 (N649, N644, N292, N417, N636);
not NOT1 (N650, N443);
and AND2 (N651, N645, N267);
not NOT1 (N652, N641);
xor XOR2 (N653, N652, N271);
and AND2 (N654, N651, N43);
nand NAND2 (N655, N653, N358);
buf BUF1 (N656, N646);
not NOT1 (N657, N633);
and AND3 (N658, N632, N151, N216);
xor XOR2 (N659, N649, N24);
not NOT1 (N660, N650);
nor NOR3 (N661, N660, N71, N44);
nand NAND2 (N662, N658, N156);
nand NAND3 (N663, N648, N404, N301);
or OR4 (N664, N656, N384, N519, N534);
or OR4 (N665, N659, N488, N196, N234);
or OR3 (N666, N654, N140, N80);
nor NOR4 (N667, N647, N211, N542, N643);
xor XOR2 (N668, N661, N8);
buf BUF1 (N669, N664);
buf BUF1 (N670, N662);
or OR4 (N671, N670, N647, N317, N148);
and AND4 (N672, N671, N302, N666, N478);
not NOT1 (N673, N83);
nand NAND3 (N674, N673, N154, N43);
nand NAND2 (N675, N663, N277);
buf BUF1 (N676, N668);
nand NAND4 (N677, N655, N163, N352, N612);
nand NAND3 (N678, N657, N39, N452);
nand NAND4 (N679, N625, N368, N296, N340);
and AND3 (N680, N669, N364, N675);
not NOT1 (N681, N464);
xor XOR2 (N682, N678, N48);
buf BUF1 (N683, N665);
nor NOR2 (N684, N676, N339);
nand NAND4 (N685, N667, N19, N172, N599);
nor NOR4 (N686, N677, N372, N49, N521);
buf BUF1 (N687, N682);
and AND3 (N688, N679, N75, N202);
not NOT1 (N689, N687);
nand NAND4 (N690, N680, N68, N519, N58);
nor NOR4 (N691, N689, N453, N679, N161);
and AND4 (N692, N685, N327, N89, N139);
xor XOR2 (N693, N691, N445);
nor NOR3 (N694, N674, N10, N164);
nand NAND3 (N695, N693, N96, N689);
and AND2 (N696, N694, N217);
not NOT1 (N697, N684);
buf BUF1 (N698, N695);
not NOT1 (N699, N698);
not NOT1 (N700, N697);
nor NOR4 (N701, N686, N582, N228, N541);
buf BUF1 (N702, N672);
nor NOR2 (N703, N700, N100);
nor NOR4 (N704, N701, N283, N615, N226);
xor XOR2 (N705, N704, N198);
nand NAND2 (N706, N705, N558);
or OR2 (N707, N688, N405);
not NOT1 (N708, N690);
xor XOR2 (N709, N708, N425);
xor XOR2 (N710, N681, N409);
not NOT1 (N711, N706);
nand NAND4 (N712, N692, N316, N202, N451);
nand NAND4 (N713, N696, N79, N10, N658);
nor NOR3 (N714, N712, N671, N155);
and AND2 (N715, N699, N493);
nand NAND4 (N716, N714, N611, N537, N361);
and AND3 (N717, N702, N335, N608);
not NOT1 (N718, N709);
buf BUF1 (N719, N715);
xor XOR2 (N720, N717, N66);
not NOT1 (N721, N683);
buf BUF1 (N722, N716);
not NOT1 (N723, N713);
xor XOR2 (N724, N718, N346);
or OR3 (N725, N703, N272, N414);
or OR4 (N726, N719, N195, N465, N54);
nor NOR4 (N727, N722, N533, N274, N12);
not NOT1 (N728, N710);
buf BUF1 (N729, N727);
xor XOR2 (N730, N725, N223);
or OR2 (N731, N721, N459);
or OR3 (N732, N723, N323, N328);
or OR2 (N733, N732, N526);
nand NAND4 (N734, N731, N645, N57, N725);
nand NAND4 (N735, N711, N380, N95, N649);
buf BUF1 (N736, N728);
nand NAND2 (N737, N736, N592);
and AND3 (N738, N737, N116, N100);
xor XOR2 (N739, N734, N281);
and AND4 (N740, N724, N76, N274, N616);
nor NOR2 (N741, N738, N616);
nor NOR4 (N742, N720, N31, N298, N660);
not NOT1 (N743, N729);
buf BUF1 (N744, N742);
nand NAND2 (N745, N739, N27);
xor XOR2 (N746, N735, N29);
buf BUF1 (N747, N744);
nor NOR3 (N748, N730, N509, N623);
or OR3 (N749, N743, N736, N234);
or OR2 (N750, N749, N567);
not NOT1 (N751, N745);
xor XOR2 (N752, N751, N84);
xor XOR2 (N753, N707, N182);
xor XOR2 (N754, N747, N185);
and AND4 (N755, N748, N281, N725, N467);
nor NOR3 (N756, N752, N337, N720);
nand NAND2 (N757, N733, N48);
xor XOR2 (N758, N753, N480);
buf BUF1 (N759, N740);
and AND2 (N760, N741, N686);
nand NAND4 (N761, N759, N402, N319, N308);
nor NOR3 (N762, N755, N719, N176);
xor XOR2 (N763, N726, N340);
nor NOR4 (N764, N746, N509, N376, N547);
xor XOR2 (N765, N756, N132);
buf BUF1 (N766, N757);
not NOT1 (N767, N750);
buf BUF1 (N768, N754);
nor NOR3 (N769, N765, N253, N468);
buf BUF1 (N770, N763);
buf BUF1 (N771, N768);
xor XOR2 (N772, N758, N542);
xor XOR2 (N773, N771, N17);
or OR3 (N774, N769, N584, N447);
not NOT1 (N775, N767);
xor XOR2 (N776, N775, N612);
nor NOR4 (N777, N766, N212, N764, N45);
buf BUF1 (N778, N335);
buf BUF1 (N779, N761);
not NOT1 (N780, N770);
xor XOR2 (N781, N760, N420);
not NOT1 (N782, N780);
or OR3 (N783, N762, N725, N147);
not NOT1 (N784, N783);
buf BUF1 (N785, N784);
nand NAND3 (N786, N777, N459, N647);
and AND3 (N787, N781, N437, N89);
nor NOR3 (N788, N772, N388, N271);
not NOT1 (N789, N773);
buf BUF1 (N790, N782);
nand NAND4 (N791, N789, N621, N293, N295);
nor NOR3 (N792, N785, N399, N579);
and AND3 (N793, N792, N702, N82);
nand NAND4 (N794, N779, N210, N311, N104);
xor XOR2 (N795, N793, N726);
nor NOR4 (N796, N790, N539, N495, N688);
and AND3 (N797, N796, N49, N748);
buf BUF1 (N798, N786);
or OR4 (N799, N774, N550, N374, N187);
and AND2 (N800, N799, N54);
not NOT1 (N801, N788);
nor NOR2 (N802, N787, N571);
and AND3 (N803, N776, N763, N182);
nor NOR3 (N804, N791, N685, N677);
buf BUF1 (N805, N803);
and AND2 (N806, N805, N485);
nand NAND3 (N807, N795, N780, N191);
nor NOR2 (N808, N801, N473);
not NOT1 (N809, N804);
buf BUF1 (N810, N808);
xor XOR2 (N811, N807, N139);
and AND2 (N812, N800, N91);
and AND4 (N813, N812, N6, N189, N735);
or OR4 (N814, N778, N228, N101, N796);
nor NOR2 (N815, N794, N421);
or OR2 (N816, N806, N482);
not NOT1 (N817, N815);
nor NOR3 (N818, N810, N175, N383);
buf BUF1 (N819, N813);
not NOT1 (N820, N798);
nor NOR4 (N821, N814, N547, N749, N160);
xor XOR2 (N822, N816, N22);
nand NAND2 (N823, N822, N91);
or OR2 (N824, N811, N588);
xor XOR2 (N825, N797, N213);
nand NAND2 (N826, N824, N137);
or OR4 (N827, N826, N655, N518, N638);
nand NAND2 (N828, N819, N248);
xor XOR2 (N829, N823, N774);
not NOT1 (N830, N809);
not NOT1 (N831, N828);
nor NOR2 (N832, N821, N427);
buf BUF1 (N833, N802);
buf BUF1 (N834, N820);
nand NAND2 (N835, N829, N93);
nor NOR3 (N836, N825, N244, N576);
buf BUF1 (N837, N834);
not NOT1 (N838, N830);
xor XOR2 (N839, N836, N377);
buf BUF1 (N840, N837);
or OR2 (N841, N835, N652);
not NOT1 (N842, N818);
not NOT1 (N843, N839);
nand NAND4 (N844, N841, N168, N219, N545);
nor NOR4 (N845, N844, N331, N319, N742);
buf BUF1 (N846, N831);
xor XOR2 (N847, N827, N576);
xor XOR2 (N848, N832, N649);
nor NOR2 (N849, N840, N681);
nor NOR2 (N850, N838, N410);
xor XOR2 (N851, N850, N433);
not NOT1 (N852, N846);
xor XOR2 (N853, N845, N149);
not NOT1 (N854, N843);
xor XOR2 (N855, N852, N12);
not NOT1 (N856, N853);
nor NOR4 (N857, N847, N158, N704, N213);
buf BUF1 (N858, N849);
not NOT1 (N859, N842);
not NOT1 (N860, N854);
nand NAND4 (N861, N817, N385, N437, N770);
xor XOR2 (N862, N851, N265);
nor NOR4 (N863, N860, N71, N269, N28);
nand NAND2 (N864, N862, N75);
or OR3 (N865, N864, N755, N316);
buf BUF1 (N866, N859);
xor XOR2 (N867, N863, N15);
nand NAND2 (N868, N857, N205);
nor NOR2 (N869, N868, N772);
or OR2 (N870, N867, N55);
nor NOR4 (N871, N866, N58, N615, N88);
not NOT1 (N872, N871);
and AND3 (N873, N858, N103, N770);
or OR3 (N874, N848, N816, N544);
nor NOR2 (N875, N855, N313);
xor XOR2 (N876, N861, N157);
not NOT1 (N877, N876);
not NOT1 (N878, N873);
nor NOR2 (N879, N872, N81);
not NOT1 (N880, N875);
and AND2 (N881, N877, N330);
buf BUF1 (N882, N856);
buf BUF1 (N883, N880);
nor NOR3 (N884, N833, N470, N101);
buf BUF1 (N885, N878);
xor XOR2 (N886, N882, N674);
nor NOR4 (N887, N870, N515, N329, N36);
buf BUF1 (N888, N885);
not NOT1 (N889, N881);
xor XOR2 (N890, N869, N367);
xor XOR2 (N891, N879, N340);
xor XOR2 (N892, N883, N776);
nand NAND3 (N893, N891, N365, N227);
and AND2 (N894, N893, N138);
nand NAND3 (N895, N865, N465, N655);
xor XOR2 (N896, N892, N218);
nor NOR3 (N897, N884, N812, N247);
and AND4 (N898, N895, N637, N612, N431);
nand NAND2 (N899, N894, N403);
xor XOR2 (N900, N874, N385);
buf BUF1 (N901, N900);
xor XOR2 (N902, N888, N696);
buf BUF1 (N903, N889);
xor XOR2 (N904, N890, N663);
buf BUF1 (N905, N887);
and AND3 (N906, N905, N610, N408);
buf BUF1 (N907, N896);
and AND2 (N908, N903, N408);
buf BUF1 (N909, N897);
not NOT1 (N910, N904);
xor XOR2 (N911, N899, N108);
nor NOR4 (N912, N906, N221, N312, N499);
or OR4 (N913, N886, N384, N318, N29);
xor XOR2 (N914, N901, N501);
and AND4 (N915, N907, N13, N117, N346);
and AND2 (N916, N909, N257);
not NOT1 (N917, N902);
xor XOR2 (N918, N911, N334);
buf BUF1 (N919, N898);
not NOT1 (N920, N910);
not NOT1 (N921, N917);
or OR3 (N922, N916, N365, N541);
or OR3 (N923, N921, N719, N552);
nor NOR2 (N924, N913, N59);
and AND2 (N925, N919, N700);
not NOT1 (N926, N918);
not NOT1 (N927, N912);
not NOT1 (N928, N915);
nand NAND3 (N929, N926, N86, N876);
not NOT1 (N930, N908);
nand NAND3 (N931, N930, N779, N659);
and AND3 (N932, N927, N57, N526);
xor XOR2 (N933, N923, N382);
or OR2 (N934, N933, N852);
nor NOR3 (N935, N914, N317, N352);
not NOT1 (N936, N922);
nand NAND4 (N937, N935, N452, N710, N709);
buf BUF1 (N938, N931);
and AND2 (N939, N929, N454);
nor NOR2 (N940, N938, N872);
buf BUF1 (N941, N932);
nand NAND4 (N942, N928, N367, N841, N529);
nand NAND4 (N943, N939, N624, N906, N867);
not NOT1 (N944, N934);
or OR3 (N945, N920, N201, N657);
xor XOR2 (N946, N936, N362);
buf BUF1 (N947, N944);
or OR2 (N948, N941, N316);
nand NAND3 (N949, N937, N258, N785);
and AND3 (N950, N946, N326, N34);
and AND4 (N951, N948, N487, N698, N421);
not NOT1 (N952, N947);
not NOT1 (N953, N951);
buf BUF1 (N954, N942);
or OR3 (N955, N954, N939, N305);
xor XOR2 (N956, N945, N598);
or OR4 (N957, N943, N729, N734, N138);
nand NAND3 (N958, N955, N369, N133);
or OR3 (N959, N953, N372, N825);
and AND4 (N960, N958, N338, N285, N776);
nand NAND3 (N961, N957, N47, N122);
xor XOR2 (N962, N952, N416);
xor XOR2 (N963, N962, N479);
nor NOR4 (N964, N949, N166, N547, N42);
not NOT1 (N965, N964);
buf BUF1 (N966, N965);
not NOT1 (N967, N963);
or OR3 (N968, N950, N666, N594);
nor NOR4 (N969, N924, N600, N749, N509);
xor XOR2 (N970, N960, N293);
buf BUF1 (N971, N970);
nor NOR3 (N972, N969, N419, N405);
and AND3 (N973, N972, N783, N149);
or OR4 (N974, N967, N369, N653, N637);
buf BUF1 (N975, N925);
or OR4 (N976, N975, N373, N921, N587);
and AND3 (N977, N961, N698, N531);
nand NAND3 (N978, N940, N646, N100);
xor XOR2 (N979, N959, N946);
nand NAND2 (N980, N968, N771);
nor NOR4 (N981, N977, N474, N616, N622);
or OR3 (N982, N966, N511, N681);
xor XOR2 (N983, N973, N888);
and AND2 (N984, N974, N945);
nor NOR2 (N985, N979, N460);
and AND2 (N986, N976, N286);
buf BUF1 (N987, N986);
nand NAND3 (N988, N982, N819, N779);
nand NAND4 (N989, N984, N578, N550, N785);
not NOT1 (N990, N988);
and AND3 (N991, N980, N42, N301);
xor XOR2 (N992, N985, N279);
not NOT1 (N993, N983);
nor NOR4 (N994, N971, N759, N46, N919);
not NOT1 (N995, N978);
nand NAND4 (N996, N981, N268, N890, N302);
xor XOR2 (N997, N987, N647);
nand NAND2 (N998, N995, N483);
xor XOR2 (N999, N989, N688);
and AND4 (N1000, N997, N405, N864, N146);
nand NAND4 (N1001, N993, N687, N513, N791);
or OR4 (N1002, N994, N888, N572, N745);
xor XOR2 (N1003, N998, N738);
buf BUF1 (N1004, N1003);
nand NAND2 (N1005, N991, N856);
xor XOR2 (N1006, N1004, N225);
nor NOR2 (N1007, N1000, N81);
not NOT1 (N1008, N990);
buf BUF1 (N1009, N996);
and AND2 (N1010, N1008, N205);
and AND4 (N1011, N1001, N829, N994, N978);
xor XOR2 (N1012, N956, N12);
nor NOR3 (N1013, N1009, N688, N868);
xor XOR2 (N1014, N1012, N744);
not NOT1 (N1015, N1002);
not NOT1 (N1016, N1014);
or OR2 (N1017, N1016, N577);
nor NOR4 (N1018, N999, N850, N709, N1011);
nor NOR2 (N1019, N993, N664);
nor NOR3 (N1020, N1015, N960, N220);
buf BUF1 (N1021, N1007);
not NOT1 (N1022, N1021);
nand NAND3 (N1023, N1013, N223, N129);
not NOT1 (N1024, N1020);
buf BUF1 (N1025, N1024);
or OR2 (N1026, N1017, N940);
buf BUF1 (N1027, N1018);
nor NOR2 (N1028, N1005, N656);
nand NAND4 (N1029, N1027, N674, N214, N790);
and AND4 (N1030, N1019, N681, N487, N726);
nor NOR3 (N1031, N1028, N170, N799);
xor XOR2 (N1032, N1026, N258);
and AND4 (N1033, N1010, N780, N785, N544);
not NOT1 (N1034, N1025);
nand NAND2 (N1035, N1030, N43);
nor NOR4 (N1036, N1033, N471, N807, N755);
not NOT1 (N1037, N1032);
nor NOR3 (N1038, N1031, N816, N601);
and AND2 (N1039, N1034, N325);
or OR4 (N1040, N1039, N406, N1019, N559);
and AND3 (N1041, N1040, N705, N51);
and AND4 (N1042, N1022, N977, N271, N127);
buf BUF1 (N1043, N1042);
buf BUF1 (N1044, N1041);
nor NOR4 (N1045, N1044, N596, N1001, N433);
not NOT1 (N1046, N1037);
nor NOR3 (N1047, N1045, N1010, N610);
and AND3 (N1048, N1036, N896, N185);
nand NAND4 (N1049, N992, N597, N870, N208);
and AND2 (N1050, N1029, N298);
buf BUF1 (N1051, N1038);
and AND2 (N1052, N1046, N420);
or OR4 (N1053, N1043, N214, N222, N905);
not NOT1 (N1054, N1035);
nand NAND4 (N1055, N1049, N211, N828, N897);
and AND2 (N1056, N1006, N995);
buf BUF1 (N1057, N1051);
nand NAND4 (N1058, N1054, N969, N890, N64);
or OR2 (N1059, N1048, N734);
nand NAND2 (N1060, N1023, N527);
xor XOR2 (N1061, N1060, N754);
and AND3 (N1062, N1053, N734, N128);
nand NAND2 (N1063, N1061, N814);
not NOT1 (N1064, N1056);
nor NOR4 (N1065, N1058, N143, N869, N718);
xor XOR2 (N1066, N1063, N819);
xor XOR2 (N1067, N1055, N312);
or OR2 (N1068, N1059, N573);
nand NAND3 (N1069, N1068, N769, N731);
and AND2 (N1070, N1050, N242);
nand NAND4 (N1071, N1065, N504, N300, N546);
not NOT1 (N1072, N1071);
buf BUF1 (N1073, N1062);
xor XOR2 (N1074, N1052, N1025);
nand NAND2 (N1075, N1070, N343);
buf BUF1 (N1076, N1067);
or OR4 (N1077, N1074, N917, N171, N170);
and AND2 (N1078, N1047, N994);
buf BUF1 (N1079, N1073);
buf BUF1 (N1080, N1078);
buf BUF1 (N1081, N1077);
buf BUF1 (N1082, N1064);
or OR3 (N1083, N1082, N598, N973);
not NOT1 (N1084, N1079);
nor NOR2 (N1085, N1057, N303);
not NOT1 (N1086, N1072);
not NOT1 (N1087, N1085);
not NOT1 (N1088, N1066);
and AND3 (N1089, N1087, N468, N805);
and AND4 (N1090, N1086, N971, N831, N673);
xor XOR2 (N1091, N1080, N337);
buf BUF1 (N1092, N1083);
buf BUF1 (N1093, N1076);
buf BUF1 (N1094, N1075);
xor XOR2 (N1095, N1089, N634);
not NOT1 (N1096, N1092);
nor NOR2 (N1097, N1088, N676);
not NOT1 (N1098, N1094);
not NOT1 (N1099, N1098);
nor NOR2 (N1100, N1099, N55);
and AND4 (N1101, N1084, N832, N18, N835);
or OR3 (N1102, N1101, N526, N1025);
not NOT1 (N1103, N1091);
nor NOR2 (N1104, N1103, N452);
and AND3 (N1105, N1093, N284, N1005);
or OR3 (N1106, N1090, N1079, N319);
nand NAND4 (N1107, N1100, N551, N103, N970);
xor XOR2 (N1108, N1096, N42);
and AND3 (N1109, N1108, N175, N1008);
not NOT1 (N1110, N1105);
and AND4 (N1111, N1095, N79, N571, N266);
nand NAND4 (N1112, N1107, N360, N709, N511);
nand NAND4 (N1113, N1111, N883, N385, N915);
not NOT1 (N1114, N1109);
or OR3 (N1115, N1114, N295, N1007);
not NOT1 (N1116, N1104);
or OR3 (N1117, N1113, N262, N898);
or OR2 (N1118, N1112, N707);
buf BUF1 (N1119, N1116);
not NOT1 (N1120, N1102);
nand NAND2 (N1121, N1115, N1118);
buf BUF1 (N1122, N1044);
or OR4 (N1123, N1097, N330, N906, N516);
or OR3 (N1124, N1110, N816, N301);
nor NOR3 (N1125, N1122, N957, N377);
xor XOR2 (N1126, N1120, N292);
nor NOR4 (N1127, N1069, N988, N218, N975);
nand NAND4 (N1128, N1126, N768, N289, N864);
xor XOR2 (N1129, N1117, N426);
nand NAND2 (N1130, N1123, N173);
nor NOR3 (N1131, N1130, N827, N138);
xor XOR2 (N1132, N1106, N1118);
or OR4 (N1133, N1132, N725, N845, N561);
buf BUF1 (N1134, N1124);
nand NAND2 (N1135, N1125, N697);
and AND3 (N1136, N1081, N13, N1033);
buf BUF1 (N1137, N1127);
xor XOR2 (N1138, N1119, N76);
not NOT1 (N1139, N1134);
not NOT1 (N1140, N1129);
nand NAND2 (N1141, N1138, N792);
or OR4 (N1142, N1139, N478, N784, N314);
nor NOR4 (N1143, N1142, N600, N488, N360);
xor XOR2 (N1144, N1136, N194);
xor XOR2 (N1145, N1143, N22);
buf BUF1 (N1146, N1145);
nor NOR2 (N1147, N1121, N1131);
xor XOR2 (N1148, N757, N742);
or OR2 (N1149, N1144, N1078);
or OR4 (N1150, N1137, N827, N196, N850);
not NOT1 (N1151, N1147);
and AND2 (N1152, N1146, N962);
and AND3 (N1153, N1150, N70, N750);
xor XOR2 (N1154, N1151, N220);
not NOT1 (N1155, N1153);
not NOT1 (N1156, N1149);
xor XOR2 (N1157, N1128, N466);
nor NOR3 (N1158, N1156, N900, N400);
nor NOR2 (N1159, N1155, N42);
and AND3 (N1160, N1159, N265, N322);
not NOT1 (N1161, N1148);
nand NAND3 (N1162, N1140, N460, N979);
or OR2 (N1163, N1135, N252);
nand NAND2 (N1164, N1154, N589);
xor XOR2 (N1165, N1141, N774);
or OR3 (N1166, N1158, N726, N574);
nor NOR2 (N1167, N1152, N1036);
nor NOR3 (N1168, N1160, N692, N795);
and AND4 (N1169, N1167, N61, N175, N203);
buf BUF1 (N1170, N1163);
buf BUF1 (N1171, N1133);
or OR2 (N1172, N1171, N89);
nor NOR2 (N1173, N1164, N699);
buf BUF1 (N1174, N1168);
and AND2 (N1175, N1157, N163);
or OR4 (N1176, N1174, N560, N836, N966);
not NOT1 (N1177, N1172);
xor XOR2 (N1178, N1162, N153);
nor NOR2 (N1179, N1166, N278);
or OR3 (N1180, N1165, N1134, N191);
nor NOR2 (N1181, N1175, N880);
nand NAND3 (N1182, N1161, N204, N273);
xor XOR2 (N1183, N1182, N209);
nand NAND3 (N1184, N1176, N721, N500);
or OR4 (N1185, N1173, N923, N330, N382);
and AND3 (N1186, N1184, N683, N596);
and AND2 (N1187, N1183, N388);
or OR2 (N1188, N1169, N544);
xor XOR2 (N1189, N1178, N191);
xor XOR2 (N1190, N1186, N951);
xor XOR2 (N1191, N1188, N647);
not NOT1 (N1192, N1177);
not NOT1 (N1193, N1190);
nand NAND3 (N1194, N1193, N222, N306);
and AND2 (N1195, N1194, N715);
not NOT1 (N1196, N1191);
or OR4 (N1197, N1189, N1118, N110, N980);
xor XOR2 (N1198, N1195, N862);
xor XOR2 (N1199, N1185, N666);
nand NAND4 (N1200, N1197, N721, N408, N976);
xor XOR2 (N1201, N1192, N1078);
not NOT1 (N1202, N1170);
nand NAND4 (N1203, N1198, N394, N89, N953);
not NOT1 (N1204, N1187);
not NOT1 (N1205, N1199);
and AND3 (N1206, N1202, N332, N182);
xor XOR2 (N1207, N1179, N470);
nand NAND3 (N1208, N1207, N908, N523);
xor XOR2 (N1209, N1206, N689);
or OR4 (N1210, N1180, N861, N921, N984);
xor XOR2 (N1211, N1208, N1003);
nor NOR3 (N1212, N1196, N728, N566);
xor XOR2 (N1213, N1181, N900);
buf BUF1 (N1214, N1200);
and AND2 (N1215, N1204, N1162);
and AND3 (N1216, N1212, N890, N528);
or OR4 (N1217, N1216, N141, N787, N308);
buf BUF1 (N1218, N1215);
or OR4 (N1219, N1203, N609, N618, N975);
and AND2 (N1220, N1201, N45);
buf BUF1 (N1221, N1217);
or OR3 (N1222, N1221, N757, N836);
and AND3 (N1223, N1220, N1106, N245);
nor NOR4 (N1224, N1210, N443, N145, N1141);
xor XOR2 (N1225, N1211, N951);
buf BUF1 (N1226, N1218);
not NOT1 (N1227, N1205);
nor NOR3 (N1228, N1225, N944, N1016);
or OR2 (N1229, N1209, N181);
or OR4 (N1230, N1219, N426, N1179, N706);
and AND3 (N1231, N1230, N395, N181);
and AND3 (N1232, N1228, N1218, N398);
xor XOR2 (N1233, N1232, N467);
and AND4 (N1234, N1226, N506, N228, N212);
buf BUF1 (N1235, N1222);
xor XOR2 (N1236, N1234, N1094);
nor NOR2 (N1237, N1214, N602);
nor NOR2 (N1238, N1231, N617);
xor XOR2 (N1239, N1227, N1086);
nand NAND3 (N1240, N1239, N246, N318);
or OR3 (N1241, N1237, N546, N782);
nor NOR4 (N1242, N1235, N253, N338, N1227);
nand NAND3 (N1243, N1223, N156, N588);
nor NOR2 (N1244, N1242, N751);
xor XOR2 (N1245, N1240, N324);
not NOT1 (N1246, N1243);
nor NOR2 (N1247, N1224, N218);
or OR3 (N1248, N1241, N600, N472);
nand NAND4 (N1249, N1248, N364, N647, N175);
nand NAND3 (N1250, N1238, N64, N838);
or OR2 (N1251, N1236, N595);
nand NAND4 (N1252, N1247, N760, N743, N1166);
nor NOR2 (N1253, N1252, N30);
and AND2 (N1254, N1244, N1114);
buf BUF1 (N1255, N1250);
nor NOR2 (N1256, N1249, N19);
and AND4 (N1257, N1253, N41, N220, N829);
xor XOR2 (N1258, N1213, N1239);
nor NOR3 (N1259, N1251, N692, N325);
nand NAND4 (N1260, N1256, N764, N371, N1065);
nor NOR2 (N1261, N1255, N596);
xor XOR2 (N1262, N1259, N1038);
xor XOR2 (N1263, N1257, N1173);
or OR2 (N1264, N1262, N990);
buf BUF1 (N1265, N1263);
or OR3 (N1266, N1254, N736, N470);
nor NOR4 (N1267, N1245, N670, N762, N819);
xor XOR2 (N1268, N1246, N1231);
or OR3 (N1269, N1264, N1168, N1165);
or OR3 (N1270, N1260, N329, N90);
xor XOR2 (N1271, N1258, N354);
nand NAND2 (N1272, N1229, N302);
nand NAND4 (N1273, N1233, N453, N728, N735);
nand NAND4 (N1274, N1273, N649, N348, N1270);
xor XOR2 (N1275, N1166, N271);
nor NOR3 (N1276, N1268, N920, N613);
or OR4 (N1277, N1261, N893, N941, N1259);
not NOT1 (N1278, N1265);
buf BUF1 (N1279, N1271);
or OR4 (N1280, N1277, N1221, N1011, N535);
xor XOR2 (N1281, N1269, N881);
or OR2 (N1282, N1272, N475);
not NOT1 (N1283, N1275);
nand NAND4 (N1284, N1282, N212, N1149, N1186);
or OR2 (N1285, N1279, N734);
nand NAND4 (N1286, N1266, N1065, N1209, N780);
and AND3 (N1287, N1280, N1201, N700);
nand NAND3 (N1288, N1278, N533, N1045);
nor NOR3 (N1289, N1284, N273, N573);
nand NAND2 (N1290, N1289, N792);
and AND4 (N1291, N1276, N1283, N559, N1259);
or OR3 (N1292, N650, N202, N167);
not NOT1 (N1293, N1274);
and AND2 (N1294, N1285, N583);
nor NOR2 (N1295, N1267, N986);
and AND2 (N1296, N1294, N469);
buf BUF1 (N1297, N1287);
nand NAND3 (N1298, N1286, N221, N264);
or OR4 (N1299, N1288, N1015, N1205, N1263);
nand NAND4 (N1300, N1292, N1292, N1291, N499);
or OR4 (N1301, N509, N1299, N1079, N484);
buf BUF1 (N1302, N1154);
xor XOR2 (N1303, N1290, N559);
not NOT1 (N1304, N1303);
nor NOR4 (N1305, N1295, N1288, N496, N18);
not NOT1 (N1306, N1297);
xor XOR2 (N1307, N1301, N948);
not NOT1 (N1308, N1302);
buf BUF1 (N1309, N1305);
xor XOR2 (N1310, N1306, N791);
not NOT1 (N1311, N1304);
not NOT1 (N1312, N1281);
nor NOR4 (N1313, N1310, N276, N37, N16);
buf BUF1 (N1314, N1300);
and AND2 (N1315, N1313, N434);
buf BUF1 (N1316, N1298);
nand NAND3 (N1317, N1296, N63, N1156);
nand NAND4 (N1318, N1317, N1076, N677, N321);
xor XOR2 (N1319, N1309, N1154);
or OR4 (N1320, N1318, N191, N702, N436);
nand NAND4 (N1321, N1308, N1155, N1246, N109);
or OR2 (N1322, N1315, N323);
nand NAND2 (N1323, N1316, N938);
nand NAND4 (N1324, N1312, N23, N930, N597);
nand NAND2 (N1325, N1319, N1112);
nand NAND3 (N1326, N1324, N160, N751);
xor XOR2 (N1327, N1314, N348);
buf BUF1 (N1328, N1321);
nand NAND3 (N1329, N1326, N297, N372);
and AND2 (N1330, N1328, N1087);
buf BUF1 (N1331, N1320);
and AND2 (N1332, N1325, N1194);
xor XOR2 (N1333, N1329, N667);
buf BUF1 (N1334, N1333);
or OR2 (N1335, N1322, N28);
and AND3 (N1336, N1330, N936, N95);
xor XOR2 (N1337, N1332, N857);
buf BUF1 (N1338, N1331);
nor NOR3 (N1339, N1338, N1033, N598);
nand NAND2 (N1340, N1334, N416);
xor XOR2 (N1341, N1323, N71);
not NOT1 (N1342, N1335);
or OR4 (N1343, N1340, N987, N1304, N895);
or OR3 (N1344, N1293, N690, N1237);
xor XOR2 (N1345, N1307, N403);
nand NAND3 (N1346, N1339, N1324, N941);
not NOT1 (N1347, N1344);
not NOT1 (N1348, N1342);
nor NOR4 (N1349, N1337, N452, N800, N620);
and AND4 (N1350, N1311, N755, N15, N160);
and AND2 (N1351, N1345, N285);
or OR2 (N1352, N1350, N866);
not NOT1 (N1353, N1327);
or OR4 (N1354, N1352, N1085, N430, N4);
buf BUF1 (N1355, N1343);
not NOT1 (N1356, N1341);
not NOT1 (N1357, N1336);
nand NAND4 (N1358, N1355, N978, N1112, N986);
or OR3 (N1359, N1348, N1066, N765);
or OR3 (N1360, N1353, N695, N213);
buf BUF1 (N1361, N1357);
not NOT1 (N1362, N1359);
not NOT1 (N1363, N1362);
buf BUF1 (N1364, N1349);
buf BUF1 (N1365, N1364);
not NOT1 (N1366, N1356);
or OR2 (N1367, N1360, N816);
nand NAND2 (N1368, N1354, N19);
or OR3 (N1369, N1358, N834, N1294);
or OR2 (N1370, N1366, N888);
or OR4 (N1371, N1369, N135, N1215, N329);
nand NAND2 (N1372, N1361, N898);
buf BUF1 (N1373, N1351);
not NOT1 (N1374, N1347);
nand NAND2 (N1375, N1374, N1297);
buf BUF1 (N1376, N1367);
not NOT1 (N1377, N1372);
nand NAND4 (N1378, N1375, N494, N592, N824);
nand NAND2 (N1379, N1370, N1170);
xor XOR2 (N1380, N1373, N565);
xor XOR2 (N1381, N1365, N1215);
nor NOR4 (N1382, N1371, N1154, N1083, N1255);
not NOT1 (N1383, N1363);
not NOT1 (N1384, N1376);
xor XOR2 (N1385, N1384, N765);
nor NOR4 (N1386, N1368, N355, N569, N439);
buf BUF1 (N1387, N1378);
or OR4 (N1388, N1346, N954, N1112, N657);
nand NAND2 (N1389, N1385, N19);
xor XOR2 (N1390, N1386, N643);
buf BUF1 (N1391, N1380);
buf BUF1 (N1392, N1390);
and AND3 (N1393, N1382, N371, N577);
xor XOR2 (N1394, N1389, N1381);
buf BUF1 (N1395, N173);
xor XOR2 (N1396, N1392, N408);
nor NOR4 (N1397, N1388, N176, N535, N1019);
nand NAND2 (N1398, N1397, N416);
nor NOR2 (N1399, N1377, N441);
or OR3 (N1400, N1399, N229, N854);
nand NAND2 (N1401, N1395, N827);
or OR3 (N1402, N1400, N563, N615);
not NOT1 (N1403, N1396);
nand NAND3 (N1404, N1387, N305, N1147);
or OR2 (N1405, N1401, N738);
nand NAND4 (N1406, N1394, N51, N1040, N918);
nor NOR3 (N1407, N1379, N41, N1163);
xor XOR2 (N1408, N1405, N1053);
buf BUF1 (N1409, N1404);
nand NAND3 (N1410, N1393, N1372, N651);
or OR4 (N1411, N1406, N996, N809, N533);
not NOT1 (N1412, N1407);
xor XOR2 (N1413, N1383, N150);
buf BUF1 (N1414, N1398);
or OR2 (N1415, N1409, N1167);
buf BUF1 (N1416, N1410);
and AND4 (N1417, N1391, N1107, N217, N941);
and AND3 (N1418, N1402, N890, N1232);
nand NAND3 (N1419, N1403, N997, N687);
nor NOR3 (N1420, N1408, N9, N953);
or OR2 (N1421, N1418, N497);
and AND4 (N1422, N1412, N1289, N667, N629);
nor NOR3 (N1423, N1419, N545, N1004);
buf BUF1 (N1424, N1413);
and AND4 (N1425, N1422, N180, N24, N1167);
nor NOR4 (N1426, N1414, N241, N1415, N1083);
or OR4 (N1427, N143, N382, N821, N126);
and AND4 (N1428, N1411, N692, N1313, N42);
not NOT1 (N1429, N1425);
nand NAND3 (N1430, N1423, N1297, N1178);
nor NOR2 (N1431, N1429, N1327);
not NOT1 (N1432, N1431);
not NOT1 (N1433, N1421);
or OR3 (N1434, N1417, N597, N1207);
or OR2 (N1435, N1430, N636);
not NOT1 (N1436, N1432);
nor NOR3 (N1437, N1420, N600, N273);
not NOT1 (N1438, N1434);
and AND2 (N1439, N1437, N748);
buf BUF1 (N1440, N1439);
and AND3 (N1441, N1426, N792, N202);
xor XOR2 (N1442, N1428, N1272);
and AND4 (N1443, N1436, N1409, N135, N1439);
nand NAND3 (N1444, N1440, N667, N1153);
not NOT1 (N1445, N1438);
or OR2 (N1446, N1424, N1381);
and AND4 (N1447, N1433, N89, N748, N851);
not NOT1 (N1448, N1416);
not NOT1 (N1449, N1435);
not NOT1 (N1450, N1427);
nor NOR2 (N1451, N1450, N1209);
xor XOR2 (N1452, N1443, N197);
buf BUF1 (N1453, N1448);
buf BUF1 (N1454, N1453);
and AND3 (N1455, N1446, N527, N1264);
xor XOR2 (N1456, N1451, N1130);
xor XOR2 (N1457, N1444, N49);
not NOT1 (N1458, N1449);
not NOT1 (N1459, N1442);
nor NOR4 (N1460, N1445, N1188, N121, N551);
buf BUF1 (N1461, N1456);
nor NOR2 (N1462, N1459, N272);
not NOT1 (N1463, N1461);
buf BUF1 (N1464, N1457);
or OR2 (N1465, N1463, N938);
buf BUF1 (N1466, N1464);
buf BUF1 (N1467, N1455);
xor XOR2 (N1468, N1452, N1098);
nor NOR3 (N1469, N1460, N662, N754);
nand NAND3 (N1470, N1468, N735, N669);
buf BUF1 (N1471, N1465);
not NOT1 (N1472, N1467);
not NOT1 (N1473, N1471);
or OR2 (N1474, N1441, N910);
or OR3 (N1475, N1473, N176, N1324);
nand NAND3 (N1476, N1466, N112, N1424);
and AND2 (N1477, N1469, N1155);
nand NAND4 (N1478, N1472, N1204, N108, N44);
nor NOR3 (N1479, N1454, N1350, N1308);
buf BUF1 (N1480, N1476);
or OR3 (N1481, N1474, N231, N425);
nor NOR4 (N1482, N1477, N1304, N145, N1401);
and AND3 (N1483, N1481, N1144, N212);
xor XOR2 (N1484, N1478, N308);
or OR3 (N1485, N1462, N318, N67);
buf BUF1 (N1486, N1484);
and AND4 (N1487, N1486, N139, N311, N1213);
xor XOR2 (N1488, N1483, N1297);
or OR4 (N1489, N1488, N909, N1168, N1427);
nand NAND2 (N1490, N1487, N85);
buf BUF1 (N1491, N1490);
nand NAND3 (N1492, N1489, N645, N118);
xor XOR2 (N1493, N1491, N101);
nand NAND3 (N1494, N1480, N873, N293);
nor NOR4 (N1495, N1485, N278, N9, N559);
and AND4 (N1496, N1479, N521, N778, N3);
nand NAND4 (N1497, N1470, N383, N856, N508);
not NOT1 (N1498, N1495);
nand NAND3 (N1499, N1475, N1430, N319);
xor XOR2 (N1500, N1493, N443);
or OR4 (N1501, N1458, N454, N1377, N1250);
buf BUF1 (N1502, N1499);
not NOT1 (N1503, N1500);
not NOT1 (N1504, N1494);
not NOT1 (N1505, N1492);
or OR4 (N1506, N1501, N1295, N1226, N105);
nor NOR2 (N1507, N1498, N945);
and AND3 (N1508, N1482, N1389, N1148);
xor XOR2 (N1509, N1497, N591);
not NOT1 (N1510, N1509);
nand NAND2 (N1511, N1503, N14);
buf BUF1 (N1512, N1507);
xor XOR2 (N1513, N1511, N66);
nand NAND4 (N1514, N1506, N1200, N534, N854);
nor NOR2 (N1515, N1510, N944);
nor NOR3 (N1516, N1496, N230, N1503);
and AND3 (N1517, N1514, N338, N1454);
nor NOR3 (N1518, N1508, N1162, N1136);
nor NOR4 (N1519, N1516, N1358, N1204, N64);
xor XOR2 (N1520, N1504, N825);
and AND2 (N1521, N1502, N528);
nor NOR2 (N1522, N1515, N727);
nand NAND2 (N1523, N1505, N1350);
or OR3 (N1524, N1447, N90, N1460);
not NOT1 (N1525, N1519);
buf BUF1 (N1526, N1512);
nor NOR3 (N1527, N1520, N1385, N986);
nand NAND3 (N1528, N1522, N16, N1153);
nor NOR3 (N1529, N1528, N1131, N22);
nand NAND3 (N1530, N1518, N1524, N370);
and AND4 (N1531, N142, N528, N1244, N96);
xor XOR2 (N1532, N1517, N1241);
nand NAND2 (N1533, N1526, N257);
nand NAND4 (N1534, N1525, N1338, N906, N1298);
nand NAND3 (N1535, N1530, N264, N1274);
xor XOR2 (N1536, N1534, N299);
nand NAND2 (N1537, N1531, N1190);
xor XOR2 (N1538, N1532, N1446);
buf BUF1 (N1539, N1536);
buf BUF1 (N1540, N1513);
nor NOR4 (N1541, N1539, N1203, N1284, N575);
or OR2 (N1542, N1537, N331);
not NOT1 (N1543, N1542);
buf BUF1 (N1544, N1543);
nand NAND3 (N1545, N1544, N594, N1120);
xor XOR2 (N1546, N1538, N359);
nand NAND3 (N1547, N1546, N517, N51);
nor NOR4 (N1548, N1521, N250, N1215, N229);
nand NAND3 (N1549, N1533, N89, N1389);
not NOT1 (N1550, N1527);
and AND3 (N1551, N1547, N1062, N1422);
and AND2 (N1552, N1540, N631);
and AND3 (N1553, N1535, N179, N480);
nand NAND2 (N1554, N1523, N80);
nand NAND3 (N1555, N1541, N283, N31);
not NOT1 (N1556, N1545);
nand NAND3 (N1557, N1549, N757, N304);
xor XOR2 (N1558, N1551, N1333);
and AND2 (N1559, N1529, N1201);
or OR4 (N1560, N1552, N1098, N351, N578);
buf BUF1 (N1561, N1560);
nor NOR2 (N1562, N1553, N775);
buf BUF1 (N1563, N1556);
buf BUF1 (N1564, N1548);
or OR2 (N1565, N1563, N1434);
not NOT1 (N1566, N1565);
nor NOR2 (N1567, N1550, N161);
xor XOR2 (N1568, N1555, N616);
buf BUF1 (N1569, N1558);
or OR2 (N1570, N1568, N735);
and AND2 (N1571, N1554, N1405);
not NOT1 (N1572, N1557);
nor NOR2 (N1573, N1559, N1508);
nand NAND3 (N1574, N1561, N1192, N1300);
nor NOR4 (N1575, N1571, N892, N684, N1014);
and AND4 (N1576, N1570, N203, N485, N238);
or OR3 (N1577, N1575, N544, N1541);
buf BUF1 (N1578, N1567);
and AND4 (N1579, N1564, N916, N543, N1188);
nand NAND2 (N1580, N1562, N307);
not NOT1 (N1581, N1574);
buf BUF1 (N1582, N1581);
not NOT1 (N1583, N1576);
and AND3 (N1584, N1580, N247, N1271);
xor XOR2 (N1585, N1566, N658);
buf BUF1 (N1586, N1578);
not NOT1 (N1587, N1573);
and AND4 (N1588, N1569, N1043, N867, N1140);
not NOT1 (N1589, N1582);
or OR3 (N1590, N1585, N1073, N330);
xor XOR2 (N1591, N1584, N52);
xor XOR2 (N1592, N1587, N1456);
xor XOR2 (N1593, N1591, N444);
and AND4 (N1594, N1583, N240, N738, N1076);
buf BUF1 (N1595, N1590);
and AND3 (N1596, N1577, N675, N955);
or OR3 (N1597, N1593, N1455, N677);
nand NAND4 (N1598, N1596, N1459, N1531, N744);
buf BUF1 (N1599, N1579);
or OR3 (N1600, N1592, N1301, N1007);
buf BUF1 (N1601, N1600);
nor NOR4 (N1602, N1597, N17, N34, N1178);
or OR3 (N1603, N1588, N581, N469);
nor NOR3 (N1604, N1601, N1432, N984);
and AND2 (N1605, N1589, N625);
nand NAND3 (N1606, N1594, N525, N369);
and AND4 (N1607, N1604, N1427, N630, N481);
nor NOR4 (N1608, N1602, N519, N1014, N982);
buf BUF1 (N1609, N1606);
nand NAND4 (N1610, N1605, N153, N14, N882);
nor NOR3 (N1611, N1599, N479, N368);
buf BUF1 (N1612, N1608);
or OR4 (N1613, N1586, N1082, N1060, N14);
or OR2 (N1614, N1612, N1397);
xor XOR2 (N1615, N1609, N1387);
buf BUF1 (N1616, N1603);
xor XOR2 (N1617, N1572, N1399);
buf BUF1 (N1618, N1614);
nor NOR2 (N1619, N1616, N1043);
nor NOR2 (N1620, N1610, N526);
nor NOR3 (N1621, N1615, N110, N409);
nor NOR2 (N1622, N1620, N1213);
buf BUF1 (N1623, N1607);
not NOT1 (N1624, N1598);
nand NAND4 (N1625, N1613, N574, N700, N523);
nand NAND3 (N1626, N1622, N198, N1455);
not NOT1 (N1627, N1618);
xor XOR2 (N1628, N1623, N1591);
nor NOR4 (N1629, N1621, N852, N492, N1426);
xor XOR2 (N1630, N1619, N885);
not NOT1 (N1631, N1595);
nand NAND4 (N1632, N1625, N527, N1572, N134);
not NOT1 (N1633, N1629);
and AND4 (N1634, N1617, N423, N1144, N1142);
or OR4 (N1635, N1631, N1279, N1260, N1005);
nor NOR4 (N1636, N1633, N594, N709, N312);
not NOT1 (N1637, N1636);
and AND3 (N1638, N1624, N700, N1038);
nor NOR3 (N1639, N1634, N736, N998);
or OR2 (N1640, N1632, N801);
not NOT1 (N1641, N1628);
nor NOR4 (N1642, N1611, N739, N644, N609);
and AND2 (N1643, N1635, N227);
and AND3 (N1644, N1640, N1292, N293);
and AND2 (N1645, N1637, N244);
nor NOR2 (N1646, N1630, N272);
and AND3 (N1647, N1643, N744, N1469);
nand NAND4 (N1648, N1638, N137, N870, N990);
not NOT1 (N1649, N1639);
nand NAND2 (N1650, N1649, N281);
buf BUF1 (N1651, N1645);
and AND4 (N1652, N1626, N1091, N903, N1312);
nand NAND3 (N1653, N1642, N1507, N1526);
nor NOR3 (N1654, N1653, N137, N376);
and AND3 (N1655, N1641, N1161, N107);
buf BUF1 (N1656, N1627);
nand NAND4 (N1657, N1654, N767, N1391, N1387);
not NOT1 (N1658, N1650);
not NOT1 (N1659, N1647);
buf BUF1 (N1660, N1655);
or OR4 (N1661, N1658, N497, N550, N96);
buf BUF1 (N1662, N1652);
nor NOR4 (N1663, N1661, N384, N752, N797);
nor NOR3 (N1664, N1660, N317, N1466);
or OR4 (N1665, N1657, N85, N1077, N775);
buf BUF1 (N1666, N1665);
and AND2 (N1667, N1666, N1514);
not NOT1 (N1668, N1648);
or OR4 (N1669, N1667, N449, N237, N338);
or OR3 (N1670, N1664, N638, N546);
and AND3 (N1671, N1651, N741, N918);
xor XOR2 (N1672, N1663, N1008);
xor XOR2 (N1673, N1659, N1350);
and AND3 (N1674, N1668, N1180, N1216);
nand NAND3 (N1675, N1662, N1205, N406);
nor NOR3 (N1676, N1656, N517, N897);
nor NOR2 (N1677, N1676, N40);
and AND4 (N1678, N1672, N311, N1336, N239);
nor NOR4 (N1679, N1646, N919, N452, N503);
or OR2 (N1680, N1674, N1386);
and AND4 (N1681, N1677, N577, N1680, N1672);
xor XOR2 (N1682, N394, N1638);
nor NOR3 (N1683, N1644, N1256, N799);
or OR2 (N1684, N1669, N428);
or OR4 (N1685, N1681, N1656, N365, N654);
buf BUF1 (N1686, N1678);
not NOT1 (N1687, N1682);
xor XOR2 (N1688, N1673, N755);
or OR2 (N1689, N1688, N103);
and AND3 (N1690, N1675, N652, N767);
nor NOR3 (N1691, N1683, N885, N1368);
nor NOR4 (N1692, N1687, N1224, N639, N682);
xor XOR2 (N1693, N1671, N544);
not NOT1 (N1694, N1679);
buf BUF1 (N1695, N1692);
and AND3 (N1696, N1686, N429, N295);
and AND2 (N1697, N1693, N883);
nor NOR2 (N1698, N1690, N508);
nor NOR2 (N1699, N1691, N723);
xor XOR2 (N1700, N1695, N490);
xor XOR2 (N1701, N1685, N1449);
not NOT1 (N1702, N1696);
nor NOR3 (N1703, N1694, N1506, N835);
nor NOR4 (N1704, N1698, N1002, N1272, N670);
and AND3 (N1705, N1702, N1469, N746);
buf BUF1 (N1706, N1689);
or OR3 (N1707, N1700, N1602, N1535);
nand NAND3 (N1708, N1699, N228, N589);
not NOT1 (N1709, N1707);
nand NAND2 (N1710, N1684, N945);
xor XOR2 (N1711, N1709, N320);
and AND3 (N1712, N1706, N477, N359);
xor XOR2 (N1713, N1701, N997);
nor NOR2 (N1714, N1708, N1178);
xor XOR2 (N1715, N1711, N1112);
nand NAND3 (N1716, N1715, N1069, N734);
or OR3 (N1717, N1714, N220, N1658);
not NOT1 (N1718, N1712);
and AND4 (N1719, N1710, N958, N365, N1197);
not NOT1 (N1720, N1719);
not NOT1 (N1721, N1704);
nand NAND3 (N1722, N1718, N535, N1308);
and AND3 (N1723, N1705, N26, N635);
nand NAND2 (N1724, N1723, N596);
or OR4 (N1725, N1716, N1342, N915, N110);
xor XOR2 (N1726, N1717, N673);
buf BUF1 (N1727, N1713);
nor NOR4 (N1728, N1724, N1312, N1084, N1718);
nor NOR4 (N1729, N1697, N724, N185, N1276);
or OR4 (N1730, N1670, N245, N1363, N1000);
nand NAND3 (N1731, N1730, N228, N766);
buf BUF1 (N1732, N1721);
nor NOR2 (N1733, N1703, N1695);
nand NAND2 (N1734, N1728, N313);
buf BUF1 (N1735, N1726);
xor XOR2 (N1736, N1727, N1162);
not NOT1 (N1737, N1729);
not NOT1 (N1738, N1734);
xor XOR2 (N1739, N1738, N755);
buf BUF1 (N1740, N1739);
and AND3 (N1741, N1737, N419, N1592);
not NOT1 (N1742, N1722);
buf BUF1 (N1743, N1725);
nand NAND3 (N1744, N1740, N839, N204);
nor NOR2 (N1745, N1731, N331);
nand NAND4 (N1746, N1732, N1468, N1181, N472);
not NOT1 (N1747, N1733);
not NOT1 (N1748, N1720);
nor NOR2 (N1749, N1746, N1296);
or OR4 (N1750, N1745, N1017, N905, N733);
nand NAND4 (N1751, N1742, N1255, N1051, N1598);
nor NOR4 (N1752, N1749, N1142, N1750, N845);
not NOT1 (N1753, N1715);
not NOT1 (N1754, N1744);
nor NOR2 (N1755, N1741, N639);
not NOT1 (N1756, N1743);
or OR4 (N1757, N1736, N457, N984, N1164);
xor XOR2 (N1758, N1751, N139);
buf BUF1 (N1759, N1757);
nand NAND4 (N1760, N1747, N1527, N769, N199);
nor NOR2 (N1761, N1754, N1746);
nor NOR3 (N1762, N1760, N1022, N1209);
or OR2 (N1763, N1759, N1637);
and AND2 (N1764, N1753, N938);
and AND4 (N1765, N1761, N1487, N1247, N1160);
and AND3 (N1766, N1735, N1461, N132);
not NOT1 (N1767, N1764);
xor XOR2 (N1768, N1765, N977);
buf BUF1 (N1769, N1762);
nor NOR3 (N1770, N1756, N521, N1401);
and AND3 (N1771, N1763, N1369, N1436);
not NOT1 (N1772, N1752);
buf BUF1 (N1773, N1766);
nor NOR3 (N1774, N1758, N448, N1707);
or OR3 (N1775, N1767, N1477, N1013);
or OR2 (N1776, N1774, N1402);
xor XOR2 (N1777, N1768, N897);
nor NOR3 (N1778, N1775, N300, N1298);
and AND4 (N1779, N1769, N191, N350, N1452);
buf BUF1 (N1780, N1748);
not NOT1 (N1781, N1755);
xor XOR2 (N1782, N1771, N428);
not NOT1 (N1783, N1777);
or OR2 (N1784, N1780, N108);
xor XOR2 (N1785, N1782, N264);
nor NOR4 (N1786, N1783, N534, N1629, N1408);
and AND2 (N1787, N1770, N1644);
or OR2 (N1788, N1772, N198);
xor XOR2 (N1789, N1784, N1007);
buf BUF1 (N1790, N1779);
buf BUF1 (N1791, N1776);
nor NOR3 (N1792, N1790, N375, N1184);
and AND2 (N1793, N1792, N354);
buf BUF1 (N1794, N1791);
and AND4 (N1795, N1787, N941, N1497, N1634);
xor XOR2 (N1796, N1778, N1194);
nand NAND3 (N1797, N1796, N1356, N893);
not NOT1 (N1798, N1781);
nor NOR4 (N1799, N1773, N1400, N449, N785);
not NOT1 (N1800, N1786);
xor XOR2 (N1801, N1797, N1481);
or OR3 (N1802, N1801, N711, N1200);
and AND2 (N1803, N1799, N1528);
or OR2 (N1804, N1793, N1454);
not NOT1 (N1805, N1802);
and AND2 (N1806, N1789, N1146);
xor XOR2 (N1807, N1806, N1345);
xor XOR2 (N1808, N1804, N40);
not NOT1 (N1809, N1800);
or OR3 (N1810, N1795, N41, N531);
or OR3 (N1811, N1805, N1493, N1343);
or OR4 (N1812, N1794, N1359, N1524, N757);
nand NAND3 (N1813, N1811, N362, N262);
xor XOR2 (N1814, N1798, N247);
and AND3 (N1815, N1814, N610, N1045);
and AND4 (N1816, N1813, N112, N1412, N533);
buf BUF1 (N1817, N1785);
xor XOR2 (N1818, N1816, N1698);
nor NOR4 (N1819, N1817, N1197, N636, N540);
and AND2 (N1820, N1818, N922);
buf BUF1 (N1821, N1819);
nor NOR3 (N1822, N1821, N105, N712);
and AND2 (N1823, N1812, N794);
and AND4 (N1824, N1803, N223, N396, N281);
and AND2 (N1825, N1824, N1765);
nor NOR2 (N1826, N1807, N1291);
and AND3 (N1827, N1788, N399, N360);
or OR3 (N1828, N1826, N804, N1294);
nand NAND2 (N1829, N1809, N909);
xor XOR2 (N1830, N1810, N1478);
nor NOR3 (N1831, N1830, N1465, N853);
not NOT1 (N1832, N1831);
or OR4 (N1833, N1828, N268, N1803, N291);
not NOT1 (N1834, N1820);
or OR3 (N1835, N1829, N1315, N1101);
xor XOR2 (N1836, N1822, N1406);
not NOT1 (N1837, N1833);
nand NAND4 (N1838, N1825, N410, N619, N1257);
nor NOR2 (N1839, N1838, N1270);
and AND4 (N1840, N1832, N1423, N1351, N17);
xor XOR2 (N1841, N1823, N1422);
not NOT1 (N1842, N1839);
nor NOR4 (N1843, N1840, N684, N1796, N1109);
xor XOR2 (N1844, N1843, N1251);
or OR3 (N1845, N1834, N17, N1404);
and AND2 (N1846, N1844, N785);
nor NOR2 (N1847, N1835, N1045);
nor NOR3 (N1848, N1827, N1074, N513);
not NOT1 (N1849, N1815);
buf BUF1 (N1850, N1846);
buf BUF1 (N1851, N1849);
and AND2 (N1852, N1808, N973);
and AND3 (N1853, N1851, N372, N1055);
nor NOR4 (N1854, N1842, N8, N711, N1731);
or OR4 (N1855, N1853, N1555, N1762, N444);
and AND4 (N1856, N1854, N798, N254, N951);
nor NOR4 (N1857, N1847, N691, N1234, N1752);
not NOT1 (N1858, N1857);
and AND2 (N1859, N1841, N1700);
and AND3 (N1860, N1856, N233, N1017);
and AND3 (N1861, N1860, N676, N1154);
buf BUF1 (N1862, N1858);
not NOT1 (N1863, N1837);
buf BUF1 (N1864, N1850);
and AND4 (N1865, N1864, N1688, N278, N1050);
nor NOR3 (N1866, N1865, N254, N316);
nor NOR2 (N1867, N1836, N1165);
not NOT1 (N1868, N1845);
and AND4 (N1869, N1855, N1328, N1251, N611);
buf BUF1 (N1870, N1863);
xor XOR2 (N1871, N1862, N286);
nand NAND2 (N1872, N1870, N1753);
and AND4 (N1873, N1872, N1211, N1499, N515);
and AND4 (N1874, N1852, N645, N253, N609);
and AND4 (N1875, N1859, N890, N1315, N39);
nand NAND2 (N1876, N1848, N1570);
xor XOR2 (N1877, N1876, N492);
buf BUF1 (N1878, N1871);
xor XOR2 (N1879, N1866, N1655);
or OR3 (N1880, N1861, N128, N1039);
nor NOR2 (N1881, N1877, N914);
not NOT1 (N1882, N1879);
xor XOR2 (N1883, N1880, N1697);
buf BUF1 (N1884, N1868);
not NOT1 (N1885, N1869);
and AND4 (N1886, N1884, N772, N1706, N567);
nand NAND4 (N1887, N1875, N1453, N367, N497);
and AND4 (N1888, N1881, N1887, N1525, N153);
nor NOR3 (N1889, N1004, N619, N927);
or OR3 (N1890, N1888, N734, N1838);
and AND2 (N1891, N1890, N441);
nor NOR3 (N1892, N1886, N1415, N1786);
nor NOR3 (N1893, N1883, N1064, N180);
not NOT1 (N1894, N1892);
not NOT1 (N1895, N1882);
nor NOR2 (N1896, N1867, N870);
xor XOR2 (N1897, N1896, N1532);
buf BUF1 (N1898, N1889);
not NOT1 (N1899, N1873);
buf BUF1 (N1900, N1878);
or OR4 (N1901, N1895, N162, N1683, N1876);
or OR4 (N1902, N1885, N1373, N663, N5);
nor NOR3 (N1903, N1891, N1343, N1133);
nor NOR3 (N1904, N1898, N82, N1784);
nand NAND3 (N1905, N1894, N1460, N641);
and AND2 (N1906, N1904, N181);
buf BUF1 (N1907, N1874);
xor XOR2 (N1908, N1900, N16);
xor XOR2 (N1909, N1897, N931);
buf BUF1 (N1910, N1902);
nand NAND2 (N1911, N1899, N416);
nand NAND2 (N1912, N1903, N484);
or OR3 (N1913, N1901, N1903, N805);
or OR2 (N1914, N1906, N484);
nor NOR2 (N1915, N1910, N1868);
nand NAND2 (N1916, N1915, N1826);
or OR3 (N1917, N1912, N1089, N363);
xor XOR2 (N1918, N1916, N256);
xor XOR2 (N1919, N1913, N1068);
buf BUF1 (N1920, N1908);
buf BUF1 (N1921, N1920);
nor NOR3 (N1922, N1919, N1849, N648);
nor NOR3 (N1923, N1918, N1523, N658);
nand NAND2 (N1924, N1914, N1103);
and AND2 (N1925, N1924, N1282);
not NOT1 (N1926, N1923);
or OR2 (N1927, N1905, N1531);
nand NAND3 (N1928, N1925, N1200, N1489);
nor NOR4 (N1929, N1909, N709, N1096, N969);
buf BUF1 (N1930, N1929);
or OR4 (N1931, N1893, N780, N1469, N72);
nor NOR4 (N1932, N1926, N729, N760, N650);
buf BUF1 (N1933, N1922);
or OR2 (N1934, N1932, N1358);
and AND4 (N1935, N1933, N208, N1919, N1177);
nor NOR4 (N1936, N1911, N155, N339, N1696);
and AND4 (N1937, N1930, N1553, N1365, N917);
buf BUF1 (N1938, N1935);
and AND4 (N1939, N1917, N944, N134, N572);
nand NAND4 (N1940, N1936, N1898, N117, N406);
and AND4 (N1941, N1927, N1890, N923, N289);
xor XOR2 (N1942, N1907, N1472);
nor NOR4 (N1943, N1940, N129, N1080, N1383);
nor NOR3 (N1944, N1928, N1158, N1873);
nor NOR4 (N1945, N1938, N916, N1881, N723);
nor NOR3 (N1946, N1937, N824, N442);
buf BUF1 (N1947, N1944);
or OR2 (N1948, N1947, N1033);
buf BUF1 (N1949, N1948);
and AND3 (N1950, N1931, N349, N526);
buf BUF1 (N1951, N1934);
or OR3 (N1952, N1949, N1127, N768);
or OR3 (N1953, N1946, N810, N1209);
nor NOR4 (N1954, N1953, N909, N684, N1057);
buf BUF1 (N1955, N1921);
xor XOR2 (N1956, N1952, N910);
not NOT1 (N1957, N1941);
nor NOR4 (N1958, N1939, N1034, N334, N531);
or OR4 (N1959, N1954, N665, N668, N1713);
nand NAND3 (N1960, N1943, N1740, N1456);
or OR3 (N1961, N1955, N1324, N854);
nor NOR3 (N1962, N1950, N1103, N142);
nand NAND4 (N1963, N1962, N1948, N1817, N521);
xor XOR2 (N1964, N1942, N1725);
or OR2 (N1965, N1945, N1625);
not NOT1 (N1966, N1963);
or OR3 (N1967, N1960, N327, N1451);
buf BUF1 (N1968, N1965);
nand NAND4 (N1969, N1961, N1529, N1295, N789);
or OR4 (N1970, N1969, N1030, N1565, N1592);
nor NOR4 (N1971, N1970, N1121, N1754, N917);
and AND2 (N1972, N1951, N306);
and AND3 (N1973, N1958, N1616, N1134);
or OR2 (N1974, N1973, N704);
nand NAND4 (N1975, N1964, N881, N805, N783);
or OR3 (N1976, N1967, N1815, N934);
or OR4 (N1977, N1956, N1726, N102, N261);
xor XOR2 (N1978, N1975, N1314);
or OR4 (N1979, N1968, N1870, N1784, N1764);
xor XOR2 (N1980, N1966, N630);
xor XOR2 (N1981, N1971, N247);
xor XOR2 (N1982, N1977, N149);
or OR4 (N1983, N1959, N407, N1211, N984);
nor NOR2 (N1984, N1972, N878);
or OR4 (N1985, N1984, N854, N7, N988);
nand NAND4 (N1986, N1982, N958, N34, N917);
or OR4 (N1987, N1974, N1014, N1357, N454);
nand NAND3 (N1988, N1978, N1569, N952);
and AND3 (N1989, N1981, N1603, N1042);
nor NOR2 (N1990, N1987, N991);
or OR3 (N1991, N1990, N1797, N669);
nand NAND3 (N1992, N1988, N1030, N931);
and AND4 (N1993, N1992, N415, N199, N880);
nand NAND4 (N1994, N1980, N490, N658, N1981);
not NOT1 (N1995, N1993);
nand NAND2 (N1996, N1983, N576);
and AND4 (N1997, N1957, N1861, N1454, N854);
nor NOR2 (N1998, N1979, N674);
and AND3 (N1999, N1997, N1597, N1204);
not NOT1 (N2000, N1999);
nor NOR4 (N2001, N1991, N1186, N1786, N223);
nand NAND3 (N2002, N1994, N997, N94);
and AND2 (N2003, N2000, N1479);
and AND4 (N2004, N1986, N319, N535, N1195);
and AND3 (N2005, N2003, N1333, N1069);
buf BUF1 (N2006, N1985);
or OR3 (N2007, N1989, N1464, N87);
xor XOR2 (N2008, N2004, N1541);
nor NOR4 (N2009, N2001, N305, N1265, N1785);
or OR3 (N2010, N1995, N617, N1732);
xor XOR2 (N2011, N1998, N484);
and AND2 (N2012, N2006, N1839);
and AND2 (N2013, N2005, N667);
buf BUF1 (N2014, N2012);
nor NOR4 (N2015, N2007, N647, N54, N1352);
buf BUF1 (N2016, N2013);
or OR4 (N2017, N1976, N1934, N818, N1221);
buf BUF1 (N2018, N2010);
or OR4 (N2019, N2002, N1795, N1224, N1276);
not NOT1 (N2020, N2014);
not NOT1 (N2021, N2020);
buf BUF1 (N2022, N2015);
or OR2 (N2023, N2021, N1670);
buf BUF1 (N2024, N2009);
and AND2 (N2025, N2019, N482);
nand NAND2 (N2026, N2018, N865);
not NOT1 (N2027, N2025);
buf BUF1 (N2028, N2016);
not NOT1 (N2029, N2011);
buf BUF1 (N2030, N1996);
buf BUF1 (N2031, N2022);
and AND3 (N2032, N2028, N550, N1121);
nor NOR2 (N2033, N2029, N871);
nor NOR3 (N2034, N2030, N1800, N1520);
and AND2 (N2035, N2024, N1023);
or OR2 (N2036, N2035, N1302);
xor XOR2 (N2037, N2008, N1247);
and AND4 (N2038, N2034, N1673, N245, N1761);
nand NAND3 (N2039, N2032, N1332, N910);
nand NAND3 (N2040, N2033, N1621, N1833);
buf BUF1 (N2041, N2037);
nor NOR3 (N2042, N2040, N59, N566);
xor XOR2 (N2043, N2041, N256);
buf BUF1 (N2044, N2027);
buf BUF1 (N2045, N2017);
not NOT1 (N2046, N2031);
nand NAND3 (N2047, N2042, N318, N1135);
and AND4 (N2048, N2047, N736, N304, N722);
xor XOR2 (N2049, N2048, N1770);
buf BUF1 (N2050, N2044);
not NOT1 (N2051, N2049);
or OR3 (N2052, N2043, N1120, N302);
nor NOR2 (N2053, N2046, N1408);
not NOT1 (N2054, N2039);
nand NAND2 (N2055, N2050, N566);
and AND4 (N2056, N2052, N1019, N368, N520);
xor XOR2 (N2057, N2056, N1627);
xor XOR2 (N2058, N2023, N1600);
nor NOR2 (N2059, N2051, N492);
nor NOR4 (N2060, N2045, N1478, N639, N740);
xor XOR2 (N2061, N2058, N1781);
xor XOR2 (N2062, N2059, N305);
buf BUF1 (N2063, N2061);
buf BUF1 (N2064, N2062);
buf BUF1 (N2065, N2038);
not NOT1 (N2066, N2054);
nand NAND2 (N2067, N2057, N86);
or OR3 (N2068, N2065, N1399, N715);
and AND4 (N2069, N2060, N1095, N725, N237);
not NOT1 (N2070, N2063);
buf BUF1 (N2071, N2068);
xor XOR2 (N2072, N2036, N1505);
nand NAND4 (N2073, N2072, N1509, N185, N1243);
and AND3 (N2074, N2066, N717, N614);
nand NAND3 (N2075, N2055, N139, N965);
buf BUF1 (N2076, N2067);
or OR3 (N2077, N2069, N1617, N1385);
nor NOR4 (N2078, N2073, N1294, N235, N1247);
or OR4 (N2079, N2064, N1870, N1106, N522);
nand NAND4 (N2080, N2079, N1663, N1798, N1305);
and AND4 (N2081, N2026, N622, N78, N703);
not NOT1 (N2082, N2081);
xor XOR2 (N2083, N2076, N1929);
and AND3 (N2084, N2077, N590, N833);
or OR2 (N2085, N2080, N1005);
or OR2 (N2086, N2071, N275);
and AND4 (N2087, N2053, N2047, N844, N1930);
not NOT1 (N2088, N2075);
or OR4 (N2089, N2074, N767, N1558, N82);
not NOT1 (N2090, N2089);
not NOT1 (N2091, N2087);
or OR2 (N2092, N2078, N370);
not NOT1 (N2093, N2091);
nand NAND2 (N2094, N2086, N738);
or OR3 (N2095, N2085, N1042, N1488);
xor XOR2 (N2096, N2070, N1601);
and AND3 (N2097, N2095, N1122, N737);
xor XOR2 (N2098, N2084, N760);
not NOT1 (N2099, N2094);
nor NOR3 (N2100, N2083, N162, N1977);
not NOT1 (N2101, N2093);
buf BUF1 (N2102, N2097);
or OR4 (N2103, N2100, N554, N1247, N2070);
or OR2 (N2104, N2092, N926);
nand NAND3 (N2105, N2099, N996, N1269);
or OR2 (N2106, N2098, N1117);
nand NAND4 (N2107, N2096, N2094, N1809, N1355);
and AND2 (N2108, N2103, N1926);
nand NAND3 (N2109, N2106, N1396, N1586);
or OR2 (N2110, N2101, N154);
nor NOR2 (N2111, N2102, N1583);
buf BUF1 (N2112, N2108);
and AND4 (N2113, N2107, N1076, N544, N765);
xor XOR2 (N2114, N2088, N766);
not NOT1 (N2115, N2111);
not NOT1 (N2116, N2114);
not NOT1 (N2117, N2082);
and AND4 (N2118, N2110, N2046, N1014, N2038);
nor NOR4 (N2119, N2109, N1064, N2083, N757);
xor XOR2 (N2120, N2116, N687);
xor XOR2 (N2121, N2113, N2045);
buf BUF1 (N2122, N2117);
nand NAND2 (N2123, N2090, N1748);
or OR2 (N2124, N2118, N1889);
and AND3 (N2125, N2112, N29, N1834);
nand NAND3 (N2126, N2119, N1542, N1789);
xor XOR2 (N2127, N2105, N883);
nor NOR3 (N2128, N2124, N1643, N1873);
xor XOR2 (N2129, N2128, N1345);
not NOT1 (N2130, N2127);
and AND3 (N2131, N2125, N798, N1077);
xor XOR2 (N2132, N2129, N665);
not NOT1 (N2133, N2132);
xor XOR2 (N2134, N2115, N1003);
and AND4 (N2135, N2134, N1841, N1077, N685);
or OR3 (N2136, N2120, N242, N385);
not NOT1 (N2137, N2123);
xor XOR2 (N2138, N2135, N1578);
or OR3 (N2139, N2126, N1230, N1826);
not NOT1 (N2140, N2137);
nor NOR2 (N2141, N2122, N993);
and AND4 (N2142, N2133, N756, N786, N335);
nand NAND4 (N2143, N2104, N298, N445, N1795);
or OR3 (N2144, N2130, N663, N1285);
xor XOR2 (N2145, N2138, N280);
nand NAND3 (N2146, N2139, N615, N10);
not NOT1 (N2147, N2144);
buf BUF1 (N2148, N2131);
buf BUF1 (N2149, N2147);
and AND2 (N2150, N2140, N1165);
and AND2 (N2151, N2148, N13);
xor XOR2 (N2152, N2145, N450);
nor NOR3 (N2153, N2142, N1628, N1170);
xor XOR2 (N2154, N2146, N1141);
xor XOR2 (N2155, N2149, N2054);
nand NAND2 (N2156, N2136, N1143);
not NOT1 (N2157, N2156);
nand NAND4 (N2158, N2155, N1977, N254, N814);
nand NAND4 (N2159, N2150, N1976, N2023, N578);
buf BUF1 (N2160, N2143);
xor XOR2 (N2161, N2121, N470);
buf BUF1 (N2162, N2157);
nor NOR2 (N2163, N2159, N737);
and AND3 (N2164, N2162, N1310, N279);
xor XOR2 (N2165, N2158, N1236);
xor XOR2 (N2166, N2153, N111);
and AND4 (N2167, N2160, N1623, N1487, N1245);
and AND2 (N2168, N2166, N1850);
or OR4 (N2169, N2154, N1514, N42, N1829);
and AND2 (N2170, N2152, N667);
and AND2 (N2171, N2167, N1850);
buf BUF1 (N2172, N2170);
nand NAND4 (N2173, N2165, N1770, N2163, N1416);
not NOT1 (N2174, N925);
xor XOR2 (N2175, N2151, N842);
and AND2 (N2176, N2161, N185);
and AND3 (N2177, N2172, N337, N364);
not NOT1 (N2178, N2164);
xor XOR2 (N2179, N2176, N403);
nor NOR4 (N2180, N2173, N1843, N293, N787);
nand NAND2 (N2181, N2177, N610);
not NOT1 (N2182, N2168);
or OR3 (N2183, N2181, N380, N532);
xor XOR2 (N2184, N2179, N90);
not NOT1 (N2185, N2184);
xor XOR2 (N2186, N2171, N214);
nand NAND4 (N2187, N2185, N1043, N472, N749);
xor XOR2 (N2188, N2187, N418);
nor NOR2 (N2189, N2180, N63);
nor NOR3 (N2190, N2174, N655, N1952);
nor NOR4 (N2191, N2178, N1661, N1181, N1077);
nand NAND3 (N2192, N2188, N1690, N1945);
not NOT1 (N2193, N2141);
and AND2 (N2194, N2186, N843);
nor NOR2 (N2195, N2190, N134);
nor NOR4 (N2196, N2194, N261, N110, N272);
nand NAND3 (N2197, N2193, N775, N1823);
nor NOR4 (N2198, N2169, N838, N1758, N2);
or OR2 (N2199, N2197, N1071);
buf BUF1 (N2200, N2198);
xor XOR2 (N2201, N2175, N546);
xor XOR2 (N2202, N2195, N174);
xor XOR2 (N2203, N2199, N1090);
not NOT1 (N2204, N2196);
or OR2 (N2205, N2201, N1502);
and AND3 (N2206, N2183, N1650, N770);
xor XOR2 (N2207, N2191, N2054);
and AND4 (N2208, N2200, N902, N1879, N1709);
buf BUF1 (N2209, N2202);
and AND4 (N2210, N2206, N1446, N103, N496);
xor XOR2 (N2211, N2182, N1948);
xor XOR2 (N2212, N2208, N1343);
and AND2 (N2213, N2205, N1041);
nor NOR4 (N2214, N2189, N1835, N646, N1294);
buf BUF1 (N2215, N2210);
xor XOR2 (N2216, N2212, N86);
xor XOR2 (N2217, N2211, N1546);
buf BUF1 (N2218, N2209);
buf BUF1 (N2219, N2217);
buf BUF1 (N2220, N2203);
nand NAND4 (N2221, N2215, N373, N1334, N1003);
nor NOR2 (N2222, N2207, N2054);
or OR3 (N2223, N2221, N2181, N408);
or OR2 (N2224, N2214, N271);
buf BUF1 (N2225, N2192);
buf BUF1 (N2226, N2224);
buf BUF1 (N2227, N2225);
nor NOR2 (N2228, N2204, N206);
or OR3 (N2229, N2219, N700, N2084);
not NOT1 (N2230, N2216);
nand NAND3 (N2231, N2222, N2, N1794);
xor XOR2 (N2232, N2213, N1228);
and AND2 (N2233, N2232, N674);
nand NAND2 (N2234, N2218, N1620);
or OR3 (N2235, N2227, N892, N311);
buf BUF1 (N2236, N2226);
nor NOR4 (N2237, N2228, N2163, N2216, N1938);
nor NOR2 (N2238, N2230, N1131);
and AND3 (N2239, N2234, N115, N1614);
and AND2 (N2240, N2236, N488);
xor XOR2 (N2241, N2231, N1060);
nor NOR2 (N2242, N2220, N785);
or OR3 (N2243, N2237, N1405, N2052);
nand NAND4 (N2244, N2229, N1963, N249, N1070);
nand NAND4 (N2245, N2238, N38, N1263, N157);
not NOT1 (N2246, N2239);
not NOT1 (N2247, N2223);
and AND4 (N2248, N2247, N756, N890, N155);
nand NAND4 (N2249, N2242, N797, N338, N630);
and AND4 (N2250, N2235, N95, N2040, N2121);
nand NAND2 (N2251, N2243, N1242);
not NOT1 (N2252, N2244);
nor NOR3 (N2253, N2245, N813, N161);
not NOT1 (N2254, N2233);
nand NAND3 (N2255, N2249, N320, N1285);
nor NOR3 (N2256, N2250, N1552, N1822);
or OR4 (N2257, N2240, N1336, N2099, N433);
and AND2 (N2258, N2241, N1142);
and AND2 (N2259, N2253, N1008);
xor XOR2 (N2260, N2258, N2139);
or OR2 (N2261, N2252, N2236);
nand NAND2 (N2262, N2259, N1749);
and AND2 (N2263, N2260, N287);
buf BUF1 (N2264, N2256);
nor NOR2 (N2265, N2261, N2238);
nand NAND4 (N2266, N2265, N1789, N433, N639);
not NOT1 (N2267, N2257);
nand NAND2 (N2268, N2262, N1384);
xor XOR2 (N2269, N2263, N427);
nor NOR2 (N2270, N2264, N2037);
nand NAND4 (N2271, N2251, N1912, N1552, N1877);
nor NOR2 (N2272, N2255, N93);
xor XOR2 (N2273, N2272, N205);
and AND2 (N2274, N2273, N2148);
not NOT1 (N2275, N2248);
xor XOR2 (N2276, N2271, N190);
and AND2 (N2277, N2267, N1521);
not NOT1 (N2278, N2276);
not NOT1 (N2279, N2254);
buf BUF1 (N2280, N2266);
not NOT1 (N2281, N2279);
not NOT1 (N2282, N2275);
and AND3 (N2283, N2281, N1415, N1297);
nand NAND3 (N2284, N2269, N1569, N1404);
xor XOR2 (N2285, N2284, N346);
nand NAND3 (N2286, N2285, N1761, N76);
and AND3 (N2287, N2274, N411, N1394);
buf BUF1 (N2288, N2286);
xor XOR2 (N2289, N2246, N852);
nand NAND4 (N2290, N2280, N1860, N248, N1832);
not NOT1 (N2291, N2290);
nor NOR3 (N2292, N2277, N2040, N2187);
and AND2 (N2293, N2287, N1095);
buf BUF1 (N2294, N2270);
not NOT1 (N2295, N2282);
nor NOR4 (N2296, N2283, N1250, N475, N392);
and AND2 (N2297, N2295, N1914);
buf BUF1 (N2298, N2288);
nor NOR3 (N2299, N2297, N1559, N824);
xor XOR2 (N2300, N2299, N1798);
buf BUF1 (N2301, N2294);
not NOT1 (N2302, N2301);
and AND4 (N2303, N2298, N1376, N1756, N1104);
nand NAND2 (N2304, N2296, N577);
nand NAND3 (N2305, N2278, N1882, N55);
or OR2 (N2306, N2305, N1221);
not NOT1 (N2307, N2306);
and AND3 (N2308, N2307, N1954, N1250);
buf BUF1 (N2309, N2303);
nand NAND4 (N2310, N2289, N1272, N2, N1477);
or OR2 (N2311, N2308, N2304);
buf BUF1 (N2312, N1971);
nand NAND3 (N2313, N2312, N1060, N1632);
buf BUF1 (N2314, N2313);
not NOT1 (N2315, N2300);
xor XOR2 (N2316, N2293, N1705);
and AND3 (N2317, N2302, N179, N688);
buf BUF1 (N2318, N2311);
xor XOR2 (N2319, N2314, N1308);
xor XOR2 (N2320, N2317, N909);
xor XOR2 (N2321, N2309, N2067);
not NOT1 (N2322, N2318);
nand NAND2 (N2323, N2315, N644);
nor NOR3 (N2324, N2310, N983, N875);
or OR4 (N2325, N2322, N1892, N1686, N1019);
or OR4 (N2326, N2291, N1415, N1377, N342);
buf BUF1 (N2327, N2321);
buf BUF1 (N2328, N2319);
nand NAND2 (N2329, N2268, N1805);
or OR3 (N2330, N2328, N1183, N630);
and AND2 (N2331, N2316, N2150);
xor XOR2 (N2332, N2320, N2331);
and AND4 (N2333, N1536, N2112, N425, N1936);
nand NAND2 (N2334, N2329, N1242);
or OR2 (N2335, N2334, N1854);
or OR2 (N2336, N2323, N1758);
xor XOR2 (N2337, N2333, N937);
buf BUF1 (N2338, N2335);
xor XOR2 (N2339, N2324, N1617);
and AND2 (N2340, N2330, N351);
xor XOR2 (N2341, N2338, N713);
and AND2 (N2342, N2332, N2065);
xor XOR2 (N2343, N2342, N992);
not NOT1 (N2344, N2292);
not NOT1 (N2345, N2340);
nor NOR4 (N2346, N2341, N1783, N1913, N2093);
nor NOR2 (N2347, N2343, N1525);
or OR3 (N2348, N2326, N1328, N1485);
nor NOR2 (N2349, N2337, N339);
xor XOR2 (N2350, N2349, N1810);
nor NOR2 (N2351, N2345, N2204);
or OR3 (N2352, N2346, N2279, N2042);
and AND2 (N2353, N2351, N605);
or OR3 (N2354, N2348, N902, N2242);
and AND2 (N2355, N2325, N817);
or OR2 (N2356, N2352, N167);
buf BUF1 (N2357, N2344);
not NOT1 (N2358, N2347);
nor NOR4 (N2359, N2350, N486, N827, N971);
nand NAND3 (N2360, N2336, N781, N128);
xor XOR2 (N2361, N2327, N1126);
xor XOR2 (N2362, N2354, N295);
nor NOR2 (N2363, N2339, N2215);
xor XOR2 (N2364, N2359, N1059);
buf BUF1 (N2365, N2355);
and AND4 (N2366, N2360, N1430, N2204, N1737);
or OR4 (N2367, N2363, N236, N760, N69);
and AND3 (N2368, N2353, N1815, N884);
nand NAND2 (N2369, N2357, N1436);
nor NOR4 (N2370, N2362, N1961, N1286, N522);
xor XOR2 (N2371, N2361, N874);
and AND4 (N2372, N2358, N286, N147, N336);
buf BUF1 (N2373, N2365);
not NOT1 (N2374, N2373);
and AND3 (N2375, N2371, N634, N843);
nand NAND2 (N2376, N2374, N738);
or OR2 (N2377, N2369, N1776);
buf BUF1 (N2378, N2367);
and AND4 (N2379, N2372, N740, N1889, N1992);
xor XOR2 (N2380, N2356, N1330);
nand NAND2 (N2381, N2368, N1612);
nor NOR4 (N2382, N2364, N1264, N1532, N862);
nor NOR2 (N2383, N2379, N2298);
nand NAND4 (N2384, N2378, N1853, N172, N223);
and AND4 (N2385, N2366, N79, N1602, N1076);
or OR3 (N2386, N2380, N930, N968);
or OR2 (N2387, N2385, N158);
and AND2 (N2388, N2381, N1295);
not NOT1 (N2389, N2370);
xor XOR2 (N2390, N2383, N96);
or OR2 (N2391, N2388, N234);
not NOT1 (N2392, N2386);
xor XOR2 (N2393, N2377, N590);
and AND2 (N2394, N2390, N166);
or OR4 (N2395, N2382, N632, N1626, N1745);
nand NAND4 (N2396, N2393, N1562, N1147, N294);
or OR3 (N2397, N2391, N1636, N1238);
nor NOR2 (N2398, N2395, N2335);
nor NOR2 (N2399, N2396, N1286);
or OR3 (N2400, N2392, N1634, N1694);
not NOT1 (N2401, N2397);
buf BUF1 (N2402, N2399);
buf BUF1 (N2403, N2401);
nand NAND4 (N2404, N2384, N736, N1427, N1291);
nor NOR3 (N2405, N2404, N2326, N1840);
buf BUF1 (N2406, N2398);
or OR3 (N2407, N2389, N1502, N1535);
or OR2 (N2408, N2375, N2045);
xor XOR2 (N2409, N2394, N1492);
or OR4 (N2410, N2403, N763, N955, N1678);
nand NAND3 (N2411, N2400, N1589, N951);
nand NAND3 (N2412, N2376, N423, N669);
or OR3 (N2413, N2407, N1709, N129);
not NOT1 (N2414, N2387);
nand NAND4 (N2415, N2413, N991, N2140, N1808);
or OR3 (N2416, N2408, N39, N1976);
not NOT1 (N2417, N2416);
or OR3 (N2418, N2411, N1646, N796);
nand NAND3 (N2419, N2412, N64, N697);
nor NOR2 (N2420, N2419, N827);
buf BUF1 (N2421, N2418);
and AND2 (N2422, N2417, N1923);
nand NAND3 (N2423, N2409, N856, N2221);
buf BUF1 (N2424, N2405);
not NOT1 (N2425, N2402);
buf BUF1 (N2426, N2415);
nor NOR3 (N2427, N2414, N868, N2101);
nor NOR4 (N2428, N2420, N766, N275, N1973);
nand NAND2 (N2429, N2425, N1151);
xor XOR2 (N2430, N2410, N697);
nor NOR3 (N2431, N2421, N773, N1060);
xor XOR2 (N2432, N2430, N1951);
or OR4 (N2433, N2429, N1853, N1717, N1771);
xor XOR2 (N2434, N2426, N1931);
xor XOR2 (N2435, N2406, N1468);
xor XOR2 (N2436, N2428, N2184);
or OR2 (N2437, N2434, N1802);
nand NAND4 (N2438, N2432, N1734, N1775, N409);
nand NAND3 (N2439, N2431, N1170, N2040);
and AND2 (N2440, N2427, N1240);
xor XOR2 (N2441, N2423, N1452);
not NOT1 (N2442, N2435);
and AND4 (N2443, N2442, N777, N2068, N213);
or OR2 (N2444, N2424, N1351);
nor NOR4 (N2445, N2441, N1976, N1360, N77);
xor XOR2 (N2446, N2443, N2069);
or OR4 (N2447, N2438, N1925, N2021, N499);
and AND3 (N2448, N2433, N1652, N363);
nor NOR4 (N2449, N2422, N1681, N1273, N1928);
nand NAND3 (N2450, N2447, N632, N2172);
xor XOR2 (N2451, N2444, N883);
and AND3 (N2452, N2437, N1657, N343);
nor NOR2 (N2453, N2449, N2201);
not NOT1 (N2454, N2450);
not NOT1 (N2455, N2440);
nand NAND2 (N2456, N2452, N65);
nor NOR3 (N2457, N2453, N563, N675);
xor XOR2 (N2458, N2446, N1175);
not NOT1 (N2459, N2451);
or OR2 (N2460, N2458, N355);
buf BUF1 (N2461, N2459);
or OR3 (N2462, N2448, N193, N1473);
not NOT1 (N2463, N2445);
not NOT1 (N2464, N2457);
or OR3 (N2465, N2439, N48, N1094);
nand NAND3 (N2466, N2436, N2182, N87);
xor XOR2 (N2467, N2465, N1868);
and AND2 (N2468, N2463, N1806);
buf BUF1 (N2469, N2466);
not NOT1 (N2470, N2460);
or OR2 (N2471, N2467, N85);
and AND3 (N2472, N2469, N377, N966);
not NOT1 (N2473, N2471);
or OR3 (N2474, N2470, N225, N986);
nor NOR3 (N2475, N2454, N1582, N888);
buf BUF1 (N2476, N2456);
nor NOR4 (N2477, N2462, N504, N71, N1964);
nand NAND3 (N2478, N2474, N267, N435);
buf BUF1 (N2479, N2478);
xor XOR2 (N2480, N2455, N1487);
and AND2 (N2481, N2475, N1766);
nand NAND2 (N2482, N2476, N886);
xor XOR2 (N2483, N2464, N1594);
nor NOR4 (N2484, N2483, N360, N1042, N869);
xor XOR2 (N2485, N2484, N582);
not NOT1 (N2486, N2473);
and AND4 (N2487, N2461, N594, N1500, N1676);
not NOT1 (N2488, N2468);
buf BUF1 (N2489, N2480);
buf BUF1 (N2490, N2472);
buf BUF1 (N2491, N2490);
and AND3 (N2492, N2489, N530, N627);
buf BUF1 (N2493, N2477);
not NOT1 (N2494, N2488);
and AND3 (N2495, N2487, N1353, N728);
xor XOR2 (N2496, N2493, N155);
and AND2 (N2497, N2481, N1076);
and AND3 (N2498, N2494, N2457, N94);
xor XOR2 (N2499, N2485, N1290);
nand NAND3 (N2500, N2486, N1518, N1297);
and AND2 (N2501, N2491, N1407);
nor NOR3 (N2502, N2495, N1445, N1344);
not NOT1 (N2503, N2502);
or OR3 (N2504, N2499, N2476, N1074);
xor XOR2 (N2505, N2504, N2435);
nor NOR3 (N2506, N2501, N2492, N2403);
nor NOR3 (N2507, N1868, N1528, N943);
xor XOR2 (N2508, N2500, N1883);
nor NOR4 (N2509, N2496, N738, N749, N1022);
buf BUF1 (N2510, N2509);
and AND4 (N2511, N2498, N66, N2202, N696);
nor NOR2 (N2512, N2505, N1625);
buf BUF1 (N2513, N2511);
and AND4 (N2514, N2510, N1320, N1195, N239);
buf BUF1 (N2515, N2497);
nor NOR2 (N2516, N2503, N126);
and AND3 (N2517, N2507, N647, N1731);
xor XOR2 (N2518, N2508, N1367);
nor NOR3 (N2519, N2516, N2153, N484);
and AND4 (N2520, N2479, N313, N951, N782);
nor NOR2 (N2521, N2517, N873);
not NOT1 (N2522, N2520);
buf BUF1 (N2523, N2519);
xor XOR2 (N2524, N2518, N1522);
nor NOR4 (N2525, N2506, N1025, N1304, N107);
nand NAND4 (N2526, N2521, N1644, N2174, N1848);
or OR4 (N2527, N2513, N1018, N159, N1291);
xor XOR2 (N2528, N2527, N2133);
buf BUF1 (N2529, N2482);
xor XOR2 (N2530, N2524, N458);
nand NAND3 (N2531, N2526, N213, N1289);
xor XOR2 (N2532, N2515, N1254);
and AND3 (N2533, N2532, N1509, N1599);
and AND2 (N2534, N2528, N1816);
xor XOR2 (N2535, N2531, N952);
nand NAND3 (N2536, N2525, N1672, N138);
or OR3 (N2537, N2512, N1947, N1701);
buf BUF1 (N2538, N2522);
xor XOR2 (N2539, N2514, N2163);
buf BUF1 (N2540, N2536);
or OR4 (N2541, N2537, N1967, N1337, N914);
and AND2 (N2542, N2541, N2219);
nor NOR2 (N2543, N2530, N1061);
or OR2 (N2544, N2534, N572);
buf BUF1 (N2545, N2538);
nor NOR3 (N2546, N2529, N1217, N258);
or OR4 (N2547, N2545, N1439, N803, N1817);
and AND4 (N2548, N2544, N1383, N1190, N2211);
buf BUF1 (N2549, N2548);
and AND2 (N2550, N2543, N171);
buf BUF1 (N2551, N2549);
buf BUF1 (N2552, N2533);
and AND4 (N2553, N2535, N2326, N1528, N1912);
xor XOR2 (N2554, N2540, N1473);
nor NOR3 (N2555, N2551, N669, N862);
buf BUF1 (N2556, N2539);
xor XOR2 (N2557, N2550, N260);
nand NAND2 (N2558, N2547, N132);
and AND3 (N2559, N2557, N1316, N2438);
xor XOR2 (N2560, N2554, N415);
nor NOR3 (N2561, N2553, N2102, N2400);
buf BUF1 (N2562, N2523);
nor NOR4 (N2563, N2560, N1573, N874, N1500);
and AND2 (N2564, N2542, N1947);
nand NAND4 (N2565, N2563, N2377, N1078, N1686);
and AND2 (N2566, N2558, N894);
not NOT1 (N2567, N2559);
and AND3 (N2568, N2552, N1719, N2484);
xor XOR2 (N2569, N2567, N2);
and AND4 (N2570, N2568, N349, N810, N1796);
or OR2 (N2571, N2562, N993);
buf BUF1 (N2572, N2570);
nor NOR2 (N2573, N2572, N477);
or OR4 (N2574, N2564, N1998, N2071, N1852);
and AND2 (N2575, N2555, N1781);
xor XOR2 (N2576, N2546, N780);
not NOT1 (N2577, N2573);
not NOT1 (N2578, N2576);
nor NOR2 (N2579, N2569, N36);
not NOT1 (N2580, N2566);
nor NOR4 (N2581, N2577, N2209, N475, N138);
or OR4 (N2582, N2556, N1073, N531, N747);
and AND4 (N2583, N2580, N92, N1142, N1331);
or OR4 (N2584, N2561, N1197, N1333, N2074);
nand NAND2 (N2585, N2565, N1976);
nand NAND3 (N2586, N2584, N2235, N2387);
not NOT1 (N2587, N2575);
buf BUF1 (N2588, N2571);
xor XOR2 (N2589, N2574, N1892);
buf BUF1 (N2590, N2582);
buf BUF1 (N2591, N2590);
xor XOR2 (N2592, N2583, N2241);
nor NOR4 (N2593, N2586, N1916, N387, N411);
and AND4 (N2594, N2591, N2055, N1968, N861);
nand NAND4 (N2595, N2592, N832, N2445, N2540);
buf BUF1 (N2596, N2581);
nand NAND4 (N2597, N2594, N784, N120, N96);
and AND2 (N2598, N2578, N2006);
buf BUF1 (N2599, N2597);
not NOT1 (N2600, N2596);
xor XOR2 (N2601, N2600, N1496);
and AND4 (N2602, N2601, N2030, N807, N1254);
buf BUF1 (N2603, N2595);
and AND2 (N2604, N2598, N918);
and AND4 (N2605, N2585, N754, N1298, N387);
buf BUF1 (N2606, N2588);
not NOT1 (N2607, N2593);
xor XOR2 (N2608, N2599, N2442);
nor NOR3 (N2609, N2602, N1558, N2448);
not NOT1 (N2610, N2607);
or OR4 (N2611, N2610, N1521, N2455, N1582);
and AND4 (N2612, N2609, N409, N2318, N2303);
or OR2 (N2613, N2608, N1111);
buf BUF1 (N2614, N2589);
nand NAND2 (N2615, N2611, N1634);
xor XOR2 (N2616, N2615, N419);
and AND4 (N2617, N2612, N1562, N2046, N2582);
or OR2 (N2618, N2604, N1153);
nand NAND2 (N2619, N2587, N2205);
nand NAND4 (N2620, N2618, N1324, N2366, N1173);
and AND3 (N2621, N2579, N439, N174);
buf BUF1 (N2622, N2613);
buf BUF1 (N2623, N2603);
and AND2 (N2624, N2614, N1459);
not NOT1 (N2625, N2617);
or OR4 (N2626, N2619, N1209, N1095, N1797);
nand NAND3 (N2627, N2623, N1565, N940);
buf BUF1 (N2628, N2625);
xor XOR2 (N2629, N2621, N914);
and AND4 (N2630, N2627, N286, N960, N2439);
nor NOR2 (N2631, N2616, N816);
nand NAND2 (N2632, N2630, N298);
not NOT1 (N2633, N2629);
nand NAND2 (N2634, N2622, N1293);
nand NAND3 (N2635, N2634, N1820, N1003);
not NOT1 (N2636, N2605);
nor NOR2 (N2637, N2620, N1577);
or OR4 (N2638, N2636, N2010, N833, N468);
xor XOR2 (N2639, N2637, N1714);
not NOT1 (N2640, N2606);
buf BUF1 (N2641, N2638);
nand NAND4 (N2642, N2639, N1171, N521, N1719);
xor XOR2 (N2643, N2640, N2596);
nand NAND4 (N2644, N2626, N1833, N1541, N527);
and AND2 (N2645, N2641, N1162);
buf BUF1 (N2646, N2624);
xor XOR2 (N2647, N2645, N728);
or OR4 (N2648, N2642, N2058, N414, N1524);
xor XOR2 (N2649, N2647, N1363);
not NOT1 (N2650, N2635);
and AND2 (N2651, N2631, N1951);
buf BUF1 (N2652, N2648);
not NOT1 (N2653, N2651);
xor XOR2 (N2654, N2633, N1387);
xor XOR2 (N2655, N2649, N216);
or OR4 (N2656, N2652, N2617, N1040, N400);
nor NOR4 (N2657, N2628, N1924, N1764, N649);
nand NAND2 (N2658, N2654, N1926);
or OR4 (N2659, N2655, N1444, N365, N2464);
buf BUF1 (N2660, N2650);
buf BUF1 (N2661, N2646);
nand NAND4 (N2662, N2643, N2435, N2447, N1302);
not NOT1 (N2663, N2656);
nand NAND4 (N2664, N2660, N2349, N1200, N2480);
buf BUF1 (N2665, N2632);
or OR2 (N2666, N2663, N1394);
not NOT1 (N2667, N2666);
nand NAND4 (N2668, N2665, N2250, N1819, N2299);
xor XOR2 (N2669, N2664, N1640);
nand NAND4 (N2670, N2668, N1577, N1969, N2569);
and AND4 (N2671, N2657, N541, N762, N1967);
nor NOR3 (N2672, N2667, N571, N2094);
or OR4 (N2673, N2653, N541, N1234, N2080);
nor NOR3 (N2674, N2671, N2039, N1762);
or OR3 (N2675, N2658, N2024, N1941);
or OR4 (N2676, N2661, N2130, N2573, N1574);
and AND4 (N2677, N2662, N2350, N2396, N87);
and AND3 (N2678, N2674, N2593, N2191);
or OR4 (N2679, N2678, N2229, N1332, N544);
and AND3 (N2680, N2673, N149, N230);
or OR3 (N2681, N2644, N1593, N2159);
or OR4 (N2682, N2670, N1014, N1861, N495);
nand NAND4 (N2683, N2675, N1324, N176, N440);
xor XOR2 (N2684, N2681, N892);
and AND2 (N2685, N2682, N217);
xor XOR2 (N2686, N2679, N1041);
nor NOR3 (N2687, N2680, N1046, N1689);
xor XOR2 (N2688, N2676, N2488);
buf BUF1 (N2689, N2677);
and AND3 (N2690, N2689, N493, N1003);
xor XOR2 (N2691, N2686, N991);
and AND3 (N2692, N2669, N1538, N1319);
and AND3 (N2693, N2684, N275, N1657);
nor NOR3 (N2694, N2687, N2002, N1621);
or OR4 (N2695, N2691, N1599, N2528, N1272);
xor XOR2 (N2696, N2672, N2680);
buf BUF1 (N2697, N2688);
not NOT1 (N2698, N2685);
nand NAND4 (N2699, N2659, N516, N2631, N1933);
nand NAND4 (N2700, N2690, N28, N2227, N679);
buf BUF1 (N2701, N2692);
and AND3 (N2702, N2693, N1248, N2355);
nor NOR3 (N2703, N2700, N801, N1965);
buf BUF1 (N2704, N2703);
buf BUF1 (N2705, N2694);
and AND3 (N2706, N2696, N407, N73);
or OR3 (N2707, N2697, N1090, N1020);
not NOT1 (N2708, N2704);
not NOT1 (N2709, N2695);
buf BUF1 (N2710, N2705);
and AND3 (N2711, N2683, N1113, N547);
xor XOR2 (N2712, N2701, N1768);
nor NOR4 (N2713, N2708, N393, N1326, N2466);
nand NAND2 (N2714, N2711, N2217);
buf BUF1 (N2715, N2702);
nor NOR3 (N2716, N2707, N1633, N2340);
nor NOR2 (N2717, N2699, N1813);
or OR2 (N2718, N2713, N1908);
nand NAND3 (N2719, N2710, N2100, N2245);
and AND3 (N2720, N2698, N728, N127);
not NOT1 (N2721, N2717);
xor XOR2 (N2722, N2721, N1296);
nand NAND3 (N2723, N2706, N943, N129);
or OR2 (N2724, N2716, N167);
nor NOR3 (N2725, N2722, N1303, N1979);
and AND2 (N2726, N2724, N827);
or OR3 (N2727, N2726, N1586, N1179);
nand NAND4 (N2728, N2727, N1266, N890, N1419);
or OR2 (N2729, N2709, N1931);
not NOT1 (N2730, N2719);
nand NAND4 (N2731, N2728, N1225, N2552, N1799);
nor NOR2 (N2732, N2712, N809);
buf BUF1 (N2733, N2718);
xor XOR2 (N2734, N2731, N659);
xor XOR2 (N2735, N2720, N2612);
buf BUF1 (N2736, N2715);
buf BUF1 (N2737, N2714);
nor NOR2 (N2738, N2734, N1124);
and AND2 (N2739, N2725, N1229);
not NOT1 (N2740, N2735);
not NOT1 (N2741, N2739);
or OR3 (N2742, N2733, N567, N1641);
not NOT1 (N2743, N2729);
and AND2 (N2744, N2741, N1063);
nand NAND2 (N2745, N2730, N2134);
or OR2 (N2746, N2742, N1357);
nor NOR4 (N2747, N2743, N220, N1459, N2168);
nor NOR4 (N2748, N2747, N1927, N619, N639);
nand NAND3 (N2749, N2748, N1926, N1403);
or OR2 (N2750, N2737, N208);
buf BUF1 (N2751, N2740);
or OR3 (N2752, N2745, N21, N778);
nand NAND2 (N2753, N2744, N782);
xor XOR2 (N2754, N2738, N2602);
or OR4 (N2755, N2746, N665, N875, N977);
or OR2 (N2756, N2752, N1780);
not NOT1 (N2757, N2754);
nand NAND3 (N2758, N2755, N2687, N1658);
nor NOR3 (N2759, N2756, N2248, N890);
and AND4 (N2760, N2759, N2254, N1454, N819);
nand NAND2 (N2761, N2753, N1863);
xor XOR2 (N2762, N2751, N148);
xor XOR2 (N2763, N2732, N2187);
xor XOR2 (N2764, N2723, N2406);
and AND3 (N2765, N2750, N612, N1351);
nand NAND3 (N2766, N2764, N1875, N1933);
buf BUF1 (N2767, N2757);
or OR4 (N2768, N2761, N1034, N145, N1831);
buf BUF1 (N2769, N2749);
xor XOR2 (N2770, N2763, N1602);
and AND2 (N2771, N2765, N2437);
nand NAND4 (N2772, N2766, N956, N114, N727);
not NOT1 (N2773, N2770);
or OR4 (N2774, N2771, N872, N1482, N2497);
nand NAND2 (N2775, N2772, N464);
nor NOR4 (N2776, N2736, N1267, N1145, N432);
and AND3 (N2777, N2767, N2496, N2285);
xor XOR2 (N2778, N2758, N1216);
and AND4 (N2779, N2768, N1255, N871, N1132);
nand NAND2 (N2780, N2762, N1773);
nor NOR3 (N2781, N2774, N1356, N1975);
nand NAND3 (N2782, N2769, N1780, N1233);
and AND3 (N2783, N2777, N731, N1665);
or OR4 (N2784, N2783, N1803, N423, N2019);
not NOT1 (N2785, N2779);
not NOT1 (N2786, N2781);
not NOT1 (N2787, N2785);
and AND4 (N2788, N2776, N1600, N1141, N1102);
buf BUF1 (N2789, N2782);
nand NAND3 (N2790, N2787, N2403, N2629);
or OR3 (N2791, N2778, N1713, N471);
nand NAND2 (N2792, N2788, N2559);
nor NOR3 (N2793, N2784, N676, N2160);
nand NAND2 (N2794, N2789, N1467);
and AND2 (N2795, N2760, N29);
nor NOR2 (N2796, N2793, N1364);
xor XOR2 (N2797, N2775, N474);
nand NAND2 (N2798, N2786, N2716);
nor NOR2 (N2799, N2795, N1649);
or OR3 (N2800, N2773, N2054, N1241);
xor XOR2 (N2801, N2796, N1133);
nand NAND3 (N2802, N2792, N1169, N594);
not NOT1 (N2803, N2801);
nand NAND4 (N2804, N2800, N2663, N1177, N2198);
nand NAND3 (N2805, N2798, N2732, N2266);
nor NOR4 (N2806, N2804, N2735, N1436, N1458);
xor XOR2 (N2807, N2805, N1269);
or OR2 (N2808, N2806, N81);
and AND4 (N2809, N2799, N956, N1509, N378);
xor XOR2 (N2810, N2807, N1663);
nand NAND2 (N2811, N2808, N2573);
and AND3 (N2812, N2810, N650, N2042);
nand NAND4 (N2813, N2802, N1472, N1630, N2411);
buf BUF1 (N2814, N2811);
buf BUF1 (N2815, N2812);
nor NOR2 (N2816, N2797, N919);
buf BUF1 (N2817, N2809);
nand NAND3 (N2818, N2791, N476, N2246);
nor NOR4 (N2819, N2815, N2785, N923, N1467);
or OR4 (N2820, N2780, N713, N1925, N454);
xor XOR2 (N2821, N2790, N1905);
nor NOR2 (N2822, N2819, N1161);
xor XOR2 (N2823, N2821, N1589);
and AND3 (N2824, N2823, N2494, N214);
nand NAND4 (N2825, N2816, N855, N1306, N604);
and AND4 (N2826, N2824, N50, N558, N1210);
buf BUF1 (N2827, N2820);
or OR3 (N2828, N2827, N890, N1982);
buf BUF1 (N2829, N2818);
and AND2 (N2830, N2825, N2177);
xor XOR2 (N2831, N2803, N1595);
not NOT1 (N2832, N2817);
nor NOR4 (N2833, N2828, N267, N458, N2260);
nand NAND2 (N2834, N2830, N1000);
not NOT1 (N2835, N2822);
buf BUF1 (N2836, N2829);
nand NAND4 (N2837, N2794, N1456, N1847, N2590);
nand NAND3 (N2838, N2835, N1497, N194);
not NOT1 (N2839, N2813);
nand NAND2 (N2840, N2836, N2768);
xor XOR2 (N2841, N2834, N1209);
and AND3 (N2842, N2833, N1035, N1406);
and AND3 (N2843, N2826, N1230, N95);
nor NOR2 (N2844, N2832, N2059);
buf BUF1 (N2845, N2841);
nor NOR2 (N2846, N2845, N1195);
or OR3 (N2847, N2838, N1132, N1665);
buf BUF1 (N2848, N2843);
nand NAND4 (N2849, N2848, N2416, N557, N1900);
and AND2 (N2850, N2839, N984);
or OR2 (N2851, N2837, N1200);
buf BUF1 (N2852, N2840);
and AND3 (N2853, N2849, N1544, N275);
or OR3 (N2854, N2814, N2526, N841);
not NOT1 (N2855, N2854);
xor XOR2 (N2856, N2851, N2192);
and AND4 (N2857, N2856, N2234, N2066, N389);
nand NAND3 (N2858, N2846, N392, N2250);
and AND3 (N2859, N2847, N1833, N1821);
and AND4 (N2860, N2857, N2224, N848, N1315);
nand NAND3 (N2861, N2859, N567, N24);
nor NOR3 (N2862, N2850, N1153, N2442);
buf BUF1 (N2863, N2862);
not NOT1 (N2864, N2860);
nor NOR3 (N2865, N2855, N667, N1254);
nand NAND2 (N2866, N2864, N2731);
nor NOR4 (N2867, N2852, N2469, N142, N2566);
xor XOR2 (N2868, N2831, N1336);
nand NAND3 (N2869, N2863, N5, N747);
nor NOR3 (N2870, N2842, N1509, N2240);
buf BUF1 (N2871, N2865);
nand NAND4 (N2872, N2853, N49, N2480, N2224);
xor XOR2 (N2873, N2858, N367);
and AND2 (N2874, N2867, N1276);
nor NOR4 (N2875, N2874, N546, N1531, N2267);
nand NAND4 (N2876, N2869, N1444, N2520, N1039);
nand NAND2 (N2877, N2871, N781);
nand NAND2 (N2878, N2877, N179);
nor NOR4 (N2879, N2876, N303, N1467, N350);
nand NAND3 (N2880, N2866, N2191, N2715);
and AND4 (N2881, N2870, N1293, N2268, N836);
buf BUF1 (N2882, N2861);
buf BUF1 (N2883, N2844);
not NOT1 (N2884, N2875);
xor XOR2 (N2885, N2881, N2281);
or OR2 (N2886, N2884, N39);
nand NAND2 (N2887, N2883, N1677);
nand NAND4 (N2888, N2878, N2548, N1942, N2217);
nand NAND2 (N2889, N2880, N1806);
nor NOR2 (N2890, N2872, N2163);
nor NOR3 (N2891, N2889, N311, N2426);
or OR3 (N2892, N2879, N1974, N2730);
buf BUF1 (N2893, N2892);
xor XOR2 (N2894, N2893, N2185);
and AND4 (N2895, N2891, N2752, N2005, N2409);
buf BUF1 (N2896, N2895);
buf BUF1 (N2897, N2887);
nor NOR2 (N2898, N2888, N2726);
xor XOR2 (N2899, N2896, N1506);
nor NOR4 (N2900, N2885, N1738, N586, N2749);
not NOT1 (N2901, N2886);
xor XOR2 (N2902, N2868, N1238);
nand NAND3 (N2903, N2873, N2773, N1988);
nor NOR4 (N2904, N2901, N1612, N1733, N1522);
nand NAND4 (N2905, N2897, N41, N2550, N1793);
buf BUF1 (N2906, N2900);
buf BUF1 (N2907, N2899);
nand NAND4 (N2908, N2906, N2238, N1294, N1511);
nand NAND2 (N2909, N2908, N1989);
not NOT1 (N2910, N2905);
xor XOR2 (N2911, N2882, N2037);
nor NOR2 (N2912, N2909, N161);
buf BUF1 (N2913, N2898);
xor XOR2 (N2914, N2903, N1102);
nand NAND2 (N2915, N2907, N1912);
and AND4 (N2916, N2915, N1545, N2278, N929);
buf BUF1 (N2917, N2916);
nand NAND3 (N2918, N2914, N64, N1541);
xor XOR2 (N2919, N2904, N2386);
xor XOR2 (N2920, N2911, N829);
xor XOR2 (N2921, N2918, N271);
not NOT1 (N2922, N2912);
and AND3 (N2923, N2921, N1521, N2757);
nand NAND4 (N2924, N2902, N2112, N508, N1177);
and AND2 (N2925, N2924, N227);
buf BUF1 (N2926, N2920);
or OR4 (N2927, N2890, N316, N660, N53);
not NOT1 (N2928, N2925);
and AND3 (N2929, N2919, N2122, N1986);
nor NOR2 (N2930, N2922, N721);
not NOT1 (N2931, N2926);
not NOT1 (N2932, N2927);
not NOT1 (N2933, N2931);
or OR2 (N2934, N2923, N1985);
nor NOR2 (N2935, N2934, N2404);
or OR4 (N2936, N2913, N1340, N1511, N2499);
and AND4 (N2937, N2917, N257, N2275, N323);
nand NAND4 (N2938, N2936, N1028, N1425, N1973);
and AND4 (N2939, N2930, N1216, N2935, N1442);
and AND2 (N2940, N237, N3);
xor XOR2 (N2941, N2940, N598);
xor XOR2 (N2942, N2910, N746);
or OR2 (N2943, N2938, N751);
not NOT1 (N2944, N2939);
not NOT1 (N2945, N2943);
and AND3 (N2946, N2944, N748, N1904);
buf BUF1 (N2947, N2946);
and AND2 (N2948, N2928, N1961);
buf BUF1 (N2949, N2933);
or OR3 (N2950, N2941, N2824, N2796);
not NOT1 (N2951, N2942);
nand NAND2 (N2952, N2948, N1894);
nor NOR2 (N2953, N2937, N2354);
nor NOR2 (N2954, N2894, N1965);
or OR2 (N2955, N2950, N2135);
nand NAND3 (N2956, N2954, N2250, N1596);
nand NAND3 (N2957, N2953, N2794, N2620);
buf BUF1 (N2958, N2932);
nand NAND2 (N2959, N2949, N50);
buf BUF1 (N2960, N2959);
xor XOR2 (N2961, N2929, N1781);
nor NOR4 (N2962, N2958, N1537, N394, N56);
buf BUF1 (N2963, N2955);
buf BUF1 (N2964, N2961);
xor XOR2 (N2965, N2963, N1346);
xor XOR2 (N2966, N2952, N2476);
nand NAND4 (N2967, N2947, N911, N2281, N666);
not NOT1 (N2968, N2945);
nand NAND3 (N2969, N2956, N245, N1180);
or OR3 (N2970, N2964, N2959, N1150);
or OR4 (N2971, N2965, N1563, N172, N215);
nor NOR3 (N2972, N2960, N1807, N1819);
nand NAND4 (N2973, N2968, N349, N249, N906);
and AND2 (N2974, N2973, N1894);
or OR4 (N2975, N2970, N1759, N2606, N303);
not NOT1 (N2976, N2971);
nand NAND3 (N2977, N2976, N751, N1918);
and AND4 (N2978, N2957, N2516, N2083, N1949);
xor XOR2 (N2979, N2972, N2040);
buf BUF1 (N2980, N2975);
not NOT1 (N2981, N2966);
buf BUF1 (N2982, N2951);
not NOT1 (N2983, N2978);
not NOT1 (N2984, N2983);
not NOT1 (N2985, N2981);
or OR2 (N2986, N2977, N1241);
xor XOR2 (N2987, N2974, N1140);
buf BUF1 (N2988, N2967);
not NOT1 (N2989, N2969);
nor NOR2 (N2990, N2980, N283);
nor NOR3 (N2991, N2990, N264, N1820);
xor XOR2 (N2992, N2989, N695);
nor NOR3 (N2993, N2979, N1042, N1357);
xor XOR2 (N2994, N2962, N2456);
xor XOR2 (N2995, N2987, N1932);
nand NAND4 (N2996, N2984, N1187, N128, N1494);
not NOT1 (N2997, N2985);
nor NOR4 (N2998, N2995, N1343, N2670, N457);
nand NAND4 (N2999, N2988, N910, N2051, N2673);
nand NAND3 (N3000, N2996, N1, N270);
nor NOR2 (N3001, N3000, N1760);
nand NAND4 (N3002, N3001, N1547, N2683, N317);
buf BUF1 (N3003, N2994);
or OR3 (N3004, N2998, N2299, N1820);
not NOT1 (N3005, N2992);
nor NOR3 (N3006, N2982, N560, N2468);
buf BUF1 (N3007, N3002);
xor XOR2 (N3008, N2993, N1495);
nor NOR3 (N3009, N2999, N2902, N258);
nand NAND3 (N3010, N3009, N127, N731);
xor XOR2 (N3011, N2997, N1760);
and AND2 (N3012, N3007, N1820);
xor XOR2 (N3013, N3012, N743);
nor NOR3 (N3014, N3006, N1475, N2710);
or OR2 (N3015, N2986, N773);
nor NOR3 (N3016, N3011, N1135, N1183);
or OR3 (N3017, N3005, N2243, N697);
not NOT1 (N3018, N3016);
and AND2 (N3019, N3018, N554);
nor NOR2 (N3020, N3013, N2507);
buf BUF1 (N3021, N3020);
buf BUF1 (N3022, N3019);
xor XOR2 (N3023, N3010, N2963);
and AND2 (N3024, N3017, N1255);
nor NOR4 (N3025, N3021, N1991, N998, N2513);
not NOT1 (N3026, N2991);
not NOT1 (N3027, N3014);
or OR3 (N3028, N3027, N1645, N845);
nor NOR2 (N3029, N3023, N573);
not NOT1 (N3030, N3015);
or OR4 (N3031, N3003, N2278, N49, N627);
not NOT1 (N3032, N3030);
and AND2 (N3033, N3031, N1241);
or OR2 (N3034, N3024, N2519);
or OR3 (N3035, N3025, N1358, N1703);
nand NAND4 (N3036, N3032, N1413, N1083, N1192);
and AND2 (N3037, N3029, N289);
xor XOR2 (N3038, N3028, N179);
nand NAND2 (N3039, N3004, N1606);
nor NOR4 (N3040, N3033, N1397, N41, N254);
buf BUF1 (N3041, N3022);
nor NOR4 (N3042, N3037, N1857, N549, N2138);
or OR2 (N3043, N3034, N174);
and AND2 (N3044, N3038, N2932);
nand NAND4 (N3045, N3043, N36, N1536, N404);
not NOT1 (N3046, N3035);
not NOT1 (N3047, N3008);
nor NOR3 (N3048, N3046, N813, N353);
not NOT1 (N3049, N3036);
and AND3 (N3050, N3042, N1492, N1121);
nand NAND4 (N3051, N3044, N2032, N2410, N1581);
nand NAND3 (N3052, N3049, N1231, N1172);
not NOT1 (N3053, N3026);
not NOT1 (N3054, N3051);
or OR4 (N3055, N3050, N455, N764, N788);
or OR2 (N3056, N3054, N677);
nand NAND2 (N3057, N3048, N965);
or OR2 (N3058, N3041, N1634);
nor NOR4 (N3059, N3040, N1901, N2857, N515);
buf BUF1 (N3060, N3053);
and AND4 (N3061, N3045, N154, N229, N2090);
not NOT1 (N3062, N3061);
nand NAND4 (N3063, N3062, N1240, N756, N99);
not NOT1 (N3064, N3047);
nand NAND3 (N3065, N3058, N253, N2120);
xor XOR2 (N3066, N3057, N1582);
xor XOR2 (N3067, N3060, N2079);
xor XOR2 (N3068, N3065, N2745);
nor NOR2 (N3069, N3055, N2378);
not NOT1 (N3070, N3066);
not NOT1 (N3071, N3052);
and AND2 (N3072, N3070, N1893);
xor XOR2 (N3073, N3069, N1818);
and AND3 (N3074, N3073, N2394, N1903);
xor XOR2 (N3075, N3067, N2408);
buf BUF1 (N3076, N3039);
not NOT1 (N3077, N3076);
not NOT1 (N3078, N3064);
xor XOR2 (N3079, N3072, N2908);
not NOT1 (N3080, N3059);
not NOT1 (N3081, N3063);
nand NAND2 (N3082, N3081, N2417);
or OR3 (N3083, N3075, N274, N2172);
not NOT1 (N3084, N3071);
xor XOR2 (N3085, N3078, N2400);
xor XOR2 (N3086, N3056, N1254);
not NOT1 (N3087, N3083);
xor XOR2 (N3088, N3087, N1033);
xor XOR2 (N3089, N3079, N270);
not NOT1 (N3090, N3088);
nand NAND2 (N3091, N3082, N209);
nor NOR4 (N3092, N3091, N292, N611, N1952);
xor XOR2 (N3093, N3084, N1498);
buf BUF1 (N3094, N3085);
or OR3 (N3095, N3080, N577, N1608);
or OR3 (N3096, N3089, N1606, N2115);
not NOT1 (N3097, N3095);
not NOT1 (N3098, N3097);
buf BUF1 (N3099, N3068);
xor XOR2 (N3100, N3092, N901);
xor XOR2 (N3101, N3100, N1090);
buf BUF1 (N3102, N3094);
not NOT1 (N3103, N3099);
or OR3 (N3104, N3101, N164, N115);
buf BUF1 (N3105, N3086);
buf BUF1 (N3106, N3105);
or OR3 (N3107, N3096, N2970, N269);
xor XOR2 (N3108, N3077, N2578);
nor NOR3 (N3109, N3106, N609, N1008);
nand NAND3 (N3110, N3102, N233, N825);
or OR2 (N3111, N3103, N2974);
and AND2 (N3112, N3098, N680);
buf BUF1 (N3113, N3112);
not NOT1 (N3114, N3104);
nor NOR3 (N3115, N3090, N2713, N177);
buf BUF1 (N3116, N3113);
nand NAND3 (N3117, N3109, N2387, N2572);
xor XOR2 (N3118, N3115, N1448);
xor XOR2 (N3119, N3108, N2010);
nor NOR4 (N3120, N3118, N18, N2127, N960);
xor XOR2 (N3121, N3119, N1504);
buf BUF1 (N3122, N3110);
not NOT1 (N3123, N3114);
not NOT1 (N3124, N3074);
or OR4 (N3125, N3123, N15, N2519, N1834);
buf BUF1 (N3126, N3121);
nand NAND2 (N3127, N3111, N2072);
nand NAND3 (N3128, N3122, N1316, N2029);
and AND3 (N3129, N3116, N1579, N1218);
nand NAND3 (N3130, N3120, N2482, N522);
not NOT1 (N3131, N3125);
xor XOR2 (N3132, N3126, N1661);
not NOT1 (N3133, N3129);
and AND2 (N3134, N3107, N2071);
buf BUF1 (N3135, N3133);
not NOT1 (N3136, N3135);
and AND2 (N3137, N3132, N2574);
buf BUF1 (N3138, N3117);
not NOT1 (N3139, N3134);
buf BUF1 (N3140, N3137);
not NOT1 (N3141, N3127);
buf BUF1 (N3142, N3139);
buf BUF1 (N3143, N3138);
and AND4 (N3144, N3093, N2503, N2432, N617);
buf BUF1 (N3145, N3142);
xor XOR2 (N3146, N3145, N2650);
and AND4 (N3147, N3140, N1666, N2490, N1914);
xor XOR2 (N3148, N3147, N194);
nor NOR3 (N3149, N3124, N34, N3134);
buf BUF1 (N3150, N3136);
nor NOR4 (N3151, N3146, N1487, N1482, N1137);
buf BUF1 (N3152, N3151);
buf BUF1 (N3153, N3130);
and AND4 (N3154, N3148, N2341, N2391, N1235);
not NOT1 (N3155, N3154);
xor XOR2 (N3156, N3143, N876);
nor NOR2 (N3157, N3144, N1165);
or OR4 (N3158, N3157, N1888, N10, N802);
nand NAND4 (N3159, N3149, N2821, N2827, N2423);
not NOT1 (N3160, N3159);
xor XOR2 (N3161, N3158, N2462);
xor XOR2 (N3162, N3161, N1871);
buf BUF1 (N3163, N3155);
or OR4 (N3164, N3150, N2937, N2786, N935);
nand NAND4 (N3165, N3128, N2638, N1510, N3103);
not NOT1 (N3166, N3152);
nor NOR2 (N3167, N3165, N2868);
xor XOR2 (N3168, N3141, N1829);
nor NOR4 (N3169, N3156, N1334, N2113, N2045);
or OR4 (N3170, N3169, N570, N1789, N2550);
nand NAND3 (N3171, N3164, N110, N2293);
not NOT1 (N3172, N3167);
buf BUF1 (N3173, N3168);
buf BUF1 (N3174, N3166);
nand NAND3 (N3175, N3160, N826, N1667);
and AND3 (N3176, N3173, N2655, N1342);
or OR3 (N3177, N3131, N2687, N111);
not NOT1 (N3178, N3153);
or OR2 (N3179, N3163, N2448);
and AND3 (N3180, N3174, N1279, N1934);
and AND4 (N3181, N3172, N795, N1394, N2510);
buf BUF1 (N3182, N3181);
buf BUF1 (N3183, N3180);
buf BUF1 (N3184, N3176);
nand NAND2 (N3185, N3177, N518);
xor XOR2 (N3186, N3185, N2959);
xor XOR2 (N3187, N3171, N2386);
and AND3 (N3188, N3183, N3145, N38);
nor NOR2 (N3189, N3170, N309);
or OR4 (N3190, N3162, N2977, N148, N2879);
or OR3 (N3191, N3182, N1960, N379);
xor XOR2 (N3192, N3188, N1537);
not NOT1 (N3193, N3186);
and AND3 (N3194, N3179, N567, N725);
or OR2 (N3195, N3187, N2508);
and AND2 (N3196, N3178, N2924);
buf BUF1 (N3197, N3190);
nand NAND4 (N3198, N3197, N2216, N2780, N1579);
or OR3 (N3199, N3196, N32, N213);
nor NOR3 (N3200, N3191, N76, N1221);
not NOT1 (N3201, N3195);
not NOT1 (N3202, N3201);
nor NOR4 (N3203, N3193, N1410, N2571, N1439);
not NOT1 (N3204, N3184);
nand NAND3 (N3205, N3198, N1949, N2246);
or OR2 (N3206, N3175, N1416);
nor NOR3 (N3207, N3202, N2483, N64);
buf BUF1 (N3208, N3194);
xor XOR2 (N3209, N3207, N2735);
nand NAND3 (N3210, N3200, N2142, N123);
not NOT1 (N3211, N3209);
or OR4 (N3212, N3203, N508, N2928, N54);
not NOT1 (N3213, N3204);
nand NAND4 (N3214, N3206, N303, N387, N1602);
or OR3 (N3215, N3211, N1484, N1956);
endmodule